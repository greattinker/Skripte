// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17;

output N415,N399,N402,N400,N407,N398,N408,N416,N412,N417;

or OR2 (N18, N9, N17);
not NOT1 (N19, N9);
buf BUF1 (N20, N7);
xor XOR2 (N21, N1, N4);
nor NOR2 (N22, N4, N12);
nor NOR3 (N23, N3, N17, N6);
or OR2 (N24, N6, N11);
nor NOR2 (N25, N23, N16);
buf BUF1 (N26, N8);
nor NOR4 (N27, N13, N12, N8, N18);
xor XOR2 (N28, N18, N20);
and AND4 (N29, N26, N26, N23, N19);
buf BUF1 (N30, N27);
not NOT1 (N31, N5);
buf BUF1 (N32, N27);
buf BUF1 (N33, N8);
and AND2 (N34, N21, N29);
nand NAND2 (N35, N22, N17);
buf BUF1 (N36, N14);
not NOT1 (N37, N34);
nand NAND4 (N38, N28, N4, N33, N20);
and AND3 (N39, N22, N7, N1);
nand NAND4 (N40, N31, N33, N15, N7);
nand NAND2 (N41, N39, N37);
or OR3 (N42, N33, N24, N34);
or OR3 (N43, N5, N40, N41);
xor XOR2 (N44, N2, N34);
nor NOR3 (N45, N13, N9, N4);
nor NOR2 (N46, N42, N32);
buf BUF1 (N47, N25);
and AND3 (N48, N43, N27, N44);
nor NOR3 (N49, N43, N28, N2);
not NOT1 (N50, N29);
nand NAND4 (N51, N47, N30, N31, N41);
nand NAND4 (N52, N18, N27, N15, N1);
not NOT1 (N53, N45);
buf BUF1 (N54, N53);
xor XOR2 (N55, N46, N45);
or OR2 (N56, N35, N28);
and AND4 (N57, N50, N20, N48, N29);
buf BUF1 (N58, N45);
xor XOR2 (N59, N49, N14);
and AND4 (N60, N38, N1, N58, N53);
and AND3 (N61, N1, N50, N37);
and AND3 (N62, N36, N31, N19);
and AND3 (N63, N52, N4, N46);
not NOT1 (N64, N61);
nand NAND4 (N65, N54, N39, N34, N8);
not NOT1 (N66, N55);
xor XOR2 (N67, N65, N43);
or OR2 (N68, N62, N63);
or OR3 (N69, N34, N13, N36);
nor NOR3 (N70, N67, N31, N22);
nor NOR3 (N71, N66, N39, N16);
xor XOR2 (N72, N68, N51);
nor NOR4 (N73, N28, N40, N66, N38);
and AND4 (N74, N59, N69, N15, N47);
xor XOR2 (N75, N17, N47);
buf BUF1 (N76, N64);
nor NOR2 (N77, N72, N68);
buf BUF1 (N78, N60);
buf BUF1 (N79, N56);
not NOT1 (N80, N70);
nor NOR4 (N81, N71, N44, N59, N65);
buf BUF1 (N82, N73);
nand NAND3 (N83, N75, N18, N34);
nand NAND4 (N84, N81, N43, N24, N22);
nand NAND2 (N85, N57, N57);
xor XOR2 (N86, N76, N74);
buf BUF1 (N87, N35);
not NOT1 (N88, N86);
xor XOR2 (N89, N78, N42);
or OR2 (N90, N87, N33);
buf BUF1 (N91, N85);
buf BUF1 (N92, N79);
buf BUF1 (N93, N91);
or OR3 (N94, N83, N14, N5);
xor XOR2 (N95, N82, N13);
nand NAND4 (N96, N92, N73, N11, N26);
xor XOR2 (N97, N94, N68);
and AND2 (N98, N88, N34);
or OR3 (N99, N97, N43, N66);
not NOT1 (N100, N98);
not NOT1 (N101, N90);
nor NOR4 (N102, N80, N25, N78, N92);
not NOT1 (N103, N100);
not NOT1 (N104, N99);
or OR3 (N105, N77, N80, N6);
nor NOR4 (N106, N96, N77, N15, N1);
not NOT1 (N107, N95);
nand NAND2 (N108, N107, N107);
or OR2 (N109, N102, N101);
xor XOR2 (N110, N77, N10);
nand NAND4 (N111, N104, N93, N3, N6);
xor XOR2 (N112, N11, N91);
not NOT1 (N113, N105);
buf BUF1 (N114, N84);
or OR2 (N115, N112, N29);
xor XOR2 (N116, N113, N58);
and AND3 (N117, N108, N77, N50);
buf BUF1 (N118, N111);
xor XOR2 (N119, N118, N101);
not NOT1 (N120, N106);
xor XOR2 (N121, N115, N17);
nor NOR3 (N122, N103, N5, N12);
nand NAND4 (N123, N117, N83, N15, N121);
nand NAND3 (N124, N95, N74, N64);
and AND4 (N125, N120, N4, N117, N72);
nor NOR4 (N126, N124, N91, N63, N101);
buf BUF1 (N127, N126);
not NOT1 (N128, N110);
and AND2 (N129, N114, N125);
not NOT1 (N130, N76);
buf BUF1 (N131, N109);
not NOT1 (N132, N89);
not NOT1 (N133, N119);
buf BUF1 (N134, N133);
and AND2 (N135, N132, N60);
nand NAND2 (N136, N122, N57);
buf BUF1 (N137, N136);
xor XOR2 (N138, N129, N38);
xor XOR2 (N139, N130, N32);
nand NAND4 (N140, N137, N107, N39, N45);
nand NAND2 (N141, N128, N125);
buf BUF1 (N142, N135);
and AND2 (N143, N123, N88);
buf BUF1 (N144, N141);
buf BUF1 (N145, N127);
nand NAND4 (N146, N138, N101, N85, N71);
not NOT1 (N147, N144);
and AND3 (N148, N146, N130, N8);
nand NAND3 (N149, N147, N77, N113);
xor XOR2 (N150, N145, N42);
or OR4 (N151, N143, N21, N92, N101);
not NOT1 (N152, N116);
buf BUF1 (N153, N140);
nor NOR2 (N154, N150, N150);
nor NOR3 (N155, N154, N139, N123);
xor XOR2 (N156, N43, N24);
or OR3 (N157, N153, N88, N4);
not NOT1 (N158, N156);
nor NOR4 (N159, N134, N136, N1, N137);
nor NOR2 (N160, N142, N39);
xor XOR2 (N161, N152, N142);
buf BUF1 (N162, N157);
nand NAND2 (N163, N162, N144);
nor NOR4 (N164, N160, N156, N163, N86);
or OR2 (N165, N161, N122);
or OR2 (N166, N78, N65);
xor XOR2 (N167, N158, N140);
xor XOR2 (N168, N131, N2);
nor NOR2 (N169, N168, N56);
xor XOR2 (N170, N165, N97);
and AND3 (N171, N155, N102, N67);
nand NAND2 (N172, N170, N81);
nor NOR3 (N173, N169, N131, N65);
nor NOR4 (N174, N167, N25, N27, N145);
not NOT1 (N175, N174);
nor NOR2 (N176, N149, N29);
xor XOR2 (N177, N173, N45);
or OR2 (N178, N164, N103);
buf BUF1 (N179, N172);
xor XOR2 (N180, N171, N103);
and AND2 (N181, N175, N130);
buf BUF1 (N182, N148);
or OR3 (N183, N151, N40, N110);
and AND2 (N184, N182, N129);
nor NOR4 (N185, N179, N80, N111, N135);
buf BUF1 (N186, N185);
and AND2 (N187, N184, N135);
nand NAND3 (N188, N183, N103, N41);
not NOT1 (N189, N187);
nand NAND3 (N190, N188, N182, N82);
or OR2 (N191, N190, N55);
or OR3 (N192, N159, N101, N165);
nor NOR3 (N193, N178, N123, N139);
or OR2 (N194, N181, N98);
buf BUF1 (N195, N194);
xor XOR2 (N196, N176, N88);
not NOT1 (N197, N195);
buf BUF1 (N198, N180);
nor NOR2 (N199, N191, N128);
and AND4 (N200, N192, N139, N115, N109);
xor XOR2 (N201, N166, N16);
not NOT1 (N202, N198);
xor XOR2 (N203, N193, N20);
nand NAND4 (N204, N189, N124, N112, N154);
xor XOR2 (N205, N197, N103);
buf BUF1 (N206, N203);
buf BUF1 (N207, N196);
xor XOR2 (N208, N202, N141);
buf BUF1 (N209, N177);
buf BUF1 (N210, N205);
nor NOR4 (N211, N206, N159, N117, N158);
or OR4 (N212, N200, N30, N210, N197);
nor NOR4 (N213, N41, N82, N50, N75);
nor NOR3 (N214, N186, N76, N20);
not NOT1 (N215, N204);
xor XOR2 (N216, N215, N166);
and AND3 (N217, N207, N101, N9);
nor NOR3 (N218, N208, N130, N184);
nand NAND4 (N219, N212, N11, N54, N170);
and AND4 (N220, N211, N183, N67, N82);
nor NOR2 (N221, N214, N94);
nand NAND3 (N222, N218, N88, N142);
and AND4 (N223, N220, N56, N160, N144);
nor NOR3 (N224, N223, N125, N48);
nand NAND2 (N225, N209, N77);
not NOT1 (N226, N219);
nand NAND4 (N227, N213, N149, N54, N38);
xor XOR2 (N228, N225, N51);
buf BUF1 (N229, N226);
and AND4 (N230, N201, N139, N105, N26);
nor NOR4 (N231, N229, N191, N191, N71);
nand NAND4 (N232, N231, N104, N193, N150);
nand NAND2 (N233, N224, N34);
nor NOR2 (N234, N217, N162);
nand NAND2 (N235, N228, N44);
or OR3 (N236, N221, N165, N140);
nand NAND2 (N237, N216, N69);
xor XOR2 (N238, N232, N221);
not NOT1 (N239, N227);
nor NOR4 (N240, N238, N87, N78, N7);
not NOT1 (N241, N199);
nor NOR4 (N242, N234, N133, N170, N96);
or OR3 (N243, N237, N174, N34);
buf BUF1 (N244, N236);
or OR4 (N245, N241, N195, N160, N3);
xor XOR2 (N246, N233, N2);
and AND4 (N247, N243, N106, N47, N74);
buf BUF1 (N248, N245);
nor NOR2 (N249, N235, N92);
or OR4 (N250, N242, N170, N204, N234);
or OR3 (N251, N247, N135, N232);
not NOT1 (N252, N251);
buf BUF1 (N253, N222);
not NOT1 (N254, N253);
xor XOR2 (N255, N240, N17);
nand NAND4 (N256, N230, N116, N74, N173);
not NOT1 (N257, N248);
buf BUF1 (N258, N256);
or OR4 (N259, N258, N35, N9, N248);
nor NOR2 (N260, N250, N57);
and AND4 (N261, N246, N173, N151, N233);
xor XOR2 (N262, N259, N78);
not NOT1 (N263, N257);
nor NOR2 (N264, N249, N30);
or OR3 (N265, N260, N19, N187);
nor NOR3 (N266, N239, N179, N79);
and AND4 (N267, N265, N14, N106, N148);
or OR3 (N268, N261, N202, N189);
xor XOR2 (N269, N254, N218);
buf BUF1 (N270, N262);
or OR2 (N271, N263, N255);
nand NAND2 (N272, N176, N86);
xor XOR2 (N273, N264, N54);
and AND2 (N274, N272, N15);
xor XOR2 (N275, N271, N25);
not NOT1 (N276, N252);
not NOT1 (N277, N270);
nand NAND4 (N278, N276, N18, N126, N169);
nand NAND4 (N279, N267, N251, N119, N219);
and AND4 (N280, N275, N131, N237, N18);
nor NOR2 (N281, N274, N50);
buf BUF1 (N282, N273);
not NOT1 (N283, N266);
and AND3 (N284, N278, N160, N14);
nor NOR2 (N285, N280, N8);
nand NAND2 (N286, N277, N259);
nor NOR2 (N287, N269, N238);
or OR4 (N288, N244, N94, N130, N138);
not NOT1 (N289, N282);
and AND2 (N290, N284, N45);
and AND2 (N291, N289, N51);
buf BUF1 (N292, N283);
and AND3 (N293, N285, N32, N96);
or OR3 (N294, N279, N266, N234);
nor NOR4 (N295, N294, N57, N220, N114);
nor NOR2 (N296, N288, N223);
nand NAND2 (N297, N290, N156);
nor NOR4 (N298, N291, N15, N195, N78);
nor NOR4 (N299, N297, N58, N40, N65);
and AND3 (N300, N287, N13, N120);
and AND4 (N301, N286, N252, N30, N50);
or OR2 (N302, N298, N59);
not NOT1 (N303, N281);
or OR2 (N304, N268, N19);
buf BUF1 (N305, N295);
buf BUF1 (N306, N304);
nand NAND4 (N307, N301, N230, N279, N265);
xor XOR2 (N308, N300, N105);
and AND3 (N309, N292, N139, N148);
buf BUF1 (N310, N293);
xor XOR2 (N311, N296, N11);
xor XOR2 (N312, N307, N207);
not NOT1 (N313, N299);
xor XOR2 (N314, N305, N15);
not NOT1 (N315, N310);
buf BUF1 (N316, N309);
or OR3 (N317, N312, N68, N273);
not NOT1 (N318, N311);
not NOT1 (N319, N313);
not NOT1 (N320, N303);
not NOT1 (N321, N302);
nand NAND3 (N322, N308, N44, N254);
not NOT1 (N323, N320);
nor NOR2 (N324, N321, N179);
buf BUF1 (N325, N316);
or OR2 (N326, N306, N204);
nor NOR2 (N327, N323, N256);
nand NAND3 (N328, N317, N105, N47);
not NOT1 (N329, N327);
nor NOR4 (N330, N314, N309, N88, N196);
nor NOR2 (N331, N330, N238);
or OR2 (N332, N322, N289);
and AND3 (N333, N318, N62, N251);
buf BUF1 (N334, N331);
or OR4 (N335, N324, N330, N94, N303);
or OR3 (N336, N315, N209, N257);
or OR2 (N337, N325, N310);
and AND2 (N338, N329, N164);
not NOT1 (N339, N328);
nand NAND4 (N340, N335, N23, N202, N76);
buf BUF1 (N341, N334);
and AND2 (N342, N319, N152);
nor NOR3 (N343, N333, N174, N2);
nor NOR3 (N344, N336, N45, N247);
nand NAND4 (N345, N326, N317, N198, N6);
and AND2 (N346, N342, N248);
nand NAND4 (N347, N343, N170, N119, N335);
or OR3 (N348, N347, N90, N57);
xor XOR2 (N349, N338, N76);
not NOT1 (N350, N337);
and AND2 (N351, N339, N157);
nand NAND2 (N352, N341, N146);
not NOT1 (N353, N340);
nor NOR3 (N354, N350, N213, N239);
nand NAND4 (N355, N348, N228, N68, N129);
xor XOR2 (N356, N345, N11);
xor XOR2 (N357, N353, N126);
xor XOR2 (N358, N346, N3);
nor NOR2 (N359, N332, N284);
not NOT1 (N360, N351);
nand NAND2 (N361, N360, N24);
or OR4 (N362, N357, N3, N50, N119);
not NOT1 (N363, N344);
and AND4 (N364, N363, N137, N144, N79);
not NOT1 (N365, N364);
buf BUF1 (N366, N361);
nor NOR4 (N367, N365, N52, N306, N245);
not NOT1 (N368, N359);
not NOT1 (N369, N367);
and AND4 (N370, N355, N259, N38, N330);
or OR3 (N371, N370, N364, N5);
buf BUF1 (N372, N358);
nor NOR3 (N373, N354, N35, N304);
not NOT1 (N374, N362);
or OR4 (N375, N374, N187, N112, N78);
nand NAND2 (N376, N368, N57);
or OR4 (N377, N372, N7, N179, N118);
nor NOR3 (N378, N373, N296, N123);
and AND4 (N379, N371, N123, N59, N310);
not NOT1 (N380, N356);
or OR2 (N381, N369, N155);
or OR3 (N382, N375, N158, N151);
or OR2 (N383, N378, N210);
nand NAND3 (N384, N366, N162, N257);
nor NOR3 (N385, N349, N59, N174);
nand NAND3 (N386, N381, N256, N309);
nand NAND2 (N387, N382, N46);
nor NOR4 (N388, N386, N83, N111, N289);
not NOT1 (N389, N377);
nand NAND3 (N390, N376, N65, N288);
buf BUF1 (N391, N388);
buf BUF1 (N392, N389);
buf BUF1 (N393, N380);
nor NOR2 (N394, N387, N83);
xor XOR2 (N395, N352, N4);
or OR2 (N396, N391, N11);
not NOT1 (N397, N393);
and AND2 (N398, N385, N16);
nor NOR4 (N399, N384, N335, N299, N278);
and AND2 (N400, N392, N19);
or OR4 (N401, N395, N397, N228, N160);
buf BUF1 (N402, N157);
not NOT1 (N403, N396);
nand NAND4 (N404, N403, N108, N200, N382);
nand NAND3 (N405, N401, N31, N342);
xor XOR2 (N406, N405, N194);
not NOT1 (N407, N390);
nor NOR2 (N408, N394, N355);
xor XOR2 (N409, N406, N157);
or OR4 (N410, N379, N221, N90, N332);
xor XOR2 (N411, N404, N22);
nor NOR3 (N412, N411, N343, N113);
buf BUF1 (N413, N383);
or OR3 (N414, N410, N298, N149);
xor XOR2 (N415, N413, N382);
nor NOR4 (N416, N409, N242, N114, N216);
xor XOR2 (N417, N414, N242);
endmodule