// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;

output N814,N816,N817,N805,N808,N803,N812,N815,N795,N818;

and AND4 (N19, N9, N16, N8, N17);
nor NOR2 (N20, N19, N19);
xor XOR2 (N21, N8, N20);
nor NOR2 (N22, N16, N11);
nor NOR3 (N23, N10, N15, N5);
and AND2 (N24, N17, N17);
nor NOR3 (N25, N19, N5, N5);
nand NAND2 (N26, N25, N19);
xor XOR2 (N27, N24, N20);
not NOT1 (N28, N19);
nand NAND3 (N29, N25, N3, N6);
or OR4 (N30, N16, N25, N6, N17);
nor NOR3 (N31, N10, N24, N12);
not NOT1 (N32, N23);
not NOT1 (N33, N22);
not NOT1 (N34, N28);
nor NOR3 (N35, N27, N21, N15);
not NOT1 (N36, N18);
nor NOR4 (N37, N8, N33, N2, N24);
not NOT1 (N38, N22);
buf BUF1 (N39, N31);
xor XOR2 (N40, N35, N17);
or OR2 (N41, N38, N16);
and AND3 (N42, N29, N14, N39);
or OR2 (N43, N8, N5);
nand NAND3 (N44, N30, N26, N30);
not NOT1 (N45, N29);
not NOT1 (N46, N43);
nand NAND3 (N47, N42, N18, N18);
nand NAND4 (N48, N46, N1, N27, N45);
and AND4 (N49, N42, N34, N7, N5);
or OR2 (N50, N13, N24);
buf BUF1 (N51, N49);
nand NAND2 (N52, N51, N22);
xor XOR2 (N53, N40, N38);
and AND2 (N54, N50, N50);
buf BUF1 (N55, N52);
not NOT1 (N56, N48);
and AND2 (N57, N41, N37);
nand NAND3 (N58, N23, N39, N33);
buf BUF1 (N59, N57);
xor XOR2 (N60, N55, N42);
not NOT1 (N61, N36);
nor NOR3 (N62, N61, N54, N35);
buf BUF1 (N63, N60);
buf BUF1 (N64, N24);
not NOT1 (N65, N53);
not NOT1 (N66, N62);
and AND2 (N67, N63, N63);
or OR2 (N68, N67, N37);
buf BUF1 (N69, N56);
or OR4 (N70, N47, N30, N2, N42);
nor NOR4 (N71, N44, N3, N7, N26);
xor XOR2 (N72, N68, N55);
xor XOR2 (N73, N58, N60);
not NOT1 (N74, N66);
or OR4 (N75, N70, N52, N37, N49);
not NOT1 (N76, N73);
nor NOR3 (N77, N76, N11, N35);
buf BUF1 (N78, N32);
not NOT1 (N79, N59);
buf BUF1 (N80, N74);
nand NAND4 (N81, N78, N72, N31, N17);
or OR2 (N82, N80, N52);
and AND3 (N83, N7, N1, N18);
or OR4 (N84, N83, N12, N42, N13);
buf BUF1 (N85, N84);
nand NAND3 (N86, N71, N70, N33);
not NOT1 (N87, N75);
nor NOR4 (N88, N82, N34, N57, N37);
nand NAND3 (N89, N86, N26, N11);
not NOT1 (N90, N85);
xor XOR2 (N91, N81, N63);
not NOT1 (N92, N91);
nand NAND2 (N93, N79, N5);
buf BUF1 (N94, N93);
nand NAND3 (N95, N94, N41, N3);
nand NAND4 (N96, N87, N43, N87, N26);
and AND2 (N97, N77, N38);
and AND3 (N98, N97, N96, N50);
nor NOR2 (N99, N27, N43);
or OR2 (N100, N69, N75);
xor XOR2 (N101, N100, N7);
nand NAND2 (N102, N92, N87);
xor XOR2 (N103, N102, N56);
buf BUF1 (N104, N103);
nor NOR3 (N105, N95, N55, N90);
not NOT1 (N106, N103);
buf BUF1 (N107, N65);
xor XOR2 (N108, N98, N21);
and AND4 (N109, N104, N49, N74, N84);
nor NOR2 (N110, N64, N24);
not NOT1 (N111, N88);
nand NAND3 (N112, N108, N65, N46);
buf BUF1 (N113, N112);
buf BUF1 (N114, N107);
nor NOR3 (N115, N109, N50, N114);
or OR3 (N116, N13, N43, N44);
not NOT1 (N117, N99);
nand NAND4 (N118, N106, N56, N15, N84);
buf BUF1 (N119, N113);
not NOT1 (N120, N110);
nand NAND2 (N121, N118, N77);
nand NAND3 (N122, N116, N70, N106);
nor NOR4 (N123, N101, N86, N64, N101);
and AND2 (N124, N121, N107);
nor NOR4 (N125, N89, N106, N85, N77);
nor NOR3 (N126, N115, N107, N84);
xor XOR2 (N127, N122, N37);
or OR4 (N128, N119, N74, N1, N14);
or OR4 (N129, N126, N93, N37, N122);
nand NAND4 (N130, N129, N39, N25, N2);
xor XOR2 (N131, N125, N35);
xor XOR2 (N132, N120, N112);
not NOT1 (N133, N124);
buf BUF1 (N134, N131);
not NOT1 (N135, N111);
and AND3 (N136, N117, N37, N59);
nor NOR2 (N137, N135, N47);
and AND2 (N138, N137, N25);
nor NOR3 (N139, N136, N85, N130);
nor NOR3 (N140, N28, N52, N26);
and AND2 (N141, N140, N79);
or OR4 (N142, N133, N90, N62, N8);
nor NOR4 (N143, N132, N138, N27, N50);
and AND2 (N144, N139, N14);
xor XOR2 (N145, N12, N127);
xor XOR2 (N146, N38, N86);
nor NOR2 (N147, N145, N55);
nor NOR4 (N148, N128, N45, N48, N26);
nor NOR4 (N149, N123, N6, N95, N116);
nand NAND4 (N150, N142, N137, N94, N7);
and AND2 (N151, N150, N4);
and AND3 (N152, N144, N75, N16);
nor NOR3 (N153, N143, N77, N64);
and AND2 (N154, N141, N91);
buf BUF1 (N155, N105);
or OR3 (N156, N134, N94, N25);
nand NAND3 (N157, N151, N21, N16);
xor XOR2 (N158, N146, N141);
xor XOR2 (N159, N153, N6);
nand NAND2 (N160, N149, N37);
nor NOR3 (N161, N148, N57, N154);
not NOT1 (N162, N121);
not NOT1 (N163, N156);
or OR4 (N164, N152, N122, N4, N155);
xor XOR2 (N165, N87, N27);
buf BUF1 (N166, N165);
xor XOR2 (N167, N162, N121);
nor NOR2 (N168, N160, N87);
buf BUF1 (N169, N157);
buf BUF1 (N170, N158);
nand NAND2 (N171, N147, N127);
nand NAND4 (N172, N159, N39, N135, N76);
nor NOR3 (N173, N167, N130, N98);
xor XOR2 (N174, N161, N33);
buf BUF1 (N175, N174);
buf BUF1 (N176, N175);
and AND3 (N177, N164, N12, N44);
nor NOR3 (N178, N170, N70, N151);
nand NAND2 (N179, N178, N95);
nand NAND4 (N180, N171, N67, N5, N71);
nand NAND4 (N181, N172, N24, N145, N2);
or OR2 (N182, N181, N59);
or OR3 (N183, N177, N53, N125);
nand NAND3 (N184, N173, N158, N100);
nor NOR4 (N185, N169, N165, N125, N129);
nor NOR2 (N186, N179, N135);
nand NAND2 (N187, N184, N170);
not NOT1 (N188, N163);
nor NOR4 (N189, N180, N36, N178, N25);
buf BUF1 (N190, N188);
and AND4 (N191, N190, N50, N38, N19);
or OR2 (N192, N176, N123);
xor XOR2 (N193, N189, N81);
or OR4 (N194, N193, N149, N31, N75);
or OR2 (N195, N187, N60);
not NOT1 (N196, N168);
not NOT1 (N197, N182);
nand NAND2 (N198, N185, N107);
not NOT1 (N199, N186);
xor XOR2 (N200, N198, N145);
or OR3 (N201, N199, N12, N86);
nand NAND4 (N202, N195, N190, N146, N74);
nor NOR3 (N203, N192, N33, N139);
not NOT1 (N204, N183);
or OR2 (N205, N203, N141);
or OR3 (N206, N200, N192, N190);
nand NAND2 (N207, N201, N76);
and AND2 (N208, N202, N153);
xor XOR2 (N209, N191, N114);
buf BUF1 (N210, N206);
not NOT1 (N211, N197);
or OR3 (N212, N210, N54, N29);
buf BUF1 (N213, N194);
buf BUF1 (N214, N213);
not NOT1 (N215, N208);
nand NAND4 (N216, N209, N212, N178, N61);
nand NAND4 (N217, N160, N186, N178, N60);
nand NAND3 (N218, N214, N62, N124);
nor NOR2 (N219, N196, N46);
nand NAND4 (N220, N215, N204, N13, N127);
xor XOR2 (N221, N55, N118);
xor XOR2 (N222, N166, N169);
nor NOR4 (N223, N218, N95, N163, N193);
nand NAND4 (N224, N219, N221, N60, N82);
and AND2 (N225, N193, N182);
not NOT1 (N226, N216);
nor NOR3 (N227, N211, N141, N146);
xor XOR2 (N228, N207, N28);
not NOT1 (N229, N217);
buf BUF1 (N230, N224);
and AND3 (N231, N205, N2, N120);
nand NAND4 (N232, N228, N93, N85, N160);
nor NOR3 (N233, N231, N18, N71);
or OR2 (N234, N223, N93);
nand NAND4 (N235, N234, N84, N61, N123);
nor NOR4 (N236, N227, N32, N43, N188);
or OR2 (N237, N225, N21);
not NOT1 (N238, N226);
xor XOR2 (N239, N233, N153);
nor NOR4 (N240, N229, N162, N130, N224);
nand NAND2 (N241, N222, N239);
and AND2 (N242, N160, N92);
xor XOR2 (N243, N237, N143);
or OR2 (N244, N242, N209);
buf BUF1 (N245, N235);
or OR3 (N246, N241, N210, N171);
or OR4 (N247, N232, N19, N124, N96);
nor NOR2 (N248, N230, N219);
and AND2 (N249, N245, N205);
nand NAND4 (N250, N247, N213, N71, N167);
nand NAND2 (N251, N249, N150);
nand NAND3 (N252, N250, N235, N40);
not NOT1 (N253, N251);
buf BUF1 (N254, N252);
not NOT1 (N255, N244);
not NOT1 (N256, N236);
and AND2 (N257, N240, N156);
and AND2 (N258, N220, N43);
not NOT1 (N259, N248);
buf BUF1 (N260, N255);
and AND3 (N261, N253, N198, N76);
or OR3 (N262, N238, N94, N79);
nand NAND3 (N263, N262, N181, N155);
and AND4 (N264, N259, N217, N83, N174);
not NOT1 (N265, N261);
not NOT1 (N266, N257);
xor XOR2 (N267, N263, N231);
buf BUF1 (N268, N266);
buf BUF1 (N269, N246);
buf BUF1 (N270, N260);
not NOT1 (N271, N256);
nor NOR4 (N272, N268, N104, N209, N243);
buf BUF1 (N273, N95);
not NOT1 (N274, N254);
not NOT1 (N275, N258);
not NOT1 (N276, N272);
and AND4 (N277, N270, N12, N167, N98);
nand NAND3 (N278, N267, N118, N220);
nand NAND4 (N279, N277, N52, N144, N209);
and AND3 (N280, N264, N94, N243);
and AND4 (N281, N276, N211, N115, N209);
nor NOR3 (N282, N275, N17, N127);
xor XOR2 (N283, N282, N28);
not NOT1 (N284, N273);
xor XOR2 (N285, N269, N229);
xor XOR2 (N286, N278, N187);
nand NAND2 (N287, N271, N168);
and AND3 (N288, N286, N107, N127);
not NOT1 (N289, N283);
or OR3 (N290, N280, N240, N208);
nor NOR3 (N291, N289, N232, N253);
nor NOR2 (N292, N281, N87);
xor XOR2 (N293, N284, N138);
or OR3 (N294, N287, N152, N93);
nor NOR3 (N295, N285, N71, N87);
xor XOR2 (N296, N265, N171);
xor XOR2 (N297, N288, N64);
xor XOR2 (N298, N294, N204);
and AND2 (N299, N295, N107);
not NOT1 (N300, N292);
not NOT1 (N301, N290);
not NOT1 (N302, N301);
nand NAND2 (N303, N300, N34);
not NOT1 (N304, N293);
or OR2 (N305, N302, N10);
nand NAND3 (N306, N299, N150, N29);
nor NOR2 (N307, N305, N240);
or OR4 (N308, N291, N133, N244, N188);
nand NAND4 (N309, N297, N67, N292, N167);
and AND3 (N310, N309, N46, N148);
nor NOR4 (N311, N298, N180, N72, N293);
nand NAND2 (N312, N308, N279);
and AND2 (N313, N114, N186);
xor XOR2 (N314, N313, N230);
or OR4 (N315, N314, N21, N36, N150);
not NOT1 (N316, N315);
and AND3 (N317, N274, N187, N253);
nand NAND3 (N318, N316, N189, N62);
not NOT1 (N319, N303);
not NOT1 (N320, N304);
nor NOR3 (N321, N311, N209, N149);
not NOT1 (N322, N296);
not NOT1 (N323, N310);
nand NAND3 (N324, N306, N113, N122);
and AND3 (N325, N322, N282, N203);
not NOT1 (N326, N325);
nor NOR2 (N327, N319, N155);
xor XOR2 (N328, N324, N193);
or OR2 (N329, N320, N69);
not NOT1 (N330, N318);
buf BUF1 (N331, N326);
or OR2 (N332, N330, N65);
buf BUF1 (N333, N323);
nand NAND4 (N334, N317, N181, N309, N99);
nor NOR2 (N335, N332, N277);
xor XOR2 (N336, N321, N105);
not NOT1 (N337, N307);
nor NOR4 (N338, N337, N196, N52, N87);
xor XOR2 (N339, N331, N158);
buf BUF1 (N340, N312);
xor XOR2 (N341, N339, N113);
nand NAND2 (N342, N334, N20);
or OR2 (N343, N342, N146);
not NOT1 (N344, N336);
or OR2 (N345, N333, N336);
nor NOR2 (N346, N343, N23);
buf BUF1 (N347, N327);
nand NAND3 (N348, N340, N298, N344);
buf BUF1 (N349, N68);
xor XOR2 (N350, N349, N317);
not NOT1 (N351, N328);
and AND4 (N352, N329, N219, N200, N175);
nor NOR4 (N353, N348, N237, N141, N312);
not NOT1 (N354, N347);
nand NAND2 (N355, N350, N138);
not NOT1 (N356, N346);
xor XOR2 (N357, N356, N49);
xor XOR2 (N358, N351, N66);
not NOT1 (N359, N352);
not NOT1 (N360, N341);
not NOT1 (N361, N355);
or OR4 (N362, N358, N238, N292, N95);
and AND4 (N363, N338, N179, N276, N246);
or OR3 (N364, N354, N212, N176);
nor NOR4 (N365, N363, N336, N96, N138);
xor XOR2 (N366, N357, N255);
or OR4 (N367, N366, N139, N192, N156);
not NOT1 (N368, N335);
nor NOR2 (N369, N362, N183);
not NOT1 (N370, N368);
buf BUF1 (N371, N345);
or OR2 (N372, N370, N316);
or OR4 (N373, N369, N114, N281, N218);
buf BUF1 (N374, N353);
not NOT1 (N375, N372);
and AND2 (N376, N365, N263);
not NOT1 (N377, N374);
nand NAND2 (N378, N367, N179);
or OR3 (N379, N364, N102, N185);
xor XOR2 (N380, N373, N128);
and AND2 (N381, N360, N369);
nand NAND3 (N382, N377, N152, N37);
buf BUF1 (N383, N379);
or OR3 (N384, N371, N172, N366);
nand NAND4 (N385, N359, N278, N144, N320);
and AND4 (N386, N361, N237, N240, N307);
not NOT1 (N387, N386);
nand NAND4 (N388, N381, N152, N351, N232);
or OR2 (N389, N385, N249);
and AND2 (N390, N384, N107);
not NOT1 (N391, N388);
buf BUF1 (N392, N376);
buf BUF1 (N393, N390);
xor XOR2 (N394, N387, N2);
nor NOR4 (N395, N393, N268, N295, N214);
nand NAND4 (N396, N378, N147, N145, N131);
not NOT1 (N397, N389);
nor NOR3 (N398, N397, N48, N40);
nand NAND4 (N399, N395, N257, N154, N88);
nand NAND4 (N400, N391, N270, N122, N337);
or OR3 (N401, N382, N205, N349);
or OR2 (N402, N400, N43);
nor NOR4 (N403, N396, N275, N89, N5);
nor NOR4 (N404, N375, N140, N40, N188);
buf BUF1 (N405, N398);
not NOT1 (N406, N380);
nor NOR4 (N407, N383, N150, N255, N49);
or OR2 (N408, N401, N258);
xor XOR2 (N409, N399, N360);
nor NOR2 (N410, N407, N340);
nand NAND3 (N411, N410, N224, N10);
nor NOR2 (N412, N405, N320);
not NOT1 (N413, N412);
nor NOR4 (N414, N392, N37, N404, N368);
not NOT1 (N415, N1);
not NOT1 (N416, N402);
buf BUF1 (N417, N409);
not NOT1 (N418, N414);
not NOT1 (N419, N413);
nor NOR3 (N420, N417, N239, N271);
not NOT1 (N421, N411);
and AND3 (N422, N416, N45, N368);
xor XOR2 (N423, N421, N219);
nand NAND4 (N424, N422, N255, N364, N300);
buf BUF1 (N425, N403);
nor NOR4 (N426, N419, N321, N148, N414);
nor NOR2 (N427, N415, N270);
nor NOR2 (N428, N418, N109);
or OR3 (N429, N427, N222, N15);
or OR2 (N430, N429, N91);
or OR2 (N431, N394, N136);
or OR3 (N432, N423, N391, N208);
nand NAND2 (N433, N426, N222);
and AND3 (N434, N430, N200, N80);
nand NAND3 (N435, N425, N398, N381);
buf BUF1 (N436, N408);
nand NAND3 (N437, N435, N227, N261);
xor XOR2 (N438, N428, N224);
buf BUF1 (N439, N434);
nor NOR2 (N440, N433, N258);
and AND4 (N441, N436, N260, N85, N335);
nor NOR3 (N442, N406, N184, N98);
or OR2 (N443, N420, N28);
buf BUF1 (N444, N438);
xor XOR2 (N445, N424, N139);
nand NAND3 (N446, N444, N288, N88);
and AND2 (N447, N431, N6);
or OR2 (N448, N432, N427);
not NOT1 (N449, N443);
buf BUF1 (N450, N448);
nor NOR3 (N451, N446, N156, N417);
not NOT1 (N452, N439);
or OR2 (N453, N450, N200);
not NOT1 (N454, N449);
nor NOR2 (N455, N447, N248);
nor NOR4 (N456, N437, N151, N112, N88);
nand NAND3 (N457, N455, N101, N320);
or OR2 (N458, N454, N159);
not NOT1 (N459, N445);
nor NOR3 (N460, N442, N83, N201);
buf BUF1 (N461, N459);
and AND2 (N462, N441, N109);
xor XOR2 (N463, N458, N374);
and AND4 (N464, N452, N250, N444, N248);
and AND2 (N465, N461, N306);
or OR2 (N466, N440, N144);
nand NAND3 (N467, N466, N395, N102);
buf BUF1 (N468, N467);
nand NAND4 (N469, N457, N129, N444, N213);
and AND2 (N470, N468, N443);
not NOT1 (N471, N460);
not NOT1 (N472, N471);
or OR4 (N473, N470, N259, N170, N334);
buf BUF1 (N474, N473);
or OR4 (N475, N465, N202, N36, N35);
xor XOR2 (N476, N456, N439);
and AND3 (N477, N472, N364, N388);
or OR4 (N478, N453, N460, N430, N452);
nand NAND4 (N479, N469, N445, N241, N123);
xor XOR2 (N480, N474, N202);
and AND3 (N481, N463, N114, N341);
not NOT1 (N482, N480);
and AND2 (N483, N481, N360);
buf BUF1 (N484, N462);
and AND2 (N485, N482, N167);
not NOT1 (N486, N485);
nor NOR2 (N487, N483, N411);
xor XOR2 (N488, N484, N37);
buf BUF1 (N489, N478);
or OR4 (N490, N489, N345, N395, N459);
buf BUF1 (N491, N477);
not NOT1 (N492, N475);
or OR4 (N493, N451, N224, N168, N384);
or OR4 (N494, N479, N128, N37, N438);
and AND2 (N495, N494, N146);
or OR4 (N496, N486, N152, N275, N203);
xor XOR2 (N497, N492, N242);
and AND4 (N498, N488, N246, N395, N466);
and AND3 (N499, N490, N328, N150);
and AND4 (N500, N491, N493, N266, N374);
xor XOR2 (N501, N389, N359);
or OR2 (N502, N496, N106);
not NOT1 (N503, N487);
xor XOR2 (N504, N495, N206);
nand NAND4 (N505, N497, N298, N456, N186);
xor XOR2 (N506, N500, N225);
nand NAND3 (N507, N498, N35, N467);
and AND2 (N508, N476, N95);
nand NAND4 (N509, N506, N222, N92, N168);
and AND3 (N510, N504, N55, N286);
nor NOR3 (N511, N502, N179, N46);
and AND4 (N512, N508, N120, N127, N56);
nor NOR4 (N513, N512, N447, N249, N361);
and AND4 (N514, N501, N123, N344, N72);
not NOT1 (N515, N514);
not NOT1 (N516, N509);
and AND2 (N517, N507, N229);
not NOT1 (N518, N511);
and AND3 (N519, N515, N290, N36);
or OR3 (N520, N505, N128, N295);
not NOT1 (N521, N513);
nand NAND4 (N522, N518, N167, N377, N258);
and AND2 (N523, N503, N4);
or OR4 (N524, N464, N74, N129, N89);
buf BUF1 (N525, N516);
xor XOR2 (N526, N523, N31);
and AND3 (N527, N525, N22, N265);
or OR4 (N528, N510, N395, N259, N253);
not NOT1 (N529, N521);
buf BUF1 (N530, N528);
buf BUF1 (N531, N529);
and AND3 (N532, N517, N237, N103);
or OR3 (N533, N524, N25, N212);
xor XOR2 (N534, N526, N395);
buf BUF1 (N535, N519);
not NOT1 (N536, N522);
not NOT1 (N537, N536);
or OR4 (N538, N527, N190, N190, N472);
nor NOR4 (N539, N534, N206, N291, N99);
and AND2 (N540, N499, N443);
or OR3 (N541, N532, N492, N179);
nor NOR4 (N542, N539, N214, N535, N304);
nand NAND2 (N543, N75, N70);
nor NOR3 (N544, N520, N193, N57);
xor XOR2 (N545, N533, N278);
nand NAND2 (N546, N544, N323);
or OR2 (N547, N530, N232);
nand NAND2 (N548, N541, N451);
xor XOR2 (N549, N538, N294);
or OR2 (N550, N543, N316);
xor XOR2 (N551, N542, N58);
nor NOR2 (N552, N540, N152);
not NOT1 (N553, N537);
nor NOR4 (N554, N548, N149, N60, N420);
xor XOR2 (N555, N553, N17);
and AND4 (N556, N545, N373, N428, N207);
nand NAND4 (N557, N556, N340, N32, N381);
or OR3 (N558, N531, N296, N213);
or OR2 (N559, N557, N103);
buf BUF1 (N560, N546);
not NOT1 (N561, N550);
buf BUF1 (N562, N554);
not NOT1 (N563, N549);
buf BUF1 (N564, N562);
nor NOR2 (N565, N547, N388);
or OR4 (N566, N559, N461, N413, N133);
or OR3 (N567, N566, N311, N213);
and AND2 (N568, N551, N378);
or OR2 (N569, N563, N270);
and AND2 (N570, N569, N351);
or OR2 (N571, N570, N478);
buf BUF1 (N572, N552);
and AND4 (N573, N561, N435, N426, N341);
buf BUF1 (N574, N573);
buf BUF1 (N575, N571);
nor NOR4 (N576, N555, N204, N484, N569);
nor NOR4 (N577, N558, N202, N183, N367);
or OR2 (N578, N575, N185);
nand NAND3 (N579, N572, N335, N568);
nor NOR4 (N580, N377, N301, N553, N174);
nand NAND4 (N581, N576, N468, N169, N470);
xor XOR2 (N582, N567, N407);
buf BUF1 (N583, N574);
not NOT1 (N584, N564);
and AND3 (N585, N580, N479, N224);
and AND4 (N586, N584, N374, N388, N351);
buf BUF1 (N587, N565);
xor XOR2 (N588, N577, N484);
not NOT1 (N589, N581);
nand NAND4 (N590, N586, N483, N326, N391);
xor XOR2 (N591, N585, N525);
nand NAND2 (N592, N587, N530);
buf BUF1 (N593, N589);
nand NAND4 (N594, N590, N342, N47, N398);
buf BUF1 (N595, N591);
and AND3 (N596, N592, N330, N399);
and AND2 (N597, N583, N439);
or OR2 (N598, N596, N532);
and AND2 (N599, N597, N43);
nor NOR4 (N600, N593, N160, N293, N108);
not NOT1 (N601, N579);
not NOT1 (N602, N588);
not NOT1 (N603, N578);
and AND2 (N604, N560, N314);
and AND2 (N605, N601, N95);
not NOT1 (N606, N605);
and AND4 (N607, N582, N219, N315, N423);
nor NOR2 (N608, N607, N149);
buf BUF1 (N609, N603);
nand NAND4 (N610, N594, N43, N50, N67);
nor NOR2 (N611, N609, N143);
not NOT1 (N612, N604);
xor XOR2 (N613, N598, N117);
buf BUF1 (N614, N612);
and AND2 (N615, N608, N553);
nor NOR3 (N616, N611, N421, N335);
nor NOR2 (N617, N599, N112);
xor XOR2 (N618, N616, N93);
nand NAND2 (N619, N606, N462);
nor NOR3 (N620, N595, N249, N105);
or OR4 (N621, N619, N271, N599, N279);
nor NOR4 (N622, N613, N520, N447, N376);
nand NAND3 (N623, N600, N19, N301);
and AND4 (N624, N621, N408, N208, N93);
nand NAND2 (N625, N620, N387);
nor NOR2 (N626, N623, N581);
buf BUF1 (N627, N618);
buf BUF1 (N628, N615);
or OR3 (N629, N625, N606, N184);
xor XOR2 (N630, N627, N575);
xor XOR2 (N631, N628, N561);
nor NOR4 (N632, N626, N145, N453, N78);
and AND3 (N633, N622, N609, N356);
nor NOR4 (N634, N602, N604, N492, N413);
or OR3 (N635, N617, N216, N450);
nor NOR2 (N636, N633, N547);
xor XOR2 (N637, N632, N624);
nand NAND3 (N638, N539, N171, N4);
nand NAND3 (N639, N610, N362, N73);
buf BUF1 (N640, N629);
buf BUF1 (N641, N640);
not NOT1 (N642, N641);
buf BUF1 (N643, N634);
buf BUF1 (N644, N630);
buf BUF1 (N645, N635);
and AND3 (N646, N636, N129, N160);
buf BUF1 (N647, N639);
xor XOR2 (N648, N642, N550);
not NOT1 (N649, N631);
nand NAND2 (N650, N644, N27);
nor NOR2 (N651, N646, N96);
nor NOR2 (N652, N643, N454);
nor NOR2 (N653, N645, N25);
or OR4 (N654, N648, N404, N95, N489);
buf BUF1 (N655, N654);
xor XOR2 (N656, N649, N449);
or OR2 (N657, N614, N66);
buf BUF1 (N658, N653);
nor NOR2 (N659, N657, N190);
xor XOR2 (N660, N655, N152);
buf BUF1 (N661, N660);
not NOT1 (N662, N650);
xor XOR2 (N663, N651, N508);
xor XOR2 (N664, N637, N588);
or OR2 (N665, N662, N517);
buf BUF1 (N666, N638);
not NOT1 (N667, N661);
nor NOR4 (N668, N652, N649, N582, N441);
not NOT1 (N669, N659);
or OR2 (N670, N663, N370);
or OR2 (N671, N669, N588);
not NOT1 (N672, N665);
nand NAND3 (N673, N671, N479, N254);
not NOT1 (N674, N668);
buf BUF1 (N675, N672);
buf BUF1 (N676, N656);
not NOT1 (N677, N647);
and AND2 (N678, N674, N306);
not NOT1 (N679, N664);
and AND4 (N680, N678, N183, N138, N51);
xor XOR2 (N681, N673, N206);
buf BUF1 (N682, N667);
nor NOR2 (N683, N658, N480);
buf BUF1 (N684, N680);
nand NAND3 (N685, N684, N573, N474);
nor NOR3 (N686, N670, N549, N282);
or OR2 (N687, N686, N227);
buf BUF1 (N688, N681);
xor XOR2 (N689, N666, N255);
or OR2 (N690, N676, N15);
not NOT1 (N691, N675);
nand NAND3 (N692, N689, N611, N415);
not NOT1 (N693, N691);
or OR3 (N694, N677, N276, N366);
nand NAND2 (N695, N690, N663);
buf BUF1 (N696, N693);
not NOT1 (N697, N695);
nand NAND2 (N698, N682, N78);
buf BUF1 (N699, N688);
not NOT1 (N700, N692);
not NOT1 (N701, N694);
xor XOR2 (N702, N679, N408);
not NOT1 (N703, N683);
and AND3 (N704, N696, N52, N109);
and AND3 (N705, N703, N499, N176);
nand NAND2 (N706, N699, N579);
or OR2 (N707, N697, N159);
nor NOR2 (N708, N702, N647);
xor XOR2 (N709, N704, N282);
or OR2 (N710, N700, N411);
or OR2 (N711, N708, N408);
nand NAND2 (N712, N698, N501);
not NOT1 (N713, N685);
not NOT1 (N714, N709);
nor NOR4 (N715, N713, N487, N547, N214);
xor XOR2 (N716, N705, N573);
xor XOR2 (N717, N687, N452);
not NOT1 (N718, N710);
xor XOR2 (N719, N701, N274);
and AND4 (N720, N712, N642, N388, N540);
and AND4 (N721, N716, N523, N82, N325);
xor XOR2 (N722, N717, N549);
xor XOR2 (N723, N720, N126);
buf BUF1 (N724, N714);
or OR2 (N725, N721, N683);
not NOT1 (N726, N724);
nand NAND3 (N727, N715, N539, N10);
or OR2 (N728, N722, N198);
and AND3 (N729, N718, N531, N47);
nand NAND2 (N730, N728, N300);
nor NOR4 (N731, N726, N579, N625, N711);
or OR3 (N732, N248, N29, N396);
not NOT1 (N733, N706);
nor NOR4 (N734, N725, N720, N522, N311);
nor NOR3 (N735, N727, N443, N287);
or OR3 (N736, N730, N309, N252);
not NOT1 (N737, N733);
nor NOR4 (N738, N707, N152, N88, N445);
not NOT1 (N739, N719);
and AND4 (N740, N739, N708, N727, N502);
and AND4 (N741, N734, N272, N478, N171);
xor XOR2 (N742, N736, N477);
nor NOR4 (N743, N732, N572, N648, N64);
or OR4 (N744, N741, N33, N443, N21);
and AND2 (N745, N737, N480);
xor XOR2 (N746, N731, N57);
or OR2 (N747, N743, N42);
not NOT1 (N748, N745);
and AND2 (N749, N740, N237);
nor NOR4 (N750, N744, N648, N332, N326);
nand NAND4 (N751, N749, N234, N123, N276);
xor XOR2 (N752, N735, N121);
buf BUF1 (N753, N751);
buf BUF1 (N754, N746);
and AND3 (N755, N754, N534, N53);
or OR4 (N756, N742, N393, N659, N465);
not NOT1 (N757, N747);
and AND3 (N758, N729, N532, N370);
xor XOR2 (N759, N750, N205);
not NOT1 (N760, N757);
xor XOR2 (N761, N748, N396);
and AND3 (N762, N756, N401, N151);
xor XOR2 (N763, N760, N213);
and AND2 (N764, N762, N47);
and AND4 (N765, N755, N647, N181, N415);
and AND4 (N766, N738, N354, N180, N709);
nand NAND2 (N767, N752, N541);
nor NOR4 (N768, N723, N477, N40, N680);
nor NOR3 (N769, N759, N426, N227);
nor NOR3 (N770, N768, N29, N604);
not NOT1 (N771, N769);
nand NAND2 (N772, N766, N214);
and AND2 (N773, N758, N472);
not NOT1 (N774, N765);
not NOT1 (N775, N770);
and AND2 (N776, N764, N655);
and AND2 (N777, N761, N46);
and AND4 (N778, N774, N214, N15, N750);
buf BUF1 (N779, N778);
not NOT1 (N780, N773);
not NOT1 (N781, N779);
or OR4 (N782, N775, N772, N493, N100);
not NOT1 (N783, N156);
nor NOR3 (N784, N771, N234, N776);
nand NAND3 (N785, N754, N736, N784);
or OR4 (N786, N700, N397, N615, N597);
not NOT1 (N787, N753);
buf BUF1 (N788, N777);
xor XOR2 (N789, N781, N551);
nand NAND2 (N790, N789, N94);
xor XOR2 (N791, N785, N264);
not NOT1 (N792, N791);
buf BUF1 (N793, N763);
xor XOR2 (N794, N790, N488);
nor NOR3 (N795, N793, N313, N290);
buf BUF1 (N796, N782);
xor XOR2 (N797, N786, N368);
not NOT1 (N798, N783);
xor XOR2 (N799, N792, N166);
and AND3 (N800, N767, N427, N510);
nor NOR2 (N801, N796, N76);
nor NOR4 (N802, N801, N379, N319, N605);
buf BUF1 (N803, N799);
xor XOR2 (N804, N802, N462);
and AND3 (N805, N804, N528, N499);
buf BUF1 (N806, N800);
or OR4 (N807, N780, N646, N617, N477);
buf BUF1 (N808, N787);
nor NOR2 (N809, N798, N542);
not NOT1 (N810, N807);
and AND2 (N811, N809, N807);
or OR3 (N812, N811, N584, N216);
or OR2 (N813, N794, N727);
and AND3 (N814, N788, N741, N416);
buf BUF1 (N815, N813);
and AND2 (N816, N806, N62);
buf BUF1 (N817, N810);
nor NOR4 (N818, N797, N251, N588, N499);
endmodule