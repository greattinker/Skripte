// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20;

output N3019,N3011,N2990,N3013,N3016,N3017,N3015,N3012,N3009,N3020;

nor NOR2 (N21, N15, N3);
and AND2 (N22, N10, N20);
or OR2 (N23, N3, N19);
not NOT1 (N24, N8);
nand NAND3 (N25, N21, N13, N20);
and AND4 (N26, N24, N17, N18, N21);
nor NOR4 (N27, N12, N19, N20, N7);
nand NAND4 (N28, N7, N3, N25, N3);
buf BUF1 (N29, N5);
not NOT1 (N30, N25);
xor XOR2 (N31, N19, N29);
not NOT1 (N32, N3);
nand NAND3 (N33, N2, N21, N27);
buf BUF1 (N34, N12);
not NOT1 (N35, N1);
buf BUF1 (N36, N32);
buf BUF1 (N37, N23);
and AND4 (N38, N33, N4, N26, N11);
or OR2 (N39, N23, N29);
nor NOR4 (N40, N22, N21, N18, N38);
xor XOR2 (N41, N37, N33);
nand NAND2 (N42, N36, N31);
nor NOR2 (N43, N1, N12);
nand NAND3 (N44, N40, N31, N41);
xor XOR2 (N45, N25, N20);
buf BUF1 (N46, N38);
xor XOR2 (N47, N35, N30);
xor XOR2 (N48, N41, N40);
nand NAND4 (N49, N45, N39, N3, N8);
nor NOR4 (N50, N4, N15, N42, N46);
nand NAND4 (N51, N38, N14, N50, N12);
or OR3 (N52, N13, N3, N10);
xor XOR2 (N53, N37, N33);
xor XOR2 (N54, N43, N18);
nand NAND4 (N55, N48, N3, N15, N52);
xor XOR2 (N56, N21, N29);
nand NAND4 (N57, N47, N29, N30, N13);
or OR4 (N58, N49, N5, N41, N52);
xor XOR2 (N59, N57, N7);
nor NOR4 (N60, N58, N4, N23, N17);
and AND4 (N61, N54, N23, N2, N24);
nor NOR2 (N62, N59, N32);
and AND3 (N63, N62, N35, N51);
xor XOR2 (N64, N42, N20);
or OR3 (N65, N34, N36, N63);
nor NOR2 (N66, N50, N11);
buf BUF1 (N67, N64);
xor XOR2 (N68, N67, N26);
not NOT1 (N69, N55);
nor NOR2 (N70, N69, N39);
nand NAND2 (N71, N56, N68);
not NOT1 (N72, N71);
buf BUF1 (N73, N18);
or OR2 (N74, N73, N32);
xor XOR2 (N75, N66, N65);
not NOT1 (N76, N16);
nor NOR4 (N77, N76, N34, N69, N3);
or OR3 (N78, N70, N6, N35);
nor NOR3 (N79, N61, N43, N59);
buf BUF1 (N80, N78);
not NOT1 (N81, N75);
and AND3 (N82, N72, N15, N71);
xor XOR2 (N83, N77, N28);
not NOT1 (N84, N44);
not NOT1 (N85, N12);
nand NAND3 (N86, N82, N10, N11);
nand NAND4 (N87, N84, N69, N36, N13);
not NOT1 (N88, N87);
not NOT1 (N89, N53);
buf BUF1 (N90, N80);
nand NAND3 (N91, N86, N43, N24);
nand NAND4 (N92, N83, N19, N74, N60);
not NOT1 (N93, N74);
buf BUF1 (N94, N3);
xor XOR2 (N95, N85, N29);
nor NOR2 (N96, N91, N56);
nand NAND3 (N97, N89, N35, N81);
buf BUF1 (N98, N80);
nor NOR2 (N99, N92, N18);
buf BUF1 (N100, N93);
xor XOR2 (N101, N90, N36);
not NOT1 (N102, N94);
xor XOR2 (N103, N100, N66);
nand NAND3 (N104, N99, N61, N83);
not NOT1 (N105, N102);
nor NOR2 (N106, N97, N31);
and AND4 (N107, N106, N36, N75, N95);
nand NAND4 (N108, N98, N67, N18, N7);
buf BUF1 (N109, N99);
not NOT1 (N110, N108);
not NOT1 (N111, N104);
nor NOR4 (N112, N103, N99, N18, N49);
buf BUF1 (N113, N111);
nand NAND4 (N114, N105, N107, N68, N14);
or OR4 (N115, N33, N83, N80, N28);
xor XOR2 (N116, N109, N57);
nor NOR2 (N117, N101, N23);
xor XOR2 (N118, N88, N53);
xor XOR2 (N119, N110, N88);
and AND2 (N120, N117, N21);
and AND2 (N121, N116, N34);
buf BUF1 (N122, N120);
nor NOR3 (N123, N112, N42, N35);
not NOT1 (N124, N122);
and AND2 (N125, N124, N56);
xor XOR2 (N126, N121, N101);
nand NAND2 (N127, N119, N117);
not NOT1 (N128, N125);
nor NOR4 (N129, N127, N33, N110, N125);
not NOT1 (N130, N115);
and AND3 (N131, N114, N98, N110);
buf BUF1 (N132, N123);
or OR3 (N133, N118, N54, N122);
nand NAND4 (N134, N79, N92, N86, N62);
nand NAND2 (N135, N129, N33);
not NOT1 (N136, N133);
nand NAND2 (N137, N131, N89);
xor XOR2 (N138, N113, N82);
or OR4 (N139, N137, N105, N20, N7);
and AND2 (N140, N132, N138);
nand NAND3 (N141, N64, N5, N125);
not NOT1 (N142, N140);
not NOT1 (N143, N139);
nand NAND4 (N144, N130, N47, N118, N53);
xor XOR2 (N145, N142, N41);
nor NOR4 (N146, N141, N86, N125, N41);
buf BUF1 (N147, N128);
buf BUF1 (N148, N96);
xor XOR2 (N149, N126, N69);
nand NAND2 (N150, N143, N84);
not NOT1 (N151, N149);
or OR3 (N152, N146, N83, N68);
nor NOR2 (N153, N147, N15);
buf BUF1 (N154, N153);
nand NAND3 (N155, N134, N73, N109);
or OR3 (N156, N154, N76, N54);
nor NOR2 (N157, N155, N18);
nand NAND2 (N158, N152, N126);
and AND3 (N159, N145, N99, N5);
and AND3 (N160, N135, N63, N121);
xor XOR2 (N161, N158, N82);
nor NOR3 (N162, N136, N71, N31);
not NOT1 (N163, N150);
or OR3 (N164, N144, N36, N73);
nand NAND4 (N165, N161, N115, N84, N68);
not NOT1 (N166, N159);
and AND2 (N167, N164, N74);
not NOT1 (N168, N151);
nand NAND4 (N169, N167, N164, N102, N113);
or OR3 (N170, N148, N6, N124);
buf BUF1 (N171, N166);
and AND2 (N172, N163, N87);
or OR4 (N173, N169, N122, N145, N96);
and AND3 (N174, N157, N26, N30);
xor XOR2 (N175, N160, N127);
and AND2 (N176, N162, N85);
xor XOR2 (N177, N170, N54);
xor XOR2 (N178, N175, N99);
buf BUF1 (N179, N165);
and AND3 (N180, N176, N100, N146);
xor XOR2 (N181, N171, N118);
xor XOR2 (N182, N156, N49);
xor XOR2 (N183, N180, N6);
or OR4 (N184, N177, N16, N155, N17);
not NOT1 (N185, N174);
nor NOR3 (N186, N181, N43, N7);
not NOT1 (N187, N168);
nor NOR4 (N188, N178, N91, N20, N108);
buf BUF1 (N189, N188);
or OR3 (N190, N179, N93, N53);
or OR3 (N191, N185, N104, N102);
or OR4 (N192, N190, N179, N175, N6);
buf BUF1 (N193, N186);
nor NOR4 (N194, N193, N156, N82, N193);
xor XOR2 (N195, N189, N89);
not NOT1 (N196, N172);
buf BUF1 (N197, N192);
not NOT1 (N198, N182);
xor XOR2 (N199, N184, N41);
and AND2 (N200, N183, N126);
and AND2 (N201, N173, N121);
or OR4 (N202, N195, N76, N136, N27);
xor XOR2 (N203, N187, N147);
nor NOR3 (N204, N199, N24, N153);
nor NOR2 (N205, N194, N182);
nor NOR4 (N206, N200, N96, N94, N67);
xor XOR2 (N207, N197, N60);
xor XOR2 (N208, N201, N186);
buf BUF1 (N209, N198);
and AND2 (N210, N207, N36);
nand NAND4 (N211, N209, N57, N3, N109);
and AND3 (N212, N210, N32, N167);
buf BUF1 (N213, N206);
and AND2 (N214, N211, N62);
nor NOR3 (N215, N204, N173, N10);
nand NAND4 (N216, N196, N167, N181, N152);
nand NAND4 (N217, N191, N10, N26, N210);
xor XOR2 (N218, N208, N87);
or OR4 (N219, N217, N36, N17, N181);
and AND3 (N220, N214, N85, N86);
not NOT1 (N221, N215);
buf BUF1 (N222, N220);
or OR2 (N223, N213, N126);
nor NOR3 (N224, N212, N184, N128);
nor NOR2 (N225, N222, N140);
xor XOR2 (N226, N202, N209);
not NOT1 (N227, N219);
not NOT1 (N228, N203);
buf BUF1 (N229, N227);
nor NOR2 (N230, N221, N186);
not NOT1 (N231, N228);
xor XOR2 (N232, N218, N7);
nand NAND3 (N233, N216, N216, N146);
xor XOR2 (N234, N223, N19);
nor NOR4 (N235, N229, N204, N215, N225);
xor XOR2 (N236, N219, N38);
or OR3 (N237, N233, N172, N219);
nor NOR2 (N238, N236, N79);
and AND4 (N239, N230, N202, N171, N155);
and AND2 (N240, N239, N206);
and AND3 (N241, N235, N159, N120);
not NOT1 (N242, N232);
nor NOR2 (N243, N240, N110);
and AND2 (N244, N238, N6);
buf BUF1 (N245, N241);
nor NOR4 (N246, N245, N142, N233, N151);
nor NOR2 (N247, N237, N50);
nand NAND3 (N248, N242, N31, N146);
nand NAND2 (N249, N226, N15);
and AND3 (N250, N249, N88, N47);
not NOT1 (N251, N244);
and AND3 (N252, N248, N218, N245);
and AND3 (N253, N252, N157, N61);
and AND2 (N254, N234, N156);
nor NOR2 (N255, N205, N192);
not NOT1 (N256, N243);
xor XOR2 (N257, N253, N103);
nor NOR4 (N258, N251, N257, N171, N161);
or OR3 (N259, N75, N238, N30);
not NOT1 (N260, N231);
or OR3 (N261, N250, N223, N111);
not NOT1 (N262, N261);
nor NOR2 (N263, N258, N262);
or OR3 (N264, N254, N246, N27);
or OR4 (N265, N228, N121, N82, N40);
xor XOR2 (N266, N96, N138);
not NOT1 (N267, N259);
nor NOR2 (N268, N247, N217);
not NOT1 (N269, N255);
not NOT1 (N270, N266);
and AND3 (N271, N260, N96, N232);
xor XOR2 (N272, N264, N137);
xor XOR2 (N273, N270, N189);
not NOT1 (N274, N272);
not NOT1 (N275, N263);
xor XOR2 (N276, N265, N236);
and AND3 (N277, N271, N128, N239);
buf BUF1 (N278, N273);
or OR2 (N279, N268, N40);
and AND2 (N280, N256, N220);
not NOT1 (N281, N276);
or OR3 (N282, N275, N127, N157);
not NOT1 (N283, N281);
nor NOR2 (N284, N280, N126);
not NOT1 (N285, N282);
xor XOR2 (N286, N284, N109);
or OR3 (N287, N224, N238, N221);
buf BUF1 (N288, N283);
or OR2 (N289, N274, N266);
and AND2 (N290, N286, N98);
nor NOR4 (N291, N277, N169, N130, N256);
buf BUF1 (N292, N267);
xor XOR2 (N293, N287, N274);
nand NAND2 (N294, N292, N276);
nand NAND4 (N295, N278, N106, N58, N6);
xor XOR2 (N296, N285, N39);
buf BUF1 (N297, N293);
buf BUF1 (N298, N291);
buf BUF1 (N299, N294);
buf BUF1 (N300, N290);
xor XOR2 (N301, N269, N163);
nor NOR3 (N302, N300, N11, N86);
or OR4 (N303, N279, N255, N290, N105);
or OR2 (N304, N296, N43);
xor XOR2 (N305, N289, N63);
and AND3 (N306, N298, N188, N195);
or OR3 (N307, N297, N97, N224);
not NOT1 (N308, N299);
or OR2 (N309, N307, N305);
not NOT1 (N310, N246);
and AND3 (N311, N309, N163, N219);
or OR4 (N312, N303, N283, N212, N255);
nor NOR2 (N313, N288, N48);
nor NOR3 (N314, N312, N112, N301);
and AND4 (N315, N131, N149, N222, N226);
or OR3 (N316, N295, N241, N152);
not NOT1 (N317, N310);
nor NOR4 (N318, N314, N280, N303, N93);
and AND4 (N319, N313, N57, N103, N120);
xor XOR2 (N320, N308, N211);
nor NOR4 (N321, N302, N247, N108, N297);
nor NOR3 (N322, N321, N303, N57);
xor XOR2 (N323, N322, N154);
xor XOR2 (N324, N318, N300);
not NOT1 (N325, N304);
and AND4 (N326, N325, N53, N193, N278);
buf BUF1 (N327, N306);
xor XOR2 (N328, N319, N107);
buf BUF1 (N329, N323);
not NOT1 (N330, N327);
xor XOR2 (N331, N315, N266);
xor XOR2 (N332, N328, N300);
nor NOR4 (N333, N316, N117, N113, N119);
and AND3 (N334, N331, N145, N320);
xor XOR2 (N335, N240, N17);
and AND3 (N336, N324, N309, N291);
buf BUF1 (N337, N326);
and AND3 (N338, N330, N231, N128);
xor XOR2 (N339, N333, N52);
nand NAND2 (N340, N311, N106);
buf BUF1 (N341, N337);
buf BUF1 (N342, N329);
buf BUF1 (N343, N317);
nor NOR2 (N344, N343, N253);
not NOT1 (N345, N341);
nand NAND4 (N346, N339, N112, N172, N257);
not NOT1 (N347, N346);
and AND3 (N348, N332, N134, N323);
xor XOR2 (N349, N342, N130);
xor XOR2 (N350, N347, N64);
nor NOR3 (N351, N350, N320, N239);
or OR2 (N352, N351, N292);
nor NOR3 (N353, N349, N104, N190);
and AND3 (N354, N345, N325, N205);
and AND3 (N355, N340, N148, N157);
and AND2 (N356, N348, N125);
xor XOR2 (N357, N344, N83);
xor XOR2 (N358, N335, N106);
and AND3 (N359, N357, N174, N135);
xor XOR2 (N360, N354, N134);
not NOT1 (N361, N352);
nor NOR3 (N362, N359, N12, N274);
not NOT1 (N363, N358);
and AND3 (N364, N353, N231, N243);
nor NOR4 (N365, N362, N124, N337, N265);
buf BUF1 (N366, N334);
or OR4 (N367, N361, N237, N179, N62);
nand NAND3 (N368, N366, N230, N226);
and AND4 (N369, N365, N289, N121, N50);
or OR3 (N370, N355, N282, N256);
buf BUF1 (N371, N336);
and AND3 (N372, N363, N199, N9);
not NOT1 (N373, N338);
not NOT1 (N374, N368);
not NOT1 (N375, N372);
buf BUF1 (N376, N364);
nor NOR2 (N377, N367, N287);
nor NOR2 (N378, N377, N314);
not NOT1 (N379, N376);
or OR2 (N380, N370, N132);
xor XOR2 (N381, N380, N68);
not NOT1 (N382, N374);
buf BUF1 (N383, N382);
or OR2 (N384, N369, N328);
and AND4 (N385, N381, N182, N384, N245);
buf BUF1 (N386, N216);
nor NOR4 (N387, N378, N310, N42, N286);
buf BUF1 (N388, N387);
buf BUF1 (N389, N375);
or OR3 (N390, N389, N187, N163);
not NOT1 (N391, N379);
not NOT1 (N392, N388);
xor XOR2 (N393, N383, N298);
xor XOR2 (N394, N356, N173);
nand NAND4 (N395, N393, N385, N168, N74);
xor XOR2 (N396, N297, N26);
xor XOR2 (N397, N373, N207);
buf BUF1 (N398, N394);
and AND2 (N399, N371, N222);
xor XOR2 (N400, N386, N304);
and AND2 (N401, N397, N263);
buf BUF1 (N402, N392);
xor XOR2 (N403, N400, N32);
not NOT1 (N404, N395);
nand NAND2 (N405, N398, N281);
not NOT1 (N406, N390);
nor NOR4 (N407, N360, N353, N177, N243);
nor NOR3 (N408, N396, N380, N348);
xor XOR2 (N409, N391, N283);
and AND2 (N410, N399, N187);
xor XOR2 (N411, N402, N385);
not NOT1 (N412, N407);
xor XOR2 (N413, N406, N287);
not NOT1 (N414, N412);
nor NOR4 (N415, N413, N118, N79, N368);
not NOT1 (N416, N405);
buf BUF1 (N417, N401);
or OR3 (N418, N414, N362, N255);
and AND3 (N419, N408, N346, N395);
xor XOR2 (N420, N419, N149);
nand NAND4 (N421, N403, N110, N67, N234);
or OR3 (N422, N409, N63, N157);
nor NOR4 (N423, N422, N268, N339, N261);
or OR3 (N424, N411, N129, N372);
nor NOR2 (N425, N420, N111);
not NOT1 (N426, N404);
xor XOR2 (N427, N410, N362);
nand NAND3 (N428, N417, N336, N378);
nor NOR3 (N429, N418, N338, N16);
xor XOR2 (N430, N428, N422);
nor NOR2 (N431, N429, N369);
not NOT1 (N432, N423);
xor XOR2 (N433, N421, N232);
or OR2 (N434, N427, N412);
or OR3 (N435, N434, N336, N88);
nand NAND3 (N436, N431, N399, N275);
buf BUF1 (N437, N415);
nor NOR4 (N438, N416, N301, N304, N119);
nand NAND2 (N439, N426, N291);
not NOT1 (N440, N433);
and AND3 (N441, N439, N308, N116);
buf BUF1 (N442, N441);
xor XOR2 (N443, N432, N222);
nand NAND3 (N444, N438, N139, N331);
and AND4 (N445, N443, N183, N116, N305);
buf BUF1 (N446, N435);
buf BUF1 (N447, N442);
buf BUF1 (N448, N447);
not NOT1 (N449, N445);
and AND3 (N450, N430, N333, N437);
or OR3 (N451, N82, N164, N364);
nor NOR2 (N452, N451, N96);
buf BUF1 (N453, N449);
not NOT1 (N454, N452);
or OR3 (N455, N444, N140, N101);
not NOT1 (N456, N453);
and AND3 (N457, N440, N199, N257);
nor NOR3 (N458, N425, N129, N428);
nor NOR4 (N459, N436, N140, N126, N106);
nor NOR2 (N460, N424, N116);
not NOT1 (N461, N456);
xor XOR2 (N462, N458, N142);
nor NOR3 (N463, N455, N445, N231);
and AND4 (N464, N457, N169, N57, N376);
xor XOR2 (N465, N450, N304);
nand NAND2 (N466, N459, N357);
nor NOR2 (N467, N466, N352);
nor NOR2 (N468, N448, N343);
nor NOR2 (N469, N454, N184);
nand NAND4 (N470, N463, N392, N329, N330);
nand NAND2 (N471, N462, N141);
and AND2 (N472, N465, N397);
buf BUF1 (N473, N467);
or OR4 (N474, N472, N289, N436, N119);
not NOT1 (N475, N471);
nor NOR2 (N476, N473, N255);
nand NAND4 (N477, N474, N123, N210, N218);
nor NOR2 (N478, N477, N143);
xor XOR2 (N479, N461, N119);
nand NAND4 (N480, N469, N109, N354, N439);
nand NAND2 (N481, N478, N202);
xor XOR2 (N482, N460, N188);
buf BUF1 (N483, N475);
xor XOR2 (N484, N468, N373);
or OR3 (N485, N480, N215, N418);
buf BUF1 (N486, N485);
or OR4 (N487, N476, N441, N37, N54);
nor NOR3 (N488, N481, N382, N82);
buf BUF1 (N489, N482);
xor XOR2 (N490, N486, N288);
nand NAND4 (N491, N464, N15, N201, N178);
xor XOR2 (N492, N488, N104);
nand NAND3 (N493, N479, N275, N90);
not NOT1 (N494, N492);
or OR4 (N495, N489, N186, N180, N471);
not NOT1 (N496, N494);
nor NOR3 (N497, N490, N248, N69);
nor NOR3 (N498, N497, N277, N389);
not NOT1 (N499, N470);
or OR2 (N500, N491, N322);
or OR3 (N501, N496, N35, N296);
and AND4 (N502, N493, N59, N176, N219);
or OR2 (N503, N484, N409);
not NOT1 (N504, N446);
not NOT1 (N505, N499);
and AND4 (N506, N487, N137, N83, N361);
xor XOR2 (N507, N504, N193);
and AND4 (N508, N501, N468, N54, N302);
and AND3 (N509, N505, N327, N55);
xor XOR2 (N510, N502, N353);
nor NOR3 (N511, N495, N498, N158);
xor XOR2 (N512, N410, N127);
and AND4 (N513, N500, N425, N421, N316);
not NOT1 (N514, N506);
nand NAND4 (N515, N512, N378, N127, N98);
nand NAND3 (N516, N508, N65, N263);
buf BUF1 (N517, N510);
and AND4 (N518, N514, N499, N485, N33);
or OR2 (N519, N515, N508);
not NOT1 (N520, N519);
nand NAND2 (N521, N503, N59);
xor XOR2 (N522, N507, N206);
xor XOR2 (N523, N516, N143);
or OR4 (N524, N523, N446, N19, N486);
nand NAND2 (N525, N511, N16);
not NOT1 (N526, N518);
buf BUF1 (N527, N509);
buf BUF1 (N528, N526);
nor NOR3 (N529, N521, N129, N112);
not NOT1 (N530, N513);
or OR4 (N531, N517, N369, N368, N409);
xor XOR2 (N532, N529, N165);
nor NOR2 (N533, N531, N419);
or OR4 (N534, N527, N13, N284, N277);
and AND3 (N535, N522, N246, N509);
buf BUF1 (N536, N520);
not NOT1 (N537, N483);
not NOT1 (N538, N525);
not NOT1 (N539, N530);
or OR4 (N540, N533, N263, N64, N497);
nand NAND3 (N541, N540, N107, N388);
nand NAND2 (N542, N534, N226);
and AND3 (N543, N524, N30, N259);
nor NOR4 (N544, N538, N414, N195, N207);
nor NOR4 (N545, N535, N394, N446, N154);
or OR2 (N546, N545, N456);
or OR3 (N547, N532, N426, N460);
or OR4 (N548, N547, N401, N255, N51);
and AND2 (N549, N543, N25);
buf BUF1 (N550, N544);
nand NAND2 (N551, N546, N237);
nand NAND4 (N552, N549, N295, N333, N337);
buf BUF1 (N553, N541);
not NOT1 (N554, N539);
and AND4 (N555, N553, N156, N354, N155);
or OR4 (N556, N554, N220, N199, N528);
and AND4 (N557, N104, N101, N184, N147);
buf BUF1 (N558, N542);
and AND4 (N559, N548, N75, N8, N201);
or OR2 (N560, N537, N177);
nand NAND4 (N561, N560, N191, N202, N269);
or OR4 (N562, N555, N374, N442, N5);
and AND3 (N563, N556, N33, N246);
and AND3 (N564, N562, N506, N535);
nor NOR2 (N565, N559, N393);
not NOT1 (N566, N563);
or OR4 (N567, N564, N131, N416, N193);
or OR2 (N568, N561, N189);
xor XOR2 (N569, N552, N485);
not NOT1 (N570, N551);
xor XOR2 (N571, N565, N59);
not NOT1 (N572, N569);
nand NAND2 (N573, N536, N402);
buf BUF1 (N574, N567);
nor NOR2 (N575, N566, N224);
or OR4 (N576, N573, N32, N187, N21);
nand NAND4 (N577, N550, N391, N416, N204);
not NOT1 (N578, N570);
nand NAND3 (N579, N557, N26, N401);
not NOT1 (N580, N577);
and AND3 (N581, N574, N371, N137);
xor XOR2 (N582, N579, N501);
or OR2 (N583, N580, N516);
nor NOR3 (N584, N582, N555, N321);
and AND4 (N585, N576, N302, N388, N197);
nand NAND4 (N586, N581, N58, N437, N398);
xor XOR2 (N587, N572, N3);
nand NAND2 (N588, N587, N481);
and AND2 (N589, N588, N16);
xor XOR2 (N590, N568, N186);
not NOT1 (N591, N589);
and AND4 (N592, N558, N50, N252, N110);
and AND4 (N593, N584, N428, N411, N555);
not NOT1 (N594, N585);
buf BUF1 (N595, N591);
and AND4 (N596, N571, N519, N378, N81);
xor XOR2 (N597, N575, N102);
nand NAND3 (N598, N595, N115, N435);
buf BUF1 (N599, N586);
buf BUF1 (N600, N596);
nand NAND2 (N601, N583, N468);
not NOT1 (N602, N598);
and AND3 (N603, N600, N328, N115);
or OR2 (N604, N599, N171);
not NOT1 (N605, N601);
not NOT1 (N606, N597);
nor NOR4 (N607, N603, N474, N261, N6);
not NOT1 (N608, N593);
and AND2 (N609, N604, N247);
not NOT1 (N610, N578);
not NOT1 (N611, N605);
xor XOR2 (N612, N611, N524);
and AND4 (N613, N607, N207, N138, N176);
and AND4 (N614, N608, N2, N61, N307);
xor XOR2 (N615, N610, N407);
nand NAND3 (N616, N609, N256, N551);
nor NOR3 (N617, N606, N483, N57);
or OR4 (N618, N594, N584, N78, N574);
and AND4 (N619, N590, N293, N602, N170);
and AND3 (N620, N20, N114, N91);
buf BUF1 (N621, N614);
nand NAND2 (N622, N615, N162);
not NOT1 (N623, N618);
xor XOR2 (N624, N622, N523);
not NOT1 (N625, N617);
buf BUF1 (N626, N620);
xor XOR2 (N627, N612, N53);
and AND4 (N628, N619, N581, N401, N91);
not NOT1 (N629, N624);
buf BUF1 (N630, N629);
nand NAND3 (N631, N592, N507, N289);
or OR3 (N632, N630, N353, N227);
and AND3 (N633, N621, N156, N294);
nor NOR4 (N634, N626, N55, N44, N299);
or OR2 (N635, N627, N388);
nand NAND4 (N636, N633, N444, N114, N418);
and AND2 (N637, N631, N406);
xor XOR2 (N638, N635, N266);
buf BUF1 (N639, N638);
and AND2 (N640, N637, N168);
nand NAND3 (N641, N632, N100, N2);
buf BUF1 (N642, N641);
nand NAND2 (N643, N623, N527);
nor NOR4 (N644, N639, N210, N495, N400);
xor XOR2 (N645, N640, N612);
nand NAND4 (N646, N628, N432, N84, N40);
not NOT1 (N647, N646);
or OR2 (N648, N647, N25);
not NOT1 (N649, N644);
or OR4 (N650, N642, N481, N106, N54);
not NOT1 (N651, N645);
nor NOR4 (N652, N643, N523, N64, N631);
or OR2 (N653, N616, N154);
nor NOR3 (N654, N649, N389, N240);
buf BUF1 (N655, N650);
and AND2 (N656, N613, N347);
not NOT1 (N657, N652);
buf BUF1 (N658, N648);
or OR2 (N659, N634, N371);
nor NOR2 (N660, N655, N486);
not NOT1 (N661, N659);
not NOT1 (N662, N651);
or OR2 (N663, N625, N654);
not NOT1 (N664, N515);
or OR2 (N665, N662, N67);
xor XOR2 (N666, N653, N256);
buf BUF1 (N667, N656);
xor XOR2 (N668, N667, N272);
and AND3 (N669, N666, N316, N98);
or OR2 (N670, N657, N22);
nor NOR4 (N671, N669, N542, N458, N218);
xor XOR2 (N672, N668, N563);
nor NOR2 (N673, N636, N211);
nor NOR4 (N674, N673, N56, N180, N399);
or OR4 (N675, N671, N366, N4, N592);
nor NOR4 (N676, N665, N197, N132, N200);
xor XOR2 (N677, N661, N625);
buf BUF1 (N678, N658);
xor XOR2 (N679, N675, N180);
xor XOR2 (N680, N679, N238);
buf BUF1 (N681, N680);
or OR2 (N682, N660, N247);
or OR4 (N683, N664, N351, N231, N543);
and AND4 (N684, N674, N195, N479, N67);
xor XOR2 (N685, N682, N162);
nand NAND2 (N686, N663, N18);
nor NOR2 (N687, N686, N640);
or OR3 (N688, N684, N495, N484);
nand NAND2 (N689, N672, N675);
not NOT1 (N690, N676);
buf BUF1 (N691, N690);
and AND3 (N692, N677, N335, N372);
xor XOR2 (N693, N689, N43);
and AND3 (N694, N681, N32, N618);
buf BUF1 (N695, N692);
nor NOR4 (N696, N691, N314, N137, N483);
nor NOR4 (N697, N695, N449, N594, N309);
and AND4 (N698, N694, N20, N336, N480);
nor NOR4 (N699, N697, N72, N79, N611);
and AND4 (N700, N685, N506, N463, N411);
nand NAND4 (N701, N678, N655, N343, N302);
buf BUF1 (N702, N670);
xor XOR2 (N703, N687, N315);
xor XOR2 (N704, N700, N139);
nor NOR4 (N705, N704, N484, N107, N671);
nor NOR2 (N706, N703, N519);
nand NAND2 (N707, N698, N618);
nor NOR2 (N708, N706, N31);
buf BUF1 (N709, N683);
buf BUF1 (N710, N696);
buf BUF1 (N711, N702);
not NOT1 (N712, N711);
nor NOR4 (N713, N705, N338, N692, N506);
nor NOR4 (N714, N709, N222, N386, N421);
or OR2 (N715, N712, N542);
and AND4 (N716, N708, N266, N258, N285);
buf BUF1 (N717, N714);
nor NOR3 (N718, N716, N121, N562);
and AND2 (N719, N693, N385);
and AND3 (N720, N707, N328, N582);
buf BUF1 (N721, N715);
not NOT1 (N722, N699);
and AND4 (N723, N701, N661, N538, N238);
and AND4 (N724, N717, N527, N686, N32);
xor XOR2 (N725, N688, N620);
nor NOR2 (N726, N723, N353);
not NOT1 (N727, N721);
or OR4 (N728, N720, N538, N488, N414);
nor NOR2 (N729, N724, N698);
xor XOR2 (N730, N726, N428);
nand NAND4 (N731, N719, N209, N588, N220);
or OR2 (N732, N728, N417);
nand NAND4 (N733, N730, N48, N466, N549);
xor XOR2 (N734, N725, N585);
or OR4 (N735, N722, N531, N76, N6);
nor NOR4 (N736, N733, N435, N443, N453);
nand NAND3 (N737, N718, N380, N120);
nand NAND3 (N738, N710, N93, N377);
nor NOR3 (N739, N731, N254, N356);
buf BUF1 (N740, N737);
nand NAND4 (N741, N729, N553, N351, N622);
and AND4 (N742, N713, N148, N381, N178);
or OR3 (N743, N738, N533, N317);
and AND2 (N744, N736, N482);
or OR2 (N745, N732, N524);
or OR2 (N746, N743, N445);
xor XOR2 (N747, N744, N321);
nor NOR4 (N748, N735, N127, N592, N246);
buf BUF1 (N749, N747);
and AND2 (N750, N745, N348);
or OR3 (N751, N749, N233, N242);
xor XOR2 (N752, N751, N91);
buf BUF1 (N753, N752);
xor XOR2 (N754, N746, N439);
and AND3 (N755, N748, N451, N230);
nand NAND3 (N756, N750, N308, N576);
or OR2 (N757, N754, N529);
nor NOR4 (N758, N727, N406, N506, N236);
nand NAND4 (N759, N742, N61, N255, N144);
and AND2 (N760, N759, N280);
xor XOR2 (N761, N755, N461);
and AND4 (N762, N758, N81, N242, N681);
xor XOR2 (N763, N739, N182);
not NOT1 (N764, N740);
xor XOR2 (N765, N756, N719);
buf BUF1 (N766, N762);
nor NOR4 (N767, N763, N394, N305, N297);
buf BUF1 (N768, N760);
or OR3 (N769, N753, N3, N325);
xor XOR2 (N770, N757, N81);
buf BUF1 (N771, N761);
nand NAND3 (N772, N770, N391, N319);
and AND3 (N773, N741, N391, N188);
and AND4 (N774, N773, N733, N136, N166);
nand NAND3 (N775, N766, N392, N512);
xor XOR2 (N776, N768, N675);
or OR2 (N777, N769, N89);
and AND3 (N778, N771, N760, N16);
or OR3 (N779, N778, N117, N745);
or OR3 (N780, N767, N115, N588);
xor XOR2 (N781, N765, N134);
or OR2 (N782, N774, N550);
not NOT1 (N783, N776);
buf BUF1 (N784, N781);
nand NAND2 (N785, N783, N221);
and AND3 (N786, N782, N154, N211);
nor NOR3 (N787, N780, N435, N104);
or OR2 (N788, N777, N145);
nand NAND2 (N789, N764, N203);
or OR3 (N790, N734, N448, N495);
nor NOR3 (N791, N775, N161, N596);
nand NAND3 (N792, N786, N596, N441);
nor NOR2 (N793, N792, N753);
or OR4 (N794, N787, N314, N49, N236);
or OR2 (N795, N793, N444);
xor XOR2 (N796, N791, N329);
xor XOR2 (N797, N789, N334);
xor XOR2 (N798, N795, N699);
buf BUF1 (N799, N796);
xor XOR2 (N800, N772, N309);
and AND3 (N801, N794, N710, N682);
not NOT1 (N802, N790);
xor XOR2 (N803, N788, N536);
and AND4 (N804, N784, N43, N479, N116);
xor XOR2 (N805, N803, N532);
buf BUF1 (N806, N785);
and AND4 (N807, N806, N494, N275, N795);
not NOT1 (N808, N805);
nor NOR4 (N809, N797, N635, N313, N326);
or OR2 (N810, N804, N656);
buf BUF1 (N811, N800);
nor NOR3 (N812, N811, N170, N761);
or OR4 (N813, N810, N214, N660, N335);
not NOT1 (N814, N808);
nor NOR2 (N815, N812, N40);
or OR2 (N816, N815, N814);
and AND2 (N817, N484, N4);
xor XOR2 (N818, N817, N508);
or OR4 (N819, N801, N528, N427, N55);
or OR2 (N820, N813, N769);
nor NOR3 (N821, N799, N233, N773);
nor NOR4 (N822, N816, N152, N754, N78);
not NOT1 (N823, N819);
xor XOR2 (N824, N820, N685);
and AND2 (N825, N824, N766);
or OR4 (N826, N802, N169, N165, N129);
nor NOR4 (N827, N807, N89, N757, N484);
nand NAND4 (N828, N826, N820, N453, N176);
xor XOR2 (N829, N798, N767);
not NOT1 (N830, N827);
nor NOR3 (N831, N809, N212, N311);
nor NOR3 (N832, N831, N395, N471);
xor XOR2 (N833, N832, N110);
or OR2 (N834, N821, N700);
nand NAND4 (N835, N829, N342, N301, N754);
not NOT1 (N836, N834);
xor XOR2 (N837, N836, N693);
xor XOR2 (N838, N825, N64);
or OR3 (N839, N833, N552, N403);
buf BUF1 (N840, N823);
and AND3 (N841, N779, N839, N105);
not NOT1 (N842, N18);
nor NOR3 (N843, N835, N459, N744);
buf BUF1 (N844, N842);
xor XOR2 (N845, N843, N194);
nor NOR4 (N846, N828, N421, N533, N577);
buf BUF1 (N847, N840);
xor XOR2 (N848, N838, N39);
xor XOR2 (N849, N822, N805);
nand NAND3 (N850, N830, N423, N542);
or OR2 (N851, N848, N715);
or OR3 (N852, N846, N797, N83);
or OR3 (N853, N847, N419, N295);
nand NAND4 (N854, N837, N230, N695, N317);
xor XOR2 (N855, N852, N676);
and AND2 (N856, N850, N103);
nand NAND3 (N857, N854, N340, N638);
buf BUF1 (N858, N841);
or OR3 (N859, N818, N442, N483);
not NOT1 (N860, N856);
nor NOR4 (N861, N855, N27, N786, N548);
not NOT1 (N862, N851);
not NOT1 (N863, N849);
not NOT1 (N864, N862);
or OR3 (N865, N853, N105, N129);
and AND4 (N866, N860, N513, N806, N134);
nor NOR4 (N867, N866, N818, N13, N412);
buf BUF1 (N868, N863);
xor XOR2 (N869, N868, N766);
xor XOR2 (N870, N867, N691);
not NOT1 (N871, N857);
nor NOR3 (N872, N864, N347, N245);
not NOT1 (N873, N861);
and AND4 (N874, N845, N19, N476, N799);
or OR4 (N875, N869, N182, N170, N874);
and AND4 (N876, N388, N512, N77, N831);
buf BUF1 (N877, N871);
buf BUF1 (N878, N872);
nor NOR3 (N879, N858, N614, N646);
nor NOR2 (N880, N870, N311);
buf BUF1 (N881, N876);
nand NAND3 (N882, N879, N353, N681);
or OR2 (N883, N865, N374);
nor NOR2 (N884, N875, N407);
or OR4 (N885, N877, N21, N863, N493);
xor XOR2 (N886, N873, N33);
buf BUF1 (N887, N886);
and AND4 (N888, N878, N37, N863, N74);
and AND3 (N889, N882, N430, N60);
or OR2 (N890, N887, N551);
or OR3 (N891, N889, N598, N58);
not NOT1 (N892, N885);
xor XOR2 (N893, N890, N217);
and AND2 (N894, N859, N305);
buf BUF1 (N895, N884);
buf BUF1 (N896, N844);
or OR3 (N897, N880, N154, N360);
and AND3 (N898, N891, N282, N145);
and AND2 (N899, N892, N152);
or OR4 (N900, N888, N414, N116, N775);
and AND2 (N901, N899, N143);
and AND4 (N902, N901, N182, N753, N469);
and AND3 (N903, N897, N406, N381);
or OR3 (N904, N902, N231, N367);
xor XOR2 (N905, N898, N183);
xor XOR2 (N906, N895, N703);
not NOT1 (N907, N904);
nand NAND2 (N908, N893, N20);
xor XOR2 (N909, N896, N682);
buf BUF1 (N910, N908);
buf BUF1 (N911, N905);
and AND4 (N912, N906, N842, N271, N417);
not NOT1 (N913, N881);
buf BUF1 (N914, N894);
not NOT1 (N915, N883);
not NOT1 (N916, N911);
not NOT1 (N917, N915);
xor XOR2 (N918, N907, N16);
xor XOR2 (N919, N909, N802);
or OR3 (N920, N900, N685, N692);
or OR2 (N921, N910, N455);
nand NAND2 (N922, N916, N751);
and AND4 (N923, N919, N308, N291, N153);
nor NOR4 (N924, N918, N115, N670, N817);
xor XOR2 (N925, N917, N785);
xor XOR2 (N926, N912, N267);
or OR2 (N927, N926, N356);
and AND4 (N928, N925, N672, N780, N846);
buf BUF1 (N929, N921);
nand NAND3 (N930, N927, N2, N112);
nor NOR4 (N931, N914, N80, N718, N621);
and AND3 (N932, N924, N227, N625);
not NOT1 (N933, N931);
xor XOR2 (N934, N929, N445);
and AND2 (N935, N933, N749);
buf BUF1 (N936, N922);
xor XOR2 (N937, N930, N921);
not NOT1 (N938, N928);
xor XOR2 (N939, N936, N347);
nand NAND2 (N940, N935, N327);
xor XOR2 (N941, N939, N399);
xor XOR2 (N942, N940, N614);
nor NOR2 (N943, N938, N592);
not NOT1 (N944, N913);
nor NOR4 (N945, N944, N560, N2, N41);
buf BUF1 (N946, N923);
buf BUF1 (N947, N934);
nand NAND3 (N948, N945, N119, N936);
nand NAND3 (N949, N947, N336, N385);
buf BUF1 (N950, N943);
and AND3 (N951, N920, N37, N599);
nand NAND4 (N952, N950, N938, N203, N323);
nor NOR4 (N953, N948, N813, N56, N748);
nor NOR2 (N954, N932, N886);
xor XOR2 (N955, N941, N886);
not NOT1 (N956, N946);
and AND4 (N957, N903, N642, N458, N51);
xor XOR2 (N958, N955, N884);
or OR4 (N959, N956, N345, N21, N8);
or OR2 (N960, N958, N740);
not NOT1 (N961, N954);
nand NAND3 (N962, N953, N254, N922);
not NOT1 (N963, N937);
nand NAND4 (N964, N957, N774, N600, N362);
and AND4 (N965, N942, N143, N406, N775);
and AND3 (N966, N952, N965, N534);
nor NOR3 (N967, N828, N851, N771);
and AND3 (N968, N959, N476, N629);
nand NAND3 (N969, N966, N580, N780);
not NOT1 (N970, N951);
or OR4 (N971, N961, N751, N809, N43);
not NOT1 (N972, N949);
buf BUF1 (N973, N968);
not NOT1 (N974, N972);
not NOT1 (N975, N973);
or OR4 (N976, N970, N77, N159, N638);
nand NAND2 (N977, N974, N25);
nor NOR2 (N978, N962, N939);
not NOT1 (N979, N976);
buf BUF1 (N980, N963);
nand NAND3 (N981, N960, N490, N910);
nand NAND3 (N982, N964, N530, N976);
nor NOR4 (N983, N977, N667, N9, N464);
xor XOR2 (N984, N983, N185);
not NOT1 (N985, N984);
and AND2 (N986, N980, N788);
not NOT1 (N987, N971);
and AND2 (N988, N969, N944);
xor XOR2 (N989, N975, N442);
nand NAND4 (N990, N986, N495, N213, N141);
not NOT1 (N991, N982);
nand NAND2 (N992, N978, N114);
buf BUF1 (N993, N979);
and AND4 (N994, N967, N347, N28, N828);
or OR3 (N995, N987, N223, N911);
xor XOR2 (N996, N995, N348);
xor XOR2 (N997, N988, N19);
and AND4 (N998, N994, N500, N151, N685);
not NOT1 (N999, N989);
and AND4 (N1000, N998, N810, N74, N385);
and AND4 (N1001, N991, N482, N213, N407);
not NOT1 (N1002, N996);
or OR4 (N1003, N985, N144, N707, N636);
and AND3 (N1004, N997, N81, N288);
and AND4 (N1005, N993, N199, N637, N532);
nor NOR3 (N1006, N1003, N952, N985);
or OR2 (N1007, N990, N60);
and AND4 (N1008, N1007, N433, N7, N586);
not NOT1 (N1009, N1002);
and AND3 (N1010, N992, N682, N397);
nor NOR4 (N1011, N1006, N618, N553, N660);
xor XOR2 (N1012, N1000, N456);
not NOT1 (N1013, N1008);
xor XOR2 (N1014, N1010, N790);
xor XOR2 (N1015, N1005, N1000);
nor NOR4 (N1016, N999, N729, N537, N645);
buf BUF1 (N1017, N1004);
buf BUF1 (N1018, N1015);
buf BUF1 (N1019, N981);
buf BUF1 (N1020, N1001);
xor XOR2 (N1021, N1020, N823);
nand NAND4 (N1022, N1012, N63, N104, N198);
or OR4 (N1023, N1011, N435, N635, N963);
not NOT1 (N1024, N1021);
or OR4 (N1025, N1023, N568, N662, N38);
nor NOR2 (N1026, N1009, N767);
not NOT1 (N1027, N1017);
not NOT1 (N1028, N1014);
not NOT1 (N1029, N1025);
or OR4 (N1030, N1019, N21, N308, N970);
not NOT1 (N1031, N1022);
and AND3 (N1032, N1013, N283, N264);
nor NOR4 (N1033, N1027, N352, N512, N62);
nor NOR2 (N1034, N1031, N131);
nand NAND3 (N1035, N1016, N834, N751);
buf BUF1 (N1036, N1034);
nand NAND3 (N1037, N1036, N691, N859);
nor NOR4 (N1038, N1028, N343, N62, N67);
and AND3 (N1039, N1030, N72, N789);
nor NOR3 (N1040, N1024, N801, N817);
nor NOR3 (N1041, N1029, N174, N845);
nor NOR4 (N1042, N1026, N544, N999, N16);
not NOT1 (N1043, N1033);
not NOT1 (N1044, N1038);
and AND3 (N1045, N1032, N346, N309);
nand NAND2 (N1046, N1042, N454);
nor NOR4 (N1047, N1037, N520, N879, N777);
and AND3 (N1048, N1045, N698, N510);
buf BUF1 (N1049, N1048);
buf BUF1 (N1050, N1040);
nand NAND2 (N1051, N1046, N640);
not NOT1 (N1052, N1039);
and AND4 (N1053, N1044, N191, N291, N362);
not NOT1 (N1054, N1035);
xor XOR2 (N1055, N1054, N233);
nand NAND4 (N1056, N1047, N1009, N561, N1023);
nand NAND4 (N1057, N1018, N783, N362, N1026);
or OR4 (N1058, N1050, N526, N5, N828);
or OR3 (N1059, N1056, N673, N254);
not NOT1 (N1060, N1043);
nor NOR2 (N1061, N1059, N328);
buf BUF1 (N1062, N1051);
nand NAND4 (N1063, N1061, N332, N240, N833);
and AND3 (N1064, N1063, N144, N470);
not NOT1 (N1065, N1064);
nor NOR3 (N1066, N1055, N625, N247);
nand NAND4 (N1067, N1041, N379, N320, N573);
and AND3 (N1068, N1049, N403, N400);
not NOT1 (N1069, N1052);
nor NOR4 (N1070, N1062, N742, N716, N372);
not NOT1 (N1071, N1068);
nor NOR4 (N1072, N1071, N780, N420, N680);
and AND4 (N1073, N1058, N1052, N973, N192);
or OR4 (N1074, N1057, N375, N543, N730);
not NOT1 (N1075, N1073);
nand NAND3 (N1076, N1053, N25, N963);
and AND4 (N1077, N1067, N288, N538, N840);
nand NAND2 (N1078, N1075, N846);
nor NOR3 (N1079, N1066, N920, N774);
buf BUF1 (N1080, N1069);
nand NAND4 (N1081, N1079, N497, N145, N515);
nand NAND2 (N1082, N1074, N846);
nand NAND4 (N1083, N1082, N966, N467, N655);
nor NOR2 (N1084, N1080, N690);
and AND2 (N1085, N1060, N62);
or OR4 (N1086, N1078, N265, N908, N896);
nor NOR2 (N1087, N1070, N792);
not NOT1 (N1088, N1087);
xor XOR2 (N1089, N1084, N996);
nor NOR2 (N1090, N1076, N380);
xor XOR2 (N1091, N1088, N98);
and AND3 (N1092, N1065, N756, N77);
nand NAND3 (N1093, N1077, N799, N84);
nor NOR2 (N1094, N1072, N782);
nor NOR2 (N1095, N1085, N296);
nor NOR4 (N1096, N1094, N409, N522, N1058);
nor NOR4 (N1097, N1095, N169, N891, N24);
nand NAND2 (N1098, N1089, N904);
xor XOR2 (N1099, N1096, N463);
or OR4 (N1100, N1083, N308, N45, N705);
buf BUF1 (N1101, N1090);
buf BUF1 (N1102, N1097);
nor NOR4 (N1103, N1102, N1000, N1058, N404);
xor XOR2 (N1104, N1091, N671);
and AND3 (N1105, N1092, N151, N710);
xor XOR2 (N1106, N1098, N514);
not NOT1 (N1107, N1099);
buf BUF1 (N1108, N1107);
xor XOR2 (N1109, N1103, N689);
nand NAND3 (N1110, N1106, N547, N119);
nand NAND3 (N1111, N1086, N233, N887);
or OR4 (N1112, N1110, N399, N1010, N891);
buf BUF1 (N1113, N1105);
buf BUF1 (N1114, N1112);
and AND2 (N1115, N1109, N789);
or OR4 (N1116, N1104, N301, N477, N813);
or OR3 (N1117, N1100, N225, N871);
not NOT1 (N1118, N1117);
not NOT1 (N1119, N1093);
nand NAND3 (N1120, N1115, N522, N852);
not NOT1 (N1121, N1116);
buf BUF1 (N1122, N1101);
nor NOR2 (N1123, N1119, N344);
or OR4 (N1124, N1113, N473, N885, N349);
nand NAND2 (N1125, N1081, N470);
not NOT1 (N1126, N1122);
not NOT1 (N1127, N1111);
or OR2 (N1128, N1123, N1116);
nor NOR4 (N1129, N1126, N1016, N1119, N775);
or OR4 (N1130, N1114, N999, N859, N280);
and AND4 (N1131, N1124, N987, N879, N234);
or OR3 (N1132, N1129, N1043, N613);
and AND2 (N1133, N1128, N896);
nand NAND2 (N1134, N1133, N336);
and AND2 (N1135, N1134, N544);
xor XOR2 (N1136, N1135, N415);
and AND3 (N1137, N1130, N483, N1027);
or OR3 (N1138, N1131, N65, N954);
nand NAND4 (N1139, N1127, N439, N918, N672);
buf BUF1 (N1140, N1108);
or OR2 (N1141, N1136, N1077);
xor XOR2 (N1142, N1140, N211);
nand NAND2 (N1143, N1138, N598);
nand NAND2 (N1144, N1137, N814);
xor XOR2 (N1145, N1144, N97);
buf BUF1 (N1146, N1132);
buf BUF1 (N1147, N1139);
not NOT1 (N1148, N1118);
buf BUF1 (N1149, N1142);
not NOT1 (N1150, N1145);
buf BUF1 (N1151, N1120);
xor XOR2 (N1152, N1149, N769);
and AND2 (N1153, N1150, N999);
nor NOR2 (N1154, N1121, N423);
buf BUF1 (N1155, N1146);
and AND2 (N1156, N1148, N781);
not NOT1 (N1157, N1143);
nand NAND4 (N1158, N1155, N160, N367, N207);
and AND3 (N1159, N1156, N849, N630);
and AND4 (N1160, N1125, N197, N951, N998);
nor NOR4 (N1161, N1157, N579, N879, N822);
not NOT1 (N1162, N1141);
or OR3 (N1163, N1162, N223, N28);
buf BUF1 (N1164, N1152);
nor NOR4 (N1165, N1159, N1045, N637, N1012);
xor XOR2 (N1166, N1160, N820);
not NOT1 (N1167, N1163);
nand NAND4 (N1168, N1153, N981, N275, N799);
and AND4 (N1169, N1154, N5, N1112, N725);
nand NAND3 (N1170, N1166, N904, N909);
or OR3 (N1171, N1170, N322, N161);
nor NOR2 (N1172, N1158, N472);
not NOT1 (N1173, N1164);
buf BUF1 (N1174, N1151);
buf BUF1 (N1175, N1172);
not NOT1 (N1176, N1175);
buf BUF1 (N1177, N1169);
nor NOR2 (N1178, N1167, N1019);
or OR4 (N1179, N1165, N202, N725, N295);
not NOT1 (N1180, N1161);
buf BUF1 (N1181, N1179);
or OR3 (N1182, N1181, N577, N19);
buf BUF1 (N1183, N1174);
or OR2 (N1184, N1147, N187);
nor NOR4 (N1185, N1182, N1003, N390, N488);
not NOT1 (N1186, N1180);
or OR2 (N1187, N1178, N313);
nand NAND2 (N1188, N1187, N241);
nor NOR3 (N1189, N1176, N345, N938);
xor XOR2 (N1190, N1185, N916);
nand NAND2 (N1191, N1168, N650);
buf BUF1 (N1192, N1188);
buf BUF1 (N1193, N1173);
nand NAND4 (N1194, N1184, N568, N798, N557);
xor XOR2 (N1195, N1183, N282);
and AND2 (N1196, N1191, N367);
nand NAND2 (N1197, N1190, N121);
nand NAND2 (N1198, N1177, N628);
xor XOR2 (N1199, N1193, N995);
buf BUF1 (N1200, N1198);
xor XOR2 (N1201, N1189, N1063);
xor XOR2 (N1202, N1194, N1078);
buf BUF1 (N1203, N1197);
xor XOR2 (N1204, N1200, N169);
xor XOR2 (N1205, N1192, N1182);
nor NOR2 (N1206, N1204, N185);
nor NOR3 (N1207, N1205, N515, N1105);
buf BUF1 (N1208, N1201);
nor NOR2 (N1209, N1208, N220);
not NOT1 (N1210, N1186);
not NOT1 (N1211, N1207);
nand NAND4 (N1212, N1202, N503, N1028, N322);
buf BUF1 (N1213, N1210);
not NOT1 (N1214, N1211);
not NOT1 (N1215, N1206);
and AND3 (N1216, N1195, N579, N97);
nand NAND3 (N1217, N1209, N1074, N1051);
not NOT1 (N1218, N1215);
buf BUF1 (N1219, N1199);
not NOT1 (N1220, N1213);
nor NOR2 (N1221, N1171, N352);
and AND3 (N1222, N1203, N625, N133);
and AND3 (N1223, N1222, N11, N385);
and AND4 (N1224, N1212, N229, N21, N401);
and AND3 (N1225, N1218, N77, N681);
and AND2 (N1226, N1225, N626);
nor NOR2 (N1227, N1214, N1127);
and AND2 (N1228, N1217, N831);
not NOT1 (N1229, N1221);
nor NOR2 (N1230, N1220, N1178);
buf BUF1 (N1231, N1230);
and AND3 (N1232, N1228, N1193, N930);
nand NAND3 (N1233, N1196, N1122, N568);
or OR2 (N1234, N1227, N164);
and AND4 (N1235, N1226, N326, N759, N104);
xor XOR2 (N1236, N1233, N106);
and AND4 (N1237, N1234, N711, N10, N497);
or OR2 (N1238, N1216, N860);
nand NAND3 (N1239, N1224, N225, N858);
buf BUF1 (N1240, N1229);
not NOT1 (N1241, N1235);
nand NAND2 (N1242, N1236, N47);
not NOT1 (N1243, N1223);
nand NAND4 (N1244, N1231, N699, N452, N555);
nand NAND4 (N1245, N1243, N614, N197, N1098);
xor XOR2 (N1246, N1237, N687);
not NOT1 (N1247, N1241);
or OR3 (N1248, N1245, N826, N919);
nor NOR2 (N1249, N1242, N1032);
nor NOR3 (N1250, N1248, N423, N488);
and AND2 (N1251, N1250, N883);
nand NAND3 (N1252, N1240, N1068, N319);
xor XOR2 (N1253, N1251, N909);
and AND2 (N1254, N1232, N947);
not NOT1 (N1255, N1247);
or OR4 (N1256, N1246, N931, N878, N1072);
not NOT1 (N1257, N1256);
not NOT1 (N1258, N1252);
nor NOR3 (N1259, N1258, N1054, N23);
nand NAND4 (N1260, N1244, N1181, N815, N116);
nand NAND3 (N1261, N1253, N629, N306);
buf BUF1 (N1262, N1261);
or OR4 (N1263, N1257, N647, N180, N826);
and AND2 (N1264, N1262, N873);
buf BUF1 (N1265, N1239);
xor XOR2 (N1266, N1254, N587);
xor XOR2 (N1267, N1238, N786);
and AND2 (N1268, N1267, N1027);
or OR2 (N1269, N1264, N783);
nor NOR4 (N1270, N1255, N1072, N149, N971);
nand NAND2 (N1271, N1260, N988);
xor XOR2 (N1272, N1271, N433);
nor NOR4 (N1273, N1272, N308, N445, N1206);
xor XOR2 (N1274, N1266, N291);
or OR4 (N1275, N1219, N500, N1128, N446);
and AND3 (N1276, N1274, N442, N332);
nor NOR2 (N1277, N1273, N1178);
buf BUF1 (N1278, N1249);
and AND3 (N1279, N1276, N937, N77);
and AND4 (N1280, N1269, N653, N288, N506);
and AND4 (N1281, N1278, N487, N763, N631);
nand NAND3 (N1282, N1268, N751, N1084);
nand NAND4 (N1283, N1265, N567, N454, N209);
and AND2 (N1284, N1277, N514);
and AND4 (N1285, N1284, N1191, N538, N1281);
nor NOR2 (N1286, N28, N813);
xor XOR2 (N1287, N1282, N714);
or OR4 (N1288, N1275, N488, N436, N101);
nand NAND3 (N1289, N1283, N827, N125);
nand NAND4 (N1290, N1287, N848, N1256, N454);
nor NOR3 (N1291, N1290, N1135, N372);
or OR2 (N1292, N1263, N526);
and AND2 (N1293, N1279, N52);
or OR2 (N1294, N1286, N69);
not NOT1 (N1295, N1259);
nand NAND4 (N1296, N1293, N545, N1056, N145);
xor XOR2 (N1297, N1289, N110);
and AND3 (N1298, N1292, N720, N779);
buf BUF1 (N1299, N1296);
nand NAND3 (N1300, N1298, N266, N1226);
nor NOR3 (N1301, N1294, N1026, N325);
buf BUF1 (N1302, N1280);
buf BUF1 (N1303, N1299);
nor NOR3 (N1304, N1270, N1239, N1295);
and AND3 (N1305, N193, N26, N748);
not NOT1 (N1306, N1302);
and AND2 (N1307, N1300, N364);
buf BUF1 (N1308, N1305);
or OR2 (N1309, N1301, N1244);
or OR2 (N1310, N1307, N1003);
and AND2 (N1311, N1308, N832);
or OR4 (N1312, N1310, N1031, N853, N6);
nand NAND3 (N1313, N1306, N740, N1149);
buf BUF1 (N1314, N1309);
and AND2 (N1315, N1314, N974);
nand NAND3 (N1316, N1285, N553, N480);
buf BUF1 (N1317, N1311);
xor XOR2 (N1318, N1313, N627);
or OR2 (N1319, N1303, N821);
and AND2 (N1320, N1291, N984);
buf BUF1 (N1321, N1304);
not NOT1 (N1322, N1320);
not NOT1 (N1323, N1321);
or OR4 (N1324, N1318, N666, N195, N162);
xor XOR2 (N1325, N1324, N152);
xor XOR2 (N1326, N1322, N794);
xor XOR2 (N1327, N1323, N1140);
buf BUF1 (N1328, N1316);
not NOT1 (N1329, N1317);
nor NOR3 (N1330, N1326, N1018, N303);
buf BUF1 (N1331, N1327);
and AND2 (N1332, N1325, N876);
nand NAND3 (N1333, N1297, N534, N358);
xor XOR2 (N1334, N1333, N1291);
buf BUF1 (N1335, N1288);
buf BUF1 (N1336, N1328);
buf BUF1 (N1337, N1315);
nor NOR4 (N1338, N1334, N1056, N545, N551);
xor XOR2 (N1339, N1319, N410);
not NOT1 (N1340, N1339);
buf BUF1 (N1341, N1332);
xor XOR2 (N1342, N1329, N918);
xor XOR2 (N1343, N1340, N679);
xor XOR2 (N1344, N1342, N721);
or OR4 (N1345, N1337, N1023, N479, N1074);
nor NOR2 (N1346, N1338, N27);
xor XOR2 (N1347, N1345, N363);
buf BUF1 (N1348, N1346);
not NOT1 (N1349, N1348);
nand NAND4 (N1350, N1330, N644, N492, N422);
or OR2 (N1351, N1344, N974);
xor XOR2 (N1352, N1335, N499);
buf BUF1 (N1353, N1351);
nor NOR2 (N1354, N1341, N113);
and AND4 (N1355, N1312, N921, N108, N573);
nand NAND3 (N1356, N1349, N896, N531);
nor NOR2 (N1357, N1352, N1132);
and AND2 (N1358, N1353, N781);
xor XOR2 (N1359, N1336, N692);
or OR2 (N1360, N1347, N180);
and AND3 (N1361, N1359, N957, N5);
not NOT1 (N1362, N1357);
and AND4 (N1363, N1361, N1012, N687, N1345);
xor XOR2 (N1364, N1355, N1169);
or OR4 (N1365, N1354, N170, N1089, N616);
nand NAND2 (N1366, N1362, N1124);
nand NAND4 (N1367, N1360, N24, N1173, N21);
not NOT1 (N1368, N1367);
buf BUF1 (N1369, N1366);
not NOT1 (N1370, N1363);
xor XOR2 (N1371, N1364, N276);
xor XOR2 (N1372, N1369, N1154);
buf BUF1 (N1373, N1371);
nor NOR4 (N1374, N1358, N1001, N989, N1065);
and AND2 (N1375, N1365, N1145);
and AND4 (N1376, N1350, N1283, N697, N332);
xor XOR2 (N1377, N1374, N446);
or OR4 (N1378, N1356, N572, N93, N1188);
buf BUF1 (N1379, N1368);
and AND3 (N1380, N1331, N788, N1245);
or OR2 (N1381, N1376, N602);
buf BUF1 (N1382, N1377);
not NOT1 (N1383, N1370);
and AND2 (N1384, N1382, N702);
xor XOR2 (N1385, N1343, N145);
xor XOR2 (N1386, N1383, N318);
buf BUF1 (N1387, N1379);
and AND3 (N1388, N1375, N1099, N1033);
xor XOR2 (N1389, N1385, N1043);
xor XOR2 (N1390, N1378, N1275);
buf BUF1 (N1391, N1388);
xor XOR2 (N1392, N1384, N872);
nor NOR4 (N1393, N1387, N537, N1010, N500);
not NOT1 (N1394, N1390);
or OR3 (N1395, N1394, N1196, N1240);
buf BUF1 (N1396, N1380);
buf BUF1 (N1397, N1392);
nor NOR2 (N1398, N1389, N922);
and AND3 (N1399, N1393, N200, N1122);
and AND2 (N1400, N1398, N523);
and AND3 (N1401, N1396, N187, N1289);
not NOT1 (N1402, N1397);
nand NAND4 (N1403, N1372, N768, N480, N872);
xor XOR2 (N1404, N1400, N308);
buf BUF1 (N1405, N1391);
xor XOR2 (N1406, N1403, N283);
or OR2 (N1407, N1405, N309);
nor NOR3 (N1408, N1373, N1008, N199);
buf BUF1 (N1409, N1402);
nand NAND2 (N1410, N1399, N832);
xor XOR2 (N1411, N1381, N80);
nor NOR2 (N1412, N1386, N355);
nor NOR2 (N1413, N1401, N79);
nand NAND4 (N1414, N1413, N910, N529, N79);
and AND2 (N1415, N1410, N960);
not NOT1 (N1416, N1407);
xor XOR2 (N1417, N1411, N1203);
nor NOR3 (N1418, N1412, N1099, N232);
not NOT1 (N1419, N1404);
and AND2 (N1420, N1395, N698);
nor NOR3 (N1421, N1415, N1405, N871);
and AND3 (N1422, N1418, N397, N471);
nor NOR4 (N1423, N1421, N389, N2, N1192);
buf BUF1 (N1424, N1417);
or OR4 (N1425, N1423, N770, N1335, N1281);
or OR4 (N1426, N1424, N266, N1105, N334);
or OR4 (N1427, N1419, N1164, N143, N597);
nor NOR2 (N1428, N1409, N1140);
and AND4 (N1429, N1420, N1423, N170, N847);
not NOT1 (N1430, N1428);
nor NOR2 (N1431, N1414, N952);
nand NAND2 (N1432, N1408, N730);
nor NOR2 (N1433, N1416, N123);
nand NAND2 (N1434, N1430, N349);
buf BUF1 (N1435, N1427);
xor XOR2 (N1436, N1431, N797);
and AND2 (N1437, N1425, N1381);
nor NOR4 (N1438, N1422, N576, N426, N1406);
xor XOR2 (N1439, N609, N1079);
nand NAND4 (N1440, N1429, N837, N290, N1275);
and AND3 (N1441, N1439, N204, N472);
and AND2 (N1442, N1426, N974);
nand NAND3 (N1443, N1442, N1127, N552);
xor XOR2 (N1444, N1441, N1279);
buf BUF1 (N1445, N1443);
and AND2 (N1446, N1440, N948);
and AND3 (N1447, N1436, N1274, N65);
or OR2 (N1448, N1444, N1342);
buf BUF1 (N1449, N1446);
not NOT1 (N1450, N1433);
and AND3 (N1451, N1432, N843, N889);
and AND2 (N1452, N1435, N16);
xor XOR2 (N1453, N1437, N1341);
and AND3 (N1454, N1448, N1389, N668);
buf BUF1 (N1455, N1438);
and AND3 (N1456, N1450, N140, N1131);
nand NAND3 (N1457, N1445, N1338, N1240);
buf BUF1 (N1458, N1456);
buf BUF1 (N1459, N1454);
not NOT1 (N1460, N1459);
and AND4 (N1461, N1434, N1256, N1209, N398);
nand NAND4 (N1462, N1458, N384, N383, N1295);
or OR4 (N1463, N1455, N1272, N1203, N970);
nor NOR4 (N1464, N1460, N816, N154, N942);
or OR3 (N1465, N1447, N476, N1165);
nor NOR4 (N1466, N1464, N1002, N658, N1464);
nand NAND2 (N1467, N1461, N976);
and AND3 (N1468, N1466, N1221, N1093);
nor NOR4 (N1469, N1468, N538, N678, N423);
not NOT1 (N1470, N1462);
or OR4 (N1471, N1451, N211, N880, N1079);
and AND3 (N1472, N1470, N200, N615);
buf BUF1 (N1473, N1452);
or OR2 (N1474, N1469, N1374);
xor XOR2 (N1475, N1449, N272);
buf BUF1 (N1476, N1471);
xor XOR2 (N1477, N1476, N16);
not NOT1 (N1478, N1473);
not NOT1 (N1479, N1463);
xor XOR2 (N1480, N1479, N899);
xor XOR2 (N1481, N1475, N127);
or OR2 (N1482, N1472, N469);
or OR4 (N1483, N1453, N701, N1233, N141);
nor NOR3 (N1484, N1482, N594, N1424);
not NOT1 (N1485, N1457);
buf BUF1 (N1486, N1483);
not NOT1 (N1487, N1474);
buf BUF1 (N1488, N1484);
buf BUF1 (N1489, N1487);
and AND2 (N1490, N1485, N1178);
nor NOR3 (N1491, N1465, N606, N877);
not NOT1 (N1492, N1478);
not NOT1 (N1493, N1490);
or OR4 (N1494, N1486, N159, N586, N274);
and AND3 (N1495, N1480, N1321, N1414);
buf BUF1 (N1496, N1491);
not NOT1 (N1497, N1493);
not NOT1 (N1498, N1489);
not NOT1 (N1499, N1496);
xor XOR2 (N1500, N1497, N121);
xor XOR2 (N1501, N1488, N703);
buf BUF1 (N1502, N1494);
buf BUF1 (N1503, N1481);
or OR4 (N1504, N1477, N952, N965, N683);
buf BUF1 (N1505, N1492);
xor XOR2 (N1506, N1503, N1101);
and AND3 (N1507, N1467, N43, N1075);
xor XOR2 (N1508, N1495, N603);
buf BUF1 (N1509, N1501);
nor NOR4 (N1510, N1499, N1414, N1428, N411);
not NOT1 (N1511, N1498);
and AND2 (N1512, N1505, N823);
buf BUF1 (N1513, N1506);
not NOT1 (N1514, N1508);
nor NOR4 (N1515, N1500, N835, N1271, N947);
and AND2 (N1516, N1509, N403);
not NOT1 (N1517, N1514);
or OR4 (N1518, N1513, N252, N356, N33);
and AND2 (N1519, N1512, N850);
nand NAND4 (N1520, N1502, N181, N726, N1507);
and AND4 (N1521, N742, N280, N493, N787);
buf BUF1 (N1522, N1520);
not NOT1 (N1523, N1518);
or OR4 (N1524, N1519, N938, N229, N1159);
or OR2 (N1525, N1504, N1403);
nand NAND2 (N1526, N1517, N663);
buf BUF1 (N1527, N1521);
xor XOR2 (N1528, N1523, N946);
nand NAND2 (N1529, N1515, N17);
not NOT1 (N1530, N1524);
or OR3 (N1531, N1528, N818, N139);
nor NOR3 (N1532, N1511, N1432, N540);
nor NOR3 (N1533, N1532, N1438, N641);
xor XOR2 (N1534, N1531, N1078);
nor NOR3 (N1535, N1529, N1162, N442);
nand NAND4 (N1536, N1535, N1004, N56, N729);
buf BUF1 (N1537, N1536);
buf BUF1 (N1538, N1522);
nor NOR3 (N1539, N1525, N255, N610);
not NOT1 (N1540, N1538);
or OR2 (N1541, N1510, N943);
or OR4 (N1542, N1539, N305, N776, N500);
and AND2 (N1543, N1541, N801);
buf BUF1 (N1544, N1543);
nor NOR3 (N1545, N1537, N1522, N520);
or OR3 (N1546, N1533, N806, N471);
not NOT1 (N1547, N1545);
buf BUF1 (N1548, N1527);
buf BUF1 (N1549, N1526);
nor NOR3 (N1550, N1549, N661, N226);
xor XOR2 (N1551, N1530, N151);
and AND3 (N1552, N1548, N484, N632);
nand NAND3 (N1553, N1546, N768, N866);
not NOT1 (N1554, N1552);
and AND2 (N1555, N1516, N1440);
buf BUF1 (N1556, N1551);
not NOT1 (N1557, N1555);
or OR4 (N1558, N1556, N1042, N774, N987);
nor NOR2 (N1559, N1534, N66);
buf BUF1 (N1560, N1559);
xor XOR2 (N1561, N1547, N902);
buf BUF1 (N1562, N1542);
xor XOR2 (N1563, N1544, N1329);
not NOT1 (N1564, N1554);
or OR2 (N1565, N1553, N33);
xor XOR2 (N1566, N1557, N287);
nand NAND2 (N1567, N1540, N417);
nor NOR4 (N1568, N1558, N1246, N141, N1095);
and AND2 (N1569, N1560, N209);
nand NAND3 (N1570, N1567, N240, N826);
and AND4 (N1571, N1550, N736, N27, N1343);
and AND2 (N1572, N1566, N693);
or OR3 (N1573, N1568, N728, N1124);
xor XOR2 (N1574, N1561, N1413);
nand NAND4 (N1575, N1564, N960, N393, N586);
not NOT1 (N1576, N1571);
or OR2 (N1577, N1565, N86);
nor NOR2 (N1578, N1574, N558);
and AND3 (N1579, N1577, N1518, N253);
not NOT1 (N1580, N1578);
xor XOR2 (N1581, N1562, N27);
nand NAND2 (N1582, N1573, N532);
xor XOR2 (N1583, N1580, N22);
and AND3 (N1584, N1572, N829, N1347);
buf BUF1 (N1585, N1570);
and AND4 (N1586, N1576, N758, N1078, N1234);
buf BUF1 (N1587, N1585);
nor NOR3 (N1588, N1584, N789, N3);
buf BUF1 (N1589, N1582);
nand NAND2 (N1590, N1569, N151);
nand NAND3 (N1591, N1579, N286, N321);
or OR3 (N1592, N1589, N938, N1494);
not NOT1 (N1593, N1588);
nand NAND2 (N1594, N1586, N33);
nor NOR3 (N1595, N1594, N1000, N630);
and AND4 (N1596, N1575, N1278, N391, N650);
not NOT1 (N1597, N1581);
not NOT1 (N1598, N1590);
xor XOR2 (N1599, N1591, N611);
buf BUF1 (N1600, N1592);
nor NOR2 (N1601, N1596, N1530);
buf BUF1 (N1602, N1598);
buf BUF1 (N1603, N1597);
and AND2 (N1604, N1603, N611);
or OR3 (N1605, N1602, N1258, N681);
nor NOR3 (N1606, N1587, N458, N704);
and AND2 (N1607, N1600, N246);
nor NOR2 (N1608, N1601, N1069);
nor NOR4 (N1609, N1604, N1016, N1606, N1191);
or OR4 (N1610, N412, N297, N477, N1226);
and AND2 (N1611, N1595, N1428);
not NOT1 (N1612, N1583);
buf BUF1 (N1613, N1563);
and AND4 (N1614, N1608, N1560, N1327, N1063);
nand NAND3 (N1615, N1614, N155, N1547);
and AND2 (N1616, N1607, N1060);
xor XOR2 (N1617, N1616, N969);
xor XOR2 (N1618, N1617, N667);
or OR3 (N1619, N1593, N1524, N1000);
or OR2 (N1620, N1610, N1334);
nand NAND2 (N1621, N1613, N1385);
nor NOR3 (N1622, N1609, N252, N1053);
buf BUF1 (N1623, N1619);
not NOT1 (N1624, N1612);
not NOT1 (N1625, N1611);
nor NOR2 (N1626, N1599, N1030);
buf BUF1 (N1627, N1620);
nor NOR3 (N1628, N1626, N649, N606);
and AND2 (N1629, N1605, N597);
xor XOR2 (N1630, N1629, N350);
or OR2 (N1631, N1630, N1539);
nor NOR4 (N1632, N1625, N1252, N306, N550);
xor XOR2 (N1633, N1631, N741);
xor XOR2 (N1634, N1621, N550);
nor NOR2 (N1635, N1618, N498);
nand NAND2 (N1636, N1624, N511);
buf BUF1 (N1637, N1636);
not NOT1 (N1638, N1633);
xor XOR2 (N1639, N1615, N1613);
nand NAND4 (N1640, N1638, N220, N311, N1269);
and AND3 (N1641, N1627, N1027, N485);
nor NOR4 (N1642, N1622, N434, N268, N286);
buf BUF1 (N1643, N1639);
or OR2 (N1644, N1628, N255);
or OR3 (N1645, N1623, N1529, N1182);
buf BUF1 (N1646, N1632);
buf BUF1 (N1647, N1645);
or OR3 (N1648, N1647, N1105, N264);
not NOT1 (N1649, N1648);
and AND2 (N1650, N1642, N1083);
or OR3 (N1651, N1637, N1618, N82);
not NOT1 (N1652, N1635);
and AND3 (N1653, N1640, N592, N390);
nor NOR3 (N1654, N1650, N120, N1326);
buf BUF1 (N1655, N1643);
nand NAND2 (N1656, N1651, N1196);
buf BUF1 (N1657, N1649);
nand NAND4 (N1658, N1634, N678, N252, N1190);
and AND3 (N1659, N1658, N722, N1603);
nand NAND2 (N1660, N1652, N1386);
not NOT1 (N1661, N1657);
buf BUF1 (N1662, N1653);
nor NOR4 (N1663, N1655, N1479, N36, N773);
buf BUF1 (N1664, N1660);
buf BUF1 (N1665, N1644);
not NOT1 (N1666, N1663);
or OR3 (N1667, N1661, N876, N1232);
nor NOR3 (N1668, N1666, N1322, N723);
or OR4 (N1669, N1641, N330, N815, N1055);
nor NOR2 (N1670, N1664, N1006);
nor NOR3 (N1671, N1654, N668, N897);
buf BUF1 (N1672, N1665);
nor NOR4 (N1673, N1646, N1309, N1041, N633);
buf BUF1 (N1674, N1672);
nor NOR4 (N1675, N1670, N1619, N356, N1571);
xor XOR2 (N1676, N1675, N886);
nand NAND3 (N1677, N1674, N635, N1507);
or OR4 (N1678, N1669, N138, N756, N1083);
or OR2 (N1679, N1668, N935);
and AND3 (N1680, N1677, N1642, N1385);
nor NOR3 (N1681, N1676, N100, N1589);
nand NAND4 (N1682, N1681, N1527, N913, N823);
nand NAND3 (N1683, N1667, N1256, N1477);
xor XOR2 (N1684, N1682, N1212);
not NOT1 (N1685, N1680);
nor NOR2 (N1686, N1685, N1608);
not NOT1 (N1687, N1662);
nor NOR2 (N1688, N1656, N1058);
not NOT1 (N1689, N1659);
nor NOR2 (N1690, N1688, N713);
nor NOR3 (N1691, N1679, N1071, N1618);
or OR2 (N1692, N1671, N140);
and AND4 (N1693, N1687, N175, N1224, N1550);
buf BUF1 (N1694, N1691);
nand NAND3 (N1695, N1690, N552, N674);
or OR4 (N1696, N1689, N772, N282, N62);
or OR3 (N1697, N1692, N1403, N904);
xor XOR2 (N1698, N1696, N650);
xor XOR2 (N1699, N1683, N1285);
xor XOR2 (N1700, N1673, N779);
nand NAND4 (N1701, N1697, N1300, N1241, N1250);
not NOT1 (N1702, N1701);
buf BUF1 (N1703, N1695);
nor NOR2 (N1704, N1702, N1230);
nor NOR2 (N1705, N1684, N208);
nor NOR4 (N1706, N1694, N1010, N1624, N362);
buf BUF1 (N1707, N1698);
xor XOR2 (N1708, N1678, N948);
buf BUF1 (N1709, N1686);
nand NAND2 (N1710, N1704, N1694);
or OR4 (N1711, N1708, N1039, N112, N1120);
or OR4 (N1712, N1703, N383, N523, N1576);
or OR4 (N1713, N1710, N501, N1278, N572);
nor NOR2 (N1714, N1711, N810);
xor XOR2 (N1715, N1712, N1261);
not NOT1 (N1716, N1706);
nand NAND2 (N1717, N1705, N710);
and AND4 (N1718, N1709, N1457, N1656, N417);
xor XOR2 (N1719, N1700, N754);
nor NOR3 (N1720, N1719, N1489, N1298);
buf BUF1 (N1721, N1717);
and AND2 (N1722, N1721, N1603);
and AND4 (N1723, N1718, N62, N985, N1163);
xor XOR2 (N1724, N1707, N1365);
and AND2 (N1725, N1720, N196);
nand NAND4 (N1726, N1715, N1214, N356, N520);
or OR2 (N1727, N1714, N7);
buf BUF1 (N1728, N1699);
xor XOR2 (N1729, N1722, N1611);
nor NOR3 (N1730, N1723, N767, N1573);
and AND3 (N1731, N1730, N421, N1518);
and AND4 (N1732, N1726, N150, N1579, N586);
or OR3 (N1733, N1725, N55, N1410);
or OR4 (N1734, N1729, N739, N903, N679);
not NOT1 (N1735, N1731);
not NOT1 (N1736, N1724);
and AND3 (N1737, N1716, N1439, N976);
buf BUF1 (N1738, N1727);
and AND3 (N1739, N1734, N754, N1593);
buf BUF1 (N1740, N1713);
xor XOR2 (N1741, N1736, N5);
and AND3 (N1742, N1741, N1031, N1388);
or OR3 (N1743, N1728, N1472, N294);
not NOT1 (N1744, N1743);
not NOT1 (N1745, N1735);
and AND3 (N1746, N1737, N1000, N1456);
nand NAND3 (N1747, N1693, N1518, N657);
nand NAND4 (N1748, N1733, N839, N61, N775);
and AND3 (N1749, N1739, N777, N390);
and AND3 (N1750, N1738, N994, N933);
buf BUF1 (N1751, N1732);
nor NOR4 (N1752, N1750, N88, N486, N379);
nor NOR3 (N1753, N1752, N1450, N1188);
or OR2 (N1754, N1744, N1559);
nand NAND3 (N1755, N1748, N15, N1370);
and AND4 (N1756, N1754, N399, N1591, N769);
xor XOR2 (N1757, N1742, N522);
xor XOR2 (N1758, N1740, N1526);
buf BUF1 (N1759, N1749);
nor NOR3 (N1760, N1753, N766, N1188);
buf BUF1 (N1761, N1747);
nor NOR4 (N1762, N1751, N1570, N1040, N1252);
buf BUF1 (N1763, N1755);
not NOT1 (N1764, N1759);
not NOT1 (N1765, N1763);
nor NOR2 (N1766, N1758, N621);
xor XOR2 (N1767, N1746, N490);
or OR2 (N1768, N1757, N838);
or OR3 (N1769, N1766, N1431, N789);
and AND2 (N1770, N1764, N739);
nor NOR2 (N1771, N1762, N1439);
nor NOR2 (N1772, N1760, N267);
nand NAND4 (N1773, N1768, N436, N724, N1516);
or OR3 (N1774, N1767, N650, N522);
not NOT1 (N1775, N1771);
not NOT1 (N1776, N1769);
xor XOR2 (N1777, N1770, N1659);
buf BUF1 (N1778, N1774);
not NOT1 (N1779, N1772);
and AND2 (N1780, N1756, N1136);
buf BUF1 (N1781, N1765);
nand NAND3 (N1782, N1778, N687, N315);
or OR3 (N1783, N1780, N915, N823);
or OR4 (N1784, N1773, N627, N148, N849);
nor NOR3 (N1785, N1783, N247, N1014);
and AND4 (N1786, N1776, N1328, N537, N1764);
nor NOR4 (N1787, N1781, N1081, N798, N83);
nand NAND3 (N1788, N1784, N1234, N1261);
or OR4 (N1789, N1745, N1231, N672, N743);
not NOT1 (N1790, N1779);
buf BUF1 (N1791, N1777);
nand NAND2 (N1792, N1775, N1597);
buf BUF1 (N1793, N1788);
and AND2 (N1794, N1789, N1008);
nor NOR2 (N1795, N1787, N83);
or OR3 (N1796, N1785, N800, N674);
and AND4 (N1797, N1795, N72, N150, N73);
nand NAND3 (N1798, N1793, N308, N367);
nand NAND4 (N1799, N1792, N1090, N1331, N682);
or OR3 (N1800, N1794, N1392, N139);
and AND3 (N1801, N1786, N1576, N1204);
or OR4 (N1802, N1790, N493, N1233, N1294);
and AND4 (N1803, N1791, N1098, N21, N587);
not NOT1 (N1804, N1782);
nor NOR2 (N1805, N1803, N271);
xor XOR2 (N1806, N1804, N615);
nor NOR3 (N1807, N1761, N95, N445);
nor NOR2 (N1808, N1806, N858);
not NOT1 (N1809, N1801);
buf BUF1 (N1810, N1805);
not NOT1 (N1811, N1802);
and AND4 (N1812, N1809, N940, N30, N201);
buf BUF1 (N1813, N1812);
and AND3 (N1814, N1808, N1436, N730);
nor NOR4 (N1815, N1798, N1137, N1665, N260);
nor NOR3 (N1816, N1811, N1158, N1427);
nand NAND3 (N1817, N1799, N577, N224);
or OR4 (N1818, N1814, N1145, N557, N221);
xor XOR2 (N1819, N1800, N1591);
xor XOR2 (N1820, N1810, N1061);
nor NOR2 (N1821, N1818, N302);
buf BUF1 (N1822, N1797);
xor XOR2 (N1823, N1821, N1597);
nor NOR4 (N1824, N1820, N291, N670, N734);
not NOT1 (N1825, N1817);
nor NOR3 (N1826, N1824, N435, N1081);
and AND4 (N1827, N1796, N157, N1799, N758);
and AND3 (N1828, N1822, N236, N41);
nand NAND4 (N1829, N1823, N1425, N800, N1362);
buf BUF1 (N1830, N1819);
not NOT1 (N1831, N1828);
buf BUF1 (N1832, N1827);
xor XOR2 (N1833, N1815, N312);
and AND4 (N1834, N1826, N855, N292, N812);
and AND3 (N1835, N1813, N300, N1780);
xor XOR2 (N1836, N1829, N996);
buf BUF1 (N1837, N1831);
nand NAND3 (N1838, N1830, N219, N276);
not NOT1 (N1839, N1832);
nor NOR3 (N1840, N1839, N1818, N525);
not NOT1 (N1841, N1840);
xor XOR2 (N1842, N1838, N423);
buf BUF1 (N1843, N1842);
or OR4 (N1844, N1833, N262, N76, N1811);
nand NAND3 (N1845, N1834, N59, N625);
not NOT1 (N1846, N1816);
xor XOR2 (N1847, N1843, N634);
and AND4 (N1848, N1846, N386, N716, N1713);
nor NOR2 (N1849, N1837, N700);
nand NAND3 (N1850, N1847, N179, N514);
nand NAND2 (N1851, N1845, N750);
and AND4 (N1852, N1835, N10, N1104, N1155);
xor XOR2 (N1853, N1850, N1135);
buf BUF1 (N1854, N1807);
xor XOR2 (N1855, N1848, N151);
xor XOR2 (N1856, N1852, N245);
nand NAND2 (N1857, N1836, N949);
and AND2 (N1858, N1841, N1050);
buf BUF1 (N1859, N1849);
or OR3 (N1860, N1855, N1566, N1664);
buf BUF1 (N1861, N1825);
xor XOR2 (N1862, N1844, N1654);
xor XOR2 (N1863, N1857, N1147);
or OR3 (N1864, N1853, N1590, N1763);
buf BUF1 (N1865, N1862);
or OR3 (N1866, N1858, N499, N1196);
nor NOR3 (N1867, N1863, N1766, N158);
and AND4 (N1868, N1864, N397, N75, N1855);
nand NAND2 (N1869, N1865, N1362);
nand NAND4 (N1870, N1867, N838, N105, N626);
and AND2 (N1871, N1869, N416);
not NOT1 (N1872, N1861);
nor NOR3 (N1873, N1868, N650, N869);
nor NOR2 (N1874, N1859, N566);
nand NAND4 (N1875, N1870, N500, N235, N633);
not NOT1 (N1876, N1866);
nand NAND4 (N1877, N1871, N419, N141, N1329);
nand NAND2 (N1878, N1873, N1010);
and AND3 (N1879, N1878, N1523, N1128);
buf BUF1 (N1880, N1876);
nand NAND4 (N1881, N1872, N993, N1400, N1517);
or OR2 (N1882, N1860, N544);
xor XOR2 (N1883, N1880, N515);
and AND4 (N1884, N1851, N1366, N1142, N989);
and AND3 (N1885, N1879, N944, N1377);
not NOT1 (N1886, N1875);
nand NAND3 (N1887, N1882, N254, N1590);
and AND3 (N1888, N1854, N22, N1667);
not NOT1 (N1889, N1886);
nor NOR3 (N1890, N1881, N1391, N1789);
xor XOR2 (N1891, N1887, N380);
nor NOR4 (N1892, N1877, N389, N1551, N1421);
or OR4 (N1893, N1884, N1643, N1144, N1142);
nand NAND4 (N1894, N1890, N1827, N1278, N580);
not NOT1 (N1895, N1856);
xor XOR2 (N1896, N1893, N429);
and AND2 (N1897, N1892, N548);
buf BUF1 (N1898, N1896);
nand NAND4 (N1899, N1889, N27, N807, N851);
xor XOR2 (N1900, N1899, N611);
or OR2 (N1901, N1900, N1510);
buf BUF1 (N1902, N1891);
nor NOR2 (N1903, N1883, N1857);
nand NAND4 (N1904, N1897, N120, N568, N1237);
and AND2 (N1905, N1898, N1779);
not NOT1 (N1906, N1874);
or OR2 (N1907, N1894, N1378);
or OR4 (N1908, N1905, N564, N1792, N1692);
nor NOR3 (N1909, N1904, N649, N896);
or OR3 (N1910, N1901, N1657, N201);
buf BUF1 (N1911, N1895);
nand NAND4 (N1912, N1911, N716, N397, N312);
or OR3 (N1913, N1910, N229, N1274);
and AND4 (N1914, N1888, N512, N1892, N981);
nand NAND4 (N1915, N1913, N73, N6, N552);
or OR2 (N1916, N1915, N1780);
nor NOR3 (N1917, N1903, N386, N325);
nand NAND3 (N1918, N1909, N212, N563);
nor NOR4 (N1919, N1906, N829, N1680, N530);
buf BUF1 (N1920, N1917);
nand NAND4 (N1921, N1919, N134, N1573, N1067);
nand NAND2 (N1922, N1914, N715);
and AND4 (N1923, N1916, N964, N1588, N1456);
and AND2 (N1924, N1920, N1020);
not NOT1 (N1925, N1907);
and AND3 (N1926, N1885, N1799, N506);
not NOT1 (N1927, N1912);
and AND2 (N1928, N1902, N199);
nor NOR4 (N1929, N1923, N204, N1438, N1579);
not NOT1 (N1930, N1929);
nor NOR2 (N1931, N1924, N1505);
and AND3 (N1932, N1922, N309, N1162);
xor XOR2 (N1933, N1925, N458);
xor XOR2 (N1934, N1926, N828);
and AND3 (N1935, N1918, N336, N576);
not NOT1 (N1936, N1933);
xor XOR2 (N1937, N1932, N309);
and AND3 (N1938, N1927, N1767, N374);
xor XOR2 (N1939, N1935, N930);
not NOT1 (N1940, N1921);
xor XOR2 (N1941, N1908, N748);
nand NAND4 (N1942, N1928, N1199, N1841, N574);
or OR3 (N1943, N1939, N789, N799);
not NOT1 (N1944, N1938);
buf BUF1 (N1945, N1930);
nand NAND2 (N1946, N1941, N868);
and AND3 (N1947, N1934, N820, N1482);
buf BUF1 (N1948, N1937);
nor NOR3 (N1949, N1947, N1767, N485);
buf BUF1 (N1950, N1944);
buf BUF1 (N1951, N1943);
buf BUF1 (N1952, N1946);
buf BUF1 (N1953, N1936);
buf BUF1 (N1954, N1950);
or OR4 (N1955, N1953, N1071, N1806, N1607);
nand NAND3 (N1956, N1954, N456, N1865);
xor XOR2 (N1957, N1949, N1061);
buf BUF1 (N1958, N1955);
not NOT1 (N1959, N1957);
xor XOR2 (N1960, N1952, N331);
xor XOR2 (N1961, N1942, N1391);
xor XOR2 (N1962, N1961, N506);
nand NAND2 (N1963, N1958, N1751);
not NOT1 (N1964, N1962);
nor NOR4 (N1965, N1959, N926, N732, N682);
not NOT1 (N1966, N1948);
and AND3 (N1967, N1964, N47, N1188);
buf BUF1 (N1968, N1967);
xor XOR2 (N1969, N1951, N602);
xor XOR2 (N1970, N1963, N1499);
buf BUF1 (N1971, N1931);
nor NOR2 (N1972, N1966, N927);
not NOT1 (N1973, N1968);
buf BUF1 (N1974, N1970);
or OR2 (N1975, N1940, N984);
buf BUF1 (N1976, N1971);
nor NOR4 (N1977, N1975, N1704, N876, N106);
or OR3 (N1978, N1969, N1565, N888);
xor XOR2 (N1979, N1976, N1017);
not NOT1 (N1980, N1979);
nand NAND4 (N1981, N1978, N680, N669, N517);
and AND2 (N1982, N1956, N1807);
nor NOR3 (N1983, N1972, N1963, N916);
xor XOR2 (N1984, N1980, N332);
xor XOR2 (N1985, N1983, N1220);
nand NAND4 (N1986, N1984, N1441, N1913, N1840);
not NOT1 (N1987, N1986);
nor NOR3 (N1988, N1985, N16, N216);
and AND4 (N1989, N1974, N1295, N24, N805);
not NOT1 (N1990, N1988);
and AND4 (N1991, N1990, N1148, N1849, N504);
xor XOR2 (N1992, N1977, N647);
and AND2 (N1993, N1945, N1188);
nand NAND2 (N1994, N1981, N355);
nand NAND4 (N1995, N1987, N1760, N1590, N980);
or OR3 (N1996, N1994, N1070, N1308);
or OR4 (N1997, N1996, N460, N1599, N1766);
nor NOR4 (N1998, N1993, N305, N836, N1287);
and AND2 (N1999, N1998, N413);
xor XOR2 (N2000, N1973, N143);
buf BUF1 (N2001, N1999);
nand NAND2 (N2002, N1991, N788);
nor NOR2 (N2003, N2001, N544);
or OR3 (N2004, N2000, N366, N728);
not NOT1 (N2005, N1960);
and AND4 (N2006, N1992, N924, N502, N1458);
nor NOR4 (N2007, N2002, N81, N1528, N875);
and AND2 (N2008, N1989, N1270);
nand NAND2 (N2009, N1997, N401);
and AND2 (N2010, N1982, N1179);
xor XOR2 (N2011, N2003, N372);
buf BUF1 (N2012, N2011);
xor XOR2 (N2013, N2009, N187);
buf BUF1 (N2014, N1965);
nand NAND4 (N2015, N1995, N930, N1983, N1993);
xor XOR2 (N2016, N2006, N1969);
nand NAND4 (N2017, N2004, N487, N1974, N70);
buf BUF1 (N2018, N2008);
nor NOR2 (N2019, N2018, N1462);
not NOT1 (N2020, N2015);
nand NAND2 (N2021, N2020, N880);
nand NAND4 (N2022, N2007, N891, N752, N1015);
buf BUF1 (N2023, N2022);
xor XOR2 (N2024, N2023, N89);
not NOT1 (N2025, N2010);
and AND3 (N2026, N2021, N1912, N848);
or OR3 (N2027, N2005, N1079, N139);
xor XOR2 (N2028, N2027, N1021);
nor NOR3 (N2029, N2016, N662, N1783);
or OR3 (N2030, N2026, N1034, N1453);
nand NAND2 (N2031, N2012, N1528);
nor NOR2 (N2032, N2019, N1465);
xor XOR2 (N2033, N2024, N1787);
or OR3 (N2034, N2028, N295, N1563);
nor NOR3 (N2035, N2017, N1079, N1665);
and AND3 (N2036, N2034, N1814, N1892);
xor XOR2 (N2037, N2029, N291);
or OR2 (N2038, N2014, N1886);
xor XOR2 (N2039, N2030, N2007);
not NOT1 (N2040, N2039);
nand NAND3 (N2041, N2033, N1307, N1033);
xor XOR2 (N2042, N2041, N1789);
buf BUF1 (N2043, N2040);
buf BUF1 (N2044, N2035);
or OR4 (N2045, N2013, N1527, N1965, N422);
and AND2 (N2046, N2036, N1957);
and AND4 (N2047, N2031, N1741, N1003, N1592);
nor NOR3 (N2048, N2045, N1322, N1708);
not NOT1 (N2049, N2047);
not NOT1 (N2050, N2042);
nor NOR3 (N2051, N2048, N1364, N1426);
and AND3 (N2052, N2046, N1986, N875);
or OR3 (N2053, N2052, N323, N748);
nor NOR3 (N2054, N2037, N252, N1395);
nor NOR3 (N2055, N2032, N1839, N1199);
and AND2 (N2056, N2043, N722);
or OR3 (N2057, N2038, N1782, N1258);
buf BUF1 (N2058, N2053);
nor NOR4 (N2059, N2057, N431, N1604, N900);
buf BUF1 (N2060, N2056);
buf BUF1 (N2061, N2051);
nand NAND2 (N2062, N2055, N722);
xor XOR2 (N2063, N2061, N264);
xor XOR2 (N2064, N2054, N685);
xor XOR2 (N2065, N2060, N1202);
nor NOR3 (N2066, N2058, N1011, N57);
nand NAND2 (N2067, N2025, N107);
and AND3 (N2068, N2064, N426, N983);
xor XOR2 (N2069, N2066, N335);
nor NOR3 (N2070, N2067, N301, N1952);
not NOT1 (N2071, N2062);
or OR2 (N2072, N2063, N566);
and AND2 (N2073, N2059, N17);
nor NOR2 (N2074, N2044, N1807);
nor NOR3 (N2075, N2070, N160, N999);
xor XOR2 (N2076, N2065, N1527);
buf BUF1 (N2077, N2073);
nand NAND3 (N2078, N2068, N231, N48);
nand NAND2 (N2079, N2075, N542);
nand NAND2 (N2080, N2076, N692);
xor XOR2 (N2081, N2074, N131);
nand NAND4 (N2082, N2069, N51, N1148, N718);
buf BUF1 (N2083, N2072);
nor NOR3 (N2084, N2080, N1465, N391);
xor XOR2 (N2085, N2084, N1440);
not NOT1 (N2086, N2083);
nand NAND2 (N2087, N2078, N1621);
nand NAND2 (N2088, N2077, N419);
not NOT1 (N2089, N2087);
nor NOR4 (N2090, N2079, N603, N1666, N268);
or OR3 (N2091, N2081, N72, N481);
or OR4 (N2092, N2091, N1063, N111, N1809);
not NOT1 (N2093, N2071);
xor XOR2 (N2094, N2088, N1614);
and AND4 (N2095, N2082, N1673, N825, N1100);
buf BUF1 (N2096, N2092);
nand NAND2 (N2097, N2094, N535);
not NOT1 (N2098, N2086);
buf BUF1 (N2099, N2098);
not NOT1 (N2100, N2097);
and AND4 (N2101, N2089, N1868, N362, N1398);
or OR2 (N2102, N2099, N1015);
and AND3 (N2103, N2050, N546, N532);
not NOT1 (N2104, N2049);
or OR4 (N2105, N2095, N1989, N600, N650);
and AND2 (N2106, N2096, N592);
and AND4 (N2107, N2103, N2065, N846, N301);
nand NAND2 (N2108, N2106, N978);
xor XOR2 (N2109, N2108, N486);
not NOT1 (N2110, N2085);
not NOT1 (N2111, N2110);
and AND3 (N2112, N2090, N1179, N1604);
nor NOR4 (N2113, N2093, N647, N712, N979);
not NOT1 (N2114, N2105);
nand NAND4 (N2115, N2112, N758, N1194, N1643);
or OR4 (N2116, N2102, N2028, N1096, N1641);
nand NAND2 (N2117, N2114, N50);
not NOT1 (N2118, N2109);
xor XOR2 (N2119, N2118, N1590);
nand NAND3 (N2120, N2100, N1004, N392);
or OR4 (N2121, N2119, N145, N2024, N30);
nor NOR3 (N2122, N2115, N496, N2021);
nand NAND2 (N2123, N2111, N1524);
or OR2 (N2124, N2116, N592);
xor XOR2 (N2125, N2124, N998);
xor XOR2 (N2126, N2107, N151);
buf BUF1 (N2127, N2113);
xor XOR2 (N2128, N2123, N361);
buf BUF1 (N2129, N2122);
nand NAND4 (N2130, N2129, N212, N1990, N646);
xor XOR2 (N2131, N2121, N751);
and AND3 (N2132, N2101, N227, N1302);
and AND4 (N2133, N2104, N1237, N1708, N229);
and AND4 (N2134, N2125, N813, N388, N1731);
nand NAND3 (N2135, N2117, N1026, N619);
or OR3 (N2136, N2131, N413, N1949);
and AND2 (N2137, N2127, N1982);
xor XOR2 (N2138, N2132, N1904);
buf BUF1 (N2139, N2137);
or OR3 (N2140, N2138, N963, N312);
nand NAND2 (N2141, N2139, N1338);
not NOT1 (N2142, N2128);
buf BUF1 (N2143, N2133);
not NOT1 (N2144, N2134);
or OR2 (N2145, N2141, N1301);
buf BUF1 (N2146, N2144);
buf BUF1 (N2147, N2142);
or OR4 (N2148, N2143, N1591, N319, N153);
or OR3 (N2149, N2135, N244, N1900);
not NOT1 (N2150, N2148);
and AND3 (N2151, N2136, N411, N1956);
xor XOR2 (N2152, N2151, N627);
or OR2 (N2153, N2130, N1646);
nor NOR4 (N2154, N2140, N1938, N657, N206);
not NOT1 (N2155, N2154);
or OR2 (N2156, N2120, N2052);
or OR3 (N2157, N2145, N25, N410);
or OR2 (N2158, N2155, N1903);
nor NOR4 (N2159, N2150, N743, N1211, N715);
not NOT1 (N2160, N2152);
xor XOR2 (N2161, N2157, N323);
and AND3 (N2162, N2149, N1587, N1560);
not NOT1 (N2163, N2146);
buf BUF1 (N2164, N2161);
nand NAND2 (N2165, N2159, N828);
xor XOR2 (N2166, N2147, N191);
or OR4 (N2167, N2160, N720, N175, N377);
nand NAND2 (N2168, N2163, N1373);
nor NOR4 (N2169, N2165, N2149, N1307, N664);
not NOT1 (N2170, N2162);
not NOT1 (N2171, N2153);
not NOT1 (N2172, N2168);
nand NAND2 (N2173, N2126, N215);
not NOT1 (N2174, N2173);
or OR4 (N2175, N2169, N1255, N37, N551);
not NOT1 (N2176, N2172);
and AND2 (N2177, N2176, N1729);
xor XOR2 (N2178, N2164, N789);
and AND3 (N2179, N2174, N1763, N527);
xor XOR2 (N2180, N2179, N1287);
not NOT1 (N2181, N2156);
xor XOR2 (N2182, N2166, N1274);
nand NAND2 (N2183, N2167, N233);
and AND4 (N2184, N2182, N1008, N1014, N1866);
xor XOR2 (N2185, N2177, N927);
nor NOR4 (N2186, N2170, N102, N1407, N919);
not NOT1 (N2187, N2178);
not NOT1 (N2188, N2181);
not NOT1 (N2189, N2183);
buf BUF1 (N2190, N2189);
nand NAND4 (N2191, N2188, N762, N2061, N870);
nor NOR2 (N2192, N2171, N1316);
and AND4 (N2193, N2158, N2055, N1340, N1427);
or OR3 (N2194, N2186, N638, N1742);
or OR3 (N2195, N2191, N1919, N1947);
nor NOR2 (N2196, N2187, N380);
buf BUF1 (N2197, N2192);
nor NOR2 (N2198, N2175, N1524);
or OR2 (N2199, N2185, N376);
not NOT1 (N2200, N2190);
nor NOR3 (N2201, N2194, N1697, N665);
not NOT1 (N2202, N2198);
or OR3 (N2203, N2193, N1599, N1229);
and AND2 (N2204, N2201, N1355);
buf BUF1 (N2205, N2199);
nor NOR4 (N2206, N2204, N1284, N1807, N948);
nor NOR3 (N2207, N2196, N2085, N1803);
xor XOR2 (N2208, N2206, N247);
not NOT1 (N2209, N2208);
and AND3 (N2210, N2209, N217, N832);
not NOT1 (N2211, N2210);
or OR3 (N2212, N2184, N2100, N100);
nor NOR4 (N2213, N2205, N1105, N14, N217);
buf BUF1 (N2214, N2195);
or OR4 (N2215, N2200, N1490, N1139, N1446);
or OR3 (N2216, N2207, N750, N342);
or OR2 (N2217, N2212, N832);
nor NOR3 (N2218, N2211, N922, N342);
or OR4 (N2219, N2213, N1020, N1246, N1614);
and AND3 (N2220, N2215, N1550, N805);
nor NOR2 (N2221, N2217, N2169);
and AND4 (N2222, N2180, N1021, N1726, N2045);
xor XOR2 (N2223, N2219, N399);
xor XOR2 (N2224, N2221, N1757);
xor XOR2 (N2225, N2218, N1629);
xor XOR2 (N2226, N2225, N1248);
not NOT1 (N2227, N2223);
not NOT1 (N2228, N2216);
and AND4 (N2229, N2214, N1530, N1164, N1285);
xor XOR2 (N2230, N2203, N312);
buf BUF1 (N2231, N2229);
xor XOR2 (N2232, N2230, N244);
nor NOR2 (N2233, N2227, N454);
or OR3 (N2234, N2232, N276, N1273);
buf BUF1 (N2235, N2226);
xor XOR2 (N2236, N2235, N1913);
or OR2 (N2237, N2222, N1274);
nor NOR4 (N2238, N2236, N13, N1784, N558);
not NOT1 (N2239, N2234);
or OR2 (N2240, N2239, N130);
not NOT1 (N2241, N2240);
and AND4 (N2242, N2228, N1749, N2065, N63);
xor XOR2 (N2243, N2237, N996);
nor NOR4 (N2244, N2241, N1190, N1104, N1259);
xor XOR2 (N2245, N2242, N1374);
xor XOR2 (N2246, N2224, N965);
nand NAND4 (N2247, N2238, N1675, N1208, N2156);
or OR3 (N2248, N2244, N819, N1498);
xor XOR2 (N2249, N2197, N1435);
buf BUF1 (N2250, N2233);
buf BUF1 (N2251, N2248);
and AND4 (N2252, N2247, N1346, N462, N95);
xor XOR2 (N2253, N2245, N1126);
buf BUF1 (N2254, N2243);
and AND3 (N2255, N2246, N1387, N574);
nor NOR3 (N2256, N2253, N730, N533);
xor XOR2 (N2257, N2255, N2127);
buf BUF1 (N2258, N2251);
and AND3 (N2259, N2254, N1270, N1069);
and AND3 (N2260, N2231, N1317, N550);
and AND3 (N2261, N2202, N366, N104);
xor XOR2 (N2262, N2259, N489);
buf BUF1 (N2263, N2250);
not NOT1 (N2264, N2257);
buf BUF1 (N2265, N2264);
not NOT1 (N2266, N2261);
or OR2 (N2267, N2258, N179);
xor XOR2 (N2268, N2249, N885);
buf BUF1 (N2269, N2265);
and AND4 (N2270, N2260, N110, N495, N544);
buf BUF1 (N2271, N2252);
not NOT1 (N2272, N2271);
or OR4 (N2273, N2256, N66, N48, N1844);
nand NAND2 (N2274, N2263, N386);
buf BUF1 (N2275, N2267);
and AND4 (N2276, N2269, N1811, N1757, N2033);
nor NOR2 (N2277, N2275, N1064);
or OR4 (N2278, N2273, N821, N386, N319);
nor NOR2 (N2279, N2262, N2146);
not NOT1 (N2280, N2268);
buf BUF1 (N2281, N2274);
and AND3 (N2282, N2266, N518, N88);
nor NOR4 (N2283, N2270, N1687, N1742, N734);
nand NAND3 (N2284, N2272, N1594, N1585);
not NOT1 (N2285, N2283);
xor XOR2 (N2286, N2276, N2147);
buf BUF1 (N2287, N2281);
buf BUF1 (N2288, N2285);
nand NAND4 (N2289, N2286, N183, N247, N2248);
or OR2 (N2290, N2289, N1200);
not NOT1 (N2291, N2220);
and AND4 (N2292, N2282, N2279, N1513, N871);
or OR2 (N2293, N1434, N1634);
xor XOR2 (N2294, N2280, N1039);
nor NOR2 (N2295, N2277, N843);
or OR3 (N2296, N2287, N752, N1635);
and AND2 (N2297, N2295, N846);
nand NAND3 (N2298, N2290, N998, N441);
and AND3 (N2299, N2296, N1211, N1333);
and AND2 (N2300, N2288, N275);
xor XOR2 (N2301, N2284, N2128);
nand NAND2 (N2302, N2301, N550);
not NOT1 (N2303, N2302);
or OR3 (N2304, N2291, N351, N1146);
and AND4 (N2305, N2299, N2290, N1839, N193);
and AND4 (N2306, N2293, N777, N1034, N1135);
nor NOR2 (N2307, N2304, N827);
not NOT1 (N2308, N2298);
buf BUF1 (N2309, N2278);
buf BUF1 (N2310, N2306);
and AND4 (N2311, N2308, N73, N1456, N2292);
buf BUF1 (N2312, N641);
buf BUF1 (N2313, N2303);
nor NOR4 (N2314, N2297, N1691, N1561, N1093);
and AND3 (N2315, N2300, N1152, N1118);
and AND4 (N2316, N2312, N1769, N1621, N503);
and AND3 (N2317, N2314, N1433, N1850);
buf BUF1 (N2318, N2294);
and AND3 (N2319, N2315, N1926, N654);
xor XOR2 (N2320, N2307, N925);
nor NOR4 (N2321, N2313, N762, N582, N720);
or OR2 (N2322, N2317, N1071);
not NOT1 (N2323, N2319);
xor XOR2 (N2324, N2311, N82);
not NOT1 (N2325, N2318);
xor XOR2 (N2326, N2323, N1072);
buf BUF1 (N2327, N2326);
and AND4 (N2328, N2310, N912, N2113, N2042);
not NOT1 (N2329, N2320);
buf BUF1 (N2330, N2322);
and AND4 (N2331, N2309, N2262, N1944, N1961);
and AND4 (N2332, N2330, N937, N1615, N733);
and AND3 (N2333, N2324, N452, N314);
and AND3 (N2334, N2316, N374, N1636);
nor NOR3 (N2335, N2334, N771, N1063);
and AND3 (N2336, N2321, N1568, N2316);
or OR4 (N2337, N2325, N2032, N268, N1879);
not NOT1 (N2338, N2337);
nand NAND3 (N2339, N2333, N1740, N2091);
nand NAND2 (N2340, N2328, N1514);
or OR2 (N2341, N2335, N1404);
nor NOR2 (N2342, N2341, N633);
buf BUF1 (N2343, N2339);
not NOT1 (N2344, N2342);
or OR2 (N2345, N2336, N1272);
nor NOR3 (N2346, N2344, N1550, N1143);
xor XOR2 (N2347, N2340, N752);
and AND3 (N2348, N2327, N2070, N1993);
nand NAND4 (N2349, N2305, N196, N69, N943);
buf BUF1 (N2350, N2345);
buf BUF1 (N2351, N2350);
buf BUF1 (N2352, N2329);
nor NOR2 (N2353, N2332, N1047);
or OR4 (N2354, N2349, N944, N1732, N2052);
nor NOR4 (N2355, N2352, N251, N1498, N348);
and AND4 (N2356, N2338, N1396, N1814, N757);
nor NOR2 (N2357, N2351, N2226);
not NOT1 (N2358, N2346);
nor NOR2 (N2359, N2353, N1687);
nor NOR3 (N2360, N2356, N1677, N1926);
buf BUF1 (N2361, N2359);
nand NAND4 (N2362, N2355, N53, N1434, N1088);
xor XOR2 (N2363, N2343, N1570);
or OR2 (N2364, N2362, N2047);
nor NOR3 (N2365, N2360, N956, N2197);
nand NAND2 (N2366, N2331, N2221);
or OR4 (N2367, N2354, N1548, N1596, N1433);
buf BUF1 (N2368, N2357);
buf BUF1 (N2369, N2368);
or OR2 (N2370, N2361, N2260);
nand NAND4 (N2371, N2367, N405, N1792, N1489);
xor XOR2 (N2372, N2348, N459);
not NOT1 (N2373, N2370);
nand NAND3 (N2374, N2358, N335, N74);
nand NAND4 (N2375, N2364, N1972, N1240, N1301);
xor XOR2 (N2376, N2366, N1697);
xor XOR2 (N2377, N2372, N694);
xor XOR2 (N2378, N2373, N1430);
or OR3 (N2379, N2363, N63, N1000);
xor XOR2 (N2380, N2374, N185);
and AND3 (N2381, N2347, N788, N2163);
nor NOR3 (N2382, N2381, N488, N78);
not NOT1 (N2383, N2377);
nor NOR3 (N2384, N2369, N1364, N1355);
or OR3 (N2385, N2375, N862, N789);
or OR3 (N2386, N2380, N1337, N1141);
or OR2 (N2387, N2385, N1472);
nand NAND2 (N2388, N2376, N134);
nand NAND4 (N2389, N2382, N1376, N728, N530);
or OR2 (N2390, N2371, N484);
nand NAND2 (N2391, N2390, N896);
and AND4 (N2392, N2391, N453, N89, N2185);
nor NOR2 (N2393, N2386, N1604);
xor XOR2 (N2394, N2389, N917);
not NOT1 (N2395, N2388);
nand NAND4 (N2396, N2387, N915, N2316, N307);
nand NAND4 (N2397, N2395, N1822, N144, N38);
buf BUF1 (N2398, N2384);
and AND4 (N2399, N2393, N1882, N564, N847);
nor NOR3 (N2400, N2383, N1676, N1368);
nand NAND4 (N2401, N2379, N439, N2349, N554);
xor XOR2 (N2402, N2378, N2090);
nor NOR2 (N2403, N2398, N1089);
buf BUF1 (N2404, N2400);
or OR3 (N2405, N2397, N824, N1565);
or OR2 (N2406, N2405, N1872);
nor NOR2 (N2407, N2404, N1726);
not NOT1 (N2408, N2407);
and AND3 (N2409, N2403, N478, N1479);
not NOT1 (N2410, N2392);
or OR4 (N2411, N2399, N1722, N1526, N1780);
nand NAND2 (N2412, N2365, N2327);
or OR2 (N2413, N2409, N1026);
nor NOR4 (N2414, N2411, N1509, N2047, N2074);
xor XOR2 (N2415, N2401, N1828);
buf BUF1 (N2416, N2402);
not NOT1 (N2417, N2415);
and AND4 (N2418, N2417, N1161, N1946, N1214);
not NOT1 (N2419, N2410);
nor NOR3 (N2420, N2396, N1866, N2103);
buf BUF1 (N2421, N2414);
not NOT1 (N2422, N2421);
xor XOR2 (N2423, N2420, N1847);
and AND3 (N2424, N2406, N2077, N1215);
xor XOR2 (N2425, N2416, N103);
xor XOR2 (N2426, N2394, N1169);
nand NAND3 (N2427, N2426, N267, N672);
not NOT1 (N2428, N2423);
xor XOR2 (N2429, N2418, N754);
not NOT1 (N2430, N2428);
or OR3 (N2431, N2424, N1025, N1006);
xor XOR2 (N2432, N2419, N682);
nand NAND4 (N2433, N2430, N87, N1747, N1893);
nor NOR2 (N2434, N2413, N174);
nand NAND4 (N2435, N2412, N330, N803, N475);
nor NOR3 (N2436, N2429, N1216, N320);
and AND2 (N2437, N2435, N1888);
buf BUF1 (N2438, N2432);
nor NOR3 (N2439, N2422, N229, N194);
nor NOR2 (N2440, N2434, N715);
xor XOR2 (N2441, N2439, N1869);
and AND4 (N2442, N2438, N703, N432, N628);
xor XOR2 (N2443, N2437, N1969);
nor NOR2 (N2444, N2431, N1393);
and AND2 (N2445, N2444, N112);
nor NOR4 (N2446, N2442, N977, N2413, N33);
nand NAND3 (N2447, N2425, N1995, N218);
nand NAND3 (N2448, N2427, N349, N54);
nand NAND4 (N2449, N2441, N1899, N1001, N552);
buf BUF1 (N2450, N2408);
nor NOR4 (N2451, N2443, N916, N1106, N59);
not NOT1 (N2452, N2451);
or OR2 (N2453, N2433, N2185);
and AND2 (N2454, N2445, N1818);
not NOT1 (N2455, N2454);
not NOT1 (N2456, N2450);
and AND4 (N2457, N2446, N1427, N2412, N695);
not NOT1 (N2458, N2456);
buf BUF1 (N2459, N2449);
buf BUF1 (N2460, N2448);
xor XOR2 (N2461, N2458, N1400);
or OR4 (N2462, N2436, N964, N1658, N605);
nand NAND4 (N2463, N2457, N488, N2057, N1133);
xor XOR2 (N2464, N2460, N2112);
nand NAND2 (N2465, N2463, N1154);
or OR2 (N2466, N2462, N2067);
nor NOR4 (N2467, N2452, N531, N1113, N1050);
and AND4 (N2468, N2464, N537, N22, N2051);
or OR3 (N2469, N2459, N1632, N46);
buf BUF1 (N2470, N2461);
or OR3 (N2471, N2440, N750, N540);
nand NAND4 (N2472, N2468, N1734, N1670, N944);
nand NAND2 (N2473, N2455, N1566);
and AND2 (N2474, N2447, N1506);
and AND2 (N2475, N2470, N92);
nor NOR4 (N2476, N2466, N383, N871, N1991);
nor NOR3 (N2477, N2472, N1251, N400);
nor NOR3 (N2478, N2467, N702, N467);
not NOT1 (N2479, N2477);
buf BUF1 (N2480, N2475);
nor NOR4 (N2481, N2471, N2260, N753, N2141);
and AND3 (N2482, N2465, N1498, N2153);
buf BUF1 (N2483, N2479);
nand NAND4 (N2484, N2483, N1301, N103, N557);
nor NOR3 (N2485, N2473, N1012, N1695);
xor XOR2 (N2486, N2481, N114);
buf BUF1 (N2487, N2453);
and AND2 (N2488, N2478, N1634);
nand NAND4 (N2489, N2482, N749, N2061, N1084);
buf BUF1 (N2490, N2476);
xor XOR2 (N2491, N2480, N1216);
xor XOR2 (N2492, N2484, N17);
not NOT1 (N2493, N2488);
buf BUF1 (N2494, N2489);
xor XOR2 (N2495, N2474, N1407);
and AND2 (N2496, N2493, N1346);
xor XOR2 (N2497, N2469, N1585);
nor NOR4 (N2498, N2496, N238, N1855, N552);
nor NOR4 (N2499, N2490, N43, N113, N150);
xor XOR2 (N2500, N2495, N1692);
nand NAND2 (N2501, N2491, N1438);
not NOT1 (N2502, N2499);
not NOT1 (N2503, N2494);
buf BUF1 (N2504, N2503);
xor XOR2 (N2505, N2485, N2189);
not NOT1 (N2506, N2504);
xor XOR2 (N2507, N2497, N829);
buf BUF1 (N2508, N2498);
or OR3 (N2509, N2486, N2152, N2421);
buf BUF1 (N2510, N2508);
xor XOR2 (N2511, N2500, N2145);
and AND2 (N2512, N2506, N1040);
xor XOR2 (N2513, N2507, N876);
nand NAND3 (N2514, N2502, N1973, N1402);
and AND4 (N2515, N2501, N545, N457, N757);
nand NAND2 (N2516, N2510, N1358);
not NOT1 (N2517, N2514);
buf BUF1 (N2518, N2509);
not NOT1 (N2519, N2515);
not NOT1 (N2520, N2519);
or OR4 (N2521, N2517, N1074, N642, N2205);
or OR4 (N2522, N2511, N184, N1368, N1028);
nand NAND3 (N2523, N2513, N915, N277);
buf BUF1 (N2524, N2520);
nor NOR4 (N2525, N2516, N1987, N110, N1786);
or OR2 (N2526, N2492, N792);
not NOT1 (N2527, N2521);
buf BUF1 (N2528, N2523);
or OR4 (N2529, N2512, N2305, N2437, N1294);
not NOT1 (N2530, N2527);
not NOT1 (N2531, N2522);
or OR4 (N2532, N2518, N1232, N2040, N1009);
not NOT1 (N2533, N2524);
xor XOR2 (N2534, N2531, N2321);
nand NAND2 (N2535, N2530, N2326);
xor XOR2 (N2536, N2487, N2266);
nand NAND3 (N2537, N2532, N964, N2423);
or OR2 (N2538, N2533, N791);
buf BUF1 (N2539, N2505);
not NOT1 (N2540, N2539);
or OR3 (N2541, N2529, N252, N727);
and AND4 (N2542, N2528, N1904, N2299, N1602);
nor NOR3 (N2543, N2526, N1306, N1980);
not NOT1 (N2544, N2542);
or OR2 (N2545, N2537, N1809);
buf BUF1 (N2546, N2545);
nor NOR2 (N2547, N2534, N2063);
xor XOR2 (N2548, N2544, N1434);
xor XOR2 (N2549, N2546, N1900);
xor XOR2 (N2550, N2541, N540);
nand NAND2 (N2551, N2543, N853);
xor XOR2 (N2552, N2548, N1944);
nor NOR4 (N2553, N2547, N2014, N2218, N1866);
nor NOR4 (N2554, N2540, N2309, N62, N891);
xor XOR2 (N2555, N2550, N843);
nor NOR2 (N2556, N2536, N190);
or OR2 (N2557, N2555, N591);
nor NOR2 (N2558, N2538, N1937);
xor XOR2 (N2559, N2553, N1643);
nand NAND4 (N2560, N2535, N1355, N1265, N1788);
xor XOR2 (N2561, N2551, N922);
or OR2 (N2562, N2554, N106);
buf BUF1 (N2563, N2557);
buf BUF1 (N2564, N2552);
buf BUF1 (N2565, N2559);
nor NOR2 (N2566, N2549, N804);
or OR3 (N2567, N2566, N1753, N1963);
and AND3 (N2568, N2560, N1683, N2244);
or OR3 (N2569, N2562, N791, N2337);
nand NAND4 (N2570, N2556, N2039, N1995, N1689);
xor XOR2 (N2571, N2561, N506);
or OR4 (N2572, N2525, N1097, N100, N995);
and AND2 (N2573, N2558, N2120);
not NOT1 (N2574, N2571);
xor XOR2 (N2575, N2568, N566);
nor NOR3 (N2576, N2565, N2066, N484);
xor XOR2 (N2577, N2575, N2230);
nand NAND3 (N2578, N2572, N2576, N35);
nor NOR2 (N2579, N835, N2457);
and AND3 (N2580, N2570, N843, N1058);
and AND2 (N2581, N2580, N186);
nor NOR4 (N2582, N2563, N1424, N1507, N322);
or OR4 (N2583, N2567, N2330, N1433, N2019);
nor NOR2 (N2584, N2574, N1427);
nor NOR2 (N2585, N2577, N1105);
nor NOR3 (N2586, N2573, N1464, N1175);
xor XOR2 (N2587, N2583, N1545);
nor NOR4 (N2588, N2586, N58, N1378, N147);
not NOT1 (N2589, N2569);
or OR3 (N2590, N2589, N285, N599);
not NOT1 (N2591, N2582);
not NOT1 (N2592, N2588);
not NOT1 (N2593, N2590);
not NOT1 (N2594, N2587);
or OR3 (N2595, N2564, N792, N2558);
nand NAND3 (N2596, N2593, N422, N2127);
buf BUF1 (N2597, N2585);
and AND4 (N2598, N2584, N2230, N1640, N75);
buf BUF1 (N2599, N2597);
and AND2 (N2600, N2578, N517);
buf BUF1 (N2601, N2600);
and AND4 (N2602, N2579, N536, N2275, N2068);
not NOT1 (N2603, N2602);
or OR2 (N2604, N2603, N2294);
and AND2 (N2605, N2604, N602);
xor XOR2 (N2606, N2601, N2155);
or OR4 (N2607, N2596, N1966, N1598, N465);
buf BUF1 (N2608, N2607);
nor NOR3 (N2609, N2599, N1524, N1218);
or OR4 (N2610, N2598, N767, N2085, N1915);
nor NOR2 (N2611, N2610, N1637);
nor NOR4 (N2612, N2611, N2072, N579, N566);
nand NAND4 (N2613, N2595, N465, N1168, N824);
nand NAND3 (N2614, N2594, N1177, N964);
buf BUF1 (N2615, N2581);
xor XOR2 (N2616, N2605, N87);
not NOT1 (N2617, N2613);
nand NAND2 (N2618, N2608, N2492);
nor NOR3 (N2619, N2606, N30, N247);
buf BUF1 (N2620, N2617);
buf BUF1 (N2621, N2616);
and AND3 (N2622, N2609, N1013, N948);
and AND4 (N2623, N2614, N1280, N2036, N1922);
or OR3 (N2624, N2619, N155, N1805);
buf BUF1 (N2625, N2615);
xor XOR2 (N2626, N2612, N2377);
or OR3 (N2627, N2625, N1245, N1380);
buf BUF1 (N2628, N2622);
not NOT1 (N2629, N2618);
not NOT1 (N2630, N2626);
not NOT1 (N2631, N2624);
buf BUF1 (N2632, N2621);
nand NAND3 (N2633, N2630, N355, N1059);
nand NAND4 (N2634, N2633, N475, N1053, N887);
nand NAND2 (N2635, N2592, N2396);
buf BUF1 (N2636, N2620);
and AND4 (N2637, N2632, N703, N1799, N127);
or OR4 (N2638, N2623, N1023, N1536, N1486);
not NOT1 (N2639, N2628);
not NOT1 (N2640, N2637);
nor NOR2 (N2641, N2635, N1244);
nand NAND2 (N2642, N2636, N2479);
and AND3 (N2643, N2629, N807, N1264);
or OR4 (N2644, N2639, N2630, N1127, N1047);
xor XOR2 (N2645, N2631, N1241);
not NOT1 (N2646, N2591);
and AND2 (N2647, N2641, N367);
buf BUF1 (N2648, N2646);
nand NAND3 (N2649, N2640, N2250, N810);
not NOT1 (N2650, N2647);
nand NAND2 (N2651, N2648, N237);
nor NOR2 (N2652, N2644, N985);
and AND3 (N2653, N2650, N847, N2399);
or OR2 (N2654, N2634, N2357);
and AND3 (N2655, N2653, N2111, N2191);
or OR3 (N2656, N2627, N738, N2633);
or OR2 (N2657, N2655, N42);
or OR4 (N2658, N2638, N1166, N1563, N1570);
nor NOR3 (N2659, N2652, N1813, N1419);
or OR4 (N2660, N2656, N1990, N2413, N544);
nand NAND2 (N2661, N2657, N337);
and AND2 (N2662, N2660, N1030);
and AND3 (N2663, N2658, N2517, N1007);
buf BUF1 (N2664, N2654);
xor XOR2 (N2665, N2664, N1954);
buf BUF1 (N2666, N2665);
and AND4 (N2667, N2659, N187, N127, N2397);
or OR4 (N2668, N2661, N523, N2458, N2284);
and AND4 (N2669, N2645, N470, N882, N1670);
xor XOR2 (N2670, N2668, N688);
nor NOR3 (N2671, N2669, N1133, N1223);
and AND3 (N2672, N2642, N1274, N2403);
xor XOR2 (N2673, N2651, N492);
nand NAND4 (N2674, N2643, N2597, N2356, N2430);
not NOT1 (N2675, N2663);
nor NOR4 (N2676, N2670, N2093, N1281, N830);
not NOT1 (N2677, N2649);
xor XOR2 (N2678, N2671, N1998);
or OR4 (N2679, N2677, N2053, N1002, N604);
nor NOR4 (N2680, N2679, N575, N302, N1483);
xor XOR2 (N2681, N2678, N1220);
nand NAND3 (N2682, N2673, N199, N1929);
and AND3 (N2683, N2681, N1231, N266);
xor XOR2 (N2684, N2682, N1569);
nand NAND2 (N2685, N2674, N2133);
buf BUF1 (N2686, N2676);
xor XOR2 (N2687, N2667, N623);
and AND3 (N2688, N2685, N1782, N1084);
xor XOR2 (N2689, N2684, N778);
nor NOR4 (N2690, N2687, N2053, N324, N377);
xor XOR2 (N2691, N2686, N2247);
buf BUF1 (N2692, N2666);
not NOT1 (N2693, N2662);
or OR3 (N2694, N2672, N1431, N1660);
buf BUF1 (N2695, N2680);
not NOT1 (N2696, N2683);
buf BUF1 (N2697, N2675);
nand NAND4 (N2698, N2696, N344, N1271, N2172);
xor XOR2 (N2699, N2693, N1556);
not NOT1 (N2700, N2690);
not NOT1 (N2701, N2695);
buf BUF1 (N2702, N2700);
and AND3 (N2703, N2692, N643, N2358);
buf BUF1 (N2704, N2698);
not NOT1 (N2705, N2689);
nor NOR2 (N2706, N2688, N675);
not NOT1 (N2707, N2691);
buf BUF1 (N2708, N2706);
or OR4 (N2709, N2702, N2357, N257, N1417);
nor NOR4 (N2710, N2697, N712, N297, N2580);
xor XOR2 (N2711, N2707, N1853);
nor NOR3 (N2712, N2699, N2670, N2451);
not NOT1 (N2713, N2710);
nor NOR2 (N2714, N2703, N2659);
or OR4 (N2715, N2708, N2100, N741, N455);
and AND4 (N2716, N2694, N750, N1108, N2437);
not NOT1 (N2717, N2715);
nand NAND4 (N2718, N2713, N1735, N370, N2416);
or OR3 (N2719, N2714, N1366, N157);
and AND3 (N2720, N2712, N1885, N1145);
nor NOR3 (N2721, N2718, N2097, N439);
and AND3 (N2722, N2720, N287, N793);
not NOT1 (N2723, N2719);
nor NOR4 (N2724, N2709, N1322, N2273, N526);
not NOT1 (N2725, N2724);
buf BUF1 (N2726, N2717);
nand NAND3 (N2727, N2705, N2544, N2667);
and AND3 (N2728, N2723, N1052, N749);
not NOT1 (N2729, N2716);
xor XOR2 (N2730, N2711, N1898);
nor NOR3 (N2731, N2727, N614, N585);
buf BUF1 (N2732, N2704);
or OR4 (N2733, N2726, N1048, N1110, N788);
nor NOR3 (N2734, N2701, N1202, N2245);
xor XOR2 (N2735, N2731, N1595);
not NOT1 (N2736, N2735);
xor XOR2 (N2737, N2728, N1601);
nand NAND4 (N2738, N2730, N1852, N123, N600);
and AND4 (N2739, N2738, N1530, N2283, N2206);
or OR4 (N2740, N2739, N1131, N1994, N1251);
buf BUF1 (N2741, N2721);
not NOT1 (N2742, N2741);
and AND3 (N2743, N2734, N112, N695);
nor NOR2 (N2744, N2737, N1447);
xor XOR2 (N2745, N2733, N1594);
and AND3 (N2746, N2736, N169, N714);
not NOT1 (N2747, N2743);
nand NAND4 (N2748, N2740, N2613, N2287, N1823);
not NOT1 (N2749, N2746);
nand NAND2 (N2750, N2747, N1996);
not NOT1 (N2751, N2744);
or OR4 (N2752, N2725, N211, N1315, N312);
nand NAND3 (N2753, N2752, N491, N1352);
xor XOR2 (N2754, N2722, N1257);
xor XOR2 (N2755, N2732, N2334);
xor XOR2 (N2756, N2754, N664);
or OR4 (N2757, N2749, N2499, N1592, N1646);
xor XOR2 (N2758, N2748, N1295);
or OR4 (N2759, N2753, N889, N919, N1787);
nand NAND2 (N2760, N2757, N2735);
or OR2 (N2761, N2758, N731);
not NOT1 (N2762, N2751);
buf BUF1 (N2763, N2762);
xor XOR2 (N2764, N2729, N2755);
or OR2 (N2765, N2312, N213);
nor NOR4 (N2766, N2764, N1946, N2123, N2658);
nor NOR4 (N2767, N2745, N282, N795, N205);
and AND2 (N2768, N2742, N711);
buf BUF1 (N2769, N2766);
or OR2 (N2770, N2765, N47);
not NOT1 (N2771, N2760);
and AND2 (N2772, N2771, N625);
not NOT1 (N2773, N2767);
and AND2 (N2774, N2761, N1942);
nor NOR3 (N2775, N2773, N2592, N1023);
not NOT1 (N2776, N2763);
not NOT1 (N2777, N2770);
and AND4 (N2778, N2775, N1693, N395, N283);
or OR3 (N2779, N2777, N1224, N1789);
buf BUF1 (N2780, N2779);
not NOT1 (N2781, N2769);
and AND4 (N2782, N2768, N1434, N1971, N477);
or OR4 (N2783, N2781, N2320, N2178, N2466);
and AND3 (N2784, N2759, N1207, N1244);
buf BUF1 (N2785, N2774);
nor NOR4 (N2786, N2756, N286, N653, N1857);
or OR3 (N2787, N2782, N1286, N1461);
and AND2 (N2788, N2750, N1424);
nor NOR3 (N2789, N2787, N1672, N1659);
nand NAND4 (N2790, N2789, N1983, N1360, N2393);
buf BUF1 (N2791, N2776);
not NOT1 (N2792, N2784);
buf BUF1 (N2793, N2788);
or OR4 (N2794, N2780, N2683, N243, N1695);
xor XOR2 (N2795, N2792, N1098);
nor NOR3 (N2796, N2793, N1187, N1431);
xor XOR2 (N2797, N2791, N66);
not NOT1 (N2798, N2783);
not NOT1 (N2799, N2798);
nor NOR2 (N2800, N2785, N802);
xor XOR2 (N2801, N2790, N280);
buf BUF1 (N2802, N2801);
xor XOR2 (N2803, N2797, N510);
nor NOR2 (N2804, N2799, N645);
and AND4 (N2805, N2795, N1420, N2069, N2383);
nand NAND4 (N2806, N2802, N1724, N130, N1247);
and AND4 (N2807, N2796, N2279, N956, N362);
not NOT1 (N2808, N2800);
nand NAND3 (N2809, N2794, N1556, N815);
and AND2 (N2810, N2806, N448);
buf BUF1 (N2811, N2808);
not NOT1 (N2812, N2807);
or OR4 (N2813, N2809, N1762, N2495, N714);
and AND3 (N2814, N2813, N18, N755);
nor NOR2 (N2815, N2778, N1554);
buf BUF1 (N2816, N2804);
xor XOR2 (N2817, N2810, N1631);
xor XOR2 (N2818, N2814, N397);
buf BUF1 (N2819, N2803);
xor XOR2 (N2820, N2815, N558);
xor XOR2 (N2821, N2817, N1803);
nand NAND2 (N2822, N2805, N275);
buf BUF1 (N2823, N2811);
nor NOR4 (N2824, N2812, N1824, N2061, N1027);
xor XOR2 (N2825, N2816, N1372);
buf BUF1 (N2826, N2786);
nand NAND4 (N2827, N2772, N2524, N66, N543);
nand NAND3 (N2828, N2826, N1893, N1765);
or OR2 (N2829, N2824, N1263);
xor XOR2 (N2830, N2821, N1375);
nand NAND2 (N2831, N2819, N2083);
xor XOR2 (N2832, N2818, N211);
nand NAND2 (N2833, N2825, N1105);
nor NOR4 (N2834, N2828, N77, N316, N121);
or OR4 (N2835, N2830, N1293, N1045, N2235);
or OR3 (N2836, N2827, N1617, N29);
nand NAND2 (N2837, N2836, N2408);
not NOT1 (N2838, N2822);
not NOT1 (N2839, N2838);
not NOT1 (N2840, N2829);
or OR2 (N2841, N2832, N273);
buf BUF1 (N2842, N2834);
xor XOR2 (N2843, N2841, N1496);
xor XOR2 (N2844, N2833, N2111);
buf BUF1 (N2845, N2842);
buf BUF1 (N2846, N2835);
xor XOR2 (N2847, N2843, N2097);
nor NOR3 (N2848, N2837, N563, N2460);
xor XOR2 (N2849, N2840, N2825);
not NOT1 (N2850, N2820);
xor XOR2 (N2851, N2844, N2324);
and AND3 (N2852, N2847, N1219, N1846);
not NOT1 (N2853, N2839);
nand NAND3 (N2854, N2850, N1350, N2673);
xor XOR2 (N2855, N2823, N195);
nor NOR2 (N2856, N2831, N1482);
not NOT1 (N2857, N2854);
or OR4 (N2858, N2846, N679, N1995, N1682);
xor XOR2 (N2859, N2856, N2752);
nand NAND3 (N2860, N2845, N781, N1653);
nand NAND4 (N2861, N2848, N2793, N1493, N2302);
nor NOR2 (N2862, N2861, N2395);
nor NOR2 (N2863, N2852, N2073);
nand NAND4 (N2864, N2860, N982, N2848, N1747);
or OR4 (N2865, N2862, N907, N1431, N2052);
not NOT1 (N2866, N2864);
and AND3 (N2867, N2866, N456, N816);
nor NOR2 (N2868, N2859, N2316);
or OR4 (N2869, N2865, N2778, N1086, N1164);
xor XOR2 (N2870, N2855, N1982);
xor XOR2 (N2871, N2863, N2676);
nor NOR2 (N2872, N2853, N1645);
or OR2 (N2873, N2868, N1023);
and AND3 (N2874, N2870, N2730, N1770);
buf BUF1 (N2875, N2857);
not NOT1 (N2876, N2873);
buf BUF1 (N2877, N2849);
and AND4 (N2878, N2872, N333, N1891, N2477);
nand NAND4 (N2879, N2867, N2202, N583, N1524);
or OR4 (N2880, N2874, N1348, N2576, N2879);
and AND3 (N2881, N2812, N488, N630);
and AND2 (N2882, N2876, N1740);
buf BUF1 (N2883, N2871);
buf BUF1 (N2884, N2882);
xor XOR2 (N2885, N2880, N1228);
nand NAND4 (N2886, N2878, N1447, N6, N194);
or OR4 (N2887, N2851, N748, N2652, N1790);
nand NAND2 (N2888, N2883, N1994);
buf BUF1 (N2889, N2877);
nor NOR3 (N2890, N2869, N2054, N301);
and AND2 (N2891, N2886, N2363);
xor XOR2 (N2892, N2887, N4);
xor XOR2 (N2893, N2858, N2756);
nand NAND2 (N2894, N2875, N427);
xor XOR2 (N2895, N2893, N2221);
nand NAND3 (N2896, N2888, N703, N1588);
nor NOR4 (N2897, N2894, N37, N2889, N1389);
buf BUF1 (N2898, N1352);
or OR2 (N2899, N2892, N754);
nand NAND3 (N2900, N2891, N2080, N1744);
nand NAND3 (N2901, N2899, N374, N2532);
nand NAND3 (N2902, N2881, N1757, N2306);
not NOT1 (N2903, N2900);
xor XOR2 (N2904, N2901, N2657);
not NOT1 (N2905, N2885);
nor NOR4 (N2906, N2890, N1550, N602, N2783);
not NOT1 (N2907, N2903);
buf BUF1 (N2908, N2898);
or OR2 (N2909, N2884, N314);
or OR3 (N2910, N2907, N1396, N2293);
nand NAND4 (N2911, N2897, N2456, N2523, N966);
nor NOR4 (N2912, N2909, N2672, N553, N2160);
xor XOR2 (N2913, N2910, N414);
nand NAND2 (N2914, N2906, N136);
nand NAND2 (N2915, N2911, N2217);
and AND2 (N2916, N2902, N2501);
and AND4 (N2917, N2913, N1884, N2138, N1084);
buf BUF1 (N2918, N2916);
nor NOR2 (N2919, N2918, N2720);
xor XOR2 (N2920, N2896, N2339);
nor NOR4 (N2921, N2905, N488, N2132, N1556);
buf BUF1 (N2922, N2904);
or OR2 (N2923, N2922, N2392);
not NOT1 (N2924, N2908);
buf BUF1 (N2925, N2895);
xor XOR2 (N2926, N2914, N868);
nand NAND3 (N2927, N2921, N2506, N1034);
not NOT1 (N2928, N2926);
and AND3 (N2929, N2927, N2843, N2437);
not NOT1 (N2930, N2923);
nor NOR3 (N2931, N2915, N1135, N1003);
and AND4 (N2932, N2931, N323, N1316, N1478);
or OR3 (N2933, N2932, N2716, N812);
and AND3 (N2934, N2924, N1513, N2812);
buf BUF1 (N2935, N2920);
nand NAND2 (N2936, N2919, N279);
xor XOR2 (N2937, N2934, N816);
not NOT1 (N2938, N2925);
nor NOR4 (N2939, N2929, N607, N1780, N562);
nor NOR2 (N2940, N2928, N2782);
nand NAND2 (N2941, N2938, N440);
nor NOR4 (N2942, N2917, N978, N1329, N693);
and AND4 (N2943, N2940, N2758, N1289, N2661);
and AND3 (N2944, N2941, N1166, N2586);
and AND2 (N2945, N2937, N2551);
and AND2 (N2946, N2945, N615);
nor NOR4 (N2947, N2912, N2817, N2246, N517);
nor NOR4 (N2948, N2933, N2573, N2153, N2652);
xor XOR2 (N2949, N2947, N2501);
nor NOR3 (N2950, N2936, N2209, N1486);
and AND4 (N2951, N2939, N1094, N2093, N2271);
or OR3 (N2952, N2951, N2509, N2603);
and AND4 (N2953, N2930, N2350, N1125, N1419);
or OR2 (N2954, N2949, N1511);
xor XOR2 (N2955, N2952, N1089);
not NOT1 (N2956, N2944);
or OR3 (N2957, N2935, N2543, N2307);
buf BUF1 (N2958, N2946);
and AND4 (N2959, N2948, N419, N2532, N261);
or OR2 (N2960, N2957, N1123);
and AND4 (N2961, N2955, N1666, N946, N1844);
nor NOR3 (N2962, N2954, N972, N47);
or OR2 (N2963, N2961, N1967);
nand NAND4 (N2964, N2953, N1278, N2770, N1327);
xor XOR2 (N2965, N2962, N237);
nor NOR3 (N2966, N2943, N1990, N1522);
and AND4 (N2967, N2958, N1881, N1941, N758);
nor NOR3 (N2968, N2965, N2741, N632);
and AND3 (N2969, N2963, N410, N114);
nand NAND4 (N2970, N2942, N1012, N2121, N1450);
not NOT1 (N2971, N2966);
xor XOR2 (N2972, N2968, N2752);
nand NAND4 (N2973, N2960, N2310, N733, N1684);
xor XOR2 (N2974, N2971, N1598);
nor NOR4 (N2975, N2967, N1227, N1437, N1669);
not NOT1 (N2976, N2972);
or OR2 (N2977, N2970, N198);
not NOT1 (N2978, N2977);
xor XOR2 (N2979, N2956, N1735);
nor NOR2 (N2980, N2979, N294);
nand NAND2 (N2981, N2964, N524);
nand NAND3 (N2982, N2976, N584, N740);
and AND3 (N2983, N2981, N39, N64);
and AND4 (N2984, N2959, N1471, N1685, N2191);
not NOT1 (N2985, N2950);
or OR3 (N2986, N2975, N84, N1864);
buf BUF1 (N2987, N2973);
xor XOR2 (N2988, N2969, N1986);
nand NAND4 (N2989, N2985, N1806, N1821, N730);
or OR4 (N2990, N2980, N1899, N2762, N1574);
buf BUF1 (N2991, N2984);
or OR4 (N2992, N2978, N1813, N165, N121);
or OR3 (N2993, N2989, N1072, N2991);
buf BUF1 (N2994, N1964);
xor XOR2 (N2995, N2986, N1546);
buf BUF1 (N2996, N2988);
nand NAND4 (N2997, N2996, N127, N2369, N1660);
buf BUF1 (N2998, N2995);
xor XOR2 (N2999, N2997, N1091);
not NOT1 (N3000, N2983);
xor XOR2 (N3001, N2994, N1163);
nor NOR2 (N3002, N3001, N983);
nand NAND3 (N3003, N2982, N608, N1796);
nand NAND2 (N3004, N3003, N433);
nand NAND3 (N3005, N3002, N2791, N1125);
and AND3 (N3006, N2992, N216, N2144);
xor XOR2 (N3007, N2993, N2525);
nand NAND4 (N3008, N3000, N994, N2564, N1149);
buf BUF1 (N3009, N3007);
nor NOR2 (N3010, N3008, N859);
xor XOR2 (N3011, N2974, N346);
not NOT1 (N3012, N3004);
xor XOR2 (N3013, N2987, N97);
nor NOR3 (N3014, N2998, N1396, N2224);
xor XOR2 (N3015, N2999, N2667);
or OR2 (N3016, N3010, N794);
buf BUF1 (N3017, N3006);
buf BUF1 (N3018, N3005);
and AND4 (N3019, N3018, N2924, N1392, N2638);
buf BUF1 (N3020, N3014);
endmodule