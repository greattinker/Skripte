// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15;

output N8002,N7994,N7993,N8013,N8005,N8011,N8004,N8014,N7999,N8015;

nand NAND2 (N16, N5, N8);
or OR4 (N17, N11, N6, N1, N5);
nor NOR4 (N18, N1, N6, N13, N16);
nand NAND2 (N19, N1, N5);
xor XOR2 (N20, N16, N14);
nor NOR4 (N21, N17, N11, N8, N12);
or OR3 (N22, N10, N1, N13);
xor XOR2 (N23, N8, N3);
nand NAND4 (N24, N19, N22, N1, N14);
and AND3 (N25, N17, N13, N2);
and AND3 (N26, N4, N5, N18);
nand NAND3 (N27, N11, N8, N16);
nor NOR3 (N28, N4, N17, N13);
buf BUF1 (N29, N23);
nor NOR3 (N30, N7, N2, N16);
not NOT1 (N31, N30);
or OR3 (N32, N23, N12, N8);
and AND3 (N33, N27, N5, N13);
and AND2 (N34, N31, N2);
buf BUF1 (N35, N34);
xor XOR2 (N36, N21, N11);
or OR2 (N37, N29, N7);
and AND4 (N38, N32, N16, N21, N23);
buf BUF1 (N39, N24);
or OR4 (N40, N39, N24, N22, N13);
xor XOR2 (N41, N40, N15);
or OR4 (N42, N37, N5, N24, N3);
not NOT1 (N43, N42);
nand NAND4 (N44, N25, N3, N42, N39);
not NOT1 (N45, N28);
and AND4 (N46, N43, N18, N21, N30);
not NOT1 (N47, N46);
or OR3 (N48, N38, N24, N26);
or OR3 (N49, N1, N41, N21);
nor NOR2 (N50, N4, N34);
buf BUF1 (N51, N47);
or OR3 (N52, N49, N8, N4);
and AND2 (N53, N33, N25);
nand NAND3 (N54, N35, N47, N32);
nand NAND4 (N55, N44, N44, N3, N9);
and AND4 (N56, N36, N52, N40, N33);
nand NAND2 (N57, N28, N29);
and AND4 (N58, N56, N1, N43, N33);
buf BUF1 (N59, N48);
and AND3 (N60, N55, N12, N42);
xor XOR2 (N61, N20, N14);
not NOT1 (N62, N50);
buf BUF1 (N63, N45);
not NOT1 (N64, N60);
nor NOR3 (N65, N64, N2, N19);
xor XOR2 (N66, N58, N25);
nand NAND2 (N67, N61, N31);
not NOT1 (N68, N59);
xor XOR2 (N69, N67, N17);
and AND4 (N70, N51, N31, N1, N36);
not NOT1 (N71, N69);
xor XOR2 (N72, N70, N7);
and AND4 (N73, N54, N6, N60, N44);
xor XOR2 (N74, N57, N31);
xor XOR2 (N75, N68, N6);
xor XOR2 (N76, N65, N66);
nand NAND2 (N77, N27, N7);
not NOT1 (N78, N71);
and AND3 (N79, N73, N72, N7);
or OR3 (N80, N26, N36, N53);
or OR2 (N81, N50, N66);
not NOT1 (N82, N79);
not NOT1 (N83, N62);
nand NAND2 (N84, N78, N56);
nand NAND2 (N85, N76, N37);
and AND4 (N86, N80, N48, N77, N12);
xor XOR2 (N87, N57, N52);
or OR4 (N88, N84, N33, N39, N14);
not NOT1 (N89, N81);
nor NOR3 (N90, N88, N28, N85);
not NOT1 (N91, N42);
or OR4 (N92, N75, N4, N83, N52);
not NOT1 (N93, N66);
xor XOR2 (N94, N86, N35);
nor NOR2 (N95, N91, N20);
or OR2 (N96, N82, N70);
buf BUF1 (N97, N95);
not NOT1 (N98, N92);
or OR2 (N99, N63, N84);
nor NOR2 (N100, N94, N30);
nor NOR2 (N101, N74, N88);
nor NOR3 (N102, N101, N38, N15);
buf BUF1 (N103, N100);
buf BUF1 (N104, N96);
nand NAND4 (N105, N90, N12, N83, N18);
xor XOR2 (N106, N89, N63);
xor XOR2 (N107, N93, N69);
not NOT1 (N108, N102);
not NOT1 (N109, N105);
and AND3 (N110, N106, N108, N42);
nor NOR3 (N111, N61, N7, N21);
and AND3 (N112, N99, N49, N4);
not NOT1 (N113, N87);
xor XOR2 (N114, N113, N99);
nor NOR4 (N115, N98, N7, N41, N61);
xor XOR2 (N116, N103, N112);
and AND2 (N117, N101, N88);
nand NAND3 (N118, N104, N55, N17);
and AND2 (N119, N116, N29);
xor XOR2 (N120, N111, N14);
xor XOR2 (N121, N97, N26);
and AND2 (N122, N114, N11);
and AND3 (N123, N122, N117, N7);
xor XOR2 (N124, N97, N68);
buf BUF1 (N125, N123);
nand NAND3 (N126, N107, N78, N56);
nor NOR3 (N127, N110, N16, N117);
nand NAND4 (N128, N125, N24, N52, N121);
buf BUF1 (N129, N124);
xor XOR2 (N130, N111, N108);
and AND3 (N131, N126, N66, N2);
not NOT1 (N132, N127);
not NOT1 (N133, N131);
nor NOR4 (N134, N115, N77, N18, N67);
and AND4 (N135, N134, N78, N26, N90);
and AND4 (N136, N133, N42, N117, N127);
buf BUF1 (N137, N130);
buf BUF1 (N138, N137);
or OR3 (N139, N109, N42, N28);
and AND2 (N140, N119, N117);
or OR3 (N141, N138, N110, N139);
nor NOR2 (N142, N26, N99);
xor XOR2 (N143, N129, N41);
nor NOR2 (N144, N135, N104);
and AND4 (N145, N136, N86, N79, N18);
not NOT1 (N146, N140);
nor NOR3 (N147, N141, N96, N141);
nor NOR3 (N148, N146, N60, N33);
xor XOR2 (N149, N147, N130);
nand NAND4 (N150, N132, N10, N43, N143);
nor NOR4 (N151, N35, N120, N44, N140);
xor XOR2 (N152, N115, N94);
or OR2 (N153, N118, N3);
xor XOR2 (N154, N145, N7);
not NOT1 (N155, N153);
and AND3 (N156, N142, N59, N89);
xor XOR2 (N157, N155, N22);
and AND4 (N158, N154, N101, N24, N113);
nand NAND3 (N159, N148, N4, N119);
and AND3 (N160, N159, N99, N121);
not NOT1 (N161, N157);
nor NOR3 (N162, N144, N32, N41);
nand NAND2 (N163, N158, N150);
and AND3 (N164, N1, N1, N40);
xor XOR2 (N165, N151, N84);
and AND2 (N166, N162, N46);
xor XOR2 (N167, N128, N98);
nand NAND4 (N168, N152, N146, N166, N1);
or OR4 (N169, N141, N9, N119, N48);
buf BUF1 (N170, N164);
buf BUF1 (N171, N167);
buf BUF1 (N172, N163);
xor XOR2 (N173, N169, N117);
or OR4 (N174, N165, N171, N49, N14);
or OR2 (N175, N81, N160);
xor XOR2 (N176, N154, N154);
not NOT1 (N177, N170);
and AND4 (N178, N156, N162, N170, N151);
xor XOR2 (N179, N178, N91);
not NOT1 (N180, N177);
or OR3 (N181, N179, N138, N25);
buf BUF1 (N182, N172);
buf BUF1 (N183, N149);
nand NAND3 (N184, N182, N36, N40);
xor XOR2 (N185, N176, N166);
or OR4 (N186, N173, N7, N104, N184);
nor NOR2 (N187, N70, N66);
and AND2 (N188, N174, N87);
xor XOR2 (N189, N186, N122);
nand NAND3 (N190, N175, N105, N56);
or OR2 (N191, N189, N144);
buf BUF1 (N192, N187);
and AND2 (N193, N190, N177);
xor XOR2 (N194, N181, N34);
and AND4 (N195, N188, N25, N20, N169);
xor XOR2 (N196, N193, N85);
and AND3 (N197, N194, N41, N183);
xor XOR2 (N198, N156, N143);
buf BUF1 (N199, N197);
not NOT1 (N200, N161);
and AND3 (N201, N192, N80, N17);
nand NAND2 (N202, N185, N137);
buf BUF1 (N203, N180);
buf BUF1 (N204, N203);
or OR4 (N205, N201, N189, N29, N122);
nor NOR4 (N206, N204, N152, N16, N182);
or OR2 (N207, N206, N90);
nor NOR3 (N208, N207, N17, N166);
not NOT1 (N209, N168);
and AND3 (N210, N195, N113, N200);
not NOT1 (N211, N187);
or OR3 (N212, N196, N35, N176);
nor NOR3 (N213, N210, N90, N62);
nand NAND2 (N214, N209, N116);
or OR3 (N215, N191, N156, N95);
and AND3 (N216, N208, N200, N95);
xor XOR2 (N217, N214, N97);
nor NOR3 (N218, N215, N65, N10);
nor NOR4 (N219, N213, N77, N140, N106);
or OR3 (N220, N199, N190, N139);
or OR3 (N221, N212, N119, N198);
xor XOR2 (N222, N64, N2);
nand NAND2 (N223, N211, N67);
and AND2 (N224, N221, N173);
buf BUF1 (N225, N224);
or OR4 (N226, N202, N101, N39, N211);
xor XOR2 (N227, N217, N191);
not NOT1 (N228, N223);
buf BUF1 (N229, N225);
buf BUF1 (N230, N228);
nand NAND3 (N231, N227, N92, N126);
not NOT1 (N232, N222);
buf BUF1 (N233, N219);
nor NOR3 (N234, N232, N231, N183);
nor NOR3 (N235, N199, N75, N52);
or OR2 (N236, N230, N186);
xor XOR2 (N237, N233, N174);
not NOT1 (N238, N216);
not NOT1 (N239, N205);
or OR3 (N240, N220, N47, N45);
and AND4 (N241, N218, N197, N71, N239);
buf BUF1 (N242, N20);
not NOT1 (N243, N241);
not NOT1 (N244, N229);
or OR3 (N245, N237, N212, N75);
buf BUF1 (N246, N236);
buf BUF1 (N247, N245);
nor NOR4 (N248, N243, N115, N101, N76);
or OR4 (N249, N226, N199, N202, N204);
and AND4 (N250, N242, N157, N205, N179);
and AND4 (N251, N240, N134, N192, N183);
xor XOR2 (N252, N234, N69);
or OR4 (N253, N247, N212, N200, N67);
not NOT1 (N254, N249);
nor NOR2 (N255, N253, N14);
xor XOR2 (N256, N255, N57);
not NOT1 (N257, N248);
xor XOR2 (N258, N238, N243);
nor NOR4 (N259, N235, N94, N67, N7);
not NOT1 (N260, N258);
buf BUF1 (N261, N244);
not NOT1 (N262, N260);
not NOT1 (N263, N262);
and AND2 (N264, N261, N75);
nand NAND4 (N265, N263, N93, N101, N139);
nand NAND4 (N266, N265, N55, N102, N152);
buf BUF1 (N267, N266);
nor NOR3 (N268, N257, N153, N179);
or OR3 (N269, N251, N81, N45);
not NOT1 (N270, N254);
nor NOR4 (N271, N246, N71, N262, N251);
nor NOR3 (N272, N252, N41, N239);
nor NOR2 (N273, N268, N54);
and AND2 (N274, N271, N101);
not NOT1 (N275, N273);
xor XOR2 (N276, N272, N60);
not NOT1 (N277, N269);
or OR3 (N278, N256, N94, N138);
and AND4 (N279, N276, N36, N177, N249);
nand NAND3 (N280, N274, N10, N208);
not NOT1 (N281, N259);
nor NOR2 (N282, N277, N209);
nand NAND2 (N283, N275, N128);
nand NAND2 (N284, N264, N233);
nand NAND2 (N285, N279, N146);
nand NAND4 (N286, N270, N253, N209, N33);
buf BUF1 (N287, N250);
not NOT1 (N288, N280);
or OR4 (N289, N284, N253, N272, N86);
xor XOR2 (N290, N288, N165);
and AND4 (N291, N285, N125, N264, N215);
xor XOR2 (N292, N281, N9);
and AND3 (N293, N286, N61, N213);
and AND4 (N294, N287, N85, N182, N204);
not NOT1 (N295, N294);
or OR4 (N296, N295, N284, N197, N87);
nor NOR2 (N297, N296, N12);
or OR2 (N298, N289, N71);
or OR4 (N299, N282, N206, N277, N198);
nor NOR3 (N300, N278, N195, N120);
xor XOR2 (N301, N300, N140);
nor NOR4 (N302, N301, N186, N250, N258);
or OR2 (N303, N302, N87);
nand NAND2 (N304, N267, N273);
nand NAND4 (N305, N297, N151, N153, N83);
not NOT1 (N306, N303);
xor XOR2 (N307, N292, N198);
buf BUF1 (N308, N293);
and AND2 (N309, N305, N241);
xor XOR2 (N310, N309, N229);
not NOT1 (N311, N298);
and AND2 (N312, N308, N50);
nand NAND2 (N313, N307, N16);
buf BUF1 (N314, N313);
nor NOR4 (N315, N283, N121, N286, N304);
and AND4 (N316, N24, N110, N46, N46);
and AND2 (N317, N310, N294);
xor XOR2 (N318, N290, N163);
nand NAND2 (N319, N317, N202);
nand NAND2 (N320, N306, N151);
or OR2 (N321, N311, N192);
and AND3 (N322, N314, N45, N308);
not NOT1 (N323, N312);
nor NOR4 (N324, N315, N154, N239, N290);
xor XOR2 (N325, N322, N79);
nor NOR2 (N326, N291, N50);
or OR3 (N327, N316, N88, N1);
xor XOR2 (N328, N299, N6);
and AND3 (N329, N324, N172, N293);
and AND4 (N330, N318, N93, N277, N275);
nand NAND4 (N331, N321, N233, N39, N81);
or OR2 (N332, N330, N102);
or OR4 (N333, N328, N331, N71, N121);
buf BUF1 (N334, N322);
xor XOR2 (N335, N319, N66);
nor NOR2 (N336, N334, N70);
buf BUF1 (N337, N333);
xor XOR2 (N338, N327, N114);
and AND4 (N339, N332, N230, N34, N266);
xor XOR2 (N340, N325, N11);
and AND4 (N341, N329, N262, N10, N241);
and AND2 (N342, N339, N293);
not NOT1 (N343, N320);
nand NAND3 (N344, N341, N288, N282);
xor XOR2 (N345, N340, N281);
and AND4 (N346, N337, N343, N314, N93);
nand NAND2 (N347, N311, N231);
nand NAND3 (N348, N323, N274, N236);
xor XOR2 (N349, N336, N163);
or OR3 (N350, N349, N124, N228);
nand NAND2 (N351, N326, N8);
buf BUF1 (N352, N345);
xor XOR2 (N353, N335, N302);
xor XOR2 (N354, N342, N182);
xor XOR2 (N355, N352, N295);
or OR4 (N356, N344, N277, N296, N74);
nor NOR4 (N357, N348, N154, N71, N83);
xor XOR2 (N358, N356, N221);
nand NAND4 (N359, N338, N68, N93, N297);
nor NOR2 (N360, N350, N246);
nand NAND4 (N361, N347, N187, N214, N251);
and AND2 (N362, N358, N177);
nand NAND4 (N363, N357, N349, N252, N40);
xor XOR2 (N364, N351, N167);
buf BUF1 (N365, N359);
or OR2 (N366, N353, N237);
or OR2 (N367, N366, N20);
and AND3 (N368, N346, N20, N175);
and AND4 (N369, N368, N305, N142, N20);
or OR2 (N370, N354, N68);
nor NOR4 (N371, N360, N301, N104, N115);
xor XOR2 (N372, N355, N272);
xor XOR2 (N373, N362, N134);
nand NAND3 (N374, N370, N372, N171);
buf BUF1 (N375, N306);
nor NOR2 (N376, N375, N121);
nand NAND3 (N377, N363, N351, N302);
buf BUF1 (N378, N361);
and AND3 (N379, N376, N142, N179);
not NOT1 (N380, N374);
not NOT1 (N381, N373);
xor XOR2 (N382, N378, N118);
and AND3 (N383, N377, N348, N121);
nand NAND2 (N384, N367, N239);
xor XOR2 (N385, N380, N80);
nor NOR3 (N386, N383, N17, N209);
nor NOR3 (N387, N386, N371, N87);
not NOT1 (N388, N266);
and AND2 (N389, N387, N65);
and AND4 (N390, N388, N381, N168, N13);
xor XOR2 (N391, N233, N2);
not NOT1 (N392, N389);
or OR3 (N393, N384, N33, N84);
not NOT1 (N394, N385);
nand NAND2 (N395, N392, N341);
nor NOR4 (N396, N382, N59, N395, N249);
nor NOR3 (N397, N356, N110, N332);
nand NAND4 (N398, N379, N167, N239, N126);
and AND4 (N399, N390, N337, N264, N46);
not NOT1 (N400, N391);
nor NOR4 (N401, N393, N126, N305, N250);
buf BUF1 (N402, N396);
and AND3 (N403, N399, N63, N395);
not NOT1 (N404, N369);
buf BUF1 (N405, N400);
buf BUF1 (N406, N364);
or OR3 (N407, N398, N207, N176);
not NOT1 (N408, N403);
nor NOR4 (N409, N394, N59, N183, N152);
xor XOR2 (N410, N409, N264);
or OR4 (N411, N408, N37, N405, N109);
not NOT1 (N412, N183);
and AND4 (N413, N412, N302, N9, N8);
not NOT1 (N414, N413);
nand NAND4 (N415, N407, N251, N295, N168);
not NOT1 (N416, N401);
and AND4 (N417, N411, N377, N304, N214);
buf BUF1 (N418, N402);
and AND3 (N419, N397, N244, N357);
or OR4 (N420, N417, N32, N121, N27);
nand NAND2 (N421, N415, N143);
nor NOR3 (N422, N421, N404, N51);
buf BUF1 (N423, N63);
or OR2 (N424, N410, N85);
nand NAND4 (N425, N422, N207, N239, N159);
and AND4 (N426, N420, N278, N15, N54);
xor XOR2 (N427, N419, N362);
nand NAND4 (N428, N427, N120, N33, N346);
nand NAND2 (N429, N424, N146);
xor XOR2 (N430, N406, N160);
xor XOR2 (N431, N425, N256);
xor XOR2 (N432, N426, N241);
xor XOR2 (N433, N423, N34);
nor NOR3 (N434, N430, N255, N180);
not NOT1 (N435, N428);
buf BUF1 (N436, N414);
nand NAND3 (N437, N429, N387, N375);
nand NAND3 (N438, N435, N257, N412);
not NOT1 (N439, N438);
nor NOR2 (N440, N431, N71);
nor NOR3 (N441, N432, N74, N202);
and AND4 (N442, N437, N24, N73, N273);
and AND3 (N443, N436, N384, N80);
buf BUF1 (N444, N418);
and AND4 (N445, N440, N400, N261, N176);
or OR4 (N446, N434, N29, N191, N310);
buf BUF1 (N447, N444);
not NOT1 (N448, N439);
buf BUF1 (N449, N448);
nand NAND2 (N450, N446, N295);
nand NAND3 (N451, N450, N58, N267);
nor NOR3 (N452, N442, N86, N202);
or OR3 (N453, N433, N84, N323);
nor NOR2 (N454, N365, N284);
xor XOR2 (N455, N449, N262);
nor NOR2 (N456, N447, N169);
or OR4 (N457, N443, N334, N75, N205);
or OR4 (N458, N457, N212, N79, N79);
and AND3 (N459, N451, N302, N52);
not NOT1 (N460, N453);
xor XOR2 (N461, N445, N125);
buf BUF1 (N462, N454);
not NOT1 (N463, N452);
and AND2 (N464, N416, N430);
buf BUF1 (N465, N464);
nor NOR2 (N466, N456, N250);
or OR2 (N467, N459, N187);
not NOT1 (N468, N466);
xor XOR2 (N469, N460, N201);
not NOT1 (N470, N458);
not NOT1 (N471, N463);
or OR4 (N472, N468, N108, N183, N402);
not NOT1 (N473, N441);
and AND4 (N474, N472, N380, N186, N330);
not NOT1 (N475, N474);
or OR4 (N476, N475, N306, N461, N67);
or OR2 (N477, N32, N148);
xor XOR2 (N478, N471, N342);
nand NAND4 (N479, N473, N129, N121, N242);
or OR2 (N480, N470, N134);
or OR4 (N481, N455, N356, N476, N288);
or OR4 (N482, N194, N306, N445, N336);
xor XOR2 (N483, N467, N104);
buf BUF1 (N484, N477);
not NOT1 (N485, N484);
or OR3 (N486, N478, N338, N6);
nand NAND2 (N487, N483, N50);
buf BUF1 (N488, N481);
nand NAND4 (N489, N487, N235, N450, N197);
nand NAND2 (N490, N485, N481);
nand NAND2 (N491, N490, N179);
not NOT1 (N492, N491);
buf BUF1 (N493, N488);
nand NAND3 (N494, N492, N220, N172);
nor NOR3 (N495, N479, N60, N404);
xor XOR2 (N496, N480, N237);
nor NOR4 (N497, N493, N325, N409, N493);
nand NAND4 (N498, N462, N377, N398, N25);
buf BUF1 (N499, N497);
and AND3 (N500, N494, N142, N447);
nor NOR2 (N501, N499, N473);
not NOT1 (N502, N486);
nor NOR3 (N503, N465, N307, N152);
buf BUF1 (N504, N503);
not NOT1 (N505, N495);
nor NOR2 (N506, N496, N282);
not NOT1 (N507, N482);
not NOT1 (N508, N506);
xor XOR2 (N509, N504, N369);
nor NOR4 (N510, N502, N352, N203, N480);
nand NAND3 (N511, N500, N441, N433);
nand NAND2 (N512, N508, N25);
nor NOR2 (N513, N511, N75);
and AND4 (N514, N509, N502, N214, N23);
or OR4 (N515, N514, N32, N205, N423);
nor NOR4 (N516, N505, N418, N269, N501);
and AND4 (N517, N83, N423, N26, N457);
nor NOR3 (N518, N513, N62, N413);
nand NAND2 (N519, N512, N383);
nand NAND4 (N520, N469, N329, N355, N244);
buf BUF1 (N521, N498);
xor XOR2 (N522, N515, N298);
not NOT1 (N523, N521);
nand NAND2 (N524, N520, N119);
and AND3 (N525, N489, N192, N471);
buf BUF1 (N526, N518);
nand NAND4 (N527, N525, N378, N68, N321);
nor NOR2 (N528, N527, N253);
nor NOR3 (N529, N519, N456, N513);
buf BUF1 (N530, N528);
xor XOR2 (N531, N517, N368);
nor NOR2 (N532, N523, N496);
nand NAND4 (N533, N532, N424, N492, N143);
nor NOR2 (N534, N522, N501);
xor XOR2 (N535, N507, N160);
and AND4 (N536, N533, N414, N138, N519);
xor XOR2 (N537, N526, N492);
xor XOR2 (N538, N531, N317);
or OR3 (N539, N529, N368, N373);
and AND4 (N540, N510, N113, N110, N56);
buf BUF1 (N541, N535);
xor XOR2 (N542, N516, N265);
or OR4 (N543, N541, N171, N441, N467);
nand NAND3 (N544, N538, N375, N471);
nand NAND3 (N545, N544, N137, N389);
and AND4 (N546, N545, N72, N180, N336);
and AND3 (N547, N543, N162, N427);
and AND3 (N548, N540, N445, N512);
and AND4 (N549, N542, N360, N415, N362);
nand NAND3 (N550, N536, N405, N70);
or OR2 (N551, N550, N125);
not NOT1 (N552, N524);
buf BUF1 (N553, N548);
nand NAND4 (N554, N551, N284, N169, N341);
nor NOR4 (N555, N547, N66, N495, N410);
buf BUF1 (N556, N546);
buf BUF1 (N557, N553);
xor XOR2 (N558, N534, N543);
nand NAND2 (N559, N549, N368);
xor XOR2 (N560, N552, N129);
nand NAND3 (N561, N558, N73, N299);
or OR4 (N562, N559, N206, N61, N218);
and AND4 (N563, N537, N470, N248, N550);
nor NOR4 (N564, N560, N451, N533, N465);
nand NAND2 (N565, N564, N207);
or OR2 (N566, N556, N333);
xor XOR2 (N567, N530, N152);
nor NOR4 (N568, N554, N281, N277, N66);
buf BUF1 (N569, N555);
not NOT1 (N570, N566);
xor XOR2 (N571, N557, N461);
nand NAND4 (N572, N562, N20, N71, N412);
nand NAND3 (N573, N565, N357, N301);
xor XOR2 (N574, N567, N222);
nand NAND3 (N575, N574, N314, N187);
and AND2 (N576, N539, N324);
not NOT1 (N577, N570);
nand NAND3 (N578, N563, N165, N472);
or OR2 (N579, N561, N455);
not NOT1 (N580, N576);
or OR3 (N581, N572, N505, N276);
nor NOR4 (N582, N580, N454, N83, N316);
xor XOR2 (N583, N577, N319);
xor XOR2 (N584, N569, N68);
and AND3 (N585, N571, N253, N568);
xor XOR2 (N586, N577, N212);
nor NOR2 (N587, N586, N182);
nand NAND2 (N588, N582, N140);
buf BUF1 (N589, N585);
or OR2 (N590, N578, N339);
xor XOR2 (N591, N573, N286);
xor XOR2 (N592, N587, N533);
nor NOR4 (N593, N579, N361, N44, N523);
nor NOR4 (N594, N583, N114, N362, N153);
and AND4 (N595, N590, N305, N410, N258);
buf BUF1 (N596, N594);
or OR3 (N597, N588, N425, N417);
and AND3 (N598, N595, N141, N106);
nor NOR4 (N599, N597, N591, N211, N5);
not NOT1 (N600, N129);
nand NAND4 (N601, N589, N222, N512, N590);
or OR2 (N602, N599, N433);
not NOT1 (N603, N598);
nand NAND4 (N604, N592, N131, N583, N462);
and AND2 (N605, N575, N275);
nor NOR4 (N606, N600, N155, N600, N77);
xor XOR2 (N607, N584, N104);
xor XOR2 (N608, N606, N171);
nand NAND3 (N609, N605, N344, N172);
nand NAND4 (N610, N602, N65, N341, N366);
or OR4 (N611, N596, N434, N92, N495);
buf BUF1 (N612, N593);
xor XOR2 (N613, N610, N530);
nand NAND3 (N614, N581, N193, N313);
buf BUF1 (N615, N601);
nand NAND3 (N616, N609, N5, N491);
nand NAND3 (N617, N613, N522, N526);
buf BUF1 (N618, N603);
nand NAND3 (N619, N612, N568, N217);
and AND2 (N620, N615, N205);
nor NOR2 (N621, N607, N409);
or OR3 (N622, N619, N446, N104);
xor XOR2 (N623, N614, N60);
nor NOR3 (N624, N608, N591, N529);
or OR3 (N625, N616, N442, N483);
and AND4 (N626, N604, N67, N447, N78);
xor XOR2 (N627, N626, N3);
nand NAND2 (N628, N623, N224);
nand NAND4 (N629, N620, N282, N452, N104);
or OR2 (N630, N618, N335);
or OR3 (N631, N630, N271, N403);
and AND2 (N632, N625, N57);
buf BUF1 (N633, N632);
or OR2 (N634, N631, N376);
and AND2 (N635, N617, N316);
buf BUF1 (N636, N621);
not NOT1 (N637, N634);
buf BUF1 (N638, N637);
xor XOR2 (N639, N629, N54);
nor NOR4 (N640, N638, N448, N409, N518);
buf BUF1 (N641, N628);
or OR4 (N642, N635, N90, N196, N577);
and AND2 (N643, N627, N352);
nand NAND4 (N644, N640, N466, N281, N488);
buf BUF1 (N645, N642);
nand NAND4 (N646, N633, N216, N432, N465);
buf BUF1 (N647, N645);
nand NAND4 (N648, N639, N578, N258, N472);
not NOT1 (N649, N644);
nand NAND4 (N650, N624, N202, N505, N299);
nand NAND2 (N651, N641, N51);
xor XOR2 (N652, N648, N588);
or OR3 (N653, N649, N144, N237);
buf BUF1 (N654, N611);
nor NOR3 (N655, N652, N462, N400);
or OR3 (N656, N650, N524, N545);
not NOT1 (N657, N656);
nand NAND2 (N658, N653, N80);
buf BUF1 (N659, N651);
xor XOR2 (N660, N658, N348);
or OR4 (N661, N647, N443, N483, N263);
nand NAND2 (N662, N636, N579);
or OR4 (N663, N657, N433, N497, N311);
or OR3 (N664, N622, N3, N79);
xor XOR2 (N665, N643, N609);
and AND4 (N666, N664, N620, N538, N215);
or OR3 (N667, N659, N515, N180);
or OR4 (N668, N663, N76, N429, N168);
nand NAND4 (N669, N655, N286, N377, N413);
not NOT1 (N670, N668);
not NOT1 (N671, N661);
buf BUF1 (N672, N671);
nor NOR2 (N673, N654, N289);
and AND4 (N674, N660, N362, N55, N158);
xor XOR2 (N675, N674, N277);
and AND3 (N676, N662, N317, N521);
or OR2 (N677, N675, N220);
not NOT1 (N678, N667);
and AND4 (N679, N672, N528, N267, N562);
nand NAND3 (N680, N676, N106, N418);
and AND4 (N681, N670, N58, N188, N398);
buf BUF1 (N682, N677);
xor XOR2 (N683, N682, N52);
buf BUF1 (N684, N681);
nor NOR2 (N685, N665, N82);
xor XOR2 (N686, N685, N599);
xor XOR2 (N687, N678, N388);
nor NOR2 (N688, N680, N449);
nor NOR2 (N689, N686, N378);
nor NOR3 (N690, N689, N131, N30);
not NOT1 (N691, N646);
nand NAND2 (N692, N679, N78);
nand NAND4 (N693, N669, N463, N443, N20);
buf BUF1 (N694, N692);
or OR4 (N695, N694, N374, N504, N651);
or OR3 (N696, N695, N318, N392);
or OR3 (N697, N666, N48, N106);
nand NAND4 (N698, N688, N263, N406, N553);
not NOT1 (N699, N696);
not NOT1 (N700, N673);
nand NAND4 (N701, N683, N169, N687, N41);
buf BUF1 (N702, N665);
not NOT1 (N703, N684);
not NOT1 (N704, N698);
nand NAND2 (N705, N697, N118);
buf BUF1 (N706, N705);
not NOT1 (N707, N701);
or OR2 (N708, N693, N460);
or OR3 (N709, N708, N524, N213);
nor NOR3 (N710, N700, N583, N250);
nor NOR2 (N711, N709, N560);
xor XOR2 (N712, N691, N8);
or OR2 (N713, N690, N347);
nor NOR4 (N714, N712, N564, N329, N381);
or OR2 (N715, N703, N513);
and AND2 (N716, N699, N294);
nand NAND2 (N717, N714, N352);
buf BUF1 (N718, N707);
or OR3 (N719, N717, N389, N698);
buf BUF1 (N720, N710);
or OR2 (N721, N720, N492);
buf BUF1 (N722, N716);
and AND3 (N723, N711, N277, N34);
nor NOR3 (N724, N718, N651, N427);
nand NAND4 (N725, N722, N720, N451, N398);
or OR4 (N726, N706, N230, N583, N123);
and AND4 (N727, N702, N184, N70, N374);
and AND2 (N728, N723, N722);
xor XOR2 (N729, N715, N63);
buf BUF1 (N730, N721);
xor XOR2 (N731, N704, N522);
or OR4 (N732, N725, N544, N319, N548);
buf BUF1 (N733, N727);
nand NAND3 (N734, N713, N174, N345);
not NOT1 (N735, N731);
xor XOR2 (N736, N734, N509);
or OR2 (N737, N726, N127);
xor XOR2 (N738, N733, N560);
xor XOR2 (N739, N719, N331);
nor NOR3 (N740, N730, N643, N177);
xor XOR2 (N741, N729, N381);
xor XOR2 (N742, N737, N170);
buf BUF1 (N743, N732);
not NOT1 (N744, N738);
xor XOR2 (N745, N744, N573);
and AND2 (N746, N735, N43);
nor NOR3 (N747, N746, N39, N593);
not NOT1 (N748, N739);
not NOT1 (N749, N740);
not NOT1 (N750, N745);
not NOT1 (N751, N736);
and AND4 (N752, N741, N741, N143, N388);
or OR2 (N753, N748, N372);
nand NAND2 (N754, N743, N183);
not NOT1 (N755, N742);
not NOT1 (N756, N753);
buf BUF1 (N757, N749);
nand NAND2 (N758, N724, N135);
or OR2 (N759, N747, N162);
nor NOR3 (N760, N759, N453, N752);
nand NAND2 (N761, N78, N488);
buf BUF1 (N762, N758);
buf BUF1 (N763, N754);
not NOT1 (N764, N750);
nor NOR3 (N765, N763, N90, N568);
and AND3 (N766, N757, N30, N360);
nor NOR2 (N767, N755, N134);
buf BUF1 (N768, N761);
buf BUF1 (N769, N751);
buf BUF1 (N770, N766);
nand NAND4 (N771, N762, N99, N696, N196);
or OR4 (N772, N728, N534, N542, N364);
nand NAND3 (N773, N760, N640, N5);
nor NOR3 (N774, N771, N552, N474);
not NOT1 (N775, N772);
nand NAND2 (N776, N773, N740);
xor XOR2 (N777, N770, N21);
or OR4 (N778, N776, N551, N481, N685);
and AND2 (N779, N765, N723);
and AND3 (N780, N768, N183, N543);
xor XOR2 (N781, N756, N222);
nor NOR4 (N782, N777, N476, N400, N319);
nor NOR3 (N783, N775, N185, N3);
nor NOR3 (N784, N774, N586, N480);
nand NAND4 (N785, N767, N42, N312, N713);
xor XOR2 (N786, N784, N225);
or OR2 (N787, N782, N691);
xor XOR2 (N788, N778, N585);
xor XOR2 (N789, N786, N781);
buf BUF1 (N790, N485);
nor NOR3 (N791, N790, N238, N10);
nand NAND3 (N792, N780, N562, N573);
nand NAND3 (N793, N791, N427, N717);
nor NOR4 (N794, N787, N50, N316, N617);
or OR4 (N795, N788, N430, N403, N83);
nor NOR4 (N796, N792, N119, N67, N668);
buf BUF1 (N797, N783);
not NOT1 (N798, N796);
nand NAND2 (N799, N789, N666);
or OR2 (N800, N798, N90);
or OR2 (N801, N779, N351);
nor NOR4 (N802, N769, N672, N775, N582);
xor XOR2 (N803, N802, N167);
or OR4 (N804, N795, N64, N535, N456);
buf BUF1 (N805, N794);
or OR2 (N806, N785, N40);
xor XOR2 (N807, N799, N199);
nor NOR3 (N808, N804, N298, N771);
or OR4 (N809, N803, N674, N408, N200);
xor XOR2 (N810, N793, N774);
buf BUF1 (N811, N800);
buf BUF1 (N812, N808);
nor NOR3 (N813, N810, N698, N564);
nor NOR4 (N814, N801, N398, N526, N561);
nand NAND3 (N815, N809, N614, N550);
nand NAND2 (N816, N812, N466);
xor XOR2 (N817, N797, N672);
not NOT1 (N818, N815);
buf BUF1 (N819, N816);
xor XOR2 (N820, N807, N134);
nor NOR4 (N821, N764, N790, N184, N539);
or OR3 (N822, N817, N562, N291);
nor NOR3 (N823, N813, N631, N691);
nor NOR3 (N824, N821, N556, N52);
nand NAND4 (N825, N811, N352, N576, N710);
and AND2 (N826, N806, N101);
xor XOR2 (N827, N824, N491);
xor XOR2 (N828, N826, N827);
xor XOR2 (N829, N158, N498);
not NOT1 (N830, N814);
nand NAND2 (N831, N820, N698);
xor XOR2 (N832, N818, N752);
nor NOR2 (N833, N825, N318);
and AND3 (N834, N823, N526, N51);
nor NOR2 (N835, N833, N681);
buf BUF1 (N836, N831);
nand NAND2 (N837, N832, N338);
nor NOR2 (N838, N834, N755);
nand NAND3 (N839, N805, N525, N85);
xor XOR2 (N840, N830, N119);
and AND3 (N841, N837, N797, N450);
nor NOR4 (N842, N819, N376, N669, N613);
buf BUF1 (N843, N838);
nor NOR4 (N844, N843, N362, N29, N209);
buf BUF1 (N845, N836);
nor NOR2 (N846, N828, N351);
nor NOR2 (N847, N829, N513);
and AND4 (N848, N835, N830, N76, N235);
not NOT1 (N849, N844);
nor NOR3 (N850, N846, N380, N751);
not NOT1 (N851, N847);
xor XOR2 (N852, N839, N157);
nor NOR2 (N853, N851, N781);
or OR2 (N854, N852, N756);
nor NOR2 (N855, N822, N774);
not NOT1 (N856, N854);
and AND3 (N857, N856, N475, N750);
or OR3 (N858, N848, N778, N741);
nand NAND3 (N859, N853, N160, N463);
xor XOR2 (N860, N850, N180);
buf BUF1 (N861, N860);
nor NOR3 (N862, N858, N252, N678);
or OR3 (N863, N845, N588, N762);
buf BUF1 (N864, N849);
or OR2 (N865, N840, N625);
xor XOR2 (N866, N864, N468);
nor NOR4 (N867, N865, N633, N188, N428);
xor XOR2 (N868, N862, N860);
and AND3 (N869, N857, N245, N107);
not NOT1 (N870, N859);
buf BUF1 (N871, N868);
nand NAND4 (N872, N867, N258, N166, N46);
nor NOR2 (N873, N870, N659);
nor NOR3 (N874, N873, N126, N667);
and AND2 (N875, N866, N723);
xor XOR2 (N876, N874, N596);
or OR3 (N877, N872, N747, N271);
nand NAND2 (N878, N841, N594);
nand NAND4 (N879, N869, N131, N29, N298);
or OR2 (N880, N855, N633);
nand NAND4 (N881, N877, N448, N121, N229);
nor NOR2 (N882, N879, N250);
and AND3 (N883, N880, N839, N287);
not NOT1 (N884, N875);
nand NAND4 (N885, N878, N114, N309, N760);
not NOT1 (N886, N881);
or OR3 (N887, N884, N494, N422);
nor NOR2 (N888, N882, N437);
not NOT1 (N889, N888);
xor XOR2 (N890, N885, N810);
not NOT1 (N891, N876);
and AND4 (N892, N889, N617, N247, N257);
nand NAND4 (N893, N892, N368, N530, N314);
buf BUF1 (N894, N842);
and AND4 (N895, N891, N787, N429, N425);
buf BUF1 (N896, N895);
xor XOR2 (N897, N861, N563);
nand NAND3 (N898, N871, N864, N176);
nor NOR2 (N899, N886, N698);
not NOT1 (N900, N897);
nor NOR4 (N901, N883, N877, N817, N575);
nand NAND2 (N902, N896, N145);
nor NOR4 (N903, N887, N628, N42, N85);
nand NAND3 (N904, N901, N667, N181);
nor NOR2 (N905, N898, N353);
buf BUF1 (N906, N903);
nor NOR4 (N907, N902, N140, N348, N286);
not NOT1 (N908, N907);
nor NOR4 (N909, N904, N376, N378, N546);
xor XOR2 (N910, N909, N284);
not NOT1 (N911, N863);
xor XOR2 (N912, N905, N28);
nor NOR4 (N913, N911, N597, N668, N285);
nand NAND4 (N914, N913, N213, N694, N281);
nor NOR2 (N915, N893, N360);
or OR3 (N916, N914, N465, N256);
xor XOR2 (N917, N890, N675);
buf BUF1 (N918, N894);
not NOT1 (N919, N912);
xor XOR2 (N920, N908, N657);
xor XOR2 (N921, N916, N358);
nand NAND4 (N922, N918, N715, N252, N811);
nand NAND4 (N923, N899, N277, N221, N7);
nor NOR3 (N924, N906, N418, N41);
not NOT1 (N925, N922);
nor NOR2 (N926, N900, N179);
buf BUF1 (N927, N924);
or OR4 (N928, N927, N309, N927, N144);
xor XOR2 (N929, N919, N370);
nand NAND2 (N930, N928, N532);
and AND2 (N931, N929, N788);
or OR4 (N932, N917, N269, N132, N693);
or OR3 (N933, N915, N37, N754);
xor XOR2 (N934, N920, N575);
buf BUF1 (N935, N925);
xor XOR2 (N936, N933, N500);
or OR4 (N937, N926, N558, N216, N620);
and AND4 (N938, N923, N610, N321, N167);
not NOT1 (N939, N921);
or OR2 (N940, N910, N374);
not NOT1 (N941, N937);
and AND2 (N942, N939, N135);
nand NAND4 (N943, N930, N832, N455, N152);
buf BUF1 (N944, N934);
not NOT1 (N945, N944);
xor XOR2 (N946, N936, N586);
or OR3 (N947, N938, N18, N330);
not NOT1 (N948, N943);
nand NAND2 (N949, N947, N469);
xor XOR2 (N950, N940, N104);
not NOT1 (N951, N946);
buf BUF1 (N952, N951);
xor XOR2 (N953, N945, N675);
nor NOR2 (N954, N949, N38);
xor XOR2 (N955, N952, N372);
and AND2 (N956, N932, N499);
xor XOR2 (N957, N931, N595);
nor NOR3 (N958, N935, N934, N747);
and AND3 (N959, N954, N154, N506);
nor NOR2 (N960, N958, N766);
nor NOR2 (N961, N955, N285);
not NOT1 (N962, N950);
and AND4 (N963, N957, N957, N571, N62);
or OR2 (N964, N963, N926);
not NOT1 (N965, N942);
or OR4 (N966, N962, N699, N9, N492);
not NOT1 (N967, N948);
not NOT1 (N968, N966);
or OR4 (N969, N967, N123, N802, N843);
or OR2 (N970, N968, N384);
nand NAND3 (N971, N956, N195, N747);
nand NAND3 (N972, N971, N633, N617);
buf BUF1 (N973, N941);
nand NAND2 (N974, N972, N366);
nand NAND3 (N975, N969, N307, N374);
buf BUF1 (N976, N973);
not NOT1 (N977, N953);
nand NAND2 (N978, N976, N916);
xor XOR2 (N979, N975, N846);
nand NAND4 (N980, N959, N233, N216, N180);
not NOT1 (N981, N978);
buf BUF1 (N982, N970);
or OR2 (N983, N977, N596);
nand NAND4 (N984, N982, N616, N340, N518);
xor XOR2 (N985, N979, N512);
not NOT1 (N986, N984);
not NOT1 (N987, N965);
xor XOR2 (N988, N981, N405);
and AND2 (N989, N960, N252);
or OR4 (N990, N987, N85, N522, N831);
or OR3 (N991, N961, N778, N51);
buf BUF1 (N992, N991);
nand NAND3 (N993, N986, N660, N363);
buf BUF1 (N994, N974);
or OR3 (N995, N994, N944, N527);
xor XOR2 (N996, N985, N331);
nor NOR3 (N997, N988, N396, N217);
buf BUF1 (N998, N992);
and AND2 (N999, N993, N771);
nand NAND3 (N1000, N983, N532, N407);
xor XOR2 (N1001, N990, N683);
xor XOR2 (N1002, N1001, N810);
nor NOR3 (N1003, N995, N162, N467);
nor NOR3 (N1004, N997, N777, N279);
nor NOR2 (N1005, N1002, N455);
nor NOR3 (N1006, N989, N474, N402);
or OR3 (N1007, N980, N612, N115);
buf BUF1 (N1008, N964);
nor NOR2 (N1009, N999, N895);
or OR3 (N1010, N1007, N225, N335);
buf BUF1 (N1011, N1004);
nand NAND2 (N1012, N1006, N884);
xor XOR2 (N1013, N1011, N765);
xor XOR2 (N1014, N1013, N960);
xor XOR2 (N1015, N1003, N780);
buf BUF1 (N1016, N1008);
nand NAND2 (N1017, N1009, N528);
not NOT1 (N1018, N996);
nand NAND3 (N1019, N1016, N576, N805);
buf BUF1 (N1020, N1005);
or OR2 (N1021, N1012, N898);
not NOT1 (N1022, N1018);
and AND4 (N1023, N1021, N48, N202, N602);
not NOT1 (N1024, N1010);
xor XOR2 (N1025, N1015, N62);
and AND4 (N1026, N1017, N709, N410, N743);
xor XOR2 (N1027, N1000, N134);
not NOT1 (N1028, N1027);
nand NAND2 (N1029, N1024, N980);
or OR4 (N1030, N1025, N886, N796, N842);
not NOT1 (N1031, N1019);
buf BUF1 (N1032, N998);
buf BUF1 (N1033, N1023);
xor XOR2 (N1034, N1028, N377);
nor NOR3 (N1035, N1033, N1004, N866);
buf BUF1 (N1036, N1032);
and AND3 (N1037, N1026, N1027, N157);
not NOT1 (N1038, N1034);
buf BUF1 (N1039, N1031);
or OR3 (N1040, N1029, N22, N533);
nor NOR4 (N1041, N1037, N874, N703, N361);
buf BUF1 (N1042, N1040);
or OR3 (N1043, N1041, N623, N271);
not NOT1 (N1044, N1014);
buf BUF1 (N1045, N1044);
not NOT1 (N1046, N1036);
nand NAND2 (N1047, N1039, N897);
nand NAND2 (N1048, N1042, N953);
and AND4 (N1049, N1048, N173, N685, N357);
nor NOR3 (N1050, N1043, N853, N564);
or OR3 (N1051, N1030, N894, N941);
buf BUF1 (N1052, N1038);
and AND3 (N1053, N1050, N738, N603);
and AND2 (N1054, N1049, N92);
or OR4 (N1055, N1054, N84, N1048, N331);
xor XOR2 (N1056, N1045, N248);
or OR3 (N1057, N1052, N450, N129);
buf BUF1 (N1058, N1056);
buf BUF1 (N1059, N1055);
nand NAND4 (N1060, N1059, N333, N142, N643);
and AND4 (N1061, N1060, N759, N271, N111);
and AND2 (N1062, N1020, N1012);
nand NAND4 (N1063, N1061, N699, N269, N515);
not NOT1 (N1064, N1047);
nand NAND3 (N1065, N1058, N967, N966);
and AND2 (N1066, N1064, N504);
buf BUF1 (N1067, N1053);
nor NOR4 (N1068, N1051, N143, N839, N24);
not NOT1 (N1069, N1063);
or OR3 (N1070, N1068, N348, N467);
buf BUF1 (N1071, N1022);
buf BUF1 (N1072, N1065);
buf BUF1 (N1073, N1072);
nor NOR2 (N1074, N1069, N145);
not NOT1 (N1075, N1070);
or OR4 (N1076, N1035, N835, N896, N742);
buf BUF1 (N1077, N1076);
xor XOR2 (N1078, N1046, N795);
not NOT1 (N1079, N1074);
and AND2 (N1080, N1057, N953);
and AND3 (N1081, N1075, N607, N223);
nand NAND2 (N1082, N1062, N491);
and AND4 (N1083, N1066, N328, N865, N822);
xor XOR2 (N1084, N1083, N808);
buf BUF1 (N1085, N1078);
and AND4 (N1086, N1081, N614, N692, N535);
and AND4 (N1087, N1085, N2, N229, N101);
buf BUF1 (N1088, N1079);
buf BUF1 (N1089, N1071);
buf BUF1 (N1090, N1080);
and AND2 (N1091, N1084, N1071);
or OR4 (N1092, N1087, N290, N904, N378);
or OR3 (N1093, N1091, N88, N728);
buf BUF1 (N1094, N1093);
buf BUF1 (N1095, N1073);
and AND3 (N1096, N1089, N61, N1013);
or OR4 (N1097, N1094, N807, N1039, N898);
nand NAND4 (N1098, N1077, N234, N338, N160);
buf BUF1 (N1099, N1086);
nand NAND2 (N1100, N1098, N673);
nand NAND4 (N1101, N1088, N939, N609, N256);
xor XOR2 (N1102, N1099, N415);
not NOT1 (N1103, N1097);
buf BUF1 (N1104, N1100);
xor XOR2 (N1105, N1104, N1039);
nor NOR4 (N1106, N1092, N534, N308, N1042);
or OR3 (N1107, N1103, N665, N294);
xor XOR2 (N1108, N1105, N783);
buf BUF1 (N1109, N1090);
xor XOR2 (N1110, N1107, N27);
or OR4 (N1111, N1082, N948, N579, N95);
nor NOR3 (N1112, N1101, N468, N180);
buf BUF1 (N1113, N1095);
nor NOR2 (N1114, N1108, N1065);
or OR3 (N1115, N1067, N622, N292);
or OR2 (N1116, N1096, N152);
nor NOR3 (N1117, N1109, N50, N415);
not NOT1 (N1118, N1116);
and AND3 (N1119, N1118, N203, N632);
nor NOR3 (N1120, N1110, N634, N139);
buf BUF1 (N1121, N1106);
and AND3 (N1122, N1114, N1072, N1115);
and AND3 (N1123, N629, N416, N214);
not NOT1 (N1124, N1121);
nand NAND3 (N1125, N1102, N303, N1102);
or OR3 (N1126, N1111, N1026, N785);
or OR3 (N1127, N1123, N600, N876);
and AND3 (N1128, N1113, N471, N424);
nand NAND2 (N1129, N1124, N893);
buf BUF1 (N1130, N1119);
xor XOR2 (N1131, N1125, N58);
and AND3 (N1132, N1122, N145, N900);
not NOT1 (N1133, N1112);
not NOT1 (N1134, N1130);
or OR4 (N1135, N1120, N739, N189, N185);
and AND4 (N1136, N1129, N755, N567, N404);
or OR2 (N1137, N1128, N806);
nand NAND4 (N1138, N1126, N1046, N1111, N826);
buf BUF1 (N1139, N1138);
or OR4 (N1140, N1137, N541, N828, N1099);
nor NOR4 (N1141, N1132, N156, N830, N404);
and AND3 (N1142, N1141, N291, N1070);
nand NAND2 (N1143, N1131, N64);
xor XOR2 (N1144, N1117, N701);
xor XOR2 (N1145, N1136, N723);
xor XOR2 (N1146, N1127, N258);
xor XOR2 (N1147, N1144, N1041);
buf BUF1 (N1148, N1135);
not NOT1 (N1149, N1147);
not NOT1 (N1150, N1133);
buf BUF1 (N1151, N1142);
nor NOR2 (N1152, N1145, N819);
nor NOR2 (N1153, N1152, N1130);
not NOT1 (N1154, N1151);
not NOT1 (N1155, N1134);
buf BUF1 (N1156, N1148);
xor XOR2 (N1157, N1140, N247);
nor NOR2 (N1158, N1139, N1049);
buf BUF1 (N1159, N1157);
buf BUF1 (N1160, N1154);
not NOT1 (N1161, N1150);
not NOT1 (N1162, N1143);
xor XOR2 (N1163, N1159, N174);
buf BUF1 (N1164, N1162);
nand NAND2 (N1165, N1161, N132);
not NOT1 (N1166, N1146);
or OR3 (N1167, N1158, N423, N150);
xor XOR2 (N1168, N1164, N1029);
nor NOR4 (N1169, N1167, N957, N896, N425);
nor NOR3 (N1170, N1160, N567, N1103);
not NOT1 (N1171, N1153);
or OR4 (N1172, N1169, N912, N605, N106);
buf BUF1 (N1173, N1168);
nor NOR3 (N1174, N1166, N912, N356);
buf BUF1 (N1175, N1149);
xor XOR2 (N1176, N1163, N922);
or OR2 (N1177, N1172, N589);
xor XOR2 (N1178, N1170, N426);
not NOT1 (N1179, N1176);
buf BUF1 (N1180, N1156);
buf BUF1 (N1181, N1177);
nand NAND4 (N1182, N1180, N151, N421, N588);
buf BUF1 (N1183, N1181);
nor NOR4 (N1184, N1165, N1152, N481, N306);
xor XOR2 (N1185, N1173, N573);
xor XOR2 (N1186, N1179, N1052);
nand NAND4 (N1187, N1184, N259, N254, N1163);
nand NAND3 (N1188, N1174, N1082, N108);
and AND2 (N1189, N1155, N837);
nand NAND3 (N1190, N1187, N255, N252);
not NOT1 (N1191, N1190);
xor XOR2 (N1192, N1182, N113);
nand NAND2 (N1193, N1185, N700);
nor NOR2 (N1194, N1188, N209);
nand NAND4 (N1195, N1193, N319, N105, N60);
xor XOR2 (N1196, N1175, N572);
or OR2 (N1197, N1192, N845);
buf BUF1 (N1198, N1183);
buf BUF1 (N1199, N1195);
or OR3 (N1200, N1178, N812, N846);
and AND3 (N1201, N1171, N1008, N587);
nor NOR2 (N1202, N1201, N674);
buf BUF1 (N1203, N1189);
and AND4 (N1204, N1203, N367, N1086, N720);
nand NAND3 (N1205, N1197, N44, N471);
nand NAND3 (N1206, N1199, N117, N222);
or OR4 (N1207, N1196, N254, N1123, N279);
nand NAND4 (N1208, N1204, N133, N5, N78);
nand NAND3 (N1209, N1198, N171, N949);
buf BUF1 (N1210, N1206);
or OR4 (N1211, N1191, N1028, N598, N150);
nand NAND4 (N1212, N1200, N21, N158, N172);
nand NAND2 (N1213, N1207, N71);
buf BUF1 (N1214, N1210);
xor XOR2 (N1215, N1213, N1144);
nand NAND2 (N1216, N1186, N644);
xor XOR2 (N1217, N1212, N775);
buf BUF1 (N1218, N1202);
and AND3 (N1219, N1214, N1008, N834);
and AND2 (N1220, N1211, N313);
or OR4 (N1221, N1219, N327, N62, N1080);
and AND4 (N1222, N1217, N701, N397, N831);
and AND4 (N1223, N1222, N460, N536, N775);
xor XOR2 (N1224, N1205, N485);
nand NAND4 (N1225, N1216, N1029, N858, N836);
nor NOR3 (N1226, N1209, N350, N272);
xor XOR2 (N1227, N1221, N1092);
nor NOR2 (N1228, N1218, N1197);
nand NAND4 (N1229, N1194, N748, N376, N1045);
not NOT1 (N1230, N1220);
nand NAND2 (N1231, N1227, N838);
nor NOR4 (N1232, N1228, N81, N122, N300);
or OR2 (N1233, N1229, N1031);
nor NOR3 (N1234, N1208, N777, N606);
xor XOR2 (N1235, N1225, N58);
nor NOR4 (N1236, N1232, N167, N700, N373);
or OR2 (N1237, N1236, N649);
or OR3 (N1238, N1234, N422, N411);
nand NAND2 (N1239, N1235, N46);
and AND4 (N1240, N1230, N39, N883, N49);
and AND2 (N1241, N1240, N119);
nor NOR4 (N1242, N1223, N447, N360, N945);
buf BUF1 (N1243, N1224);
xor XOR2 (N1244, N1239, N420);
xor XOR2 (N1245, N1226, N831);
or OR4 (N1246, N1243, N1215, N897, N1079);
nand NAND3 (N1247, N1222, N855, N193);
or OR2 (N1248, N1241, N203);
nor NOR3 (N1249, N1237, N9, N1144);
buf BUF1 (N1250, N1249);
not NOT1 (N1251, N1233);
not NOT1 (N1252, N1250);
nand NAND3 (N1253, N1248, N241, N249);
xor XOR2 (N1254, N1246, N434);
not NOT1 (N1255, N1244);
xor XOR2 (N1256, N1251, N884);
or OR4 (N1257, N1242, N999, N1142, N1004);
xor XOR2 (N1258, N1253, N1077);
and AND2 (N1259, N1255, N1062);
not NOT1 (N1260, N1257);
not NOT1 (N1261, N1256);
or OR3 (N1262, N1260, N517, N153);
or OR4 (N1263, N1254, N42, N237, N680);
or OR2 (N1264, N1261, N188);
xor XOR2 (N1265, N1262, N724);
nand NAND2 (N1266, N1247, N755);
and AND2 (N1267, N1238, N1097);
nand NAND2 (N1268, N1263, N100);
nand NAND2 (N1269, N1258, N1248);
or OR4 (N1270, N1267, N987, N1025, N389);
buf BUF1 (N1271, N1266);
xor XOR2 (N1272, N1231, N435);
xor XOR2 (N1273, N1259, N686);
not NOT1 (N1274, N1252);
nand NAND3 (N1275, N1271, N1073, N598);
or OR2 (N1276, N1273, N1204);
or OR4 (N1277, N1270, N61, N1152, N1025);
or OR2 (N1278, N1268, N1038);
nor NOR3 (N1279, N1278, N1164, N40);
nand NAND4 (N1280, N1277, N704, N547, N404);
xor XOR2 (N1281, N1276, N814);
nor NOR2 (N1282, N1280, N1078);
or OR2 (N1283, N1281, N992);
or OR4 (N1284, N1274, N1205, N567, N772);
nor NOR3 (N1285, N1283, N1242, N1257);
nor NOR4 (N1286, N1275, N195, N708, N713);
or OR3 (N1287, N1285, N1029, N521);
nand NAND2 (N1288, N1264, N777);
nand NAND2 (N1289, N1287, N740);
or OR4 (N1290, N1288, N830, N930, N293);
not NOT1 (N1291, N1265);
buf BUF1 (N1292, N1289);
or OR3 (N1293, N1290, N104, N748);
buf BUF1 (N1294, N1293);
xor XOR2 (N1295, N1272, N573);
nand NAND4 (N1296, N1282, N935, N637, N917);
nand NAND2 (N1297, N1291, N1292);
nor NOR3 (N1298, N1185, N932, N505);
and AND2 (N1299, N1286, N1037);
buf BUF1 (N1300, N1295);
nand NAND4 (N1301, N1284, N1279, N495, N775);
not NOT1 (N1302, N767);
xor XOR2 (N1303, N1297, N657);
and AND2 (N1304, N1296, N155);
not NOT1 (N1305, N1302);
and AND3 (N1306, N1305, N1029, N408);
nand NAND2 (N1307, N1298, N384);
not NOT1 (N1308, N1269);
nor NOR4 (N1309, N1303, N1149, N1034, N659);
or OR4 (N1310, N1245, N114, N386, N934);
nand NAND4 (N1311, N1301, N275, N306, N102);
nor NOR4 (N1312, N1306, N1073, N540, N791);
xor XOR2 (N1313, N1309, N867);
xor XOR2 (N1314, N1310, N898);
nor NOR2 (N1315, N1304, N1263);
buf BUF1 (N1316, N1294);
xor XOR2 (N1317, N1314, N365);
nor NOR2 (N1318, N1308, N1163);
xor XOR2 (N1319, N1315, N583);
and AND3 (N1320, N1313, N822, N677);
xor XOR2 (N1321, N1299, N468);
not NOT1 (N1322, N1317);
nand NAND4 (N1323, N1318, N216, N562, N1132);
and AND2 (N1324, N1300, N1237);
or OR2 (N1325, N1307, N643);
and AND3 (N1326, N1325, N265, N434);
not NOT1 (N1327, N1319);
nor NOR2 (N1328, N1321, N1081);
nor NOR3 (N1329, N1327, N438, N40);
xor XOR2 (N1330, N1316, N246);
nor NOR4 (N1331, N1328, N1000, N360, N848);
and AND4 (N1332, N1312, N634, N47, N675);
not NOT1 (N1333, N1322);
nand NAND2 (N1334, N1329, N1044);
nand NAND3 (N1335, N1331, N611, N47);
and AND3 (N1336, N1330, N601, N329);
xor XOR2 (N1337, N1311, N937);
or OR4 (N1338, N1332, N298, N357, N608);
buf BUF1 (N1339, N1333);
buf BUF1 (N1340, N1336);
buf BUF1 (N1341, N1340);
and AND3 (N1342, N1341, N945, N1090);
nand NAND3 (N1343, N1342, N1316, N583);
and AND2 (N1344, N1324, N160);
and AND2 (N1345, N1334, N564);
xor XOR2 (N1346, N1337, N510);
not NOT1 (N1347, N1339);
nand NAND2 (N1348, N1343, N148);
xor XOR2 (N1349, N1348, N841);
not NOT1 (N1350, N1349);
buf BUF1 (N1351, N1344);
xor XOR2 (N1352, N1347, N581);
nor NOR2 (N1353, N1351, N1015);
xor XOR2 (N1354, N1346, N830);
or OR4 (N1355, N1354, N1243, N9, N59);
or OR2 (N1356, N1326, N31);
nor NOR3 (N1357, N1352, N163, N389);
buf BUF1 (N1358, N1323);
not NOT1 (N1359, N1353);
and AND4 (N1360, N1338, N782, N495, N1132);
nand NAND2 (N1361, N1356, N1042);
buf BUF1 (N1362, N1355);
and AND4 (N1363, N1320, N261, N1327, N639);
and AND4 (N1364, N1363, N436, N1194, N953);
buf BUF1 (N1365, N1362);
buf BUF1 (N1366, N1361);
not NOT1 (N1367, N1364);
and AND2 (N1368, N1366, N802);
nand NAND3 (N1369, N1345, N401, N690);
nor NOR4 (N1370, N1367, N500, N389, N918);
not NOT1 (N1371, N1357);
not NOT1 (N1372, N1335);
not NOT1 (N1373, N1372);
not NOT1 (N1374, N1365);
not NOT1 (N1375, N1358);
not NOT1 (N1376, N1370);
and AND4 (N1377, N1373, N950, N1019, N634);
and AND3 (N1378, N1368, N410, N847);
buf BUF1 (N1379, N1359);
xor XOR2 (N1380, N1374, N437);
and AND3 (N1381, N1369, N236, N353);
buf BUF1 (N1382, N1360);
buf BUF1 (N1383, N1350);
xor XOR2 (N1384, N1380, N453);
or OR3 (N1385, N1381, N1276, N1298);
nand NAND3 (N1386, N1385, N283, N1284);
or OR2 (N1387, N1376, N660);
xor XOR2 (N1388, N1384, N74);
and AND2 (N1389, N1375, N803);
xor XOR2 (N1390, N1387, N420);
or OR3 (N1391, N1378, N1330, N1368);
nor NOR3 (N1392, N1379, N134, N584);
nor NOR2 (N1393, N1382, N102);
not NOT1 (N1394, N1371);
nand NAND3 (N1395, N1389, N214, N1004);
nand NAND4 (N1396, N1386, N1389, N313, N413);
nor NOR2 (N1397, N1396, N565);
and AND4 (N1398, N1397, N1154, N1281, N843);
and AND4 (N1399, N1394, N1367, N746, N152);
nand NAND3 (N1400, N1398, N639, N1360);
xor XOR2 (N1401, N1383, N835);
nand NAND2 (N1402, N1399, N9);
xor XOR2 (N1403, N1390, N68);
and AND4 (N1404, N1401, N919, N234, N122);
xor XOR2 (N1405, N1393, N1303);
xor XOR2 (N1406, N1388, N936);
nand NAND2 (N1407, N1403, N301);
not NOT1 (N1408, N1405);
and AND4 (N1409, N1392, N237, N762, N1096);
and AND4 (N1410, N1391, N11, N735, N521);
buf BUF1 (N1411, N1408);
or OR2 (N1412, N1400, N1398);
or OR4 (N1413, N1395, N698, N1312, N345);
and AND4 (N1414, N1377, N801, N592, N89);
or OR3 (N1415, N1404, N34, N744);
and AND2 (N1416, N1407, N1169);
buf BUF1 (N1417, N1415);
not NOT1 (N1418, N1411);
or OR4 (N1419, N1412, N776, N470, N185);
not NOT1 (N1420, N1414);
xor XOR2 (N1421, N1409, N656);
and AND2 (N1422, N1419, N54);
xor XOR2 (N1423, N1413, N648);
not NOT1 (N1424, N1402);
nor NOR2 (N1425, N1420, N1156);
nor NOR2 (N1426, N1410, N269);
and AND3 (N1427, N1424, N507, N164);
nor NOR2 (N1428, N1416, N108);
nor NOR3 (N1429, N1426, N1007, N573);
not NOT1 (N1430, N1422);
and AND2 (N1431, N1418, N974);
not NOT1 (N1432, N1421);
or OR3 (N1433, N1425, N786, N1073);
xor XOR2 (N1434, N1406, N737);
buf BUF1 (N1435, N1431);
xor XOR2 (N1436, N1435, N60);
and AND4 (N1437, N1417, N870, N1089, N414);
buf BUF1 (N1438, N1427);
nand NAND2 (N1439, N1430, N962);
and AND4 (N1440, N1434, N396, N893, N1041);
nand NAND4 (N1441, N1437, N300, N1021, N1116);
or OR4 (N1442, N1440, N1347, N1111, N587);
buf BUF1 (N1443, N1428);
or OR4 (N1444, N1443, N301, N1436, N931);
nor NOR4 (N1445, N439, N334, N1005, N50);
or OR3 (N1446, N1445, N1249, N598);
buf BUF1 (N1447, N1441);
buf BUF1 (N1448, N1439);
and AND2 (N1449, N1429, N1322);
nor NOR4 (N1450, N1432, N912, N324, N1327);
or OR3 (N1451, N1442, N17, N1151);
nand NAND4 (N1452, N1433, N1019, N1060, N829);
buf BUF1 (N1453, N1448);
buf BUF1 (N1454, N1447);
nand NAND2 (N1455, N1453, N818);
not NOT1 (N1456, N1444);
nand NAND2 (N1457, N1451, N1157);
not NOT1 (N1458, N1454);
or OR2 (N1459, N1438, N1415);
and AND3 (N1460, N1458, N838, N581);
and AND2 (N1461, N1460, N637);
buf BUF1 (N1462, N1449);
xor XOR2 (N1463, N1457, N126);
buf BUF1 (N1464, N1456);
or OR4 (N1465, N1423, N755, N1056, N575);
and AND4 (N1466, N1461, N33, N598, N1410);
nand NAND4 (N1467, N1455, N402, N806, N513);
or OR4 (N1468, N1450, N512, N790, N990);
and AND4 (N1469, N1467, N1210, N418, N143);
buf BUF1 (N1470, N1446);
nor NOR2 (N1471, N1465, N217);
nand NAND2 (N1472, N1466, N1351);
nand NAND4 (N1473, N1462, N730, N223, N1440);
not NOT1 (N1474, N1468);
buf BUF1 (N1475, N1464);
nand NAND4 (N1476, N1463, N1137, N1164, N1416);
xor XOR2 (N1477, N1452, N1265);
xor XOR2 (N1478, N1474, N1100);
nor NOR2 (N1479, N1469, N1162);
nor NOR2 (N1480, N1478, N724);
buf BUF1 (N1481, N1475);
or OR2 (N1482, N1470, N474);
or OR2 (N1483, N1479, N856);
nand NAND3 (N1484, N1471, N342, N797);
xor XOR2 (N1485, N1484, N1017);
buf BUF1 (N1486, N1477);
nor NOR3 (N1487, N1472, N288, N966);
not NOT1 (N1488, N1473);
xor XOR2 (N1489, N1482, N1240);
xor XOR2 (N1490, N1489, N871);
xor XOR2 (N1491, N1486, N633);
buf BUF1 (N1492, N1476);
nor NOR2 (N1493, N1490, N527);
nand NAND2 (N1494, N1487, N1392);
buf BUF1 (N1495, N1481);
nand NAND2 (N1496, N1493, N206);
or OR3 (N1497, N1491, N177, N807);
buf BUF1 (N1498, N1495);
or OR3 (N1499, N1480, N1178, N902);
buf BUF1 (N1500, N1497);
or OR3 (N1501, N1494, N1222, N124);
xor XOR2 (N1502, N1488, N1497);
xor XOR2 (N1503, N1459, N138);
and AND4 (N1504, N1492, N280, N1195, N730);
buf BUF1 (N1505, N1501);
xor XOR2 (N1506, N1505, N40);
nor NOR4 (N1507, N1498, N327, N1159, N690);
not NOT1 (N1508, N1502);
and AND4 (N1509, N1507, N458, N792, N587);
buf BUF1 (N1510, N1509);
or OR2 (N1511, N1485, N506);
and AND3 (N1512, N1496, N1477, N440);
and AND4 (N1513, N1508, N604, N385, N960);
nand NAND2 (N1514, N1512, N848);
nor NOR3 (N1515, N1506, N452, N283);
nor NOR3 (N1516, N1503, N1088, N787);
not NOT1 (N1517, N1483);
nor NOR4 (N1518, N1516, N564, N1, N148);
nand NAND2 (N1519, N1500, N48);
nand NAND4 (N1520, N1513, N609, N244, N252);
nand NAND3 (N1521, N1511, N110, N1170);
not NOT1 (N1522, N1515);
not NOT1 (N1523, N1519);
xor XOR2 (N1524, N1514, N1153);
buf BUF1 (N1525, N1499);
and AND3 (N1526, N1522, N430, N670);
or OR2 (N1527, N1520, N974);
nand NAND2 (N1528, N1527, N1107);
not NOT1 (N1529, N1523);
nor NOR2 (N1530, N1518, N1511);
or OR2 (N1531, N1526, N1400);
nor NOR4 (N1532, N1531, N1435, N13, N1096);
nor NOR3 (N1533, N1525, N377, N690);
and AND4 (N1534, N1532, N607, N923, N1064);
xor XOR2 (N1535, N1510, N201);
not NOT1 (N1536, N1530);
buf BUF1 (N1537, N1504);
nand NAND3 (N1538, N1533, N271, N221);
and AND4 (N1539, N1529, N857, N830, N1195);
or OR3 (N1540, N1536, N1323, N690);
nor NOR3 (N1541, N1540, N1040, N621);
not NOT1 (N1542, N1521);
buf BUF1 (N1543, N1538);
not NOT1 (N1544, N1534);
nand NAND2 (N1545, N1528, N1339);
or OR3 (N1546, N1535, N124, N1143);
buf BUF1 (N1547, N1517);
not NOT1 (N1548, N1539);
nand NAND4 (N1549, N1545, N1485, N1041, N1462);
and AND4 (N1550, N1549, N1513, N77, N61);
nor NOR2 (N1551, N1524, N866);
nor NOR4 (N1552, N1551, N1302, N899, N185);
xor XOR2 (N1553, N1537, N582);
xor XOR2 (N1554, N1546, N713);
and AND4 (N1555, N1542, N1126, N161, N12);
not NOT1 (N1556, N1555);
or OR2 (N1557, N1547, N401);
xor XOR2 (N1558, N1543, N1092);
not NOT1 (N1559, N1544);
nand NAND3 (N1560, N1552, N1203, N26);
buf BUF1 (N1561, N1550);
nand NAND4 (N1562, N1548, N713, N1007, N11);
buf BUF1 (N1563, N1554);
not NOT1 (N1564, N1541);
buf BUF1 (N1565, N1561);
nand NAND3 (N1566, N1557, N1039, N680);
xor XOR2 (N1567, N1559, N928);
nand NAND4 (N1568, N1567, N1262, N305, N862);
nand NAND3 (N1569, N1565, N234, N1101);
nand NAND4 (N1570, N1562, N1208, N1477, N110);
xor XOR2 (N1571, N1563, N1006);
not NOT1 (N1572, N1558);
buf BUF1 (N1573, N1553);
nand NAND2 (N1574, N1573, N214);
not NOT1 (N1575, N1564);
or OR4 (N1576, N1571, N169, N1377, N1408);
nor NOR3 (N1577, N1575, N1079, N693);
nor NOR2 (N1578, N1568, N866);
nor NOR2 (N1579, N1577, N717);
not NOT1 (N1580, N1560);
nor NOR2 (N1581, N1566, N1396);
not NOT1 (N1582, N1580);
xor XOR2 (N1583, N1569, N371);
buf BUF1 (N1584, N1576);
xor XOR2 (N1585, N1572, N657);
or OR3 (N1586, N1584, N591, N1113);
and AND4 (N1587, N1585, N758, N1330, N939);
not NOT1 (N1588, N1587);
buf BUF1 (N1589, N1588);
not NOT1 (N1590, N1556);
or OR2 (N1591, N1590, N456);
nor NOR2 (N1592, N1570, N1171);
xor XOR2 (N1593, N1583, N936);
buf BUF1 (N1594, N1591);
xor XOR2 (N1595, N1592, N34);
nand NAND4 (N1596, N1593, N481, N287, N1530);
buf BUF1 (N1597, N1596);
and AND3 (N1598, N1579, N971, N978);
nand NAND2 (N1599, N1574, N11);
and AND4 (N1600, N1597, N1121, N490, N1229);
and AND2 (N1601, N1598, N602);
nor NOR3 (N1602, N1600, N1533, N437);
nand NAND3 (N1603, N1594, N1268, N1279);
xor XOR2 (N1604, N1581, N451);
nand NAND4 (N1605, N1603, N266, N525, N1269);
buf BUF1 (N1606, N1595);
nand NAND4 (N1607, N1604, N1462, N522, N1176);
or OR4 (N1608, N1599, N1220, N22, N218);
or OR4 (N1609, N1601, N539, N268, N1540);
buf BUF1 (N1610, N1582);
or OR3 (N1611, N1606, N1272, N1457);
nor NOR2 (N1612, N1611, N480);
not NOT1 (N1613, N1586);
and AND3 (N1614, N1610, N761, N644);
nor NOR2 (N1615, N1602, N197);
buf BUF1 (N1616, N1613);
or OR3 (N1617, N1616, N1134, N1017);
nand NAND2 (N1618, N1617, N413);
xor XOR2 (N1619, N1605, N636);
nand NAND2 (N1620, N1615, N622);
not NOT1 (N1621, N1589);
and AND3 (N1622, N1620, N341, N170);
xor XOR2 (N1623, N1607, N964);
nor NOR4 (N1624, N1621, N990, N592, N1147);
nor NOR3 (N1625, N1578, N990, N980);
nor NOR2 (N1626, N1609, N199);
or OR4 (N1627, N1626, N1557, N1073, N1574);
buf BUF1 (N1628, N1622);
buf BUF1 (N1629, N1624);
buf BUF1 (N1630, N1629);
nor NOR3 (N1631, N1614, N36, N1357);
or OR4 (N1632, N1608, N661, N868, N1219);
nand NAND2 (N1633, N1632, N403);
nand NAND3 (N1634, N1628, N908, N186);
not NOT1 (N1635, N1630);
and AND4 (N1636, N1612, N102, N632, N144);
buf BUF1 (N1637, N1619);
buf BUF1 (N1638, N1618);
or OR3 (N1639, N1633, N1069, N1395);
not NOT1 (N1640, N1636);
buf BUF1 (N1641, N1627);
nor NOR3 (N1642, N1639, N1369, N684);
nor NOR3 (N1643, N1641, N316, N703);
not NOT1 (N1644, N1623);
not NOT1 (N1645, N1643);
not NOT1 (N1646, N1637);
xor XOR2 (N1647, N1645, N244);
xor XOR2 (N1648, N1638, N629);
buf BUF1 (N1649, N1631);
buf BUF1 (N1650, N1648);
xor XOR2 (N1651, N1635, N211);
xor XOR2 (N1652, N1642, N1308);
and AND4 (N1653, N1646, N891, N870, N802);
nand NAND2 (N1654, N1644, N633);
and AND4 (N1655, N1653, N734, N1200, N1506);
buf BUF1 (N1656, N1649);
nand NAND3 (N1657, N1625, N1375, N1484);
buf BUF1 (N1658, N1652);
nand NAND3 (N1659, N1656, N1358, N579);
buf BUF1 (N1660, N1654);
and AND4 (N1661, N1657, N993, N1474, N1386);
or OR2 (N1662, N1650, N1256);
xor XOR2 (N1663, N1659, N782);
and AND2 (N1664, N1662, N1451);
not NOT1 (N1665, N1658);
nand NAND2 (N1666, N1660, N1606);
and AND3 (N1667, N1665, N693, N120);
or OR4 (N1668, N1661, N593, N1405, N1451);
or OR3 (N1669, N1647, N32, N21);
nand NAND2 (N1670, N1668, N905);
or OR2 (N1671, N1651, N564);
nor NOR2 (N1672, N1671, N1019);
not NOT1 (N1673, N1663);
buf BUF1 (N1674, N1664);
nor NOR4 (N1675, N1670, N621, N1579, N68);
buf BUF1 (N1676, N1669);
buf BUF1 (N1677, N1675);
buf BUF1 (N1678, N1666);
nand NAND3 (N1679, N1676, N230, N67);
not NOT1 (N1680, N1672);
not NOT1 (N1681, N1634);
buf BUF1 (N1682, N1679);
nor NOR3 (N1683, N1655, N873, N1079);
nand NAND3 (N1684, N1677, N375, N145);
nand NAND4 (N1685, N1682, N402, N1327, N986);
buf BUF1 (N1686, N1684);
not NOT1 (N1687, N1681);
and AND3 (N1688, N1673, N766, N234);
nand NAND3 (N1689, N1687, N1501, N937);
nand NAND4 (N1690, N1674, N1450, N685, N1245);
not NOT1 (N1691, N1686);
nor NOR2 (N1692, N1683, N402);
buf BUF1 (N1693, N1692);
buf BUF1 (N1694, N1667);
and AND3 (N1695, N1691, N1096, N908);
nor NOR4 (N1696, N1678, N897, N407, N1671);
xor XOR2 (N1697, N1690, N822);
and AND4 (N1698, N1689, N1536, N377, N999);
nand NAND4 (N1699, N1696, N502, N318, N295);
not NOT1 (N1700, N1688);
buf BUF1 (N1701, N1685);
nor NOR2 (N1702, N1698, N586);
buf BUF1 (N1703, N1640);
and AND3 (N1704, N1699, N493, N703);
nor NOR3 (N1705, N1680, N64, N619);
xor XOR2 (N1706, N1697, N1619);
xor XOR2 (N1707, N1693, N558);
buf BUF1 (N1708, N1700);
buf BUF1 (N1709, N1694);
and AND3 (N1710, N1695, N960, N1547);
not NOT1 (N1711, N1702);
buf BUF1 (N1712, N1707);
xor XOR2 (N1713, N1711, N672);
buf BUF1 (N1714, N1705);
and AND3 (N1715, N1712, N954, N1278);
or OR3 (N1716, N1715, N420, N528);
nor NOR2 (N1717, N1716, N1078);
buf BUF1 (N1718, N1709);
xor XOR2 (N1719, N1701, N48);
or OR2 (N1720, N1719, N289);
and AND4 (N1721, N1720, N672, N921, N956);
buf BUF1 (N1722, N1721);
nor NOR4 (N1723, N1714, N1292, N1529, N741);
xor XOR2 (N1724, N1704, N1449);
and AND4 (N1725, N1724, N244, N813, N11);
nand NAND2 (N1726, N1706, N422);
buf BUF1 (N1727, N1718);
nor NOR3 (N1728, N1710, N280, N929);
not NOT1 (N1729, N1703);
nand NAND3 (N1730, N1728, N620, N91);
or OR4 (N1731, N1729, N1635, N26, N202);
not NOT1 (N1732, N1725);
xor XOR2 (N1733, N1730, N1005);
not NOT1 (N1734, N1727);
nand NAND3 (N1735, N1732, N528, N1042);
or OR3 (N1736, N1717, N1444, N1397);
buf BUF1 (N1737, N1722);
nand NAND4 (N1738, N1734, N1670, N1130, N1687);
xor XOR2 (N1739, N1737, N1281);
not NOT1 (N1740, N1713);
nand NAND2 (N1741, N1726, N1417);
xor XOR2 (N1742, N1738, N1329);
not NOT1 (N1743, N1723);
and AND2 (N1744, N1742, N516);
and AND3 (N1745, N1736, N266, N1269);
not NOT1 (N1746, N1740);
not NOT1 (N1747, N1733);
not NOT1 (N1748, N1744);
and AND3 (N1749, N1741, N335, N61);
xor XOR2 (N1750, N1731, N171);
not NOT1 (N1751, N1748);
and AND4 (N1752, N1746, N76, N1050, N305);
nor NOR4 (N1753, N1745, N536, N906, N1193);
xor XOR2 (N1754, N1752, N1118);
or OR2 (N1755, N1754, N906);
or OR2 (N1756, N1753, N663);
xor XOR2 (N1757, N1756, N391);
xor XOR2 (N1758, N1755, N1693);
buf BUF1 (N1759, N1747);
or OR3 (N1760, N1749, N1258, N595);
nand NAND3 (N1761, N1739, N333, N553);
not NOT1 (N1762, N1760);
or OR2 (N1763, N1761, N1067);
not NOT1 (N1764, N1762);
nor NOR3 (N1765, N1759, N590, N752);
not NOT1 (N1766, N1751);
and AND3 (N1767, N1757, N994, N1690);
and AND2 (N1768, N1765, N623);
not NOT1 (N1769, N1758);
buf BUF1 (N1770, N1769);
xor XOR2 (N1771, N1766, N1326);
or OR3 (N1772, N1764, N870, N1308);
not NOT1 (N1773, N1763);
or OR3 (N1774, N1767, N860, N1532);
not NOT1 (N1775, N1772);
or OR2 (N1776, N1743, N1593);
or OR2 (N1777, N1708, N1485);
not NOT1 (N1778, N1750);
xor XOR2 (N1779, N1777, N861);
buf BUF1 (N1780, N1771);
or OR3 (N1781, N1735, N808, N1086);
buf BUF1 (N1782, N1781);
and AND4 (N1783, N1774, N131, N694, N1111);
nand NAND4 (N1784, N1782, N59, N1528, N641);
not NOT1 (N1785, N1773);
xor XOR2 (N1786, N1780, N942);
nor NOR3 (N1787, N1776, N103, N861);
not NOT1 (N1788, N1784);
nor NOR3 (N1789, N1787, N416, N1640);
not NOT1 (N1790, N1785);
xor XOR2 (N1791, N1790, N521);
or OR2 (N1792, N1778, N510);
nand NAND3 (N1793, N1775, N539, N1731);
nor NOR4 (N1794, N1783, N1527, N775, N1530);
nor NOR2 (N1795, N1779, N25);
or OR4 (N1796, N1788, N1401, N2, N377);
not NOT1 (N1797, N1794);
nor NOR2 (N1798, N1795, N907);
nand NAND2 (N1799, N1793, N620);
nor NOR2 (N1800, N1791, N776);
buf BUF1 (N1801, N1800);
or OR3 (N1802, N1792, N1601, N786);
not NOT1 (N1803, N1770);
and AND2 (N1804, N1802, N328);
and AND2 (N1805, N1789, N1078);
buf BUF1 (N1806, N1768);
and AND4 (N1807, N1803, N1373, N1627, N810);
nor NOR4 (N1808, N1807, N874, N926, N100);
xor XOR2 (N1809, N1804, N412);
not NOT1 (N1810, N1786);
and AND4 (N1811, N1798, N1163, N285, N1261);
nor NOR2 (N1812, N1801, N195);
buf BUF1 (N1813, N1811);
xor XOR2 (N1814, N1797, N1284);
nor NOR3 (N1815, N1796, N161, N963);
nand NAND3 (N1816, N1814, N269, N1304);
buf BUF1 (N1817, N1805);
and AND2 (N1818, N1815, N1520);
nor NOR3 (N1819, N1808, N669, N91);
nand NAND3 (N1820, N1809, N496, N802);
xor XOR2 (N1821, N1816, N1155);
xor XOR2 (N1822, N1812, N991);
and AND2 (N1823, N1820, N1135);
or OR3 (N1824, N1817, N1175, N1268);
xor XOR2 (N1825, N1822, N179);
xor XOR2 (N1826, N1799, N1457);
not NOT1 (N1827, N1819);
buf BUF1 (N1828, N1827);
nand NAND3 (N1829, N1810, N294, N338);
or OR3 (N1830, N1818, N1502, N1794);
nand NAND3 (N1831, N1823, N522, N952);
and AND2 (N1832, N1829, N210);
nand NAND2 (N1833, N1832, N539);
nor NOR3 (N1834, N1824, N249, N95);
nor NOR4 (N1835, N1834, N761, N30, N952);
and AND2 (N1836, N1813, N363);
nand NAND3 (N1837, N1830, N479, N1302);
or OR2 (N1838, N1836, N1448);
and AND3 (N1839, N1806, N493, N1427);
not NOT1 (N1840, N1826);
not NOT1 (N1841, N1825);
xor XOR2 (N1842, N1833, N1135);
buf BUF1 (N1843, N1837);
and AND4 (N1844, N1821, N424, N585, N350);
buf BUF1 (N1845, N1838);
nand NAND2 (N1846, N1843, N1016);
xor XOR2 (N1847, N1846, N1564);
or OR4 (N1848, N1841, N499, N724, N1572);
nor NOR3 (N1849, N1828, N1708, N167);
and AND2 (N1850, N1848, N1505);
nor NOR4 (N1851, N1847, N370, N1416, N1462);
nor NOR4 (N1852, N1839, N944, N641, N1061);
and AND3 (N1853, N1842, N105, N1009);
or OR2 (N1854, N1845, N1656);
buf BUF1 (N1855, N1852);
nor NOR2 (N1856, N1853, N1758);
buf BUF1 (N1857, N1840);
or OR2 (N1858, N1857, N1851);
buf BUF1 (N1859, N1180);
nor NOR4 (N1860, N1856, N347, N781, N1233);
buf BUF1 (N1861, N1844);
buf BUF1 (N1862, N1860);
xor XOR2 (N1863, N1850, N1395);
and AND3 (N1864, N1855, N320, N415);
xor XOR2 (N1865, N1831, N1235);
not NOT1 (N1866, N1865);
or OR2 (N1867, N1861, N1758);
buf BUF1 (N1868, N1867);
and AND4 (N1869, N1849, N1770, N926, N36);
nor NOR2 (N1870, N1866, N199);
nand NAND4 (N1871, N1870, N1070, N593, N1853);
xor XOR2 (N1872, N1869, N1638);
nand NAND2 (N1873, N1862, N1837);
nand NAND3 (N1874, N1858, N1757, N622);
not NOT1 (N1875, N1835);
not NOT1 (N1876, N1859);
and AND3 (N1877, N1873, N180, N447);
or OR2 (N1878, N1864, N537);
nor NOR3 (N1879, N1874, N1827, N725);
nor NOR3 (N1880, N1871, N219, N95);
not NOT1 (N1881, N1880);
nor NOR3 (N1882, N1881, N1705, N131);
xor XOR2 (N1883, N1863, N1465);
nand NAND2 (N1884, N1882, N355);
xor XOR2 (N1885, N1875, N657);
and AND2 (N1886, N1885, N1655);
or OR2 (N1887, N1883, N418);
or OR4 (N1888, N1854, N1574, N907, N1811);
buf BUF1 (N1889, N1879);
xor XOR2 (N1890, N1872, N984);
nor NOR2 (N1891, N1889, N389);
nor NOR4 (N1892, N1878, N1811, N1835, N1456);
xor XOR2 (N1893, N1876, N794);
nor NOR3 (N1894, N1884, N1421, N1424);
buf BUF1 (N1895, N1893);
not NOT1 (N1896, N1887);
xor XOR2 (N1897, N1892, N721);
and AND4 (N1898, N1868, N179, N298, N303);
or OR2 (N1899, N1897, N782);
and AND2 (N1900, N1886, N1804);
xor XOR2 (N1901, N1895, N928);
xor XOR2 (N1902, N1899, N786);
buf BUF1 (N1903, N1890);
or OR2 (N1904, N1898, N874);
xor XOR2 (N1905, N1896, N1596);
or OR3 (N1906, N1901, N591, N937);
xor XOR2 (N1907, N1894, N1892);
xor XOR2 (N1908, N1900, N1850);
nor NOR4 (N1909, N1907, N810, N1131, N1442);
nand NAND4 (N1910, N1903, N479, N1566, N466);
or OR4 (N1911, N1888, N268, N495, N977);
buf BUF1 (N1912, N1911);
or OR2 (N1913, N1910, N1531);
or OR2 (N1914, N1909, N1705);
buf BUF1 (N1915, N1913);
nand NAND2 (N1916, N1902, N1828);
not NOT1 (N1917, N1916);
or OR4 (N1918, N1904, N1037, N1296, N455);
nor NOR4 (N1919, N1905, N979, N294, N72);
buf BUF1 (N1920, N1912);
nor NOR4 (N1921, N1906, N270, N1268, N872);
and AND2 (N1922, N1915, N859);
or OR4 (N1923, N1920, N1214, N609, N1211);
or OR3 (N1924, N1877, N179, N765);
buf BUF1 (N1925, N1924);
buf BUF1 (N1926, N1922);
xor XOR2 (N1927, N1917, N787);
not NOT1 (N1928, N1921);
and AND2 (N1929, N1914, N554);
buf BUF1 (N1930, N1923);
nor NOR4 (N1931, N1928, N154, N1170, N1315);
or OR2 (N1932, N1929, N1134);
and AND2 (N1933, N1930, N317);
nor NOR4 (N1934, N1933, N1180, N1196, N906);
nand NAND3 (N1935, N1891, N1862, N786);
or OR4 (N1936, N1908, N1564, N36, N422);
or OR4 (N1937, N1932, N979, N1479, N366);
buf BUF1 (N1938, N1935);
xor XOR2 (N1939, N1925, N903);
nand NAND3 (N1940, N1927, N917, N1074);
or OR3 (N1941, N1919, N199, N1295);
not NOT1 (N1942, N1918);
xor XOR2 (N1943, N1934, N1002);
not NOT1 (N1944, N1936);
not NOT1 (N1945, N1942);
nor NOR3 (N1946, N1938, N459, N406);
xor XOR2 (N1947, N1926, N670);
or OR4 (N1948, N1944, N1089, N1859, N148);
xor XOR2 (N1949, N1939, N310);
buf BUF1 (N1950, N1937);
or OR2 (N1951, N1946, N703);
nand NAND2 (N1952, N1947, N651);
nand NAND2 (N1953, N1945, N75);
and AND4 (N1954, N1943, N1796, N1796, N161);
nor NOR2 (N1955, N1941, N569);
not NOT1 (N1956, N1931);
and AND3 (N1957, N1948, N1669, N158);
nor NOR2 (N1958, N1953, N1269);
nand NAND4 (N1959, N1952, N777, N1461, N1882);
buf BUF1 (N1960, N1958);
xor XOR2 (N1961, N1960, N1704);
xor XOR2 (N1962, N1950, N1312);
not NOT1 (N1963, N1951);
not NOT1 (N1964, N1959);
and AND3 (N1965, N1961, N724, N131);
nor NOR2 (N1966, N1955, N742);
and AND2 (N1967, N1956, N1086);
and AND3 (N1968, N1949, N24, N1785);
nor NOR4 (N1969, N1954, N1614, N510, N1387);
or OR3 (N1970, N1968, N76, N918);
not NOT1 (N1971, N1964);
or OR4 (N1972, N1966, N836, N758, N830);
nor NOR4 (N1973, N1965, N869, N291, N174);
not NOT1 (N1974, N1957);
nor NOR2 (N1975, N1969, N732);
buf BUF1 (N1976, N1963);
buf BUF1 (N1977, N1962);
not NOT1 (N1978, N1973);
not NOT1 (N1979, N1977);
buf BUF1 (N1980, N1975);
xor XOR2 (N1981, N1974, N1526);
buf BUF1 (N1982, N1970);
or OR2 (N1983, N1972, N1804);
nor NOR3 (N1984, N1983, N1354, N1542);
buf BUF1 (N1985, N1984);
or OR2 (N1986, N1940, N347);
and AND4 (N1987, N1979, N1361, N702, N1638);
nor NOR2 (N1988, N1981, N32);
not NOT1 (N1989, N1986);
not NOT1 (N1990, N1989);
buf BUF1 (N1991, N1987);
xor XOR2 (N1992, N1988, N850);
nand NAND4 (N1993, N1990, N633, N1218, N1979);
not NOT1 (N1994, N1982);
buf BUF1 (N1995, N1976);
and AND3 (N1996, N1971, N189, N61);
and AND4 (N1997, N1995, N1362, N97, N645);
xor XOR2 (N1998, N1985, N504);
not NOT1 (N1999, N1992);
nand NAND3 (N2000, N1993, N665, N286);
nand NAND2 (N2001, N1978, N286);
or OR4 (N2002, N1997, N1814, N1230, N1855);
nand NAND4 (N2003, N1994, N536, N395, N154);
or OR3 (N2004, N1980, N1901, N1975);
nor NOR3 (N2005, N2003, N148, N827);
or OR3 (N2006, N1967, N1951, N1692);
or OR2 (N2007, N2004, N842);
nor NOR3 (N2008, N2005, N1831, N728);
nor NOR4 (N2009, N2000, N1861, N1665, N1832);
nor NOR2 (N2010, N2002, N676);
and AND3 (N2011, N1998, N1162, N78);
and AND4 (N2012, N2007, N345, N1652, N1249);
nor NOR2 (N2013, N2008, N1268);
or OR2 (N2014, N2009, N1376);
buf BUF1 (N2015, N2014);
nor NOR4 (N2016, N1999, N84, N132, N1619);
buf BUF1 (N2017, N2001);
nor NOR3 (N2018, N2012, N1437, N1020);
nor NOR4 (N2019, N1996, N1572, N300, N1541);
and AND4 (N2020, N1991, N713, N1050, N830);
nand NAND4 (N2021, N2016, N1385, N1874, N1813);
or OR2 (N2022, N2010, N541);
or OR3 (N2023, N2006, N1614, N306);
or OR3 (N2024, N2015, N388, N1008);
buf BUF1 (N2025, N2018);
xor XOR2 (N2026, N2011, N1705);
nand NAND4 (N2027, N2019, N190, N1609, N130);
nor NOR2 (N2028, N2017, N227);
nor NOR2 (N2029, N2020, N1864);
or OR3 (N2030, N2024, N1918, N1910);
and AND2 (N2031, N2025, N588);
or OR3 (N2032, N2031, N329, N100);
and AND4 (N2033, N2022, N1698, N1437, N1675);
nor NOR3 (N2034, N2023, N2033, N562);
not NOT1 (N2035, N1610);
nor NOR2 (N2036, N2013, N1681);
nor NOR4 (N2037, N2027, N1802, N1036, N751);
not NOT1 (N2038, N2037);
nor NOR2 (N2039, N2026, N579);
and AND4 (N2040, N2038, N1966, N1772, N463);
nor NOR4 (N2041, N2021, N1333, N324, N484);
not NOT1 (N2042, N2041);
or OR4 (N2043, N2035, N690, N1037, N857);
nand NAND4 (N2044, N2028, N1824, N1977, N118);
and AND2 (N2045, N2029, N1288);
not NOT1 (N2046, N2036);
xor XOR2 (N2047, N2030, N10);
nand NAND4 (N2048, N2034, N378, N1895, N2006);
or OR3 (N2049, N2039, N383, N687);
not NOT1 (N2050, N2043);
not NOT1 (N2051, N2046);
nor NOR2 (N2052, N2042, N127);
and AND4 (N2053, N2052, N1417, N965, N1409);
or OR3 (N2054, N2049, N1996, N477);
and AND2 (N2055, N2044, N1108);
and AND3 (N2056, N2040, N1411, N1604);
and AND2 (N2057, N2055, N1249);
not NOT1 (N2058, N2053);
xor XOR2 (N2059, N2045, N1207);
or OR4 (N2060, N2048, N178, N1996, N570);
or OR2 (N2061, N2058, N394);
nor NOR3 (N2062, N2056, N1924, N1727);
and AND3 (N2063, N2050, N1994, N410);
or OR2 (N2064, N2051, N662);
xor XOR2 (N2065, N2060, N222);
buf BUF1 (N2066, N2047);
xor XOR2 (N2067, N2059, N1459);
and AND3 (N2068, N2061, N1104, N3);
or OR3 (N2069, N2068, N863, N1439);
buf BUF1 (N2070, N2066);
or OR4 (N2071, N2069, N2005, N1076, N697);
or OR4 (N2072, N2054, N1633, N344, N982);
and AND3 (N2073, N2057, N1881, N2030);
or OR2 (N2074, N2064, N267);
xor XOR2 (N2075, N2071, N885);
buf BUF1 (N2076, N2062);
buf BUF1 (N2077, N2065);
nor NOR4 (N2078, N2077, N879, N376, N1038);
nand NAND3 (N2079, N2032, N1757, N1980);
not NOT1 (N2080, N2063);
xor XOR2 (N2081, N2070, N728);
nor NOR2 (N2082, N2072, N339);
nor NOR3 (N2083, N2080, N132, N166);
and AND4 (N2084, N2079, N740, N669, N1377);
nand NAND3 (N2085, N2082, N762, N100);
and AND3 (N2086, N2075, N1653, N1614);
or OR3 (N2087, N2085, N1113, N1043);
nand NAND3 (N2088, N2087, N1030, N1833);
xor XOR2 (N2089, N2076, N1037);
or OR4 (N2090, N2067, N64, N1205, N112);
nand NAND3 (N2091, N2073, N417, N1513);
not NOT1 (N2092, N2086);
and AND4 (N2093, N2078, N68, N946, N250);
buf BUF1 (N2094, N2092);
nor NOR2 (N2095, N2093, N934);
nand NAND4 (N2096, N2081, N1335, N744, N165);
nor NOR3 (N2097, N2095, N82, N27);
or OR3 (N2098, N2097, N1192, N640);
and AND2 (N2099, N2091, N1195);
or OR4 (N2100, N2074, N139, N1964, N732);
or OR4 (N2101, N2090, N1220, N982, N656);
buf BUF1 (N2102, N2098);
xor XOR2 (N2103, N2083, N2041);
buf BUF1 (N2104, N2089);
or OR4 (N2105, N2099, N153, N389, N1967);
not NOT1 (N2106, N2084);
or OR2 (N2107, N2106, N1505);
xor XOR2 (N2108, N2105, N463);
and AND2 (N2109, N2107, N514);
buf BUF1 (N2110, N2101);
xor XOR2 (N2111, N2100, N546);
nand NAND2 (N2112, N2109, N1105);
and AND4 (N2113, N2110, N50, N1929, N1106);
not NOT1 (N2114, N2111);
buf BUF1 (N2115, N2108);
nand NAND4 (N2116, N2094, N458, N1541, N1588);
xor XOR2 (N2117, N2096, N93);
buf BUF1 (N2118, N2114);
not NOT1 (N2119, N2116);
xor XOR2 (N2120, N2088, N1000);
xor XOR2 (N2121, N2103, N57);
nor NOR3 (N2122, N2115, N180, N1418);
and AND4 (N2123, N2113, N82, N1343, N1116);
buf BUF1 (N2124, N2123);
nand NAND4 (N2125, N2122, N498, N2060, N898);
xor XOR2 (N2126, N2117, N1656);
and AND4 (N2127, N2118, N1161, N1431, N757);
xor XOR2 (N2128, N2102, N814);
nor NOR3 (N2129, N2119, N288, N241);
not NOT1 (N2130, N2104);
buf BUF1 (N2131, N2126);
xor XOR2 (N2132, N2120, N37);
and AND4 (N2133, N2127, N1375, N1079, N1663);
buf BUF1 (N2134, N2133);
and AND2 (N2135, N2125, N1668);
nand NAND3 (N2136, N2131, N176, N685);
nor NOR3 (N2137, N2134, N413, N1807);
not NOT1 (N2138, N2124);
or OR2 (N2139, N2129, N327);
buf BUF1 (N2140, N2128);
or OR2 (N2141, N2136, N1800);
or OR2 (N2142, N2130, N1062);
xor XOR2 (N2143, N2142, N859);
not NOT1 (N2144, N2141);
or OR4 (N2145, N2144, N1987, N968, N2094);
xor XOR2 (N2146, N2135, N306);
nand NAND4 (N2147, N2132, N1640, N1760, N7);
nor NOR4 (N2148, N2147, N1488, N1199, N1543);
not NOT1 (N2149, N2121);
not NOT1 (N2150, N2148);
or OR4 (N2151, N2143, N1989, N1023, N1548);
not NOT1 (N2152, N2137);
nand NAND4 (N2153, N2140, N1126, N914, N492);
and AND2 (N2154, N2150, N1751);
and AND4 (N2155, N2145, N855, N1704, N511);
and AND4 (N2156, N2152, N508, N1265, N1449);
xor XOR2 (N2157, N2112, N1814);
xor XOR2 (N2158, N2156, N1257);
or OR2 (N2159, N2138, N1522);
or OR3 (N2160, N2146, N209, N1938);
nor NOR3 (N2161, N2153, N538, N159);
nand NAND2 (N2162, N2155, N2057);
buf BUF1 (N2163, N2157);
xor XOR2 (N2164, N2149, N830);
buf BUF1 (N2165, N2151);
nor NOR3 (N2166, N2161, N830, N1974);
buf BUF1 (N2167, N2158);
xor XOR2 (N2168, N2159, N1606);
nor NOR3 (N2169, N2154, N1045, N955);
buf BUF1 (N2170, N2162);
or OR3 (N2171, N2166, N2084, N2044);
not NOT1 (N2172, N2171);
xor XOR2 (N2173, N2160, N576);
not NOT1 (N2174, N2172);
or OR4 (N2175, N2139, N447, N138, N1454);
xor XOR2 (N2176, N2170, N658);
or OR4 (N2177, N2175, N1274, N465, N1877);
buf BUF1 (N2178, N2169);
and AND3 (N2179, N2173, N915, N1483);
or OR4 (N2180, N2164, N2122, N225, N2082);
or OR3 (N2181, N2167, N1794, N1558);
nand NAND4 (N2182, N2176, N1137, N1042, N281);
and AND2 (N2183, N2174, N1621);
buf BUF1 (N2184, N2180);
or OR2 (N2185, N2178, N837);
buf BUF1 (N2186, N2179);
buf BUF1 (N2187, N2181);
xor XOR2 (N2188, N2182, N874);
or OR2 (N2189, N2177, N1256);
buf BUF1 (N2190, N2186);
nor NOR3 (N2191, N2168, N1240, N1221);
xor XOR2 (N2192, N2187, N1162);
or OR2 (N2193, N2192, N185);
nand NAND4 (N2194, N2163, N1340, N1359, N420);
buf BUF1 (N2195, N2191);
xor XOR2 (N2196, N2185, N880);
or OR2 (N2197, N2188, N950);
buf BUF1 (N2198, N2197);
and AND2 (N2199, N2195, N944);
and AND2 (N2200, N2184, N528);
xor XOR2 (N2201, N2189, N1450);
not NOT1 (N2202, N2196);
not NOT1 (N2203, N2165);
nand NAND4 (N2204, N2198, N1735, N1220, N1805);
nor NOR2 (N2205, N2199, N939);
xor XOR2 (N2206, N2200, N1151);
nor NOR4 (N2207, N2206, N1698, N432, N1901);
or OR4 (N2208, N2205, N1702, N1646, N1205);
nand NAND2 (N2209, N2208, N2134);
or OR3 (N2210, N2193, N1842, N1595);
or OR3 (N2211, N2210, N870, N321);
and AND3 (N2212, N2201, N830, N325);
xor XOR2 (N2213, N2183, N1547);
nand NAND4 (N2214, N2203, N1825, N1260, N173);
buf BUF1 (N2215, N2202);
nand NAND3 (N2216, N2207, N2112, N2125);
not NOT1 (N2217, N2213);
and AND2 (N2218, N2190, N884);
or OR4 (N2219, N2212, N184, N545, N1680);
nor NOR2 (N2220, N2214, N478);
nor NOR4 (N2221, N2219, N1935, N1043, N1847);
nand NAND4 (N2222, N2209, N1713, N450, N535);
or OR2 (N2223, N2194, N1052);
not NOT1 (N2224, N2211);
nand NAND3 (N2225, N2222, N1000, N1650);
or OR4 (N2226, N2220, N1254, N939, N1498);
and AND3 (N2227, N2223, N1328, N835);
buf BUF1 (N2228, N2224);
not NOT1 (N2229, N2228);
not NOT1 (N2230, N2227);
or OR2 (N2231, N2215, N501);
not NOT1 (N2232, N2226);
and AND4 (N2233, N2232, N679, N1678, N757);
nor NOR2 (N2234, N2233, N95);
nand NAND4 (N2235, N2225, N1224, N2127, N37);
buf BUF1 (N2236, N2218);
xor XOR2 (N2237, N2229, N122);
xor XOR2 (N2238, N2235, N1739);
nor NOR4 (N2239, N2217, N2231, N1190, N658);
or OR3 (N2240, N803, N1008, N956);
nand NAND3 (N2241, N2237, N2006, N700);
or OR4 (N2242, N2204, N1467, N1823, N1246);
not NOT1 (N2243, N2230);
or OR3 (N2244, N2238, N1425, N1543);
nand NAND2 (N2245, N2240, N725);
or OR4 (N2246, N2244, N862, N767, N191);
nand NAND4 (N2247, N2221, N435, N920, N1688);
and AND3 (N2248, N2216, N2134, N251);
and AND2 (N2249, N2239, N1339);
and AND4 (N2250, N2247, N460, N1622, N1083);
nand NAND3 (N2251, N2243, N2154, N989);
or OR3 (N2252, N2245, N610, N262);
nand NAND4 (N2253, N2249, N1480, N54, N296);
nor NOR3 (N2254, N2234, N335, N1697);
nand NAND4 (N2255, N2250, N870, N27, N261);
nor NOR2 (N2256, N2255, N175);
not NOT1 (N2257, N2248);
xor XOR2 (N2258, N2251, N765);
xor XOR2 (N2259, N2253, N1714);
not NOT1 (N2260, N2241);
nand NAND4 (N2261, N2256, N1605, N1947, N391);
not NOT1 (N2262, N2252);
buf BUF1 (N2263, N2261);
xor XOR2 (N2264, N2254, N117);
or OR2 (N2265, N2257, N207);
or OR3 (N2266, N2259, N1719, N1320);
nor NOR2 (N2267, N2264, N858);
not NOT1 (N2268, N2265);
buf BUF1 (N2269, N2267);
not NOT1 (N2270, N2246);
or OR4 (N2271, N2262, N1307, N1777, N1808);
buf BUF1 (N2272, N2260);
xor XOR2 (N2273, N2263, N996);
nand NAND2 (N2274, N2268, N2056);
buf BUF1 (N2275, N2273);
not NOT1 (N2276, N2272);
buf BUF1 (N2277, N2270);
or OR2 (N2278, N2276, N331);
nor NOR3 (N2279, N2236, N1483, N2271);
xor XOR2 (N2280, N1463, N1668);
or OR3 (N2281, N2269, N1756, N1583);
and AND4 (N2282, N2258, N464, N1125, N868);
xor XOR2 (N2283, N2279, N133);
or OR3 (N2284, N2275, N1688, N318);
and AND2 (N2285, N2282, N987);
not NOT1 (N2286, N2281);
and AND2 (N2287, N2278, N2095);
and AND2 (N2288, N2286, N1123);
or OR3 (N2289, N2285, N938, N234);
or OR2 (N2290, N2277, N1528);
not NOT1 (N2291, N2280);
nor NOR3 (N2292, N2284, N1174, N1236);
nor NOR4 (N2293, N2242, N2207, N1523, N1720);
nand NAND3 (N2294, N2292, N2207, N2237);
nand NAND4 (N2295, N2291, N922, N1220, N931);
nor NOR3 (N2296, N2295, N1464, N165);
not NOT1 (N2297, N2287);
nor NOR4 (N2298, N2290, N733, N1954, N875);
nor NOR3 (N2299, N2266, N561, N743);
and AND3 (N2300, N2296, N675, N692);
or OR3 (N2301, N2299, N707, N655);
not NOT1 (N2302, N2293);
or OR3 (N2303, N2288, N1227, N152);
xor XOR2 (N2304, N2302, N693);
buf BUF1 (N2305, N2303);
nor NOR3 (N2306, N2300, N775, N1211);
nor NOR2 (N2307, N2306, N1552);
buf BUF1 (N2308, N2301);
xor XOR2 (N2309, N2307, N1130);
and AND2 (N2310, N2297, N346);
buf BUF1 (N2311, N2294);
buf BUF1 (N2312, N2310);
buf BUF1 (N2313, N2298);
not NOT1 (N2314, N2308);
nand NAND3 (N2315, N2289, N1905, N1803);
xor XOR2 (N2316, N2309, N89);
or OR4 (N2317, N2283, N306, N1466, N891);
xor XOR2 (N2318, N2312, N655);
not NOT1 (N2319, N2305);
nand NAND3 (N2320, N2318, N1373, N1156);
nand NAND2 (N2321, N2315, N1210);
and AND2 (N2322, N2311, N2144);
xor XOR2 (N2323, N2319, N1614);
or OR4 (N2324, N2314, N2251, N2227, N2194);
or OR4 (N2325, N2304, N2053, N1515, N557);
buf BUF1 (N2326, N2321);
buf BUF1 (N2327, N2274);
nand NAND3 (N2328, N2327, N1104, N572);
nor NOR3 (N2329, N2316, N1001, N391);
xor XOR2 (N2330, N2326, N1343);
buf BUF1 (N2331, N2329);
xor XOR2 (N2332, N2328, N1701);
buf BUF1 (N2333, N2317);
or OR4 (N2334, N2331, N1355, N138, N359);
xor XOR2 (N2335, N2334, N1314);
nor NOR3 (N2336, N2332, N1487, N1489);
and AND2 (N2337, N2325, N1069);
and AND3 (N2338, N2330, N1462, N626);
not NOT1 (N2339, N2335);
buf BUF1 (N2340, N2333);
not NOT1 (N2341, N2322);
or OR4 (N2342, N2340, N1127, N1664, N320);
and AND4 (N2343, N2336, N377, N288, N1471);
buf BUF1 (N2344, N2343);
buf BUF1 (N2345, N2313);
buf BUF1 (N2346, N2320);
buf BUF1 (N2347, N2337);
xor XOR2 (N2348, N2346, N948);
or OR3 (N2349, N2324, N1204, N945);
nor NOR4 (N2350, N2323, N1165, N2066, N1523);
buf BUF1 (N2351, N2344);
nor NOR3 (N2352, N2351, N805, N281);
not NOT1 (N2353, N2349);
and AND4 (N2354, N2350, N1722, N1357, N868);
not NOT1 (N2355, N2347);
xor XOR2 (N2356, N2342, N1135);
and AND2 (N2357, N2353, N332);
not NOT1 (N2358, N2339);
and AND3 (N2359, N2345, N2046, N1338);
or OR3 (N2360, N2356, N1980, N2052);
buf BUF1 (N2361, N2352);
not NOT1 (N2362, N2357);
nor NOR2 (N2363, N2362, N46);
or OR2 (N2364, N2338, N56);
not NOT1 (N2365, N2355);
buf BUF1 (N2366, N2358);
nand NAND2 (N2367, N2366, N1037);
and AND4 (N2368, N2348, N2244, N218, N1677);
nor NOR4 (N2369, N2341, N556, N788, N107);
buf BUF1 (N2370, N2367);
and AND4 (N2371, N2368, N498, N2304, N1826);
xor XOR2 (N2372, N2363, N2105);
nand NAND2 (N2373, N2370, N1011);
nor NOR3 (N2374, N2359, N1009, N1974);
nand NAND4 (N2375, N2374, N1607, N1055, N2042);
buf BUF1 (N2376, N2365);
buf BUF1 (N2377, N2354);
nand NAND4 (N2378, N2369, N245, N1448, N1204);
and AND4 (N2379, N2364, N1380, N274, N586);
and AND2 (N2380, N2376, N1276);
xor XOR2 (N2381, N2380, N2039);
nor NOR4 (N2382, N2373, N477, N857, N130);
not NOT1 (N2383, N2360);
xor XOR2 (N2384, N2383, N588);
nand NAND3 (N2385, N2381, N882, N453);
nor NOR3 (N2386, N2382, N1261, N1669);
not NOT1 (N2387, N2386);
nor NOR4 (N2388, N2375, N319, N1317, N1190);
and AND3 (N2389, N2378, N1160, N342);
nand NAND4 (N2390, N2361, N453, N89, N2240);
or OR2 (N2391, N2388, N1498);
xor XOR2 (N2392, N2377, N2105);
buf BUF1 (N2393, N2379);
nand NAND4 (N2394, N2384, N788, N2332, N1824);
not NOT1 (N2395, N2394);
and AND3 (N2396, N2387, N1058, N1807);
not NOT1 (N2397, N2385);
and AND4 (N2398, N2372, N150, N1625, N2095);
and AND3 (N2399, N2392, N1485, N1176);
and AND4 (N2400, N2396, N1376, N440, N346);
nand NAND2 (N2401, N2393, N2227);
xor XOR2 (N2402, N2400, N2056);
buf BUF1 (N2403, N2402);
not NOT1 (N2404, N2371);
or OR2 (N2405, N2399, N578);
buf BUF1 (N2406, N2403);
not NOT1 (N2407, N2390);
buf BUF1 (N2408, N2405);
xor XOR2 (N2409, N2391, N137);
nor NOR3 (N2410, N2409, N2044, N655);
xor XOR2 (N2411, N2406, N1822);
and AND3 (N2412, N2397, N1864, N10);
or OR4 (N2413, N2407, N1896, N176, N1331);
xor XOR2 (N2414, N2413, N2214);
nand NAND4 (N2415, N2410, N1784, N296, N1924);
or OR2 (N2416, N2411, N2033);
xor XOR2 (N2417, N2415, N289);
buf BUF1 (N2418, N2417);
buf BUF1 (N2419, N2398);
buf BUF1 (N2420, N2401);
buf BUF1 (N2421, N2420);
and AND4 (N2422, N2395, N1969, N1369, N191);
buf BUF1 (N2423, N2414);
xor XOR2 (N2424, N2418, N1180);
buf BUF1 (N2425, N2424);
nand NAND4 (N2426, N2412, N1138, N931, N908);
buf BUF1 (N2427, N2389);
or OR3 (N2428, N2421, N1327, N2195);
nor NOR2 (N2429, N2427, N877);
not NOT1 (N2430, N2429);
and AND4 (N2431, N2425, N1900, N1461, N491);
nor NOR3 (N2432, N2408, N1062, N2105);
or OR3 (N2433, N2431, N1106, N132);
nand NAND2 (N2434, N2422, N2216);
and AND2 (N2435, N2432, N2328);
nand NAND3 (N2436, N2426, N202, N961);
nor NOR2 (N2437, N2435, N1027);
buf BUF1 (N2438, N2437);
buf BUF1 (N2439, N2430);
nand NAND4 (N2440, N2433, N1014, N1590, N451);
xor XOR2 (N2441, N2440, N173);
nor NOR2 (N2442, N2439, N1265);
nand NAND2 (N2443, N2434, N2297);
not NOT1 (N2444, N2416);
nand NAND3 (N2445, N2444, N1560, N2321);
or OR2 (N2446, N2445, N1329);
nand NAND4 (N2447, N2442, N1616, N1984, N2116);
or OR4 (N2448, N2443, N2226, N1953, N959);
xor XOR2 (N2449, N2446, N1543);
or OR3 (N2450, N2447, N1357, N1788);
buf BUF1 (N2451, N2436);
and AND3 (N2452, N2448, N71, N1277);
nand NAND2 (N2453, N2438, N1739);
nor NOR3 (N2454, N2451, N1842, N2013);
nor NOR4 (N2455, N2404, N1299, N2138, N741);
nor NOR3 (N2456, N2449, N1091, N457);
and AND3 (N2457, N2454, N2366, N1128);
xor XOR2 (N2458, N2452, N71);
nor NOR2 (N2459, N2458, N1);
and AND2 (N2460, N2457, N1847);
nand NAND2 (N2461, N2423, N307);
nand NAND3 (N2462, N2453, N1090, N147);
or OR4 (N2463, N2455, N2024, N716, N2416);
not NOT1 (N2464, N2450);
nand NAND4 (N2465, N2460, N2460, N1631, N206);
nand NAND3 (N2466, N2464, N245, N1052);
xor XOR2 (N2467, N2465, N1174);
buf BUF1 (N2468, N2428);
or OR3 (N2469, N2456, N928, N2068);
and AND2 (N2470, N2419, N1200);
xor XOR2 (N2471, N2466, N1952);
nor NOR3 (N2472, N2461, N107, N1231);
or OR2 (N2473, N2469, N537);
buf BUF1 (N2474, N2441);
nor NOR4 (N2475, N2472, N641, N1783, N922);
buf BUF1 (N2476, N2471);
and AND4 (N2477, N2462, N524, N1478, N1777);
nor NOR2 (N2478, N2475, N1646);
nand NAND3 (N2479, N2468, N1259, N1528);
or OR2 (N2480, N2478, N280);
nor NOR4 (N2481, N2473, N968, N1485, N1657);
buf BUF1 (N2482, N2474);
buf BUF1 (N2483, N2477);
buf BUF1 (N2484, N2459);
buf BUF1 (N2485, N2484);
and AND4 (N2486, N2485, N1263, N291, N2471);
and AND3 (N2487, N2480, N1247, N785);
nor NOR3 (N2488, N2467, N694, N2034);
xor XOR2 (N2489, N2487, N2461);
not NOT1 (N2490, N2488);
not NOT1 (N2491, N2479);
and AND3 (N2492, N2491, N510, N1076);
nor NOR3 (N2493, N2463, N304, N1450);
and AND4 (N2494, N2490, N181, N788, N1108);
xor XOR2 (N2495, N2470, N1014);
or OR2 (N2496, N2492, N1122);
not NOT1 (N2497, N2481);
or OR3 (N2498, N2497, N1307, N1360);
xor XOR2 (N2499, N2495, N609);
or OR2 (N2500, N2482, N620);
nand NAND4 (N2501, N2499, N119, N1610, N1533);
not NOT1 (N2502, N2496);
or OR4 (N2503, N2493, N692, N581, N1173);
buf BUF1 (N2504, N2489);
or OR2 (N2505, N2500, N1600);
buf BUF1 (N2506, N2501);
xor XOR2 (N2507, N2504, N876);
or OR2 (N2508, N2494, N1165);
and AND2 (N2509, N2502, N115);
nand NAND3 (N2510, N2509, N195, N924);
and AND4 (N2511, N2498, N1391, N1219, N434);
nor NOR2 (N2512, N2508, N1151);
not NOT1 (N2513, N2507);
or OR3 (N2514, N2506, N612, N660);
nor NOR3 (N2515, N2503, N1080, N936);
not NOT1 (N2516, N2511);
or OR4 (N2517, N2515, N1683, N245, N1973);
and AND4 (N2518, N2516, N360, N1198, N2338);
nand NAND3 (N2519, N2486, N2020, N561);
not NOT1 (N2520, N2510);
nor NOR2 (N2521, N2518, N1017);
buf BUF1 (N2522, N2512);
xor XOR2 (N2523, N2505, N2088);
not NOT1 (N2524, N2517);
nand NAND4 (N2525, N2519, N619, N1000, N1423);
not NOT1 (N2526, N2523);
and AND4 (N2527, N2514, N2149, N964, N1890);
nand NAND3 (N2528, N2524, N1303, N978);
and AND2 (N2529, N2521, N1382);
not NOT1 (N2530, N2483);
and AND2 (N2531, N2527, N314);
or OR4 (N2532, N2531, N1301, N1198, N1712);
nand NAND4 (N2533, N2522, N148, N83, N580);
buf BUF1 (N2534, N2529);
nand NAND3 (N2535, N2528, N1697, N2279);
nor NOR3 (N2536, N2526, N1581, N1044);
and AND3 (N2537, N2534, N2215, N2029);
xor XOR2 (N2538, N2532, N881);
or OR2 (N2539, N2530, N2162);
xor XOR2 (N2540, N2538, N1344);
or OR4 (N2541, N2540, N405, N1911, N829);
or OR2 (N2542, N2536, N1265);
or OR4 (N2543, N2513, N2124, N718, N2156);
nand NAND3 (N2544, N2543, N185, N1682);
and AND3 (N2545, N2539, N620, N1);
nand NAND4 (N2546, N2533, N1078, N219, N795);
and AND3 (N2547, N2542, N165, N1706);
and AND3 (N2548, N2541, N1753, N2317);
xor XOR2 (N2549, N2535, N2156);
or OR3 (N2550, N2520, N1357, N538);
buf BUF1 (N2551, N2525);
xor XOR2 (N2552, N2537, N2280);
and AND3 (N2553, N2549, N913, N364);
or OR4 (N2554, N2544, N978, N669, N1925);
xor XOR2 (N2555, N2545, N2008);
buf BUF1 (N2556, N2554);
or OR2 (N2557, N2556, N954);
buf BUF1 (N2558, N2551);
xor XOR2 (N2559, N2558, N2000);
buf BUF1 (N2560, N2559);
not NOT1 (N2561, N2552);
nor NOR3 (N2562, N2557, N1777, N2298);
nand NAND3 (N2563, N2561, N1348, N967);
nor NOR4 (N2564, N2555, N198, N2152, N398);
nor NOR2 (N2565, N2562, N2551);
nor NOR3 (N2566, N2546, N2449, N1696);
not NOT1 (N2567, N2476);
and AND3 (N2568, N2550, N2126, N1694);
nor NOR2 (N2569, N2548, N1847);
nor NOR2 (N2570, N2547, N1403);
or OR3 (N2571, N2567, N1753, N243);
or OR2 (N2572, N2563, N2045);
nor NOR2 (N2573, N2564, N564);
buf BUF1 (N2574, N2553);
buf BUF1 (N2575, N2566);
xor XOR2 (N2576, N2573, N290);
buf BUF1 (N2577, N2574);
or OR3 (N2578, N2572, N54, N1826);
buf BUF1 (N2579, N2560);
xor XOR2 (N2580, N2568, N375);
not NOT1 (N2581, N2577);
or OR3 (N2582, N2579, N1166, N2126);
not NOT1 (N2583, N2576);
and AND4 (N2584, N2582, N919, N2498, N414);
buf BUF1 (N2585, N2575);
nand NAND4 (N2586, N2581, N717, N2375, N1704);
or OR2 (N2587, N2584, N825);
buf BUF1 (N2588, N2580);
nand NAND3 (N2589, N2569, N1301, N772);
not NOT1 (N2590, N2583);
or OR4 (N2591, N2565, N66, N1000, N1378);
or OR2 (N2592, N2588, N1122);
nor NOR4 (N2593, N2590, N987, N684, N817);
nor NOR4 (N2594, N2586, N1348, N1628, N654);
buf BUF1 (N2595, N2570);
and AND3 (N2596, N2594, N1200, N138);
not NOT1 (N2597, N2592);
nand NAND4 (N2598, N2595, N1116, N588, N2063);
nor NOR3 (N2599, N2571, N2313, N1890);
and AND2 (N2600, N2598, N389);
not NOT1 (N2601, N2596);
not NOT1 (N2602, N2601);
xor XOR2 (N2603, N2600, N2465);
xor XOR2 (N2604, N2591, N1000);
and AND3 (N2605, N2587, N1557, N2293);
nand NAND2 (N2606, N2585, N572);
xor XOR2 (N2607, N2593, N2350);
xor XOR2 (N2608, N2597, N2219);
not NOT1 (N2609, N2607);
nand NAND4 (N2610, N2608, N602, N2246, N2469);
nor NOR3 (N2611, N2589, N771, N1236);
buf BUF1 (N2612, N2602);
nor NOR4 (N2613, N2604, N571, N2279, N950);
buf BUF1 (N2614, N2609);
buf BUF1 (N2615, N2612);
nor NOR2 (N2616, N2611, N20);
nor NOR2 (N2617, N2606, N1706);
not NOT1 (N2618, N2599);
or OR3 (N2619, N2615, N254, N2324);
and AND4 (N2620, N2603, N2525, N776, N1609);
and AND3 (N2621, N2578, N382, N61);
and AND3 (N2622, N2618, N1879, N600);
nor NOR3 (N2623, N2619, N2530, N177);
nand NAND4 (N2624, N2621, N2030, N1766, N1291);
not NOT1 (N2625, N2623);
not NOT1 (N2626, N2616);
nand NAND2 (N2627, N2617, N2200);
xor XOR2 (N2628, N2605, N161);
buf BUF1 (N2629, N2613);
nand NAND2 (N2630, N2622, N581);
and AND2 (N2631, N2627, N735);
buf BUF1 (N2632, N2620);
nor NOR3 (N2633, N2614, N1070, N650);
xor XOR2 (N2634, N2631, N2556);
xor XOR2 (N2635, N2634, N1135);
not NOT1 (N2636, N2628);
xor XOR2 (N2637, N2630, N1297);
nand NAND3 (N2638, N2610, N378, N1048);
nand NAND4 (N2639, N2637, N1684, N1987, N594);
xor XOR2 (N2640, N2632, N1770);
or OR3 (N2641, N2635, N2139, N54);
nor NOR4 (N2642, N2633, N1040, N1493, N2351);
nand NAND2 (N2643, N2629, N2558);
or OR2 (N2644, N2640, N2377);
xor XOR2 (N2645, N2642, N1431);
nand NAND3 (N2646, N2626, N363, N1032);
not NOT1 (N2647, N2639);
nor NOR2 (N2648, N2624, N2544);
xor XOR2 (N2649, N2645, N1937);
nand NAND4 (N2650, N2649, N416, N2316, N1343);
not NOT1 (N2651, N2638);
nor NOR2 (N2652, N2625, N1009);
xor XOR2 (N2653, N2647, N69);
xor XOR2 (N2654, N2646, N420);
or OR2 (N2655, N2652, N2083);
or OR2 (N2656, N2648, N1942);
or OR2 (N2657, N2650, N497);
xor XOR2 (N2658, N2654, N2429);
buf BUF1 (N2659, N2655);
nor NOR2 (N2660, N2659, N949);
and AND2 (N2661, N2651, N2334);
or OR3 (N2662, N2644, N2111, N479);
nor NOR3 (N2663, N2643, N101, N532);
xor XOR2 (N2664, N2661, N2492);
or OR2 (N2665, N2641, N1028);
nand NAND3 (N2666, N2653, N2528, N1032);
buf BUF1 (N2667, N2662);
buf BUF1 (N2668, N2667);
xor XOR2 (N2669, N2636, N1630);
nor NOR4 (N2670, N2656, N2067, N1919, N2187);
nand NAND2 (N2671, N2666, N2619);
nand NAND3 (N2672, N2669, N1647, N2229);
and AND3 (N2673, N2668, N2189, N2355);
not NOT1 (N2674, N2665);
or OR3 (N2675, N2671, N486, N828);
or OR4 (N2676, N2672, N2271, N1791, N312);
nand NAND3 (N2677, N2657, N480, N2187);
and AND2 (N2678, N2673, N1886);
xor XOR2 (N2679, N2670, N2414);
xor XOR2 (N2680, N2674, N2122);
or OR4 (N2681, N2679, N1497, N2264, N1027);
nor NOR4 (N2682, N2678, N626, N466, N620);
nor NOR2 (N2683, N2675, N2196);
xor XOR2 (N2684, N2663, N476);
not NOT1 (N2685, N2658);
nor NOR4 (N2686, N2681, N79, N2051, N1276);
and AND4 (N2687, N2683, N2434, N1690, N1983);
or OR4 (N2688, N2686, N972, N701, N902);
nor NOR2 (N2689, N2685, N1014);
nand NAND2 (N2690, N2680, N2067);
or OR3 (N2691, N2676, N2594, N2182);
or OR3 (N2692, N2690, N2006, N905);
nand NAND3 (N2693, N2682, N288, N2552);
not NOT1 (N2694, N2688);
and AND3 (N2695, N2689, N973, N1748);
xor XOR2 (N2696, N2677, N1856);
nand NAND4 (N2697, N2684, N1637, N1902, N137);
buf BUF1 (N2698, N2696);
nor NOR4 (N2699, N2691, N534, N885, N828);
or OR4 (N2700, N2692, N1035, N886, N1771);
buf BUF1 (N2701, N2694);
nand NAND2 (N2702, N2697, N1525);
nor NOR3 (N2703, N2687, N2605, N1800);
nor NOR4 (N2704, N2660, N1621, N1027, N53);
nor NOR3 (N2705, N2702, N1486, N50);
and AND4 (N2706, N2664, N1882, N1255, N953);
or OR3 (N2707, N2700, N186, N1504);
or OR3 (N2708, N2703, N2491, N1888);
buf BUF1 (N2709, N2706);
not NOT1 (N2710, N2701);
nand NAND3 (N2711, N2707, N1360, N1887);
or OR4 (N2712, N2695, N323, N884, N1565);
buf BUF1 (N2713, N2708);
nor NOR4 (N2714, N2705, N290, N281, N254);
nor NOR4 (N2715, N2710, N1898, N327, N969);
xor XOR2 (N2716, N2709, N192);
or OR4 (N2717, N2712, N230, N230, N253);
not NOT1 (N2718, N2698);
xor XOR2 (N2719, N2713, N113);
or OR4 (N2720, N2719, N2387, N496, N905);
or OR2 (N2721, N2699, N1786);
not NOT1 (N2722, N2715);
not NOT1 (N2723, N2721);
nand NAND2 (N2724, N2711, N84);
nand NAND3 (N2725, N2723, N555, N2161);
nand NAND3 (N2726, N2716, N497, N1865);
nor NOR3 (N2727, N2720, N643, N2672);
not NOT1 (N2728, N2693);
buf BUF1 (N2729, N2727);
nand NAND4 (N2730, N2722, N1651, N1698, N2481);
and AND3 (N2731, N2724, N1364, N1523);
or OR2 (N2732, N2718, N547);
or OR2 (N2733, N2732, N1797);
buf BUF1 (N2734, N2726);
not NOT1 (N2735, N2725);
and AND2 (N2736, N2735, N12);
xor XOR2 (N2737, N2728, N2557);
nor NOR4 (N2738, N2729, N1786, N961, N15);
and AND2 (N2739, N2714, N1684);
xor XOR2 (N2740, N2738, N919);
nor NOR2 (N2741, N2730, N1512);
or OR3 (N2742, N2739, N1149, N83);
and AND3 (N2743, N2734, N1240, N967);
buf BUF1 (N2744, N2737);
xor XOR2 (N2745, N2736, N1398);
buf BUF1 (N2746, N2740);
and AND2 (N2747, N2731, N1447);
nand NAND2 (N2748, N2704, N168);
xor XOR2 (N2749, N2741, N1356);
xor XOR2 (N2750, N2747, N1595);
buf BUF1 (N2751, N2748);
not NOT1 (N2752, N2743);
nand NAND3 (N2753, N2751, N473, N2080);
nand NAND3 (N2754, N2750, N677, N1572);
buf BUF1 (N2755, N2754);
nor NOR4 (N2756, N2749, N2344, N1383, N2239);
and AND2 (N2757, N2717, N920);
not NOT1 (N2758, N2742);
nor NOR4 (N2759, N2758, N648, N1625, N721);
nand NAND3 (N2760, N2752, N299, N797);
not NOT1 (N2761, N2753);
and AND4 (N2762, N2745, N2298, N2048, N1470);
nor NOR2 (N2763, N2759, N1496);
buf BUF1 (N2764, N2746);
or OR4 (N2765, N2755, N2212, N1895, N1413);
or OR3 (N2766, N2761, N1973, N1380);
not NOT1 (N2767, N2763);
xor XOR2 (N2768, N2756, N783);
nor NOR2 (N2769, N2744, N75);
nor NOR3 (N2770, N2766, N2066, N489);
nor NOR4 (N2771, N2757, N214, N2687, N1017);
and AND2 (N2772, N2765, N1372);
buf BUF1 (N2773, N2762);
xor XOR2 (N2774, N2733, N330);
not NOT1 (N2775, N2773);
and AND2 (N2776, N2768, N1240);
or OR3 (N2777, N2776, N896, N2728);
buf BUF1 (N2778, N2775);
or OR4 (N2779, N2772, N1898, N2747, N1877);
buf BUF1 (N2780, N2769);
nor NOR2 (N2781, N2778, N1852);
xor XOR2 (N2782, N2777, N1512);
nor NOR4 (N2783, N2767, N1785, N1259, N745);
buf BUF1 (N2784, N2764);
xor XOR2 (N2785, N2779, N1481);
and AND3 (N2786, N2784, N1134, N2049);
or OR3 (N2787, N2780, N2518, N1845);
buf BUF1 (N2788, N2781);
nor NOR3 (N2789, N2783, N437, N912);
or OR4 (N2790, N2770, N916, N1363, N527);
buf BUF1 (N2791, N2788);
or OR2 (N2792, N2787, N560);
or OR3 (N2793, N2786, N1446, N1717);
xor XOR2 (N2794, N2771, N38);
or OR3 (N2795, N2794, N1020, N2350);
buf BUF1 (N2796, N2793);
buf BUF1 (N2797, N2791);
or OR3 (N2798, N2774, N719, N1120);
or OR2 (N2799, N2785, N948);
nor NOR3 (N2800, N2799, N2565, N1492);
and AND2 (N2801, N2790, N2586);
nand NAND2 (N2802, N2760, N313);
nand NAND4 (N2803, N2797, N1964, N2170, N157);
and AND3 (N2804, N2800, N1762, N2135);
nand NAND2 (N2805, N2802, N1888);
not NOT1 (N2806, N2803);
or OR4 (N2807, N2782, N776, N1925, N1267);
nand NAND4 (N2808, N2798, N354, N1229, N2673);
and AND3 (N2809, N2792, N2135, N1350);
nand NAND2 (N2810, N2796, N2684);
nor NOR3 (N2811, N2804, N104, N1809);
not NOT1 (N2812, N2811);
nor NOR3 (N2813, N2801, N1520, N2010);
or OR3 (N2814, N2813, N2168, N2465);
and AND3 (N2815, N2807, N1166, N1150);
xor XOR2 (N2816, N2808, N2241);
not NOT1 (N2817, N2809);
nand NAND2 (N2818, N2795, N368);
and AND4 (N2819, N2815, N1984, N1752, N1457);
not NOT1 (N2820, N2812);
nand NAND3 (N2821, N2806, N2583, N2371);
xor XOR2 (N2822, N2814, N659);
buf BUF1 (N2823, N2822);
not NOT1 (N2824, N2821);
xor XOR2 (N2825, N2818, N1322);
buf BUF1 (N2826, N2817);
xor XOR2 (N2827, N2825, N2202);
xor XOR2 (N2828, N2816, N1322);
or OR4 (N2829, N2828, N235, N1123, N1940);
nor NOR3 (N2830, N2826, N459, N1162);
or OR4 (N2831, N2824, N2193, N2530, N1639);
and AND2 (N2832, N2829, N2577);
not NOT1 (N2833, N2810);
buf BUF1 (N2834, N2827);
and AND4 (N2835, N2820, N2281, N1711, N458);
xor XOR2 (N2836, N2835, N1398);
and AND2 (N2837, N2823, N1753);
nand NAND4 (N2838, N2789, N1621, N2013, N15);
xor XOR2 (N2839, N2838, N56);
nor NOR2 (N2840, N2830, N2224);
or OR4 (N2841, N2831, N560, N784, N2000);
or OR2 (N2842, N2833, N1591);
not NOT1 (N2843, N2836);
not NOT1 (N2844, N2837);
or OR3 (N2845, N2844, N159, N2443);
and AND3 (N2846, N2842, N781, N286);
nand NAND2 (N2847, N2819, N1366);
not NOT1 (N2848, N2834);
xor XOR2 (N2849, N2847, N706);
nand NAND4 (N2850, N2845, N552, N1090, N1943);
nand NAND2 (N2851, N2850, N2464);
buf BUF1 (N2852, N2843);
and AND2 (N2853, N2848, N2585);
nor NOR2 (N2854, N2846, N1695);
nand NAND2 (N2855, N2840, N2786);
and AND2 (N2856, N2805, N1588);
nor NOR2 (N2857, N2853, N2708);
buf BUF1 (N2858, N2849);
nor NOR3 (N2859, N2854, N1980, N41);
or OR2 (N2860, N2858, N2337);
xor XOR2 (N2861, N2860, N2399);
or OR4 (N2862, N2857, N915, N1048, N1311);
xor XOR2 (N2863, N2856, N410);
not NOT1 (N2864, N2832);
buf BUF1 (N2865, N2863);
buf BUF1 (N2866, N2852);
nand NAND2 (N2867, N2841, N1290);
xor XOR2 (N2868, N2866, N1536);
and AND3 (N2869, N2862, N654, N1564);
not NOT1 (N2870, N2855);
nor NOR3 (N2871, N2851, N1394, N2706);
not NOT1 (N2872, N2864);
and AND4 (N2873, N2839, N1562, N1039, N821);
or OR3 (N2874, N2869, N1503, N97);
xor XOR2 (N2875, N2871, N1209);
buf BUF1 (N2876, N2865);
buf BUF1 (N2877, N2872);
and AND2 (N2878, N2868, N666);
nor NOR4 (N2879, N2859, N1947, N1002, N1542);
nand NAND3 (N2880, N2873, N1107, N292);
xor XOR2 (N2881, N2878, N457);
or OR3 (N2882, N2875, N198, N288);
buf BUF1 (N2883, N2879);
nand NAND2 (N2884, N2880, N2442);
nor NOR2 (N2885, N2882, N433);
xor XOR2 (N2886, N2885, N1970);
nand NAND4 (N2887, N2881, N2551, N2409, N1262);
xor XOR2 (N2888, N2876, N1677);
xor XOR2 (N2889, N2877, N2549);
nand NAND2 (N2890, N2867, N439);
and AND2 (N2891, N2861, N2471);
xor XOR2 (N2892, N2874, N1562);
or OR3 (N2893, N2892, N2878, N475);
or OR2 (N2894, N2884, N540);
and AND3 (N2895, N2888, N355, N1999);
not NOT1 (N2896, N2887);
nand NAND3 (N2897, N2870, N1999, N362);
buf BUF1 (N2898, N2893);
nand NAND4 (N2899, N2898, N995, N1803, N1656);
not NOT1 (N2900, N2889);
not NOT1 (N2901, N2883);
and AND3 (N2902, N2896, N1447, N2801);
buf BUF1 (N2903, N2901);
xor XOR2 (N2904, N2886, N2306);
nor NOR3 (N2905, N2900, N2731, N2422);
not NOT1 (N2906, N2890);
and AND3 (N2907, N2891, N2485, N1853);
buf BUF1 (N2908, N2907);
nor NOR2 (N2909, N2895, N1593);
nor NOR3 (N2910, N2903, N2352, N2158);
not NOT1 (N2911, N2906);
or OR4 (N2912, N2904, N1874, N2786, N1655);
nor NOR2 (N2913, N2902, N1572);
nor NOR4 (N2914, N2911, N262, N672, N2265);
buf BUF1 (N2915, N2897);
nand NAND4 (N2916, N2913, N1449, N2197, N1429);
nor NOR4 (N2917, N2894, N1949, N616, N801);
or OR2 (N2918, N2912, N2788);
nand NAND3 (N2919, N2915, N1295, N2699);
and AND2 (N2920, N2917, N792);
or OR3 (N2921, N2909, N2042, N285);
nand NAND2 (N2922, N2905, N672);
and AND2 (N2923, N2919, N2661);
not NOT1 (N2924, N2918);
nor NOR3 (N2925, N2908, N1107, N2013);
nor NOR4 (N2926, N2899, N504, N456, N1428);
nand NAND4 (N2927, N2926, N835, N1362, N2372);
not NOT1 (N2928, N2914);
xor XOR2 (N2929, N2910, N1274);
or OR4 (N2930, N2924, N1358, N1763, N1525);
nand NAND4 (N2931, N2922, N2572, N1910, N2881);
and AND2 (N2932, N2925, N1863);
nor NOR3 (N2933, N2928, N440, N1929);
not NOT1 (N2934, N2932);
buf BUF1 (N2935, N2934);
not NOT1 (N2936, N2923);
not NOT1 (N2937, N2927);
xor XOR2 (N2938, N2921, N1717);
nand NAND3 (N2939, N2937, N2295, N1355);
or OR3 (N2940, N2920, N289, N301);
or OR3 (N2941, N2935, N702, N636);
and AND2 (N2942, N2931, N1843);
nor NOR2 (N2943, N2938, N1216);
nand NAND3 (N2944, N2933, N2128, N2571);
and AND4 (N2945, N2939, N167, N366, N569);
xor XOR2 (N2946, N2941, N2895);
nand NAND4 (N2947, N2916, N961, N2809, N1634);
xor XOR2 (N2948, N2930, N447);
buf BUF1 (N2949, N2940);
buf BUF1 (N2950, N2936);
or OR3 (N2951, N2948, N1536, N1967);
or OR2 (N2952, N2945, N42);
buf BUF1 (N2953, N2929);
not NOT1 (N2954, N2949);
not NOT1 (N2955, N2953);
xor XOR2 (N2956, N2946, N1648);
nand NAND4 (N2957, N2950, N163, N2572, N1939);
nand NAND2 (N2958, N2943, N1976);
buf BUF1 (N2959, N2952);
not NOT1 (N2960, N2951);
nand NAND2 (N2961, N2944, N1418);
xor XOR2 (N2962, N2954, N762);
or OR4 (N2963, N2955, N114, N121, N657);
or OR3 (N2964, N2962, N2078, N1574);
nor NOR3 (N2965, N2942, N452, N195);
or OR4 (N2966, N2958, N1900, N2002, N2913);
and AND2 (N2967, N2957, N1146);
buf BUF1 (N2968, N2967);
or OR4 (N2969, N2964, N111, N1764, N1218);
or OR3 (N2970, N2969, N2691, N2132);
nand NAND4 (N2971, N2963, N2546, N201, N935);
and AND4 (N2972, N2966, N670, N53, N562);
or OR4 (N2973, N2965, N365, N1204, N2962);
buf BUF1 (N2974, N2970);
nand NAND2 (N2975, N2947, N1334);
or OR4 (N2976, N2973, N2766, N2957, N2073);
and AND3 (N2977, N2975, N1849, N2256);
not NOT1 (N2978, N2960);
buf BUF1 (N2979, N2976);
buf BUF1 (N2980, N2977);
and AND4 (N2981, N2979, N503, N2486, N1131);
and AND4 (N2982, N2971, N2137, N2446, N703);
and AND2 (N2983, N2980, N1564);
xor XOR2 (N2984, N2983, N17);
not NOT1 (N2985, N2981);
xor XOR2 (N2986, N2956, N2361);
xor XOR2 (N2987, N2959, N873);
xor XOR2 (N2988, N2978, N2025);
xor XOR2 (N2989, N2985, N291);
xor XOR2 (N2990, N2972, N2776);
and AND4 (N2991, N2968, N2589, N1327, N610);
buf BUF1 (N2992, N2990);
or OR3 (N2993, N2986, N769, N127);
and AND4 (N2994, N2988, N2193, N2002, N24);
not NOT1 (N2995, N2991);
or OR3 (N2996, N2994, N2722, N1076);
or OR3 (N2997, N2982, N1005, N2214);
and AND2 (N2998, N2989, N390);
xor XOR2 (N2999, N2984, N950);
and AND3 (N3000, N2961, N1131, N2239);
not NOT1 (N3001, N2995);
nor NOR2 (N3002, N2996, N50);
and AND3 (N3003, N2998, N2519, N713);
not NOT1 (N3004, N2987);
nand NAND3 (N3005, N2992, N470, N603);
nand NAND4 (N3006, N3003, N248, N1091, N939);
nand NAND2 (N3007, N2974, N1219);
nand NAND4 (N3008, N2997, N375, N1116, N1763);
or OR3 (N3009, N3008, N1184, N335);
xor XOR2 (N3010, N3006, N1194);
not NOT1 (N3011, N2993);
not NOT1 (N3012, N3004);
xor XOR2 (N3013, N3009, N2088);
xor XOR2 (N3014, N3011, N2038);
nand NAND4 (N3015, N3012, N1328, N1545, N644);
nand NAND3 (N3016, N3015, N2995, N1151);
or OR4 (N3017, N3000, N1983, N2886, N1924);
xor XOR2 (N3018, N3007, N165);
nand NAND3 (N3019, N3010, N69, N2881);
not NOT1 (N3020, N3016);
and AND4 (N3021, N3017, N1207, N1596, N1698);
nor NOR2 (N3022, N3021, N2050);
buf BUF1 (N3023, N3022);
buf BUF1 (N3024, N3005);
not NOT1 (N3025, N3020);
and AND2 (N3026, N3025, N1462);
xor XOR2 (N3027, N3026, N2195);
xor XOR2 (N3028, N3024, N2113);
buf BUF1 (N3029, N3013);
nor NOR3 (N3030, N3029, N1451, N1975);
or OR2 (N3031, N3027, N1789);
and AND4 (N3032, N3001, N82, N854, N1792);
nand NAND3 (N3033, N3018, N2073, N1920);
or OR3 (N3034, N3014, N77, N2014);
nand NAND3 (N3035, N3032, N2406, N1966);
nand NAND2 (N3036, N3028, N2715);
buf BUF1 (N3037, N3019);
nor NOR2 (N3038, N3030, N952);
not NOT1 (N3039, N2999);
buf BUF1 (N3040, N3031);
or OR2 (N3041, N3039, N1403);
nor NOR2 (N3042, N3023, N833);
or OR4 (N3043, N3042, N405, N1916, N2597);
or OR4 (N3044, N3002, N1233, N356, N765);
or OR3 (N3045, N3043, N1777, N550);
nand NAND4 (N3046, N3041, N429, N848, N2502);
nor NOR2 (N3047, N3034, N2462);
nor NOR4 (N3048, N3045, N1216, N540, N376);
xor XOR2 (N3049, N3033, N269);
nand NAND4 (N3050, N3046, N2908, N483, N2562);
nand NAND3 (N3051, N3044, N175, N1714);
nand NAND4 (N3052, N3037, N446, N1222, N1922);
nor NOR4 (N3053, N3040, N635, N1870, N2976);
xor XOR2 (N3054, N3048, N2845);
buf BUF1 (N3055, N3052);
nor NOR4 (N3056, N3050, N2332, N959, N902);
and AND4 (N3057, N3053, N2589, N258, N2405);
not NOT1 (N3058, N3035);
or OR3 (N3059, N3051, N2931, N874);
and AND2 (N3060, N3049, N2692);
not NOT1 (N3061, N3056);
nor NOR2 (N3062, N3059, N757);
xor XOR2 (N3063, N3036, N631);
xor XOR2 (N3064, N3061, N858);
nor NOR2 (N3065, N3060, N309);
nor NOR2 (N3066, N3063, N1313);
buf BUF1 (N3067, N3055);
buf BUF1 (N3068, N3057);
nor NOR4 (N3069, N3064, N1159, N371, N1304);
and AND2 (N3070, N3062, N3011);
not NOT1 (N3071, N3054);
not NOT1 (N3072, N3038);
xor XOR2 (N3073, N3065, N1057);
xor XOR2 (N3074, N3070, N2007);
and AND2 (N3075, N3066, N620);
nor NOR4 (N3076, N3073, N1020, N669, N124);
nor NOR4 (N3077, N3058, N214, N367, N1196);
not NOT1 (N3078, N3047);
not NOT1 (N3079, N3077);
not NOT1 (N3080, N3075);
xor XOR2 (N3081, N3068, N468);
buf BUF1 (N3082, N3079);
nand NAND4 (N3083, N3081, N987, N2706, N2539);
nand NAND3 (N3084, N3074, N413, N1064);
not NOT1 (N3085, N3069);
buf BUF1 (N3086, N3072);
and AND4 (N3087, N3084, N2530, N2408, N799);
nand NAND3 (N3088, N3071, N1678, N1015);
and AND2 (N3089, N3083, N2554);
not NOT1 (N3090, N3089);
xor XOR2 (N3091, N3085, N2881);
nand NAND3 (N3092, N3088, N986, N1067);
xor XOR2 (N3093, N3067, N414);
nand NAND4 (N3094, N3093, N2329, N1151, N2560);
buf BUF1 (N3095, N3082);
nor NOR4 (N3096, N3086, N1094, N2646, N2177);
and AND4 (N3097, N3078, N1460, N2443, N2701);
not NOT1 (N3098, N3076);
buf BUF1 (N3099, N3087);
xor XOR2 (N3100, N3080, N2735);
nor NOR2 (N3101, N3090, N885);
buf BUF1 (N3102, N3092);
nand NAND3 (N3103, N3097, N245, N1731);
buf BUF1 (N3104, N3102);
nand NAND2 (N3105, N3103, N1298);
buf BUF1 (N3106, N3095);
xor XOR2 (N3107, N3100, N1885);
and AND2 (N3108, N3104, N49);
not NOT1 (N3109, N3094);
nand NAND2 (N3110, N3107, N481);
not NOT1 (N3111, N3091);
nand NAND4 (N3112, N3109, N3068, N2982, N529);
nor NOR4 (N3113, N3108, N2157, N918, N3035);
and AND2 (N3114, N3096, N3027);
nor NOR2 (N3115, N3113, N206);
or OR3 (N3116, N3111, N965, N1444);
nand NAND3 (N3117, N3110, N2693, N1620);
and AND2 (N3118, N3115, N536);
nand NAND2 (N3119, N3101, N1785);
nor NOR2 (N3120, N3106, N2288);
and AND4 (N3121, N3114, N104, N966, N222);
not NOT1 (N3122, N3105);
or OR2 (N3123, N3118, N2713);
buf BUF1 (N3124, N3117);
not NOT1 (N3125, N3119);
nand NAND3 (N3126, N3120, N1665, N151);
nand NAND2 (N3127, N3112, N1668);
buf BUF1 (N3128, N3116);
buf BUF1 (N3129, N3127);
not NOT1 (N3130, N3128);
nand NAND3 (N3131, N3098, N1601, N1736);
not NOT1 (N3132, N3129);
xor XOR2 (N3133, N3131, N1091);
not NOT1 (N3134, N3124);
buf BUF1 (N3135, N3123);
and AND3 (N3136, N3099, N864, N1561);
nor NOR4 (N3137, N3135, N1434, N1099, N546);
not NOT1 (N3138, N3136);
buf BUF1 (N3139, N3137);
xor XOR2 (N3140, N3130, N1455);
nand NAND4 (N3141, N3132, N2604, N2533, N1520);
not NOT1 (N3142, N3138);
not NOT1 (N3143, N3140);
and AND4 (N3144, N3134, N2951, N99, N14);
and AND3 (N3145, N3141, N314, N2563);
xor XOR2 (N3146, N3122, N731);
nand NAND4 (N3147, N3121, N2593, N313, N970);
xor XOR2 (N3148, N3139, N1396);
not NOT1 (N3149, N3144);
nand NAND4 (N3150, N3148, N2486, N2100, N2931);
xor XOR2 (N3151, N3126, N1100);
nor NOR2 (N3152, N3151, N2760);
and AND3 (N3153, N3146, N3032, N2245);
or OR4 (N3154, N3152, N295, N2623, N2139);
and AND4 (N3155, N3150, N1144, N1630, N1421);
not NOT1 (N3156, N3143);
xor XOR2 (N3157, N3155, N2477);
or OR3 (N3158, N3147, N2428, N1253);
buf BUF1 (N3159, N3142);
nand NAND3 (N3160, N3159, N2486, N1824);
nand NAND4 (N3161, N3149, N257, N988, N2020);
and AND2 (N3162, N3158, N558);
and AND2 (N3163, N3154, N2954);
nor NOR2 (N3164, N3157, N529);
not NOT1 (N3165, N3161);
not NOT1 (N3166, N3163);
xor XOR2 (N3167, N3160, N2065);
or OR4 (N3168, N3167, N2825, N736, N2928);
or OR3 (N3169, N3133, N507, N118);
nand NAND4 (N3170, N3125, N1856, N2961, N759);
nor NOR2 (N3171, N3165, N2841);
or OR4 (N3172, N3145, N505, N803, N1373);
xor XOR2 (N3173, N3171, N1309);
xor XOR2 (N3174, N3162, N864);
xor XOR2 (N3175, N3166, N3134);
or OR4 (N3176, N3169, N1241, N2015, N2242);
not NOT1 (N3177, N3172);
buf BUF1 (N3178, N3168);
xor XOR2 (N3179, N3156, N684);
buf BUF1 (N3180, N3164);
or OR2 (N3181, N3174, N2087);
not NOT1 (N3182, N3173);
nand NAND4 (N3183, N3176, N2177, N402, N1889);
nor NOR3 (N3184, N3178, N2224, N2968);
or OR4 (N3185, N3180, N1787, N3179, N2864);
or OR4 (N3186, N1696, N3119, N2477, N846);
or OR2 (N3187, N3175, N2614);
nand NAND4 (N3188, N3183, N2035, N3163, N1197);
not NOT1 (N3189, N3181);
not NOT1 (N3190, N3187);
nor NOR3 (N3191, N3189, N1293, N74);
nor NOR3 (N3192, N3186, N1612, N2951);
buf BUF1 (N3193, N3190);
nor NOR4 (N3194, N3185, N2275, N277, N1232);
xor XOR2 (N3195, N3193, N2351);
buf BUF1 (N3196, N3170);
nor NOR3 (N3197, N3191, N756, N1766);
nand NAND3 (N3198, N3153, N2593, N660);
nor NOR3 (N3199, N3182, N1607, N1955);
or OR3 (N3200, N3177, N3116, N268);
nor NOR3 (N3201, N3198, N854, N861);
or OR3 (N3202, N3192, N1365, N2631);
buf BUF1 (N3203, N3188);
and AND4 (N3204, N3195, N501, N2467, N2087);
nand NAND2 (N3205, N3197, N1885);
and AND4 (N3206, N3202, N2631, N1900, N3091);
and AND2 (N3207, N3200, N852);
and AND4 (N3208, N3196, N457, N2354, N2073);
nand NAND4 (N3209, N3207, N286, N567, N2416);
buf BUF1 (N3210, N3194);
nor NOR4 (N3211, N3205, N3025, N972, N2195);
not NOT1 (N3212, N3203);
nor NOR3 (N3213, N3204, N602, N2610);
nand NAND2 (N3214, N3210, N1819);
buf BUF1 (N3215, N3199);
xor XOR2 (N3216, N3214, N1998);
nor NOR2 (N3217, N3208, N2690);
and AND3 (N3218, N3217, N1705, N2141);
not NOT1 (N3219, N3209);
xor XOR2 (N3220, N3215, N652);
and AND4 (N3221, N3212, N446, N2510, N960);
nor NOR4 (N3222, N3220, N2136, N541, N866);
buf BUF1 (N3223, N3206);
and AND3 (N3224, N3219, N319, N231);
buf BUF1 (N3225, N3221);
buf BUF1 (N3226, N3211);
or OR4 (N3227, N3226, N1967, N2754, N2828);
nor NOR4 (N3228, N3223, N1660, N83, N1207);
not NOT1 (N3229, N3213);
or OR4 (N3230, N3222, N444, N2247, N2463);
or OR4 (N3231, N3229, N119, N134, N3149);
or OR3 (N3232, N3218, N2136, N2906);
not NOT1 (N3233, N3227);
xor XOR2 (N3234, N3231, N373);
xor XOR2 (N3235, N3224, N2551);
xor XOR2 (N3236, N3201, N565);
and AND4 (N3237, N3234, N527, N2591, N2449);
or OR3 (N3238, N3230, N1396, N2151);
nor NOR4 (N3239, N3216, N1143, N2769, N2554);
nor NOR4 (N3240, N3225, N69, N852, N2819);
nand NAND2 (N3241, N3184, N2693);
nand NAND3 (N3242, N3228, N880, N1092);
not NOT1 (N3243, N3236);
buf BUF1 (N3244, N3243);
buf BUF1 (N3245, N3233);
buf BUF1 (N3246, N3238);
or OR3 (N3247, N3244, N2047, N1993);
and AND2 (N3248, N3239, N688);
not NOT1 (N3249, N3245);
or OR2 (N3250, N3232, N2806);
buf BUF1 (N3251, N3249);
nand NAND2 (N3252, N3237, N3215);
not NOT1 (N3253, N3240);
xor XOR2 (N3254, N3250, N1744);
xor XOR2 (N3255, N3253, N1103);
buf BUF1 (N3256, N3246);
buf BUF1 (N3257, N3255);
or OR2 (N3258, N3256, N2651);
buf BUF1 (N3259, N3242);
nor NOR2 (N3260, N3248, N2150);
and AND2 (N3261, N3260, N27);
buf BUF1 (N3262, N3251);
nor NOR2 (N3263, N3254, N1939);
nand NAND3 (N3264, N3263, N2648, N2332);
buf BUF1 (N3265, N3262);
nand NAND4 (N3266, N3247, N2353, N1333, N87);
not NOT1 (N3267, N3259);
not NOT1 (N3268, N3265);
nor NOR4 (N3269, N3241, N1595, N228, N2007);
nor NOR4 (N3270, N3266, N1854, N2265, N1808);
nand NAND2 (N3271, N3261, N2134);
xor XOR2 (N3272, N3267, N3254);
nand NAND3 (N3273, N3264, N1234, N75);
and AND2 (N3274, N3258, N3161);
or OR3 (N3275, N3274, N314, N964);
buf BUF1 (N3276, N3252);
not NOT1 (N3277, N3235);
or OR2 (N3278, N3273, N3111);
nor NOR2 (N3279, N3277, N2996);
and AND3 (N3280, N3257, N2264, N572);
xor XOR2 (N3281, N3280, N1916);
nor NOR2 (N3282, N3270, N1016);
nand NAND2 (N3283, N3269, N1587);
xor XOR2 (N3284, N3283, N692);
nand NAND3 (N3285, N3268, N3268, N842);
or OR2 (N3286, N3278, N939);
nor NOR2 (N3287, N3285, N1338);
nand NAND2 (N3288, N3271, N1205);
buf BUF1 (N3289, N3287);
buf BUF1 (N3290, N3289);
not NOT1 (N3291, N3288);
or OR4 (N3292, N3275, N2443, N789, N2214);
and AND3 (N3293, N3279, N30, N876);
nor NOR2 (N3294, N3284, N3135);
xor XOR2 (N3295, N3286, N743);
nor NOR3 (N3296, N3276, N762, N197);
not NOT1 (N3297, N3295);
or OR3 (N3298, N3293, N2653, N1315);
nand NAND3 (N3299, N3297, N1516, N1067);
or OR2 (N3300, N3292, N879);
and AND4 (N3301, N3291, N1204, N1872, N1753);
and AND2 (N3302, N3290, N2811);
not NOT1 (N3303, N3301);
or OR2 (N3304, N3299, N3184);
nor NOR2 (N3305, N3298, N2586);
not NOT1 (N3306, N3302);
xor XOR2 (N3307, N3296, N2977);
and AND2 (N3308, N3304, N2227);
or OR2 (N3309, N3294, N837);
nand NAND3 (N3310, N3307, N2721, N735);
nor NOR4 (N3311, N3305, N298, N583, N2102);
xor XOR2 (N3312, N3281, N148);
or OR2 (N3313, N3300, N1835);
not NOT1 (N3314, N3282);
buf BUF1 (N3315, N3310);
buf BUF1 (N3316, N3315);
and AND3 (N3317, N3303, N4, N1240);
or OR3 (N3318, N3312, N120, N1619);
nand NAND2 (N3319, N3316, N1561);
xor XOR2 (N3320, N3308, N2396);
nor NOR2 (N3321, N3318, N844);
xor XOR2 (N3322, N3321, N1816);
nand NAND2 (N3323, N3272, N2034);
or OR4 (N3324, N3313, N415, N1414, N1760);
xor XOR2 (N3325, N3324, N1391);
nand NAND3 (N3326, N3325, N290, N1345);
not NOT1 (N3327, N3314);
nand NAND4 (N3328, N3322, N102, N2658, N274);
not NOT1 (N3329, N3320);
and AND3 (N3330, N3319, N115, N976);
or OR4 (N3331, N3326, N469, N1789, N649);
buf BUF1 (N3332, N3331);
nor NOR2 (N3333, N3328, N2126);
nand NAND2 (N3334, N3327, N2758);
or OR4 (N3335, N3309, N42, N2896, N3323);
or OR4 (N3336, N2459, N2793, N399, N3307);
xor XOR2 (N3337, N3330, N145);
nor NOR3 (N3338, N3333, N3211, N2446);
not NOT1 (N3339, N3329);
nor NOR4 (N3340, N3332, N536, N3029, N2037);
nand NAND4 (N3341, N3335, N1386, N2502, N3338);
and AND2 (N3342, N2587, N820);
and AND3 (N3343, N3334, N407, N403);
xor XOR2 (N3344, N3336, N426);
nor NOR3 (N3345, N3317, N37, N2091);
nand NAND2 (N3346, N3341, N1927);
xor XOR2 (N3347, N3344, N1548);
nor NOR3 (N3348, N3340, N451, N656);
buf BUF1 (N3349, N3311);
xor XOR2 (N3350, N3347, N468);
or OR4 (N3351, N3346, N1564, N982, N2241);
xor XOR2 (N3352, N3349, N1468);
and AND2 (N3353, N3339, N132);
xor XOR2 (N3354, N3306, N2723);
and AND2 (N3355, N3345, N1057);
buf BUF1 (N3356, N3355);
buf BUF1 (N3357, N3343);
xor XOR2 (N3358, N3352, N1296);
xor XOR2 (N3359, N3351, N2126);
or OR3 (N3360, N3356, N2273, N446);
or OR4 (N3361, N3348, N845, N2458, N3253);
xor XOR2 (N3362, N3361, N2373);
nor NOR4 (N3363, N3353, N2781, N299, N2005);
nand NAND2 (N3364, N3357, N2968);
not NOT1 (N3365, N3363);
nor NOR4 (N3366, N3360, N1160, N1267, N2145);
not NOT1 (N3367, N3342);
or OR4 (N3368, N3366, N2531, N1467, N681);
not NOT1 (N3369, N3354);
xor XOR2 (N3370, N3364, N648);
xor XOR2 (N3371, N3350, N626);
nand NAND4 (N3372, N3368, N856, N2746, N469);
xor XOR2 (N3373, N3370, N1596);
not NOT1 (N3374, N3372);
and AND4 (N3375, N3374, N1846, N313, N2681);
and AND2 (N3376, N3358, N676);
not NOT1 (N3377, N3362);
not NOT1 (N3378, N3365);
and AND4 (N3379, N3359, N371, N2639, N2654);
and AND4 (N3380, N3375, N1781, N1360, N409);
or OR2 (N3381, N3377, N1326);
or OR4 (N3382, N3373, N2866, N3164, N3178);
not NOT1 (N3383, N3369);
or OR2 (N3384, N3382, N319);
and AND3 (N3385, N3380, N2165, N3203);
nand NAND3 (N3386, N3367, N1700, N1213);
nor NOR2 (N3387, N3385, N3078);
and AND4 (N3388, N3381, N975, N935, N1978);
nor NOR4 (N3389, N3378, N2979, N86, N3);
nor NOR4 (N3390, N3384, N3231, N1566, N864);
or OR2 (N3391, N3383, N2424);
or OR4 (N3392, N3376, N994, N445, N3324);
or OR2 (N3393, N3388, N1447);
nor NOR3 (N3394, N3389, N249, N1739);
and AND3 (N3395, N3393, N1142, N11);
nor NOR3 (N3396, N3390, N3395, N3065);
and AND2 (N3397, N1516, N1373);
not NOT1 (N3398, N3386);
not NOT1 (N3399, N3396);
buf BUF1 (N3400, N3394);
not NOT1 (N3401, N3391);
or OR3 (N3402, N3371, N3287, N284);
nor NOR2 (N3403, N3401, N2824);
or OR2 (N3404, N3400, N2341);
and AND2 (N3405, N3403, N2797);
or OR4 (N3406, N3402, N2930, N3190, N2316);
xor XOR2 (N3407, N3379, N2324);
nand NAND3 (N3408, N3398, N2732, N2081);
not NOT1 (N3409, N3387);
nor NOR4 (N3410, N3397, N1437, N3105, N444);
nor NOR3 (N3411, N3406, N243, N2413);
or OR4 (N3412, N3411, N927, N1119, N158);
buf BUF1 (N3413, N3410);
or OR4 (N3414, N3409, N3197, N380, N2993);
nor NOR3 (N3415, N3404, N3176, N2500);
buf BUF1 (N3416, N3337);
buf BUF1 (N3417, N3399);
or OR4 (N3418, N3414, N1719, N1130, N67);
not NOT1 (N3419, N3405);
nand NAND3 (N3420, N3419, N3105, N2489);
and AND3 (N3421, N3415, N2609, N2851);
and AND4 (N3422, N3407, N2243, N45, N2746);
nand NAND4 (N3423, N3416, N2079, N3005, N2912);
nor NOR2 (N3424, N3423, N1866);
nand NAND2 (N3425, N3422, N1582);
nor NOR4 (N3426, N3418, N819, N2678, N1373);
xor XOR2 (N3427, N3426, N846);
not NOT1 (N3428, N3427);
nor NOR4 (N3429, N3425, N2873, N1166, N1147);
nand NAND3 (N3430, N3408, N755, N2898);
buf BUF1 (N3431, N3412);
nand NAND3 (N3432, N3429, N2135, N375);
not NOT1 (N3433, N3417);
or OR4 (N3434, N3430, N3051, N1486, N1874);
xor XOR2 (N3435, N3420, N2863);
and AND3 (N3436, N3421, N2428, N2934);
and AND3 (N3437, N3435, N1201, N1515);
xor XOR2 (N3438, N3432, N2498);
xor XOR2 (N3439, N3437, N3429);
and AND2 (N3440, N3431, N1252);
nand NAND3 (N3441, N3438, N2945, N2749);
buf BUF1 (N3442, N3434);
or OR2 (N3443, N3413, N2215);
xor XOR2 (N3444, N3441, N2124);
not NOT1 (N3445, N3439);
xor XOR2 (N3446, N3428, N1225);
not NOT1 (N3447, N3444);
and AND2 (N3448, N3442, N3137);
buf BUF1 (N3449, N3445);
nand NAND2 (N3450, N3448, N1486);
or OR4 (N3451, N3446, N1380, N436, N1444);
or OR4 (N3452, N3436, N2935, N876, N1019);
nand NAND2 (N3453, N3440, N3020);
buf BUF1 (N3454, N3452);
and AND4 (N3455, N3392, N2659, N2047, N1957);
and AND2 (N3456, N3450, N1706);
and AND2 (N3457, N3424, N1946);
buf BUF1 (N3458, N3451);
nand NAND2 (N3459, N3455, N1293);
or OR4 (N3460, N3456, N2703, N2305, N573);
buf BUF1 (N3461, N3458);
nor NOR4 (N3462, N3453, N465, N570, N2337);
nor NOR4 (N3463, N3460, N1056, N2868, N2951);
and AND3 (N3464, N3461, N600, N1918);
buf BUF1 (N3465, N3457);
not NOT1 (N3466, N3459);
or OR4 (N3467, N3449, N354, N119, N1925);
buf BUF1 (N3468, N3433);
xor XOR2 (N3469, N3465, N2895);
not NOT1 (N3470, N3468);
xor XOR2 (N3471, N3462, N2185);
or OR2 (N3472, N3466, N123);
xor XOR2 (N3473, N3467, N2411);
buf BUF1 (N3474, N3454);
nor NOR2 (N3475, N3469, N3431);
and AND4 (N3476, N3475, N479, N1452, N1765);
buf BUF1 (N3477, N3472);
not NOT1 (N3478, N3470);
or OR3 (N3479, N3474, N2242, N2769);
buf BUF1 (N3480, N3464);
or OR4 (N3481, N3480, N2011, N326, N2279);
and AND3 (N3482, N3477, N355, N1766);
xor XOR2 (N3483, N3471, N2423);
and AND3 (N3484, N3479, N622, N2679);
buf BUF1 (N3485, N3447);
buf BUF1 (N3486, N3481);
or OR3 (N3487, N3484, N2081, N2977);
nor NOR3 (N3488, N3485, N2068, N3310);
nor NOR3 (N3489, N3476, N339, N1990);
nand NAND2 (N3490, N3463, N2211);
and AND4 (N3491, N3483, N927, N1224, N1715);
and AND3 (N3492, N3487, N1004, N2925);
xor XOR2 (N3493, N3490, N1646);
nor NOR4 (N3494, N3482, N1632, N9, N2733);
buf BUF1 (N3495, N3492);
buf BUF1 (N3496, N3473);
xor XOR2 (N3497, N3496, N3277);
and AND4 (N3498, N3478, N1098, N1175, N518);
xor XOR2 (N3499, N3495, N2681);
not NOT1 (N3500, N3486);
or OR3 (N3501, N3494, N1461, N3307);
nand NAND3 (N3502, N3500, N1552, N218);
or OR3 (N3503, N3499, N642, N2105);
buf BUF1 (N3504, N3488);
or OR4 (N3505, N3497, N2301, N748, N2940);
nor NOR3 (N3506, N3493, N97, N137);
nand NAND4 (N3507, N3489, N3241, N1508, N2809);
nand NAND3 (N3508, N3491, N977, N1750);
nor NOR3 (N3509, N3505, N2950, N3012);
not NOT1 (N3510, N3507);
and AND4 (N3511, N3503, N1343, N1252, N869);
buf BUF1 (N3512, N3510);
not NOT1 (N3513, N3501);
nand NAND4 (N3514, N3509, N2051, N508, N3049);
buf BUF1 (N3515, N3502);
nand NAND4 (N3516, N3513, N1443, N2935, N3267);
nor NOR2 (N3517, N3514, N2456);
or OR4 (N3518, N3508, N2953, N2179, N1125);
and AND3 (N3519, N3498, N458, N3457);
nand NAND4 (N3520, N3511, N50, N1926, N159);
xor XOR2 (N3521, N3519, N3150);
buf BUF1 (N3522, N3516);
not NOT1 (N3523, N3518);
nand NAND3 (N3524, N3523, N2525, N598);
and AND2 (N3525, N3521, N67);
not NOT1 (N3526, N3520);
nor NOR2 (N3527, N3504, N1035);
not NOT1 (N3528, N3524);
and AND3 (N3529, N3506, N818, N1249);
buf BUF1 (N3530, N3512);
buf BUF1 (N3531, N3530);
xor XOR2 (N3532, N3515, N1262);
or OR3 (N3533, N3532, N1992, N2239);
or OR3 (N3534, N3533, N482, N776);
nor NOR2 (N3535, N3528, N353);
xor XOR2 (N3536, N3443, N843);
buf BUF1 (N3537, N3525);
nand NAND2 (N3538, N3536, N2388);
nand NAND3 (N3539, N3538, N2902, N218);
not NOT1 (N3540, N3522);
and AND2 (N3541, N3526, N3473);
and AND2 (N3542, N3527, N2287);
nor NOR2 (N3543, N3540, N2588);
not NOT1 (N3544, N3534);
nand NAND4 (N3545, N3544, N866, N2062, N474);
nor NOR2 (N3546, N3542, N415);
or OR3 (N3547, N3535, N2351, N2147);
or OR3 (N3548, N3543, N3259, N2657);
buf BUF1 (N3549, N3531);
and AND4 (N3550, N3545, N1336, N1076, N1430);
or OR4 (N3551, N3541, N2106, N1056, N1109);
or OR4 (N3552, N3549, N2559, N1848, N2693);
nor NOR4 (N3553, N3550, N3313, N3024, N1670);
nor NOR2 (N3554, N3529, N2285);
or OR2 (N3555, N3554, N255);
or OR2 (N3556, N3548, N2268);
nand NAND3 (N3557, N3551, N77, N1355);
buf BUF1 (N3558, N3517);
xor XOR2 (N3559, N3558, N39);
buf BUF1 (N3560, N3547);
or OR3 (N3561, N3559, N1577, N461);
not NOT1 (N3562, N3555);
and AND3 (N3563, N3552, N2869, N2405);
xor XOR2 (N3564, N3557, N724);
nand NAND2 (N3565, N3563, N1054);
xor XOR2 (N3566, N3562, N1744);
nor NOR2 (N3567, N3566, N1569);
xor XOR2 (N3568, N3560, N518);
and AND3 (N3569, N3564, N3137, N187);
and AND3 (N3570, N3556, N1544, N966);
buf BUF1 (N3571, N3537);
or OR4 (N3572, N3553, N3236, N1908, N2720);
nand NAND4 (N3573, N3569, N2693, N3466, N1154);
nor NOR4 (N3574, N3565, N937, N2630, N683);
xor XOR2 (N3575, N3572, N3535);
nor NOR3 (N3576, N3574, N1475, N1304);
nand NAND2 (N3577, N3575, N1866);
or OR3 (N3578, N3539, N1633, N2975);
and AND2 (N3579, N3568, N627);
or OR4 (N3580, N3546, N1811, N1137, N2556);
or OR3 (N3581, N3578, N806, N59);
or OR2 (N3582, N3577, N2224);
or OR3 (N3583, N3581, N2190, N1454);
nor NOR4 (N3584, N3570, N2018, N2730, N1348);
xor XOR2 (N3585, N3573, N1502);
buf BUF1 (N3586, N3585);
buf BUF1 (N3587, N3579);
not NOT1 (N3588, N3582);
nor NOR2 (N3589, N3588, N2604);
nor NOR2 (N3590, N3571, N1754);
nor NOR3 (N3591, N3583, N3374, N2865);
and AND2 (N3592, N3567, N180);
not NOT1 (N3593, N3576);
nand NAND3 (N3594, N3584, N2671, N1863);
nor NOR3 (N3595, N3587, N1815, N155);
nand NAND3 (N3596, N3561, N3111, N139);
nor NOR4 (N3597, N3595, N2968, N331, N493);
or OR4 (N3598, N3597, N636, N878, N1055);
nand NAND2 (N3599, N3589, N2460);
buf BUF1 (N3600, N3591);
nor NOR3 (N3601, N3594, N701, N2268);
or OR4 (N3602, N3599, N3579, N3314, N3198);
and AND4 (N3603, N3586, N2981, N1822, N3448);
xor XOR2 (N3604, N3590, N1443);
nand NAND3 (N3605, N3593, N1169, N854);
and AND3 (N3606, N3598, N2633, N1629);
nor NOR2 (N3607, N3596, N3176);
nor NOR4 (N3608, N3603, N2463, N64, N2899);
xor XOR2 (N3609, N3608, N1600);
nand NAND2 (N3610, N3601, N1659);
buf BUF1 (N3611, N3610);
buf BUF1 (N3612, N3602);
not NOT1 (N3613, N3600);
not NOT1 (N3614, N3613);
not NOT1 (N3615, N3604);
buf BUF1 (N3616, N3580);
and AND3 (N3617, N3606, N1952, N2636);
xor XOR2 (N3618, N3592, N2485);
or OR2 (N3619, N3616, N2793);
nor NOR3 (N3620, N3605, N798, N737);
nand NAND4 (N3621, N3615, N3479, N3377, N1368);
not NOT1 (N3622, N3619);
xor XOR2 (N3623, N3614, N2213);
nor NOR2 (N3624, N3622, N2832);
or OR3 (N3625, N3612, N93, N3510);
nand NAND3 (N3626, N3618, N2085, N325);
not NOT1 (N3627, N3620);
nor NOR3 (N3628, N3623, N999, N1425);
buf BUF1 (N3629, N3628);
not NOT1 (N3630, N3611);
nand NAND3 (N3631, N3607, N399, N713);
buf BUF1 (N3632, N3629);
or OR3 (N3633, N3621, N808, N1338);
nor NOR2 (N3634, N3627, N3471);
nand NAND2 (N3635, N3626, N1615);
buf BUF1 (N3636, N3633);
xor XOR2 (N3637, N3609, N3431);
nand NAND2 (N3638, N3635, N1756);
and AND2 (N3639, N3631, N1395);
and AND4 (N3640, N3625, N886, N110, N3325);
or OR4 (N3641, N3638, N2342, N1524, N2416);
nand NAND3 (N3642, N3617, N2125, N3457);
buf BUF1 (N3643, N3630);
nor NOR4 (N3644, N3640, N2210, N2896, N1707);
nor NOR4 (N3645, N3644, N1062, N598, N2796);
not NOT1 (N3646, N3636);
nor NOR4 (N3647, N3643, N1058, N1870, N1640);
not NOT1 (N3648, N3641);
xor XOR2 (N3649, N3639, N1202);
xor XOR2 (N3650, N3624, N1113);
xor XOR2 (N3651, N3649, N2195);
and AND4 (N3652, N3646, N914, N180, N3545);
buf BUF1 (N3653, N3647);
or OR2 (N3654, N3645, N2513);
buf BUF1 (N3655, N3651);
not NOT1 (N3656, N3654);
buf BUF1 (N3657, N3656);
not NOT1 (N3658, N3632);
and AND2 (N3659, N3655, N2515);
or OR4 (N3660, N3653, N587, N2758, N3195);
nor NOR2 (N3661, N3659, N226);
xor XOR2 (N3662, N3634, N1867);
nor NOR2 (N3663, N3657, N2564);
and AND3 (N3664, N3650, N660, N1745);
and AND3 (N3665, N3648, N568, N10);
and AND3 (N3666, N3637, N1398, N3500);
and AND2 (N3667, N3664, N1584);
and AND2 (N3668, N3666, N2483);
or OR3 (N3669, N3662, N3188, N2374);
not NOT1 (N3670, N3668);
or OR3 (N3671, N3652, N50, N1110);
and AND3 (N3672, N3665, N1091, N3172);
or OR4 (N3673, N3672, N1472, N1951, N1827);
nand NAND3 (N3674, N3661, N20, N2142);
buf BUF1 (N3675, N3642);
xor XOR2 (N3676, N3673, N3134);
and AND4 (N3677, N3670, N472, N1606, N2018);
nor NOR4 (N3678, N3674, N529, N709, N1798);
and AND3 (N3679, N3671, N6, N1901);
xor XOR2 (N3680, N3658, N1747);
nor NOR4 (N3681, N3677, N2499, N2318, N24);
xor XOR2 (N3682, N3679, N3024);
nand NAND2 (N3683, N3663, N385);
buf BUF1 (N3684, N3676);
or OR3 (N3685, N3669, N2473, N3551);
and AND2 (N3686, N3667, N1468);
or OR4 (N3687, N3675, N1579, N3661, N1869);
xor XOR2 (N3688, N3681, N536);
or OR2 (N3689, N3660, N1360);
xor XOR2 (N3690, N3686, N409);
nor NOR4 (N3691, N3680, N583, N368, N1640);
buf BUF1 (N3692, N3683);
nor NOR4 (N3693, N3684, N3548, N2282, N2556);
not NOT1 (N3694, N3692);
nand NAND3 (N3695, N3693, N2799, N929);
and AND2 (N3696, N3694, N2345);
and AND2 (N3697, N3688, N2915);
and AND2 (N3698, N3690, N3341);
buf BUF1 (N3699, N3691);
buf BUF1 (N3700, N3696);
buf BUF1 (N3701, N3698);
and AND2 (N3702, N3685, N1903);
and AND4 (N3703, N3699, N3142, N495, N1948);
and AND3 (N3704, N3700, N2016, N747);
or OR3 (N3705, N3682, N3378, N504);
xor XOR2 (N3706, N3678, N3701);
nor NOR3 (N3707, N2523, N159, N1107);
and AND3 (N3708, N3702, N3115, N1246);
nand NAND4 (N3709, N3697, N350, N1098, N2250);
nor NOR2 (N3710, N3695, N1437);
and AND3 (N3711, N3710, N11, N3487);
not NOT1 (N3712, N3704);
xor XOR2 (N3713, N3709, N2550);
not NOT1 (N3714, N3707);
or OR4 (N3715, N3706, N3449, N2585, N1124);
nor NOR4 (N3716, N3714, N2776, N1324, N1482);
or OR3 (N3717, N3716, N696, N3099);
not NOT1 (N3718, N3689);
nor NOR2 (N3719, N3718, N3441);
xor XOR2 (N3720, N3687, N3297);
nor NOR4 (N3721, N3703, N1392, N3241, N639);
not NOT1 (N3722, N3719);
not NOT1 (N3723, N3717);
or OR4 (N3724, N3720, N718, N1862, N1946);
buf BUF1 (N3725, N3708);
and AND4 (N3726, N3711, N1607, N1450, N1680);
nand NAND4 (N3727, N3712, N2586, N1414, N1193);
or OR3 (N3728, N3725, N319, N3550);
or OR3 (N3729, N3727, N1754, N2647);
nand NAND3 (N3730, N3722, N3292, N74);
or OR4 (N3731, N3713, N211, N3260, N1550);
nor NOR3 (N3732, N3730, N516, N32);
buf BUF1 (N3733, N3715);
or OR3 (N3734, N3732, N865, N925);
nand NAND3 (N3735, N3726, N3289, N2425);
nor NOR2 (N3736, N3728, N1402);
xor XOR2 (N3737, N3724, N3702);
or OR4 (N3738, N3735, N2006, N354, N137);
xor XOR2 (N3739, N3737, N1519);
nand NAND4 (N3740, N3723, N2575, N2226, N1782);
not NOT1 (N3741, N3705);
buf BUF1 (N3742, N3734);
nand NAND2 (N3743, N3739, N3206);
xor XOR2 (N3744, N3740, N2267);
buf BUF1 (N3745, N3733);
and AND2 (N3746, N3736, N3719);
nand NAND3 (N3747, N3742, N195, N653);
xor XOR2 (N3748, N3743, N1590);
xor XOR2 (N3749, N3747, N2861);
buf BUF1 (N3750, N3738);
not NOT1 (N3751, N3750);
not NOT1 (N3752, N3748);
nor NOR3 (N3753, N3749, N1691, N388);
buf BUF1 (N3754, N3746);
not NOT1 (N3755, N3753);
or OR2 (N3756, N3755, N1968);
and AND4 (N3757, N3731, N929, N1157, N2873);
and AND4 (N3758, N3752, N2247, N1248, N3152);
or OR2 (N3759, N3756, N3451);
buf BUF1 (N3760, N3757);
or OR2 (N3761, N3754, N2283);
xor XOR2 (N3762, N3745, N2681);
not NOT1 (N3763, N3729);
nand NAND3 (N3764, N3758, N2308, N3045);
nand NAND2 (N3765, N3762, N2840);
not NOT1 (N3766, N3764);
not NOT1 (N3767, N3766);
and AND2 (N3768, N3721, N1532);
not NOT1 (N3769, N3768);
xor XOR2 (N3770, N3760, N2252);
or OR4 (N3771, N3761, N1136, N3606, N3148);
not NOT1 (N3772, N3767);
or OR4 (N3773, N3759, N1709, N2131, N574);
buf BUF1 (N3774, N3772);
buf BUF1 (N3775, N3744);
not NOT1 (N3776, N3771);
and AND3 (N3777, N3765, N3423, N3124);
nor NOR3 (N3778, N3777, N1868, N1743);
not NOT1 (N3779, N3751);
buf BUF1 (N3780, N3779);
and AND2 (N3781, N3780, N2506);
nand NAND2 (N3782, N3776, N2902);
or OR4 (N3783, N3769, N1182, N2010, N1026);
and AND3 (N3784, N3783, N3521, N1004);
or OR2 (N3785, N3773, N1987);
nor NOR3 (N3786, N3778, N1832, N2871);
nand NAND4 (N3787, N3786, N1886, N1720, N1711);
nand NAND2 (N3788, N3787, N1297);
and AND2 (N3789, N3763, N452);
nor NOR3 (N3790, N3789, N866, N1175);
nor NOR3 (N3791, N3775, N1101, N54);
or OR3 (N3792, N3781, N3075, N1241);
nor NOR2 (N3793, N3788, N1847);
and AND3 (N3794, N3790, N2118, N2790);
nor NOR3 (N3795, N3793, N1905, N1746);
buf BUF1 (N3796, N3741);
nand NAND4 (N3797, N3796, N3009, N3158, N2954);
or OR2 (N3798, N3792, N1058);
nor NOR2 (N3799, N3774, N770);
xor XOR2 (N3800, N3770, N1292);
xor XOR2 (N3801, N3791, N2227);
not NOT1 (N3802, N3782);
buf BUF1 (N3803, N3785);
buf BUF1 (N3804, N3801);
xor XOR2 (N3805, N3784, N3130);
or OR3 (N3806, N3804, N2871, N2924);
not NOT1 (N3807, N3799);
and AND2 (N3808, N3806, N1417);
or OR4 (N3809, N3803, N2671, N2363, N3575);
and AND2 (N3810, N3800, N713);
nand NAND2 (N3811, N3798, N90);
or OR4 (N3812, N3794, N2420, N1564, N1077);
nor NOR4 (N3813, N3795, N2544, N282, N3107);
buf BUF1 (N3814, N3805);
nand NAND3 (N3815, N3812, N260, N811);
xor XOR2 (N3816, N3802, N844);
nand NAND2 (N3817, N3815, N689);
nor NOR3 (N3818, N3808, N2957, N1795);
nand NAND3 (N3819, N3814, N144, N2912);
or OR2 (N3820, N3816, N1890);
nor NOR3 (N3821, N3797, N1530, N1027);
buf BUF1 (N3822, N3807);
nor NOR3 (N3823, N3813, N2415, N1606);
or OR3 (N3824, N3822, N1062, N3404);
not NOT1 (N3825, N3824);
not NOT1 (N3826, N3821);
or OR4 (N3827, N3820, N1685, N2493, N1111);
nor NOR3 (N3828, N3809, N1398, N1558);
buf BUF1 (N3829, N3818);
and AND2 (N3830, N3819, N1369);
nand NAND2 (N3831, N3825, N2043);
not NOT1 (N3832, N3829);
and AND3 (N3833, N3832, N2604, N3683);
and AND2 (N3834, N3810, N167);
nor NOR2 (N3835, N3817, N786);
and AND2 (N3836, N3833, N2970);
nor NOR2 (N3837, N3830, N1792);
not NOT1 (N3838, N3811);
not NOT1 (N3839, N3831);
buf BUF1 (N3840, N3836);
and AND2 (N3841, N3835, N2177);
buf BUF1 (N3842, N3839);
nor NOR4 (N3843, N3837, N2357, N3163, N3240);
nand NAND2 (N3844, N3823, N1445);
buf BUF1 (N3845, N3842);
or OR2 (N3846, N3841, N3776);
not NOT1 (N3847, N3846);
nand NAND4 (N3848, N3838, N3575, N771, N270);
not NOT1 (N3849, N3843);
buf BUF1 (N3850, N3844);
nand NAND4 (N3851, N3827, N1097, N3340, N848);
and AND4 (N3852, N3834, N2087, N1398, N2341);
or OR3 (N3853, N3847, N1788, N920);
nand NAND2 (N3854, N3845, N514);
and AND3 (N3855, N3854, N3015, N2050);
nand NAND2 (N3856, N3826, N3041);
not NOT1 (N3857, N3851);
buf BUF1 (N3858, N3857);
xor XOR2 (N3859, N3855, N2307);
not NOT1 (N3860, N3852);
nor NOR3 (N3861, N3840, N2060, N2742);
not NOT1 (N3862, N3858);
and AND4 (N3863, N3850, N2438, N2203, N3523);
or OR4 (N3864, N3849, N3191, N1153, N216);
nand NAND4 (N3865, N3853, N3585, N140, N2159);
nor NOR2 (N3866, N3863, N286);
xor XOR2 (N3867, N3848, N282);
nand NAND3 (N3868, N3861, N2266, N1923);
or OR3 (N3869, N3864, N3841, N2021);
and AND4 (N3870, N3860, N2925, N1449, N2925);
or OR2 (N3871, N3870, N1414);
nand NAND2 (N3872, N3868, N32);
nand NAND4 (N3873, N3867, N3785, N1459, N2089);
xor XOR2 (N3874, N3862, N3848);
and AND3 (N3875, N3871, N3601, N2121);
nand NAND2 (N3876, N3875, N611);
not NOT1 (N3877, N3873);
xor XOR2 (N3878, N3866, N2287);
or OR4 (N3879, N3876, N2947, N3330, N1274);
nor NOR3 (N3880, N3865, N3216, N1475);
and AND3 (N3881, N3828, N3235, N982);
nand NAND3 (N3882, N3856, N1456, N826);
nor NOR2 (N3883, N3869, N614);
or OR2 (N3884, N3879, N670);
buf BUF1 (N3885, N3859);
nand NAND4 (N3886, N3874, N2122, N743, N3324);
nand NAND3 (N3887, N3886, N1007, N3157);
nor NOR3 (N3888, N3872, N880, N3458);
xor XOR2 (N3889, N3881, N1546);
nand NAND4 (N3890, N3885, N691, N3722, N3669);
and AND4 (N3891, N3890, N94, N1772, N845);
or OR3 (N3892, N3883, N2743, N169);
or OR3 (N3893, N3887, N2415, N1943);
nor NOR4 (N3894, N3880, N2247, N2611, N2844);
or OR3 (N3895, N3878, N2394, N1789);
not NOT1 (N3896, N3895);
and AND4 (N3897, N3892, N420, N1266, N3426);
and AND3 (N3898, N3891, N522, N1022);
buf BUF1 (N3899, N3889);
not NOT1 (N3900, N3882);
and AND2 (N3901, N3877, N524);
buf BUF1 (N3902, N3894);
buf BUF1 (N3903, N3888);
and AND3 (N3904, N3903, N422, N731);
xor XOR2 (N3905, N3901, N923);
nor NOR3 (N3906, N3893, N3282, N3876);
nand NAND3 (N3907, N3897, N607, N1820);
nor NOR4 (N3908, N3898, N912, N1501, N3511);
or OR3 (N3909, N3899, N1631, N2670);
buf BUF1 (N3910, N3909);
nor NOR4 (N3911, N3906, N1797, N1981, N3517);
nand NAND2 (N3912, N3900, N31);
buf BUF1 (N3913, N3904);
not NOT1 (N3914, N3884);
nand NAND2 (N3915, N3905, N3890);
buf BUF1 (N3916, N3896);
or OR2 (N3917, N3916, N1304);
buf BUF1 (N3918, N3911);
not NOT1 (N3919, N3902);
and AND2 (N3920, N3918, N3323);
not NOT1 (N3921, N3908);
or OR4 (N3922, N3913, N1645, N1648, N963);
buf BUF1 (N3923, N3907);
nand NAND2 (N3924, N3917, N1918);
and AND2 (N3925, N3915, N3522);
nor NOR4 (N3926, N3919, N828, N2111, N2450);
and AND4 (N3927, N3926, N142, N2433, N2289);
xor XOR2 (N3928, N3922, N2168);
nand NAND4 (N3929, N3923, N576, N1968, N1577);
buf BUF1 (N3930, N3927);
nand NAND3 (N3931, N3920, N3050, N2977);
buf BUF1 (N3932, N3928);
nor NOR4 (N3933, N3914, N3469, N3618, N176);
buf BUF1 (N3934, N3932);
and AND4 (N3935, N3929, N3304, N759, N699);
nand NAND4 (N3936, N3924, N2316, N3112, N3495);
xor XOR2 (N3937, N3933, N1004);
and AND2 (N3938, N3921, N684);
and AND4 (N3939, N3935, N2974, N3039, N3238);
or OR4 (N3940, N3931, N487, N2960, N397);
buf BUF1 (N3941, N3910);
buf BUF1 (N3942, N3925);
not NOT1 (N3943, N3938);
and AND4 (N3944, N3912, N665, N3190, N859);
not NOT1 (N3945, N3937);
buf BUF1 (N3946, N3934);
nand NAND2 (N3947, N3930, N2019);
not NOT1 (N3948, N3939);
xor XOR2 (N3949, N3941, N567);
or OR2 (N3950, N3942, N561);
not NOT1 (N3951, N3949);
nand NAND2 (N3952, N3948, N3458);
buf BUF1 (N3953, N3947);
and AND3 (N3954, N3950, N1741, N491);
nor NOR2 (N3955, N3953, N580);
and AND3 (N3956, N3943, N839, N2234);
and AND3 (N3957, N3944, N2334, N2678);
not NOT1 (N3958, N3957);
and AND2 (N3959, N3940, N531);
and AND4 (N3960, N3946, N1049, N1446, N22);
or OR2 (N3961, N3952, N1152);
and AND3 (N3962, N3958, N337, N2104);
or OR4 (N3963, N3951, N1135, N2169, N1291);
nor NOR3 (N3964, N3954, N1735, N131);
xor XOR2 (N3965, N3962, N3650);
nand NAND3 (N3966, N3963, N2481, N1429);
nand NAND2 (N3967, N3955, N2440);
or OR2 (N3968, N3961, N3293);
and AND3 (N3969, N3964, N1110, N3950);
buf BUF1 (N3970, N3969);
xor XOR2 (N3971, N3967, N2186);
not NOT1 (N3972, N3970);
nor NOR2 (N3973, N3968, N1132);
xor XOR2 (N3974, N3959, N748);
buf BUF1 (N3975, N3972);
nor NOR4 (N3976, N3960, N599, N2315, N2319);
not NOT1 (N3977, N3965);
or OR3 (N3978, N3966, N1809, N2668);
xor XOR2 (N3979, N3936, N1021);
or OR3 (N3980, N3971, N331, N2923);
and AND4 (N3981, N3974, N2828, N1685, N441);
buf BUF1 (N3982, N3976);
buf BUF1 (N3983, N3945);
xor XOR2 (N3984, N3973, N1053);
buf BUF1 (N3985, N3984);
not NOT1 (N3986, N3956);
not NOT1 (N3987, N3981);
and AND4 (N3988, N3977, N2145, N2461, N2364);
not NOT1 (N3989, N3987);
buf BUF1 (N3990, N3989);
or OR4 (N3991, N3985, N2751, N3577, N3933);
nand NAND4 (N3992, N3982, N3975, N40, N2039);
not NOT1 (N3993, N1514);
buf BUF1 (N3994, N3978);
xor XOR2 (N3995, N3980, N3074);
and AND3 (N3996, N3992, N820, N1873);
and AND4 (N3997, N3994, N462, N2688, N388);
buf BUF1 (N3998, N3979);
nand NAND2 (N3999, N3997, N1139);
not NOT1 (N4000, N3999);
not NOT1 (N4001, N3983);
or OR3 (N4002, N3995, N1439, N620);
nand NAND2 (N4003, N4001, N3961);
nand NAND2 (N4004, N3996, N3028);
not NOT1 (N4005, N3991);
nand NAND4 (N4006, N3988, N2598, N3485, N1616);
xor XOR2 (N4007, N4002, N998);
xor XOR2 (N4008, N3998, N998);
or OR4 (N4009, N4000, N2097, N3747, N1959);
buf BUF1 (N4010, N4008);
xor XOR2 (N4011, N4010, N1785);
nand NAND2 (N4012, N4007, N433);
nor NOR2 (N4013, N3990, N3374);
or OR4 (N4014, N3993, N1140, N1794, N2245);
buf BUF1 (N4015, N4003);
and AND3 (N4016, N4009, N593, N1009);
and AND4 (N4017, N4016, N15, N2392, N2490);
or OR4 (N4018, N4005, N945, N3928, N1043);
xor XOR2 (N4019, N4012, N3161);
or OR3 (N4020, N4014, N3143, N3283);
and AND3 (N4021, N4015, N2409, N107);
or OR2 (N4022, N4011, N2500);
nor NOR3 (N4023, N4017, N2710, N1609);
nor NOR4 (N4024, N4019, N3100, N1245, N2808);
buf BUF1 (N4025, N4021);
nor NOR2 (N4026, N4024, N2748);
and AND4 (N4027, N4006, N842, N231, N2711);
and AND4 (N4028, N4018, N196, N1999, N1032);
not NOT1 (N4029, N4027);
and AND4 (N4030, N4022, N2475, N2399, N3841);
or OR2 (N4031, N4030, N1856);
xor XOR2 (N4032, N4023, N1194);
nor NOR3 (N4033, N4026, N2403, N2590);
or OR3 (N4034, N4032, N1740, N3004);
nor NOR3 (N4035, N4025, N1307, N1603);
xor XOR2 (N4036, N4013, N1445);
xor XOR2 (N4037, N4031, N111);
buf BUF1 (N4038, N4037);
nand NAND2 (N4039, N3986, N58);
buf BUF1 (N4040, N4038);
nand NAND3 (N4041, N4036, N2086, N609);
and AND4 (N4042, N4029, N1148, N1250, N1716);
and AND2 (N4043, N4035, N2854);
nor NOR4 (N4044, N4033, N3548, N1082, N1230);
and AND2 (N4045, N4044, N3057);
xor XOR2 (N4046, N4004, N1036);
nand NAND4 (N4047, N4041, N821, N50, N1668);
buf BUF1 (N4048, N4028);
nand NAND4 (N4049, N4040, N1787, N2123, N2358);
xor XOR2 (N4050, N4039, N3132);
nand NAND2 (N4051, N4048, N3264);
buf BUF1 (N4052, N4050);
nor NOR3 (N4053, N4052, N523, N674);
and AND2 (N4054, N4053, N2294);
nand NAND2 (N4055, N4020, N3406);
not NOT1 (N4056, N4043);
nor NOR4 (N4057, N4054, N3008, N1064, N110);
and AND3 (N4058, N4047, N893, N645);
or OR4 (N4059, N4051, N3364, N920, N2046);
nor NOR3 (N4060, N4034, N4049, N1875);
or OR4 (N4061, N2843, N3862, N1335, N3576);
xor XOR2 (N4062, N4046, N202);
or OR2 (N4063, N4057, N1871);
nor NOR2 (N4064, N4063, N1960);
or OR3 (N4065, N4064, N3325, N2746);
or OR3 (N4066, N4045, N638, N514);
or OR3 (N4067, N4058, N2719, N1776);
nand NAND4 (N4068, N4042, N2251, N3638, N2728);
or OR4 (N4069, N4056, N2500, N3123, N2816);
not NOT1 (N4070, N4069);
nand NAND3 (N4071, N4065, N2889, N245);
nand NAND3 (N4072, N4068, N1658, N886);
not NOT1 (N4073, N4060);
nor NOR4 (N4074, N4071, N693, N3763, N1284);
and AND3 (N4075, N4073, N971, N2376);
and AND2 (N4076, N4062, N2940);
or OR3 (N4077, N4055, N2838, N1978);
and AND2 (N4078, N4074, N2399);
buf BUF1 (N4079, N4076);
or OR4 (N4080, N4059, N935, N4053, N2470);
not NOT1 (N4081, N4066);
buf BUF1 (N4082, N4070);
and AND2 (N4083, N4080, N3012);
nand NAND2 (N4084, N4075, N919);
and AND3 (N4085, N4082, N956, N1221);
and AND3 (N4086, N4079, N800, N2542);
and AND3 (N4087, N4084, N1831, N1940);
buf BUF1 (N4088, N4083);
not NOT1 (N4089, N4087);
xor XOR2 (N4090, N4072, N191);
not NOT1 (N4091, N4078);
xor XOR2 (N4092, N4077, N1564);
nor NOR4 (N4093, N4061, N4005, N524, N1877);
not NOT1 (N4094, N4067);
nor NOR4 (N4095, N4092, N3863, N56, N2982);
nor NOR4 (N4096, N4091, N1335, N2944, N2377);
or OR2 (N4097, N4085, N2171);
nand NAND2 (N4098, N4095, N1986);
or OR4 (N4099, N4097, N2146, N3489, N294);
buf BUF1 (N4100, N4089);
nor NOR4 (N4101, N4088, N1339, N347, N2327);
and AND3 (N4102, N4096, N144, N1787);
nor NOR3 (N4103, N4098, N1856, N1878);
buf BUF1 (N4104, N4086);
nor NOR4 (N4105, N4081, N3594, N827, N1139);
or OR2 (N4106, N4103, N3842);
or OR3 (N4107, N4094, N589, N702);
xor XOR2 (N4108, N4100, N836);
and AND3 (N4109, N4105, N4068, N1891);
nand NAND3 (N4110, N4101, N337, N924);
or OR2 (N4111, N4099, N822);
nor NOR4 (N4112, N4093, N3790, N985, N1869);
buf BUF1 (N4113, N4112);
not NOT1 (N4114, N4104);
nor NOR3 (N4115, N4113, N665, N1367);
xor XOR2 (N4116, N4107, N3066);
xor XOR2 (N4117, N4114, N793);
nand NAND4 (N4118, N4115, N539, N1787, N2621);
and AND3 (N4119, N4118, N2107, N2329);
xor XOR2 (N4120, N4111, N1047);
xor XOR2 (N4121, N4110, N3902);
not NOT1 (N4122, N4117);
or OR2 (N4123, N4122, N1309);
nor NOR2 (N4124, N4108, N2729);
nor NOR4 (N4125, N4116, N2049, N403, N2536);
or OR3 (N4126, N4123, N1873, N1791);
or OR2 (N4127, N4125, N3822);
buf BUF1 (N4128, N4102);
or OR3 (N4129, N4126, N3119, N3501);
not NOT1 (N4130, N4106);
buf BUF1 (N4131, N4129);
not NOT1 (N4132, N4124);
or OR2 (N4133, N4120, N3232);
not NOT1 (N4134, N4131);
nand NAND2 (N4135, N4109, N1704);
nor NOR2 (N4136, N4090, N803);
xor XOR2 (N4137, N4128, N576);
nor NOR3 (N4138, N4137, N3809, N1231);
nand NAND4 (N4139, N4135, N3345, N2910, N3441);
xor XOR2 (N4140, N4121, N3148);
and AND3 (N4141, N4127, N3587, N1158);
xor XOR2 (N4142, N4138, N807);
buf BUF1 (N4143, N4142);
buf BUF1 (N4144, N4140);
not NOT1 (N4145, N4139);
and AND2 (N4146, N4136, N131);
nor NOR3 (N4147, N4133, N854, N3258);
nor NOR4 (N4148, N4134, N1539, N221, N1475);
nor NOR2 (N4149, N4132, N2521);
buf BUF1 (N4150, N4119);
and AND4 (N4151, N4144, N1715, N3361, N440);
not NOT1 (N4152, N4143);
nor NOR2 (N4153, N4151, N1078);
or OR2 (N4154, N4145, N3547);
nand NAND3 (N4155, N4147, N3392, N354);
buf BUF1 (N4156, N4152);
or OR3 (N4157, N4148, N953, N109);
nand NAND4 (N4158, N4155, N2011, N211, N978);
nand NAND2 (N4159, N4158, N989);
not NOT1 (N4160, N4149);
not NOT1 (N4161, N4150);
nand NAND3 (N4162, N4146, N1974, N3783);
nor NOR2 (N4163, N4153, N3219);
nor NOR3 (N4164, N4162, N3964, N2678);
nand NAND4 (N4165, N4156, N3488, N3301, N1046);
and AND3 (N4166, N4130, N822, N3430);
and AND2 (N4167, N4141, N1651);
or OR4 (N4168, N4165, N3416, N2283, N3516);
or OR4 (N4169, N4161, N869, N2788, N876);
nand NAND2 (N4170, N4168, N1771);
not NOT1 (N4171, N4160);
buf BUF1 (N4172, N4166);
and AND4 (N4173, N4169, N3019, N2472, N3933);
xor XOR2 (N4174, N4171, N3486);
xor XOR2 (N4175, N4163, N1760);
not NOT1 (N4176, N4170);
or OR2 (N4177, N4176, N1417);
not NOT1 (N4178, N4173);
or OR2 (N4179, N4172, N2292);
xor XOR2 (N4180, N4174, N616);
and AND3 (N4181, N4179, N1463, N101);
or OR4 (N4182, N4178, N2051, N155, N213);
nor NOR2 (N4183, N4159, N930);
nand NAND2 (N4184, N4177, N815);
and AND4 (N4185, N4167, N639, N1305, N2275);
not NOT1 (N4186, N4164);
buf BUF1 (N4187, N4183);
or OR4 (N4188, N4186, N2358, N2030, N3132);
or OR4 (N4189, N4184, N3671, N1040, N196);
xor XOR2 (N4190, N4157, N242);
or OR2 (N4191, N4188, N2196);
and AND2 (N4192, N4180, N1791);
not NOT1 (N4193, N4185);
nand NAND2 (N4194, N4189, N3669);
xor XOR2 (N4195, N4175, N2271);
not NOT1 (N4196, N4190);
or OR3 (N4197, N4192, N505, N974);
or OR3 (N4198, N4196, N2362, N3659);
not NOT1 (N4199, N4181);
buf BUF1 (N4200, N4182);
nand NAND2 (N4201, N4197, N1679);
or OR2 (N4202, N4187, N1756);
nor NOR4 (N4203, N4199, N1078, N1379, N942);
not NOT1 (N4204, N4201);
buf BUF1 (N4205, N4200);
nor NOR3 (N4206, N4203, N3393, N312);
not NOT1 (N4207, N4191);
nand NAND3 (N4208, N4193, N883, N2313);
or OR4 (N4209, N4204, N897, N38, N3185);
or OR3 (N4210, N4195, N2520, N685);
or OR3 (N4211, N4207, N565, N1023);
and AND3 (N4212, N4211, N1262, N3440);
nor NOR2 (N4213, N4212, N2323);
or OR3 (N4214, N4206, N130, N2191);
or OR3 (N4215, N4208, N3202, N2178);
and AND4 (N4216, N4202, N3025, N1343, N2857);
not NOT1 (N4217, N4213);
buf BUF1 (N4218, N4215);
not NOT1 (N4219, N4218);
nand NAND2 (N4220, N4210, N2385);
not NOT1 (N4221, N4217);
nand NAND3 (N4222, N4219, N627, N2271);
and AND4 (N4223, N4220, N2095, N429, N1839);
not NOT1 (N4224, N4216);
xor XOR2 (N4225, N4209, N4163);
and AND3 (N4226, N4221, N504, N2102);
not NOT1 (N4227, N4223);
not NOT1 (N4228, N4224);
nand NAND4 (N4229, N4225, N3797, N1087, N2838);
or OR2 (N4230, N4194, N1994);
or OR4 (N4231, N4227, N1248, N4223, N261);
xor XOR2 (N4232, N4222, N776);
nand NAND2 (N4233, N4198, N1279);
nor NOR2 (N4234, N4154, N550);
buf BUF1 (N4235, N4214);
nor NOR3 (N4236, N4231, N3587, N1958);
xor XOR2 (N4237, N4205, N83);
buf BUF1 (N4238, N4226);
xor XOR2 (N4239, N4230, N659);
and AND3 (N4240, N4239, N1898, N2064);
nor NOR2 (N4241, N4240, N1896);
not NOT1 (N4242, N4229);
and AND2 (N4243, N4234, N1465);
nand NAND4 (N4244, N4238, N1795, N766, N3395);
not NOT1 (N4245, N4228);
and AND3 (N4246, N4245, N345, N2617);
buf BUF1 (N4247, N4242);
nand NAND4 (N4248, N4243, N2522, N1225, N3902);
xor XOR2 (N4249, N4237, N2933);
nand NAND3 (N4250, N4249, N1028, N1125);
buf BUF1 (N4251, N4241);
nor NOR4 (N4252, N4232, N2926, N578, N3143);
or OR4 (N4253, N4236, N1776, N2972, N4205);
buf BUF1 (N4254, N4250);
xor XOR2 (N4255, N4244, N2859);
or OR4 (N4256, N4251, N683, N1049, N1725);
not NOT1 (N4257, N4255);
or OR4 (N4258, N4254, N1158, N1409, N1630);
and AND3 (N4259, N4246, N252, N896);
and AND2 (N4260, N4259, N2875);
nand NAND4 (N4261, N4257, N915, N1842, N1217);
nor NOR4 (N4262, N4247, N2968, N4133, N2027);
or OR4 (N4263, N4261, N406, N2747, N196);
buf BUF1 (N4264, N4263);
xor XOR2 (N4265, N4260, N1965);
not NOT1 (N4266, N4235);
nand NAND4 (N4267, N4262, N2193, N253, N1276);
nor NOR4 (N4268, N4264, N2658, N3067, N620);
not NOT1 (N4269, N4256);
and AND4 (N4270, N4248, N3310, N4043, N813);
xor XOR2 (N4271, N4267, N213);
or OR3 (N4272, N4253, N837, N2284);
and AND4 (N4273, N4258, N3157, N2983, N1864);
xor XOR2 (N4274, N4272, N900);
and AND4 (N4275, N4265, N2761, N3738, N3817);
or OR4 (N4276, N4233, N3206, N54, N4011);
nand NAND3 (N4277, N4271, N3182, N3394);
nand NAND2 (N4278, N4270, N2205);
xor XOR2 (N4279, N4268, N1921);
or OR3 (N4280, N4275, N4170, N3494);
buf BUF1 (N4281, N4269);
nand NAND2 (N4282, N4277, N2497);
xor XOR2 (N4283, N4273, N1164);
and AND2 (N4284, N4252, N3950);
not NOT1 (N4285, N4281);
or OR4 (N4286, N4276, N4166, N3613, N4217);
xor XOR2 (N4287, N4282, N763);
xor XOR2 (N4288, N4287, N1571);
buf BUF1 (N4289, N4274);
xor XOR2 (N4290, N4286, N2679);
xor XOR2 (N4291, N4288, N1714);
xor XOR2 (N4292, N4283, N900);
nand NAND2 (N4293, N4289, N1108);
xor XOR2 (N4294, N4278, N1530);
and AND2 (N4295, N4292, N336);
and AND2 (N4296, N4293, N401);
or OR2 (N4297, N4285, N297);
nand NAND3 (N4298, N4296, N2961, N755);
xor XOR2 (N4299, N4280, N3798);
not NOT1 (N4300, N4295);
not NOT1 (N4301, N4298);
and AND2 (N4302, N4297, N2767);
nor NOR2 (N4303, N4301, N1070);
buf BUF1 (N4304, N4299);
buf BUF1 (N4305, N4290);
nor NOR3 (N4306, N4303, N3951, N3923);
and AND3 (N4307, N4284, N809, N1060);
xor XOR2 (N4308, N4279, N1725);
not NOT1 (N4309, N4294);
not NOT1 (N4310, N4302);
nor NOR3 (N4311, N4300, N1307, N3839);
and AND3 (N4312, N4309, N3753, N86);
xor XOR2 (N4313, N4308, N3682);
not NOT1 (N4314, N4313);
nor NOR4 (N4315, N4305, N1735, N3453, N4244);
or OR4 (N4316, N4310, N2342, N814, N2088);
nor NOR2 (N4317, N4307, N2968);
or OR3 (N4318, N4314, N3516, N3354);
buf BUF1 (N4319, N4315);
buf BUF1 (N4320, N4318);
and AND3 (N4321, N4291, N2553, N3692);
or OR4 (N4322, N4312, N312, N2940, N3397);
nor NOR2 (N4323, N4322, N2536);
and AND4 (N4324, N4266, N3688, N3525, N783);
nor NOR3 (N4325, N4316, N1478, N3812);
or OR4 (N4326, N4325, N2610, N1636, N859);
buf BUF1 (N4327, N4326);
nand NAND2 (N4328, N4320, N2784);
nor NOR2 (N4329, N4324, N4026);
nor NOR4 (N4330, N4327, N3641, N2729, N1762);
xor XOR2 (N4331, N4323, N730);
nand NAND2 (N4332, N4329, N2454);
and AND2 (N4333, N4306, N2632);
or OR2 (N4334, N4317, N1615);
or OR2 (N4335, N4311, N1622);
or OR3 (N4336, N4330, N1562, N1261);
buf BUF1 (N4337, N4304);
buf BUF1 (N4338, N4331);
xor XOR2 (N4339, N4338, N98);
xor XOR2 (N4340, N4321, N3714);
nor NOR3 (N4341, N4328, N1072, N4102);
xor XOR2 (N4342, N4319, N1277);
or OR2 (N4343, N4342, N1615);
or OR4 (N4344, N4341, N1292, N3053, N3513);
not NOT1 (N4345, N4344);
and AND3 (N4346, N4345, N2373, N4286);
xor XOR2 (N4347, N4343, N3716);
not NOT1 (N4348, N4346);
not NOT1 (N4349, N4339);
buf BUF1 (N4350, N4333);
and AND2 (N4351, N4347, N1066);
or OR2 (N4352, N4351, N4219);
or OR4 (N4353, N4332, N3320, N3356, N3898);
or OR4 (N4354, N4352, N237, N3043, N63);
or OR3 (N4355, N4350, N1902, N2367);
nor NOR4 (N4356, N4336, N986, N463, N2164);
xor XOR2 (N4357, N4354, N2798);
nand NAND3 (N4358, N4353, N2596, N4049);
buf BUF1 (N4359, N4356);
nand NAND3 (N4360, N4340, N2170, N1293);
nand NAND2 (N4361, N4334, N709);
buf BUF1 (N4362, N4358);
and AND3 (N4363, N4360, N3083, N1652);
and AND4 (N4364, N4363, N3233, N3981, N771);
not NOT1 (N4365, N4361);
nand NAND4 (N4366, N4359, N2042, N1474, N3938);
nand NAND3 (N4367, N4357, N4144, N2373);
nor NOR3 (N4368, N4337, N1236, N1478);
or OR2 (N4369, N4349, N2169);
nand NAND4 (N4370, N4355, N831, N2367, N252);
and AND2 (N4371, N4368, N3344);
xor XOR2 (N4372, N4369, N1899);
xor XOR2 (N4373, N4365, N3317);
nor NOR2 (N4374, N4370, N3013);
xor XOR2 (N4375, N4366, N3623);
nand NAND2 (N4376, N4335, N1010);
buf BUF1 (N4377, N4364);
buf BUF1 (N4378, N4371);
not NOT1 (N4379, N4362);
or OR4 (N4380, N4367, N4132, N2035, N3309);
nand NAND2 (N4381, N4374, N3493);
or OR4 (N4382, N4378, N177, N2268, N2759);
nand NAND2 (N4383, N4379, N341);
xor XOR2 (N4384, N4373, N1871);
xor XOR2 (N4385, N4375, N1390);
not NOT1 (N4386, N4380);
or OR2 (N4387, N4381, N1282);
not NOT1 (N4388, N4377);
xor XOR2 (N4389, N4385, N3844);
not NOT1 (N4390, N4383);
and AND2 (N4391, N4387, N2022);
nor NOR3 (N4392, N4372, N1142, N1142);
buf BUF1 (N4393, N4382);
xor XOR2 (N4394, N4392, N1359);
not NOT1 (N4395, N4390);
and AND4 (N4396, N4386, N3298, N2591, N691);
xor XOR2 (N4397, N4393, N1566);
and AND3 (N4398, N4348, N4380, N352);
nor NOR2 (N4399, N4396, N3627);
buf BUF1 (N4400, N4391);
not NOT1 (N4401, N4400);
and AND2 (N4402, N4384, N1456);
not NOT1 (N4403, N4389);
and AND2 (N4404, N4395, N4094);
xor XOR2 (N4405, N4376, N1347);
and AND4 (N4406, N4405, N3540, N150, N162);
nand NAND3 (N4407, N4403, N1125, N2607);
xor XOR2 (N4408, N4398, N1025);
and AND2 (N4409, N4407, N473);
not NOT1 (N4410, N4406);
not NOT1 (N4411, N4409);
nand NAND3 (N4412, N4399, N3978, N2213);
and AND3 (N4413, N4410, N106, N1260);
buf BUF1 (N4414, N4402);
buf BUF1 (N4415, N4404);
or OR2 (N4416, N4401, N517);
nand NAND4 (N4417, N4414, N291, N2729, N2342);
nand NAND4 (N4418, N4411, N1686, N1085, N843);
buf BUF1 (N4419, N4408);
xor XOR2 (N4420, N4416, N2242);
or OR3 (N4421, N4417, N2320, N3849);
xor XOR2 (N4422, N4413, N2413);
or OR4 (N4423, N4418, N3729, N1268, N4397);
not NOT1 (N4424, N140);
nor NOR2 (N4425, N4394, N2634);
or OR2 (N4426, N4421, N2715);
nor NOR4 (N4427, N4415, N2490, N1023, N2384);
xor XOR2 (N4428, N4419, N2521);
nor NOR3 (N4429, N4420, N3474, N2967);
buf BUF1 (N4430, N4424);
buf BUF1 (N4431, N4422);
and AND4 (N4432, N4388, N2332, N1689, N1292);
buf BUF1 (N4433, N4431);
nor NOR3 (N4434, N4430, N2821, N2121);
and AND2 (N4435, N4434, N2217);
nand NAND4 (N4436, N4426, N2861, N1407, N1008);
and AND2 (N4437, N4435, N2549);
not NOT1 (N4438, N4432);
xor XOR2 (N4439, N4436, N3053);
not NOT1 (N4440, N4412);
xor XOR2 (N4441, N4433, N4321);
not NOT1 (N4442, N4423);
nand NAND4 (N4443, N4438, N3375, N2328, N1698);
or OR3 (N4444, N4437, N1986, N2044);
or OR3 (N4445, N4440, N1202, N3311);
buf BUF1 (N4446, N4441);
xor XOR2 (N4447, N4445, N870);
xor XOR2 (N4448, N4442, N1955);
xor XOR2 (N4449, N4439, N2040);
buf BUF1 (N4450, N4443);
nand NAND3 (N4451, N4427, N1913, N2813);
not NOT1 (N4452, N4447);
xor XOR2 (N4453, N4425, N223);
xor XOR2 (N4454, N4450, N3246);
or OR2 (N4455, N4454, N1591);
buf BUF1 (N4456, N4428);
nor NOR4 (N4457, N4429, N4059, N3444, N859);
and AND2 (N4458, N4457, N709);
nor NOR4 (N4459, N4452, N3815, N3443, N2300);
xor XOR2 (N4460, N4444, N1732);
nand NAND3 (N4461, N4449, N2314, N532);
or OR4 (N4462, N4448, N2371, N3103, N33);
nor NOR3 (N4463, N4453, N3694, N281);
nand NAND4 (N4464, N4462, N2480, N4200, N1375);
not NOT1 (N4465, N4456);
xor XOR2 (N4466, N4455, N1167);
xor XOR2 (N4467, N4451, N1032);
and AND4 (N4468, N4459, N282, N1093, N2959);
xor XOR2 (N4469, N4460, N4390);
not NOT1 (N4470, N4463);
or OR3 (N4471, N4466, N3053, N1722);
or OR3 (N4472, N4470, N3027, N643);
nor NOR2 (N4473, N4472, N1824);
nand NAND4 (N4474, N4467, N3470, N1124, N1562);
not NOT1 (N4475, N4458);
or OR4 (N4476, N4468, N3378, N2287, N2185);
nand NAND4 (N4477, N4465, N2238, N1497, N3857);
xor XOR2 (N4478, N4446, N44);
buf BUF1 (N4479, N4475);
or OR3 (N4480, N4473, N1245, N4117);
nor NOR4 (N4481, N4461, N576, N2372, N4302);
not NOT1 (N4482, N4471);
buf BUF1 (N4483, N4480);
and AND3 (N4484, N4469, N4094, N631);
nor NOR4 (N4485, N4484, N2176, N206, N879);
or OR2 (N4486, N4474, N509);
and AND3 (N4487, N4485, N541, N324);
nand NAND4 (N4488, N4482, N3976, N3749, N1225);
not NOT1 (N4489, N4479);
nand NAND3 (N4490, N4483, N4324, N3828);
xor XOR2 (N4491, N4489, N2933);
or OR4 (N4492, N4491, N534, N902, N1071);
xor XOR2 (N4493, N4476, N3527);
nor NOR4 (N4494, N4492, N3661, N1507, N552);
and AND4 (N4495, N4490, N1677, N3924, N1997);
or OR4 (N4496, N4481, N378, N2062, N1756);
nand NAND4 (N4497, N4477, N2821, N1595, N1055);
not NOT1 (N4498, N4486);
not NOT1 (N4499, N4494);
and AND2 (N4500, N4464, N2387);
or OR2 (N4501, N4495, N369);
xor XOR2 (N4502, N4501, N4320);
and AND3 (N4503, N4502, N1196, N1467);
xor XOR2 (N4504, N4503, N19);
nand NAND4 (N4505, N4500, N3738, N43, N1417);
xor XOR2 (N4506, N4488, N2438);
not NOT1 (N4507, N4493);
and AND3 (N4508, N4504, N1570, N3686);
nor NOR3 (N4509, N4478, N987, N2548);
nand NAND4 (N4510, N4508, N209, N3317, N4040);
nand NAND2 (N4511, N4497, N2383);
or OR4 (N4512, N4496, N668, N1440, N1302);
buf BUF1 (N4513, N4506);
nor NOR3 (N4514, N4498, N864, N727);
not NOT1 (N4515, N4512);
and AND4 (N4516, N4505, N3739, N2213, N3100);
xor XOR2 (N4517, N4499, N1894);
xor XOR2 (N4518, N4515, N3584);
xor XOR2 (N4519, N4517, N3454);
buf BUF1 (N4520, N4509);
not NOT1 (N4521, N4516);
buf BUF1 (N4522, N4487);
xor XOR2 (N4523, N4519, N2386);
not NOT1 (N4524, N4514);
buf BUF1 (N4525, N4521);
and AND3 (N4526, N4525, N3772, N331);
and AND4 (N4527, N4507, N70, N1851, N2999);
nand NAND2 (N4528, N4527, N213);
not NOT1 (N4529, N4511);
nor NOR2 (N4530, N4523, N4064);
nand NAND2 (N4531, N4520, N1451);
nor NOR2 (N4532, N4531, N1027);
and AND4 (N4533, N4526, N3884, N1612, N2019);
buf BUF1 (N4534, N4524);
nor NOR2 (N4535, N4510, N2970);
and AND2 (N4536, N4535, N3662);
not NOT1 (N4537, N4518);
xor XOR2 (N4538, N4536, N462);
or OR3 (N4539, N4529, N603, N427);
xor XOR2 (N4540, N4530, N3429);
or OR4 (N4541, N4513, N3949, N1960, N3550);
not NOT1 (N4542, N4534);
not NOT1 (N4543, N4538);
nand NAND2 (N4544, N4537, N2652);
and AND4 (N4545, N4528, N942, N1963, N1636);
buf BUF1 (N4546, N4544);
buf BUF1 (N4547, N4545);
nor NOR3 (N4548, N4532, N4075, N3835);
xor XOR2 (N4549, N4547, N1243);
xor XOR2 (N4550, N4548, N2395);
xor XOR2 (N4551, N4542, N3365);
xor XOR2 (N4552, N4551, N942);
not NOT1 (N4553, N4541);
nor NOR4 (N4554, N4539, N4230, N1863, N434);
nand NAND3 (N4555, N4554, N929, N2844);
and AND3 (N4556, N4546, N4092, N1569);
buf BUF1 (N4557, N4556);
not NOT1 (N4558, N4553);
xor XOR2 (N4559, N4550, N635);
and AND4 (N4560, N4559, N3030, N1132, N2527);
or OR4 (N4561, N4533, N969, N3308, N787);
not NOT1 (N4562, N4543);
not NOT1 (N4563, N4552);
not NOT1 (N4564, N4563);
and AND3 (N4565, N4557, N848, N2708);
nand NAND2 (N4566, N4565, N3312);
buf BUF1 (N4567, N4549);
nand NAND4 (N4568, N4561, N4397, N1709, N347);
not NOT1 (N4569, N4560);
or OR3 (N4570, N4566, N4433, N1569);
xor XOR2 (N4571, N4569, N567);
buf BUF1 (N4572, N4540);
not NOT1 (N4573, N4567);
buf BUF1 (N4574, N4572);
xor XOR2 (N4575, N4564, N1455);
nor NOR2 (N4576, N4571, N726);
nor NOR2 (N4577, N4555, N3448);
nor NOR3 (N4578, N4522, N3819, N3446);
buf BUF1 (N4579, N4578);
and AND4 (N4580, N4562, N1856, N580, N4334);
or OR2 (N4581, N4577, N1191);
nor NOR3 (N4582, N4574, N439, N1155);
nand NAND3 (N4583, N4576, N1131, N189);
buf BUF1 (N4584, N4579);
or OR2 (N4585, N4584, N1149);
xor XOR2 (N4586, N4570, N3137);
not NOT1 (N4587, N4580);
or OR2 (N4588, N4581, N339);
xor XOR2 (N4589, N4558, N3321);
buf BUF1 (N4590, N4585);
or OR2 (N4591, N4568, N2980);
nand NAND2 (N4592, N4591, N272);
or OR4 (N4593, N4587, N2795, N3085, N1921);
nand NAND2 (N4594, N4590, N3854);
and AND2 (N4595, N4588, N1821);
and AND2 (N4596, N4583, N3547);
xor XOR2 (N4597, N4596, N3812);
not NOT1 (N4598, N4593);
nor NOR4 (N4599, N4573, N199, N2785, N4301);
xor XOR2 (N4600, N4589, N3299);
and AND4 (N4601, N4594, N727, N3382, N793);
and AND4 (N4602, N4600, N39, N1882, N2898);
not NOT1 (N4603, N4601);
or OR3 (N4604, N4597, N3944, N713);
nand NAND4 (N4605, N4592, N2631, N2052, N624);
xor XOR2 (N4606, N4575, N2349);
and AND4 (N4607, N4595, N2730, N3513, N344);
nand NAND4 (N4608, N4602, N4580, N151, N3860);
xor XOR2 (N4609, N4603, N2486);
xor XOR2 (N4610, N4582, N1655);
buf BUF1 (N4611, N4607);
nand NAND2 (N4612, N4606, N4327);
nand NAND2 (N4613, N4611, N1442);
xor XOR2 (N4614, N4610, N1673);
nand NAND3 (N4615, N4586, N792, N1435);
and AND2 (N4616, N4605, N1245);
and AND2 (N4617, N4614, N3369);
xor XOR2 (N4618, N4616, N203);
xor XOR2 (N4619, N4613, N1413);
or OR4 (N4620, N4604, N3329, N1508, N3098);
or OR3 (N4621, N4598, N3098, N715);
and AND3 (N4622, N4612, N1608, N4568);
not NOT1 (N4623, N4618);
nor NOR3 (N4624, N4615, N2889, N544);
nand NAND4 (N4625, N4621, N3953, N1185, N4427);
and AND3 (N4626, N4624, N2791, N2235);
xor XOR2 (N4627, N4626, N2058);
nand NAND2 (N4628, N4620, N3554);
not NOT1 (N4629, N4627);
not NOT1 (N4630, N4619);
nor NOR3 (N4631, N4617, N2185, N1931);
or OR3 (N4632, N4628, N2676, N2442);
xor XOR2 (N4633, N4609, N1108);
nand NAND3 (N4634, N4608, N730, N1564);
and AND4 (N4635, N4629, N328, N689, N2354);
xor XOR2 (N4636, N4633, N3919);
nand NAND2 (N4637, N4599, N1636);
not NOT1 (N4638, N4636);
and AND2 (N4639, N4630, N1768);
not NOT1 (N4640, N4637);
nand NAND4 (N4641, N4623, N1245, N3682, N4231);
xor XOR2 (N4642, N4622, N862);
or OR3 (N4643, N4642, N907, N2171);
or OR2 (N4644, N4638, N1884);
nor NOR2 (N4645, N4634, N4224);
and AND4 (N4646, N4625, N4282, N697, N2813);
or OR3 (N4647, N4645, N719, N1510);
nand NAND3 (N4648, N4635, N3422, N3899);
and AND4 (N4649, N4639, N2954, N3915, N2265);
nor NOR3 (N4650, N4643, N175, N310);
not NOT1 (N4651, N4640);
nor NOR3 (N4652, N4631, N1867, N1699);
not NOT1 (N4653, N4648);
or OR3 (N4654, N4652, N1866, N2925);
nor NOR3 (N4655, N4646, N387, N20);
or OR3 (N4656, N4650, N109, N1208);
and AND2 (N4657, N4649, N1498);
and AND2 (N4658, N4641, N1687);
nand NAND4 (N4659, N4653, N3424, N2153, N1789);
or OR2 (N4660, N4647, N2639);
not NOT1 (N4661, N4659);
nand NAND4 (N4662, N4661, N769, N4151, N4095);
buf BUF1 (N4663, N4644);
nor NOR4 (N4664, N4656, N3206, N4425, N2777);
xor XOR2 (N4665, N4654, N1700);
xor XOR2 (N4666, N4664, N2977);
buf BUF1 (N4667, N4658);
and AND3 (N4668, N4662, N438, N245);
nand NAND2 (N4669, N4668, N3020);
nand NAND2 (N4670, N4655, N1997);
nor NOR4 (N4671, N4666, N1461, N2703, N3649);
xor XOR2 (N4672, N4651, N2134);
buf BUF1 (N4673, N4672);
xor XOR2 (N4674, N4670, N385);
buf BUF1 (N4675, N4632);
not NOT1 (N4676, N4669);
not NOT1 (N4677, N4667);
not NOT1 (N4678, N4677);
and AND3 (N4679, N4673, N1092, N4568);
nand NAND2 (N4680, N4674, N542);
and AND3 (N4681, N4679, N421, N1661);
buf BUF1 (N4682, N4676);
and AND2 (N4683, N4665, N2252);
or OR3 (N4684, N4680, N34, N2238);
not NOT1 (N4685, N4663);
or OR4 (N4686, N4681, N4094, N232, N1231);
nor NOR4 (N4687, N4675, N3491, N3496, N3507);
and AND4 (N4688, N4682, N2181, N659, N2427);
not NOT1 (N4689, N4687);
not NOT1 (N4690, N4671);
not NOT1 (N4691, N4660);
or OR2 (N4692, N4683, N3903);
and AND3 (N4693, N4686, N1666, N1705);
buf BUF1 (N4694, N4690);
nand NAND4 (N4695, N4691, N642, N1434, N782);
nand NAND3 (N4696, N4693, N2528, N4450);
nand NAND3 (N4697, N4678, N1837, N1815);
or OR4 (N4698, N4685, N1240, N739, N2617);
not NOT1 (N4699, N4688);
buf BUF1 (N4700, N4698);
not NOT1 (N4701, N4692);
nand NAND2 (N4702, N4657, N3180);
nand NAND3 (N4703, N4689, N4470, N1462);
xor XOR2 (N4704, N4700, N658);
nor NOR3 (N4705, N4697, N2211, N4059);
or OR4 (N4706, N4694, N3741, N3703, N827);
nor NOR4 (N4707, N4684, N2840, N3582, N4483);
and AND3 (N4708, N4702, N1381, N769);
xor XOR2 (N4709, N4703, N2336);
not NOT1 (N4710, N4699);
not NOT1 (N4711, N4705);
not NOT1 (N4712, N4710);
xor XOR2 (N4713, N4708, N1466);
nand NAND2 (N4714, N4712, N2405);
not NOT1 (N4715, N4714);
and AND3 (N4716, N4696, N2773, N215);
nor NOR3 (N4717, N4711, N2873, N2013);
nand NAND2 (N4718, N4706, N3378);
buf BUF1 (N4719, N4718);
or OR3 (N4720, N4709, N4531, N1054);
xor XOR2 (N4721, N4707, N1087);
nand NAND2 (N4722, N4721, N4686);
buf BUF1 (N4723, N4720);
xor XOR2 (N4724, N4717, N2370);
nor NOR2 (N4725, N4723, N2942);
nand NAND2 (N4726, N4713, N4235);
not NOT1 (N4727, N4716);
nand NAND3 (N4728, N4724, N2762, N463);
and AND2 (N4729, N4725, N839);
nor NOR4 (N4730, N4727, N576, N3121, N3146);
not NOT1 (N4731, N4726);
or OR2 (N4732, N4715, N1331);
or OR4 (N4733, N4701, N4030, N3897, N3231);
and AND3 (N4734, N4733, N2993, N1670);
xor XOR2 (N4735, N4732, N1600);
and AND3 (N4736, N4730, N1779, N2138);
xor XOR2 (N4737, N4722, N3058);
or OR2 (N4738, N4728, N4102);
nor NOR4 (N4739, N4695, N2582, N2980, N2933);
xor XOR2 (N4740, N4734, N4486);
or OR3 (N4741, N4737, N1945, N2114);
nand NAND3 (N4742, N4729, N256, N2259);
not NOT1 (N4743, N4740);
buf BUF1 (N4744, N4735);
nand NAND3 (N4745, N4744, N3714, N2670);
nor NOR2 (N4746, N4739, N1045);
or OR3 (N4747, N4745, N603, N862);
and AND2 (N4748, N4719, N237);
and AND3 (N4749, N4748, N181, N2242);
or OR2 (N4750, N4741, N2469);
or OR3 (N4751, N4747, N1986, N4450);
xor XOR2 (N4752, N4731, N121);
and AND3 (N4753, N4742, N57, N1382);
buf BUF1 (N4754, N4738);
and AND2 (N4755, N4743, N3811);
xor XOR2 (N4756, N4752, N3284);
not NOT1 (N4757, N4704);
xor XOR2 (N4758, N4749, N4550);
or OR2 (N4759, N4750, N3984);
and AND2 (N4760, N4758, N3024);
not NOT1 (N4761, N4755);
nand NAND2 (N4762, N4759, N1216);
or OR4 (N4763, N4746, N3051, N4415, N4100);
xor XOR2 (N4764, N4754, N708);
buf BUF1 (N4765, N4757);
and AND3 (N4766, N4765, N3717, N1562);
buf BUF1 (N4767, N4751);
and AND4 (N4768, N4761, N4571, N4177, N1916);
nand NAND4 (N4769, N4767, N1319, N2612, N1567);
buf BUF1 (N4770, N4768);
not NOT1 (N4771, N4769);
xor XOR2 (N4772, N4764, N1926);
not NOT1 (N4773, N4772);
nor NOR3 (N4774, N4753, N3225, N1035);
nand NAND4 (N4775, N4773, N2525, N1708, N1657);
and AND4 (N4776, N4766, N650, N2296, N4570);
nand NAND4 (N4777, N4770, N2678, N1573, N3752);
or OR2 (N4778, N4777, N1201);
nor NOR4 (N4779, N4762, N1002, N3651, N3751);
nor NOR2 (N4780, N4760, N2731);
nor NOR4 (N4781, N4778, N1055, N2441, N3239);
xor XOR2 (N4782, N4781, N4378);
not NOT1 (N4783, N4763);
xor XOR2 (N4784, N4774, N3843);
xor XOR2 (N4785, N4779, N3800);
not NOT1 (N4786, N4775);
or OR4 (N4787, N4736, N3155, N2806, N332);
or OR3 (N4788, N4783, N307, N2509);
and AND3 (N4789, N4784, N4464, N4113);
not NOT1 (N4790, N4771);
or OR3 (N4791, N4789, N4379, N909);
and AND2 (N4792, N4776, N918);
nor NOR3 (N4793, N4792, N380, N2712);
and AND3 (N4794, N4790, N1883, N2364);
xor XOR2 (N4795, N4780, N4003);
not NOT1 (N4796, N4786);
buf BUF1 (N4797, N4791);
xor XOR2 (N4798, N4787, N4193);
nor NOR4 (N4799, N4798, N2840, N1355, N2774);
not NOT1 (N4800, N4794);
not NOT1 (N4801, N4756);
xor XOR2 (N4802, N4785, N3025);
and AND2 (N4803, N4795, N2210);
buf BUF1 (N4804, N4788);
xor XOR2 (N4805, N4797, N132);
and AND4 (N4806, N4793, N3882, N1907, N4198);
buf BUF1 (N4807, N4800);
nand NAND4 (N4808, N4782, N2175, N4178, N146);
nor NOR3 (N4809, N4803, N2735, N635);
or OR3 (N4810, N4799, N1812, N4346);
nand NAND3 (N4811, N4804, N884, N4704);
buf BUF1 (N4812, N4796);
and AND3 (N4813, N4801, N876, N3268);
and AND3 (N4814, N4806, N1342, N1614);
or OR3 (N4815, N4807, N769, N4498);
and AND4 (N4816, N4810, N1106, N4062, N3708);
or OR3 (N4817, N4814, N1473, N2980);
not NOT1 (N4818, N4802);
not NOT1 (N4819, N4815);
buf BUF1 (N4820, N4816);
nand NAND2 (N4821, N4805, N609);
and AND2 (N4822, N4813, N196);
not NOT1 (N4823, N4809);
nand NAND2 (N4824, N4821, N3014);
not NOT1 (N4825, N4812);
not NOT1 (N4826, N4825);
buf BUF1 (N4827, N4822);
or OR3 (N4828, N4818, N4713, N1373);
or OR3 (N4829, N4828, N3504, N2840);
and AND4 (N4830, N4826, N1324, N2426, N3407);
and AND2 (N4831, N4817, N4152);
not NOT1 (N4832, N4808);
or OR4 (N4833, N4829, N3245, N238, N963);
not NOT1 (N4834, N4827);
or OR2 (N4835, N4832, N4020);
buf BUF1 (N4836, N4830);
nor NOR2 (N4837, N4823, N3716);
or OR2 (N4838, N4834, N1620);
xor XOR2 (N4839, N4811, N2935);
xor XOR2 (N4840, N4839, N510);
not NOT1 (N4841, N4831);
xor XOR2 (N4842, N4841, N1241);
xor XOR2 (N4843, N4837, N1368);
and AND3 (N4844, N4836, N3813, N4352);
nor NOR3 (N4845, N4819, N655, N2251);
or OR4 (N4846, N4842, N2293, N4791, N130);
nor NOR2 (N4847, N4844, N1802);
nand NAND4 (N4848, N4835, N4246, N556, N1487);
not NOT1 (N4849, N4847);
buf BUF1 (N4850, N4824);
and AND2 (N4851, N4838, N1196);
nor NOR4 (N4852, N4820, N692, N3711, N850);
and AND2 (N4853, N4840, N3326);
buf BUF1 (N4854, N4843);
nor NOR4 (N4855, N4848, N2149, N2885, N3677);
nand NAND2 (N4856, N4853, N4639);
buf BUF1 (N4857, N4845);
and AND3 (N4858, N4857, N1420, N964);
buf BUF1 (N4859, N4854);
or OR2 (N4860, N4858, N726);
nand NAND2 (N4861, N4846, N2480);
buf BUF1 (N4862, N4851);
nor NOR4 (N4863, N4862, N1217, N3381, N2921);
nor NOR3 (N4864, N4850, N1348, N4819);
buf BUF1 (N4865, N4852);
and AND4 (N4866, N4861, N2482, N23, N1417);
not NOT1 (N4867, N4855);
and AND4 (N4868, N4860, N4569, N4189, N4494);
not NOT1 (N4869, N4864);
not NOT1 (N4870, N4833);
nand NAND2 (N4871, N4849, N3255);
buf BUF1 (N4872, N4865);
not NOT1 (N4873, N4856);
not NOT1 (N4874, N4871);
nor NOR2 (N4875, N4873, N2324);
and AND4 (N4876, N4870, N4391, N4315, N2859);
not NOT1 (N4877, N4867);
not NOT1 (N4878, N4863);
xor XOR2 (N4879, N4869, N215);
buf BUF1 (N4880, N4874);
buf BUF1 (N4881, N4876);
or OR4 (N4882, N4868, N81, N2980, N2146);
not NOT1 (N4883, N4877);
buf BUF1 (N4884, N4880);
nand NAND3 (N4885, N4883, N3190, N2672);
not NOT1 (N4886, N4878);
nor NOR4 (N4887, N4885, N4065, N2494, N3438);
nor NOR3 (N4888, N4887, N965, N1661);
not NOT1 (N4889, N4888);
xor XOR2 (N4890, N4889, N4240);
nand NAND4 (N4891, N4879, N3417, N4658, N1775);
buf BUF1 (N4892, N4891);
buf BUF1 (N4893, N4890);
not NOT1 (N4894, N4875);
not NOT1 (N4895, N4894);
nand NAND2 (N4896, N4884, N2905);
nor NOR2 (N4897, N4886, N4281);
nand NAND4 (N4898, N4896, N3802, N2577, N4571);
not NOT1 (N4899, N4898);
not NOT1 (N4900, N4866);
xor XOR2 (N4901, N4892, N1688);
nand NAND3 (N4902, N4859, N709, N110);
nand NAND4 (N4903, N4899, N4456, N4173, N2970);
not NOT1 (N4904, N4901);
buf BUF1 (N4905, N4872);
not NOT1 (N4906, N4881);
buf BUF1 (N4907, N4902);
or OR2 (N4908, N4900, N2947);
xor XOR2 (N4909, N4893, N850);
nand NAND4 (N4910, N4882, N4308, N1810, N2758);
nor NOR3 (N4911, N4897, N1347, N4511);
xor XOR2 (N4912, N4907, N1487);
nand NAND2 (N4913, N4912, N1817);
buf BUF1 (N4914, N4904);
xor XOR2 (N4915, N4909, N926);
buf BUF1 (N4916, N4910);
or OR3 (N4917, N4915, N898, N3327);
or OR2 (N4918, N4913, N2272);
buf BUF1 (N4919, N4918);
xor XOR2 (N4920, N4914, N1490);
buf BUF1 (N4921, N4920);
or OR3 (N4922, N4895, N3987, N3238);
xor XOR2 (N4923, N4911, N1669);
nand NAND3 (N4924, N4916, N1769, N2452);
or OR2 (N4925, N4906, N4842);
buf BUF1 (N4926, N4903);
nor NOR3 (N4927, N4905, N3191, N661);
or OR4 (N4928, N4921, N2461, N4834, N4848);
nor NOR4 (N4929, N4928, N249, N3943, N3131);
nor NOR2 (N4930, N4908, N725);
or OR4 (N4931, N4925, N709, N1087, N1845);
nand NAND2 (N4932, N4923, N1964);
nor NOR2 (N4933, N4930, N4831);
not NOT1 (N4934, N4924);
or OR3 (N4935, N4922, N2370, N4400);
and AND4 (N4936, N4933, N597, N1146, N3436);
nor NOR3 (N4937, N4934, N1306, N2436);
buf BUF1 (N4938, N4937);
not NOT1 (N4939, N4927);
nor NOR2 (N4940, N4931, N3840);
xor XOR2 (N4941, N4917, N1909);
not NOT1 (N4942, N4932);
buf BUF1 (N4943, N4941);
nor NOR2 (N4944, N4935, N255);
and AND3 (N4945, N4940, N66, N4932);
and AND3 (N4946, N4945, N3997, N3920);
nor NOR3 (N4947, N4943, N3450, N1809);
nor NOR2 (N4948, N4919, N189);
and AND4 (N4949, N4938, N1835, N1095, N1802);
nor NOR3 (N4950, N4948, N3631, N1223);
buf BUF1 (N4951, N4950);
nor NOR2 (N4952, N4951, N2316);
xor XOR2 (N4953, N4936, N4653);
nor NOR2 (N4954, N4949, N1340);
nor NOR3 (N4955, N4952, N853, N2779);
buf BUF1 (N4956, N4942);
and AND4 (N4957, N4926, N3692, N2065, N907);
nor NOR2 (N4958, N4929, N1293);
and AND4 (N4959, N4953, N3274, N1624, N1300);
nor NOR4 (N4960, N4946, N2757, N1845, N4909);
nand NAND3 (N4961, N4957, N4681, N2779);
and AND2 (N4962, N4947, N4377);
or OR2 (N4963, N4956, N4492);
nand NAND4 (N4964, N4959, N3183, N1527, N852);
buf BUF1 (N4965, N4954);
xor XOR2 (N4966, N4963, N1897);
nor NOR4 (N4967, N4965, N3148, N1831, N4584);
xor XOR2 (N4968, N4960, N1364);
nand NAND2 (N4969, N4962, N1833);
nor NOR3 (N4970, N4967, N3463, N456);
nor NOR2 (N4971, N4939, N1461);
not NOT1 (N4972, N4968);
or OR3 (N4973, N4964, N3937, N3960);
buf BUF1 (N4974, N4944);
nor NOR3 (N4975, N4970, N4651, N3808);
nand NAND3 (N4976, N4955, N1547, N279);
not NOT1 (N4977, N4971);
xor XOR2 (N4978, N4974, N2661);
nor NOR3 (N4979, N4976, N3926, N2765);
nand NAND3 (N4980, N4977, N3021, N1247);
xor XOR2 (N4981, N4978, N1406);
xor XOR2 (N4982, N4979, N1697);
and AND2 (N4983, N4958, N1102);
xor XOR2 (N4984, N4983, N473);
and AND2 (N4985, N4980, N4647);
nand NAND2 (N4986, N4961, N4538);
or OR4 (N4987, N4982, N1113, N2322, N3102);
not NOT1 (N4988, N4966);
nor NOR2 (N4989, N4988, N2511);
or OR4 (N4990, N4987, N961, N4961, N2167);
or OR2 (N4991, N4984, N530);
and AND3 (N4992, N4975, N2089, N4494);
nor NOR3 (N4993, N4985, N4090, N4886);
nand NAND3 (N4994, N4973, N43, N2500);
not NOT1 (N4995, N4994);
xor XOR2 (N4996, N4981, N3276);
xor XOR2 (N4997, N4992, N4169);
buf BUF1 (N4998, N4969);
xor XOR2 (N4999, N4997, N390);
nor NOR2 (N5000, N4995, N837);
and AND4 (N5001, N4993, N1199, N4098, N1758);
nand NAND2 (N5002, N4996, N4476);
nand NAND3 (N5003, N5000, N1659, N3785);
nand NAND2 (N5004, N4990, N1947);
xor XOR2 (N5005, N4998, N2854);
buf BUF1 (N5006, N5002);
xor XOR2 (N5007, N5001, N72);
nor NOR3 (N5008, N4989, N2865, N1914);
and AND2 (N5009, N4972, N4698);
and AND4 (N5010, N5007, N1319, N2192, N2080);
not NOT1 (N5011, N4991);
not NOT1 (N5012, N5010);
nor NOR4 (N5013, N5008, N3737, N2694, N3523);
buf BUF1 (N5014, N4999);
buf BUF1 (N5015, N5009);
nand NAND3 (N5016, N5012, N2044, N1252);
not NOT1 (N5017, N5003);
or OR2 (N5018, N5011, N1045);
and AND4 (N5019, N5017, N204, N533, N2939);
or OR3 (N5020, N5014, N3178, N2308);
not NOT1 (N5021, N5016);
xor XOR2 (N5022, N5015, N2723);
not NOT1 (N5023, N5020);
or OR2 (N5024, N5006, N4351);
or OR2 (N5025, N5004, N1561);
nor NOR2 (N5026, N5019, N1638);
not NOT1 (N5027, N5024);
xor XOR2 (N5028, N5021, N3909);
or OR4 (N5029, N5028, N4141, N698, N3036);
nor NOR4 (N5030, N5026, N3924, N4621, N2914);
not NOT1 (N5031, N5027);
or OR2 (N5032, N5023, N1283);
nand NAND4 (N5033, N4986, N2194, N4825, N1360);
or OR2 (N5034, N5005, N2632);
buf BUF1 (N5035, N5034);
and AND4 (N5036, N5013, N4662, N4016, N220);
or OR2 (N5037, N5033, N70);
xor XOR2 (N5038, N5031, N610);
and AND2 (N5039, N5037, N1235);
or OR3 (N5040, N5038, N1381, N4810);
nand NAND4 (N5041, N5035, N3537, N478, N629);
and AND4 (N5042, N5040, N2434, N4240, N1238);
not NOT1 (N5043, N5029);
not NOT1 (N5044, N5025);
buf BUF1 (N5045, N5041);
and AND2 (N5046, N5018, N1652);
xor XOR2 (N5047, N5045, N1146);
and AND3 (N5048, N5047, N1078, N2840);
or OR3 (N5049, N5042, N4995, N1827);
not NOT1 (N5050, N5044);
not NOT1 (N5051, N5032);
nor NOR2 (N5052, N5050, N694);
and AND3 (N5053, N5039, N135, N1853);
buf BUF1 (N5054, N5030);
and AND3 (N5055, N5046, N604, N508);
nor NOR4 (N5056, N5049, N4846, N624, N4512);
not NOT1 (N5057, N5056);
not NOT1 (N5058, N5055);
not NOT1 (N5059, N5053);
nand NAND4 (N5060, N5051, N1478, N2761, N586);
not NOT1 (N5061, N5059);
buf BUF1 (N5062, N5036);
or OR3 (N5063, N5043, N1294, N5001);
or OR2 (N5064, N5054, N864);
buf BUF1 (N5065, N5022);
or OR3 (N5066, N5052, N676, N513);
nor NOR2 (N5067, N5057, N2636);
and AND2 (N5068, N5061, N2944);
nand NAND2 (N5069, N5064, N2135);
xor XOR2 (N5070, N5068, N1496);
buf BUF1 (N5071, N5062);
and AND3 (N5072, N5063, N2928, N708);
and AND3 (N5073, N5058, N2566, N1707);
nor NOR4 (N5074, N5048, N2238, N4980, N3889);
buf BUF1 (N5075, N5070);
nor NOR4 (N5076, N5065, N2704, N796, N1419);
buf BUF1 (N5077, N5075);
and AND3 (N5078, N5076, N3466, N4122);
xor XOR2 (N5079, N5078, N3312);
or OR3 (N5080, N5077, N4474, N796);
nand NAND4 (N5081, N5074, N4136, N3649, N3159);
and AND3 (N5082, N5080, N1284, N266);
and AND2 (N5083, N5066, N2261);
xor XOR2 (N5084, N5079, N4572);
or OR4 (N5085, N5084, N3836, N3911, N425);
xor XOR2 (N5086, N5083, N3545);
nor NOR4 (N5087, N5081, N5002, N174, N3112);
nor NOR4 (N5088, N5086, N2105, N4320, N633);
nor NOR4 (N5089, N5073, N627, N1042, N1760);
nand NAND4 (N5090, N5089, N5068, N1911, N344);
nor NOR4 (N5091, N5071, N2273, N4263, N4799);
nor NOR2 (N5092, N5067, N4081);
and AND3 (N5093, N5090, N4799, N1020);
or OR3 (N5094, N5069, N5026, N3221);
or OR3 (N5095, N5088, N2948, N2248);
nand NAND2 (N5096, N5072, N2647);
or OR2 (N5097, N5092, N4984);
nand NAND4 (N5098, N5095, N1055, N911, N291);
not NOT1 (N5099, N5060);
buf BUF1 (N5100, N5087);
xor XOR2 (N5101, N5097, N4472);
nand NAND3 (N5102, N5101, N3716, N625);
nand NAND4 (N5103, N5100, N4279, N3561, N3873);
nor NOR2 (N5104, N5096, N2355);
nand NAND2 (N5105, N5082, N2248);
nor NOR3 (N5106, N5094, N2446, N1755);
buf BUF1 (N5107, N5085);
not NOT1 (N5108, N5099);
and AND4 (N5109, N5103, N4043, N254, N2836);
not NOT1 (N5110, N5109);
and AND2 (N5111, N5107, N3307);
xor XOR2 (N5112, N5091, N3427);
nor NOR2 (N5113, N5106, N415);
and AND3 (N5114, N5102, N274, N3691);
nor NOR3 (N5115, N5112, N3902, N1764);
nor NOR4 (N5116, N5114, N1458, N1845, N1620);
not NOT1 (N5117, N5111);
buf BUF1 (N5118, N5117);
nor NOR4 (N5119, N5098, N2119, N2679, N2396);
nor NOR2 (N5120, N5115, N374);
nand NAND4 (N5121, N5118, N2798, N1154, N3641);
and AND2 (N5122, N5105, N2133);
not NOT1 (N5123, N5113);
xor XOR2 (N5124, N5116, N1652);
xor XOR2 (N5125, N5120, N3660);
and AND3 (N5126, N5104, N2718, N3113);
or OR4 (N5127, N5119, N875, N4668, N2045);
nor NOR3 (N5128, N5108, N3475, N3178);
buf BUF1 (N5129, N5093);
xor XOR2 (N5130, N5128, N3712);
nor NOR2 (N5131, N5110, N3937);
buf BUF1 (N5132, N5126);
not NOT1 (N5133, N5132);
or OR3 (N5134, N5129, N1409, N3020);
or OR3 (N5135, N5123, N3413, N4306);
buf BUF1 (N5136, N5122);
or OR4 (N5137, N5131, N4836, N1971, N767);
nand NAND3 (N5138, N5134, N2323, N2917);
nor NOR3 (N5139, N5133, N5130, N3937);
nand NAND3 (N5140, N4945, N2451, N754);
nand NAND3 (N5141, N5127, N1765, N1284);
buf BUF1 (N5142, N5135);
and AND2 (N5143, N5141, N2574);
nand NAND3 (N5144, N5142, N3743, N91);
xor XOR2 (N5145, N5125, N2045);
nor NOR3 (N5146, N5139, N1288, N4869);
and AND2 (N5147, N5143, N1783);
not NOT1 (N5148, N5147);
buf BUF1 (N5149, N5136);
buf BUF1 (N5150, N5121);
and AND3 (N5151, N5138, N2049, N3844);
or OR3 (N5152, N5144, N497, N1185);
and AND2 (N5153, N5152, N1668);
and AND3 (N5154, N5153, N2426, N732);
xor XOR2 (N5155, N5149, N4907);
nor NOR4 (N5156, N5137, N2916, N2437, N2460);
and AND4 (N5157, N5124, N2758, N82, N2281);
buf BUF1 (N5158, N5155);
or OR3 (N5159, N5140, N3248, N2928);
or OR4 (N5160, N5146, N3080, N3345, N3247);
and AND3 (N5161, N5154, N444, N1632);
buf BUF1 (N5162, N5145);
or OR4 (N5163, N5156, N3564, N1867, N1920);
buf BUF1 (N5164, N5158);
xor XOR2 (N5165, N5157, N2035);
or OR4 (N5166, N5163, N1452, N7, N2993);
nor NOR4 (N5167, N5165, N124, N972, N2815);
nor NOR2 (N5168, N5159, N560);
and AND3 (N5169, N5151, N1850, N2632);
nor NOR3 (N5170, N5167, N4313, N663);
xor XOR2 (N5171, N5169, N2252);
xor XOR2 (N5172, N5168, N2131);
or OR3 (N5173, N5172, N424, N2719);
and AND4 (N5174, N5166, N3913, N1126, N3663);
buf BUF1 (N5175, N5173);
and AND2 (N5176, N5160, N2607);
or OR3 (N5177, N5176, N4678, N3160);
buf BUF1 (N5178, N5162);
and AND3 (N5179, N5177, N2904, N47);
or OR3 (N5180, N5171, N3367, N3474);
nand NAND2 (N5181, N5178, N1019);
nor NOR4 (N5182, N5174, N4867, N2711, N2381);
nand NAND2 (N5183, N5150, N4726);
and AND2 (N5184, N5179, N3636);
nand NAND2 (N5185, N5175, N1751);
and AND3 (N5186, N5170, N4581, N3930);
nor NOR2 (N5187, N5181, N3093);
nand NAND4 (N5188, N5148, N1726, N3811, N2127);
not NOT1 (N5189, N5183);
or OR4 (N5190, N5180, N281, N2898, N435);
or OR4 (N5191, N5186, N2536, N2869, N2236);
xor XOR2 (N5192, N5161, N488);
xor XOR2 (N5193, N5184, N3521);
nand NAND3 (N5194, N5185, N86, N3930);
not NOT1 (N5195, N5194);
buf BUF1 (N5196, N5188);
buf BUF1 (N5197, N5164);
nand NAND3 (N5198, N5196, N3810, N3704);
buf BUF1 (N5199, N5182);
or OR3 (N5200, N5195, N5009, N4105);
and AND2 (N5201, N5189, N4067);
buf BUF1 (N5202, N5198);
not NOT1 (N5203, N5199);
nand NAND3 (N5204, N5187, N4978, N3778);
or OR2 (N5205, N5193, N125);
not NOT1 (N5206, N5200);
not NOT1 (N5207, N5203);
nand NAND3 (N5208, N5197, N1708, N2081);
xor XOR2 (N5209, N5208, N895);
nor NOR3 (N5210, N5206, N3588, N321);
and AND4 (N5211, N5205, N2831, N741, N1309);
not NOT1 (N5212, N5191);
and AND3 (N5213, N5192, N1515, N3268);
nand NAND4 (N5214, N5209, N2118, N753, N459);
buf BUF1 (N5215, N5214);
not NOT1 (N5216, N5210);
nor NOR4 (N5217, N5211, N4422, N471, N2747);
xor XOR2 (N5218, N5204, N4161);
or OR2 (N5219, N5216, N1226);
buf BUF1 (N5220, N5219);
or OR4 (N5221, N5213, N538, N1322, N1468);
buf BUF1 (N5222, N5220);
xor XOR2 (N5223, N5190, N4867);
not NOT1 (N5224, N5218);
xor XOR2 (N5225, N5202, N2174);
or OR3 (N5226, N5223, N3891, N2513);
and AND4 (N5227, N5222, N2233, N4472, N3499);
not NOT1 (N5228, N5224);
nor NOR2 (N5229, N5207, N170);
or OR3 (N5230, N5229, N583, N3065);
nand NAND2 (N5231, N5201, N2742);
xor XOR2 (N5232, N5226, N4757);
buf BUF1 (N5233, N5232);
xor XOR2 (N5234, N5217, N1265);
buf BUF1 (N5235, N5215);
xor XOR2 (N5236, N5235, N1070);
nor NOR3 (N5237, N5236, N4116, N3156);
not NOT1 (N5238, N5227);
nor NOR2 (N5239, N5233, N2794);
nor NOR3 (N5240, N5237, N2267, N88);
and AND4 (N5241, N5212, N3116, N5100, N5229);
and AND3 (N5242, N5221, N2253, N2485);
buf BUF1 (N5243, N5234);
xor XOR2 (N5244, N5230, N235);
nor NOR4 (N5245, N5244, N2248, N614, N1834);
and AND3 (N5246, N5242, N2966, N3800);
buf BUF1 (N5247, N5240);
buf BUF1 (N5248, N5239);
and AND2 (N5249, N5243, N3165);
and AND4 (N5250, N5225, N3909, N3665, N590);
and AND4 (N5251, N5241, N3421, N2035, N832);
xor XOR2 (N5252, N5246, N4187);
not NOT1 (N5253, N5247);
xor XOR2 (N5254, N5251, N3140);
nor NOR4 (N5255, N5250, N3446, N3212, N1719);
xor XOR2 (N5256, N5245, N2007);
nand NAND3 (N5257, N5228, N1702, N342);
nand NAND2 (N5258, N5254, N891);
nor NOR4 (N5259, N5256, N1708, N4276, N1953);
not NOT1 (N5260, N5257);
nor NOR2 (N5261, N5249, N3565);
nand NAND2 (N5262, N5260, N1352);
buf BUF1 (N5263, N5259);
nor NOR3 (N5264, N5252, N4877, N4532);
or OR2 (N5265, N5255, N2007);
nand NAND3 (N5266, N5253, N4874, N3391);
xor XOR2 (N5267, N5248, N3284);
buf BUF1 (N5268, N5238);
not NOT1 (N5269, N5267);
buf BUF1 (N5270, N5268);
nand NAND4 (N5271, N5263, N2345, N3994, N4175);
nor NOR4 (N5272, N5270, N4643, N3424, N3619);
xor XOR2 (N5273, N5264, N2562);
nor NOR4 (N5274, N5262, N5057, N3574, N1735);
buf BUF1 (N5275, N5265);
or OR3 (N5276, N5274, N3967, N1909);
nand NAND4 (N5277, N5273, N3879, N2555, N1635);
or OR2 (N5278, N5266, N665);
buf BUF1 (N5279, N5271);
nand NAND2 (N5280, N5276, N1615);
or OR3 (N5281, N5275, N5275, N1130);
nor NOR2 (N5282, N5269, N4431);
nand NAND2 (N5283, N5261, N5035);
or OR3 (N5284, N5231, N4680, N329);
xor XOR2 (N5285, N5284, N4938);
not NOT1 (N5286, N5285);
or OR2 (N5287, N5258, N3343);
and AND4 (N5288, N5283, N3316, N3324, N2927);
and AND3 (N5289, N5281, N4363, N1878);
buf BUF1 (N5290, N5288);
buf BUF1 (N5291, N5280);
nor NOR2 (N5292, N5277, N2292);
not NOT1 (N5293, N5290);
or OR4 (N5294, N5289, N4443, N3039, N463);
or OR2 (N5295, N5272, N1495);
and AND2 (N5296, N5287, N5201);
nor NOR3 (N5297, N5286, N244, N5255);
nor NOR2 (N5298, N5294, N1343);
nand NAND3 (N5299, N5291, N2209, N4536);
nand NAND2 (N5300, N5295, N4577);
nand NAND2 (N5301, N5292, N5192);
nand NAND4 (N5302, N5278, N936, N658, N188);
buf BUF1 (N5303, N5299);
buf BUF1 (N5304, N5279);
nor NOR2 (N5305, N5304, N5082);
nor NOR2 (N5306, N5303, N685);
nor NOR4 (N5307, N5298, N3265, N5, N3460);
buf BUF1 (N5308, N5307);
xor XOR2 (N5309, N5293, N1977);
buf BUF1 (N5310, N5297);
xor XOR2 (N5311, N5308, N5283);
nand NAND2 (N5312, N5282, N408);
buf BUF1 (N5313, N5302);
not NOT1 (N5314, N5312);
xor XOR2 (N5315, N5309, N2538);
buf BUF1 (N5316, N5314);
and AND4 (N5317, N5310, N3628, N2, N1599);
and AND4 (N5318, N5305, N5205, N1452, N4489);
or OR3 (N5319, N5317, N2538, N431);
xor XOR2 (N5320, N5318, N3282);
nand NAND3 (N5321, N5301, N4759, N3776);
not NOT1 (N5322, N5296);
or OR2 (N5323, N5321, N3508);
or OR3 (N5324, N5313, N5081, N3009);
or OR2 (N5325, N5306, N533);
not NOT1 (N5326, N5319);
and AND3 (N5327, N5324, N1903, N1909);
not NOT1 (N5328, N5300);
not NOT1 (N5329, N5328);
nor NOR3 (N5330, N5326, N4835, N1368);
nand NAND2 (N5331, N5316, N3377);
or OR2 (N5332, N5311, N2390);
nor NOR3 (N5333, N5329, N4149, N979);
nor NOR2 (N5334, N5325, N2255);
not NOT1 (N5335, N5332);
nor NOR3 (N5336, N5335, N2027, N3380);
nor NOR3 (N5337, N5327, N1179, N3274);
xor XOR2 (N5338, N5334, N697);
buf BUF1 (N5339, N5331);
nor NOR3 (N5340, N5315, N4100, N2528);
not NOT1 (N5341, N5337);
xor XOR2 (N5342, N5322, N2057);
or OR4 (N5343, N5342, N806, N1865, N3151);
nand NAND4 (N5344, N5339, N2668, N3221, N111);
buf BUF1 (N5345, N5343);
nand NAND4 (N5346, N5341, N4983, N1282, N5223);
nor NOR2 (N5347, N5323, N726);
nor NOR4 (N5348, N5347, N2519, N4203, N1509);
buf BUF1 (N5349, N5336);
not NOT1 (N5350, N5333);
and AND4 (N5351, N5349, N2505, N4142, N3426);
buf BUF1 (N5352, N5350);
nand NAND3 (N5353, N5340, N5271, N1178);
nor NOR4 (N5354, N5351, N1856, N1788, N545);
nor NOR2 (N5355, N5348, N1643);
buf BUF1 (N5356, N5344);
and AND2 (N5357, N5356, N5229);
not NOT1 (N5358, N5352);
and AND2 (N5359, N5330, N1932);
buf BUF1 (N5360, N5354);
buf BUF1 (N5361, N5358);
and AND2 (N5362, N5355, N1006);
xor XOR2 (N5363, N5357, N4712);
not NOT1 (N5364, N5361);
or OR3 (N5365, N5346, N521, N188);
and AND3 (N5366, N5338, N3963, N2318);
or OR2 (N5367, N5360, N246);
xor XOR2 (N5368, N5345, N4712);
nor NOR4 (N5369, N5365, N4106, N356, N4049);
buf BUF1 (N5370, N5359);
xor XOR2 (N5371, N5369, N353);
or OR4 (N5372, N5366, N5346, N1040, N685);
nor NOR4 (N5373, N5353, N4682, N2718, N288);
or OR4 (N5374, N5362, N4795, N1668, N2856);
xor XOR2 (N5375, N5374, N3863);
and AND3 (N5376, N5370, N332, N4479);
nor NOR3 (N5377, N5371, N217, N4808);
nand NAND2 (N5378, N5363, N1065);
and AND2 (N5379, N5320, N3546);
buf BUF1 (N5380, N5364);
xor XOR2 (N5381, N5367, N3184);
or OR3 (N5382, N5380, N5145, N4007);
buf BUF1 (N5383, N5376);
buf BUF1 (N5384, N5368);
nand NAND3 (N5385, N5373, N36, N1912);
nand NAND3 (N5386, N5379, N4822, N2284);
or OR2 (N5387, N5383, N2631);
not NOT1 (N5388, N5382);
or OR3 (N5389, N5387, N1154, N3073);
nand NAND4 (N5390, N5378, N5035, N3014, N3342);
nor NOR3 (N5391, N5375, N2443, N4798);
buf BUF1 (N5392, N5391);
not NOT1 (N5393, N5389);
and AND4 (N5394, N5381, N4652, N4049, N5031);
nor NOR3 (N5395, N5372, N1161, N818);
xor XOR2 (N5396, N5390, N4562);
or OR2 (N5397, N5393, N3087);
buf BUF1 (N5398, N5385);
xor XOR2 (N5399, N5396, N2701);
or OR2 (N5400, N5394, N1859);
or OR4 (N5401, N5386, N1791, N3028, N1015);
xor XOR2 (N5402, N5400, N4755);
nor NOR3 (N5403, N5397, N1276, N4869);
xor XOR2 (N5404, N5402, N1123);
nor NOR4 (N5405, N5404, N1949, N3206, N4578);
xor XOR2 (N5406, N5388, N3236);
nand NAND4 (N5407, N5384, N5097, N4441, N3279);
nor NOR4 (N5408, N5405, N4147, N2200, N2322);
nand NAND4 (N5409, N5395, N5146, N29, N48);
not NOT1 (N5410, N5377);
or OR2 (N5411, N5410, N4055);
not NOT1 (N5412, N5401);
not NOT1 (N5413, N5407);
nor NOR4 (N5414, N5399, N3, N2545, N5181);
nor NOR3 (N5415, N5413, N1931, N3082);
or OR4 (N5416, N5398, N1185, N3591, N5104);
not NOT1 (N5417, N5415);
nor NOR4 (N5418, N5412, N815, N5326, N2996);
or OR2 (N5419, N5418, N3559);
xor XOR2 (N5420, N5411, N5063);
not NOT1 (N5421, N5409);
xor XOR2 (N5422, N5406, N3553);
or OR4 (N5423, N5392, N432, N5328, N2198);
nand NAND3 (N5424, N5420, N4697, N1282);
buf BUF1 (N5425, N5416);
and AND4 (N5426, N5421, N764, N954, N234);
nand NAND3 (N5427, N5426, N1046, N4564);
buf BUF1 (N5428, N5403);
xor XOR2 (N5429, N5427, N1017);
xor XOR2 (N5430, N5414, N3836);
or OR4 (N5431, N5422, N152, N2159, N342);
xor XOR2 (N5432, N5429, N5351);
nor NOR4 (N5433, N5425, N4436, N2889, N3678);
nor NOR2 (N5434, N5431, N4914);
nand NAND4 (N5435, N5424, N3544, N2370, N4571);
and AND2 (N5436, N5430, N25);
not NOT1 (N5437, N5408);
buf BUF1 (N5438, N5435);
or OR4 (N5439, N5417, N1859, N5391, N4254);
not NOT1 (N5440, N5434);
or OR3 (N5441, N5432, N118, N3079);
buf BUF1 (N5442, N5440);
and AND2 (N5443, N5423, N4875);
nor NOR3 (N5444, N5419, N1199, N2322);
nand NAND2 (N5445, N5436, N1551);
nor NOR3 (N5446, N5444, N3633, N4873);
nor NOR3 (N5447, N5441, N168, N3207);
buf BUF1 (N5448, N5439);
not NOT1 (N5449, N5433);
buf BUF1 (N5450, N5442);
not NOT1 (N5451, N5446);
and AND2 (N5452, N5449, N1234);
or OR3 (N5453, N5451, N2057, N5240);
xor XOR2 (N5454, N5443, N2420);
and AND3 (N5455, N5454, N3255, N3249);
and AND3 (N5456, N5453, N2865, N4204);
or OR4 (N5457, N5448, N1964, N4915, N4631);
or OR4 (N5458, N5438, N236, N933, N2318);
xor XOR2 (N5459, N5458, N775);
nor NOR2 (N5460, N5447, N4426);
xor XOR2 (N5461, N5457, N711);
and AND2 (N5462, N5428, N4910);
buf BUF1 (N5463, N5462);
buf BUF1 (N5464, N5452);
and AND2 (N5465, N5456, N1205);
or OR2 (N5466, N5461, N3934);
and AND4 (N5467, N5466, N4897, N2503, N3556);
nand NAND3 (N5468, N5459, N4204, N4861);
and AND3 (N5469, N5463, N2804, N4831);
not NOT1 (N5470, N5467);
not NOT1 (N5471, N5464);
not NOT1 (N5472, N5468);
nand NAND2 (N5473, N5460, N26);
or OR2 (N5474, N5455, N2947);
nand NAND4 (N5475, N5437, N1548, N1212, N3133);
buf BUF1 (N5476, N5471);
nand NAND2 (N5477, N5450, N4875);
or OR2 (N5478, N5477, N2380);
not NOT1 (N5479, N5475);
buf BUF1 (N5480, N5474);
nor NOR4 (N5481, N5469, N982, N3292, N1682);
or OR3 (N5482, N5465, N4999, N5385);
xor XOR2 (N5483, N5478, N3032);
xor XOR2 (N5484, N5480, N3672);
not NOT1 (N5485, N5476);
nor NOR2 (N5486, N5482, N123);
xor XOR2 (N5487, N5483, N402);
or OR2 (N5488, N5470, N3478);
buf BUF1 (N5489, N5481);
buf BUF1 (N5490, N5488);
buf BUF1 (N5491, N5472);
not NOT1 (N5492, N5484);
xor XOR2 (N5493, N5492, N4850);
xor XOR2 (N5494, N5486, N5061);
buf BUF1 (N5495, N5473);
and AND3 (N5496, N5485, N4295, N1482);
xor XOR2 (N5497, N5489, N2123);
not NOT1 (N5498, N5493);
or OR3 (N5499, N5494, N3620, N2271);
or OR3 (N5500, N5487, N2900, N2829);
xor XOR2 (N5501, N5497, N799);
not NOT1 (N5502, N5500);
nand NAND4 (N5503, N5491, N3386, N1171, N4015);
and AND4 (N5504, N5495, N2195, N1931, N573);
and AND4 (N5505, N5503, N3121, N4034, N216);
xor XOR2 (N5506, N5496, N2844);
nand NAND3 (N5507, N5506, N3776, N4257);
buf BUF1 (N5508, N5445);
or OR4 (N5509, N5501, N2544, N4377, N4904);
or OR2 (N5510, N5504, N3918);
or OR2 (N5511, N5507, N3360);
xor XOR2 (N5512, N5510, N411);
or OR2 (N5513, N5490, N1702);
buf BUF1 (N5514, N5498);
nand NAND4 (N5515, N5502, N4971, N5400, N678);
or OR4 (N5516, N5499, N2661, N4323, N3679);
xor XOR2 (N5517, N5512, N3422);
buf BUF1 (N5518, N5517);
and AND3 (N5519, N5511, N357, N1616);
not NOT1 (N5520, N5519);
and AND3 (N5521, N5509, N2096, N3222);
nor NOR4 (N5522, N5521, N3388, N126, N1844);
not NOT1 (N5523, N5518);
nor NOR4 (N5524, N5514, N1059, N4473, N221);
xor XOR2 (N5525, N5479, N1083);
nor NOR3 (N5526, N5505, N1817, N3428);
xor XOR2 (N5527, N5513, N659);
nor NOR2 (N5528, N5527, N3522);
or OR4 (N5529, N5516, N2342, N2304, N5337);
nand NAND3 (N5530, N5525, N1473, N4137);
not NOT1 (N5531, N5528);
and AND3 (N5532, N5524, N4808, N2284);
or OR2 (N5533, N5520, N2080);
buf BUF1 (N5534, N5522);
nand NAND3 (N5535, N5515, N1794, N2796);
or OR2 (N5536, N5535, N5507);
buf BUF1 (N5537, N5536);
nor NOR3 (N5538, N5508, N910, N993);
not NOT1 (N5539, N5531);
buf BUF1 (N5540, N5529);
nand NAND2 (N5541, N5539, N2631);
buf BUF1 (N5542, N5538);
nand NAND4 (N5543, N5532, N5023, N1534, N4134);
buf BUF1 (N5544, N5526);
or OR2 (N5545, N5544, N886);
not NOT1 (N5546, N5545);
not NOT1 (N5547, N5541);
xor XOR2 (N5548, N5546, N2480);
nor NOR4 (N5549, N5547, N2390, N1531, N4557);
not NOT1 (N5550, N5537);
nor NOR4 (N5551, N5530, N1871, N4844, N241);
not NOT1 (N5552, N5542);
and AND4 (N5553, N5551, N4899, N3629, N4850);
and AND3 (N5554, N5552, N4128, N4650);
nand NAND4 (N5555, N5543, N1155, N3643, N5032);
and AND2 (N5556, N5523, N5511);
and AND4 (N5557, N5533, N2825, N1217, N5534);
nor NOR2 (N5558, N651, N3613);
nand NAND4 (N5559, N5548, N3940, N4917, N4051);
or OR3 (N5560, N5556, N3607, N3729);
buf BUF1 (N5561, N5559);
or OR2 (N5562, N5553, N3403);
nand NAND2 (N5563, N5549, N4948);
buf BUF1 (N5564, N5557);
buf BUF1 (N5565, N5558);
not NOT1 (N5566, N5554);
nand NAND3 (N5567, N5562, N1126, N3746);
xor XOR2 (N5568, N5566, N74);
xor XOR2 (N5569, N5563, N3783);
or OR4 (N5570, N5569, N4941, N4023, N4981);
nor NOR4 (N5571, N5555, N105, N3196, N1717);
not NOT1 (N5572, N5571);
buf BUF1 (N5573, N5564);
nor NOR2 (N5574, N5570, N1484);
nand NAND2 (N5575, N5567, N2818);
not NOT1 (N5576, N5560);
xor XOR2 (N5577, N5576, N4622);
nand NAND3 (N5578, N5575, N731, N5531);
or OR3 (N5579, N5578, N2356, N4027);
nor NOR2 (N5580, N5572, N2718);
nor NOR4 (N5581, N5579, N923, N4258, N2632);
or OR4 (N5582, N5581, N4073, N3593, N4583);
nand NAND2 (N5583, N5580, N3639);
and AND3 (N5584, N5577, N406, N3616);
buf BUF1 (N5585, N5582);
or OR3 (N5586, N5573, N3980, N149);
not NOT1 (N5587, N5583);
nand NAND4 (N5588, N5587, N86, N4061, N715);
nor NOR2 (N5589, N5588, N2958);
nand NAND3 (N5590, N5589, N1021, N1346);
buf BUF1 (N5591, N5565);
xor XOR2 (N5592, N5550, N3767);
nand NAND3 (N5593, N5574, N4482, N111);
nand NAND4 (N5594, N5585, N4392, N4765, N4176);
or OR3 (N5595, N5593, N3574, N4947);
nor NOR3 (N5596, N5594, N5590, N3778);
or OR3 (N5597, N3299, N4164, N4851);
xor XOR2 (N5598, N5592, N2664);
or OR4 (N5599, N5595, N2094, N2064, N2647);
xor XOR2 (N5600, N5586, N4283);
or OR4 (N5601, N5584, N1534, N1271, N5135);
not NOT1 (N5602, N5596);
or OR2 (N5603, N5598, N2828);
nor NOR2 (N5604, N5602, N2317);
nand NAND4 (N5605, N5591, N239, N1995, N1596);
not NOT1 (N5606, N5605);
buf BUF1 (N5607, N5599);
and AND3 (N5608, N5561, N5287, N3438);
nor NOR4 (N5609, N5540, N708, N233, N2079);
or OR2 (N5610, N5607, N3908);
nor NOR2 (N5611, N5608, N4518);
buf BUF1 (N5612, N5597);
nor NOR2 (N5613, N5606, N609);
not NOT1 (N5614, N5613);
xor XOR2 (N5615, N5603, N5325);
nand NAND4 (N5616, N5612, N4930, N3967, N3381);
xor XOR2 (N5617, N5614, N1022);
not NOT1 (N5618, N5616);
xor XOR2 (N5619, N5604, N4305);
nor NOR3 (N5620, N5568, N4746, N719);
nor NOR4 (N5621, N5617, N3393, N2930, N5378);
nor NOR3 (N5622, N5601, N1090, N5555);
or OR4 (N5623, N5611, N4026, N567, N4044);
xor XOR2 (N5624, N5619, N2908);
and AND2 (N5625, N5624, N800);
xor XOR2 (N5626, N5620, N4755);
or OR3 (N5627, N5615, N2560, N2425);
or OR3 (N5628, N5623, N1412, N5350);
and AND4 (N5629, N5621, N2920, N4450, N3792);
xor XOR2 (N5630, N5627, N4743);
or OR2 (N5631, N5610, N75);
and AND2 (N5632, N5609, N193);
nor NOR2 (N5633, N5618, N2509);
not NOT1 (N5634, N5622);
nor NOR4 (N5635, N5632, N3053, N4783, N1186);
nand NAND2 (N5636, N5628, N2571);
nand NAND3 (N5637, N5600, N3078, N1012);
not NOT1 (N5638, N5637);
nor NOR4 (N5639, N5630, N3919, N2197, N1331);
not NOT1 (N5640, N5638);
nand NAND2 (N5641, N5636, N3657);
nand NAND4 (N5642, N5631, N1218, N3508, N4007);
nand NAND2 (N5643, N5642, N2887);
not NOT1 (N5644, N5641);
nor NOR3 (N5645, N5634, N4869, N69);
nand NAND3 (N5646, N5639, N4283, N3499);
nand NAND4 (N5647, N5645, N56, N5103, N5002);
and AND2 (N5648, N5626, N1464);
and AND2 (N5649, N5648, N5383);
xor XOR2 (N5650, N5647, N4222);
xor XOR2 (N5651, N5643, N1934);
not NOT1 (N5652, N5635);
buf BUF1 (N5653, N5640);
buf BUF1 (N5654, N5633);
xor XOR2 (N5655, N5653, N5270);
or OR4 (N5656, N5651, N2891, N5242, N1107);
or OR3 (N5657, N5644, N2364, N1644);
and AND2 (N5658, N5646, N4153);
buf BUF1 (N5659, N5657);
xor XOR2 (N5660, N5656, N3015);
nor NOR2 (N5661, N5650, N5124);
or OR4 (N5662, N5625, N5062, N3975, N2357);
nor NOR4 (N5663, N5629, N5191, N491, N3953);
and AND4 (N5664, N5655, N2556, N4031, N2448);
not NOT1 (N5665, N5652);
xor XOR2 (N5666, N5658, N2639);
nand NAND4 (N5667, N5662, N3603, N914, N4595);
nor NOR2 (N5668, N5664, N538);
buf BUF1 (N5669, N5654);
buf BUF1 (N5670, N5666);
buf BUF1 (N5671, N5660);
xor XOR2 (N5672, N5649, N4738);
xor XOR2 (N5673, N5663, N3957);
buf BUF1 (N5674, N5672);
nor NOR2 (N5675, N5665, N685);
or OR2 (N5676, N5661, N3387);
buf BUF1 (N5677, N5669);
nand NAND2 (N5678, N5659, N1568);
not NOT1 (N5679, N5667);
or OR3 (N5680, N5674, N3301, N3175);
nor NOR4 (N5681, N5677, N4632, N5624, N283);
or OR2 (N5682, N5675, N3409);
xor XOR2 (N5683, N5682, N5343);
nand NAND2 (N5684, N5679, N423);
nand NAND4 (N5685, N5670, N5047, N1898, N754);
buf BUF1 (N5686, N5676);
not NOT1 (N5687, N5683);
and AND3 (N5688, N5687, N3866, N3519);
not NOT1 (N5689, N5673);
not NOT1 (N5690, N5688);
buf BUF1 (N5691, N5689);
xor XOR2 (N5692, N5680, N2512);
nand NAND2 (N5693, N5692, N4588);
xor XOR2 (N5694, N5686, N3296);
or OR4 (N5695, N5681, N3307, N3795, N629);
nor NOR2 (N5696, N5691, N3719);
nor NOR2 (N5697, N5694, N4944);
and AND2 (N5698, N5678, N1885);
nand NAND4 (N5699, N5668, N5179, N1053, N3362);
nand NAND2 (N5700, N5690, N4376);
buf BUF1 (N5701, N5693);
not NOT1 (N5702, N5685);
nand NAND3 (N5703, N5698, N5543, N3067);
and AND4 (N5704, N5671, N265, N2394, N2489);
xor XOR2 (N5705, N5697, N2969);
buf BUF1 (N5706, N5700);
nor NOR3 (N5707, N5701, N1361, N2361);
and AND2 (N5708, N5705, N5128);
buf BUF1 (N5709, N5706);
and AND3 (N5710, N5695, N373, N2370);
buf BUF1 (N5711, N5710);
nand NAND3 (N5712, N5709, N488, N1814);
and AND3 (N5713, N5703, N5468, N5050);
buf BUF1 (N5714, N5707);
not NOT1 (N5715, N5696);
nand NAND4 (N5716, N5704, N3662, N5675, N2781);
xor XOR2 (N5717, N5716, N1420);
nor NOR2 (N5718, N5712, N4945);
nor NOR3 (N5719, N5714, N2552, N4576);
nor NOR4 (N5720, N5719, N2188, N4003, N1956);
buf BUF1 (N5721, N5717);
nor NOR4 (N5722, N5699, N4146, N573, N5186);
xor XOR2 (N5723, N5715, N1772);
or OR2 (N5724, N5720, N63);
and AND2 (N5725, N5713, N4981);
buf BUF1 (N5726, N5708);
xor XOR2 (N5727, N5724, N1447);
or OR2 (N5728, N5725, N1501);
nor NOR2 (N5729, N5727, N2982);
nand NAND2 (N5730, N5721, N4607);
nor NOR3 (N5731, N5722, N5367, N2319);
or OR4 (N5732, N5726, N2261, N2750, N1077);
xor XOR2 (N5733, N5684, N3910);
or OR2 (N5734, N5732, N236);
not NOT1 (N5735, N5731);
or OR2 (N5736, N5735, N3430);
or OR4 (N5737, N5723, N1616, N1838, N1056);
nor NOR3 (N5738, N5737, N4453, N4425);
nand NAND2 (N5739, N5729, N187);
nor NOR3 (N5740, N5702, N5045, N3841);
buf BUF1 (N5741, N5728);
or OR3 (N5742, N5718, N3176, N2237);
or OR3 (N5743, N5741, N196, N4359);
or OR2 (N5744, N5740, N5062);
not NOT1 (N5745, N5736);
nor NOR2 (N5746, N5742, N392);
not NOT1 (N5747, N5730);
nor NOR2 (N5748, N5747, N4035);
or OR2 (N5749, N5711, N2940);
buf BUF1 (N5750, N5739);
and AND3 (N5751, N5749, N2064, N1803);
buf BUF1 (N5752, N5738);
nor NOR3 (N5753, N5750, N5371, N2245);
buf BUF1 (N5754, N5734);
or OR4 (N5755, N5733, N3611, N5752, N2475);
nand NAND3 (N5756, N3523, N5722, N1186);
nor NOR4 (N5757, N5756, N5528, N3382, N367);
and AND2 (N5758, N5757, N5209);
and AND2 (N5759, N5753, N600);
buf BUF1 (N5760, N5744);
and AND2 (N5761, N5755, N4429);
nand NAND3 (N5762, N5746, N3288, N294);
nand NAND4 (N5763, N5758, N5272, N1366, N2495);
buf BUF1 (N5764, N5761);
buf BUF1 (N5765, N5760);
or OR2 (N5766, N5765, N598);
not NOT1 (N5767, N5748);
nor NOR3 (N5768, N5762, N3339, N5592);
and AND4 (N5769, N5759, N4560, N868, N3417);
or OR4 (N5770, N5767, N1013, N4969, N5374);
not NOT1 (N5771, N5745);
nand NAND4 (N5772, N5766, N686, N3166, N309);
not NOT1 (N5773, N5754);
nor NOR4 (N5774, N5773, N2004, N5539, N1523);
nor NOR3 (N5775, N5751, N3437, N5118);
nor NOR3 (N5776, N5768, N2954, N1652);
and AND2 (N5777, N5771, N4476);
not NOT1 (N5778, N5770);
not NOT1 (N5779, N5776);
not NOT1 (N5780, N5779);
and AND3 (N5781, N5777, N1960, N2196);
xor XOR2 (N5782, N5743, N3715);
or OR2 (N5783, N5774, N1417);
nand NAND4 (N5784, N5781, N3819, N4530, N334);
buf BUF1 (N5785, N5769);
not NOT1 (N5786, N5785);
nor NOR2 (N5787, N5763, N1569);
or OR2 (N5788, N5786, N1785);
xor XOR2 (N5789, N5784, N5069);
nand NAND2 (N5790, N5778, N746);
and AND2 (N5791, N5782, N236);
and AND2 (N5792, N5764, N1125);
and AND3 (N5793, N5791, N2972, N2037);
or OR3 (N5794, N5793, N2435, N5415);
buf BUF1 (N5795, N5780);
xor XOR2 (N5796, N5775, N4257);
or OR2 (N5797, N5789, N4893);
xor XOR2 (N5798, N5788, N3575);
xor XOR2 (N5799, N5792, N2995);
and AND2 (N5800, N5798, N3207);
and AND4 (N5801, N5783, N2800, N5213, N673);
nand NAND2 (N5802, N5790, N4105);
xor XOR2 (N5803, N5796, N2892);
not NOT1 (N5804, N5799);
nand NAND3 (N5805, N5801, N2659, N1067);
or OR2 (N5806, N5794, N2690);
nand NAND3 (N5807, N5806, N480, N4773);
not NOT1 (N5808, N5805);
nand NAND2 (N5809, N5803, N844);
buf BUF1 (N5810, N5772);
or OR4 (N5811, N5809, N4293, N2352, N1584);
nand NAND3 (N5812, N5804, N5522, N851);
xor XOR2 (N5813, N5812, N4539);
nor NOR2 (N5814, N5797, N88);
or OR2 (N5815, N5808, N2404);
not NOT1 (N5816, N5814);
xor XOR2 (N5817, N5810, N3352);
and AND3 (N5818, N5787, N5561, N3538);
or OR4 (N5819, N5816, N827, N2854, N1737);
not NOT1 (N5820, N5802);
buf BUF1 (N5821, N5813);
or OR4 (N5822, N5800, N4574, N1299, N2606);
nor NOR3 (N5823, N5815, N5059, N2888);
not NOT1 (N5824, N5822);
nand NAND3 (N5825, N5821, N785, N204);
or OR3 (N5826, N5825, N3337, N4966);
buf BUF1 (N5827, N5818);
not NOT1 (N5828, N5827);
and AND3 (N5829, N5828, N1805, N181);
and AND3 (N5830, N5811, N424, N809);
nor NOR4 (N5831, N5820, N2522, N377, N5090);
xor XOR2 (N5832, N5795, N2350);
nand NAND2 (N5833, N5819, N3799);
not NOT1 (N5834, N5833);
nor NOR4 (N5835, N5832, N4100, N748, N4230);
xor XOR2 (N5836, N5834, N2512);
or OR4 (N5837, N5830, N3669, N201, N5644);
not NOT1 (N5838, N5829);
xor XOR2 (N5839, N5823, N4324);
xor XOR2 (N5840, N5826, N5802);
nand NAND3 (N5841, N5835, N2652, N818);
not NOT1 (N5842, N5831);
buf BUF1 (N5843, N5839);
not NOT1 (N5844, N5843);
nand NAND4 (N5845, N5824, N3686, N1653, N5432);
not NOT1 (N5846, N5841);
and AND4 (N5847, N5837, N4966, N607, N1574);
nand NAND3 (N5848, N5807, N4074, N2118);
nand NAND3 (N5849, N5840, N1666, N4630);
nand NAND3 (N5850, N5836, N1351, N4711);
xor XOR2 (N5851, N5847, N485);
and AND2 (N5852, N5838, N2124);
and AND2 (N5853, N5844, N4570);
and AND2 (N5854, N5853, N425);
or OR4 (N5855, N5817, N5194, N4066, N4704);
not NOT1 (N5856, N5850);
not NOT1 (N5857, N5855);
xor XOR2 (N5858, N5848, N1043);
or OR3 (N5859, N5856, N2029, N5663);
and AND2 (N5860, N5859, N3322);
xor XOR2 (N5861, N5857, N1362);
and AND2 (N5862, N5861, N2711);
not NOT1 (N5863, N5842);
and AND3 (N5864, N5862, N2679, N5231);
nor NOR2 (N5865, N5863, N4736);
buf BUF1 (N5866, N5846);
xor XOR2 (N5867, N5854, N3483);
nor NOR4 (N5868, N5864, N5084, N4286, N5203);
nand NAND2 (N5869, N5860, N795);
not NOT1 (N5870, N5865);
buf BUF1 (N5871, N5869);
not NOT1 (N5872, N5871);
buf BUF1 (N5873, N5870);
nand NAND3 (N5874, N5849, N4775, N5284);
or OR2 (N5875, N5868, N2892);
nor NOR2 (N5876, N5852, N977);
xor XOR2 (N5877, N5867, N3625);
xor XOR2 (N5878, N5874, N4242);
and AND3 (N5879, N5866, N511, N4857);
nor NOR3 (N5880, N5845, N2168, N3009);
and AND4 (N5881, N5877, N2681, N676, N4465);
nand NAND4 (N5882, N5880, N3703, N3354, N2722);
or OR3 (N5883, N5875, N105, N1070);
and AND3 (N5884, N5881, N712, N1171);
nand NAND3 (N5885, N5879, N647, N3711);
or OR3 (N5886, N5876, N5311, N1790);
nand NAND2 (N5887, N5885, N3937);
not NOT1 (N5888, N5878);
and AND4 (N5889, N5887, N1341, N5395, N3807);
buf BUF1 (N5890, N5888);
nand NAND4 (N5891, N5886, N919, N2410, N5890);
nand NAND3 (N5892, N4498, N277, N1255);
not NOT1 (N5893, N5892);
not NOT1 (N5894, N5882);
not NOT1 (N5895, N5873);
or OR4 (N5896, N5851, N3832, N3723, N1873);
nand NAND3 (N5897, N5883, N3544, N928);
buf BUF1 (N5898, N5889);
not NOT1 (N5899, N5858);
buf BUF1 (N5900, N5896);
nor NOR3 (N5901, N5900, N5169, N1551);
nor NOR4 (N5902, N5884, N791, N5725, N2828);
xor XOR2 (N5903, N5897, N1414);
nand NAND3 (N5904, N5894, N3387, N5672);
buf BUF1 (N5905, N5898);
nor NOR4 (N5906, N5904, N5788, N609, N1804);
not NOT1 (N5907, N5872);
xor XOR2 (N5908, N5895, N2337);
and AND4 (N5909, N5906, N5595, N2421, N5461);
not NOT1 (N5910, N5891);
xor XOR2 (N5911, N5901, N2726);
nor NOR3 (N5912, N5905, N836, N3653);
or OR3 (N5913, N5908, N1960, N1144);
nor NOR4 (N5914, N5899, N1570, N1372, N1009);
nor NOR2 (N5915, N5909, N5887);
or OR3 (N5916, N5893, N628, N4241);
or OR2 (N5917, N5912, N2752);
and AND4 (N5918, N5917, N4627, N206, N1466);
or OR3 (N5919, N5910, N5608, N1194);
nor NOR2 (N5920, N5913, N1528);
or OR4 (N5921, N5916, N5471, N1370, N5262);
buf BUF1 (N5922, N5915);
not NOT1 (N5923, N5903);
nor NOR4 (N5924, N5918, N1061, N5051, N870);
nor NOR3 (N5925, N5914, N3099, N842);
and AND3 (N5926, N5907, N3431, N4321);
not NOT1 (N5927, N5925);
not NOT1 (N5928, N5911);
xor XOR2 (N5929, N5923, N4351);
and AND3 (N5930, N5919, N47, N1147);
or OR3 (N5931, N5920, N5648, N5247);
nand NAND4 (N5932, N5930, N4916, N1082, N2156);
and AND3 (N5933, N5926, N1126, N5239);
not NOT1 (N5934, N5932);
nor NOR2 (N5935, N5927, N2687);
xor XOR2 (N5936, N5935, N2925);
or OR3 (N5937, N5902, N4550, N4697);
buf BUF1 (N5938, N5922);
buf BUF1 (N5939, N5933);
not NOT1 (N5940, N5924);
buf BUF1 (N5941, N5928);
and AND3 (N5942, N5929, N3717, N3995);
xor XOR2 (N5943, N5942, N1269);
and AND2 (N5944, N5943, N5932);
nand NAND2 (N5945, N5938, N4123);
nand NAND4 (N5946, N5937, N4602, N1959, N3510);
nor NOR2 (N5947, N5934, N4127);
nand NAND3 (N5948, N5921, N4674, N1942);
nor NOR3 (N5949, N5940, N2032, N314);
and AND4 (N5950, N5949, N3703, N1488, N3930);
or OR2 (N5951, N5941, N2153);
buf BUF1 (N5952, N5931);
buf BUF1 (N5953, N5950);
or OR4 (N5954, N5952, N1750, N5814, N5704);
xor XOR2 (N5955, N5947, N764);
and AND4 (N5956, N5939, N5620, N5253, N3260);
xor XOR2 (N5957, N5951, N4615);
xor XOR2 (N5958, N5956, N3319);
nand NAND4 (N5959, N5946, N3582, N2196, N5721);
xor XOR2 (N5960, N5945, N3782);
nor NOR3 (N5961, N5953, N4251, N3982);
and AND3 (N5962, N5959, N2454, N4828);
nor NOR2 (N5963, N5948, N5475);
nand NAND4 (N5964, N5954, N798, N5238, N3137);
not NOT1 (N5965, N5963);
or OR3 (N5966, N5964, N2212, N3940);
and AND2 (N5967, N5960, N4551);
nor NOR4 (N5968, N5944, N2264, N4787, N1954);
xor XOR2 (N5969, N5955, N104);
or OR2 (N5970, N5957, N601);
xor XOR2 (N5971, N5965, N5325);
xor XOR2 (N5972, N5968, N5771);
nand NAND2 (N5973, N5966, N5187);
and AND2 (N5974, N5958, N717);
xor XOR2 (N5975, N5962, N3251);
or OR4 (N5976, N5973, N5881, N4547, N1786);
or OR3 (N5977, N5969, N2003, N5263);
buf BUF1 (N5978, N5936);
buf BUF1 (N5979, N5961);
xor XOR2 (N5980, N5979, N4365);
nor NOR4 (N5981, N5974, N3087, N3615, N3125);
not NOT1 (N5982, N5975);
not NOT1 (N5983, N5982);
or OR4 (N5984, N5972, N102, N3651, N2108);
xor XOR2 (N5985, N5980, N3596);
nand NAND2 (N5986, N5971, N4926);
nor NOR3 (N5987, N5970, N2051, N415);
nand NAND3 (N5988, N5977, N2536, N3242);
and AND2 (N5989, N5987, N5702);
or OR4 (N5990, N5967, N3925, N2174, N325);
or OR3 (N5991, N5984, N466, N3017);
and AND2 (N5992, N5990, N3990);
buf BUF1 (N5993, N5988);
and AND2 (N5994, N5993, N763);
xor XOR2 (N5995, N5978, N891);
and AND4 (N5996, N5989, N4067, N2628, N4838);
buf BUF1 (N5997, N5985);
buf BUF1 (N5998, N5994);
buf BUF1 (N5999, N5997);
and AND4 (N6000, N5992, N2275, N5287, N373);
nand NAND2 (N6001, N5976, N322);
or OR2 (N6002, N6001, N2129);
or OR4 (N6003, N6000, N2600, N4440, N5224);
not NOT1 (N6004, N5986);
nor NOR4 (N6005, N6002, N4865, N3607, N4622);
or OR2 (N6006, N5991, N950);
not NOT1 (N6007, N6005);
buf BUF1 (N6008, N5983);
not NOT1 (N6009, N6007);
not NOT1 (N6010, N5998);
nor NOR2 (N6011, N5996, N3927);
not NOT1 (N6012, N6004);
nand NAND3 (N6013, N6010, N452, N4220);
xor XOR2 (N6014, N6013, N490);
nor NOR3 (N6015, N6008, N1994, N5744);
or OR4 (N6016, N5981, N5627, N1313, N5096);
xor XOR2 (N6017, N6014, N5955);
not NOT1 (N6018, N6006);
xor XOR2 (N6019, N6003, N5176);
buf BUF1 (N6020, N6012);
nand NAND3 (N6021, N6015, N2251, N71);
or OR2 (N6022, N6020, N5456);
buf BUF1 (N6023, N6017);
and AND4 (N6024, N6011, N5977, N3173, N2798);
or OR3 (N6025, N6016, N1519, N1999);
nand NAND3 (N6026, N6019, N3244, N605);
not NOT1 (N6027, N6024);
nor NOR3 (N6028, N6009, N3344, N820);
nor NOR3 (N6029, N6022, N2539, N3378);
not NOT1 (N6030, N6029);
and AND4 (N6031, N6027, N555, N5713, N252);
or OR4 (N6032, N6023, N1150, N5052, N1028);
or OR2 (N6033, N5999, N577);
or OR4 (N6034, N6026, N3255, N2582, N883);
nor NOR4 (N6035, N6028, N2240, N1711, N4854);
nand NAND2 (N6036, N6030, N1141);
not NOT1 (N6037, N6031);
xor XOR2 (N6038, N6037, N5018);
xor XOR2 (N6039, N6036, N7);
buf BUF1 (N6040, N6035);
nand NAND3 (N6041, N6025, N784, N5725);
not NOT1 (N6042, N6021);
not NOT1 (N6043, N6033);
nand NAND3 (N6044, N6043, N4584, N3214);
or OR3 (N6045, N6039, N3561, N6037);
nor NOR2 (N6046, N6041, N5593);
not NOT1 (N6047, N6040);
nand NAND3 (N6048, N6047, N3029, N3284);
or OR4 (N6049, N6048, N1359, N1460, N5423);
or OR2 (N6050, N6042, N4637);
or OR3 (N6051, N6038, N5808, N729);
nor NOR4 (N6052, N6050, N3363, N3361, N664);
buf BUF1 (N6053, N5995);
xor XOR2 (N6054, N6045, N297);
or OR3 (N6055, N6052, N393, N3593);
xor XOR2 (N6056, N6053, N5999);
not NOT1 (N6057, N6054);
nor NOR4 (N6058, N6018, N222, N4145, N694);
nor NOR3 (N6059, N6055, N733, N2935);
xor XOR2 (N6060, N6049, N5857);
buf BUF1 (N6061, N6044);
nor NOR4 (N6062, N6061, N1942, N3585, N964);
or OR4 (N6063, N6060, N2652, N319, N3914);
not NOT1 (N6064, N6056);
and AND2 (N6065, N6058, N676);
and AND4 (N6066, N6046, N3367, N3029, N3884);
not NOT1 (N6067, N6062);
nor NOR4 (N6068, N6065, N825, N5998, N1779);
nor NOR3 (N6069, N6068, N5059, N1363);
nor NOR3 (N6070, N6067, N2241, N2133);
nand NAND4 (N6071, N6066, N223, N1295, N1638);
nand NAND2 (N6072, N6034, N4666);
xor XOR2 (N6073, N6072, N1606);
not NOT1 (N6074, N6073);
xor XOR2 (N6075, N6063, N5581);
xor XOR2 (N6076, N6051, N4427);
or OR4 (N6077, N6070, N3612, N3719, N3657);
or OR3 (N6078, N6069, N2172, N1560);
or OR2 (N6079, N6077, N399);
nor NOR4 (N6080, N6078, N747, N1074, N4553);
nand NAND3 (N6081, N6076, N13, N2548);
or OR4 (N6082, N6081, N3961, N2918, N2555);
buf BUF1 (N6083, N6032);
or OR3 (N6084, N6071, N1339, N5448);
nor NOR3 (N6085, N6074, N52, N84);
and AND3 (N6086, N6057, N4143, N3457);
buf BUF1 (N6087, N6079);
and AND3 (N6088, N6080, N3954, N4376);
buf BUF1 (N6089, N6086);
nand NAND4 (N6090, N6089, N3204, N2013, N763);
and AND2 (N6091, N6084, N4242);
buf BUF1 (N6092, N6064);
nand NAND4 (N6093, N6059, N1343, N1731, N3541);
and AND3 (N6094, N6082, N1668, N3847);
nand NAND2 (N6095, N6083, N352);
and AND2 (N6096, N6087, N2690);
or OR4 (N6097, N6075, N1481, N372, N641);
xor XOR2 (N6098, N6096, N2401);
or OR4 (N6099, N6095, N1010, N2074, N411);
nand NAND4 (N6100, N6090, N3743, N76, N768);
buf BUF1 (N6101, N6098);
buf BUF1 (N6102, N6093);
nand NAND3 (N6103, N6092, N4662, N2517);
not NOT1 (N6104, N6100);
buf BUF1 (N6105, N6091);
nor NOR2 (N6106, N6102, N590);
and AND4 (N6107, N6085, N4868, N2824, N2359);
xor XOR2 (N6108, N6099, N1183);
or OR4 (N6109, N6108, N1067, N2391, N5550);
nand NAND4 (N6110, N6101, N5634, N3602, N4563);
not NOT1 (N6111, N6104);
and AND3 (N6112, N6088, N3386, N2635);
or OR4 (N6113, N6097, N3648, N3092, N3324);
nand NAND3 (N6114, N6113, N825, N4635);
not NOT1 (N6115, N6105);
xor XOR2 (N6116, N6107, N3857);
buf BUF1 (N6117, N6109);
xor XOR2 (N6118, N6094, N5055);
xor XOR2 (N6119, N6111, N430);
buf BUF1 (N6120, N6103);
and AND4 (N6121, N6106, N5803, N1094, N5933);
nor NOR3 (N6122, N6115, N1627, N5026);
nand NAND2 (N6123, N6114, N1543);
nand NAND3 (N6124, N6122, N4531, N2148);
buf BUF1 (N6125, N6120);
or OR3 (N6126, N6125, N2254, N6);
xor XOR2 (N6127, N6116, N5497);
and AND2 (N6128, N6119, N2337);
or OR2 (N6129, N6124, N146);
nand NAND4 (N6130, N6129, N1177, N2870, N4093);
and AND2 (N6131, N6110, N5926);
or OR4 (N6132, N6117, N2352, N373, N2741);
and AND2 (N6133, N6128, N383);
or OR2 (N6134, N6127, N3902);
nand NAND3 (N6135, N6112, N3152, N2856);
and AND3 (N6136, N6132, N582, N2833);
not NOT1 (N6137, N6118);
xor XOR2 (N6138, N6126, N6054);
nand NAND3 (N6139, N6130, N815, N3437);
nand NAND4 (N6140, N6135, N4898, N373, N1629);
or OR4 (N6141, N6140, N1876, N1624, N5099);
and AND3 (N6142, N6134, N3100, N2571);
xor XOR2 (N6143, N6123, N58);
nor NOR4 (N6144, N6136, N4214, N4451, N5393);
xor XOR2 (N6145, N6139, N3701);
xor XOR2 (N6146, N6121, N2645);
and AND4 (N6147, N6141, N5834, N5336, N359);
nand NAND4 (N6148, N6131, N4441, N4899, N1830);
not NOT1 (N6149, N6146);
nor NOR3 (N6150, N6149, N160, N1635);
not NOT1 (N6151, N6137);
and AND4 (N6152, N6148, N2407, N1718, N4353);
or OR4 (N6153, N6152, N3294, N4503, N2107);
not NOT1 (N6154, N6133);
xor XOR2 (N6155, N6138, N4847);
nand NAND4 (N6156, N6143, N784, N1131, N1469);
buf BUF1 (N6157, N6144);
or OR3 (N6158, N6157, N4207, N4534);
buf BUF1 (N6159, N6145);
xor XOR2 (N6160, N6154, N4150);
and AND4 (N6161, N6159, N691, N185, N2626);
not NOT1 (N6162, N6150);
nor NOR2 (N6163, N6153, N5641);
xor XOR2 (N6164, N6160, N5689);
nand NAND4 (N6165, N6156, N3886, N749, N1242);
xor XOR2 (N6166, N6142, N4659);
buf BUF1 (N6167, N6158);
or OR4 (N6168, N6167, N1117, N5922, N2823);
xor XOR2 (N6169, N6161, N4993);
xor XOR2 (N6170, N6147, N322);
or OR4 (N6171, N6169, N2368, N4706, N3377);
or OR4 (N6172, N6164, N597, N3402, N3);
and AND4 (N6173, N6166, N5375, N1317, N5914);
nor NOR3 (N6174, N6151, N364, N1322);
buf BUF1 (N6175, N6170);
nor NOR2 (N6176, N6175, N3796);
or OR4 (N6177, N6176, N5534, N1898, N2655);
not NOT1 (N6178, N6155);
xor XOR2 (N6179, N6178, N49);
xor XOR2 (N6180, N6162, N395);
nand NAND2 (N6181, N6163, N2568);
buf BUF1 (N6182, N6174);
nand NAND3 (N6183, N6177, N3837, N903);
nand NAND4 (N6184, N6168, N1018, N5607, N3768);
or OR3 (N6185, N6173, N212, N839);
buf BUF1 (N6186, N6182);
buf BUF1 (N6187, N6180);
or OR2 (N6188, N6183, N913);
not NOT1 (N6189, N6181);
not NOT1 (N6190, N6184);
buf BUF1 (N6191, N6165);
not NOT1 (N6192, N6185);
not NOT1 (N6193, N6190);
xor XOR2 (N6194, N6191, N4287);
buf BUF1 (N6195, N6171);
and AND4 (N6196, N6194, N5066, N2594, N5741);
nor NOR3 (N6197, N6188, N747, N5690);
not NOT1 (N6198, N6195);
and AND2 (N6199, N6179, N3683);
and AND2 (N6200, N6193, N1113);
or OR3 (N6201, N6192, N5946, N280);
buf BUF1 (N6202, N6201);
nor NOR2 (N6203, N6172, N4612);
nor NOR4 (N6204, N6199, N5049, N3144, N16);
not NOT1 (N6205, N6197);
nor NOR4 (N6206, N6196, N2556, N4759, N5007);
buf BUF1 (N6207, N6204);
and AND4 (N6208, N6206, N4152, N5599, N3077);
buf BUF1 (N6209, N6205);
xor XOR2 (N6210, N6198, N6019);
xor XOR2 (N6211, N6186, N1580);
or OR3 (N6212, N6211, N3142, N3514);
buf BUF1 (N6213, N6189);
nor NOR3 (N6214, N6187, N5499, N5914);
or OR2 (N6215, N6200, N2419);
buf BUF1 (N6216, N6203);
and AND3 (N6217, N6212, N3047, N5930);
buf BUF1 (N6218, N6202);
buf BUF1 (N6219, N6210);
and AND4 (N6220, N6213, N2640, N414, N5729);
nor NOR2 (N6221, N6207, N2954);
buf BUF1 (N6222, N6219);
nand NAND4 (N6223, N6215, N933, N323, N6215);
nor NOR3 (N6224, N6221, N3027, N65);
xor XOR2 (N6225, N6224, N386);
nand NAND3 (N6226, N6214, N2600, N3198);
xor XOR2 (N6227, N6209, N5376);
nand NAND2 (N6228, N6218, N3607);
nand NAND2 (N6229, N6222, N4736);
nor NOR4 (N6230, N6216, N1985, N6135, N2486);
and AND4 (N6231, N6208, N4013, N2565, N1711);
nor NOR2 (N6232, N6223, N390);
or OR3 (N6233, N6229, N1256, N6196);
xor XOR2 (N6234, N6230, N3466);
xor XOR2 (N6235, N6231, N3690);
xor XOR2 (N6236, N6220, N632);
xor XOR2 (N6237, N6217, N856);
not NOT1 (N6238, N6233);
or OR2 (N6239, N6234, N3074);
nor NOR3 (N6240, N6228, N4035, N4398);
xor XOR2 (N6241, N6227, N6083);
nor NOR2 (N6242, N6241, N2744);
not NOT1 (N6243, N6238);
buf BUF1 (N6244, N6232);
nand NAND2 (N6245, N6225, N2768);
and AND2 (N6246, N6236, N1177);
or OR2 (N6247, N6235, N6110);
and AND3 (N6248, N6243, N1941, N1404);
nor NOR2 (N6249, N6237, N3221);
nor NOR3 (N6250, N6240, N2906, N4299);
or OR3 (N6251, N6249, N1221, N4341);
not NOT1 (N6252, N6248);
nand NAND3 (N6253, N6247, N1499, N5207);
xor XOR2 (N6254, N6251, N1924);
nor NOR2 (N6255, N6239, N1591);
or OR3 (N6256, N6253, N1519, N2090);
not NOT1 (N6257, N6255);
nor NOR3 (N6258, N6250, N1499, N3412);
nand NAND2 (N6259, N6226, N6077);
not NOT1 (N6260, N6256);
or OR2 (N6261, N6254, N4412);
nor NOR2 (N6262, N6260, N2631);
nor NOR3 (N6263, N6259, N3807, N886);
nand NAND3 (N6264, N6261, N4129, N3793);
buf BUF1 (N6265, N6244);
or OR4 (N6266, N6245, N3776, N3229, N1384);
nand NAND3 (N6267, N6246, N1600, N1352);
not NOT1 (N6268, N6267);
not NOT1 (N6269, N6266);
xor XOR2 (N6270, N6263, N3286);
and AND2 (N6271, N6268, N3491);
buf BUF1 (N6272, N6270);
nor NOR3 (N6273, N6271, N5360, N6072);
nand NAND4 (N6274, N6258, N9, N5697, N5841);
xor XOR2 (N6275, N6257, N467);
not NOT1 (N6276, N6265);
nand NAND2 (N6277, N6275, N6060);
nor NOR3 (N6278, N6274, N3582, N3908);
xor XOR2 (N6279, N6273, N5980);
nor NOR4 (N6280, N6279, N3112, N2417, N2724);
not NOT1 (N6281, N6272);
and AND3 (N6282, N6264, N1416, N1053);
buf BUF1 (N6283, N6252);
and AND4 (N6284, N6278, N593, N5715, N4876);
nor NOR2 (N6285, N6277, N3534);
nand NAND4 (N6286, N6276, N5028, N4485, N3004);
buf BUF1 (N6287, N6281);
buf BUF1 (N6288, N6280);
nor NOR4 (N6289, N6282, N3202, N2925, N1986);
not NOT1 (N6290, N6242);
not NOT1 (N6291, N6269);
nand NAND2 (N6292, N6287, N4113);
and AND3 (N6293, N6289, N2486, N1857);
nor NOR2 (N6294, N6292, N666);
xor XOR2 (N6295, N6294, N3645);
buf BUF1 (N6296, N6283);
not NOT1 (N6297, N6262);
or OR4 (N6298, N6286, N5151, N3556, N5490);
nor NOR2 (N6299, N6284, N3594);
buf BUF1 (N6300, N6299);
xor XOR2 (N6301, N6288, N2775);
or OR2 (N6302, N6300, N124);
not NOT1 (N6303, N6291);
or OR3 (N6304, N6302, N1941, N3589);
buf BUF1 (N6305, N6297);
buf BUF1 (N6306, N6293);
buf BUF1 (N6307, N6301);
not NOT1 (N6308, N6303);
nor NOR3 (N6309, N6296, N3582, N1477);
buf BUF1 (N6310, N6304);
xor XOR2 (N6311, N6290, N4809);
and AND2 (N6312, N6305, N5823);
buf BUF1 (N6313, N6308);
not NOT1 (N6314, N6311);
buf BUF1 (N6315, N6312);
not NOT1 (N6316, N6315);
nand NAND3 (N6317, N6298, N770, N6192);
buf BUF1 (N6318, N6295);
nor NOR4 (N6319, N6317, N4337, N467, N2544);
not NOT1 (N6320, N6316);
buf BUF1 (N6321, N6310);
buf BUF1 (N6322, N6306);
and AND2 (N6323, N6319, N77);
not NOT1 (N6324, N6320);
and AND3 (N6325, N6324, N925, N2856);
nor NOR4 (N6326, N6318, N5842, N5454, N5854);
and AND4 (N6327, N6325, N5366, N4936, N53);
nor NOR2 (N6328, N6323, N399);
and AND3 (N6329, N6326, N3199, N2091);
nor NOR4 (N6330, N6285, N6208, N3961, N4159);
nor NOR4 (N6331, N6309, N5888, N1001, N5950);
buf BUF1 (N6332, N6322);
buf BUF1 (N6333, N6329);
buf BUF1 (N6334, N6321);
nand NAND4 (N6335, N6313, N4946, N1385, N4746);
nor NOR2 (N6336, N6307, N2656);
not NOT1 (N6337, N6333);
or OR2 (N6338, N6314, N2770);
buf BUF1 (N6339, N6338);
and AND3 (N6340, N6327, N5586, N5616);
not NOT1 (N6341, N6336);
nand NAND4 (N6342, N6330, N5789, N4805, N3369);
and AND2 (N6343, N6335, N1182);
not NOT1 (N6344, N6331);
not NOT1 (N6345, N6332);
nor NOR2 (N6346, N6334, N5491);
nand NAND4 (N6347, N6340, N440, N3290, N2985);
nand NAND2 (N6348, N6342, N2282);
not NOT1 (N6349, N6343);
and AND4 (N6350, N6337, N2471, N2019, N5517);
nor NOR4 (N6351, N6346, N5926, N1758, N4148);
or OR3 (N6352, N6350, N3959, N2923);
or OR3 (N6353, N6349, N5952, N3075);
and AND3 (N6354, N6352, N4882, N421);
and AND4 (N6355, N6328, N5330, N4318, N874);
nand NAND2 (N6356, N6347, N248);
xor XOR2 (N6357, N6344, N3163);
or OR2 (N6358, N6339, N3413);
and AND3 (N6359, N6351, N4291, N211);
nor NOR4 (N6360, N6358, N3029, N1494, N5935);
buf BUF1 (N6361, N6360);
buf BUF1 (N6362, N6348);
nand NAND4 (N6363, N6355, N2401, N878, N6011);
not NOT1 (N6364, N6363);
nand NAND4 (N6365, N6354, N4529, N4657, N2493);
buf BUF1 (N6366, N6353);
nand NAND4 (N6367, N6359, N2607, N5784, N1069);
nand NAND2 (N6368, N6345, N5799);
nor NOR4 (N6369, N6366, N669, N2739, N5215);
buf BUF1 (N6370, N6365);
nor NOR3 (N6371, N6361, N4318, N3245);
and AND4 (N6372, N6368, N962, N4687, N5465);
and AND4 (N6373, N6367, N6304, N4065, N2857);
nor NOR3 (N6374, N6362, N281, N2486);
xor XOR2 (N6375, N6364, N3254);
and AND2 (N6376, N6375, N5621);
or OR3 (N6377, N6356, N1237, N2741);
buf BUF1 (N6378, N6357);
or OR4 (N6379, N6374, N1544, N127, N1489);
buf BUF1 (N6380, N6370);
xor XOR2 (N6381, N6377, N5000);
nand NAND4 (N6382, N6341, N4933, N1912, N3371);
xor XOR2 (N6383, N6373, N958);
buf BUF1 (N6384, N6381);
nor NOR2 (N6385, N6382, N3282);
nand NAND4 (N6386, N6371, N1993, N3123, N1693);
buf BUF1 (N6387, N6376);
and AND3 (N6388, N6387, N3290, N4049);
not NOT1 (N6389, N6369);
or OR2 (N6390, N6383, N4462);
nand NAND3 (N6391, N6372, N1462, N112);
xor XOR2 (N6392, N6391, N4757);
or OR3 (N6393, N6385, N6053, N504);
buf BUF1 (N6394, N6386);
xor XOR2 (N6395, N6388, N2961);
nand NAND3 (N6396, N6389, N1338, N1563);
xor XOR2 (N6397, N6378, N2379);
buf BUF1 (N6398, N6397);
nand NAND3 (N6399, N6392, N4921, N1387);
xor XOR2 (N6400, N6380, N4579);
xor XOR2 (N6401, N6400, N2848);
buf BUF1 (N6402, N6393);
or OR3 (N6403, N6399, N3349, N746);
and AND3 (N6404, N6396, N395, N4362);
and AND3 (N6405, N6384, N2986, N5352);
and AND4 (N6406, N6402, N1567, N2547, N2772);
nand NAND4 (N6407, N6401, N900, N783, N5661);
or OR3 (N6408, N6398, N3269, N3862);
or OR2 (N6409, N6404, N1744);
buf BUF1 (N6410, N6408);
xor XOR2 (N6411, N6395, N2576);
not NOT1 (N6412, N6411);
or OR3 (N6413, N6407, N2234, N6370);
not NOT1 (N6414, N6412);
buf BUF1 (N6415, N6406);
buf BUF1 (N6416, N6379);
buf BUF1 (N6417, N6415);
buf BUF1 (N6418, N6417);
not NOT1 (N6419, N6394);
xor XOR2 (N6420, N6410, N3804);
or OR4 (N6421, N6409, N5121, N3349, N5676);
buf BUF1 (N6422, N6416);
xor XOR2 (N6423, N6421, N5119);
or OR4 (N6424, N6414, N1535, N5320, N4168);
nor NOR4 (N6425, N6418, N2997, N1764, N3730);
and AND2 (N6426, N6423, N1608);
and AND2 (N6427, N6422, N1898);
xor XOR2 (N6428, N6403, N6045);
not NOT1 (N6429, N6419);
buf BUF1 (N6430, N6425);
or OR4 (N6431, N6429, N4153, N3047, N428);
and AND4 (N6432, N6413, N6013, N6216, N570);
and AND2 (N6433, N6420, N6193);
nand NAND4 (N6434, N6390, N1692, N3033, N5135);
or OR2 (N6435, N6428, N894);
xor XOR2 (N6436, N6433, N4057);
buf BUF1 (N6437, N6405);
xor XOR2 (N6438, N6427, N623);
nand NAND3 (N6439, N6431, N3789, N6380);
xor XOR2 (N6440, N6438, N3177);
nor NOR2 (N6441, N6439, N1130);
buf BUF1 (N6442, N6435);
not NOT1 (N6443, N6432);
or OR4 (N6444, N6441, N1174, N1215, N4600);
and AND4 (N6445, N6430, N4148, N3719, N5240);
or OR3 (N6446, N6442, N4359, N1987);
or OR4 (N6447, N6424, N4642, N2514, N2577);
and AND3 (N6448, N6446, N1912, N1216);
xor XOR2 (N6449, N6434, N4033);
not NOT1 (N6450, N6445);
buf BUF1 (N6451, N6449);
xor XOR2 (N6452, N6443, N3876);
nor NOR4 (N6453, N6426, N1671, N5233, N5371);
nor NOR2 (N6454, N6453, N5097);
nand NAND4 (N6455, N6437, N2551, N3421, N11);
nand NAND4 (N6456, N6454, N240, N708, N3187);
xor XOR2 (N6457, N6452, N47);
xor XOR2 (N6458, N6455, N1431);
nand NAND2 (N6459, N6450, N6191);
xor XOR2 (N6460, N6436, N2647);
or OR4 (N6461, N6451, N5095, N84, N1308);
xor XOR2 (N6462, N6458, N3265);
nor NOR4 (N6463, N6457, N6455, N3886, N2512);
nor NOR4 (N6464, N6447, N5933, N3870, N5361);
nor NOR3 (N6465, N6440, N6013, N1745);
not NOT1 (N6466, N6456);
buf BUF1 (N6467, N6462);
not NOT1 (N6468, N6464);
xor XOR2 (N6469, N6466, N3309);
or OR3 (N6470, N6459, N4796, N6129);
nand NAND3 (N6471, N6467, N4653, N6175);
xor XOR2 (N6472, N6444, N4454);
or OR2 (N6473, N6470, N4078);
xor XOR2 (N6474, N6468, N2112);
nor NOR2 (N6475, N6469, N1532);
nor NOR3 (N6476, N6463, N1221, N4412);
or OR4 (N6477, N6476, N3678, N2257, N2985);
not NOT1 (N6478, N6461);
buf BUF1 (N6479, N6475);
buf BUF1 (N6480, N6477);
and AND2 (N6481, N6448, N235);
nor NOR3 (N6482, N6478, N776, N4507);
nand NAND2 (N6483, N6460, N266);
and AND2 (N6484, N6483, N4643);
not NOT1 (N6485, N6471);
not NOT1 (N6486, N6482);
or OR3 (N6487, N6472, N3824, N5397);
and AND3 (N6488, N6484, N1270, N5883);
nand NAND2 (N6489, N6473, N3375);
nand NAND2 (N6490, N6481, N3588);
or OR2 (N6491, N6479, N1555);
nor NOR2 (N6492, N6491, N5507);
or OR3 (N6493, N6485, N5967, N5567);
nand NAND2 (N6494, N6465, N3205);
buf BUF1 (N6495, N6492);
and AND3 (N6496, N6489, N5749, N2843);
nor NOR2 (N6497, N6494, N1298);
or OR2 (N6498, N6488, N5068);
nor NOR3 (N6499, N6498, N4315, N2816);
or OR4 (N6500, N6497, N3488, N591, N6246);
buf BUF1 (N6501, N6493);
nand NAND4 (N6502, N6496, N1649, N4932, N5295);
nand NAND4 (N6503, N6495, N5899, N4908, N458);
and AND4 (N6504, N6480, N450, N6295, N1590);
nor NOR4 (N6505, N6504, N569, N3612, N5839);
or OR3 (N6506, N6490, N6084, N5347);
not NOT1 (N6507, N6487);
and AND3 (N6508, N6502, N1805, N1891);
and AND3 (N6509, N6505, N108, N4315);
nor NOR4 (N6510, N6506, N359, N4844, N5996);
buf BUF1 (N6511, N6507);
not NOT1 (N6512, N6503);
not NOT1 (N6513, N6501);
buf BUF1 (N6514, N6508);
xor XOR2 (N6515, N6513, N3860);
xor XOR2 (N6516, N6474, N1999);
and AND2 (N6517, N6486, N2253);
nor NOR2 (N6518, N6514, N2028);
not NOT1 (N6519, N6515);
nand NAND3 (N6520, N6517, N5169, N3715);
nor NOR3 (N6521, N6520, N5538, N4186);
not NOT1 (N6522, N6516);
and AND4 (N6523, N6512, N2394, N6359, N2403);
nand NAND2 (N6524, N6510, N20);
nor NOR2 (N6525, N6523, N2549);
nor NOR4 (N6526, N6521, N4649, N5692, N5647);
and AND4 (N6527, N6522, N1393, N5667, N1190);
nor NOR2 (N6528, N6519, N833);
nand NAND2 (N6529, N6509, N1546);
not NOT1 (N6530, N6524);
nand NAND4 (N6531, N6527, N2549, N3238, N4798);
and AND3 (N6532, N6529, N3141, N2373);
xor XOR2 (N6533, N6531, N5181);
not NOT1 (N6534, N6530);
not NOT1 (N6535, N6532);
not NOT1 (N6536, N6534);
or OR2 (N6537, N6533, N2248);
nor NOR4 (N6538, N6528, N3530, N5342, N6506);
nand NAND2 (N6539, N6518, N221);
buf BUF1 (N6540, N6499);
xor XOR2 (N6541, N6538, N509);
nor NOR4 (N6542, N6539, N561, N1322, N5046);
nor NOR3 (N6543, N6525, N839, N2538);
not NOT1 (N6544, N6541);
and AND2 (N6545, N6537, N43);
not NOT1 (N6546, N6536);
and AND2 (N6547, N6511, N4616);
nor NOR3 (N6548, N6535, N3945, N5856);
nor NOR4 (N6549, N6526, N5370, N5087, N5309);
buf BUF1 (N6550, N6540);
not NOT1 (N6551, N6545);
or OR2 (N6552, N6547, N3206);
or OR4 (N6553, N6551, N2312, N3502, N2813);
nand NAND4 (N6554, N6544, N748, N1140, N3590);
buf BUF1 (N6555, N6553);
xor XOR2 (N6556, N6555, N3471);
nand NAND2 (N6557, N6542, N5629);
buf BUF1 (N6558, N6549);
and AND2 (N6559, N6552, N2426);
xor XOR2 (N6560, N6500, N2176);
and AND4 (N6561, N6543, N3070, N4396, N3078);
buf BUF1 (N6562, N6546);
buf BUF1 (N6563, N6558);
xor XOR2 (N6564, N6563, N3688);
or OR4 (N6565, N6560, N229, N2897, N4587);
buf BUF1 (N6566, N6562);
buf BUF1 (N6567, N6561);
nor NOR4 (N6568, N6556, N4526, N1493, N5087);
nor NOR3 (N6569, N6567, N5519, N220);
and AND4 (N6570, N6559, N3920, N1466, N4017);
and AND4 (N6571, N6566, N1717, N385, N3251);
buf BUF1 (N6572, N6554);
xor XOR2 (N6573, N6568, N1240);
and AND3 (N6574, N6570, N338, N4344);
not NOT1 (N6575, N6573);
nor NOR4 (N6576, N6571, N4256, N6516, N4194);
nand NAND3 (N6577, N6548, N5687, N6125);
xor XOR2 (N6578, N6564, N2414);
nor NOR4 (N6579, N6575, N260, N5429, N410);
buf BUF1 (N6580, N6557);
xor XOR2 (N6581, N6572, N4659);
or OR4 (N6582, N6574, N3712, N3519, N5619);
nand NAND2 (N6583, N6582, N5657);
nand NAND3 (N6584, N6579, N2682, N1296);
or OR4 (N6585, N6550, N1769, N2629, N3037);
xor XOR2 (N6586, N6580, N4317);
or OR4 (N6587, N6584, N3956, N6094, N196);
not NOT1 (N6588, N6565);
or OR3 (N6589, N6577, N5691, N2829);
not NOT1 (N6590, N6587);
buf BUF1 (N6591, N6569);
or OR3 (N6592, N6589, N5308, N4260);
nand NAND3 (N6593, N6576, N3146, N2878);
nand NAND2 (N6594, N6591, N1614);
xor XOR2 (N6595, N6581, N897);
nor NOR3 (N6596, N6578, N184, N1915);
and AND3 (N6597, N6585, N4556, N5423);
buf BUF1 (N6598, N6592);
or OR4 (N6599, N6593, N4327, N2893, N6470);
xor XOR2 (N6600, N6594, N6506);
nor NOR2 (N6601, N6596, N4710);
and AND4 (N6602, N6598, N4169, N1828, N533);
and AND2 (N6603, N6586, N5519);
or OR3 (N6604, N6595, N2450, N229);
buf BUF1 (N6605, N6597);
or OR2 (N6606, N6600, N4249);
buf BUF1 (N6607, N6583);
not NOT1 (N6608, N6603);
not NOT1 (N6609, N6608);
xor XOR2 (N6610, N6590, N2548);
or OR4 (N6611, N6610, N4836, N4923, N6169);
not NOT1 (N6612, N6607);
buf BUF1 (N6613, N6612);
and AND4 (N6614, N6588, N5576, N3410, N2214);
or OR3 (N6615, N6605, N770, N5645);
and AND3 (N6616, N6604, N5131, N5675);
and AND3 (N6617, N6615, N6050, N3487);
not NOT1 (N6618, N6611);
and AND4 (N6619, N6602, N4553, N4070, N1562);
buf BUF1 (N6620, N6613);
not NOT1 (N6621, N6620);
or OR2 (N6622, N6618, N3318);
or OR2 (N6623, N6616, N4606);
nand NAND3 (N6624, N6621, N1203, N1514);
or OR2 (N6625, N6617, N5345);
xor XOR2 (N6626, N6623, N5948);
buf BUF1 (N6627, N6625);
and AND3 (N6628, N6624, N6499, N3646);
or OR3 (N6629, N6628, N1666, N111);
not NOT1 (N6630, N6622);
xor XOR2 (N6631, N6619, N2949);
buf BUF1 (N6632, N6609);
xor XOR2 (N6633, N6599, N5603);
nand NAND4 (N6634, N6631, N5662, N390, N4231);
or OR4 (N6635, N6634, N3043, N5686, N1103);
not NOT1 (N6636, N6626);
buf BUF1 (N6637, N6627);
not NOT1 (N6638, N6635);
not NOT1 (N6639, N6606);
or OR2 (N6640, N6633, N2758);
nand NAND2 (N6641, N6636, N6613);
or OR2 (N6642, N6601, N6534);
nand NAND2 (N6643, N6640, N47);
nand NAND2 (N6644, N6630, N1140);
nand NAND2 (N6645, N6638, N2552);
buf BUF1 (N6646, N6643);
xor XOR2 (N6647, N6641, N902);
and AND3 (N6648, N6632, N235, N1095);
and AND4 (N6649, N6644, N5692, N2466, N3619);
xor XOR2 (N6650, N6637, N4784);
xor XOR2 (N6651, N6648, N2947);
xor XOR2 (N6652, N6645, N860);
and AND4 (N6653, N6629, N4071, N3978, N4785);
nand NAND3 (N6654, N6646, N883, N427);
not NOT1 (N6655, N6654);
or OR3 (N6656, N6649, N1123, N1557);
nand NAND4 (N6657, N6652, N6117, N4153, N105);
and AND2 (N6658, N6642, N5338);
xor XOR2 (N6659, N6651, N2908);
and AND3 (N6660, N6656, N5359, N2730);
buf BUF1 (N6661, N6660);
buf BUF1 (N6662, N6614);
or OR3 (N6663, N6639, N4654, N2373);
nor NOR2 (N6664, N6650, N337);
nor NOR4 (N6665, N6664, N4216, N3688, N3221);
xor XOR2 (N6666, N6647, N1203);
nand NAND4 (N6667, N6665, N4401, N1830, N5541);
buf BUF1 (N6668, N6666);
buf BUF1 (N6669, N6667);
buf BUF1 (N6670, N6655);
and AND4 (N6671, N6659, N2671, N6028, N5720);
nor NOR2 (N6672, N6668, N4492);
buf BUF1 (N6673, N6669);
or OR3 (N6674, N6657, N2644, N418);
xor XOR2 (N6675, N6670, N6070);
or OR4 (N6676, N6662, N31, N5089, N3736);
and AND2 (N6677, N6675, N5832);
and AND2 (N6678, N6673, N331);
and AND2 (N6679, N6676, N5397);
not NOT1 (N6680, N6663);
nor NOR3 (N6681, N6671, N805, N3551);
xor XOR2 (N6682, N6681, N2860);
and AND3 (N6683, N6653, N3716, N1558);
and AND2 (N6684, N6672, N1196);
or OR3 (N6685, N6684, N6247, N5118);
and AND4 (N6686, N6678, N6130, N5089, N6180);
xor XOR2 (N6687, N6682, N2063);
not NOT1 (N6688, N6683);
or OR3 (N6689, N6687, N1343, N1617);
buf BUF1 (N6690, N6679);
buf BUF1 (N6691, N6690);
and AND2 (N6692, N6661, N5283);
buf BUF1 (N6693, N6680);
not NOT1 (N6694, N6686);
or OR2 (N6695, N6688, N5926);
nor NOR3 (N6696, N6674, N6085, N4375);
nor NOR3 (N6697, N6677, N5310, N579);
nor NOR3 (N6698, N6689, N727, N5044);
nand NAND2 (N6699, N6697, N3411);
or OR4 (N6700, N6695, N2094, N4271, N3672);
xor XOR2 (N6701, N6693, N119);
buf BUF1 (N6702, N6696);
nor NOR2 (N6703, N6700, N4551);
buf BUF1 (N6704, N6685);
or OR2 (N6705, N6704, N1664);
buf BUF1 (N6706, N6694);
nand NAND2 (N6707, N6698, N963);
and AND2 (N6708, N6702, N3733);
and AND3 (N6709, N6706, N2357, N3298);
nand NAND2 (N6710, N6701, N6041);
or OR2 (N6711, N6703, N4672);
or OR4 (N6712, N6709, N264, N2504, N5527);
xor XOR2 (N6713, N6708, N4905);
or OR2 (N6714, N6711, N567);
buf BUF1 (N6715, N6705);
buf BUF1 (N6716, N6714);
buf BUF1 (N6717, N6692);
nand NAND2 (N6718, N6710, N1375);
buf BUF1 (N6719, N6691);
and AND2 (N6720, N6712, N3037);
not NOT1 (N6721, N6699);
not NOT1 (N6722, N6721);
buf BUF1 (N6723, N6715);
not NOT1 (N6724, N6658);
nand NAND3 (N6725, N6722, N2209, N4639);
not NOT1 (N6726, N6725);
buf BUF1 (N6727, N6716);
not NOT1 (N6728, N6717);
nor NOR4 (N6729, N6718, N1263, N4998, N1584);
not NOT1 (N6730, N6724);
not NOT1 (N6731, N6728);
nor NOR2 (N6732, N6707, N4162);
and AND4 (N6733, N6720, N4552, N3262, N2352);
nand NAND4 (N6734, N6733, N5644, N5699, N1401);
buf BUF1 (N6735, N6719);
nand NAND4 (N6736, N6734, N932, N3750, N6463);
buf BUF1 (N6737, N6726);
xor XOR2 (N6738, N6731, N5054);
nand NAND2 (N6739, N6729, N3577);
nand NAND2 (N6740, N6730, N2481);
nor NOR2 (N6741, N6736, N1754);
nor NOR4 (N6742, N6740, N2032, N4100, N2329);
nand NAND2 (N6743, N6723, N1778);
or OR2 (N6744, N6739, N3919);
nand NAND2 (N6745, N6738, N193);
buf BUF1 (N6746, N6745);
nand NAND2 (N6747, N6735, N5563);
nand NAND3 (N6748, N6732, N1129, N5655);
nor NOR4 (N6749, N6741, N2178, N829, N478);
and AND2 (N6750, N6713, N5748);
buf BUF1 (N6751, N6748);
buf BUF1 (N6752, N6737);
nor NOR2 (N6753, N6751, N4146);
xor XOR2 (N6754, N6743, N5539);
or OR2 (N6755, N6727, N1609);
xor XOR2 (N6756, N6754, N4432);
nand NAND3 (N6757, N6749, N5043, N6320);
buf BUF1 (N6758, N6755);
not NOT1 (N6759, N6744);
nand NAND3 (N6760, N6742, N2428, N3154);
xor XOR2 (N6761, N6758, N224);
nor NOR2 (N6762, N6750, N3233);
or OR4 (N6763, N6760, N6372, N485, N4223);
nor NOR3 (N6764, N6746, N5695, N1816);
or OR3 (N6765, N6756, N5727, N3527);
and AND2 (N6766, N6747, N3128);
xor XOR2 (N6767, N6759, N362);
xor XOR2 (N6768, N6766, N3311);
xor XOR2 (N6769, N6762, N131);
buf BUF1 (N6770, N6757);
or OR2 (N6771, N6768, N770);
or OR4 (N6772, N6761, N6061, N4884, N3885);
nand NAND2 (N6773, N6771, N3978);
not NOT1 (N6774, N6772);
buf BUF1 (N6775, N6752);
not NOT1 (N6776, N6775);
xor XOR2 (N6777, N6773, N5826);
nor NOR4 (N6778, N6770, N205, N538, N332);
nor NOR3 (N6779, N6777, N4566, N2198);
not NOT1 (N6780, N6753);
nand NAND4 (N6781, N6765, N3245, N5569, N5974);
nor NOR4 (N6782, N6769, N3662, N2015, N835);
not NOT1 (N6783, N6780);
nor NOR2 (N6784, N6776, N3173);
nand NAND2 (N6785, N6763, N4984);
not NOT1 (N6786, N6783);
not NOT1 (N6787, N6774);
and AND4 (N6788, N6781, N26, N1307, N2557);
nand NAND4 (N6789, N6764, N4971, N394, N3417);
or OR2 (N6790, N6788, N1592);
nand NAND3 (N6791, N6787, N1524, N5550);
nor NOR3 (N6792, N6784, N4022, N4658);
nand NAND2 (N6793, N6792, N5902);
not NOT1 (N6794, N6785);
and AND4 (N6795, N6782, N2881, N5584, N5360);
or OR2 (N6796, N6779, N5720);
xor XOR2 (N6797, N6796, N4870);
buf BUF1 (N6798, N6767);
not NOT1 (N6799, N6790);
nand NAND2 (N6800, N6799, N2092);
buf BUF1 (N6801, N6800);
and AND4 (N6802, N6797, N11, N1427, N6449);
xor XOR2 (N6803, N6786, N2222);
xor XOR2 (N6804, N6803, N6554);
xor XOR2 (N6805, N6794, N1222);
buf BUF1 (N6806, N6778);
or OR3 (N6807, N6798, N6147, N527);
and AND3 (N6808, N6801, N1174, N704);
xor XOR2 (N6809, N6795, N5897);
buf BUF1 (N6810, N6807);
nor NOR4 (N6811, N6806, N5196, N3116, N1872);
nand NAND4 (N6812, N6804, N3539, N5103, N6605);
xor XOR2 (N6813, N6791, N4988);
xor XOR2 (N6814, N6812, N2753);
or OR2 (N6815, N6811, N2409);
nand NAND2 (N6816, N6793, N4910);
nand NAND4 (N6817, N6815, N995, N6416, N5909);
and AND3 (N6818, N6809, N1171, N5896);
buf BUF1 (N6819, N6814);
xor XOR2 (N6820, N6802, N4890);
not NOT1 (N6821, N6820);
xor XOR2 (N6822, N6805, N6161);
nand NAND4 (N6823, N6810, N236, N2873, N1877);
buf BUF1 (N6824, N6816);
not NOT1 (N6825, N6822);
nor NOR2 (N6826, N6821, N5381);
xor XOR2 (N6827, N6825, N4781);
not NOT1 (N6828, N6827);
and AND3 (N6829, N6819, N2126, N1407);
nor NOR4 (N6830, N6824, N1484, N6806, N3503);
nand NAND4 (N6831, N6813, N4231, N5323, N5072);
or OR2 (N6832, N6831, N2265);
nor NOR4 (N6833, N6823, N2924, N3866, N5590);
nand NAND4 (N6834, N6829, N3709, N634, N18);
or OR2 (N6835, N6833, N3077);
buf BUF1 (N6836, N6789);
buf BUF1 (N6837, N6834);
or OR3 (N6838, N6817, N2031, N5321);
not NOT1 (N6839, N6828);
buf BUF1 (N6840, N6818);
nand NAND4 (N6841, N6830, N2542, N6388, N6600);
or OR3 (N6842, N6835, N1438, N6291);
buf BUF1 (N6843, N6840);
nand NAND4 (N6844, N6837, N2367, N1140, N2277);
nand NAND3 (N6845, N6842, N4360, N2609);
not NOT1 (N6846, N6839);
or OR3 (N6847, N6826, N1270, N3179);
xor XOR2 (N6848, N6841, N835);
nor NOR2 (N6849, N6845, N5190);
xor XOR2 (N6850, N6847, N2105);
buf BUF1 (N6851, N6846);
xor XOR2 (N6852, N6849, N6690);
or OR3 (N6853, N6836, N6562, N3348);
xor XOR2 (N6854, N6832, N1818);
not NOT1 (N6855, N6838);
nor NOR2 (N6856, N6808, N3204);
xor XOR2 (N6857, N6848, N678);
xor XOR2 (N6858, N6853, N5699);
nand NAND4 (N6859, N6857, N5237, N2962, N926);
nand NAND3 (N6860, N6844, N954, N5008);
and AND3 (N6861, N6852, N5129, N436);
buf BUF1 (N6862, N6851);
xor XOR2 (N6863, N6856, N6114);
nor NOR2 (N6864, N6858, N2452);
buf BUF1 (N6865, N6850);
and AND3 (N6866, N6865, N28, N6341);
or OR4 (N6867, N6859, N1453, N4548, N1816);
and AND4 (N6868, N6863, N5969, N687, N2286);
or OR3 (N6869, N6861, N5886, N6299);
nor NOR4 (N6870, N6864, N6308, N5977, N2937);
not NOT1 (N6871, N6854);
not NOT1 (N6872, N6855);
and AND4 (N6873, N6843, N217, N3060, N4873);
and AND3 (N6874, N6860, N3547, N5233);
xor XOR2 (N6875, N6868, N1532);
not NOT1 (N6876, N6874);
buf BUF1 (N6877, N6869);
buf BUF1 (N6878, N6876);
nor NOR2 (N6879, N6870, N2446);
not NOT1 (N6880, N6872);
and AND3 (N6881, N6878, N4448, N3009);
buf BUF1 (N6882, N6880);
and AND3 (N6883, N6877, N4144, N4579);
and AND2 (N6884, N6866, N818);
xor XOR2 (N6885, N6867, N2123);
xor XOR2 (N6886, N6881, N839);
nor NOR2 (N6887, N6886, N6707);
nand NAND3 (N6888, N6887, N1316, N1002);
nand NAND3 (N6889, N6862, N1191, N2322);
xor XOR2 (N6890, N6889, N5754);
nor NOR2 (N6891, N6871, N3364);
and AND2 (N6892, N6875, N1789);
not NOT1 (N6893, N6883);
or OR3 (N6894, N6890, N2236, N3695);
not NOT1 (N6895, N6894);
or OR4 (N6896, N6892, N2272, N4470, N3887);
and AND3 (N6897, N6888, N5756, N5562);
xor XOR2 (N6898, N6885, N2211);
or OR4 (N6899, N6895, N2415, N6767, N2200);
and AND4 (N6900, N6898, N584, N90, N1855);
not NOT1 (N6901, N6900);
or OR4 (N6902, N6891, N2675, N3919, N3032);
not NOT1 (N6903, N6882);
nor NOR4 (N6904, N6903, N2372, N1303, N5858);
xor XOR2 (N6905, N6873, N111);
and AND3 (N6906, N6901, N1316, N393);
and AND4 (N6907, N6893, N5975, N6502, N809);
or OR4 (N6908, N6896, N184, N372, N3985);
nand NAND2 (N6909, N6905, N2329);
and AND3 (N6910, N6909, N5267, N4128);
buf BUF1 (N6911, N6899);
nand NAND2 (N6912, N6907, N5906);
nor NOR3 (N6913, N6908, N560, N6360);
not NOT1 (N6914, N6879);
buf BUF1 (N6915, N6906);
buf BUF1 (N6916, N6915);
nor NOR3 (N6917, N6884, N6551, N2066);
xor XOR2 (N6918, N6914, N2534);
and AND3 (N6919, N6916, N6783, N4210);
nand NAND2 (N6920, N6912, N4377);
not NOT1 (N6921, N6918);
nand NAND4 (N6922, N6913, N6115, N6067, N329);
nor NOR4 (N6923, N6919, N3082, N1254, N4649);
nand NAND4 (N6924, N6904, N3277, N4255, N2590);
not NOT1 (N6925, N6902);
or OR4 (N6926, N6924, N6889, N5100, N6290);
nor NOR3 (N6927, N6923, N6288, N6408);
buf BUF1 (N6928, N6897);
nor NOR4 (N6929, N6922, N6125, N1888, N295);
or OR2 (N6930, N6910, N2591);
nor NOR4 (N6931, N6911, N881, N4672, N3307);
xor XOR2 (N6932, N6930, N3824);
xor XOR2 (N6933, N6920, N6588);
nand NAND4 (N6934, N6928, N4096, N6763, N418);
buf BUF1 (N6935, N6925);
and AND3 (N6936, N6934, N3661, N3621);
xor XOR2 (N6937, N6921, N498);
not NOT1 (N6938, N6917);
and AND4 (N6939, N6933, N3298, N4458, N5214);
buf BUF1 (N6940, N6939);
nor NOR4 (N6941, N6938, N5650, N4055, N6041);
nand NAND2 (N6942, N6927, N2714);
not NOT1 (N6943, N6937);
and AND3 (N6944, N6940, N6188, N3865);
xor XOR2 (N6945, N6942, N6258);
nand NAND2 (N6946, N6941, N2597);
nand NAND3 (N6947, N6944, N3413, N1956);
not NOT1 (N6948, N6932);
buf BUF1 (N6949, N6936);
nand NAND2 (N6950, N6945, N6770);
and AND2 (N6951, N6947, N2432);
nor NOR4 (N6952, N6931, N195, N384, N945);
nor NOR4 (N6953, N6948, N6738, N2321, N938);
nor NOR3 (N6954, N6943, N4567, N3135);
nor NOR4 (N6955, N6954, N3672, N4699, N1851);
nand NAND4 (N6956, N6953, N2615, N3717, N6412);
not NOT1 (N6957, N6949);
xor XOR2 (N6958, N6957, N394);
nor NOR4 (N6959, N6951, N4065, N4046, N3743);
nand NAND3 (N6960, N6946, N1924, N4916);
or OR2 (N6961, N6926, N2984);
not NOT1 (N6962, N6955);
buf BUF1 (N6963, N6962);
xor XOR2 (N6964, N6959, N685);
xor XOR2 (N6965, N6935, N5207);
xor XOR2 (N6966, N6961, N3285);
and AND2 (N6967, N6966, N6679);
nand NAND3 (N6968, N6958, N3261, N2318);
nor NOR3 (N6969, N6960, N4715, N709);
nand NAND4 (N6970, N6968, N6462, N3251, N1924);
buf BUF1 (N6971, N6965);
nor NOR3 (N6972, N6970, N4541, N1972);
or OR4 (N6973, N6952, N2478, N2643, N1709);
buf BUF1 (N6974, N6969);
nor NOR4 (N6975, N6972, N4823, N1182, N2053);
not NOT1 (N6976, N6975);
or OR2 (N6977, N6976, N1135);
not NOT1 (N6978, N6950);
nor NOR2 (N6979, N6929, N1134);
xor XOR2 (N6980, N6967, N5395);
and AND4 (N6981, N6978, N6145, N6892, N688);
buf BUF1 (N6982, N6956);
nor NOR3 (N6983, N6964, N2085, N5977);
not NOT1 (N6984, N6971);
not NOT1 (N6985, N6984);
or OR4 (N6986, N6981, N2234, N1513, N3974);
buf BUF1 (N6987, N6980);
nor NOR3 (N6988, N6983, N3177, N6500);
not NOT1 (N6989, N6977);
nor NOR2 (N6990, N6987, N323);
xor XOR2 (N6991, N6985, N2003);
nand NAND3 (N6992, N6988, N6239, N5019);
buf BUF1 (N6993, N6979);
buf BUF1 (N6994, N6990);
xor XOR2 (N6995, N6973, N4034);
not NOT1 (N6996, N6986);
not NOT1 (N6997, N6992);
and AND2 (N6998, N6989, N1334);
buf BUF1 (N6999, N6997);
buf BUF1 (N7000, N6998);
nor NOR3 (N7001, N6996, N5978, N5366);
nand NAND4 (N7002, N6999, N773, N2330, N601);
nand NAND4 (N7003, N6963, N2519, N160, N1823);
nand NAND4 (N7004, N6993, N4272, N5031, N1876);
buf BUF1 (N7005, N7004);
nor NOR3 (N7006, N6994, N6720, N1335);
and AND4 (N7007, N6974, N2995, N1405, N1305);
buf BUF1 (N7008, N7001);
xor XOR2 (N7009, N6991, N1161);
and AND2 (N7010, N7009, N6201);
nor NOR3 (N7011, N7010, N2314, N5827);
buf BUF1 (N7012, N7006);
or OR3 (N7013, N7002, N571, N2646);
nor NOR3 (N7014, N6982, N6747, N3515);
buf BUF1 (N7015, N7008);
nor NOR4 (N7016, N7012, N5088, N3873, N4880);
or OR4 (N7017, N7003, N722, N1524, N2333);
not NOT1 (N7018, N7017);
nor NOR4 (N7019, N7013, N301, N6237, N3350);
xor XOR2 (N7020, N7011, N3632);
nand NAND4 (N7021, N6995, N6954, N128, N5840);
buf BUF1 (N7022, N7005);
not NOT1 (N7023, N7020);
or OR2 (N7024, N7016, N5861);
or OR2 (N7025, N7021, N2610);
and AND2 (N7026, N7022, N4734);
and AND3 (N7027, N7014, N1340, N1946);
nor NOR3 (N7028, N7026, N1717, N6451);
or OR2 (N7029, N7019, N4203);
and AND2 (N7030, N7015, N3075);
or OR3 (N7031, N7029, N2100, N1531);
buf BUF1 (N7032, N7028);
nor NOR4 (N7033, N7018, N4173, N6686, N5008);
nor NOR4 (N7034, N7024, N497, N4075, N4989);
and AND2 (N7035, N7027, N6295);
nor NOR4 (N7036, N7033, N761, N3078, N3543);
nand NAND2 (N7037, N7007, N4234);
buf BUF1 (N7038, N7031);
and AND2 (N7039, N7000, N3684);
buf BUF1 (N7040, N7023);
not NOT1 (N7041, N7034);
nand NAND2 (N7042, N7025, N5874);
nor NOR2 (N7043, N7032, N6953);
nor NOR4 (N7044, N7043, N837, N6369, N6614);
not NOT1 (N7045, N7040);
not NOT1 (N7046, N7037);
and AND2 (N7047, N7041, N222);
nor NOR2 (N7048, N7045, N6085);
nor NOR3 (N7049, N7048, N2021, N380);
buf BUF1 (N7050, N7038);
xor XOR2 (N7051, N7046, N5823);
nand NAND2 (N7052, N7050, N1841);
xor XOR2 (N7053, N7044, N5326);
nor NOR2 (N7054, N7049, N5178);
not NOT1 (N7055, N7053);
nor NOR3 (N7056, N7047, N2107, N6899);
and AND4 (N7057, N7052, N6150, N2847, N1301);
xor XOR2 (N7058, N7039, N908);
xor XOR2 (N7059, N7057, N2444);
nor NOR2 (N7060, N7036, N312);
and AND3 (N7061, N7030, N2877, N1974);
xor XOR2 (N7062, N7054, N4119);
nand NAND4 (N7063, N7060, N2991, N2158, N4071);
nand NAND4 (N7064, N7035, N6904, N2108, N1142);
buf BUF1 (N7065, N7055);
xor XOR2 (N7066, N7061, N4830);
or OR3 (N7067, N7059, N364, N2063);
nand NAND3 (N7068, N7064, N1451, N5979);
xor XOR2 (N7069, N7062, N187);
nor NOR4 (N7070, N7051, N5069, N5811, N5287);
xor XOR2 (N7071, N7067, N2012);
buf BUF1 (N7072, N7065);
xor XOR2 (N7073, N7058, N1733);
xor XOR2 (N7074, N7073, N4861);
not NOT1 (N7075, N7074);
nor NOR4 (N7076, N7075, N2855, N3804, N5452);
nand NAND4 (N7077, N7072, N4742, N2152, N5339);
nand NAND3 (N7078, N7063, N4748, N3218);
nor NOR2 (N7079, N7077, N6817);
not NOT1 (N7080, N7076);
buf BUF1 (N7081, N7069);
or OR4 (N7082, N7081, N4703, N4698, N4975);
buf BUF1 (N7083, N7068);
nand NAND2 (N7084, N7070, N490);
and AND4 (N7085, N7082, N1726, N1658, N6804);
nand NAND2 (N7086, N7085, N3104);
or OR3 (N7087, N7066, N5675, N5780);
and AND3 (N7088, N7084, N1523, N810);
nand NAND2 (N7089, N7080, N6768);
and AND3 (N7090, N7078, N3375, N3361);
buf BUF1 (N7091, N7088);
or OR4 (N7092, N7087, N249, N2822, N5358);
not NOT1 (N7093, N7091);
or OR2 (N7094, N7090, N337);
or OR4 (N7095, N7094, N6341, N6662, N3163);
and AND4 (N7096, N7086, N1354, N5067, N2618);
nor NOR2 (N7097, N7089, N4439);
not NOT1 (N7098, N7096);
not NOT1 (N7099, N7093);
buf BUF1 (N7100, N7097);
or OR2 (N7101, N7056, N4279);
nand NAND3 (N7102, N7099, N6691, N4263);
not NOT1 (N7103, N7102);
buf BUF1 (N7104, N7101);
not NOT1 (N7105, N7071);
not NOT1 (N7106, N7103);
nor NOR2 (N7107, N7079, N562);
or OR3 (N7108, N7095, N3414, N6523);
or OR4 (N7109, N7083, N3404, N6025, N5552);
xor XOR2 (N7110, N7106, N142);
buf BUF1 (N7111, N7092);
buf BUF1 (N7112, N7111);
buf BUF1 (N7113, N7105);
not NOT1 (N7114, N7110);
or OR2 (N7115, N7109, N2438);
xor XOR2 (N7116, N7113, N2785);
nor NOR2 (N7117, N7042, N3279);
nor NOR3 (N7118, N7107, N4933, N2558);
nand NAND2 (N7119, N7104, N5480);
not NOT1 (N7120, N7114);
or OR3 (N7121, N7100, N4191, N2945);
or OR3 (N7122, N7118, N2516, N6104);
xor XOR2 (N7123, N7115, N2434);
nor NOR3 (N7124, N7119, N1612, N5404);
not NOT1 (N7125, N7121);
nand NAND3 (N7126, N7123, N1692, N3401);
and AND3 (N7127, N7125, N1112, N3984);
buf BUF1 (N7128, N7126);
nor NOR4 (N7129, N7116, N5445, N4297, N2026);
or OR2 (N7130, N7120, N4345);
nor NOR3 (N7131, N7124, N3023, N6782);
not NOT1 (N7132, N7098);
nand NAND3 (N7133, N7117, N505, N2552);
nand NAND4 (N7134, N7132, N2791, N5217, N602);
xor XOR2 (N7135, N7130, N5296);
not NOT1 (N7136, N7134);
nor NOR4 (N7137, N7131, N5809, N4631, N699);
nand NAND4 (N7138, N7129, N6614, N2340, N6359);
nor NOR3 (N7139, N7135, N6806, N2787);
and AND3 (N7140, N7127, N3645, N337);
nand NAND4 (N7141, N7108, N800, N6873, N5776);
nor NOR4 (N7142, N7138, N5841, N6053, N4725);
nor NOR2 (N7143, N7133, N649);
nand NAND3 (N7144, N7122, N1927, N8);
buf BUF1 (N7145, N7144);
nor NOR3 (N7146, N7139, N2185, N6740);
not NOT1 (N7147, N7145);
buf BUF1 (N7148, N7141);
xor XOR2 (N7149, N7136, N6722);
nor NOR3 (N7150, N7149, N403, N4443);
or OR2 (N7151, N7128, N3780);
nand NAND2 (N7152, N7137, N2113);
and AND3 (N7153, N7147, N1141, N1286);
or OR3 (N7154, N7151, N3138, N376);
and AND3 (N7155, N7150, N4131, N2347);
and AND4 (N7156, N7155, N5520, N513, N4378);
xor XOR2 (N7157, N7140, N365);
and AND2 (N7158, N7152, N4087);
nor NOR4 (N7159, N7148, N1678, N5382, N1560);
nand NAND4 (N7160, N7156, N7128, N7074, N4821);
xor XOR2 (N7161, N7112, N239);
nor NOR2 (N7162, N7142, N5508);
xor XOR2 (N7163, N7160, N1834);
nand NAND3 (N7164, N7154, N6069, N2917);
nor NOR4 (N7165, N7159, N2297, N2323, N4498);
xor XOR2 (N7166, N7165, N924);
or OR2 (N7167, N7161, N1143);
not NOT1 (N7168, N7143);
xor XOR2 (N7169, N7164, N3783);
nand NAND4 (N7170, N7146, N3876, N2578, N3338);
and AND4 (N7171, N7170, N5934, N1937, N2711);
xor XOR2 (N7172, N7168, N193);
nand NAND3 (N7173, N7171, N6538, N5915);
or OR2 (N7174, N7158, N4917);
and AND2 (N7175, N7153, N6082);
buf BUF1 (N7176, N7166);
and AND3 (N7177, N7175, N6329, N6685);
nor NOR3 (N7178, N7172, N7089, N5098);
nor NOR4 (N7179, N7178, N1397, N3037, N3227);
or OR4 (N7180, N7169, N2330, N4120, N6374);
xor XOR2 (N7181, N7167, N4510);
not NOT1 (N7182, N7176);
nand NAND2 (N7183, N7177, N3430);
or OR4 (N7184, N7173, N5437, N4446, N697);
buf BUF1 (N7185, N7183);
and AND2 (N7186, N7162, N2492);
and AND4 (N7187, N7174, N6614, N7119, N5800);
or OR4 (N7188, N7185, N1273, N3360, N6437);
and AND4 (N7189, N7163, N3939, N4691, N4268);
or OR4 (N7190, N7157, N5591, N4796, N1599);
and AND4 (N7191, N7187, N627, N6194, N5166);
nand NAND4 (N7192, N7184, N637, N3231, N1883);
nor NOR4 (N7193, N7188, N525, N5612, N3834);
nor NOR4 (N7194, N7193, N3748, N2912, N2767);
or OR4 (N7195, N7189, N2117, N6049, N6834);
xor XOR2 (N7196, N7191, N5539);
nand NAND4 (N7197, N7180, N1770, N4336, N2814);
xor XOR2 (N7198, N7186, N5611);
buf BUF1 (N7199, N7195);
nor NOR2 (N7200, N7194, N119);
buf BUF1 (N7201, N7192);
xor XOR2 (N7202, N7179, N4255);
or OR3 (N7203, N7199, N4778, N3345);
buf BUF1 (N7204, N7198);
not NOT1 (N7205, N7197);
and AND2 (N7206, N7196, N3226);
or OR4 (N7207, N7203, N2541, N5702, N5568);
not NOT1 (N7208, N7204);
xor XOR2 (N7209, N7182, N2837);
nor NOR2 (N7210, N7209, N4508);
buf BUF1 (N7211, N7190);
or OR3 (N7212, N7181, N5126, N6929);
xor XOR2 (N7213, N7202, N1237);
buf BUF1 (N7214, N7205);
nor NOR2 (N7215, N7200, N4522);
or OR2 (N7216, N7214, N1461);
nand NAND3 (N7217, N7215, N1993, N1366);
buf BUF1 (N7218, N7217);
nor NOR3 (N7219, N7207, N4500, N4798);
not NOT1 (N7220, N7211);
and AND3 (N7221, N7212, N894, N2599);
not NOT1 (N7222, N7206);
nor NOR4 (N7223, N7222, N4605, N4062, N8);
and AND3 (N7224, N7220, N3623, N7141);
buf BUF1 (N7225, N7221);
nor NOR3 (N7226, N7213, N5215, N4956);
buf BUF1 (N7227, N7225);
or OR2 (N7228, N7201, N1261);
not NOT1 (N7229, N7228);
or OR3 (N7230, N7216, N1995, N2513);
or OR3 (N7231, N7210, N4588, N3658);
or OR2 (N7232, N7224, N5100);
not NOT1 (N7233, N7230);
xor XOR2 (N7234, N7232, N3425);
xor XOR2 (N7235, N7233, N4688);
nand NAND3 (N7236, N7229, N5508, N5852);
nand NAND2 (N7237, N7226, N1590);
buf BUF1 (N7238, N7235);
nand NAND4 (N7239, N7236, N1074, N5825, N6670);
buf BUF1 (N7240, N7219);
or OR4 (N7241, N7227, N5715, N4490, N6633);
buf BUF1 (N7242, N7237);
buf BUF1 (N7243, N7208);
buf BUF1 (N7244, N7231);
nor NOR2 (N7245, N7238, N6849);
and AND4 (N7246, N7218, N75, N7209, N1590);
nor NOR4 (N7247, N7240, N3955, N2474, N6264);
nor NOR2 (N7248, N7245, N6927);
nand NAND3 (N7249, N7244, N644, N4389);
and AND2 (N7250, N7247, N4170);
nor NOR2 (N7251, N7248, N2345);
and AND2 (N7252, N7239, N1873);
not NOT1 (N7253, N7243);
and AND4 (N7254, N7252, N6553, N5448, N4336);
nor NOR4 (N7255, N7246, N3708, N4851, N4105);
buf BUF1 (N7256, N7242);
and AND4 (N7257, N7251, N5000, N6223, N5785);
or OR4 (N7258, N7254, N7183, N4487, N2153);
not NOT1 (N7259, N7253);
buf BUF1 (N7260, N7223);
and AND3 (N7261, N7257, N1749, N6367);
xor XOR2 (N7262, N7249, N6620);
buf BUF1 (N7263, N7256);
nor NOR2 (N7264, N7261, N5950);
and AND4 (N7265, N7262, N5152, N1159, N6574);
nand NAND3 (N7266, N7260, N4368, N705);
nand NAND2 (N7267, N7259, N5594);
and AND2 (N7268, N7250, N3258);
not NOT1 (N7269, N7263);
nor NOR3 (N7270, N7267, N5848, N3518);
and AND2 (N7271, N7265, N4233);
nand NAND3 (N7272, N7271, N5578, N4466);
nand NAND2 (N7273, N7270, N7188);
xor XOR2 (N7274, N7273, N1647);
and AND2 (N7275, N7272, N138);
buf BUF1 (N7276, N7264);
not NOT1 (N7277, N7258);
nor NOR4 (N7278, N7266, N852, N756, N418);
nor NOR4 (N7279, N7241, N5238, N2167, N4257);
nor NOR4 (N7280, N7276, N2196, N3224, N5305);
xor XOR2 (N7281, N7278, N114);
buf BUF1 (N7282, N7234);
xor XOR2 (N7283, N7275, N6127);
xor XOR2 (N7284, N7269, N2238);
nand NAND3 (N7285, N7281, N4309, N6613);
buf BUF1 (N7286, N7283);
and AND4 (N7287, N7280, N2086, N6605, N6110);
buf BUF1 (N7288, N7282);
not NOT1 (N7289, N7274);
buf BUF1 (N7290, N7255);
nor NOR2 (N7291, N7284, N1978);
xor XOR2 (N7292, N7290, N2797);
not NOT1 (N7293, N7289);
xor XOR2 (N7294, N7268, N2300);
xor XOR2 (N7295, N7286, N703);
and AND4 (N7296, N7295, N5923, N3174, N1639);
and AND3 (N7297, N7293, N924, N330);
buf BUF1 (N7298, N7292);
and AND2 (N7299, N7288, N2318);
buf BUF1 (N7300, N7291);
nor NOR4 (N7301, N7279, N4857, N3643, N6542);
xor XOR2 (N7302, N7300, N2553);
nand NAND4 (N7303, N7287, N6305, N4742, N3406);
buf BUF1 (N7304, N7296);
nand NAND3 (N7305, N7303, N2715, N1178);
not NOT1 (N7306, N7297);
nand NAND4 (N7307, N7277, N5699, N3070, N4259);
nand NAND2 (N7308, N7298, N103);
nor NOR4 (N7309, N7299, N3432, N4211, N7125);
buf BUF1 (N7310, N7306);
not NOT1 (N7311, N7308);
nor NOR4 (N7312, N7304, N5912, N1963, N4831);
xor XOR2 (N7313, N7301, N4554);
not NOT1 (N7314, N7311);
buf BUF1 (N7315, N7294);
or OR4 (N7316, N7309, N7118, N6138, N4671);
or OR3 (N7317, N7316, N6352, N1249);
or OR2 (N7318, N7310, N4437);
nand NAND3 (N7319, N7315, N6839, N6538);
nand NAND3 (N7320, N7317, N6798, N6508);
or OR2 (N7321, N7318, N6252);
or OR3 (N7322, N7302, N2969, N6826);
not NOT1 (N7323, N7319);
xor XOR2 (N7324, N7313, N6557);
xor XOR2 (N7325, N7323, N3283);
buf BUF1 (N7326, N7307);
xor XOR2 (N7327, N7312, N1485);
nand NAND2 (N7328, N7325, N2441);
or OR3 (N7329, N7314, N6495, N1188);
or OR2 (N7330, N7320, N935);
or OR2 (N7331, N7329, N595);
buf BUF1 (N7332, N7328);
nand NAND2 (N7333, N7321, N4854);
and AND3 (N7334, N7331, N4915, N5370);
nand NAND3 (N7335, N7322, N3875, N6195);
nand NAND2 (N7336, N7285, N7226);
nor NOR4 (N7337, N7335, N7052, N397, N5730);
nor NOR2 (N7338, N7333, N1510);
not NOT1 (N7339, N7324);
buf BUF1 (N7340, N7332);
nor NOR3 (N7341, N7337, N1012, N5846);
xor XOR2 (N7342, N7327, N4579);
not NOT1 (N7343, N7334);
buf BUF1 (N7344, N7339);
not NOT1 (N7345, N7336);
not NOT1 (N7346, N7338);
not NOT1 (N7347, N7340);
or OR2 (N7348, N7346, N4752);
not NOT1 (N7349, N7344);
xor XOR2 (N7350, N7330, N4850);
or OR3 (N7351, N7342, N6020, N944);
nor NOR2 (N7352, N7326, N6696);
xor XOR2 (N7353, N7305, N1412);
nor NOR4 (N7354, N7349, N6729, N5967, N6808);
nand NAND4 (N7355, N7348, N4878, N1157, N1132);
buf BUF1 (N7356, N7353);
nor NOR4 (N7357, N7355, N3533, N2349, N4941);
nor NOR4 (N7358, N7350, N2745, N2951, N4595);
xor XOR2 (N7359, N7354, N1823);
or OR4 (N7360, N7359, N1152, N1804, N4638);
nand NAND3 (N7361, N7358, N7075, N5130);
buf BUF1 (N7362, N7360);
nand NAND3 (N7363, N7356, N3260, N3368);
nand NAND4 (N7364, N7343, N3598, N5914, N45);
nor NOR2 (N7365, N7362, N6287);
xor XOR2 (N7366, N7364, N4403);
nor NOR4 (N7367, N7361, N1358, N602, N6545);
nand NAND2 (N7368, N7366, N653);
not NOT1 (N7369, N7363);
or OR4 (N7370, N7365, N2970, N382, N5065);
and AND3 (N7371, N7367, N7095, N2115);
or OR2 (N7372, N7368, N6895);
and AND2 (N7373, N7369, N3779);
nor NOR2 (N7374, N7352, N3139);
or OR3 (N7375, N7351, N6201, N1307);
or OR3 (N7376, N7345, N5934, N7232);
buf BUF1 (N7377, N7357);
nand NAND4 (N7378, N7377, N334, N5352, N2747);
and AND3 (N7379, N7378, N4630, N2215);
not NOT1 (N7380, N7347);
or OR2 (N7381, N7371, N6243);
buf BUF1 (N7382, N7379);
not NOT1 (N7383, N7372);
and AND3 (N7384, N7382, N2396, N5138);
nand NAND3 (N7385, N7374, N3237, N3823);
xor XOR2 (N7386, N7341, N3339);
not NOT1 (N7387, N7370);
not NOT1 (N7388, N7387);
not NOT1 (N7389, N7383);
not NOT1 (N7390, N7381);
nand NAND2 (N7391, N7384, N5699);
and AND3 (N7392, N7376, N444, N3787);
or OR2 (N7393, N7373, N105);
not NOT1 (N7394, N7385);
nand NAND2 (N7395, N7392, N4679);
nand NAND4 (N7396, N7386, N1060, N2187, N7220);
nand NAND3 (N7397, N7375, N7163, N6504);
buf BUF1 (N7398, N7390);
or OR4 (N7399, N7396, N4804, N5100, N6323);
buf BUF1 (N7400, N7394);
or OR2 (N7401, N7391, N2608);
buf BUF1 (N7402, N7401);
xor XOR2 (N7403, N7393, N3114);
not NOT1 (N7404, N7389);
or OR2 (N7405, N7399, N5744);
nand NAND2 (N7406, N7400, N4380);
xor XOR2 (N7407, N7395, N6161);
nor NOR2 (N7408, N7407, N1038);
and AND4 (N7409, N7408, N5251, N5804, N6186);
buf BUF1 (N7410, N7404);
nand NAND3 (N7411, N7388, N2562, N4183);
not NOT1 (N7412, N7398);
buf BUF1 (N7413, N7402);
xor XOR2 (N7414, N7413, N6737);
buf BUF1 (N7415, N7411);
buf BUF1 (N7416, N7405);
not NOT1 (N7417, N7403);
or OR4 (N7418, N7406, N6598, N3251, N4625);
not NOT1 (N7419, N7416);
xor XOR2 (N7420, N7410, N6980);
not NOT1 (N7421, N7414);
xor XOR2 (N7422, N7415, N57);
and AND4 (N7423, N7422, N881, N6557, N5887);
not NOT1 (N7424, N7420);
xor XOR2 (N7425, N7417, N852);
buf BUF1 (N7426, N7421);
not NOT1 (N7427, N7419);
or OR3 (N7428, N7409, N4020, N5409);
nand NAND3 (N7429, N7412, N1586, N6907);
nor NOR4 (N7430, N7423, N1389, N6677, N4208);
or OR2 (N7431, N7427, N5155);
and AND3 (N7432, N7380, N1243, N4616);
not NOT1 (N7433, N7432);
nor NOR2 (N7434, N7430, N1766);
buf BUF1 (N7435, N7397);
xor XOR2 (N7436, N7429, N4870);
xor XOR2 (N7437, N7435, N4066);
xor XOR2 (N7438, N7428, N429);
and AND4 (N7439, N7431, N3507, N7014, N6886);
nand NAND3 (N7440, N7433, N245, N3637);
buf BUF1 (N7441, N7434);
nor NOR3 (N7442, N7440, N2012, N2783);
and AND3 (N7443, N7425, N584, N2341);
and AND4 (N7444, N7441, N2691, N2531, N4456);
nand NAND4 (N7445, N7424, N2059, N7110, N3370);
and AND2 (N7446, N7426, N4536);
nor NOR4 (N7447, N7443, N753, N5962, N5254);
nor NOR2 (N7448, N7439, N2593);
nor NOR2 (N7449, N7444, N5781);
not NOT1 (N7450, N7437);
nor NOR3 (N7451, N7438, N4444, N972);
xor XOR2 (N7452, N7450, N3293);
or OR4 (N7453, N7452, N92, N2766, N2858);
or OR4 (N7454, N7418, N6655, N5444, N6957);
not NOT1 (N7455, N7445);
and AND3 (N7456, N7436, N558, N7014);
not NOT1 (N7457, N7453);
nand NAND4 (N7458, N7449, N6965, N1247, N4134);
xor XOR2 (N7459, N7446, N1705);
nor NOR3 (N7460, N7458, N565, N260);
or OR3 (N7461, N7456, N2591, N4103);
and AND3 (N7462, N7461, N7146, N6414);
buf BUF1 (N7463, N7460);
buf BUF1 (N7464, N7447);
buf BUF1 (N7465, N7462);
nand NAND4 (N7466, N7465, N5510, N3148, N6403);
xor XOR2 (N7467, N7451, N1700);
or OR2 (N7468, N7448, N6246);
nand NAND3 (N7469, N7467, N6697, N5751);
or OR2 (N7470, N7442, N3578);
nor NOR4 (N7471, N7466, N1537, N1928, N2713);
nor NOR4 (N7472, N7463, N994, N1009, N3914);
buf BUF1 (N7473, N7464);
buf BUF1 (N7474, N7457);
or OR2 (N7475, N7455, N6836);
not NOT1 (N7476, N7474);
and AND3 (N7477, N7454, N5053, N4850);
and AND4 (N7478, N7469, N6163, N1965, N2663);
xor XOR2 (N7479, N7468, N2988);
not NOT1 (N7480, N7477);
buf BUF1 (N7481, N7480);
xor XOR2 (N7482, N7470, N7344);
nand NAND4 (N7483, N7481, N804, N1236, N2713);
and AND3 (N7484, N7482, N5979, N3715);
buf BUF1 (N7485, N7459);
not NOT1 (N7486, N7473);
nor NOR3 (N7487, N7476, N5715, N4411);
nor NOR4 (N7488, N7471, N7059, N259, N280);
or OR2 (N7489, N7479, N6134);
and AND4 (N7490, N7484, N85, N5272, N357);
and AND4 (N7491, N7490, N1143, N2986, N3528);
nand NAND4 (N7492, N7475, N4427, N3730, N94);
not NOT1 (N7493, N7485);
not NOT1 (N7494, N7478);
or OR3 (N7495, N7494, N5229, N4623);
xor XOR2 (N7496, N7492, N5402);
and AND3 (N7497, N7486, N4101, N3151);
buf BUF1 (N7498, N7472);
or OR4 (N7499, N7483, N427, N4108, N2171);
and AND2 (N7500, N7487, N7201);
and AND4 (N7501, N7498, N969, N816, N1281);
nand NAND3 (N7502, N7493, N7228, N5749);
not NOT1 (N7503, N7496);
and AND4 (N7504, N7489, N6861, N438, N2340);
nor NOR3 (N7505, N7504, N3314, N7093);
nor NOR3 (N7506, N7501, N5686, N2325);
nor NOR3 (N7507, N7491, N7172, N409);
or OR2 (N7508, N7495, N5119);
and AND3 (N7509, N7497, N4625, N3407);
xor XOR2 (N7510, N7506, N5396);
not NOT1 (N7511, N7508);
not NOT1 (N7512, N7511);
nand NAND4 (N7513, N7503, N4593, N5829, N1843);
or OR4 (N7514, N7510, N1568, N1675, N6463);
buf BUF1 (N7515, N7509);
buf BUF1 (N7516, N7512);
and AND4 (N7517, N7488, N4490, N1585, N163);
nor NOR4 (N7518, N7507, N5015, N3110, N5022);
xor XOR2 (N7519, N7518, N2830);
and AND3 (N7520, N7499, N1209, N6812);
and AND4 (N7521, N7519, N2861, N3212, N3148);
xor XOR2 (N7522, N7521, N2139);
xor XOR2 (N7523, N7517, N5471);
nand NAND2 (N7524, N7515, N610);
or OR3 (N7525, N7514, N7282, N4680);
xor XOR2 (N7526, N7520, N1559);
or OR4 (N7527, N7505, N5640, N1339, N5674);
buf BUF1 (N7528, N7525);
nand NAND4 (N7529, N7528, N3122, N6080, N350);
xor XOR2 (N7530, N7523, N3079);
and AND3 (N7531, N7500, N966, N524);
and AND4 (N7532, N7531, N1958, N6152, N2219);
nor NOR4 (N7533, N7524, N818, N3098, N5315);
and AND4 (N7534, N7532, N110, N5163, N4941);
nor NOR4 (N7535, N7522, N2262, N6857, N4741);
buf BUF1 (N7536, N7513);
and AND4 (N7537, N7534, N4206, N353, N4211);
buf BUF1 (N7538, N7516);
nor NOR3 (N7539, N7526, N2107, N6419);
or OR4 (N7540, N7530, N5331, N390, N3966);
not NOT1 (N7541, N7539);
buf BUF1 (N7542, N7537);
nand NAND3 (N7543, N7529, N5031, N4277);
not NOT1 (N7544, N7540);
xor XOR2 (N7545, N7535, N671);
nand NAND3 (N7546, N7533, N5943, N4263);
buf BUF1 (N7547, N7527);
buf BUF1 (N7548, N7541);
nor NOR4 (N7549, N7547, N5546, N2030, N292);
xor XOR2 (N7550, N7543, N2281);
not NOT1 (N7551, N7550);
nor NOR4 (N7552, N7536, N6964, N4116, N4393);
nor NOR3 (N7553, N7538, N6331, N5966);
not NOT1 (N7554, N7545);
and AND2 (N7555, N7542, N1106);
nor NOR2 (N7556, N7553, N4588);
not NOT1 (N7557, N7546);
nor NOR3 (N7558, N7544, N525, N4679);
xor XOR2 (N7559, N7502, N33);
buf BUF1 (N7560, N7551);
nor NOR2 (N7561, N7556, N6348);
and AND4 (N7562, N7560, N5209, N1689, N4535);
not NOT1 (N7563, N7549);
and AND4 (N7564, N7562, N5769, N3118, N6796);
buf BUF1 (N7565, N7552);
buf BUF1 (N7566, N7558);
nor NOR2 (N7567, N7566, N3420);
xor XOR2 (N7568, N7565, N4818);
or OR4 (N7569, N7557, N5151, N579, N5985);
nor NOR2 (N7570, N7561, N902);
and AND2 (N7571, N7564, N1101);
and AND3 (N7572, N7571, N6062, N2921);
not NOT1 (N7573, N7554);
nand NAND2 (N7574, N7548, N4364);
xor XOR2 (N7575, N7563, N3661);
or OR4 (N7576, N7570, N3527, N1841, N5874);
nor NOR3 (N7577, N7573, N214, N6633);
or OR3 (N7578, N7577, N3262, N3685);
nand NAND3 (N7579, N7574, N3094, N5118);
and AND2 (N7580, N7575, N3459);
nor NOR3 (N7581, N7576, N3052, N713);
buf BUF1 (N7582, N7572);
and AND4 (N7583, N7555, N2260, N4088, N4292);
or OR4 (N7584, N7578, N845, N2399, N45);
and AND2 (N7585, N7584, N894);
not NOT1 (N7586, N7569);
nor NOR2 (N7587, N7567, N3565);
xor XOR2 (N7588, N7581, N2410);
nor NOR3 (N7589, N7579, N2534, N1373);
buf BUF1 (N7590, N7588);
nor NOR4 (N7591, N7580, N4040, N7567, N6974);
xor XOR2 (N7592, N7568, N4085);
nand NAND3 (N7593, N7587, N5631, N7197);
not NOT1 (N7594, N7592);
and AND4 (N7595, N7585, N4018, N2148, N6791);
not NOT1 (N7596, N7594);
xor XOR2 (N7597, N7589, N6991);
nand NAND3 (N7598, N7597, N6961, N5723);
buf BUF1 (N7599, N7596);
nand NAND3 (N7600, N7583, N1938, N6451);
buf BUF1 (N7601, N7591);
nor NOR3 (N7602, N7600, N100, N7409);
nand NAND2 (N7603, N7595, N854);
nand NAND2 (N7604, N7586, N76);
xor XOR2 (N7605, N7559, N3341);
xor XOR2 (N7606, N7599, N1814);
not NOT1 (N7607, N7604);
buf BUF1 (N7608, N7601);
not NOT1 (N7609, N7582);
nand NAND4 (N7610, N7607, N4310, N941, N2714);
xor XOR2 (N7611, N7609, N725);
nor NOR3 (N7612, N7608, N2115, N2975);
nand NAND2 (N7613, N7611, N3973);
nand NAND3 (N7614, N7593, N1581, N2402);
and AND3 (N7615, N7602, N3744, N4868);
not NOT1 (N7616, N7605);
buf BUF1 (N7617, N7614);
not NOT1 (N7618, N7590);
nand NAND4 (N7619, N7617, N5962, N2382, N6384);
or OR4 (N7620, N7618, N2083, N2772, N1335);
nor NOR4 (N7621, N7619, N1925, N2491, N6895);
or OR4 (N7622, N7603, N675, N7326, N6776);
buf BUF1 (N7623, N7622);
nand NAND4 (N7624, N7615, N3286, N5525, N1089);
buf BUF1 (N7625, N7623);
not NOT1 (N7626, N7625);
and AND4 (N7627, N7606, N3423, N4094, N1169);
nor NOR3 (N7628, N7624, N6038, N5620);
or OR4 (N7629, N7621, N286, N1325, N2818);
xor XOR2 (N7630, N7598, N575);
nor NOR4 (N7631, N7620, N1548, N3014, N6985);
nor NOR4 (N7632, N7631, N654, N3252, N1607);
or OR3 (N7633, N7616, N5937, N5511);
xor XOR2 (N7634, N7627, N3339);
not NOT1 (N7635, N7626);
buf BUF1 (N7636, N7610);
xor XOR2 (N7637, N7632, N4754);
nor NOR2 (N7638, N7628, N2412);
nand NAND4 (N7639, N7636, N4733, N3599, N6838);
and AND3 (N7640, N7637, N4053, N4863);
xor XOR2 (N7641, N7639, N4561);
and AND3 (N7642, N7633, N2396, N3515);
nor NOR4 (N7643, N7613, N3366, N3476, N7392);
nand NAND4 (N7644, N7643, N7017, N1335, N7567);
or OR2 (N7645, N7635, N3645);
not NOT1 (N7646, N7640);
or OR4 (N7647, N7638, N1216, N6806, N2075);
not NOT1 (N7648, N7634);
and AND3 (N7649, N7642, N3447, N4322);
and AND2 (N7650, N7612, N6517);
nand NAND2 (N7651, N7641, N1709);
or OR4 (N7652, N7646, N6345, N5849, N539);
or OR2 (N7653, N7644, N1776);
not NOT1 (N7654, N7648);
xor XOR2 (N7655, N7654, N1979);
buf BUF1 (N7656, N7629);
nand NAND3 (N7657, N7630, N6546, N6427);
and AND4 (N7658, N7649, N351, N210, N7108);
xor XOR2 (N7659, N7650, N5947);
not NOT1 (N7660, N7659);
nand NAND4 (N7661, N7657, N4664, N6423, N5085);
or OR2 (N7662, N7652, N6652);
or OR3 (N7663, N7647, N2055, N5273);
nand NAND4 (N7664, N7663, N4087, N2840, N4275);
buf BUF1 (N7665, N7655);
xor XOR2 (N7666, N7660, N1442);
xor XOR2 (N7667, N7666, N1719);
xor XOR2 (N7668, N7664, N3224);
xor XOR2 (N7669, N7662, N2908);
xor XOR2 (N7670, N7665, N2200);
nor NOR2 (N7671, N7667, N1676);
nand NAND4 (N7672, N7658, N6677, N274, N2104);
not NOT1 (N7673, N7668);
buf BUF1 (N7674, N7645);
or OR4 (N7675, N7669, N1888, N3210, N3079);
nor NOR3 (N7676, N7672, N3698, N2906);
buf BUF1 (N7677, N7675);
and AND4 (N7678, N7656, N577, N7608, N5917);
not NOT1 (N7679, N7676);
or OR3 (N7680, N7677, N6620, N2528);
buf BUF1 (N7681, N7673);
not NOT1 (N7682, N7671);
buf BUF1 (N7683, N7651);
nor NOR4 (N7684, N7679, N3194, N222, N7452);
xor XOR2 (N7685, N7683, N4367);
and AND4 (N7686, N7678, N5450, N7153, N1038);
not NOT1 (N7687, N7684);
buf BUF1 (N7688, N7686);
xor XOR2 (N7689, N7680, N2473);
not NOT1 (N7690, N7670);
nand NAND4 (N7691, N7685, N5471, N5931, N6742);
xor XOR2 (N7692, N7674, N3247);
nor NOR4 (N7693, N7653, N4895, N458, N2520);
nand NAND4 (N7694, N7692, N4196, N369, N6749);
nor NOR4 (N7695, N7691, N4186, N5656, N2138);
nand NAND4 (N7696, N7693, N5437, N6219, N5238);
nor NOR3 (N7697, N7682, N3422, N5543);
xor XOR2 (N7698, N7687, N5807);
nor NOR3 (N7699, N7694, N2808, N1239);
buf BUF1 (N7700, N7689);
nor NOR2 (N7701, N7696, N6861);
not NOT1 (N7702, N7699);
nor NOR3 (N7703, N7681, N1714, N4542);
nor NOR4 (N7704, N7701, N3467, N3925, N6642);
or OR3 (N7705, N7697, N5806, N3476);
xor XOR2 (N7706, N7700, N3646);
nor NOR2 (N7707, N7661, N7234);
nand NAND3 (N7708, N7690, N994, N3975);
not NOT1 (N7709, N7702);
or OR3 (N7710, N7705, N557, N843);
or OR3 (N7711, N7709, N3608, N218);
nor NOR3 (N7712, N7688, N1848, N1951);
xor XOR2 (N7713, N7707, N4091);
xor XOR2 (N7714, N7698, N433);
not NOT1 (N7715, N7713);
buf BUF1 (N7716, N7714);
nand NAND3 (N7717, N7716, N2440, N2803);
not NOT1 (N7718, N7704);
not NOT1 (N7719, N7711);
xor XOR2 (N7720, N7695, N2454);
nand NAND2 (N7721, N7710, N4122);
not NOT1 (N7722, N7720);
nand NAND4 (N7723, N7717, N4718, N102, N7603);
or OR2 (N7724, N7722, N6602);
nor NOR2 (N7725, N7703, N3781);
nor NOR4 (N7726, N7723, N3519, N2313, N7026);
or OR2 (N7727, N7708, N4665);
not NOT1 (N7728, N7718);
or OR4 (N7729, N7725, N1868, N3221, N6246);
nand NAND4 (N7730, N7715, N4050, N6216, N7067);
xor XOR2 (N7731, N7728, N924);
nand NAND2 (N7732, N7719, N25);
nand NAND2 (N7733, N7731, N2093);
xor XOR2 (N7734, N7712, N1719);
or OR4 (N7735, N7729, N1282, N1354, N3539);
not NOT1 (N7736, N7721);
nand NAND3 (N7737, N7724, N1156, N5269);
xor XOR2 (N7738, N7733, N6622);
not NOT1 (N7739, N7735);
or OR3 (N7740, N7739, N3815, N2851);
nand NAND2 (N7741, N7738, N6431);
nand NAND3 (N7742, N7737, N4354, N3642);
and AND3 (N7743, N7726, N248, N7692);
nor NOR2 (N7744, N7740, N14);
or OR2 (N7745, N7741, N6858);
xor XOR2 (N7746, N7744, N223);
and AND3 (N7747, N7746, N7614, N4291);
xor XOR2 (N7748, N7706, N5585);
and AND4 (N7749, N7743, N4622, N3909, N6442);
buf BUF1 (N7750, N7730);
nor NOR2 (N7751, N7745, N4778);
or OR3 (N7752, N7749, N3560, N4282);
nor NOR2 (N7753, N7742, N7662);
and AND2 (N7754, N7727, N5934);
buf BUF1 (N7755, N7750);
or OR3 (N7756, N7747, N4143, N6970);
nand NAND2 (N7757, N7734, N1068);
nor NOR2 (N7758, N7754, N6126);
not NOT1 (N7759, N7757);
or OR3 (N7760, N7755, N7141, N2478);
xor XOR2 (N7761, N7748, N7639);
not NOT1 (N7762, N7732);
nor NOR2 (N7763, N7753, N5279);
nand NAND4 (N7764, N7751, N7614, N4260, N1354);
not NOT1 (N7765, N7762);
or OR3 (N7766, N7758, N2583, N5707);
not NOT1 (N7767, N7759);
nor NOR2 (N7768, N7756, N742);
nor NOR2 (N7769, N7767, N1041);
not NOT1 (N7770, N7760);
nand NAND4 (N7771, N7766, N1509, N405, N7356);
or OR2 (N7772, N7770, N1777);
nor NOR4 (N7773, N7763, N6716, N7766, N1377);
buf BUF1 (N7774, N7771);
not NOT1 (N7775, N7772);
or OR2 (N7776, N7774, N1366);
nor NOR4 (N7777, N7769, N7400, N1869, N2505);
nand NAND4 (N7778, N7777, N4039, N4124, N3300);
not NOT1 (N7779, N7752);
or OR3 (N7780, N7773, N3173, N402);
not NOT1 (N7781, N7736);
not NOT1 (N7782, N7781);
not NOT1 (N7783, N7778);
and AND3 (N7784, N7780, N6384, N4326);
nor NOR4 (N7785, N7783, N5980, N3496, N7095);
or OR4 (N7786, N7764, N3136, N6673, N3832);
or OR3 (N7787, N7784, N4881, N7420);
buf BUF1 (N7788, N7761);
nand NAND3 (N7789, N7787, N6796, N3127);
and AND3 (N7790, N7788, N3680, N15);
nand NAND2 (N7791, N7785, N4320);
nand NAND2 (N7792, N7775, N894);
nand NAND3 (N7793, N7776, N1124, N2661);
xor XOR2 (N7794, N7779, N447);
not NOT1 (N7795, N7768);
xor XOR2 (N7796, N7765, N7668);
not NOT1 (N7797, N7789);
xor XOR2 (N7798, N7791, N6141);
nand NAND2 (N7799, N7786, N1885);
buf BUF1 (N7800, N7795);
buf BUF1 (N7801, N7793);
nand NAND3 (N7802, N7782, N6949, N2679);
nand NAND2 (N7803, N7792, N1051);
xor XOR2 (N7804, N7797, N1121);
nor NOR3 (N7805, N7790, N4904, N919);
nand NAND2 (N7806, N7794, N4934);
buf BUF1 (N7807, N7804);
and AND3 (N7808, N7806, N3515, N6279);
not NOT1 (N7809, N7805);
or OR2 (N7810, N7802, N6103);
or OR4 (N7811, N7809, N2213, N7743, N2403);
not NOT1 (N7812, N7798);
xor XOR2 (N7813, N7801, N5163);
and AND3 (N7814, N7803, N4430, N7254);
and AND2 (N7815, N7799, N1401);
or OR4 (N7816, N7807, N1911, N180, N6619);
and AND2 (N7817, N7813, N6908);
or OR2 (N7818, N7808, N7126);
nand NAND3 (N7819, N7812, N3188, N5511);
nor NOR3 (N7820, N7811, N4005, N5959);
nand NAND2 (N7821, N7796, N4228);
or OR4 (N7822, N7815, N6313, N7054, N1057);
buf BUF1 (N7823, N7814);
and AND3 (N7824, N7822, N1143, N4321);
xor XOR2 (N7825, N7823, N5826);
nor NOR4 (N7826, N7818, N3384, N4413, N1980);
nand NAND3 (N7827, N7810, N2506, N5522);
or OR2 (N7828, N7820, N7396);
nor NOR3 (N7829, N7817, N5098, N5038);
nor NOR3 (N7830, N7819, N6745, N849);
xor XOR2 (N7831, N7828, N396);
xor XOR2 (N7832, N7826, N1477);
xor XOR2 (N7833, N7827, N408);
xor XOR2 (N7834, N7832, N1368);
nor NOR2 (N7835, N7821, N4331);
and AND3 (N7836, N7835, N905, N2156);
xor XOR2 (N7837, N7824, N4353);
nand NAND4 (N7838, N7837, N3869, N6583, N4512);
nand NAND3 (N7839, N7829, N5052, N5665);
nor NOR3 (N7840, N7838, N7322, N7021);
buf BUF1 (N7841, N7836);
not NOT1 (N7842, N7800);
nand NAND4 (N7843, N7834, N7495, N1313, N1738);
nor NOR3 (N7844, N7839, N5566, N6850);
nand NAND3 (N7845, N7840, N549, N5955);
buf BUF1 (N7846, N7831);
nand NAND4 (N7847, N7833, N7725, N1759, N11);
and AND2 (N7848, N7842, N2540);
or OR3 (N7849, N7847, N710, N231);
or OR4 (N7850, N7849, N1819, N109, N7238);
and AND4 (N7851, N7846, N3664, N5808, N5421);
xor XOR2 (N7852, N7841, N411);
xor XOR2 (N7853, N7843, N3257);
and AND4 (N7854, N7851, N6925, N394, N5588);
xor XOR2 (N7855, N7825, N2358);
buf BUF1 (N7856, N7848);
buf BUF1 (N7857, N7816);
xor XOR2 (N7858, N7830, N97);
nand NAND2 (N7859, N7858, N163);
or OR3 (N7860, N7844, N2733, N7832);
buf BUF1 (N7861, N7856);
buf BUF1 (N7862, N7852);
and AND2 (N7863, N7854, N6348);
nor NOR2 (N7864, N7861, N6329);
not NOT1 (N7865, N7853);
or OR2 (N7866, N7863, N7259);
or OR3 (N7867, N7865, N2315, N273);
not NOT1 (N7868, N7867);
nor NOR3 (N7869, N7862, N3390, N7627);
xor XOR2 (N7870, N7864, N602);
xor XOR2 (N7871, N7850, N1122);
and AND2 (N7872, N7855, N1721);
not NOT1 (N7873, N7857);
not NOT1 (N7874, N7845);
nor NOR2 (N7875, N7872, N3719);
nor NOR4 (N7876, N7873, N1228, N6364, N3684);
xor XOR2 (N7877, N7871, N5445);
and AND4 (N7878, N7870, N5440, N4151, N5310);
nor NOR2 (N7879, N7860, N561);
buf BUF1 (N7880, N7866);
buf BUF1 (N7881, N7869);
xor XOR2 (N7882, N7868, N4822);
and AND2 (N7883, N7879, N1925);
xor XOR2 (N7884, N7882, N3079);
nand NAND4 (N7885, N7880, N2557, N3427, N7114);
nand NAND2 (N7886, N7885, N3704);
xor XOR2 (N7887, N7883, N3731);
and AND4 (N7888, N7875, N4232, N1741, N7040);
or OR3 (N7889, N7881, N6859, N6725);
not NOT1 (N7890, N7889);
nand NAND4 (N7891, N7888, N7596, N1576, N6484);
buf BUF1 (N7892, N7876);
not NOT1 (N7893, N7859);
buf BUF1 (N7894, N7877);
nor NOR2 (N7895, N7890, N3252);
not NOT1 (N7896, N7887);
xor XOR2 (N7897, N7895, N182);
xor XOR2 (N7898, N7892, N1009);
nand NAND4 (N7899, N7891, N4097, N2215, N4002);
nor NOR4 (N7900, N7896, N802, N3637, N3868);
not NOT1 (N7901, N7898);
and AND3 (N7902, N7894, N742, N2458);
not NOT1 (N7903, N7902);
buf BUF1 (N7904, N7900);
not NOT1 (N7905, N7893);
or OR4 (N7906, N7878, N7081, N220, N1859);
xor XOR2 (N7907, N7905, N3828);
and AND4 (N7908, N7874, N7326, N673, N1251);
nand NAND4 (N7909, N7886, N206, N4678, N6297);
xor XOR2 (N7910, N7909, N1200);
xor XOR2 (N7911, N7897, N1778);
xor XOR2 (N7912, N7907, N6624);
buf BUF1 (N7913, N7912);
buf BUF1 (N7914, N7913);
or OR4 (N7915, N7906, N1479, N2768, N6221);
buf BUF1 (N7916, N7914);
and AND4 (N7917, N7903, N973, N2967, N2720);
buf BUF1 (N7918, N7901);
or OR4 (N7919, N7916, N964, N4817, N5807);
buf BUF1 (N7920, N7910);
nand NAND4 (N7921, N7884, N7385, N5516, N3424);
or OR2 (N7922, N7917, N2017);
xor XOR2 (N7923, N7908, N1176);
buf BUF1 (N7924, N7918);
not NOT1 (N7925, N7922);
nor NOR4 (N7926, N7911, N3450, N1194, N1809);
nor NOR3 (N7927, N7924, N5416, N4663);
or OR3 (N7928, N7920, N2855, N5168);
nand NAND3 (N7929, N7923, N1308, N1881);
xor XOR2 (N7930, N7921, N7909);
and AND4 (N7931, N7928, N2283, N266, N7676);
nand NAND3 (N7932, N7931, N7332, N5509);
nand NAND2 (N7933, N7925, N7438);
not NOT1 (N7934, N7929);
buf BUF1 (N7935, N7932);
buf BUF1 (N7936, N7930);
nand NAND4 (N7937, N7899, N5356, N2458, N6330);
nor NOR4 (N7938, N7936, N2978, N3500, N5984);
and AND2 (N7939, N7926, N7290);
nand NAND2 (N7940, N7933, N1213);
or OR3 (N7941, N7904, N4833, N4153);
not NOT1 (N7942, N7941);
buf BUF1 (N7943, N7919);
nor NOR2 (N7944, N7937, N4941);
or OR2 (N7945, N7935, N7821);
and AND2 (N7946, N7940, N2639);
buf BUF1 (N7947, N7944);
and AND4 (N7948, N7915, N1988, N2516, N3966);
xor XOR2 (N7949, N7939, N2119);
not NOT1 (N7950, N7934);
nor NOR2 (N7951, N7938, N7852);
or OR4 (N7952, N7949, N2617, N5066, N2786);
buf BUF1 (N7953, N7948);
and AND2 (N7954, N7950, N7271);
and AND4 (N7955, N7946, N2705, N5271, N4031);
xor XOR2 (N7956, N7955, N3159);
or OR2 (N7957, N7942, N627);
buf BUF1 (N7958, N7945);
nand NAND4 (N7959, N7952, N4482, N848, N5521);
xor XOR2 (N7960, N7958, N1412);
nor NOR4 (N7961, N7956, N4065, N7609, N3230);
or OR2 (N7962, N7953, N4560);
nand NAND3 (N7963, N7927, N6757, N143);
buf BUF1 (N7964, N7960);
and AND2 (N7965, N7961, N63);
buf BUF1 (N7966, N7947);
buf BUF1 (N7967, N7959);
buf BUF1 (N7968, N7951);
not NOT1 (N7969, N7962);
nand NAND3 (N7970, N7963, N5946, N217);
not NOT1 (N7971, N7966);
nor NOR2 (N7972, N7969, N3926);
and AND3 (N7973, N7967, N2551, N3022);
and AND3 (N7974, N7943, N6241, N3205);
buf BUF1 (N7975, N7968);
nand NAND2 (N7976, N7973, N3126);
xor XOR2 (N7977, N7954, N4801);
nand NAND3 (N7978, N7965, N2103, N7373);
nor NOR4 (N7979, N7977, N5108, N41, N2220);
not NOT1 (N7980, N7957);
or OR3 (N7981, N7974, N4727, N4994);
nand NAND4 (N7982, N7972, N4373, N4106, N7354);
nor NOR4 (N7983, N7981, N5818, N994, N5457);
buf BUF1 (N7984, N7983);
nor NOR4 (N7985, N7980, N7610, N7789, N2929);
and AND3 (N7986, N7984, N7516, N358);
buf BUF1 (N7987, N7976);
xor XOR2 (N7988, N7986, N2960);
nand NAND3 (N7989, N7975, N2363, N4760);
not NOT1 (N7990, N7987);
nand NAND4 (N7991, N7970, N2196, N2749, N5055);
buf BUF1 (N7992, N7985);
nand NAND3 (N7993, N7979, N7922, N5415);
xor XOR2 (N7994, N7978, N4860);
and AND3 (N7995, N7982, N5384, N5041);
xor XOR2 (N7996, N7988, N1132);
and AND2 (N7997, N7989, N5453);
and AND3 (N7998, N7995, N6090, N4384);
nand NAND2 (N7999, N7964, N4329);
xor XOR2 (N8000, N7991, N984);
not NOT1 (N8001, N7992);
xor XOR2 (N8002, N8000, N7524);
nor NOR3 (N8003, N7990, N5994, N2387);
buf BUF1 (N8004, N7996);
nor NOR2 (N8005, N8001, N6885);
buf BUF1 (N8006, N8003);
xor XOR2 (N8007, N7997, N6828);
buf BUF1 (N8008, N8006);
nand NAND2 (N8009, N8008, N6774);
nand NAND4 (N8010, N7971, N5557, N761, N826);
nor NOR4 (N8011, N7998, N7417, N7569, N2852);
or OR4 (N8012, N8009, N42, N5971, N4246);
nor NOR2 (N8013, N8007, N3391);
nand NAND2 (N8014, N8012, N3683);
or OR4 (N8015, N8010, N998, N2062, N302);
endmodule