// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15;

output N2000,N1995,N2010,N2011,N2005,N1996,N2014,N2003,N2012,N2015;

or OR3 (N16, N1, N10, N6);
not NOT1 (N17, N3);
nor NOR2 (N18, N13, N8);
nor NOR2 (N19, N7, N16);
nand NAND3 (N20, N6, N14, N1);
nor NOR2 (N21, N7, N4);
and AND2 (N22, N13, N7);
buf BUF1 (N23, N16);
buf BUF1 (N24, N15);
not NOT1 (N25, N13);
not NOT1 (N26, N1);
nor NOR4 (N27, N20, N9, N14, N20);
and AND4 (N28, N17, N1, N27, N5);
nor NOR3 (N29, N18, N25, N13);
buf BUF1 (N30, N24);
buf BUF1 (N31, N23);
or OR3 (N32, N21, N28, N10);
xor XOR2 (N33, N27, N31);
or OR3 (N34, N31, N6, N4);
buf BUF1 (N35, N24);
buf BUF1 (N36, N9);
xor XOR2 (N37, N22, N14);
not NOT1 (N38, N33);
nand NAND3 (N39, N37, N27, N19);
buf BUF1 (N40, N5);
nor NOR4 (N41, N40, N13, N33, N19);
xor XOR2 (N42, N41, N5);
xor XOR2 (N43, N35, N28);
not NOT1 (N44, N43);
not NOT1 (N45, N30);
or OR3 (N46, N34, N22, N27);
and AND2 (N47, N45, N36);
nand NAND4 (N48, N8, N28, N8, N37);
not NOT1 (N49, N46);
nor NOR3 (N50, N29, N25, N10);
nand NAND3 (N51, N32, N29, N21);
and AND2 (N52, N48, N26);
nand NAND4 (N53, N28, N14, N6, N33);
nor NOR2 (N54, N39, N45);
or OR2 (N55, N44, N19);
nor NOR2 (N56, N55, N24);
and AND4 (N57, N47, N9, N24, N8);
buf BUF1 (N58, N53);
and AND3 (N59, N38, N5, N24);
xor XOR2 (N60, N42, N49);
not NOT1 (N61, N32);
nand NAND4 (N62, N52, N11, N49, N5);
not NOT1 (N63, N54);
not NOT1 (N64, N60);
or OR2 (N65, N57, N9);
or OR3 (N66, N59, N49, N54);
xor XOR2 (N67, N51, N42);
and AND3 (N68, N61, N7, N10);
nand NAND3 (N69, N64, N20, N7);
or OR3 (N70, N67, N29, N1);
or OR3 (N71, N69, N61, N9);
nand NAND2 (N72, N65, N23);
nor NOR4 (N73, N70, N57, N5, N38);
and AND2 (N74, N68, N7);
xor XOR2 (N75, N62, N47);
nor NOR3 (N76, N73, N41, N39);
or OR2 (N77, N56, N30);
buf BUF1 (N78, N75);
or OR4 (N79, N50, N6, N38, N11);
or OR4 (N80, N66, N21, N41, N6);
and AND4 (N81, N79, N46, N42, N20);
buf BUF1 (N82, N72);
xor XOR2 (N83, N81, N77);
and AND2 (N84, N12, N36);
nor NOR4 (N85, N83, N34, N24, N14);
or OR3 (N86, N82, N53, N62);
and AND4 (N87, N58, N33, N82, N55);
xor XOR2 (N88, N84, N82);
or OR3 (N89, N80, N12, N66);
or OR2 (N90, N85, N56);
xor XOR2 (N91, N90, N15);
xor XOR2 (N92, N89, N90);
not NOT1 (N93, N76);
nand NAND2 (N94, N91, N41);
nand NAND3 (N95, N63, N14, N14);
nand NAND4 (N96, N92, N17, N1, N39);
not NOT1 (N97, N78);
not NOT1 (N98, N71);
nor NOR4 (N99, N88, N6, N50, N36);
or OR2 (N100, N95, N53);
nor NOR2 (N101, N93, N92);
nor NOR2 (N102, N87, N55);
nor NOR3 (N103, N96, N91, N54);
or OR4 (N104, N74, N80, N48, N5);
buf BUF1 (N105, N86);
nand NAND3 (N106, N97, N36, N46);
nor NOR2 (N107, N106, N43);
xor XOR2 (N108, N99, N35);
nor NOR3 (N109, N107, N106, N39);
xor XOR2 (N110, N100, N44);
buf BUF1 (N111, N102);
nor NOR2 (N112, N110, N2);
and AND4 (N113, N111, N57, N18, N43);
buf BUF1 (N114, N105);
nor NOR4 (N115, N94, N34, N3, N64);
nand NAND4 (N116, N103, N22, N48, N7);
nand NAND3 (N117, N108, N104, N53);
or OR3 (N118, N39, N25, N99);
nor NOR4 (N119, N112, N87, N85, N102);
or OR3 (N120, N101, N74, N74);
nor NOR2 (N121, N119, N116);
nor NOR2 (N122, N43, N110);
buf BUF1 (N123, N114);
nor NOR3 (N124, N98, N7, N1);
nor NOR4 (N125, N109, N50, N2, N121);
and AND2 (N126, N22, N72);
nand NAND4 (N127, N113, N59, N119, N70);
or OR4 (N128, N115, N33, N40, N79);
nand NAND2 (N129, N127, N126);
not NOT1 (N130, N129);
xor XOR2 (N131, N117, N11);
buf BUF1 (N132, N47);
xor XOR2 (N133, N123, N75);
xor XOR2 (N134, N124, N94);
not NOT1 (N135, N118);
xor XOR2 (N136, N135, N70);
buf BUF1 (N137, N133);
and AND3 (N138, N122, N35, N43);
or OR2 (N139, N136, N110);
xor XOR2 (N140, N139, N17);
xor XOR2 (N141, N134, N77);
xor XOR2 (N142, N128, N22);
not NOT1 (N143, N125);
and AND4 (N144, N120, N96, N70, N111);
or OR4 (N145, N144, N93, N11, N61);
buf BUF1 (N146, N137);
not NOT1 (N147, N132);
nor NOR2 (N148, N140, N136);
and AND4 (N149, N145, N47, N93, N148);
xor XOR2 (N150, N44, N47);
nand NAND2 (N151, N131, N141);
nand NAND3 (N152, N36, N82, N103);
xor XOR2 (N153, N151, N101);
or OR3 (N154, N149, N150, N32);
not NOT1 (N155, N100);
nor NOR4 (N156, N143, N132, N51, N153);
or OR3 (N157, N45, N25, N59);
xor XOR2 (N158, N138, N72);
not NOT1 (N159, N142);
buf BUF1 (N160, N146);
or OR2 (N161, N160, N144);
xor XOR2 (N162, N147, N101);
xor XOR2 (N163, N162, N93);
or OR2 (N164, N154, N60);
nand NAND2 (N165, N161, N38);
nand NAND4 (N166, N152, N117, N154, N82);
buf BUF1 (N167, N156);
nor NOR3 (N168, N166, N51, N44);
or OR3 (N169, N167, N66, N100);
buf BUF1 (N170, N164);
buf BUF1 (N171, N155);
not NOT1 (N172, N159);
nand NAND2 (N173, N171, N137);
or OR3 (N174, N165, N82, N151);
buf BUF1 (N175, N168);
buf BUF1 (N176, N172);
or OR4 (N177, N175, N153, N120, N157);
nor NOR2 (N178, N37, N62);
nand NAND2 (N179, N177, N141);
and AND3 (N180, N176, N12, N11);
nand NAND4 (N181, N180, N177, N18, N179);
nor NOR4 (N182, N101, N160, N53, N81);
and AND2 (N183, N163, N51);
or OR4 (N184, N169, N27, N134, N6);
not NOT1 (N185, N178);
and AND4 (N186, N185, N105, N19, N166);
or OR2 (N187, N173, N130);
nand NAND2 (N188, N162, N63);
xor XOR2 (N189, N181, N57);
nand NAND3 (N190, N188, N22, N137);
nand NAND2 (N191, N183, N73);
nand NAND2 (N192, N174, N116);
xor XOR2 (N193, N189, N165);
not NOT1 (N194, N191);
nand NAND3 (N195, N194, N9, N99);
and AND4 (N196, N170, N14, N54, N111);
xor XOR2 (N197, N193, N155);
xor XOR2 (N198, N158, N16);
not NOT1 (N199, N192);
not NOT1 (N200, N182);
buf BUF1 (N201, N199);
xor XOR2 (N202, N196, N108);
and AND2 (N203, N190, N157);
and AND4 (N204, N200, N140, N34, N75);
nand NAND4 (N205, N202, N79, N149, N136);
not NOT1 (N206, N205);
nor NOR3 (N207, N201, N128, N154);
nand NAND4 (N208, N203, N114, N120, N107);
nor NOR3 (N209, N197, N71, N124);
nor NOR4 (N210, N187, N9, N199, N50);
nand NAND4 (N211, N204, N7, N160, N88);
and AND3 (N212, N211, N46, N6);
buf BUF1 (N213, N209);
or OR4 (N214, N208, N55, N29, N13);
buf BUF1 (N215, N184);
nor NOR4 (N216, N206, N107, N82, N141);
xor XOR2 (N217, N207, N204);
xor XOR2 (N218, N212, N211);
or OR3 (N219, N210, N83, N36);
nor NOR2 (N220, N198, N109);
nand NAND3 (N221, N217, N173, N54);
and AND2 (N222, N214, N29);
nand NAND3 (N223, N213, N15, N134);
and AND2 (N224, N222, N56);
not NOT1 (N225, N221);
or OR3 (N226, N186, N11, N8);
xor XOR2 (N227, N220, N166);
and AND2 (N228, N227, N28);
xor XOR2 (N229, N225, N183);
xor XOR2 (N230, N195, N183);
not NOT1 (N231, N228);
or OR2 (N232, N229, N63);
and AND3 (N233, N215, N76, N170);
or OR2 (N234, N224, N212);
xor XOR2 (N235, N218, N206);
and AND3 (N236, N216, N45, N145);
xor XOR2 (N237, N232, N164);
nand NAND2 (N238, N236, N76);
or OR2 (N239, N219, N29);
xor XOR2 (N240, N237, N167);
xor XOR2 (N241, N238, N205);
not NOT1 (N242, N226);
or OR4 (N243, N242, N46, N36, N241);
xor XOR2 (N244, N46, N158);
nor NOR2 (N245, N233, N100);
nand NAND4 (N246, N231, N143, N176, N14);
nor NOR4 (N247, N234, N212, N242, N157);
nand NAND4 (N248, N235, N69, N18, N221);
not NOT1 (N249, N239);
buf BUF1 (N250, N245);
xor XOR2 (N251, N240, N82);
and AND2 (N252, N223, N16);
nor NOR3 (N253, N250, N8, N249);
nor NOR4 (N254, N146, N113, N120, N88);
xor XOR2 (N255, N247, N56);
and AND3 (N256, N255, N36, N159);
nand NAND2 (N257, N252, N38);
buf BUF1 (N258, N253);
buf BUF1 (N259, N257);
or OR3 (N260, N254, N101, N238);
or OR4 (N261, N246, N225, N32, N9);
buf BUF1 (N262, N248);
nor NOR2 (N263, N256, N7);
buf BUF1 (N264, N230);
or OR2 (N265, N262, N48);
nor NOR2 (N266, N244, N109);
nor NOR3 (N267, N265, N9, N246);
xor XOR2 (N268, N264, N161);
and AND2 (N269, N258, N114);
nand NAND2 (N270, N259, N232);
and AND2 (N271, N268, N224);
nor NOR3 (N272, N267, N98, N4);
or OR3 (N273, N272, N121, N132);
or OR4 (N274, N270, N145, N69, N257);
or OR3 (N275, N243, N3, N181);
and AND2 (N276, N271, N107);
nand NAND4 (N277, N269, N188, N244, N74);
nor NOR4 (N278, N261, N36, N35, N248);
nand NAND4 (N279, N278, N246, N7, N20);
xor XOR2 (N280, N266, N231);
and AND2 (N281, N273, N233);
not NOT1 (N282, N263);
not NOT1 (N283, N277);
xor XOR2 (N284, N275, N230);
nor NOR4 (N285, N274, N47, N202, N223);
buf BUF1 (N286, N279);
not NOT1 (N287, N286);
and AND2 (N288, N284, N71);
buf BUF1 (N289, N285);
nor NOR4 (N290, N260, N236, N251, N285);
or OR2 (N291, N236, N117);
nor NOR3 (N292, N291, N139, N239);
xor XOR2 (N293, N288, N273);
or OR4 (N294, N282, N81, N259, N128);
and AND3 (N295, N293, N116, N38);
nor NOR2 (N296, N287, N36);
or OR3 (N297, N289, N16, N245);
nand NAND4 (N298, N281, N45, N84, N107);
nand NAND4 (N299, N290, N218, N114, N185);
and AND4 (N300, N292, N74, N60, N90);
nand NAND2 (N301, N298, N296);
buf BUF1 (N302, N40);
xor XOR2 (N303, N295, N30);
nand NAND4 (N304, N276, N253, N244, N66);
or OR2 (N305, N280, N186);
and AND3 (N306, N297, N231, N288);
and AND2 (N307, N300, N219);
buf BUF1 (N308, N306);
xor XOR2 (N309, N294, N294);
not NOT1 (N310, N309);
nand NAND2 (N311, N307, N198);
nand NAND2 (N312, N301, N145);
or OR3 (N313, N283, N240, N53);
or OR3 (N314, N303, N57, N175);
and AND3 (N315, N313, N143, N39);
buf BUF1 (N316, N311);
and AND3 (N317, N302, N87, N33);
and AND3 (N318, N314, N208, N57);
buf BUF1 (N319, N310);
nor NOR4 (N320, N316, N43, N64, N296);
nand NAND3 (N321, N305, N83, N253);
nand NAND4 (N322, N315, N10, N269, N16);
and AND2 (N323, N322, N258);
and AND3 (N324, N312, N40, N291);
nand NAND3 (N325, N318, N53, N119);
nand NAND4 (N326, N299, N208, N190, N304);
buf BUF1 (N327, N95);
nand NAND3 (N328, N308, N134, N73);
or OR4 (N329, N327, N240, N81, N296);
buf BUF1 (N330, N326);
or OR2 (N331, N329, N138);
xor XOR2 (N332, N319, N237);
nand NAND4 (N333, N320, N308, N28, N18);
nor NOR2 (N334, N330, N158);
xor XOR2 (N335, N331, N190);
buf BUF1 (N336, N323);
and AND2 (N337, N336, N90);
nand NAND3 (N338, N334, N170, N183);
nand NAND4 (N339, N338, N186, N303, N3);
nor NOR3 (N340, N333, N170, N114);
xor XOR2 (N341, N332, N145);
xor XOR2 (N342, N341, N200);
buf BUF1 (N343, N337);
not NOT1 (N344, N339);
and AND2 (N345, N328, N111);
nand NAND2 (N346, N345, N241);
xor XOR2 (N347, N317, N17);
not NOT1 (N348, N342);
nand NAND4 (N349, N325, N172, N105, N218);
or OR4 (N350, N335, N64, N180, N336);
and AND4 (N351, N347, N178, N135, N284);
or OR4 (N352, N344, N3, N276, N260);
nand NAND4 (N353, N324, N16, N207, N217);
nand NAND2 (N354, N353, N310);
not NOT1 (N355, N351);
nor NOR4 (N356, N346, N289, N13, N11);
not NOT1 (N357, N354);
nand NAND4 (N358, N343, N102, N207, N35);
nand NAND3 (N359, N340, N204, N121);
not NOT1 (N360, N356);
xor XOR2 (N361, N352, N94);
nor NOR2 (N362, N359, N205);
buf BUF1 (N363, N361);
or OR3 (N364, N355, N269, N157);
xor XOR2 (N365, N364, N266);
buf BUF1 (N366, N363);
nand NAND2 (N367, N348, N132);
xor XOR2 (N368, N365, N45);
xor XOR2 (N369, N350, N211);
and AND3 (N370, N358, N325, N182);
nand NAND4 (N371, N360, N191, N25, N113);
nor NOR3 (N372, N370, N203, N94);
nand NAND4 (N373, N362, N167, N352, N6);
and AND2 (N374, N372, N353);
xor XOR2 (N375, N321, N67);
nor NOR3 (N376, N375, N22, N18);
nand NAND2 (N377, N376, N49);
not NOT1 (N378, N368);
xor XOR2 (N379, N349, N99);
not NOT1 (N380, N369);
nor NOR4 (N381, N367, N146, N169, N247);
xor XOR2 (N382, N357, N171);
and AND2 (N383, N371, N270);
and AND2 (N384, N374, N24);
or OR3 (N385, N377, N192, N149);
buf BUF1 (N386, N385);
nand NAND3 (N387, N380, N203, N258);
nand NAND3 (N388, N378, N262, N260);
not NOT1 (N389, N388);
nand NAND2 (N390, N373, N300);
or OR3 (N391, N381, N301, N3);
nand NAND4 (N392, N390, N160, N147, N363);
nand NAND4 (N393, N386, N290, N311, N342);
not NOT1 (N394, N392);
xor XOR2 (N395, N379, N223);
not NOT1 (N396, N395);
nand NAND2 (N397, N382, N58);
nand NAND3 (N398, N384, N112, N171);
not NOT1 (N399, N398);
buf BUF1 (N400, N397);
buf BUF1 (N401, N366);
and AND4 (N402, N396, N393, N8, N338);
not NOT1 (N403, N120);
and AND3 (N404, N401, N18, N27);
or OR3 (N405, N383, N145, N327);
nand NAND4 (N406, N405, N396, N263, N286);
or OR4 (N407, N394, N229, N16, N349);
nand NAND2 (N408, N391, N365);
nor NOR4 (N409, N404, N402, N330, N165);
and AND2 (N410, N18, N342);
not NOT1 (N411, N403);
buf BUF1 (N412, N389);
and AND4 (N413, N400, N112, N63, N149);
not NOT1 (N414, N413);
not NOT1 (N415, N409);
not NOT1 (N416, N387);
and AND2 (N417, N411, N138);
or OR3 (N418, N415, N188, N72);
nor NOR2 (N419, N410, N73);
xor XOR2 (N420, N417, N158);
nand NAND4 (N421, N419, N210, N359, N67);
buf BUF1 (N422, N407);
xor XOR2 (N423, N406, N36);
nand NAND3 (N424, N399, N122, N37);
buf BUF1 (N425, N424);
and AND2 (N426, N425, N196);
not NOT1 (N427, N414);
and AND2 (N428, N420, N259);
nand NAND2 (N429, N426, N242);
and AND3 (N430, N416, N417, N98);
and AND3 (N431, N418, N185, N261);
or OR2 (N432, N430, N290);
and AND4 (N433, N431, N274, N356, N360);
xor XOR2 (N434, N422, N106);
or OR4 (N435, N434, N103, N217, N145);
not NOT1 (N436, N429);
xor XOR2 (N437, N435, N388);
xor XOR2 (N438, N433, N311);
nor NOR3 (N439, N421, N73, N35);
xor XOR2 (N440, N432, N386);
xor XOR2 (N441, N412, N3);
and AND4 (N442, N437, N103, N319, N86);
and AND3 (N443, N438, N190, N238);
buf BUF1 (N444, N440);
nand NAND2 (N445, N444, N322);
not NOT1 (N446, N423);
and AND2 (N447, N442, N204);
or OR3 (N448, N428, N430, N343);
nor NOR2 (N449, N447, N313);
nand NAND2 (N450, N427, N6);
xor XOR2 (N451, N441, N368);
xor XOR2 (N452, N450, N52);
nand NAND3 (N453, N452, N115, N141);
buf BUF1 (N454, N443);
not NOT1 (N455, N449);
and AND2 (N456, N453, N210);
nand NAND4 (N457, N454, N332, N99, N378);
nor NOR2 (N458, N436, N195);
buf BUF1 (N459, N439);
buf BUF1 (N460, N448);
xor XOR2 (N461, N451, N437);
and AND2 (N462, N446, N250);
nor NOR4 (N463, N456, N79, N18, N289);
not NOT1 (N464, N461);
nand NAND4 (N465, N445, N317, N77, N39);
nand NAND3 (N466, N408, N30, N43);
and AND3 (N467, N466, N47, N98);
buf BUF1 (N468, N455);
buf BUF1 (N469, N457);
and AND2 (N470, N469, N320);
and AND2 (N471, N462, N447);
buf BUF1 (N472, N458);
and AND2 (N473, N472, N266);
and AND3 (N474, N465, N241, N92);
nor NOR4 (N475, N468, N473, N150, N452);
nand NAND2 (N476, N447, N357);
nand NAND2 (N477, N474, N451);
not NOT1 (N478, N471);
not NOT1 (N479, N464);
not NOT1 (N480, N463);
and AND3 (N481, N470, N283, N299);
buf BUF1 (N482, N481);
xor XOR2 (N483, N459, N284);
nor NOR4 (N484, N479, N107, N207, N15);
nand NAND3 (N485, N484, N324, N418);
nor NOR2 (N486, N476, N8);
nor NOR2 (N487, N475, N175);
and AND4 (N488, N485, N384, N185, N397);
xor XOR2 (N489, N488, N85);
nor NOR2 (N490, N482, N87);
buf BUF1 (N491, N489);
or OR4 (N492, N477, N115, N399, N33);
or OR3 (N493, N460, N361, N314);
nand NAND2 (N494, N486, N180);
nand NAND4 (N495, N487, N42, N138, N3);
and AND3 (N496, N480, N399, N147);
nand NAND3 (N497, N478, N199, N241);
nor NOR3 (N498, N497, N235, N234);
not NOT1 (N499, N490);
buf BUF1 (N500, N496);
buf BUF1 (N501, N495);
xor XOR2 (N502, N491, N429);
or OR2 (N503, N467, N488);
xor XOR2 (N504, N503, N203);
or OR4 (N505, N502, N9, N92, N269);
and AND4 (N506, N493, N234, N278, N127);
xor XOR2 (N507, N501, N70);
or OR3 (N508, N505, N400, N369);
nand NAND2 (N509, N492, N319);
nor NOR4 (N510, N494, N378, N32, N287);
nor NOR2 (N511, N508, N266);
and AND2 (N512, N510, N152);
buf BUF1 (N513, N506);
or OR2 (N514, N509, N179);
nand NAND2 (N515, N499, N18);
nor NOR3 (N516, N500, N64, N301);
not NOT1 (N517, N516);
or OR3 (N518, N498, N317, N473);
nor NOR3 (N519, N507, N404, N270);
xor XOR2 (N520, N512, N230);
nand NAND4 (N521, N513, N81, N104, N396);
xor XOR2 (N522, N483, N14);
xor XOR2 (N523, N521, N349);
nor NOR4 (N524, N517, N28, N58, N456);
buf BUF1 (N525, N522);
nand NAND2 (N526, N523, N517);
nand NAND4 (N527, N511, N32, N20, N162);
not NOT1 (N528, N515);
buf BUF1 (N529, N519);
nand NAND2 (N530, N520, N342);
not NOT1 (N531, N529);
not NOT1 (N532, N514);
xor XOR2 (N533, N504, N363);
and AND4 (N534, N528, N523, N238, N103);
xor XOR2 (N535, N525, N202);
nand NAND4 (N536, N527, N443, N385, N44);
nand NAND2 (N537, N518, N163);
or OR4 (N538, N537, N358, N203, N109);
xor XOR2 (N539, N524, N317);
not NOT1 (N540, N539);
and AND3 (N541, N530, N204, N428);
or OR3 (N542, N533, N168, N9);
and AND2 (N543, N536, N399);
nand NAND2 (N544, N531, N243);
nor NOR4 (N545, N541, N307, N201, N47);
nand NAND4 (N546, N540, N166, N386, N15);
nand NAND4 (N547, N543, N312, N319, N229);
and AND2 (N548, N545, N41);
buf BUF1 (N549, N542);
xor XOR2 (N550, N546, N1);
and AND2 (N551, N547, N57);
buf BUF1 (N552, N535);
nand NAND4 (N553, N552, N542, N182, N314);
and AND2 (N554, N526, N46);
nor NOR4 (N555, N551, N518, N413, N459);
nand NAND4 (N556, N544, N60, N260, N423);
not NOT1 (N557, N534);
buf BUF1 (N558, N553);
xor XOR2 (N559, N550, N146);
xor XOR2 (N560, N532, N110);
nand NAND3 (N561, N558, N274, N190);
buf BUF1 (N562, N556);
buf BUF1 (N563, N559);
or OR3 (N564, N562, N179, N287);
and AND4 (N565, N555, N15, N470, N468);
or OR3 (N566, N549, N316, N49);
nand NAND3 (N567, N561, N258, N198);
or OR4 (N568, N565, N30, N30, N488);
and AND2 (N569, N560, N95);
or OR4 (N570, N564, N61, N369, N68);
or OR3 (N571, N566, N150, N327);
not NOT1 (N572, N569);
or OR3 (N573, N572, N50, N465);
buf BUF1 (N574, N570);
nand NAND2 (N575, N574, N339);
not NOT1 (N576, N548);
buf BUF1 (N577, N568);
xor XOR2 (N578, N563, N87);
nor NOR3 (N579, N557, N382, N396);
or OR2 (N580, N575, N391);
buf BUF1 (N581, N554);
xor XOR2 (N582, N577, N163);
nor NOR2 (N583, N538, N506);
xor XOR2 (N584, N571, N275);
nand NAND4 (N585, N582, N191, N543, N402);
xor XOR2 (N586, N578, N440);
xor XOR2 (N587, N573, N162);
or OR4 (N588, N576, N404, N581, N152);
nor NOR3 (N589, N1, N554, N162);
nor NOR4 (N590, N586, N458, N97, N435);
xor XOR2 (N591, N585, N462);
xor XOR2 (N592, N589, N447);
and AND4 (N593, N579, N395, N129, N379);
nand NAND4 (N594, N584, N53, N514, N280);
not NOT1 (N595, N567);
or OR4 (N596, N583, N75, N393, N318);
not NOT1 (N597, N594);
or OR3 (N598, N590, N208, N414);
or OR3 (N599, N592, N573, N415);
or OR4 (N600, N588, N212, N254, N542);
not NOT1 (N601, N599);
nor NOR4 (N602, N593, N177, N128, N109);
not NOT1 (N603, N601);
xor XOR2 (N604, N580, N394);
nand NAND3 (N605, N603, N157, N304);
buf BUF1 (N606, N604);
nand NAND2 (N607, N600, N22);
xor XOR2 (N608, N607, N298);
nand NAND4 (N609, N587, N2, N418, N331);
xor XOR2 (N610, N608, N537);
and AND4 (N611, N598, N548, N82, N145);
and AND2 (N612, N606, N440);
or OR4 (N613, N597, N508, N521, N136);
nand NAND3 (N614, N602, N222, N154);
nor NOR2 (N615, N605, N326);
and AND4 (N616, N595, N220, N328, N536);
or OR3 (N617, N613, N421, N451);
not NOT1 (N618, N616);
nor NOR3 (N619, N610, N516, N119);
xor XOR2 (N620, N609, N434);
not NOT1 (N621, N619);
nand NAND2 (N622, N596, N220);
buf BUF1 (N623, N620);
xor XOR2 (N624, N618, N1);
xor XOR2 (N625, N591, N176);
or OR2 (N626, N621, N174);
nor NOR3 (N627, N611, N248, N487);
buf BUF1 (N628, N626);
not NOT1 (N629, N612);
nor NOR3 (N630, N627, N394, N339);
buf BUF1 (N631, N614);
nand NAND2 (N632, N625, N258);
not NOT1 (N633, N630);
not NOT1 (N634, N624);
xor XOR2 (N635, N633, N448);
nand NAND3 (N636, N632, N230, N297);
or OR4 (N637, N635, N175, N193, N355);
xor XOR2 (N638, N631, N625);
buf BUF1 (N639, N628);
buf BUF1 (N640, N637);
xor XOR2 (N641, N622, N152);
nor NOR3 (N642, N634, N277, N359);
nand NAND3 (N643, N623, N160, N39);
nand NAND3 (N644, N617, N236, N24);
nor NOR3 (N645, N639, N33, N161);
or OR2 (N646, N642, N199);
nor NOR4 (N647, N638, N552, N176, N333);
or OR3 (N648, N646, N601, N336);
and AND3 (N649, N629, N384, N106);
nor NOR2 (N650, N643, N145);
xor XOR2 (N651, N650, N266);
buf BUF1 (N652, N649);
buf BUF1 (N653, N640);
buf BUF1 (N654, N644);
buf BUF1 (N655, N651);
and AND4 (N656, N645, N521, N571, N547);
xor XOR2 (N657, N656, N441);
not NOT1 (N658, N636);
nand NAND4 (N659, N657, N77, N403, N531);
or OR4 (N660, N648, N408, N373, N573);
nand NAND3 (N661, N659, N421, N471);
buf BUF1 (N662, N655);
xor XOR2 (N663, N654, N375);
not NOT1 (N664, N662);
and AND4 (N665, N664, N302, N400, N514);
not NOT1 (N666, N647);
xor XOR2 (N667, N658, N305);
or OR3 (N668, N666, N147, N309);
nand NAND2 (N669, N663, N259);
not NOT1 (N670, N667);
and AND2 (N671, N653, N231);
and AND4 (N672, N670, N365, N554, N246);
nor NOR3 (N673, N641, N448, N236);
not NOT1 (N674, N673);
not NOT1 (N675, N661);
nor NOR4 (N676, N675, N153, N411, N57);
or OR3 (N677, N669, N184, N549);
xor XOR2 (N678, N668, N547);
and AND3 (N679, N676, N342, N66);
and AND4 (N680, N672, N656, N77, N489);
and AND4 (N681, N615, N658, N654, N171);
xor XOR2 (N682, N671, N383);
nand NAND2 (N683, N678, N356);
not NOT1 (N684, N674);
xor XOR2 (N685, N683, N412);
nand NAND4 (N686, N682, N479, N671, N409);
or OR2 (N687, N677, N399);
not NOT1 (N688, N680);
buf BUF1 (N689, N679);
nor NOR4 (N690, N660, N401, N650, N242);
and AND4 (N691, N688, N188, N359, N158);
xor XOR2 (N692, N690, N546);
nor NOR3 (N693, N691, N637, N665);
nand NAND4 (N694, N488, N509, N185, N499);
or OR4 (N695, N692, N270, N82, N496);
and AND4 (N696, N687, N101, N624, N337);
xor XOR2 (N697, N685, N555);
and AND4 (N698, N681, N90, N167, N638);
buf BUF1 (N699, N652);
not NOT1 (N700, N698);
xor XOR2 (N701, N689, N578);
xor XOR2 (N702, N693, N686);
or OR3 (N703, N48, N109, N166);
nor NOR4 (N704, N699, N267, N386, N148);
buf BUF1 (N705, N697);
xor XOR2 (N706, N696, N399);
nor NOR2 (N707, N700, N592);
not NOT1 (N708, N701);
nand NAND2 (N709, N702, N75);
nor NOR2 (N710, N708, N501);
and AND3 (N711, N695, N323, N655);
nand NAND3 (N712, N710, N316, N111);
nor NOR2 (N713, N684, N96);
or OR2 (N714, N704, N307);
nor NOR4 (N715, N709, N676, N220, N602);
not NOT1 (N716, N714);
nor NOR2 (N717, N712, N418);
nand NAND4 (N718, N715, N366, N423, N571);
not NOT1 (N719, N707);
not NOT1 (N720, N706);
nand NAND4 (N721, N717, N495, N375, N573);
not NOT1 (N722, N713);
and AND3 (N723, N703, N469, N408);
xor XOR2 (N724, N720, N628);
nor NOR3 (N725, N721, N490, N354);
nand NAND4 (N726, N723, N452, N260, N18);
not NOT1 (N727, N724);
nand NAND3 (N728, N711, N310, N506);
xor XOR2 (N729, N727, N567);
and AND3 (N730, N694, N27, N672);
not NOT1 (N731, N722);
and AND4 (N732, N731, N401, N152, N578);
and AND2 (N733, N726, N586);
and AND4 (N734, N718, N387, N340, N164);
or OR3 (N735, N734, N338, N90);
buf BUF1 (N736, N719);
xor XOR2 (N737, N736, N682);
nor NOR4 (N738, N732, N595, N461, N181);
nand NAND4 (N739, N737, N410, N305, N32);
buf BUF1 (N740, N705);
and AND4 (N741, N730, N515, N396, N245);
not NOT1 (N742, N733);
and AND3 (N743, N735, N285, N521);
buf BUF1 (N744, N741);
xor XOR2 (N745, N742, N740);
nand NAND2 (N746, N350, N667);
nand NAND3 (N747, N746, N381, N297);
nor NOR4 (N748, N738, N471, N39, N292);
nor NOR2 (N749, N744, N100);
and AND4 (N750, N739, N406, N659, N173);
and AND4 (N751, N728, N126, N40, N23);
or OR3 (N752, N725, N224, N230);
xor XOR2 (N753, N743, N385);
and AND2 (N754, N716, N44);
and AND2 (N755, N747, N449);
nor NOR3 (N756, N749, N503, N562);
buf BUF1 (N757, N750);
nand NAND2 (N758, N729, N742);
xor XOR2 (N759, N751, N73);
or OR4 (N760, N754, N530, N568, N463);
not NOT1 (N761, N755);
buf BUF1 (N762, N752);
not NOT1 (N763, N745);
and AND2 (N764, N757, N443);
xor XOR2 (N765, N753, N598);
buf BUF1 (N766, N759);
buf BUF1 (N767, N758);
nand NAND4 (N768, N767, N264, N471, N82);
xor XOR2 (N769, N762, N272);
not NOT1 (N770, N763);
nor NOR3 (N771, N769, N58, N88);
and AND4 (N772, N765, N674, N272, N610);
xor XOR2 (N773, N770, N77);
nand NAND3 (N774, N748, N509, N12);
xor XOR2 (N775, N766, N364);
xor XOR2 (N776, N756, N451);
nand NAND3 (N777, N774, N292, N469);
not NOT1 (N778, N768);
and AND4 (N779, N772, N403, N361, N367);
or OR4 (N780, N760, N245, N588, N673);
xor XOR2 (N781, N771, N220);
xor XOR2 (N782, N773, N67);
xor XOR2 (N783, N777, N73);
and AND2 (N784, N776, N242);
and AND2 (N785, N775, N628);
not NOT1 (N786, N778);
not NOT1 (N787, N785);
or OR4 (N788, N761, N172, N365, N771);
nand NAND4 (N789, N781, N122, N336, N361);
nand NAND4 (N790, N764, N260, N765, N499);
buf BUF1 (N791, N789);
or OR3 (N792, N790, N485, N469);
not NOT1 (N793, N784);
not NOT1 (N794, N782);
and AND2 (N795, N791, N424);
not NOT1 (N796, N787);
nand NAND2 (N797, N786, N363);
xor XOR2 (N798, N793, N361);
nand NAND4 (N799, N780, N544, N765, N117);
nor NOR2 (N800, N796, N463);
not NOT1 (N801, N792);
xor XOR2 (N802, N798, N582);
xor XOR2 (N803, N783, N784);
or OR3 (N804, N799, N146, N699);
nand NAND3 (N805, N803, N168, N164);
nand NAND3 (N806, N794, N49, N250);
nand NAND4 (N807, N804, N388, N51, N753);
buf BUF1 (N808, N800);
xor XOR2 (N809, N801, N274);
xor XOR2 (N810, N795, N10);
or OR3 (N811, N808, N179, N549);
or OR4 (N812, N788, N773, N683, N90);
not NOT1 (N813, N797);
and AND2 (N814, N802, N82);
not NOT1 (N815, N805);
or OR4 (N816, N814, N25, N288, N434);
not NOT1 (N817, N816);
nand NAND3 (N818, N806, N527, N300);
or OR2 (N819, N779, N40);
not NOT1 (N820, N815);
and AND3 (N821, N807, N309, N816);
xor XOR2 (N822, N821, N537);
buf BUF1 (N823, N810);
buf BUF1 (N824, N809);
nand NAND2 (N825, N818, N178);
nor NOR3 (N826, N820, N491, N669);
or OR4 (N827, N823, N808, N709, N143);
or OR4 (N828, N813, N88, N186, N22);
not NOT1 (N829, N827);
and AND3 (N830, N811, N95, N765);
and AND3 (N831, N819, N136, N628);
nor NOR3 (N832, N829, N237, N11);
xor XOR2 (N833, N828, N620);
nor NOR4 (N834, N831, N407, N263, N527);
and AND3 (N835, N822, N124, N702);
or OR4 (N836, N833, N162, N592, N710);
or OR3 (N837, N830, N577, N357);
and AND2 (N838, N836, N45);
and AND4 (N839, N838, N347, N136, N259);
and AND3 (N840, N825, N156, N624);
nor NOR2 (N841, N824, N618);
and AND3 (N842, N839, N794, N686);
buf BUF1 (N843, N812);
buf BUF1 (N844, N842);
xor XOR2 (N845, N832, N137);
and AND3 (N846, N826, N616, N724);
xor XOR2 (N847, N841, N252);
or OR3 (N848, N846, N602, N501);
xor XOR2 (N849, N847, N215);
and AND4 (N850, N835, N387, N431, N94);
nor NOR3 (N851, N843, N683, N151);
not NOT1 (N852, N834);
xor XOR2 (N853, N844, N378);
not NOT1 (N854, N851);
buf BUF1 (N855, N850);
nand NAND2 (N856, N840, N43);
not NOT1 (N857, N854);
and AND4 (N858, N857, N56, N433, N485);
or OR3 (N859, N845, N291, N816);
and AND2 (N860, N858, N655);
xor XOR2 (N861, N852, N315);
not NOT1 (N862, N859);
or OR3 (N863, N855, N799, N583);
not NOT1 (N864, N863);
xor XOR2 (N865, N861, N728);
or OR2 (N866, N853, N279);
not NOT1 (N867, N860);
and AND4 (N868, N817, N10, N341, N545);
buf BUF1 (N869, N856);
not NOT1 (N870, N867);
nand NAND3 (N871, N868, N219, N158);
and AND2 (N872, N865, N741);
buf BUF1 (N873, N872);
nor NOR3 (N874, N849, N655, N130);
not NOT1 (N875, N862);
and AND3 (N876, N870, N473, N217);
and AND2 (N877, N876, N847);
xor XOR2 (N878, N874, N173);
and AND3 (N879, N878, N655, N39);
nand NAND4 (N880, N864, N795, N795, N66);
and AND3 (N881, N873, N47, N513);
buf BUF1 (N882, N837);
and AND4 (N883, N882, N556, N723, N335);
not NOT1 (N884, N877);
and AND3 (N885, N879, N84, N866);
buf BUF1 (N886, N324);
nand NAND2 (N887, N871, N680);
buf BUF1 (N888, N887);
buf BUF1 (N889, N888);
nor NOR3 (N890, N869, N123, N275);
buf BUF1 (N891, N885);
nand NAND2 (N892, N883, N529);
nor NOR2 (N893, N890, N804);
buf BUF1 (N894, N884);
buf BUF1 (N895, N891);
and AND3 (N896, N848, N211, N139);
or OR2 (N897, N875, N890);
buf BUF1 (N898, N880);
nor NOR4 (N899, N897, N409, N40, N800);
nand NAND2 (N900, N889, N757);
not NOT1 (N901, N900);
or OR2 (N902, N881, N48);
xor XOR2 (N903, N886, N858);
xor XOR2 (N904, N894, N496);
buf BUF1 (N905, N896);
nand NAND2 (N906, N905, N548);
or OR3 (N907, N899, N380, N173);
not NOT1 (N908, N902);
and AND2 (N909, N901, N581);
and AND4 (N910, N895, N631, N820, N19);
not NOT1 (N911, N906);
or OR3 (N912, N903, N56, N776);
nor NOR4 (N913, N907, N901, N415, N563);
buf BUF1 (N914, N898);
xor XOR2 (N915, N909, N57);
nor NOR3 (N916, N911, N646, N772);
nand NAND4 (N917, N892, N566, N53, N882);
nor NOR3 (N918, N893, N323, N460);
nand NAND2 (N919, N904, N141);
or OR3 (N920, N915, N534, N130);
nand NAND4 (N921, N908, N764, N784, N136);
or OR2 (N922, N910, N122);
nand NAND3 (N923, N922, N522, N823);
or OR2 (N924, N918, N893);
not NOT1 (N925, N921);
xor XOR2 (N926, N924, N734);
xor XOR2 (N927, N919, N104);
not NOT1 (N928, N913);
and AND2 (N929, N912, N279);
nor NOR3 (N930, N914, N885, N837);
nand NAND3 (N931, N916, N682, N823);
or OR4 (N932, N930, N202, N313, N114);
nor NOR3 (N933, N931, N753, N515);
buf BUF1 (N934, N929);
nor NOR2 (N935, N923, N300);
nand NAND4 (N936, N920, N744, N144, N244);
not NOT1 (N937, N933);
nor NOR2 (N938, N934, N69);
and AND4 (N939, N927, N192, N266, N794);
and AND4 (N940, N917, N322, N410, N403);
xor XOR2 (N941, N937, N285);
buf BUF1 (N942, N938);
and AND4 (N943, N940, N12, N671, N113);
nor NOR4 (N944, N925, N474, N204, N17);
buf BUF1 (N945, N941);
xor XOR2 (N946, N935, N160);
nand NAND2 (N947, N932, N859);
not NOT1 (N948, N943);
or OR4 (N949, N947, N789, N220, N492);
not NOT1 (N950, N936);
xor XOR2 (N951, N942, N58);
nor NOR3 (N952, N951, N731, N150);
nor NOR4 (N953, N939, N157, N854, N859);
nor NOR4 (N954, N945, N370, N588, N928);
nor NOR2 (N955, N456, N239);
nor NOR2 (N956, N944, N929);
xor XOR2 (N957, N926, N950);
nand NAND3 (N958, N413, N207, N328);
not NOT1 (N959, N946);
nand NAND4 (N960, N954, N264, N419, N443);
nor NOR2 (N961, N948, N498);
buf BUF1 (N962, N952);
or OR4 (N963, N953, N655, N722, N866);
nor NOR2 (N964, N958, N431);
nor NOR4 (N965, N962, N328, N328, N850);
or OR4 (N966, N959, N48, N77, N812);
or OR2 (N967, N949, N1);
and AND2 (N968, N956, N366);
not NOT1 (N969, N968);
nand NAND4 (N970, N966, N370, N369, N761);
xor XOR2 (N971, N955, N863);
xor XOR2 (N972, N960, N323);
nor NOR3 (N973, N969, N720, N799);
buf BUF1 (N974, N961);
nor NOR4 (N975, N970, N851, N588, N800);
nand NAND3 (N976, N972, N146, N747);
xor XOR2 (N977, N976, N592);
and AND4 (N978, N977, N833, N954, N696);
and AND2 (N979, N965, N695);
buf BUF1 (N980, N971);
not NOT1 (N981, N980);
not NOT1 (N982, N981);
or OR4 (N983, N974, N74, N613, N366);
or OR2 (N984, N967, N807);
xor XOR2 (N985, N964, N320);
and AND4 (N986, N984, N611, N717, N275);
nor NOR2 (N987, N983, N94);
and AND2 (N988, N982, N171);
nor NOR3 (N989, N985, N969, N338);
and AND4 (N990, N986, N384, N640, N757);
buf BUF1 (N991, N978);
nand NAND3 (N992, N990, N922, N8);
nor NOR4 (N993, N957, N528, N412, N63);
or OR3 (N994, N975, N535, N964);
nor NOR2 (N995, N991, N154);
xor XOR2 (N996, N993, N261);
not NOT1 (N997, N992);
and AND3 (N998, N987, N734, N575);
xor XOR2 (N999, N989, N595);
or OR4 (N1000, N973, N706, N759, N819);
not NOT1 (N1001, N998);
nand NAND4 (N1002, N996, N674, N387, N715);
buf BUF1 (N1003, N963);
buf BUF1 (N1004, N999);
buf BUF1 (N1005, N1003);
nand NAND4 (N1006, N995, N418, N927, N966);
or OR2 (N1007, N1006, N434);
or OR3 (N1008, N1001, N140, N156);
not NOT1 (N1009, N1007);
nand NAND3 (N1010, N988, N36, N682);
nor NOR2 (N1011, N997, N872);
xor XOR2 (N1012, N1009, N559);
nand NAND2 (N1013, N1008, N878);
not NOT1 (N1014, N1011);
xor XOR2 (N1015, N1013, N110);
nor NOR3 (N1016, N1015, N770, N690);
not NOT1 (N1017, N1016);
xor XOR2 (N1018, N1010, N716);
buf BUF1 (N1019, N1002);
xor XOR2 (N1020, N1018, N830);
or OR2 (N1021, N1000, N253);
nor NOR2 (N1022, N994, N821);
not NOT1 (N1023, N1019);
buf BUF1 (N1024, N1023);
nand NAND2 (N1025, N1005, N826);
xor XOR2 (N1026, N1017, N813);
not NOT1 (N1027, N1026);
nand NAND4 (N1028, N1004, N547, N372, N325);
and AND4 (N1029, N1027, N211, N827, N927);
nor NOR3 (N1030, N1014, N909, N105);
and AND3 (N1031, N1020, N608, N1015);
or OR3 (N1032, N1012, N733, N589);
or OR4 (N1033, N1022, N495, N1026, N959);
not NOT1 (N1034, N1028);
nor NOR2 (N1035, N1034, N814);
nand NAND3 (N1036, N1029, N811, N359);
and AND3 (N1037, N979, N78, N915);
or OR4 (N1038, N1036, N153, N225, N887);
xor XOR2 (N1039, N1021, N372);
nor NOR2 (N1040, N1024, N399);
not NOT1 (N1041, N1032);
nor NOR2 (N1042, N1039, N276);
and AND3 (N1043, N1025, N379, N137);
and AND2 (N1044, N1040, N324);
buf BUF1 (N1045, N1038);
or OR2 (N1046, N1043, N1025);
xor XOR2 (N1047, N1046, N317);
and AND3 (N1048, N1047, N953, N326);
and AND2 (N1049, N1045, N262);
and AND3 (N1050, N1037, N309, N1048);
nand NAND3 (N1051, N800, N230, N865);
xor XOR2 (N1052, N1031, N139);
nand NAND2 (N1053, N1033, N325);
nand NAND3 (N1054, N1049, N821, N889);
xor XOR2 (N1055, N1041, N853);
and AND3 (N1056, N1042, N870, N649);
xor XOR2 (N1057, N1050, N445);
nand NAND4 (N1058, N1052, N183, N807, N958);
not NOT1 (N1059, N1051);
nor NOR2 (N1060, N1055, N210);
nor NOR3 (N1061, N1053, N987, N1011);
not NOT1 (N1062, N1056);
xor XOR2 (N1063, N1044, N282);
nand NAND4 (N1064, N1057, N798, N373, N220);
and AND4 (N1065, N1035, N497, N545, N656);
or OR4 (N1066, N1054, N89, N217, N492);
buf BUF1 (N1067, N1065);
not NOT1 (N1068, N1066);
not NOT1 (N1069, N1058);
xor XOR2 (N1070, N1068, N619);
nor NOR4 (N1071, N1064, N780, N60, N542);
nor NOR4 (N1072, N1063, N283, N934, N550);
not NOT1 (N1073, N1072);
or OR4 (N1074, N1073, N899, N708, N405);
buf BUF1 (N1075, N1059);
or OR4 (N1076, N1071, N412, N361, N477);
and AND4 (N1077, N1030, N343, N828, N459);
nor NOR4 (N1078, N1075, N83, N563, N265);
and AND4 (N1079, N1077, N999, N424, N490);
and AND4 (N1080, N1069, N84, N335, N873);
buf BUF1 (N1081, N1067);
nor NOR3 (N1082, N1061, N905, N676);
xor XOR2 (N1083, N1081, N1076);
and AND2 (N1084, N1023, N947);
not NOT1 (N1085, N1082);
buf BUF1 (N1086, N1085);
nand NAND3 (N1087, N1083, N317, N904);
buf BUF1 (N1088, N1078);
nand NAND2 (N1089, N1086, N752);
buf BUF1 (N1090, N1070);
buf BUF1 (N1091, N1080);
not NOT1 (N1092, N1088);
nor NOR2 (N1093, N1087, N188);
nor NOR4 (N1094, N1079, N969, N68, N161);
or OR2 (N1095, N1093, N78);
and AND3 (N1096, N1084, N25, N408);
buf BUF1 (N1097, N1060);
or OR2 (N1098, N1096, N400);
or OR4 (N1099, N1074, N331, N941, N282);
nand NAND3 (N1100, N1089, N929, N22);
and AND4 (N1101, N1092, N244, N539, N854);
not NOT1 (N1102, N1090);
buf BUF1 (N1103, N1102);
nor NOR2 (N1104, N1095, N978);
or OR2 (N1105, N1101, N577);
and AND3 (N1106, N1104, N1051, N148);
or OR4 (N1107, N1094, N184, N389, N1096);
not NOT1 (N1108, N1105);
nand NAND2 (N1109, N1108, N923);
not NOT1 (N1110, N1062);
or OR3 (N1111, N1099, N569, N841);
xor XOR2 (N1112, N1109, N1046);
nor NOR4 (N1113, N1091, N937, N910, N810);
or OR4 (N1114, N1107, N30, N310, N342);
not NOT1 (N1115, N1111);
not NOT1 (N1116, N1113);
xor XOR2 (N1117, N1103, N167);
buf BUF1 (N1118, N1110);
nor NOR4 (N1119, N1114, N385, N674, N837);
buf BUF1 (N1120, N1117);
not NOT1 (N1121, N1115);
buf BUF1 (N1122, N1120);
not NOT1 (N1123, N1112);
or OR3 (N1124, N1106, N300, N922);
and AND3 (N1125, N1124, N48, N838);
not NOT1 (N1126, N1098);
buf BUF1 (N1127, N1119);
nor NOR2 (N1128, N1100, N625);
not NOT1 (N1129, N1122);
nor NOR4 (N1130, N1121, N1103, N634, N639);
xor XOR2 (N1131, N1129, N940);
nand NAND4 (N1132, N1118, N1050, N699, N470);
or OR4 (N1133, N1130, N353, N128, N90);
xor XOR2 (N1134, N1097, N552);
xor XOR2 (N1135, N1123, N805);
and AND3 (N1136, N1126, N127, N466);
not NOT1 (N1137, N1127);
nand NAND4 (N1138, N1136, N496, N274, N190);
not NOT1 (N1139, N1131);
or OR2 (N1140, N1133, N814);
not NOT1 (N1141, N1139);
buf BUF1 (N1142, N1128);
and AND2 (N1143, N1137, N639);
or OR2 (N1144, N1142, N269);
not NOT1 (N1145, N1135);
nor NOR2 (N1146, N1145, N462);
xor XOR2 (N1147, N1144, N1125);
nand NAND3 (N1148, N436, N618, N157);
or OR4 (N1149, N1146, N693, N205, N219);
nand NAND3 (N1150, N1134, N624, N197);
xor XOR2 (N1151, N1147, N706);
nor NOR2 (N1152, N1141, N324);
not NOT1 (N1153, N1152);
xor XOR2 (N1154, N1151, N841);
nor NOR2 (N1155, N1153, N478);
xor XOR2 (N1156, N1154, N897);
or OR4 (N1157, N1148, N800, N34, N928);
nand NAND3 (N1158, N1157, N705, N1133);
buf BUF1 (N1159, N1138);
nand NAND2 (N1160, N1155, N287);
nand NAND4 (N1161, N1150, N749, N586, N749);
and AND4 (N1162, N1158, N462, N39, N859);
or OR2 (N1163, N1116, N473);
or OR4 (N1164, N1161, N258, N599, N355);
or OR2 (N1165, N1132, N65);
not NOT1 (N1166, N1156);
buf BUF1 (N1167, N1149);
nand NAND4 (N1168, N1140, N265, N55, N189);
not NOT1 (N1169, N1164);
xor XOR2 (N1170, N1159, N391);
not NOT1 (N1171, N1167);
xor XOR2 (N1172, N1169, N138);
nor NOR3 (N1173, N1170, N175, N526);
not NOT1 (N1174, N1143);
not NOT1 (N1175, N1160);
nand NAND3 (N1176, N1172, N948, N1110);
nor NOR4 (N1177, N1173, N1122, N548, N1094);
nor NOR2 (N1178, N1165, N1089);
not NOT1 (N1179, N1168);
nor NOR3 (N1180, N1162, N945, N611);
xor XOR2 (N1181, N1175, N1119);
buf BUF1 (N1182, N1179);
xor XOR2 (N1183, N1177, N913);
buf BUF1 (N1184, N1180);
xor XOR2 (N1185, N1176, N22);
buf BUF1 (N1186, N1178);
nor NOR4 (N1187, N1182, N774, N985, N554);
nand NAND4 (N1188, N1163, N365, N1047, N889);
and AND3 (N1189, N1186, N552, N208);
nor NOR2 (N1190, N1174, N1173);
and AND2 (N1191, N1171, N964);
not NOT1 (N1192, N1188);
nor NOR4 (N1193, N1191, N356, N1125, N732);
not NOT1 (N1194, N1181);
xor XOR2 (N1195, N1183, N750);
not NOT1 (N1196, N1194);
or OR2 (N1197, N1189, N478);
not NOT1 (N1198, N1196);
or OR3 (N1199, N1190, N426, N885);
nor NOR2 (N1200, N1187, N688);
or OR2 (N1201, N1195, N377);
not NOT1 (N1202, N1184);
nor NOR2 (N1203, N1185, N1051);
xor XOR2 (N1204, N1197, N559);
or OR3 (N1205, N1200, N154, N635);
and AND4 (N1206, N1203, N411, N769, N853);
nor NOR4 (N1207, N1199, N1014, N525, N853);
or OR2 (N1208, N1192, N228);
not NOT1 (N1209, N1207);
nor NOR4 (N1210, N1204, N512, N1105, N944);
and AND2 (N1211, N1202, N913);
or OR3 (N1212, N1166, N1078, N515);
not NOT1 (N1213, N1193);
not NOT1 (N1214, N1201);
nand NAND2 (N1215, N1198, N1116);
xor XOR2 (N1216, N1208, N1114);
not NOT1 (N1217, N1205);
not NOT1 (N1218, N1214);
nor NOR4 (N1219, N1210, N1167, N525, N99);
nor NOR2 (N1220, N1206, N295);
nand NAND3 (N1221, N1209, N304, N21);
nand NAND2 (N1222, N1219, N1139);
xor XOR2 (N1223, N1218, N153);
or OR4 (N1224, N1220, N559, N149, N582);
or OR4 (N1225, N1213, N63, N1203, N1183);
and AND3 (N1226, N1224, N579, N720);
buf BUF1 (N1227, N1225);
and AND2 (N1228, N1216, N785);
nor NOR2 (N1229, N1228, N616);
or OR4 (N1230, N1223, N1030, N77, N941);
nor NOR4 (N1231, N1211, N358, N1032, N1049);
not NOT1 (N1232, N1227);
xor XOR2 (N1233, N1215, N163);
nand NAND4 (N1234, N1221, N19, N433, N686);
or OR4 (N1235, N1231, N665, N458, N809);
or OR3 (N1236, N1230, N680, N620);
nor NOR2 (N1237, N1236, N893);
and AND2 (N1238, N1226, N994);
buf BUF1 (N1239, N1234);
nand NAND2 (N1240, N1238, N597);
and AND4 (N1241, N1232, N237, N145, N929);
and AND4 (N1242, N1222, N546, N74, N843);
and AND3 (N1243, N1217, N566, N120);
xor XOR2 (N1244, N1242, N314);
and AND4 (N1245, N1212, N415, N247, N798);
xor XOR2 (N1246, N1244, N829);
and AND4 (N1247, N1246, N859, N199, N36);
xor XOR2 (N1248, N1237, N332);
buf BUF1 (N1249, N1235);
buf BUF1 (N1250, N1249);
and AND4 (N1251, N1240, N765, N782, N853);
xor XOR2 (N1252, N1245, N851);
xor XOR2 (N1253, N1252, N647);
and AND3 (N1254, N1233, N1237, N291);
and AND3 (N1255, N1239, N1001, N500);
and AND2 (N1256, N1253, N648);
or OR2 (N1257, N1251, N273);
nand NAND2 (N1258, N1243, N220);
nand NAND4 (N1259, N1256, N997, N1124, N1159);
buf BUF1 (N1260, N1258);
buf BUF1 (N1261, N1229);
buf BUF1 (N1262, N1257);
nor NOR4 (N1263, N1260, N304, N99, N627);
xor XOR2 (N1264, N1254, N1149);
xor XOR2 (N1265, N1248, N799);
xor XOR2 (N1266, N1250, N594);
nand NAND3 (N1267, N1262, N342, N809);
not NOT1 (N1268, N1255);
nand NAND2 (N1269, N1261, N508);
and AND4 (N1270, N1247, N1115, N99, N722);
not NOT1 (N1271, N1266);
nand NAND2 (N1272, N1271, N1068);
and AND2 (N1273, N1267, N7);
buf BUF1 (N1274, N1264);
nor NOR3 (N1275, N1241, N862, N731);
xor XOR2 (N1276, N1259, N771);
xor XOR2 (N1277, N1276, N779);
xor XOR2 (N1278, N1277, N940);
and AND3 (N1279, N1263, N750, N551);
buf BUF1 (N1280, N1269);
nor NOR2 (N1281, N1274, N292);
buf BUF1 (N1282, N1270);
buf BUF1 (N1283, N1265);
and AND3 (N1284, N1279, N643, N1113);
and AND2 (N1285, N1273, N1028);
xor XOR2 (N1286, N1282, N269);
or OR2 (N1287, N1286, N93);
nor NOR2 (N1288, N1280, N1242);
xor XOR2 (N1289, N1287, N1154);
not NOT1 (N1290, N1268);
nor NOR2 (N1291, N1288, N200);
nor NOR2 (N1292, N1278, N1212);
not NOT1 (N1293, N1292);
buf BUF1 (N1294, N1272);
nand NAND2 (N1295, N1281, N1161);
not NOT1 (N1296, N1284);
nand NAND4 (N1297, N1296, N1118, N892, N1125);
buf BUF1 (N1298, N1285);
nor NOR2 (N1299, N1291, N245);
buf BUF1 (N1300, N1293);
nor NOR2 (N1301, N1295, N883);
buf BUF1 (N1302, N1299);
and AND2 (N1303, N1289, N1198);
nor NOR4 (N1304, N1294, N585, N931, N715);
buf BUF1 (N1305, N1300);
xor XOR2 (N1306, N1298, N976);
xor XOR2 (N1307, N1283, N896);
not NOT1 (N1308, N1307);
nand NAND4 (N1309, N1297, N424, N965, N584);
not NOT1 (N1310, N1304);
or OR4 (N1311, N1275, N638, N22, N386);
buf BUF1 (N1312, N1302);
nand NAND3 (N1313, N1312, N1014, N1140);
not NOT1 (N1314, N1308);
xor XOR2 (N1315, N1310, N819);
buf BUF1 (N1316, N1290);
and AND2 (N1317, N1303, N1058);
nor NOR2 (N1318, N1305, N1128);
or OR3 (N1319, N1306, N568, N48);
xor XOR2 (N1320, N1311, N250);
nand NAND2 (N1321, N1318, N134);
nand NAND2 (N1322, N1301, N384);
or OR3 (N1323, N1317, N817, N365);
nand NAND4 (N1324, N1309, N1139, N1200, N1105);
nand NAND4 (N1325, N1316, N1202, N685, N976);
nor NOR4 (N1326, N1322, N1189, N1127, N992);
buf BUF1 (N1327, N1315);
xor XOR2 (N1328, N1327, N91);
xor XOR2 (N1329, N1314, N456);
and AND2 (N1330, N1320, N280);
xor XOR2 (N1331, N1313, N500);
and AND2 (N1332, N1324, N459);
and AND3 (N1333, N1329, N1220, N388);
nor NOR4 (N1334, N1326, N171, N955, N60);
and AND3 (N1335, N1323, N636, N265);
or OR3 (N1336, N1332, N959, N120);
and AND4 (N1337, N1334, N855, N963, N1253);
not NOT1 (N1338, N1319);
or OR2 (N1339, N1337, N138);
nor NOR3 (N1340, N1325, N594, N1142);
or OR2 (N1341, N1328, N298);
not NOT1 (N1342, N1321);
xor XOR2 (N1343, N1338, N1037);
xor XOR2 (N1344, N1336, N243);
nand NAND4 (N1345, N1344, N718, N345, N719);
and AND3 (N1346, N1340, N694, N324);
xor XOR2 (N1347, N1342, N344);
or OR4 (N1348, N1341, N226, N241, N341);
nor NOR4 (N1349, N1330, N393, N362, N127);
nor NOR4 (N1350, N1347, N1236, N44, N1004);
or OR4 (N1351, N1345, N40, N839, N796);
xor XOR2 (N1352, N1350, N883);
or OR3 (N1353, N1346, N1073, N925);
buf BUF1 (N1354, N1339);
nor NOR4 (N1355, N1333, N1240, N963, N819);
or OR3 (N1356, N1353, N1145, N893);
or OR3 (N1357, N1348, N1033, N795);
and AND4 (N1358, N1357, N1145, N260, N141);
nand NAND3 (N1359, N1335, N1135, N1125);
nor NOR4 (N1360, N1349, N1152, N615, N1056);
or OR3 (N1361, N1354, N865, N28);
nand NAND2 (N1362, N1355, N386);
xor XOR2 (N1363, N1352, N471);
nor NOR3 (N1364, N1358, N947, N794);
not NOT1 (N1365, N1363);
nand NAND3 (N1366, N1331, N709, N1343);
and AND3 (N1367, N1042, N676, N880);
xor XOR2 (N1368, N1367, N243);
buf BUF1 (N1369, N1359);
buf BUF1 (N1370, N1351);
buf BUF1 (N1371, N1362);
or OR4 (N1372, N1371, N1337, N632, N1218);
nor NOR3 (N1373, N1365, N23, N1033);
nor NOR2 (N1374, N1366, N1106);
nor NOR2 (N1375, N1374, N1283);
xor XOR2 (N1376, N1360, N3);
and AND4 (N1377, N1368, N52, N86, N787);
buf BUF1 (N1378, N1361);
not NOT1 (N1379, N1370);
and AND2 (N1380, N1369, N175);
or OR2 (N1381, N1376, N1283);
buf BUF1 (N1382, N1380);
and AND3 (N1383, N1381, N38, N412);
or OR3 (N1384, N1356, N200, N128);
xor XOR2 (N1385, N1383, N1265);
buf BUF1 (N1386, N1372);
nor NOR3 (N1387, N1364, N1066, N142);
or OR2 (N1388, N1377, N1170);
and AND2 (N1389, N1384, N396);
and AND4 (N1390, N1375, N606, N173, N254);
nand NAND3 (N1391, N1389, N695, N887);
nand NAND4 (N1392, N1386, N1020, N1026, N1058);
nor NOR2 (N1393, N1392, N487);
xor XOR2 (N1394, N1391, N887);
nand NAND2 (N1395, N1382, N480);
buf BUF1 (N1396, N1394);
nand NAND4 (N1397, N1385, N360, N1290, N5);
or OR2 (N1398, N1393, N574);
xor XOR2 (N1399, N1396, N1131);
or OR4 (N1400, N1395, N930, N1363, N697);
nor NOR2 (N1401, N1373, N1063);
and AND2 (N1402, N1401, N1223);
xor XOR2 (N1403, N1400, N1098);
nor NOR4 (N1404, N1388, N1347, N748, N662);
nor NOR2 (N1405, N1399, N452);
nand NAND4 (N1406, N1397, N1124, N1008, N1050);
not NOT1 (N1407, N1378);
buf BUF1 (N1408, N1402);
or OR3 (N1409, N1398, N1013, N444);
or OR2 (N1410, N1390, N1276);
xor XOR2 (N1411, N1405, N391);
buf BUF1 (N1412, N1406);
and AND4 (N1413, N1403, N268, N1345, N1371);
xor XOR2 (N1414, N1404, N485);
and AND2 (N1415, N1387, N272);
and AND4 (N1416, N1409, N1057, N1387, N1393);
or OR4 (N1417, N1379, N902, N304, N178);
xor XOR2 (N1418, N1416, N847);
nand NAND3 (N1419, N1407, N1223, N951);
not NOT1 (N1420, N1412);
nand NAND3 (N1421, N1411, N409, N193);
nor NOR3 (N1422, N1418, N210, N52);
nand NAND3 (N1423, N1420, N578, N662);
xor XOR2 (N1424, N1419, N991);
nor NOR2 (N1425, N1424, N1011);
nor NOR2 (N1426, N1410, N1405);
nor NOR2 (N1427, N1423, N533);
nand NAND2 (N1428, N1421, N589);
and AND4 (N1429, N1413, N1064, N1381, N1303);
not NOT1 (N1430, N1417);
buf BUF1 (N1431, N1430);
nand NAND2 (N1432, N1422, N408);
or OR4 (N1433, N1414, N822, N684, N971);
or OR3 (N1434, N1427, N839, N499);
and AND2 (N1435, N1415, N1210);
and AND3 (N1436, N1434, N384, N111);
and AND3 (N1437, N1431, N891, N808);
nand NAND4 (N1438, N1428, N970, N1398, N16);
buf BUF1 (N1439, N1435);
or OR4 (N1440, N1432, N445, N1232, N392);
nand NAND3 (N1441, N1437, N1379, N138);
not NOT1 (N1442, N1441);
nand NAND4 (N1443, N1429, N353, N1186, N1011);
and AND2 (N1444, N1442, N1302);
xor XOR2 (N1445, N1426, N638);
not NOT1 (N1446, N1433);
or OR3 (N1447, N1446, N623, N1207);
or OR3 (N1448, N1444, N457, N1160);
nand NAND2 (N1449, N1436, N550);
nor NOR3 (N1450, N1408, N133, N625);
nor NOR2 (N1451, N1450, N797);
buf BUF1 (N1452, N1449);
nor NOR4 (N1453, N1438, N616, N574, N521);
and AND4 (N1454, N1439, N1093, N865, N599);
or OR2 (N1455, N1451, N308);
xor XOR2 (N1456, N1447, N1431);
not NOT1 (N1457, N1448);
nor NOR4 (N1458, N1453, N704, N1274, N141);
buf BUF1 (N1459, N1452);
buf BUF1 (N1460, N1457);
nand NAND3 (N1461, N1455, N923, N230);
buf BUF1 (N1462, N1454);
or OR3 (N1463, N1456, N841, N454);
xor XOR2 (N1464, N1440, N64);
and AND4 (N1465, N1464, N1230, N916, N1148);
nor NOR3 (N1466, N1461, N1369, N11);
buf BUF1 (N1467, N1445);
and AND3 (N1468, N1462, N1071, N690);
xor XOR2 (N1469, N1443, N1071);
nand NAND4 (N1470, N1459, N1135, N1443, N648);
or OR4 (N1471, N1425, N1064, N1378, N509);
xor XOR2 (N1472, N1470, N368);
not NOT1 (N1473, N1468);
xor XOR2 (N1474, N1458, N269);
not NOT1 (N1475, N1472);
and AND2 (N1476, N1473, N989);
buf BUF1 (N1477, N1467);
nand NAND3 (N1478, N1469, N1155, N37);
xor XOR2 (N1479, N1460, N1305);
not NOT1 (N1480, N1479);
nor NOR4 (N1481, N1475, N671, N695, N1336);
or OR3 (N1482, N1476, N686, N718);
nor NOR3 (N1483, N1477, N1124, N1103);
not NOT1 (N1484, N1482);
nor NOR2 (N1485, N1471, N243);
and AND2 (N1486, N1465, N20);
or OR3 (N1487, N1480, N549, N135);
or OR3 (N1488, N1478, N817, N1149);
and AND3 (N1489, N1485, N1211, N1425);
not NOT1 (N1490, N1463);
xor XOR2 (N1491, N1484, N235);
nor NOR2 (N1492, N1488, N1413);
xor XOR2 (N1493, N1486, N498);
and AND2 (N1494, N1466, N1382);
buf BUF1 (N1495, N1494);
xor XOR2 (N1496, N1492, N287);
buf BUF1 (N1497, N1489);
or OR3 (N1498, N1495, N778, N857);
nand NAND3 (N1499, N1483, N26, N844);
not NOT1 (N1500, N1497);
or OR3 (N1501, N1499, N112, N310);
buf BUF1 (N1502, N1491);
nor NOR4 (N1503, N1502, N971, N163, N872);
not NOT1 (N1504, N1481);
buf BUF1 (N1505, N1498);
and AND4 (N1506, N1503, N962, N15, N1442);
or OR2 (N1507, N1496, N1470);
and AND4 (N1508, N1507, N295, N218, N93);
not NOT1 (N1509, N1490);
or OR4 (N1510, N1509, N29, N873, N946);
or OR4 (N1511, N1504, N786, N68, N518);
nand NAND4 (N1512, N1501, N1291, N159, N1);
and AND3 (N1513, N1511, N1326, N734);
not NOT1 (N1514, N1505);
nor NOR3 (N1515, N1487, N951, N744);
nand NAND2 (N1516, N1500, N561);
nor NOR2 (N1517, N1514, N542);
nand NAND2 (N1518, N1512, N910);
not NOT1 (N1519, N1506);
nand NAND2 (N1520, N1510, N828);
not NOT1 (N1521, N1515);
buf BUF1 (N1522, N1520);
not NOT1 (N1523, N1516);
xor XOR2 (N1524, N1518, N781);
and AND3 (N1525, N1523, N1047, N941);
or OR2 (N1526, N1474, N164);
xor XOR2 (N1527, N1522, N35);
buf BUF1 (N1528, N1525);
nor NOR4 (N1529, N1528, N33, N1528, N55);
nor NOR4 (N1530, N1493, N260, N39, N193);
or OR3 (N1531, N1519, N995, N568);
not NOT1 (N1532, N1508);
nand NAND3 (N1533, N1527, N1100, N1168);
nand NAND3 (N1534, N1533, N1231, N789);
xor XOR2 (N1535, N1526, N567);
xor XOR2 (N1536, N1532, N960);
buf BUF1 (N1537, N1513);
nor NOR2 (N1538, N1535, N567);
and AND3 (N1539, N1521, N996, N1479);
nand NAND3 (N1540, N1530, N434, N708);
buf BUF1 (N1541, N1531);
or OR3 (N1542, N1529, N342, N1000);
nand NAND3 (N1543, N1517, N446, N415);
nand NAND2 (N1544, N1524, N1030);
buf BUF1 (N1545, N1539);
nand NAND4 (N1546, N1536, N162, N455, N310);
or OR3 (N1547, N1537, N170, N1244);
and AND4 (N1548, N1546, N554, N26, N888);
buf BUF1 (N1549, N1540);
nor NOR2 (N1550, N1541, N635);
and AND2 (N1551, N1548, N1106);
and AND2 (N1552, N1544, N392);
nor NOR2 (N1553, N1550, N1490);
not NOT1 (N1554, N1538);
and AND2 (N1555, N1543, N905);
or OR3 (N1556, N1547, N1291, N1472);
not NOT1 (N1557, N1556);
nor NOR2 (N1558, N1542, N1106);
nand NAND4 (N1559, N1558, N1156, N1333, N550);
nand NAND2 (N1560, N1534, N1373);
nor NOR2 (N1561, N1545, N247);
buf BUF1 (N1562, N1561);
nor NOR3 (N1563, N1551, N41, N1393);
and AND3 (N1564, N1549, N795, N185);
and AND3 (N1565, N1552, N67, N450);
and AND2 (N1566, N1559, N818);
buf BUF1 (N1567, N1564);
nor NOR4 (N1568, N1563, N208, N1086, N1476);
and AND4 (N1569, N1566, N571, N677, N1386);
not NOT1 (N1570, N1555);
nand NAND4 (N1571, N1553, N905, N912, N458);
and AND2 (N1572, N1567, N940);
xor XOR2 (N1573, N1571, N1028);
nor NOR4 (N1574, N1565, N546, N1300, N359);
not NOT1 (N1575, N1562);
buf BUF1 (N1576, N1569);
or OR4 (N1577, N1568, N47, N940, N805);
or OR2 (N1578, N1575, N422);
xor XOR2 (N1579, N1572, N1514);
and AND2 (N1580, N1573, N505);
buf BUF1 (N1581, N1554);
not NOT1 (N1582, N1570);
xor XOR2 (N1583, N1576, N147);
nor NOR3 (N1584, N1557, N1536, N932);
nor NOR4 (N1585, N1578, N1528, N370, N573);
nor NOR2 (N1586, N1584, N831);
or OR4 (N1587, N1580, N1025, N703, N651);
or OR2 (N1588, N1583, N308);
buf BUF1 (N1589, N1579);
not NOT1 (N1590, N1587);
or OR2 (N1591, N1588, N321);
nor NOR3 (N1592, N1590, N1450, N1478);
not NOT1 (N1593, N1582);
xor XOR2 (N1594, N1593, N35);
not NOT1 (N1595, N1592);
xor XOR2 (N1596, N1591, N1574);
or OR2 (N1597, N1543, N909);
not NOT1 (N1598, N1596);
nor NOR3 (N1599, N1581, N677, N864);
buf BUF1 (N1600, N1577);
not NOT1 (N1601, N1597);
not NOT1 (N1602, N1600);
not NOT1 (N1603, N1602);
xor XOR2 (N1604, N1585, N927);
xor XOR2 (N1605, N1598, N1388);
xor XOR2 (N1606, N1603, N1426);
xor XOR2 (N1607, N1599, N920);
nand NAND3 (N1608, N1601, N1533, N486);
buf BUF1 (N1609, N1560);
and AND4 (N1610, N1609, N938, N1350, N27);
nand NAND3 (N1611, N1604, N193, N660);
and AND2 (N1612, N1608, N450);
or OR3 (N1613, N1611, N1281, N689);
nor NOR3 (N1614, N1605, N880, N106);
xor XOR2 (N1615, N1586, N607);
or OR2 (N1616, N1606, N1077);
and AND3 (N1617, N1614, N1372, N1110);
buf BUF1 (N1618, N1616);
nor NOR4 (N1619, N1594, N1511, N331, N387);
nor NOR3 (N1620, N1613, N871, N841);
xor XOR2 (N1621, N1607, N1338);
or OR3 (N1622, N1621, N1428, N236);
buf BUF1 (N1623, N1612);
nor NOR3 (N1624, N1622, N1460, N1490);
nor NOR3 (N1625, N1620, N1564, N706);
or OR3 (N1626, N1624, N729, N1584);
xor XOR2 (N1627, N1626, N805);
or OR3 (N1628, N1617, N1448, N1009);
or OR3 (N1629, N1625, N889, N536);
nor NOR3 (N1630, N1615, N1161, N467);
or OR2 (N1631, N1628, N326);
nor NOR4 (N1632, N1623, N1151, N936, N172);
nand NAND3 (N1633, N1610, N586, N1383);
nand NAND3 (N1634, N1595, N1550, N912);
or OR3 (N1635, N1619, N1174, N404);
or OR4 (N1636, N1629, N1166, N229, N667);
or OR2 (N1637, N1633, N972);
buf BUF1 (N1638, N1632);
and AND4 (N1639, N1631, N641, N1400, N624);
or OR3 (N1640, N1630, N937, N1460);
xor XOR2 (N1641, N1638, N1375);
nor NOR4 (N1642, N1639, N194, N1361, N1618);
nand NAND2 (N1643, N452, N1304);
xor XOR2 (N1644, N1641, N1563);
nand NAND4 (N1645, N1627, N418, N1268, N204);
and AND3 (N1646, N1643, N679, N627);
not NOT1 (N1647, N1636);
buf BUF1 (N1648, N1646);
and AND4 (N1649, N1637, N1469, N1476, N8);
not NOT1 (N1650, N1648);
not NOT1 (N1651, N1645);
buf BUF1 (N1652, N1651);
or OR2 (N1653, N1649, N853);
or OR3 (N1654, N1642, N1542, N1632);
nand NAND3 (N1655, N1647, N1024, N821);
xor XOR2 (N1656, N1589, N1199);
nor NOR2 (N1657, N1644, N74);
not NOT1 (N1658, N1655);
or OR2 (N1659, N1656, N92);
and AND4 (N1660, N1654, N1176, N442, N1236);
or OR2 (N1661, N1650, N428);
not NOT1 (N1662, N1660);
buf BUF1 (N1663, N1657);
xor XOR2 (N1664, N1640, N833);
or OR4 (N1665, N1658, N1008, N71, N49);
buf BUF1 (N1666, N1664);
buf BUF1 (N1667, N1634);
buf BUF1 (N1668, N1665);
not NOT1 (N1669, N1661);
nand NAND2 (N1670, N1667, N1534);
and AND3 (N1671, N1668, N1387, N187);
and AND3 (N1672, N1662, N448, N125);
nand NAND4 (N1673, N1671, N1020, N834, N822);
xor XOR2 (N1674, N1666, N1225);
xor XOR2 (N1675, N1673, N1252);
buf BUF1 (N1676, N1670);
nand NAND3 (N1677, N1653, N589, N1630);
and AND4 (N1678, N1676, N940, N1421, N43);
nor NOR4 (N1679, N1675, N1518, N1187, N73);
not NOT1 (N1680, N1679);
nor NOR2 (N1681, N1635, N1380);
xor XOR2 (N1682, N1677, N797);
nand NAND4 (N1683, N1669, N1224, N430, N1113);
buf BUF1 (N1684, N1652);
buf BUF1 (N1685, N1672);
not NOT1 (N1686, N1663);
buf BUF1 (N1687, N1685);
and AND2 (N1688, N1682, N1472);
and AND2 (N1689, N1688, N1078);
xor XOR2 (N1690, N1678, N126);
nor NOR2 (N1691, N1681, N1670);
not NOT1 (N1692, N1686);
nand NAND4 (N1693, N1674, N552, N1142, N1464);
or OR3 (N1694, N1690, N48, N919);
and AND3 (N1695, N1689, N158, N385);
buf BUF1 (N1696, N1680);
buf BUF1 (N1697, N1684);
not NOT1 (N1698, N1694);
xor XOR2 (N1699, N1696, N339);
not NOT1 (N1700, N1687);
xor XOR2 (N1701, N1683, N594);
nor NOR4 (N1702, N1699, N1001, N994, N937);
xor XOR2 (N1703, N1692, N1168);
nand NAND3 (N1704, N1697, N80, N428);
xor XOR2 (N1705, N1698, N1615);
not NOT1 (N1706, N1700);
and AND4 (N1707, N1705, N105, N477, N1301);
nor NOR3 (N1708, N1659, N1304, N570);
or OR2 (N1709, N1695, N1608);
nand NAND2 (N1710, N1701, N566);
nor NOR4 (N1711, N1710, N1379, N14, N503);
buf BUF1 (N1712, N1711);
buf BUF1 (N1713, N1708);
buf BUF1 (N1714, N1706);
and AND4 (N1715, N1693, N1377, N67, N1701);
nand NAND3 (N1716, N1712, N1240, N972);
nor NOR3 (N1717, N1713, N1343, N539);
or OR2 (N1718, N1714, N1329);
nor NOR3 (N1719, N1703, N727, N1424);
nand NAND4 (N1720, N1717, N1266, N899, N1337);
buf BUF1 (N1721, N1720);
or OR2 (N1722, N1719, N399);
or OR3 (N1723, N1721, N1411, N318);
nor NOR4 (N1724, N1715, N667, N734, N1180);
buf BUF1 (N1725, N1716);
xor XOR2 (N1726, N1724, N1605);
nor NOR3 (N1727, N1702, N318, N842);
nand NAND3 (N1728, N1726, N906, N1653);
nand NAND3 (N1729, N1718, N814, N80);
buf BUF1 (N1730, N1727);
nand NAND2 (N1731, N1704, N1388);
not NOT1 (N1732, N1707);
nor NOR2 (N1733, N1730, N1580);
not NOT1 (N1734, N1723);
xor XOR2 (N1735, N1734, N1654);
xor XOR2 (N1736, N1735, N511);
buf BUF1 (N1737, N1728);
and AND2 (N1738, N1733, N974);
buf BUF1 (N1739, N1736);
nand NAND4 (N1740, N1739, N803, N964, N1199);
or OR4 (N1741, N1737, N1245, N1225, N66);
buf BUF1 (N1742, N1732);
nor NOR3 (N1743, N1722, N128, N545);
xor XOR2 (N1744, N1740, N253);
nand NAND2 (N1745, N1709, N412);
or OR2 (N1746, N1738, N1268);
nand NAND4 (N1747, N1743, N869, N405, N369);
xor XOR2 (N1748, N1725, N1222);
not NOT1 (N1749, N1729);
xor XOR2 (N1750, N1745, N965);
and AND3 (N1751, N1731, N647, N372);
or OR4 (N1752, N1742, N1007, N1686, N1169);
nand NAND3 (N1753, N1744, N1582, N161);
not NOT1 (N1754, N1691);
or OR2 (N1755, N1753, N955);
nor NOR3 (N1756, N1752, N404, N270);
xor XOR2 (N1757, N1746, N571);
buf BUF1 (N1758, N1755);
nand NAND4 (N1759, N1748, N386, N773, N151);
and AND2 (N1760, N1757, N1713);
or OR3 (N1761, N1749, N636, N1478);
nand NAND3 (N1762, N1760, N296, N893);
or OR3 (N1763, N1741, N1513, N68);
nand NAND2 (N1764, N1747, N1535);
nor NOR4 (N1765, N1761, N1072, N508, N785);
not NOT1 (N1766, N1763);
nand NAND4 (N1767, N1759, N1145, N498, N428);
or OR2 (N1768, N1767, N1559);
or OR3 (N1769, N1758, N1381, N361);
and AND3 (N1770, N1754, N1652, N1341);
buf BUF1 (N1771, N1756);
or OR2 (N1772, N1751, N1469);
and AND4 (N1773, N1766, N1616, N636, N48);
not NOT1 (N1774, N1768);
nand NAND2 (N1775, N1771, N760);
and AND4 (N1776, N1773, N29, N1567, N1046);
xor XOR2 (N1777, N1762, N715);
or OR4 (N1778, N1774, N1706, N258, N1150);
nand NAND2 (N1779, N1764, N1639);
xor XOR2 (N1780, N1775, N54);
not NOT1 (N1781, N1780);
xor XOR2 (N1782, N1779, N778);
and AND4 (N1783, N1782, N277, N1353, N731);
nand NAND2 (N1784, N1776, N776);
nand NAND2 (N1785, N1777, N812);
and AND2 (N1786, N1750, N1104);
nand NAND4 (N1787, N1769, N23, N1268, N1108);
buf BUF1 (N1788, N1781);
or OR4 (N1789, N1785, N417, N1690, N397);
xor XOR2 (N1790, N1783, N269);
nand NAND2 (N1791, N1784, N1307);
and AND4 (N1792, N1789, N1188, N375, N198);
buf BUF1 (N1793, N1788);
and AND4 (N1794, N1791, N1743, N926, N1724);
or OR4 (N1795, N1786, N1083, N1391, N1316);
nor NOR3 (N1796, N1778, N1252, N935);
and AND4 (N1797, N1796, N1414, N1233, N640);
xor XOR2 (N1798, N1772, N629);
or OR2 (N1799, N1795, N528);
nor NOR3 (N1800, N1790, N1406, N775);
nor NOR3 (N1801, N1770, N1059, N1075);
xor XOR2 (N1802, N1801, N781);
or OR2 (N1803, N1797, N1229);
nand NAND4 (N1804, N1792, N753, N591, N1324);
xor XOR2 (N1805, N1802, N1652);
nor NOR3 (N1806, N1787, N1255, N1070);
xor XOR2 (N1807, N1805, N95);
nor NOR3 (N1808, N1794, N666, N788);
or OR4 (N1809, N1765, N1199, N1483, N90);
nand NAND3 (N1810, N1798, N657, N1389);
nor NOR2 (N1811, N1810, N423);
and AND3 (N1812, N1807, N1044, N728);
nor NOR2 (N1813, N1812, N1757);
xor XOR2 (N1814, N1808, N1673);
or OR4 (N1815, N1800, N1586, N566, N701);
xor XOR2 (N1816, N1806, N95);
xor XOR2 (N1817, N1811, N963);
and AND4 (N1818, N1814, N1592, N941, N1020);
and AND3 (N1819, N1793, N1503, N244);
and AND3 (N1820, N1816, N1440, N928);
buf BUF1 (N1821, N1803);
not NOT1 (N1822, N1817);
not NOT1 (N1823, N1804);
not NOT1 (N1824, N1820);
nor NOR3 (N1825, N1809, N177, N165);
buf BUF1 (N1826, N1819);
nor NOR3 (N1827, N1821, N1561, N1396);
not NOT1 (N1828, N1815);
or OR3 (N1829, N1818, N400, N347);
nand NAND4 (N1830, N1829, N165, N6, N102);
xor XOR2 (N1831, N1827, N1141);
nand NAND2 (N1832, N1824, N1623);
buf BUF1 (N1833, N1823);
buf BUF1 (N1834, N1831);
and AND3 (N1835, N1822, N1421, N441);
not NOT1 (N1836, N1835);
nor NOR2 (N1837, N1826, N1019);
xor XOR2 (N1838, N1834, N139);
and AND3 (N1839, N1833, N1370, N233);
not NOT1 (N1840, N1838);
nor NOR2 (N1841, N1830, N108);
xor XOR2 (N1842, N1840, N1550);
and AND2 (N1843, N1825, N939);
or OR4 (N1844, N1839, N263, N558, N745);
and AND4 (N1845, N1813, N65, N1727, N256);
nor NOR4 (N1846, N1844, N554, N680, N1616);
and AND4 (N1847, N1845, N1534, N726, N852);
not NOT1 (N1848, N1799);
xor XOR2 (N1849, N1842, N998);
xor XOR2 (N1850, N1843, N1432);
buf BUF1 (N1851, N1828);
xor XOR2 (N1852, N1832, N1801);
nand NAND2 (N1853, N1846, N768);
nor NOR2 (N1854, N1836, N1369);
or OR2 (N1855, N1854, N1839);
or OR4 (N1856, N1852, N915, N289, N146);
nand NAND3 (N1857, N1847, N595, N1511);
or OR2 (N1858, N1851, N996);
not NOT1 (N1859, N1850);
nand NAND4 (N1860, N1837, N1858, N268, N826);
not NOT1 (N1861, N325);
buf BUF1 (N1862, N1849);
nand NAND2 (N1863, N1859, N357);
or OR4 (N1864, N1856, N964, N74, N802);
nand NAND2 (N1865, N1861, N1374);
nand NAND3 (N1866, N1860, N257, N1069);
xor XOR2 (N1867, N1857, N1095);
nor NOR4 (N1868, N1862, N1137, N1459, N45);
xor XOR2 (N1869, N1864, N1789);
nor NOR3 (N1870, N1867, N753, N1495);
nand NAND2 (N1871, N1869, N195);
and AND2 (N1872, N1870, N1567);
nand NAND4 (N1873, N1863, N637, N327, N1669);
nor NOR3 (N1874, N1873, N1007, N407);
or OR2 (N1875, N1874, N292);
not NOT1 (N1876, N1865);
or OR2 (N1877, N1872, N1230);
buf BUF1 (N1878, N1848);
or OR4 (N1879, N1871, N822, N1372, N1379);
nor NOR2 (N1880, N1875, N258);
nor NOR2 (N1881, N1868, N534);
or OR3 (N1882, N1881, N1334, N1594);
and AND3 (N1883, N1877, N1240, N567);
buf BUF1 (N1884, N1876);
nand NAND4 (N1885, N1878, N1023, N1840, N395);
and AND3 (N1886, N1885, N1030, N1454);
nand NAND4 (N1887, N1853, N441, N1162, N841);
buf BUF1 (N1888, N1880);
nand NAND4 (N1889, N1879, N1746, N1331, N1870);
or OR2 (N1890, N1884, N1517);
nor NOR4 (N1891, N1882, N1811, N1324, N419);
nor NOR2 (N1892, N1855, N1588);
xor XOR2 (N1893, N1888, N773);
nand NAND3 (N1894, N1841, N73, N1844);
nand NAND4 (N1895, N1892, N864, N999, N799);
xor XOR2 (N1896, N1891, N101);
and AND3 (N1897, N1886, N1356, N1880);
not NOT1 (N1898, N1893);
buf BUF1 (N1899, N1898);
nand NAND2 (N1900, N1895, N659);
nor NOR2 (N1901, N1887, N1545);
and AND3 (N1902, N1900, N1193, N1264);
nand NAND3 (N1903, N1866, N1578, N144);
xor XOR2 (N1904, N1889, N1777);
nor NOR3 (N1905, N1890, N84, N1609);
and AND2 (N1906, N1901, N1716);
xor XOR2 (N1907, N1905, N1146);
or OR4 (N1908, N1896, N512, N768, N890);
xor XOR2 (N1909, N1904, N311);
nor NOR2 (N1910, N1894, N1850);
or OR3 (N1911, N1907, N1779, N62);
nor NOR2 (N1912, N1897, N1326);
and AND2 (N1913, N1911, N519);
or OR4 (N1914, N1908, N1368, N140, N934);
not NOT1 (N1915, N1883);
xor XOR2 (N1916, N1914, N590);
buf BUF1 (N1917, N1910);
and AND2 (N1918, N1906, N1016);
buf BUF1 (N1919, N1903);
or OR3 (N1920, N1909, N481, N1196);
and AND3 (N1921, N1902, N87, N345);
not NOT1 (N1922, N1918);
not NOT1 (N1923, N1921);
or OR2 (N1924, N1915, N1915);
and AND2 (N1925, N1913, N438);
or OR3 (N1926, N1916, N110, N791);
or OR2 (N1927, N1924, N749);
and AND2 (N1928, N1927, N523);
and AND3 (N1929, N1917, N352, N164);
nor NOR2 (N1930, N1912, N1483);
not NOT1 (N1931, N1929);
not NOT1 (N1932, N1925);
nor NOR3 (N1933, N1932, N167, N1002);
not NOT1 (N1934, N1930);
buf BUF1 (N1935, N1926);
xor XOR2 (N1936, N1935, N1366);
nand NAND4 (N1937, N1933, N781, N2, N1838);
not NOT1 (N1938, N1934);
or OR4 (N1939, N1928, N1136, N135, N1574);
not NOT1 (N1940, N1919);
buf BUF1 (N1941, N1937);
not NOT1 (N1942, N1936);
not NOT1 (N1943, N1938);
nand NAND2 (N1944, N1931, N94);
nor NOR2 (N1945, N1942, N522);
nand NAND3 (N1946, N1939, N1916, N1362);
and AND3 (N1947, N1945, N1145, N1250);
nand NAND4 (N1948, N1923, N193, N1604, N1294);
xor XOR2 (N1949, N1946, N373);
buf BUF1 (N1950, N1922);
or OR3 (N1951, N1948, N125, N1624);
buf BUF1 (N1952, N1899);
nand NAND2 (N1953, N1949, N1199);
nand NAND3 (N1954, N1941, N907, N879);
and AND4 (N1955, N1953, N1239, N435, N937);
nand NAND3 (N1956, N1950, N1807, N1360);
or OR4 (N1957, N1952, N1277, N554, N832);
nand NAND2 (N1958, N1955, N320);
not NOT1 (N1959, N1920);
xor XOR2 (N1960, N1940, N1005);
not NOT1 (N1961, N1957);
and AND3 (N1962, N1951, N459, N1117);
and AND2 (N1963, N1944, N851);
nand NAND3 (N1964, N1960, N1165, N1139);
xor XOR2 (N1965, N1947, N897);
nor NOR3 (N1966, N1943, N578, N583);
buf BUF1 (N1967, N1958);
xor XOR2 (N1968, N1965, N1456);
nand NAND2 (N1969, N1963, N1361);
and AND3 (N1970, N1966, N992, N1470);
nand NAND3 (N1971, N1968, N180, N768);
xor XOR2 (N1972, N1967, N414);
and AND4 (N1973, N1961, N1825, N1874, N1428);
nand NAND4 (N1974, N1959, N1416, N1809, N1040);
or OR4 (N1975, N1956, N1566, N1941, N1654);
buf BUF1 (N1976, N1969);
nor NOR3 (N1977, N1975, N1308, N149);
buf BUF1 (N1978, N1977);
nor NOR2 (N1979, N1954, N1350);
and AND4 (N1980, N1971, N1568, N1870, N421);
buf BUF1 (N1981, N1980);
nand NAND2 (N1982, N1976, N720);
nand NAND4 (N1983, N1981, N1319, N1178, N1905);
or OR3 (N1984, N1973, N1586, N671);
buf BUF1 (N1985, N1970);
not NOT1 (N1986, N1978);
nor NOR3 (N1987, N1974, N1777, N954);
or OR3 (N1988, N1987, N1441, N1857);
or OR4 (N1989, N1979, N1171, N1777, N1875);
buf BUF1 (N1990, N1983);
nand NAND4 (N1991, N1988, N860, N1896, N843);
or OR2 (N1992, N1982, N1885);
xor XOR2 (N1993, N1991, N868);
or OR2 (N1994, N1964, N18);
and AND2 (N1995, N1985, N888);
and AND3 (N1996, N1972, N742, N161);
nor NOR3 (N1997, N1993, N1798, N629);
xor XOR2 (N1998, N1992, N839);
not NOT1 (N1999, N1994);
or OR2 (N2000, N1997, N1300);
nor NOR3 (N2001, N1989, N94, N810);
buf BUF1 (N2002, N1984);
nand NAND2 (N2003, N1998, N1896);
nand NAND4 (N2004, N1962, N273, N819, N1584);
nand NAND3 (N2005, N1990, N364, N118);
nor NOR3 (N2006, N2004, N1767, N12);
nand NAND3 (N2007, N2002, N715, N643);
xor XOR2 (N2008, N2001, N1370);
nor NOR3 (N2009, N2007, N272, N230);
or OR3 (N2010, N2006, N291, N1499);
nor NOR4 (N2011, N2008, N629, N96, N1016);
nand NAND2 (N2012, N2009, N1339);
nor NOR3 (N2013, N1999, N275, N1335);
xor XOR2 (N2014, N1986, N1855);
nand NAND4 (N2015, N2013, N1268, N208, N326);
endmodule