// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20;

output N410,N417,N418,N413,N414,N416,N395,N415,N419,N420;

nor NOR4 (N21, N20, N3, N20, N13);
or OR2 (N22, N8, N7);
and AND2 (N23, N22, N15);
xor XOR2 (N24, N13, N16);
or OR2 (N25, N18, N7);
xor XOR2 (N26, N11, N15);
and AND2 (N27, N1, N6);
not NOT1 (N28, N10);
and AND4 (N29, N10, N9, N23, N21);
and AND2 (N30, N15, N3);
xor XOR2 (N31, N25, N24);
buf BUF1 (N32, N30);
and AND4 (N33, N11, N13, N7, N14);
nor NOR3 (N34, N20, N15, N31);
nor NOR3 (N35, N6, N10, N28);
buf BUF1 (N36, N25);
nand NAND3 (N37, N12, N30, N19);
xor XOR2 (N38, N20, N8);
xor XOR2 (N39, N38, N32);
or OR3 (N40, N3, N13, N4);
and AND4 (N41, N27, N34, N31, N37);
and AND3 (N42, N12, N13, N41);
not NOT1 (N43, N27);
nand NAND4 (N44, N24, N12, N14, N3);
and AND3 (N45, N42, N17, N11);
or OR3 (N46, N26, N6, N30);
xor XOR2 (N47, N29, N33);
or OR2 (N48, N20, N30);
and AND2 (N49, N36, N33);
and AND3 (N50, N35, N14, N6);
xor XOR2 (N51, N49, N17);
xor XOR2 (N52, N51, N15);
not NOT1 (N53, N47);
or OR4 (N54, N52, N16, N50, N17);
buf BUF1 (N55, N37);
not NOT1 (N56, N53);
or OR4 (N57, N44, N38, N21, N36);
nor NOR2 (N58, N45, N38);
or OR4 (N59, N40, N51, N27, N19);
or OR2 (N60, N56, N27);
and AND3 (N61, N58, N29, N22);
nor NOR2 (N62, N48, N53);
nand NAND4 (N63, N59, N4, N11, N25);
buf BUF1 (N64, N54);
buf BUF1 (N65, N55);
nand NAND4 (N66, N39, N7, N55, N36);
not NOT1 (N67, N66);
nand NAND2 (N68, N60, N59);
buf BUF1 (N69, N64);
nand NAND2 (N70, N68, N68);
nand NAND3 (N71, N57, N34, N29);
or OR3 (N72, N63, N58, N32);
not NOT1 (N73, N46);
xor XOR2 (N74, N71, N48);
and AND2 (N75, N70, N5);
xor XOR2 (N76, N69, N10);
or OR3 (N77, N75, N58, N76);
or OR2 (N78, N49, N27);
nand NAND4 (N79, N65, N76, N29, N67);
not NOT1 (N80, N8);
or OR3 (N81, N61, N53, N25);
nor NOR3 (N82, N77, N72, N3);
nor NOR4 (N83, N48, N5, N66, N2);
not NOT1 (N84, N62);
or OR3 (N85, N80, N50, N8);
xor XOR2 (N86, N78, N20);
nand NAND3 (N87, N86, N26, N29);
nor NOR4 (N88, N79, N31, N28, N47);
and AND2 (N89, N87, N37);
and AND2 (N90, N89, N82);
buf BUF1 (N91, N87);
or OR3 (N92, N43, N14, N55);
and AND4 (N93, N81, N38, N16, N45);
and AND3 (N94, N73, N36, N90);
xor XOR2 (N95, N59, N87);
xor XOR2 (N96, N88, N41);
and AND4 (N97, N91, N93, N36, N39);
nand NAND3 (N98, N52, N71, N68);
not NOT1 (N99, N97);
or OR2 (N100, N96, N62);
nor NOR3 (N101, N83, N64, N27);
nor NOR2 (N102, N98, N18);
xor XOR2 (N103, N94, N65);
buf BUF1 (N104, N102);
buf BUF1 (N105, N74);
or OR4 (N106, N105, N90, N38, N45);
buf BUF1 (N107, N106);
xor XOR2 (N108, N107, N101);
not NOT1 (N109, N87);
xor XOR2 (N110, N100, N60);
xor XOR2 (N111, N110, N92);
buf BUF1 (N112, N78);
buf BUF1 (N113, N95);
xor XOR2 (N114, N103, N25);
buf BUF1 (N115, N114);
xor XOR2 (N116, N115, N50);
buf BUF1 (N117, N116);
nor NOR4 (N118, N84, N39, N85, N31);
nor NOR4 (N119, N70, N10, N107, N90);
nand NAND4 (N120, N109, N42, N61, N66);
nor NOR4 (N121, N119, N56, N51, N70);
nand NAND3 (N122, N108, N32, N48);
buf BUF1 (N123, N120);
not NOT1 (N124, N121);
and AND3 (N125, N124, N35, N37);
or OR3 (N126, N99, N75, N47);
or OR3 (N127, N125, N108, N96);
nand NAND3 (N128, N127, N38, N88);
or OR4 (N129, N117, N100, N113, N81);
xor XOR2 (N130, N54, N88);
and AND4 (N131, N126, N99, N96, N120);
buf BUF1 (N132, N111);
or OR2 (N133, N118, N63);
nand NAND2 (N134, N132, N129);
nor NOR3 (N135, N32, N45, N27);
not NOT1 (N136, N133);
buf BUF1 (N137, N135);
not NOT1 (N138, N112);
or OR4 (N139, N130, N94, N6, N131);
xor XOR2 (N140, N89, N37);
buf BUF1 (N141, N134);
nand NAND3 (N142, N104, N108, N136);
nor NOR2 (N143, N55, N111);
and AND2 (N144, N122, N122);
nor NOR3 (N145, N123, N17, N111);
nand NAND4 (N146, N140, N95, N5, N122);
not NOT1 (N147, N144);
xor XOR2 (N148, N147, N15);
or OR2 (N149, N146, N78);
nand NAND4 (N150, N142, N54, N46, N135);
buf BUF1 (N151, N139);
or OR2 (N152, N141, N133);
nand NAND2 (N153, N150, N41);
and AND2 (N154, N148, N106);
buf BUF1 (N155, N151);
buf BUF1 (N156, N138);
xor XOR2 (N157, N156, N140);
and AND2 (N158, N143, N22);
or OR4 (N159, N155, N3, N56, N2);
buf BUF1 (N160, N128);
not NOT1 (N161, N152);
xor XOR2 (N162, N161, N64);
xor XOR2 (N163, N159, N36);
nand NAND4 (N164, N157, N17, N74, N98);
not NOT1 (N165, N154);
not NOT1 (N166, N145);
nand NAND2 (N167, N162, N36);
or OR3 (N168, N137, N84, N140);
nor NOR3 (N169, N164, N56, N94);
buf BUF1 (N170, N169);
nor NOR4 (N171, N163, N141, N108, N85);
buf BUF1 (N172, N165);
xor XOR2 (N173, N168, N142);
and AND4 (N174, N173, N146, N93, N156);
and AND3 (N175, N167, N30, N55);
nand NAND2 (N176, N171, N116);
nor NOR3 (N177, N176, N21, N139);
nand NAND4 (N178, N172, N163, N39, N36);
and AND2 (N179, N177, N149);
or OR3 (N180, N159, N119, N140);
nand NAND2 (N181, N175, N60);
or OR4 (N182, N181, N151, N29, N94);
and AND3 (N183, N166, N53, N144);
or OR4 (N184, N182, N120, N56, N89);
buf BUF1 (N185, N180);
or OR2 (N186, N160, N10);
nor NOR2 (N187, N158, N107);
xor XOR2 (N188, N183, N154);
and AND3 (N189, N153, N65, N183);
xor XOR2 (N190, N185, N77);
xor XOR2 (N191, N187, N132);
nor NOR3 (N192, N174, N120, N177);
xor XOR2 (N193, N184, N187);
not NOT1 (N194, N179);
not NOT1 (N195, N170);
xor XOR2 (N196, N194, N39);
xor XOR2 (N197, N186, N2);
xor XOR2 (N198, N197, N173);
xor XOR2 (N199, N188, N35);
nand NAND4 (N200, N196, N100, N163, N99);
nand NAND4 (N201, N195, N16, N116, N42);
nor NOR3 (N202, N190, N3, N195);
xor XOR2 (N203, N200, N171);
nor NOR4 (N204, N203, N61, N101, N123);
not NOT1 (N205, N202);
nand NAND2 (N206, N192, N118);
xor XOR2 (N207, N193, N79);
not NOT1 (N208, N205);
not NOT1 (N209, N206);
nor NOR2 (N210, N191, N137);
nand NAND2 (N211, N189, N3);
xor XOR2 (N212, N209, N129);
or OR4 (N213, N208, N148, N14, N94);
not NOT1 (N214, N210);
or OR4 (N215, N212, N116, N106, N48);
or OR2 (N216, N215, N76);
nand NAND2 (N217, N213, N124);
nor NOR4 (N218, N211, N215, N59, N177);
buf BUF1 (N219, N216);
nor NOR2 (N220, N207, N108);
and AND4 (N221, N219, N11, N155, N102);
buf BUF1 (N222, N220);
xor XOR2 (N223, N222, N205);
not NOT1 (N224, N221);
not NOT1 (N225, N224);
or OR4 (N226, N214, N217, N159, N66);
xor XOR2 (N227, N24, N28);
or OR2 (N228, N198, N143);
or OR2 (N229, N178, N194);
and AND2 (N230, N226, N56);
and AND4 (N231, N218, N9, N142, N105);
nor NOR2 (N232, N230, N159);
not NOT1 (N233, N227);
nand NAND4 (N234, N228, N45, N183, N74);
and AND4 (N235, N225, N86, N6, N44);
nand NAND3 (N236, N223, N201, N105);
not NOT1 (N237, N235);
not NOT1 (N238, N176);
not NOT1 (N239, N238);
nand NAND3 (N240, N204, N119, N154);
or OR3 (N241, N240, N114, N211);
and AND3 (N242, N233, N135, N132);
and AND2 (N243, N232, N231);
buf BUF1 (N244, N60);
or OR2 (N245, N229, N201);
not NOT1 (N246, N241);
buf BUF1 (N247, N245);
not NOT1 (N248, N237);
buf BUF1 (N249, N248);
and AND3 (N250, N247, N201, N105);
buf BUF1 (N251, N239);
or OR2 (N252, N199, N83);
nand NAND4 (N253, N242, N66, N215, N228);
and AND4 (N254, N250, N115, N133, N105);
and AND4 (N255, N236, N46, N154, N120);
nand NAND2 (N256, N251, N46);
or OR2 (N257, N234, N9);
and AND3 (N258, N253, N76, N177);
nor NOR4 (N259, N244, N150, N92, N184);
not NOT1 (N260, N259);
xor XOR2 (N261, N257, N7);
and AND2 (N262, N255, N143);
and AND2 (N263, N252, N65);
not NOT1 (N264, N246);
nor NOR3 (N265, N260, N13, N220);
nor NOR3 (N266, N261, N183, N217);
nor NOR3 (N267, N263, N247, N94);
buf BUF1 (N268, N254);
and AND2 (N269, N268, N185);
or OR4 (N270, N266, N110, N63, N213);
xor XOR2 (N271, N269, N17);
nand NAND3 (N272, N262, N181, N265);
nand NAND2 (N273, N4, N238);
buf BUF1 (N274, N264);
xor XOR2 (N275, N272, N65);
xor XOR2 (N276, N258, N268);
nor NOR4 (N277, N267, N163, N172, N64);
and AND4 (N278, N274, N260, N211, N204);
nor NOR2 (N279, N243, N222);
or OR4 (N280, N273, N113, N237, N211);
xor XOR2 (N281, N249, N93);
and AND3 (N282, N277, N44, N27);
and AND2 (N283, N282, N236);
xor XOR2 (N284, N279, N14);
xor XOR2 (N285, N283, N13);
and AND2 (N286, N276, N257);
nor NOR3 (N287, N270, N186, N248);
nand NAND2 (N288, N281, N200);
not NOT1 (N289, N256);
nand NAND4 (N290, N280, N234, N192, N178);
and AND3 (N291, N288, N239, N171);
buf BUF1 (N292, N285);
or OR3 (N293, N278, N18, N76);
nand NAND3 (N294, N271, N182, N55);
nor NOR4 (N295, N293, N291, N249, N224);
or OR2 (N296, N150, N281);
or OR2 (N297, N289, N185);
buf BUF1 (N298, N292);
or OR4 (N299, N295, N146, N273, N149);
buf BUF1 (N300, N284);
nor NOR2 (N301, N296, N24);
nor NOR2 (N302, N301, N262);
buf BUF1 (N303, N298);
not NOT1 (N304, N303);
and AND3 (N305, N290, N243, N201);
nand NAND2 (N306, N294, N304);
xor XOR2 (N307, N150, N79);
xor XOR2 (N308, N287, N118);
or OR2 (N309, N275, N136);
nand NAND3 (N310, N299, N162, N224);
nor NOR4 (N311, N300, N299, N53, N304);
buf BUF1 (N312, N310);
nand NAND4 (N313, N286, N108, N67, N214);
nand NAND3 (N314, N306, N99, N230);
or OR2 (N315, N305, N21);
or OR2 (N316, N313, N290);
xor XOR2 (N317, N308, N176);
or OR3 (N318, N309, N87, N133);
nand NAND4 (N319, N312, N240, N23, N267);
buf BUF1 (N320, N297);
nand NAND3 (N321, N315, N102, N236);
xor XOR2 (N322, N307, N128);
not NOT1 (N323, N321);
nor NOR2 (N324, N317, N221);
buf BUF1 (N325, N316);
not NOT1 (N326, N325);
or OR3 (N327, N320, N241, N174);
or OR3 (N328, N318, N129, N175);
xor XOR2 (N329, N322, N69);
nand NAND2 (N330, N319, N9);
and AND2 (N331, N323, N325);
or OR2 (N332, N324, N183);
buf BUF1 (N333, N329);
xor XOR2 (N334, N314, N36);
nor NOR3 (N335, N328, N17, N14);
and AND2 (N336, N330, N16);
nand NAND3 (N337, N332, N208, N55);
or OR3 (N338, N335, N273, N29);
nor NOR2 (N339, N311, N140);
buf BUF1 (N340, N339);
not NOT1 (N341, N338);
and AND4 (N342, N340, N160, N316, N182);
or OR3 (N343, N302, N333, N132);
or OR3 (N344, N240, N25, N132);
and AND3 (N345, N336, N249, N341);
and AND4 (N346, N83, N241, N51, N275);
xor XOR2 (N347, N342, N318);
nor NOR4 (N348, N345, N13, N35, N108);
not NOT1 (N349, N326);
or OR4 (N350, N347, N111, N121, N41);
and AND4 (N351, N344, N86, N332, N179);
nor NOR4 (N352, N346, N249, N125, N284);
and AND4 (N353, N349, N88, N276, N338);
buf BUF1 (N354, N350);
buf BUF1 (N355, N352);
nand NAND2 (N356, N337, N232);
nand NAND4 (N357, N351, N39, N119, N27);
nor NOR2 (N358, N334, N218);
nor NOR4 (N359, N348, N70, N62, N47);
nand NAND4 (N360, N354, N16, N202, N10);
or OR3 (N361, N357, N303, N22);
nor NOR3 (N362, N353, N335, N232);
xor XOR2 (N363, N355, N270);
not NOT1 (N364, N358);
or OR2 (N365, N360, N83);
and AND2 (N366, N359, N246);
xor XOR2 (N367, N365, N68);
nor NOR3 (N368, N343, N17, N61);
buf BUF1 (N369, N363);
not NOT1 (N370, N361);
or OR4 (N371, N356, N216, N169, N50);
nand NAND2 (N372, N368, N184);
or OR3 (N373, N331, N364, N179);
buf BUF1 (N374, N149);
buf BUF1 (N375, N370);
buf BUF1 (N376, N372);
not NOT1 (N377, N375);
or OR4 (N378, N376, N341, N345, N96);
buf BUF1 (N379, N362);
and AND3 (N380, N379, N250, N121);
nor NOR2 (N381, N367, N316);
buf BUF1 (N382, N369);
buf BUF1 (N383, N378);
or OR2 (N384, N383, N142);
or OR3 (N385, N371, N185, N130);
buf BUF1 (N386, N382);
buf BUF1 (N387, N327);
nor NOR2 (N388, N381, N351);
buf BUF1 (N389, N373);
or OR3 (N390, N380, N249, N354);
nor NOR3 (N391, N386, N32, N142);
or OR2 (N392, N374, N7);
xor XOR2 (N393, N384, N344);
xor XOR2 (N394, N377, N145);
nand NAND2 (N395, N389, N300);
nor NOR2 (N396, N387, N336);
xor XOR2 (N397, N390, N91);
nand NAND3 (N398, N366, N282, N371);
buf BUF1 (N399, N394);
xor XOR2 (N400, N399, N86);
nand NAND3 (N401, N393, N267, N260);
nand NAND4 (N402, N400, N97, N365, N329);
or OR3 (N403, N396, N142, N252);
and AND2 (N404, N402, N328);
not NOT1 (N405, N401);
xor XOR2 (N406, N385, N262);
buf BUF1 (N407, N392);
nor NOR4 (N408, N405, N152, N243, N125);
not NOT1 (N409, N407);
not NOT1 (N410, N398);
nand NAND2 (N411, N397, N95);
nor NOR2 (N412, N403, N362);
and AND2 (N413, N406, N41);
nand NAND2 (N414, N408, N222);
or OR4 (N415, N404, N13, N40, N88);
buf BUF1 (N416, N411);
nor NOR3 (N417, N412, N305, N116);
buf BUF1 (N418, N391);
buf BUF1 (N419, N388);
or OR3 (N420, N409, N283, N356);
endmodule