// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13;

output N390,N398,N409,N407,N410,N402,N404,N412,N396,N413;

nand NAND4 (N14, N3, N10, N8, N8);
or OR2 (N15, N3, N2);
nand NAND4 (N16, N6, N11, N13, N8);
or OR3 (N17, N16, N5, N8);
not NOT1 (N18, N12);
xor XOR2 (N19, N4, N18);
xor XOR2 (N20, N16, N7);
nand NAND2 (N21, N4, N3);
buf BUF1 (N22, N18);
not NOT1 (N23, N1);
buf BUF1 (N24, N10);
buf BUF1 (N25, N12);
or OR4 (N26, N15, N7, N20, N2);
or OR4 (N27, N20, N14, N15, N15);
or OR4 (N28, N7, N13, N23, N17);
nor NOR2 (N29, N12, N3);
xor XOR2 (N30, N24, N26);
nor NOR4 (N31, N27, N17, N20, N2);
buf BUF1 (N32, N16);
not NOT1 (N33, N5);
and AND2 (N34, N30, N27);
xor XOR2 (N35, N31, N21);
or OR2 (N36, N3, N31);
or OR4 (N37, N33, N20, N12, N25);
buf BUF1 (N38, N25);
and AND3 (N39, N28, N10, N15);
nand NAND2 (N40, N37, N29);
not NOT1 (N41, N16);
xor XOR2 (N42, N19, N12);
not NOT1 (N43, N32);
nand NAND3 (N44, N42, N26, N17);
nor NOR4 (N45, N39, N39, N11, N31);
not NOT1 (N46, N38);
and AND2 (N47, N40, N7);
buf BUF1 (N48, N43);
not NOT1 (N49, N35);
or OR2 (N50, N46, N13);
nand NAND3 (N51, N49, N39, N25);
nor NOR4 (N52, N45, N1, N11, N48);
nor NOR3 (N53, N38, N10, N41);
nor NOR3 (N54, N26, N38, N26);
and AND2 (N55, N51, N16);
xor XOR2 (N56, N55, N37);
nand NAND4 (N57, N22, N43, N28, N55);
or OR3 (N58, N53, N28, N23);
buf BUF1 (N59, N56);
or OR3 (N60, N47, N41, N37);
xor XOR2 (N61, N57, N40);
nor NOR3 (N62, N44, N56, N10);
not NOT1 (N63, N58);
and AND3 (N64, N60, N3, N28);
or OR4 (N65, N61, N60, N36, N59);
buf BUF1 (N66, N56);
or OR2 (N67, N20, N47);
nor NOR2 (N68, N66, N57);
and AND3 (N69, N63, N31, N17);
and AND3 (N70, N52, N41, N56);
or OR3 (N71, N64, N51, N29);
or OR2 (N72, N69, N68);
xor XOR2 (N73, N63, N27);
nand NAND4 (N74, N70, N35, N71, N52);
xor XOR2 (N75, N13, N38);
nand NAND2 (N76, N73, N51);
nand NAND2 (N77, N65, N53);
xor XOR2 (N78, N62, N49);
or OR3 (N79, N54, N1, N25);
or OR2 (N80, N67, N55);
nor NOR4 (N81, N34, N18, N77, N23);
nor NOR3 (N82, N4, N30, N24);
xor XOR2 (N83, N80, N59);
nand NAND3 (N84, N82, N83, N17);
nand NAND3 (N85, N12, N6, N78);
buf BUF1 (N86, N64);
xor XOR2 (N87, N50, N60);
and AND2 (N88, N86, N65);
nand NAND4 (N89, N74, N51, N26, N88);
nor NOR3 (N90, N56, N4, N18);
nand NAND3 (N91, N84, N72, N58);
and AND2 (N92, N5, N26);
nand NAND3 (N93, N87, N46, N68);
not NOT1 (N94, N91);
and AND3 (N95, N85, N66, N7);
or OR2 (N96, N76, N19);
and AND2 (N97, N95, N48);
and AND4 (N98, N94, N55, N65, N76);
buf BUF1 (N99, N79);
nand NAND4 (N100, N81, N53, N97, N47);
and AND2 (N101, N21, N87);
or OR2 (N102, N98, N94);
and AND2 (N103, N93, N51);
or OR2 (N104, N102, N32);
nand NAND4 (N105, N99, N80, N68, N36);
and AND2 (N106, N101, N4);
not NOT1 (N107, N92);
buf BUF1 (N108, N106);
or OR2 (N109, N107, N99);
buf BUF1 (N110, N90);
not NOT1 (N111, N96);
buf BUF1 (N112, N89);
nand NAND4 (N113, N112, N84, N76, N67);
or OR3 (N114, N104, N67, N89);
xor XOR2 (N115, N100, N66);
and AND3 (N116, N109, N63, N77);
xor XOR2 (N117, N116, N63);
not NOT1 (N118, N103);
nor NOR4 (N119, N118, N57, N113, N42);
xor XOR2 (N120, N63, N41);
nor NOR3 (N121, N110, N59, N9);
not NOT1 (N122, N115);
nor NOR2 (N123, N114, N6);
and AND2 (N124, N108, N51);
and AND3 (N125, N120, N84, N34);
not NOT1 (N126, N105);
nor NOR2 (N127, N75, N108);
or OR2 (N128, N124, N45);
not NOT1 (N129, N111);
not NOT1 (N130, N121);
not NOT1 (N131, N125);
nor NOR2 (N132, N123, N107);
nor NOR4 (N133, N128, N75, N73, N106);
nor NOR4 (N134, N132, N36, N43, N14);
buf BUF1 (N135, N129);
nor NOR3 (N136, N131, N107, N105);
nor NOR3 (N137, N117, N2, N82);
not NOT1 (N138, N137);
not NOT1 (N139, N126);
not NOT1 (N140, N133);
and AND2 (N141, N136, N64);
nand NAND2 (N142, N140, N20);
buf BUF1 (N143, N127);
xor XOR2 (N144, N142, N104);
or OR4 (N145, N143, N114, N37, N144);
nor NOR3 (N146, N84, N9, N98);
or OR2 (N147, N146, N22);
xor XOR2 (N148, N147, N134);
nand NAND4 (N149, N104, N59, N23, N45);
xor XOR2 (N150, N139, N55);
buf BUF1 (N151, N130);
nor NOR3 (N152, N135, N62, N83);
buf BUF1 (N153, N150);
not NOT1 (N154, N145);
xor XOR2 (N155, N119, N114);
buf BUF1 (N156, N151);
not NOT1 (N157, N138);
xor XOR2 (N158, N148, N131);
not NOT1 (N159, N154);
xor XOR2 (N160, N155, N90);
not NOT1 (N161, N141);
or OR2 (N162, N158, N98);
not NOT1 (N163, N149);
nand NAND3 (N164, N153, N48, N124);
buf BUF1 (N165, N157);
buf BUF1 (N166, N160);
nor NOR3 (N167, N165, N157, N163);
nand NAND4 (N168, N152, N98, N54, N103);
or OR3 (N169, N109, N62, N26);
or OR3 (N170, N169, N164, N108);
not NOT1 (N171, N39);
buf BUF1 (N172, N159);
buf BUF1 (N173, N170);
nor NOR4 (N174, N173, N24, N158, N128);
and AND2 (N175, N172, N4);
nor NOR3 (N176, N175, N120, N148);
nand NAND3 (N177, N166, N61, N104);
not NOT1 (N178, N174);
not NOT1 (N179, N171);
not NOT1 (N180, N179);
nor NOR3 (N181, N180, N89, N39);
or OR2 (N182, N178, N161);
nor NOR2 (N183, N122, N79);
and AND3 (N184, N47, N158, N37);
not NOT1 (N185, N162);
buf BUF1 (N186, N168);
not NOT1 (N187, N181);
xor XOR2 (N188, N182, N114);
xor XOR2 (N189, N186, N78);
buf BUF1 (N190, N185);
or OR3 (N191, N183, N32, N180);
xor XOR2 (N192, N167, N89);
not NOT1 (N193, N176);
xor XOR2 (N194, N192, N20);
and AND3 (N195, N156, N43, N18);
nor NOR3 (N196, N190, N163, N187);
not NOT1 (N197, N163);
not NOT1 (N198, N184);
not NOT1 (N199, N194);
nand NAND2 (N200, N198, N65);
nand NAND4 (N201, N188, N74, N15, N63);
buf BUF1 (N202, N197);
buf BUF1 (N203, N191);
nor NOR3 (N204, N203, N73, N132);
nand NAND3 (N205, N177, N38, N121);
or OR2 (N206, N195, N165);
nor NOR4 (N207, N200, N24, N169, N167);
and AND4 (N208, N196, N18, N41, N206);
and AND4 (N209, N58, N137, N125, N99);
or OR4 (N210, N193, N30, N151, N198);
or OR2 (N211, N201, N18);
buf BUF1 (N212, N207);
or OR3 (N213, N212, N24, N128);
nand NAND3 (N214, N205, N152, N167);
nand NAND3 (N215, N208, N158, N85);
and AND2 (N216, N189, N77);
nand NAND3 (N217, N213, N85, N209);
nor NOR2 (N218, N3, N82);
and AND4 (N219, N217, N6, N164, N56);
nor NOR2 (N220, N215, N154);
not NOT1 (N221, N214);
or OR3 (N222, N220, N125, N172);
buf BUF1 (N223, N218);
nand NAND3 (N224, N223, N110, N94);
nor NOR3 (N225, N221, N82, N6);
not NOT1 (N226, N202);
or OR2 (N227, N224, N219);
nor NOR2 (N228, N37, N33);
buf BUF1 (N229, N228);
not NOT1 (N230, N216);
or OR4 (N231, N199, N135, N64, N12);
nand NAND3 (N232, N210, N101, N156);
nor NOR4 (N233, N232, N152, N112, N131);
nand NAND4 (N234, N229, N34, N161, N40);
and AND2 (N235, N231, N115);
not NOT1 (N236, N234);
nand NAND2 (N237, N226, N28);
or OR4 (N238, N222, N235, N214, N97);
or OR3 (N239, N171, N169, N8);
nor NOR4 (N240, N230, N204, N13, N91);
xor XOR2 (N241, N39, N188);
nor NOR2 (N242, N237, N66);
or OR2 (N243, N233, N31);
or OR4 (N244, N225, N31, N52, N140);
buf BUF1 (N245, N211);
nand NAND2 (N246, N227, N136);
not NOT1 (N247, N238);
xor XOR2 (N248, N239, N26);
nand NAND3 (N249, N247, N167, N178);
and AND4 (N250, N242, N7, N210, N5);
nand NAND2 (N251, N241, N54);
not NOT1 (N252, N246);
nor NOR3 (N253, N245, N171, N200);
buf BUF1 (N254, N252);
and AND4 (N255, N248, N47, N203, N131);
and AND3 (N256, N255, N66, N236);
xor XOR2 (N257, N76, N248);
or OR4 (N258, N243, N14, N60, N209);
nor NOR2 (N259, N250, N52);
nand NAND2 (N260, N254, N21);
buf BUF1 (N261, N249);
nand NAND3 (N262, N256, N146, N80);
and AND4 (N263, N257, N201, N129, N193);
or OR2 (N264, N251, N191);
not NOT1 (N265, N261);
nand NAND3 (N266, N253, N52, N131);
nand NAND4 (N267, N263, N144, N250, N154);
nor NOR4 (N268, N264, N198, N122, N237);
nand NAND4 (N269, N260, N53, N39, N5);
or OR2 (N270, N244, N147);
xor XOR2 (N271, N258, N200);
or OR2 (N272, N259, N146);
nand NAND4 (N273, N240, N130, N38, N17);
and AND2 (N274, N273, N26);
and AND2 (N275, N274, N115);
not NOT1 (N276, N267);
not NOT1 (N277, N270);
xor XOR2 (N278, N276, N66);
xor XOR2 (N279, N265, N92);
nor NOR3 (N280, N279, N172, N64);
nor NOR3 (N281, N271, N169, N82);
buf BUF1 (N282, N262);
nand NAND4 (N283, N266, N203, N117, N272);
xor XOR2 (N284, N160, N56);
or OR3 (N285, N280, N107, N82);
or OR2 (N286, N282, N18);
and AND3 (N287, N275, N12, N151);
xor XOR2 (N288, N268, N259);
nor NOR4 (N289, N286, N28, N158, N27);
buf BUF1 (N290, N269);
nor NOR3 (N291, N287, N46, N157);
not NOT1 (N292, N284);
and AND3 (N293, N288, N34, N41);
buf BUF1 (N294, N277);
nor NOR2 (N295, N285, N66);
nor NOR3 (N296, N295, N241, N288);
nand NAND3 (N297, N278, N196, N226);
not NOT1 (N298, N293);
xor XOR2 (N299, N281, N40);
buf BUF1 (N300, N290);
xor XOR2 (N301, N300, N145);
buf BUF1 (N302, N294);
nand NAND3 (N303, N292, N235, N197);
not NOT1 (N304, N302);
nor NOR3 (N305, N297, N75, N59);
nand NAND3 (N306, N291, N7, N251);
xor XOR2 (N307, N301, N111);
or OR4 (N308, N306, N64, N273, N51);
buf BUF1 (N309, N305);
not NOT1 (N310, N283);
nor NOR3 (N311, N303, N145, N112);
or OR3 (N312, N310, N192, N84);
not NOT1 (N313, N289);
buf BUF1 (N314, N298);
xor XOR2 (N315, N308, N239);
nand NAND4 (N316, N315, N82, N168, N38);
buf BUF1 (N317, N314);
not NOT1 (N318, N313);
xor XOR2 (N319, N304, N89);
nand NAND2 (N320, N296, N188);
xor XOR2 (N321, N319, N169);
not NOT1 (N322, N312);
and AND2 (N323, N299, N118);
nand NAND3 (N324, N309, N160, N43);
not NOT1 (N325, N320);
nand NAND3 (N326, N307, N168, N162);
xor XOR2 (N327, N325, N324);
nand NAND4 (N328, N234, N213, N145, N232);
nor NOR3 (N329, N323, N186, N137);
and AND4 (N330, N321, N107, N224, N78);
not NOT1 (N331, N326);
nor NOR2 (N332, N322, N118);
and AND3 (N333, N317, N167, N305);
or OR4 (N334, N333, N112, N275, N260);
and AND4 (N335, N316, N38, N75, N30);
xor XOR2 (N336, N328, N299);
nand NAND3 (N337, N336, N189, N255);
xor XOR2 (N338, N334, N14);
not NOT1 (N339, N337);
or OR3 (N340, N338, N200, N318);
nand NAND4 (N341, N248, N252, N175, N271);
buf BUF1 (N342, N332);
nor NOR2 (N343, N340, N165);
xor XOR2 (N344, N329, N256);
not NOT1 (N345, N335);
and AND4 (N346, N341, N73, N156, N6);
buf BUF1 (N347, N346);
nand NAND3 (N348, N347, N85, N194);
nor NOR4 (N349, N339, N184, N336, N289);
nand NAND3 (N350, N331, N333, N290);
nor NOR2 (N351, N343, N49);
buf BUF1 (N352, N348);
buf BUF1 (N353, N327);
or OR2 (N354, N311, N337);
nor NOR4 (N355, N354, N167, N218, N292);
or OR4 (N356, N342, N155, N318, N229);
buf BUF1 (N357, N350);
nand NAND2 (N358, N351, N312);
and AND4 (N359, N330, N252, N38, N186);
or OR4 (N360, N349, N245, N182, N284);
buf BUF1 (N361, N353);
and AND3 (N362, N359, N153, N283);
nand NAND2 (N363, N345, N145);
nand NAND4 (N364, N362, N98, N124, N171);
xor XOR2 (N365, N364, N209);
buf BUF1 (N366, N365);
xor XOR2 (N367, N356, N17);
nand NAND3 (N368, N344, N230, N236);
xor XOR2 (N369, N368, N362);
not NOT1 (N370, N369);
xor XOR2 (N371, N357, N9);
and AND2 (N372, N358, N119);
not NOT1 (N373, N363);
buf BUF1 (N374, N360);
nor NOR3 (N375, N373, N324, N272);
and AND2 (N376, N352, N100);
and AND3 (N377, N372, N365, N172);
or OR3 (N378, N370, N104, N21);
xor XOR2 (N379, N376, N166);
and AND3 (N380, N377, N110, N160);
not NOT1 (N381, N375);
and AND4 (N382, N380, N206, N227, N376);
buf BUF1 (N383, N374);
nand NAND4 (N384, N361, N326, N41, N341);
buf BUF1 (N385, N382);
nand NAND4 (N386, N381, N322, N124, N182);
nand NAND2 (N387, N366, N86);
nand NAND3 (N388, N383, N63, N283);
not NOT1 (N389, N387);
or OR4 (N390, N385, N319, N339, N175);
buf BUF1 (N391, N378);
xor XOR2 (N392, N371, N28);
not NOT1 (N393, N384);
xor XOR2 (N394, N392, N220);
nand NAND3 (N395, N389, N98, N175);
buf BUF1 (N396, N379);
buf BUF1 (N397, N394);
xor XOR2 (N398, N397, N58);
and AND2 (N399, N355, N244);
xor XOR2 (N400, N393, N248);
not NOT1 (N401, N367);
xor XOR2 (N402, N400, N244);
nor NOR2 (N403, N401, N133);
xor XOR2 (N404, N386, N319);
or OR3 (N405, N388, N40, N170);
and AND3 (N406, N405, N240, N248);
nor NOR2 (N407, N406, N312);
and AND3 (N408, N403, N178, N155);
buf BUF1 (N409, N395);
and AND2 (N410, N408, N345);
not NOT1 (N411, N399);
or OR3 (N412, N391, N306, N150);
not NOT1 (N413, N411);
endmodule