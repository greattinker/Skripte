// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11;

output N4008,N4002,N4010,N4006,N4007,N4005,N3985,N4009,N4001,N4011;

nor NOR3 (N12, N10, N8, N3);
buf BUF1 (N13, N11);
and AND2 (N14, N13, N6);
and AND3 (N15, N1, N14, N5);
not NOT1 (N16, N12);
not NOT1 (N17, N11);
nand NAND4 (N18, N6, N10, N16, N4);
or OR3 (N19, N13, N4, N10);
nand NAND2 (N20, N18, N3);
nor NOR2 (N21, N17, N1);
and AND2 (N22, N16, N8);
nor NOR4 (N23, N1, N8, N12, N8);
nand NAND4 (N24, N10, N23, N9, N18);
not NOT1 (N25, N13);
nor NOR2 (N26, N15, N19);
xor XOR2 (N27, N1, N1);
or OR2 (N28, N26, N19);
not NOT1 (N29, N2);
or OR4 (N30, N12, N25, N29, N3);
buf BUF1 (N31, N24);
xor XOR2 (N32, N1, N16);
xor XOR2 (N33, N20, N5);
nor NOR2 (N34, N4, N20);
buf BUF1 (N35, N13);
or OR2 (N36, N28, N3);
nor NOR2 (N37, N21, N34);
nor NOR2 (N38, N27, N22);
nand NAND3 (N39, N28, N26, N13);
nor NOR2 (N40, N28, N23);
and AND4 (N41, N40, N31, N5, N22);
xor XOR2 (N42, N4, N34);
buf BUF1 (N43, N38);
and AND4 (N44, N41, N18, N41, N24);
not NOT1 (N45, N32);
and AND3 (N46, N39, N37, N14);
or OR2 (N47, N32, N11);
not NOT1 (N48, N47);
nand NAND4 (N49, N48, N30, N35, N33);
buf BUF1 (N50, N32);
and AND2 (N51, N2, N2);
nand NAND4 (N52, N12, N16, N25, N36);
not NOT1 (N53, N47);
nor NOR2 (N54, N50, N1);
xor XOR2 (N55, N43, N17);
and AND2 (N56, N44, N19);
or OR2 (N57, N45, N46);
xor XOR2 (N58, N16, N42);
not NOT1 (N59, N26);
or OR3 (N60, N59, N59, N44);
not NOT1 (N61, N57);
or OR2 (N62, N61, N21);
buf BUF1 (N63, N58);
nand NAND2 (N64, N62, N36);
nand NAND4 (N65, N56, N24, N33, N46);
and AND4 (N66, N51, N34, N62, N48);
not NOT1 (N67, N49);
nand NAND3 (N68, N67, N53, N46);
xor XOR2 (N69, N25, N55);
nand NAND4 (N70, N31, N25, N26, N19);
and AND3 (N71, N65, N58, N31);
xor XOR2 (N72, N66, N38);
nand NAND4 (N73, N71, N15, N41, N26);
and AND4 (N74, N69, N61, N61, N63);
and AND2 (N75, N8, N62);
buf BUF1 (N76, N72);
not NOT1 (N77, N68);
or OR2 (N78, N73, N8);
nand NAND3 (N79, N78, N24, N6);
or OR2 (N80, N60, N76);
and AND2 (N81, N58, N2);
nor NOR3 (N82, N81, N19, N24);
nor NOR4 (N83, N77, N73, N19, N1);
buf BUF1 (N84, N74);
and AND2 (N85, N64, N79);
nor NOR2 (N86, N39, N48);
nor NOR2 (N87, N52, N52);
nor NOR2 (N88, N80, N22);
and AND3 (N89, N84, N56, N68);
nand NAND2 (N90, N85, N16);
and AND2 (N91, N89, N85);
xor XOR2 (N92, N91, N44);
buf BUF1 (N93, N90);
xor XOR2 (N94, N87, N61);
nor NOR4 (N95, N94, N89, N4, N8);
not NOT1 (N96, N93);
and AND4 (N97, N86, N89, N40, N17);
nand NAND3 (N98, N75, N97, N65);
and AND2 (N99, N46, N11);
or OR2 (N100, N54, N40);
xor XOR2 (N101, N83, N41);
nand NAND4 (N102, N96, N25, N13, N13);
nor NOR4 (N103, N99, N11, N39, N86);
nand NAND2 (N104, N103, N42);
nor NOR4 (N105, N100, N96, N103, N24);
or OR2 (N106, N104, N69);
nor NOR2 (N107, N95, N51);
xor XOR2 (N108, N88, N20);
or OR3 (N109, N92, N99, N41);
and AND4 (N110, N108, N73, N18, N94);
not NOT1 (N111, N109);
buf BUF1 (N112, N102);
or OR4 (N113, N98, N112, N17, N14);
not NOT1 (N114, N5);
nand NAND3 (N115, N105, N61, N60);
not NOT1 (N116, N82);
or OR4 (N117, N114, N61, N69, N25);
or OR4 (N118, N106, N59, N16, N86);
buf BUF1 (N119, N115);
and AND3 (N120, N117, N59, N80);
not NOT1 (N121, N118);
not NOT1 (N122, N70);
not NOT1 (N123, N107);
nand NAND4 (N124, N120, N59, N13, N41);
xor XOR2 (N125, N121, N7);
nand NAND3 (N126, N119, N17, N23);
not NOT1 (N127, N126);
buf BUF1 (N128, N101);
not NOT1 (N129, N111);
xor XOR2 (N130, N122, N129);
xor XOR2 (N131, N5, N74);
or OR4 (N132, N131, N22, N56, N32);
not NOT1 (N133, N124);
nor NOR3 (N134, N127, N124, N86);
xor XOR2 (N135, N125, N108);
xor XOR2 (N136, N128, N123);
or OR4 (N137, N100, N95, N123, N121);
nor NOR4 (N138, N136, N60, N17, N1);
nand NAND3 (N139, N135, N111, N75);
and AND2 (N140, N134, N7);
or OR4 (N141, N116, N117, N114, N97);
and AND3 (N142, N133, N29, N36);
xor XOR2 (N143, N130, N53);
or OR4 (N144, N142, N130, N30, N78);
not NOT1 (N145, N110);
and AND2 (N146, N144, N89);
nand NAND4 (N147, N137, N72, N59, N13);
or OR4 (N148, N147, N135, N71, N37);
nor NOR3 (N149, N132, N108, N104);
and AND4 (N150, N113, N90, N74, N130);
xor XOR2 (N151, N138, N10);
and AND4 (N152, N143, N1, N80, N8);
buf BUF1 (N153, N151);
nand NAND2 (N154, N141, N87);
buf BUF1 (N155, N152);
buf BUF1 (N156, N146);
xor XOR2 (N157, N156, N144);
nor NOR4 (N158, N145, N140, N1, N144);
nor NOR3 (N159, N98, N92, N101);
xor XOR2 (N160, N157, N16);
not NOT1 (N161, N149);
not NOT1 (N162, N155);
nand NAND4 (N163, N161, N11, N5, N3);
nand NAND4 (N164, N163, N66, N161, N122);
and AND3 (N165, N148, N33, N122);
or OR3 (N166, N159, N34, N165);
nand NAND2 (N167, N139, N150);
xor XOR2 (N168, N140, N121);
not NOT1 (N169, N122);
xor XOR2 (N170, N158, N112);
xor XOR2 (N171, N166, N112);
nor NOR2 (N172, N160, N68);
nor NOR3 (N173, N169, N72, N17);
not NOT1 (N174, N153);
xor XOR2 (N175, N171, N102);
not NOT1 (N176, N167);
xor XOR2 (N177, N168, N104);
and AND4 (N178, N170, N150, N46, N93);
buf BUF1 (N179, N178);
and AND2 (N180, N176, N40);
buf BUF1 (N181, N172);
or OR4 (N182, N179, N84, N153, N13);
and AND3 (N183, N180, N56, N48);
nor NOR3 (N184, N162, N21, N94);
nor NOR2 (N185, N164, N26);
or OR3 (N186, N175, N109, N155);
not NOT1 (N187, N182);
nand NAND3 (N188, N174, N72, N59);
nand NAND4 (N189, N181, N98, N22, N76);
buf BUF1 (N190, N183);
xor XOR2 (N191, N187, N76);
buf BUF1 (N192, N177);
and AND2 (N193, N154, N166);
xor XOR2 (N194, N193, N154);
nor NOR4 (N195, N184, N98, N106, N61);
nor NOR3 (N196, N188, N120, N40);
xor XOR2 (N197, N195, N91);
xor XOR2 (N198, N186, N57);
and AND2 (N199, N198, N34);
nand NAND3 (N200, N191, N166, N194);
nor NOR4 (N201, N161, N62, N155, N154);
and AND4 (N202, N201, N147, N57, N75);
not NOT1 (N203, N192);
nand NAND4 (N204, N200, N195, N68, N202);
xor XOR2 (N205, N109, N138);
nand NAND2 (N206, N173, N39);
xor XOR2 (N207, N196, N109);
and AND3 (N208, N205, N71, N153);
nor NOR3 (N209, N203, N64, N200);
not NOT1 (N210, N207);
or OR4 (N211, N197, N93, N127, N81);
xor XOR2 (N212, N185, N66);
buf BUF1 (N213, N204);
xor XOR2 (N214, N213, N183);
not NOT1 (N215, N206);
or OR4 (N216, N189, N6, N19, N50);
or OR3 (N217, N208, N68, N89);
nand NAND4 (N218, N210, N72, N208, N176);
buf BUF1 (N219, N209);
nor NOR3 (N220, N218, N66, N20);
nor NOR2 (N221, N219, N15);
and AND4 (N222, N220, N15, N55, N200);
nor NOR4 (N223, N217, N92, N129, N74);
or OR3 (N224, N212, N38, N204);
buf BUF1 (N225, N190);
xor XOR2 (N226, N222, N18);
nor NOR2 (N227, N216, N142);
nor NOR2 (N228, N223, N68);
or OR3 (N229, N214, N113, N167);
nor NOR2 (N230, N211, N110);
or OR4 (N231, N226, N50, N95, N205);
not NOT1 (N232, N230);
or OR4 (N233, N225, N175, N7, N53);
nand NAND3 (N234, N224, N104, N158);
and AND2 (N235, N234, N106);
nor NOR2 (N236, N233, N147);
nand NAND3 (N237, N199, N132, N15);
buf BUF1 (N238, N231);
xor XOR2 (N239, N221, N122);
xor XOR2 (N240, N237, N99);
nand NAND2 (N241, N235, N144);
nor NOR2 (N242, N238, N95);
nor NOR4 (N243, N215, N7, N228, N239);
or OR2 (N244, N168, N200);
not NOT1 (N245, N21);
nand NAND3 (N246, N243, N6, N232);
not NOT1 (N247, N10);
buf BUF1 (N248, N246);
xor XOR2 (N249, N247, N142);
buf BUF1 (N250, N227);
and AND4 (N251, N236, N76, N181, N107);
and AND4 (N252, N250, N228, N58, N249);
nand NAND2 (N253, N52, N124);
not NOT1 (N254, N241);
buf BUF1 (N255, N253);
buf BUF1 (N256, N229);
buf BUF1 (N257, N240);
buf BUF1 (N258, N244);
or OR4 (N259, N252, N45, N11, N159);
xor XOR2 (N260, N256, N214);
nor NOR2 (N261, N259, N42);
nor NOR4 (N262, N261, N79, N103, N178);
buf BUF1 (N263, N248);
xor XOR2 (N264, N263, N250);
xor XOR2 (N265, N254, N129);
not NOT1 (N266, N258);
and AND3 (N267, N264, N176, N71);
nor NOR3 (N268, N266, N177, N12);
xor XOR2 (N269, N268, N173);
or OR2 (N270, N245, N246);
xor XOR2 (N271, N270, N62);
nand NAND3 (N272, N260, N26, N57);
or OR4 (N273, N271, N97, N227, N263);
xor XOR2 (N274, N242, N189);
and AND3 (N275, N269, N251, N153);
and AND2 (N276, N40, N148);
not NOT1 (N277, N262);
buf BUF1 (N278, N275);
buf BUF1 (N279, N257);
xor XOR2 (N280, N267, N261);
and AND4 (N281, N278, N190, N161, N82);
buf BUF1 (N282, N280);
not NOT1 (N283, N274);
xor XOR2 (N284, N283, N150);
or OR3 (N285, N255, N148, N58);
xor XOR2 (N286, N273, N127);
nand NAND3 (N287, N286, N94, N153);
and AND4 (N288, N272, N6, N67, N110);
nor NOR3 (N289, N287, N152, N210);
and AND4 (N290, N277, N245, N259, N214);
nand NAND2 (N291, N279, N220);
not NOT1 (N292, N288);
and AND3 (N293, N285, N128, N83);
or OR2 (N294, N292, N194);
and AND3 (N295, N276, N90, N245);
or OR3 (N296, N291, N25, N205);
nand NAND4 (N297, N293, N3, N218, N16);
and AND3 (N298, N289, N60, N124);
and AND3 (N299, N284, N84, N273);
nand NAND2 (N300, N299, N46);
buf BUF1 (N301, N294);
nand NAND3 (N302, N298, N42, N204);
and AND4 (N303, N296, N205, N171, N245);
buf BUF1 (N304, N302);
buf BUF1 (N305, N301);
or OR3 (N306, N290, N155, N157);
nor NOR3 (N307, N300, N134, N285);
xor XOR2 (N308, N297, N198);
and AND3 (N309, N304, N278, N85);
buf BUF1 (N310, N308);
not NOT1 (N311, N306);
and AND3 (N312, N281, N280, N126);
not NOT1 (N313, N307);
buf BUF1 (N314, N311);
nand NAND3 (N315, N313, N308, N38);
and AND4 (N316, N303, N99, N29, N284);
xor XOR2 (N317, N295, N273);
nor NOR4 (N318, N309, N119, N104, N173);
nand NAND2 (N319, N314, N110);
or OR4 (N320, N282, N13, N99, N162);
nand NAND2 (N321, N310, N88);
nand NAND2 (N322, N320, N144);
or OR4 (N323, N316, N307, N218, N262);
not NOT1 (N324, N305);
and AND2 (N325, N324, N246);
not NOT1 (N326, N322);
nor NOR4 (N327, N265, N290, N18, N131);
not NOT1 (N328, N317);
not NOT1 (N329, N326);
or OR4 (N330, N325, N327, N314, N281);
nor NOR4 (N331, N328, N236, N227, N131);
xor XOR2 (N332, N124, N50);
nor NOR2 (N333, N315, N15);
nand NAND3 (N334, N332, N136, N206);
not NOT1 (N335, N321);
nand NAND3 (N336, N333, N278, N238);
and AND4 (N337, N336, N187, N73, N192);
nand NAND4 (N338, N323, N243, N172, N47);
buf BUF1 (N339, N338);
buf BUF1 (N340, N335);
and AND2 (N341, N319, N140);
xor XOR2 (N342, N312, N297);
xor XOR2 (N343, N330, N122);
or OR3 (N344, N342, N269, N101);
buf BUF1 (N345, N331);
or OR4 (N346, N329, N120, N333, N45);
and AND3 (N347, N337, N335, N13);
not NOT1 (N348, N340);
xor XOR2 (N349, N347, N10);
xor XOR2 (N350, N348, N137);
or OR3 (N351, N346, N252, N163);
buf BUF1 (N352, N349);
nand NAND2 (N353, N339, N42);
buf BUF1 (N354, N353);
not NOT1 (N355, N350);
and AND3 (N356, N351, N26, N231);
not NOT1 (N357, N352);
nand NAND2 (N358, N344, N182);
or OR4 (N359, N343, N226, N217, N134);
or OR2 (N360, N359, N55);
buf BUF1 (N361, N357);
or OR4 (N362, N354, N59, N180, N3);
nand NAND4 (N363, N356, N300, N161, N250);
and AND3 (N364, N361, N16, N176);
not NOT1 (N365, N345);
or OR2 (N366, N355, N357);
buf BUF1 (N367, N362);
nor NOR2 (N368, N318, N38);
or OR4 (N369, N360, N122, N48, N156);
buf BUF1 (N370, N358);
xor XOR2 (N371, N364, N359);
not NOT1 (N372, N370);
and AND2 (N373, N365, N191);
not NOT1 (N374, N363);
nand NAND3 (N375, N373, N154, N263);
xor XOR2 (N376, N341, N6);
xor XOR2 (N377, N334, N6);
xor XOR2 (N378, N374, N40);
nand NAND4 (N379, N372, N254, N279, N353);
nand NAND2 (N380, N366, N41);
xor XOR2 (N381, N380, N291);
or OR4 (N382, N376, N216, N124, N62);
buf BUF1 (N383, N381);
nor NOR4 (N384, N367, N355, N5, N26);
or OR3 (N385, N371, N352, N48);
buf BUF1 (N386, N383);
nand NAND3 (N387, N382, N370, N196);
buf BUF1 (N388, N369);
or OR2 (N389, N377, N266);
buf BUF1 (N390, N379);
or OR4 (N391, N368, N227, N221, N220);
not NOT1 (N392, N388);
not NOT1 (N393, N389);
nand NAND4 (N394, N392, N139, N351, N245);
and AND4 (N395, N386, N308, N252, N45);
xor XOR2 (N396, N394, N95);
buf BUF1 (N397, N375);
and AND4 (N398, N397, N337, N263, N84);
and AND2 (N399, N391, N151);
or OR4 (N400, N399, N164, N291, N12);
buf BUF1 (N401, N398);
nand NAND3 (N402, N378, N253, N186);
nor NOR4 (N403, N385, N36, N72, N95);
and AND2 (N404, N402, N334);
nor NOR4 (N405, N393, N289, N90, N107);
xor XOR2 (N406, N403, N286);
nand NAND4 (N407, N387, N251, N384, N85);
and AND4 (N408, N46, N115, N279, N265);
xor XOR2 (N409, N390, N56);
or OR3 (N410, N408, N51, N106);
and AND2 (N411, N410, N158);
nand NAND3 (N412, N404, N12, N275);
nand NAND3 (N413, N400, N274, N340);
nor NOR4 (N414, N409, N75, N244, N354);
nor NOR2 (N415, N401, N83);
nor NOR4 (N416, N415, N2, N143, N153);
or OR3 (N417, N406, N22, N135);
not NOT1 (N418, N396);
xor XOR2 (N419, N405, N151);
nand NAND2 (N420, N416, N245);
nand NAND2 (N421, N420, N28);
nor NOR4 (N422, N407, N230, N216, N344);
not NOT1 (N423, N412);
not NOT1 (N424, N422);
not NOT1 (N425, N419);
or OR3 (N426, N414, N182, N332);
or OR2 (N427, N418, N312);
xor XOR2 (N428, N411, N20);
nand NAND3 (N429, N428, N275, N114);
not NOT1 (N430, N423);
buf BUF1 (N431, N395);
nor NOR3 (N432, N426, N429, N7);
and AND3 (N433, N178, N49, N365);
nor NOR4 (N434, N413, N256, N276, N172);
or OR4 (N435, N417, N122, N291, N103);
not NOT1 (N436, N434);
nand NAND3 (N437, N431, N148, N89);
not NOT1 (N438, N424);
not NOT1 (N439, N433);
nand NAND3 (N440, N435, N20, N142);
and AND3 (N441, N438, N438, N155);
not NOT1 (N442, N432);
and AND4 (N443, N437, N325, N184, N301);
nor NOR3 (N444, N441, N68, N15);
xor XOR2 (N445, N443, N371);
nand NAND4 (N446, N427, N101, N39, N427);
nor NOR4 (N447, N444, N162, N27, N7);
and AND3 (N448, N440, N238, N247);
and AND2 (N449, N421, N250);
nand NAND3 (N450, N442, N67, N334);
xor XOR2 (N451, N445, N410);
buf BUF1 (N452, N451);
nor NOR2 (N453, N446, N97);
buf BUF1 (N454, N452);
and AND4 (N455, N436, N201, N141, N391);
nand NAND3 (N456, N447, N342, N210);
nand NAND2 (N457, N453, N295);
nor NOR2 (N458, N425, N116);
not NOT1 (N459, N430);
not NOT1 (N460, N439);
buf BUF1 (N461, N457);
or OR4 (N462, N454, N144, N94, N387);
and AND3 (N463, N460, N345, N12);
or OR2 (N464, N456, N283);
not NOT1 (N465, N449);
nor NOR3 (N466, N463, N285, N313);
and AND4 (N467, N461, N455, N434, N179);
or OR3 (N468, N326, N332, N171);
nand NAND4 (N469, N462, N309, N240, N329);
xor XOR2 (N470, N458, N375);
not NOT1 (N471, N448);
nand NAND4 (N472, N469, N279, N67, N303);
or OR4 (N473, N465, N184, N208, N192);
nand NAND3 (N474, N466, N359, N295);
nand NAND3 (N475, N468, N203, N291);
nor NOR2 (N476, N467, N331);
nor NOR4 (N477, N450, N152, N470, N341);
or OR2 (N478, N361, N263);
nand NAND3 (N479, N471, N158, N417);
nor NOR3 (N480, N464, N228, N337);
nor NOR4 (N481, N476, N397, N444, N453);
or OR2 (N482, N472, N241);
buf BUF1 (N483, N478);
and AND4 (N484, N475, N182, N410, N85);
and AND4 (N485, N480, N76, N166, N439);
or OR3 (N486, N483, N328, N307);
and AND3 (N487, N481, N376, N218);
xor XOR2 (N488, N484, N293);
and AND4 (N489, N479, N236, N24, N246);
or OR3 (N490, N473, N313, N341);
not NOT1 (N491, N482);
buf BUF1 (N492, N491);
nand NAND3 (N493, N490, N485, N361);
xor XOR2 (N494, N481, N181);
buf BUF1 (N495, N474);
nand NAND2 (N496, N494, N92);
nor NOR3 (N497, N488, N136, N219);
nand NAND3 (N498, N489, N433, N421);
xor XOR2 (N499, N487, N421);
xor XOR2 (N500, N477, N285);
and AND3 (N501, N492, N462, N28);
not NOT1 (N502, N496);
not NOT1 (N503, N493);
buf BUF1 (N504, N495);
or OR3 (N505, N498, N430, N165);
nor NOR2 (N506, N502, N418);
xor XOR2 (N507, N459, N375);
and AND2 (N508, N505, N161);
buf BUF1 (N509, N497);
or OR2 (N510, N500, N335);
and AND2 (N511, N509, N330);
or OR2 (N512, N503, N170);
nor NOR3 (N513, N506, N272, N269);
or OR3 (N514, N510, N264, N394);
or OR2 (N515, N513, N42);
or OR3 (N516, N501, N71, N79);
nand NAND3 (N517, N507, N268, N222);
xor XOR2 (N518, N499, N198);
nor NOR2 (N519, N486, N396);
not NOT1 (N520, N519);
buf BUF1 (N521, N520);
nand NAND2 (N522, N516, N484);
buf BUF1 (N523, N508);
nor NOR4 (N524, N523, N150, N318, N141);
nor NOR4 (N525, N512, N195, N223, N333);
xor XOR2 (N526, N515, N512);
or OR3 (N527, N517, N198, N492);
and AND4 (N528, N526, N114, N93, N489);
and AND3 (N529, N522, N283, N421);
nor NOR2 (N530, N511, N171);
xor XOR2 (N531, N525, N203);
nor NOR3 (N532, N528, N323, N531);
not NOT1 (N533, N118);
nor NOR2 (N534, N533, N532);
nor NOR3 (N535, N504, N301, N144);
not NOT1 (N536, N104);
not NOT1 (N537, N527);
not NOT1 (N538, N534);
and AND3 (N539, N530, N406, N307);
nor NOR3 (N540, N535, N268, N18);
nor NOR4 (N541, N518, N199, N14, N370);
or OR3 (N542, N524, N50, N539);
not NOT1 (N543, N174);
buf BUF1 (N544, N514);
buf BUF1 (N545, N529);
nor NOR4 (N546, N537, N512, N242, N230);
xor XOR2 (N547, N540, N364);
not NOT1 (N548, N542);
buf BUF1 (N549, N538);
xor XOR2 (N550, N545, N262);
nand NAND3 (N551, N521, N472, N430);
and AND4 (N552, N548, N248, N384, N303);
buf BUF1 (N553, N543);
nand NAND4 (N554, N549, N118, N62, N126);
buf BUF1 (N555, N536);
xor XOR2 (N556, N551, N369);
and AND2 (N557, N550, N372);
buf BUF1 (N558, N544);
nor NOR4 (N559, N552, N317, N325, N476);
not NOT1 (N560, N559);
buf BUF1 (N561, N556);
nor NOR4 (N562, N547, N33, N318, N199);
buf BUF1 (N563, N557);
nand NAND2 (N564, N561, N463);
or OR2 (N565, N563, N7);
nand NAND2 (N566, N553, N268);
and AND3 (N567, N558, N322, N304);
buf BUF1 (N568, N565);
and AND2 (N569, N567, N325);
nor NOR3 (N570, N569, N299, N515);
or OR3 (N571, N568, N496, N405);
not NOT1 (N572, N541);
not NOT1 (N573, N571);
and AND3 (N574, N555, N16, N20);
xor XOR2 (N575, N566, N227);
buf BUF1 (N576, N574);
xor XOR2 (N577, N573, N379);
xor XOR2 (N578, N564, N259);
and AND4 (N579, N554, N109, N79, N249);
nand NAND4 (N580, N560, N83, N357, N464);
buf BUF1 (N581, N577);
not NOT1 (N582, N581);
nor NOR4 (N583, N580, N17, N24, N344);
nand NAND4 (N584, N572, N290, N161, N296);
xor XOR2 (N585, N578, N27);
and AND4 (N586, N585, N118, N78, N217);
buf BUF1 (N587, N576);
xor XOR2 (N588, N562, N334);
nand NAND4 (N589, N582, N495, N281, N420);
nor NOR2 (N590, N575, N478);
nor NOR2 (N591, N584, N439);
nor NOR4 (N592, N546, N414, N485, N135);
buf BUF1 (N593, N583);
buf BUF1 (N594, N586);
or OR3 (N595, N579, N155, N64);
xor XOR2 (N596, N589, N285);
nor NOR2 (N597, N595, N182);
xor XOR2 (N598, N587, N541);
and AND3 (N599, N591, N120, N477);
and AND2 (N600, N598, N88);
nand NAND4 (N601, N594, N266, N21, N288);
xor XOR2 (N602, N570, N599);
nand NAND4 (N603, N343, N324, N27, N319);
and AND2 (N604, N596, N239);
and AND3 (N605, N601, N570, N41);
buf BUF1 (N606, N597);
and AND2 (N607, N600, N71);
not NOT1 (N608, N604);
xor XOR2 (N609, N607, N95);
xor XOR2 (N610, N603, N115);
xor XOR2 (N611, N608, N430);
nand NAND2 (N612, N611, N30);
and AND3 (N613, N609, N164, N275);
not NOT1 (N614, N592);
and AND3 (N615, N590, N575, N419);
buf BUF1 (N616, N606);
or OR2 (N617, N612, N215);
nor NOR2 (N618, N615, N56);
or OR2 (N619, N588, N32);
not NOT1 (N620, N593);
or OR4 (N621, N610, N483, N413, N130);
nand NAND3 (N622, N614, N153, N600);
and AND3 (N623, N605, N248, N161);
nor NOR3 (N624, N620, N427, N512);
xor XOR2 (N625, N622, N245);
nor NOR2 (N626, N623, N435);
and AND2 (N627, N602, N178);
not NOT1 (N628, N616);
xor XOR2 (N629, N617, N363);
nor NOR4 (N630, N613, N17, N454, N179);
xor XOR2 (N631, N630, N45);
not NOT1 (N632, N619);
nor NOR2 (N633, N629, N348);
buf BUF1 (N634, N625);
xor XOR2 (N635, N628, N110);
not NOT1 (N636, N632);
nor NOR2 (N637, N636, N541);
nor NOR2 (N638, N618, N300);
not NOT1 (N639, N638);
or OR2 (N640, N634, N382);
nand NAND4 (N641, N639, N286, N562, N337);
and AND2 (N642, N621, N600);
nor NOR3 (N643, N624, N83, N465);
nor NOR3 (N644, N642, N231, N264);
and AND3 (N645, N635, N591, N218);
not NOT1 (N646, N641);
nand NAND2 (N647, N646, N226);
buf BUF1 (N648, N637);
nor NOR4 (N649, N626, N144, N436, N302);
and AND3 (N650, N644, N96, N473);
xor XOR2 (N651, N650, N126);
xor XOR2 (N652, N633, N269);
buf BUF1 (N653, N648);
nor NOR3 (N654, N643, N136, N274);
buf BUF1 (N655, N640);
or OR4 (N656, N649, N77, N90, N66);
buf BUF1 (N657, N647);
not NOT1 (N658, N655);
not NOT1 (N659, N656);
xor XOR2 (N660, N654, N590);
nor NOR4 (N661, N645, N537, N321, N256);
and AND3 (N662, N660, N395, N214);
or OR2 (N663, N651, N240);
xor XOR2 (N664, N661, N180);
nor NOR4 (N665, N662, N134, N8, N363);
and AND2 (N666, N631, N247);
nand NAND3 (N667, N666, N373, N600);
nor NOR4 (N668, N657, N168, N454, N324);
xor XOR2 (N669, N663, N410);
nand NAND3 (N670, N665, N352, N633);
buf BUF1 (N671, N627);
nand NAND3 (N672, N667, N186, N83);
and AND3 (N673, N671, N218, N250);
or OR4 (N674, N672, N45, N163, N30);
nand NAND4 (N675, N673, N104, N579, N344);
not NOT1 (N676, N653);
xor XOR2 (N677, N658, N290);
xor XOR2 (N678, N670, N268);
nor NOR3 (N679, N676, N645, N643);
buf BUF1 (N680, N652);
xor XOR2 (N681, N659, N109);
not NOT1 (N682, N664);
nand NAND3 (N683, N682, N50, N79);
nand NAND2 (N684, N669, N67);
nand NAND3 (N685, N678, N634, N661);
not NOT1 (N686, N683);
or OR4 (N687, N668, N479, N482, N479);
nor NOR2 (N688, N685, N484);
or OR4 (N689, N687, N475, N535, N215);
and AND4 (N690, N684, N571, N194, N407);
not NOT1 (N691, N690);
or OR4 (N692, N689, N389, N675, N376);
nor NOR3 (N693, N580, N249, N170);
or OR2 (N694, N681, N114);
not NOT1 (N695, N688);
not NOT1 (N696, N691);
buf BUF1 (N697, N674);
not NOT1 (N698, N692);
xor XOR2 (N699, N679, N427);
xor XOR2 (N700, N686, N315);
nand NAND4 (N701, N697, N686, N295, N561);
nor NOR3 (N702, N698, N33, N237);
nor NOR3 (N703, N694, N170, N583);
and AND4 (N704, N702, N49, N472, N323);
and AND2 (N705, N677, N503);
nor NOR2 (N706, N703, N644);
buf BUF1 (N707, N695);
buf BUF1 (N708, N704);
buf BUF1 (N709, N696);
xor XOR2 (N710, N701, N634);
not NOT1 (N711, N700);
buf BUF1 (N712, N680);
and AND3 (N713, N712, N609, N420);
nand NAND3 (N714, N707, N574, N712);
and AND3 (N715, N710, N676, N31);
not NOT1 (N716, N714);
nor NOR4 (N717, N716, N654, N169, N666);
buf BUF1 (N718, N693);
and AND2 (N719, N717, N502);
nand NAND3 (N720, N719, N145, N553);
nor NOR4 (N721, N709, N580, N119, N666);
xor XOR2 (N722, N718, N664);
buf BUF1 (N723, N715);
nand NAND2 (N724, N713, N332);
and AND4 (N725, N721, N230, N541, N539);
and AND4 (N726, N722, N258, N693, N644);
xor XOR2 (N727, N726, N599);
and AND3 (N728, N711, N62, N172);
buf BUF1 (N729, N724);
buf BUF1 (N730, N708);
xor XOR2 (N731, N730, N594);
buf BUF1 (N732, N725);
buf BUF1 (N733, N732);
nand NAND4 (N734, N706, N431, N705, N558);
buf BUF1 (N735, N138);
and AND4 (N736, N728, N576, N708, N436);
buf BUF1 (N737, N723);
nor NOR4 (N738, N731, N514, N723, N441);
or OR4 (N739, N734, N473, N569, N647);
buf BUF1 (N740, N720);
xor XOR2 (N741, N735, N474);
buf BUF1 (N742, N739);
buf BUF1 (N743, N727);
or OR3 (N744, N743, N307, N140);
and AND4 (N745, N744, N163, N299, N456);
nor NOR2 (N746, N733, N369);
not NOT1 (N747, N741);
not NOT1 (N748, N742);
nand NAND3 (N749, N699, N454, N413);
not NOT1 (N750, N729);
nand NAND3 (N751, N748, N512, N499);
xor XOR2 (N752, N749, N26);
xor XOR2 (N753, N738, N238);
xor XOR2 (N754, N750, N401);
and AND3 (N755, N754, N67, N526);
buf BUF1 (N756, N737);
not NOT1 (N757, N740);
buf BUF1 (N758, N736);
nand NAND4 (N759, N755, N163, N78, N312);
buf BUF1 (N760, N752);
and AND2 (N761, N757, N662);
xor XOR2 (N762, N753, N541);
not NOT1 (N763, N761);
nor NOR2 (N764, N745, N258);
nand NAND2 (N765, N747, N152);
nand NAND4 (N766, N759, N549, N227, N181);
xor XOR2 (N767, N764, N469);
nand NAND2 (N768, N765, N603);
and AND4 (N769, N766, N282, N639, N2);
not NOT1 (N770, N768);
or OR2 (N771, N756, N83);
not NOT1 (N772, N760);
xor XOR2 (N773, N762, N123);
xor XOR2 (N774, N763, N55);
nor NOR3 (N775, N767, N16, N150);
or OR3 (N776, N772, N259, N250);
and AND2 (N777, N774, N256);
nor NOR3 (N778, N769, N269, N59);
buf BUF1 (N779, N775);
nand NAND2 (N780, N771, N441);
not NOT1 (N781, N751);
not NOT1 (N782, N758);
nor NOR4 (N783, N770, N160, N775, N106);
nor NOR2 (N784, N778, N574);
buf BUF1 (N785, N776);
xor XOR2 (N786, N783, N460);
nand NAND4 (N787, N779, N311, N703, N272);
xor XOR2 (N788, N746, N288);
xor XOR2 (N789, N780, N566);
nor NOR3 (N790, N788, N73, N602);
buf BUF1 (N791, N781);
not NOT1 (N792, N789);
nand NAND2 (N793, N782, N221);
buf BUF1 (N794, N790);
not NOT1 (N795, N791);
xor XOR2 (N796, N785, N537);
xor XOR2 (N797, N795, N324);
not NOT1 (N798, N792);
buf BUF1 (N799, N786);
or OR3 (N800, N796, N283, N680);
not NOT1 (N801, N794);
nand NAND4 (N802, N787, N738, N325, N64);
not NOT1 (N803, N793);
and AND2 (N804, N799, N425);
buf BUF1 (N805, N773);
nor NOR3 (N806, N805, N719, N316);
not NOT1 (N807, N804);
and AND3 (N808, N801, N231, N636);
not NOT1 (N809, N807);
and AND4 (N810, N802, N94, N795, N732);
xor XOR2 (N811, N810, N701);
xor XOR2 (N812, N806, N399);
buf BUF1 (N813, N809);
not NOT1 (N814, N797);
and AND4 (N815, N784, N177, N169, N229);
or OR3 (N816, N815, N496, N432);
and AND4 (N817, N798, N110, N327, N595);
nand NAND3 (N818, N816, N271, N498);
not NOT1 (N819, N777);
xor XOR2 (N820, N803, N80);
and AND4 (N821, N820, N628, N183, N157);
and AND2 (N822, N819, N20);
or OR4 (N823, N812, N126, N578, N172);
xor XOR2 (N824, N808, N209);
nand NAND2 (N825, N800, N600);
not NOT1 (N826, N811);
or OR4 (N827, N826, N216, N448, N565);
xor XOR2 (N828, N822, N195);
nand NAND4 (N829, N814, N789, N57, N273);
nor NOR4 (N830, N823, N777, N565, N179);
nand NAND3 (N831, N824, N166, N677);
nor NOR3 (N832, N830, N454, N659);
and AND2 (N833, N828, N180);
nor NOR3 (N834, N821, N35, N302);
or OR2 (N835, N833, N442);
not NOT1 (N836, N818);
and AND4 (N837, N835, N22, N94, N254);
not NOT1 (N838, N836);
buf BUF1 (N839, N837);
nor NOR4 (N840, N817, N342, N90, N830);
xor XOR2 (N841, N829, N597);
buf BUF1 (N842, N841);
xor XOR2 (N843, N834, N244);
buf BUF1 (N844, N842);
nor NOR4 (N845, N839, N589, N775, N799);
buf BUF1 (N846, N832);
nor NOR3 (N847, N827, N562, N272);
buf BUF1 (N848, N846);
nor NOR2 (N849, N838, N683);
buf BUF1 (N850, N840);
or OR4 (N851, N848, N384, N489, N141);
xor XOR2 (N852, N847, N78);
nor NOR2 (N853, N831, N798);
or OR2 (N854, N852, N652);
buf BUF1 (N855, N843);
or OR3 (N856, N855, N810, N370);
and AND2 (N857, N845, N134);
buf BUF1 (N858, N849);
buf BUF1 (N859, N813);
and AND4 (N860, N854, N309, N16, N184);
or OR2 (N861, N850, N411);
nor NOR4 (N862, N858, N153, N741, N399);
buf BUF1 (N863, N844);
buf BUF1 (N864, N853);
nand NAND3 (N865, N859, N550, N516);
buf BUF1 (N866, N860);
buf BUF1 (N867, N866);
xor XOR2 (N868, N857, N189);
or OR2 (N869, N867, N529);
nand NAND4 (N870, N865, N193, N134, N821);
or OR3 (N871, N862, N711, N339);
buf BUF1 (N872, N868);
xor XOR2 (N873, N825, N228);
xor XOR2 (N874, N870, N693);
nand NAND2 (N875, N863, N578);
nor NOR4 (N876, N864, N152, N639, N383);
xor XOR2 (N877, N875, N535);
nand NAND4 (N878, N873, N193, N276, N393);
nand NAND3 (N879, N869, N200, N84);
xor XOR2 (N880, N856, N682);
nand NAND2 (N881, N872, N770);
xor XOR2 (N882, N879, N816);
and AND3 (N883, N874, N381, N881);
nor NOR3 (N884, N868, N696, N464);
or OR3 (N885, N861, N826, N614);
not NOT1 (N886, N884);
buf BUF1 (N887, N882);
xor XOR2 (N888, N887, N435);
nand NAND3 (N889, N851, N868, N572);
not NOT1 (N890, N883);
or OR2 (N891, N886, N491);
nor NOR4 (N892, N888, N323, N856, N877);
nor NOR3 (N893, N606, N372, N865);
nor NOR3 (N894, N890, N721, N95);
not NOT1 (N895, N892);
xor XOR2 (N896, N894, N87);
nor NOR4 (N897, N878, N527, N45, N182);
xor XOR2 (N898, N895, N787);
buf BUF1 (N899, N893);
not NOT1 (N900, N885);
and AND4 (N901, N889, N125, N790, N155);
not NOT1 (N902, N891);
nor NOR3 (N903, N900, N585, N581);
not NOT1 (N904, N902);
xor XOR2 (N905, N880, N36);
not NOT1 (N906, N901);
buf BUF1 (N907, N898);
nor NOR2 (N908, N899, N645);
xor XOR2 (N909, N903, N318);
not NOT1 (N910, N905);
xor XOR2 (N911, N896, N179);
xor XOR2 (N912, N904, N57);
nor NOR2 (N913, N876, N784);
not NOT1 (N914, N908);
nand NAND3 (N915, N911, N799, N419);
buf BUF1 (N916, N910);
buf BUF1 (N917, N909);
not NOT1 (N918, N871);
buf BUF1 (N919, N915);
and AND3 (N920, N912, N648, N12);
or OR2 (N921, N906, N560);
nor NOR4 (N922, N920, N683, N517, N239);
nand NAND2 (N923, N921, N316);
and AND4 (N924, N922, N99, N231, N896);
nor NOR2 (N925, N897, N324);
nor NOR3 (N926, N913, N604, N53);
and AND2 (N927, N914, N712);
xor XOR2 (N928, N919, N112);
nor NOR4 (N929, N926, N908, N683, N601);
buf BUF1 (N930, N916);
buf BUF1 (N931, N927);
nor NOR2 (N932, N918, N562);
buf BUF1 (N933, N931);
buf BUF1 (N934, N929);
xor XOR2 (N935, N907, N714);
buf BUF1 (N936, N935);
xor XOR2 (N937, N930, N475);
not NOT1 (N938, N924);
xor XOR2 (N939, N932, N934);
buf BUF1 (N940, N216);
nand NAND3 (N941, N923, N353, N412);
buf BUF1 (N942, N936);
nor NOR3 (N943, N938, N281, N346);
or OR4 (N944, N937, N480, N4, N334);
nand NAND3 (N945, N933, N166, N226);
and AND2 (N946, N917, N500);
and AND3 (N947, N943, N179, N116);
buf BUF1 (N948, N946);
nor NOR2 (N949, N947, N329);
and AND3 (N950, N941, N17, N150);
or OR3 (N951, N940, N633, N525);
buf BUF1 (N952, N942);
not NOT1 (N953, N948);
nor NOR3 (N954, N950, N464, N814);
and AND4 (N955, N952, N256, N786, N460);
nand NAND4 (N956, N944, N502, N663, N365);
buf BUF1 (N957, N939);
and AND2 (N958, N945, N646);
buf BUF1 (N959, N928);
and AND4 (N960, N953, N807, N536, N317);
xor XOR2 (N961, N957, N322);
or OR3 (N962, N955, N601, N734);
xor XOR2 (N963, N956, N892);
and AND4 (N964, N960, N156, N186, N845);
xor XOR2 (N965, N949, N71);
and AND3 (N966, N962, N803, N7);
nand NAND2 (N967, N966, N455);
not NOT1 (N968, N951);
or OR2 (N969, N963, N220);
or OR2 (N970, N958, N793);
or OR3 (N971, N961, N769, N457);
and AND3 (N972, N925, N88, N43);
not NOT1 (N973, N959);
not NOT1 (N974, N970);
xor XOR2 (N975, N971, N44);
or OR3 (N976, N967, N688, N443);
buf BUF1 (N977, N954);
or OR2 (N978, N977, N811);
buf BUF1 (N979, N974);
buf BUF1 (N980, N969);
not NOT1 (N981, N975);
xor XOR2 (N982, N979, N399);
buf BUF1 (N983, N980);
or OR3 (N984, N981, N963, N264);
and AND4 (N985, N982, N563, N521, N820);
nor NOR2 (N986, N965, N611);
buf BUF1 (N987, N986);
xor XOR2 (N988, N983, N572);
and AND4 (N989, N968, N330, N279, N856);
and AND4 (N990, N978, N232, N59, N97);
and AND4 (N991, N990, N119, N499, N156);
nand NAND3 (N992, N964, N708, N188);
and AND4 (N993, N992, N758, N860, N710);
nor NOR3 (N994, N985, N230, N717);
and AND4 (N995, N991, N31, N788, N831);
xor XOR2 (N996, N993, N359);
xor XOR2 (N997, N994, N60);
and AND3 (N998, N989, N523, N153);
and AND3 (N999, N995, N536, N3);
buf BUF1 (N1000, N988);
buf BUF1 (N1001, N996);
not NOT1 (N1002, N976);
xor XOR2 (N1003, N987, N936);
nor NOR4 (N1004, N997, N215, N178, N847);
xor XOR2 (N1005, N973, N180);
or OR3 (N1006, N998, N795, N555);
nand NAND3 (N1007, N1004, N260, N944);
buf BUF1 (N1008, N1003);
xor XOR2 (N1009, N1005, N346);
not NOT1 (N1010, N999);
nor NOR4 (N1011, N984, N793, N770, N902);
nor NOR2 (N1012, N972, N975);
buf BUF1 (N1013, N1006);
xor XOR2 (N1014, N1001, N969);
or OR3 (N1015, N1008, N388, N461);
or OR4 (N1016, N1000, N336, N766, N378);
and AND4 (N1017, N1009, N100, N833, N678);
or OR3 (N1018, N1002, N734, N389);
or OR2 (N1019, N1015, N986);
xor XOR2 (N1020, N1007, N477);
not NOT1 (N1021, N1018);
buf BUF1 (N1022, N1013);
or OR4 (N1023, N1012, N317, N226, N697);
buf BUF1 (N1024, N1010);
buf BUF1 (N1025, N1019);
or OR3 (N1026, N1025, N793, N181);
buf BUF1 (N1027, N1021);
not NOT1 (N1028, N1027);
and AND4 (N1029, N1017, N687, N392, N209);
or OR2 (N1030, N1011, N296);
nor NOR4 (N1031, N1022, N746, N571, N447);
or OR2 (N1032, N1026, N487);
or OR3 (N1033, N1028, N968, N708);
buf BUF1 (N1034, N1020);
not NOT1 (N1035, N1023);
nand NAND3 (N1036, N1031, N222, N962);
or OR3 (N1037, N1024, N471, N918);
nor NOR4 (N1038, N1037, N259, N728, N221);
nand NAND3 (N1039, N1036, N525, N720);
nand NAND4 (N1040, N1030, N1028, N668, N3);
and AND3 (N1041, N1032, N91, N7);
nand NAND2 (N1042, N1041, N593);
or OR3 (N1043, N1038, N531, N881);
nor NOR4 (N1044, N1035, N697, N512, N555);
or OR3 (N1045, N1039, N71, N211);
xor XOR2 (N1046, N1040, N928);
xor XOR2 (N1047, N1016, N491);
xor XOR2 (N1048, N1045, N150);
or OR2 (N1049, N1048, N94);
not NOT1 (N1050, N1046);
and AND4 (N1051, N1033, N517, N236, N757);
buf BUF1 (N1052, N1042);
not NOT1 (N1053, N1043);
nand NAND3 (N1054, N1053, N38, N436);
nand NAND2 (N1055, N1051, N195);
not NOT1 (N1056, N1049);
nand NAND2 (N1057, N1050, N278);
nor NOR2 (N1058, N1047, N1019);
xor XOR2 (N1059, N1057, N662);
buf BUF1 (N1060, N1056);
nand NAND4 (N1061, N1034, N976, N442, N287);
nand NAND2 (N1062, N1061, N524);
or OR4 (N1063, N1055, N753, N306, N859);
xor XOR2 (N1064, N1062, N850);
not NOT1 (N1065, N1052);
xor XOR2 (N1066, N1064, N649);
nor NOR3 (N1067, N1054, N1012, N388);
nand NAND2 (N1068, N1065, N573);
and AND2 (N1069, N1029, N1005);
nand NAND3 (N1070, N1067, N1008, N1011);
nor NOR3 (N1071, N1058, N9, N253);
nor NOR4 (N1072, N1071, N917, N702, N542);
nor NOR4 (N1073, N1060, N300, N579, N177);
not NOT1 (N1074, N1070);
or OR2 (N1075, N1044, N303);
and AND3 (N1076, N1069, N902, N524);
buf BUF1 (N1077, N1014);
nor NOR4 (N1078, N1073, N221, N460, N322);
xor XOR2 (N1079, N1078, N43);
xor XOR2 (N1080, N1075, N653);
nand NAND4 (N1081, N1059, N727, N564, N1073);
nand NAND3 (N1082, N1076, N277, N728);
nand NAND3 (N1083, N1068, N952, N907);
or OR3 (N1084, N1080, N177, N988);
xor XOR2 (N1085, N1083, N74);
not NOT1 (N1086, N1063);
nand NAND2 (N1087, N1066, N297);
not NOT1 (N1088, N1085);
or OR4 (N1089, N1088, N183, N672, N666);
xor XOR2 (N1090, N1079, N856);
nand NAND2 (N1091, N1077, N789);
buf BUF1 (N1092, N1074);
xor XOR2 (N1093, N1082, N865);
or OR4 (N1094, N1090, N901, N466, N168);
buf BUF1 (N1095, N1081);
xor XOR2 (N1096, N1091, N876);
nand NAND2 (N1097, N1089, N541);
nor NOR4 (N1098, N1087, N280, N1005, N589);
and AND2 (N1099, N1098, N720);
not NOT1 (N1100, N1096);
not NOT1 (N1101, N1097);
and AND2 (N1102, N1084, N972);
nand NAND4 (N1103, N1095, N340, N468, N118);
nand NAND3 (N1104, N1072, N485, N12);
not NOT1 (N1105, N1086);
nor NOR3 (N1106, N1099, N682, N479);
xor XOR2 (N1107, N1101, N259);
nor NOR4 (N1108, N1104, N580, N102, N89);
nand NAND3 (N1109, N1093, N832, N711);
xor XOR2 (N1110, N1106, N768);
not NOT1 (N1111, N1108);
nand NAND2 (N1112, N1094, N718);
nor NOR4 (N1113, N1111, N640, N815, N721);
and AND3 (N1114, N1110, N596, N874);
buf BUF1 (N1115, N1109);
xor XOR2 (N1116, N1092, N540);
buf BUF1 (N1117, N1103);
and AND3 (N1118, N1107, N663, N63);
nand NAND2 (N1119, N1105, N923);
nand NAND3 (N1120, N1115, N91, N484);
xor XOR2 (N1121, N1119, N871);
or OR3 (N1122, N1121, N28, N685);
nor NOR2 (N1123, N1120, N594);
and AND3 (N1124, N1118, N490, N319);
nor NOR3 (N1125, N1114, N721, N1112);
or OR2 (N1126, N1075, N326);
and AND3 (N1127, N1100, N1075, N901);
and AND3 (N1128, N1125, N512, N954);
buf BUF1 (N1129, N1122);
buf BUF1 (N1130, N1123);
buf BUF1 (N1131, N1128);
nor NOR2 (N1132, N1102, N200);
nor NOR3 (N1133, N1126, N84, N327);
nor NOR2 (N1134, N1124, N421);
or OR4 (N1135, N1131, N527, N498, N676);
nand NAND4 (N1136, N1135, N96, N188, N618);
buf BUF1 (N1137, N1133);
or OR3 (N1138, N1117, N290, N632);
and AND3 (N1139, N1138, N370, N190);
nand NAND4 (N1140, N1113, N319, N661, N950);
nand NAND3 (N1141, N1134, N683, N605);
buf BUF1 (N1142, N1141);
xor XOR2 (N1143, N1127, N1114);
or OR3 (N1144, N1129, N1118, N1039);
not NOT1 (N1145, N1116);
nand NAND3 (N1146, N1130, N903, N631);
or OR3 (N1147, N1140, N339, N93);
nand NAND4 (N1148, N1142, N1020, N538, N1004);
nor NOR4 (N1149, N1143, N505, N866, N227);
nand NAND4 (N1150, N1132, N226, N704, N960);
buf BUF1 (N1151, N1136);
and AND2 (N1152, N1137, N1040);
nand NAND3 (N1153, N1146, N1018, N364);
nand NAND4 (N1154, N1152, N323, N613, N77);
buf BUF1 (N1155, N1154);
or OR4 (N1156, N1150, N681, N1023, N766);
and AND2 (N1157, N1139, N890);
or OR3 (N1158, N1145, N344, N455);
or OR4 (N1159, N1144, N980, N472, N191);
nor NOR4 (N1160, N1153, N967, N736, N431);
or OR3 (N1161, N1159, N1058, N974);
xor XOR2 (N1162, N1156, N1053);
and AND2 (N1163, N1148, N986);
nor NOR4 (N1164, N1162, N169, N1159, N503);
and AND2 (N1165, N1157, N1000);
and AND3 (N1166, N1149, N731, N679);
xor XOR2 (N1167, N1166, N943);
buf BUF1 (N1168, N1161);
or OR4 (N1169, N1147, N1021, N20, N696);
and AND4 (N1170, N1165, N287, N157, N18);
nor NOR2 (N1171, N1158, N6);
xor XOR2 (N1172, N1167, N38);
not NOT1 (N1173, N1169);
and AND4 (N1174, N1155, N1079, N684, N1142);
buf BUF1 (N1175, N1174);
or OR2 (N1176, N1168, N1072);
not NOT1 (N1177, N1176);
xor XOR2 (N1178, N1160, N46);
buf BUF1 (N1179, N1164);
nand NAND2 (N1180, N1175, N949);
xor XOR2 (N1181, N1179, N732);
xor XOR2 (N1182, N1173, N949);
nor NOR3 (N1183, N1181, N191, N346);
or OR2 (N1184, N1182, N110);
not NOT1 (N1185, N1170);
buf BUF1 (N1186, N1163);
buf BUF1 (N1187, N1172);
and AND4 (N1188, N1178, N77, N875, N147);
buf BUF1 (N1189, N1183);
not NOT1 (N1190, N1186);
not NOT1 (N1191, N1187);
nand NAND3 (N1192, N1180, N942, N287);
buf BUF1 (N1193, N1185);
nand NAND2 (N1194, N1177, N486);
not NOT1 (N1195, N1184);
buf BUF1 (N1196, N1151);
or OR4 (N1197, N1192, N843, N157, N419);
xor XOR2 (N1198, N1189, N266);
nand NAND2 (N1199, N1197, N1046);
nor NOR4 (N1200, N1193, N548, N36, N39);
buf BUF1 (N1201, N1198);
not NOT1 (N1202, N1171);
not NOT1 (N1203, N1202);
or OR4 (N1204, N1195, N730, N990, N1175);
buf BUF1 (N1205, N1200);
buf BUF1 (N1206, N1188);
or OR2 (N1207, N1196, N44);
not NOT1 (N1208, N1191);
and AND4 (N1209, N1194, N7, N324, N2);
buf BUF1 (N1210, N1207);
xor XOR2 (N1211, N1209, N329);
nand NAND2 (N1212, N1211, N234);
nor NOR3 (N1213, N1212, N999, N23);
and AND4 (N1214, N1203, N591, N826, N562);
nand NAND4 (N1215, N1214, N757, N739, N329);
nor NOR2 (N1216, N1199, N947);
nor NOR4 (N1217, N1215, N745, N720, N1158);
nand NAND2 (N1218, N1213, N371);
and AND3 (N1219, N1201, N258, N1115);
buf BUF1 (N1220, N1217);
and AND2 (N1221, N1206, N362);
xor XOR2 (N1222, N1205, N586);
xor XOR2 (N1223, N1190, N1116);
not NOT1 (N1224, N1222);
buf BUF1 (N1225, N1224);
xor XOR2 (N1226, N1208, N986);
and AND4 (N1227, N1223, N360, N1, N575);
nor NOR4 (N1228, N1218, N1155, N699, N419);
nor NOR4 (N1229, N1221, N759, N830, N999);
nand NAND4 (N1230, N1216, N553, N1076, N990);
nand NAND4 (N1231, N1230, N572, N403, N895);
xor XOR2 (N1232, N1229, N1060);
buf BUF1 (N1233, N1228);
nand NAND2 (N1234, N1225, N897);
not NOT1 (N1235, N1210);
not NOT1 (N1236, N1233);
or OR2 (N1237, N1234, N664);
and AND3 (N1238, N1219, N374, N462);
or OR3 (N1239, N1237, N1181, N73);
nor NOR2 (N1240, N1227, N110);
not NOT1 (N1241, N1235);
nor NOR3 (N1242, N1232, N461, N726);
not NOT1 (N1243, N1241);
or OR4 (N1244, N1240, N767, N309, N347);
not NOT1 (N1245, N1231);
or OR2 (N1246, N1245, N186);
not NOT1 (N1247, N1239);
nor NOR3 (N1248, N1226, N465, N563);
and AND4 (N1249, N1244, N91, N168, N1014);
not NOT1 (N1250, N1248);
nor NOR4 (N1251, N1250, N178, N1149, N392);
nor NOR4 (N1252, N1238, N1036, N607, N701);
nor NOR2 (N1253, N1204, N1123);
nor NOR4 (N1254, N1253, N1013, N1161, N587);
nand NAND3 (N1255, N1220, N804, N215);
and AND4 (N1256, N1252, N565, N663, N331);
and AND4 (N1257, N1246, N742, N864, N965);
or OR2 (N1258, N1251, N524);
xor XOR2 (N1259, N1249, N1249);
xor XOR2 (N1260, N1255, N1101);
or OR3 (N1261, N1259, N1123, N1115);
xor XOR2 (N1262, N1257, N1015);
buf BUF1 (N1263, N1247);
buf BUF1 (N1264, N1260);
not NOT1 (N1265, N1262);
xor XOR2 (N1266, N1236, N235);
nand NAND2 (N1267, N1243, N254);
buf BUF1 (N1268, N1256);
or OR3 (N1269, N1261, N322, N812);
xor XOR2 (N1270, N1266, N672);
xor XOR2 (N1271, N1263, N690);
nor NOR4 (N1272, N1270, N1205, N141, N494);
xor XOR2 (N1273, N1271, N163);
buf BUF1 (N1274, N1264);
nand NAND3 (N1275, N1267, N478, N916);
xor XOR2 (N1276, N1254, N140);
xor XOR2 (N1277, N1258, N1016);
and AND2 (N1278, N1272, N348);
or OR2 (N1279, N1277, N603);
nand NAND4 (N1280, N1242, N103, N833, N481);
or OR3 (N1281, N1265, N1027, N314);
and AND4 (N1282, N1279, N775, N1028, N637);
and AND3 (N1283, N1281, N564, N833);
buf BUF1 (N1284, N1278);
and AND4 (N1285, N1283, N627, N343, N621);
or OR4 (N1286, N1274, N488, N892, N1025);
nand NAND4 (N1287, N1273, N928, N885, N1231);
nor NOR4 (N1288, N1268, N277, N511, N1265);
nor NOR2 (N1289, N1269, N893);
not NOT1 (N1290, N1288);
xor XOR2 (N1291, N1276, N1138);
not NOT1 (N1292, N1284);
or OR2 (N1293, N1289, N790);
and AND3 (N1294, N1282, N1050, N440);
and AND3 (N1295, N1292, N439, N1286);
and AND3 (N1296, N618, N36, N865);
buf BUF1 (N1297, N1290);
xor XOR2 (N1298, N1275, N1015);
xor XOR2 (N1299, N1294, N1140);
buf BUF1 (N1300, N1291);
nor NOR4 (N1301, N1296, N83, N1112, N1167);
nor NOR3 (N1302, N1280, N135, N259);
nand NAND4 (N1303, N1302, N421, N437, N722);
buf BUF1 (N1304, N1295);
not NOT1 (N1305, N1297);
xor XOR2 (N1306, N1304, N167);
and AND2 (N1307, N1299, N577);
and AND2 (N1308, N1303, N681);
or OR2 (N1309, N1306, N484);
nand NAND4 (N1310, N1307, N996, N688, N309);
not NOT1 (N1311, N1308);
nor NOR3 (N1312, N1305, N414, N222);
buf BUF1 (N1313, N1309);
nor NOR4 (N1314, N1301, N101, N377, N1071);
not NOT1 (N1315, N1314);
and AND2 (N1316, N1285, N1289);
buf BUF1 (N1317, N1298);
and AND3 (N1318, N1315, N1286, N466);
xor XOR2 (N1319, N1313, N1008);
nor NOR2 (N1320, N1318, N978);
and AND4 (N1321, N1310, N1081, N708, N925);
not NOT1 (N1322, N1287);
nor NOR4 (N1323, N1317, N581, N472, N1304);
or OR2 (N1324, N1320, N44);
or OR3 (N1325, N1322, N998, N733);
or OR4 (N1326, N1323, N506, N394, N1147);
or OR3 (N1327, N1311, N1130, N621);
not NOT1 (N1328, N1321);
not NOT1 (N1329, N1327);
and AND2 (N1330, N1326, N510);
nand NAND2 (N1331, N1324, N439);
nand NAND3 (N1332, N1329, N647, N1016);
buf BUF1 (N1333, N1312);
nand NAND2 (N1334, N1328, N141);
buf BUF1 (N1335, N1330);
or OR2 (N1336, N1319, N53);
buf BUF1 (N1337, N1336);
not NOT1 (N1338, N1316);
and AND4 (N1339, N1333, N261, N1300, N963);
xor XOR2 (N1340, N241, N393);
buf BUF1 (N1341, N1293);
buf BUF1 (N1342, N1334);
or OR3 (N1343, N1331, N492, N11);
nor NOR2 (N1344, N1335, N34);
xor XOR2 (N1345, N1342, N394);
nor NOR4 (N1346, N1345, N384, N321, N397);
xor XOR2 (N1347, N1346, N1235);
buf BUF1 (N1348, N1338);
and AND3 (N1349, N1325, N857, N1142);
and AND3 (N1350, N1349, N562, N1297);
buf BUF1 (N1351, N1332);
or OR2 (N1352, N1339, N675);
or OR2 (N1353, N1350, N1195);
not NOT1 (N1354, N1351);
buf BUF1 (N1355, N1341);
not NOT1 (N1356, N1355);
xor XOR2 (N1357, N1354, N1317);
or OR3 (N1358, N1337, N245, N1179);
nor NOR4 (N1359, N1353, N743, N235, N172);
not NOT1 (N1360, N1357);
not NOT1 (N1361, N1356);
nand NAND4 (N1362, N1360, N305, N507, N866);
xor XOR2 (N1363, N1359, N1013);
xor XOR2 (N1364, N1361, N51);
buf BUF1 (N1365, N1363);
nand NAND4 (N1366, N1340, N838, N431, N1317);
and AND3 (N1367, N1364, N947, N62);
buf BUF1 (N1368, N1358);
not NOT1 (N1369, N1368);
or OR3 (N1370, N1348, N15, N148);
or OR4 (N1371, N1362, N201, N873, N538);
nor NOR2 (N1372, N1370, N581);
nor NOR4 (N1373, N1365, N472, N629, N1156);
nand NAND3 (N1374, N1372, N309, N1351);
or OR2 (N1375, N1347, N1312);
xor XOR2 (N1376, N1343, N555);
xor XOR2 (N1377, N1366, N1091);
not NOT1 (N1378, N1367);
nor NOR2 (N1379, N1371, N241);
not NOT1 (N1380, N1369);
or OR3 (N1381, N1380, N1007, N890);
xor XOR2 (N1382, N1378, N220);
or OR2 (N1383, N1374, N1316);
xor XOR2 (N1384, N1379, N1294);
not NOT1 (N1385, N1384);
buf BUF1 (N1386, N1344);
or OR2 (N1387, N1383, N299);
buf BUF1 (N1388, N1376);
or OR3 (N1389, N1381, N366, N1243);
or OR4 (N1390, N1389, N1146, N1021, N1279);
nor NOR4 (N1391, N1388, N213, N1112, N1184);
nand NAND3 (N1392, N1377, N394, N1239);
nor NOR3 (N1393, N1386, N1078, N715);
not NOT1 (N1394, N1391);
buf BUF1 (N1395, N1394);
nor NOR4 (N1396, N1385, N509, N153, N639);
xor XOR2 (N1397, N1352, N1209);
nor NOR4 (N1398, N1373, N75, N269, N448);
nor NOR2 (N1399, N1398, N933);
or OR2 (N1400, N1390, N757);
buf BUF1 (N1401, N1397);
or OR4 (N1402, N1392, N650, N1217, N956);
nor NOR2 (N1403, N1382, N695);
xor XOR2 (N1404, N1403, N89);
and AND2 (N1405, N1387, N608);
nand NAND2 (N1406, N1400, N597);
nor NOR3 (N1407, N1405, N1104, N283);
nand NAND3 (N1408, N1396, N1267, N42);
nor NOR2 (N1409, N1402, N427);
or OR3 (N1410, N1395, N1354, N1306);
not NOT1 (N1411, N1399);
or OR4 (N1412, N1410, N631, N195, N752);
buf BUF1 (N1413, N1408);
and AND2 (N1414, N1413, N1142);
and AND2 (N1415, N1412, N702);
xor XOR2 (N1416, N1411, N420);
or OR3 (N1417, N1406, N58, N163);
nor NOR3 (N1418, N1375, N975, N183);
nor NOR4 (N1419, N1404, N273, N1128, N1095);
or OR4 (N1420, N1407, N85, N1291, N1338);
and AND3 (N1421, N1420, N330, N761);
and AND3 (N1422, N1416, N1158, N828);
or OR4 (N1423, N1419, N754, N59, N1048);
buf BUF1 (N1424, N1417);
not NOT1 (N1425, N1393);
or OR4 (N1426, N1418, N904, N65, N1398);
nand NAND2 (N1427, N1424, N567);
buf BUF1 (N1428, N1409);
not NOT1 (N1429, N1422);
and AND3 (N1430, N1429, N593, N319);
nand NAND4 (N1431, N1426, N1140, N457, N946);
nand NAND3 (N1432, N1421, N1415, N1350);
nand NAND3 (N1433, N1346, N611, N212);
nand NAND3 (N1434, N1428, N872, N1378);
or OR3 (N1435, N1401, N937, N1047);
nor NOR4 (N1436, N1435, N777, N393, N182);
nor NOR3 (N1437, N1414, N1208, N948);
xor XOR2 (N1438, N1427, N614);
xor XOR2 (N1439, N1423, N297);
and AND4 (N1440, N1438, N62, N325, N907);
nor NOR4 (N1441, N1432, N701, N287, N931);
nand NAND4 (N1442, N1434, N1070, N1171, N769);
nand NAND4 (N1443, N1430, N1108, N759, N421);
or OR2 (N1444, N1431, N644);
or OR4 (N1445, N1425, N149, N354, N433);
buf BUF1 (N1446, N1441);
or OR4 (N1447, N1445, N343, N130, N737);
nand NAND4 (N1448, N1442, N636, N28, N528);
nand NAND2 (N1449, N1448, N518);
nor NOR3 (N1450, N1437, N1170, N1331);
nand NAND3 (N1451, N1449, N1077, N111);
not NOT1 (N1452, N1433);
buf BUF1 (N1453, N1446);
nand NAND4 (N1454, N1443, N1080, N1044, N1302);
or OR3 (N1455, N1436, N526, N123);
nand NAND3 (N1456, N1451, N905, N913);
and AND2 (N1457, N1452, N799);
and AND4 (N1458, N1444, N444, N279, N41);
buf BUF1 (N1459, N1458);
nor NOR4 (N1460, N1455, N1128, N1126, N1128);
nor NOR3 (N1461, N1450, N772, N725);
or OR3 (N1462, N1457, N1139, N974);
or OR2 (N1463, N1440, N110);
not NOT1 (N1464, N1461);
and AND3 (N1465, N1447, N508, N31);
nor NOR3 (N1466, N1453, N627, N39);
nor NOR2 (N1467, N1462, N1441);
not NOT1 (N1468, N1454);
nor NOR3 (N1469, N1439, N677, N1031);
nor NOR4 (N1470, N1469, N758, N347, N508);
nor NOR4 (N1471, N1456, N839, N1062, N506);
nand NAND2 (N1472, N1468, N914);
or OR4 (N1473, N1472, N207, N219, N1336);
or OR4 (N1474, N1467, N1246, N825, N466);
xor XOR2 (N1475, N1474, N778);
and AND2 (N1476, N1473, N1405);
or OR4 (N1477, N1465, N674, N230, N632);
and AND4 (N1478, N1471, N391, N1328, N706);
xor XOR2 (N1479, N1464, N983);
nand NAND2 (N1480, N1475, N84);
not NOT1 (N1481, N1480);
xor XOR2 (N1482, N1477, N1126);
or OR4 (N1483, N1460, N455, N725, N1425);
xor XOR2 (N1484, N1466, N1073);
buf BUF1 (N1485, N1479);
xor XOR2 (N1486, N1482, N874);
xor XOR2 (N1487, N1485, N646);
buf BUF1 (N1488, N1476);
and AND4 (N1489, N1484, N493, N109, N1403);
buf BUF1 (N1490, N1463);
nor NOR4 (N1491, N1488, N918, N12, N287);
or OR4 (N1492, N1487, N666, N1202, N781);
buf BUF1 (N1493, N1490);
buf BUF1 (N1494, N1483);
buf BUF1 (N1495, N1489);
and AND3 (N1496, N1459, N825, N5);
xor XOR2 (N1497, N1496, N733);
and AND2 (N1498, N1470, N85);
and AND2 (N1499, N1481, N1051);
or OR2 (N1500, N1493, N1165);
or OR2 (N1501, N1495, N368);
not NOT1 (N1502, N1491);
and AND4 (N1503, N1478, N542, N701, N1184);
nand NAND4 (N1504, N1501, N847, N35, N670);
xor XOR2 (N1505, N1503, N1429);
and AND3 (N1506, N1500, N827, N1157);
or OR3 (N1507, N1505, N472, N1379);
not NOT1 (N1508, N1486);
buf BUF1 (N1509, N1499);
xor XOR2 (N1510, N1506, N532);
not NOT1 (N1511, N1494);
nand NAND2 (N1512, N1502, N559);
buf BUF1 (N1513, N1511);
buf BUF1 (N1514, N1509);
or OR3 (N1515, N1497, N1411, N1063);
nand NAND4 (N1516, N1514, N790, N357, N1181);
buf BUF1 (N1517, N1516);
nor NOR4 (N1518, N1513, N775, N1385, N421);
and AND4 (N1519, N1492, N182, N1407, N903);
or OR2 (N1520, N1518, N416);
xor XOR2 (N1521, N1507, N82);
buf BUF1 (N1522, N1517);
and AND4 (N1523, N1521, N980, N586, N792);
or OR3 (N1524, N1510, N441, N654);
or OR3 (N1525, N1523, N1335, N508);
xor XOR2 (N1526, N1508, N1137);
xor XOR2 (N1527, N1525, N918);
xor XOR2 (N1528, N1504, N686);
nor NOR4 (N1529, N1520, N690, N417, N1003);
xor XOR2 (N1530, N1527, N1140);
and AND4 (N1531, N1528, N40, N1189, N778);
and AND3 (N1532, N1512, N1238, N345);
nand NAND3 (N1533, N1532, N1132, N431);
nor NOR3 (N1534, N1519, N719, N1156);
nor NOR3 (N1535, N1534, N482, N263);
not NOT1 (N1536, N1522);
nor NOR3 (N1537, N1531, N1415, N397);
xor XOR2 (N1538, N1530, N1204);
or OR2 (N1539, N1529, N920);
nand NAND4 (N1540, N1539, N474, N926, N1529);
buf BUF1 (N1541, N1524);
nand NAND2 (N1542, N1541, N266);
not NOT1 (N1543, N1540);
not NOT1 (N1544, N1537);
nand NAND3 (N1545, N1526, N702, N306);
nor NOR3 (N1546, N1536, N1017, N1340);
nor NOR4 (N1547, N1535, N721, N1054, N158);
and AND4 (N1548, N1498, N1466, N281, N1125);
nand NAND4 (N1549, N1546, N1055, N937, N1119);
nor NOR4 (N1550, N1548, N1429, N524, N1227);
not NOT1 (N1551, N1550);
not NOT1 (N1552, N1538);
or OR3 (N1553, N1549, N1171, N77);
nor NOR2 (N1554, N1547, N321);
nand NAND2 (N1555, N1551, N783);
not NOT1 (N1556, N1544);
not NOT1 (N1557, N1555);
nor NOR2 (N1558, N1552, N174);
not NOT1 (N1559, N1542);
not NOT1 (N1560, N1545);
or OR2 (N1561, N1533, N368);
nand NAND3 (N1562, N1543, N711, N1546);
nand NAND2 (N1563, N1556, N990);
buf BUF1 (N1564, N1557);
nand NAND2 (N1565, N1554, N1004);
xor XOR2 (N1566, N1563, N1501);
buf BUF1 (N1567, N1561);
not NOT1 (N1568, N1565);
buf BUF1 (N1569, N1558);
not NOT1 (N1570, N1562);
and AND3 (N1571, N1568, N380, N344);
or OR2 (N1572, N1566, N730);
xor XOR2 (N1573, N1559, N1199);
buf BUF1 (N1574, N1572);
nor NOR4 (N1575, N1564, N223, N671, N685);
and AND4 (N1576, N1574, N203, N1096, N211);
xor XOR2 (N1577, N1567, N219);
xor XOR2 (N1578, N1576, N174);
nor NOR3 (N1579, N1571, N417, N311);
and AND3 (N1580, N1560, N119, N1050);
not NOT1 (N1581, N1553);
xor XOR2 (N1582, N1570, N1392);
nand NAND2 (N1583, N1582, N421);
nand NAND3 (N1584, N1580, N1392, N1092);
nand NAND3 (N1585, N1581, N31, N527);
not NOT1 (N1586, N1575);
and AND2 (N1587, N1583, N516);
xor XOR2 (N1588, N1587, N804);
nor NOR4 (N1589, N1586, N1358, N19, N572);
nor NOR3 (N1590, N1589, N783, N1318);
xor XOR2 (N1591, N1569, N1089);
nor NOR2 (N1592, N1585, N200);
or OR3 (N1593, N1588, N688, N398);
not NOT1 (N1594, N1590);
buf BUF1 (N1595, N1594);
xor XOR2 (N1596, N1592, N1494);
nand NAND4 (N1597, N1593, N947, N1524, N1101);
buf BUF1 (N1598, N1579);
nor NOR4 (N1599, N1573, N683, N1362, N769);
or OR4 (N1600, N1599, N1159, N725, N501);
not NOT1 (N1601, N1597);
xor XOR2 (N1602, N1601, N121);
buf BUF1 (N1603, N1515);
buf BUF1 (N1604, N1603);
and AND4 (N1605, N1591, N818, N1167, N1417);
nand NAND2 (N1606, N1602, N192);
nand NAND3 (N1607, N1600, N942, N116);
buf BUF1 (N1608, N1606);
or OR3 (N1609, N1578, N455, N1090);
not NOT1 (N1610, N1577);
not NOT1 (N1611, N1609);
nand NAND3 (N1612, N1607, N491, N764);
nor NOR3 (N1613, N1584, N471, N631);
xor XOR2 (N1614, N1596, N666);
nand NAND4 (N1615, N1604, N45, N1254, N460);
nor NOR2 (N1616, N1605, N135);
buf BUF1 (N1617, N1613);
not NOT1 (N1618, N1608);
and AND4 (N1619, N1612, N958, N1343, N323);
nor NOR3 (N1620, N1617, N1553, N86);
xor XOR2 (N1621, N1618, N906);
not NOT1 (N1622, N1598);
nand NAND3 (N1623, N1615, N508, N193);
not NOT1 (N1624, N1611);
or OR2 (N1625, N1595, N708);
not NOT1 (N1626, N1621);
nor NOR4 (N1627, N1614, N72, N536, N1167);
not NOT1 (N1628, N1627);
not NOT1 (N1629, N1625);
buf BUF1 (N1630, N1628);
xor XOR2 (N1631, N1626, N1496);
or OR4 (N1632, N1610, N1234, N1196, N1431);
buf BUF1 (N1633, N1630);
and AND2 (N1634, N1623, N1427);
nand NAND4 (N1635, N1634, N456, N1013, N1094);
or OR2 (N1636, N1619, N840);
and AND2 (N1637, N1629, N919);
xor XOR2 (N1638, N1624, N498);
xor XOR2 (N1639, N1631, N621);
not NOT1 (N1640, N1620);
and AND3 (N1641, N1639, N71, N331);
and AND2 (N1642, N1633, N1484);
nand NAND3 (N1643, N1641, N463, N221);
nand NAND3 (N1644, N1640, N147, N264);
or OR3 (N1645, N1636, N775, N1491);
xor XOR2 (N1646, N1638, N792);
or OR4 (N1647, N1637, N934, N1371, N37);
nor NOR3 (N1648, N1645, N292, N1070);
and AND2 (N1649, N1648, N193);
nand NAND2 (N1650, N1622, N364);
xor XOR2 (N1651, N1650, N419);
not NOT1 (N1652, N1643);
not NOT1 (N1653, N1616);
or OR4 (N1654, N1642, N798, N1187, N634);
and AND3 (N1655, N1654, N326, N19);
xor XOR2 (N1656, N1635, N788);
buf BUF1 (N1657, N1649);
and AND4 (N1658, N1646, N427, N1276, N1525);
xor XOR2 (N1659, N1653, N1490);
and AND2 (N1660, N1658, N427);
or OR2 (N1661, N1660, N1289);
nor NOR3 (N1662, N1659, N1624, N646);
nand NAND4 (N1663, N1655, N101, N993, N1204);
nand NAND4 (N1664, N1656, N894, N1265, N548);
and AND3 (N1665, N1663, N587, N1132);
xor XOR2 (N1666, N1644, N1111);
nor NOR4 (N1667, N1651, N975, N1168, N1637);
xor XOR2 (N1668, N1666, N1434);
or OR4 (N1669, N1632, N1634, N1234, N14);
not NOT1 (N1670, N1669);
nand NAND4 (N1671, N1657, N966, N52, N1494);
xor XOR2 (N1672, N1664, N953);
buf BUF1 (N1673, N1671);
or OR3 (N1674, N1661, N42, N747);
xor XOR2 (N1675, N1673, N828);
buf BUF1 (N1676, N1652);
nand NAND4 (N1677, N1662, N355, N1054, N925);
or OR4 (N1678, N1677, N1259, N442, N1341);
not NOT1 (N1679, N1647);
nor NOR2 (N1680, N1676, N483);
buf BUF1 (N1681, N1670);
and AND2 (N1682, N1680, N777);
not NOT1 (N1683, N1681);
and AND2 (N1684, N1674, N1227);
xor XOR2 (N1685, N1665, N1127);
xor XOR2 (N1686, N1682, N556);
buf BUF1 (N1687, N1678);
not NOT1 (N1688, N1687);
or OR3 (N1689, N1672, N1422, N1684);
xor XOR2 (N1690, N1208, N1175);
or OR4 (N1691, N1690, N1646, N1502, N361);
nand NAND4 (N1692, N1668, N1104, N919, N1165);
nor NOR4 (N1693, N1689, N669, N779, N891);
nand NAND4 (N1694, N1686, N1656, N1640, N102);
and AND2 (N1695, N1693, N245);
and AND3 (N1696, N1679, N86, N456);
not NOT1 (N1697, N1688);
xor XOR2 (N1698, N1691, N94);
not NOT1 (N1699, N1685);
or OR2 (N1700, N1698, N86);
nand NAND2 (N1701, N1700, N1700);
not NOT1 (N1702, N1695);
or OR3 (N1703, N1697, N1424, N327);
or OR2 (N1704, N1699, N68);
or OR2 (N1705, N1675, N387);
and AND3 (N1706, N1704, N978, N829);
nand NAND4 (N1707, N1696, N1679, N1220, N304);
not NOT1 (N1708, N1692);
not NOT1 (N1709, N1683);
not NOT1 (N1710, N1702);
nand NAND2 (N1711, N1667, N749);
nor NOR2 (N1712, N1694, N1175);
nor NOR2 (N1713, N1710, N444);
or OR3 (N1714, N1703, N615, N51);
not NOT1 (N1715, N1714);
nor NOR3 (N1716, N1705, N541, N19);
not NOT1 (N1717, N1715);
not NOT1 (N1718, N1709);
or OR2 (N1719, N1708, N1654);
or OR4 (N1720, N1707, N891, N110, N1281);
and AND2 (N1721, N1717, N751);
or OR3 (N1722, N1720, N1216, N1662);
xor XOR2 (N1723, N1721, N1411);
and AND4 (N1724, N1713, N1404, N344, N714);
nand NAND4 (N1725, N1716, N1623, N1139, N272);
and AND2 (N1726, N1718, N1359);
and AND3 (N1727, N1725, N810, N1238);
not NOT1 (N1728, N1723);
and AND2 (N1729, N1726, N1704);
xor XOR2 (N1730, N1724, N1054);
not NOT1 (N1731, N1729);
xor XOR2 (N1732, N1731, N854);
nand NAND2 (N1733, N1719, N426);
buf BUF1 (N1734, N1727);
not NOT1 (N1735, N1712);
xor XOR2 (N1736, N1711, N578);
xor XOR2 (N1737, N1735, N1566);
xor XOR2 (N1738, N1737, N607);
buf BUF1 (N1739, N1734);
nor NOR4 (N1740, N1730, N1339, N482, N961);
or OR3 (N1741, N1722, N338, N552);
buf BUF1 (N1742, N1738);
buf BUF1 (N1743, N1706);
buf BUF1 (N1744, N1701);
and AND3 (N1745, N1742, N192, N298);
nand NAND3 (N1746, N1728, N240, N582);
buf BUF1 (N1747, N1736);
nor NOR2 (N1748, N1744, N137);
nand NAND3 (N1749, N1747, N1301, N393);
xor XOR2 (N1750, N1741, N1190);
and AND4 (N1751, N1750, N1720, N91, N1588);
or OR4 (N1752, N1748, N452, N745, N114);
nor NOR2 (N1753, N1740, N1188);
nor NOR4 (N1754, N1749, N1472, N231, N1383);
nand NAND2 (N1755, N1754, N757);
or OR4 (N1756, N1732, N963, N980, N487);
buf BUF1 (N1757, N1755);
and AND3 (N1758, N1733, N768, N402);
not NOT1 (N1759, N1757);
or OR3 (N1760, N1753, N1626, N1587);
nor NOR2 (N1761, N1739, N1198);
xor XOR2 (N1762, N1759, N1615);
and AND2 (N1763, N1746, N429);
nand NAND4 (N1764, N1743, N913, N13, N412);
or OR4 (N1765, N1751, N1215, N228, N118);
not NOT1 (N1766, N1752);
nand NAND4 (N1767, N1760, N1430, N235, N723);
or OR4 (N1768, N1758, N1617, N525, N556);
nor NOR3 (N1769, N1762, N945, N1304);
or OR4 (N1770, N1745, N154, N1582, N908);
nand NAND4 (N1771, N1769, N1315, N1351, N127);
and AND2 (N1772, N1761, N886);
not NOT1 (N1773, N1764);
nand NAND2 (N1774, N1773, N335);
nor NOR4 (N1775, N1756, N96, N1693, N585);
or OR3 (N1776, N1767, N1263, N1273);
or OR3 (N1777, N1776, N1066, N918);
xor XOR2 (N1778, N1775, N1489);
or OR3 (N1779, N1766, N1087, N1261);
not NOT1 (N1780, N1774);
nor NOR4 (N1781, N1779, N54, N1273, N986);
and AND4 (N1782, N1765, N1653, N943, N1090);
and AND3 (N1783, N1763, N1593, N1470);
nor NOR3 (N1784, N1778, N26, N178);
buf BUF1 (N1785, N1772);
or OR2 (N1786, N1784, N284);
not NOT1 (N1787, N1783);
and AND2 (N1788, N1777, N911);
nor NOR4 (N1789, N1771, N1182, N814, N1550);
nor NOR3 (N1790, N1770, N1147, N574);
nand NAND3 (N1791, N1787, N153, N1235);
nand NAND2 (N1792, N1790, N1620);
or OR3 (N1793, N1780, N164, N32);
buf BUF1 (N1794, N1788);
nor NOR4 (N1795, N1768, N326, N227, N1461);
nor NOR2 (N1796, N1785, N1723);
or OR4 (N1797, N1792, N32, N1437, N93);
buf BUF1 (N1798, N1794);
buf BUF1 (N1799, N1782);
buf BUF1 (N1800, N1797);
nor NOR3 (N1801, N1795, N296, N1540);
not NOT1 (N1802, N1791);
and AND4 (N1803, N1801, N1164, N1365, N1241);
or OR4 (N1804, N1781, N631, N1000, N1741);
and AND2 (N1805, N1800, N1233);
and AND2 (N1806, N1789, N1289);
nor NOR4 (N1807, N1806, N1502, N1706, N240);
and AND2 (N1808, N1796, N913);
and AND2 (N1809, N1793, N414);
nand NAND2 (N1810, N1799, N1588);
not NOT1 (N1811, N1808);
nor NOR3 (N1812, N1786, N1672, N26);
and AND2 (N1813, N1811, N653);
or OR3 (N1814, N1812, N1262, N1135);
not NOT1 (N1815, N1805);
xor XOR2 (N1816, N1813, N1118);
and AND4 (N1817, N1803, N271, N113, N895);
nor NOR4 (N1818, N1798, N274, N955, N50);
not NOT1 (N1819, N1804);
and AND3 (N1820, N1818, N275, N274);
nor NOR2 (N1821, N1807, N1820);
not NOT1 (N1822, N1628);
or OR4 (N1823, N1822, N283, N1144, N671);
or OR3 (N1824, N1802, N548, N977);
nand NAND3 (N1825, N1809, N1394, N1255);
nor NOR3 (N1826, N1815, N388, N1050);
nand NAND3 (N1827, N1819, N110, N1189);
nand NAND2 (N1828, N1817, N1646);
not NOT1 (N1829, N1826);
buf BUF1 (N1830, N1824);
buf BUF1 (N1831, N1829);
and AND3 (N1832, N1814, N276, N258);
or OR4 (N1833, N1825, N1618, N892, N979);
nor NOR3 (N1834, N1830, N1351, N164);
nand NAND4 (N1835, N1831, N653, N390, N440);
xor XOR2 (N1836, N1810, N909);
or OR2 (N1837, N1821, N625);
nand NAND2 (N1838, N1828, N369);
nand NAND2 (N1839, N1835, N1049);
nor NOR3 (N1840, N1832, N438, N1178);
xor XOR2 (N1841, N1833, N833);
or OR2 (N1842, N1839, N1667);
buf BUF1 (N1843, N1816);
nor NOR2 (N1844, N1823, N1219);
or OR3 (N1845, N1843, N1279, N1234);
or OR3 (N1846, N1827, N1358, N806);
buf BUF1 (N1847, N1840);
nor NOR3 (N1848, N1847, N1657, N1560);
and AND3 (N1849, N1834, N1738, N37);
not NOT1 (N1850, N1836);
nor NOR4 (N1851, N1838, N1719, N368, N1206);
or OR2 (N1852, N1846, N1005);
xor XOR2 (N1853, N1848, N1687);
and AND2 (N1854, N1853, N494);
or OR2 (N1855, N1844, N1494);
nand NAND2 (N1856, N1837, N1248);
nand NAND4 (N1857, N1849, N1747, N723, N1366);
and AND3 (N1858, N1852, N708, N127);
buf BUF1 (N1859, N1858);
nand NAND4 (N1860, N1856, N1091, N1748, N199);
and AND4 (N1861, N1851, N1735, N1308, N546);
nor NOR4 (N1862, N1860, N342, N1781, N959);
and AND3 (N1863, N1862, N534, N82);
or OR2 (N1864, N1841, N311);
not NOT1 (N1865, N1855);
nand NAND3 (N1866, N1857, N1423, N469);
xor XOR2 (N1867, N1859, N1217);
and AND2 (N1868, N1842, N902);
buf BUF1 (N1869, N1865);
or OR4 (N1870, N1861, N1124, N152, N407);
and AND3 (N1871, N1850, N1837, N877);
buf BUF1 (N1872, N1866);
buf BUF1 (N1873, N1845);
not NOT1 (N1874, N1863);
not NOT1 (N1875, N1873);
buf BUF1 (N1876, N1874);
buf BUF1 (N1877, N1871);
buf BUF1 (N1878, N1869);
buf BUF1 (N1879, N1867);
not NOT1 (N1880, N1870);
xor XOR2 (N1881, N1879, N184);
xor XOR2 (N1882, N1877, N1716);
nor NOR2 (N1883, N1868, N727);
not NOT1 (N1884, N1854);
nand NAND3 (N1885, N1876, N347, N965);
nor NOR4 (N1886, N1881, N412, N569, N1120);
and AND3 (N1887, N1864, N391, N1842);
buf BUF1 (N1888, N1875);
or OR2 (N1889, N1884, N742);
not NOT1 (N1890, N1880);
buf BUF1 (N1891, N1889);
or OR4 (N1892, N1882, N583, N372, N1745);
and AND3 (N1893, N1883, N727, N1065);
and AND3 (N1894, N1885, N1833, N14);
nor NOR2 (N1895, N1891, N1437);
buf BUF1 (N1896, N1895);
and AND2 (N1897, N1893, N860);
and AND4 (N1898, N1872, N102, N195, N429);
nor NOR2 (N1899, N1887, N1740);
buf BUF1 (N1900, N1894);
nor NOR2 (N1901, N1899, N663);
and AND2 (N1902, N1898, N676);
or OR3 (N1903, N1896, N1148, N845);
not NOT1 (N1904, N1886);
buf BUF1 (N1905, N1904);
and AND2 (N1906, N1905, N1094);
nor NOR4 (N1907, N1890, N731, N1375, N449);
nor NOR2 (N1908, N1903, N1632);
or OR2 (N1909, N1878, N31);
nor NOR3 (N1910, N1909, N326, N1056);
not NOT1 (N1911, N1910);
nand NAND3 (N1912, N1911, N246, N211);
and AND3 (N1913, N1897, N949, N1440);
xor XOR2 (N1914, N1908, N889);
and AND3 (N1915, N1914, N727, N1093);
xor XOR2 (N1916, N1901, N1714);
buf BUF1 (N1917, N1900);
nor NOR4 (N1918, N1907, N859, N1247, N194);
nand NAND3 (N1919, N1913, N520, N1162);
nand NAND4 (N1920, N1917, N1691, N807, N1149);
or OR2 (N1921, N1920, N334);
xor XOR2 (N1922, N1888, N965);
nor NOR2 (N1923, N1892, N1689);
or OR2 (N1924, N1906, N289);
buf BUF1 (N1925, N1918);
nor NOR2 (N1926, N1924, N1200);
or OR4 (N1927, N1922, N293, N236, N449);
nor NOR2 (N1928, N1926, N1183);
not NOT1 (N1929, N1916);
not NOT1 (N1930, N1929);
and AND4 (N1931, N1919, N1512, N1632, N319);
xor XOR2 (N1932, N1902, N911);
nor NOR4 (N1933, N1930, N1383, N1143, N818);
xor XOR2 (N1934, N1915, N75);
or OR2 (N1935, N1925, N302);
nand NAND2 (N1936, N1921, N734);
and AND3 (N1937, N1923, N456, N473);
nand NAND4 (N1938, N1927, N1661, N1744, N1742);
xor XOR2 (N1939, N1928, N381);
or OR3 (N1940, N1938, N261, N1613);
or OR2 (N1941, N1939, N1024);
or OR4 (N1942, N1934, N754, N733, N1268);
nand NAND4 (N1943, N1940, N266, N1470, N1130);
not NOT1 (N1944, N1943);
not NOT1 (N1945, N1912);
and AND3 (N1946, N1935, N1853, N1371);
and AND3 (N1947, N1932, N1234, N416);
xor XOR2 (N1948, N1931, N1506);
and AND3 (N1949, N1942, N1185, N760);
and AND2 (N1950, N1937, N1267);
and AND4 (N1951, N1946, N1445, N1802, N1225);
xor XOR2 (N1952, N1933, N875);
or OR3 (N1953, N1947, N1767, N308);
nor NOR3 (N1954, N1949, N1650, N604);
buf BUF1 (N1955, N1944);
nand NAND3 (N1956, N1955, N473, N1124);
xor XOR2 (N1957, N1951, N1293);
xor XOR2 (N1958, N1954, N1293);
or OR2 (N1959, N1936, N509);
not NOT1 (N1960, N1956);
not NOT1 (N1961, N1948);
and AND3 (N1962, N1960, N1845, N1183);
not NOT1 (N1963, N1950);
not NOT1 (N1964, N1957);
nand NAND4 (N1965, N1941, N364, N516, N738);
buf BUF1 (N1966, N1952);
and AND4 (N1967, N1962, N468, N1952, N692);
nand NAND4 (N1968, N1959, N497, N647, N1612);
nand NAND2 (N1969, N1958, N1848);
or OR4 (N1970, N1967, N730, N865, N1031);
not NOT1 (N1971, N1963);
nand NAND2 (N1972, N1953, N937);
and AND2 (N1973, N1966, N189);
nor NOR4 (N1974, N1968, N38, N3, N253);
nand NAND4 (N1975, N1973, N887, N1408, N647);
not NOT1 (N1976, N1965);
nand NAND2 (N1977, N1970, N1376);
nor NOR4 (N1978, N1964, N425, N1919, N1381);
not NOT1 (N1979, N1975);
nor NOR4 (N1980, N1976, N749, N1346, N317);
xor XOR2 (N1981, N1961, N1322);
and AND4 (N1982, N1977, N1687, N1417, N124);
or OR2 (N1983, N1981, N568);
nor NOR4 (N1984, N1969, N1310, N1816, N1013);
or OR3 (N1985, N1984, N818, N1771);
buf BUF1 (N1986, N1945);
not NOT1 (N1987, N1982);
buf BUF1 (N1988, N1978);
not NOT1 (N1989, N1971);
xor XOR2 (N1990, N1989, N335);
xor XOR2 (N1991, N1988, N546);
and AND2 (N1992, N1983, N1924);
and AND2 (N1993, N1974, N1107);
not NOT1 (N1994, N1991);
buf BUF1 (N1995, N1990);
xor XOR2 (N1996, N1986, N1913);
nand NAND3 (N1997, N1979, N1433, N1859);
nand NAND3 (N1998, N1972, N156, N1697);
buf BUF1 (N1999, N1998);
xor XOR2 (N2000, N1980, N168);
not NOT1 (N2001, N1987);
and AND2 (N2002, N1995, N1763);
or OR3 (N2003, N2001, N1988, N1611);
and AND2 (N2004, N1993, N1075);
buf BUF1 (N2005, N1997);
or OR2 (N2006, N2002, N268);
xor XOR2 (N2007, N1992, N1643);
and AND2 (N2008, N2003, N494);
nand NAND2 (N2009, N1994, N892);
nor NOR4 (N2010, N1996, N1848, N1457, N58);
xor XOR2 (N2011, N2000, N967);
and AND3 (N2012, N2007, N1957, N1036);
not NOT1 (N2013, N2009);
nor NOR2 (N2014, N2010, N1605);
not NOT1 (N2015, N2011);
buf BUF1 (N2016, N1999);
xor XOR2 (N2017, N2004, N1885);
or OR4 (N2018, N2008, N734, N167, N1765);
or OR2 (N2019, N2012, N1402);
nor NOR3 (N2020, N1985, N1883, N1218);
not NOT1 (N2021, N2020);
xor XOR2 (N2022, N2021, N180);
nor NOR2 (N2023, N2022, N894);
and AND2 (N2024, N2014, N1253);
or OR2 (N2025, N2017, N1884);
or OR2 (N2026, N2018, N1373);
nand NAND4 (N2027, N2013, N403, N671, N1959);
nand NAND2 (N2028, N2006, N626);
and AND3 (N2029, N2025, N730, N162);
nor NOR2 (N2030, N2023, N122);
xor XOR2 (N2031, N2024, N1860);
not NOT1 (N2032, N2019);
buf BUF1 (N2033, N2026);
not NOT1 (N2034, N2031);
not NOT1 (N2035, N2034);
not NOT1 (N2036, N2015);
buf BUF1 (N2037, N2036);
or OR3 (N2038, N2029, N1194, N640);
not NOT1 (N2039, N2038);
xor XOR2 (N2040, N2037, N15);
buf BUF1 (N2041, N2035);
nand NAND2 (N2042, N2028, N46);
not NOT1 (N2043, N2027);
nor NOR2 (N2044, N2041, N21);
buf BUF1 (N2045, N2032);
buf BUF1 (N2046, N2016);
not NOT1 (N2047, N2040);
buf BUF1 (N2048, N2030);
or OR2 (N2049, N2033, N1920);
and AND2 (N2050, N2049, N759);
xor XOR2 (N2051, N2045, N733);
nor NOR3 (N2052, N2046, N540, N1294);
buf BUF1 (N2053, N2052);
buf BUF1 (N2054, N2039);
and AND3 (N2055, N2051, N1942, N1916);
and AND2 (N2056, N2047, N982);
xor XOR2 (N2057, N2044, N583);
buf BUF1 (N2058, N2054);
and AND2 (N2059, N2043, N299);
not NOT1 (N2060, N2055);
not NOT1 (N2061, N2058);
nor NOR2 (N2062, N2053, N137);
and AND2 (N2063, N2062, N426);
or OR3 (N2064, N2061, N666, N455);
not NOT1 (N2065, N2063);
and AND3 (N2066, N2056, N596, N1325);
not NOT1 (N2067, N2048);
not NOT1 (N2068, N2064);
nor NOR4 (N2069, N2060, N520, N1263, N1754);
not NOT1 (N2070, N2059);
and AND4 (N2071, N2066, N277, N1986, N898);
xor XOR2 (N2072, N2068, N52);
buf BUF1 (N2073, N2005);
and AND3 (N2074, N2072, N98, N1870);
and AND3 (N2075, N2057, N1241, N856);
and AND2 (N2076, N2067, N1353);
and AND3 (N2077, N2065, N830, N316);
not NOT1 (N2078, N2042);
or OR3 (N2079, N2077, N1714, N143);
and AND4 (N2080, N2050, N361, N693, N1488);
and AND3 (N2081, N2080, N22, N509);
buf BUF1 (N2082, N2076);
nor NOR3 (N2083, N2081, N1718, N1087);
or OR2 (N2084, N2082, N207);
xor XOR2 (N2085, N2069, N1196);
xor XOR2 (N2086, N2078, N814);
not NOT1 (N2087, N2085);
xor XOR2 (N2088, N2086, N129);
xor XOR2 (N2089, N2083, N1131);
nor NOR2 (N2090, N2089, N1771);
nand NAND3 (N2091, N2079, N193, N1452);
not NOT1 (N2092, N2087);
nor NOR2 (N2093, N2070, N1757);
xor XOR2 (N2094, N2073, N431);
nand NAND3 (N2095, N2088, N1076, N1326);
and AND4 (N2096, N2084, N1170, N309, N1401);
or OR4 (N2097, N2075, N357, N754, N179);
xor XOR2 (N2098, N2092, N1491);
and AND4 (N2099, N2098, N709, N1783, N828);
not NOT1 (N2100, N2097);
not NOT1 (N2101, N2096);
not NOT1 (N2102, N2094);
or OR3 (N2103, N2101, N770, N743);
not NOT1 (N2104, N2074);
not NOT1 (N2105, N2071);
nor NOR3 (N2106, N2090, N1894, N421);
nand NAND2 (N2107, N2093, N1460);
and AND3 (N2108, N2091, N1493, N781);
not NOT1 (N2109, N2102);
buf BUF1 (N2110, N2108);
buf BUF1 (N2111, N2103);
and AND3 (N2112, N2105, N1841, N226);
and AND3 (N2113, N2104, N680, N1103);
buf BUF1 (N2114, N2113);
buf BUF1 (N2115, N2107);
not NOT1 (N2116, N2100);
nand NAND4 (N2117, N2112, N502, N42, N1434);
nand NAND4 (N2118, N2111, N13, N1462, N658);
and AND2 (N2119, N2114, N1033);
nand NAND4 (N2120, N2116, N652, N127, N1663);
nor NOR3 (N2121, N2099, N1709, N688);
or OR3 (N2122, N2120, N1497, N1314);
or OR4 (N2123, N2121, N1962, N465, N1091);
nor NOR2 (N2124, N2119, N1756);
or OR4 (N2125, N2106, N2073, N373, N479);
and AND2 (N2126, N2124, N963);
or OR2 (N2127, N2115, N1836);
nand NAND4 (N2128, N2117, N103, N79, N1434);
not NOT1 (N2129, N2127);
and AND2 (N2130, N2126, N24);
not NOT1 (N2131, N2125);
and AND4 (N2132, N2129, N1231, N2125, N666);
not NOT1 (N2133, N2109);
xor XOR2 (N2134, N2128, N875);
or OR2 (N2135, N2132, N1580);
or OR4 (N2136, N2134, N2110, N1632, N980);
and AND3 (N2137, N234, N325, N1294);
xor XOR2 (N2138, N2137, N907);
or OR3 (N2139, N2130, N108, N1302);
not NOT1 (N2140, N2133);
xor XOR2 (N2141, N2135, N2017);
buf BUF1 (N2142, N2095);
not NOT1 (N2143, N2140);
or OR4 (N2144, N2118, N333, N1488, N2030);
not NOT1 (N2145, N2136);
buf BUF1 (N2146, N2142);
xor XOR2 (N2147, N2144, N405);
or OR2 (N2148, N2139, N568);
and AND3 (N2149, N2131, N633, N625);
xor XOR2 (N2150, N2146, N1043);
xor XOR2 (N2151, N2150, N1228);
xor XOR2 (N2152, N2147, N1514);
and AND4 (N2153, N2141, N1217, N1487, N1317);
or OR2 (N2154, N2149, N1709);
buf BUF1 (N2155, N2148);
nor NOR3 (N2156, N2155, N1130, N982);
and AND4 (N2157, N2154, N670, N1838, N909);
buf BUF1 (N2158, N2138);
buf BUF1 (N2159, N2151);
or OR4 (N2160, N2157, N122, N1177, N789);
buf BUF1 (N2161, N2156);
not NOT1 (N2162, N2159);
nor NOR3 (N2163, N2145, N504, N1946);
or OR4 (N2164, N2123, N131, N1276, N803);
not NOT1 (N2165, N2163);
nor NOR4 (N2166, N2160, N1127, N897, N406);
or OR2 (N2167, N2122, N1989);
nor NOR3 (N2168, N2166, N1328, N1993);
xor XOR2 (N2169, N2153, N544);
or OR2 (N2170, N2161, N1249);
nor NOR2 (N2171, N2158, N1472);
nor NOR3 (N2172, N2170, N711, N981);
nand NAND4 (N2173, N2165, N824, N1814, N1698);
buf BUF1 (N2174, N2171);
nor NOR2 (N2175, N2143, N835);
buf BUF1 (N2176, N2167);
not NOT1 (N2177, N2169);
and AND3 (N2178, N2174, N2010, N930);
nor NOR3 (N2179, N2172, N2172, N628);
or OR3 (N2180, N2179, N736, N200);
nor NOR3 (N2181, N2173, N1624, N1917);
and AND2 (N2182, N2177, N1836);
buf BUF1 (N2183, N2178);
and AND3 (N2184, N2152, N1628, N1285);
xor XOR2 (N2185, N2175, N1962);
buf BUF1 (N2186, N2176);
xor XOR2 (N2187, N2168, N1065);
xor XOR2 (N2188, N2162, N592);
xor XOR2 (N2189, N2188, N1805);
and AND3 (N2190, N2180, N494, N197);
and AND3 (N2191, N2189, N1336, N1948);
buf BUF1 (N2192, N2164);
nor NOR2 (N2193, N2183, N1828);
nor NOR4 (N2194, N2186, N1357, N1999, N16);
buf BUF1 (N2195, N2181);
not NOT1 (N2196, N2187);
or OR3 (N2197, N2185, N994, N944);
buf BUF1 (N2198, N2197);
and AND3 (N2199, N2193, N912, N1366);
nor NOR2 (N2200, N2198, N583);
nand NAND3 (N2201, N2190, N1732, N1548);
and AND4 (N2202, N2199, N1862, N1569, N1116);
buf BUF1 (N2203, N2192);
or OR3 (N2204, N2203, N1866, N1100);
nand NAND4 (N2205, N2196, N2185, N609, N735);
nand NAND2 (N2206, N2202, N699);
and AND3 (N2207, N2195, N1064, N1079);
nor NOR3 (N2208, N2184, N1115, N1898);
xor XOR2 (N2209, N2194, N1635);
nor NOR3 (N2210, N2201, N583, N2071);
and AND4 (N2211, N2208, N1819, N888, N830);
and AND4 (N2212, N2200, N300, N1616, N2031);
and AND2 (N2213, N2205, N1300);
nand NAND4 (N2214, N2209, N201, N1134, N85);
or OR2 (N2215, N2214, N532);
xor XOR2 (N2216, N2191, N1319);
nand NAND3 (N2217, N2206, N1363, N1310);
xor XOR2 (N2218, N2210, N749);
xor XOR2 (N2219, N2182, N1281);
nand NAND3 (N2220, N2216, N892, N492);
buf BUF1 (N2221, N2211);
and AND2 (N2222, N2218, N1759);
and AND4 (N2223, N2213, N87, N49, N796);
or OR4 (N2224, N2215, N655, N2009, N924);
nor NOR3 (N2225, N2219, N647, N1727);
and AND2 (N2226, N2207, N810);
and AND3 (N2227, N2225, N1280, N1180);
nand NAND4 (N2228, N2221, N1027, N1093, N1038);
or OR3 (N2229, N2228, N2172, N158);
not NOT1 (N2230, N2227);
and AND3 (N2231, N2224, N1329, N1125);
buf BUF1 (N2232, N2204);
nor NOR2 (N2233, N2220, N1556);
xor XOR2 (N2234, N2231, N302);
buf BUF1 (N2235, N2226);
xor XOR2 (N2236, N2232, N1220);
and AND4 (N2237, N2233, N1344, N914, N1458);
and AND2 (N2238, N2237, N1391);
or OR4 (N2239, N2223, N1689, N2176, N1809);
and AND2 (N2240, N2236, N2113);
xor XOR2 (N2241, N2217, N1742);
nand NAND3 (N2242, N2239, N1780, N1134);
and AND4 (N2243, N2229, N1990, N549, N1333);
xor XOR2 (N2244, N2234, N264);
or OR4 (N2245, N2235, N1671, N1670, N950);
buf BUF1 (N2246, N2230);
buf BUF1 (N2247, N2238);
buf BUF1 (N2248, N2242);
or OR2 (N2249, N2247, N1461);
xor XOR2 (N2250, N2244, N1888);
buf BUF1 (N2251, N2246);
nor NOR3 (N2252, N2251, N1597, N1977);
nand NAND2 (N2253, N2212, N864);
or OR3 (N2254, N2249, N53, N2125);
or OR3 (N2255, N2240, N1290, N705);
nand NAND2 (N2256, N2243, N1195);
or OR4 (N2257, N2252, N1949, N717, N407);
nor NOR2 (N2258, N2222, N1920);
nand NAND2 (N2259, N2253, N697);
and AND3 (N2260, N2258, N1940, N2128);
nor NOR4 (N2261, N2260, N1201, N1024, N554);
or OR3 (N2262, N2250, N1751, N441);
xor XOR2 (N2263, N2245, N1029);
xor XOR2 (N2264, N2256, N146);
not NOT1 (N2265, N2261);
not NOT1 (N2266, N2265);
xor XOR2 (N2267, N2263, N34);
buf BUF1 (N2268, N2255);
nor NOR3 (N2269, N2266, N1052, N858);
xor XOR2 (N2270, N2264, N1465);
not NOT1 (N2271, N2262);
not NOT1 (N2272, N2241);
xor XOR2 (N2273, N2272, N612);
or OR4 (N2274, N2269, N1883, N1154, N1257);
xor XOR2 (N2275, N2270, N2176);
and AND2 (N2276, N2275, N525);
xor XOR2 (N2277, N2257, N2187);
nor NOR2 (N2278, N2254, N1669);
nor NOR4 (N2279, N2273, N2150, N2212, N223);
xor XOR2 (N2280, N2248, N744);
nand NAND2 (N2281, N2268, N1282);
xor XOR2 (N2282, N2278, N1894);
nand NAND3 (N2283, N2274, N564, N780);
nand NAND4 (N2284, N2281, N294, N1547, N2161);
buf BUF1 (N2285, N2279);
buf BUF1 (N2286, N2282);
buf BUF1 (N2287, N2283);
and AND2 (N2288, N2276, N1394);
xor XOR2 (N2289, N2286, N1166);
nand NAND3 (N2290, N2289, N805, N1205);
not NOT1 (N2291, N2271);
buf BUF1 (N2292, N2290);
or OR4 (N2293, N2267, N2168, N638, N699);
xor XOR2 (N2294, N2277, N1692);
buf BUF1 (N2295, N2284);
not NOT1 (N2296, N2280);
not NOT1 (N2297, N2285);
nor NOR2 (N2298, N2292, N876);
and AND4 (N2299, N2287, N1839, N1874, N883);
not NOT1 (N2300, N2296);
buf BUF1 (N2301, N2300);
nand NAND3 (N2302, N2295, N1461, N2293);
nand NAND3 (N2303, N15, N223, N1480);
nand NAND4 (N2304, N2302, N556, N1142, N2301);
xor XOR2 (N2305, N1927, N865);
buf BUF1 (N2306, N2294);
or OR4 (N2307, N2297, N279, N527, N60);
nand NAND3 (N2308, N2307, N1451, N1539);
or OR4 (N2309, N2291, N1442, N1970, N697);
buf BUF1 (N2310, N2303);
nor NOR2 (N2311, N2259, N1289);
nand NAND2 (N2312, N2299, N471);
or OR3 (N2313, N2309, N1227, N1238);
not NOT1 (N2314, N2312);
and AND2 (N2315, N2313, N1033);
xor XOR2 (N2316, N2306, N1465);
nand NAND3 (N2317, N2305, N466, N1324);
nor NOR2 (N2318, N2310, N1611);
not NOT1 (N2319, N2316);
and AND3 (N2320, N2288, N2034, N211);
or OR4 (N2321, N2314, N2243, N63, N2266);
not NOT1 (N2322, N2308);
not NOT1 (N2323, N2317);
and AND2 (N2324, N2318, N1173);
buf BUF1 (N2325, N2324);
nand NAND4 (N2326, N2298, N1081, N2224, N2262);
nor NOR3 (N2327, N2304, N1776, N1338);
or OR4 (N2328, N2326, N1621, N1692, N1991);
or OR2 (N2329, N2328, N1357);
not NOT1 (N2330, N2327);
and AND2 (N2331, N2325, N1592);
xor XOR2 (N2332, N2311, N1531);
not NOT1 (N2333, N2321);
nand NAND2 (N2334, N2320, N1396);
nand NAND2 (N2335, N2333, N129);
not NOT1 (N2336, N2334);
and AND2 (N2337, N2315, N287);
nand NAND3 (N2338, N2322, N1012, N1931);
xor XOR2 (N2339, N2319, N2098);
buf BUF1 (N2340, N2332);
nor NOR3 (N2341, N2330, N1154, N151);
xor XOR2 (N2342, N2336, N1272);
nor NOR4 (N2343, N2338, N875, N803, N1883);
buf BUF1 (N2344, N2340);
buf BUF1 (N2345, N2335);
nor NOR3 (N2346, N2337, N967, N689);
buf BUF1 (N2347, N2323);
nand NAND3 (N2348, N2345, N1805, N179);
and AND2 (N2349, N2331, N1177);
and AND2 (N2350, N2346, N1665);
and AND3 (N2351, N2349, N1795, N825);
xor XOR2 (N2352, N2339, N1768);
buf BUF1 (N2353, N2341);
buf BUF1 (N2354, N2353);
xor XOR2 (N2355, N2348, N2203);
nand NAND4 (N2356, N2352, N72, N1888, N1351);
or OR4 (N2357, N2344, N54, N724, N2038);
or OR3 (N2358, N2350, N247, N1149);
buf BUF1 (N2359, N2355);
not NOT1 (N2360, N2359);
not NOT1 (N2361, N2354);
buf BUF1 (N2362, N2343);
buf BUF1 (N2363, N2361);
nor NOR4 (N2364, N2363, N1837, N517, N1289);
buf BUF1 (N2365, N2364);
xor XOR2 (N2366, N2351, N2210);
and AND4 (N2367, N2347, N1639, N1203, N1849);
buf BUF1 (N2368, N2360);
nand NAND3 (N2369, N2356, N2330, N154);
xor XOR2 (N2370, N2362, N2364);
and AND3 (N2371, N2357, N1278, N1983);
or OR3 (N2372, N2365, N1368, N622);
nor NOR2 (N2373, N2369, N1805);
xor XOR2 (N2374, N2366, N2012);
and AND2 (N2375, N2329, N1941);
nor NOR4 (N2376, N2342, N2154, N185, N699);
nand NAND2 (N2377, N2375, N1742);
and AND3 (N2378, N2373, N1270, N1899);
buf BUF1 (N2379, N2374);
and AND2 (N2380, N2368, N1314);
and AND3 (N2381, N2370, N84, N1314);
nand NAND2 (N2382, N2379, N2194);
not NOT1 (N2383, N2371);
xor XOR2 (N2384, N2377, N1451);
xor XOR2 (N2385, N2378, N388);
nor NOR3 (N2386, N2367, N2145, N1981);
xor XOR2 (N2387, N2383, N122);
xor XOR2 (N2388, N2382, N551);
nand NAND3 (N2389, N2381, N1185, N2387);
or OR3 (N2390, N1388, N1545, N872);
or OR4 (N2391, N2372, N1549, N64, N18);
and AND4 (N2392, N2389, N1809, N2017, N238);
nand NAND2 (N2393, N2390, N1324);
not NOT1 (N2394, N2391);
xor XOR2 (N2395, N2392, N1536);
nand NAND4 (N2396, N2380, N1573, N1147, N1716);
buf BUF1 (N2397, N2358);
buf BUF1 (N2398, N2376);
xor XOR2 (N2399, N2385, N1668);
not NOT1 (N2400, N2393);
not NOT1 (N2401, N2386);
nand NAND3 (N2402, N2394, N505, N236);
nor NOR3 (N2403, N2397, N5, N1099);
or OR2 (N2404, N2384, N253);
xor XOR2 (N2405, N2398, N2293);
buf BUF1 (N2406, N2400);
nor NOR3 (N2407, N2405, N1905, N1956);
nand NAND4 (N2408, N2396, N1857, N1339, N1843);
xor XOR2 (N2409, N2388, N1192);
nor NOR2 (N2410, N2401, N346);
xor XOR2 (N2411, N2406, N1094);
not NOT1 (N2412, N2399);
or OR3 (N2413, N2403, N360, N609);
nand NAND2 (N2414, N2412, N238);
nor NOR4 (N2415, N2413, N512, N1007, N2018);
xor XOR2 (N2416, N2395, N1797);
or OR4 (N2417, N2404, N441, N1037, N2212);
not NOT1 (N2418, N2417);
nor NOR3 (N2419, N2411, N385, N1049);
and AND2 (N2420, N2418, N1115);
and AND3 (N2421, N2420, N45, N2162);
nor NOR2 (N2422, N2421, N1670);
or OR2 (N2423, N2408, N1851);
nand NAND2 (N2424, N2419, N1159);
xor XOR2 (N2425, N2409, N1520);
or OR2 (N2426, N2423, N1841);
and AND3 (N2427, N2414, N1724, N1308);
nor NOR2 (N2428, N2407, N1806);
and AND2 (N2429, N2428, N1918);
xor XOR2 (N2430, N2410, N1959);
not NOT1 (N2431, N2424);
buf BUF1 (N2432, N2422);
nand NAND4 (N2433, N2430, N781, N2303, N957);
or OR3 (N2434, N2427, N2082, N355);
and AND4 (N2435, N2432, N738, N2183, N1108);
and AND2 (N2436, N2435, N878);
or OR3 (N2437, N2431, N2163, N264);
nand NAND3 (N2438, N2429, N1284, N1477);
nor NOR2 (N2439, N2425, N2287);
and AND2 (N2440, N2438, N1870);
xor XOR2 (N2441, N2436, N1580);
buf BUF1 (N2442, N2437);
not NOT1 (N2443, N2442);
buf BUF1 (N2444, N2416);
and AND4 (N2445, N2443, N11, N2296, N1845);
nand NAND3 (N2446, N2440, N1813, N413);
xor XOR2 (N2447, N2402, N1633);
and AND4 (N2448, N2444, N1822, N983, N1427);
nor NOR4 (N2449, N2434, N1621, N1085, N1797);
and AND2 (N2450, N2448, N1897);
xor XOR2 (N2451, N2441, N1474);
and AND2 (N2452, N2439, N448);
nor NOR2 (N2453, N2452, N2139);
nor NOR4 (N2454, N2450, N1976, N2178, N2284);
not NOT1 (N2455, N2447);
not NOT1 (N2456, N2426);
and AND2 (N2457, N2433, N1047);
xor XOR2 (N2458, N2449, N844);
xor XOR2 (N2459, N2457, N582);
and AND4 (N2460, N2415, N918, N2173, N10);
buf BUF1 (N2461, N2458);
nand NAND4 (N2462, N2445, N27, N937, N1330);
buf BUF1 (N2463, N2461);
xor XOR2 (N2464, N2462, N1548);
buf BUF1 (N2465, N2454);
nand NAND2 (N2466, N2464, N795);
buf BUF1 (N2467, N2460);
nand NAND2 (N2468, N2455, N1503);
nand NAND3 (N2469, N2463, N1399, N2198);
nand NAND2 (N2470, N2456, N1728);
nand NAND2 (N2471, N2466, N2217);
nor NOR3 (N2472, N2467, N1436, N78);
or OR3 (N2473, N2459, N581, N77);
not NOT1 (N2474, N2471);
buf BUF1 (N2475, N2465);
nand NAND3 (N2476, N2472, N978, N2312);
buf BUF1 (N2477, N2446);
and AND2 (N2478, N2474, N1263);
xor XOR2 (N2479, N2478, N374);
or OR3 (N2480, N2476, N2118, N318);
nand NAND4 (N2481, N2477, N2412, N1944, N1455);
or OR4 (N2482, N2475, N1210, N1579, N74);
or OR2 (N2483, N2453, N2426);
not NOT1 (N2484, N2479);
nor NOR2 (N2485, N2484, N2153);
and AND4 (N2486, N2483, N1782, N1187, N2180);
not NOT1 (N2487, N2473);
and AND2 (N2488, N2451, N2378);
not NOT1 (N2489, N2470);
nand NAND2 (N2490, N2482, N1054);
not NOT1 (N2491, N2485);
and AND3 (N2492, N2491, N1945, N122);
buf BUF1 (N2493, N2492);
and AND3 (N2494, N2468, N515, N2154);
nor NOR4 (N2495, N2486, N1328, N396, N1038);
or OR2 (N2496, N2481, N231);
or OR2 (N2497, N2488, N846);
and AND4 (N2498, N2480, N487, N992, N224);
or OR4 (N2499, N2489, N982, N327, N347);
and AND3 (N2500, N2490, N1711, N2050);
not NOT1 (N2501, N2498);
not NOT1 (N2502, N2495);
xor XOR2 (N2503, N2469, N1439);
and AND4 (N2504, N2503, N861, N496, N1024);
nand NAND4 (N2505, N2504, N2328, N1626, N142);
and AND3 (N2506, N2500, N353, N92);
buf BUF1 (N2507, N2502);
or OR4 (N2508, N2493, N1660, N196, N1034);
nor NOR2 (N2509, N2501, N349);
and AND3 (N2510, N2509, N2188, N2410);
xor XOR2 (N2511, N2496, N1318);
buf BUF1 (N2512, N2506);
not NOT1 (N2513, N2494);
nor NOR3 (N2514, N2497, N1389, N1774);
nor NOR4 (N2515, N2514, N419, N1569, N2158);
and AND4 (N2516, N2515, N1392, N1142, N2347);
and AND2 (N2517, N2507, N1562);
or OR4 (N2518, N2513, N810, N2486, N2421);
xor XOR2 (N2519, N2499, N2319);
nor NOR4 (N2520, N2505, N1821, N1304, N1139);
xor XOR2 (N2521, N2518, N2216);
and AND2 (N2522, N2510, N1063);
xor XOR2 (N2523, N2521, N2349);
buf BUF1 (N2524, N2487);
or OR2 (N2525, N2520, N2086);
and AND3 (N2526, N2524, N2254, N578);
buf BUF1 (N2527, N2516);
and AND2 (N2528, N2512, N627);
nor NOR3 (N2529, N2522, N1177, N1693);
or OR4 (N2530, N2519, N1114, N831, N802);
xor XOR2 (N2531, N2530, N2402);
or OR2 (N2532, N2511, N1349);
nand NAND3 (N2533, N2528, N838, N609);
or OR4 (N2534, N2508, N661, N697, N2240);
buf BUF1 (N2535, N2523);
buf BUF1 (N2536, N2525);
buf BUF1 (N2537, N2517);
or OR4 (N2538, N2537, N1279, N435, N261);
nand NAND3 (N2539, N2527, N1969, N1446);
and AND4 (N2540, N2538, N2093, N833, N1621);
or OR3 (N2541, N2540, N2136, N1292);
buf BUF1 (N2542, N2535);
nand NAND3 (N2543, N2533, N542, N1101);
nor NOR2 (N2544, N2543, N2516);
nor NOR2 (N2545, N2529, N276);
nand NAND4 (N2546, N2544, N761, N194, N500);
buf BUF1 (N2547, N2539);
buf BUF1 (N2548, N2546);
buf BUF1 (N2549, N2531);
xor XOR2 (N2550, N2541, N2186);
nand NAND2 (N2551, N2526, N2264);
not NOT1 (N2552, N2549);
nand NAND4 (N2553, N2532, N2141, N601, N1840);
xor XOR2 (N2554, N2542, N871);
and AND4 (N2555, N2534, N1075, N743, N2230);
nand NAND3 (N2556, N2545, N18, N599);
buf BUF1 (N2557, N2547);
or OR4 (N2558, N2536, N367, N474, N512);
not NOT1 (N2559, N2558);
or OR2 (N2560, N2551, N1438);
and AND4 (N2561, N2552, N50, N374, N994);
not NOT1 (N2562, N2553);
nand NAND4 (N2563, N2554, N784, N1352, N1241);
nor NOR3 (N2564, N2561, N735, N1565);
not NOT1 (N2565, N2555);
or OR4 (N2566, N2556, N1078, N823, N1106);
and AND3 (N2567, N2560, N524, N1412);
nand NAND2 (N2568, N2557, N648);
or OR3 (N2569, N2565, N1400, N1126);
and AND3 (N2570, N2569, N1986, N813);
or OR4 (N2571, N2564, N1835, N82, N1980);
nand NAND4 (N2572, N2568, N758, N2428, N1613);
xor XOR2 (N2573, N2548, N2309);
xor XOR2 (N2574, N2571, N1956);
not NOT1 (N2575, N2567);
not NOT1 (N2576, N2566);
xor XOR2 (N2577, N2572, N275);
not NOT1 (N2578, N2576);
buf BUF1 (N2579, N2577);
buf BUF1 (N2580, N2562);
not NOT1 (N2581, N2575);
buf BUF1 (N2582, N2574);
xor XOR2 (N2583, N2550, N456);
nor NOR3 (N2584, N2579, N1542, N2172);
nor NOR2 (N2585, N2563, N2531);
and AND3 (N2586, N2583, N1714, N1332);
nand NAND4 (N2587, N2580, N948, N549, N1824);
nor NOR2 (N2588, N2585, N1327);
and AND3 (N2589, N2570, N347, N1514);
nand NAND3 (N2590, N2582, N801, N841);
or OR2 (N2591, N2578, N1191);
nor NOR2 (N2592, N2559, N1271);
nor NOR4 (N2593, N2592, N1772, N2373, N546);
xor XOR2 (N2594, N2586, N751);
or OR4 (N2595, N2594, N2128, N1091, N419);
nand NAND4 (N2596, N2591, N2071, N936, N255);
nand NAND4 (N2597, N2584, N431, N769, N2299);
and AND3 (N2598, N2573, N1152, N1778);
nand NAND3 (N2599, N2595, N2179, N595);
nand NAND3 (N2600, N2587, N692, N1024);
nor NOR2 (N2601, N2597, N2595);
or OR4 (N2602, N2596, N2132, N491, N2036);
buf BUF1 (N2603, N2589);
not NOT1 (N2604, N2598);
or OR3 (N2605, N2602, N1517, N1742);
buf BUF1 (N2606, N2605);
xor XOR2 (N2607, N2601, N2132);
or OR2 (N2608, N2581, N1254);
nand NAND4 (N2609, N2607, N1773, N2495, N707);
and AND2 (N2610, N2599, N1979);
not NOT1 (N2611, N2590);
or OR3 (N2612, N2593, N1358, N1926);
or OR3 (N2613, N2588, N215, N2373);
or OR4 (N2614, N2613, N2122, N2250, N1104);
nor NOR2 (N2615, N2612, N153);
not NOT1 (N2616, N2614);
buf BUF1 (N2617, N2616);
xor XOR2 (N2618, N2617, N984);
or OR2 (N2619, N2608, N1098);
or OR2 (N2620, N2615, N1050);
xor XOR2 (N2621, N2603, N344);
not NOT1 (N2622, N2604);
nand NAND3 (N2623, N2619, N1520, N670);
and AND2 (N2624, N2620, N1747);
or OR2 (N2625, N2621, N1313);
or OR4 (N2626, N2609, N1996, N1430, N1959);
xor XOR2 (N2627, N2606, N1217);
nand NAND3 (N2628, N2600, N2600, N567);
not NOT1 (N2629, N2625);
not NOT1 (N2630, N2629);
and AND4 (N2631, N2618, N802, N1525, N2445);
and AND2 (N2632, N2623, N2061);
and AND2 (N2633, N2632, N800);
buf BUF1 (N2634, N2628);
nand NAND4 (N2635, N2633, N520, N384, N1358);
not NOT1 (N2636, N2626);
nand NAND3 (N2637, N2627, N1067, N736);
buf BUF1 (N2638, N2610);
nand NAND4 (N2639, N2635, N2254, N1043, N324);
nand NAND3 (N2640, N2637, N1244, N1488);
xor XOR2 (N2641, N2634, N51);
buf BUF1 (N2642, N2624);
nor NOR2 (N2643, N2630, N1818);
and AND4 (N2644, N2642, N832, N1650, N402);
or OR2 (N2645, N2641, N1423);
xor XOR2 (N2646, N2639, N251);
not NOT1 (N2647, N2611);
nand NAND3 (N2648, N2631, N1554, N127);
or OR3 (N2649, N2644, N1493, N129);
xor XOR2 (N2650, N2648, N2472);
not NOT1 (N2651, N2622);
nand NAND4 (N2652, N2640, N372, N102, N2224);
nor NOR4 (N2653, N2645, N2453, N783, N2493);
nand NAND3 (N2654, N2651, N852, N1666);
or OR2 (N2655, N2650, N139);
xor XOR2 (N2656, N2647, N1297);
xor XOR2 (N2657, N2649, N660);
buf BUF1 (N2658, N2657);
and AND3 (N2659, N2643, N1790, N2509);
or OR4 (N2660, N2653, N2631, N1331, N82);
nand NAND4 (N2661, N2646, N1645, N2314, N241);
xor XOR2 (N2662, N2660, N1343);
buf BUF1 (N2663, N2636);
or OR3 (N2664, N2654, N2234, N1533);
nor NOR4 (N2665, N2655, N830, N1623, N1881);
buf BUF1 (N2666, N2665);
buf BUF1 (N2667, N2658);
nand NAND2 (N2668, N2667, N1141);
nand NAND2 (N2669, N2663, N1633);
nand NAND3 (N2670, N2668, N1039, N1661);
or OR4 (N2671, N2662, N619, N2615, N1505);
or OR2 (N2672, N2666, N179);
buf BUF1 (N2673, N2671);
not NOT1 (N2674, N2661);
buf BUF1 (N2675, N2672);
xor XOR2 (N2676, N2674, N465);
xor XOR2 (N2677, N2676, N467);
xor XOR2 (N2678, N2656, N12);
xor XOR2 (N2679, N2669, N423);
nor NOR3 (N2680, N2670, N517, N148);
buf BUF1 (N2681, N2652);
or OR2 (N2682, N2664, N2533);
buf BUF1 (N2683, N2680);
nor NOR3 (N2684, N2678, N462, N1889);
buf BUF1 (N2685, N2682);
and AND3 (N2686, N2638, N2339, N1512);
buf BUF1 (N2687, N2659);
buf BUF1 (N2688, N2685);
xor XOR2 (N2689, N2673, N1956);
xor XOR2 (N2690, N2679, N1558);
xor XOR2 (N2691, N2689, N2102);
xor XOR2 (N2692, N2684, N1809);
nor NOR4 (N2693, N2675, N61, N393, N2168);
buf BUF1 (N2694, N2686);
xor XOR2 (N2695, N2692, N1114);
and AND4 (N2696, N2694, N1373, N494, N2381);
not NOT1 (N2697, N2687);
nor NOR3 (N2698, N2690, N2109, N2083);
nor NOR3 (N2699, N2697, N1007, N760);
xor XOR2 (N2700, N2696, N11);
not NOT1 (N2701, N2681);
nor NOR4 (N2702, N2699, N108, N919, N688);
xor XOR2 (N2703, N2701, N1465);
or OR2 (N2704, N2703, N811);
or OR4 (N2705, N2691, N1687, N427, N1728);
not NOT1 (N2706, N2695);
nand NAND2 (N2707, N2702, N2013);
or OR2 (N2708, N2707, N1919);
or OR2 (N2709, N2688, N430);
xor XOR2 (N2710, N2677, N144);
not NOT1 (N2711, N2700);
not NOT1 (N2712, N2705);
and AND4 (N2713, N2710, N1931, N696, N691);
not NOT1 (N2714, N2712);
nand NAND3 (N2715, N2693, N2089, N557);
not NOT1 (N2716, N2706);
xor XOR2 (N2717, N2714, N294);
or OR2 (N2718, N2704, N2202);
buf BUF1 (N2719, N2709);
nor NOR2 (N2720, N2717, N1628);
nor NOR3 (N2721, N2698, N425, N459);
xor XOR2 (N2722, N2715, N1260);
or OR4 (N2723, N2719, N1993, N1987, N2095);
and AND3 (N2724, N2722, N1675, N2445);
or OR2 (N2725, N2683, N1263);
nor NOR2 (N2726, N2716, N2113);
or OR4 (N2727, N2725, N996, N238, N882);
and AND3 (N2728, N2713, N2248, N2163);
nand NAND4 (N2729, N2724, N641, N1763, N550);
nor NOR3 (N2730, N2721, N2475, N1430);
not NOT1 (N2731, N2726);
not NOT1 (N2732, N2718);
xor XOR2 (N2733, N2723, N1881);
or OR4 (N2734, N2708, N598, N1710, N661);
nand NAND4 (N2735, N2733, N2251, N1607, N2522);
nor NOR2 (N2736, N2732, N884);
xor XOR2 (N2737, N2734, N2001);
buf BUF1 (N2738, N2735);
nand NAND2 (N2739, N2730, N2366);
nor NOR2 (N2740, N2731, N550);
and AND2 (N2741, N2737, N1083);
nor NOR2 (N2742, N2740, N112);
nor NOR4 (N2743, N2739, N2443, N648, N1006);
buf BUF1 (N2744, N2742);
buf BUF1 (N2745, N2729);
and AND2 (N2746, N2736, N1635);
or OR4 (N2747, N2744, N1271, N1541, N69);
buf BUF1 (N2748, N2720);
xor XOR2 (N2749, N2743, N2168);
buf BUF1 (N2750, N2745);
buf BUF1 (N2751, N2741);
nor NOR4 (N2752, N2711, N2676, N2310, N1085);
xor XOR2 (N2753, N2738, N143);
buf BUF1 (N2754, N2747);
and AND4 (N2755, N2751, N1126, N1765, N194);
xor XOR2 (N2756, N2746, N458);
not NOT1 (N2757, N2750);
or OR3 (N2758, N2756, N2102, N905);
xor XOR2 (N2759, N2749, N2530);
buf BUF1 (N2760, N2754);
not NOT1 (N2761, N2759);
or OR2 (N2762, N2748, N317);
not NOT1 (N2763, N2752);
nor NOR4 (N2764, N2753, N2131, N224, N113);
buf BUF1 (N2765, N2728);
or OR4 (N2766, N2762, N552, N1476, N1490);
and AND3 (N2767, N2764, N28, N2004);
xor XOR2 (N2768, N2766, N774);
not NOT1 (N2769, N2765);
buf BUF1 (N2770, N2768);
and AND3 (N2771, N2767, N1142, N565);
nor NOR2 (N2772, N2727, N2291);
nor NOR4 (N2773, N2769, N1562, N699, N161);
nor NOR2 (N2774, N2772, N1275);
and AND2 (N2775, N2760, N2489);
nor NOR3 (N2776, N2771, N1737, N516);
nor NOR2 (N2777, N2758, N493);
or OR3 (N2778, N2774, N2490, N1253);
or OR2 (N2779, N2777, N907);
xor XOR2 (N2780, N2763, N1839);
and AND3 (N2781, N2775, N636, N2230);
or OR2 (N2782, N2780, N2738);
nor NOR3 (N2783, N2773, N2704, N2359);
and AND2 (N2784, N2781, N660);
or OR3 (N2785, N2757, N968, N1988);
not NOT1 (N2786, N2785);
nand NAND4 (N2787, N2755, N1459, N2264, N547);
xor XOR2 (N2788, N2770, N693);
and AND3 (N2789, N2788, N1293, N890);
or OR3 (N2790, N2779, N2244, N1764);
not NOT1 (N2791, N2790);
buf BUF1 (N2792, N2776);
nand NAND3 (N2793, N2783, N1316, N261);
buf BUF1 (N2794, N2793);
xor XOR2 (N2795, N2791, N1224);
xor XOR2 (N2796, N2782, N397);
or OR3 (N2797, N2794, N2417, N2406);
nand NAND3 (N2798, N2792, N2277, N2716);
nand NAND4 (N2799, N2789, N978, N297, N753);
nor NOR4 (N2800, N2796, N373, N204, N1936);
nor NOR4 (N2801, N2761, N2105, N1502, N2553);
xor XOR2 (N2802, N2797, N1331);
or OR2 (N2803, N2800, N1344);
nand NAND3 (N2804, N2801, N191, N649);
xor XOR2 (N2805, N2799, N2218);
not NOT1 (N2806, N2778);
nand NAND2 (N2807, N2786, N691);
nor NOR4 (N2808, N2803, N1520, N977, N1887);
nand NAND2 (N2809, N2784, N1840);
buf BUF1 (N2810, N2802);
buf BUF1 (N2811, N2808);
xor XOR2 (N2812, N2809, N710);
nor NOR3 (N2813, N2810, N1516, N788);
buf BUF1 (N2814, N2798);
buf BUF1 (N2815, N2787);
nor NOR4 (N2816, N2805, N2028, N781, N976);
or OR2 (N2817, N2812, N1791);
buf BUF1 (N2818, N2811);
nand NAND4 (N2819, N2795, N1610, N407, N851);
not NOT1 (N2820, N2804);
buf BUF1 (N2821, N2813);
buf BUF1 (N2822, N2821);
nor NOR3 (N2823, N2816, N2275, N433);
and AND3 (N2824, N2806, N2029, N757);
and AND3 (N2825, N2824, N113, N2651);
buf BUF1 (N2826, N2819);
xor XOR2 (N2827, N2823, N2385);
xor XOR2 (N2828, N2825, N2388);
not NOT1 (N2829, N2826);
buf BUF1 (N2830, N2815);
or OR3 (N2831, N2814, N1269, N1465);
nand NAND3 (N2832, N2820, N2750, N1862);
nand NAND2 (N2833, N2830, N188);
buf BUF1 (N2834, N2818);
xor XOR2 (N2835, N2834, N1453);
nor NOR3 (N2836, N2822, N1287, N1324);
nor NOR2 (N2837, N2817, N780);
nor NOR2 (N2838, N2807, N860);
nor NOR2 (N2839, N2831, N519);
and AND3 (N2840, N2839, N1687, N153);
or OR2 (N2841, N2828, N1266);
not NOT1 (N2842, N2833);
buf BUF1 (N2843, N2837);
xor XOR2 (N2844, N2836, N484);
or OR2 (N2845, N2829, N1112);
nor NOR2 (N2846, N2842, N363);
not NOT1 (N2847, N2835);
xor XOR2 (N2848, N2827, N591);
not NOT1 (N2849, N2848);
not NOT1 (N2850, N2841);
nor NOR3 (N2851, N2849, N2672, N133);
nand NAND4 (N2852, N2846, N1506, N129, N2632);
or OR4 (N2853, N2832, N726, N421, N950);
nor NOR2 (N2854, N2838, N982);
xor XOR2 (N2855, N2840, N2651);
and AND4 (N2856, N2851, N1417, N219, N678);
not NOT1 (N2857, N2856);
buf BUF1 (N2858, N2857);
nor NOR3 (N2859, N2858, N1319, N993);
buf BUF1 (N2860, N2845);
nor NOR4 (N2861, N2852, N1151, N2032, N2220);
or OR4 (N2862, N2859, N246, N2416, N2349);
nand NAND3 (N2863, N2847, N1554, N272);
xor XOR2 (N2864, N2855, N286);
and AND4 (N2865, N2854, N1323, N1264, N38);
and AND3 (N2866, N2861, N1574, N1192);
not NOT1 (N2867, N2865);
or OR4 (N2868, N2867, N1459, N2613, N1302);
or OR2 (N2869, N2866, N276);
or OR3 (N2870, N2843, N1241, N747);
buf BUF1 (N2871, N2870);
buf BUF1 (N2872, N2844);
not NOT1 (N2873, N2860);
or OR4 (N2874, N2868, N2476, N2715, N965);
xor XOR2 (N2875, N2850, N1625);
xor XOR2 (N2876, N2853, N550);
or OR3 (N2877, N2864, N1004, N2468);
buf BUF1 (N2878, N2874);
xor XOR2 (N2879, N2873, N1705);
nand NAND3 (N2880, N2878, N567, N1483);
not NOT1 (N2881, N2876);
nand NAND4 (N2882, N2875, N2088, N2808, N2758);
nor NOR4 (N2883, N2863, N1543, N2439, N1141);
nand NAND3 (N2884, N2862, N2740, N1365);
buf BUF1 (N2885, N2872);
nor NOR3 (N2886, N2882, N1274, N1910);
not NOT1 (N2887, N2869);
not NOT1 (N2888, N2883);
not NOT1 (N2889, N2888);
xor XOR2 (N2890, N2889, N2787);
or OR2 (N2891, N2879, N501);
buf BUF1 (N2892, N2884);
nand NAND4 (N2893, N2887, N553, N349, N578);
or OR3 (N2894, N2881, N2316, N319);
or OR3 (N2895, N2885, N1103, N1510);
and AND4 (N2896, N2893, N2316, N1467, N1994);
nor NOR3 (N2897, N2890, N908, N2542);
not NOT1 (N2898, N2892);
and AND4 (N2899, N2897, N456, N117, N2233);
nand NAND2 (N2900, N2899, N1885);
xor XOR2 (N2901, N2871, N2068);
buf BUF1 (N2902, N2895);
or OR4 (N2903, N2880, N2395, N2017, N1027);
and AND2 (N2904, N2877, N222);
not NOT1 (N2905, N2886);
and AND3 (N2906, N2901, N404, N1676);
not NOT1 (N2907, N2902);
or OR2 (N2908, N2906, N111);
not NOT1 (N2909, N2907);
buf BUF1 (N2910, N2905);
and AND3 (N2911, N2900, N2692, N2866);
nor NOR3 (N2912, N2898, N2749, N209);
or OR4 (N2913, N2912, N1786, N2348, N1697);
or OR3 (N2914, N2896, N971, N1797);
xor XOR2 (N2915, N2913, N708);
nand NAND4 (N2916, N2908, N1485, N2034, N569);
xor XOR2 (N2917, N2904, N2792);
or OR2 (N2918, N2909, N1301);
and AND4 (N2919, N2917, N1081, N2063, N2271);
nor NOR4 (N2920, N2910, N745, N1445, N2605);
nor NOR4 (N2921, N2903, N2404, N224, N1947);
and AND4 (N2922, N2920, N7, N336, N184);
and AND3 (N2923, N2914, N59, N1030);
nand NAND4 (N2924, N2894, N500, N2535, N1149);
xor XOR2 (N2925, N2923, N571);
or OR2 (N2926, N2918, N485);
or OR3 (N2927, N2924, N1030, N2300);
and AND3 (N2928, N2919, N1530, N1518);
buf BUF1 (N2929, N2926);
not NOT1 (N2930, N2927);
nor NOR2 (N2931, N2915, N362);
buf BUF1 (N2932, N2931);
nand NAND3 (N2933, N2932, N2142, N2420);
xor XOR2 (N2934, N2922, N2328);
not NOT1 (N2935, N2929);
nor NOR2 (N2936, N2925, N1318);
nor NOR3 (N2937, N2916, N2451, N2742);
and AND2 (N2938, N2934, N2050);
nand NAND2 (N2939, N2936, N1346);
nand NAND2 (N2940, N2935, N699);
xor XOR2 (N2941, N2933, N279);
xor XOR2 (N2942, N2937, N2208);
not NOT1 (N2943, N2940);
or OR4 (N2944, N2928, N2340, N1993, N2383);
and AND4 (N2945, N2911, N186, N1402, N2158);
and AND2 (N2946, N2938, N2403);
nand NAND2 (N2947, N2921, N428);
buf BUF1 (N2948, N2942);
nor NOR4 (N2949, N2946, N862, N1184, N1894);
not NOT1 (N2950, N2943);
and AND4 (N2951, N2939, N137, N332, N998);
or OR2 (N2952, N2951, N2396);
not NOT1 (N2953, N2930);
buf BUF1 (N2954, N2941);
nand NAND4 (N2955, N2953, N291, N1324, N595);
nor NOR4 (N2956, N2947, N2281, N406, N1770);
not NOT1 (N2957, N2944);
nor NOR3 (N2958, N2956, N553, N1668);
not NOT1 (N2959, N2891);
buf BUF1 (N2960, N2952);
and AND3 (N2961, N2954, N2903, N2597);
buf BUF1 (N2962, N2960);
nor NOR4 (N2963, N2961, N2638, N367, N331);
buf BUF1 (N2964, N2945);
or OR2 (N2965, N2958, N514);
buf BUF1 (N2966, N2964);
nand NAND4 (N2967, N2962, N2014, N1795, N2422);
nand NAND2 (N2968, N2949, N933);
buf BUF1 (N2969, N2968);
or OR4 (N2970, N2955, N2816, N478, N2455);
buf BUF1 (N2971, N2950);
nand NAND4 (N2972, N2963, N1037, N2805, N356);
xor XOR2 (N2973, N2969, N690);
buf BUF1 (N2974, N2959);
nor NOR3 (N2975, N2965, N128, N1171);
nor NOR2 (N2976, N2972, N2743);
buf BUF1 (N2977, N2975);
not NOT1 (N2978, N2971);
nor NOR3 (N2979, N2977, N1575, N1936);
and AND3 (N2980, N2967, N2973, N2910);
and AND3 (N2981, N2741, N541, N848);
not NOT1 (N2982, N2948);
nor NOR2 (N2983, N2970, N2436);
and AND4 (N2984, N2982, N1018, N1787, N1386);
xor XOR2 (N2985, N2981, N1487);
nor NOR2 (N2986, N2984, N2407);
and AND2 (N2987, N2979, N2426);
nand NAND2 (N2988, N2957, N2738);
not NOT1 (N2989, N2978);
xor XOR2 (N2990, N2974, N255);
nand NAND4 (N2991, N2990, N815, N2128, N958);
and AND3 (N2992, N2976, N135, N1638);
nand NAND3 (N2993, N2987, N900, N342);
or OR3 (N2994, N2986, N2775, N2716);
buf BUF1 (N2995, N2992);
and AND2 (N2996, N2995, N2960);
buf BUF1 (N2997, N2988);
xor XOR2 (N2998, N2983, N1927);
and AND4 (N2999, N2966, N304, N202, N594);
nor NOR4 (N3000, N2985, N1553, N2055, N2588);
xor XOR2 (N3001, N2980, N2521);
or OR3 (N3002, N2994, N656, N2153);
xor XOR2 (N3003, N2993, N296);
buf BUF1 (N3004, N3002);
xor XOR2 (N3005, N3000, N2811);
buf BUF1 (N3006, N2997);
nor NOR3 (N3007, N3006, N864, N404);
nor NOR4 (N3008, N3007, N2712, N267, N970);
nand NAND4 (N3009, N3001, N2605, N617, N2631);
and AND3 (N3010, N3009, N2424, N2105);
nor NOR2 (N3011, N2999, N1177);
buf BUF1 (N3012, N2991);
buf BUF1 (N3013, N2989);
and AND4 (N3014, N3012, N713, N250, N47);
nor NOR3 (N3015, N3011, N1817, N1939);
xor XOR2 (N3016, N2998, N275);
not NOT1 (N3017, N3003);
nand NAND3 (N3018, N3015, N285, N841);
not NOT1 (N3019, N3013);
nand NAND4 (N3020, N3010, N2341, N1253, N1010);
nor NOR2 (N3021, N3019, N2630);
not NOT1 (N3022, N3008);
nor NOR4 (N3023, N3017, N237, N443, N1221);
buf BUF1 (N3024, N2996);
nor NOR4 (N3025, N3020, N1375, N961, N2573);
nor NOR2 (N3026, N3024, N1784);
and AND3 (N3027, N3004, N2116, N788);
xor XOR2 (N3028, N3027, N1196);
or OR3 (N3029, N3028, N1721, N2292);
or OR2 (N3030, N3005, N174);
nand NAND2 (N3031, N3030, N3006);
or OR3 (N3032, N3025, N1778, N675);
nand NAND4 (N3033, N3032, N35, N2006, N924);
buf BUF1 (N3034, N3031);
and AND3 (N3035, N3022, N28, N1533);
nand NAND4 (N3036, N3033, N1036, N2097, N1546);
buf BUF1 (N3037, N3034);
buf BUF1 (N3038, N3021);
not NOT1 (N3039, N3018);
nor NOR4 (N3040, N3014, N666, N2805, N292);
xor XOR2 (N3041, N3037, N1813);
buf BUF1 (N3042, N3016);
or OR4 (N3043, N3040, N2707, N1274, N935);
not NOT1 (N3044, N3036);
and AND4 (N3045, N3042, N2233, N1441, N2658);
buf BUF1 (N3046, N3023);
or OR4 (N3047, N3045, N2658, N1038, N852);
not NOT1 (N3048, N3046);
nand NAND2 (N3049, N3044, N1667);
nor NOR3 (N3050, N3049, N367, N2766);
buf BUF1 (N3051, N3038);
and AND2 (N3052, N3041, N30);
or OR2 (N3053, N3039, N1109);
nand NAND2 (N3054, N3035, N556);
buf BUF1 (N3055, N3052);
nor NOR2 (N3056, N3029, N971);
and AND2 (N3057, N3056, N2919);
nor NOR2 (N3058, N3053, N1850);
nor NOR3 (N3059, N3050, N1, N1273);
not NOT1 (N3060, N3055);
nor NOR2 (N3061, N3048, N1110);
not NOT1 (N3062, N3026);
buf BUF1 (N3063, N3054);
nor NOR2 (N3064, N3060, N2355);
nor NOR2 (N3065, N3051, N593);
nor NOR3 (N3066, N3061, N2283, N1096);
nand NAND3 (N3067, N3062, N1768, N911);
and AND4 (N3068, N3064, N1331, N1883, N2237);
nand NAND4 (N3069, N3043, N724, N1000, N1218);
nand NAND2 (N3070, N3057, N2767);
buf BUF1 (N3071, N3067);
nor NOR4 (N3072, N3047, N334, N637, N664);
not NOT1 (N3073, N3066);
or OR3 (N3074, N3063, N1533, N1078);
buf BUF1 (N3075, N3068);
and AND3 (N3076, N3072, N92, N184);
and AND2 (N3077, N3075, N2229);
and AND2 (N3078, N3071, N677);
nand NAND2 (N3079, N3069, N2935);
or OR3 (N3080, N3077, N3032, N2979);
or OR2 (N3081, N3070, N2723);
buf BUF1 (N3082, N3076);
nor NOR3 (N3083, N3059, N2503, N2458);
buf BUF1 (N3084, N3073);
buf BUF1 (N3085, N3079);
and AND3 (N3086, N3082, N689, N1308);
not NOT1 (N3087, N3081);
xor XOR2 (N3088, N3085, N1803);
and AND3 (N3089, N3086, N1351, N1118);
and AND2 (N3090, N3089, N2273);
xor XOR2 (N3091, N3080, N377);
xor XOR2 (N3092, N3088, N2155);
not NOT1 (N3093, N3087);
xor XOR2 (N3094, N3078, N1268);
nand NAND3 (N3095, N3083, N477, N3093);
nor NOR3 (N3096, N2850, N1196, N1095);
not NOT1 (N3097, N3091);
or OR2 (N3098, N3095, N168);
and AND2 (N3099, N3090, N1868);
xor XOR2 (N3100, N3099, N2912);
nand NAND2 (N3101, N3084, N1718);
xor XOR2 (N3102, N3101, N2563);
not NOT1 (N3103, N3102);
not NOT1 (N3104, N3074);
nor NOR3 (N3105, N3092, N545, N703);
and AND4 (N3106, N3104, N616, N267, N2052);
nor NOR4 (N3107, N3106, N657, N2195, N2030);
or OR2 (N3108, N3105, N2623);
nor NOR3 (N3109, N3065, N469, N1334);
or OR3 (N3110, N3096, N2060, N2059);
and AND3 (N3111, N3097, N2841, N3026);
nor NOR3 (N3112, N3094, N2908, N507);
nand NAND4 (N3113, N3112, N449, N987, N1136);
or OR3 (N3114, N3111, N248, N1291);
buf BUF1 (N3115, N3108);
not NOT1 (N3116, N3103);
not NOT1 (N3117, N3098);
nor NOR3 (N3118, N3117, N1388, N567);
nor NOR2 (N3119, N3118, N2873);
buf BUF1 (N3120, N3119);
buf BUF1 (N3121, N3114);
not NOT1 (N3122, N3115);
nand NAND3 (N3123, N3109, N2004, N2342);
nor NOR3 (N3124, N3110, N2806, N1641);
or OR2 (N3125, N3124, N117);
xor XOR2 (N3126, N3116, N1240);
xor XOR2 (N3127, N3126, N789);
nor NOR2 (N3128, N3121, N2291);
buf BUF1 (N3129, N3122);
nor NOR4 (N3130, N3128, N789, N1641, N1917);
xor XOR2 (N3131, N3100, N888);
xor XOR2 (N3132, N3131, N1181);
nor NOR2 (N3133, N3127, N2714);
and AND2 (N3134, N3058, N2204);
not NOT1 (N3135, N3125);
nor NOR3 (N3136, N3107, N3091, N1983);
not NOT1 (N3137, N3120);
or OR3 (N3138, N3123, N190, N2300);
nor NOR3 (N3139, N3129, N3079, N1310);
nor NOR4 (N3140, N3130, N280, N935, N2362);
xor XOR2 (N3141, N3135, N2474);
not NOT1 (N3142, N3141);
or OR3 (N3143, N3142, N1560, N2711);
xor XOR2 (N3144, N3132, N1089);
nand NAND4 (N3145, N3137, N1877, N799, N2085);
buf BUF1 (N3146, N3139);
xor XOR2 (N3147, N3143, N1245);
nand NAND2 (N3148, N3144, N1327);
not NOT1 (N3149, N3133);
buf BUF1 (N3150, N3138);
buf BUF1 (N3151, N3113);
and AND3 (N3152, N3146, N1560, N280);
xor XOR2 (N3153, N3148, N1444);
nand NAND3 (N3154, N3150, N3089, N586);
nand NAND3 (N3155, N3152, N2697, N1724);
or OR4 (N3156, N3140, N139, N777, N1947);
not NOT1 (N3157, N3136);
and AND4 (N3158, N3156, N1150, N1882, N2233);
xor XOR2 (N3159, N3145, N2927);
buf BUF1 (N3160, N3147);
xor XOR2 (N3161, N3134, N2411);
buf BUF1 (N3162, N3151);
not NOT1 (N3163, N3157);
or OR2 (N3164, N3163, N2869);
not NOT1 (N3165, N3153);
nor NOR2 (N3166, N3155, N2464);
not NOT1 (N3167, N3149);
not NOT1 (N3168, N3160);
and AND4 (N3169, N3166, N2447, N606, N2262);
nor NOR2 (N3170, N3159, N1659);
nand NAND3 (N3171, N3164, N1628, N636);
not NOT1 (N3172, N3170);
nand NAND2 (N3173, N3161, N2231);
not NOT1 (N3174, N3173);
nor NOR2 (N3175, N3158, N2230);
nor NOR3 (N3176, N3174, N422, N3010);
nand NAND3 (N3177, N3162, N463, N2081);
xor XOR2 (N3178, N3165, N3124);
and AND2 (N3179, N3154, N3081);
buf BUF1 (N3180, N3179);
nor NOR2 (N3181, N3168, N2706);
and AND3 (N3182, N3177, N2077, N1232);
or OR2 (N3183, N3181, N2027);
or OR2 (N3184, N3180, N562);
nor NOR4 (N3185, N3182, N799, N2929, N2670);
buf BUF1 (N3186, N3169);
nor NOR3 (N3187, N3178, N765, N2227);
nand NAND3 (N3188, N3175, N1658, N1560);
buf BUF1 (N3189, N3187);
not NOT1 (N3190, N3172);
or OR3 (N3191, N3189, N1097, N606);
nand NAND4 (N3192, N3185, N3016, N662, N45);
buf BUF1 (N3193, N3167);
not NOT1 (N3194, N3190);
xor XOR2 (N3195, N3188, N2162);
not NOT1 (N3196, N3191);
xor XOR2 (N3197, N3193, N3186);
not NOT1 (N3198, N1353);
and AND2 (N3199, N3184, N849);
buf BUF1 (N3200, N3196);
nand NAND2 (N3201, N3171, N144);
buf BUF1 (N3202, N3198);
nand NAND3 (N3203, N3197, N2410, N2639);
or OR2 (N3204, N3202, N1956);
and AND2 (N3205, N3176, N3143);
xor XOR2 (N3206, N3203, N2672);
not NOT1 (N3207, N3194);
not NOT1 (N3208, N3195);
buf BUF1 (N3209, N3206);
buf BUF1 (N3210, N3183);
or OR4 (N3211, N3192, N1819, N516, N1100);
not NOT1 (N3212, N3200);
buf BUF1 (N3213, N3212);
nand NAND2 (N3214, N3213, N35);
buf BUF1 (N3215, N3214);
and AND2 (N3216, N3210, N493);
not NOT1 (N3217, N3207);
nand NAND2 (N3218, N3216, N1600);
buf BUF1 (N3219, N3209);
xor XOR2 (N3220, N3199, N1063);
and AND2 (N3221, N3219, N481);
and AND2 (N3222, N3218, N1144);
nor NOR4 (N3223, N3215, N2742, N2804, N87);
not NOT1 (N3224, N3217);
buf BUF1 (N3225, N3220);
nand NAND4 (N3226, N3222, N1384, N406, N2288);
or OR2 (N3227, N3223, N2249);
or OR2 (N3228, N3225, N2342);
nand NAND4 (N3229, N3226, N2450, N142, N1305);
and AND3 (N3230, N3208, N2865, N2762);
xor XOR2 (N3231, N3227, N216);
nand NAND3 (N3232, N3228, N1691, N1041);
not NOT1 (N3233, N3229);
nand NAND4 (N3234, N3221, N3170, N1477, N2622);
not NOT1 (N3235, N3224);
nand NAND2 (N3236, N3235, N845);
nor NOR2 (N3237, N3236, N843);
not NOT1 (N3238, N3232);
nor NOR3 (N3239, N3230, N1840, N1706);
not NOT1 (N3240, N3238);
nor NOR3 (N3241, N3231, N610, N632);
or OR3 (N3242, N3205, N3238, N197);
and AND2 (N3243, N3241, N205);
or OR3 (N3244, N3242, N1771, N62);
and AND3 (N3245, N3243, N1201, N1279);
nand NAND2 (N3246, N3234, N1581);
not NOT1 (N3247, N3245);
nor NOR2 (N3248, N3237, N1775);
nand NAND3 (N3249, N3248, N1513, N1846);
nor NOR4 (N3250, N3249, N1562, N2785, N915);
buf BUF1 (N3251, N3233);
or OR3 (N3252, N3246, N2109, N1465);
and AND4 (N3253, N3252, N2439, N2440, N1807);
buf BUF1 (N3254, N3253);
or OR3 (N3255, N3244, N1299, N1899);
nor NOR2 (N3256, N3255, N802);
xor XOR2 (N3257, N3240, N363);
nor NOR3 (N3258, N3256, N775, N130);
nor NOR3 (N3259, N3257, N2712, N973);
and AND4 (N3260, N3211, N1584, N397, N834);
xor XOR2 (N3261, N3251, N479);
nor NOR4 (N3262, N3254, N2535, N310, N2767);
xor XOR2 (N3263, N3259, N2095);
nor NOR2 (N3264, N3201, N98);
nand NAND2 (N3265, N3258, N832);
buf BUF1 (N3266, N3260);
and AND2 (N3267, N3204, N2866);
xor XOR2 (N3268, N3239, N3211);
nor NOR2 (N3269, N3261, N334);
or OR4 (N3270, N3266, N1429, N636, N1876);
and AND2 (N3271, N3262, N933);
xor XOR2 (N3272, N3263, N2424);
and AND3 (N3273, N3268, N2623, N1813);
nor NOR3 (N3274, N3250, N2603, N2220);
nand NAND4 (N3275, N3269, N371, N3208, N1399);
nor NOR3 (N3276, N3264, N1247, N1594);
or OR3 (N3277, N3272, N2313, N1091);
and AND3 (N3278, N3247, N2206, N1369);
nand NAND2 (N3279, N3277, N216);
nor NOR4 (N3280, N3279, N14, N141, N1518);
not NOT1 (N3281, N3265);
and AND3 (N3282, N3273, N1387, N2932);
and AND3 (N3283, N3276, N1668, N4);
nand NAND2 (N3284, N3270, N1361);
or OR4 (N3285, N3284, N2874, N3020, N1029);
nand NAND4 (N3286, N3275, N2554, N1777, N3047);
nand NAND3 (N3287, N3285, N2859, N1369);
and AND3 (N3288, N3278, N1505, N2020);
xor XOR2 (N3289, N3280, N366);
nor NOR2 (N3290, N3267, N3005);
not NOT1 (N3291, N3288);
buf BUF1 (N3292, N3291);
nor NOR2 (N3293, N3271, N2889);
nor NOR2 (N3294, N3286, N2943);
nor NOR3 (N3295, N3290, N1737, N2318);
nor NOR4 (N3296, N3293, N3249, N987, N1103);
buf BUF1 (N3297, N3281);
nand NAND3 (N3298, N3297, N3107, N3106);
and AND3 (N3299, N3295, N1902, N2331);
buf BUF1 (N3300, N3287);
or OR4 (N3301, N3298, N2548, N3183, N3192);
or OR3 (N3302, N3282, N780, N2477);
not NOT1 (N3303, N3274);
nand NAND3 (N3304, N3300, N3003, N2048);
xor XOR2 (N3305, N3292, N356);
or OR2 (N3306, N3302, N2301);
or OR4 (N3307, N3299, N3306, N1237, N2386);
buf BUF1 (N3308, N1);
nor NOR2 (N3309, N3296, N856);
nand NAND3 (N3310, N3294, N2755, N541);
xor XOR2 (N3311, N3301, N1836);
buf BUF1 (N3312, N3304);
buf BUF1 (N3313, N3305);
not NOT1 (N3314, N3283);
and AND3 (N3315, N3309, N720, N2353);
and AND4 (N3316, N3308, N456, N589, N590);
or OR4 (N3317, N3315, N2177, N977, N1009);
or OR4 (N3318, N3307, N1102, N81, N820);
and AND3 (N3319, N3318, N1394, N463);
xor XOR2 (N3320, N3303, N987);
not NOT1 (N3321, N3316);
nand NAND3 (N3322, N3311, N2962, N2276);
nor NOR2 (N3323, N3310, N1915);
nor NOR2 (N3324, N3317, N1269);
xor XOR2 (N3325, N3314, N2343);
nand NAND4 (N3326, N3323, N1388, N3307, N1498);
not NOT1 (N3327, N3313);
and AND3 (N3328, N3325, N1105, N1502);
xor XOR2 (N3329, N3322, N747);
xor XOR2 (N3330, N3324, N3245);
nand NAND2 (N3331, N3328, N3214);
or OR2 (N3332, N3320, N2532);
nor NOR4 (N3333, N3319, N2100, N3204, N427);
buf BUF1 (N3334, N3289);
buf BUF1 (N3335, N3321);
nand NAND2 (N3336, N3329, N31);
xor XOR2 (N3337, N3334, N2309);
xor XOR2 (N3338, N3332, N1422);
and AND2 (N3339, N3338, N1666);
nor NOR4 (N3340, N3330, N2823, N2250, N233);
or OR2 (N3341, N3333, N498);
nor NOR4 (N3342, N3331, N729, N1428, N2399);
not NOT1 (N3343, N3312);
nand NAND4 (N3344, N3336, N3077, N967, N1263);
not NOT1 (N3345, N3339);
and AND4 (N3346, N3344, N1211, N841, N1176);
or OR3 (N3347, N3340, N1798, N2641);
nand NAND2 (N3348, N3342, N2998);
and AND4 (N3349, N3326, N2929, N1691, N1529);
nor NOR3 (N3350, N3349, N1122, N530);
buf BUF1 (N3351, N3337);
and AND3 (N3352, N3351, N1147, N2779);
nor NOR4 (N3353, N3327, N3220, N666, N1743);
xor XOR2 (N3354, N3343, N22);
xor XOR2 (N3355, N3354, N2506);
buf BUF1 (N3356, N3353);
buf BUF1 (N3357, N3335);
or OR4 (N3358, N3352, N2619, N3171, N1446);
nor NOR3 (N3359, N3348, N2695, N1652);
not NOT1 (N3360, N3355);
or OR3 (N3361, N3345, N2546, N2490);
nor NOR3 (N3362, N3359, N404, N3340);
nor NOR4 (N3363, N3361, N528, N123, N1903);
xor XOR2 (N3364, N3356, N1885);
not NOT1 (N3365, N3350);
xor XOR2 (N3366, N3347, N1604);
buf BUF1 (N3367, N3341);
not NOT1 (N3368, N3358);
buf BUF1 (N3369, N3360);
buf BUF1 (N3370, N3365);
nand NAND2 (N3371, N3363, N3019);
xor XOR2 (N3372, N3369, N2350);
and AND2 (N3373, N3367, N1903);
not NOT1 (N3374, N3364);
xor XOR2 (N3375, N3357, N530);
and AND3 (N3376, N3373, N3221, N459);
or OR3 (N3377, N3366, N679, N1966);
nand NAND3 (N3378, N3370, N3251, N1451);
and AND4 (N3379, N3375, N898, N431, N2437);
xor XOR2 (N3380, N3377, N1990);
nand NAND3 (N3381, N3374, N2679, N362);
nor NOR4 (N3382, N3379, N159, N217, N571);
buf BUF1 (N3383, N3371);
nor NOR4 (N3384, N3381, N1614, N152, N2478);
nand NAND2 (N3385, N3383, N1565);
xor XOR2 (N3386, N3385, N1337);
or OR3 (N3387, N3384, N2838, N949);
or OR3 (N3388, N3380, N11, N1823);
not NOT1 (N3389, N3378);
not NOT1 (N3390, N3387);
or OR4 (N3391, N3386, N3119, N609, N445);
xor XOR2 (N3392, N3390, N261);
nor NOR4 (N3393, N3372, N3141, N2098, N2000);
buf BUF1 (N3394, N3391);
xor XOR2 (N3395, N3382, N2679);
buf BUF1 (N3396, N3388);
and AND2 (N3397, N3389, N3035);
xor XOR2 (N3398, N3376, N1757);
and AND2 (N3399, N3398, N1027);
or OR4 (N3400, N3394, N2491, N2009, N360);
nor NOR3 (N3401, N3346, N3124, N2126);
and AND2 (N3402, N3401, N1082);
and AND4 (N3403, N3362, N2364, N2339, N2913);
nor NOR3 (N3404, N3403, N1427, N2377);
not NOT1 (N3405, N3368);
nor NOR3 (N3406, N3402, N1929, N513);
buf BUF1 (N3407, N3396);
nand NAND2 (N3408, N3397, N2516);
or OR2 (N3409, N3400, N125);
and AND4 (N3410, N3399, N1730, N2195, N2368);
nor NOR3 (N3411, N3393, N724, N2755);
buf BUF1 (N3412, N3408);
xor XOR2 (N3413, N3392, N975);
xor XOR2 (N3414, N3410, N3301);
or OR4 (N3415, N3412, N1091, N1725, N523);
xor XOR2 (N3416, N3407, N3118);
nor NOR3 (N3417, N3413, N2808, N1891);
and AND3 (N3418, N3409, N2245, N892);
xor XOR2 (N3419, N3417, N309);
or OR2 (N3420, N3419, N648);
or OR3 (N3421, N3420, N383, N2878);
xor XOR2 (N3422, N3395, N2112);
buf BUF1 (N3423, N3406);
or OR4 (N3424, N3421, N280, N2430, N2692);
nand NAND4 (N3425, N3424, N764, N565, N82);
buf BUF1 (N3426, N3418);
nor NOR3 (N3427, N3423, N2378, N2413);
and AND4 (N3428, N3416, N302, N1461, N2085);
nor NOR3 (N3429, N3425, N2423, N263);
and AND4 (N3430, N3411, N349, N384, N3291);
and AND3 (N3431, N3426, N2404, N816);
buf BUF1 (N3432, N3415);
or OR2 (N3433, N3428, N541);
or OR4 (N3434, N3414, N2959, N1340, N2117);
nor NOR3 (N3435, N3405, N1045, N1283);
buf BUF1 (N3436, N3429);
or OR2 (N3437, N3434, N1810);
nand NAND2 (N3438, N3404, N1354);
nor NOR4 (N3439, N3436, N2081, N2268, N2906);
or OR3 (N3440, N3439, N922, N102);
nor NOR2 (N3441, N3438, N2567);
nand NAND4 (N3442, N3437, N2035, N2552, N1248);
buf BUF1 (N3443, N3442);
not NOT1 (N3444, N3433);
and AND3 (N3445, N3443, N884, N521);
buf BUF1 (N3446, N3441);
nor NOR3 (N3447, N3444, N2788, N1132);
and AND2 (N3448, N3432, N1844);
or OR3 (N3449, N3446, N2241, N2074);
nor NOR4 (N3450, N3445, N856, N2309, N3173);
nand NAND3 (N3451, N3450, N1474, N1701);
nor NOR2 (N3452, N3435, N335);
nand NAND4 (N3453, N3451, N3402, N3152, N1665);
buf BUF1 (N3454, N3430);
buf BUF1 (N3455, N3422);
not NOT1 (N3456, N3427);
nor NOR4 (N3457, N3455, N1182, N2557, N1722);
and AND4 (N3458, N3447, N1518, N2981, N2294);
and AND3 (N3459, N3452, N3369, N1251);
not NOT1 (N3460, N3457);
buf BUF1 (N3461, N3453);
not NOT1 (N3462, N3454);
or OR4 (N3463, N3448, N109, N92, N2971);
and AND2 (N3464, N3458, N7);
nor NOR4 (N3465, N3462, N2995, N622, N3141);
nand NAND3 (N3466, N3460, N3285, N860);
xor XOR2 (N3467, N3465, N1381);
nor NOR4 (N3468, N3459, N51, N1454, N909);
and AND2 (N3469, N3456, N1735);
nand NAND3 (N3470, N3461, N497, N636);
xor XOR2 (N3471, N3470, N1811);
and AND2 (N3472, N3468, N3383);
nor NOR3 (N3473, N3471, N2575, N1616);
or OR3 (N3474, N3469, N588, N178);
and AND3 (N3475, N3464, N1826, N2893);
buf BUF1 (N3476, N3431);
or OR2 (N3477, N3440, N305);
or OR4 (N3478, N3449, N158, N2490, N727);
nor NOR2 (N3479, N3463, N2732);
not NOT1 (N3480, N3477);
nor NOR2 (N3481, N3479, N3098);
nor NOR2 (N3482, N3478, N2426);
nand NAND2 (N3483, N3466, N2361);
not NOT1 (N3484, N3472);
or OR4 (N3485, N3474, N2030, N3470, N1059);
not NOT1 (N3486, N3485);
xor XOR2 (N3487, N3484, N437);
xor XOR2 (N3488, N3482, N523);
buf BUF1 (N3489, N3480);
and AND4 (N3490, N3489, N1709, N3312, N2686);
and AND2 (N3491, N3476, N2938);
not NOT1 (N3492, N3481);
nor NOR4 (N3493, N3490, N2309, N791, N241);
nor NOR2 (N3494, N3473, N1399);
and AND2 (N3495, N3491, N1301);
nand NAND3 (N3496, N3494, N403, N786);
or OR3 (N3497, N3488, N2027, N3072);
nor NOR2 (N3498, N3497, N1140);
not NOT1 (N3499, N3475);
nand NAND3 (N3500, N3486, N1188, N670);
nand NAND2 (N3501, N3495, N2267);
xor XOR2 (N3502, N3483, N3227);
or OR2 (N3503, N3498, N719);
xor XOR2 (N3504, N3492, N70);
nand NAND2 (N3505, N3504, N776);
or OR4 (N3506, N3493, N608, N348, N619);
and AND4 (N3507, N3496, N2491, N3042, N1617);
nor NOR2 (N3508, N3506, N3257);
not NOT1 (N3509, N3500);
nor NOR4 (N3510, N3505, N3139, N2636, N1484);
nor NOR2 (N3511, N3499, N100);
or OR4 (N3512, N3509, N1792, N3217, N2635);
buf BUF1 (N3513, N3508);
nor NOR4 (N3514, N3507, N3231, N127, N1091);
not NOT1 (N3515, N3487);
buf BUF1 (N3516, N3513);
nor NOR3 (N3517, N3502, N873, N3491);
or OR3 (N3518, N3510, N1476, N2205);
nor NOR4 (N3519, N3518, N1743, N1196, N760);
nand NAND2 (N3520, N3515, N2111);
and AND2 (N3521, N3467, N1900);
and AND2 (N3522, N3514, N925);
buf BUF1 (N3523, N3512);
and AND2 (N3524, N3511, N649);
nand NAND3 (N3525, N3519, N91, N3464);
buf BUF1 (N3526, N3503);
not NOT1 (N3527, N3516);
xor XOR2 (N3528, N3501, N2952);
xor XOR2 (N3529, N3522, N1017);
xor XOR2 (N3530, N3521, N3308);
nor NOR4 (N3531, N3530, N1893, N282, N2967);
buf BUF1 (N3532, N3526);
xor XOR2 (N3533, N3527, N573);
and AND3 (N3534, N3532, N545, N888);
and AND4 (N3535, N3531, N333, N2920, N206);
nand NAND2 (N3536, N3534, N3533);
nand NAND4 (N3537, N2458, N2503, N2459, N1103);
not NOT1 (N3538, N3537);
not NOT1 (N3539, N3520);
and AND4 (N3540, N3528, N724, N1117, N98);
not NOT1 (N3541, N3538);
nor NOR3 (N3542, N3524, N1965, N1922);
xor XOR2 (N3543, N3523, N2715);
nand NAND3 (N3544, N3529, N1477, N1887);
buf BUF1 (N3545, N3542);
not NOT1 (N3546, N3539);
nor NOR4 (N3547, N3535, N2971, N2264, N1808);
not NOT1 (N3548, N3540);
not NOT1 (N3549, N3547);
and AND2 (N3550, N3545, N2036);
nand NAND2 (N3551, N3543, N2520);
buf BUF1 (N3552, N3548);
buf BUF1 (N3553, N3552);
nor NOR4 (N3554, N3517, N3366, N845, N3482);
nand NAND2 (N3555, N3553, N3205);
buf BUF1 (N3556, N3555);
xor XOR2 (N3557, N3525, N1959);
buf BUF1 (N3558, N3550);
buf BUF1 (N3559, N3544);
xor XOR2 (N3560, N3554, N2965);
and AND2 (N3561, N3556, N248);
or OR3 (N3562, N3541, N1284, N1350);
nor NOR2 (N3563, N3549, N1002);
nor NOR3 (N3564, N3563, N438, N2857);
buf BUF1 (N3565, N3536);
nand NAND3 (N3566, N3557, N1245, N2813);
and AND3 (N3567, N3564, N2382, N3268);
and AND2 (N3568, N3560, N1636);
and AND4 (N3569, N3559, N2420, N35, N1251);
not NOT1 (N3570, N3558);
not NOT1 (N3571, N3568);
buf BUF1 (N3572, N3562);
nor NOR3 (N3573, N3572, N2473, N569);
not NOT1 (N3574, N3573);
nor NOR2 (N3575, N3567, N2400);
or OR2 (N3576, N3569, N3547);
buf BUF1 (N3577, N3566);
or OR4 (N3578, N3574, N1328, N740, N41);
buf BUF1 (N3579, N3575);
not NOT1 (N3580, N3570);
nor NOR4 (N3581, N3551, N3140, N816, N498);
nand NAND3 (N3582, N3580, N1730, N3336);
nor NOR2 (N3583, N3577, N1465);
not NOT1 (N3584, N3565);
nand NAND3 (N3585, N3581, N1185, N203);
not NOT1 (N3586, N3578);
and AND2 (N3587, N3584, N153);
nand NAND4 (N3588, N3587, N725, N730, N1130);
buf BUF1 (N3589, N3576);
xor XOR2 (N3590, N3585, N263);
buf BUF1 (N3591, N3571);
and AND3 (N3592, N3588, N3538, N102);
or OR2 (N3593, N3561, N3211);
buf BUF1 (N3594, N3579);
and AND3 (N3595, N3591, N2982, N216);
not NOT1 (N3596, N3546);
and AND2 (N3597, N3583, N3026);
not NOT1 (N3598, N3590);
not NOT1 (N3599, N3598);
not NOT1 (N3600, N3582);
not NOT1 (N3601, N3596);
nand NAND4 (N3602, N3601, N2515, N2025, N3477);
not NOT1 (N3603, N3586);
buf BUF1 (N3604, N3599);
and AND2 (N3605, N3595, N1573);
nand NAND4 (N3606, N3592, N3444, N968, N628);
and AND3 (N3607, N3605, N2485, N2318);
nor NOR2 (N3608, N3606, N2979);
nor NOR3 (N3609, N3589, N1096, N2488);
nand NAND4 (N3610, N3594, N2548, N720, N1791);
buf BUF1 (N3611, N3610);
and AND3 (N3612, N3602, N1664, N254);
xor XOR2 (N3613, N3609, N1760);
nand NAND3 (N3614, N3593, N1591, N1337);
buf BUF1 (N3615, N3613);
xor XOR2 (N3616, N3612, N218);
or OR4 (N3617, N3607, N615, N169, N533);
xor XOR2 (N3618, N3614, N444);
nor NOR4 (N3619, N3615, N3560, N1012, N570);
and AND4 (N3620, N3616, N2443, N2989, N1163);
nor NOR3 (N3621, N3620, N3347, N1013);
nand NAND2 (N3622, N3604, N895);
xor XOR2 (N3623, N3597, N3126);
buf BUF1 (N3624, N3600);
nor NOR4 (N3625, N3618, N1428, N3022, N1346);
buf BUF1 (N3626, N3611);
nand NAND3 (N3627, N3619, N2112, N713);
or OR3 (N3628, N3623, N2710, N2119);
not NOT1 (N3629, N3625);
nand NAND3 (N3630, N3622, N1251, N3129);
and AND3 (N3631, N3630, N3199, N231);
nor NOR2 (N3632, N3608, N2658);
nor NOR3 (N3633, N3617, N3044, N2994);
not NOT1 (N3634, N3629);
or OR2 (N3635, N3631, N2256);
buf BUF1 (N3636, N3635);
and AND3 (N3637, N3632, N2775, N2687);
or OR2 (N3638, N3624, N3150);
nor NOR3 (N3639, N3621, N2195, N1377);
buf BUF1 (N3640, N3636);
and AND3 (N3641, N3628, N3240, N210);
or OR2 (N3642, N3640, N2925);
or OR2 (N3643, N3638, N1804);
nor NOR3 (N3644, N3627, N2967, N3092);
nand NAND4 (N3645, N3642, N387, N2216, N2793);
and AND3 (N3646, N3634, N219, N2793);
nor NOR3 (N3647, N3641, N1572, N1211);
nand NAND4 (N3648, N3646, N2422, N20, N951);
or OR4 (N3649, N3633, N3589, N2623, N60);
or OR2 (N3650, N3647, N2926);
not NOT1 (N3651, N3637);
nand NAND4 (N3652, N3639, N1259, N2616, N1580);
nor NOR2 (N3653, N3650, N903);
xor XOR2 (N3654, N3651, N1576);
not NOT1 (N3655, N3653);
or OR4 (N3656, N3652, N1062, N1474, N3149);
not NOT1 (N3657, N3644);
xor XOR2 (N3658, N3648, N3301);
not NOT1 (N3659, N3649);
xor XOR2 (N3660, N3656, N1026);
not NOT1 (N3661, N3645);
or OR2 (N3662, N3643, N1010);
buf BUF1 (N3663, N3654);
nor NOR2 (N3664, N3659, N2268);
not NOT1 (N3665, N3658);
xor XOR2 (N3666, N3661, N1276);
xor XOR2 (N3667, N3626, N2674);
or OR4 (N3668, N3657, N2644, N2009, N152);
buf BUF1 (N3669, N3664);
xor XOR2 (N3670, N3667, N1691);
nor NOR4 (N3671, N3669, N727, N1981, N2015);
not NOT1 (N3672, N3603);
not NOT1 (N3673, N3666);
buf BUF1 (N3674, N3665);
buf BUF1 (N3675, N3662);
or OR2 (N3676, N3675, N1188);
or OR4 (N3677, N3674, N3417, N897, N2481);
and AND4 (N3678, N3671, N3559, N514, N460);
buf BUF1 (N3679, N3676);
buf BUF1 (N3680, N3663);
nand NAND3 (N3681, N3668, N2714, N1656);
not NOT1 (N3682, N3660);
not NOT1 (N3683, N3681);
or OR3 (N3684, N3679, N2499, N1829);
and AND4 (N3685, N3682, N726, N1632, N3544);
and AND3 (N3686, N3684, N1277, N3264);
not NOT1 (N3687, N3685);
and AND3 (N3688, N3672, N1302, N2669);
nand NAND2 (N3689, N3687, N3432);
nor NOR3 (N3690, N3686, N1233, N3603);
not NOT1 (N3691, N3677);
nand NAND4 (N3692, N3688, N2122, N3355, N1541);
and AND2 (N3693, N3689, N3376);
and AND2 (N3694, N3692, N1786);
and AND3 (N3695, N3670, N2654, N1904);
buf BUF1 (N3696, N3690);
or OR4 (N3697, N3695, N1378, N1053, N1547);
nand NAND3 (N3698, N3697, N229, N3172);
nand NAND4 (N3699, N3655, N896, N1811, N2096);
nand NAND4 (N3700, N3696, N699, N171, N2301);
nand NAND2 (N3701, N3680, N3153);
buf BUF1 (N3702, N3698);
nand NAND2 (N3703, N3673, N1104);
xor XOR2 (N3704, N3703, N2407);
buf BUF1 (N3705, N3693);
buf BUF1 (N3706, N3705);
nand NAND4 (N3707, N3699, N1986, N1363, N3664);
nor NOR2 (N3708, N3707, N2757);
buf BUF1 (N3709, N3691);
xor XOR2 (N3710, N3704, N2983);
not NOT1 (N3711, N3709);
nor NOR4 (N3712, N3700, N3277, N154, N3246);
nor NOR3 (N3713, N3694, N978, N8);
buf BUF1 (N3714, N3702);
and AND4 (N3715, N3713, N1071, N1204, N2320);
buf BUF1 (N3716, N3712);
xor XOR2 (N3717, N3716, N1890);
or OR3 (N3718, N3706, N3247, N1023);
and AND4 (N3719, N3715, N1390, N1577, N1127);
or OR3 (N3720, N3701, N123, N1935);
xor XOR2 (N3721, N3711, N2967);
nor NOR4 (N3722, N3683, N2059, N2639, N1176);
and AND4 (N3723, N3721, N1113, N3700, N3288);
not NOT1 (N3724, N3708);
not NOT1 (N3725, N3718);
xor XOR2 (N3726, N3717, N54);
buf BUF1 (N3727, N3724);
or OR2 (N3728, N3678, N35);
nor NOR3 (N3729, N3722, N1914, N2099);
nor NOR3 (N3730, N3726, N1745, N377);
nand NAND3 (N3731, N3719, N2683, N2346);
buf BUF1 (N3732, N3727);
buf BUF1 (N3733, N3725);
buf BUF1 (N3734, N3723);
buf BUF1 (N3735, N3731);
not NOT1 (N3736, N3720);
buf BUF1 (N3737, N3728);
nor NOR2 (N3738, N3737, N2760);
nand NAND2 (N3739, N3714, N2518);
nor NOR2 (N3740, N3730, N2213);
or OR3 (N3741, N3732, N2600, N1578);
buf BUF1 (N3742, N3739);
buf BUF1 (N3743, N3734);
buf BUF1 (N3744, N3741);
nand NAND4 (N3745, N3736, N3711, N614, N2276);
not NOT1 (N3746, N3740);
nand NAND2 (N3747, N3742, N1693);
buf BUF1 (N3748, N3746);
buf BUF1 (N3749, N3729);
nand NAND2 (N3750, N3744, N2954);
nor NOR3 (N3751, N3733, N1480, N2072);
nand NAND2 (N3752, N3743, N3036);
xor XOR2 (N3753, N3710, N2430);
nand NAND4 (N3754, N3752, N1818, N2776, N3441);
and AND3 (N3755, N3735, N1887, N2251);
nand NAND4 (N3756, N3748, N1396, N2783, N2251);
nand NAND3 (N3757, N3751, N3404, N2079);
nand NAND4 (N3758, N3747, N3627, N771, N2888);
xor XOR2 (N3759, N3758, N2778);
or OR3 (N3760, N3753, N823, N1809);
not NOT1 (N3761, N3760);
nor NOR4 (N3762, N3738, N3156, N246, N3449);
and AND3 (N3763, N3749, N2881, N1658);
buf BUF1 (N3764, N3756);
nand NAND4 (N3765, N3755, N3550, N3411, N2917);
nand NAND3 (N3766, N3764, N1136, N415);
nand NAND3 (N3767, N3754, N718, N731);
nor NOR3 (N3768, N3759, N762, N2205);
not NOT1 (N3769, N3766);
or OR4 (N3770, N3763, N259, N2744, N1451);
nor NOR2 (N3771, N3765, N1079);
xor XOR2 (N3772, N3768, N2323);
and AND3 (N3773, N3745, N3062, N985);
xor XOR2 (N3774, N3769, N2816);
not NOT1 (N3775, N3771);
nor NOR4 (N3776, N3750, N495, N2601, N1643);
not NOT1 (N3777, N3770);
and AND4 (N3778, N3762, N1499, N1986, N2691);
nand NAND3 (N3779, N3778, N324, N67);
xor XOR2 (N3780, N3761, N2900);
not NOT1 (N3781, N3779);
not NOT1 (N3782, N3767);
or OR2 (N3783, N3773, N3625);
nand NAND3 (N3784, N3780, N557, N2060);
xor XOR2 (N3785, N3777, N97);
nor NOR2 (N3786, N3783, N2946);
or OR3 (N3787, N3775, N3075, N2953);
buf BUF1 (N3788, N3781);
or OR2 (N3789, N3784, N2463);
not NOT1 (N3790, N3772);
xor XOR2 (N3791, N3757, N1266);
nor NOR4 (N3792, N3787, N1021, N2858, N2479);
xor XOR2 (N3793, N3790, N1439);
xor XOR2 (N3794, N3774, N1847);
xor XOR2 (N3795, N3776, N3327);
xor XOR2 (N3796, N3795, N1824);
nand NAND2 (N3797, N3788, N1197);
nor NOR4 (N3798, N3792, N2313, N821, N2426);
xor XOR2 (N3799, N3794, N3215);
buf BUF1 (N3800, N3786);
nand NAND3 (N3801, N3798, N1752, N1213);
nor NOR3 (N3802, N3791, N1225, N3167);
buf BUF1 (N3803, N3782);
or OR3 (N3804, N3785, N286, N1714);
nand NAND2 (N3805, N3803, N2965);
nand NAND3 (N3806, N3797, N2405, N1156);
not NOT1 (N3807, N3805);
xor XOR2 (N3808, N3793, N846);
buf BUF1 (N3809, N3800);
nand NAND4 (N3810, N3799, N621, N497, N2550);
buf BUF1 (N3811, N3809);
and AND2 (N3812, N3807, N878);
not NOT1 (N3813, N3810);
and AND4 (N3814, N3813, N3551, N1491, N1999);
and AND2 (N3815, N3801, N3140);
and AND4 (N3816, N3811, N407, N2591, N1611);
buf BUF1 (N3817, N3804);
and AND4 (N3818, N3808, N703, N2280, N1388);
not NOT1 (N3819, N3818);
and AND4 (N3820, N3812, N1969, N2522, N691);
buf BUF1 (N3821, N3820);
not NOT1 (N3822, N3802);
not NOT1 (N3823, N3814);
not NOT1 (N3824, N3821);
nand NAND3 (N3825, N3789, N415, N2237);
and AND3 (N3826, N3815, N2092, N121);
nor NOR3 (N3827, N3823, N3539, N1127);
or OR2 (N3828, N3796, N3443);
not NOT1 (N3829, N3816);
and AND2 (N3830, N3827, N3058);
buf BUF1 (N3831, N3806);
xor XOR2 (N3832, N3822, N626);
nand NAND3 (N3833, N3831, N948, N2014);
nand NAND4 (N3834, N3825, N554, N3512, N1388);
nand NAND2 (N3835, N3829, N2166);
or OR3 (N3836, N3835, N186, N46);
nand NAND2 (N3837, N3824, N252);
xor XOR2 (N3838, N3819, N1098);
not NOT1 (N3839, N3837);
or OR4 (N3840, N3834, N3062, N2629, N1172);
not NOT1 (N3841, N3817);
and AND3 (N3842, N3839, N3839, N2786);
or OR3 (N3843, N3842, N1661, N1240);
or OR4 (N3844, N3836, N3046, N3105, N528);
or OR2 (N3845, N3844, N3252);
buf BUF1 (N3846, N3833);
or OR4 (N3847, N3843, N3317, N635, N3696);
not NOT1 (N3848, N3845);
buf BUF1 (N3849, N3838);
or OR2 (N3850, N3840, N1245);
not NOT1 (N3851, N3826);
xor XOR2 (N3852, N3849, N2705);
and AND4 (N3853, N3841, N3209, N2295, N3413);
buf BUF1 (N3854, N3853);
nand NAND4 (N3855, N3846, N3042, N3333, N2608);
xor XOR2 (N3856, N3850, N2549);
nand NAND4 (N3857, N3856, N298, N1346, N1121);
nand NAND3 (N3858, N3852, N1432, N3660);
buf BUF1 (N3859, N3832);
nand NAND2 (N3860, N3847, N273);
or OR3 (N3861, N3854, N2237, N236);
and AND3 (N3862, N3860, N1667, N2280);
or OR2 (N3863, N3848, N531);
buf BUF1 (N3864, N3851);
nor NOR2 (N3865, N3858, N1205);
not NOT1 (N3866, N3862);
or OR3 (N3867, N3864, N1799, N3832);
xor XOR2 (N3868, N3859, N3761);
not NOT1 (N3869, N3830);
and AND4 (N3870, N3857, N831, N923, N2991);
xor XOR2 (N3871, N3868, N991);
nand NAND2 (N3872, N3855, N578);
nor NOR2 (N3873, N3865, N3604);
not NOT1 (N3874, N3870);
nor NOR2 (N3875, N3874, N3641);
and AND3 (N3876, N3828, N1229, N2085);
nor NOR4 (N3877, N3871, N1947, N2477, N1721);
not NOT1 (N3878, N3861);
not NOT1 (N3879, N3867);
not NOT1 (N3880, N3875);
buf BUF1 (N3881, N3872);
or OR2 (N3882, N3869, N2503);
buf BUF1 (N3883, N3881);
not NOT1 (N3884, N3876);
nor NOR4 (N3885, N3866, N1485, N2986, N577);
not NOT1 (N3886, N3884);
nor NOR4 (N3887, N3877, N896, N1515, N542);
and AND2 (N3888, N3883, N65);
and AND2 (N3889, N3878, N988);
nand NAND2 (N3890, N3873, N671);
xor XOR2 (N3891, N3882, N1648);
xor XOR2 (N3892, N3863, N1332);
nand NAND4 (N3893, N3889, N972, N2803, N3146);
buf BUF1 (N3894, N3888);
xor XOR2 (N3895, N3885, N2310);
nor NOR3 (N3896, N3894, N724, N2432);
buf BUF1 (N3897, N3896);
buf BUF1 (N3898, N3880);
or OR3 (N3899, N3897, N1666, N1104);
buf BUF1 (N3900, N3886);
nand NAND3 (N3901, N3890, N1746, N3806);
xor XOR2 (N3902, N3879, N2989);
and AND3 (N3903, N3892, N3527, N437);
buf BUF1 (N3904, N3898);
not NOT1 (N3905, N3893);
nand NAND4 (N3906, N3901, N3597, N3614, N2447);
or OR2 (N3907, N3887, N2586);
nor NOR2 (N3908, N3895, N1520);
not NOT1 (N3909, N3902);
nor NOR2 (N3910, N3906, N1735);
xor XOR2 (N3911, N3909, N2647);
xor XOR2 (N3912, N3905, N2240);
nand NAND2 (N3913, N3912, N3456);
nor NOR2 (N3914, N3907, N695);
not NOT1 (N3915, N3910);
nand NAND2 (N3916, N3911, N2750);
buf BUF1 (N3917, N3891);
buf BUF1 (N3918, N3903);
not NOT1 (N3919, N3899);
nand NAND4 (N3920, N3908, N3311, N3747, N628);
nand NAND2 (N3921, N3919, N1605);
nor NOR4 (N3922, N3900, N1268, N3840, N3075);
nand NAND2 (N3923, N3915, N1648);
nand NAND3 (N3924, N3917, N734, N265);
not NOT1 (N3925, N3921);
xor XOR2 (N3926, N3918, N2494);
nor NOR2 (N3927, N3924, N356);
or OR2 (N3928, N3925, N2926);
and AND3 (N3929, N3928, N561, N3863);
nand NAND4 (N3930, N3913, N1848, N3304, N727);
nor NOR4 (N3931, N3916, N3290, N1965, N1910);
nor NOR4 (N3932, N3914, N3244, N1512, N3183);
and AND3 (N3933, N3930, N71, N2952);
not NOT1 (N3934, N3926);
buf BUF1 (N3935, N3929);
and AND4 (N3936, N3922, N2827, N2289, N3905);
not NOT1 (N3937, N3936);
nor NOR4 (N3938, N3933, N91, N3655, N2583);
nand NAND3 (N3939, N3931, N3272, N640);
buf BUF1 (N3940, N3934);
not NOT1 (N3941, N3937);
and AND4 (N3942, N3941, N1321, N1114, N1724);
and AND3 (N3943, N3939, N781, N457);
and AND4 (N3944, N3923, N1578, N1419, N532);
and AND2 (N3945, N3927, N995);
xor XOR2 (N3946, N3940, N3427);
and AND4 (N3947, N3932, N71, N1380, N1462);
not NOT1 (N3948, N3920);
not NOT1 (N3949, N3943);
or OR3 (N3950, N3935, N3217, N3359);
or OR3 (N3951, N3944, N2848, N1966);
xor XOR2 (N3952, N3951, N113);
xor XOR2 (N3953, N3938, N1762);
buf BUF1 (N3954, N3904);
not NOT1 (N3955, N3947);
or OR3 (N3956, N3945, N780, N3057);
and AND2 (N3957, N3949, N1860);
or OR2 (N3958, N3946, N3155);
and AND3 (N3959, N3950, N47, N1356);
not NOT1 (N3960, N3955);
xor XOR2 (N3961, N3960, N1504);
nor NOR3 (N3962, N3953, N1548, N3817);
buf BUF1 (N3963, N3958);
or OR4 (N3964, N3948, N933, N1086, N3961);
not NOT1 (N3965, N2246);
and AND2 (N3966, N3965, N2910);
nand NAND3 (N3967, N3952, N22, N505);
xor XOR2 (N3968, N3942, N1458);
or OR3 (N3969, N3963, N2917, N1335);
not NOT1 (N3970, N3969);
nor NOR2 (N3971, N3957, N1333);
and AND3 (N3972, N3968, N1813, N1892);
or OR4 (N3973, N3962, N1325, N3142, N1553);
and AND4 (N3974, N3964, N2597, N1586, N2793);
xor XOR2 (N3975, N3966, N2534);
nor NOR4 (N3976, N3971, N296, N1314, N1788);
xor XOR2 (N3977, N3954, N711);
not NOT1 (N3978, N3977);
buf BUF1 (N3979, N3975);
xor XOR2 (N3980, N3972, N3252);
or OR3 (N3981, N3980, N3688, N1870);
nand NAND3 (N3982, N3981, N3456, N742);
and AND4 (N3983, N3979, N1621, N221, N51);
nor NOR2 (N3984, N3974, N720);
nor NOR4 (N3985, N3973, N808, N1651, N2142);
not NOT1 (N3986, N3982);
or OR2 (N3987, N3970, N1470);
or OR2 (N3988, N3986, N3689);
nand NAND3 (N3989, N3987, N1378, N2276);
and AND4 (N3990, N3983, N2064, N1522, N709);
xor XOR2 (N3991, N3990, N2519);
nor NOR2 (N3992, N3988, N2771);
nor NOR2 (N3993, N3989, N1577);
buf BUF1 (N3994, N3993);
nand NAND3 (N3995, N3976, N1990, N86);
nor NOR2 (N3996, N3984, N343);
not NOT1 (N3997, N3994);
nor NOR4 (N3998, N3996, N79, N983, N1054);
xor XOR2 (N3999, N3992, N1580);
nor NOR3 (N4000, N3959, N2483, N3928);
buf BUF1 (N4001, N3967);
xor XOR2 (N4002, N3978, N963);
or OR2 (N4003, N3998, N227);
not NOT1 (N4004, N4000);
nor NOR2 (N4005, N4004, N1533);
and AND4 (N4006, N3956, N908, N1169, N2120);
not NOT1 (N4007, N3997);
nor NOR3 (N4008, N3999, N2008, N1747);
or OR4 (N4009, N4003, N2341, N3069, N3658);
xor XOR2 (N4010, N3995, N1605);
nor NOR4 (N4011, N3991, N1256, N707, N780);
endmodule