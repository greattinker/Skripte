// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11;

output N595,N607,N602,N609,N603,N610,N605,N608,N593,N611;

nor NOR4 (N12, N2, N1, N6, N7);
nor NOR4 (N13, N6, N4, N2, N5);
not NOT1 (N14, N2);
or OR4 (N15, N12, N11, N2, N13);
buf BUF1 (N16, N12);
nor NOR2 (N17, N1, N12);
or OR2 (N18, N11, N16);
or OR2 (N19, N9, N3);
nor NOR2 (N20, N10, N3);
not NOT1 (N21, N4);
nand NAND3 (N22, N1, N18, N2);
not NOT1 (N23, N17);
and AND3 (N24, N8, N16, N2);
or OR3 (N25, N21, N23, N10);
and AND2 (N26, N11, N5);
and AND2 (N27, N23, N13);
buf BUF1 (N28, N23);
xor XOR2 (N29, N24, N7);
not NOT1 (N30, N15);
or OR4 (N31, N29, N17, N23, N14);
nand NAND2 (N32, N3, N12);
nand NAND2 (N33, N20, N26);
and AND4 (N34, N3, N23, N16, N21);
buf BUF1 (N35, N32);
or OR2 (N36, N27, N35);
buf BUF1 (N37, N31);
nor NOR3 (N38, N37, N4, N20);
nand NAND3 (N39, N38, N29, N9);
buf BUF1 (N40, N5);
and AND3 (N41, N40, N6, N39);
and AND4 (N42, N1, N1, N20, N19);
not NOT1 (N43, N12);
and AND3 (N44, N36, N40, N7);
xor XOR2 (N45, N30, N12);
or OR3 (N46, N34, N34, N38);
and AND2 (N47, N43, N26);
nor NOR3 (N48, N33, N28, N10);
or OR2 (N49, N42, N13);
and AND3 (N50, N6, N41, N41);
xor XOR2 (N51, N12, N48);
nand NAND3 (N52, N12, N11, N27);
not NOT1 (N53, N47);
nor NOR4 (N54, N45, N36, N4, N20);
and AND2 (N55, N25, N34);
buf BUF1 (N56, N46);
or OR2 (N57, N44, N25);
nand NAND4 (N58, N57, N44, N45, N15);
and AND4 (N59, N52, N58, N35, N40);
and AND4 (N60, N42, N17, N50, N21);
and AND4 (N61, N29, N30, N46, N17);
and AND2 (N62, N59, N4);
nand NAND4 (N63, N55, N61, N23, N57);
nand NAND2 (N64, N4, N61);
buf BUF1 (N65, N63);
buf BUF1 (N66, N53);
nor NOR4 (N67, N62, N23, N9, N33);
buf BUF1 (N68, N54);
xor XOR2 (N69, N60, N30);
xor XOR2 (N70, N22, N39);
nand NAND4 (N71, N49, N35, N26, N20);
xor XOR2 (N72, N64, N41);
buf BUF1 (N73, N70);
or OR3 (N74, N66, N71, N40);
nand NAND4 (N75, N15, N6, N13, N29);
buf BUF1 (N76, N65);
buf BUF1 (N77, N51);
or OR3 (N78, N69, N27, N28);
xor XOR2 (N79, N76, N74);
nand NAND4 (N80, N23, N65, N62, N75);
buf BUF1 (N81, N61);
buf BUF1 (N82, N77);
or OR2 (N83, N67, N22);
nand NAND2 (N84, N83, N8);
nor NOR4 (N85, N73, N18, N24, N9);
nand NAND3 (N86, N79, N80, N38);
buf BUF1 (N87, N31);
and AND2 (N88, N82, N73);
and AND3 (N89, N85, N21, N22);
or OR3 (N90, N86, N70, N77);
nand NAND2 (N91, N78, N27);
not NOT1 (N92, N72);
or OR4 (N93, N87, N65, N92, N1);
nand NAND3 (N94, N23, N41, N9);
xor XOR2 (N95, N90, N32);
and AND2 (N96, N88, N44);
and AND3 (N97, N84, N91, N95);
xor XOR2 (N98, N3, N81);
nand NAND3 (N99, N22, N58, N1);
not NOT1 (N100, N51);
xor XOR2 (N101, N93, N44);
or OR4 (N102, N94, N74, N73, N85);
or OR4 (N103, N101, N8, N75, N23);
not NOT1 (N104, N89);
xor XOR2 (N105, N97, N79);
nor NOR2 (N106, N103, N62);
nor NOR3 (N107, N102, N84, N47);
buf BUF1 (N108, N104);
nor NOR4 (N109, N99, N33, N64, N65);
or OR3 (N110, N100, N68, N27);
and AND3 (N111, N35, N22, N18);
not NOT1 (N112, N105);
nand NAND3 (N113, N110, N33, N94);
nand NAND2 (N114, N111, N65);
or OR4 (N115, N113, N112, N37, N90);
nand NAND3 (N116, N55, N95, N81);
nand NAND3 (N117, N106, N55, N17);
or OR4 (N118, N108, N27, N99, N101);
buf BUF1 (N119, N114);
xor XOR2 (N120, N109, N91);
buf BUF1 (N121, N116);
nand NAND4 (N122, N120, N34, N115, N116);
and AND2 (N123, N45, N121);
nand NAND3 (N124, N49, N20, N20);
not NOT1 (N125, N124);
not NOT1 (N126, N98);
not NOT1 (N127, N117);
nor NOR3 (N128, N122, N30, N66);
not NOT1 (N129, N123);
not NOT1 (N130, N56);
nand NAND3 (N131, N96, N10, N29);
nor NOR2 (N132, N129, N130);
not NOT1 (N133, N48);
not NOT1 (N134, N128);
and AND3 (N135, N125, N59, N133);
nand NAND2 (N136, N63, N9);
not NOT1 (N137, N126);
not NOT1 (N138, N136);
xor XOR2 (N139, N134, N85);
buf BUF1 (N140, N138);
nand NAND2 (N141, N135, N125);
buf BUF1 (N142, N118);
or OR3 (N143, N131, N64, N85);
and AND2 (N144, N127, N127);
nor NOR3 (N145, N137, N21, N56);
nor NOR2 (N146, N143, N96);
nand NAND4 (N147, N146, N72, N79, N137);
and AND4 (N148, N144, N115, N25, N28);
buf BUF1 (N149, N141);
xor XOR2 (N150, N119, N2);
and AND4 (N151, N148, N3, N104, N96);
xor XOR2 (N152, N142, N76);
not NOT1 (N153, N151);
or OR4 (N154, N132, N132, N141, N97);
nor NOR3 (N155, N150, N45, N1);
or OR3 (N156, N149, N123, N105);
and AND3 (N157, N147, N29, N10);
or OR2 (N158, N152, N86);
nor NOR3 (N159, N107, N130, N48);
nand NAND4 (N160, N156, N72, N99, N157);
or OR3 (N161, N8, N72, N55);
not NOT1 (N162, N158);
buf BUF1 (N163, N145);
nand NAND2 (N164, N155, N65);
xor XOR2 (N165, N159, N10);
buf BUF1 (N166, N165);
or OR4 (N167, N140, N26, N136, N97);
nor NOR4 (N168, N160, N18, N87, N138);
buf BUF1 (N169, N154);
nor NOR2 (N170, N167, N156);
and AND2 (N171, N166, N93);
or OR4 (N172, N168, N84, N17, N169);
buf BUF1 (N173, N165);
xor XOR2 (N174, N164, N61);
xor XOR2 (N175, N171, N2);
not NOT1 (N176, N139);
and AND4 (N177, N174, N25, N28, N17);
or OR4 (N178, N173, N15, N30, N97);
buf BUF1 (N179, N162);
nand NAND2 (N180, N163, N155);
or OR4 (N181, N177, N81, N157, N33);
buf BUF1 (N182, N161);
not NOT1 (N183, N182);
nand NAND2 (N184, N172, N51);
nand NAND4 (N185, N181, N35, N82, N56);
nor NOR2 (N186, N184, N130);
and AND3 (N187, N175, N85, N105);
nor NOR4 (N188, N176, N98, N181, N60);
buf BUF1 (N189, N153);
buf BUF1 (N190, N179);
not NOT1 (N191, N170);
or OR2 (N192, N180, N12);
nand NAND2 (N193, N189, N117);
buf BUF1 (N194, N183);
nor NOR4 (N195, N178, N117, N168, N31);
nor NOR4 (N196, N188, N128, N161, N195);
not NOT1 (N197, N2);
xor XOR2 (N198, N192, N53);
nor NOR3 (N199, N198, N65, N148);
and AND4 (N200, N190, N32, N13, N32);
not NOT1 (N201, N185);
nor NOR3 (N202, N193, N13, N26);
not NOT1 (N203, N196);
nand NAND4 (N204, N202, N159, N65, N59);
nor NOR3 (N205, N191, N131, N73);
and AND2 (N206, N186, N12);
xor XOR2 (N207, N199, N118);
nand NAND2 (N208, N205, N53);
and AND2 (N209, N207, N197);
not NOT1 (N210, N71);
nand NAND2 (N211, N209, N177);
nor NOR2 (N212, N206, N168);
and AND4 (N213, N194, N140, N119, N136);
buf BUF1 (N214, N201);
not NOT1 (N215, N203);
xor XOR2 (N216, N213, N119);
nand NAND3 (N217, N210, N186, N197);
nor NOR3 (N218, N216, N70, N80);
xor XOR2 (N219, N200, N77);
buf BUF1 (N220, N217);
xor XOR2 (N221, N218, N19);
and AND4 (N222, N220, N157, N107, N127);
or OR4 (N223, N219, N44, N195, N115);
and AND3 (N224, N215, N43, N174);
or OR3 (N225, N214, N198, N74);
or OR4 (N226, N224, N211, N40, N211);
nor NOR4 (N227, N156, N126, N25, N192);
xor XOR2 (N228, N221, N124);
nor NOR3 (N229, N187, N78, N195);
or OR3 (N230, N204, N119, N95);
buf BUF1 (N231, N228);
buf BUF1 (N232, N222);
and AND2 (N233, N225, N40);
and AND3 (N234, N229, N39, N199);
buf BUF1 (N235, N234);
nand NAND3 (N236, N232, N118, N86);
nor NOR3 (N237, N227, N202, N19);
and AND3 (N238, N208, N54, N171);
xor XOR2 (N239, N236, N93);
not NOT1 (N240, N238);
nor NOR4 (N241, N226, N6, N41, N151);
and AND2 (N242, N239, N64);
or OR4 (N243, N233, N14, N52, N191);
nor NOR2 (N244, N230, N24);
not NOT1 (N245, N244);
and AND4 (N246, N223, N192, N36, N12);
nor NOR4 (N247, N242, N174, N69, N126);
not NOT1 (N248, N246);
or OR3 (N249, N235, N184, N222);
or OR3 (N250, N249, N53, N11);
nor NOR3 (N251, N250, N167, N121);
buf BUF1 (N252, N241);
nor NOR4 (N253, N247, N127, N250, N18);
xor XOR2 (N254, N251, N204);
and AND3 (N255, N243, N13, N29);
and AND4 (N256, N245, N243, N172, N128);
not NOT1 (N257, N212);
xor XOR2 (N258, N252, N231);
not NOT1 (N259, N154);
not NOT1 (N260, N254);
xor XOR2 (N261, N255, N85);
and AND4 (N262, N237, N192, N129, N223);
xor XOR2 (N263, N253, N244);
nor NOR3 (N264, N262, N103, N71);
and AND2 (N265, N261, N48);
nand NAND2 (N266, N248, N139);
or OR4 (N267, N260, N14, N113, N246);
xor XOR2 (N268, N264, N44);
or OR2 (N269, N263, N255);
or OR2 (N270, N265, N90);
buf BUF1 (N271, N258);
buf BUF1 (N272, N271);
xor XOR2 (N273, N257, N217);
nand NAND2 (N274, N266, N116);
nor NOR3 (N275, N259, N67, N158);
buf BUF1 (N276, N275);
nor NOR2 (N277, N274, N99);
nor NOR4 (N278, N240, N238, N52, N63);
nor NOR3 (N279, N267, N167, N50);
or OR4 (N280, N272, N272, N129, N262);
xor XOR2 (N281, N268, N58);
nor NOR2 (N282, N256, N230);
or OR2 (N283, N280, N147);
nand NAND2 (N284, N270, N267);
and AND4 (N285, N278, N186, N45, N159);
not NOT1 (N286, N273);
nor NOR3 (N287, N286, N39, N261);
buf BUF1 (N288, N269);
xor XOR2 (N289, N288, N19);
and AND3 (N290, N279, N170, N278);
and AND2 (N291, N276, N18);
not NOT1 (N292, N283);
nor NOR4 (N293, N285, N124, N93, N283);
and AND2 (N294, N277, N11);
and AND4 (N295, N292, N52, N31, N40);
nand NAND2 (N296, N291, N128);
xor XOR2 (N297, N296, N188);
buf BUF1 (N298, N287);
not NOT1 (N299, N282);
nand NAND3 (N300, N281, N39, N49);
xor XOR2 (N301, N289, N32);
buf BUF1 (N302, N300);
buf BUF1 (N303, N293);
buf BUF1 (N304, N299);
buf BUF1 (N305, N284);
buf BUF1 (N306, N297);
not NOT1 (N307, N303);
buf BUF1 (N308, N295);
xor XOR2 (N309, N290, N95);
buf BUF1 (N310, N298);
nand NAND2 (N311, N308, N67);
xor XOR2 (N312, N311, N309);
or OR2 (N313, N210, N46);
xor XOR2 (N314, N312, N99);
and AND3 (N315, N302, N140, N260);
nand NAND4 (N316, N314, N120, N18, N309);
nor NOR2 (N317, N294, N149);
and AND3 (N318, N305, N26, N19);
nand NAND3 (N319, N313, N301, N174);
buf BUF1 (N320, N153);
nand NAND2 (N321, N317, N135);
or OR3 (N322, N310, N202, N25);
not NOT1 (N323, N306);
buf BUF1 (N324, N316);
not NOT1 (N325, N319);
xor XOR2 (N326, N324, N260);
or OR4 (N327, N326, N130, N38, N16);
xor XOR2 (N328, N321, N230);
or OR2 (N329, N325, N170);
and AND3 (N330, N322, N160, N164);
nand NAND3 (N331, N315, N6, N234);
nor NOR3 (N332, N328, N60, N83);
nand NAND3 (N333, N332, N30, N311);
and AND4 (N334, N304, N39, N43, N146);
nor NOR3 (N335, N323, N26, N201);
or OR2 (N336, N329, N308);
nor NOR4 (N337, N335, N326, N165, N88);
not NOT1 (N338, N336);
not NOT1 (N339, N334);
nor NOR3 (N340, N333, N287, N99);
xor XOR2 (N341, N339, N186);
xor XOR2 (N342, N331, N261);
nor NOR2 (N343, N307, N43);
or OR4 (N344, N343, N204, N240, N49);
nand NAND2 (N345, N320, N237);
nand NAND3 (N346, N342, N59, N274);
not NOT1 (N347, N338);
or OR2 (N348, N337, N108);
xor XOR2 (N349, N341, N111);
and AND2 (N350, N344, N1);
and AND2 (N351, N327, N325);
not NOT1 (N352, N350);
and AND4 (N353, N346, N49, N89, N87);
xor XOR2 (N354, N340, N154);
not NOT1 (N355, N330);
nand NAND2 (N356, N354, N145);
not NOT1 (N357, N349);
and AND2 (N358, N318, N313);
nor NOR2 (N359, N355, N57);
nand NAND4 (N360, N345, N221, N9, N14);
not NOT1 (N361, N359);
nor NOR4 (N362, N353, N43, N359, N77);
buf BUF1 (N363, N348);
and AND3 (N364, N352, N343, N80);
nand NAND3 (N365, N362, N110, N318);
or OR2 (N366, N360, N29);
xor XOR2 (N367, N363, N114);
or OR3 (N368, N364, N90, N330);
buf BUF1 (N369, N351);
and AND4 (N370, N367, N51, N309, N226);
nor NOR4 (N371, N356, N318, N302, N359);
and AND4 (N372, N365, N119, N117, N157);
not NOT1 (N373, N366);
or OR4 (N374, N357, N68, N215, N57);
and AND3 (N375, N374, N213, N282);
buf BUF1 (N376, N369);
not NOT1 (N377, N371);
and AND3 (N378, N361, N123, N347);
or OR2 (N379, N108, N284);
xor XOR2 (N380, N372, N332);
not NOT1 (N381, N375);
xor XOR2 (N382, N373, N56);
or OR3 (N383, N358, N376, N9);
buf BUF1 (N384, N207);
not NOT1 (N385, N383);
buf BUF1 (N386, N381);
nand NAND3 (N387, N370, N349, N324);
nand NAND2 (N388, N377, N243);
buf BUF1 (N389, N380);
or OR3 (N390, N382, N295, N13);
or OR3 (N391, N387, N32, N99);
buf BUF1 (N392, N390);
or OR4 (N393, N386, N277, N40, N115);
xor XOR2 (N394, N389, N193);
nand NAND4 (N395, N394, N217, N323, N343);
or OR3 (N396, N395, N342, N338);
not NOT1 (N397, N388);
or OR4 (N398, N378, N336, N187, N62);
nand NAND2 (N399, N397, N146);
or OR2 (N400, N385, N372);
nand NAND4 (N401, N398, N301, N123, N384);
buf BUF1 (N402, N224);
nand NAND4 (N403, N400, N298, N223, N82);
nand NAND4 (N404, N379, N345, N284, N63);
and AND2 (N405, N402, N196);
not NOT1 (N406, N368);
and AND2 (N407, N396, N229);
nor NOR2 (N408, N393, N287);
or OR3 (N409, N407, N122, N72);
buf BUF1 (N410, N409);
or OR3 (N411, N403, N343, N238);
or OR4 (N412, N408, N305, N335, N298);
buf BUF1 (N413, N401);
or OR2 (N414, N404, N108);
nor NOR2 (N415, N410, N1);
and AND4 (N416, N406, N409, N331, N87);
and AND3 (N417, N413, N4, N77);
xor XOR2 (N418, N392, N170);
xor XOR2 (N419, N414, N418);
and AND3 (N420, N192, N120, N51);
buf BUF1 (N421, N419);
not NOT1 (N422, N416);
xor XOR2 (N423, N421, N412);
buf BUF1 (N424, N223);
buf BUF1 (N425, N424);
buf BUF1 (N426, N411);
or OR3 (N427, N425, N413, N106);
buf BUF1 (N428, N415);
nand NAND3 (N429, N417, N391, N29);
buf BUF1 (N430, N375);
buf BUF1 (N431, N405);
nor NOR4 (N432, N427, N70, N353, N168);
nor NOR3 (N433, N429, N380, N339);
or OR4 (N434, N432, N44, N330, N284);
nand NAND2 (N435, N434, N108);
buf BUF1 (N436, N433);
xor XOR2 (N437, N431, N332);
xor XOR2 (N438, N428, N375);
or OR3 (N439, N438, N35, N424);
and AND4 (N440, N430, N396, N84, N406);
not NOT1 (N441, N426);
nand NAND2 (N442, N420, N411);
buf BUF1 (N443, N423);
nor NOR4 (N444, N436, N397, N276, N132);
nor NOR4 (N445, N440, N39, N306, N136);
nand NAND4 (N446, N439, N208, N400, N345);
nand NAND4 (N447, N441, N144, N161, N190);
xor XOR2 (N448, N443, N225);
nand NAND4 (N449, N448, N43, N259, N109);
not NOT1 (N450, N437);
or OR2 (N451, N447, N130);
xor XOR2 (N452, N435, N38);
and AND2 (N453, N422, N34);
buf BUF1 (N454, N450);
and AND2 (N455, N449, N177);
or OR2 (N456, N445, N252);
and AND4 (N457, N452, N179, N60, N165);
xor XOR2 (N458, N453, N87);
or OR3 (N459, N456, N6, N175);
nand NAND4 (N460, N459, N120, N385, N349);
buf BUF1 (N461, N458);
buf BUF1 (N462, N399);
nor NOR2 (N463, N446, N88);
nand NAND4 (N464, N460, N413, N72, N188);
not NOT1 (N465, N461);
not NOT1 (N466, N444);
and AND4 (N467, N466, N183, N287, N208);
and AND4 (N468, N451, N159, N461, N395);
and AND3 (N469, N442, N458, N427);
nand NAND2 (N470, N465, N205);
buf BUF1 (N471, N455);
xor XOR2 (N472, N463, N12);
buf BUF1 (N473, N464);
nand NAND4 (N474, N468, N70, N147, N118);
nand NAND2 (N475, N474, N292);
and AND2 (N476, N472, N332);
or OR4 (N477, N467, N157, N224, N414);
nand NAND2 (N478, N469, N138);
not NOT1 (N479, N473);
and AND4 (N480, N462, N257, N96, N108);
buf BUF1 (N481, N475);
nor NOR4 (N482, N478, N137, N65, N443);
buf BUF1 (N483, N470);
or OR2 (N484, N457, N82);
nor NOR3 (N485, N471, N105, N127);
nand NAND4 (N486, N484, N150, N363, N364);
or OR4 (N487, N479, N58, N380, N126);
not NOT1 (N488, N482);
or OR4 (N489, N488, N144, N342, N322);
and AND3 (N490, N481, N45, N49);
buf BUF1 (N491, N454);
nor NOR3 (N492, N490, N476, N134);
or OR4 (N493, N262, N59, N334, N348);
nand NAND2 (N494, N493, N59);
and AND3 (N495, N477, N221, N1);
buf BUF1 (N496, N483);
buf BUF1 (N497, N485);
xor XOR2 (N498, N496, N230);
buf BUF1 (N499, N492);
buf BUF1 (N500, N487);
nor NOR2 (N501, N499, N49);
xor XOR2 (N502, N486, N227);
nand NAND3 (N503, N495, N159, N191);
nand NAND4 (N504, N502, N449, N284, N303);
not NOT1 (N505, N501);
nor NOR3 (N506, N494, N112, N52);
xor XOR2 (N507, N491, N492);
nor NOR4 (N508, N504, N189, N31, N462);
or OR4 (N509, N489, N188, N288, N444);
nand NAND3 (N510, N498, N18, N363);
and AND3 (N511, N510, N33, N358);
buf BUF1 (N512, N508);
not NOT1 (N513, N509);
not NOT1 (N514, N506);
and AND4 (N515, N500, N405, N326, N437);
and AND4 (N516, N503, N82, N24, N296);
not NOT1 (N517, N515);
xor XOR2 (N518, N516, N429);
nand NAND2 (N519, N517, N479);
or OR4 (N520, N514, N316, N110, N342);
nand NAND4 (N521, N505, N104, N437, N493);
xor XOR2 (N522, N513, N478);
or OR2 (N523, N520, N94);
nand NAND4 (N524, N519, N77, N391, N140);
nand NAND2 (N525, N507, N162);
and AND4 (N526, N518, N160, N256, N3);
nand NAND4 (N527, N526, N141, N254, N407);
buf BUF1 (N528, N497);
not NOT1 (N529, N523);
not NOT1 (N530, N511);
not NOT1 (N531, N528);
buf BUF1 (N532, N512);
xor XOR2 (N533, N480, N453);
not NOT1 (N534, N525);
nand NAND2 (N535, N533, N264);
nand NAND2 (N536, N529, N298);
xor XOR2 (N537, N532, N199);
and AND2 (N538, N527, N471);
or OR3 (N539, N536, N496, N153);
not NOT1 (N540, N531);
xor XOR2 (N541, N540, N344);
buf BUF1 (N542, N530);
or OR2 (N543, N541, N291);
xor XOR2 (N544, N534, N415);
buf BUF1 (N545, N537);
nor NOR3 (N546, N538, N285, N59);
xor XOR2 (N547, N524, N199);
and AND2 (N548, N542, N133);
or OR2 (N549, N535, N132);
or OR2 (N550, N539, N497);
nor NOR2 (N551, N549, N300);
nand NAND2 (N552, N548, N477);
nor NOR3 (N553, N545, N248, N416);
or OR3 (N554, N522, N117, N145);
or OR3 (N555, N553, N231, N539);
xor XOR2 (N556, N552, N246);
xor XOR2 (N557, N551, N37);
and AND4 (N558, N554, N249, N145, N72);
nor NOR4 (N559, N547, N251, N131, N481);
nand NAND4 (N560, N543, N84, N299, N336);
buf BUF1 (N561, N558);
nand NAND3 (N562, N559, N305, N268);
nand NAND2 (N563, N546, N214);
buf BUF1 (N564, N556);
not NOT1 (N565, N555);
nor NOR2 (N566, N565, N504);
and AND2 (N567, N566, N529);
not NOT1 (N568, N564);
not NOT1 (N569, N562);
nand NAND2 (N570, N550, N424);
nand NAND2 (N571, N561, N16);
xor XOR2 (N572, N557, N521);
xor XOR2 (N573, N518, N274);
nor NOR4 (N574, N560, N293, N494, N269);
and AND3 (N575, N567, N124, N43);
and AND2 (N576, N572, N307);
xor XOR2 (N577, N575, N47);
nor NOR4 (N578, N544, N500, N19, N126);
or OR2 (N579, N571, N428);
and AND4 (N580, N573, N393, N455, N317);
nand NAND3 (N581, N577, N52, N191);
nor NOR3 (N582, N574, N170, N230);
nor NOR4 (N583, N578, N399, N106, N375);
not NOT1 (N584, N576);
nand NAND2 (N585, N563, N352);
or OR3 (N586, N584, N334, N401);
nor NOR4 (N587, N579, N264, N220, N467);
xor XOR2 (N588, N581, N23);
buf BUF1 (N589, N585);
nand NAND2 (N590, N568, N367);
or OR2 (N591, N582, N233);
nand NAND3 (N592, N587, N311, N84);
nor NOR3 (N593, N570, N63, N364);
or OR3 (N594, N583, N423, N142);
xor XOR2 (N595, N588, N75);
nor NOR2 (N596, N580, N448);
buf BUF1 (N597, N569);
and AND3 (N598, N596, N180, N171);
nand NAND2 (N599, N597, N322);
and AND3 (N600, N589, N221, N397);
or OR3 (N601, N600, N206, N344);
not NOT1 (N602, N591);
not NOT1 (N603, N594);
nor NOR3 (N604, N601, N581, N528);
not NOT1 (N605, N599);
buf BUF1 (N606, N598);
nor NOR2 (N607, N606, N463);
buf BUF1 (N608, N590);
buf BUF1 (N609, N586);
and AND2 (N610, N592, N36);
and AND2 (N611, N604, N132);
endmodule