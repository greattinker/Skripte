// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23;

output N512,N522,N521,N503,N506,N519,N520,N511,N509,N523;

xor XOR2 (N24, N14, N11);
nand NAND4 (N25, N16, N8, N19, N19);
nor NOR3 (N26, N18, N25, N15);
buf BUF1 (N27, N16);
or OR4 (N28, N23, N12, N4, N17);
nand NAND3 (N29, N23, N19, N28);
not NOT1 (N30, N13);
xor XOR2 (N31, N22, N21);
and AND2 (N32, N25, N6);
buf BUF1 (N33, N31);
or OR2 (N34, N18, N30);
nand NAND4 (N35, N26, N9, N21, N18);
nor NOR2 (N36, N5, N1);
not NOT1 (N37, N16);
or OR2 (N38, N17, N9);
nand NAND3 (N39, N36, N35, N37);
not NOT1 (N40, N13);
or OR2 (N41, N13, N2);
buf BUF1 (N42, N29);
nand NAND4 (N43, N24, N25, N28, N10);
not NOT1 (N44, N41);
or OR2 (N45, N34, N31);
nor NOR2 (N46, N39, N30);
nand NAND3 (N47, N38, N42, N4);
xor XOR2 (N48, N6, N21);
not NOT1 (N49, N43);
or OR2 (N50, N32, N4);
nand NAND3 (N51, N49, N9, N6);
nor NOR4 (N52, N48, N15, N16, N44);
or OR3 (N53, N31, N43, N34);
nor NOR4 (N54, N45, N40, N31, N14);
nor NOR2 (N55, N23, N48);
or OR3 (N56, N50, N36, N45);
nand NAND3 (N57, N54, N50, N43);
not NOT1 (N58, N47);
and AND3 (N59, N55, N17, N50);
or OR3 (N60, N33, N47, N3);
not NOT1 (N61, N60);
and AND2 (N62, N52, N38);
not NOT1 (N63, N59);
and AND2 (N64, N56, N29);
and AND3 (N65, N51, N48, N3);
not NOT1 (N66, N57);
and AND2 (N67, N46, N20);
and AND4 (N68, N27, N28, N50, N59);
and AND2 (N69, N53, N35);
not NOT1 (N70, N68);
buf BUF1 (N71, N65);
not NOT1 (N72, N64);
xor XOR2 (N73, N67, N19);
nor NOR4 (N74, N66, N53, N26, N7);
buf BUF1 (N75, N71);
buf BUF1 (N76, N69);
nor NOR4 (N77, N63, N3, N29, N57);
or OR2 (N78, N75, N31);
not NOT1 (N79, N77);
nor NOR2 (N80, N74, N2);
xor XOR2 (N81, N80, N73);
nand NAND2 (N82, N44, N3);
xor XOR2 (N83, N61, N42);
nand NAND2 (N84, N79, N69);
nor NOR4 (N85, N58, N33, N84, N4);
nand NAND3 (N86, N84, N9, N52);
not NOT1 (N87, N78);
and AND2 (N88, N76, N79);
and AND3 (N89, N86, N26, N39);
not NOT1 (N90, N87);
or OR2 (N91, N70, N64);
nand NAND4 (N92, N82, N77, N78, N13);
nor NOR4 (N93, N90, N9, N3, N3);
xor XOR2 (N94, N93, N6);
nand NAND2 (N95, N89, N64);
nor NOR3 (N96, N85, N5, N9);
xor XOR2 (N97, N91, N67);
buf BUF1 (N98, N72);
or OR3 (N99, N92, N9, N37);
xor XOR2 (N100, N94, N54);
nor NOR2 (N101, N62, N87);
buf BUF1 (N102, N95);
xor XOR2 (N103, N83, N53);
nor NOR4 (N104, N102, N81, N97, N78);
xor XOR2 (N105, N18, N76);
not NOT1 (N106, N87);
not NOT1 (N107, N104);
and AND2 (N108, N99, N22);
xor XOR2 (N109, N96, N64);
and AND2 (N110, N100, N76);
or OR2 (N111, N106, N96);
xor XOR2 (N112, N111, N97);
nor NOR2 (N113, N109, N13);
buf BUF1 (N114, N103);
buf BUF1 (N115, N114);
not NOT1 (N116, N115);
nand NAND3 (N117, N107, N29, N13);
nand NAND2 (N118, N117, N2);
nor NOR4 (N119, N113, N10, N41, N104);
nor NOR4 (N120, N119, N72, N63, N56);
nand NAND4 (N121, N101, N39, N79, N39);
or OR2 (N122, N108, N60);
buf BUF1 (N123, N116);
or OR2 (N124, N88, N96);
or OR4 (N125, N123, N74, N29, N100);
nor NOR3 (N126, N121, N61, N33);
or OR3 (N127, N110, N95, N117);
not NOT1 (N128, N112);
nor NOR3 (N129, N125, N60, N5);
buf BUF1 (N130, N98);
nand NAND3 (N131, N128, N80, N61);
buf BUF1 (N132, N122);
nor NOR4 (N133, N126, N11, N127, N74);
nand NAND3 (N134, N113, N4, N130);
xor XOR2 (N135, N90, N102);
buf BUF1 (N136, N129);
nand NAND2 (N137, N134, N31);
nor NOR2 (N138, N132, N134);
buf BUF1 (N139, N120);
buf BUF1 (N140, N133);
not NOT1 (N141, N118);
nand NAND3 (N142, N141, N78, N9);
and AND3 (N143, N139, N92, N5);
or OR3 (N144, N105, N97, N113);
nor NOR4 (N145, N131, N41, N114, N37);
nor NOR4 (N146, N142, N92, N102, N67);
and AND2 (N147, N145, N131);
or OR3 (N148, N138, N64, N13);
buf BUF1 (N149, N148);
nor NOR4 (N150, N124, N88, N115, N103);
not NOT1 (N151, N146);
and AND3 (N152, N150, N26, N5);
and AND2 (N153, N135, N107);
and AND3 (N154, N144, N111, N110);
not NOT1 (N155, N136);
or OR2 (N156, N152, N90);
nand NAND3 (N157, N155, N17, N129);
buf BUF1 (N158, N140);
and AND3 (N159, N149, N9, N31);
not NOT1 (N160, N137);
buf BUF1 (N161, N147);
and AND3 (N162, N160, N10, N135);
not NOT1 (N163, N156);
nor NOR2 (N164, N158, N104);
and AND2 (N165, N163, N27);
buf BUF1 (N166, N143);
xor XOR2 (N167, N166, N18);
xor XOR2 (N168, N157, N50);
or OR2 (N169, N153, N150);
or OR4 (N170, N154, N80, N70, N22);
nor NOR4 (N171, N164, N86, N51, N35);
or OR2 (N172, N159, N75);
xor XOR2 (N173, N171, N157);
buf BUF1 (N174, N172);
not NOT1 (N175, N170);
xor XOR2 (N176, N174, N55);
buf BUF1 (N177, N169);
or OR2 (N178, N151, N7);
not NOT1 (N179, N168);
nor NOR2 (N180, N162, N3);
xor XOR2 (N181, N176, N20);
and AND4 (N182, N181, N68, N73, N112);
and AND4 (N183, N175, N62, N148, N118);
nor NOR3 (N184, N177, N133, N139);
nor NOR4 (N185, N182, N102, N119, N70);
nor NOR3 (N186, N184, N38, N151);
xor XOR2 (N187, N185, N46);
and AND4 (N188, N179, N46, N57, N162);
not NOT1 (N189, N187);
buf BUF1 (N190, N183);
and AND3 (N191, N186, N189, N42);
buf BUF1 (N192, N161);
and AND4 (N193, N138, N91, N166, N188);
or OR3 (N194, N89, N155, N71);
or OR3 (N195, N193, N154, N184);
and AND4 (N196, N191, N10, N62, N78);
not NOT1 (N197, N192);
nand NAND4 (N198, N197, N79, N142, N98);
or OR2 (N199, N173, N177);
or OR3 (N200, N180, N166, N106);
xor XOR2 (N201, N195, N146);
xor XOR2 (N202, N167, N128);
and AND3 (N203, N198, N128, N188);
buf BUF1 (N204, N190);
nor NOR3 (N205, N165, N182, N163);
buf BUF1 (N206, N200);
nor NOR4 (N207, N205, N176, N162, N145);
not NOT1 (N208, N194);
and AND2 (N209, N202, N90);
buf BUF1 (N210, N206);
and AND2 (N211, N209, N163);
or OR2 (N212, N203, N181);
or OR3 (N213, N212, N14, N208);
and AND3 (N214, N183, N133, N160);
buf BUF1 (N215, N201);
not NOT1 (N216, N178);
nor NOR2 (N217, N199, N158);
and AND2 (N218, N211, N113);
and AND2 (N219, N207, N116);
or OR3 (N220, N219, N62, N203);
buf BUF1 (N221, N217);
and AND3 (N222, N196, N100, N195);
nor NOR4 (N223, N214, N111, N101, N39);
and AND4 (N224, N223, N41, N60, N69);
nand NAND3 (N225, N213, N210, N96);
not NOT1 (N226, N48);
buf BUF1 (N227, N216);
or OR2 (N228, N225, N216);
not NOT1 (N229, N215);
or OR4 (N230, N204, N140, N197, N200);
nor NOR4 (N231, N221, N143, N30, N5);
nand NAND4 (N232, N228, N11, N9, N116);
and AND3 (N233, N220, N146, N71);
buf BUF1 (N234, N226);
xor XOR2 (N235, N227, N63);
nor NOR3 (N236, N235, N210, N57);
xor XOR2 (N237, N232, N213);
or OR4 (N238, N231, N197, N217, N214);
xor XOR2 (N239, N218, N51);
buf BUF1 (N240, N236);
not NOT1 (N241, N229);
and AND2 (N242, N222, N60);
and AND4 (N243, N233, N179, N214, N138);
or OR3 (N244, N237, N64, N28);
nand NAND2 (N245, N230, N209);
or OR3 (N246, N238, N137, N120);
xor XOR2 (N247, N224, N46);
not NOT1 (N248, N240);
nand NAND3 (N249, N244, N116, N246);
and AND2 (N250, N222, N186);
nor NOR4 (N251, N250, N50, N86, N121);
xor XOR2 (N252, N251, N231);
buf BUF1 (N253, N245);
buf BUF1 (N254, N243);
or OR3 (N255, N252, N142, N67);
nand NAND3 (N256, N242, N7, N76);
buf BUF1 (N257, N254);
and AND3 (N258, N257, N241, N215);
not NOT1 (N259, N59);
nand NAND2 (N260, N256, N229);
buf BUF1 (N261, N234);
nand NAND4 (N262, N259, N227, N8, N107);
or OR2 (N263, N239, N217);
not NOT1 (N264, N249);
and AND3 (N265, N264, N65, N35);
nor NOR4 (N266, N247, N171, N163, N225);
nor NOR3 (N267, N253, N57, N103);
and AND4 (N268, N248, N122, N246, N29);
or OR3 (N269, N265, N97, N183);
or OR2 (N270, N268, N266);
or OR2 (N271, N244, N38);
nand NAND3 (N272, N271, N185, N248);
buf BUF1 (N273, N262);
and AND4 (N274, N260, N173, N26, N69);
xor XOR2 (N275, N272, N259);
or OR3 (N276, N275, N203, N45);
buf BUF1 (N277, N261);
nor NOR4 (N278, N276, N80, N10, N39);
buf BUF1 (N279, N278);
xor XOR2 (N280, N267, N262);
xor XOR2 (N281, N270, N196);
not NOT1 (N282, N269);
xor XOR2 (N283, N280, N43);
nand NAND4 (N284, N258, N7, N113, N255);
not NOT1 (N285, N186);
buf BUF1 (N286, N284);
not NOT1 (N287, N274);
buf BUF1 (N288, N263);
nor NOR3 (N289, N279, N215, N194);
nor NOR4 (N290, N286, N106, N250, N43);
xor XOR2 (N291, N282, N253);
buf BUF1 (N292, N273);
xor XOR2 (N293, N285, N288);
nor NOR2 (N294, N240, N255);
or OR4 (N295, N281, N3, N37, N88);
and AND3 (N296, N291, N261, N183);
buf BUF1 (N297, N287);
nand NAND2 (N298, N294, N166);
xor XOR2 (N299, N283, N248);
or OR3 (N300, N295, N171, N200);
nand NAND2 (N301, N277, N143);
xor XOR2 (N302, N290, N20);
and AND3 (N303, N298, N103, N90);
nor NOR2 (N304, N300, N293);
buf BUF1 (N305, N297);
and AND3 (N306, N87, N48, N8);
nor NOR2 (N307, N299, N177);
buf BUF1 (N308, N292);
nand NAND4 (N309, N289, N104, N119, N87);
and AND2 (N310, N302, N171);
and AND3 (N311, N310, N83, N290);
buf BUF1 (N312, N301);
xor XOR2 (N313, N312, N277);
nand NAND4 (N314, N309, N139, N222, N174);
and AND3 (N315, N305, N31, N38);
xor XOR2 (N316, N314, N104);
xor XOR2 (N317, N311, N55);
xor XOR2 (N318, N317, N287);
nor NOR2 (N319, N315, N8);
or OR3 (N320, N319, N4, N131);
xor XOR2 (N321, N316, N63);
and AND2 (N322, N306, N18);
nor NOR4 (N323, N303, N36, N43, N188);
and AND4 (N324, N307, N146, N235, N68);
nor NOR2 (N325, N313, N19);
and AND3 (N326, N325, N71, N70);
not NOT1 (N327, N326);
xor XOR2 (N328, N323, N298);
or OR2 (N329, N322, N226);
nor NOR2 (N330, N324, N256);
and AND4 (N331, N321, N199, N239, N60);
not NOT1 (N332, N329);
xor XOR2 (N333, N296, N328);
xor XOR2 (N334, N132, N147);
or OR4 (N335, N332, N231, N245, N317);
not NOT1 (N336, N320);
not NOT1 (N337, N333);
buf BUF1 (N338, N334);
nand NAND3 (N339, N338, N188, N268);
and AND2 (N340, N318, N66);
and AND4 (N341, N330, N253, N79, N14);
buf BUF1 (N342, N304);
or OR2 (N343, N335, N253);
and AND4 (N344, N342, N66, N193, N36);
or OR2 (N345, N331, N71);
buf BUF1 (N346, N327);
nand NAND3 (N347, N343, N342, N21);
xor XOR2 (N348, N346, N199);
not NOT1 (N349, N339);
buf BUF1 (N350, N341);
not NOT1 (N351, N350);
or OR4 (N352, N308, N323, N66, N163);
not NOT1 (N353, N345);
buf BUF1 (N354, N351);
and AND4 (N355, N349, N123, N276, N298);
xor XOR2 (N356, N348, N99);
or OR3 (N357, N354, N161, N138);
buf BUF1 (N358, N355);
or OR3 (N359, N337, N19, N181);
xor XOR2 (N360, N336, N278);
nor NOR4 (N361, N344, N241, N169, N240);
or OR3 (N362, N361, N98, N292);
or OR4 (N363, N340, N194, N345, N309);
nor NOR4 (N364, N359, N4, N331, N278);
nand NAND4 (N365, N352, N260, N341, N162);
buf BUF1 (N366, N353);
xor XOR2 (N367, N360, N90);
xor XOR2 (N368, N367, N241);
xor XOR2 (N369, N366, N120);
not NOT1 (N370, N365);
nor NOR2 (N371, N370, N19);
nand NAND2 (N372, N363, N74);
xor XOR2 (N373, N369, N194);
nand NAND3 (N374, N357, N104, N181);
nand NAND2 (N375, N362, N292);
nand NAND2 (N376, N372, N266);
buf BUF1 (N377, N373);
and AND2 (N378, N377, N7);
nand NAND3 (N379, N374, N289, N25);
xor XOR2 (N380, N358, N305);
or OR4 (N381, N368, N148, N212, N249);
or OR2 (N382, N347, N306);
not NOT1 (N383, N381);
nor NOR4 (N384, N375, N19, N285, N135);
nand NAND4 (N385, N356, N22, N2, N12);
nor NOR2 (N386, N364, N24);
not NOT1 (N387, N380);
nor NOR3 (N388, N384, N170, N136);
buf BUF1 (N389, N388);
nor NOR4 (N390, N379, N51, N18, N94);
nand NAND2 (N391, N378, N31);
and AND3 (N392, N382, N107, N169);
or OR4 (N393, N385, N129, N282, N350);
and AND2 (N394, N387, N191);
buf BUF1 (N395, N386);
nand NAND2 (N396, N371, N153);
xor XOR2 (N397, N391, N60);
and AND4 (N398, N390, N237, N347, N318);
and AND4 (N399, N395, N107, N61, N309);
xor XOR2 (N400, N389, N47);
or OR4 (N401, N399, N205, N398, N217);
or OR4 (N402, N274, N292, N367, N322);
xor XOR2 (N403, N402, N157);
xor XOR2 (N404, N392, N326);
buf BUF1 (N405, N400);
or OR4 (N406, N404, N302, N7, N95);
nand NAND4 (N407, N394, N160, N342, N55);
or OR4 (N408, N406, N163, N307, N355);
nor NOR4 (N409, N383, N181, N337, N137);
nand NAND4 (N410, N403, N68, N244, N368);
not NOT1 (N411, N409);
xor XOR2 (N412, N401, N362);
buf BUF1 (N413, N393);
buf BUF1 (N414, N410);
nand NAND3 (N415, N405, N19, N382);
not NOT1 (N416, N396);
not NOT1 (N417, N412);
not NOT1 (N418, N417);
or OR2 (N419, N411, N22);
nor NOR3 (N420, N418, N29, N367);
not NOT1 (N421, N416);
not NOT1 (N422, N420);
not NOT1 (N423, N415);
nand NAND4 (N424, N407, N114, N230, N281);
not NOT1 (N425, N421);
and AND3 (N426, N425, N280, N199);
or OR4 (N427, N419, N193, N354, N139);
nor NOR4 (N428, N408, N198, N188, N308);
nor NOR4 (N429, N423, N373, N142, N6);
buf BUF1 (N430, N397);
buf BUF1 (N431, N376);
nand NAND2 (N432, N428, N196);
and AND2 (N433, N430, N369);
nor NOR3 (N434, N427, N416, N20);
buf BUF1 (N435, N433);
buf BUF1 (N436, N426);
nand NAND4 (N437, N432, N208, N233, N252);
not NOT1 (N438, N434);
or OR3 (N439, N438, N395, N35);
nor NOR4 (N440, N422, N154, N310, N85);
not NOT1 (N441, N431);
buf BUF1 (N442, N436);
xor XOR2 (N443, N429, N220);
or OR2 (N444, N435, N191);
or OR2 (N445, N443, N423);
and AND2 (N446, N442, N297);
nor NOR3 (N447, N437, N372, N48);
nand NAND2 (N448, N445, N210);
xor XOR2 (N449, N414, N58);
nand NAND4 (N450, N441, N6, N208, N323);
nor NOR3 (N451, N424, N263, N128);
buf BUF1 (N452, N450);
xor XOR2 (N453, N448, N31);
and AND2 (N454, N446, N329);
nor NOR4 (N455, N447, N260, N432, N300);
xor XOR2 (N456, N444, N444);
not NOT1 (N457, N452);
buf BUF1 (N458, N454);
not NOT1 (N459, N458);
or OR2 (N460, N439, N152);
buf BUF1 (N461, N460);
or OR4 (N462, N459, N298, N236, N251);
xor XOR2 (N463, N461, N437);
and AND2 (N464, N455, N369);
nand NAND3 (N465, N440, N278, N395);
or OR2 (N466, N456, N143);
xor XOR2 (N467, N449, N370);
or OR4 (N468, N465, N433, N307, N416);
and AND3 (N469, N451, N449, N9);
nand NAND3 (N470, N453, N468, N393);
nand NAND4 (N471, N36, N438, N33, N179);
buf BUF1 (N472, N471);
nand NAND2 (N473, N466, N453);
xor XOR2 (N474, N473, N408);
buf BUF1 (N475, N462);
xor XOR2 (N476, N469, N187);
not NOT1 (N477, N470);
xor XOR2 (N478, N413, N37);
or OR4 (N479, N476, N351, N236, N203);
or OR4 (N480, N479, N133, N288, N429);
buf BUF1 (N481, N474);
buf BUF1 (N482, N467);
not NOT1 (N483, N482);
nor NOR2 (N484, N457, N89);
or OR2 (N485, N472, N191);
or OR2 (N486, N463, N47);
and AND2 (N487, N485, N293);
nor NOR4 (N488, N481, N415, N127, N180);
or OR3 (N489, N486, N345, N122);
not NOT1 (N490, N478);
and AND2 (N491, N475, N218);
or OR4 (N492, N489, N89, N155, N266);
nor NOR4 (N493, N488, N93, N414, N348);
nor NOR3 (N494, N464, N422, N175);
buf BUF1 (N495, N483);
xor XOR2 (N496, N487, N147);
buf BUF1 (N497, N491);
or OR3 (N498, N496, N76, N65);
buf BUF1 (N499, N477);
nand NAND3 (N500, N494, N347, N455);
or OR4 (N501, N500, N317, N203, N466);
nand NAND2 (N502, N492, N62);
nor NOR2 (N503, N480, N7);
buf BUF1 (N504, N502);
and AND4 (N505, N504, N231, N408, N445);
nand NAND4 (N506, N505, N7, N324, N191);
and AND2 (N507, N501, N323);
buf BUF1 (N508, N507);
or OR3 (N509, N484, N75, N206);
and AND2 (N510, N497, N273);
nor NOR4 (N511, N510, N449, N343, N160);
nand NAND3 (N512, N508, N44, N307);
xor XOR2 (N513, N498, N215);
or OR3 (N514, N493, N402, N368);
and AND4 (N515, N514, N477, N276, N187);
nand NAND3 (N516, N499, N22, N457);
and AND4 (N517, N515, N28, N316, N20);
nor NOR4 (N518, N495, N266, N187, N104);
not NOT1 (N519, N517);
nand NAND4 (N520, N513, N312, N148, N489);
buf BUF1 (N521, N490);
and AND4 (N522, N518, N179, N84, N418);
buf BUF1 (N523, N516);
endmodule