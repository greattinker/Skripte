// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15;

output N25914,N25911,N25894,N25898,N25885,N25902,N25912,N25906,N25913,N25915;

nor NOR3 (N16, N10, N5, N9);
xor XOR2 (N17, N8, N16);
nor NOR3 (N18, N11, N1, N16);
nor NOR2 (N19, N14, N14);
nor NOR2 (N20, N14, N9);
or OR3 (N21, N8, N6, N5);
buf BUF1 (N22, N4);
and AND4 (N23, N19, N14, N22, N20);
or OR3 (N24, N21, N14, N11);
not NOT1 (N25, N24);
and AND2 (N26, N13, N15);
not NOT1 (N27, N21);
nor NOR4 (N28, N13, N24, N10, N2);
or OR2 (N29, N15, N3);
not NOT1 (N30, N17);
buf BUF1 (N31, N26);
nand NAND4 (N32, N10, N19, N19, N2);
nand NAND4 (N33, N6, N27, N24, N21);
buf BUF1 (N34, N2);
and AND3 (N35, N34, N18, N11);
nand NAND4 (N36, N15, N30, N11, N8);
nor NOR4 (N37, N32, N17, N12, N32);
buf BUF1 (N38, N8);
or OR4 (N39, N38, N34, N9, N33);
not NOT1 (N40, N3);
and AND4 (N41, N37, N4, N15, N11);
or OR4 (N42, N40, N30, N18, N2);
xor XOR2 (N43, N39, N10);
not NOT1 (N44, N43);
or OR2 (N45, N41, N6);
not NOT1 (N46, N35);
nand NAND3 (N47, N36, N26, N14);
and AND2 (N48, N42, N30);
or OR2 (N49, N25, N19);
nand NAND3 (N50, N44, N39, N2);
buf BUF1 (N51, N45);
nor NOR2 (N52, N29, N45);
xor XOR2 (N53, N51, N10);
xor XOR2 (N54, N49, N39);
not NOT1 (N55, N31);
buf BUF1 (N56, N28);
buf BUF1 (N57, N48);
or OR4 (N58, N23, N25, N5, N26);
not NOT1 (N59, N50);
or OR3 (N60, N47, N52, N44);
nand NAND2 (N61, N30, N50);
xor XOR2 (N62, N56, N57);
and AND3 (N63, N38, N58, N21);
buf BUF1 (N64, N44);
nand NAND4 (N65, N59, N6, N44, N51);
buf BUF1 (N66, N55);
nand NAND4 (N67, N63, N33, N36, N25);
nor NOR4 (N68, N62, N65, N27, N54);
and AND4 (N69, N5, N36, N58, N45);
nand NAND2 (N70, N60, N24);
xor XOR2 (N71, N10, N17);
not NOT1 (N72, N61);
nand NAND2 (N73, N72, N67);
xor XOR2 (N74, N33, N11);
nand NAND3 (N75, N69, N7, N45);
not NOT1 (N76, N74);
nand NAND3 (N77, N53, N63, N70);
not NOT1 (N78, N60);
not NOT1 (N79, N78);
not NOT1 (N80, N75);
and AND3 (N81, N79, N7, N2);
nand NAND3 (N82, N80, N49, N25);
buf BUF1 (N83, N77);
nor NOR2 (N84, N66, N36);
not NOT1 (N85, N73);
nand NAND2 (N86, N81, N60);
buf BUF1 (N87, N83);
buf BUF1 (N88, N84);
xor XOR2 (N89, N86, N29);
or OR3 (N90, N68, N3, N4);
and AND2 (N91, N88, N86);
buf BUF1 (N92, N87);
buf BUF1 (N93, N46);
and AND4 (N94, N76, N38, N90, N92);
nor NOR4 (N95, N16, N58, N72, N14);
xor XOR2 (N96, N49, N55);
nor NOR2 (N97, N89, N45);
nand NAND3 (N98, N91, N60, N41);
or OR3 (N99, N94, N97, N93);
nor NOR4 (N100, N39, N69, N14, N69);
nor NOR3 (N101, N37, N7, N53);
not NOT1 (N102, N82);
or OR4 (N103, N99, N102, N74, N84);
nand NAND2 (N104, N62, N96);
nor NOR2 (N105, N87, N49);
and AND2 (N106, N101, N103);
nor NOR3 (N107, N41, N45, N58);
nand NAND2 (N108, N106, N100);
buf BUF1 (N109, N93);
buf BUF1 (N110, N108);
nand NAND2 (N111, N85, N18);
not NOT1 (N112, N64);
xor XOR2 (N113, N105, N35);
not NOT1 (N114, N111);
and AND4 (N115, N109, N63, N88, N82);
xor XOR2 (N116, N104, N30);
and AND2 (N117, N115, N90);
nand NAND4 (N118, N98, N101, N108, N20);
buf BUF1 (N119, N113);
nor NOR4 (N120, N117, N79, N92, N110);
xor XOR2 (N121, N12, N29);
nor NOR2 (N122, N120, N33);
xor XOR2 (N123, N118, N96);
and AND4 (N124, N123, N78, N107, N89);
or OR2 (N125, N109, N65);
not NOT1 (N126, N95);
buf BUF1 (N127, N122);
xor XOR2 (N128, N124, N26);
and AND4 (N129, N126, N69, N83, N36);
nand NAND3 (N130, N71, N4, N129);
or OR2 (N131, N129, N113);
xor XOR2 (N132, N119, N32);
or OR2 (N133, N132, N63);
and AND4 (N134, N125, N42, N35, N92);
and AND4 (N135, N128, N31, N126, N55);
buf BUF1 (N136, N130);
nor NOR4 (N137, N133, N96, N87, N52);
and AND2 (N138, N116, N126);
nor NOR4 (N139, N134, N120, N25, N3);
not NOT1 (N140, N139);
xor XOR2 (N141, N127, N94);
and AND4 (N142, N121, N105, N63, N15);
or OR3 (N143, N140, N20, N102);
nor NOR2 (N144, N135, N101);
nor NOR2 (N145, N144, N121);
buf BUF1 (N146, N112);
nor NOR4 (N147, N145, N118, N101, N48);
buf BUF1 (N148, N137);
xor XOR2 (N149, N148, N38);
nor NOR4 (N150, N141, N27, N108, N118);
nor NOR3 (N151, N147, N45, N148);
nand NAND4 (N152, N114, N87, N144, N18);
or OR2 (N153, N136, N55);
xor XOR2 (N154, N143, N6);
buf BUF1 (N155, N138);
nand NAND2 (N156, N151, N53);
nand NAND4 (N157, N150, N68, N78, N51);
not NOT1 (N158, N142);
buf BUF1 (N159, N152);
xor XOR2 (N160, N131, N81);
or OR3 (N161, N159, N136, N116);
xor XOR2 (N162, N153, N4);
nand NAND4 (N163, N162, N41, N132, N67);
nand NAND2 (N164, N160, N134);
and AND2 (N165, N156, N63);
or OR2 (N166, N146, N3);
buf BUF1 (N167, N157);
buf BUF1 (N168, N158);
xor XOR2 (N169, N161, N131);
nand NAND3 (N170, N169, N9, N92);
xor XOR2 (N171, N163, N104);
not NOT1 (N172, N170);
buf BUF1 (N173, N164);
and AND2 (N174, N173, N51);
xor XOR2 (N175, N168, N21);
and AND3 (N176, N171, N86, N51);
nor NOR2 (N177, N167, N92);
nand NAND4 (N178, N174, N157, N29, N9);
not NOT1 (N179, N172);
nor NOR4 (N180, N154, N139, N21, N92);
nor NOR3 (N181, N179, N78, N108);
nand NAND4 (N182, N165, N178, N72, N66);
not NOT1 (N183, N135);
nor NOR2 (N184, N176, N123);
not NOT1 (N185, N184);
xor XOR2 (N186, N183, N169);
not NOT1 (N187, N181);
nand NAND2 (N188, N182, N152);
not NOT1 (N189, N187);
buf BUF1 (N190, N185);
nand NAND3 (N191, N190, N28, N68);
xor XOR2 (N192, N155, N158);
or OR3 (N193, N186, N57, N169);
nand NAND3 (N194, N192, N171, N52);
xor XOR2 (N195, N175, N33);
nor NOR4 (N196, N149, N134, N179, N51);
and AND2 (N197, N166, N114);
buf BUF1 (N198, N180);
nor NOR3 (N199, N189, N15, N188);
and AND2 (N200, N50, N159);
nand NAND2 (N201, N193, N27);
nor NOR4 (N202, N197, N84, N190, N139);
or OR4 (N203, N195, N2, N166, N35);
nand NAND4 (N204, N202, N124, N127, N141);
nor NOR4 (N205, N191, N87, N75, N128);
nand NAND2 (N206, N194, N129);
and AND4 (N207, N203, N73, N74, N90);
buf BUF1 (N208, N207);
buf BUF1 (N209, N206);
or OR2 (N210, N208, N22);
nand NAND2 (N211, N210, N122);
buf BUF1 (N212, N205);
nand NAND3 (N213, N196, N112, N29);
xor XOR2 (N214, N199, N196);
and AND2 (N215, N201, N18);
xor XOR2 (N216, N200, N200);
and AND3 (N217, N216, N73, N102);
not NOT1 (N218, N211);
and AND2 (N219, N213, N86);
buf BUF1 (N220, N217);
nand NAND4 (N221, N212, N48, N111, N6);
nor NOR2 (N222, N218, N78);
and AND2 (N223, N222, N1);
or OR2 (N224, N198, N28);
and AND4 (N225, N215, N176, N175, N23);
nand NAND4 (N226, N224, N125, N170, N36);
nor NOR3 (N227, N214, N155, N89);
nand NAND3 (N228, N226, N174, N76);
not NOT1 (N229, N220);
nor NOR3 (N230, N219, N46, N53);
xor XOR2 (N231, N177, N180);
nand NAND2 (N232, N221, N118);
or OR2 (N233, N209, N141);
nand NAND4 (N234, N229, N221, N66, N26);
nand NAND4 (N235, N227, N164, N117, N99);
nand NAND2 (N236, N234, N7);
buf BUF1 (N237, N204);
buf BUF1 (N238, N225);
nor NOR4 (N239, N236, N109, N207, N124);
nand NAND2 (N240, N239, N235);
buf BUF1 (N241, N207);
nand NAND3 (N242, N230, N175, N227);
xor XOR2 (N243, N223, N47);
and AND4 (N244, N240, N176, N1, N171);
nand NAND4 (N245, N244, N220, N53, N211);
or OR4 (N246, N231, N176, N243, N39);
nand NAND2 (N247, N136, N89);
xor XOR2 (N248, N245, N2);
xor XOR2 (N249, N248, N17);
buf BUF1 (N250, N232);
buf BUF1 (N251, N242);
buf BUF1 (N252, N247);
and AND4 (N253, N249, N100, N25, N155);
xor XOR2 (N254, N238, N114);
nand NAND4 (N255, N233, N93, N186, N165);
not NOT1 (N256, N241);
nor NOR3 (N257, N237, N81, N157);
buf BUF1 (N258, N251);
and AND3 (N259, N252, N213, N199);
not NOT1 (N260, N256);
nand NAND4 (N261, N257, N34, N68, N242);
and AND3 (N262, N260, N4, N6);
nand NAND2 (N263, N261, N209);
nand NAND4 (N264, N255, N241, N232, N152);
buf BUF1 (N265, N264);
buf BUF1 (N266, N262);
or OR2 (N267, N259, N4);
xor XOR2 (N268, N265, N131);
nor NOR3 (N269, N268, N30, N227);
buf BUF1 (N270, N250);
nand NAND4 (N271, N270, N35, N12, N200);
buf BUF1 (N272, N246);
nand NAND2 (N273, N228, N36);
not NOT1 (N274, N269);
and AND3 (N275, N253, N274, N232);
and AND4 (N276, N235, N202, N253, N193);
and AND2 (N277, N271, N148);
or OR3 (N278, N266, N271, N227);
and AND2 (N279, N275, N202);
xor XOR2 (N280, N258, N22);
buf BUF1 (N281, N267);
not NOT1 (N282, N280);
nand NAND4 (N283, N282, N46, N271, N133);
nor NOR4 (N284, N272, N22, N191, N229);
xor XOR2 (N285, N276, N41);
nand NAND3 (N286, N277, N259, N200);
nand NAND3 (N287, N285, N276, N278);
and AND2 (N288, N178, N226);
nand NAND3 (N289, N281, N101, N5);
xor XOR2 (N290, N263, N128);
nor NOR3 (N291, N284, N25, N140);
and AND3 (N292, N289, N150, N236);
xor XOR2 (N293, N273, N248);
nor NOR4 (N294, N292, N188, N208, N220);
buf BUF1 (N295, N286);
not NOT1 (N296, N283);
nor NOR4 (N297, N287, N107, N167, N209);
nor NOR3 (N298, N291, N190, N6);
xor XOR2 (N299, N295, N252);
nor NOR2 (N300, N297, N228);
or OR2 (N301, N254, N56);
or OR4 (N302, N300, N108, N137, N298);
or OR2 (N303, N5, N221);
not NOT1 (N304, N296);
buf BUF1 (N305, N294);
nor NOR4 (N306, N305, N199, N266, N209);
nand NAND4 (N307, N279, N142, N128, N241);
buf BUF1 (N308, N293);
nor NOR4 (N309, N304, N86, N166, N215);
not NOT1 (N310, N290);
xor XOR2 (N311, N302, N87);
nand NAND2 (N312, N311, N206);
or OR3 (N313, N310, N36, N186);
not NOT1 (N314, N309);
xor XOR2 (N315, N307, N166);
or OR2 (N316, N313, N117);
buf BUF1 (N317, N308);
and AND2 (N318, N316, N152);
not NOT1 (N319, N303);
nand NAND2 (N320, N318, N175);
nor NOR4 (N321, N319, N318, N168, N264);
or OR4 (N322, N317, N220, N63, N233);
and AND4 (N323, N299, N56, N209, N43);
or OR4 (N324, N312, N29, N314, N252);
or OR3 (N325, N269, N217, N171);
nor NOR2 (N326, N325, N153);
not NOT1 (N327, N320);
xor XOR2 (N328, N321, N187);
buf BUF1 (N329, N324);
buf BUF1 (N330, N288);
buf BUF1 (N331, N323);
not NOT1 (N332, N322);
buf BUF1 (N333, N330);
nand NAND2 (N334, N331, N150);
not NOT1 (N335, N333);
buf BUF1 (N336, N327);
nand NAND3 (N337, N301, N166, N269);
not NOT1 (N338, N335);
nor NOR2 (N339, N332, N72);
xor XOR2 (N340, N336, N198);
or OR3 (N341, N339, N117, N12);
nand NAND3 (N342, N315, N195, N208);
nand NAND4 (N343, N340, N323, N250, N267);
nor NOR4 (N344, N329, N333, N249, N189);
or OR2 (N345, N337, N272);
or OR2 (N346, N345, N88);
not NOT1 (N347, N344);
nor NOR2 (N348, N346, N210);
not NOT1 (N349, N306);
nand NAND3 (N350, N326, N317, N254);
and AND4 (N351, N349, N350, N166, N182);
nor NOR3 (N352, N40, N263, N312);
nor NOR2 (N353, N348, N201);
not NOT1 (N354, N338);
or OR2 (N355, N343, N44);
not NOT1 (N356, N334);
nand NAND3 (N357, N353, N211, N113);
xor XOR2 (N358, N355, N154);
nand NAND3 (N359, N341, N289, N77);
buf BUF1 (N360, N347);
or OR2 (N361, N356, N38);
not NOT1 (N362, N358);
nand NAND3 (N363, N328, N133, N82);
not NOT1 (N364, N342);
nand NAND4 (N365, N351, N103, N49, N277);
and AND3 (N366, N354, N205, N153);
and AND3 (N367, N360, N267, N280);
nand NAND3 (N368, N361, N254, N46);
not NOT1 (N369, N368);
and AND2 (N370, N367, N151);
nor NOR3 (N371, N366, N363, N58);
buf BUF1 (N372, N273);
buf BUF1 (N373, N370);
xor XOR2 (N374, N359, N7);
or OR4 (N375, N364, N372, N269, N92);
nor NOR2 (N376, N251, N310);
and AND2 (N377, N373, N54);
xor XOR2 (N378, N357, N368);
not NOT1 (N379, N365);
nand NAND2 (N380, N374, N121);
and AND3 (N381, N378, N86, N228);
or OR3 (N382, N371, N358, N181);
and AND4 (N383, N352, N116, N288, N104);
or OR3 (N384, N379, N273, N345);
buf BUF1 (N385, N381);
nor NOR2 (N386, N380, N92);
nor NOR3 (N387, N375, N82, N34);
xor XOR2 (N388, N384, N355);
xor XOR2 (N389, N369, N326);
and AND2 (N390, N362, N338);
xor XOR2 (N391, N388, N134);
nand NAND2 (N392, N390, N146);
or OR2 (N393, N383, N365);
buf BUF1 (N394, N376);
buf BUF1 (N395, N386);
and AND3 (N396, N391, N252, N99);
not NOT1 (N397, N389);
nor NOR2 (N398, N394, N383);
xor XOR2 (N399, N385, N124);
nand NAND3 (N400, N397, N78, N38);
nor NOR2 (N401, N398, N10);
buf BUF1 (N402, N377);
not NOT1 (N403, N395);
buf BUF1 (N404, N401);
buf BUF1 (N405, N402);
nand NAND2 (N406, N393, N289);
xor XOR2 (N407, N399, N202);
nand NAND2 (N408, N400, N104);
nor NOR2 (N409, N392, N376);
nand NAND4 (N410, N406, N113, N289, N296);
not NOT1 (N411, N396);
and AND4 (N412, N405, N57, N396, N199);
nor NOR3 (N413, N411, N291, N403);
xor XOR2 (N414, N383, N355);
not NOT1 (N415, N414);
buf BUF1 (N416, N409);
not NOT1 (N417, N382);
not NOT1 (N418, N412);
and AND2 (N419, N387, N363);
xor XOR2 (N420, N416, N158);
not NOT1 (N421, N420);
nor NOR3 (N422, N408, N135, N136);
buf BUF1 (N423, N421);
nand NAND3 (N424, N422, N308, N92);
not NOT1 (N425, N417);
not NOT1 (N426, N410);
buf BUF1 (N427, N413);
or OR4 (N428, N423, N274, N87, N36);
not NOT1 (N429, N407);
or OR4 (N430, N427, N13, N85, N62);
or OR2 (N431, N428, N145);
xor XOR2 (N432, N429, N120);
nor NOR2 (N433, N431, N322);
nor NOR3 (N434, N419, N156, N105);
not NOT1 (N435, N430);
and AND4 (N436, N435, N410, N253, N121);
and AND3 (N437, N426, N423, N205);
or OR3 (N438, N436, N7, N66);
or OR2 (N439, N438, N46);
nor NOR4 (N440, N415, N198, N51, N387);
and AND3 (N441, N440, N269, N341);
nand NAND4 (N442, N424, N352, N182, N5);
nor NOR4 (N443, N441, N122, N302, N279);
buf BUF1 (N444, N442);
or OR2 (N445, N404, N32);
not NOT1 (N446, N432);
or OR2 (N447, N437, N371);
nand NAND2 (N448, N445, N354);
not NOT1 (N449, N443);
or OR3 (N450, N434, N284, N110);
or OR3 (N451, N444, N447, N365);
and AND3 (N452, N358, N255, N130);
nor NOR4 (N453, N448, N129, N174, N387);
and AND3 (N454, N452, N414, N35);
or OR4 (N455, N451, N233, N93, N395);
not NOT1 (N456, N450);
xor XOR2 (N457, N455, N66);
buf BUF1 (N458, N446);
nor NOR4 (N459, N457, N224, N287, N164);
xor XOR2 (N460, N454, N421);
nor NOR2 (N461, N458, N209);
nand NAND4 (N462, N418, N263, N382, N40);
not NOT1 (N463, N433);
xor XOR2 (N464, N460, N131);
buf BUF1 (N465, N449);
or OR3 (N466, N456, N134, N41);
nor NOR4 (N467, N425, N290, N231, N27);
nor NOR4 (N468, N463, N328, N291, N83);
nand NAND2 (N469, N439, N163);
nand NAND3 (N470, N469, N286, N370);
nor NOR4 (N471, N470, N63, N413, N41);
nor NOR4 (N472, N464, N267, N365, N410);
and AND2 (N473, N468, N63);
or OR4 (N474, N472, N204, N192, N129);
xor XOR2 (N475, N474, N411);
and AND4 (N476, N465, N214, N409, N2);
nand NAND4 (N477, N467, N84, N354, N142);
nor NOR3 (N478, N459, N331, N145);
not NOT1 (N479, N462);
and AND3 (N480, N476, N265, N411);
buf BUF1 (N481, N453);
nor NOR4 (N482, N475, N331, N411, N426);
and AND2 (N483, N482, N277);
or OR2 (N484, N478, N428);
or OR4 (N485, N483, N309, N107, N226);
nor NOR2 (N486, N477, N356);
not NOT1 (N487, N461);
nand NAND2 (N488, N486, N310);
nand NAND2 (N489, N488, N55);
nor NOR4 (N490, N480, N272, N319, N377);
and AND2 (N491, N479, N336);
or OR4 (N492, N473, N96, N350, N317);
xor XOR2 (N493, N471, N250);
and AND4 (N494, N484, N234, N48, N148);
not NOT1 (N495, N492);
buf BUF1 (N496, N495);
nand NAND4 (N497, N494, N151, N44, N493);
or OR3 (N498, N397, N197, N80);
not NOT1 (N499, N487);
buf BUF1 (N500, N489);
nor NOR4 (N501, N496, N285, N444, N416);
xor XOR2 (N502, N490, N45);
nor NOR2 (N503, N481, N423);
xor XOR2 (N504, N498, N121);
nor NOR2 (N505, N503, N51);
not NOT1 (N506, N485);
or OR3 (N507, N505, N220, N406);
buf BUF1 (N508, N504);
not NOT1 (N509, N501);
and AND3 (N510, N507, N10, N276);
buf BUF1 (N511, N510);
nand NAND3 (N512, N499, N490, N88);
xor XOR2 (N513, N509, N191);
and AND4 (N514, N466, N322, N374, N321);
not NOT1 (N515, N511);
not NOT1 (N516, N514);
or OR4 (N517, N515, N78, N356, N465);
and AND3 (N518, N516, N257, N147);
not NOT1 (N519, N508);
or OR3 (N520, N519, N407, N282);
nor NOR2 (N521, N517, N374);
and AND2 (N522, N513, N162);
not NOT1 (N523, N497);
nand NAND3 (N524, N522, N359, N280);
nand NAND2 (N525, N518, N204);
and AND4 (N526, N500, N330, N366, N44);
xor XOR2 (N527, N526, N240);
nand NAND2 (N528, N527, N51);
xor XOR2 (N529, N502, N246);
or OR2 (N530, N491, N260);
nor NOR4 (N531, N523, N264, N492, N398);
and AND3 (N532, N521, N291, N233);
nand NAND4 (N533, N524, N397, N125, N66);
xor XOR2 (N534, N520, N253);
and AND4 (N535, N528, N360, N81, N262);
xor XOR2 (N536, N512, N494);
and AND4 (N537, N535, N293, N14, N113);
and AND4 (N538, N530, N231, N280, N93);
nand NAND4 (N539, N533, N355, N333, N431);
and AND3 (N540, N534, N220, N482);
xor XOR2 (N541, N537, N63);
nor NOR4 (N542, N506, N449, N110, N174);
nand NAND2 (N543, N536, N220);
not NOT1 (N544, N540);
nor NOR2 (N545, N541, N157);
or OR4 (N546, N539, N466, N514, N428);
nand NAND4 (N547, N542, N160, N456, N453);
nand NAND3 (N548, N525, N105, N294);
or OR4 (N549, N544, N31, N164, N299);
nor NOR3 (N550, N546, N540, N412);
buf BUF1 (N551, N547);
and AND3 (N552, N532, N489, N400);
or OR3 (N553, N550, N35, N164);
buf BUF1 (N554, N549);
buf BUF1 (N555, N551);
buf BUF1 (N556, N531);
xor XOR2 (N557, N555, N400);
and AND2 (N558, N553, N178);
nand NAND3 (N559, N529, N520, N49);
buf BUF1 (N560, N556);
buf BUF1 (N561, N558);
not NOT1 (N562, N543);
xor XOR2 (N563, N559, N171);
buf BUF1 (N564, N552);
and AND4 (N565, N548, N442, N241, N290);
not NOT1 (N566, N554);
buf BUF1 (N567, N538);
buf BUF1 (N568, N557);
nand NAND2 (N569, N560, N293);
not NOT1 (N570, N566);
or OR4 (N571, N565, N559, N192, N68);
nor NOR4 (N572, N570, N218, N433, N532);
xor XOR2 (N573, N568, N168);
nand NAND4 (N574, N563, N418, N75, N325);
xor XOR2 (N575, N564, N340);
nand NAND3 (N576, N567, N95, N433);
or OR4 (N577, N575, N10, N228, N397);
nand NAND3 (N578, N569, N102, N15);
not NOT1 (N579, N561);
nand NAND2 (N580, N574, N244);
or OR2 (N581, N545, N373);
nand NAND3 (N582, N580, N145, N371);
xor XOR2 (N583, N572, N324);
xor XOR2 (N584, N583, N372);
and AND2 (N585, N573, N330);
or OR3 (N586, N585, N166, N178);
nand NAND3 (N587, N584, N479, N300);
xor XOR2 (N588, N581, N341);
and AND4 (N589, N562, N49, N556, N83);
buf BUF1 (N590, N588);
nand NAND2 (N591, N579, N72);
nor NOR3 (N592, N591, N587, N196);
nand NAND4 (N593, N283, N7, N444, N255);
or OR2 (N594, N593, N202);
nor NOR3 (N595, N577, N480, N518);
buf BUF1 (N596, N582);
nor NOR4 (N597, N571, N478, N277, N439);
or OR2 (N598, N596, N204);
not NOT1 (N599, N586);
not NOT1 (N600, N597);
xor XOR2 (N601, N576, N436);
xor XOR2 (N602, N589, N570);
not NOT1 (N603, N592);
buf BUF1 (N604, N594);
nand NAND3 (N605, N578, N194, N228);
buf BUF1 (N606, N595);
and AND2 (N607, N606, N49);
nand NAND3 (N608, N599, N506, N460);
nand NAND2 (N609, N604, N340);
buf BUF1 (N610, N603);
and AND2 (N611, N600, N181);
nand NAND4 (N612, N611, N521, N475, N152);
nand NAND4 (N613, N602, N351, N419, N444);
buf BUF1 (N614, N605);
nor NOR2 (N615, N590, N433);
or OR3 (N616, N612, N295, N588);
and AND4 (N617, N598, N461, N143, N506);
buf BUF1 (N618, N601);
and AND2 (N619, N615, N569);
and AND4 (N620, N613, N560, N22, N102);
not NOT1 (N621, N617);
or OR4 (N622, N610, N615, N525, N295);
nor NOR4 (N623, N608, N442, N544, N590);
and AND4 (N624, N614, N309, N74, N50);
nor NOR4 (N625, N624, N244, N329, N425);
and AND3 (N626, N619, N359, N580);
or OR3 (N627, N618, N211, N560);
and AND2 (N628, N620, N246);
xor XOR2 (N629, N607, N615);
not NOT1 (N630, N626);
xor XOR2 (N631, N630, N74);
or OR3 (N632, N629, N596, N182);
or OR3 (N633, N631, N468, N9);
xor XOR2 (N634, N628, N468);
and AND2 (N635, N621, N411);
buf BUF1 (N636, N616);
buf BUF1 (N637, N636);
buf BUF1 (N638, N622);
or OR4 (N639, N633, N125, N85, N152);
and AND2 (N640, N639, N384);
or OR4 (N641, N635, N84, N351, N440);
nor NOR3 (N642, N632, N283, N440);
xor XOR2 (N643, N634, N552);
nand NAND3 (N644, N627, N382, N198);
xor XOR2 (N645, N642, N393);
xor XOR2 (N646, N645, N35);
or OR2 (N647, N643, N512);
nand NAND3 (N648, N644, N580, N512);
nand NAND4 (N649, N638, N47, N152, N14);
xor XOR2 (N650, N623, N161);
xor XOR2 (N651, N609, N199);
and AND2 (N652, N637, N636);
xor XOR2 (N653, N650, N632);
and AND4 (N654, N641, N259, N478, N453);
or OR3 (N655, N649, N180, N83);
not NOT1 (N656, N654);
buf BUF1 (N657, N640);
xor XOR2 (N658, N647, N41);
not NOT1 (N659, N658);
buf BUF1 (N660, N651);
nand NAND3 (N661, N660, N61, N276);
and AND2 (N662, N659, N214);
xor XOR2 (N663, N655, N130);
or OR3 (N664, N652, N517, N44);
xor XOR2 (N665, N656, N233);
or OR4 (N666, N657, N417, N583, N627);
and AND3 (N667, N646, N156, N197);
not NOT1 (N668, N648);
not NOT1 (N669, N666);
or OR2 (N670, N664, N486);
buf BUF1 (N671, N667);
buf BUF1 (N672, N669);
or OR2 (N673, N663, N345);
not NOT1 (N674, N671);
and AND2 (N675, N625, N668);
or OR4 (N676, N248, N647, N160, N514);
buf BUF1 (N677, N662);
or OR2 (N678, N675, N301);
buf BUF1 (N679, N673);
xor XOR2 (N680, N677, N209);
not NOT1 (N681, N674);
and AND3 (N682, N672, N479, N140);
nand NAND4 (N683, N676, N548, N638, N35);
not NOT1 (N684, N678);
and AND2 (N685, N680, N332);
not NOT1 (N686, N653);
buf BUF1 (N687, N665);
or OR3 (N688, N687, N79, N297);
nor NOR4 (N689, N683, N436, N242, N636);
not NOT1 (N690, N681);
nor NOR4 (N691, N661, N605, N263, N614);
nor NOR3 (N692, N691, N151, N563);
or OR2 (N693, N688, N586);
xor XOR2 (N694, N685, N631);
buf BUF1 (N695, N694);
and AND4 (N696, N682, N679, N547, N113);
and AND2 (N697, N239, N39);
nand NAND4 (N698, N692, N367, N100, N76);
xor XOR2 (N699, N684, N323);
not NOT1 (N700, N693);
xor XOR2 (N701, N686, N171);
buf BUF1 (N702, N699);
buf BUF1 (N703, N700);
nand NAND4 (N704, N697, N23, N183, N616);
and AND4 (N705, N689, N47, N36, N90);
nand NAND3 (N706, N670, N389, N44);
nor NOR3 (N707, N703, N633, N141);
and AND4 (N708, N706, N71, N612, N176);
and AND2 (N709, N696, N473);
xor XOR2 (N710, N709, N70);
or OR2 (N711, N695, N641);
buf BUF1 (N712, N702);
not NOT1 (N713, N708);
xor XOR2 (N714, N712, N377);
xor XOR2 (N715, N704, N495);
not NOT1 (N716, N714);
xor XOR2 (N717, N707, N134);
nand NAND3 (N718, N690, N235, N354);
xor XOR2 (N719, N713, N243);
buf BUF1 (N720, N719);
buf BUF1 (N721, N718);
nand NAND4 (N722, N715, N17, N83, N444);
xor XOR2 (N723, N705, N18);
nor NOR4 (N724, N721, N368, N187, N688);
not NOT1 (N725, N701);
nor NOR3 (N726, N723, N210, N191);
nor NOR3 (N727, N698, N183, N30);
and AND4 (N728, N724, N554, N334, N258);
buf BUF1 (N729, N722);
or OR4 (N730, N716, N647, N414, N281);
xor XOR2 (N731, N728, N540);
nor NOR3 (N732, N731, N4, N133);
or OR3 (N733, N711, N219, N725);
and AND3 (N734, N730, N353, N259);
buf BUF1 (N735, N723);
not NOT1 (N736, N729);
or OR3 (N737, N736, N237, N534);
nor NOR3 (N738, N727, N704, N218);
not NOT1 (N739, N733);
xor XOR2 (N740, N717, N195);
not NOT1 (N741, N739);
xor XOR2 (N742, N741, N288);
buf BUF1 (N743, N710);
xor XOR2 (N744, N740, N83);
or OR4 (N745, N744, N179, N244, N40);
nor NOR4 (N746, N742, N131, N412, N543);
nand NAND3 (N747, N746, N320, N7);
not NOT1 (N748, N743);
buf BUF1 (N749, N737);
xor XOR2 (N750, N749, N402);
nand NAND3 (N751, N738, N135, N83);
or OR4 (N752, N745, N378, N548, N699);
nand NAND4 (N753, N752, N174, N536, N614);
nand NAND3 (N754, N750, N719, N537);
or OR2 (N755, N734, N271);
buf BUF1 (N756, N747);
nor NOR3 (N757, N732, N627, N381);
buf BUF1 (N758, N753);
or OR3 (N759, N755, N625, N458);
buf BUF1 (N760, N720);
buf BUF1 (N761, N754);
xor XOR2 (N762, N756, N618);
or OR3 (N763, N762, N371, N108);
and AND3 (N764, N760, N304, N301);
nor NOR2 (N765, N751, N94);
buf BUF1 (N766, N765);
or OR3 (N767, N766, N271, N626);
and AND3 (N768, N748, N254, N201);
buf BUF1 (N769, N761);
nor NOR2 (N770, N763, N653);
or OR2 (N771, N757, N10);
or OR4 (N772, N768, N503, N56, N47);
xor XOR2 (N773, N769, N306);
or OR2 (N774, N735, N528);
or OR3 (N775, N773, N221, N416);
xor XOR2 (N776, N758, N308);
and AND4 (N777, N772, N587, N211, N66);
nand NAND4 (N778, N776, N383, N634, N61);
nor NOR2 (N779, N774, N173);
buf BUF1 (N780, N764);
nor NOR2 (N781, N771, N271);
xor XOR2 (N782, N781, N150);
nor NOR2 (N783, N777, N764);
or OR2 (N784, N726, N232);
buf BUF1 (N785, N770);
or OR4 (N786, N783, N232, N575, N614);
and AND3 (N787, N779, N628, N576);
not NOT1 (N788, N775);
buf BUF1 (N789, N767);
or OR2 (N790, N780, N558);
and AND3 (N791, N786, N156, N130);
buf BUF1 (N792, N789);
nor NOR4 (N793, N784, N535, N368, N168);
nor NOR2 (N794, N792, N417);
buf BUF1 (N795, N790);
xor XOR2 (N796, N794, N171);
xor XOR2 (N797, N782, N267);
and AND3 (N798, N759, N54, N649);
buf BUF1 (N799, N785);
nand NAND4 (N800, N793, N545, N496, N263);
nor NOR2 (N801, N787, N199);
not NOT1 (N802, N778);
xor XOR2 (N803, N802, N412);
and AND4 (N804, N799, N357, N334, N433);
buf BUF1 (N805, N796);
not NOT1 (N806, N805);
not NOT1 (N807, N798);
nor NOR4 (N808, N807, N73, N803, N682);
xor XOR2 (N809, N508, N540);
buf BUF1 (N810, N800);
nand NAND2 (N811, N795, N567);
xor XOR2 (N812, N808, N267);
or OR4 (N813, N788, N86, N515, N811);
not NOT1 (N814, N654);
buf BUF1 (N815, N797);
buf BUF1 (N816, N815);
and AND4 (N817, N806, N547, N587, N648);
not NOT1 (N818, N817);
not NOT1 (N819, N812);
nand NAND4 (N820, N801, N614, N567, N88);
not NOT1 (N821, N818);
buf BUF1 (N822, N814);
xor XOR2 (N823, N813, N331);
nand NAND4 (N824, N804, N334, N217, N126);
nand NAND3 (N825, N809, N219, N548);
nor NOR2 (N826, N810, N714);
nand NAND3 (N827, N825, N768, N583);
nor NOR2 (N828, N816, N730);
xor XOR2 (N829, N821, N556);
or OR2 (N830, N829, N511);
nand NAND4 (N831, N826, N803, N45, N729);
nor NOR3 (N832, N824, N370, N85);
and AND3 (N833, N822, N764, N816);
xor XOR2 (N834, N830, N811);
nand NAND2 (N835, N834, N784);
not NOT1 (N836, N835);
or OR4 (N837, N827, N148, N497, N63);
xor XOR2 (N838, N791, N112);
not NOT1 (N839, N832);
buf BUF1 (N840, N831);
and AND2 (N841, N840, N699);
not NOT1 (N842, N838);
nand NAND4 (N843, N839, N395, N77, N137);
nand NAND3 (N844, N841, N579, N183);
buf BUF1 (N845, N820);
or OR2 (N846, N845, N397);
xor XOR2 (N847, N836, N735);
nor NOR2 (N848, N843, N794);
nor NOR3 (N849, N844, N108, N330);
and AND3 (N850, N842, N498, N747);
and AND2 (N851, N850, N758);
or OR3 (N852, N848, N734, N704);
or OR2 (N853, N849, N610);
not NOT1 (N854, N853);
not NOT1 (N855, N837);
nor NOR2 (N856, N851, N175);
not NOT1 (N857, N819);
nor NOR4 (N858, N854, N373, N558, N828);
buf BUF1 (N859, N341);
and AND2 (N860, N856, N227);
nor NOR3 (N861, N858, N806, N745);
buf BUF1 (N862, N833);
and AND3 (N863, N823, N226, N242);
buf BUF1 (N864, N857);
xor XOR2 (N865, N861, N791);
nand NAND4 (N866, N855, N93, N17, N498);
or OR2 (N867, N865, N116);
nor NOR3 (N868, N847, N136, N274);
xor XOR2 (N869, N864, N517);
not NOT1 (N870, N867);
or OR2 (N871, N868, N471);
nor NOR3 (N872, N860, N870, N791);
nor NOR2 (N873, N62, N362);
and AND4 (N874, N862, N496, N850, N542);
nand NAND3 (N875, N873, N459, N719);
nand NAND3 (N876, N872, N123, N679);
or OR4 (N877, N846, N177, N20, N847);
nor NOR4 (N878, N869, N587, N629, N229);
not NOT1 (N879, N859);
nor NOR2 (N880, N875, N461);
not NOT1 (N881, N863);
nand NAND2 (N882, N866, N860);
nor NOR2 (N883, N881, N200);
buf BUF1 (N884, N882);
buf BUF1 (N885, N878);
or OR4 (N886, N884, N142, N475, N431);
nand NAND2 (N887, N874, N201);
nand NAND4 (N888, N885, N19, N287, N777);
nor NOR2 (N889, N888, N321);
not NOT1 (N890, N852);
buf BUF1 (N891, N890);
nand NAND3 (N892, N891, N818, N787);
nor NOR3 (N893, N871, N419, N217);
nor NOR2 (N894, N893, N228);
xor XOR2 (N895, N880, N89);
or OR4 (N896, N877, N18, N736, N456);
xor XOR2 (N897, N886, N855);
nor NOR4 (N898, N876, N281, N87, N694);
xor XOR2 (N899, N895, N530);
nand NAND3 (N900, N889, N615, N417);
not NOT1 (N901, N892);
buf BUF1 (N902, N896);
nand NAND3 (N903, N894, N169, N384);
or OR2 (N904, N887, N882);
and AND2 (N905, N902, N438);
and AND4 (N906, N897, N394, N587, N234);
buf BUF1 (N907, N898);
and AND4 (N908, N904, N292, N571, N797);
buf BUF1 (N909, N883);
nand NAND3 (N910, N899, N657, N626);
xor XOR2 (N911, N879, N638);
and AND3 (N912, N901, N787, N686);
nor NOR4 (N913, N911, N37, N157, N23);
nand NAND3 (N914, N913, N534, N463);
buf BUF1 (N915, N907);
and AND2 (N916, N908, N593);
nand NAND2 (N917, N916, N512);
nor NOR3 (N918, N905, N432, N737);
and AND2 (N919, N910, N720);
not NOT1 (N920, N912);
buf BUF1 (N921, N914);
buf BUF1 (N922, N903);
not NOT1 (N923, N906);
nand NAND2 (N924, N923, N835);
xor XOR2 (N925, N917, N515);
or OR3 (N926, N920, N54, N33);
nand NAND2 (N927, N909, N500);
not NOT1 (N928, N915);
not NOT1 (N929, N924);
nand NAND3 (N930, N919, N224, N774);
nor NOR4 (N931, N921, N772, N73, N508);
nand NAND2 (N932, N931, N620);
and AND4 (N933, N926, N461, N467, N350);
nand NAND4 (N934, N927, N478, N405, N647);
buf BUF1 (N935, N922);
not NOT1 (N936, N933);
nor NOR3 (N937, N929, N770, N225);
or OR3 (N938, N932, N68, N792);
nand NAND3 (N939, N936, N691, N515);
nand NAND3 (N940, N928, N164, N894);
nand NAND4 (N941, N939, N745, N633, N709);
buf BUF1 (N942, N938);
buf BUF1 (N943, N940);
not NOT1 (N944, N937);
or OR4 (N945, N941, N540, N139, N738);
xor XOR2 (N946, N944, N280);
nor NOR3 (N947, N945, N873, N70);
xor XOR2 (N948, N946, N198);
and AND2 (N949, N947, N204);
buf BUF1 (N950, N934);
nor NOR3 (N951, N918, N640, N571);
not NOT1 (N952, N900);
nor NOR2 (N953, N949, N68);
and AND3 (N954, N943, N918, N126);
not NOT1 (N955, N935);
nor NOR4 (N956, N925, N709, N5, N289);
not NOT1 (N957, N955);
xor XOR2 (N958, N930, N812);
and AND4 (N959, N948, N776, N649, N860);
nand NAND4 (N960, N958, N109, N561, N242);
not NOT1 (N961, N942);
nor NOR2 (N962, N953, N569);
buf BUF1 (N963, N951);
or OR2 (N964, N961, N363);
buf BUF1 (N965, N959);
xor XOR2 (N966, N960, N428);
not NOT1 (N967, N963);
and AND2 (N968, N957, N443);
buf BUF1 (N969, N965);
buf BUF1 (N970, N967);
not NOT1 (N971, N969);
or OR3 (N972, N971, N724, N205);
not NOT1 (N973, N956);
nand NAND2 (N974, N968, N241);
or OR4 (N975, N974, N211, N168, N29);
nand NAND4 (N976, N966, N356, N598, N916);
and AND4 (N977, N972, N199, N345, N510);
and AND4 (N978, N970, N585, N647, N282);
nor NOR2 (N979, N977, N670);
and AND4 (N980, N964, N682, N628, N529);
or OR4 (N981, N952, N606, N499, N696);
not NOT1 (N982, N980);
buf BUF1 (N983, N950);
or OR4 (N984, N983, N887, N512, N656);
not NOT1 (N985, N981);
buf BUF1 (N986, N982);
buf BUF1 (N987, N979);
xor XOR2 (N988, N976, N38);
or OR4 (N989, N988, N636, N789, N746);
not NOT1 (N990, N987);
buf BUF1 (N991, N990);
not NOT1 (N992, N973);
nor NOR2 (N993, N975, N385);
not NOT1 (N994, N962);
nor NOR2 (N995, N994, N67);
nand NAND3 (N996, N995, N5, N426);
nor NOR3 (N997, N993, N873, N815);
and AND3 (N998, N989, N758, N42);
nor NOR2 (N999, N984, N413);
or OR3 (N1000, N985, N339, N752);
nand NAND3 (N1001, N954, N804, N513);
xor XOR2 (N1002, N986, N392);
nand NAND3 (N1003, N992, N193, N123);
or OR2 (N1004, N978, N959);
nor NOR3 (N1005, N1002, N706, N631);
and AND4 (N1006, N998, N793, N107, N566);
nand NAND4 (N1007, N1000, N738, N729, N793);
buf BUF1 (N1008, N1001);
nor NOR2 (N1009, N1004, N375);
xor XOR2 (N1010, N1008, N739);
and AND4 (N1011, N1003, N806, N472, N391);
nand NAND4 (N1012, N996, N773, N806, N684);
nand NAND4 (N1013, N1011, N1002, N648, N827);
nor NOR2 (N1014, N1009, N423);
nand NAND3 (N1015, N1014, N599, N784);
buf BUF1 (N1016, N1006);
xor XOR2 (N1017, N997, N152);
and AND3 (N1018, N1012, N693, N939);
nand NAND3 (N1019, N1016, N521, N960);
not NOT1 (N1020, N1018);
buf BUF1 (N1021, N991);
or OR3 (N1022, N1005, N609, N698);
buf BUF1 (N1023, N1017);
nand NAND2 (N1024, N1022, N523);
xor XOR2 (N1025, N1007, N175);
nand NAND2 (N1026, N1021, N184);
nand NAND4 (N1027, N1023, N583, N149, N225);
nor NOR2 (N1028, N1026, N787);
nor NOR2 (N1029, N1010, N385);
nor NOR4 (N1030, N1020, N549, N783, N894);
nand NAND3 (N1031, N1015, N327, N192);
buf BUF1 (N1032, N1029);
not NOT1 (N1033, N1024);
and AND2 (N1034, N1027, N846);
xor XOR2 (N1035, N1033, N347);
nand NAND2 (N1036, N1034, N819);
xor XOR2 (N1037, N1028, N431);
or OR3 (N1038, N1036, N578, N602);
nor NOR3 (N1039, N1031, N753, N626);
and AND4 (N1040, N1032, N57, N933, N102);
nor NOR4 (N1041, N1037, N192, N749, N728);
nor NOR4 (N1042, N1039, N208, N530, N673);
nor NOR4 (N1043, N1013, N491, N128, N548);
nand NAND4 (N1044, N1019, N594, N893, N176);
buf BUF1 (N1045, N1038);
nor NOR3 (N1046, N1041, N899, N161);
buf BUF1 (N1047, N1035);
nor NOR3 (N1048, N1047, N98, N593);
not NOT1 (N1049, N1043);
and AND2 (N1050, N1049, N375);
nand NAND3 (N1051, N1025, N907, N690);
xor XOR2 (N1052, N1042, N489);
nor NOR2 (N1053, N1046, N525);
buf BUF1 (N1054, N1044);
xor XOR2 (N1055, N1045, N788);
buf BUF1 (N1056, N1048);
and AND4 (N1057, N999, N331, N130, N439);
nand NAND4 (N1058, N1055, N459, N387, N919);
or OR4 (N1059, N1056, N1032, N836, N784);
nor NOR2 (N1060, N1040, N828);
or OR3 (N1061, N1057, N55, N171);
nand NAND2 (N1062, N1059, N531);
nor NOR4 (N1063, N1050, N926, N29, N133);
and AND2 (N1064, N1061, N214);
xor XOR2 (N1065, N1054, N717);
xor XOR2 (N1066, N1058, N551);
nand NAND4 (N1067, N1062, N153, N337, N891);
buf BUF1 (N1068, N1051);
nor NOR4 (N1069, N1063, N229, N519, N398);
nand NAND2 (N1070, N1060, N783);
not NOT1 (N1071, N1069);
and AND2 (N1072, N1067, N505);
not NOT1 (N1073, N1072);
nand NAND2 (N1074, N1053, N784);
not NOT1 (N1075, N1065);
nor NOR4 (N1076, N1030, N897, N152, N442);
nor NOR4 (N1077, N1066, N211, N126, N746);
nor NOR3 (N1078, N1076, N246, N990);
or OR3 (N1079, N1077, N461, N381);
buf BUF1 (N1080, N1071);
nand NAND3 (N1081, N1073, N736, N278);
and AND4 (N1082, N1070, N335, N444, N441);
not NOT1 (N1083, N1078);
xor XOR2 (N1084, N1079, N488);
not NOT1 (N1085, N1084);
and AND4 (N1086, N1082, N351, N725, N340);
xor XOR2 (N1087, N1052, N140);
nand NAND3 (N1088, N1083, N879, N685);
and AND2 (N1089, N1081, N718);
nor NOR2 (N1090, N1089, N796);
not NOT1 (N1091, N1068);
or OR2 (N1092, N1080, N71);
xor XOR2 (N1093, N1064, N844);
xor XOR2 (N1094, N1075, N461);
and AND3 (N1095, N1074, N741, N423);
nor NOR3 (N1096, N1090, N1020, N737);
nor NOR3 (N1097, N1087, N430, N851);
nand NAND2 (N1098, N1092, N621);
not NOT1 (N1099, N1086);
nand NAND4 (N1100, N1099, N110, N409, N186);
not NOT1 (N1101, N1085);
nor NOR4 (N1102, N1100, N675, N128, N840);
xor XOR2 (N1103, N1098, N459);
xor XOR2 (N1104, N1102, N890);
buf BUF1 (N1105, N1096);
nand NAND3 (N1106, N1104, N285, N841);
buf BUF1 (N1107, N1094);
nand NAND2 (N1108, N1103, N400);
nor NOR2 (N1109, N1108, N1060);
buf BUF1 (N1110, N1106);
buf BUF1 (N1111, N1101);
nor NOR3 (N1112, N1095, N774, N686);
nand NAND4 (N1113, N1091, N796, N876, N18);
xor XOR2 (N1114, N1097, N467);
buf BUF1 (N1115, N1113);
not NOT1 (N1116, N1115);
xor XOR2 (N1117, N1105, N589);
nand NAND2 (N1118, N1111, N241);
buf BUF1 (N1119, N1088);
not NOT1 (N1120, N1093);
nor NOR3 (N1121, N1118, N505, N357);
nor NOR3 (N1122, N1107, N771, N562);
xor XOR2 (N1123, N1121, N1076);
buf BUF1 (N1124, N1117);
or OR2 (N1125, N1120, N271);
nor NOR2 (N1126, N1114, N795);
not NOT1 (N1127, N1123);
or OR2 (N1128, N1112, N986);
xor XOR2 (N1129, N1127, N976);
or OR3 (N1130, N1126, N773, N892);
xor XOR2 (N1131, N1130, N1050);
buf BUF1 (N1132, N1131);
and AND4 (N1133, N1132, N753, N939, N178);
or OR2 (N1134, N1125, N517);
nor NOR2 (N1135, N1109, N549);
xor XOR2 (N1136, N1122, N207);
nor NOR4 (N1137, N1134, N798, N744, N451);
xor XOR2 (N1138, N1128, N240);
and AND3 (N1139, N1135, N990, N444);
nand NAND2 (N1140, N1136, N359);
xor XOR2 (N1141, N1133, N982);
buf BUF1 (N1142, N1139);
buf BUF1 (N1143, N1137);
not NOT1 (N1144, N1129);
and AND3 (N1145, N1141, N173, N1125);
xor XOR2 (N1146, N1140, N624);
or OR2 (N1147, N1110, N347);
not NOT1 (N1148, N1147);
and AND4 (N1149, N1148, N541, N117, N609);
or OR2 (N1150, N1119, N533);
not NOT1 (N1151, N1145);
or OR3 (N1152, N1149, N1034, N166);
nand NAND3 (N1153, N1116, N13, N1042);
nand NAND3 (N1154, N1143, N843, N981);
or OR4 (N1155, N1142, N534, N300, N818);
or OR3 (N1156, N1124, N211, N1142);
xor XOR2 (N1157, N1144, N150);
xor XOR2 (N1158, N1138, N212);
not NOT1 (N1159, N1154);
not NOT1 (N1160, N1155);
and AND3 (N1161, N1150, N260, N524);
not NOT1 (N1162, N1151);
and AND2 (N1163, N1162, N584);
buf BUF1 (N1164, N1158);
buf BUF1 (N1165, N1152);
buf BUF1 (N1166, N1161);
nor NOR4 (N1167, N1146, N299, N95, N445);
not NOT1 (N1168, N1165);
xor XOR2 (N1169, N1164, N821);
not NOT1 (N1170, N1169);
buf BUF1 (N1171, N1153);
xor XOR2 (N1172, N1163, N293);
not NOT1 (N1173, N1166);
or OR3 (N1174, N1168, N818, N70);
nor NOR2 (N1175, N1173, N337);
nor NOR3 (N1176, N1159, N55, N1072);
and AND3 (N1177, N1156, N275, N406);
and AND2 (N1178, N1167, N1035);
xor XOR2 (N1179, N1171, N147);
and AND4 (N1180, N1178, N723, N1126, N418);
xor XOR2 (N1181, N1180, N309);
xor XOR2 (N1182, N1175, N24);
nand NAND4 (N1183, N1172, N352, N804, N294);
xor XOR2 (N1184, N1160, N439);
or OR4 (N1185, N1157, N634, N1164, N235);
or OR3 (N1186, N1174, N863, N905);
and AND3 (N1187, N1184, N1002, N931);
nand NAND2 (N1188, N1181, N1117);
xor XOR2 (N1189, N1187, N355);
buf BUF1 (N1190, N1177);
nor NOR3 (N1191, N1189, N507, N458);
buf BUF1 (N1192, N1182);
nand NAND2 (N1193, N1192, N898);
and AND4 (N1194, N1170, N899, N475, N360);
or OR3 (N1195, N1194, N550, N473);
nand NAND2 (N1196, N1185, N163);
and AND2 (N1197, N1195, N246);
not NOT1 (N1198, N1190);
xor XOR2 (N1199, N1198, N65);
nor NOR3 (N1200, N1176, N843, N74);
and AND4 (N1201, N1193, N414, N1062, N795);
and AND2 (N1202, N1191, N500);
and AND4 (N1203, N1179, N623, N748, N964);
xor XOR2 (N1204, N1203, N134);
nor NOR4 (N1205, N1201, N72, N505, N1183);
buf BUF1 (N1206, N1153);
not NOT1 (N1207, N1199);
buf BUF1 (N1208, N1205);
buf BUF1 (N1209, N1188);
nand NAND2 (N1210, N1206, N397);
buf BUF1 (N1211, N1186);
xor XOR2 (N1212, N1211, N33);
nor NOR4 (N1213, N1204, N380, N1047, N92);
nor NOR2 (N1214, N1209, N1030);
nor NOR3 (N1215, N1196, N282, N935);
not NOT1 (N1216, N1202);
nand NAND3 (N1217, N1207, N791, N698);
nor NOR3 (N1218, N1216, N643, N461);
buf BUF1 (N1219, N1212);
not NOT1 (N1220, N1210);
not NOT1 (N1221, N1213);
xor XOR2 (N1222, N1217, N917);
and AND2 (N1223, N1197, N1183);
nor NOR2 (N1224, N1219, N344);
buf BUF1 (N1225, N1215);
xor XOR2 (N1226, N1200, N643);
and AND4 (N1227, N1226, N1041, N416, N663);
buf BUF1 (N1228, N1225);
nor NOR3 (N1229, N1223, N953, N354);
buf BUF1 (N1230, N1229);
xor XOR2 (N1231, N1230, N665);
xor XOR2 (N1232, N1221, N686);
xor XOR2 (N1233, N1227, N164);
not NOT1 (N1234, N1218);
xor XOR2 (N1235, N1224, N1066);
and AND2 (N1236, N1232, N456);
nand NAND4 (N1237, N1233, N1104, N1182, N534);
not NOT1 (N1238, N1220);
and AND4 (N1239, N1222, N1137, N320, N870);
nand NAND4 (N1240, N1234, N1227, N183, N799);
or OR3 (N1241, N1214, N1084, N171);
nand NAND4 (N1242, N1228, N589, N664, N670);
and AND2 (N1243, N1242, N653);
buf BUF1 (N1244, N1235);
nor NOR3 (N1245, N1244, N270, N1136);
nor NOR2 (N1246, N1241, N354);
nand NAND2 (N1247, N1245, N1121);
nand NAND4 (N1248, N1246, N160, N718, N540);
not NOT1 (N1249, N1239);
buf BUF1 (N1250, N1243);
or OR2 (N1251, N1249, N814);
and AND2 (N1252, N1247, N970);
nand NAND2 (N1253, N1251, N116);
nor NOR3 (N1254, N1250, N830, N510);
not NOT1 (N1255, N1254);
and AND2 (N1256, N1253, N645);
buf BUF1 (N1257, N1240);
or OR2 (N1258, N1238, N918);
and AND4 (N1259, N1236, N352, N549, N574);
nand NAND4 (N1260, N1208, N797, N221, N1198);
buf BUF1 (N1261, N1257);
nor NOR2 (N1262, N1248, N1133);
not NOT1 (N1263, N1237);
nand NAND2 (N1264, N1258, N152);
nand NAND4 (N1265, N1264, N205, N1153, N703);
nand NAND2 (N1266, N1262, N800);
xor XOR2 (N1267, N1252, N1088);
or OR4 (N1268, N1231, N1228, N489, N1161);
nand NAND4 (N1269, N1265, N879, N259, N923);
or OR4 (N1270, N1267, N522, N303, N1098);
xor XOR2 (N1271, N1263, N293);
buf BUF1 (N1272, N1256);
nor NOR2 (N1273, N1269, N332);
nand NAND3 (N1274, N1259, N1164, N1210);
nand NAND3 (N1275, N1273, N1212, N914);
xor XOR2 (N1276, N1261, N439);
and AND4 (N1277, N1266, N776, N86, N9);
xor XOR2 (N1278, N1275, N272);
and AND2 (N1279, N1272, N152);
nor NOR2 (N1280, N1271, N543);
not NOT1 (N1281, N1279);
buf BUF1 (N1282, N1281);
and AND2 (N1283, N1278, N91);
not NOT1 (N1284, N1270);
not NOT1 (N1285, N1274);
nor NOR2 (N1286, N1280, N60);
and AND3 (N1287, N1260, N808, N957);
and AND3 (N1288, N1276, N1212, N222);
nor NOR3 (N1289, N1287, N328, N1264);
or OR2 (N1290, N1268, N130);
and AND3 (N1291, N1277, N515, N456);
buf BUF1 (N1292, N1291);
buf BUF1 (N1293, N1282);
xor XOR2 (N1294, N1284, N66);
xor XOR2 (N1295, N1290, N1281);
not NOT1 (N1296, N1288);
buf BUF1 (N1297, N1293);
buf BUF1 (N1298, N1296);
xor XOR2 (N1299, N1285, N1133);
nor NOR3 (N1300, N1294, N444, N62);
or OR4 (N1301, N1297, N741, N535, N1216);
nor NOR3 (N1302, N1286, N712, N320);
buf BUF1 (N1303, N1292);
buf BUF1 (N1304, N1283);
and AND3 (N1305, N1299, N592, N304);
or OR2 (N1306, N1298, N450);
or OR4 (N1307, N1302, N434, N913, N77);
nand NAND2 (N1308, N1303, N19);
buf BUF1 (N1309, N1301);
xor XOR2 (N1310, N1308, N1132);
and AND4 (N1311, N1289, N798, N871, N242);
not NOT1 (N1312, N1309);
or OR4 (N1313, N1306, N820, N829, N346);
xor XOR2 (N1314, N1307, N213);
or OR4 (N1315, N1305, N761, N241, N680);
nand NAND2 (N1316, N1310, N140);
not NOT1 (N1317, N1312);
xor XOR2 (N1318, N1311, N1177);
not NOT1 (N1319, N1295);
xor XOR2 (N1320, N1304, N726);
nor NOR4 (N1321, N1313, N106, N565, N268);
nor NOR2 (N1322, N1314, N71);
not NOT1 (N1323, N1316);
nor NOR2 (N1324, N1319, N616);
or OR4 (N1325, N1321, N470, N676, N634);
not NOT1 (N1326, N1323);
xor XOR2 (N1327, N1300, N99);
or OR3 (N1328, N1326, N729, N1001);
not NOT1 (N1329, N1315);
nor NOR2 (N1330, N1317, N922);
nand NAND2 (N1331, N1328, N983);
and AND2 (N1332, N1255, N273);
xor XOR2 (N1333, N1330, N959);
or OR4 (N1334, N1332, N730, N391, N806);
not NOT1 (N1335, N1318);
and AND3 (N1336, N1324, N54, N1081);
xor XOR2 (N1337, N1327, N602);
xor XOR2 (N1338, N1320, N1311);
or OR3 (N1339, N1336, N249, N36);
buf BUF1 (N1340, N1331);
xor XOR2 (N1341, N1335, N1005);
nand NAND4 (N1342, N1334, N895, N309, N847);
not NOT1 (N1343, N1341);
nand NAND4 (N1344, N1329, N825, N771, N521);
or OR4 (N1345, N1337, N1056, N1041, N784);
nor NOR4 (N1346, N1322, N174, N556, N514);
xor XOR2 (N1347, N1340, N22);
buf BUF1 (N1348, N1347);
or OR2 (N1349, N1333, N93);
buf BUF1 (N1350, N1345);
nor NOR3 (N1351, N1339, N1173, N1008);
nand NAND3 (N1352, N1350, N344, N784);
nor NOR3 (N1353, N1348, N1155, N1058);
and AND2 (N1354, N1325, N632);
xor XOR2 (N1355, N1342, N915);
xor XOR2 (N1356, N1353, N885);
nand NAND2 (N1357, N1338, N723);
buf BUF1 (N1358, N1357);
not NOT1 (N1359, N1343);
nand NAND2 (N1360, N1351, N745);
and AND2 (N1361, N1346, N995);
buf BUF1 (N1362, N1361);
not NOT1 (N1363, N1344);
not NOT1 (N1364, N1362);
nor NOR4 (N1365, N1359, N731, N88, N764);
xor XOR2 (N1366, N1352, N29);
xor XOR2 (N1367, N1355, N355);
buf BUF1 (N1368, N1365);
not NOT1 (N1369, N1358);
or OR2 (N1370, N1349, N253);
xor XOR2 (N1371, N1369, N186);
and AND4 (N1372, N1368, N234, N575, N1082);
nand NAND2 (N1373, N1367, N357);
buf BUF1 (N1374, N1356);
buf BUF1 (N1375, N1360);
not NOT1 (N1376, N1373);
and AND3 (N1377, N1374, N1252, N1171);
or OR4 (N1378, N1372, N1149, N17, N1353);
and AND4 (N1379, N1375, N359, N607, N927);
nor NOR4 (N1380, N1379, N1331, N475, N785);
and AND4 (N1381, N1371, N1082, N294, N813);
nor NOR4 (N1382, N1370, N237, N852, N979);
and AND3 (N1383, N1380, N1304, N171);
xor XOR2 (N1384, N1381, N1333);
or OR2 (N1385, N1384, N516);
nand NAND2 (N1386, N1366, N77);
and AND3 (N1387, N1385, N838, N807);
xor XOR2 (N1388, N1382, N803);
or OR3 (N1389, N1386, N518, N646);
and AND3 (N1390, N1354, N88, N38);
nor NOR2 (N1391, N1389, N1133);
buf BUF1 (N1392, N1388);
not NOT1 (N1393, N1377);
nand NAND3 (N1394, N1363, N260, N379);
or OR2 (N1395, N1390, N562);
and AND4 (N1396, N1364, N1176, N932, N1314);
or OR3 (N1397, N1396, N252, N1235);
nand NAND2 (N1398, N1378, N1325);
not NOT1 (N1399, N1376);
buf BUF1 (N1400, N1392);
or OR3 (N1401, N1383, N171, N32);
nor NOR2 (N1402, N1397, N492);
and AND2 (N1403, N1393, N518);
nand NAND4 (N1404, N1395, N240, N57, N575);
or OR3 (N1405, N1391, N528, N494);
or OR4 (N1406, N1403, N872, N1275, N483);
xor XOR2 (N1407, N1394, N991);
not NOT1 (N1408, N1400);
buf BUF1 (N1409, N1407);
nand NAND3 (N1410, N1399, N1077, N1128);
not NOT1 (N1411, N1402);
and AND2 (N1412, N1411, N1272);
nor NOR2 (N1413, N1401, N261);
xor XOR2 (N1414, N1412, N1320);
not NOT1 (N1415, N1408);
not NOT1 (N1416, N1414);
xor XOR2 (N1417, N1398, N1391);
not NOT1 (N1418, N1415);
nand NAND2 (N1419, N1404, N1110);
and AND3 (N1420, N1413, N740, N499);
nand NAND4 (N1421, N1405, N317, N617, N195);
or OR2 (N1422, N1418, N88);
nor NOR3 (N1423, N1419, N937, N449);
xor XOR2 (N1424, N1387, N605);
nor NOR3 (N1425, N1421, N911, N11);
and AND4 (N1426, N1417, N725, N123, N1177);
buf BUF1 (N1427, N1422);
and AND2 (N1428, N1425, N244);
nand NAND2 (N1429, N1428, N211);
nand NAND2 (N1430, N1429, N245);
buf BUF1 (N1431, N1423);
buf BUF1 (N1432, N1416);
nand NAND2 (N1433, N1426, N774);
xor XOR2 (N1434, N1424, N1122);
xor XOR2 (N1435, N1430, N214);
buf BUF1 (N1436, N1434);
and AND2 (N1437, N1432, N541);
nand NAND2 (N1438, N1410, N471);
or OR2 (N1439, N1437, N847);
not NOT1 (N1440, N1436);
xor XOR2 (N1441, N1406, N536);
or OR2 (N1442, N1438, N889);
nand NAND4 (N1443, N1409, N1174, N699, N996);
buf BUF1 (N1444, N1427);
xor XOR2 (N1445, N1440, N488);
or OR3 (N1446, N1431, N1010, N1433);
nor NOR4 (N1447, N781, N903, N625, N552);
not NOT1 (N1448, N1447);
and AND2 (N1449, N1439, N566);
nand NAND3 (N1450, N1448, N512, N559);
and AND4 (N1451, N1420, N196, N851, N1360);
and AND3 (N1452, N1450, N76, N845);
not NOT1 (N1453, N1446);
not NOT1 (N1454, N1449);
not NOT1 (N1455, N1453);
and AND2 (N1456, N1442, N876);
buf BUF1 (N1457, N1454);
nor NOR4 (N1458, N1435, N1190, N1041, N988);
and AND4 (N1459, N1452, N688, N1284, N1393);
nor NOR4 (N1460, N1457, N340, N1015, N700);
nor NOR4 (N1461, N1455, N572, N1294, N1005);
or OR4 (N1462, N1443, N599, N124, N222);
nor NOR2 (N1463, N1461, N505);
nand NAND4 (N1464, N1460, N1334, N679, N550);
or OR4 (N1465, N1463, N1036, N889, N1122);
buf BUF1 (N1466, N1444);
or OR3 (N1467, N1464, N932, N772);
nor NOR3 (N1468, N1467, N1013, N464);
and AND4 (N1469, N1441, N1060, N795, N1023);
and AND4 (N1470, N1465, N1357, N68, N401);
nor NOR2 (N1471, N1456, N644);
buf BUF1 (N1472, N1459);
xor XOR2 (N1473, N1445, N777);
and AND4 (N1474, N1462, N538, N1152, N548);
and AND4 (N1475, N1473, N388, N1341, N1161);
or OR3 (N1476, N1475, N277, N1102);
and AND4 (N1477, N1476, N1111, N804, N1088);
nand NAND4 (N1478, N1451, N471, N283, N258);
buf BUF1 (N1479, N1474);
xor XOR2 (N1480, N1471, N45);
or OR2 (N1481, N1472, N465);
nand NAND4 (N1482, N1477, N1372, N1252, N988);
and AND2 (N1483, N1458, N1465);
nand NAND2 (N1484, N1480, N629);
nor NOR2 (N1485, N1482, N1452);
not NOT1 (N1486, N1478);
xor XOR2 (N1487, N1466, N1185);
not NOT1 (N1488, N1487);
buf BUF1 (N1489, N1479);
buf BUF1 (N1490, N1486);
xor XOR2 (N1491, N1481, N138);
nor NOR3 (N1492, N1488, N179, N1343);
buf BUF1 (N1493, N1485);
buf BUF1 (N1494, N1470);
and AND3 (N1495, N1483, N13, N341);
xor XOR2 (N1496, N1493, N855);
xor XOR2 (N1497, N1468, N1308);
nor NOR3 (N1498, N1489, N1453, N1377);
and AND4 (N1499, N1491, N1289, N617, N1408);
and AND4 (N1500, N1497, N537, N1082, N1214);
xor XOR2 (N1501, N1484, N1109);
buf BUF1 (N1502, N1492);
nand NAND4 (N1503, N1496, N522, N163, N496);
buf BUF1 (N1504, N1495);
nor NOR3 (N1505, N1501, N227, N74);
not NOT1 (N1506, N1500);
not NOT1 (N1507, N1505);
nor NOR3 (N1508, N1498, N1370, N673);
or OR3 (N1509, N1503, N165, N411);
and AND2 (N1510, N1502, N303);
nor NOR2 (N1511, N1499, N1302);
not NOT1 (N1512, N1510);
xor XOR2 (N1513, N1490, N491);
or OR2 (N1514, N1513, N1173);
and AND3 (N1515, N1511, N765, N998);
xor XOR2 (N1516, N1509, N1092);
nand NAND4 (N1517, N1508, N1347, N377, N965);
nand NAND3 (N1518, N1517, N1185, N160);
nor NOR3 (N1519, N1469, N1397, N600);
xor XOR2 (N1520, N1506, N821);
not NOT1 (N1521, N1518);
or OR3 (N1522, N1516, N1357, N679);
nand NAND3 (N1523, N1514, N1356, N707);
nor NOR3 (N1524, N1515, N754, N1391);
nand NAND4 (N1525, N1494, N756, N485, N456);
or OR3 (N1526, N1504, N172, N1436);
not NOT1 (N1527, N1526);
not NOT1 (N1528, N1524);
nand NAND3 (N1529, N1507, N1229, N309);
nand NAND2 (N1530, N1523, N825);
xor XOR2 (N1531, N1530, N877);
nor NOR4 (N1532, N1520, N737, N1354, N1365);
or OR4 (N1533, N1512, N73, N1338, N1446);
not NOT1 (N1534, N1531);
not NOT1 (N1535, N1521);
and AND4 (N1536, N1519, N1139, N205, N84);
not NOT1 (N1537, N1534);
buf BUF1 (N1538, N1529);
and AND3 (N1539, N1537, N37, N456);
and AND4 (N1540, N1538, N924, N134, N283);
or OR4 (N1541, N1532, N482, N814, N23);
nand NAND2 (N1542, N1522, N633);
or OR4 (N1543, N1540, N1401, N666, N1367);
or OR4 (N1544, N1525, N817, N626, N1474);
buf BUF1 (N1545, N1528);
xor XOR2 (N1546, N1533, N431);
nand NAND3 (N1547, N1542, N291, N1330);
buf BUF1 (N1548, N1544);
and AND2 (N1549, N1536, N1159);
buf BUF1 (N1550, N1543);
xor XOR2 (N1551, N1546, N48);
and AND3 (N1552, N1548, N611, N109);
and AND3 (N1553, N1541, N897, N1423);
and AND2 (N1554, N1551, N58);
buf BUF1 (N1555, N1539);
xor XOR2 (N1556, N1554, N211);
nand NAND2 (N1557, N1527, N1241);
xor XOR2 (N1558, N1553, N273);
or OR2 (N1559, N1550, N185);
nand NAND3 (N1560, N1547, N49, N199);
nand NAND4 (N1561, N1549, N715, N724, N1329);
nand NAND2 (N1562, N1556, N1082);
and AND4 (N1563, N1555, N1149, N213, N66);
buf BUF1 (N1564, N1558);
and AND4 (N1565, N1557, N194, N477, N320);
buf BUF1 (N1566, N1563);
or OR3 (N1567, N1560, N1166, N956);
nand NAND4 (N1568, N1535, N1304, N1153, N745);
and AND3 (N1569, N1566, N397, N492);
not NOT1 (N1570, N1568);
buf BUF1 (N1571, N1561);
not NOT1 (N1572, N1564);
nor NOR2 (N1573, N1567, N162);
nor NOR2 (N1574, N1573, N1320);
nand NAND2 (N1575, N1552, N352);
not NOT1 (N1576, N1545);
nor NOR3 (N1577, N1576, N695, N1161);
or OR3 (N1578, N1565, N293, N1038);
buf BUF1 (N1579, N1562);
xor XOR2 (N1580, N1577, N722);
not NOT1 (N1581, N1572);
xor XOR2 (N1582, N1581, N678);
and AND4 (N1583, N1569, N1347, N271, N962);
and AND4 (N1584, N1559, N414, N715, N528);
xor XOR2 (N1585, N1579, N349);
xor XOR2 (N1586, N1584, N503);
nand NAND2 (N1587, N1574, N1399);
nand NAND3 (N1588, N1571, N637, N751);
nor NOR4 (N1589, N1575, N497, N1358, N826);
nor NOR2 (N1590, N1587, N258);
nor NOR2 (N1591, N1570, N1500);
or OR3 (N1592, N1583, N818, N507);
xor XOR2 (N1593, N1590, N1590);
and AND2 (N1594, N1580, N179);
nand NAND2 (N1595, N1594, N870);
nand NAND4 (N1596, N1593, N879, N156, N494);
and AND2 (N1597, N1591, N1253);
xor XOR2 (N1598, N1597, N985);
and AND3 (N1599, N1588, N616, N488);
or OR2 (N1600, N1586, N583);
xor XOR2 (N1601, N1599, N1579);
buf BUF1 (N1602, N1578);
buf BUF1 (N1603, N1601);
xor XOR2 (N1604, N1582, N745);
xor XOR2 (N1605, N1602, N1494);
nand NAND3 (N1606, N1604, N819, N967);
or OR2 (N1607, N1603, N840);
not NOT1 (N1608, N1598);
buf BUF1 (N1609, N1607);
nor NOR3 (N1610, N1605, N140, N1109);
xor XOR2 (N1611, N1595, N711);
xor XOR2 (N1612, N1600, N1579);
and AND2 (N1613, N1589, N606);
buf BUF1 (N1614, N1592);
nor NOR2 (N1615, N1609, N956);
nand NAND3 (N1616, N1608, N932, N1497);
nor NOR4 (N1617, N1585, N929, N216, N974);
or OR2 (N1618, N1612, N799);
not NOT1 (N1619, N1617);
and AND4 (N1620, N1610, N1103, N851, N1328);
nor NOR3 (N1621, N1614, N1452, N745);
nand NAND4 (N1622, N1613, N1031, N483, N375);
xor XOR2 (N1623, N1621, N603);
or OR3 (N1624, N1606, N789, N821);
not NOT1 (N1625, N1615);
not NOT1 (N1626, N1624);
buf BUF1 (N1627, N1626);
buf BUF1 (N1628, N1616);
not NOT1 (N1629, N1628);
xor XOR2 (N1630, N1623, N608);
and AND2 (N1631, N1622, N682);
xor XOR2 (N1632, N1618, N1502);
xor XOR2 (N1633, N1596, N230);
buf BUF1 (N1634, N1629);
xor XOR2 (N1635, N1634, N1036);
nor NOR3 (N1636, N1631, N392, N7);
xor XOR2 (N1637, N1630, N1340);
nor NOR4 (N1638, N1637, N839, N650, N1528);
and AND3 (N1639, N1633, N1532, N1305);
nand NAND4 (N1640, N1611, N750, N847, N1207);
and AND3 (N1641, N1625, N872, N555);
nor NOR2 (N1642, N1638, N1266);
buf BUF1 (N1643, N1635);
not NOT1 (N1644, N1639);
and AND3 (N1645, N1627, N169, N114);
xor XOR2 (N1646, N1620, N959);
or OR2 (N1647, N1632, N1315);
nand NAND2 (N1648, N1647, N68);
nor NOR2 (N1649, N1640, N904);
xor XOR2 (N1650, N1648, N462);
and AND3 (N1651, N1619, N1218, N54);
and AND2 (N1652, N1644, N623);
not NOT1 (N1653, N1642);
not NOT1 (N1654, N1636);
nand NAND4 (N1655, N1651, N1048, N1190, N955);
nor NOR4 (N1656, N1643, N699, N1267, N891);
and AND3 (N1657, N1645, N1014, N614);
or OR3 (N1658, N1641, N22, N1068);
and AND4 (N1659, N1656, N1020, N1477, N95);
and AND2 (N1660, N1649, N596);
xor XOR2 (N1661, N1646, N281);
nor NOR3 (N1662, N1652, N1263, N52);
nand NAND4 (N1663, N1662, N1616, N121, N1412);
not NOT1 (N1664, N1660);
nor NOR3 (N1665, N1663, N1521, N1346);
buf BUF1 (N1666, N1665);
and AND4 (N1667, N1659, N317, N165, N1061);
nor NOR2 (N1668, N1666, N771);
not NOT1 (N1669, N1661);
or OR4 (N1670, N1667, N1123, N506, N328);
buf BUF1 (N1671, N1654);
or OR4 (N1672, N1657, N266, N317, N843);
buf BUF1 (N1673, N1671);
nor NOR4 (N1674, N1670, N892, N1112, N14);
xor XOR2 (N1675, N1672, N1260);
nor NOR3 (N1676, N1650, N377, N1015);
xor XOR2 (N1677, N1664, N461);
and AND3 (N1678, N1676, N292, N1151);
buf BUF1 (N1679, N1674);
nand NAND2 (N1680, N1673, N615);
or OR3 (N1681, N1653, N117, N756);
not NOT1 (N1682, N1655);
nand NAND2 (N1683, N1669, N1172);
xor XOR2 (N1684, N1680, N1446);
nand NAND4 (N1685, N1677, N195, N584, N639);
buf BUF1 (N1686, N1678);
buf BUF1 (N1687, N1685);
nor NOR2 (N1688, N1684, N501);
xor XOR2 (N1689, N1668, N1286);
buf BUF1 (N1690, N1675);
nand NAND3 (N1691, N1682, N517, N1352);
or OR4 (N1692, N1691, N1403, N1035, N814);
not NOT1 (N1693, N1681);
nand NAND3 (N1694, N1687, N1160, N756);
nand NAND2 (N1695, N1658, N815);
nand NAND3 (N1696, N1688, N364, N400);
and AND3 (N1697, N1695, N971, N1529);
nor NOR3 (N1698, N1694, N303, N373);
or OR2 (N1699, N1690, N779);
and AND2 (N1700, N1686, N825);
not NOT1 (N1701, N1700);
and AND4 (N1702, N1701, N374, N1516, N979);
and AND2 (N1703, N1693, N723);
nand NAND4 (N1704, N1689, N1296, N1000, N56);
nor NOR3 (N1705, N1698, N766, N348);
xor XOR2 (N1706, N1683, N1158);
and AND2 (N1707, N1703, N967);
buf BUF1 (N1708, N1679);
xor XOR2 (N1709, N1696, N1362);
buf BUF1 (N1710, N1706);
nor NOR3 (N1711, N1702, N1445, N1049);
xor XOR2 (N1712, N1692, N469);
buf BUF1 (N1713, N1707);
or OR4 (N1714, N1697, N1324, N1267, N841);
xor XOR2 (N1715, N1714, N458);
not NOT1 (N1716, N1711);
and AND2 (N1717, N1699, N390);
nor NOR4 (N1718, N1709, N111, N872, N48);
nor NOR3 (N1719, N1717, N191, N1072);
or OR2 (N1720, N1704, N1155);
buf BUF1 (N1721, N1710);
and AND2 (N1722, N1715, N1090);
buf BUF1 (N1723, N1712);
not NOT1 (N1724, N1718);
nand NAND3 (N1725, N1716, N1033, N271);
not NOT1 (N1726, N1720);
buf BUF1 (N1727, N1705);
nor NOR2 (N1728, N1723, N75);
nor NOR3 (N1729, N1724, N632, N1115);
nand NAND3 (N1730, N1727, N1559, N1054);
nor NOR4 (N1731, N1730, N1443, N523, N23);
buf BUF1 (N1732, N1726);
and AND2 (N1733, N1721, N357);
not NOT1 (N1734, N1725);
xor XOR2 (N1735, N1732, N1618);
xor XOR2 (N1736, N1729, N791);
xor XOR2 (N1737, N1731, N625);
not NOT1 (N1738, N1734);
or OR4 (N1739, N1733, N1348, N379, N148);
or OR2 (N1740, N1708, N1270);
not NOT1 (N1741, N1728);
nor NOR4 (N1742, N1740, N65, N187, N679);
or OR3 (N1743, N1739, N473, N506);
buf BUF1 (N1744, N1719);
nand NAND2 (N1745, N1744, N247);
or OR2 (N1746, N1738, N919);
xor XOR2 (N1747, N1741, N1702);
xor XOR2 (N1748, N1735, N315);
not NOT1 (N1749, N1713);
buf BUF1 (N1750, N1722);
nor NOR2 (N1751, N1737, N612);
not NOT1 (N1752, N1748);
nand NAND3 (N1753, N1745, N355, N243);
xor XOR2 (N1754, N1751, N1493);
buf BUF1 (N1755, N1746);
and AND2 (N1756, N1742, N350);
xor XOR2 (N1757, N1750, N773);
xor XOR2 (N1758, N1749, N70);
xor XOR2 (N1759, N1736, N1708);
xor XOR2 (N1760, N1759, N531);
nor NOR3 (N1761, N1743, N782, N792);
nor NOR4 (N1762, N1755, N1632, N138, N945);
xor XOR2 (N1763, N1753, N1579);
xor XOR2 (N1764, N1762, N1655);
and AND4 (N1765, N1764, N855, N205, N1309);
not NOT1 (N1766, N1754);
xor XOR2 (N1767, N1752, N1282);
not NOT1 (N1768, N1767);
xor XOR2 (N1769, N1763, N923);
or OR3 (N1770, N1756, N877, N804);
nor NOR4 (N1771, N1765, N1408, N824, N385);
nand NAND3 (N1772, N1768, N206, N1624);
nand NAND3 (N1773, N1761, N1016, N1270);
or OR2 (N1774, N1757, N1295);
and AND4 (N1775, N1760, N1627, N935, N817);
not NOT1 (N1776, N1766);
buf BUF1 (N1777, N1758);
and AND2 (N1778, N1775, N1355);
xor XOR2 (N1779, N1772, N940);
and AND3 (N1780, N1773, N1066, N1590);
not NOT1 (N1781, N1780);
nor NOR3 (N1782, N1747, N935, N518);
and AND3 (N1783, N1781, N630, N1041);
xor XOR2 (N1784, N1782, N1535);
not NOT1 (N1785, N1777);
buf BUF1 (N1786, N1774);
or OR3 (N1787, N1785, N287, N592);
nor NOR4 (N1788, N1776, N685, N1148, N471);
or OR2 (N1789, N1786, N858);
and AND3 (N1790, N1783, N1433, N1451);
nand NAND3 (N1791, N1787, N126, N1391);
nand NAND3 (N1792, N1769, N207, N1103);
buf BUF1 (N1793, N1779);
not NOT1 (N1794, N1788);
buf BUF1 (N1795, N1792);
xor XOR2 (N1796, N1794, N1519);
nor NOR3 (N1797, N1790, N1171, N808);
xor XOR2 (N1798, N1796, N514);
buf BUF1 (N1799, N1784);
xor XOR2 (N1800, N1797, N1488);
not NOT1 (N1801, N1778);
nand NAND4 (N1802, N1795, N294, N345, N754);
xor XOR2 (N1803, N1791, N1562);
and AND4 (N1804, N1799, N694, N1666, N182);
or OR2 (N1805, N1771, N1049);
nor NOR2 (N1806, N1802, N538);
nor NOR3 (N1807, N1803, N233, N511);
buf BUF1 (N1808, N1789);
not NOT1 (N1809, N1807);
xor XOR2 (N1810, N1806, N252);
nand NAND4 (N1811, N1793, N315, N1061, N112);
nor NOR3 (N1812, N1805, N1567, N403);
and AND4 (N1813, N1770, N332, N632, N296);
xor XOR2 (N1814, N1811, N1040);
and AND2 (N1815, N1814, N640);
or OR3 (N1816, N1808, N724, N1202);
nor NOR3 (N1817, N1810, N558, N664);
and AND2 (N1818, N1816, N1204);
or OR3 (N1819, N1813, N957, N89);
xor XOR2 (N1820, N1804, N168);
buf BUF1 (N1821, N1798);
or OR2 (N1822, N1815, N611);
xor XOR2 (N1823, N1821, N1117);
xor XOR2 (N1824, N1800, N1106);
nor NOR3 (N1825, N1818, N1089, N510);
buf BUF1 (N1826, N1825);
and AND2 (N1827, N1809, N916);
not NOT1 (N1828, N1823);
xor XOR2 (N1829, N1824, N819);
not NOT1 (N1830, N1820);
or OR2 (N1831, N1826, N861);
nor NOR4 (N1832, N1812, N1116, N1649, N46);
nand NAND4 (N1833, N1819, N1307, N667, N1146);
and AND3 (N1834, N1822, N1804, N744);
not NOT1 (N1835, N1827);
nand NAND3 (N1836, N1801, N1603, N1083);
xor XOR2 (N1837, N1835, N562);
nor NOR2 (N1838, N1828, N138);
nor NOR3 (N1839, N1838, N1157, N615);
not NOT1 (N1840, N1830);
xor XOR2 (N1841, N1832, N527);
not NOT1 (N1842, N1841);
not NOT1 (N1843, N1834);
and AND2 (N1844, N1840, N557);
xor XOR2 (N1845, N1843, N82);
nand NAND4 (N1846, N1839, N1647, N878, N1707);
and AND2 (N1847, N1831, N1768);
buf BUF1 (N1848, N1829);
buf BUF1 (N1849, N1845);
not NOT1 (N1850, N1842);
not NOT1 (N1851, N1844);
nor NOR2 (N1852, N1837, N556);
xor XOR2 (N1853, N1836, N1580);
not NOT1 (N1854, N1849);
nor NOR2 (N1855, N1850, N461);
buf BUF1 (N1856, N1855);
and AND2 (N1857, N1852, N603);
xor XOR2 (N1858, N1848, N623);
nand NAND2 (N1859, N1817, N309);
nand NAND2 (N1860, N1856, N126);
or OR2 (N1861, N1851, N600);
xor XOR2 (N1862, N1860, N377);
and AND3 (N1863, N1846, N956, N363);
nor NOR4 (N1864, N1861, N594, N688, N1672);
and AND3 (N1865, N1847, N302, N1321);
xor XOR2 (N1866, N1833, N1697);
or OR4 (N1867, N1857, N1274, N1686, N1356);
xor XOR2 (N1868, N1862, N672);
xor XOR2 (N1869, N1867, N1416);
buf BUF1 (N1870, N1859);
buf BUF1 (N1871, N1863);
nor NOR2 (N1872, N1865, N644);
not NOT1 (N1873, N1869);
nand NAND3 (N1874, N1873, N198, N491);
and AND2 (N1875, N1858, N1680);
nor NOR4 (N1876, N1864, N567, N880, N48);
xor XOR2 (N1877, N1872, N1057);
nand NAND2 (N1878, N1870, N1875);
buf BUF1 (N1879, N461);
buf BUF1 (N1880, N1878);
xor XOR2 (N1881, N1880, N1796);
nand NAND4 (N1882, N1879, N288, N1762, N373);
nor NOR4 (N1883, N1868, N571, N1766, N1305);
xor XOR2 (N1884, N1854, N563);
xor XOR2 (N1885, N1884, N1716);
buf BUF1 (N1886, N1874);
buf BUF1 (N1887, N1882);
and AND2 (N1888, N1866, N807);
buf BUF1 (N1889, N1887);
xor XOR2 (N1890, N1886, N1092);
buf BUF1 (N1891, N1890);
xor XOR2 (N1892, N1885, N1766);
buf BUF1 (N1893, N1892);
nor NOR2 (N1894, N1883, N674);
and AND4 (N1895, N1877, N1119, N852, N39);
nand NAND2 (N1896, N1888, N552);
not NOT1 (N1897, N1881);
not NOT1 (N1898, N1893);
xor XOR2 (N1899, N1853, N38);
not NOT1 (N1900, N1891);
and AND2 (N1901, N1889, N504);
buf BUF1 (N1902, N1901);
nand NAND2 (N1903, N1900, N1745);
nand NAND2 (N1904, N1903, N778);
and AND2 (N1905, N1897, N525);
or OR2 (N1906, N1898, N1303);
not NOT1 (N1907, N1871);
nor NOR3 (N1908, N1895, N816, N1876);
nand NAND4 (N1909, N1642, N1053, N1807, N1562);
or OR3 (N1910, N1894, N417, N47);
and AND4 (N1911, N1904, N511, N1584, N96);
nand NAND2 (N1912, N1902, N409);
and AND4 (N1913, N1899, N656, N525, N461);
xor XOR2 (N1914, N1912, N555);
nand NAND2 (N1915, N1914, N521);
not NOT1 (N1916, N1910);
and AND2 (N1917, N1906, N1398);
nand NAND3 (N1918, N1896, N1142, N734);
or OR3 (N1919, N1909, N1760, N1109);
and AND3 (N1920, N1919, N445, N147);
not NOT1 (N1921, N1917);
xor XOR2 (N1922, N1921, N366);
or OR3 (N1923, N1920, N1774, N923);
and AND3 (N1924, N1922, N833, N1278);
nor NOR3 (N1925, N1923, N1733, N98);
buf BUF1 (N1926, N1924);
or OR2 (N1927, N1925, N1568);
or OR4 (N1928, N1907, N1224, N662, N1447);
and AND2 (N1929, N1905, N1577);
not NOT1 (N1930, N1929);
not NOT1 (N1931, N1913);
or OR3 (N1932, N1927, N1343, N1731);
or OR4 (N1933, N1916, N23, N1853, N687);
buf BUF1 (N1934, N1918);
not NOT1 (N1935, N1908);
or OR2 (N1936, N1928, N1299);
nand NAND2 (N1937, N1926, N1373);
nor NOR2 (N1938, N1932, N1114);
buf BUF1 (N1939, N1931);
and AND3 (N1940, N1933, N396, N1046);
not NOT1 (N1941, N1934);
and AND4 (N1942, N1935, N1638, N1568, N350);
and AND2 (N1943, N1936, N514);
xor XOR2 (N1944, N1938, N1197);
nand NAND2 (N1945, N1943, N1339);
nand NAND2 (N1946, N1940, N1936);
and AND4 (N1947, N1944, N211, N603, N1311);
buf BUF1 (N1948, N1947);
not NOT1 (N1949, N1941);
not NOT1 (N1950, N1915);
nand NAND2 (N1951, N1911, N280);
xor XOR2 (N1952, N1949, N1332);
nand NAND4 (N1953, N1946, N1488, N1494, N1895);
buf BUF1 (N1954, N1951);
nand NAND4 (N1955, N1950, N1250, N829, N69);
and AND4 (N1956, N1942, N1885, N261, N140);
or OR3 (N1957, N1955, N1663, N532);
nand NAND4 (N1958, N1945, N786, N1844, N1639);
buf BUF1 (N1959, N1930);
buf BUF1 (N1960, N1959);
or OR3 (N1961, N1960, N660, N1404);
not NOT1 (N1962, N1948);
xor XOR2 (N1963, N1957, N1281);
nand NAND2 (N1964, N1954, N1645);
and AND3 (N1965, N1952, N867, N1535);
xor XOR2 (N1966, N1937, N805);
xor XOR2 (N1967, N1953, N1161);
buf BUF1 (N1968, N1965);
and AND4 (N1969, N1962, N301, N839, N1423);
nand NAND4 (N1970, N1963, N647, N356, N1780);
buf BUF1 (N1971, N1966);
not NOT1 (N1972, N1967);
not NOT1 (N1973, N1968);
nand NAND3 (N1974, N1971, N1355, N1639);
or OR4 (N1975, N1939, N1780, N299, N1972);
or OR4 (N1976, N957, N225, N1504, N1135);
not NOT1 (N1977, N1974);
nand NAND2 (N1978, N1969, N68);
not NOT1 (N1979, N1977);
nand NAND3 (N1980, N1956, N1772, N1246);
buf BUF1 (N1981, N1964);
not NOT1 (N1982, N1979);
or OR3 (N1983, N1973, N440, N1285);
buf BUF1 (N1984, N1982);
xor XOR2 (N1985, N1961, N412);
or OR2 (N1986, N1983, N1848);
and AND3 (N1987, N1986, N58, N1812);
nor NOR4 (N1988, N1978, N1529, N278, N1346);
xor XOR2 (N1989, N1981, N1044);
xor XOR2 (N1990, N1988, N927);
and AND4 (N1991, N1990, N1757, N742, N1569);
xor XOR2 (N1992, N1985, N1732);
and AND4 (N1993, N1984, N692, N1561, N1435);
or OR2 (N1994, N1958, N1682);
not NOT1 (N1995, N1994);
not NOT1 (N1996, N1975);
xor XOR2 (N1997, N1996, N795);
nand NAND3 (N1998, N1997, N888, N333);
nand NAND3 (N1999, N1995, N620, N1212);
nand NAND3 (N2000, N1976, N984, N1963);
xor XOR2 (N2001, N1989, N1440);
not NOT1 (N2002, N1970);
and AND3 (N2003, N1980, N1554, N104);
not NOT1 (N2004, N1999);
buf BUF1 (N2005, N2003);
or OR4 (N2006, N2000, N1981, N1930, N966);
nand NAND2 (N2007, N2005, N1951);
buf BUF1 (N2008, N2007);
buf BUF1 (N2009, N2004);
or OR3 (N2010, N1998, N394, N1545);
not NOT1 (N2011, N2008);
nand NAND4 (N2012, N2002, N432, N871, N906);
not NOT1 (N2013, N1992);
buf BUF1 (N2014, N1987);
or OR3 (N2015, N1993, N178, N1777);
and AND4 (N2016, N2013, N1635, N445, N888);
not NOT1 (N2017, N2014);
buf BUF1 (N2018, N2017);
buf BUF1 (N2019, N2010);
or OR4 (N2020, N2015, N51, N658, N333);
and AND2 (N2021, N2020, N1662);
buf BUF1 (N2022, N2019);
nand NAND3 (N2023, N2001, N395, N993);
nor NOR4 (N2024, N2006, N394, N1302, N366);
xor XOR2 (N2025, N1991, N1234);
nand NAND2 (N2026, N2022, N938);
xor XOR2 (N2027, N2023, N959);
buf BUF1 (N2028, N2012);
or OR2 (N2029, N2016, N1761);
nand NAND2 (N2030, N2028, N1614);
nor NOR4 (N2031, N2030, N952, N540, N1460);
not NOT1 (N2032, N2024);
and AND3 (N2033, N2029, N1142, N1395);
nor NOR3 (N2034, N2011, N1801, N1825);
nand NAND4 (N2035, N2026, N822, N1162, N1572);
nor NOR4 (N2036, N2018, N763, N1003, N1026);
xor XOR2 (N2037, N2032, N1898);
nor NOR3 (N2038, N2036, N1601, N51);
nand NAND3 (N2039, N2031, N181, N1380);
or OR4 (N2040, N2021, N1479, N7, N208);
and AND2 (N2041, N2037, N1394);
and AND2 (N2042, N2038, N458);
or OR3 (N2043, N2039, N140, N1287);
buf BUF1 (N2044, N2040);
nand NAND4 (N2045, N2044, N744, N528, N1405);
and AND2 (N2046, N2009, N1720);
or OR3 (N2047, N2042, N1112, N1422);
xor XOR2 (N2048, N2027, N1085);
not NOT1 (N2049, N2041);
not NOT1 (N2050, N2034);
and AND4 (N2051, N2025, N2015, N255, N2021);
nand NAND2 (N2052, N2049, N1105);
nand NAND3 (N2053, N2048, N537, N685);
nor NOR4 (N2054, N2043, N1448, N508, N1767);
nor NOR2 (N2055, N2035, N451);
not NOT1 (N2056, N2045);
not NOT1 (N2057, N2033);
buf BUF1 (N2058, N2047);
buf BUF1 (N2059, N2046);
and AND2 (N2060, N2057, N1439);
nand NAND4 (N2061, N2060, N1182, N886, N248);
not NOT1 (N2062, N2054);
and AND4 (N2063, N2053, N1645, N432, N1941);
nor NOR4 (N2064, N2059, N18, N722, N714);
xor XOR2 (N2065, N2051, N1657);
not NOT1 (N2066, N2058);
buf BUF1 (N2067, N2062);
buf BUF1 (N2068, N2055);
and AND3 (N2069, N2066, N919, N404);
nand NAND3 (N2070, N2068, N1966, N1344);
xor XOR2 (N2071, N2063, N334);
nor NOR4 (N2072, N2065, N127, N1347, N931);
nand NAND3 (N2073, N2052, N870, N721);
not NOT1 (N2074, N2073);
or OR3 (N2075, N2069, N1340, N1742);
not NOT1 (N2076, N2056);
xor XOR2 (N2077, N2072, N500);
and AND2 (N2078, N2067, N263);
not NOT1 (N2079, N2074);
nand NAND2 (N2080, N2079, N474);
and AND3 (N2081, N2080, N1987, N1182);
and AND2 (N2082, N2064, N795);
and AND3 (N2083, N2071, N1799, N982);
nand NAND4 (N2084, N2082, N2026, N467, N1977);
xor XOR2 (N2085, N2084, N160);
nor NOR3 (N2086, N2078, N2040, N2017);
or OR4 (N2087, N2081, N1011, N343, N482);
xor XOR2 (N2088, N2086, N1233);
nand NAND4 (N2089, N2087, N730, N1058, N1897);
not NOT1 (N2090, N2050);
buf BUF1 (N2091, N2085);
xor XOR2 (N2092, N2076, N1312);
nand NAND2 (N2093, N2070, N1128);
not NOT1 (N2094, N2093);
nand NAND4 (N2095, N2091, N1740, N1410, N1258);
xor XOR2 (N2096, N2095, N1988);
buf BUF1 (N2097, N2061);
and AND2 (N2098, N2088, N694);
nor NOR4 (N2099, N2097, N2039, N563, N1817);
nand NAND3 (N2100, N2089, N1898, N910);
buf BUF1 (N2101, N2075);
xor XOR2 (N2102, N2092, N1675);
or OR4 (N2103, N2094, N1634, N658, N221);
and AND4 (N2104, N2100, N1494, N696, N2087);
nor NOR2 (N2105, N2098, N1580);
or OR4 (N2106, N2077, N1002, N373, N1941);
or OR4 (N2107, N2099, N1211, N1746, N696);
nor NOR2 (N2108, N2090, N1239);
nor NOR3 (N2109, N2096, N632, N1656);
xor XOR2 (N2110, N2105, N1036);
and AND3 (N2111, N2106, N1437, N1821);
nand NAND4 (N2112, N2083, N41, N1491, N128);
buf BUF1 (N2113, N2110);
and AND3 (N2114, N2109, N279, N1512);
nor NOR2 (N2115, N2113, N226);
or OR4 (N2116, N2111, N538, N1788, N1063);
buf BUF1 (N2117, N2116);
not NOT1 (N2118, N2112);
buf BUF1 (N2119, N2102);
nor NOR3 (N2120, N2115, N2098, N1772);
and AND4 (N2121, N2119, N1316, N1323, N208);
or OR2 (N2122, N2101, N1601);
not NOT1 (N2123, N2103);
or OR4 (N2124, N2120, N1917, N180, N1238);
nand NAND3 (N2125, N2114, N905, N1013);
xor XOR2 (N2126, N2125, N748);
not NOT1 (N2127, N2122);
nor NOR2 (N2128, N2127, N174);
xor XOR2 (N2129, N2118, N1537);
or OR3 (N2130, N2108, N707, N1676);
not NOT1 (N2131, N2128);
buf BUF1 (N2132, N2129);
nand NAND3 (N2133, N2131, N1611, N764);
xor XOR2 (N2134, N2117, N1888);
and AND3 (N2135, N2126, N239, N1145);
not NOT1 (N2136, N2135);
and AND2 (N2137, N2121, N706);
xor XOR2 (N2138, N2132, N1152);
buf BUF1 (N2139, N2136);
not NOT1 (N2140, N2104);
nand NAND3 (N2141, N2134, N1577, N1830);
nor NOR4 (N2142, N2123, N525, N1601, N361);
or OR4 (N2143, N2141, N1411, N617, N1552);
and AND2 (N2144, N2124, N2045);
and AND2 (N2145, N2130, N943);
buf BUF1 (N2146, N2143);
buf BUF1 (N2147, N2146);
xor XOR2 (N2148, N2139, N1058);
xor XOR2 (N2149, N2107, N20);
and AND4 (N2150, N2140, N352, N67, N1019);
not NOT1 (N2151, N2150);
xor XOR2 (N2152, N2149, N29);
or OR4 (N2153, N2148, N1209, N669, N147);
nand NAND4 (N2154, N2152, N346, N1634, N122);
or OR2 (N2155, N2144, N626);
or OR2 (N2156, N2147, N820);
nor NOR4 (N2157, N2145, N914, N576, N50);
nand NAND2 (N2158, N2151, N772);
buf BUF1 (N2159, N2157);
buf BUF1 (N2160, N2156);
nor NOR4 (N2161, N2138, N1038, N26, N468);
or OR2 (N2162, N2158, N1050);
nor NOR2 (N2163, N2160, N875);
or OR4 (N2164, N2133, N1881, N880, N1574);
not NOT1 (N2165, N2153);
and AND4 (N2166, N2155, N1955, N209, N1811);
or OR2 (N2167, N2163, N1267);
not NOT1 (N2168, N2154);
nand NAND4 (N2169, N2166, N471, N895, N1324);
and AND4 (N2170, N2167, N1873, N1942, N356);
and AND3 (N2171, N2168, N326, N934);
or OR4 (N2172, N2137, N1858, N1907, N795);
nor NOR2 (N2173, N2159, N2116);
nor NOR4 (N2174, N2171, N603, N1194, N555);
and AND3 (N2175, N2161, N25, N2068);
nor NOR3 (N2176, N2142, N2117, N1460);
nor NOR3 (N2177, N2162, N178, N619);
xor XOR2 (N2178, N2164, N1969);
or OR4 (N2179, N2174, N321, N1007, N882);
not NOT1 (N2180, N2173);
and AND3 (N2181, N2175, N1378, N328);
and AND3 (N2182, N2165, N1864, N1718);
and AND3 (N2183, N2176, N1251, N2130);
and AND2 (N2184, N2179, N1132);
or OR2 (N2185, N2182, N989);
buf BUF1 (N2186, N2177);
nor NOR3 (N2187, N2170, N646, N407);
nand NAND3 (N2188, N2181, N1271, N1981);
nor NOR3 (N2189, N2187, N35, N721);
nor NOR3 (N2190, N2189, N2152, N182);
buf BUF1 (N2191, N2184);
nor NOR2 (N2192, N2186, N1678);
nand NAND3 (N2193, N2183, N284, N2097);
nor NOR4 (N2194, N2185, N1035, N417, N1616);
or OR2 (N2195, N2191, N414);
nand NAND2 (N2196, N2190, N2072);
xor XOR2 (N2197, N2192, N734);
not NOT1 (N2198, N2172);
and AND3 (N2199, N2197, N804, N1936);
nand NAND2 (N2200, N2198, N532);
buf BUF1 (N2201, N2188);
nor NOR4 (N2202, N2194, N311, N898, N488);
nor NOR3 (N2203, N2180, N115, N1797);
and AND2 (N2204, N2199, N1139);
and AND3 (N2205, N2196, N691, N1909);
not NOT1 (N2206, N2169);
nand NAND3 (N2207, N2202, N2060, N1272);
buf BUF1 (N2208, N2201);
and AND4 (N2209, N2203, N2161, N526, N956);
and AND2 (N2210, N2206, N654);
nand NAND3 (N2211, N2208, N147, N527);
not NOT1 (N2212, N2210);
and AND2 (N2213, N2211, N1577);
nor NOR3 (N2214, N2209, N2167, N1212);
nor NOR3 (N2215, N2195, N886, N1502);
and AND2 (N2216, N2213, N1322);
xor XOR2 (N2217, N2200, N371);
not NOT1 (N2218, N2212);
nor NOR4 (N2219, N2215, N1514, N1686, N1762);
or OR2 (N2220, N2218, N1202);
or OR2 (N2221, N2204, N1852);
xor XOR2 (N2222, N2217, N966);
not NOT1 (N2223, N2216);
nand NAND4 (N2224, N2205, N1499, N474, N1898);
buf BUF1 (N2225, N2223);
or OR3 (N2226, N2214, N1882, N1854);
or OR4 (N2227, N2222, N1211, N1063, N466);
not NOT1 (N2228, N2220);
xor XOR2 (N2229, N2226, N1384);
buf BUF1 (N2230, N2227);
or OR4 (N2231, N2193, N1075, N2128, N149);
xor XOR2 (N2232, N2178, N394);
not NOT1 (N2233, N2228);
nand NAND3 (N2234, N2231, N156, N993);
buf BUF1 (N2235, N2234);
or OR2 (N2236, N2230, N2010);
not NOT1 (N2237, N2207);
or OR4 (N2238, N2232, N1131, N1560, N1051);
nand NAND2 (N2239, N2238, N1879);
and AND4 (N2240, N2229, N565, N2164, N73);
not NOT1 (N2241, N2224);
or OR2 (N2242, N2235, N1068);
or OR3 (N2243, N2237, N508, N1721);
nor NOR2 (N2244, N2240, N1082);
nand NAND2 (N2245, N2233, N1459);
nand NAND3 (N2246, N2241, N210, N2217);
not NOT1 (N2247, N2236);
or OR3 (N2248, N2242, N1003, N229);
nand NAND3 (N2249, N2248, N194, N606);
not NOT1 (N2250, N2247);
and AND3 (N2251, N2246, N2058, N1475);
and AND4 (N2252, N2245, N86, N1823, N796);
nor NOR3 (N2253, N2243, N1371, N926);
and AND2 (N2254, N2239, N247);
xor XOR2 (N2255, N2221, N499);
and AND3 (N2256, N2253, N687, N2190);
and AND3 (N2257, N2254, N1614, N2229);
nand NAND2 (N2258, N2255, N1550);
not NOT1 (N2259, N2219);
nor NOR2 (N2260, N2251, N2150);
xor XOR2 (N2261, N2256, N1293);
xor XOR2 (N2262, N2244, N538);
xor XOR2 (N2263, N2225, N17);
buf BUF1 (N2264, N2262);
nand NAND4 (N2265, N2263, N1113, N449, N1518);
xor XOR2 (N2266, N2257, N2201);
nor NOR4 (N2267, N2266, N439, N1483, N1057);
and AND4 (N2268, N2250, N2250, N2001, N1288);
and AND2 (N2269, N2249, N1822);
xor XOR2 (N2270, N2268, N274);
nor NOR4 (N2271, N2265, N1450, N1174, N1527);
xor XOR2 (N2272, N2271, N810);
not NOT1 (N2273, N2252);
and AND3 (N2274, N2267, N994, N235);
and AND2 (N2275, N2272, N765);
and AND2 (N2276, N2259, N567);
xor XOR2 (N2277, N2274, N635);
not NOT1 (N2278, N2277);
or OR2 (N2279, N2273, N811);
not NOT1 (N2280, N2278);
or OR4 (N2281, N2276, N1058, N883, N2067);
not NOT1 (N2282, N2258);
nand NAND4 (N2283, N2275, N1056, N1388, N2279);
not NOT1 (N2284, N1396);
nand NAND4 (N2285, N2269, N605, N1385, N2069);
nor NOR4 (N2286, N2281, N674, N1582, N939);
buf BUF1 (N2287, N2261);
buf BUF1 (N2288, N2284);
nor NOR2 (N2289, N2260, N1608);
or OR2 (N2290, N2285, N1072);
nand NAND4 (N2291, N2270, N1147, N26, N1908);
or OR2 (N2292, N2283, N20);
or OR2 (N2293, N2288, N135);
and AND2 (N2294, N2282, N1475);
nor NOR4 (N2295, N2289, N2151, N421, N1692);
or OR2 (N2296, N2292, N439);
and AND4 (N2297, N2295, N529, N1681, N1099);
buf BUF1 (N2298, N2290);
and AND2 (N2299, N2296, N764);
and AND4 (N2300, N2264, N1781, N1039, N1274);
and AND4 (N2301, N2287, N1467, N1840, N270);
nand NAND3 (N2302, N2294, N1709, N1664);
and AND4 (N2303, N2286, N1193, N648, N1788);
and AND2 (N2304, N2299, N626);
buf BUF1 (N2305, N2301);
not NOT1 (N2306, N2303);
nand NAND3 (N2307, N2298, N1886, N1777);
and AND4 (N2308, N2280, N1596, N224, N876);
nor NOR4 (N2309, N2306, N407, N1229, N185);
and AND2 (N2310, N2305, N1649);
not NOT1 (N2311, N2307);
nor NOR4 (N2312, N2291, N2049, N2286, N2056);
xor XOR2 (N2313, N2312, N304);
buf BUF1 (N2314, N2297);
or OR4 (N2315, N2310, N1561, N76, N855);
nor NOR2 (N2316, N2311, N87);
xor XOR2 (N2317, N2313, N1388);
buf BUF1 (N2318, N2304);
xor XOR2 (N2319, N2300, N440);
and AND3 (N2320, N2315, N664, N700);
xor XOR2 (N2321, N2319, N2277);
nor NOR3 (N2322, N2314, N1607, N337);
and AND3 (N2323, N2302, N2030, N960);
or OR3 (N2324, N2308, N390, N1315);
or OR3 (N2325, N2324, N1055, N2021);
and AND2 (N2326, N2325, N376);
nor NOR2 (N2327, N2318, N934);
xor XOR2 (N2328, N2323, N119);
or OR3 (N2329, N2328, N1790, N1474);
nand NAND3 (N2330, N2321, N1792, N1491);
not NOT1 (N2331, N2326);
nand NAND3 (N2332, N2327, N1363, N2147);
and AND4 (N2333, N2330, N840, N321, N477);
nand NAND3 (N2334, N2309, N457, N1435);
nor NOR3 (N2335, N2332, N1815, N1485);
xor XOR2 (N2336, N2334, N2003);
nor NOR4 (N2337, N2333, N1330, N1486, N1163);
not NOT1 (N2338, N2320);
nand NAND4 (N2339, N2322, N1172, N1112, N1941);
not NOT1 (N2340, N2316);
or OR3 (N2341, N2335, N1347, N405);
and AND3 (N2342, N2331, N745, N1595);
and AND2 (N2343, N2317, N1881);
nand NAND4 (N2344, N2336, N565, N1607, N738);
buf BUF1 (N2345, N2341);
and AND3 (N2346, N2340, N883, N1499);
and AND2 (N2347, N2329, N1071);
nor NOR4 (N2348, N2345, N1962, N375, N2106);
or OR3 (N2349, N2337, N1551, N2054);
buf BUF1 (N2350, N2344);
nand NAND2 (N2351, N2349, N2168);
and AND2 (N2352, N2346, N1458);
and AND3 (N2353, N2339, N156, N483);
nor NOR3 (N2354, N2350, N2079, N399);
buf BUF1 (N2355, N2338);
not NOT1 (N2356, N2343);
buf BUF1 (N2357, N2347);
nor NOR3 (N2358, N2356, N979, N2085);
not NOT1 (N2359, N2351);
nor NOR3 (N2360, N2352, N140, N2111);
not NOT1 (N2361, N2348);
buf BUF1 (N2362, N2360);
buf BUF1 (N2363, N2353);
xor XOR2 (N2364, N2361, N2158);
xor XOR2 (N2365, N2293, N1227);
nand NAND3 (N2366, N2355, N2176, N1001);
buf BUF1 (N2367, N2363);
buf BUF1 (N2368, N2342);
not NOT1 (N2369, N2354);
or OR4 (N2370, N2365, N1603, N914, N279);
nand NAND2 (N2371, N2367, N1698);
or OR2 (N2372, N2357, N540);
and AND2 (N2373, N2358, N2123);
xor XOR2 (N2374, N2359, N906);
not NOT1 (N2375, N2373);
nand NAND2 (N2376, N2372, N1544);
not NOT1 (N2377, N2369);
or OR3 (N2378, N2362, N2041, N482);
not NOT1 (N2379, N2366);
xor XOR2 (N2380, N2375, N1659);
and AND2 (N2381, N2378, N655);
or OR2 (N2382, N2377, N261);
xor XOR2 (N2383, N2370, N1671);
xor XOR2 (N2384, N2380, N1600);
nor NOR2 (N2385, N2368, N1883);
nand NAND4 (N2386, N2371, N135, N1067, N398);
and AND2 (N2387, N2383, N611);
buf BUF1 (N2388, N2386);
nor NOR4 (N2389, N2387, N1255, N222, N1785);
and AND3 (N2390, N2388, N1728, N1248);
buf BUF1 (N2391, N2389);
or OR4 (N2392, N2374, N2357, N145, N1397);
and AND3 (N2393, N2392, N1298, N1934);
or OR3 (N2394, N2390, N1335, N756);
or OR3 (N2395, N2393, N208, N1912);
buf BUF1 (N2396, N2394);
buf BUF1 (N2397, N2379);
not NOT1 (N2398, N2382);
or OR3 (N2399, N2376, N2086, N1998);
xor XOR2 (N2400, N2384, N657);
or OR4 (N2401, N2395, N2049, N2285, N2068);
and AND2 (N2402, N2396, N640);
buf BUF1 (N2403, N2401);
buf BUF1 (N2404, N2403);
and AND3 (N2405, N2399, N1201, N1506);
nand NAND2 (N2406, N2405, N1132);
or OR4 (N2407, N2402, N606, N839, N561);
or OR3 (N2408, N2381, N1131, N1934);
nand NAND4 (N2409, N2385, N1786, N1235, N257);
nor NOR2 (N2410, N2404, N951);
xor XOR2 (N2411, N2407, N602);
xor XOR2 (N2412, N2398, N1010);
nand NAND3 (N2413, N2364, N1953, N1202);
and AND2 (N2414, N2409, N1395);
nor NOR2 (N2415, N2406, N1536);
buf BUF1 (N2416, N2411);
or OR3 (N2417, N2410, N2240, N1136);
or OR4 (N2418, N2416, N130, N358, N345);
xor XOR2 (N2419, N2412, N2348);
xor XOR2 (N2420, N2408, N1825);
xor XOR2 (N2421, N2414, N2242);
not NOT1 (N2422, N2417);
nand NAND4 (N2423, N2421, N1053, N1738, N1276);
nand NAND4 (N2424, N2420, N2165, N654, N1964);
or OR3 (N2425, N2423, N2291, N1540);
and AND3 (N2426, N2400, N791, N1851);
not NOT1 (N2427, N2425);
and AND4 (N2428, N2419, N649, N1240, N2242);
nor NOR4 (N2429, N2397, N1696, N1302, N1749);
xor XOR2 (N2430, N2428, N229);
nand NAND3 (N2431, N2422, N2064, N1545);
not NOT1 (N2432, N2430);
and AND2 (N2433, N2432, N495);
buf BUF1 (N2434, N2418);
nor NOR2 (N2435, N2431, N938);
nor NOR3 (N2436, N2435, N2214, N1639);
nand NAND4 (N2437, N2434, N55, N1392, N2385);
nor NOR2 (N2438, N2413, N239);
nand NAND4 (N2439, N2391, N196, N1917, N105);
xor XOR2 (N2440, N2437, N2298);
or OR3 (N2441, N2440, N579, N1320);
nand NAND2 (N2442, N2439, N827);
nor NOR4 (N2443, N2436, N174, N73, N445);
and AND2 (N2444, N2429, N760);
not NOT1 (N2445, N2415);
buf BUF1 (N2446, N2442);
nor NOR4 (N2447, N2446, N2100, N323, N1934);
and AND4 (N2448, N2441, N14, N2379, N188);
nor NOR3 (N2449, N2445, N961, N2115);
xor XOR2 (N2450, N2447, N2129);
buf BUF1 (N2451, N2424);
not NOT1 (N2452, N2433);
or OR4 (N2453, N2450, N469, N998, N1071);
and AND3 (N2454, N2452, N1180, N1598);
xor XOR2 (N2455, N2449, N268);
buf BUF1 (N2456, N2444);
not NOT1 (N2457, N2454);
or OR3 (N2458, N2426, N2112, N1027);
not NOT1 (N2459, N2455);
and AND2 (N2460, N2443, N1589);
xor XOR2 (N2461, N2451, N173);
nor NOR3 (N2462, N2460, N323, N354);
xor XOR2 (N2463, N2453, N1027);
nor NOR4 (N2464, N2463, N2425, N117, N880);
and AND2 (N2465, N2461, N832);
or OR4 (N2466, N2456, N1718, N1725, N2266);
or OR3 (N2467, N2457, N1866, N1166);
not NOT1 (N2468, N2459);
and AND4 (N2469, N2448, N2245, N2426, N1019);
nor NOR4 (N2470, N2467, N1786, N2170, N428);
not NOT1 (N2471, N2470);
nor NOR3 (N2472, N2468, N2230, N1499);
xor XOR2 (N2473, N2427, N957);
xor XOR2 (N2474, N2464, N675);
and AND2 (N2475, N2458, N1887);
buf BUF1 (N2476, N2472);
nor NOR2 (N2477, N2465, N2402);
nand NAND2 (N2478, N2473, N1428);
not NOT1 (N2479, N2475);
xor XOR2 (N2480, N2478, N958);
nor NOR2 (N2481, N2471, N1698);
buf BUF1 (N2482, N2479);
xor XOR2 (N2483, N2469, N1575);
nor NOR3 (N2484, N2462, N194, N403);
nor NOR2 (N2485, N2482, N2180);
and AND3 (N2486, N2481, N2260, N1078);
and AND2 (N2487, N2477, N1185);
and AND4 (N2488, N2483, N2145, N1568, N2341);
or OR4 (N2489, N2476, N1835, N1726, N534);
nand NAND3 (N2490, N2466, N972, N1301);
or OR4 (N2491, N2438, N2075, N2482, N830);
buf BUF1 (N2492, N2491);
nor NOR3 (N2493, N2486, N2429, N430);
nand NAND2 (N2494, N2492, N1890);
and AND4 (N2495, N2494, N1685, N1190, N1784);
or OR2 (N2496, N2474, N1848);
nor NOR4 (N2497, N2484, N61, N12, N236);
or OR2 (N2498, N2497, N1357);
or OR2 (N2499, N2488, N741);
or OR2 (N2500, N2495, N1696);
xor XOR2 (N2501, N2480, N1838);
or OR4 (N2502, N2496, N1509, N1213, N305);
and AND3 (N2503, N2493, N5, N288);
nor NOR2 (N2504, N2490, N2495);
xor XOR2 (N2505, N2500, N1292);
nor NOR4 (N2506, N2487, N2289, N1338, N667);
nand NAND4 (N2507, N2489, N1009, N1216, N1669);
nand NAND2 (N2508, N2485, N406);
nor NOR2 (N2509, N2499, N1845);
xor XOR2 (N2510, N2503, N2147);
and AND2 (N2511, N2505, N2206);
xor XOR2 (N2512, N2504, N2505);
nor NOR3 (N2513, N2501, N1147, N918);
or OR4 (N2514, N2513, N1805, N755, N1715);
nand NAND3 (N2515, N2510, N817, N1977);
xor XOR2 (N2516, N2511, N1367);
xor XOR2 (N2517, N2508, N1905);
and AND3 (N2518, N2509, N1873, N2141);
xor XOR2 (N2519, N2512, N48);
not NOT1 (N2520, N2514);
buf BUF1 (N2521, N2506);
not NOT1 (N2522, N2521);
nor NOR4 (N2523, N2518, N2276, N41, N6);
or OR2 (N2524, N2502, N1486);
or OR3 (N2525, N2515, N1060, N380);
xor XOR2 (N2526, N2523, N1289);
buf BUF1 (N2527, N2517);
and AND4 (N2528, N2519, N709, N438, N1966);
nor NOR3 (N2529, N2527, N1545, N1750);
or OR3 (N2530, N2522, N2021, N1239);
not NOT1 (N2531, N2525);
nand NAND3 (N2532, N2498, N2193, N1528);
or OR4 (N2533, N2524, N592, N715, N315);
xor XOR2 (N2534, N2526, N146);
xor XOR2 (N2535, N2520, N1718);
and AND4 (N2536, N2530, N2020, N1717, N971);
or OR3 (N2537, N2535, N33, N1451);
xor XOR2 (N2538, N2516, N2015);
xor XOR2 (N2539, N2532, N309);
and AND2 (N2540, N2533, N1153);
xor XOR2 (N2541, N2537, N2167);
nand NAND4 (N2542, N2534, N829, N1590, N422);
and AND3 (N2543, N2531, N2525, N813);
and AND4 (N2544, N2540, N478, N1586, N1966);
nand NAND3 (N2545, N2528, N251, N1297);
nand NAND3 (N2546, N2539, N59, N424);
buf BUF1 (N2547, N2543);
nor NOR2 (N2548, N2546, N164);
buf BUF1 (N2549, N2547);
xor XOR2 (N2550, N2541, N134);
or OR4 (N2551, N2538, N2369, N2374, N519);
not NOT1 (N2552, N2544);
nor NOR2 (N2553, N2545, N654);
or OR3 (N2554, N2549, N1318, N56);
nor NOR3 (N2555, N2548, N2474, N759);
nor NOR4 (N2556, N2554, N1012, N1966, N733);
xor XOR2 (N2557, N2529, N1935);
nor NOR4 (N2558, N2555, N1177, N2344, N1238);
or OR4 (N2559, N2556, N1713, N524, N1582);
or OR4 (N2560, N2552, N2219, N1701, N667);
or OR2 (N2561, N2536, N1059);
and AND3 (N2562, N2558, N1396, N1505);
or OR4 (N2563, N2507, N1860, N1783, N2548);
nand NAND2 (N2564, N2563, N2092);
not NOT1 (N2565, N2550);
not NOT1 (N2566, N2559);
nor NOR3 (N2567, N2562, N214, N2431);
nor NOR3 (N2568, N2567, N1052, N1015);
nand NAND3 (N2569, N2557, N551, N198);
nor NOR4 (N2570, N2569, N388, N2017, N2527);
nand NAND3 (N2571, N2561, N2118, N1241);
nor NOR3 (N2572, N2568, N1891, N37);
and AND2 (N2573, N2570, N1611);
or OR3 (N2574, N2551, N965, N1903);
nand NAND3 (N2575, N2560, N462, N2017);
xor XOR2 (N2576, N2564, N768);
and AND4 (N2577, N2542, N13, N339, N1131);
nand NAND3 (N2578, N2575, N1636, N1934);
nor NOR4 (N2579, N2576, N226, N2272, N1541);
and AND3 (N2580, N2572, N271, N2077);
xor XOR2 (N2581, N2579, N170);
nand NAND4 (N2582, N2565, N1171, N1881, N941);
or OR3 (N2583, N2553, N1585, N841);
or OR2 (N2584, N2574, N1707);
nand NAND3 (N2585, N2581, N804, N558);
or OR3 (N2586, N2582, N1524, N2366);
xor XOR2 (N2587, N2580, N2468);
nand NAND3 (N2588, N2577, N940, N2518);
xor XOR2 (N2589, N2586, N1864);
nand NAND4 (N2590, N2583, N974, N684, N397);
xor XOR2 (N2591, N2571, N1366);
xor XOR2 (N2592, N2591, N635);
buf BUF1 (N2593, N2573);
nand NAND4 (N2594, N2593, N1808, N1983, N477);
buf BUF1 (N2595, N2587);
buf BUF1 (N2596, N2590);
or OR4 (N2597, N2589, N2452, N297, N411);
xor XOR2 (N2598, N2592, N148);
not NOT1 (N2599, N2595);
or OR2 (N2600, N2584, N2000);
not NOT1 (N2601, N2566);
nor NOR2 (N2602, N2594, N137);
not NOT1 (N2603, N2588);
xor XOR2 (N2604, N2585, N411);
not NOT1 (N2605, N2604);
buf BUF1 (N2606, N2603);
nand NAND2 (N2607, N2596, N377);
nand NAND3 (N2608, N2607, N237, N2123);
buf BUF1 (N2609, N2597);
not NOT1 (N2610, N2606);
or OR3 (N2611, N2609, N541, N6);
and AND4 (N2612, N2611, N2002, N2369, N1929);
not NOT1 (N2613, N2578);
or OR2 (N2614, N2602, N1275);
or OR3 (N2615, N2599, N246, N293);
buf BUF1 (N2616, N2605);
nor NOR2 (N2617, N2601, N1357);
xor XOR2 (N2618, N2613, N2366);
buf BUF1 (N2619, N2616);
and AND3 (N2620, N2617, N2156, N2083);
or OR3 (N2621, N2608, N137, N1554);
buf BUF1 (N2622, N2619);
xor XOR2 (N2623, N2615, N601);
and AND2 (N2624, N2622, N2201);
not NOT1 (N2625, N2623);
or OR3 (N2626, N2598, N16, N243);
not NOT1 (N2627, N2618);
buf BUF1 (N2628, N2624);
nand NAND2 (N2629, N2628, N1043);
and AND2 (N2630, N2600, N1847);
xor XOR2 (N2631, N2625, N1661);
nand NAND4 (N2632, N2630, N2167, N1303, N2095);
and AND4 (N2633, N2621, N2148, N509, N90);
or OR4 (N2634, N2612, N975, N2251, N430);
not NOT1 (N2635, N2614);
nand NAND4 (N2636, N2632, N18, N1034, N2326);
and AND4 (N2637, N2636, N71, N2379, N934);
buf BUF1 (N2638, N2634);
nand NAND2 (N2639, N2635, N2269);
nand NAND3 (N2640, N2639, N164, N1027);
buf BUF1 (N2641, N2627);
not NOT1 (N2642, N2640);
buf BUF1 (N2643, N2633);
and AND2 (N2644, N2610, N2539);
xor XOR2 (N2645, N2641, N747);
xor XOR2 (N2646, N2642, N2452);
nor NOR2 (N2647, N2626, N2251);
xor XOR2 (N2648, N2643, N2153);
xor XOR2 (N2649, N2631, N1464);
or OR4 (N2650, N2646, N438, N1569, N621);
nor NOR4 (N2651, N2638, N267, N1142, N1312);
or OR2 (N2652, N2645, N2507);
xor XOR2 (N2653, N2652, N502);
xor XOR2 (N2654, N2620, N1021);
buf BUF1 (N2655, N2644);
buf BUF1 (N2656, N2649);
or OR2 (N2657, N2656, N2583);
nand NAND3 (N2658, N2653, N2488, N213);
nor NOR3 (N2659, N2647, N68, N773);
nand NAND3 (N2660, N2650, N2131, N744);
buf BUF1 (N2661, N2657);
xor XOR2 (N2662, N2629, N637);
and AND3 (N2663, N2655, N1258, N160);
not NOT1 (N2664, N2660);
nor NOR2 (N2665, N2654, N2057);
xor XOR2 (N2666, N2651, N1428);
not NOT1 (N2667, N2659);
not NOT1 (N2668, N2667);
buf BUF1 (N2669, N2664);
buf BUF1 (N2670, N2669);
or OR2 (N2671, N2666, N1617);
nand NAND3 (N2672, N2648, N1417, N2248);
nand NAND4 (N2673, N2670, N2361, N125, N646);
nand NAND4 (N2674, N2662, N1323, N1472, N692);
or OR2 (N2675, N2658, N35);
and AND4 (N2676, N2672, N36, N1211, N856);
or OR2 (N2677, N2665, N547);
buf BUF1 (N2678, N2637);
buf BUF1 (N2679, N2674);
nor NOR3 (N2680, N2675, N747, N2405);
nand NAND4 (N2681, N2680, N1333, N1807, N1866);
and AND2 (N2682, N2668, N1409);
buf BUF1 (N2683, N2681);
not NOT1 (N2684, N2683);
buf BUF1 (N2685, N2684);
or OR4 (N2686, N2671, N91, N420, N2510);
nand NAND4 (N2687, N2661, N2500, N2211, N2514);
nand NAND3 (N2688, N2682, N1114, N1586);
and AND2 (N2689, N2686, N1449);
nand NAND3 (N2690, N2679, N1977, N2632);
nor NOR4 (N2691, N2678, N1194, N966, N1456);
buf BUF1 (N2692, N2673);
nor NOR3 (N2693, N2690, N1341, N1269);
and AND4 (N2694, N2676, N798, N1037, N635);
nor NOR3 (N2695, N2677, N1981, N1745);
buf BUF1 (N2696, N2687);
buf BUF1 (N2697, N2692);
nor NOR2 (N2698, N2689, N859);
buf BUF1 (N2699, N2688);
not NOT1 (N2700, N2685);
not NOT1 (N2701, N2699);
buf BUF1 (N2702, N2663);
not NOT1 (N2703, N2700);
buf BUF1 (N2704, N2696);
and AND4 (N2705, N2704, N1722, N1295, N1287);
nor NOR2 (N2706, N2705, N1761);
and AND3 (N2707, N2706, N562, N2223);
buf BUF1 (N2708, N2698);
nor NOR3 (N2709, N2695, N353, N887);
nand NAND3 (N2710, N2694, N2079, N1339);
buf BUF1 (N2711, N2703);
not NOT1 (N2712, N2701);
nand NAND2 (N2713, N2702, N1283);
nor NOR3 (N2714, N2711, N953, N1521);
not NOT1 (N2715, N2707);
xor XOR2 (N2716, N2708, N20);
or OR2 (N2717, N2716, N851);
or OR2 (N2718, N2697, N138);
not NOT1 (N2719, N2709);
nor NOR2 (N2720, N2714, N1712);
nor NOR3 (N2721, N2710, N2203, N445);
xor XOR2 (N2722, N2715, N1093);
not NOT1 (N2723, N2691);
not NOT1 (N2724, N2721);
or OR2 (N2725, N2724, N2173);
not NOT1 (N2726, N2713);
not NOT1 (N2727, N2719);
not NOT1 (N2728, N2725);
buf BUF1 (N2729, N2722);
xor XOR2 (N2730, N2729, N1064);
nand NAND2 (N2731, N2718, N2196);
or OR4 (N2732, N2723, N766, N886, N220);
or OR4 (N2733, N2728, N14, N1526, N2136);
buf BUF1 (N2734, N2730);
and AND4 (N2735, N2693, N111, N742, N1303);
and AND3 (N2736, N2731, N112, N797);
nor NOR3 (N2737, N2717, N880, N1130);
and AND4 (N2738, N2712, N753, N2614, N122);
and AND2 (N2739, N2726, N1399);
xor XOR2 (N2740, N2739, N2462);
or OR4 (N2741, N2737, N1732, N2707, N2241);
or OR3 (N2742, N2738, N1327, N844);
and AND4 (N2743, N2736, N2679, N260, N2271);
xor XOR2 (N2744, N2740, N2686);
and AND3 (N2745, N2744, N142, N1379);
not NOT1 (N2746, N2735);
xor XOR2 (N2747, N2743, N1853);
and AND4 (N2748, N2720, N2744, N1646, N761);
not NOT1 (N2749, N2746);
buf BUF1 (N2750, N2747);
nor NOR4 (N2751, N2734, N1090, N1496, N346);
or OR4 (N2752, N2727, N2452, N1771, N2256);
not NOT1 (N2753, N2745);
not NOT1 (N2754, N2748);
xor XOR2 (N2755, N2733, N2633);
xor XOR2 (N2756, N2755, N2050);
nor NOR3 (N2757, N2749, N1736, N316);
buf BUF1 (N2758, N2741);
not NOT1 (N2759, N2732);
not NOT1 (N2760, N2754);
nor NOR4 (N2761, N2752, N369, N1015, N2562);
nand NAND2 (N2762, N2750, N888);
xor XOR2 (N2763, N2742, N153);
or OR4 (N2764, N2762, N630, N294, N248);
nor NOR2 (N2765, N2753, N229);
and AND3 (N2766, N2756, N279, N1889);
xor XOR2 (N2767, N2766, N1121);
nand NAND2 (N2768, N2760, N1466);
buf BUF1 (N2769, N2759);
and AND4 (N2770, N2768, N1274, N2578, N146);
or OR3 (N2771, N2761, N1232, N994);
or OR3 (N2772, N2769, N1015, N1370);
nand NAND3 (N2773, N2765, N184, N1257);
or OR2 (N2774, N2758, N2640);
or OR3 (N2775, N2763, N1007, N2087);
not NOT1 (N2776, N2774);
or OR4 (N2777, N2773, N2272, N1097, N1875);
nand NAND4 (N2778, N2757, N50, N771, N1449);
not NOT1 (N2779, N2751);
xor XOR2 (N2780, N2779, N135);
or OR3 (N2781, N2770, N2777, N255);
not NOT1 (N2782, N1152);
not NOT1 (N2783, N2782);
nand NAND3 (N2784, N2767, N130, N1468);
buf BUF1 (N2785, N2776);
or OR2 (N2786, N2775, N2556);
nand NAND2 (N2787, N2781, N2544);
xor XOR2 (N2788, N2785, N1785);
buf BUF1 (N2789, N2772);
or OR2 (N2790, N2780, N1785);
nor NOR4 (N2791, N2786, N1329, N2523, N63);
xor XOR2 (N2792, N2784, N88);
nand NAND4 (N2793, N2789, N1607, N1108, N1661);
xor XOR2 (N2794, N2792, N196);
or OR3 (N2795, N2790, N272, N458);
not NOT1 (N2796, N2764);
xor XOR2 (N2797, N2791, N1279);
nand NAND3 (N2798, N2771, N1391, N348);
buf BUF1 (N2799, N2788);
not NOT1 (N2800, N2795);
buf BUF1 (N2801, N2797);
not NOT1 (N2802, N2793);
not NOT1 (N2803, N2800);
buf BUF1 (N2804, N2787);
nor NOR2 (N2805, N2778, N2145);
or OR3 (N2806, N2783, N279, N777);
buf BUF1 (N2807, N2802);
not NOT1 (N2808, N2798);
not NOT1 (N2809, N2806);
not NOT1 (N2810, N2799);
xor XOR2 (N2811, N2805, N1988);
xor XOR2 (N2812, N2801, N613);
not NOT1 (N2813, N2810);
or OR3 (N2814, N2809, N1362, N2099);
buf BUF1 (N2815, N2808);
buf BUF1 (N2816, N2813);
or OR3 (N2817, N2814, N824, N1598);
xor XOR2 (N2818, N2816, N2610);
or OR4 (N2819, N2812, N2312, N2414, N396);
nor NOR3 (N2820, N2796, N224, N219);
or OR3 (N2821, N2818, N2105, N1671);
not NOT1 (N2822, N2821);
nor NOR3 (N2823, N2804, N1327, N2430);
buf BUF1 (N2824, N2815);
and AND4 (N2825, N2824, N83, N1976, N396);
nand NAND2 (N2826, N2825, N1928);
not NOT1 (N2827, N2820);
nor NOR2 (N2828, N2794, N1337);
xor XOR2 (N2829, N2823, N1626);
not NOT1 (N2830, N2803);
xor XOR2 (N2831, N2822, N1473);
nand NAND4 (N2832, N2828, N2357, N2446, N499);
buf BUF1 (N2833, N2827);
not NOT1 (N2834, N2811);
nor NOR3 (N2835, N2831, N1586, N2217);
xor XOR2 (N2836, N2807, N1691);
xor XOR2 (N2837, N2826, N2635);
and AND2 (N2838, N2834, N628);
nor NOR4 (N2839, N2830, N722, N569, N1840);
nor NOR4 (N2840, N2819, N866, N469, N1951);
buf BUF1 (N2841, N2829);
nor NOR4 (N2842, N2835, N1046, N2008, N1686);
or OR3 (N2843, N2839, N1600, N1774);
buf BUF1 (N2844, N2832);
xor XOR2 (N2845, N2838, N1985);
nand NAND4 (N2846, N2837, N843, N840, N242);
or OR4 (N2847, N2840, N2518, N242, N2275);
and AND4 (N2848, N2846, N2404, N1102, N2580);
or OR2 (N2849, N2833, N2688);
xor XOR2 (N2850, N2843, N385);
or OR4 (N2851, N2841, N328, N679, N2114);
nand NAND2 (N2852, N2849, N2524);
not NOT1 (N2853, N2851);
nand NAND4 (N2854, N2845, N670, N1164, N2024);
and AND3 (N2855, N2854, N544, N214);
nand NAND4 (N2856, N2853, N1840, N1579, N669);
not NOT1 (N2857, N2856);
nor NOR2 (N2858, N2857, N1987);
not NOT1 (N2859, N2855);
nand NAND3 (N2860, N2848, N2741, N2491);
and AND4 (N2861, N2836, N517, N2503, N2561);
buf BUF1 (N2862, N2847);
not NOT1 (N2863, N2852);
not NOT1 (N2864, N2859);
nor NOR4 (N2865, N2862, N2525, N729, N1286);
or OR2 (N2866, N2858, N301);
nor NOR2 (N2867, N2842, N1853);
xor XOR2 (N2868, N2864, N1106);
or OR3 (N2869, N2861, N1952, N1744);
and AND2 (N2870, N2863, N775);
xor XOR2 (N2871, N2865, N1125);
or OR4 (N2872, N2869, N2594, N1506, N1580);
nand NAND2 (N2873, N2850, N2163);
and AND4 (N2874, N2870, N1576, N83, N1760);
nor NOR4 (N2875, N2868, N2116, N1931, N998);
or OR3 (N2876, N2874, N538, N2105);
nor NOR2 (N2877, N2872, N1676);
or OR3 (N2878, N2860, N2580, N1415);
nor NOR3 (N2879, N2877, N336, N351);
buf BUF1 (N2880, N2875);
and AND2 (N2881, N2871, N2371);
nor NOR4 (N2882, N2879, N2513, N1361, N2226);
and AND3 (N2883, N2817, N472, N1973);
not NOT1 (N2884, N2878);
nor NOR2 (N2885, N2873, N1763);
nand NAND2 (N2886, N2880, N2017);
nor NOR3 (N2887, N2885, N1426, N2393);
nand NAND3 (N2888, N2887, N1832, N2665);
buf BUF1 (N2889, N2884);
and AND2 (N2890, N2882, N1374);
nand NAND2 (N2891, N2890, N669);
buf BUF1 (N2892, N2844);
and AND3 (N2893, N2866, N28, N1008);
not NOT1 (N2894, N2893);
nand NAND4 (N2895, N2867, N2734, N460, N2792);
not NOT1 (N2896, N2889);
and AND2 (N2897, N2876, N1000);
xor XOR2 (N2898, N2883, N492);
nor NOR4 (N2899, N2898, N2400, N1774, N2050);
nand NAND2 (N2900, N2899, N2268);
or OR3 (N2901, N2896, N676, N2069);
or OR4 (N2902, N2886, N1852, N687, N1714);
buf BUF1 (N2903, N2891);
and AND3 (N2904, N2902, N2118, N250);
nand NAND3 (N2905, N2894, N916, N2374);
buf BUF1 (N2906, N2897);
xor XOR2 (N2907, N2904, N52);
buf BUF1 (N2908, N2888);
and AND4 (N2909, N2906, N2637, N999, N2347);
buf BUF1 (N2910, N2907);
or OR2 (N2911, N2881, N333);
not NOT1 (N2912, N2908);
nor NOR3 (N2913, N2909, N1242, N1292);
nor NOR3 (N2914, N2903, N919, N468);
and AND3 (N2915, N2913, N1967, N2260);
buf BUF1 (N2916, N2900);
buf BUF1 (N2917, N2895);
xor XOR2 (N2918, N2914, N2473);
or OR3 (N2919, N2892, N1373, N1627);
not NOT1 (N2920, N2910);
or OR4 (N2921, N2918, N2705, N101, N1562);
nand NAND3 (N2922, N2919, N689, N1265);
or OR3 (N2923, N2921, N2212, N2180);
nand NAND2 (N2924, N2920, N2764);
nand NAND4 (N2925, N2922, N1869, N705, N1547);
or OR2 (N2926, N2916, N2620);
nand NAND3 (N2927, N2915, N2721, N1212);
nand NAND2 (N2928, N2926, N514);
or OR4 (N2929, N2911, N2601, N2113, N760);
not NOT1 (N2930, N2905);
not NOT1 (N2931, N2923);
buf BUF1 (N2932, N2924);
buf BUF1 (N2933, N2932);
not NOT1 (N2934, N2927);
nand NAND2 (N2935, N2928, N1788);
and AND3 (N2936, N2917, N33, N2812);
not NOT1 (N2937, N2925);
buf BUF1 (N2938, N2935);
nand NAND4 (N2939, N2901, N2336, N51, N1258);
nor NOR3 (N2940, N2939, N2738, N250);
buf BUF1 (N2941, N2929);
not NOT1 (N2942, N2931);
buf BUF1 (N2943, N2936);
xor XOR2 (N2944, N2912, N622);
and AND3 (N2945, N2942, N2101, N853);
nor NOR4 (N2946, N2937, N1331, N950, N1100);
nand NAND4 (N2947, N2943, N1351, N192, N1401);
not NOT1 (N2948, N2930);
or OR4 (N2949, N2940, N811, N1848, N1621);
nor NOR2 (N2950, N2949, N1661);
buf BUF1 (N2951, N2947);
or OR2 (N2952, N2951, N771);
xor XOR2 (N2953, N2933, N2662);
xor XOR2 (N2954, N2945, N616);
nor NOR4 (N2955, N2948, N2642, N653, N1040);
nor NOR4 (N2956, N2934, N2668, N2229, N1049);
or OR3 (N2957, N2944, N389, N463);
or OR3 (N2958, N2954, N69, N2380);
nand NAND2 (N2959, N2953, N2853);
xor XOR2 (N2960, N2955, N1227);
and AND2 (N2961, N2959, N1912);
nor NOR2 (N2962, N2950, N2908);
nand NAND4 (N2963, N2962, N1350, N1704, N825);
buf BUF1 (N2964, N2938);
buf BUF1 (N2965, N2952);
nor NOR3 (N2966, N2961, N2403, N2560);
and AND4 (N2967, N2958, N1867, N1050, N2748);
xor XOR2 (N2968, N2965, N708);
not NOT1 (N2969, N2963);
or OR3 (N2970, N2960, N2847, N2745);
nand NAND2 (N2971, N2967, N967);
and AND4 (N2972, N2957, N1675, N2753, N803);
and AND3 (N2973, N2970, N1890, N1629);
xor XOR2 (N2974, N2956, N2109);
or OR3 (N2975, N2966, N2471, N42);
not NOT1 (N2976, N2968);
nor NOR3 (N2977, N2969, N2165, N1251);
or OR4 (N2978, N2975, N2506, N1929, N356);
buf BUF1 (N2979, N2941);
buf BUF1 (N2980, N2976);
not NOT1 (N2981, N2971);
xor XOR2 (N2982, N2980, N2258);
or OR2 (N2983, N2974, N1653);
and AND2 (N2984, N2978, N64);
or OR3 (N2985, N2977, N880, N658);
and AND2 (N2986, N2985, N960);
nor NOR4 (N2987, N2972, N212, N1981, N2837);
buf BUF1 (N2988, N2986);
nor NOR3 (N2989, N2983, N1440, N60);
nand NAND2 (N2990, N2973, N245);
or OR3 (N2991, N2989, N2628, N2646);
xor XOR2 (N2992, N2946, N1661);
nand NAND2 (N2993, N2991, N322);
and AND2 (N2994, N2982, N2817);
buf BUF1 (N2995, N2984);
nor NOR2 (N2996, N2964, N2349);
xor XOR2 (N2997, N2996, N2221);
buf BUF1 (N2998, N2987);
and AND4 (N2999, N2979, N1039, N2583, N2724);
nand NAND3 (N3000, N2993, N1565, N2571);
not NOT1 (N3001, N2992);
xor XOR2 (N3002, N2998, N2473);
nor NOR3 (N3003, N2988, N1502, N62);
buf BUF1 (N3004, N3000);
nand NAND4 (N3005, N2981, N1367, N2391, N2026);
or OR3 (N3006, N3002, N223, N404);
not NOT1 (N3007, N3003);
xor XOR2 (N3008, N2999, N888);
and AND3 (N3009, N2997, N1162, N162);
not NOT1 (N3010, N3005);
and AND4 (N3011, N2990, N242, N2797, N1404);
nand NAND2 (N3012, N3007, N110);
nand NAND3 (N3013, N3012, N686, N1018);
or OR2 (N3014, N2995, N1626);
nor NOR3 (N3015, N3013, N1636, N1276);
xor XOR2 (N3016, N3004, N2360);
nand NAND3 (N3017, N3006, N514, N2631);
and AND2 (N3018, N3010, N1420);
and AND2 (N3019, N3001, N2473);
and AND3 (N3020, N3019, N2536, N2482);
xor XOR2 (N3021, N3014, N260);
nor NOR2 (N3022, N3015, N2903);
nand NAND4 (N3023, N3017, N3001, N576, N1110);
not NOT1 (N3024, N3009);
nand NAND2 (N3025, N3008, N1588);
xor XOR2 (N3026, N3021, N2326);
not NOT1 (N3027, N3016);
not NOT1 (N3028, N3023);
and AND2 (N3029, N3026, N2492);
not NOT1 (N3030, N3018);
not NOT1 (N3031, N3028);
nand NAND4 (N3032, N3020, N1598, N822, N1259);
or OR3 (N3033, N3024, N120, N56);
nand NAND4 (N3034, N3011, N1530, N2872, N1344);
nor NOR4 (N3035, N3022, N210, N1063, N2174);
not NOT1 (N3036, N3030);
not NOT1 (N3037, N3029);
or OR4 (N3038, N3031, N1799, N1135, N2433);
nor NOR3 (N3039, N3034, N398, N447);
or OR2 (N3040, N3025, N1037);
xor XOR2 (N3041, N3040, N2509);
nor NOR2 (N3042, N3038, N1803);
nand NAND4 (N3043, N3042, N2595, N1058, N1189);
buf BUF1 (N3044, N3035);
and AND3 (N3045, N3041, N1485, N791);
nor NOR4 (N3046, N3027, N1599, N2351, N61);
and AND2 (N3047, N3039, N2731);
not NOT1 (N3048, N3033);
xor XOR2 (N3049, N3048, N2478);
buf BUF1 (N3050, N3032);
or OR4 (N3051, N3050, N613, N913, N771);
xor XOR2 (N3052, N3046, N1348);
nand NAND3 (N3053, N3043, N2821, N1209);
buf BUF1 (N3054, N3051);
or OR3 (N3055, N3052, N7, N1383);
xor XOR2 (N3056, N3045, N324);
not NOT1 (N3057, N2994);
and AND3 (N3058, N3053, N2808, N337);
nand NAND4 (N3059, N3049, N898, N190, N521);
nand NAND2 (N3060, N3054, N2440);
nand NAND2 (N3061, N3056, N169);
not NOT1 (N3062, N3061);
or OR3 (N3063, N3058, N2925, N2651);
nor NOR4 (N3064, N3057, N2470, N1677, N1042);
or OR4 (N3065, N3063, N1443, N1962, N1700);
not NOT1 (N3066, N3055);
buf BUF1 (N3067, N3044);
and AND2 (N3068, N3047, N182);
not NOT1 (N3069, N3060);
nand NAND3 (N3070, N3069, N1429, N3026);
buf BUF1 (N3071, N3064);
not NOT1 (N3072, N3036);
or OR2 (N3073, N3062, N2353);
buf BUF1 (N3074, N3067);
or OR2 (N3075, N3074, N767);
and AND3 (N3076, N3075, N125, N260);
buf BUF1 (N3077, N3073);
buf BUF1 (N3078, N3059);
not NOT1 (N3079, N3037);
or OR3 (N3080, N3077, N304, N2021);
or OR3 (N3081, N3071, N47, N1729);
or OR3 (N3082, N3070, N993, N2473);
nand NAND3 (N3083, N3079, N724, N196);
nand NAND3 (N3084, N3076, N1022, N866);
nand NAND2 (N3085, N3072, N1466);
buf BUF1 (N3086, N3078);
or OR2 (N3087, N3081, N461);
buf BUF1 (N3088, N3080);
nor NOR2 (N3089, N3086, N1032);
not NOT1 (N3090, N3089);
and AND3 (N3091, N3083, N2587, N2804);
nor NOR3 (N3092, N3090, N26, N177);
and AND4 (N3093, N3092, N3083, N376, N2231);
nor NOR2 (N3094, N3087, N2964);
nand NAND3 (N3095, N3091, N1432, N1468);
buf BUF1 (N3096, N3094);
not NOT1 (N3097, N3093);
xor XOR2 (N3098, N3096, N2074);
or OR4 (N3099, N3066, N1731, N117, N1227);
not NOT1 (N3100, N3082);
and AND4 (N3101, N3100, N1215, N2860, N76);
not NOT1 (N3102, N3095);
or OR4 (N3103, N3099, N605, N2883, N1706);
or OR2 (N3104, N3103, N349);
nor NOR4 (N3105, N3085, N2374, N2072, N1902);
or OR4 (N3106, N3105, N1864, N2464, N75);
and AND2 (N3107, N3097, N580);
not NOT1 (N3108, N3102);
or OR2 (N3109, N3107, N231);
and AND3 (N3110, N3108, N1237, N2295);
not NOT1 (N3111, N3110);
not NOT1 (N3112, N3106);
and AND3 (N3113, N3065, N2519, N2958);
nor NOR3 (N3114, N3088, N1989, N484);
xor XOR2 (N3115, N3113, N2534);
and AND3 (N3116, N3068, N2769, N914);
not NOT1 (N3117, N3114);
xor XOR2 (N3118, N3109, N2723);
and AND3 (N3119, N3116, N1244, N2230);
xor XOR2 (N3120, N3118, N2553);
not NOT1 (N3121, N3101);
buf BUF1 (N3122, N3098);
xor XOR2 (N3123, N3120, N617);
and AND4 (N3124, N3112, N2019, N1345, N704);
or OR2 (N3125, N3121, N2686);
not NOT1 (N3126, N3104);
nor NOR3 (N3127, N3084, N1411, N2425);
or OR3 (N3128, N3123, N499, N691);
nor NOR2 (N3129, N3117, N664);
and AND2 (N3130, N3126, N654);
xor XOR2 (N3131, N3127, N1613);
buf BUF1 (N3132, N3122);
not NOT1 (N3133, N3111);
not NOT1 (N3134, N3131);
buf BUF1 (N3135, N3125);
not NOT1 (N3136, N3132);
nor NOR4 (N3137, N3130, N1948, N1388, N571);
nand NAND3 (N3138, N3137, N1053, N871);
and AND4 (N3139, N3124, N1844, N184, N1212);
not NOT1 (N3140, N3129);
nand NAND3 (N3141, N3140, N1119, N2835);
nand NAND3 (N3142, N3136, N2091, N1753);
buf BUF1 (N3143, N3142);
nand NAND2 (N3144, N3119, N2041);
not NOT1 (N3145, N3144);
not NOT1 (N3146, N3128);
buf BUF1 (N3147, N3115);
nand NAND2 (N3148, N3138, N252);
and AND2 (N3149, N3133, N842);
nor NOR4 (N3150, N3143, N2871, N461, N1378);
buf BUF1 (N3151, N3141);
or OR4 (N3152, N3148, N1756, N1047, N2547);
nand NAND4 (N3153, N3146, N214, N1916, N2871);
buf BUF1 (N3154, N3149);
xor XOR2 (N3155, N3151, N1075);
buf BUF1 (N3156, N3153);
nand NAND3 (N3157, N3134, N504, N2491);
buf BUF1 (N3158, N3139);
not NOT1 (N3159, N3147);
xor XOR2 (N3160, N3158, N1251);
and AND4 (N3161, N3154, N2990, N2616, N2453);
xor XOR2 (N3162, N3161, N2545);
and AND4 (N3163, N3152, N2590, N2902, N2629);
or OR3 (N3164, N3159, N697, N249);
buf BUF1 (N3165, N3135);
not NOT1 (N3166, N3156);
buf BUF1 (N3167, N3162);
nand NAND2 (N3168, N3165, N2580);
nor NOR3 (N3169, N3167, N2723, N1122);
buf BUF1 (N3170, N3155);
or OR2 (N3171, N3164, N2814);
and AND4 (N3172, N3157, N2397, N1194, N2191);
and AND2 (N3173, N3166, N2111);
nor NOR4 (N3174, N3170, N1325, N1157, N524);
xor XOR2 (N3175, N3172, N2137);
nor NOR3 (N3176, N3168, N1706, N2532);
not NOT1 (N3177, N3171);
and AND4 (N3178, N3160, N1927, N1527, N1447);
not NOT1 (N3179, N3175);
and AND3 (N3180, N3178, N1930, N2057);
nor NOR2 (N3181, N3163, N182);
and AND3 (N3182, N3169, N2946, N665);
not NOT1 (N3183, N3174);
and AND3 (N3184, N3145, N500, N2196);
nor NOR4 (N3185, N3182, N2120, N2415, N947);
nor NOR3 (N3186, N3179, N1277, N2568);
xor XOR2 (N3187, N3150, N330);
xor XOR2 (N3188, N3187, N1438);
buf BUF1 (N3189, N3184);
nor NOR4 (N3190, N3173, N3016, N29, N1320);
not NOT1 (N3191, N3189);
and AND4 (N3192, N3177, N934, N603, N376);
xor XOR2 (N3193, N3180, N915);
buf BUF1 (N3194, N3176);
buf BUF1 (N3195, N3183);
and AND2 (N3196, N3188, N3005);
buf BUF1 (N3197, N3181);
xor XOR2 (N3198, N3186, N1493);
buf BUF1 (N3199, N3196);
nand NAND4 (N3200, N3199, N2698, N2170, N2431);
nor NOR4 (N3201, N3194, N1092, N866, N519);
and AND3 (N3202, N3200, N1602, N2558);
not NOT1 (N3203, N3190);
not NOT1 (N3204, N3193);
and AND2 (N3205, N3204, N802);
not NOT1 (N3206, N3192);
and AND4 (N3207, N3202, N74, N2081, N3181);
xor XOR2 (N3208, N3205, N1109);
xor XOR2 (N3209, N3207, N1162);
and AND3 (N3210, N3203, N704, N793);
nor NOR3 (N3211, N3191, N1888, N2065);
not NOT1 (N3212, N3211);
buf BUF1 (N3213, N3198);
nor NOR3 (N3214, N3206, N1548, N186);
not NOT1 (N3215, N3201);
nand NAND4 (N3216, N3210, N690, N3203, N1043);
xor XOR2 (N3217, N3212, N2163);
not NOT1 (N3218, N3214);
nand NAND3 (N3219, N3218, N2794, N1910);
nand NAND3 (N3220, N3185, N2322, N1873);
and AND4 (N3221, N3213, N1360, N3079, N2112);
xor XOR2 (N3222, N3208, N2506);
buf BUF1 (N3223, N3222);
and AND3 (N3224, N3223, N1347, N2853);
nand NAND2 (N3225, N3219, N1426);
nand NAND3 (N3226, N3220, N2629, N247);
xor XOR2 (N3227, N3226, N1014);
buf BUF1 (N3228, N3227);
buf BUF1 (N3229, N3228);
xor XOR2 (N3230, N3225, N858);
not NOT1 (N3231, N3224);
not NOT1 (N3232, N3216);
xor XOR2 (N3233, N3217, N1812);
nor NOR2 (N3234, N3221, N1663);
and AND4 (N3235, N3215, N940, N101, N528);
or OR2 (N3236, N3231, N2916);
not NOT1 (N3237, N3197);
nand NAND3 (N3238, N3235, N1139, N2035);
or OR3 (N3239, N3232, N282, N1046);
buf BUF1 (N3240, N3233);
nor NOR3 (N3241, N3240, N1542, N2652);
nand NAND4 (N3242, N3238, N1522, N1019, N2395);
not NOT1 (N3243, N3237);
xor XOR2 (N3244, N3241, N439);
xor XOR2 (N3245, N3195, N2277);
and AND3 (N3246, N3230, N3007, N1581);
nand NAND4 (N3247, N3234, N927, N1498, N2726);
buf BUF1 (N3248, N3245);
xor XOR2 (N3249, N3247, N668);
not NOT1 (N3250, N3248);
and AND4 (N3251, N3209, N1529, N2892, N620);
nand NAND3 (N3252, N3242, N1971, N1289);
xor XOR2 (N3253, N3239, N2855);
nor NOR2 (N3254, N3251, N1974);
nand NAND4 (N3255, N3252, N1576, N322, N612);
xor XOR2 (N3256, N3249, N294);
nand NAND3 (N3257, N3243, N2016, N2855);
buf BUF1 (N3258, N3254);
and AND4 (N3259, N3258, N2645, N936, N3056);
nor NOR3 (N3260, N3250, N1000, N2024);
or OR4 (N3261, N3244, N292, N792, N1709);
nor NOR4 (N3262, N3253, N2256, N1358, N3237);
not NOT1 (N3263, N3257);
buf BUF1 (N3264, N3236);
buf BUF1 (N3265, N3262);
nand NAND2 (N3266, N3260, N1870);
or OR3 (N3267, N3261, N126, N1782);
nand NAND3 (N3268, N3256, N1724, N12);
not NOT1 (N3269, N3266);
buf BUF1 (N3270, N3269);
not NOT1 (N3271, N3268);
or OR2 (N3272, N3265, N27);
not NOT1 (N3273, N3263);
or OR3 (N3274, N3255, N1434, N1097);
xor XOR2 (N3275, N3246, N1256);
not NOT1 (N3276, N3270);
or OR3 (N3277, N3273, N1309, N758);
buf BUF1 (N3278, N3277);
and AND4 (N3279, N3276, N2360, N2864, N1442);
nand NAND3 (N3280, N3278, N1969, N2594);
not NOT1 (N3281, N3274);
nand NAND2 (N3282, N3259, N1088);
not NOT1 (N3283, N3282);
buf BUF1 (N3284, N3281);
nor NOR2 (N3285, N3283, N2647);
or OR4 (N3286, N3272, N102, N519, N287);
or OR2 (N3287, N3286, N1584);
nor NOR2 (N3288, N3267, N1238);
xor XOR2 (N3289, N3285, N1303);
not NOT1 (N3290, N3264);
or OR4 (N3291, N3229, N2015, N420, N1610);
or OR4 (N3292, N3271, N1172, N1873, N2139);
nand NAND4 (N3293, N3290, N947, N312, N935);
and AND3 (N3294, N3280, N1498, N1063);
and AND4 (N3295, N3294, N1658, N2892, N2403);
xor XOR2 (N3296, N3279, N428);
and AND4 (N3297, N3288, N2052, N1741, N127);
buf BUF1 (N3298, N3297);
buf BUF1 (N3299, N3298);
nand NAND3 (N3300, N3291, N2037, N2480);
or OR4 (N3301, N3296, N729, N2667, N2575);
or OR2 (N3302, N3287, N1210);
xor XOR2 (N3303, N3293, N2605);
or OR3 (N3304, N3303, N2094, N1009);
or OR2 (N3305, N3275, N2);
xor XOR2 (N3306, N3305, N1220);
nor NOR4 (N3307, N3300, N698, N2496, N2339);
xor XOR2 (N3308, N3289, N1775);
nand NAND2 (N3309, N3284, N430);
or OR4 (N3310, N3304, N812, N2825, N3248);
or OR3 (N3311, N3301, N910, N669);
nor NOR3 (N3312, N3292, N1395, N1688);
and AND2 (N3313, N3295, N2572);
xor XOR2 (N3314, N3309, N2723);
and AND3 (N3315, N3314, N1043, N1121);
nor NOR4 (N3316, N3313, N2029, N950, N606);
or OR4 (N3317, N3299, N1521, N526, N2847);
or OR2 (N3318, N3311, N2633);
xor XOR2 (N3319, N3318, N1521);
nand NAND4 (N3320, N3308, N1477, N1816, N2453);
not NOT1 (N3321, N3312);
nor NOR4 (N3322, N3316, N726, N3236, N2705);
and AND2 (N3323, N3302, N2240);
and AND3 (N3324, N3322, N97, N277);
not NOT1 (N3325, N3320);
nor NOR2 (N3326, N3321, N2144);
not NOT1 (N3327, N3307);
or OR2 (N3328, N3326, N3121);
nor NOR2 (N3329, N3328, N687);
nor NOR3 (N3330, N3319, N3106, N3224);
buf BUF1 (N3331, N3306);
and AND2 (N3332, N3315, N1381);
xor XOR2 (N3333, N3332, N935);
nand NAND4 (N3334, N3317, N2108, N3194, N3306);
or OR2 (N3335, N3323, N2606);
buf BUF1 (N3336, N3330);
and AND2 (N3337, N3329, N62);
nand NAND2 (N3338, N3337, N2717);
nand NAND2 (N3339, N3336, N1409);
nor NOR3 (N3340, N3324, N403, N76);
nand NAND3 (N3341, N3327, N1300, N2335);
xor XOR2 (N3342, N3341, N2581);
not NOT1 (N3343, N3334);
buf BUF1 (N3344, N3331);
and AND3 (N3345, N3344, N2581, N1636);
not NOT1 (N3346, N3325);
xor XOR2 (N3347, N3339, N1825);
xor XOR2 (N3348, N3338, N2067);
or OR4 (N3349, N3348, N2602, N2963, N981);
and AND2 (N3350, N3333, N729);
buf BUF1 (N3351, N3335);
not NOT1 (N3352, N3351);
nand NAND3 (N3353, N3349, N2790, N2897);
and AND4 (N3354, N3342, N3080, N730, N369);
and AND4 (N3355, N3343, N1932, N406, N492);
not NOT1 (N3356, N3345);
nor NOR4 (N3357, N3340, N2859, N2491, N3023);
and AND3 (N3358, N3354, N1026, N1148);
and AND4 (N3359, N3357, N1086, N169, N2811);
and AND2 (N3360, N3353, N2987);
nor NOR2 (N3361, N3356, N3106);
buf BUF1 (N3362, N3360);
nor NOR4 (N3363, N3347, N3245, N1690, N2769);
buf BUF1 (N3364, N3359);
nor NOR2 (N3365, N3355, N1282);
xor XOR2 (N3366, N3361, N3174);
buf BUF1 (N3367, N3350);
buf BUF1 (N3368, N3365);
or OR3 (N3369, N3366, N3113, N147);
nand NAND4 (N3370, N3368, N3043, N2069, N372);
not NOT1 (N3371, N3346);
not NOT1 (N3372, N3367);
not NOT1 (N3373, N3363);
nor NOR3 (N3374, N3370, N1718, N2145);
and AND4 (N3375, N3369, N2885, N1752, N2178);
not NOT1 (N3376, N3358);
or OR2 (N3377, N3371, N2308);
xor XOR2 (N3378, N3376, N2742);
or OR3 (N3379, N3362, N268, N349);
xor XOR2 (N3380, N3375, N539);
or OR2 (N3381, N3352, N2830);
or OR3 (N3382, N3374, N3140, N333);
not NOT1 (N3383, N3310);
or OR3 (N3384, N3364, N2812, N395);
nand NAND4 (N3385, N3384, N299, N1841, N2387);
nand NAND3 (N3386, N3380, N2003, N188);
or OR4 (N3387, N3373, N3174, N488, N2543);
nand NAND2 (N3388, N3378, N2777);
xor XOR2 (N3389, N3386, N3321);
nor NOR3 (N3390, N3379, N1326, N2631);
not NOT1 (N3391, N3390);
or OR2 (N3392, N3377, N1233);
nor NOR2 (N3393, N3388, N1729);
or OR2 (N3394, N3385, N1833);
not NOT1 (N3395, N3372);
not NOT1 (N3396, N3382);
nor NOR3 (N3397, N3392, N454, N638);
not NOT1 (N3398, N3381);
buf BUF1 (N3399, N3391);
nor NOR3 (N3400, N3399, N87, N2591);
or OR4 (N3401, N3387, N217, N2524, N3156);
nand NAND4 (N3402, N3383, N1623, N1658, N1189);
nand NAND3 (N3403, N3398, N2412, N1143);
or OR3 (N3404, N3397, N990, N2539);
xor XOR2 (N3405, N3403, N404);
buf BUF1 (N3406, N3401);
nand NAND2 (N3407, N3400, N1946);
nor NOR4 (N3408, N3395, N3094, N2504, N18);
buf BUF1 (N3409, N3404);
and AND3 (N3410, N3406, N2033, N3209);
not NOT1 (N3411, N3410);
nor NOR3 (N3412, N3408, N2522, N53);
and AND2 (N3413, N3393, N1345);
nand NAND4 (N3414, N3409, N1487, N2693, N2567);
xor XOR2 (N3415, N3414, N2547);
or OR4 (N3416, N3402, N1604, N1477, N1773);
or OR2 (N3417, N3413, N1036);
buf BUF1 (N3418, N3412);
nand NAND2 (N3419, N3417, N2715);
buf BUF1 (N3420, N3411);
buf BUF1 (N3421, N3420);
or OR3 (N3422, N3389, N2097, N378);
not NOT1 (N3423, N3418);
buf BUF1 (N3424, N3396);
nor NOR3 (N3425, N3422, N1424, N1579);
and AND4 (N3426, N3394, N2972, N2905, N3320);
xor XOR2 (N3427, N3421, N132);
not NOT1 (N3428, N3427);
or OR3 (N3429, N3426, N1015, N2269);
nand NAND4 (N3430, N3428, N1140, N1117, N2282);
and AND2 (N3431, N3405, N340);
xor XOR2 (N3432, N3430, N1781);
nand NAND2 (N3433, N3432, N2324);
nor NOR2 (N3434, N3431, N300);
buf BUF1 (N3435, N3424);
or OR2 (N3436, N3407, N2358);
and AND4 (N3437, N3433, N1833, N1536, N1955);
or OR2 (N3438, N3415, N2960);
buf BUF1 (N3439, N3437);
nand NAND4 (N3440, N3423, N3076, N2611, N697);
not NOT1 (N3441, N3435);
and AND2 (N3442, N3439, N2354);
not NOT1 (N3443, N3440);
xor XOR2 (N3444, N3441, N2620);
not NOT1 (N3445, N3444);
or OR2 (N3446, N3445, N1635);
not NOT1 (N3447, N3443);
xor XOR2 (N3448, N3425, N3117);
or OR3 (N3449, N3447, N2353, N713);
not NOT1 (N3450, N3446);
or OR4 (N3451, N3429, N1195, N1349, N34);
nand NAND3 (N3452, N3436, N304, N2616);
nor NOR3 (N3453, N3442, N225, N3346);
not NOT1 (N3454, N3452);
or OR4 (N3455, N3453, N161, N2559, N3145);
or OR2 (N3456, N3450, N2761);
or OR4 (N3457, N3434, N1739, N982, N323);
or OR3 (N3458, N3448, N383, N660);
and AND4 (N3459, N3457, N902, N1491, N1287);
not NOT1 (N3460, N3454);
and AND3 (N3461, N3458, N1519, N172);
not NOT1 (N3462, N3461);
not NOT1 (N3463, N3460);
or OR4 (N3464, N3416, N649, N922, N3126);
not NOT1 (N3465, N3438);
nand NAND3 (N3466, N3449, N1536, N939);
and AND4 (N3467, N3455, N2100, N1520, N1262);
not NOT1 (N3468, N3466);
or OR3 (N3469, N3459, N1861, N2209);
and AND4 (N3470, N3456, N1469, N809, N714);
and AND2 (N3471, N3419, N2200);
or OR4 (N3472, N3467, N1814, N2726, N1205);
and AND4 (N3473, N3472, N2505, N383, N2921);
buf BUF1 (N3474, N3465);
nand NAND4 (N3475, N3468, N3006, N2909, N2740);
not NOT1 (N3476, N3471);
nand NAND2 (N3477, N3451, N1661);
or OR4 (N3478, N3464, N2917, N730, N768);
xor XOR2 (N3479, N3473, N2334);
xor XOR2 (N3480, N3469, N149);
nor NOR3 (N3481, N3475, N1107, N1526);
not NOT1 (N3482, N3476);
not NOT1 (N3483, N3482);
or OR2 (N3484, N3470, N1329);
not NOT1 (N3485, N3483);
nand NAND2 (N3486, N3463, N2552);
xor XOR2 (N3487, N3481, N2915);
or OR4 (N3488, N3479, N801, N386, N3025);
and AND2 (N3489, N3484, N193);
or OR2 (N3490, N3478, N1360);
or OR2 (N3491, N3474, N1827);
or OR2 (N3492, N3462, N2283);
xor XOR2 (N3493, N3490, N2026);
buf BUF1 (N3494, N3485);
and AND4 (N3495, N3480, N2708, N536, N3375);
or OR2 (N3496, N3493, N2093);
nand NAND4 (N3497, N3495, N2878, N783, N1117);
and AND3 (N3498, N3494, N942, N1303);
not NOT1 (N3499, N3489);
xor XOR2 (N3500, N3498, N1345);
buf BUF1 (N3501, N3497);
not NOT1 (N3502, N3488);
nor NOR3 (N3503, N3492, N2682, N384);
and AND4 (N3504, N3502, N2784, N1161, N2939);
nor NOR2 (N3505, N3477, N2616);
not NOT1 (N3506, N3505);
or OR3 (N3507, N3500, N467, N1132);
and AND2 (N3508, N3496, N2384);
and AND2 (N3509, N3507, N2866);
xor XOR2 (N3510, N3491, N2550);
buf BUF1 (N3511, N3508);
or OR3 (N3512, N3487, N3058, N691);
or OR2 (N3513, N3499, N2118);
nand NAND3 (N3514, N3503, N2728, N2572);
nor NOR4 (N3515, N3512, N724, N709, N2560);
or OR2 (N3516, N3513, N1199);
and AND4 (N3517, N3510, N1283, N257, N1964);
or OR4 (N3518, N3509, N2985, N22, N2291);
not NOT1 (N3519, N3515);
nand NAND2 (N3520, N3516, N2698);
buf BUF1 (N3521, N3511);
nand NAND2 (N3522, N3486, N114);
buf BUF1 (N3523, N3520);
xor XOR2 (N3524, N3506, N337);
buf BUF1 (N3525, N3522);
not NOT1 (N3526, N3523);
xor XOR2 (N3527, N3524, N1424);
nand NAND3 (N3528, N3526, N3340, N2069);
nor NOR4 (N3529, N3519, N1893, N842, N2261);
xor XOR2 (N3530, N3517, N342);
or OR2 (N3531, N3527, N378);
and AND3 (N3532, N3514, N1537, N306);
or OR2 (N3533, N3501, N2799);
buf BUF1 (N3534, N3533);
and AND3 (N3535, N3534, N161, N68);
not NOT1 (N3536, N3521);
nand NAND2 (N3537, N3529, N394);
and AND4 (N3538, N3504, N2818, N449, N2348);
xor XOR2 (N3539, N3525, N1169);
xor XOR2 (N3540, N3530, N762);
nand NAND2 (N3541, N3536, N2672);
buf BUF1 (N3542, N3518);
xor XOR2 (N3543, N3535, N547);
and AND4 (N3544, N3537, N2668, N2702, N1467);
and AND3 (N3545, N3532, N1409, N8);
nor NOR3 (N3546, N3541, N1919, N1577);
xor XOR2 (N3547, N3546, N2629);
nand NAND2 (N3548, N3545, N1041);
nand NAND4 (N3549, N3542, N1598, N2071, N2591);
nand NAND4 (N3550, N3544, N447, N2003, N2599);
buf BUF1 (N3551, N3540);
or OR3 (N3552, N3531, N1756, N3137);
or OR4 (N3553, N3547, N733, N1790, N1433);
nand NAND2 (N3554, N3543, N1232);
nor NOR4 (N3555, N3552, N1491, N1256, N238);
nand NAND3 (N3556, N3551, N945, N1189);
buf BUF1 (N3557, N3548);
not NOT1 (N3558, N3528);
or OR2 (N3559, N3555, N3496);
nand NAND4 (N3560, N3554, N1528, N2997, N252);
xor XOR2 (N3561, N3539, N2207);
nor NOR2 (N3562, N3538, N3016);
buf BUF1 (N3563, N3556);
not NOT1 (N3564, N3563);
nor NOR4 (N3565, N3562, N1857, N2432, N1145);
not NOT1 (N3566, N3559);
nor NOR4 (N3567, N3560, N1178, N2509, N3239);
nor NOR4 (N3568, N3567, N3447, N3171, N81);
xor XOR2 (N3569, N3566, N383);
nor NOR3 (N3570, N3557, N1536, N92);
nor NOR3 (N3571, N3553, N966, N1885);
nor NOR2 (N3572, N3569, N1065);
not NOT1 (N3573, N3570);
or OR4 (N3574, N3549, N3001, N1726, N2481);
or OR2 (N3575, N3561, N3303);
xor XOR2 (N3576, N3558, N1890);
not NOT1 (N3577, N3575);
nand NAND3 (N3578, N3565, N927, N1585);
buf BUF1 (N3579, N3571);
or OR4 (N3580, N3572, N1567, N2246, N1173);
or OR4 (N3581, N3573, N664, N2019, N1212);
or OR4 (N3582, N3577, N191, N2122, N786);
not NOT1 (N3583, N3580);
not NOT1 (N3584, N3576);
xor XOR2 (N3585, N3584, N2649);
not NOT1 (N3586, N3550);
and AND3 (N3587, N3583, N2229, N217);
or OR4 (N3588, N3581, N2757, N542, N3344);
and AND3 (N3589, N3587, N2867, N3323);
buf BUF1 (N3590, N3589);
xor XOR2 (N3591, N3586, N1460);
not NOT1 (N3592, N3564);
not NOT1 (N3593, N3568);
nand NAND4 (N3594, N3578, N448, N1810, N1036);
nand NAND4 (N3595, N3574, N1210, N3380, N101);
not NOT1 (N3596, N3582);
nand NAND4 (N3597, N3588, N751, N1973, N2916);
nand NAND4 (N3598, N3579, N889, N1942, N1223);
nand NAND2 (N3599, N3596, N2097);
buf BUF1 (N3600, N3595);
not NOT1 (N3601, N3591);
not NOT1 (N3602, N3592);
xor XOR2 (N3603, N3601, N25);
and AND4 (N3604, N3593, N3143, N2623, N2407);
buf BUF1 (N3605, N3590);
not NOT1 (N3606, N3602);
or OR3 (N3607, N3606, N3221, N1267);
nand NAND2 (N3608, N3599, N1756);
buf BUF1 (N3609, N3603);
not NOT1 (N3610, N3609);
xor XOR2 (N3611, N3600, N2212);
or OR4 (N3612, N3604, N3583, N1071, N271);
not NOT1 (N3613, N3605);
xor XOR2 (N3614, N3594, N2992);
or OR3 (N3615, N3608, N2019, N1793);
and AND4 (N3616, N3615, N2247, N3370, N1125);
nor NOR3 (N3617, N3616, N429, N2023);
nor NOR2 (N3618, N3612, N342);
buf BUF1 (N3619, N3610);
xor XOR2 (N3620, N3619, N321);
and AND4 (N3621, N3620, N3071, N2551, N2008);
xor XOR2 (N3622, N3614, N596);
nand NAND4 (N3623, N3618, N3363, N193, N3098);
nor NOR3 (N3624, N3617, N1656, N1599);
nand NAND3 (N3625, N3623, N1969, N270);
and AND4 (N3626, N3585, N633, N2302, N855);
nand NAND3 (N3627, N3607, N3616, N1092);
and AND3 (N3628, N3598, N1889, N2604);
or OR4 (N3629, N3611, N2947, N2263, N2194);
not NOT1 (N3630, N3629);
xor XOR2 (N3631, N3625, N3568);
not NOT1 (N3632, N3622);
buf BUF1 (N3633, N3631);
nand NAND3 (N3634, N3627, N2217, N1029);
xor XOR2 (N3635, N3628, N630);
and AND4 (N3636, N3635, N2059, N1584, N1499);
buf BUF1 (N3637, N3633);
or OR2 (N3638, N3597, N3483);
xor XOR2 (N3639, N3632, N3210);
nand NAND4 (N3640, N3637, N448, N3357, N544);
buf BUF1 (N3641, N3639);
nor NOR3 (N3642, N3630, N2055, N928);
not NOT1 (N3643, N3640);
xor XOR2 (N3644, N3636, N3240);
nand NAND2 (N3645, N3624, N1178);
and AND4 (N3646, N3644, N461, N2510, N3205);
nor NOR2 (N3647, N3646, N938);
nor NOR2 (N3648, N3621, N2529);
and AND3 (N3649, N3642, N872, N3346);
or OR2 (N3650, N3626, N606);
nor NOR3 (N3651, N3638, N54, N1852);
xor XOR2 (N3652, N3643, N978);
and AND2 (N3653, N3651, N2758);
nand NAND4 (N3654, N3648, N843, N3486, N2592);
nor NOR3 (N3655, N3649, N2547, N6);
not NOT1 (N3656, N3634);
or OR3 (N3657, N3653, N3176, N1357);
not NOT1 (N3658, N3654);
xor XOR2 (N3659, N3650, N1835);
nor NOR4 (N3660, N3647, N2701, N2105, N1632);
nor NOR4 (N3661, N3656, N3086, N604, N1714);
not NOT1 (N3662, N3613);
nor NOR4 (N3663, N3662, N3586, N2757, N912);
and AND4 (N3664, N3658, N1604, N1932, N399);
buf BUF1 (N3665, N3659);
not NOT1 (N3666, N3665);
not NOT1 (N3667, N3652);
xor XOR2 (N3668, N3661, N2561);
or OR3 (N3669, N3663, N3562, N2756);
xor XOR2 (N3670, N3669, N795);
nand NAND3 (N3671, N3666, N3554, N845);
nor NOR4 (N3672, N3664, N3349, N2892, N314);
or OR3 (N3673, N3657, N569, N2419);
not NOT1 (N3674, N3645);
xor XOR2 (N3675, N3641, N3332);
nor NOR4 (N3676, N3655, N3315, N696, N1479);
or OR4 (N3677, N3671, N3602, N975, N901);
not NOT1 (N3678, N3674);
and AND4 (N3679, N3660, N2626, N1330, N3472);
and AND3 (N3680, N3675, N1040, N2604);
nor NOR4 (N3681, N3667, N2561, N3500, N3547);
and AND3 (N3682, N3679, N1680, N2791);
nand NAND4 (N3683, N3673, N1905, N3226, N912);
or OR3 (N3684, N3680, N212, N3039);
or OR2 (N3685, N3677, N1730);
nor NOR3 (N3686, N3668, N3522, N847);
not NOT1 (N3687, N3684);
and AND2 (N3688, N3676, N1471);
and AND4 (N3689, N3672, N2929, N1888, N925);
nor NOR4 (N3690, N3689, N794, N3269, N759);
or OR3 (N3691, N3687, N3057, N1955);
not NOT1 (N3692, N3691);
nor NOR2 (N3693, N3692, N1891);
nand NAND4 (N3694, N3683, N1043, N3538, N3095);
and AND2 (N3695, N3693, N1910);
xor XOR2 (N3696, N3694, N2346);
xor XOR2 (N3697, N3685, N302);
buf BUF1 (N3698, N3696);
not NOT1 (N3699, N3670);
and AND4 (N3700, N3698, N214, N2979, N2897);
nor NOR4 (N3701, N3695, N2013, N1977, N2075);
xor XOR2 (N3702, N3682, N2743);
not NOT1 (N3703, N3678);
nand NAND2 (N3704, N3703, N1094);
nand NAND3 (N3705, N3699, N983, N2088);
or OR4 (N3706, N3704, N2573, N505, N2742);
buf BUF1 (N3707, N3697);
or OR4 (N3708, N3686, N3121, N392, N104);
xor XOR2 (N3709, N3688, N3589);
nand NAND3 (N3710, N3690, N721, N1458);
buf BUF1 (N3711, N3709);
buf BUF1 (N3712, N3702);
not NOT1 (N3713, N3701);
and AND3 (N3714, N3711, N890, N219);
nor NOR4 (N3715, N3713, N2107, N580, N1856);
nor NOR3 (N3716, N3700, N267, N2101);
xor XOR2 (N3717, N3712, N348);
nand NAND2 (N3718, N3707, N1324);
buf BUF1 (N3719, N3716);
nand NAND4 (N3720, N3710, N1438, N2087, N3419);
not NOT1 (N3721, N3717);
and AND2 (N3722, N3708, N357);
nand NAND4 (N3723, N3705, N2821, N144, N2647);
xor XOR2 (N3724, N3706, N1009);
buf BUF1 (N3725, N3722);
nor NOR2 (N3726, N3718, N2795);
xor XOR2 (N3727, N3719, N1267);
nand NAND4 (N3728, N3723, N3059, N1096, N3720);
not NOT1 (N3729, N3531);
xor XOR2 (N3730, N3715, N2498);
nand NAND3 (N3731, N3729, N3308, N2185);
not NOT1 (N3732, N3721);
or OR2 (N3733, N3724, N3497);
or OR4 (N3734, N3732, N2080, N2902, N1661);
buf BUF1 (N3735, N3727);
and AND2 (N3736, N3714, N2904);
nand NAND4 (N3737, N3733, N2518, N2792, N501);
xor XOR2 (N3738, N3725, N2353);
nor NOR2 (N3739, N3681, N282);
buf BUF1 (N3740, N3737);
buf BUF1 (N3741, N3739);
and AND2 (N3742, N3730, N3723);
and AND2 (N3743, N3734, N2846);
and AND3 (N3744, N3741, N609, N401);
nand NAND4 (N3745, N3743, N1648, N3034, N3442);
not NOT1 (N3746, N3745);
not NOT1 (N3747, N3744);
not NOT1 (N3748, N3740);
xor XOR2 (N3749, N3728, N3410);
buf BUF1 (N3750, N3748);
nor NOR2 (N3751, N3749, N2777);
not NOT1 (N3752, N3742);
or OR4 (N3753, N3735, N3214, N1763, N1822);
and AND3 (N3754, N3726, N3149, N547);
nand NAND2 (N3755, N3750, N3286);
xor XOR2 (N3756, N3754, N3219);
not NOT1 (N3757, N3751);
or OR4 (N3758, N3731, N126, N2702, N960);
not NOT1 (N3759, N3738);
or OR4 (N3760, N3753, N148, N142, N1313);
buf BUF1 (N3761, N3759);
xor XOR2 (N3762, N3747, N1003);
nor NOR2 (N3763, N3746, N1632);
nand NAND2 (N3764, N3762, N1232);
xor XOR2 (N3765, N3756, N2961);
nor NOR2 (N3766, N3763, N2643);
not NOT1 (N3767, N3757);
nand NAND2 (N3768, N3752, N1984);
buf BUF1 (N3769, N3765);
or OR4 (N3770, N3755, N2151, N281, N677);
or OR4 (N3771, N3767, N953, N1658, N2387);
buf BUF1 (N3772, N3760);
buf BUF1 (N3773, N3769);
nor NOR3 (N3774, N3761, N3308, N2968);
xor XOR2 (N3775, N3772, N1299);
xor XOR2 (N3776, N3770, N2973);
buf BUF1 (N3777, N3764);
nor NOR3 (N3778, N3777, N1053, N2444);
not NOT1 (N3779, N3776);
nand NAND2 (N3780, N3766, N3715);
buf BUF1 (N3781, N3780);
buf BUF1 (N3782, N3768);
buf BUF1 (N3783, N3771);
buf BUF1 (N3784, N3779);
nand NAND4 (N3785, N3774, N139, N726, N3617);
not NOT1 (N3786, N3781);
not NOT1 (N3787, N3783);
not NOT1 (N3788, N3787);
and AND4 (N3789, N3782, N3148, N1293, N3609);
or OR3 (N3790, N3785, N295, N178);
and AND4 (N3791, N3789, N572, N3589, N1039);
and AND2 (N3792, N3790, N254);
not NOT1 (N3793, N3773);
and AND2 (N3794, N3784, N1807);
or OR2 (N3795, N3794, N573);
buf BUF1 (N3796, N3786);
xor XOR2 (N3797, N3792, N3211);
and AND4 (N3798, N3797, N1066, N3525, N2623);
or OR3 (N3799, N3788, N1669, N1287);
nor NOR2 (N3800, N3791, N2465);
nand NAND3 (N3801, N3793, N2733, N2298);
xor XOR2 (N3802, N3736, N2072);
nor NOR4 (N3803, N3795, N2557, N133, N1531);
buf BUF1 (N3804, N3801);
nor NOR2 (N3805, N3758, N3614);
nor NOR2 (N3806, N3778, N444);
buf BUF1 (N3807, N3802);
not NOT1 (N3808, N3796);
or OR2 (N3809, N3799, N3045);
buf BUF1 (N3810, N3809);
buf BUF1 (N3811, N3803);
or OR3 (N3812, N3806, N1654, N2087);
not NOT1 (N3813, N3798);
not NOT1 (N3814, N3810);
and AND2 (N3815, N3808, N1312);
nand NAND2 (N3816, N3813, N3588);
nor NOR3 (N3817, N3775, N847, N3373);
not NOT1 (N3818, N3800);
nand NAND2 (N3819, N3804, N54);
buf BUF1 (N3820, N3816);
xor XOR2 (N3821, N3807, N1729);
xor XOR2 (N3822, N3821, N684);
nor NOR2 (N3823, N3819, N1582);
xor XOR2 (N3824, N3812, N428);
not NOT1 (N3825, N3805);
nand NAND4 (N3826, N3815, N1631, N2271, N664);
nand NAND3 (N3827, N3822, N3770, N1688);
or OR2 (N3828, N3826, N3323);
nor NOR4 (N3829, N3823, N2571, N454, N1575);
and AND3 (N3830, N3818, N3457, N523);
not NOT1 (N3831, N3814);
nor NOR2 (N3832, N3830, N3427);
nor NOR4 (N3833, N3824, N255, N428, N1935);
and AND4 (N3834, N3832, N508, N2083, N2715);
and AND2 (N3835, N3829, N2564);
buf BUF1 (N3836, N3835);
not NOT1 (N3837, N3831);
buf BUF1 (N3838, N3828);
not NOT1 (N3839, N3825);
not NOT1 (N3840, N3836);
and AND4 (N3841, N3811, N1941, N1279, N3140);
and AND3 (N3842, N3827, N3564, N711);
nand NAND4 (N3843, N3842, N1906, N3530, N2993);
and AND4 (N3844, N3839, N2200, N1023, N42);
and AND2 (N3845, N3834, N1022);
or OR3 (N3846, N3817, N245, N2225);
nand NAND4 (N3847, N3837, N1360, N961, N1769);
not NOT1 (N3848, N3846);
nor NOR3 (N3849, N3833, N2987, N2585);
nor NOR3 (N3850, N3840, N3833, N1956);
xor XOR2 (N3851, N3847, N3131);
nor NOR2 (N3852, N3849, N2368);
or OR2 (N3853, N3843, N3442);
nor NOR4 (N3854, N3844, N3501, N1633, N3648);
nor NOR3 (N3855, N3853, N1619, N1647);
nor NOR2 (N3856, N3855, N3062);
buf BUF1 (N3857, N3841);
nand NAND2 (N3858, N3820, N3005);
buf BUF1 (N3859, N3845);
nor NOR4 (N3860, N3858, N2447, N3289, N2452);
xor XOR2 (N3861, N3851, N3673);
and AND4 (N3862, N3856, N234, N1068, N3125);
not NOT1 (N3863, N3854);
not NOT1 (N3864, N3848);
buf BUF1 (N3865, N3859);
xor XOR2 (N3866, N3863, N3130);
or OR3 (N3867, N3864, N1937, N1324);
not NOT1 (N3868, N3860);
not NOT1 (N3869, N3857);
nor NOR3 (N3870, N3865, N774, N3739);
xor XOR2 (N3871, N3850, N2178);
and AND3 (N3872, N3861, N217, N1155);
buf BUF1 (N3873, N3838);
or OR2 (N3874, N3862, N1702);
nor NOR2 (N3875, N3852, N1932);
xor XOR2 (N3876, N3874, N3300);
buf BUF1 (N3877, N3867);
nor NOR4 (N3878, N3868, N802, N3250, N1917);
not NOT1 (N3879, N3873);
nand NAND2 (N3880, N3875, N483);
buf BUF1 (N3881, N3872);
not NOT1 (N3882, N3881);
nand NAND2 (N3883, N3882, N2775);
buf BUF1 (N3884, N3883);
xor XOR2 (N3885, N3877, N3025);
not NOT1 (N3886, N3884);
buf BUF1 (N3887, N3871);
buf BUF1 (N3888, N3880);
and AND4 (N3889, N3878, N3637, N1029, N1670);
not NOT1 (N3890, N3866);
and AND2 (N3891, N3869, N2887);
or OR4 (N3892, N3887, N1163, N2824, N300);
or OR3 (N3893, N3890, N1258, N2018);
nand NAND2 (N3894, N3888, N3566);
nand NAND3 (N3895, N3886, N2459, N211);
buf BUF1 (N3896, N3891);
buf BUF1 (N3897, N3896);
nand NAND4 (N3898, N3897, N2680, N1308, N3768);
xor XOR2 (N3899, N3870, N2084);
xor XOR2 (N3900, N3885, N2708);
nor NOR4 (N3901, N3889, N1087, N2538, N2551);
buf BUF1 (N3902, N3879);
not NOT1 (N3903, N3902);
and AND3 (N3904, N3898, N2504, N1956);
or OR4 (N3905, N3901, N2352, N1570, N116);
buf BUF1 (N3906, N3899);
xor XOR2 (N3907, N3903, N2016);
buf BUF1 (N3908, N3895);
not NOT1 (N3909, N3892);
not NOT1 (N3910, N3907);
buf BUF1 (N3911, N3905);
xor XOR2 (N3912, N3900, N3863);
xor XOR2 (N3913, N3909, N1883);
buf BUF1 (N3914, N3913);
xor XOR2 (N3915, N3906, N3292);
nand NAND2 (N3916, N3911, N2065);
buf BUF1 (N3917, N3894);
xor XOR2 (N3918, N3908, N235);
and AND2 (N3919, N3893, N2783);
or OR2 (N3920, N3917, N2698);
nor NOR2 (N3921, N3912, N1339);
and AND4 (N3922, N3876, N2473, N1003, N3812);
nand NAND3 (N3923, N3919, N1763, N1209);
and AND3 (N3924, N3921, N2963, N402);
nand NAND3 (N3925, N3915, N1342, N1556);
or OR4 (N3926, N3914, N3637, N2557, N1502);
buf BUF1 (N3927, N3910);
and AND3 (N3928, N3916, N904, N2313);
and AND3 (N3929, N3904, N1924, N2991);
nand NAND4 (N3930, N3923, N3192, N2, N1354);
or OR3 (N3931, N3929, N1148, N3068);
nand NAND3 (N3932, N3924, N2203, N3763);
not NOT1 (N3933, N3918);
xor XOR2 (N3934, N3930, N2738);
xor XOR2 (N3935, N3933, N3003);
or OR4 (N3936, N3925, N3825, N3717, N1197);
buf BUF1 (N3937, N3935);
xor XOR2 (N3938, N3926, N1645);
and AND3 (N3939, N3931, N1776, N3198);
nand NAND4 (N3940, N3939, N2186, N1823, N2506);
and AND3 (N3941, N3940, N2936, N841);
nand NAND2 (N3942, N3922, N3505);
not NOT1 (N3943, N3937);
nor NOR2 (N3944, N3920, N52);
xor XOR2 (N3945, N3944, N3747);
not NOT1 (N3946, N3945);
xor XOR2 (N3947, N3928, N3680);
nand NAND2 (N3948, N3934, N3327);
and AND2 (N3949, N3943, N941);
buf BUF1 (N3950, N3941);
xor XOR2 (N3951, N3947, N1450);
nor NOR3 (N3952, N3932, N1301, N560);
nand NAND3 (N3953, N3949, N1751, N1075);
or OR2 (N3954, N3948, N1869);
xor XOR2 (N3955, N3946, N50);
and AND4 (N3956, N3951, N3675, N3240, N2367);
xor XOR2 (N3957, N3942, N1410);
and AND4 (N3958, N3954, N3082, N906, N2285);
xor XOR2 (N3959, N3958, N2147);
or OR4 (N3960, N3927, N3506, N1045, N1851);
nor NOR3 (N3961, N3938, N3100, N2394);
and AND3 (N3962, N3950, N3902, N694);
nand NAND4 (N3963, N3952, N2440, N2046, N2252);
or OR2 (N3964, N3960, N3662);
and AND2 (N3965, N3962, N261);
or OR2 (N3966, N3965, N2209);
buf BUF1 (N3967, N3955);
xor XOR2 (N3968, N3966, N3611);
buf BUF1 (N3969, N3968);
and AND4 (N3970, N3959, N3465, N1519, N3174);
buf BUF1 (N3971, N3956);
not NOT1 (N3972, N3971);
buf BUF1 (N3973, N3972);
buf BUF1 (N3974, N3969);
and AND4 (N3975, N3970, N3051, N3427, N3651);
or OR2 (N3976, N3957, N1661);
not NOT1 (N3977, N3961);
not NOT1 (N3978, N3974);
xor XOR2 (N3979, N3978, N268);
and AND4 (N3980, N3975, N3591, N2213, N892);
buf BUF1 (N3981, N3936);
buf BUF1 (N3982, N3979);
or OR4 (N3983, N3963, N871, N1238, N749);
not NOT1 (N3984, N3983);
not NOT1 (N3985, N3984);
nand NAND4 (N3986, N3973, N3469, N3600, N3186);
xor XOR2 (N3987, N3964, N1967);
xor XOR2 (N3988, N3986, N384);
xor XOR2 (N3989, N3987, N928);
or OR2 (N3990, N3980, N3771);
or OR4 (N3991, N3977, N2540, N1426, N1928);
or OR3 (N3992, N3976, N517, N2578);
xor XOR2 (N3993, N3989, N2578);
nand NAND4 (N3994, N3981, N1937, N2700, N3541);
and AND2 (N3995, N3953, N219);
nor NOR3 (N3996, N3992, N3945, N1698);
xor XOR2 (N3997, N3993, N1065);
and AND3 (N3998, N3988, N3476, N2574);
xor XOR2 (N3999, N3996, N2382);
nor NOR4 (N4000, N3982, N3377, N273, N2436);
and AND2 (N4001, N3998, N445);
nand NAND2 (N4002, N3997, N705);
nor NOR3 (N4003, N4002, N3203, N1576);
xor XOR2 (N4004, N3994, N3835);
and AND3 (N4005, N3967, N2493, N347);
xor XOR2 (N4006, N3990, N2790);
or OR2 (N4007, N4001, N3563);
or OR2 (N4008, N4004, N316);
or OR4 (N4009, N4003, N3509, N2189, N3888);
buf BUF1 (N4010, N3985);
or OR4 (N4011, N4009, N3728, N1013, N1661);
and AND3 (N4012, N4011, N1530, N1852);
xor XOR2 (N4013, N4006, N3953);
buf BUF1 (N4014, N3995);
nor NOR4 (N4015, N4010, N182, N2564, N1035);
nand NAND2 (N4016, N4005, N1657);
nor NOR3 (N4017, N4000, N2519, N205);
buf BUF1 (N4018, N4016);
nand NAND3 (N4019, N4014, N1068, N1407);
or OR2 (N4020, N4018, N1113);
and AND4 (N4021, N4012, N651, N367, N3799);
xor XOR2 (N4022, N3999, N3337);
buf BUF1 (N4023, N4020);
or OR3 (N4024, N4017, N1953, N2008);
not NOT1 (N4025, N3991);
and AND4 (N4026, N4008, N2073, N2885, N672);
not NOT1 (N4027, N4015);
xor XOR2 (N4028, N4025, N807);
and AND3 (N4029, N4023, N678, N1072);
or OR4 (N4030, N4027, N2682, N3884, N1838);
nand NAND3 (N4031, N4022, N1937, N1803);
not NOT1 (N4032, N4028);
or OR2 (N4033, N4013, N2912);
nor NOR4 (N4034, N4026, N3630, N3706, N1153);
nor NOR3 (N4035, N4024, N1342, N3850);
or OR4 (N4036, N4029, N2981, N217, N1003);
nand NAND2 (N4037, N4033, N327);
nand NAND4 (N4038, N4007, N1501, N2077, N3850);
buf BUF1 (N4039, N4019);
or OR4 (N4040, N4039, N564, N2619, N1485);
not NOT1 (N4041, N4037);
xor XOR2 (N4042, N4021, N3721);
not NOT1 (N4043, N4034);
xor XOR2 (N4044, N4031, N2808);
buf BUF1 (N4045, N4035);
buf BUF1 (N4046, N4042);
nand NAND4 (N4047, N4046, N2548, N3647, N3410);
nor NOR3 (N4048, N4043, N785, N351);
xor XOR2 (N4049, N4030, N2507);
and AND2 (N4050, N4044, N48);
xor XOR2 (N4051, N4032, N1024);
nand NAND2 (N4052, N4040, N3799);
buf BUF1 (N4053, N4047);
nand NAND2 (N4054, N4051, N4042);
or OR4 (N4055, N4054, N1080, N317, N1021);
nand NAND3 (N4056, N4041, N2915, N123);
buf BUF1 (N4057, N4048);
not NOT1 (N4058, N4045);
nand NAND4 (N4059, N4056, N1354, N1941, N1622);
nor NOR4 (N4060, N4036, N3839, N1569, N880);
not NOT1 (N4061, N4057);
buf BUF1 (N4062, N4055);
nand NAND4 (N4063, N4061, N169, N1315, N3652);
nand NAND2 (N4064, N4063, N428);
buf BUF1 (N4065, N4062);
buf BUF1 (N4066, N4052);
nor NOR4 (N4067, N4049, N276, N1665, N2097);
nor NOR3 (N4068, N4059, N2804, N1101);
or OR3 (N4069, N4065, N3825, N489);
nor NOR4 (N4070, N4068, N835, N3925, N3031);
buf BUF1 (N4071, N4064);
or OR2 (N4072, N4053, N2491);
xor XOR2 (N4073, N4072, N4);
and AND4 (N4074, N4069, N1559, N1315, N1898);
nor NOR4 (N4075, N4067, N3345, N2898, N3890);
buf BUF1 (N4076, N4074);
and AND4 (N4077, N4076, N10, N1297, N1246);
xor XOR2 (N4078, N4050, N3937);
xor XOR2 (N4079, N4066, N1765);
not NOT1 (N4080, N4038);
xor XOR2 (N4081, N4075, N2942);
buf BUF1 (N4082, N4079);
nor NOR2 (N4083, N4080, N1158);
nor NOR3 (N4084, N4078, N166, N2606);
buf BUF1 (N4085, N4058);
nor NOR4 (N4086, N4083, N722, N3364, N1282);
not NOT1 (N4087, N4086);
or OR4 (N4088, N4087, N108, N2320, N982);
xor XOR2 (N4089, N4088, N3209);
buf BUF1 (N4090, N4085);
nor NOR3 (N4091, N4071, N1125, N1154);
or OR4 (N4092, N4089, N1902, N3570, N360);
or OR2 (N4093, N4081, N3518);
buf BUF1 (N4094, N4093);
xor XOR2 (N4095, N4070, N3946);
xor XOR2 (N4096, N4090, N1658);
nand NAND4 (N4097, N4060, N2586, N548, N1796);
nand NAND2 (N4098, N4082, N138);
nand NAND2 (N4099, N4084, N23);
and AND2 (N4100, N4097, N2733);
buf BUF1 (N4101, N4077);
xor XOR2 (N4102, N4099, N3982);
buf BUF1 (N4103, N4101);
nand NAND3 (N4104, N4098, N438, N4057);
buf BUF1 (N4105, N4104);
not NOT1 (N4106, N4094);
and AND4 (N4107, N4073, N3778, N3850, N1970);
nand NAND2 (N4108, N4092, N2632);
not NOT1 (N4109, N4106);
buf BUF1 (N4110, N4091);
xor XOR2 (N4111, N4110, N358);
and AND2 (N4112, N4109, N2421);
nor NOR4 (N4113, N4105, N626, N1298, N367);
nand NAND4 (N4114, N4107, N2615, N3640, N1802);
nand NAND3 (N4115, N4113, N3537, N2016);
buf BUF1 (N4116, N4108);
nor NOR3 (N4117, N4114, N1318, N3771);
nand NAND2 (N4118, N4096, N283);
buf BUF1 (N4119, N4103);
and AND3 (N4120, N4118, N971, N9);
xor XOR2 (N4121, N4111, N2428);
not NOT1 (N4122, N4112);
buf BUF1 (N4123, N4122);
nand NAND2 (N4124, N4121, N2388);
or OR2 (N4125, N4123, N2317);
nor NOR4 (N4126, N4115, N2927, N3059, N3455);
xor XOR2 (N4127, N4126, N740);
or OR3 (N4128, N4124, N1740, N1099);
xor XOR2 (N4129, N4127, N201);
nand NAND4 (N4130, N4102, N460, N3966, N2280);
buf BUF1 (N4131, N4130);
and AND4 (N4132, N4131, N2851, N2797, N680);
and AND3 (N4133, N4129, N1701, N4048);
or OR2 (N4134, N4128, N1302);
nand NAND2 (N4135, N4117, N4105);
not NOT1 (N4136, N4095);
xor XOR2 (N4137, N4116, N1374);
buf BUF1 (N4138, N4119);
and AND2 (N4139, N4134, N3890);
nand NAND2 (N4140, N4132, N583);
nor NOR4 (N4141, N4139, N936, N2328, N2823);
nor NOR2 (N4142, N4135, N3303);
nor NOR3 (N4143, N4120, N2788, N3435);
nand NAND3 (N4144, N4100, N219, N3539);
or OR2 (N4145, N4137, N905);
or OR3 (N4146, N4142, N2632, N95);
buf BUF1 (N4147, N4125);
buf BUF1 (N4148, N4147);
nand NAND3 (N4149, N4140, N3235, N2192);
and AND4 (N4150, N4149, N3420, N3868, N330);
or OR4 (N4151, N4150, N2586, N298, N1638);
nor NOR3 (N4152, N4151, N2267, N538);
nand NAND3 (N4153, N4144, N2497, N2471);
xor XOR2 (N4154, N4138, N2759);
nor NOR3 (N4155, N4154, N393, N2650);
xor XOR2 (N4156, N4153, N1350);
or OR2 (N4157, N4143, N3078);
nor NOR4 (N4158, N4148, N1195, N1369, N985);
or OR2 (N4159, N4158, N283);
nor NOR2 (N4160, N4155, N581);
nand NAND2 (N4161, N4152, N2956);
nor NOR3 (N4162, N4160, N306, N2623);
nor NOR4 (N4163, N4159, N3318, N159, N2779);
and AND3 (N4164, N4145, N80, N237);
or OR3 (N4165, N4136, N4031, N534);
and AND3 (N4166, N4156, N971, N2601);
nand NAND4 (N4167, N4133, N2214, N3673, N1627);
nand NAND4 (N4168, N4165, N2184, N1216, N2552);
not NOT1 (N4169, N4161);
xor XOR2 (N4170, N4141, N409);
not NOT1 (N4171, N4157);
xor XOR2 (N4172, N4164, N432);
or OR4 (N4173, N4171, N4015, N2057, N3958);
xor XOR2 (N4174, N4162, N1119);
xor XOR2 (N4175, N4169, N2367);
not NOT1 (N4176, N4163);
and AND4 (N4177, N4174, N3546, N2949, N3267);
or OR2 (N4178, N4176, N1331);
or OR4 (N4179, N4146, N4040, N466, N202);
buf BUF1 (N4180, N4177);
nor NOR2 (N4181, N4168, N204);
nor NOR4 (N4182, N4172, N4075, N1281, N94);
buf BUF1 (N4183, N4173);
nand NAND2 (N4184, N4167, N850);
nor NOR2 (N4185, N4166, N1723);
not NOT1 (N4186, N4183);
and AND3 (N4187, N4180, N1906, N2000);
or OR4 (N4188, N4175, N3817, N2072, N997);
buf BUF1 (N4189, N4184);
and AND4 (N4190, N4188, N1263, N2054, N208);
buf BUF1 (N4191, N4179);
buf BUF1 (N4192, N4191);
not NOT1 (N4193, N4182);
or OR2 (N4194, N4181, N3478);
or OR3 (N4195, N4192, N30, N1078);
xor XOR2 (N4196, N4189, N2466);
or OR4 (N4197, N4186, N348, N1685, N2192);
nand NAND2 (N4198, N4196, N3444);
nand NAND3 (N4199, N4178, N4096, N3258);
xor XOR2 (N4200, N4194, N3822);
nand NAND2 (N4201, N4170, N952);
and AND4 (N4202, N4187, N943, N4065, N1965);
or OR3 (N4203, N4201, N1860, N1862);
or OR4 (N4204, N4190, N3434, N2996, N816);
nand NAND2 (N4205, N4185, N2891);
buf BUF1 (N4206, N4200);
not NOT1 (N4207, N4197);
nand NAND3 (N4208, N4198, N2737, N3204);
xor XOR2 (N4209, N4206, N2792);
nand NAND2 (N4210, N4208, N2568);
buf BUF1 (N4211, N4199);
not NOT1 (N4212, N4204);
nand NAND4 (N4213, N4210, N365, N3616, N2330);
buf BUF1 (N4214, N4202);
buf BUF1 (N4215, N4209);
or OR2 (N4216, N4212, N2807);
nor NOR4 (N4217, N4216, N95, N2026, N963);
buf BUF1 (N4218, N4213);
not NOT1 (N4219, N4203);
xor XOR2 (N4220, N4215, N1750);
nor NOR2 (N4221, N4195, N585);
or OR2 (N4222, N4193, N1552);
and AND2 (N4223, N4211, N1666);
and AND2 (N4224, N4223, N3708);
xor XOR2 (N4225, N4217, N3526);
or OR2 (N4226, N4225, N3785);
nor NOR2 (N4227, N4220, N1107);
nor NOR3 (N4228, N4218, N1011, N3571);
or OR3 (N4229, N4219, N2611, N577);
buf BUF1 (N4230, N4224);
or OR2 (N4231, N4207, N4207);
xor XOR2 (N4232, N4221, N3333);
nand NAND3 (N4233, N4226, N50, N3145);
xor XOR2 (N4234, N4205, N2492);
xor XOR2 (N4235, N4229, N2306);
not NOT1 (N4236, N4214);
nand NAND4 (N4237, N4233, N4209, N2112, N2017);
xor XOR2 (N4238, N4230, N1455);
or OR2 (N4239, N4227, N1770);
buf BUF1 (N4240, N4232);
or OR3 (N4241, N4240, N3839, N1459);
buf BUF1 (N4242, N4222);
nor NOR3 (N4243, N4231, N1006, N204);
xor XOR2 (N4244, N4236, N2791);
xor XOR2 (N4245, N4237, N920);
nor NOR2 (N4246, N4241, N2694);
nor NOR2 (N4247, N4234, N3404);
nor NOR3 (N4248, N4242, N2710, N2932);
buf BUF1 (N4249, N4245);
not NOT1 (N4250, N4235);
and AND4 (N4251, N4228, N1171, N1040, N587);
nor NOR3 (N4252, N4238, N767, N697);
xor XOR2 (N4253, N4252, N2977);
not NOT1 (N4254, N4244);
nor NOR2 (N4255, N4247, N2020);
or OR4 (N4256, N4255, N1432, N1867, N76);
nand NAND3 (N4257, N4248, N75, N3176);
nor NOR4 (N4258, N4239, N2176, N800, N2047);
xor XOR2 (N4259, N4258, N2139);
nand NAND3 (N4260, N4257, N966, N3358);
buf BUF1 (N4261, N4253);
or OR2 (N4262, N4254, N42);
not NOT1 (N4263, N4256);
not NOT1 (N4264, N4261);
nand NAND3 (N4265, N4262, N753, N3969);
nor NOR3 (N4266, N4243, N3950, N186);
nor NOR2 (N4267, N4251, N3378);
xor XOR2 (N4268, N4265, N818);
nor NOR4 (N4269, N4264, N3512, N3700, N228);
and AND3 (N4270, N4250, N509, N3349);
not NOT1 (N4271, N4246);
nand NAND2 (N4272, N4266, N4093);
and AND4 (N4273, N4260, N2688, N2807, N2723);
and AND4 (N4274, N4271, N826, N2957, N2079);
and AND2 (N4275, N4267, N3934);
not NOT1 (N4276, N4272);
not NOT1 (N4277, N4259);
nand NAND2 (N4278, N4263, N2847);
nor NOR4 (N4279, N4277, N777, N253, N1873);
buf BUF1 (N4280, N4276);
nand NAND2 (N4281, N4268, N1557);
not NOT1 (N4282, N4274);
nor NOR3 (N4283, N4249, N2079, N2554);
buf BUF1 (N4284, N4273);
and AND3 (N4285, N4275, N1198, N2529);
nand NAND2 (N4286, N4282, N608);
buf BUF1 (N4287, N4270);
or OR3 (N4288, N4283, N1973, N3744);
and AND2 (N4289, N4269, N1057);
nor NOR4 (N4290, N4289, N3785, N3425, N2378);
nor NOR3 (N4291, N4284, N4173, N1391);
not NOT1 (N4292, N4286);
not NOT1 (N4293, N4285);
buf BUF1 (N4294, N4281);
nand NAND3 (N4295, N4288, N3871, N1477);
nand NAND4 (N4296, N4294, N1704, N2925, N3990);
nand NAND2 (N4297, N4293, N4011);
and AND4 (N4298, N4297, N2557, N3341, N1096);
xor XOR2 (N4299, N4292, N789);
nand NAND2 (N4300, N4298, N2468);
nand NAND3 (N4301, N4280, N441, N269);
not NOT1 (N4302, N4279);
or OR2 (N4303, N4300, N1203);
or OR2 (N4304, N4291, N748);
buf BUF1 (N4305, N4303);
nor NOR2 (N4306, N4296, N2750);
buf BUF1 (N4307, N4278);
not NOT1 (N4308, N4301);
not NOT1 (N4309, N4307);
xor XOR2 (N4310, N4304, N2300);
not NOT1 (N4311, N4309);
nand NAND3 (N4312, N4295, N1926, N3626);
or OR2 (N4313, N4310, N3443);
nor NOR3 (N4314, N4287, N2270, N1350);
buf BUF1 (N4315, N4311);
xor XOR2 (N4316, N4306, N1902);
or OR2 (N4317, N4313, N3589);
not NOT1 (N4318, N4314);
nand NAND3 (N4319, N4299, N132, N4290);
and AND4 (N4320, N1368, N1702, N3631, N465);
nand NAND4 (N4321, N4305, N2854, N3198, N1918);
not NOT1 (N4322, N4316);
not NOT1 (N4323, N4321);
nor NOR4 (N4324, N4308, N2739, N2604, N2724);
buf BUF1 (N4325, N4302);
xor XOR2 (N4326, N4318, N142);
not NOT1 (N4327, N4326);
or OR2 (N4328, N4319, N1601);
nor NOR2 (N4329, N4320, N3249);
nor NOR3 (N4330, N4312, N572, N884);
and AND3 (N4331, N4315, N1426, N2419);
nor NOR2 (N4332, N4325, N2014);
buf BUF1 (N4333, N4329);
xor XOR2 (N4334, N4327, N625);
and AND4 (N4335, N4331, N4254, N3669, N3517);
nor NOR2 (N4336, N4317, N2144);
nor NOR3 (N4337, N4332, N3558, N1280);
xor XOR2 (N4338, N4336, N4093);
and AND4 (N4339, N4338, N2934, N2045, N2988);
and AND2 (N4340, N4323, N3288);
and AND3 (N4341, N4330, N3534, N1181);
and AND2 (N4342, N4334, N1611);
or OR2 (N4343, N4340, N679);
not NOT1 (N4344, N4339);
not NOT1 (N4345, N4322);
nand NAND2 (N4346, N4337, N1490);
xor XOR2 (N4347, N4333, N2604);
and AND2 (N4348, N4345, N4058);
and AND4 (N4349, N4324, N1850, N3513, N1179);
not NOT1 (N4350, N4335);
and AND3 (N4351, N4348, N139, N3803);
or OR2 (N4352, N4346, N1667);
and AND2 (N4353, N4343, N213);
or OR3 (N4354, N4350, N2183, N2261);
or OR2 (N4355, N4349, N1665);
xor XOR2 (N4356, N4347, N3842);
not NOT1 (N4357, N4354);
nand NAND4 (N4358, N4355, N273, N207, N4343);
or OR3 (N4359, N4358, N2214, N3967);
buf BUF1 (N4360, N4351);
xor XOR2 (N4361, N4360, N613);
or OR2 (N4362, N4352, N2375);
buf BUF1 (N4363, N4328);
not NOT1 (N4364, N4353);
not NOT1 (N4365, N4356);
not NOT1 (N4366, N4342);
buf BUF1 (N4367, N4341);
buf BUF1 (N4368, N4367);
xor XOR2 (N4369, N4363, N1322);
nand NAND4 (N4370, N4365, N3562, N1214, N3639);
nand NAND2 (N4371, N4362, N2544);
nand NAND4 (N4372, N4371, N1585, N4143, N1310);
nor NOR3 (N4373, N4368, N2006, N590);
nand NAND2 (N4374, N4372, N909);
and AND4 (N4375, N4359, N2651, N3406, N2267);
nand NAND2 (N4376, N4344, N1817);
not NOT1 (N4377, N4369);
and AND4 (N4378, N4361, N723, N3218, N3350);
xor XOR2 (N4379, N4366, N2613);
xor XOR2 (N4380, N4379, N3677);
xor XOR2 (N4381, N4373, N1502);
or OR4 (N4382, N4374, N3859, N1171, N82);
and AND4 (N4383, N4380, N2935, N628, N230);
nor NOR2 (N4384, N4357, N3687);
buf BUF1 (N4385, N4375);
or OR2 (N4386, N4385, N1569);
not NOT1 (N4387, N4377);
or OR4 (N4388, N4384, N1738, N2752, N343);
nor NOR3 (N4389, N4370, N164, N2014);
xor XOR2 (N4390, N4382, N3659);
not NOT1 (N4391, N4388);
not NOT1 (N4392, N4389);
buf BUF1 (N4393, N4383);
xor XOR2 (N4394, N4387, N2363);
not NOT1 (N4395, N4376);
nor NOR3 (N4396, N4392, N3735, N2374);
nand NAND2 (N4397, N4391, N3478);
buf BUF1 (N4398, N4364);
and AND2 (N4399, N4393, N3118);
buf BUF1 (N4400, N4386);
buf BUF1 (N4401, N4378);
and AND2 (N4402, N4381, N4133);
or OR3 (N4403, N4400, N3266, N1667);
buf BUF1 (N4404, N4394);
nor NOR2 (N4405, N4395, N4313);
buf BUF1 (N4406, N4402);
nor NOR4 (N4407, N4401, N2156, N3005, N3108);
not NOT1 (N4408, N4390);
buf BUF1 (N4409, N4399);
xor XOR2 (N4410, N4405, N549);
nand NAND3 (N4411, N4409, N838, N1171);
nor NOR3 (N4412, N4407, N4263, N2849);
nor NOR2 (N4413, N4411, N237);
nand NAND3 (N4414, N4406, N1423, N2354);
nand NAND3 (N4415, N4398, N485, N3147);
xor XOR2 (N4416, N4403, N1693);
or OR2 (N4417, N4414, N841);
and AND3 (N4418, N4404, N3819, N3782);
and AND4 (N4419, N4412, N2, N1482, N3274);
nand NAND3 (N4420, N4415, N2185, N1917);
or OR4 (N4421, N4416, N2129, N2293, N2913);
nand NAND2 (N4422, N4408, N1360);
not NOT1 (N4423, N4410);
xor XOR2 (N4424, N4420, N2502);
buf BUF1 (N4425, N4424);
buf BUF1 (N4426, N4419);
xor XOR2 (N4427, N4426, N1841);
xor XOR2 (N4428, N4397, N976);
and AND2 (N4429, N4396, N3727);
nor NOR3 (N4430, N4422, N1362, N823);
buf BUF1 (N4431, N4423);
nor NOR3 (N4432, N4413, N115, N651);
buf BUF1 (N4433, N4428);
nand NAND2 (N4434, N4427, N2495);
nand NAND3 (N4435, N4417, N3388, N2661);
xor XOR2 (N4436, N4418, N1638);
or OR3 (N4437, N4421, N1532, N3931);
buf BUF1 (N4438, N4437);
xor XOR2 (N4439, N4431, N307);
not NOT1 (N4440, N4435);
xor XOR2 (N4441, N4438, N2679);
nand NAND3 (N4442, N4432, N1642, N2529);
nand NAND2 (N4443, N4433, N474);
and AND3 (N4444, N4436, N1266, N2531);
and AND4 (N4445, N4430, N2682, N2254, N473);
nand NAND4 (N4446, N4425, N1232, N919, N1197);
buf BUF1 (N4447, N4439);
or OR3 (N4448, N4443, N709, N1857);
nor NOR4 (N4449, N4448, N1424, N61, N364);
not NOT1 (N4450, N4429);
nor NOR3 (N4451, N4450, N1317, N913);
and AND3 (N4452, N4440, N3189, N3692);
not NOT1 (N4453, N4452);
or OR4 (N4454, N4445, N1241, N2050, N4350);
nand NAND3 (N4455, N4444, N292, N3376);
and AND4 (N4456, N4434, N885, N1199, N1813);
and AND3 (N4457, N4455, N3380, N3710);
and AND4 (N4458, N4442, N2145, N2714, N715);
xor XOR2 (N4459, N4449, N3018);
buf BUF1 (N4460, N4446);
or OR3 (N4461, N4460, N3603, N3224);
xor XOR2 (N4462, N4451, N391);
nor NOR3 (N4463, N4458, N3294, N263);
or OR3 (N4464, N4461, N4237, N1209);
nor NOR2 (N4465, N4462, N1338);
nand NAND2 (N4466, N4454, N31);
not NOT1 (N4467, N4463);
or OR4 (N4468, N4457, N1786, N1893, N316);
nand NAND4 (N4469, N4459, N3870, N927, N1839);
and AND4 (N4470, N4469, N1605, N3881, N1314);
not NOT1 (N4471, N4468);
nand NAND2 (N4472, N4456, N3308);
and AND2 (N4473, N4453, N316);
xor XOR2 (N4474, N4464, N2090);
nand NAND3 (N4475, N4465, N1389, N1893);
xor XOR2 (N4476, N4470, N2355);
nor NOR4 (N4477, N4475, N1157, N4170, N2432);
nor NOR3 (N4478, N4441, N1999, N4436);
or OR4 (N4479, N4472, N603, N785, N3693);
buf BUF1 (N4480, N4467);
nor NOR4 (N4481, N4466, N2391, N2944, N41);
nand NAND3 (N4482, N4476, N3234, N1867);
nand NAND2 (N4483, N4477, N4306);
not NOT1 (N4484, N4474);
nor NOR2 (N4485, N4447, N2966);
or OR2 (N4486, N4471, N335);
nand NAND2 (N4487, N4478, N3808);
and AND4 (N4488, N4485, N4017, N1773, N1991);
nor NOR4 (N4489, N4484, N2756, N2831, N1359);
nor NOR4 (N4490, N4473, N2170, N4158, N661);
buf BUF1 (N4491, N4479);
not NOT1 (N4492, N4490);
or OR4 (N4493, N4488, N464, N429, N2451);
not NOT1 (N4494, N4493);
buf BUF1 (N4495, N4486);
not NOT1 (N4496, N4483);
nor NOR3 (N4497, N4487, N2550, N4005);
nor NOR3 (N4498, N4495, N1612, N2100);
buf BUF1 (N4499, N4489);
and AND2 (N4500, N4492, N1307);
xor XOR2 (N4501, N4491, N610);
nor NOR4 (N4502, N4482, N861, N2002, N4068);
not NOT1 (N4503, N4496);
buf BUF1 (N4504, N4498);
and AND4 (N4505, N4502, N28, N2386, N1449);
buf BUF1 (N4506, N4494);
nor NOR4 (N4507, N4500, N1939, N3016, N633);
nand NAND4 (N4508, N4506, N1570, N1463, N2660);
and AND4 (N4509, N4497, N1089, N3465, N1535);
nor NOR4 (N4510, N4507, N923, N1242, N2723);
buf BUF1 (N4511, N4510);
buf BUF1 (N4512, N4509);
xor XOR2 (N4513, N4512, N2982);
or OR2 (N4514, N4513, N2238);
xor XOR2 (N4515, N4511, N1818);
nor NOR2 (N4516, N4480, N4271);
buf BUF1 (N4517, N4503);
not NOT1 (N4518, N4508);
nor NOR4 (N4519, N4504, N116, N1539, N3005);
nor NOR3 (N4520, N4519, N3352, N3099);
nand NAND3 (N4521, N4514, N1034, N3513);
and AND3 (N4522, N4501, N2888, N776);
not NOT1 (N4523, N4499);
and AND3 (N4524, N4520, N1079, N917);
not NOT1 (N4525, N4517);
xor XOR2 (N4526, N4481, N4000);
nand NAND2 (N4527, N4505, N2331);
xor XOR2 (N4528, N4527, N179);
not NOT1 (N4529, N4524);
nor NOR2 (N4530, N4525, N541);
nand NAND3 (N4531, N4515, N776, N145);
or OR3 (N4532, N4516, N1528, N1502);
xor XOR2 (N4533, N4530, N532);
or OR3 (N4534, N4521, N2415, N1216);
nand NAND4 (N4535, N4526, N1394, N2447, N1069);
and AND4 (N4536, N4518, N2535, N942, N1299);
nand NAND3 (N4537, N4536, N1269, N1821);
buf BUF1 (N4538, N4537);
and AND2 (N4539, N4531, N857);
and AND2 (N4540, N4522, N2114);
nand NAND3 (N4541, N4540, N2169, N2390);
and AND3 (N4542, N4534, N818, N3918);
or OR3 (N4543, N4541, N384, N4071);
nand NAND3 (N4544, N4533, N97, N3620);
nor NOR3 (N4545, N4528, N182, N2816);
and AND3 (N4546, N4523, N3492, N3282);
or OR2 (N4547, N4542, N1611);
and AND2 (N4548, N4546, N2265);
xor XOR2 (N4549, N4548, N3924);
buf BUF1 (N4550, N4529);
not NOT1 (N4551, N4549);
nand NAND3 (N4552, N4532, N4531, N786);
xor XOR2 (N4553, N4547, N2805);
and AND4 (N4554, N4551, N1629, N4477, N3480);
not NOT1 (N4555, N4544);
buf BUF1 (N4556, N4543);
buf BUF1 (N4557, N4545);
not NOT1 (N4558, N4553);
nor NOR2 (N4559, N4558, N3360);
xor XOR2 (N4560, N4554, N3133);
not NOT1 (N4561, N4550);
nor NOR3 (N4562, N4556, N3659, N663);
buf BUF1 (N4563, N4560);
nand NAND3 (N4564, N4535, N1291, N1667);
buf BUF1 (N4565, N4561);
xor XOR2 (N4566, N4562, N3953);
nand NAND2 (N4567, N4565, N3993);
buf BUF1 (N4568, N4552);
xor XOR2 (N4569, N4568, N113);
buf BUF1 (N4570, N4538);
or OR2 (N4571, N4563, N963);
and AND4 (N4572, N4557, N1799, N4457, N1231);
nor NOR4 (N4573, N4566, N2416, N1482, N3165);
nor NOR4 (N4574, N4571, N1667, N4385, N3917);
nor NOR3 (N4575, N4569, N193, N3786);
nand NAND2 (N4576, N4567, N2584);
and AND4 (N4577, N4576, N3506, N1144, N1658);
nor NOR4 (N4578, N4555, N1324, N4551, N1509);
not NOT1 (N4579, N4564);
not NOT1 (N4580, N4570);
xor XOR2 (N4581, N4578, N2398);
nor NOR3 (N4582, N4579, N828, N1015);
and AND3 (N4583, N4574, N2277, N2974);
xor XOR2 (N4584, N4580, N3652);
buf BUF1 (N4585, N4583);
and AND4 (N4586, N4585, N221, N2901, N4441);
nor NOR4 (N4587, N4573, N2772, N2456, N2895);
or OR4 (N4588, N4539, N3526, N103, N2793);
not NOT1 (N4589, N4587);
not NOT1 (N4590, N4588);
buf BUF1 (N4591, N4581);
xor XOR2 (N4592, N4572, N4296);
xor XOR2 (N4593, N4559, N1082);
nor NOR3 (N4594, N4586, N2645, N160);
xor XOR2 (N4595, N4590, N4500);
or OR4 (N4596, N4592, N3028, N2299, N3675);
not NOT1 (N4597, N4589);
buf BUF1 (N4598, N4596);
nor NOR2 (N4599, N4598, N4478);
nor NOR2 (N4600, N4594, N4469);
and AND4 (N4601, N4582, N2865, N214, N362);
and AND4 (N4602, N4599, N1568, N4570, N2612);
or OR3 (N4603, N4575, N4428, N921);
xor XOR2 (N4604, N4577, N2797);
or OR2 (N4605, N4593, N210);
nand NAND3 (N4606, N4591, N3568, N4477);
buf BUF1 (N4607, N4584);
buf BUF1 (N4608, N4595);
or OR4 (N4609, N4602, N2055, N1002, N1774);
xor XOR2 (N4610, N4603, N4555);
or OR3 (N4611, N4609, N1799, N4021);
or OR3 (N4612, N4604, N1431, N175);
and AND2 (N4613, N4610, N2491);
and AND2 (N4614, N4601, N2992);
and AND3 (N4615, N4606, N7, N1330);
nor NOR2 (N4616, N4615, N1655);
or OR4 (N4617, N4600, N2300, N276, N3001);
and AND4 (N4618, N4608, N2548, N1872, N1467);
nor NOR3 (N4619, N4612, N3326, N2353);
xor XOR2 (N4620, N4618, N506);
not NOT1 (N4621, N4619);
not NOT1 (N4622, N4607);
or OR2 (N4623, N4617, N3120);
nand NAND2 (N4624, N4616, N2948);
or OR4 (N4625, N4624, N3276, N3892, N112);
nand NAND2 (N4626, N4622, N4390);
nor NOR3 (N4627, N4605, N3417, N209);
buf BUF1 (N4628, N4597);
or OR2 (N4629, N4620, N89);
nand NAND2 (N4630, N4623, N1747);
nor NOR2 (N4631, N4626, N3682);
and AND2 (N4632, N4629, N3172);
or OR4 (N4633, N4614, N4169, N2280, N3501);
xor XOR2 (N4634, N4630, N2170);
nand NAND4 (N4635, N4627, N1199, N1775, N4090);
nand NAND4 (N4636, N4628, N4214, N1586, N929);
and AND3 (N4637, N4634, N1061, N2257);
buf BUF1 (N4638, N4625);
xor XOR2 (N4639, N4632, N2610);
xor XOR2 (N4640, N4621, N4268);
not NOT1 (N4641, N4640);
nand NAND3 (N4642, N4613, N1760, N2062);
nand NAND2 (N4643, N4633, N2495);
buf BUF1 (N4644, N4631);
nor NOR4 (N4645, N4635, N3311, N507, N4510);
and AND4 (N4646, N4642, N135, N62, N919);
or OR2 (N4647, N4638, N180);
xor XOR2 (N4648, N4645, N4);
or OR4 (N4649, N4643, N2908, N3603, N1822);
and AND3 (N4650, N4636, N827, N1881);
nor NOR2 (N4651, N4649, N4408);
and AND4 (N4652, N4650, N816, N1585, N2626);
buf BUF1 (N4653, N4652);
and AND4 (N4654, N4611, N3959, N1209, N1578);
nand NAND4 (N4655, N4653, N862, N3184, N1093);
or OR2 (N4656, N4654, N4105);
nor NOR4 (N4657, N4641, N2058, N2381, N1337);
and AND4 (N4658, N4639, N1633, N4463, N36);
nor NOR3 (N4659, N4655, N58, N3913);
or OR2 (N4660, N4646, N3148);
xor XOR2 (N4661, N4656, N3524);
or OR2 (N4662, N4648, N1087);
not NOT1 (N4663, N4657);
nand NAND4 (N4664, N4647, N1109, N4308, N325);
nand NAND2 (N4665, N4664, N2752);
or OR2 (N4666, N4660, N2690);
nor NOR3 (N4667, N4662, N4320, N4311);
or OR4 (N4668, N4658, N247, N877, N4531);
xor XOR2 (N4669, N4644, N4587);
or OR4 (N4670, N4668, N4651, N3115, N1559);
nand NAND4 (N4671, N503, N1278, N854, N1475);
nand NAND2 (N4672, N4666, N4627);
xor XOR2 (N4673, N4661, N4624);
and AND2 (N4674, N4670, N3439);
xor XOR2 (N4675, N4659, N42);
not NOT1 (N4676, N4665);
nand NAND3 (N4677, N4676, N1859, N1678);
and AND2 (N4678, N4673, N872);
buf BUF1 (N4679, N4674);
buf BUF1 (N4680, N4671);
nor NOR4 (N4681, N4680, N2949, N4258, N184);
xor XOR2 (N4682, N4675, N4334);
and AND3 (N4683, N4667, N149, N3749);
nand NAND4 (N4684, N4663, N3838, N4182, N1592);
nor NOR3 (N4685, N4684, N1723, N49);
and AND4 (N4686, N4669, N2429, N382, N4404);
nor NOR4 (N4687, N4686, N2518, N1369, N881);
buf BUF1 (N4688, N4681);
or OR2 (N4689, N4677, N4535);
not NOT1 (N4690, N4672);
nor NOR3 (N4691, N4689, N1525, N1848);
not NOT1 (N4692, N4688);
not NOT1 (N4693, N4683);
nand NAND4 (N4694, N4690, N740, N2247, N48);
xor XOR2 (N4695, N4687, N2662);
nand NAND2 (N4696, N4678, N2956);
not NOT1 (N4697, N4693);
not NOT1 (N4698, N4679);
and AND4 (N4699, N4691, N3424, N3295, N2350);
nand NAND4 (N4700, N4699, N1730, N3374, N3837);
or OR2 (N4701, N4697, N1920);
or OR4 (N4702, N4637, N2352, N2390, N1893);
not NOT1 (N4703, N4701);
nand NAND2 (N4704, N4685, N694);
or OR4 (N4705, N4692, N3422, N3577, N2220);
buf BUF1 (N4706, N4696);
xor XOR2 (N4707, N4706, N4290);
and AND4 (N4708, N4698, N2794, N1483, N705);
not NOT1 (N4709, N4704);
or OR3 (N4710, N4700, N4528, N1840);
xor XOR2 (N4711, N4682, N1603);
buf BUF1 (N4712, N4710);
and AND3 (N4713, N4712, N357, N437);
buf BUF1 (N4714, N4695);
not NOT1 (N4715, N4702);
nor NOR2 (N4716, N4709, N3890);
not NOT1 (N4717, N4714);
not NOT1 (N4718, N4717);
or OR2 (N4719, N4708, N3392);
buf BUF1 (N4720, N4713);
not NOT1 (N4721, N4694);
and AND2 (N4722, N4711, N4397);
nor NOR4 (N4723, N4703, N2685, N2282, N1452);
buf BUF1 (N4724, N4715);
not NOT1 (N4725, N4716);
and AND2 (N4726, N4720, N4107);
and AND4 (N4727, N4723, N1974, N462, N887);
and AND3 (N4728, N4725, N600, N4558);
not NOT1 (N4729, N4728);
or OR3 (N4730, N4707, N1806, N2901);
buf BUF1 (N4731, N4727);
not NOT1 (N4732, N4724);
or OR3 (N4733, N4718, N3676, N3590);
nor NOR2 (N4734, N4729, N4032);
nand NAND2 (N4735, N4721, N3898);
or OR2 (N4736, N4731, N606);
xor XOR2 (N4737, N4735, N2837);
nor NOR3 (N4738, N4719, N2047, N3547);
nor NOR4 (N4739, N4732, N2150, N3763, N2414);
buf BUF1 (N4740, N4736);
and AND4 (N4741, N4739, N2258, N3999, N809);
nand NAND4 (N4742, N4734, N670, N3030, N8);
or OR3 (N4743, N4738, N4016, N3692);
buf BUF1 (N4744, N4726);
or OR4 (N4745, N4740, N1218, N687, N3634);
and AND2 (N4746, N4743, N2261);
nor NOR2 (N4747, N4730, N3980);
or OR3 (N4748, N4733, N3910, N283);
xor XOR2 (N4749, N4748, N3571);
not NOT1 (N4750, N4737);
xor XOR2 (N4751, N4750, N2993);
not NOT1 (N4752, N4746);
buf BUF1 (N4753, N4742);
nand NAND2 (N4754, N4753, N2728);
xor XOR2 (N4755, N4722, N1);
not NOT1 (N4756, N4752);
xor XOR2 (N4757, N4749, N2043);
xor XOR2 (N4758, N4755, N507);
xor XOR2 (N4759, N4745, N4295);
buf BUF1 (N4760, N4756);
buf BUF1 (N4761, N4760);
and AND4 (N4762, N4751, N4341, N1193, N2881);
or OR2 (N4763, N4744, N378);
or OR3 (N4764, N4705, N3234, N4351);
not NOT1 (N4765, N4762);
nor NOR3 (N4766, N4757, N3989, N12);
nand NAND2 (N4767, N4763, N2820);
and AND4 (N4768, N4741, N2732, N4449, N769);
nor NOR2 (N4769, N4768, N4149);
or OR3 (N4770, N4766, N1935, N292);
nor NOR4 (N4771, N4759, N418, N4033, N17);
not NOT1 (N4772, N4765);
not NOT1 (N4773, N4764);
not NOT1 (N4774, N4754);
nand NAND3 (N4775, N4758, N3015, N3468);
and AND2 (N4776, N4772, N2633);
buf BUF1 (N4777, N4771);
xor XOR2 (N4778, N4777, N2501);
nor NOR3 (N4779, N4761, N928, N4022);
and AND2 (N4780, N4769, N4131);
buf BUF1 (N4781, N4770);
buf BUF1 (N4782, N4767);
or OR2 (N4783, N4778, N2413);
nor NOR2 (N4784, N4775, N1093);
xor XOR2 (N4785, N4783, N2224);
nor NOR4 (N4786, N4784, N412, N2916, N1729);
buf BUF1 (N4787, N4782);
xor XOR2 (N4788, N4774, N1739);
not NOT1 (N4789, N4776);
nand NAND2 (N4790, N4747, N3626);
nand NAND3 (N4791, N4786, N4155, N4182);
xor XOR2 (N4792, N4790, N1364);
nand NAND4 (N4793, N4787, N3695, N1065, N1847);
or OR4 (N4794, N4781, N2717, N4694, N2702);
and AND4 (N4795, N4780, N688, N1375, N4743);
not NOT1 (N4796, N4794);
and AND4 (N4797, N4779, N2085, N882, N1588);
xor XOR2 (N4798, N4785, N3035);
xor XOR2 (N4799, N4793, N247);
xor XOR2 (N4800, N4797, N277);
or OR4 (N4801, N4791, N934, N8, N652);
or OR2 (N4802, N4799, N198);
nor NOR3 (N4803, N4800, N1288, N1490);
not NOT1 (N4804, N4795);
not NOT1 (N4805, N4802);
or OR3 (N4806, N4788, N1743, N1058);
and AND3 (N4807, N4792, N3938, N3539);
buf BUF1 (N4808, N4789);
xor XOR2 (N4809, N4803, N4737);
nand NAND3 (N4810, N4796, N1296, N4071);
and AND3 (N4811, N4806, N1286, N130);
nor NOR3 (N4812, N4773, N3855, N4211);
buf BUF1 (N4813, N4801);
not NOT1 (N4814, N4807);
not NOT1 (N4815, N4805);
buf BUF1 (N4816, N4813);
nand NAND3 (N4817, N4809, N1512, N3211);
nor NOR4 (N4818, N4814, N371, N2471, N1929);
and AND3 (N4819, N4811, N2936, N2318);
nor NOR3 (N4820, N4816, N2633, N4514);
nand NAND3 (N4821, N4810, N3626, N1667);
nand NAND2 (N4822, N4820, N2746);
or OR2 (N4823, N4818, N245);
nand NAND4 (N4824, N4822, N735, N4571, N1960);
buf BUF1 (N4825, N4823);
nor NOR4 (N4826, N4817, N3634, N29, N4199);
not NOT1 (N4827, N4815);
nor NOR3 (N4828, N4825, N2960, N4503);
xor XOR2 (N4829, N4828, N4578);
not NOT1 (N4830, N4827);
nand NAND4 (N4831, N4819, N754, N4062, N1388);
xor XOR2 (N4832, N4831, N1167);
nor NOR2 (N4833, N4824, N1203);
xor XOR2 (N4834, N4808, N240);
buf BUF1 (N4835, N4812);
not NOT1 (N4836, N4826);
or OR3 (N4837, N4830, N648, N1208);
buf BUF1 (N4838, N4821);
not NOT1 (N4839, N4837);
nand NAND2 (N4840, N4839, N1592);
buf BUF1 (N4841, N4836);
and AND4 (N4842, N4833, N3862, N2013, N144);
buf BUF1 (N4843, N4804);
nand NAND4 (N4844, N4832, N4201, N4095, N471);
nand NAND2 (N4845, N4840, N2799);
xor XOR2 (N4846, N4844, N2126);
buf BUF1 (N4847, N4843);
xor XOR2 (N4848, N4838, N46);
not NOT1 (N4849, N4798);
and AND3 (N4850, N4849, N616, N3622);
nor NOR3 (N4851, N4829, N962, N3040);
nor NOR3 (N4852, N4835, N4377, N4514);
xor XOR2 (N4853, N4850, N3659);
xor XOR2 (N4854, N4851, N2161);
nand NAND4 (N4855, N4848, N418, N3434, N2228);
nand NAND4 (N4856, N4845, N2295, N3574, N1004);
buf BUF1 (N4857, N4834);
xor XOR2 (N4858, N4854, N969);
and AND2 (N4859, N4852, N262);
and AND3 (N4860, N4847, N2882, N687);
nor NOR4 (N4861, N4858, N269, N4356, N275);
and AND2 (N4862, N4856, N4074);
and AND4 (N4863, N4857, N2817, N1426, N2993);
and AND4 (N4864, N4861, N4648, N1134, N2817);
and AND3 (N4865, N4846, N1936, N2621);
nor NOR3 (N4866, N4862, N1981, N4773);
not NOT1 (N4867, N4853);
buf BUF1 (N4868, N4867);
and AND2 (N4869, N4842, N2499);
buf BUF1 (N4870, N4868);
and AND3 (N4871, N4860, N189, N3672);
nor NOR4 (N4872, N4869, N4362, N855, N1439);
xor XOR2 (N4873, N4841, N811);
not NOT1 (N4874, N4863);
or OR3 (N4875, N4874, N1696, N1725);
xor XOR2 (N4876, N4864, N240);
nand NAND4 (N4877, N4872, N2078, N3421, N4608);
nor NOR4 (N4878, N4875, N4394, N584, N3681);
and AND3 (N4879, N4855, N2641, N2298);
xor XOR2 (N4880, N4876, N1739);
and AND4 (N4881, N4878, N659, N3251, N3426);
buf BUF1 (N4882, N4866);
buf BUF1 (N4883, N4879);
nand NAND2 (N4884, N4882, N980);
nor NOR2 (N4885, N4871, N4309);
nand NAND3 (N4886, N4885, N3299, N1178);
not NOT1 (N4887, N4865);
buf BUF1 (N4888, N4873);
nor NOR3 (N4889, N4859, N3073, N2057);
not NOT1 (N4890, N4880);
or OR4 (N4891, N4888, N4125, N1102, N35);
not NOT1 (N4892, N4889);
or OR2 (N4893, N4870, N4493);
buf BUF1 (N4894, N4890);
xor XOR2 (N4895, N4877, N1246);
buf BUF1 (N4896, N4886);
nor NOR3 (N4897, N4884, N1381, N3457);
xor XOR2 (N4898, N4897, N4685);
or OR3 (N4899, N4893, N4303, N4621);
not NOT1 (N4900, N4892);
not NOT1 (N4901, N4900);
nor NOR4 (N4902, N4895, N2795, N4502, N3734);
xor XOR2 (N4903, N4898, N4674);
xor XOR2 (N4904, N4902, N3000);
buf BUF1 (N4905, N4887);
nor NOR2 (N4906, N4881, N901);
buf BUF1 (N4907, N4904);
and AND4 (N4908, N4906, N2041, N1150, N188);
not NOT1 (N4909, N4908);
xor XOR2 (N4910, N4909, N4510);
nor NOR3 (N4911, N4901, N1245, N3699);
xor XOR2 (N4912, N4883, N4313);
not NOT1 (N4913, N4899);
nor NOR2 (N4914, N4894, N1824);
not NOT1 (N4915, N4911);
nor NOR4 (N4916, N4905, N827, N13, N4671);
xor XOR2 (N4917, N4907, N898);
or OR3 (N4918, N4912, N393, N4432);
or OR2 (N4919, N4916, N1390);
xor XOR2 (N4920, N4917, N3719);
buf BUF1 (N4921, N4903);
nand NAND2 (N4922, N4918, N4093);
xor XOR2 (N4923, N4896, N3990);
nand NAND4 (N4924, N4920, N2059, N2662, N2364);
not NOT1 (N4925, N4923);
and AND2 (N4926, N4914, N1141);
and AND3 (N4927, N4925, N4043, N1206);
nand NAND4 (N4928, N4921, N605, N3144, N816);
nor NOR3 (N4929, N4915, N4641, N3505);
not NOT1 (N4930, N4924);
nand NAND2 (N4931, N4910, N4253);
not NOT1 (N4932, N4929);
nor NOR2 (N4933, N4926, N4665);
buf BUF1 (N4934, N4891);
and AND2 (N4935, N4913, N4745);
xor XOR2 (N4936, N4931, N3990);
or OR2 (N4937, N4932, N4342);
nand NAND4 (N4938, N4934, N421, N1232, N2812);
nor NOR2 (N4939, N4938, N3254);
or OR2 (N4940, N4928, N4909);
or OR2 (N4941, N4933, N2827);
and AND4 (N4942, N4919, N3376, N1630, N4418);
buf BUF1 (N4943, N4937);
and AND4 (N4944, N4943, N3683, N1502, N3378);
buf BUF1 (N4945, N4940);
not NOT1 (N4946, N4930);
or OR4 (N4947, N4927, N2470, N4584, N1437);
or OR3 (N4948, N4922, N1223, N1742);
or OR4 (N4949, N4941, N1530, N1453, N4087);
xor XOR2 (N4950, N4939, N1330);
nand NAND3 (N4951, N4948, N197, N485);
or OR3 (N4952, N4946, N4868, N1048);
nor NOR3 (N4953, N4942, N2913, N395);
and AND3 (N4954, N4945, N4666, N4927);
nor NOR4 (N4955, N4954, N3508, N1336, N1336);
buf BUF1 (N4956, N4947);
not NOT1 (N4957, N4955);
not NOT1 (N4958, N4957);
buf BUF1 (N4959, N4951);
nand NAND4 (N4960, N4958, N4544, N4876, N4599);
nor NOR4 (N4961, N4936, N4506, N4051, N1936);
xor XOR2 (N4962, N4961, N1400);
and AND3 (N4963, N4952, N3760, N2463);
nor NOR2 (N4964, N4963, N1652);
nor NOR3 (N4965, N4964, N4915, N3895);
not NOT1 (N4966, N4935);
or OR2 (N4967, N4962, N3956);
and AND4 (N4968, N4959, N3550, N4597, N2543);
xor XOR2 (N4969, N4956, N2303);
buf BUF1 (N4970, N4953);
nand NAND2 (N4971, N4970, N3336);
or OR4 (N4972, N4949, N788, N4400, N4309);
xor XOR2 (N4973, N4969, N564);
not NOT1 (N4974, N4968);
xor XOR2 (N4975, N4950, N3067);
not NOT1 (N4976, N4960);
nor NOR2 (N4977, N4966, N4937);
xor XOR2 (N4978, N4967, N4798);
nor NOR2 (N4979, N4978, N2716);
or OR2 (N4980, N4972, N1826);
and AND4 (N4981, N4980, N880, N311, N3265);
not NOT1 (N4982, N4944);
not NOT1 (N4983, N4981);
nor NOR4 (N4984, N4974, N3081, N2026, N856);
nor NOR3 (N4985, N4983, N4659, N3221);
or OR4 (N4986, N4979, N4775, N1737, N2708);
not NOT1 (N4987, N4986);
buf BUF1 (N4988, N4982);
nor NOR3 (N4989, N4973, N954, N1983);
not NOT1 (N4990, N4987);
xor XOR2 (N4991, N4965, N1132);
not NOT1 (N4992, N4990);
buf BUF1 (N4993, N4992);
nor NOR2 (N4994, N4976, N3475);
or OR3 (N4995, N4988, N4046, N4);
nand NAND3 (N4996, N4971, N3658, N668);
not NOT1 (N4997, N4995);
nand NAND3 (N4998, N4993, N4240, N3485);
xor XOR2 (N4999, N4996, N2472);
or OR3 (N5000, N4997, N12, N2348);
and AND2 (N5001, N4994, N4066);
xor XOR2 (N5002, N4977, N2436);
and AND4 (N5003, N4999, N43, N2203, N2134);
nand NAND4 (N5004, N4975, N3219, N924, N4255);
not NOT1 (N5005, N4989);
xor XOR2 (N5006, N5003, N3327);
nand NAND3 (N5007, N4984, N1512, N4037);
and AND2 (N5008, N4998, N3859);
or OR3 (N5009, N5006, N204, N3306);
nand NAND2 (N5010, N5004, N3064);
xor XOR2 (N5011, N5005, N1409);
xor XOR2 (N5012, N5001, N4147);
xor XOR2 (N5013, N5011, N4540);
xor XOR2 (N5014, N5013, N3426);
nor NOR3 (N5015, N5000, N1121, N4309);
buf BUF1 (N5016, N5014);
or OR4 (N5017, N4985, N3823, N1894, N2045);
nand NAND2 (N5018, N5015, N2892);
xor XOR2 (N5019, N5002, N3286);
and AND3 (N5020, N5019, N2842, N221);
nand NAND4 (N5021, N5009, N655, N466, N65);
and AND3 (N5022, N5016, N3861, N2918);
buf BUF1 (N5023, N5008);
nor NOR4 (N5024, N5022, N4791, N2710, N2198);
and AND2 (N5025, N5023, N3570);
or OR2 (N5026, N5024, N3838);
nor NOR2 (N5027, N5026, N4348);
or OR2 (N5028, N5010, N780);
nand NAND2 (N5029, N5012, N3705);
not NOT1 (N5030, N5018);
and AND2 (N5031, N5021, N3196);
and AND4 (N5032, N5030, N3672, N1215, N2389);
xor XOR2 (N5033, N5032, N4734);
xor XOR2 (N5034, N5007, N811);
and AND2 (N5035, N5031, N4560);
not NOT1 (N5036, N5035);
or OR2 (N5037, N5033, N931);
or OR3 (N5038, N5029, N2094, N2300);
nor NOR3 (N5039, N5037, N2038, N1923);
and AND4 (N5040, N5034, N1999, N641, N3243);
and AND2 (N5041, N5040, N1143);
or OR2 (N5042, N5041, N367);
xor XOR2 (N5043, N5025, N162);
buf BUF1 (N5044, N5043);
buf BUF1 (N5045, N5020);
and AND4 (N5046, N5039, N4527, N3613, N344);
nand NAND2 (N5047, N5028, N92);
buf BUF1 (N5048, N5042);
not NOT1 (N5049, N5027);
buf BUF1 (N5050, N5045);
and AND4 (N5051, N5017, N327, N819, N4358);
nor NOR4 (N5052, N5046, N3896, N1665, N267);
nor NOR2 (N5053, N5050, N208);
xor XOR2 (N5054, N5051, N4164);
buf BUF1 (N5055, N5049);
or OR2 (N5056, N5036, N773);
not NOT1 (N5057, N5055);
and AND2 (N5058, N5052, N236);
nor NOR2 (N5059, N5058, N1157);
or OR3 (N5060, N5048, N347, N4117);
not NOT1 (N5061, N5047);
nor NOR2 (N5062, N5056, N629);
nor NOR4 (N5063, N5054, N3841, N1905, N18);
or OR2 (N5064, N5059, N1148);
or OR4 (N5065, N5063, N3197, N721, N5009);
not NOT1 (N5066, N5061);
and AND3 (N5067, N5057, N4423, N4302);
nor NOR3 (N5068, N5062, N1748, N600);
xor XOR2 (N5069, N5065, N2195);
not NOT1 (N5070, N5066);
nand NAND4 (N5071, N5060, N4135, N3169, N3966);
and AND4 (N5072, N5044, N1499, N2723, N4713);
nand NAND4 (N5073, N5069, N3225, N2412, N1503);
not NOT1 (N5074, N5053);
and AND3 (N5075, N5073, N4958, N3870);
nand NAND3 (N5076, N5064, N3386, N3276);
buf BUF1 (N5077, N5072);
xor XOR2 (N5078, N5070, N1536);
not NOT1 (N5079, N5077);
or OR4 (N5080, N5068, N4816, N3939, N3024);
buf BUF1 (N5081, N5071);
xor XOR2 (N5082, N5067, N3421);
buf BUF1 (N5083, N5078);
or OR4 (N5084, N5075, N4967, N3198, N5005);
xor XOR2 (N5085, N5074, N1590);
nand NAND3 (N5086, N5076, N1601, N3445);
and AND2 (N5087, N5086, N4100);
nor NOR2 (N5088, N5081, N3410);
xor XOR2 (N5089, N5083, N2835);
nor NOR4 (N5090, N4991, N365, N3855, N3398);
nand NAND2 (N5091, N5084, N987);
nand NAND4 (N5092, N5091, N461, N505, N1453);
not NOT1 (N5093, N5090);
nand NAND3 (N5094, N5038, N1918, N3142);
and AND2 (N5095, N5085, N1529);
nand NAND3 (N5096, N5092, N1016, N1538);
not NOT1 (N5097, N5080);
nor NOR2 (N5098, N5093, N3297);
or OR3 (N5099, N5094, N890, N3350);
or OR3 (N5100, N5096, N3115, N1105);
and AND4 (N5101, N5082, N824, N4446, N115);
nand NAND2 (N5102, N5089, N2985);
nor NOR4 (N5103, N5087, N2216, N1690, N2378);
xor XOR2 (N5104, N5103, N3124);
buf BUF1 (N5105, N5079);
nor NOR2 (N5106, N5104, N4929);
nor NOR3 (N5107, N5095, N3629, N1166);
xor XOR2 (N5108, N5101, N2267);
xor XOR2 (N5109, N5100, N3211);
and AND2 (N5110, N5099, N603);
or OR2 (N5111, N5109, N4338);
nor NOR4 (N5112, N5111, N4546, N63, N2010);
not NOT1 (N5113, N5106);
or OR3 (N5114, N5112, N2690, N3668);
and AND4 (N5115, N5107, N734, N2845, N309);
buf BUF1 (N5116, N5114);
nor NOR4 (N5117, N5116, N1851, N581, N1087);
buf BUF1 (N5118, N5097);
buf BUF1 (N5119, N5098);
and AND3 (N5120, N5115, N2653, N1173);
nand NAND3 (N5121, N5108, N1425, N2773);
or OR2 (N5122, N5088, N2886);
and AND2 (N5123, N5113, N1522);
nand NAND2 (N5124, N5117, N1050);
and AND2 (N5125, N5124, N2111);
and AND2 (N5126, N5123, N2497);
and AND2 (N5127, N5121, N3048);
nand NAND4 (N5128, N5122, N2288, N4443, N4661);
nor NOR4 (N5129, N5105, N4869, N4572, N1754);
and AND4 (N5130, N5128, N3747, N894, N2121);
nor NOR2 (N5131, N5127, N2579);
nand NAND4 (N5132, N5126, N1951, N797, N140);
nor NOR2 (N5133, N5129, N2860);
buf BUF1 (N5134, N5133);
xor XOR2 (N5135, N5125, N4432);
xor XOR2 (N5136, N5131, N2263);
or OR4 (N5137, N5134, N1317, N4334, N270);
nand NAND3 (N5138, N5118, N2806, N2021);
buf BUF1 (N5139, N5110);
xor XOR2 (N5140, N5119, N2379);
not NOT1 (N5141, N5138);
not NOT1 (N5142, N5140);
buf BUF1 (N5143, N5136);
not NOT1 (N5144, N5142);
or OR3 (N5145, N5135, N4531, N4791);
and AND3 (N5146, N5141, N418, N1528);
or OR4 (N5147, N5143, N4783, N420, N636);
xor XOR2 (N5148, N5144, N4693);
or OR3 (N5149, N5145, N933, N4821);
and AND4 (N5150, N5149, N789, N4801, N3735);
nand NAND2 (N5151, N5102, N4978);
or OR4 (N5152, N5130, N108, N2340, N640);
nor NOR3 (N5153, N5139, N2261, N301);
not NOT1 (N5154, N5152);
buf BUF1 (N5155, N5132);
xor XOR2 (N5156, N5150, N433);
and AND3 (N5157, N5147, N75, N2121);
and AND3 (N5158, N5148, N2128, N59);
buf BUF1 (N5159, N5157);
nor NOR2 (N5160, N5156, N1590);
nand NAND2 (N5161, N5159, N2600);
and AND4 (N5162, N5120, N2540, N3149, N2539);
or OR2 (N5163, N5158, N611);
xor XOR2 (N5164, N5137, N4826);
and AND2 (N5165, N5153, N4417);
nand NAND4 (N5166, N5146, N4813, N4686, N791);
nor NOR4 (N5167, N5155, N4361, N285, N4259);
and AND4 (N5168, N5161, N4618, N1998, N3205);
nand NAND2 (N5169, N5160, N859);
and AND2 (N5170, N5167, N3390);
buf BUF1 (N5171, N5164);
or OR4 (N5172, N5169, N366, N5042, N3135);
and AND3 (N5173, N5168, N2019, N4669);
xor XOR2 (N5174, N5163, N1220);
nor NOR4 (N5175, N5154, N4203, N3788, N1222);
or OR3 (N5176, N5170, N4089, N1714);
not NOT1 (N5177, N5172);
buf BUF1 (N5178, N5176);
or OR2 (N5179, N5166, N3439);
buf BUF1 (N5180, N5173);
buf BUF1 (N5181, N5180);
or OR4 (N5182, N5165, N3889, N752, N1226);
xor XOR2 (N5183, N5177, N3940);
not NOT1 (N5184, N5183);
buf BUF1 (N5185, N5181);
and AND3 (N5186, N5175, N2816, N2623);
or OR2 (N5187, N5182, N4866);
buf BUF1 (N5188, N5178);
buf BUF1 (N5189, N5187);
or OR4 (N5190, N5186, N3236, N3558, N4129);
nor NOR3 (N5191, N5171, N4505, N2001);
not NOT1 (N5192, N5151);
not NOT1 (N5193, N5179);
and AND4 (N5194, N5188, N2291, N2654, N3636);
or OR4 (N5195, N5174, N3131, N3746, N2870);
xor XOR2 (N5196, N5190, N3973);
not NOT1 (N5197, N5193);
or OR3 (N5198, N5185, N1801, N1297);
nor NOR2 (N5199, N5196, N3468);
not NOT1 (N5200, N5189);
xor XOR2 (N5201, N5191, N1815);
or OR2 (N5202, N5194, N2034);
and AND3 (N5203, N5197, N5098, N1488);
or OR3 (N5204, N5200, N3676, N1590);
buf BUF1 (N5205, N5198);
not NOT1 (N5206, N5204);
or OR4 (N5207, N5195, N993, N2481, N1517);
nor NOR2 (N5208, N5192, N3398);
buf BUF1 (N5209, N5205);
or OR3 (N5210, N5199, N2019, N1031);
buf BUF1 (N5211, N5207);
not NOT1 (N5212, N5162);
nor NOR2 (N5213, N5203, N3010);
not NOT1 (N5214, N5184);
nand NAND4 (N5215, N5210, N2353, N3975, N3250);
buf BUF1 (N5216, N5208);
nor NOR3 (N5217, N5209, N483, N1150);
nor NOR2 (N5218, N5211, N4211);
or OR2 (N5219, N5201, N896);
or OR4 (N5220, N5218, N4674, N410, N1191);
not NOT1 (N5221, N5212);
xor XOR2 (N5222, N5216, N1255);
xor XOR2 (N5223, N5213, N2909);
buf BUF1 (N5224, N5220);
xor XOR2 (N5225, N5206, N4971);
and AND4 (N5226, N5215, N3575, N4587, N1991);
and AND3 (N5227, N5224, N5115, N3200);
nor NOR4 (N5228, N5225, N4854, N4987, N3775);
or OR2 (N5229, N5228, N2454);
not NOT1 (N5230, N5221);
and AND2 (N5231, N5217, N4688);
buf BUF1 (N5232, N5202);
xor XOR2 (N5233, N5214, N1497);
or OR2 (N5234, N5223, N3182);
nand NAND4 (N5235, N5229, N347, N1721, N1630);
xor XOR2 (N5236, N5235, N68);
not NOT1 (N5237, N5230);
or OR3 (N5238, N5227, N4913, N194);
nor NOR3 (N5239, N5222, N2824, N706);
nor NOR3 (N5240, N5234, N1572, N5150);
not NOT1 (N5241, N5233);
xor XOR2 (N5242, N5238, N2125);
or OR2 (N5243, N5232, N1346);
or OR3 (N5244, N5242, N1260, N4001);
nand NAND3 (N5245, N5243, N4803, N5142);
buf BUF1 (N5246, N5226);
not NOT1 (N5247, N5241);
nor NOR2 (N5248, N5236, N5057);
not NOT1 (N5249, N5244);
nand NAND2 (N5250, N5231, N822);
nand NAND4 (N5251, N5219, N4606, N5128, N2039);
not NOT1 (N5252, N5246);
or OR4 (N5253, N5237, N325, N2649, N784);
xor XOR2 (N5254, N5249, N422);
or OR3 (N5255, N5251, N704, N2405);
not NOT1 (N5256, N5255);
xor XOR2 (N5257, N5253, N2978);
xor XOR2 (N5258, N5248, N829);
nor NOR2 (N5259, N5254, N2146);
nor NOR3 (N5260, N5256, N2951, N3971);
and AND3 (N5261, N5239, N511, N1324);
or OR4 (N5262, N5258, N2186, N3041, N4758);
nor NOR4 (N5263, N5259, N4831, N4361, N2710);
buf BUF1 (N5264, N5247);
nor NOR2 (N5265, N5240, N4768);
not NOT1 (N5266, N5261);
or OR4 (N5267, N5266, N3212, N1171, N3911);
xor XOR2 (N5268, N5250, N2132);
and AND4 (N5269, N5245, N2209, N2357, N4706);
xor XOR2 (N5270, N5269, N4602);
buf BUF1 (N5271, N5252);
nor NOR3 (N5272, N5271, N1730, N1924);
and AND3 (N5273, N5272, N5005, N2452);
not NOT1 (N5274, N5260);
buf BUF1 (N5275, N5257);
nor NOR3 (N5276, N5262, N1628, N2106);
or OR3 (N5277, N5274, N230, N4567);
nor NOR3 (N5278, N5275, N5093, N4915);
buf BUF1 (N5279, N5265);
or OR4 (N5280, N5277, N1649, N2421, N3540);
buf BUF1 (N5281, N5278);
or OR3 (N5282, N5264, N2097, N3077);
not NOT1 (N5283, N5276);
xor XOR2 (N5284, N5280, N2277);
buf BUF1 (N5285, N5279);
nand NAND2 (N5286, N5267, N3160);
nand NAND3 (N5287, N5284, N3356, N1995);
xor XOR2 (N5288, N5285, N1978);
xor XOR2 (N5289, N5268, N1406);
and AND4 (N5290, N5283, N4256, N5263, N3448);
and AND4 (N5291, N1774, N4678, N933, N1272);
not NOT1 (N5292, N5290);
nor NOR3 (N5293, N5291, N1443, N1099);
not NOT1 (N5294, N5286);
buf BUF1 (N5295, N5288);
not NOT1 (N5296, N5287);
buf BUF1 (N5297, N5282);
buf BUF1 (N5298, N5273);
xor XOR2 (N5299, N5270, N2421);
buf BUF1 (N5300, N5297);
xor XOR2 (N5301, N5295, N1557);
or OR4 (N5302, N5300, N1755, N3044, N3296);
and AND3 (N5303, N5289, N1601, N711);
nor NOR4 (N5304, N5298, N712, N4446, N5220);
nand NAND3 (N5305, N5292, N1154, N3380);
nand NAND2 (N5306, N5303, N3193);
xor XOR2 (N5307, N5306, N5185);
buf BUF1 (N5308, N5299);
xor XOR2 (N5309, N5281, N509);
nand NAND4 (N5310, N5304, N3751, N1251, N648);
buf BUF1 (N5311, N5302);
and AND4 (N5312, N5301, N373, N848, N2414);
xor XOR2 (N5313, N5312, N959);
and AND2 (N5314, N5293, N4446);
buf BUF1 (N5315, N5311);
nor NOR2 (N5316, N5294, N678);
nand NAND3 (N5317, N5310, N1816, N3383);
or OR2 (N5318, N5317, N3943);
nand NAND2 (N5319, N5313, N682);
or OR3 (N5320, N5318, N3577, N1946);
nand NAND4 (N5321, N5308, N4517, N2355, N3662);
xor XOR2 (N5322, N5307, N5045);
nand NAND2 (N5323, N5316, N1697);
buf BUF1 (N5324, N5320);
or OR3 (N5325, N5315, N2698, N3573);
nand NAND4 (N5326, N5305, N4785, N1899, N1246);
nor NOR2 (N5327, N5325, N4899);
or OR2 (N5328, N5324, N916);
buf BUF1 (N5329, N5327);
nand NAND3 (N5330, N5328, N2506, N2355);
nor NOR2 (N5331, N5326, N3291);
xor XOR2 (N5332, N5314, N4410);
nand NAND4 (N5333, N5309, N4018, N3405, N3395);
xor XOR2 (N5334, N5322, N3941);
buf BUF1 (N5335, N5330);
xor XOR2 (N5336, N5329, N4930);
xor XOR2 (N5337, N5335, N3121);
not NOT1 (N5338, N5336);
xor XOR2 (N5339, N5338, N1785);
buf BUF1 (N5340, N5332);
not NOT1 (N5341, N5296);
not NOT1 (N5342, N5331);
nand NAND3 (N5343, N5323, N3024, N3431);
xor XOR2 (N5344, N5319, N3733);
not NOT1 (N5345, N5321);
buf BUF1 (N5346, N5337);
or OR2 (N5347, N5341, N836);
buf BUF1 (N5348, N5333);
xor XOR2 (N5349, N5342, N1309);
nor NOR4 (N5350, N5344, N2998, N2004, N3141);
nand NAND2 (N5351, N5343, N4589);
and AND4 (N5352, N5346, N4054, N700, N3672);
xor XOR2 (N5353, N5348, N20);
or OR2 (N5354, N5349, N749);
nand NAND3 (N5355, N5350, N2768, N5141);
nor NOR2 (N5356, N5355, N350);
xor XOR2 (N5357, N5345, N4266);
and AND2 (N5358, N5351, N2622);
nor NOR4 (N5359, N5353, N1097, N3543, N4844);
and AND4 (N5360, N5359, N3729, N4535, N1715);
nor NOR3 (N5361, N5352, N5127, N3384);
or OR3 (N5362, N5354, N441, N2404);
buf BUF1 (N5363, N5356);
nand NAND3 (N5364, N5357, N2506, N4562);
and AND2 (N5365, N5358, N2217);
nor NOR3 (N5366, N5361, N781, N844);
xor XOR2 (N5367, N5339, N4495);
xor XOR2 (N5368, N5347, N879);
or OR4 (N5369, N5340, N360, N1884, N1440);
not NOT1 (N5370, N5368);
and AND3 (N5371, N5367, N3443, N1307);
or OR3 (N5372, N5365, N4535, N5291);
and AND2 (N5373, N5371, N3540);
nor NOR2 (N5374, N5373, N92);
nor NOR2 (N5375, N5364, N4199);
xor XOR2 (N5376, N5366, N4338);
xor XOR2 (N5377, N5370, N4196);
nor NOR3 (N5378, N5360, N4836, N2345);
or OR3 (N5379, N5369, N2443, N737);
nor NOR3 (N5380, N5378, N3635, N4463);
nand NAND4 (N5381, N5374, N2357, N2187, N4182);
or OR2 (N5382, N5372, N4772);
buf BUF1 (N5383, N5376);
xor XOR2 (N5384, N5375, N3094);
buf BUF1 (N5385, N5382);
not NOT1 (N5386, N5384);
and AND4 (N5387, N5381, N5021, N820, N1564);
buf BUF1 (N5388, N5383);
buf BUF1 (N5389, N5377);
buf BUF1 (N5390, N5380);
nand NAND4 (N5391, N5385, N4903, N872, N4453);
nor NOR4 (N5392, N5334, N750, N1772, N4835);
or OR3 (N5393, N5379, N2919, N4250);
and AND4 (N5394, N5388, N492, N4144, N2264);
and AND3 (N5395, N5391, N494, N92);
and AND3 (N5396, N5395, N353, N4992);
or OR4 (N5397, N5389, N597, N344, N1378);
and AND3 (N5398, N5397, N5210, N799);
nand NAND2 (N5399, N5390, N612);
not NOT1 (N5400, N5363);
not NOT1 (N5401, N5399);
or OR4 (N5402, N5393, N930, N1292, N2374);
buf BUF1 (N5403, N5401);
or OR2 (N5404, N5386, N3883);
nand NAND2 (N5405, N5394, N4824);
buf BUF1 (N5406, N5405);
xor XOR2 (N5407, N5362, N442);
xor XOR2 (N5408, N5404, N3346);
nor NOR2 (N5409, N5392, N3478);
or OR2 (N5410, N5408, N947);
nand NAND2 (N5411, N5410, N5382);
not NOT1 (N5412, N5396);
nor NOR2 (N5413, N5409, N5283);
buf BUF1 (N5414, N5407);
buf BUF1 (N5415, N5412);
xor XOR2 (N5416, N5402, N1971);
buf BUF1 (N5417, N5411);
and AND3 (N5418, N5387, N5294, N2974);
or OR4 (N5419, N5398, N4644, N572, N3205);
or OR4 (N5420, N5403, N1719, N1723, N1296);
nor NOR3 (N5421, N5400, N4800, N2774);
buf BUF1 (N5422, N5406);
nor NOR4 (N5423, N5414, N1115, N2963, N1302);
or OR3 (N5424, N5419, N3732, N4247);
not NOT1 (N5425, N5423);
nand NAND3 (N5426, N5425, N4744, N3062);
and AND4 (N5427, N5415, N2626, N1008, N2464);
and AND4 (N5428, N5418, N1106, N1179, N3586);
and AND2 (N5429, N5413, N4917);
or OR4 (N5430, N5420, N4213, N2833, N1751);
buf BUF1 (N5431, N5429);
not NOT1 (N5432, N5424);
or OR2 (N5433, N5421, N4417);
not NOT1 (N5434, N5417);
nand NAND2 (N5435, N5431, N799);
xor XOR2 (N5436, N5432, N2055);
xor XOR2 (N5437, N5426, N369);
and AND3 (N5438, N5428, N3681, N1271);
or OR2 (N5439, N5416, N3763);
not NOT1 (N5440, N5438);
nand NAND2 (N5441, N5435, N3998);
or OR2 (N5442, N5439, N2316);
and AND3 (N5443, N5440, N4302, N2331);
or OR3 (N5444, N5442, N4766, N1209);
nor NOR3 (N5445, N5430, N3207, N5162);
and AND3 (N5446, N5444, N1237, N4391);
nor NOR3 (N5447, N5443, N1720, N388);
buf BUF1 (N5448, N5434);
or OR2 (N5449, N5446, N3132);
or OR2 (N5450, N5436, N1429);
nor NOR2 (N5451, N5437, N1815);
nor NOR3 (N5452, N5441, N4328, N2137);
not NOT1 (N5453, N5447);
and AND2 (N5454, N5450, N2108);
or OR3 (N5455, N5453, N4991, N1058);
buf BUF1 (N5456, N5427);
not NOT1 (N5457, N5452);
and AND4 (N5458, N5454, N3366, N2938, N2991);
nand NAND2 (N5459, N5433, N303);
not NOT1 (N5460, N5449);
not NOT1 (N5461, N5455);
nor NOR4 (N5462, N5445, N5241, N1979, N4833);
nand NAND2 (N5463, N5458, N968);
nor NOR2 (N5464, N5457, N1058);
nor NOR4 (N5465, N5461, N171, N4389, N219);
and AND4 (N5466, N5463, N4242, N843, N1619);
nor NOR2 (N5467, N5451, N3332);
nor NOR3 (N5468, N5465, N2816, N3645);
and AND2 (N5469, N5448, N578);
nor NOR3 (N5470, N5422, N1293, N4641);
not NOT1 (N5471, N5464);
nor NOR3 (N5472, N5466, N3136, N2475);
buf BUF1 (N5473, N5469);
nand NAND2 (N5474, N5473, N3970);
not NOT1 (N5475, N5467);
or OR4 (N5476, N5462, N4642, N1479, N2727);
nor NOR4 (N5477, N5468, N668, N4180, N2737);
or OR3 (N5478, N5475, N4643, N2039);
or OR3 (N5479, N5476, N540, N4897);
or OR3 (N5480, N5479, N1898, N1778);
not NOT1 (N5481, N5474);
buf BUF1 (N5482, N5478);
nand NAND4 (N5483, N5471, N5087, N3304, N171);
not NOT1 (N5484, N5482);
and AND4 (N5485, N5459, N3907, N1, N3150);
nor NOR4 (N5486, N5485, N5050, N4607, N1739);
xor XOR2 (N5487, N5480, N1591);
or OR2 (N5488, N5481, N2947);
nand NAND3 (N5489, N5487, N1820, N709);
and AND3 (N5490, N5456, N2015, N3622);
or OR2 (N5491, N5470, N3075);
not NOT1 (N5492, N5460);
and AND2 (N5493, N5483, N4523);
buf BUF1 (N5494, N5492);
and AND3 (N5495, N5484, N797, N1056);
nor NOR2 (N5496, N5495, N1751);
and AND2 (N5497, N5490, N984);
nor NOR4 (N5498, N5497, N4387, N3514, N5254);
xor XOR2 (N5499, N5472, N868);
buf BUF1 (N5500, N5489);
and AND2 (N5501, N5486, N3004);
nand NAND3 (N5502, N5499, N2055, N1047);
nand NAND2 (N5503, N5477, N1993);
nand NAND4 (N5504, N5488, N648, N1181, N805);
not NOT1 (N5505, N5500);
buf BUF1 (N5506, N5493);
xor XOR2 (N5507, N5496, N485);
nor NOR2 (N5508, N5506, N1774);
or OR3 (N5509, N5498, N610, N4162);
nand NAND2 (N5510, N5504, N3112);
buf BUF1 (N5511, N5503);
nor NOR3 (N5512, N5494, N894, N3894);
nor NOR3 (N5513, N5505, N5172, N197);
nor NOR4 (N5514, N5491, N4705, N4026, N1134);
nand NAND3 (N5515, N5510, N4376, N656);
and AND2 (N5516, N5502, N3911);
and AND3 (N5517, N5516, N2255, N4467);
not NOT1 (N5518, N5511);
or OR3 (N5519, N5517, N618, N2213);
or OR3 (N5520, N5512, N3451, N5253);
not NOT1 (N5521, N5509);
not NOT1 (N5522, N5515);
nor NOR2 (N5523, N5501, N3536);
or OR3 (N5524, N5518, N1429, N3410);
not NOT1 (N5525, N5519);
buf BUF1 (N5526, N5513);
nor NOR2 (N5527, N5507, N2091);
nand NAND2 (N5528, N5520, N2852);
and AND3 (N5529, N5524, N3309, N2597);
buf BUF1 (N5530, N5529);
and AND2 (N5531, N5523, N2408);
xor XOR2 (N5532, N5531, N2262);
buf BUF1 (N5533, N5514);
xor XOR2 (N5534, N5508, N3111);
not NOT1 (N5535, N5521);
and AND4 (N5536, N5525, N4148, N428, N2816);
and AND2 (N5537, N5526, N3721);
nor NOR3 (N5538, N5530, N2354, N2357);
nand NAND2 (N5539, N5537, N2244);
buf BUF1 (N5540, N5528);
or OR2 (N5541, N5540, N3679);
xor XOR2 (N5542, N5532, N1362);
nor NOR4 (N5543, N5533, N4115, N4382, N4563);
nor NOR2 (N5544, N5538, N3613);
xor XOR2 (N5545, N5543, N2616);
not NOT1 (N5546, N5522);
and AND3 (N5547, N5539, N5281, N2698);
nand NAND4 (N5548, N5542, N2565, N1763, N2699);
not NOT1 (N5549, N5547);
not NOT1 (N5550, N5548);
nand NAND2 (N5551, N5541, N5059);
or OR2 (N5552, N5535, N3359);
nor NOR2 (N5553, N5545, N251);
not NOT1 (N5554, N5536);
nand NAND2 (N5555, N5552, N3854);
buf BUF1 (N5556, N5555);
or OR3 (N5557, N5556, N5140, N4885);
nand NAND3 (N5558, N5553, N276, N3594);
or OR2 (N5559, N5534, N2900);
buf BUF1 (N5560, N5527);
nand NAND3 (N5561, N5544, N2675, N1411);
and AND4 (N5562, N5550, N5091, N2442, N286);
nand NAND2 (N5563, N5559, N3380);
xor XOR2 (N5564, N5563, N4224);
buf BUF1 (N5565, N5546);
xor XOR2 (N5566, N5558, N2628);
and AND4 (N5567, N5565, N1843, N3026, N1089);
xor XOR2 (N5568, N5549, N803);
xor XOR2 (N5569, N5561, N2344);
not NOT1 (N5570, N5564);
and AND3 (N5571, N5570, N2019, N2301);
and AND4 (N5572, N5568, N1280, N4193, N167);
or OR2 (N5573, N5562, N935);
xor XOR2 (N5574, N5554, N4965);
nand NAND4 (N5575, N5557, N4367, N4466, N1749);
nand NAND2 (N5576, N5567, N2991);
or OR4 (N5577, N5560, N4119, N3312, N382);
nand NAND3 (N5578, N5551, N4637, N5213);
not NOT1 (N5579, N5566);
xor XOR2 (N5580, N5575, N5056);
buf BUF1 (N5581, N5574);
xor XOR2 (N5582, N5580, N4210);
xor XOR2 (N5583, N5578, N1019);
nand NAND2 (N5584, N5573, N5149);
and AND3 (N5585, N5579, N1564, N3207);
nand NAND3 (N5586, N5577, N272, N2154);
not NOT1 (N5587, N5571);
nor NOR3 (N5588, N5587, N397, N4242);
not NOT1 (N5589, N5584);
or OR4 (N5590, N5582, N884, N3821, N1023);
nand NAND2 (N5591, N5586, N759);
nand NAND3 (N5592, N5590, N1836, N1618);
not NOT1 (N5593, N5581);
nand NAND4 (N5594, N5591, N4597, N439, N2175);
nand NAND2 (N5595, N5585, N347);
or OR2 (N5596, N5589, N1168);
xor XOR2 (N5597, N5594, N1720);
or OR3 (N5598, N5576, N258, N2050);
and AND2 (N5599, N5572, N4285);
nand NAND2 (N5600, N5599, N3850);
xor XOR2 (N5601, N5598, N764);
not NOT1 (N5602, N5569);
buf BUF1 (N5603, N5597);
not NOT1 (N5604, N5588);
and AND2 (N5605, N5583, N896);
xor XOR2 (N5606, N5595, N2533);
or OR4 (N5607, N5592, N967, N3832, N4114);
and AND2 (N5608, N5606, N4070);
nor NOR4 (N5609, N5604, N1507, N832, N4306);
not NOT1 (N5610, N5605);
or OR2 (N5611, N5602, N1108);
buf BUF1 (N5612, N5603);
not NOT1 (N5613, N5611);
xor XOR2 (N5614, N5612, N4051);
xor XOR2 (N5615, N5607, N4095);
buf BUF1 (N5616, N5600);
xor XOR2 (N5617, N5613, N2690);
nand NAND3 (N5618, N5610, N4858, N2194);
xor XOR2 (N5619, N5608, N2110);
not NOT1 (N5620, N5618);
nand NAND4 (N5621, N5616, N3984, N1642, N650);
and AND2 (N5622, N5601, N5107);
not NOT1 (N5623, N5621);
xor XOR2 (N5624, N5609, N4136);
not NOT1 (N5625, N5620);
xor XOR2 (N5626, N5622, N3460);
nor NOR3 (N5627, N5624, N2708, N1507);
xor XOR2 (N5628, N5617, N4968);
xor XOR2 (N5629, N5593, N3237);
or OR2 (N5630, N5619, N2879);
and AND4 (N5631, N5630, N4097, N1360, N3016);
and AND3 (N5632, N5628, N5197, N1281);
nor NOR2 (N5633, N5632, N2995);
buf BUF1 (N5634, N5596);
nand NAND3 (N5635, N5627, N708, N4145);
xor XOR2 (N5636, N5635, N2725);
not NOT1 (N5637, N5615);
xor XOR2 (N5638, N5625, N229);
and AND3 (N5639, N5633, N1441, N4157);
or OR2 (N5640, N5614, N4415);
xor XOR2 (N5641, N5626, N2334);
and AND4 (N5642, N5637, N4678, N2958, N4269);
or OR3 (N5643, N5636, N3271, N1958);
nand NAND3 (N5644, N5629, N154, N3409);
not NOT1 (N5645, N5643);
nand NAND2 (N5646, N5638, N4586);
nand NAND3 (N5647, N5641, N3902, N2589);
buf BUF1 (N5648, N5645);
or OR2 (N5649, N5647, N1733);
buf BUF1 (N5650, N5640);
and AND4 (N5651, N5634, N3830, N2840, N5077);
buf BUF1 (N5652, N5631);
buf BUF1 (N5653, N5639);
or OR3 (N5654, N5652, N1412, N2499);
nand NAND4 (N5655, N5649, N4201, N1875, N4260);
xor XOR2 (N5656, N5646, N2785);
buf BUF1 (N5657, N5651);
and AND2 (N5658, N5655, N1054);
xor XOR2 (N5659, N5644, N2266);
nor NOR3 (N5660, N5658, N3614, N5409);
not NOT1 (N5661, N5648);
xor XOR2 (N5662, N5642, N4946);
nand NAND2 (N5663, N5662, N1427);
buf BUF1 (N5664, N5661);
not NOT1 (N5665, N5664);
nor NOR4 (N5666, N5650, N1795, N5207, N2071);
buf BUF1 (N5667, N5660);
or OR3 (N5668, N5663, N4855, N3780);
or OR3 (N5669, N5653, N2017, N1941);
and AND2 (N5670, N5659, N4454);
nand NAND4 (N5671, N5667, N5518, N2468, N445);
nand NAND3 (N5672, N5670, N5144, N437);
not NOT1 (N5673, N5669);
nand NAND2 (N5674, N5665, N169);
nand NAND4 (N5675, N5673, N5672, N2384, N2905);
buf BUF1 (N5676, N1003);
and AND2 (N5677, N5654, N5376);
xor XOR2 (N5678, N5623, N5194);
nand NAND3 (N5679, N5668, N4720, N212);
xor XOR2 (N5680, N5679, N4318);
or OR2 (N5681, N5657, N5134);
nor NOR2 (N5682, N5676, N1350);
buf BUF1 (N5683, N5682);
not NOT1 (N5684, N5674);
and AND2 (N5685, N5680, N2088);
not NOT1 (N5686, N5677);
xor XOR2 (N5687, N5671, N2738);
buf BUF1 (N5688, N5685);
nand NAND2 (N5689, N5684, N1469);
nor NOR3 (N5690, N5686, N4216, N5306);
or OR2 (N5691, N5688, N5215);
nand NAND2 (N5692, N5666, N201);
or OR3 (N5693, N5690, N596, N5294);
buf BUF1 (N5694, N5683);
not NOT1 (N5695, N5692);
not NOT1 (N5696, N5693);
nand NAND2 (N5697, N5694, N4774);
buf BUF1 (N5698, N5681);
and AND3 (N5699, N5675, N3064, N2351);
and AND2 (N5700, N5687, N1614);
nor NOR3 (N5701, N5678, N1695, N3948);
and AND4 (N5702, N5698, N2581, N3526, N718);
or OR4 (N5703, N5689, N2532, N626, N240);
or OR3 (N5704, N5703, N3507, N4443);
not NOT1 (N5705, N5701);
not NOT1 (N5706, N5700);
buf BUF1 (N5707, N5656);
or OR3 (N5708, N5704, N1417, N810);
or OR3 (N5709, N5705, N1251, N3655);
and AND2 (N5710, N5707, N2486);
buf BUF1 (N5711, N5696);
not NOT1 (N5712, N5709);
buf BUF1 (N5713, N5712);
nor NOR3 (N5714, N5708, N3429, N4599);
not NOT1 (N5715, N5697);
nor NOR3 (N5716, N5715, N4358, N658);
buf BUF1 (N5717, N5714);
nand NAND4 (N5718, N5706, N3764, N4041, N5685);
not NOT1 (N5719, N5691);
and AND3 (N5720, N5717, N2730, N3674);
buf BUF1 (N5721, N5713);
xor XOR2 (N5722, N5702, N2459);
nand NAND3 (N5723, N5695, N2005, N1327);
nand NAND4 (N5724, N5711, N5355, N590, N3381);
or OR3 (N5725, N5721, N1438, N201);
xor XOR2 (N5726, N5720, N5224);
buf BUF1 (N5727, N5710);
or OR3 (N5728, N5723, N939, N26);
or OR3 (N5729, N5727, N2598, N4200);
buf BUF1 (N5730, N5716);
xor XOR2 (N5731, N5726, N1195);
nor NOR4 (N5732, N5731, N1402, N2821, N3276);
nor NOR2 (N5733, N5730, N3880);
xor XOR2 (N5734, N5733, N4897);
or OR2 (N5735, N5725, N2565);
not NOT1 (N5736, N5732);
not NOT1 (N5737, N5718);
or OR3 (N5738, N5724, N5549, N285);
and AND4 (N5739, N5738, N1825, N3075, N501);
nand NAND4 (N5740, N5736, N757, N4469, N4453);
xor XOR2 (N5741, N5735, N5607);
nor NOR2 (N5742, N5699, N2041);
buf BUF1 (N5743, N5728);
not NOT1 (N5744, N5739);
and AND3 (N5745, N5743, N4659, N418);
not NOT1 (N5746, N5737);
buf BUF1 (N5747, N5744);
nand NAND4 (N5748, N5747, N3204, N4716, N3196);
and AND2 (N5749, N5748, N3040);
buf BUF1 (N5750, N5719);
nand NAND3 (N5751, N5745, N5390, N2907);
not NOT1 (N5752, N5749);
nand NAND4 (N5753, N5740, N2254, N4376, N3010);
xor XOR2 (N5754, N5751, N1981);
or OR4 (N5755, N5742, N1689, N2989, N4917);
xor XOR2 (N5756, N5750, N5504);
not NOT1 (N5757, N5756);
nand NAND2 (N5758, N5734, N1800);
xor XOR2 (N5759, N5752, N2054);
and AND4 (N5760, N5746, N5253, N4819, N45);
xor XOR2 (N5761, N5758, N1269);
not NOT1 (N5762, N5755);
nor NOR4 (N5763, N5753, N2813, N5417, N629);
or OR4 (N5764, N5759, N711, N119, N1091);
nor NOR2 (N5765, N5741, N2381);
nand NAND3 (N5766, N5757, N650, N1376);
xor XOR2 (N5767, N5763, N4851);
and AND4 (N5768, N5762, N3625, N723, N1817);
not NOT1 (N5769, N5760);
nor NOR4 (N5770, N5761, N4062, N206, N2479);
nand NAND3 (N5771, N5766, N1580, N287);
or OR3 (N5772, N5729, N1364, N4869);
buf BUF1 (N5773, N5765);
not NOT1 (N5774, N5772);
and AND3 (N5775, N5774, N352, N1574);
nand NAND2 (N5776, N5768, N2947);
not NOT1 (N5777, N5776);
or OR2 (N5778, N5775, N3949);
xor XOR2 (N5779, N5770, N4467);
xor XOR2 (N5780, N5764, N158);
or OR3 (N5781, N5771, N143, N1319);
buf BUF1 (N5782, N5780);
or OR4 (N5783, N5782, N2874, N2090, N1144);
nor NOR4 (N5784, N5778, N1383, N3325, N5466);
nor NOR2 (N5785, N5779, N134);
and AND2 (N5786, N5785, N5291);
not NOT1 (N5787, N5783);
nor NOR2 (N5788, N5767, N4200);
nor NOR4 (N5789, N5781, N76, N1720, N635);
and AND4 (N5790, N5784, N1791, N3949, N3550);
nor NOR2 (N5791, N5722, N4061);
not NOT1 (N5792, N5754);
not NOT1 (N5793, N5788);
buf BUF1 (N5794, N5769);
nor NOR2 (N5795, N5790, N2486);
and AND2 (N5796, N5791, N5140);
xor XOR2 (N5797, N5796, N5376);
and AND4 (N5798, N5773, N1676, N3150, N3159);
not NOT1 (N5799, N5786);
xor XOR2 (N5800, N5799, N1316);
buf BUF1 (N5801, N5777);
or OR2 (N5802, N5787, N3420);
not NOT1 (N5803, N5793);
nand NAND2 (N5804, N5802, N1368);
or OR2 (N5805, N5792, N5521);
or OR2 (N5806, N5797, N4570);
not NOT1 (N5807, N5806);
nand NAND4 (N5808, N5801, N5398, N3308, N5409);
not NOT1 (N5809, N5800);
nor NOR3 (N5810, N5789, N5218, N3095);
and AND4 (N5811, N5808, N4988, N2905, N972);
xor XOR2 (N5812, N5803, N5592);
buf BUF1 (N5813, N5809);
and AND3 (N5814, N5810, N1072, N2569);
xor XOR2 (N5815, N5794, N4662);
nor NOR4 (N5816, N5804, N2829, N4149, N5807);
nor NOR4 (N5817, N2053, N365, N5773, N4453);
nor NOR3 (N5818, N5815, N4131, N2257);
not NOT1 (N5819, N5798);
xor XOR2 (N5820, N5812, N2556);
nand NAND3 (N5821, N5819, N2464, N3765);
nor NOR3 (N5822, N5795, N5151, N5548);
xor XOR2 (N5823, N5811, N4506);
and AND2 (N5824, N5814, N681);
buf BUF1 (N5825, N5813);
xor XOR2 (N5826, N5816, N2894);
and AND4 (N5827, N5826, N808, N4566, N997);
nand NAND4 (N5828, N5820, N3519, N11, N748);
not NOT1 (N5829, N5821);
nand NAND3 (N5830, N5828, N3439, N757);
nand NAND4 (N5831, N5818, N632, N3867, N3863);
or OR3 (N5832, N5827, N476, N4113);
or OR4 (N5833, N5824, N1829, N3482, N4819);
buf BUF1 (N5834, N5805);
or OR3 (N5835, N5829, N4606, N4889);
not NOT1 (N5836, N5830);
xor XOR2 (N5837, N5831, N1276);
and AND3 (N5838, N5834, N2079, N502);
not NOT1 (N5839, N5833);
nor NOR2 (N5840, N5832, N3779);
or OR3 (N5841, N5823, N853, N1200);
not NOT1 (N5842, N5825);
or OR4 (N5843, N5841, N667, N4369, N4613);
buf BUF1 (N5844, N5842);
not NOT1 (N5845, N5840);
nand NAND4 (N5846, N5837, N3965, N4573, N4323);
buf BUF1 (N5847, N5844);
buf BUF1 (N5848, N5822);
not NOT1 (N5849, N5847);
nand NAND2 (N5850, N5838, N1312);
buf BUF1 (N5851, N5848);
nand NAND4 (N5852, N5835, N4453, N2660, N2240);
nand NAND3 (N5853, N5852, N3634, N478);
or OR4 (N5854, N5851, N4884, N5816, N3378);
nand NAND4 (N5855, N5836, N1077, N1590, N4839);
or OR3 (N5856, N5853, N4318, N1577);
buf BUF1 (N5857, N5845);
nand NAND3 (N5858, N5854, N3865, N94);
buf BUF1 (N5859, N5849);
nand NAND4 (N5860, N5855, N145, N4743, N1823);
not NOT1 (N5861, N5850);
not NOT1 (N5862, N5846);
or OR4 (N5863, N5856, N3346, N1363, N1943);
xor XOR2 (N5864, N5860, N831);
or OR2 (N5865, N5817, N1970);
and AND2 (N5866, N5839, N4794);
xor XOR2 (N5867, N5858, N5420);
nor NOR4 (N5868, N5861, N1221, N3271, N4069);
nor NOR2 (N5869, N5868, N594);
not NOT1 (N5870, N5867);
buf BUF1 (N5871, N5857);
not NOT1 (N5872, N5871);
buf BUF1 (N5873, N5862);
nor NOR4 (N5874, N5873, N683, N3747, N4917);
nor NOR3 (N5875, N5874, N3268, N5572);
and AND2 (N5876, N5843, N4484);
or OR4 (N5877, N5876, N3332, N2280, N139);
not NOT1 (N5878, N5875);
and AND2 (N5879, N5866, N5164);
xor XOR2 (N5880, N5859, N2489);
nand NAND2 (N5881, N5879, N2036);
nor NOR3 (N5882, N5878, N2268, N5509);
or OR4 (N5883, N5869, N973, N669, N3186);
buf BUF1 (N5884, N5872);
not NOT1 (N5885, N5877);
nand NAND2 (N5886, N5865, N1246);
nand NAND4 (N5887, N5886, N627, N515, N2384);
buf BUF1 (N5888, N5887);
nor NOR4 (N5889, N5863, N5074, N4562, N354);
xor XOR2 (N5890, N5884, N5295);
not NOT1 (N5891, N5882);
nor NOR2 (N5892, N5889, N2706);
not NOT1 (N5893, N5888);
buf BUF1 (N5894, N5892);
not NOT1 (N5895, N5894);
and AND2 (N5896, N5864, N2054);
nor NOR2 (N5897, N5880, N5660);
xor XOR2 (N5898, N5893, N5558);
or OR2 (N5899, N5885, N1462);
not NOT1 (N5900, N5881);
not NOT1 (N5901, N5900);
or OR3 (N5902, N5891, N3724, N5822);
nor NOR4 (N5903, N5901, N5054, N3540, N1725);
nand NAND2 (N5904, N5870, N1369);
or OR2 (N5905, N5902, N2215);
nor NOR3 (N5906, N5904, N857, N344);
and AND3 (N5907, N5890, N3654, N3907);
nand NAND2 (N5908, N5898, N1750);
or OR3 (N5909, N5908, N5588, N4365);
nand NAND4 (N5910, N5896, N1585, N4066, N1637);
nand NAND2 (N5911, N5903, N1673);
buf BUF1 (N5912, N5907);
or OR2 (N5913, N5883, N5841);
buf BUF1 (N5914, N5913);
buf BUF1 (N5915, N5909);
and AND4 (N5916, N5915, N2687, N4782, N1110);
not NOT1 (N5917, N5906);
not NOT1 (N5918, N5917);
nand NAND2 (N5919, N5910, N5491);
nand NAND2 (N5920, N5895, N5184);
nor NOR4 (N5921, N5912, N2664, N465, N2418);
nor NOR2 (N5922, N5911, N1687);
nor NOR2 (N5923, N5921, N3228);
xor XOR2 (N5924, N5922, N1296);
nand NAND2 (N5925, N5914, N5906);
xor XOR2 (N5926, N5899, N983);
nand NAND3 (N5927, N5919, N4371, N719);
or OR2 (N5928, N5926, N2857);
and AND2 (N5929, N5920, N3116);
xor XOR2 (N5930, N5928, N1276);
not NOT1 (N5931, N5930);
nor NOR4 (N5932, N5916, N4308, N1242, N390);
xor XOR2 (N5933, N5924, N1160);
nor NOR2 (N5934, N5918, N4100);
nand NAND4 (N5935, N5933, N2319, N4741, N4451);
xor XOR2 (N5936, N5932, N5709);
buf BUF1 (N5937, N5905);
buf BUF1 (N5938, N5929);
and AND2 (N5939, N5936, N5521);
nand NAND4 (N5940, N5934, N3846, N4991, N3531);
not NOT1 (N5941, N5935);
not NOT1 (N5942, N5927);
nand NAND4 (N5943, N5941, N1278, N2423, N1390);
and AND3 (N5944, N5940, N3288, N1594);
or OR4 (N5945, N5937, N2941, N3893, N1662);
nor NOR2 (N5946, N5938, N1994);
and AND3 (N5947, N5944, N198, N1566);
nand NAND2 (N5948, N5939, N928);
nor NOR2 (N5949, N5942, N2861);
buf BUF1 (N5950, N5948);
nand NAND2 (N5951, N5945, N3217);
not NOT1 (N5952, N5947);
buf BUF1 (N5953, N5950);
buf BUF1 (N5954, N5953);
nand NAND3 (N5955, N5946, N2702, N4899);
nor NOR3 (N5956, N5954, N437, N5719);
and AND2 (N5957, N5952, N5331);
or OR2 (N5958, N5955, N5115);
nor NOR4 (N5959, N5949, N5618, N3350, N5618);
xor XOR2 (N5960, N5956, N3004);
not NOT1 (N5961, N5957);
and AND4 (N5962, N5960, N1918, N2469, N2605);
and AND2 (N5963, N5961, N5414);
and AND2 (N5964, N5958, N4053);
not NOT1 (N5965, N5962);
or OR4 (N5966, N5925, N5056, N2581, N4007);
nor NOR4 (N5967, N5966, N773, N4830, N1723);
xor XOR2 (N5968, N5897, N1408);
and AND3 (N5969, N5968, N5362, N4195);
and AND2 (N5970, N5943, N471);
nor NOR2 (N5971, N5951, N1679);
nor NOR3 (N5972, N5923, N2319, N3771);
or OR2 (N5973, N5967, N1264);
and AND3 (N5974, N5969, N4640, N4894);
not NOT1 (N5975, N5964);
and AND4 (N5976, N5965, N954, N566, N746);
nor NOR2 (N5977, N5972, N2987);
not NOT1 (N5978, N5963);
buf BUF1 (N5979, N5976);
buf BUF1 (N5980, N5959);
nand NAND3 (N5981, N5980, N4847, N1466);
or OR4 (N5982, N5974, N3288, N2451, N5783);
nor NOR3 (N5983, N5971, N4371, N2732);
and AND4 (N5984, N5931, N1320, N4112, N921);
buf BUF1 (N5985, N5982);
xor XOR2 (N5986, N5981, N1499);
nand NAND2 (N5987, N5986, N5281);
not NOT1 (N5988, N5987);
nand NAND3 (N5989, N5973, N2493, N4271);
or OR4 (N5990, N5979, N1462, N5196, N1695);
xor XOR2 (N5991, N5978, N1840);
and AND4 (N5992, N5983, N1823, N4671, N256);
and AND3 (N5993, N5989, N887, N697);
and AND3 (N5994, N5991, N274, N4759);
not NOT1 (N5995, N5990);
xor XOR2 (N5996, N5977, N3834);
buf BUF1 (N5997, N5975);
nor NOR2 (N5998, N5995, N2681);
not NOT1 (N5999, N5998);
and AND2 (N6000, N5992, N5392);
xor XOR2 (N6001, N5997, N3694);
xor XOR2 (N6002, N5984, N5468);
buf BUF1 (N6003, N5994);
nand NAND2 (N6004, N5993, N3142);
and AND3 (N6005, N6003, N4655, N5029);
buf BUF1 (N6006, N5985);
nor NOR4 (N6007, N6000, N2494, N3344, N2531);
buf BUF1 (N6008, N6002);
buf BUF1 (N6009, N5996);
and AND3 (N6010, N6001, N1652, N3333);
nor NOR3 (N6011, N6007, N1578, N2752);
nand NAND3 (N6012, N6010, N226, N1893);
nand NAND2 (N6013, N6011, N2828);
buf BUF1 (N6014, N5999);
xor XOR2 (N6015, N6013, N2145);
nand NAND4 (N6016, N6014, N2202, N4357, N5237);
not NOT1 (N6017, N6009);
not NOT1 (N6018, N6004);
xor XOR2 (N6019, N6012, N1995);
or OR4 (N6020, N6017, N3747, N3992, N4381);
and AND4 (N6021, N6016, N2650, N3834, N3938);
nor NOR4 (N6022, N6008, N5383, N3074, N1510);
or OR4 (N6023, N6021, N2082, N5124, N5569);
nor NOR2 (N6024, N6019, N5015);
buf BUF1 (N6025, N6018);
or OR3 (N6026, N6006, N4139, N1719);
buf BUF1 (N6027, N6025);
and AND2 (N6028, N6024, N3238);
nor NOR2 (N6029, N6027, N2612);
buf BUF1 (N6030, N6029);
not NOT1 (N6031, N6023);
nand NAND3 (N6032, N6020, N3076, N5950);
not NOT1 (N6033, N6030);
nand NAND4 (N6034, N6031, N4269, N1278, N649);
and AND2 (N6035, N6026, N1490);
xor XOR2 (N6036, N6022, N4721);
xor XOR2 (N6037, N5988, N5074);
nand NAND2 (N6038, N6028, N1110);
and AND4 (N6039, N6005, N4857, N477, N2489);
xor XOR2 (N6040, N6038, N4651);
nor NOR4 (N6041, N6039, N2141, N3886, N1594);
or OR2 (N6042, N6037, N405);
and AND2 (N6043, N5970, N5006);
nand NAND2 (N6044, N6036, N3567);
nand NAND4 (N6045, N6040, N5846, N214, N2507);
xor XOR2 (N6046, N6033, N5625);
not NOT1 (N6047, N6041);
nand NAND2 (N6048, N6035, N1917);
nor NOR3 (N6049, N6045, N396, N3797);
and AND4 (N6050, N6046, N256, N152, N5190);
nand NAND3 (N6051, N6047, N2038, N368);
nand NAND3 (N6052, N6032, N4006, N5374);
buf BUF1 (N6053, N6044);
or OR3 (N6054, N6043, N1796, N437);
or OR3 (N6055, N6054, N1664, N3162);
or OR3 (N6056, N6052, N5029, N3637);
not NOT1 (N6057, N6042);
or OR3 (N6058, N6057, N2368, N5151);
nand NAND4 (N6059, N6015, N2860, N3349, N4054);
xor XOR2 (N6060, N6059, N5133);
and AND2 (N6061, N6034, N5624);
and AND3 (N6062, N6049, N4478, N2125);
nand NAND4 (N6063, N6050, N3144, N1619, N4942);
xor XOR2 (N6064, N6058, N4844);
buf BUF1 (N6065, N6051);
nor NOR4 (N6066, N6060, N4112, N565, N4270);
not NOT1 (N6067, N6062);
or OR2 (N6068, N6067, N3570);
nand NAND3 (N6069, N6065, N5037, N624);
or OR2 (N6070, N6064, N2881);
nor NOR4 (N6071, N6063, N2524, N4928, N4595);
and AND4 (N6072, N6055, N4278, N1428, N4571);
nand NAND4 (N6073, N6069, N5388, N4933, N4832);
buf BUF1 (N6074, N6048);
not NOT1 (N6075, N6056);
xor XOR2 (N6076, N6075, N199);
xor XOR2 (N6077, N6070, N213);
xor XOR2 (N6078, N6068, N3221);
buf BUF1 (N6079, N6074);
or OR3 (N6080, N6077, N1086, N5388);
xor XOR2 (N6081, N6073, N3398);
and AND3 (N6082, N6072, N566, N1209);
nor NOR3 (N6083, N6081, N3927, N5271);
nor NOR4 (N6084, N6066, N4301, N4752, N2156);
not NOT1 (N6085, N6071);
and AND2 (N6086, N6076, N3494);
nand NAND2 (N6087, N6082, N3916);
buf BUF1 (N6088, N6080);
nor NOR2 (N6089, N6088, N4832);
or OR2 (N6090, N6053, N4397);
not NOT1 (N6091, N6078);
xor XOR2 (N6092, N6087, N844);
or OR3 (N6093, N6084, N5827, N5994);
nand NAND3 (N6094, N6085, N1923, N3995);
and AND2 (N6095, N6094, N3776);
nand NAND3 (N6096, N6091, N3448, N5593);
nor NOR2 (N6097, N6096, N564);
xor XOR2 (N6098, N6093, N3725);
buf BUF1 (N6099, N6089);
not NOT1 (N6100, N6098);
xor XOR2 (N6101, N6061, N4554);
nor NOR3 (N6102, N6101, N3624, N2334);
nand NAND3 (N6103, N6079, N3486, N2176);
or OR4 (N6104, N6090, N4245, N4588, N2739);
xor XOR2 (N6105, N6086, N2315);
or OR2 (N6106, N6099, N2347);
nand NAND2 (N6107, N6103, N3464);
nand NAND3 (N6108, N6104, N59, N4219);
nand NAND2 (N6109, N6105, N1431);
nor NOR4 (N6110, N6100, N4865, N1593, N349);
nand NAND3 (N6111, N6109, N2938, N109);
nand NAND4 (N6112, N6110, N5501, N2004, N1895);
or OR3 (N6113, N6107, N2835, N5200);
and AND4 (N6114, N6092, N3083, N1263, N5028);
nor NOR2 (N6115, N6113, N2546);
and AND4 (N6116, N6114, N4360, N2311, N5673);
and AND3 (N6117, N6116, N847, N4245);
xor XOR2 (N6118, N6097, N5234);
nand NAND2 (N6119, N6115, N5025);
nand NAND2 (N6120, N6108, N4310);
not NOT1 (N6121, N6118);
or OR2 (N6122, N6111, N1213);
or OR4 (N6123, N6106, N5255, N5558, N5252);
not NOT1 (N6124, N6123);
not NOT1 (N6125, N6119);
nand NAND2 (N6126, N6095, N1627);
nand NAND4 (N6127, N6120, N1210, N6112, N1778);
xor XOR2 (N6128, N4797, N5374);
buf BUF1 (N6129, N6125);
or OR2 (N6130, N6128, N554);
and AND4 (N6131, N6130, N3262, N5176, N554);
nand NAND4 (N6132, N6131, N1975, N5606, N1205);
and AND4 (N6133, N6129, N4730, N4733, N1836);
xor XOR2 (N6134, N6133, N5958);
xor XOR2 (N6135, N6126, N5058);
not NOT1 (N6136, N6135);
nor NOR3 (N6137, N6136, N652, N734);
or OR4 (N6138, N6122, N5357, N3012, N4143);
or OR2 (N6139, N6132, N5716);
buf BUF1 (N6140, N6138);
or OR3 (N6141, N6134, N2561, N5803);
buf BUF1 (N6142, N6141);
or OR3 (N6143, N6102, N6086, N2525);
buf BUF1 (N6144, N6137);
nor NOR4 (N6145, N6143, N5992, N5903, N4464);
or OR2 (N6146, N6139, N1633);
and AND3 (N6147, N6146, N3164, N5296);
nor NOR4 (N6148, N6127, N2371, N3111, N3683);
or OR2 (N6149, N6147, N4619);
nand NAND3 (N6150, N6148, N2638, N1377);
not NOT1 (N6151, N6145);
nand NAND4 (N6152, N6150, N1331, N3961, N5943);
nand NAND2 (N6153, N6142, N2929);
nand NAND4 (N6154, N6117, N4235, N1289, N5587);
nor NOR3 (N6155, N6124, N6056, N4081);
nor NOR2 (N6156, N6155, N2105);
nor NOR4 (N6157, N6149, N1955, N852, N5814);
nand NAND4 (N6158, N6140, N4015, N4911, N5532);
xor XOR2 (N6159, N6083, N6119);
and AND4 (N6160, N6154, N2302, N536, N1676);
buf BUF1 (N6161, N6157);
nand NAND4 (N6162, N6156, N455, N2448, N4705);
xor XOR2 (N6163, N6160, N2570);
and AND2 (N6164, N6151, N1876);
nand NAND4 (N6165, N6164, N3261, N5497, N2211);
and AND2 (N6166, N6161, N6148);
and AND3 (N6167, N6163, N1416, N3105);
nor NOR4 (N6168, N6167, N1414, N3637, N1548);
nand NAND2 (N6169, N6158, N5706);
xor XOR2 (N6170, N6121, N5732);
buf BUF1 (N6171, N6144);
not NOT1 (N6172, N6152);
xor XOR2 (N6173, N6166, N4785);
xor XOR2 (N6174, N6171, N4690);
not NOT1 (N6175, N6168);
buf BUF1 (N6176, N6153);
nor NOR4 (N6177, N6174, N3018, N2262, N4297);
buf BUF1 (N6178, N6173);
or OR2 (N6179, N6162, N4968);
nor NOR2 (N6180, N6177, N410);
nor NOR2 (N6181, N6179, N274);
xor XOR2 (N6182, N6175, N3268);
xor XOR2 (N6183, N6165, N2288);
xor XOR2 (N6184, N6169, N2746);
buf BUF1 (N6185, N6176);
and AND2 (N6186, N6159, N5057);
xor XOR2 (N6187, N6172, N2698);
buf BUF1 (N6188, N6180);
buf BUF1 (N6189, N6185);
or OR4 (N6190, N6187, N2053, N425, N5880);
buf BUF1 (N6191, N6170);
not NOT1 (N6192, N6191);
nor NOR2 (N6193, N6178, N223);
buf BUF1 (N6194, N6183);
or OR2 (N6195, N6189, N5557);
nand NAND3 (N6196, N6181, N5194, N5975);
or OR4 (N6197, N6192, N3717, N5225, N5255);
or OR3 (N6198, N6184, N5192, N913);
or OR4 (N6199, N6193, N3977, N2736, N4140);
xor XOR2 (N6200, N6199, N1565);
or OR2 (N6201, N6200, N607);
nor NOR3 (N6202, N6194, N2536, N2909);
nand NAND4 (N6203, N6182, N1060, N1854, N5250);
nand NAND4 (N6204, N6198, N2459, N3102, N3206);
and AND3 (N6205, N6203, N5876, N5626);
xor XOR2 (N6206, N6197, N2208);
not NOT1 (N6207, N6190);
buf BUF1 (N6208, N6196);
not NOT1 (N6209, N6195);
and AND3 (N6210, N6206, N1434, N2806);
not NOT1 (N6211, N6188);
xor XOR2 (N6212, N6211, N3995);
buf BUF1 (N6213, N6207);
xor XOR2 (N6214, N6186, N5331);
not NOT1 (N6215, N6213);
nor NOR2 (N6216, N6208, N1531);
not NOT1 (N6217, N6212);
nor NOR3 (N6218, N6215, N510, N3813);
xor XOR2 (N6219, N6210, N899);
or OR3 (N6220, N6209, N44, N3950);
buf BUF1 (N6221, N6204);
xor XOR2 (N6222, N6221, N4363);
nand NAND4 (N6223, N6217, N2058, N2629, N5681);
not NOT1 (N6224, N6216);
xor XOR2 (N6225, N6202, N1187);
and AND2 (N6226, N6225, N3706);
nand NAND2 (N6227, N6220, N3561);
and AND4 (N6228, N6205, N4334, N2512, N4056);
and AND4 (N6229, N6223, N16, N2523, N526);
nor NOR3 (N6230, N6219, N4871, N2290);
xor XOR2 (N6231, N6218, N4487);
nor NOR3 (N6232, N6224, N376, N6066);
or OR4 (N6233, N6229, N5530, N292, N4446);
or OR4 (N6234, N6226, N4521, N502, N6103);
and AND3 (N6235, N6232, N5860, N5164);
or OR2 (N6236, N6222, N2084);
or OR2 (N6237, N6233, N4203);
nand NAND4 (N6238, N6231, N4112, N102, N3827);
and AND3 (N6239, N6237, N495, N494);
nor NOR3 (N6240, N6239, N3932, N2785);
and AND4 (N6241, N6238, N2624, N3098, N824);
and AND4 (N6242, N6201, N707, N432, N5954);
not NOT1 (N6243, N6242);
xor XOR2 (N6244, N6227, N1686);
buf BUF1 (N6245, N6235);
not NOT1 (N6246, N6234);
xor XOR2 (N6247, N6230, N3780);
nand NAND4 (N6248, N6245, N3701, N6115, N1947);
not NOT1 (N6249, N6240);
nor NOR3 (N6250, N6249, N4318, N940);
buf BUF1 (N6251, N6214);
nor NOR2 (N6252, N6246, N87);
or OR2 (N6253, N6243, N3396);
nor NOR4 (N6254, N6253, N4717, N5675, N2052);
nor NOR2 (N6255, N6241, N3729);
buf BUF1 (N6256, N6247);
not NOT1 (N6257, N6254);
and AND3 (N6258, N6255, N1648, N4688);
nand NAND2 (N6259, N6258, N4032);
not NOT1 (N6260, N6251);
xor XOR2 (N6261, N6259, N993);
and AND4 (N6262, N6252, N5417, N6130, N2149);
or OR2 (N6263, N6236, N42);
buf BUF1 (N6264, N6257);
not NOT1 (N6265, N6261);
nor NOR3 (N6266, N6248, N5500, N659);
and AND2 (N6267, N6266, N5247);
and AND3 (N6268, N6256, N458, N5804);
xor XOR2 (N6269, N6264, N3415);
buf BUF1 (N6270, N6263);
not NOT1 (N6271, N6270);
and AND2 (N6272, N6267, N271);
nor NOR3 (N6273, N6260, N1677, N5308);
not NOT1 (N6274, N6265);
xor XOR2 (N6275, N6273, N5876);
not NOT1 (N6276, N6274);
nor NOR3 (N6277, N6244, N3543, N1363);
or OR2 (N6278, N6271, N5804);
or OR4 (N6279, N6275, N5627, N4109, N5812);
nor NOR4 (N6280, N6276, N4656, N2393, N4365);
buf BUF1 (N6281, N6228);
and AND3 (N6282, N6280, N236, N5202);
not NOT1 (N6283, N6279);
xor XOR2 (N6284, N6269, N2771);
xor XOR2 (N6285, N6282, N4237);
and AND2 (N6286, N6250, N2999);
xor XOR2 (N6287, N6285, N2893);
or OR2 (N6288, N6277, N5697);
xor XOR2 (N6289, N6286, N4680);
nor NOR3 (N6290, N6262, N3250, N4138);
and AND2 (N6291, N6283, N4707);
nor NOR3 (N6292, N6291, N3297, N4530);
nor NOR4 (N6293, N6287, N1718, N2685, N1906);
and AND2 (N6294, N6289, N851);
not NOT1 (N6295, N6281);
nor NOR4 (N6296, N6288, N4394, N2079, N4589);
nand NAND4 (N6297, N6284, N2606, N1087, N6204);
buf BUF1 (N6298, N6278);
nor NOR3 (N6299, N6292, N1646, N5515);
not NOT1 (N6300, N6293);
and AND3 (N6301, N6272, N3210, N1417);
and AND3 (N6302, N6299, N1672, N5300);
buf BUF1 (N6303, N6302);
not NOT1 (N6304, N6295);
and AND3 (N6305, N6298, N3570, N5217);
nor NOR4 (N6306, N6304, N222, N6155, N1308);
nor NOR2 (N6307, N6300, N786);
nor NOR3 (N6308, N6307, N1119, N537);
and AND4 (N6309, N6305, N972, N2506, N1825);
not NOT1 (N6310, N6308);
or OR2 (N6311, N6296, N5444);
and AND2 (N6312, N6294, N835);
not NOT1 (N6313, N6290);
and AND2 (N6314, N6313, N1436);
and AND3 (N6315, N6303, N6243, N5649);
not NOT1 (N6316, N6306);
nand NAND3 (N6317, N6309, N5068, N3378);
not NOT1 (N6318, N6315);
buf BUF1 (N6319, N6311);
buf BUF1 (N6320, N6319);
xor XOR2 (N6321, N6320, N5980);
buf BUF1 (N6322, N6318);
buf BUF1 (N6323, N6310);
buf BUF1 (N6324, N6317);
nor NOR3 (N6325, N6321, N1799, N3195);
nand NAND4 (N6326, N6323, N3794, N1806, N432);
not NOT1 (N6327, N6268);
and AND2 (N6328, N6325, N2908);
not NOT1 (N6329, N6328);
nor NOR3 (N6330, N6301, N3392, N5290);
nand NAND2 (N6331, N6314, N5511);
not NOT1 (N6332, N6331);
not NOT1 (N6333, N6327);
or OR4 (N6334, N6330, N6278, N4763, N4672);
xor XOR2 (N6335, N6333, N194);
xor XOR2 (N6336, N6326, N4013);
buf BUF1 (N6337, N6329);
buf BUF1 (N6338, N6337);
not NOT1 (N6339, N6316);
and AND3 (N6340, N6297, N4581, N1982);
xor XOR2 (N6341, N6324, N3947);
buf BUF1 (N6342, N6338);
buf BUF1 (N6343, N6334);
not NOT1 (N6344, N6341);
and AND4 (N6345, N6342, N5262, N4597, N968);
nor NOR2 (N6346, N6343, N1247);
xor XOR2 (N6347, N6339, N327);
and AND4 (N6348, N6345, N1363, N6318, N4133);
or OR2 (N6349, N6312, N939);
or OR3 (N6350, N6340, N6097, N4306);
xor XOR2 (N6351, N6346, N1673);
or OR2 (N6352, N6348, N5719);
xor XOR2 (N6353, N6336, N3662);
nand NAND2 (N6354, N6352, N3951);
nand NAND2 (N6355, N6351, N2884);
nand NAND4 (N6356, N6322, N5856, N1687, N4482);
nand NAND2 (N6357, N6354, N4055);
and AND4 (N6358, N6332, N1413, N4546, N1001);
and AND4 (N6359, N6347, N2105, N1269, N4435);
nor NOR4 (N6360, N6335, N2922, N2623, N1568);
xor XOR2 (N6361, N6356, N5568);
and AND3 (N6362, N6361, N1630, N5919);
xor XOR2 (N6363, N6358, N6194);
nand NAND3 (N6364, N6349, N2117, N4726);
buf BUF1 (N6365, N6362);
nand NAND4 (N6366, N6363, N6308, N4304, N3954);
nor NOR2 (N6367, N6366, N4395);
nor NOR2 (N6368, N6355, N496);
nand NAND4 (N6369, N6357, N3072, N5153, N3199);
nor NOR2 (N6370, N6365, N5217);
nor NOR4 (N6371, N6353, N5188, N5491, N2116);
xor XOR2 (N6372, N6350, N4725);
nor NOR4 (N6373, N6344, N5269, N702, N3898);
and AND3 (N6374, N6369, N3497, N3965);
and AND3 (N6375, N6360, N1727, N2892);
nor NOR4 (N6376, N6371, N370, N4648, N1188);
nand NAND4 (N6377, N6367, N1416, N801, N5267);
and AND4 (N6378, N6373, N4175, N6119, N3073);
buf BUF1 (N6379, N6376);
xor XOR2 (N6380, N6374, N2187);
buf BUF1 (N6381, N6359);
and AND2 (N6382, N6364, N1308);
or OR2 (N6383, N6368, N6071);
nand NAND2 (N6384, N6375, N5169);
or OR3 (N6385, N6377, N4996, N1551);
or OR3 (N6386, N6380, N81, N266);
or OR4 (N6387, N6383, N5942, N4642, N2008);
not NOT1 (N6388, N6382);
xor XOR2 (N6389, N6384, N4969);
and AND2 (N6390, N6386, N105);
not NOT1 (N6391, N6372);
nand NAND2 (N6392, N6370, N243);
nand NAND3 (N6393, N6389, N2618, N4997);
or OR3 (N6394, N6379, N508, N1202);
not NOT1 (N6395, N6394);
and AND3 (N6396, N6390, N5579, N2063);
and AND3 (N6397, N6391, N269, N5671);
or OR4 (N6398, N6381, N5390, N2625, N6217);
nor NOR4 (N6399, N6393, N3471, N6352, N5412);
and AND3 (N6400, N6398, N5709, N1484);
not NOT1 (N6401, N6385);
buf BUF1 (N6402, N6387);
not NOT1 (N6403, N6400);
or OR4 (N6404, N6388, N4562, N4864, N5155);
xor XOR2 (N6405, N6401, N2810);
or OR4 (N6406, N6404, N4949, N4424, N4705);
and AND4 (N6407, N6402, N5386, N1997, N300);
buf BUF1 (N6408, N6406);
nor NOR2 (N6409, N6403, N3774);
nor NOR2 (N6410, N6405, N1806);
nor NOR2 (N6411, N6409, N572);
nand NAND3 (N6412, N6408, N2273, N890);
and AND3 (N6413, N6378, N2455, N5696);
buf BUF1 (N6414, N6399);
nor NOR2 (N6415, N6397, N4462);
and AND4 (N6416, N6412, N30, N6065, N6175);
and AND2 (N6417, N6411, N806);
buf BUF1 (N6418, N6415);
or OR2 (N6419, N6392, N6008);
nand NAND4 (N6420, N6416, N2562, N1224, N320);
or OR3 (N6421, N6413, N1988, N3421);
not NOT1 (N6422, N6421);
not NOT1 (N6423, N6418);
or OR3 (N6424, N6420, N2031, N5313);
or OR4 (N6425, N6422, N2440, N4740, N3833);
and AND2 (N6426, N6396, N654);
buf BUF1 (N6427, N6424);
and AND4 (N6428, N6426, N4974, N5816, N3792);
and AND4 (N6429, N6419, N255, N5951, N1352);
not NOT1 (N6430, N6425);
nor NOR2 (N6431, N6414, N1202);
not NOT1 (N6432, N6431);
and AND4 (N6433, N6410, N648, N5280, N4446);
nor NOR2 (N6434, N6407, N3151);
nor NOR2 (N6435, N6417, N6259);
or OR4 (N6436, N6435, N4711, N6359, N947);
not NOT1 (N6437, N6436);
buf BUF1 (N6438, N6429);
xor XOR2 (N6439, N6438, N5463);
buf BUF1 (N6440, N6432);
and AND4 (N6441, N6423, N5091, N4104, N1571);
and AND2 (N6442, N6440, N2365);
not NOT1 (N6443, N6428);
or OR3 (N6444, N6434, N4060, N1500);
xor XOR2 (N6445, N6442, N2778);
or OR2 (N6446, N6444, N5521);
and AND2 (N6447, N6443, N3014);
and AND2 (N6448, N6439, N5181);
xor XOR2 (N6449, N6430, N2098);
nand NAND4 (N6450, N6448, N3757, N5525, N2957);
xor XOR2 (N6451, N6445, N3615);
nor NOR4 (N6452, N6441, N4409, N4186, N1359);
and AND3 (N6453, N6452, N83, N4204);
and AND3 (N6454, N6450, N3626, N760);
xor XOR2 (N6455, N6433, N2822);
not NOT1 (N6456, N6395);
nor NOR3 (N6457, N6446, N1687, N3167);
buf BUF1 (N6458, N6454);
and AND4 (N6459, N6447, N1379, N6230, N3471);
nor NOR2 (N6460, N6427, N2654);
and AND2 (N6461, N6459, N601);
and AND2 (N6462, N6451, N170);
nand NAND3 (N6463, N6455, N4845, N2839);
nor NOR2 (N6464, N6457, N3278);
nand NAND2 (N6465, N6462, N6102);
not NOT1 (N6466, N6464);
xor XOR2 (N6467, N6465, N6248);
buf BUF1 (N6468, N6461);
nor NOR2 (N6469, N6467, N3091);
nand NAND2 (N6470, N6449, N5315);
buf BUF1 (N6471, N6466);
nor NOR2 (N6472, N6453, N5325);
and AND3 (N6473, N6472, N750, N3995);
buf BUF1 (N6474, N6437);
nor NOR2 (N6475, N6460, N3491);
buf BUF1 (N6476, N6471);
or OR4 (N6477, N6475, N1662, N762, N5539);
xor XOR2 (N6478, N6470, N4062);
buf BUF1 (N6479, N6474);
nor NOR4 (N6480, N6477, N2759, N804, N3764);
and AND3 (N6481, N6468, N3580, N630);
buf BUF1 (N6482, N6469);
and AND3 (N6483, N6481, N4435, N6461);
buf BUF1 (N6484, N6483);
and AND4 (N6485, N6456, N330, N1114, N3312);
or OR2 (N6486, N6479, N710);
or OR2 (N6487, N6486, N5425);
xor XOR2 (N6488, N6478, N6152);
not NOT1 (N6489, N6485);
not NOT1 (N6490, N6458);
buf BUF1 (N6491, N6482);
not NOT1 (N6492, N6473);
and AND3 (N6493, N6488, N6332, N1271);
xor XOR2 (N6494, N6463, N5185);
xor XOR2 (N6495, N6491, N3881);
xor XOR2 (N6496, N6476, N411);
nand NAND2 (N6497, N6487, N5816);
or OR4 (N6498, N6496, N2568, N6086, N2361);
buf BUF1 (N6499, N6493);
buf BUF1 (N6500, N6494);
buf BUF1 (N6501, N6484);
nand NAND3 (N6502, N6490, N2948, N347);
nand NAND2 (N6503, N6489, N3880);
not NOT1 (N6504, N6499);
or OR4 (N6505, N6504, N5139, N362, N1202);
or OR4 (N6506, N6502, N6157, N1588, N4957);
nor NOR2 (N6507, N6501, N2936);
nor NOR4 (N6508, N6495, N6402, N2329, N240);
nand NAND3 (N6509, N6507, N5943, N2690);
not NOT1 (N6510, N6492);
buf BUF1 (N6511, N6509);
nand NAND3 (N6512, N6505, N3932, N225);
and AND4 (N6513, N6500, N4774, N4864, N4809);
and AND3 (N6514, N6511, N3846, N831);
buf BUF1 (N6515, N6497);
buf BUF1 (N6516, N6503);
and AND4 (N6517, N6480, N2821, N2829, N2318);
or OR3 (N6518, N6498, N5884, N2422);
not NOT1 (N6519, N6510);
nor NOR3 (N6520, N6518, N6032, N490);
buf BUF1 (N6521, N6513);
not NOT1 (N6522, N6517);
nand NAND4 (N6523, N6522, N2011, N5075, N4183);
nand NAND3 (N6524, N6523, N5405, N1993);
or OR4 (N6525, N6515, N2133, N47, N4549);
or OR2 (N6526, N6520, N5517);
buf BUF1 (N6527, N6525);
nand NAND2 (N6528, N6514, N5467);
nand NAND4 (N6529, N6527, N196, N522, N4530);
or OR4 (N6530, N6516, N1825, N4482, N5091);
or OR4 (N6531, N6508, N6510, N6188, N2574);
nor NOR4 (N6532, N6531, N4342, N4801, N4614);
buf BUF1 (N6533, N6521);
buf BUF1 (N6534, N6529);
or OR2 (N6535, N6524, N562);
not NOT1 (N6536, N6526);
nand NAND4 (N6537, N6512, N3243, N869, N5711);
nor NOR4 (N6538, N6528, N5435, N3025, N2652);
buf BUF1 (N6539, N6530);
xor XOR2 (N6540, N6533, N466);
nand NAND2 (N6541, N6519, N5910);
not NOT1 (N6542, N6537);
not NOT1 (N6543, N6538);
nor NOR3 (N6544, N6539, N2783, N3444);
xor XOR2 (N6545, N6532, N4863);
buf BUF1 (N6546, N6535);
xor XOR2 (N6547, N6544, N3997);
nand NAND4 (N6548, N6540, N4421, N3875, N5553);
xor XOR2 (N6549, N6541, N3737);
or OR3 (N6550, N6506, N4422, N4835);
not NOT1 (N6551, N6546);
nor NOR2 (N6552, N6542, N3000);
nor NOR2 (N6553, N6534, N2533);
xor XOR2 (N6554, N6553, N2915);
buf BUF1 (N6555, N6536);
buf BUF1 (N6556, N6549);
buf BUF1 (N6557, N6548);
and AND2 (N6558, N6556, N2919);
xor XOR2 (N6559, N6554, N3499);
or OR3 (N6560, N6545, N4740, N625);
or OR4 (N6561, N6559, N6258, N4106, N3976);
or OR3 (N6562, N6555, N4470, N6474);
buf BUF1 (N6563, N6560);
nor NOR4 (N6564, N6547, N4311, N3871, N852);
not NOT1 (N6565, N6550);
and AND3 (N6566, N6564, N3892, N3601);
or OR3 (N6567, N6565, N5196, N5528);
buf BUF1 (N6568, N6562);
xor XOR2 (N6569, N6566, N6385);
or OR4 (N6570, N6558, N2175, N1056, N5114);
buf BUF1 (N6571, N6568);
and AND3 (N6572, N6551, N5364, N4652);
xor XOR2 (N6573, N6561, N4719);
nor NOR2 (N6574, N6572, N3136);
nand NAND2 (N6575, N6571, N630);
nand NAND3 (N6576, N6563, N5286, N6430);
buf BUF1 (N6577, N6574);
nand NAND2 (N6578, N6575, N4772);
nand NAND3 (N6579, N6573, N5695, N3807);
nor NOR2 (N6580, N6557, N4447);
not NOT1 (N6581, N6576);
or OR4 (N6582, N6579, N5484, N3169, N1241);
and AND2 (N6583, N6552, N5402);
not NOT1 (N6584, N6569);
nand NAND3 (N6585, N6543, N6083, N2053);
and AND2 (N6586, N6581, N1015);
xor XOR2 (N6587, N6580, N3880);
or OR4 (N6588, N6584, N4235, N5161, N1302);
buf BUF1 (N6589, N6570);
xor XOR2 (N6590, N6578, N1073);
and AND4 (N6591, N6585, N5217, N4640, N156);
xor XOR2 (N6592, N6587, N1812);
not NOT1 (N6593, N6583);
nand NAND3 (N6594, N6591, N6364, N5396);
xor XOR2 (N6595, N6588, N1811);
xor XOR2 (N6596, N6593, N98);
nor NOR3 (N6597, N6594, N324, N1931);
nor NOR2 (N6598, N6586, N5875);
or OR2 (N6599, N6598, N3324);
nor NOR2 (N6600, N6577, N695);
or OR2 (N6601, N6600, N2506);
not NOT1 (N6602, N6589);
or OR4 (N6603, N6597, N4850, N1178, N4243);
nor NOR3 (N6604, N6582, N4931, N1047);
nor NOR3 (N6605, N6567, N3728, N4775);
not NOT1 (N6606, N6590);
or OR4 (N6607, N6592, N379, N896, N6449);
buf BUF1 (N6608, N6605);
buf BUF1 (N6609, N6607);
and AND3 (N6610, N6603, N5072, N1877);
buf BUF1 (N6611, N6601);
buf BUF1 (N6612, N6609);
nor NOR3 (N6613, N6604, N1869, N3964);
or OR2 (N6614, N6613, N3162);
buf BUF1 (N6615, N6606);
not NOT1 (N6616, N6614);
buf BUF1 (N6617, N6610);
buf BUF1 (N6618, N6595);
buf BUF1 (N6619, N6608);
nand NAND3 (N6620, N6616, N3100, N6171);
buf BUF1 (N6621, N6611);
xor XOR2 (N6622, N6615, N3359);
not NOT1 (N6623, N6602);
nand NAND2 (N6624, N6618, N6182);
and AND2 (N6625, N6599, N722);
buf BUF1 (N6626, N6619);
and AND3 (N6627, N6621, N2714, N6228);
xor XOR2 (N6628, N6627, N3531);
nor NOR3 (N6629, N6596, N5853, N3159);
not NOT1 (N6630, N6628);
xor XOR2 (N6631, N6622, N1499);
and AND3 (N6632, N6620, N425, N2530);
nand NAND4 (N6633, N6629, N6310, N6126, N5341);
and AND2 (N6634, N6625, N4813);
buf BUF1 (N6635, N6626);
or OR3 (N6636, N6624, N4639, N1253);
xor XOR2 (N6637, N6630, N2411);
or OR4 (N6638, N6636, N5439, N518, N6447);
xor XOR2 (N6639, N6633, N1131);
and AND2 (N6640, N6635, N4578);
xor XOR2 (N6641, N6637, N3201);
or OR4 (N6642, N6641, N3610, N5582, N614);
not NOT1 (N6643, N6639);
nand NAND2 (N6644, N6632, N4468);
not NOT1 (N6645, N6643);
or OR3 (N6646, N6623, N1795, N1842);
not NOT1 (N6647, N6642);
not NOT1 (N6648, N6631);
xor XOR2 (N6649, N6634, N3355);
not NOT1 (N6650, N6646);
or OR2 (N6651, N6638, N6367);
or OR2 (N6652, N6617, N4248);
not NOT1 (N6653, N6650);
and AND4 (N6654, N6653, N3117, N6598, N1109);
not NOT1 (N6655, N6648);
nand NAND4 (N6656, N6612, N1567, N1908, N4273);
xor XOR2 (N6657, N6649, N2601);
or OR4 (N6658, N6657, N3726, N3137, N6299);
xor XOR2 (N6659, N6645, N2227);
and AND4 (N6660, N6658, N5890, N5468, N643);
and AND3 (N6661, N6644, N5214, N2431);
and AND2 (N6662, N6656, N2165);
nor NOR2 (N6663, N6654, N5296);
not NOT1 (N6664, N6655);
nor NOR3 (N6665, N6647, N6507, N454);
not NOT1 (N6666, N6661);
nand NAND2 (N6667, N6659, N1474);
or OR4 (N6668, N6664, N5470, N2387, N806);
xor XOR2 (N6669, N6640, N5326);
not NOT1 (N6670, N6652);
or OR4 (N6671, N6662, N994, N6630, N144);
buf BUF1 (N6672, N6667);
xor XOR2 (N6673, N6668, N2362);
nand NAND3 (N6674, N6651, N4890, N2457);
not NOT1 (N6675, N6674);
not NOT1 (N6676, N6669);
xor XOR2 (N6677, N6673, N387);
or OR4 (N6678, N6675, N3145, N3048, N1697);
nand NAND2 (N6679, N6671, N2202);
nor NOR3 (N6680, N6676, N252, N2553);
and AND3 (N6681, N6663, N4224, N4071);
nor NOR4 (N6682, N6672, N3655, N3600, N2035);
buf BUF1 (N6683, N6678);
and AND4 (N6684, N6683, N3888, N5646, N788);
and AND3 (N6685, N6665, N5511, N2150);
nor NOR3 (N6686, N6681, N1039, N2651);
and AND2 (N6687, N6684, N5821);
xor XOR2 (N6688, N6666, N2579);
or OR4 (N6689, N6670, N779, N3852, N1076);
and AND4 (N6690, N6660, N2197, N4488, N6380);
nand NAND2 (N6691, N6687, N5657);
buf BUF1 (N6692, N6688);
xor XOR2 (N6693, N6685, N3490);
nand NAND4 (N6694, N6692, N6044, N2129, N5583);
buf BUF1 (N6695, N6689);
nand NAND3 (N6696, N6679, N3537, N1956);
buf BUF1 (N6697, N6680);
and AND3 (N6698, N6693, N5150, N3427);
nand NAND4 (N6699, N6698, N4642, N4287, N5578);
xor XOR2 (N6700, N6690, N2450);
buf BUF1 (N6701, N6700);
buf BUF1 (N6702, N6701);
buf BUF1 (N6703, N6677);
and AND3 (N6704, N6682, N3637, N1528);
nor NOR4 (N6705, N6703, N3205, N354, N1324);
xor XOR2 (N6706, N6699, N4318);
or OR2 (N6707, N6697, N2780);
not NOT1 (N6708, N6704);
nand NAND3 (N6709, N6694, N6335, N2670);
or OR3 (N6710, N6708, N4845, N4950);
nand NAND2 (N6711, N6710, N4933);
not NOT1 (N6712, N6686);
not NOT1 (N6713, N6712);
or OR2 (N6714, N6711, N1077);
and AND4 (N6715, N6713, N4544, N4024, N233);
and AND3 (N6716, N6695, N5191, N370);
nand NAND3 (N6717, N6709, N6664, N5137);
or OR4 (N6718, N6714, N2016, N6540, N6074);
nor NOR3 (N6719, N6696, N182, N480);
not NOT1 (N6720, N6719);
or OR2 (N6721, N6717, N3913);
or OR4 (N6722, N6691, N2921, N811, N96);
nor NOR3 (N6723, N6716, N5349, N2743);
and AND4 (N6724, N6722, N510, N6677, N4184);
nand NAND4 (N6725, N6715, N1745, N1846, N2351);
xor XOR2 (N6726, N6707, N4759);
nor NOR3 (N6727, N6706, N5249, N986);
buf BUF1 (N6728, N6725);
not NOT1 (N6729, N6705);
nor NOR4 (N6730, N6728, N2789, N6367, N6236);
nor NOR3 (N6731, N6721, N6051, N1670);
nor NOR3 (N6732, N6724, N5920, N6257);
xor XOR2 (N6733, N6720, N2302);
xor XOR2 (N6734, N6729, N307);
and AND3 (N6735, N6727, N109, N4204);
not NOT1 (N6736, N6734);
and AND2 (N6737, N6731, N3462);
nor NOR2 (N6738, N6702, N4354);
nand NAND4 (N6739, N6737, N6458, N2093, N1688);
xor XOR2 (N6740, N6730, N3661);
nand NAND2 (N6741, N6732, N71);
xor XOR2 (N6742, N6733, N3872);
buf BUF1 (N6743, N6739);
nor NOR2 (N6744, N6736, N4156);
nand NAND4 (N6745, N6718, N1320, N4807, N1947);
nand NAND3 (N6746, N6743, N1091, N1102);
nor NOR4 (N6747, N6735, N4437, N4475, N332);
buf BUF1 (N6748, N6738);
nand NAND3 (N6749, N6740, N2278, N5771);
nand NAND3 (N6750, N6742, N3381, N4390);
nand NAND3 (N6751, N6723, N1982, N5763);
nor NOR3 (N6752, N6750, N5344, N4363);
nor NOR4 (N6753, N6749, N3227, N831, N244);
or OR4 (N6754, N6745, N1903, N4697, N2771);
xor XOR2 (N6755, N6741, N2840);
nor NOR2 (N6756, N6744, N4816);
nor NOR4 (N6757, N6748, N1330, N3483, N969);
not NOT1 (N6758, N6756);
nand NAND2 (N6759, N6758, N2267);
nor NOR2 (N6760, N6755, N5339);
and AND4 (N6761, N6751, N5185, N2544, N5930);
nor NOR4 (N6762, N6746, N3207, N6743, N38);
nor NOR3 (N6763, N6761, N145, N2338);
xor XOR2 (N6764, N6726, N3646);
nor NOR2 (N6765, N6764, N2845);
and AND3 (N6766, N6752, N836, N2638);
buf BUF1 (N6767, N6766);
nor NOR2 (N6768, N6754, N2917);
or OR2 (N6769, N6763, N6408);
not NOT1 (N6770, N6769);
not NOT1 (N6771, N6759);
buf BUF1 (N6772, N6762);
or OR3 (N6773, N6753, N1840, N471);
buf BUF1 (N6774, N6767);
or OR2 (N6775, N6774, N5966);
or OR4 (N6776, N6765, N4520, N4993, N2769);
xor XOR2 (N6777, N6747, N2343);
xor XOR2 (N6778, N6772, N404);
not NOT1 (N6779, N6776);
and AND3 (N6780, N6779, N1981, N3664);
buf BUF1 (N6781, N6771);
or OR3 (N6782, N6757, N5535, N2757);
xor XOR2 (N6783, N6768, N2139);
and AND3 (N6784, N6777, N3905, N5541);
or OR2 (N6785, N6781, N5988);
and AND4 (N6786, N6760, N166, N5106, N3274);
not NOT1 (N6787, N6775);
nand NAND2 (N6788, N6782, N1081);
nor NOR2 (N6789, N6773, N97);
nor NOR3 (N6790, N6789, N4764, N4290);
buf BUF1 (N6791, N6788);
not NOT1 (N6792, N6790);
buf BUF1 (N6793, N6780);
or OR3 (N6794, N6784, N2797, N584);
not NOT1 (N6795, N6785);
not NOT1 (N6796, N6794);
nor NOR2 (N6797, N6770, N2659);
buf BUF1 (N6798, N6791);
and AND3 (N6799, N6786, N1910, N5310);
nor NOR3 (N6800, N6797, N1403, N2626);
or OR4 (N6801, N6793, N6648, N1639, N2711);
not NOT1 (N6802, N6796);
buf BUF1 (N6803, N6783);
not NOT1 (N6804, N6802);
nand NAND4 (N6805, N6795, N5312, N5948, N6309);
buf BUF1 (N6806, N6798);
not NOT1 (N6807, N6799);
nand NAND2 (N6808, N6801, N2381);
and AND4 (N6809, N6803, N1066, N6269, N734);
and AND4 (N6810, N6800, N2867, N3469, N3857);
nand NAND2 (N6811, N6805, N737);
nor NOR3 (N6812, N6804, N2094, N4229);
buf BUF1 (N6813, N6810);
nand NAND3 (N6814, N6778, N3441, N3024);
nor NOR2 (N6815, N6814, N2710);
buf BUF1 (N6816, N6812);
not NOT1 (N6817, N6808);
buf BUF1 (N6818, N6809);
or OR4 (N6819, N6811, N726, N6335, N1311);
nand NAND2 (N6820, N6813, N157);
or OR3 (N6821, N6806, N2681, N6067);
nor NOR4 (N6822, N6821, N4829, N4657, N6353);
not NOT1 (N6823, N6787);
nand NAND3 (N6824, N6815, N372, N5072);
nand NAND4 (N6825, N6792, N2615, N3367, N6564);
not NOT1 (N6826, N6825);
buf BUF1 (N6827, N6817);
xor XOR2 (N6828, N6822, N3088);
nand NAND4 (N6829, N6826, N2832, N5305, N6006);
buf BUF1 (N6830, N6827);
nor NOR4 (N6831, N6829, N3914, N4421, N6095);
and AND4 (N6832, N6823, N5460, N4706, N1960);
or OR4 (N6833, N6818, N5665, N2653, N4128);
not NOT1 (N6834, N6831);
not NOT1 (N6835, N6816);
buf BUF1 (N6836, N6824);
and AND2 (N6837, N6834, N3535);
nor NOR4 (N6838, N6820, N3770, N1592, N5059);
nand NAND3 (N6839, N6807, N1905, N6653);
buf BUF1 (N6840, N6833);
and AND4 (N6841, N6838, N1156, N520, N4368);
not NOT1 (N6842, N6836);
buf BUF1 (N6843, N6819);
buf BUF1 (N6844, N6841);
and AND2 (N6845, N6830, N6337);
nor NOR4 (N6846, N6837, N1705, N401, N479);
not NOT1 (N6847, N6844);
buf BUF1 (N6848, N6842);
nor NOR3 (N6849, N6839, N365, N1731);
buf BUF1 (N6850, N6845);
nand NAND3 (N6851, N6847, N109, N1718);
and AND2 (N6852, N6846, N4462);
nand NAND4 (N6853, N6850, N1360, N2989, N5140);
or OR4 (N6854, N6843, N6472, N3617, N2111);
nand NAND2 (N6855, N6840, N4120);
buf BUF1 (N6856, N6849);
nand NAND4 (N6857, N6855, N2587, N421, N6367);
nand NAND3 (N6858, N6853, N5597, N3677);
or OR4 (N6859, N6854, N5409, N4665, N696);
xor XOR2 (N6860, N6856, N2405);
not NOT1 (N6861, N6859);
nor NOR2 (N6862, N6835, N3859);
or OR3 (N6863, N6860, N4447, N720);
nor NOR3 (N6864, N6861, N2462, N2598);
or OR3 (N6865, N6832, N102, N3851);
and AND3 (N6866, N6848, N5627, N5304);
not NOT1 (N6867, N6864);
and AND4 (N6868, N6867, N1537, N5446, N4109);
not NOT1 (N6869, N6863);
xor XOR2 (N6870, N6869, N4839);
buf BUF1 (N6871, N6858);
nand NAND4 (N6872, N6852, N5815, N1178, N288);
and AND2 (N6873, N6862, N2871);
and AND4 (N6874, N6871, N193, N6733, N5958);
buf BUF1 (N6875, N6828);
nand NAND3 (N6876, N6868, N4892, N2106);
nor NOR4 (N6877, N6874, N3745, N29, N5257);
buf BUF1 (N6878, N6851);
nand NAND3 (N6879, N6875, N5941, N3748);
not NOT1 (N6880, N6878);
not NOT1 (N6881, N6876);
not NOT1 (N6882, N6865);
nand NAND3 (N6883, N6870, N4998, N4332);
not NOT1 (N6884, N6880);
and AND3 (N6885, N6866, N5418, N2327);
nor NOR4 (N6886, N6885, N6745, N32, N6551);
and AND2 (N6887, N6857, N1200);
buf BUF1 (N6888, N6873);
not NOT1 (N6889, N6888);
and AND4 (N6890, N6886, N6227, N2809, N1226);
buf BUF1 (N6891, N6884);
nand NAND2 (N6892, N6889, N4309);
nand NAND4 (N6893, N6891, N2232, N535, N4138);
buf BUF1 (N6894, N6893);
buf BUF1 (N6895, N6892);
xor XOR2 (N6896, N6881, N5393);
xor XOR2 (N6897, N6882, N131);
not NOT1 (N6898, N6890);
nor NOR4 (N6899, N6887, N1126, N2311, N4638);
and AND4 (N6900, N6899, N5362, N4292, N5816);
buf BUF1 (N6901, N6895);
buf BUF1 (N6902, N6898);
xor XOR2 (N6903, N6879, N4248);
xor XOR2 (N6904, N6883, N1600);
buf BUF1 (N6905, N6903);
buf BUF1 (N6906, N6894);
xor XOR2 (N6907, N6900, N431);
nor NOR3 (N6908, N6907, N4404, N3216);
and AND4 (N6909, N6897, N4154, N2696, N6038);
xor XOR2 (N6910, N6902, N3297);
nand NAND2 (N6911, N6906, N4595);
nand NAND4 (N6912, N6872, N2374, N3172, N6106);
nand NAND3 (N6913, N6911, N1932, N3204);
not NOT1 (N6914, N6877);
not NOT1 (N6915, N6901);
nor NOR2 (N6916, N6912, N2448);
nor NOR4 (N6917, N6908, N1132, N3309, N4524);
buf BUF1 (N6918, N6904);
buf BUF1 (N6919, N6913);
xor XOR2 (N6920, N6910, N3007);
not NOT1 (N6921, N6920);
and AND3 (N6922, N6919, N5733, N3574);
nor NOR4 (N6923, N6918, N1790, N2966, N6249);
and AND2 (N6924, N6917, N3830);
nor NOR3 (N6925, N6924, N585, N4913);
nand NAND2 (N6926, N6896, N315);
not NOT1 (N6927, N6915);
or OR4 (N6928, N6926, N5117, N1518, N5445);
xor XOR2 (N6929, N6914, N5715);
nand NAND2 (N6930, N6927, N2825);
nor NOR3 (N6931, N6923, N1107, N615);
nor NOR3 (N6932, N6909, N129, N4554);
buf BUF1 (N6933, N6921);
nand NAND4 (N6934, N6916, N3800, N4607, N5671);
and AND4 (N6935, N6930, N3808, N2285, N5018);
not NOT1 (N6936, N6933);
xor XOR2 (N6937, N6934, N4436);
and AND2 (N6938, N6932, N3013);
and AND2 (N6939, N6929, N2287);
and AND3 (N6940, N6937, N5587, N3776);
nand NAND4 (N6941, N6905, N4053, N3259, N3962);
and AND3 (N6942, N6931, N974, N272);
or OR3 (N6943, N6938, N6406, N234);
nor NOR2 (N6944, N6922, N4905);
buf BUF1 (N6945, N6941);
nor NOR4 (N6946, N6935, N2551, N424, N4543);
xor XOR2 (N6947, N6936, N1413);
nand NAND3 (N6948, N6925, N5584, N6233);
xor XOR2 (N6949, N6948, N3556);
buf BUF1 (N6950, N6940);
buf BUF1 (N6951, N6942);
nor NOR2 (N6952, N6951, N3903);
buf BUF1 (N6953, N6939);
or OR2 (N6954, N6953, N877);
nor NOR3 (N6955, N6950, N2258, N5147);
nor NOR3 (N6956, N6944, N5954, N4071);
buf BUF1 (N6957, N6955);
nor NOR4 (N6958, N6946, N725, N1905, N1727);
nor NOR3 (N6959, N6958, N1962, N3089);
and AND2 (N6960, N6956, N4305);
xor XOR2 (N6961, N6945, N2490);
buf BUF1 (N6962, N6928);
or OR3 (N6963, N6957, N2508, N3546);
not NOT1 (N6964, N6954);
nor NOR4 (N6965, N6962, N161, N1816, N3893);
or OR3 (N6966, N6960, N2014, N4815);
not NOT1 (N6967, N6966);
or OR3 (N6968, N6961, N1799, N2568);
not NOT1 (N6969, N6947);
or OR3 (N6970, N6964, N6197, N6634);
nand NAND3 (N6971, N6970, N600, N6412);
nor NOR2 (N6972, N6952, N755);
and AND4 (N6973, N6968, N1691, N2441, N5897);
and AND4 (N6974, N6949, N4907, N220, N198);
xor XOR2 (N6975, N6959, N277);
or OR3 (N6976, N6975, N5984, N1548);
xor XOR2 (N6977, N6973, N6490);
not NOT1 (N6978, N6977);
not NOT1 (N6979, N6969);
nand NAND4 (N6980, N6963, N6055, N3420, N5145);
or OR2 (N6981, N6976, N1896);
xor XOR2 (N6982, N6972, N5838);
and AND2 (N6983, N6971, N5153);
or OR4 (N6984, N6943, N583, N4596, N5154);
and AND4 (N6985, N6983, N5613, N6672, N6611);
and AND3 (N6986, N6965, N5788, N1098);
nor NOR3 (N6987, N6967, N3037, N2293);
not NOT1 (N6988, N6986);
nand NAND4 (N6989, N6979, N4750, N2481, N4315);
nor NOR3 (N6990, N6981, N2777, N2444);
or OR2 (N6991, N6989, N3067);
xor XOR2 (N6992, N6990, N523);
nor NOR3 (N6993, N6991, N418, N6966);
nand NAND4 (N6994, N6982, N2450, N2555, N2909);
xor XOR2 (N6995, N6980, N4798);
or OR4 (N6996, N6993, N6783, N5299, N3932);
nand NAND3 (N6997, N6985, N262, N1189);
buf BUF1 (N6998, N6974);
not NOT1 (N6999, N6984);
xor XOR2 (N7000, N6995, N5842);
and AND4 (N7001, N6997, N6277, N931, N4641);
or OR4 (N7002, N6987, N1866, N5184, N3481);
nand NAND2 (N7003, N6988, N541);
not NOT1 (N7004, N6998);
not NOT1 (N7005, N7002);
nand NAND2 (N7006, N7001, N5886);
buf BUF1 (N7007, N7000);
nand NAND3 (N7008, N7007, N4308, N4072);
nor NOR3 (N7009, N7005, N4294, N4377);
nand NAND3 (N7010, N7006, N5036, N4059);
or OR3 (N7011, N7003, N6965, N2226);
and AND3 (N7012, N7009, N3825, N1340);
and AND2 (N7013, N7008, N1765);
and AND2 (N7014, N7013, N4062);
and AND3 (N7015, N6992, N1657, N6136);
nand NAND2 (N7016, N6978, N882);
nand NAND3 (N7017, N6999, N1795, N6548);
buf BUF1 (N7018, N7015);
buf BUF1 (N7019, N6996);
not NOT1 (N7020, N7016);
not NOT1 (N7021, N7020);
xor XOR2 (N7022, N7012, N3862);
buf BUF1 (N7023, N7017);
and AND4 (N7024, N6994, N6042, N5669, N4651);
or OR2 (N7025, N7014, N1799);
not NOT1 (N7026, N7019);
not NOT1 (N7027, N7022);
or OR4 (N7028, N7027, N2854, N5540, N4308);
or OR3 (N7029, N7028, N3239, N4770);
and AND3 (N7030, N7026, N4141, N3301);
not NOT1 (N7031, N7011);
or OR3 (N7032, N7021, N4328, N5478);
nand NAND2 (N7033, N7018, N3761);
buf BUF1 (N7034, N7032);
nand NAND2 (N7035, N7024, N6173);
nand NAND4 (N7036, N7031, N4747, N6738, N1462);
buf BUF1 (N7037, N7033);
nor NOR4 (N7038, N7004, N1436, N4909, N3477);
xor XOR2 (N7039, N7036, N3040);
or OR4 (N7040, N7038, N2648, N2480, N3135);
and AND4 (N7041, N7025, N7024, N4704, N1841);
or OR2 (N7042, N7034, N4398);
and AND3 (N7043, N7042, N5359, N1678);
or OR2 (N7044, N7040, N6315);
nand NAND2 (N7045, N7044, N328);
and AND2 (N7046, N7010, N1429);
nor NOR2 (N7047, N7041, N3574);
not NOT1 (N7048, N7035);
nor NOR2 (N7049, N7029, N6485);
and AND3 (N7050, N7043, N311, N1537);
buf BUF1 (N7051, N7047);
nand NAND3 (N7052, N7049, N2561, N2967);
or OR2 (N7053, N7030, N6578);
nand NAND2 (N7054, N7046, N997);
and AND3 (N7055, N7037, N5402, N3325);
xor XOR2 (N7056, N7048, N2473);
not NOT1 (N7057, N7051);
nand NAND4 (N7058, N7054, N4275, N3484, N2933);
not NOT1 (N7059, N7050);
or OR2 (N7060, N7055, N4875);
xor XOR2 (N7061, N7060, N6648);
and AND2 (N7062, N7039, N910);
nor NOR3 (N7063, N7058, N3643, N6644);
xor XOR2 (N7064, N7063, N5072);
not NOT1 (N7065, N7064);
xor XOR2 (N7066, N7062, N3329);
not NOT1 (N7067, N7053);
xor XOR2 (N7068, N7023, N2964);
and AND3 (N7069, N7065, N5003, N1875);
and AND3 (N7070, N7061, N798, N672);
and AND3 (N7071, N7069, N655, N5614);
nand NAND2 (N7072, N7056, N882);
buf BUF1 (N7073, N7057);
or OR4 (N7074, N7066, N5636, N2282, N1790);
not NOT1 (N7075, N7052);
not NOT1 (N7076, N7074);
nor NOR3 (N7077, N7072, N839, N3730);
not NOT1 (N7078, N7073);
and AND2 (N7079, N7078, N313);
nand NAND4 (N7080, N7079, N3899, N119, N5158);
and AND4 (N7081, N7080, N4018, N6353, N6419);
nor NOR3 (N7082, N7070, N1389, N299);
nand NAND4 (N7083, N7067, N6972, N6525, N5330);
and AND3 (N7084, N7082, N986, N6000);
not NOT1 (N7085, N7077);
or OR2 (N7086, N7083, N4433);
nor NOR3 (N7087, N7085, N5032, N6335);
not NOT1 (N7088, N7068);
nor NOR3 (N7089, N7081, N6888, N6092);
and AND3 (N7090, N7076, N2948, N1810);
buf BUF1 (N7091, N7088);
buf BUF1 (N7092, N7084);
nand NAND3 (N7093, N7089, N349, N1221);
nor NOR4 (N7094, N7091, N6037, N3511, N1405);
or OR4 (N7095, N7045, N2081, N4612, N3963);
and AND3 (N7096, N7094, N6265, N1547);
nand NAND2 (N7097, N7090, N399);
not NOT1 (N7098, N7097);
not NOT1 (N7099, N7098);
and AND2 (N7100, N7087, N5248);
and AND3 (N7101, N7096, N4095, N5978);
nand NAND3 (N7102, N7075, N1370, N5254);
not NOT1 (N7103, N7099);
not NOT1 (N7104, N7102);
nor NOR2 (N7105, N7095, N1971);
and AND2 (N7106, N7101, N2299);
xor XOR2 (N7107, N7100, N4244);
and AND3 (N7108, N7059, N4559, N7045);
xor XOR2 (N7109, N7103, N566);
or OR4 (N7110, N7109, N614, N1181, N2084);
and AND2 (N7111, N7092, N3045);
or OR3 (N7112, N7104, N3649, N471);
not NOT1 (N7113, N7108);
nor NOR4 (N7114, N7086, N1025, N2615, N3657);
nor NOR4 (N7115, N7114, N2165, N6529, N5203);
buf BUF1 (N7116, N7093);
nor NOR3 (N7117, N7106, N3561, N6273);
xor XOR2 (N7118, N7071, N1160);
nand NAND3 (N7119, N7118, N1314, N4702);
and AND3 (N7120, N7112, N6758, N4023);
or OR4 (N7121, N7107, N3958, N2674, N2904);
xor XOR2 (N7122, N7111, N4950);
and AND3 (N7123, N7117, N4542, N1166);
nor NOR2 (N7124, N7119, N6891);
xor XOR2 (N7125, N7120, N3283);
not NOT1 (N7126, N7124);
nor NOR4 (N7127, N7113, N762, N5951, N5246);
or OR4 (N7128, N7125, N4981, N1114, N1898);
nor NOR2 (N7129, N7115, N3623);
buf BUF1 (N7130, N7126);
and AND3 (N7131, N7110, N2997, N6346);
not NOT1 (N7132, N7116);
xor XOR2 (N7133, N7129, N3976);
not NOT1 (N7134, N7130);
buf BUF1 (N7135, N7105);
xor XOR2 (N7136, N7132, N2022);
xor XOR2 (N7137, N7123, N6206);
buf BUF1 (N7138, N7131);
buf BUF1 (N7139, N7135);
buf BUF1 (N7140, N7133);
nor NOR2 (N7141, N7128, N5603);
xor XOR2 (N7142, N7122, N5711);
xor XOR2 (N7143, N7136, N5437);
buf BUF1 (N7144, N7121);
nand NAND3 (N7145, N7140, N1979, N1228);
nand NAND3 (N7146, N7142, N1492, N610);
nor NOR2 (N7147, N7134, N5124);
buf BUF1 (N7148, N7147);
or OR4 (N7149, N7137, N2661, N7072, N1590);
buf BUF1 (N7150, N7146);
or OR4 (N7151, N7149, N4994, N3776, N3850);
nand NAND2 (N7152, N7145, N5331);
not NOT1 (N7153, N7144);
xor XOR2 (N7154, N7138, N2358);
xor XOR2 (N7155, N7139, N6101);
nor NOR4 (N7156, N7141, N6724, N6086, N2380);
buf BUF1 (N7157, N7152);
xor XOR2 (N7158, N7155, N164);
nand NAND3 (N7159, N7153, N5121, N2424);
not NOT1 (N7160, N7156);
or OR4 (N7161, N7143, N213, N1038, N2609);
nand NAND3 (N7162, N7148, N691, N4183);
buf BUF1 (N7163, N7150);
and AND3 (N7164, N7158, N2396, N3500);
and AND2 (N7165, N7164, N5364);
and AND2 (N7166, N7154, N484);
nor NOR4 (N7167, N7166, N5380, N1909, N1662);
or OR2 (N7168, N7165, N1683);
xor XOR2 (N7169, N7167, N6254);
not NOT1 (N7170, N7159);
nand NAND4 (N7171, N7160, N2965, N397, N653);
nor NOR3 (N7172, N7168, N1617, N2931);
nand NAND4 (N7173, N7170, N5168, N6491, N3840);
and AND4 (N7174, N7173, N4005, N1730, N6799);
and AND3 (N7175, N7162, N3098, N6021);
buf BUF1 (N7176, N7172);
buf BUF1 (N7177, N7163);
or OR2 (N7178, N7177, N4331);
buf BUF1 (N7179, N7171);
or OR3 (N7180, N7174, N5274, N4897);
buf BUF1 (N7181, N7151);
and AND2 (N7182, N7179, N2790);
nand NAND3 (N7183, N7176, N685, N3837);
xor XOR2 (N7184, N7127, N3747);
or OR2 (N7185, N7169, N1195);
or OR4 (N7186, N7181, N4683, N5985, N3539);
and AND2 (N7187, N7185, N5637);
buf BUF1 (N7188, N7183);
xor XOR2 (N7189, N7175, N3506);
nor NOR2 (N7190, N7189, N3001);
or OR4 (N7191, N7188, N5113, N1558, N1332);
buf BUF1 (N7192, N7191);
or OR2 (N7193, N7184, N6262);
not NOT1 (N7194, N7190);
or OR4 (N7195, N7161, N6525, N6134, N2104);
or OR4 (N7196, N7192, N7111, N5512, N1811);
nor NOR4 (N7197, N7182, N3515, N1905, N3456);
or OR2 (N7198, N7157, N5920);
xor XOR2 (N7199, N7180, N7037);
buf BUF1 (N7200, N7194);
and AND4 (N7201, N7199, N3177, N1215, N873);
xor XOR2 (N7202, N7201, N1350);
not NOT1 (N7203, N7178);
not NOT1 (N7204, N7202);
not NOT1 (N7205, N7200);
not NOT1 (N7206, N7197);
or OR3 (N7207, N7205, N6973, N4212);
and AND3 (N7208, N7193, N1979, N4979);
xor XOR2 (N7209, N7208, N5489);
not NOT1 (N7210, N7203);
or OR4 (N7211, N7207, N4077, N4156, N3746);
nor NOR3 (N7212, N7187, N1936, N4468);
not NOT1 (N7213, N7212);
buf BUF1 (N7214, N7196);
nand NAND4 (N7215, N7204, N1929, N1385, N2035);
and AND2 (N7216, N7198, N4551);
buf BUF1 (N7217, N7210);
not NOT1 (N7218, N7216);
or OR3 (N7219, N7195, N358, N4629);
xor XOR2 (N7220, N7186, N4696);
and AND2 (N7221, N7206, N22);
xor XOR2 (N7222, N7217, N2181);
nand NAND2 (N7223, N7209, N339);
and AND4 (N7224, N7222, N1612, N370, N7090);
not NOT1 (N7225, N7223);
or OR2 (N7226, N7220, N2762);
nand NAND4 (N7227, N7211, N4479, N5249, N3170);
xor XOR2 (N7228, N7219, N694);
not NOT1 (N7229, N7227);
and AND2 (N7230, N7226, N3658);
nor NOR4 (N7231, N7218, N6274, N1057, N4676);
buf BUF1 (N7232, N7214);
nor NOR4 (N7233, N7230, N377, N1335, N5452);
nor NOR3 (N7234, N7232, N2933, N215);
nand NAND3 (N7235, N7229, N795, N883);
or OR2 (N7236, N7213, N6527);
xor XOR2 (N7237, N7225, N1167);
nand NAND3 (N7238, N7221, N5605, N4902);
nand NAND2 (N7239, N7233, N1057);
nor NOR2 (N7240, N7235, N30);
or OR2 (N7241, N7238, N5034);
not NOT1 (N7242, N7231);
or OR4 (N7243, N7234, N36, N314, N5804);
and AND3 (N7244, N7241, N988, N684);
xor XOR2 (N7245, N7236, N2779);
xor XOR2 (N7246, N7240, N2048);
nor NOR4 (N7247, N7215, N120, N6922, N5737);
and AND2 (N7248, N7243, N5216);
not NOT1 (N7249, N7247);
buf BUF1 (N7250, N7249);
and AND3 (N7251, N7245, N3701, N650);
not NOT1 (N7252, N7244);
nand NAND3 (N7253, N7248, N6662, N6549);
buf BUF1 (N7254, N7246);
not NOT1 (N7255, N7251);
buf BUF1 (N7256, N7242);
nor NOR2 (N7257, N7252, N5717);
nand NAND2 (N7258, N7253, N1500);
xor XOR2 (N7259, N7228, N6648);
buf BUF1 (N7260, N7237);
buf BUF1 (N7261, N7258);
nand NAND4 (N7262, N7254, N4004, N1556, N4913);
nor NOR4 (N7263, N7224, N3393, N2189, N6190);
xor XOR2 (N7264, N7263, N1470);
or OR2 (N7265, N7256, N355);
not NOT1 (N7266, N7257);
and AND3 (N7267, N7255, N105, N1107);
or OR4 (N7268, N7250, N2279, N683, N6838);
nor NOR2 (N7269, N7262, N1050);
or OR4 (N7270, N7239, N2010, N5557, N42);
and AND3 (N7271, N7268, N4786, N5241);
buf BUF1 (N7272, N7259);
or OR2 (N7273, N7267, N4613);
and AND3 (N7274, N7265, N5870, N906);
and AND4 (N7275, N7260, N998, N5131, N1950);
xor XOR2 (N7276, N7270, N5411);
nand NAND3 (N7277, N7276, N3314, N104);
and AND4 (N7278, N7264, N2540, N2624, N2501);
not NOT1 (N7279, N7277);
not NOT1 (N7280, N7279);
or OR4 (N7281, N7269, N6141, N2366, N5585);
nor NOR3 (N7282, N7272, N333, N2451);
or OR2 (N7283, N7281, N4351);
and AND2 (N7284, N7280, N6763);
nand NAND3 (N7285, N7274, N2419, N719);
not NOT1 (N7286, N7284);
not NOT1 (N7287, N7275);
or OR2 (N7288, N7266, N3869);
nand NAND4 (N7289, N7282, N5048, N2774, N1928);
and AND2 (N7290, N7288, N2661);
not NOT1 (N7291, N7287);
and AND3 (N7292, N7291, N2808, N3403);
or OR2 (N7293, N7285, N4473);
nor NOR3 (N7294, N7289, N5434, N287);
nor NOR4 (N7295, N7273, N4153, N2185, N6317);
nand NAND3 (N7296, N7261, N3087, N5416);
and AND3 (N7297, N7295, N4087, N6092);
buf BUF1 (N7298, N7283);
nand NAND3 (N7299, N7286, N3661, N2000);
and AND3 (N7300, N7293, N2032, N5688);
not NOT1 (N7301, N7278);
nand NAND2 (N7302, N7297, N1010);
xor XOR2 (N7303, N7296, N6970);
xor XOR2 (N7304, N7300, N5474);
buf BUF1 (N7305, N7292);
or OR3 (N7306, N7290, N6776, N1092);
xor XOR2 (N7307, N7298, N38);
not NOT1 (N7308, N7306);
nor NOR2 (N7309, N7304, N4113);
nand NAND2 (N7310, N7308, N4305);
nor NOR4 (N7311, N7299, N1629, N3767, N5698);
and AND2 (N7312, N7307, N1111);
not NOT1 (N7313, N7303);
nand NAND4 (N7314, N7294, N1591, N2377, N5120);
nor NOR4 (N7315, N7314, N5777, N5415, N6416);
nor NOR4 (N7316, N7313, N4777, N3030, N6747);
buf BUF1 (N7317, N7301);
and AND3 (N7318, N7311, N5991, N4402);
xor XOR2 (N7319, N7315, N1617);
nor NOR3 (N7320, N7319, N3923, N538);
not NOT1 (N7321, N7316);
nand NAND2 (N7322, N7317, N5258);
and AND4 (N7323, N7302, N5943, N5154, N2885);
not NOT1 (N7324, N7305);
nor NOR3 (N7325, N7312, N3110, N2373);
nand NAND4 (N7326, N7322, N2077, N6705, N5374);
nand NAND3 (N7327, N7318, N6798, N1608);
buf BUF1 (N7328, N7323);
xor XOR2 (N7329, N7310, N2141);
xor XOR2 (N7330, N7309, N700);
nor NOR2 (N7331, N7271, N2220);
nor NOR2 (N7332, N7331, N7017);
xor XOR2 (N7333, N7330, N6760);
nand NAND2 (N7334, N7321, N2726);
nand NAND2 (N7335, N7325, N1283);
xor XOR2 (N7336, N7324, N3590);
not NOT1 (N7337, N7320);
nand NAND3 (N7338, N7329, N2167, N1861);
nor NOR4 (N7339, N7336, N4391, N4128, N2257);
and AND4 (N7340, N7334, N3382, N3341, N982);
nand NAND4 (N7341, N7338, N6505, N1985, N6255);
nor NOR3 (N7342, N7328, N4552, N5690);
and AND4 (N7343, N7342, N4432, N6597, N781);
buf BUF1 (N7344, N7337);
nand NAND3 (N7345, N7326, N635, N5602);
nor NOR2 (N7346, N7333, N6793);
and AND4 (N7347, N7339, N2240, N6059, N2156);
not NOT1 (N7348, N7327);
and AND2 (N7349, N7345, N5475);
and AND4 (N7350, N7340, N6717, N6635, N6113);
and AND4 (N7351, N7347, N944, N4264, N5271);
and AND3 (N7352, N7341, N6279, N3635);
xor XOR2 (N7353, N7352, N6228);
buf BUF1 (N7354, N7335);
nor NOR2 (N7355, N7343, N356);
nor NOR4 (N7356, N7351, N6930, N3560, N4278);
and AND4 (N7357, N7353, N2638, N5581, N5057);
nand NAND2 (N7358, N7356, N1524);
not NOT1 (N7359, N7332);
not NOT1 (N7360, N7344);
nand NAND2 (N7361, N7357, N748);
and AND2 (N7362, N7350, N1705);
nor NOR2 (N7363, N7360, N4662);
or OR3 (N7364, N7361, N5731, N6439);
nor NOR4 (N7365, N7346, N7073, N3799, N2778);
nor NOR2 (N7366, N7364, N7219);
not NOT1 (N7367, N7359);
xor XOR2 (N7368, N7365, N1506);
and AND2 (N7369, N7355, N6394);
and AND4 (N7370, N7368, N2889, N67, N1227);
xor XOR2 (N7371, N7363, N1591);
or OR4 (N7372, N7348, N3040, N806, N4214);
nand NAND3 (N7373, N7362, N932, N3751);
not NOT1 (N7374, N7373);
xor XOR2 (N7375, N7367, N6223);
nand NAND4 (N7376, N7372, N5887, N2691, N1952);
or OR4 (N7377, N7376, N4188, N2810, N4599);
and AND2 (N7378, N7369, N3091);
or OR4 (N7379, N7371, N6960, N7216, N7335);
nor NOR3 (N7380, N7366, N1818, N526);
xor XOR2 (N7381, N7378, N4463);
and AND2 (N7382, N7358, N6926);
not NOT1 (N7383, N7377);
buf BUF1 (N7384, N7354);
buf BUF1 (N7385, N7380);
nor NOR4 (N7386, N7349, N2254, N3897, N2315);
nand NAND4 (N7387, N7370, N47, N3306, N2462);
and AND2 (N7388, N7375, N6303);
nand NAND4 (N7389, N7388, N2170, N1810, N5400);
not NOT1 (N7390, N7385);
or OR4 (N7391, N7389, N4492, N3742, N4242);
xor XOR2 (N7392, N7390, N681);
nand NAND2 (N7393, N7379, N4123);
or OR3 (N7394, N7392, N1739, N4596);
nor NOR2 (N7395, N7383, N631);
buf BUF1 (N7396, N7391);
nand NAND4 (N7397, N7393, N1696, N5722, N1576);
nand NAND3 (N7398, N7395, N4324, N5598);
or OR4 (N7399, N7387, N4609, N5807, N219);
nor NOR3 (N7400, N7398, N1962, N6017);
and AND3 (N7401, N7399, N252, N649);
nand NAND2 (N7402, N7394, N1138);
not NOT1 (N7403, N7396);
and AND4 (N7404, N7401, N7216, N7399, N3970);
xor XOR2 (N7405, N7382, N3895);
not NOT1 (N7406, N7402);
nand NAND2 (N7407, N7406, N4981);
or OR3 (N7408, N7400, N6204, N6823);
nor NOR2 (N7409, N7374, N4429);
or OR4 (N7410, N7397, N416, N6971, N6840);
buf BUF1 (N7411, N7408);
or OR4 (N7412, N7411, N1214, N3301, N6031);
and AND4 (N7413, N7405, N2128, N7100, N1453);
and AND3 (N7414, N7381, N6801, N70);
and AND4 (N7415, N7414, N5208, N6317, N4615);
not NOT1 (N7416, N7415);
or OR2 (N7417, N7404, N7288);
or OR4 (N7418, N7410, N186, N5528, N2685);
xor XOR2 (N7419, N7418, N5904);
buf BUF1 (N7420, N7409);
buf BUF1 (N7421, N7386);
nand NAND4 (N7422, N7417, N7261, N4092, N7210);
buf BUF1 (N7423, N7421);
nor NOR3 (N7424, N7384, N757, N3075);
nor NOR2 (N7425, N7416, N5851);
or OR2 (N7426, N7413, N5909);
and AND2 (N7427, N7425, N6218);
buf BUF1 (N7428, N7427);
nand NAND3 (N7429, N7422, N7303, N245);
and AND3 (N7430, N7403, N447, N4534);
nor NOR4 (N7431, N7407, N2991, N5793, N5950);
buf BUF1 (N7432, N7420);
nor NOR4 (N7433, N7429, N4900, N1871, N1281);
buf BUF1 (N7434, N7431);
nand NAND3 (N7435, N7412, N7011, N3205);
xor XOR2 (N7436, N7419, N6587);
nand NAND3 (N7437, N7423, N4018, N2402);
not NOT1 (N7438, N7436);
or OR4 (N7439, N7438, N2821, N45, N7240);
nor NOR2 (N7440, N7430, N6217);
nor NOR2 (N7441, N7424, N5541);
or OR4 (N7442, N7432, N6636, N3229, N6293);
nand NAND3 (N7443, N7437, N5072, N3882);
and AND2 (N7444, N7435, N4089);
not NOT1 (N7445, N7433);
nand NAND2 (N7446, N7442, N4609);
buf BUF1 (N7447, N7440);
buf BUF1 (N7448, N7443);
nor NOR2 (N7449, N7446, N6961);
buf BUF1 (N7450, N7449);
xor XOR2 (N7451, N7441, N2103);
and AND2 (N7452, N7428, N3161);
nor NOR2 (N7453, N7448, N2384);
not NOT1 (N7454, N7445);
nor NOR3 (N7455, N7434, N5676, N1143);
xor XOR2 (N7456, N7453, N6320);
buf BUF1 (N7457, N7456);
buf BUF1 (N7458, N7439);
not NOT1 (N7459, N7444);
and AND2 (N7460, N7426, N529);
nor NOR4 (N7461, N7457, N3388, N6779, N1818);
nand NAND3 (N7462, N7458, N5412, N1372);
buf BUF1 (N7463, N7461);
or OR4 (N7464, N7454, N4315, N1776, N1799);
buf BUF1 (N7465, N7452);
or OR2 (N7466, N7447, N2385);
or OR2 (N7467, N7450, N1203);
nor NOR2 (N7468, N7467, N744);
nor NOR2 (N7469, N7468, N5383);
or OR3 (N7470, N7460, N198, N6901);
nor NOR3 (N7471, N7464, N6039, N6457);
xor XOR2 (N7472, N7462, N3062);
not NOT1 (N7473, N7472);
xor XOR2 (N7474, N7463, N502);
buf BUF1 (N7475, N7470);
buf BUF1 (N7476, N7469);
or OR2 (N7477, N7455, N182);
buf BUF1 (N7478, N7474);
or OR3 (N7479, N7478, N1850, N984);
or OR3 (N7480, N7473, N5765, N4765);
and AND4 (N7481, N7475, N4929, N7177, N4749);
or OR4 (N7482, N7471, N2604, N193, N1480);
xor XOR2 (N7483, N7459, N5107);
buf BUF1 (N7484, N7465);
and AND2 (N7485, N7476, N6089);
not NOT1 (N7486, N7484);
buf BUF1 (N7487, N7480);
or OR3 (N7488, N7487, N2961, N4506);
or OR2 (N7489, N7483, N3762);
nor NOR4 (N7490, N7479, N5460, N7371, N4027);
or OR4 (N7491, N7490, N2816, N2758, N5720);
buf BUF1 (N7492, N7485);
xor XOR2 (N7493, N7482, N4626);
nand NAND3 (N7494, N7492, N5316, N5298);
nor NOR4 (N7495, N7493, N5184, N6769, N5531);
not NOT1 (N7496, N7486);
and AND4 (N7497, N7489, N1801, N5446, N1125);
not NOT1 (N7498, N7477);
and AND4 (N7499, N7488, N3106, N7036, N85);
buf BUF1 (N7500, N7494);
xor XOR2 (N7501, N7495, N2639);
xor XOR2 (N7502, N7496, N2540);
xor XOR2 (N7503, N7497, N4979);
buf BUF1 (N7504, N7481);
or OR3 (N7505, N7498, N6779, N6102);
and AND4 (N7506, N7500, N4175, N4791, N3047);
or OR3 (N7507, N7499, N5307, N3848);
and AND4 (N7508, N7491, N5911, N2755, N5881);
nor NOR2 (N7509, N7505, N1962);
nor NOR3 (N7510, N7501, N4989, N1607);
or OR3 (N7511, N7504, N4350, N83);
buf BUF1 (N7512, N7502);
not NOT1 (N7513, N7509);
nor NOR4 (N7514, N7511, N3416, N701, N5026);
not NOT1 (N7515, N7503);
nand NAND2 (N7516, N7512, N3779);
not NOT1 (N7517, N7451);
or OR2 (N7518, N7513, N5875);
or OR4 (N7519, N7508, N7256, N5588, N1489);
and AND4 (N7520, N7514, N7038, N873, N1260);
and AND3 (N7521, N7506, N4765, N3108);
nand NAND4 (N7522, N7515, N1909, N1363, N2001);
nor NOR3 (N7523, N7521, N5527, N5005);
xor XOR2 (N7524, N7518, N4242);
and AND2 (N7525, N7523, N1587);
or OR3 (N7526, N7516, N2151, N1141);
and AND2 (N7527, N7526, N3572);
or OR4 (N7528, N7527, N2080, N2927, N2601);
not NOT1 (N7529, N7519);
buf BUF1 (N7530, N7466);
xor XOR2 (N7531, N7525, N7073);
and AND3 (N7532, N7507, N5876, N1402);
nand NAND2 (N7533, N7531, N6328);
and AND2 (N7534, N7517, N7447);
not NOT1 (N7535, N7520);
or OR4 (N7536, N7524, N4267, N4702, N3898);
xor XOR2 (N7537, N7533, N4228);
nand NAND4 (N7538, N7510, N6866, N730, N4740);
buf BUF1 (N7539, N7536);
or OR4 (N7540, N7530, N2308, N4587, N5404);
nand NAND4 (N7541, N7538, N289, N6564, N5351);
xor XOR2 (N7542, N7535, N5890);
nand NAND2 (N7543, N7528, N7344);
nor NOR2 (N7544, N7542, N1752);
xor XOR2 (N7545, N7522, N7445);
not NOT1 (N7546, N7529);
nand NAND3 (N7547, N7532, N2197, N6201);
and AND4 (N7548, N7540, N5245, N2874, N4097);
not NOT1 (N7549, N7544);
xor XOR2 (N7550, N7534, N5803);
not NOT1 (N7551, N7541);
not NOT1 (N7552, N7537);
buf BUF1 (N7553, N7550);
and AND4 (N7554, N7543, N624, N5014, N587);
and AND4 (N7555, N7545, N5812, N6541, N4460);
not NOT1 (N7556, N7551);
nor NOR3 (N7557, N7554, N5274, N4083);
and AND2 (N7558, N7556, N2150);
nor NOR2 (N7559, N7548, N5711);
nor NOR2 (N7560, N7547, N3353);
not NOT1 (N7561, N7557);
nor NOR4 (N7562, N7558, N300, N5993, N5409);
buf BUF1 (N7563, N7546);
xor XOR2 (N7564, N7562, N4164);
or OR3 (N7565, N7553, N127, N2393);
nand NAND2 (N7566, N7552, N1915);
buf BUF1 (N7567, N7565);
or OR4 (N7568, N7559, N3386, N5824, N6020);
not NOT1 (N7569, N7549);
and AND2 (N7570, N7564, N7342);
or OR2 (N7571, N7568, N4031);
or OR2 (N7572, N7571, N5310);
nor NOR3 (N7573, N7569, N6489, N1914);
not NOT1 (N7574, N7561);
or OR3 (N7575, N7563, N2877, N1205);
xor XOR2 (N7576, N7560, N2059);
and AND4 (N7577, N7576, N2687, N1642, N2733);
not NOT1 (N7578, N7572);
and AND2 (N7579, N7570, N2325);
nand NAND2 (N7580, N7573, N937);
nand NAND4 (N7581, N7555, N2307, N2793, N6456);
xor XOR2 (N7582, N7581, N4032);
nor NOR4 (N7583, N7566, N1408, N3820, N3587);
nand NAND2 (N7584, N7574, N1969);
and AND3 (N7585, N7539, N4226, N7244);
nand NAND3 (N7586, N7585, N3768, N1472);
or OR4 (N7587, N7586, N5220, N4259, N2075);
nand NAND2 (N7588, N7578, N494);
nor NOR2 (N7589, N7583, N3374);
nor NOR3 (N7590, N7589, N5372, N297);
xor XOR2 (N7591, N7577, N224);
nor NOR2 (N7592, N7582, N4407);
not NOT1 (N7593, N7575);
xor XOR2 (N7594, N7590, N7257);
buf BUF1 (N7595, N7567);
not NOT1 (N7596, N7580);
or OR3 (N7597, N7595, N468, N5925);
nor NOR4 (N7598, N7587, N6352, N3067, N3606);
nand NAND4 (N7599, N7593, N2679, N1013, N6098);
or OR3 (N7600, N7598, N6873, N5312);
and AND3 (N7601, N7594, N546, N4802);
xor XOR2 (N7602, N7596, N6196);
xor XOR2 (N7603, N7602, N5319);
nand NAND2 (N7604, N7591, N277);
and AND3 (N7605, N7592, N5395, N7035);
xor XOR2 (N7606, N7597, N6591);
nor NOR2 (N7607, N7603, N2351);
nand NAND2 (N7608, N7588, N7515);
or OR2 (N7609, N7601, N1532);
xor XOR2 (N7610, N7584, N918);
and AND4 (N7611, N7609, N3586, N5804, N2902);
or OR3 (N7612, N7599, N5872, N7513);
buf BUF1 (N7613, N7605);
or OR3 (N7614, N7606, N5968, N4805);
nor NOR4 (N7615, N7600, N2582, N5934, N458);
nor NOR3 (N7616, N7614, N7461, N1383);
not NOT1 (N7617, N7607);
xor XOR2 (N7618, N7610, N3732);
not NOT1 (N7619, N7615);
not NOT1 (N7620, N7579);
not NOT1 (N7621, N7608);
not NOT1 (N7622, N7617);
nand NAND4 (N7623, N7620, N4317, N1665, N7095);
and AND4 (N7624, N7622, N655, N2163, N6884);
not NOT1 (N7625, N7611);
or OR3 (N7626, N7621, N5208, N6432);
not NOT1 (N7627, N7604);
buf BUF1 (N7628, N7623);
xor XOR2 (N7629, N7624, N923);
nor NOR3 (N7630, N7625, N5765, N4320);
nor NOR2 (N7631, N7627, N5848);
and AND2 (N7632, N7628, N7062);
nand NAND2 (N7633, N7626, N895);
not NOT1 (N7634, N7612);
xor XOR2 (N7635, N7632, N5915);
nand NAND4 (N7636, N7635, N5496, N2504, N162);
nor NOR2 (N7637, N7634, N3681);
or OR2 (N7638, N7636, N4791);
nor NOR4 (N7639, N7633, N6068, N1918, N33);
nand NAND4 (N7640, N7629, N5505, N110, N4631);
or OR2 (N7641, N7640, N6046);
or OR4 (N7642, N7639, N7148, N5542, N7171);
nor NOR4 (N7643, N7616, N2339, N7135, N1367);
and AND3 (N7644, N7619, N4497, N872);
xor XOR2 (N7645, N7638, N5950);
xor XOR2 (N7646, N7613, N4598);
xor XOR2 (N7647, N7646, N1424);
or OR4 (N7648, N7641, N3543, N3762, N2097);
buf BUF1 (N7649, N7643);
nand NAND4 (N7650, N7645, N7281, N4265, N4675);
buf BUF1 (N7651, N7648);
or OR3 (N7652, N7650, N4644, N3641);
nor NOR3 (N7653, N7651, N3729, N7151);
not NOT1 (N7654, N7618);
xor XOR2 (N7655, N7631, N1745);
nand NAND3 (N7656, N7655, N2501, N5649);
buf BUF1 (N7657, N7654);
xor XOR2 (N7658, N7630, N7634);
nor NOR4 (N7659, N7649, N84, N6716, N551);
nand NAND2 (N7660, N7653, N943);
buf BUF1 (N7661, N7659);
nand NAND4 (N7662, N7637, N7315, N3688, N5670);
xor XOR2 (N7663, N7642, N2070);
buf BUF1 (N7664, N7647);
xor XOR2 (N7665, N7664, N4201);
nor NOR4 (N7666, N7665, N3480, N2224, N5521);
nand NAND2 (N7667, N7661, N2186);
nand NAND4 (N7668, N7662, N1314, N4525, N7006);
nor NOR4 (N7669, N7663, N3041, N1974, N7107);
xor XOR2 (N7670, N7644, N7274);
nor NOR3 (N7671, N7658, N6382, N3006);
buf BUF1 (N7672, N7670);
not NOT1 (N7673, N7667);
xor XOR2 (N7674, N7660, N3523);
xor XOR2 (N7675, N7668, N6012);
and AND3 (N7676, N7652, N1453, N7098);
not NOT1 (N7677, N7673);
not NOT1 (N7678, N7672);
not NOT1 (N7679, N7676);
nor NOR3 (N7680, N7671, N2564, N7667);
not NOT1 (N7681, N7678);
buf BUF1 (N7682, N7669);
nand NAND3 (N7683, N7679, N5797, N7252);
nand NAND2 (N7684, N7656, N4577);
and AND3 (N7685, N7682, N3114, N6150);
not NOT1 (N7686, N7677);
nor NOR4 (N7687, N7681, N858, N2638, N5239);
xor XOR2 (N7688, N7674, N6394);
and AND2 (N7689, N7686, N5964);
buf BUF1 (N7690, N7688);
xor XOR2 (N7691, N7675, N1169);
nand NAND3 (N7692, N7691, N3576, N4372);
and AND3 (N7693, N7680, N314, N4836);
not NOT1 (N7694, N7692);
and AND2 (N7695, N7657, N7020);
nand NAND4 (N7696, N7690, N7551, N3877, N4077);
buf BUF1 (N7697, N7695);
and AND3 (N7698, N7666, N5439, N2768);
or OR4 (N7699, N7693, N2350, N4032, N1918);
not NOT1 (N7700, N7699);
nand NAND2 (N7701, N7697, N7120);
nand NAND3 (N7702, N7684, N6580, N7635);
not NOT1 (N7703, N7698);
not NOT1 (N7704, N7694);
xor XOR2 (N7705, N7704, N744);
nor NOR4 (N7706, N7689, N1694, N5446, N7390);
or OR3 (N7707, N7706, N133, N2390);
nor NOR4 (N7708, N7696, N4525, N3634, N4540);
buf BUF1 (N7709, N7700);
not NOT1 (N7710, N7683);
buf BUF1 (N7711, N7708);
or OR2 (N7712, N7685, N1249);
not NOT1 (N7713, N7701);
buf BUF1 (N7714, N7703);
not NOT1 (N7715, N7709);
buf BUF1 (N7716, N7687);
buf BUF1 (N7717, N7702);
and AND2 (N7718, N7715, N2436);
nor NOR3 (N7719, N7713, N81, N1441);
nand NAND2 (N7720, N7714, N3789);
or OR4 (N7721, N7712, N4701, N6278, N1435);
or OR2 (N7722, N7710, N1103);
nor NOR3 (N7723, N7717, N7119, N2046);
not NOT1 (N7724, N7711);
or OR2 (N7725, N7707, N2646);
xor XOR2 (N7726, N7720, N6521);
and AND4 (N7727, N7718, N1712, N1671, N7419);
buf BUF1 (N7728, N7722);
nand NAND3 (N7729, N7716, N3151, N3210);
or OR3 (N7730, N7723, N7303, N7172);
xor XOR2 (N7731, N7705, N227);
nand NAND4 (N7732, N7731, N4775, N6753, N4947);
nand NAND4 (N7733, N7730, N1300, N1858, N93);
and AND2 (N7734, N7732, N2297);
not NOT1 (N7735, N7729);
buf BUF1 (N7736, N7724);
or OR4 (N7737, N7721, N6786, N7567, N1811);
and AND2 (N7738, N7727, N6867);
and AND3 (N7739, N7734, N1194, N3991);
xor XOR2 (N7740, N7719, N6901);
nor NOR3 (N7741, N7737, N4152, N6142);
xor XOR2 (N7742, N7740, N5312);
or OR3 (N7743, N7736, N4818, N4123);
nor NOR4 (N7744, N7739, N1339, N3202, N4912);
and AND3 (N7745, N7726, N5670, N6960);
nor NOR3 (N7746, N7743, N6056, N5777);
xor XOR2 (N7747, N7725, N7277);
nand NAND2 (N7748, N7746, N2367);
nand NAND2 (N7749, N7741, N2693);
not NOT1 (N7750, N7742);
nor NOR4 (N7751, N7745, N5462, N2652, N6720);
and AND2 (N7752, N7728, N7061);
or OR4 (N7753, N7747, N1433, N5207, N4634);
or OR3 (N7754, N7735, N4619, N4779);
not NOT1 (N7755, N7748);
buf BUF1 (N7756, N7750);
nor NOR3 (N7757, N7754, N5338, N2469);
xor XOR2 (N7758, N7756, N268);
buf BUF1 (N7759, N7758);
buf BUF1 (N7760, N7751);
nand NAND2 (N7761, N7744, N3674);
nor NOR4 (N7762, N7761, N1605, N6595, N3800);
or OR2 (N7763, N7755, N5331);
and AND2 (N7764, N7749, N944);
nand NAND3 (N7765, N7738, N52, N1718);
nor NOR4 (N7766, N7757, N370, N5404, N2441);
buf BUF1 (N7767, N7752);
and AND2 (N7768, N7753, N959);
nor NOR2 (N7769, N7767, N2801);
nor NOR2 (N7770, N7760, N1666);
nor NOR4 (N7771, N7733, N5987, N359, N3447);
buf BUF1 (N7772, N7762);
or OR2 (N7773, N7770, N5029);
and AND4 (N7774, N7769, N5826, N301, N796);
and AND2 (N7775, N7771, N7312);
buf BUF1 (N7776, N7765);
buf BUF1 (N7777, N7776);
and AND2 (N7778, N7774, N4003);
nand NAND3 (N7779, N7766, N1532, N6839);
and AND3 (N7780, N7768, N7204, N2915);
nor NOR2 (N7781, N7759, N6825);
or OR4 (N7782, N7764, N4842, N2774, N5118);
and AND4 (N7783, N7778, N5897, N2931, N7729);
or OR2 (N7784, N7763, N1060);
or OR2 (N7785, N7773, N2160);
buf BUF1 (N7786, N7784);
not NOT1 (N7787, N7781);
or OR3 (N7788, N7772, N4714, N3707);
buf BUF1 (N7789, N7777);
not NOT1 (N7790, N7775);
xor XOR2 (N7791, N7790, N2558);
buf BUF1 (N7792, N7791);
nand NAND4 (N7793, N7787, N3939, N4459, N2761);
not NOT1 (N7794, N7780);
nand NAND4 (N7795, N7786, N5692, N7567, N5042);
or OR2 (N7796, N7779, N5601);
not NOT1 (N7797, N7792);
and AND2 (N7798, N7785, N3334);
buf BUF1 (N7799, N7782);
and AND2 (N7800, N7795, N280);
or OR2 (N7801, N7789, N350);
not NOT1 (N7802, N7799);
xor XOR2 (N7803, N7798, N3590);
xor XOR2 (N7804, N7801, N4997);
nor NOR3 (N7805, N7800, N1413, N7349);
nand NAND2 (N7806, N7804, N4094);
and AND3 (N7807, N7794, N3186, N4456);
buf BUF1 (N7808, N7802);
nor NOR3 (N7809, N7807, N7054, N7030);
buf BUF1 (N7810, N7783);
nor NOR3 (N7811, N7788, N5456, N7071);
nor NOR3 (N7812, N7810, N6055, N1558);
buf BUF1 (N7813, N7806);
not NOT1 (N7814, N7809);
xor XOR2 (N7815, N7813, N1814);
or OR4 (N7816, N7814, N2002, N1029, N7813);
and AND3 (N7817, N7815, N5029, N7587);
xor XOR2 (N7818, N7808, N7344);
nand NAND2 (N7819, N7797, N2706);
and AND4 (N7820, N7796, N2642, N3851, N4972);
buf BUF1 (N7821, N7819);
xor XOR2 (N7822, N7812, N5132);
or OR2 (N7823, N7817, N2465);
or OR3 (N7824, N7818, N3075, N5609);
buf BUF1 (N7825, N7820);
buf BUF1 (N7826, N7823);
not NOT1 (N7827, N7826);
or OR2 (N7828, N7824, N6126);
and AND2 (N7829, N7828, N3615);
and AND2 (N7830, N7822, N7703);
buf BUF1 (N7831, N7827);
not NOT1 (N7832, N7829);
xor XOR2 (N7833, N7825, N3174);
not NOT1 (N7834, N7831);
buf BUF1 (N7835, N7816);
and AND2 (N7836, N7830, N6610);
and AND3 (N7837, N7821, N397, N494);
xor XOR2 (N7838, N7803, N5131);
nand NAND2 (N7839, N7811, N2934);
nand NAND2 (N7840, N7793, N7538);
buf BUF1 (N7841, N7832);
not NOT1 (N7842, N7834);
nor NOR2 (N7843, N7805, N5527);
nor NOR4 (N7844, N7841, N7100, N4087, N6342);
not NOT1 (N7845, N7844);
xor XOR2 (N7846, N7835, N4323);
nand NAND3 (N7847, N7838, N729, N5031);
and AND2 (N7848, N7836, N5528);
buf BUF1 (N7849, N7837);
or OR4 (N7850, N7843, N7781, N4246, N1668);
nor NOR4 (N7851, N7847, N157, N5295, N443);
buf BUF1 (N7852, N7840);
nand NAND3 (N7853, N7848, N2567, N6229);
nand NAND4 (N7854, N7852, N3657, N3367, N1653);
nand NAND4 (N7855, N7839, N807, N4291, N5614);
xor XOR2 (N7856, N7851, N3578);
not NOT1 (N7857, N7850);
nand NAND3 (N7858, N7856, N3398, N3797);
buf BUF1 (N7859, N7842);
buf BUF1 (N7860, N7846);
and AND3 (N7861, N7860, N7762, N366);
buf BUF1 (N7862, N7853);
and AND4 (N7863, N7861, N6651, N7612, N2737);
not NOT1 (N7864, N7833);
nand NAND3 (N7865, N7854, N6314, N1306);
nand NAND4 (N7866, N7863, N5194, N6021, N39);
nand NAND3 (N7867, N7858, N914, N534);
buf BUF1 (N7868, N7866);
and AND2 (N7869, N7865, N7156);
or OR3 (N7870, N7869, N6382, N6066);
nor NOR3 (N7871, N7857, N4072, N838);
not NOT1 (N7872, N7868);
nor NOR4 (N7873, N7871, N3751, N2246, N7478);
xor XOR2 (N7874, N7859, N3726);
buf BUF1 (N7875, N7870);
xor XOR2 (N7876, N7875, N2302);
nand NAND2 (N7877, N7872, N7385);
or OR3 (N7878, N7874, N6573, N341);
buf BUF1 (N7879, N7876);
not NOT1 (N7880, N7849);
xor XOR2 (N7881, N7862, N4478);
xor XOR2 (N7882, N7880, N4658);
nor NOR2 (N7883, N7845, N7034);
nand NAND4 (N7884, N7878, N866, N3899, N6825);
xor XOR2 (N7885, N7867, N425);
xor XOR2 (N7886, N7879, N7828);
xor XOR2 (N7887, N7881, N5291);
xor XOR2 (N7888, N7883, N2756);
or OR3 (N7889, N7888, N7062, N3122);
nor NOR3 (N7890, N7873, N1207, N3347);
and AND2 (N7891, N7877, N4536);
nand NAND2 (N7892, N7864, N670);
buf BUF1 (N7893, N7891);
not NOT1 (N7894, N7892);
nor NOR2 (N7895, N7855, N4783);
nand NAND3 (N7896, N7895, N7651, N4162);
nor NOR3 (N7897, N7889, N4899, N6240);
xor XOR2 (N7898, N7896, N7155);
not NOT1 (N7899, N7887);
nand NAND4 (N7900, N7890, N3684, N6960, N1128);
xor XOR2 (N7901, N7894, N4855);
and AND4 (N7902, N7900, N274, N7053, N5526);
or OR4 (N7903, N7901, N1130, N3787, N4457);
and AND2 (N7904, N7899, N160);
not NOT1 (N7905, N7897);
and AND3 (N7906, N7905, N7239, N4600);
xor XOR2 (N7907, N7886, N5718);
nand NAND4 (N7908, N7884, N7723, N2112, N3476);
or OR4 (N7909, N7903, N2966, N57, N2321);
xor XOR2 (N7910, N7885, N2400);
buf BUF1 (N7911, N7908);
xor XOR2 (N7912, N7907, N6465);
or OR3 (N7913, N7909, N2658, N5793);
buf BUF1 (N7914, N7911);
xor XOR2 (N7915, N7912, N1226);
and AND4 (N7916, N7902, N7189, N1176, N5397);
nand NAND3 (N7917, N7906, N7707, N2259);
xor XOR2 (N7918, N7893, N4051);
buf BUF1 (N7919, N7914);
nand NAND3 (N7920, N7918, N2122, N4301);
xor XOR2 (N7921, N7898, N1407);
or OR3 (N7922, N7915, N5931, N1832);
or OR3 (N7923, N7904, N1333, N1108);
or OR3 (N7924, N7916, N902, N1030);
not NOT1 (N7925, N7913);
xor XOR2 (N7926, N7882, N5016);
nand NAND3 (N7927, N7919, N1125, N5462);
or OR4 (N7928, N7925, N6706, N98, N1773);
not NOT1 (N7929, N7924);
nand NAND4 (N7930, N7921, N5278, N2772, N6394);
and AND3 (N7931, N7922, N6765, N5637);
or OR2 (N7932, N7910, N4936);
nor NOR2 (N7933, N7923, N7632);
nand NAND2 (N7934, N7930, N2631);
buf BUF1 (N7935, N7932);
nor NOR3 (N7936, N7928, N7776, N7618);
nand NAND3 (N7937, N7935, N2186, N1874);
or OR3 (N7938, N7937, N2337, N664);
nand NAND2 (N7939, N7934, N4428);
not NOT1 (N7940, N7936);
and AND2 (N7941, N7939, N772);
nand NAND3 (N7942, N7940, N4801, N6403);
or OR2 (N7943, N7933, N4989);
buf BUF1 (N7944, N7929);
not NOT1 (N7945, N7931);
and AND3 (N7946, N7943, N6379, N3159);
or OR3 (N7947, N7941, N5055, N1887);
xor XOR2 (N7948, N7926, N3852);
or OR4 (N7949, N7945, N4621, N526, N6084);
nand NAND2 (N7950, N7917, N6093);
nand NAND4 (N7951, N7944, N932, N5764, N5561);
nor NOR2 (N7952, N7951, N3890);
and AND4 (N7953, N7949, N1916, N1347, N3002);
buf BUF1 (N7954, N7947);
not NOT1 (N7955, N7920);
nand NAND2 (N7956, N7952, N4960);
xor XOR2 (N7957, N7953, N633);
not NOT1 (N7958, N7927);
nor NOR3 (N7959, N7950, N133, N6248);
or OR3 (N7960, N7956, N1695, N3303);
buf BUF1 (N7961, N7938);
and AND2 (N7962, N7958, N2894);
xor XOR2 (N7963, N7942, N7391);
nor NOR2 (N7964, N7960, N1411);
nor NOR4 (N7965, N7948, N6945, N265, N3081);
nand NAND4 (N7966, N7963, N7950, N177, N7350);
and AND4 (N7967, N7955, N920, N6967, N1174);
xor XOR2 (N7968, N7946, N1749);
not NOT1 (N7969, N7954);
or OR3 (N7970, N7957, N2752, N1237);
nor NOR3 (N7971, N7959, N4627, N1127);
nor NOR4 (N7972, N7968, N7614, N7550, N203);
not NOT1 (N7973, N7965);
xor XOR2 (N7974, N7961, N6073);
xor XOR2 (N7975, N7972, N6117);
buf BUF1 (N7976, N7966);
or OR4 (N7977, N7964, N5934, N3718, N7780);
not NOT1 (N7978, N7975);
not NOT1 (N7979, N7974);
nand NAND2 (N7980, N7976, N6296);
nor NOR2 (N7981, N7973, N5291);
and AND2 (N7982, N7962, N474);
or OR3 (N7983, N7978, N301, N3636);
nand NAND3 (N7984, N7970, N2570, N3036);
and AND2 (N7985, N7981, N1982);
or OR4 (N7986, N7971, N1135, N7794, N7325);
nor NOR3 (N7987, N7985, N5402, N5833);
nand NAND3 (N7988, N7986, N4638, N1541);
nand NAND2 (N7989, N7979, N448);
and AND2 (N7990, N7989, N6584);
nor NOR4 (N7991, N7969, N1510, N6889, N7893);
buf BUF1 (N7992, N7988);
xor XOR2 (N7993, N7980, N2456);
nor NOR4 (N7994, N7993, N476, N6894, N6018);
not NOT1 (N7995, N7994);
nor NOR2 (N7996, N7991, N4129);
or OR3 (N7997, N7992, N5702, N4466);
buf BUF1 (N7998, N7987);
nor NOR3 (N7999, N7997, N2120, N1834);
nand NAND3 (N8000, N7977, N2546, N4067);
buf BUF1 (N8001, N8000);
xor XOR2 (N8002, N8001, N1531);
nor NOR2 (N8003, N7982, N275);
nand NAND2 (N8004, N7983, N1920);
and AND3 (N8005, N7967, N5191, N6080);
and AND4 (N8006, N8003, N1949, N690, N3428);
nand NAND4 (N8007, N8002, N728, N6480, N2802);
buf BUF1 (N8008, N7990);
buf BUF1 (N8009, N7995);
nand NAND3 (N8010, N8009, N4835, N2198);
nand NAND3 (N8011, N8010, N997, N2038);
xor XOR2 (N8012, N8011, N244);
xor XOR2 (N8013, N8006, N4588);
or OR3 (N8014, N7984, N5265, N5506);
not NOT1 (N8015, N8007);
xor XOR2 (N8016, N8004, N5855);
or OR2 (N8017, N8008, N2535);
xor XOR2 (N8018, N8015, N4624);
xor XOR2 (N8019, N7999, N5574);
xor XOR2 (N8020, N8017, N7398);
and AND3 (N8021, N8014, N4291, N7807);
not NOT1 (N8022, N7998);
or OR3 (N8023, N8020, N1959, N5369);
buf BUF1 (N8024, N8019);
or OR4 (N8025, N8013, N2879, N995, N1621);
nand NAND2 (N8026, N8012, N7013);
buf BUF1 (N8027, N8018);
xor XOR2 (N8028, N8021, N3363);
nor NOR3 (N8029, N7996, N632, N3770);
nor NOR2 (N8030, N8024, N5129);
buf BUF1 (N8031, N8023);
buf BUF1 (N8032, N8028);
and AND2 (N8033, N8029, N7618);
not NOT1 (N8034, N8032);
nand NAND3 (N8035, N8034, N4568, N2170);
nor NOR2 (N8036, N8035, N7388);
nand NAND3 (N8037, N8033, N4255, N7805);
nand NAND3 (N8038, N8022, N5588, N94);
not NOT1 (N8039, N8037);
and AND2 (N8040, N8016, N2373);
nand NAND3 (N8041, N8026, N1020, N35);
and AND2 (N8042, N8036, N7192);
and AND4 (N8043, N8038, N5807, N6611, N2529);
or OR3 (N8044, N8027, N2889, N7423);
or OR2 (N8045, N8030, N3835);
and AND4 (N8046, N8025, N5173, N4398, N5302);
or OR3 (N8047, N8031, N6232, N124);
buf BUF1 (N8048, N8005);
or OR3 (N8049, N8045, N4111, N4713);
not NOT1 (N8050, N8042);
nand NAND2 (N8051, N8039, N1620);
buf BUF1 (N8052, N8043);
nand NAND4 (N8053, N8041, N7941, N6604, N2263);
or OR3 (N8054, N8048, N5436, N5895);
nand NAND4 (N8055, N8052, N5512, N1419, N966);
nand NAND4 (N8056, N8040, N7082, N462, N2125);
not NOT1 (N8057, N8044);
nor NOR2 (N8058, N8046, N2546);
or OR4 (N8059, N8057, N5644, N4036, N4082);
and AND2 (N8060, N8049, N2239);
or OR4 (N8061, N8047, N2803, N4013, N4217);
or OR3 (N8062, N8056, N1055, N6399);
buf BUF1 (N8063, N8051);
nor NOR3 (N8064, N8050, N444, N1612);
xor XOR2 (N8065, N8064, N1120);
not NOT1 (N8066, N8055);
nor NOR3 (N8067, N8059, N3107, N3024);
nor NOR4 (N8068, N8062, N2544, N7272, N2329);
nor NOR2 (N8069, N8068, N7835);
buf BUF1 (N8070, N8054);
nor NOR2 (N8071, N8060, N2901);
nor NOR4 (N8072, N8065, N7854, N4963, N4883);
and AND4 (N8073, N8071, N6538, N7009, N678);
nand NAND3 (N8074, N8073, N1516, N1373);
buf BUF1 (N8075, N8070);
buf BUF1 (N8076, N8066);
nor NOR3 (N8077, N8072, N103, N5330);
xor XOR2 (N8078, N8069, N3488);
xor XOR2 (N8079, N8076, N2006);
or OR4 (N8080, N8063, N1024, N3614, N6210);
not NOT1 (N8081, N8080);
xor XOR2 (N8082, N8074, N3165);
and AND3 (N8083, N8067, N973, N5186);
and AND2 (N8084, N8077, N6050);
not NOT1 (N8085, N8084);
and AND3 (N8086, N8053, N3460, N4917);
not NOT1 (N8087, N8078);
nor NOR2 (N8088, N8082, N1957);
or OR4 (N8089, N8079, N2080, N3532, N7951);
buf BUF1 (N8090, N8089);
nor NOR4 (N8091, N8083, N7580, N6582, N3291);
or OR3 (N8092, N8081, N5353, N2876);
nor NOR4 (N8093, N8086, N3916, N5557, N6862);
or OR3 (N8094, N8093, N6390, N5527);
nand NAND4 (N8095, N8061, N6327, N5737, N7865);
not NOT1 (N8096, N8094);
nor NOR3 (N8097, N8075, N1844, N3880);
nor NOR3 (N8098, N8096, N6442, N5249);
not NOT1 (N8099, N8097);
nand NAND3 (N8100, N8099, N6291, N485);
and AND4 (N8101, N8088, N5488, N6980, N3458);
and AND3 (N8102, N8090, N2180, N4783);
buf BUF1 (N8103, N8058);
and AND2 (N8104, N8101, N2913);
xor XOR2 (N8105, N8100, N862);
not NOT1 (N8106, N8095);
buf BUF1 (N8107, N8085);
not NOT1 (N8108, N8106);
not NOT1 (N8109, N8087);
or OR4 (N8110, N8103, N5564, N6469, N5946);
nand NAND4 (N8111, N8102, N5709, N4898, N7020);
buf BUF1 (N8112, N8108);
nor NOR4 (N8113, N8109, N6456, N823, N1128);
not NOT1 (N8114, N8092);
nor NOR4 (N8115, N8104, N6521, N1237, N2595);
nor NOR3 (N8116, N8113, N5143, N2041);
not NOT1 (N8117, N8098);
buf BUF1 (N8118, N8091);
or OR4 (N8119, N8114, N3941, N5095, N3818);
buf BUF1 (N8120, N8110);
nand NAND3 (N8121, N8112, N7483, N1010);
not NOT1 (N8122, N8105);
and AND3 (N8123, N8117, N7459, N2565);
or OR4 (N8124, N8120, N1284, N6911, N1005);
and AND3 (N8125, N8123, N4190, N2078);
not NOT1 (N8126, N8122);
or OR2 (N8127, N8125, N1796);
not NOT1 (N8128, N8116);
buf BUF1 (N8129, N8118);
buf BUF1 (N8130, N8124);
nor NOR2 (N8131, N8121, N5301);
nand NAND2 (N8132, N8130, N868);
not NOT1 (N8133, N8129);
nor NOR3 (N8134, N8119, N5567, N3110);
buf BUF1 (N8135, N8134);
buf BUF1 (N8136, N8131);
not NOT1 (N8137, N8128);
buf BUF1 (N8138, N8127);
buf BUF1 (N8139, N8136);
and AND3 (N8140, N8132, N4300, N1280);
nor NOR4 (N8141, N8138, N1962, N4460, N7825);
not NOT1 (N8142, N8141);
not NOT1 (N8143, N8140);
nand NAND3 (N8144, N8133, N7380, N5024);
or OR2 (N8145, N8139, N4188);
nand NAND4 (N8146, N8126, N6989, N516, N3084);
not NOT1 (N8147, N8111);
not NOT1 (N8148, N8107);
nor NOR3 (N8149, N8115, N1051, N315);
not NOT1 (N8150, N8144);
xor XOR2 (N8151, N8146, N6412);
or OR3 (N8152, N8150, N432, N4901);
or OR3 (N8153, N8135, N7714, N1362);
buf BUF1 (N8154, N8153);
and AND2 (N8155, N8152, N6263);
and AND2 (N8156, N8148, N3936);
xor XOR2 (N8157, N8155, N1929);
nor NOR3 (N8158, N8143, N4167, N2353);
xor XOR2 (N8159, N8156, N6225);
not NOT1 (N8160, N8159);
or OR2 (N8161, N8154, N756);
xor XOR2 (N8162, N8158, N6106);
xor XOR2 (N8163, N8162, N3162);
xor XOR2 (N8164, N8149, N634);
nand NAND3 (N8165, N8137, N6990, N5032);
xor XOR2 (N8166, N8165, N2602);
and AND2 (N8167, N8145, N8012);
nor NOR3 (N8168, N8164, N5898, N6559);
or OR2 (N8169, N8147, N4980);
nor NOR4 (N8170, N8166, N6968, N2552, N841);
not NOT1 (N8171, N8169);
not NOT1 (N8172, N8171);
and AND4 (N8173, N8163, N5330, N7334, N5200);
or OR3 (N8174, N8170, N4767, N464);
nand NAND4 (N8175, N8168, N7927, N5707, N3556);
and AND2 (N8176, N8172, N2932);
xor XOR2 (N8177, N8174, N6419);
nand NAND3 (N8178, N8175, N1434, N7468);
not NOT1 (N8179, N8160);
not NOT1 (N8180, N8173);
and AND2 (N8181, N8142, N5469);
and AND4 (N8182, N8151, N4252, N3462, N2762);
nand NAND2 (N8183, N8177, N1498);
and AND4 (N8184, N8161, N3269, N6176, N8061);
buf BUF1 (N8185, N8183);
xor XOR2 (N8186, N8185, N1594);
not NOT1 (N8187, N8182);
not NOT1 (N8188, N8157);
nand NAND3 (N8189, N8186, N135, N6568);
nor NOR4 (N8190, N8179, N1762, N325, N5892);
nand NAND2 (N8191, N8189, N7722);
xor XOR2 (N8192, N8184, N711);
nor NOR4 (N8193, N8191, N6650, N2371, N6148);
and AND2 (N8194, N8192, N7310);
nand NAND3 (N8195, N8190, N5771, N3960);
buf BUF1 (N8196, N8180);
and AND4 (N8197, N8178, N5911, N6371, N7341);
nand NAND3 (N8198, N8195, N1120, N6963);
buf BUF1 (N8199, N8198);
buf BUF1 (N8200, N8196);
xor XOR2 (N8201, N8197, N3196);
and AND3 (N8202, N8201, N1649, N1472);
nor NOR3 (N8203, N8193, N4822, N6947);
or OR4 (N8204, N8199, N1470, N2355, N2312);
nand NAND2 (N8205, N8203, N5482);
or OR4 (N8206, N8167, N7341, N5023, N6171);
xor XOR2 (N8207, N8176, N1172);
nor NOR4 (N8208, N8181, N7292, N7681, N6798);
buf BUF1 (N8209, N8188);
buf BUF1 (N8210, N8209);
or OR4 (N8211, N8207, N8022, N8169, N552);
not NOT1 (N8212, N8194);
buf BUF1 (N8213, N8205);
or OR3 (N8214, N8187, N3102, N4434);
nand NAND4 (N8215, N8200, N7626, N5207, N4754);
xor XOR2 (N8216, N8208, N6019);
and AND4 (N8217, N8210, N7451, N7296, N4340);
or OR4 (N8218, N8216, N3731, N3479, N4061);
or OR2 (N8219, N8214, N5060);
xor XOR2 (N8220, N8218, N6683);
not NOT1 (N8221, N8219);
or OR3 (N8222, N8212, N6864, N4448);
nand NAND4 (N8223, N8220, N4168, N7946, N5615);
buf BUF1 (N8224, N8223);
xor XOR2 (N8225, N8202, N7729);
and AND3 (N8226, N8222, N2047, N7599);
xor XOR2 (N8227, N8204, N3250);
nor NOR3 (N8228, N8225, N6472, N4394);
or OR4 (N8229, N8224, N6564, N3459, N8131);
not NOT1 (N8230, N8221);
nand NAND2 (N8231, N8217, N3331);
or OR3 (N8232, N8226, N1160, N7244);
and AND3 (N8233, N8227, N434, N3653);
nor NOR3 (N8234, N8230, N1461, N6240);
not NOT1 (N8235, N8211);
xor XOR2 (N8236, N8206, N8079);
or OR4 (N8237, N8235, N6946, N1513, N5625);
buf BUF1 (N8238, N8234);
and AND3 (N8239, N8229, N3639, N3969);
buf BUF1 (N8240, N8238);
or OR3 (N8241, N8231, N2463, N2839);
and AND2 (N8242, N8213, N4926);
buf BUF1 (N8243, N8239);
buf BUF1 (N8244, N8242);
nor NOR3 (N8245, N8236, N5756, N3261);
nand NAND2 (N8246, N8237, N2505);
not NOT1 (N8247, N8228);
buf BUF1 (N8248, N8240);
nand NAND2 (N8249, N8246, N4151);
nand NAND3 (N8250, N8248, N2295, N3331);
and AND3 (N8251, N8233, N2277, N3529);
nand NAND2 (N8252, N8241, N5968);
nor NOR2 (N8253, N8215, N5887);
nand NAND4 (N8254, N8244, N243, N7347, N2408);
not NOT1 (N8255, N8252);
and AND3 (N8256, N8253, N8171, N2471);
and AND3 (N8257, N8245, N6624, N3291);
nor NOR3 (N8258, N8247, N94, N2331);
buf BUF1 (N8259, N8258);
xor XOR2 (N8260, N8254, N3821);
xor XOR2 (N8261, N8249, N5644);
buf BUF1 (N8262, N8259);
not NOT1 (N8263, N8250);
nor NOR2 (N8264, N8243, N2690);
and AND2 (N8265, N8263, N7235);
nand NAND4 (N8266, N8265, N365, N7084, N3590);
or OR3 (N8267, N8257, N3588, N3012);
nand NAND3 (N8268, N8261, N4340, N3033);
nor NOR4 (N8269, N8255, N6897, N2967, N4841);
nor NOR2 (N8270, N8266, N3730);
not NOT1 (N8271, N8262);
xor XOR2 (N8272, N8267, N4459);
nor NOR3 (N8273, N8260, N1767, N6228);
buf BUF1 (N8274, N8271);
nand NAND3 (N8275, N8268, N7268, N3621);
buf BUF1 (N8276, N8275);
not NOT1 (N8277, N8273);
not NOT1 (N8278, N8270);
or OR3 (N8279, N8264, N5829, N6803);
nor NOR4 (N8280, N8276, N8265, N3687, N2230);
buf BUF1 (N8281, N8256);
nand NAND2 (N8282, N8281, N5468);
nand NAND3 (N8283, N8278, N3138, N2615);
and AND2 (N8284, N8277, N681);
buf BUF1 (N8285, N8269);
xor XOR2 (N8286, N8274, N3735);
and AND2 (N8287, N8232, N1615);
buf BUF1 (N8288, N8284);
buf BUF1 (N8289, N8280);
and AND4 (N8290, N8285, N5631, N4794, N40);
nand NAND2 (N8291, N8290, N696);
nand NAND4 (N8292, N8288, N5549, N4216, N6256);
buf BUF1 (N8293, N8286);
and AND2 (N8294, N8291, N1634);
and AND2 (N8295, N8294, N5762);
nand NAND3 (N8296, N8287, N4666, N8038);
nand NAND3 (N8297, N8289, N1330, N582);
xor XOR2 (N8298, N8295, N3748);
nor NOR4 (N8299, N8292, N1827, N2106, N4066);
nand NAND2 (N8300, N8297, N6430);
or OR4 (N8301, N8296, N4466, N2390, N3244);
nand NAND3 (N8302, N8300, N7629, N6650);
xor XOR2 (N8303, N8251, N5890);
and AND4 (N8304, N8283, N2153, N2645, N5058);
and AND3 (N8305, N8302, N4968, N6161);
not NOT1 (N8306, N8305);
not NOT1 (N8307, N8298);
or OR2 (N8308, N8299, N2271);
xor XOR2 (N8309, N8293, N2513);
not NOT1 (N8310, N8304);
or OR4 (N8311, N8310, N2080, N6070, N8085);
xor XOR2 (N8312, N8308, N2203);
and AND4 (N8313, N8303, N5874, N3736, N3747);
nor NOR2 (N8314, N8279, N954);
not NOT1 (N8315, N8307);
buf BUF1 (N8316, N8272);
or OR2 (N8317, N8311, N7409);
nand NAND2 (N8318, N8282, N3215);
or OR3 (N8319, N8312, N7615, N6551);
nand NAND3 (N8320, N8318, N153, N2659);
not NOT1 (N8321, N8306);
not NOT1 (N8322, N8314);
and AND3 (N8323, N8322, N4635, N3368);
xor XOR2 (N8324, N8301, N1875);
nand NAND4 (N8325, N8321, N6485, N6108, N3353);
xor XOR2 (N8326, N8309, N6434);
nor NOR3 (N8327, N8326, N5330, N3193);
xor XOR2 (N8328, N8317, N5329);
xor XOR2 (N8329, N8328, N4832);
and AND3 (N8330, N8324, N2440, N7439);
not NOT1 (N8331, N8329);
xor XOR2 (N8332, N8313, N902);
nand NAND4 (N8333, N8320, N6777, N4804, N1385);
xor XOR2 (N8334, N8330, N3327);
nor NOR3 (N8335, N8315, N2996, N980);
xor XOR2 (N8336, N8331, N2908);
not NOT1 (N8337, N8327);
nor NOR3 (N8338, N8333, N6237, N6217);
or OR4 (N8339, N8335, N3787, N2943, N7091);
and AND2 (N8340, N8323, N2574);
and AND3 (N8341, N8339, N6649, N450);
buf BUF1 (N8342, N8325);
nand NAND4 (N8343, N8319, N390, N883, N7594);
nand NAND2 (N8344, N8341, N3008);
xor XOR2 (N8345, N8344, N7648);
or OR3 (N8346, N8337, N1379, N2669);
xor XOR2 (N8347, N8334, N5221);
or OR4 (N8348, N8346, N3432, N2070, N5466);
buf BUF1 (N8349, N8348);
xor XOR2 (N8350, N8316, N7473);
and AND2 (N8351, N8332, N3539);
and AND3 (N8352, N8340, N2866, N1227);
nand NAND4 (N8353, N8349, N4273, N2673, N3698);
not NOT1 (N8354, N8345);
nor NOR4 (N8355, N8347, N5829, N7436, N2989);
or OR3 (N8356, N8342, N8048, N1460);
xor XOR2 (N8357, N8350, N2680);
and AND2 (N8358, N8351, N3168);
not NOT1 (N8359, N8336);
xor XOR2 (N8360, N8343, N2402);
and AND3 (N8361, N8360, N6641, N3251);
nor NOR3 (N8362, N8358, N975, N3044);
and AND3 (N8363, N8357, N844, N2423);
not NOT1 (N8364, N8363);
buf BUF1 (N8365, N8364);
nand NAND2 (N8366, N8353, N1646);
not NOT1 (N8367, N8355);
nand NAND3 (N8368, N8365, N3751, N60);
not NOT1 (N8369, N8352);
and AND4 (N8370, N8368, N4254, N4263, N2046);
and AND3 (N8371, N8361, N5611, N5097);
and AND2 (N8372, N8366, N445);
not NOT1 (N8373, N8369);
xor XOR2 (N8374, N8372, N4165);
or OR4 (N8375, N8370, N304, N3179, N5524);
xor XOR2 (N8376, N8375, N1014);
buf BUF1 (N8377, N8354);
nor NOR3 (N8378, N8377, N7711, N2554);
xor XOR2 (N8379, N8371, N1925);
and AND3 (N8380, N8379, N2677, N1210);
buf BUF1 (N8381, N8338);
xor XOR2 (N8382, N8362, N2815);
buf BUF1 (N8383, N8378);
nor NOR3 (N8384, N8376, N8007, N2821);
xor XOR2 (N8385, N8373, N6092);
nand NAND2 (N8386, N8367, N5727);
or OR3 (N8387, N8374, N567, N7171);
nand NAND4 (N8388, N8387, N776, N6431, N3406);
buf BUF1 (N8389, N8359);
nor NOR4 (N8390, N8385, N275, N5436, N5608);
xor XOR2 (N8391, N8380, N478);
and AND3 (N8392, N8390, N4039, N3017);
buf BUF1 (N8393, N8389);
and AND2 (N8394, N8393, N5119);
nor NOR2 (N8395, N8384, N3317);
and AND3 (N8396, N8391, N4261, N2399);
xor XOR2 (N8397, N8392, N6912);
or OR4 (N8398, N8396, N6174, N57, N7072);
or OR4 (N8399, N8395, N5496, N7623, N3132);
and AND3 (N8400, N8381, N3440, N265);
or OR2 (N8401, N8397, N8087);
buf BUF1 (N8402, N8401);
not NOT1 (N8403, N8394);
or OR3 (N8404, N8386, N7794, N8070);
not NOT1 (N8405, N8388);
nor NOR3 (N8406, N8405, N21, N8379);
or OR3 (N8407, N8404, N4745, N1085);
not NOT1 (N8408, N8400);
not NOT1 (N8409, N8402);
or OR4 (N8410, N8409, N6602, N1064, N7255);
nand NAND4 (N8411, N8403, N684, N7945, N765);
nor NOR2 (N8412, N8356, N2270);
buf BUF1 (N8413, N8382);
nor NOR3 (N8414, N8410, N2256, N522);
nand NAND4 (N8415, N8414, N821, N4553, N1719);
xor XOR2 (N8416, N8411, N7323);
xor XOR2 (N8417, N8406, N7322);
xor XOR2 (N8418, N8415, N1591);
buf BUF1 (N8419, N8417);
xor XOR2 (N8420, N8416, N4689);
buf BUF1 (N8421, N8412);
or OR2 (N8422, N8413, N2806);
buf BUF1 (N8423, N8398);
nand NAND2 (N8424, N8383, N4899);
and AND2 (N8425, N8421, N958);
and AND4 (N8426, N8418, N2392, N4268, N4601);
buf BUF1 (N8427, N8423);
nor NOR2 (N8428, N8422, N586);
nor NOR3 (N8429, N8420, N723, N3060);
or OR2 (N8430, N8427, N8219);
xor XOR2 (N8431, N8407, N6163);
not NOT1 (N8432, N8424);
not NOT1 (N8433, N8431);
nand NAND4 (N8434, N8408, N1979, N3660, N2929);
xor XOR2 (N8435, N8429, N73);
nor NOR2 (N8436, N8434, N71);
not NOT1 (N8437, N8432);
and AND4 (N8438, N8419, N2638, N7917, N6675);
nor NOR4 (N8439, N8433, N1128, N1324, N2319);
nand NAND4 (N8440, N8436, N7788, N8023, N945);
and AND2 (N8441, N8438, N696);
xor XOR2 (N8442, N8440, N498);
and AND2 (N8443, N8426, N3175);
nand NAND2 (N8444, N8443, N6406);
not NOT1 (N8445, N8428);
buf BUF1 (N8446, N8445);
buf BUF1 (N8447, N8439);
nand NAND4 (N8448, N8442, N2874, N8122, N4043);
buf BUF1 (N8449, N8441);
nand NAND4 (N8450, N8435, N1996, N7777, N2215);
and AND3 (N8451, N8450, N6179, N5501);
nand NAND2 (N8452, N8446, N8051);
nor NOR4 (N8453, N8444, N7448, N7125, N8139);
not NOT1 (N8454, N8447);
and AND3 (N8455, N8448, N4037, N2966);
or OR4 (N8456, N8437, N7593, N15, N8158);
buf BUF1 (N8457, N8453);
nor NOR3 (N8458, N8457, N8220, N8248);
not NOT1 (N8459, N8456);
nor NOR4 (N8460, N8449, N7286, N1628, N3203);
nor NOR2 (N8461, N8458, N3352);
buf BUF1 (N8462, N8430);
and AND2 (N8463, N8455, N371);
xor XOR2 (N8464, N8451, N1893);
xor XOR2 (N8465, N8452, N1354);
xor XOR2 (N8466, N8460, N1208);
buf BUF1 (N8467, N8464);
xor XOR2 (N8468, N8461, N2528);
or OR3 (N8469, N8466, N5550, N718);
xor XOR2 (N8470, N8462, N6233);
nand NAND3 (N8471, N8465, N8444, N1507);
and AND4 (N8472, N8399, N7769, N6098, N6153);
and AND3 (N8473, N8472, N7586, N1133);
xor XOR2 (N8474, N8467, N3631);
buf BUF1 (N8475, N8469);
or OR2 (N8476, N8468, N7752);
not NOT1 (N8477, N8475);
nand NAND3 (N8478, N8470, N6913, N4685);
buf BUF1 (N8479, N8454);
xor XOR2 (N8480, N8478, N950);
nor NOR4 (N8481, N8473, N3250, N2001, N4235);
not NOT1 (N8482, N8474);
and AND3 (N8483, N8471, N3570, N7712);
buf BUF1 (N8484, N8483);
nor NOR3 (N8485, N8480, N6252, N7928);
nand NAND2 (N8486, N8485, N3589);
or OR3 (N8487, N8459, N4968, N2260);
nor NOR4 (N8488, N8481, N3644, N3501, N3916);
and AND4 (N8489, N8484, N5538, N6928, N4456);
nor NOR4 (N8490, N8488, N4186, N1626, N7900);
nor NOR4 (N8491, N8477, N261, N6424, N5263);
and AND4 (N8492, N8491, N3334, N1771, N3628);
buf BUF1 (N8493, N8482);
buf BUF1 (N8494, N8492);
or OR2 (N8495, N8490, N3947);
buf BUF1 (N8496, N8493);
buf BUF1 (N8497, N8487);
and AND3 (N8498, N8495, N8206, N2120);
buf BUF1 (N8499, N8489);
and AND2 (N8500, N8496, N2108);
and AND3 (N8501, N8463, N1580, N7676);
not NOT1 (N8502, N8479);
nor NOR3 (N8503, N8501, N1182, N2973);
buf BUF1 (N8504, N8486);
nand NAND2 (N8505, N8503, N113);
nor NOR4 (N8506, N8499, N5344, N5069, N7941);
xor XOR2 (N8507, N8500, N849);
nand NAND4 (N8508, N8504, N1114, N3259, N7182);
nor NOR2 (N8509, N8502, N4494);
or OR3 (N8510, N8509, N8134, N4909);
buf BUF1 (N8511, N8425);
xor XOR2 (N8512, N8494, N4608);
and AND2 (N8513, N8508, N6590);
not NOT1 (N8514, N8511);
buf BUF1 (N8515, N8507);
and AND3 (N8516, N8505, N8190, N1520);
nand NAND2 (N8517, N8515, N3606);
xor XOR2 (N8518, N8476, N6819);
buf BUF1 (N8519, N8498);
nand NAND2 (N8520, N8510, N5545);
nand NAND3 (N8521, N8497, N3785, N1676);
nand NAND3 (N8522, N8517, N5945, N5297);
buf BUF1 (N8523, N8512);
buf BUF1 (N8524, N8513);
buf BUF1 (N8525, N8522);
nor NOR4 (N8526, N8525, N4872, N2250, N8408);
buf BUF1 (N8527, N8519);
and AND3 (N8528, N8516, N3720, N3558);
and AND3 (N8529, N8518, N4207, N6832);
not NOT1 (N8530, N8526);
nor NOR2 (N8531, N8506, N5984);
or OR2 (N8532, N8523, N5565);
xor XOR2 (N8533, N8521, N1522);
and AND4 (N8534, N8524, N6163, N5305, N2983);
or OR2 (N8535, N8529, N7325);
buf BUF1 (N8536, N8520);
xor XOR2 (N8537, N8531, N1627);
and AND3 (N8538, N8527, N3065, N1090);
and AND2 (N8539, N8537, N2351);
and AND3 (N8540, N8534, N1490, N5684);
or OR4 (N8541, N8528, N1272, N2876, N1271);
not NOT1 (N8542, N8536);
and AND2 (N8543, N8538, N3960);
or OR3 (N8544, N8543, N8407, N4462);
nor NOR3 (N8545, N8514, N260, N702);
and AND4 (N8546, N8539, N7975, N4656, N1273);
buf BUF1 (N8547, N8545);
or OR2 (N8548, N8533, N5037);
nor NOR4 (N8549, N8546, N5786, N2238, N5068);
or OR4 (N8550, N8530, N550, N164, N7683);
or OR3 (N8551, N8542, N4581, N5004);
or OR4 (N8552, N8548, N7082, N8530, N2963);
and AND4 (N8553, N8550, N6768, N7353, N4749);
buf BUF1 (N8554, N8535);
buf BUF1 (N8555, N8554);
xor XOR2 (N8556, N8549, N1687);
buf BUF1 (N8557, N8544);
nand NAND3 (N8558, N8547, N4740, N4612);
or OR3 (N8559, N8552, N6848, N4924);
and AND2 (N8560, N8559, N182);
and AND2 (N8561, N8560, N3067);
and AND3 (N8562, N8551, N7369, N5355);
nor NOR4 (N8563, N8557, N4736, N6009, N7218);
nand NAND4 (N8564, N8556, N8087, N4337, N3120);
not NOT1 (N8565, N8564);
nor NOR3 (N8566, N8562, N8138, N7496);
not NOT1 (N8567, N8555);
and AND3 (N8568, N8532, N1042, N5608);
xor XOR2 (N8569, N8553, N5704);
buf BUF1 (N8570, N8561);
and AND4 (N8571, N8565, N5006, N5426, N2339);
and AND2 (N8572, N8558, N1863);
or OR4 (N8573, N8568, N7127, N7152, N1832);
or OR3 (N8574, N8541, N7081, N8143);
buf BUF1 (N8575, N8571);
xor XOR2 (N8576, N8567, N4375);
xor XOR2 (N8577, N8575, N8026);
buf BUF1 (N8578, N8572);
buf BUF1 (N8579, N8570);
or OR2 (N8580, N8569, N4881);
xor XOR2 (N8581, N8580, N8350);
xor XOR2 (N8582, N8574, N2896);
nand NAND4 (N8583, N8577, N15, N5147, N6545);
nor NOR3 (N8584, N8581, N1593, N3787);
nor NOR3 (N8585, N8540, N4390, N6222);
nor NOR4 (N8586, N8582, N2181, N4933, N7413);
and AND2 (N8587, N8585, N2412);
xor XOR2 (N8588, N8579, N7745);
nand NAND3 (N8589, N8587, N802, N610);
and AND4 (N8590, N8589, N5101, N4467, N1449);
and AND3 (N8591, N8578, N3318, N7177);
not NOT1 (N8592, N8584);
nand NAND3 (N8593, N8586, N413, N5018);
buf BUF1 (N8594, N8576);
not NOT1 (N8595, N8594);
xor XOR2 (N8596, N8583, N3466);
or OR3 (N8597, N8588, N7340, N1351);
or OR2 (N8598, N8597, N4537);
buf BUF1 (N8599, N8573);
not NOT1 (N8600, N8566);
nor NOR4 (N8601, N8593, N6245, N3772, N1440);
nor NOR4 (N8602, N8598, N8446, N4177, N63);
buf BUF1 (N8603, N8592);
nor NOR3 (N8604, N8591, N7118, N7847);
xor XOR2 (N8605, N8590, N720);
nand NAND3 (N8606, N8605, N2796, N1253);
nand NAND2 (N8607, N8606, N7466);
xor XOR2 (N8608, N8563, N8440);
not NOT1 (N8609, N8601);
buf BUF1 (N8610, N8596);
or OR3 (N8611, N8610, N2142, N1501);
and AND2 (N8612, N8604, N2952);
xor XOR2 (N8613, N8600, N6441);
and AND4 (N8614, N8602, N6838, N5336, N2248);
and AND2 (N8615, N8608, N1677);
and AND4 (N8616, N8611, N3053, N2275, N3201);
or OR4 (N8617, N8615, N6012, N2364, N2305);
and AND4 (N8618, N8603, N7085, N7434, N4751);
xor XOR2 (N8619, N8616, N2439);
xor XOR2 (N8620, N8599, N4990);
and AND4 (N8621, N8613, N48, N2461, N3236);
nand NAND3 (N8622, N8614, N7170, N4998);
xor XOR2 (N8623, N8622, N1614);
and AND3 (N8624, N8619, N3046, N346);
xor XOR2 (N8625, N8620, N1766);
nor NOR4 (N8626, N8621, N469, N6617, N3808);
xor XOR2 (N8627, N8595, N737);
and AND2 (N8628, N8627, N2064);
buf BUF1 (N8629, N8626);
not NOT1 (N8630, N8607);
nand NAND4 (N8631, N8628, N3979, N5621, N178);
nand NAND2 (N8632, N8630, N1608);
xor XOR2 (N8633, N8618, N8171);
or OR3 (N8634, N8629, N7047, N4896);
xor XOR2 (N8635, N8623, N5541);
not NOT1 (N8636, N8633);
and AND2 (N8637, N8631, N8564);
nor NOR4 (N8638, N8632, N3172, N6221, N4316);
and AND2 (N8639, N8617, N1080);
buf BUF1 (N8640, N8612);
and AND4 (N8641, N8624, N883, N7964, N3435);
or OR3 (N8642, N8625, N7696, N2748);
not NOT1 (N8643, N8642);
nand NAND3 (N8644, N8640, N7258, N2002);
or OR3 (N8645, N8636, N5437, N7687);
buf BUF1 (N8646, N8634);
xor XOR2 (N8647, N8646, N2129);
buf BUF1 (N8648, N8645);
nor NOR4 (N8649, N8647, N8158, N2960, N1854);
or OR3 (N8650, N8641, N4196, N5484);
or OR4 (N8651, N8644, N273, N7670, N6792);
not NOT1 (N8652, N8649);
and AND4 (N8653, N8643, N3832, N5799, N8108);
nand NAND3 (N8654, N8609, N5662, N6896);
not NOT1 (N8655, N8652);
xor XOR2 (N8656, N8635, N7198);
buf BUF1 (N8657, N8654);
and AND3 (N8658, N8638, N422, N8038);
nor NOR3 (N8659, N8657, N166, N3011);
and AND2 (N8660, N8639, N975);
or OR2 (N8661, N8655, N8652);
xor XOR2 (N8662, N8660, N6948);
buf BUF1 (N8663, N8661);
nand NAND4 (N8664, N8650, N8399, N2858, N6493);
and AND2 (N8665, N8663, N4399);
nand NAND3 (N8666, N8662, N3442, N205);
or OR3 (N8667, N8648, N7069, N8570);
xor XOR2 (N8668, N8653, N4563);
or OR3 (N8669, N8666, N6837, N177);
and AND2 (N8670, N8637, N4232);
and AND2 (N8671, N8651, N8399);
nor NOR3 (N8672, N8669, N79, N1562);
nor NOR3 (N8673, N8668, N7661, N6693);
and AND2 (N8674, N8671, N3351);
nor NOR4 (N8675, N8656, N5683, N2867, N4753);
and AND2 (N8676, N8673, N3735);
or OR3 (N8677, N8675, N3082, N7049);
not NOT1 (N8678, N8664);
xor XOR2 (N8679, N8678, N3139);
xor XOR2 (N8680, N8674, N4247);
nand NAND4 (N8681, N8677, N980, N4459, N1536);
nor NOR3 (N8682, N8670, N6958, N4937);
xor XOR2 (N8683, N8679, N7206);
or OR3 (N8684, N8672, N2568, N2148);
not NOT1 (N8685, N8676);
or OR3 (N8686, N8658, N8233, N657);
xor XOR2 (N8687, N8659, N2307);
or OR3 (N8688, N8681, N3776, N8290);
and AND4 (N8689, N8665, N2414, N4556, N6698);
nor NOR3 (N8690, N8683, N2386, N7020);
or OR3 (N8691, N8667, N1713, N6886);
and AND4 (N8692, N8688, N2078, N4034, N7265);
xor XOR2 (N8693, N8682, N4715);
xor XOR2 (N8694, N8680, N7492);
xor XOR2 (N8695, N8694, N4305);
buf BUF1 (N8696, N8692);
and AND2 (N8697, N8689, N7912);
and AND3 (N8698, N8685, N8424, N6247);
xor XOR2 (N8699, N8698, N8280);
not NOT1 (N8700, N8697);
buf BUF1 (N8701, N8699);
and AND3 (N8702, N8687, N5651, N5029);
nand NAND2 (N8703, N8693, N7186);
xor XOR2 (N8704, N8690, N1101);
and AND2 (N8705, N8686, N1286);
buf BUF1 (N8706, N8704);
nand NAND3 (N8707, N8705, N3898, N8424);
not NOT1 (N8708, N8695);
or OR3 (N8709, N8684, N5088, N5642);
not NOT1 (N8710, N8703);
buf BUF1 (N8711, N8708);
not NOT1 (N8712, N8701);
buf BUF1 (N8713, N8700);
and AND3 (N8714, N8710, N6475, N5324);
xor XOR2 (N8715, N8706, N8549);
buf BUF1 (N8716, N8707);
and AND3 (N8717, N8715, N6348, N6528);
nand NAND2 (N8718, N8702, N4129);
not NOT1 (N8719, N8711);
not NOT1 (N8720, N8719);
nor NOR4 (N8721, N8713, N5054, N2806, N239);
nor NOR4 (N8722, N8717, N6019, N6463, N2293);
nor NOR2 (N8723, N8716, N4933);
and AND4 (N8724, N8720, N8150, N6793, N1244);
not NOT1 (N8725, N8724);
not NOT1 (N8726, N8696);
buf BUF1 (N8727, N8691);
not NOT1 (N8728, N8727);
xor XOR2 (N8729, N8726, N4571);
and AND3 (N8730, N8729, N3638, N6598);
xor XOR2 (N8731, N8728, N6407);
or OR3 (N8732, N8721, N4575, N3982);
and AND2 (N8733, N8718, N3994);
nor NOR2 (N8734, N8731, N8576);
xor XOR2 (N8735, N8714, N3572);
or OR3 (N8736, N8723, N821, N6443);
or OR4 (N8737, N8732, N150, N6893, N4235);
and AND3 (N8738, N8709, N964, N5345);
not NOT1 (N8739, N8737);
and AND3 (N8740, N8722, N5704, N1705);
buf BUF1 (N8741, N8736);
and AND4 (N8742, N8725, N4850, N4800, N7689);
and AND3 (N8743, N8730, N7459, N914);
buf BUF1 (N8744, N8738);
xor XOR2 (N8745, N8742, N3370);
or OR2 (N8746, N8741, N481);
nor NOR2 (N8747, N8744, N2942);
or OR3 (N8748, N8747, N6745, N6495);
nor NOR4 (N8749, N8739, N5144, N964, N7733);
not NOT1 (N8750, N8745);
xor XOR2 (N8751, N8735, N3983);
xor XOR2 (N8752, N8751, N3275);
and AND3 (N8753, N8746, N6637, N4472);
xor XOR2 (N8754, N8750, N1505);
and AND4 (N8755, N8749, N1166, N5104, N110);
not NOT1 (N8756, N8712);
nand NAND4 (N8757, N8754, N708, N5157, N6546);
nand NAND4 (N8758, N8756, N2960, N4048, N6815);
buf BUF1 (N8759, N8748);
xor XOR2 (N8760, N8740, N3052);
buf BUF1 (N8761, N8753);
nand NAND2 (N8762, N8759, N7393);
and AND3 (N8763, N8761, N4464, N4697);
nor NOR4 (N8764, N8755, N194, N6577, N1672);
and AND3 (N8765, N8743, N2949, N1563);
and AND4 (N8766, N8757, N8725, N5104, N5779);
nor NOR4 (N8767, N8734, N925, N2596, N3147);
xor XOR2 (N8768, N8766, N6880);
nand NAND3 (N8769, N8764, N7116, N6593);
nor NOR4 (N8770, N8752, N8109, N2003, N6014);
buf BUF1 (N8771, N8763);
xor XOR2 (N8772, N8767, N5059);
xor XOR2 (N8773, N8769, N229);
xor XOR2 (N8774, N8733, N5270);
nand NAND2 (N8775, N8762, N7582);
nand NAND4 (N8776, N8760, N6405, N1621, N1246);
nor NOR3 (N8777, N8771, N6173, N4063);
nor NOR4 (N8778, N8776, N8358, N3571, N3255);
and AND4 (N8779, N8758, N3469, N4339, N7400);
buf BUF1 (N8780, N8778);
and AND3 (N8781, N8772, N5147, N7815);
and AND2 (N8782, N8768, N2391);
xor XOR2 (N8783, N8765, N3723);
nor NOR4 (N8784, N8770, N6877, N274, N4330);
or OR2 (N8785, N8780, N50);
nor NOR2 (N8786, N8782, N6395);
or OR2 (N8787, N8784, N1128);
buf BUF1 (N8788, N8774);
or OR4 (N8789, N8786, N8441, N4820, N2575);
or OR2 (N8790, N8788, N6958);
and AND3 (N8791, N8789, N4524, N2266);
xor XOR2 (N8792, N8775, N8333);
or OR4 (N8793, N8781, N1917, N3422, N8492);
xor XOR2 (N8794, N8773, N1569);
buf BUF1 (N8795, N8791);
buf BUF1 (N8796, N8793);
not NOT1 (N8797, N8790);
and AND4 (N8798, N8787, N7082, N3526, N5462);
nand NAND3 (N8799, N8779, N4540, N5402);
nor NOR2 (N8800, N8783, N3941);
nor NOR2 (N8801, N8798, N7637);
nor NOR4 (N8802, N8785, N2512, N8028, N7873);
and AND4 (N8803, N8796, N3799, N5974, N4672);
xor XOR2 (N8804, N8792, N5391);
nor NOR2 (N8805, N8795, N8361);
or OR2 (N8806, N8803, N219);
not NOT1 (N8807, N8799);
not NOT1 (N8808, N8801);
not NOT1 (N8809, N8777);
buf BUF1 (N8810, N8809);
and AND3 (N8811, N8802, N3887, N2339);
not NOT1 (N8812, N8811);
not NOT1 (N8813, N8807);
and AND3 (N8814, N8794, N2444, N1214);
nand NAND3 (N8815, N8797, N4220, N4121);
nor NOR3 (N8816, N8813, N4445, N2523);
buf BUF1 (N8817, N8816);
and AND4 (N8818, N8812, N3657, N5572, N3267);
or OR3 (N8819, N8817, N5195, N498);
nand NAND2 (N8820, N8818, N855);
or OR2 (N8821, N8810, N4678);
or OR3 (N8822, N8821, N1920, N3300);
not NOT1 (N8823, N8808);
buf BUF1 (N8824, N8805);
and AND3 (N8825, N8814, N4260, N2510);
nand NAND3 (N8826, N8824, N8670, N5318);
xor XOR2 (N8827, N8806, N4764);
or OR3 (N8828, N8800, N888, N5195);
nand NAND4 (N8829, N8826, N5152, N6001, N7458);
nand NAND4 (N8830, N8819, N1351, N6734, N5109);
nor NOR3 (N8831, N8815, N4635, N927);
not NOT1 (N8832, N8829);
nor NOR4 (N8833, N8823, N7246, N7645, N6363);
or OR3 (N8834, N8830, N4335, N6656);
not NOT1 (N8835, N8831);
buf BUF1 (N8836, N8832);
buf BUF1 (N8837, N8822);
xor XOR2 (N8838, N8834, N1331);
not NOT1 (N8839, N8828);
nand NAND3 (N8840, N8804, N2691, N1762);
not NOT1 (N8841, N8839);
nand NAND3 (N8842, N8841, N6888, N5173);
nand NAND3 (N8843, N8820, N7563, N4916);
nand NAND4 (N8844, N8827, N5570, N447, N3629);
and AND4 (N8845, N8843, N2981, N6029, N5701);
or OR4 (N8846, N8833, N1404, N2148, N6415);
nor NOR3 (N8847, N8845, N5179, N2409);
buf BUF1 (N8848, N8844);
buf BUF1 (N8849, N8825);
xor XOR2 (N8850, N8846, N3248);
nor NOR4 (N8851, N8842, N8844, N8398, N6246);
not NOT1 (N8852, N8840);
nand NAND4 (N8853, N8848, N8365, N8237, N4235);
buf BUF1 (N8854, N8838);
xor XOR2 (N8855, N8850, N8412);
buf BUF1 (N8856, N8852);
or OR3 (N8857, N8837, N6300, N3844);
buf BUF1 (N8858, N8855);
buf BUF1 (N8859, N8847);
not NOT1 (N8860, N8858);
nor NOR2 (N8861, N8853, N6368);
or OR2 (N8862, N8854, N8377);
buf BUF1 (N8863, N8836);
not NOT1 (N8864, N8859);
and AND2 (N8865, N8861, N5763);
and AND3 (N8866, N8849, N4958, N2742);
not NOT1 (N8867, N8865);
nand NAND2 (N8868, N8856, N1076);
or OR2 (N8869, N8867, N2322);
nor NOR2 (N8870, N8863, N2224);
nand NAND3 (N8871, N8862, N6608, N2161);
xor XOR2 (N8872, N8864, N3394);
not NOT1 (N8873, N8866);
nor NOR3 (N8874, N8869, N3738, N6597);
nor NOR3 (N8875, N8873, N888, N321);
not NOT1 (N8876, N8871);
nor NOR2 (N8877, N8851, N3743);
and AND2 (N8878, N8872, N1675);
or OR2 (N8879, N8835, N2872);
nor NOR2 (N8880, N8876, N7807);
buf BUF1 (N8881, N8870);
nand NAND4 (N8882, N8875, N2423, N3283, N428);
buf BUF1 (N8883, N8880);
xor XOR2 (N8884, N8874, N6599);
and AND4 (N8885, N8860, N3376, N8572, N3533);
nand NAND4 (N8886, N8883, N8049, N6623, N1528);
nor NOR3 (N8887, N8886, N5039, N4382);
not NOT1 (N8888, N8857);
or OR3 (N8889, N8868, N2073, N6234);
and AND4 (N8890, N8882, N242, N8641, N2316);
nor NOR4 (N8891, N8890, N6217, N2275, N3385);
or OR3 (N8892, N8887, N7556, N8239);
nand NAND4 (N8893, N8879, N398, N5684, N2230);
nor NOR2 (N8894, N8878, N5466);
xor XOR2 (N8895, N8892, N452);
nor NOR2 (N8896, N8881, N2202);
buf BUF1 (N8897, N8885);
or OR4 (N8898, N8884, N3715, N3436, N326);
buf BUF1 (N8899, N8888);
buf BUF1 (N8900, N8891);
and AND2 (N8901, N8899, N403);
xor XOR2 (N8902, N8889, N3388);
nand NAND3 (N8903, N8901, N2832, N8022);
nand NAND4 (N8904, N8895, N243, N192, N404);
not NOT1 (N8905, N8898);
nand NAND4 (N8906, N8903, N2515, N1264, N4156);
or OR4 (N8907, N8902, N7816, N1803, N4582);
xor XOR2 (N8908, N8905, N7031);
nand NAND2 (N8909, N8908, N2156);
or OR2 (N8910, N8897, N5219);
nor NOR3 (N8911, N8900, N5979, N8150);
nand NAND3 (N8912, N8877, N949, N7760);
nand NAND2 (N8913, N8911, N8327);
and AND4 (N8914, N8893, N4606, N6933, N2670);
nor NOR3 (N8915, N8894, N6894, N458);
xor XOR2 (N8916, N8910, N3694);
nand NAND4 (N8917, N8913, N7396, N859, N3125);
xor XOR2 (N8918, N8907, N8265);
nor NOR2 (N8919, N8896, N7447);
nand NAND3 (N8920, N8914, N2834, N5223);
nor NOR2 (N8921, N8904, N6359);
or OR2 (N8922, N8917, N7167);
nand NAND2 (N8923, N8919, N6702);
xor XOR2 (N8924, N8920, N7759);
nor NOR4 (N8925, N8912, N729, N5160, N3266);
or OR3 (N8926, N8909, N6359, N414);
or OR3 (N8927, N8922, N7021, N6036);
nor NOR3 (N8928, N8916, N2235, N2057);
nor NOR2 (N8929, N8926, N2912);
and AND3 (N8930, N8923, N4000, N2741);
and AND3 (N8931, N8918, N783, N8891);
nor NOR2 (N8932, N8921, N1934);
and AND2 (N8933, N8925, N3936);
nor NOR3 (N8934, N8932, N6332, N2704);
or OR4 (N8935, N8931, N8849, N5749, N6130);
nand NAND3 (N8936, N8934, N1970, N8276);
not NOT1 (N8937, N8906);
nand NAND2 (N8938, N8927, N3791);
nor NOR4 (N8939, N8937, N853, N8894, N4286);
not NOT1 (N8940, N8930);
nand NAND2 (N8941, N8935, N8637);
nor NOR3 (N8942, N8936, N3353, N1123);
or OR4 (N8943, N8928, N431, N1086, N2589);
nand NAND2 (N8944, N8929, N4933);
nor NOR3 (N8945, N8940, N401, N6391);
and AND3 (N8946, N8915, N794, N7242);
buf BUF1 (N8947, N8942);
or OR4 (N8948, N8938, N7884, N745, N6850);
xor XOR2 (N8949, N8947, N1727);
or OR4 (N8950, N8949, N8932, N1283, N1376);
xor XOR2 (N8951, N8941, N2663);
nand NAND4 (N8952, N8939, N246, N2623, N6118);
xor XOR2 (N8953, N8943, N8460);
nor NOR4 (N8954, N8948, N5416, N4075, N7684);
nor NOR3 (N8955, N8951, N7743, N3057);
nor NOR3 (N8956, N8955, N5619, N5858);
nor NOR3 (N8957, N8933, N4194, N8717);
nor NOR4 (N8958, N8957, N1116, N2267, N1637);
or OR3 (N8959, N8953, N4949, N216);
buf BUF1 (N8960, N8946);
nand NAND2 (N8961, N8924, N6313);
nand NAND2 (N8962, N8944, N3015);
xor XOR2 (N8963, N8956, N3711);
and AND2 (N8964, N8958, N3179);
not NOT1 (N8965, N8952);
nand NAND4 (N8966, N8962, N7572, N2797, N4708);
not NOT1 (N8967, N8959);
xor XOR2 (N8968, N8965, N7436);
nor NOR3 (N8969, N8964, N5819, N6459);
not NOT1 (N8970, N8950);
buf BUF1 (N8971, N8969);
nor NOR3 (N8972, N8967, N750, N4661);
or OR4 (N8973, N8963, N376, N1022, N513);
buf BUF1 (N8974, N8968);
xor XOR2 (N8975, N8972, N1305);
xor XOR2 (N8976, N8966, N979);
not NOT1 (N8977, N8971);
buf BUF1 (N8978, N8976);
xor XOR2 (N8979, N8954, N1180);
and AND3 (N8980, N8979, N1972, N7286);
xor XOR2 (N8981, N8980, N142);
xor XOR2 (N8982, N8970, N1462);
nand NAND4 (N8983, N8981, N1992, N495, N8744);
not NOT1 (N8984, N8973);
nor NOR4 (N8985, N8984, N3065, N921, N3050);
nand NAND3 (N8986, N8974, N1120, N916);
or OR2 (N8987, N8945, N1119);
and AND3 (N8988, N8987, N2009, N5702);
nand NAND3 (N8989, N8960, N981, N8293);
nor NOR3 (N8990, N8988, N2969, N6301);
and AND2 (N8991, N8977, N2359);
and AND3 (N8992, N8985, N1054, N368);
nand NAND2 (N8993, N8992, N8698);
nor NOR4 (N8994, N8986, N1060, N5530, N2676);
xor XOR2 (N8995, N8982, N3634);
not NOT1 (N8996, N8990);
nand NAND3 (N8997, N8983, N2389, N4517);
buf BUF1 (N8998, N8997);
nand NAND4 (N8999, N8993, N5981, N8541, N3372);
not NOT1 (N9000, N8994);
buf BUF1 (N9001, N8995);
not NOT1 (N9002, N8999);
xor XOR2 (N9003, N8998, N4081);
or OR3 (N9004, N8975, N1157, N385);
or OR4 (N9005, N8961, N2203, N6335, N1524);
and AND4 (N9006, N9004, N8909, N5088, N3040);
and AND3 (N9007, N9006, N7849, N3208);
xor XOR2 (N9008, N8989, N5206);
buf BUF1 (N9009, N9008);
or OR2 (N9010, N9007, N7047);
xor XOR2 (N9011, N9001, N8269);
buf BUF1 (N9012, N8996);
nand NAND2 (N9013, N9011, N6646);
nor NOR2 (N9014, N9009, N1339);
buf BUF1 (N9015, N9002);
nand NAND3 (N9016, N9013, N4196, N6972);
nor NOR3 (N9017, N9014, N5366, N6056);
and AND4 (N9018, N9016, N1965, N8746, N6101);
or OR3 (N9019, N9010, N4373, N1078);
buf BUF1 (N9020, N9012);
nand NAND2 (N9021, N9019, N1301);
and AND3 (N9022, N9021, N3232, N8154);
nor NOR2 (N9023, N9018, N1918);
nand NAND3 (N9024, N9003, N93, N8120);
xor XOR2 (N9025, N9017, N5766);
nand NAND3 (N9026, N8991, N4888, N235);
nor NOR4 (N9027, N9022, N2723, N437, N6191);
xor XOR2 (N9028, N9000, N4650);
buf BUF1 (N9029, N8978);
nand NAND4 (N9030, N9023, N5676, N6640, N5981);
nand NAND3 (N9031, N9030, N6016, N5098);
not NOT1 (N9032, N9027);
buf BUF1 (N9033, N9032);
nand NAND3 (N9034, N9026, N5497, N8175);
not NOT1 (N9035, N9033);
not NOT1 (N9036, N9024);
nor NOR3 (N9037, N9020, N3365, N4799);
nor NOR4 (N9038, N9028, N8341, N5662, N2342);
xor XOR2 (N9039, N9025, N4845);
nand NAND4 (N9040, N9029, N7747, N8399, N6886);
or OR3 (N9041, N9035, N8890, N5417);
nand NAND3 (N9042, N9040, N1281, N1661);
not NOT1 (N9043, N9038);
nand NAND4 (N9044, N9042, N4433, N6989, N3253);
xor XOR2 (N9045, N9037, N5970);
buf BUF1 (N9046, N9039);
xor XOR2 (N9047, N9036, N1449);
not NOT1 (N9048, N9046);
buf BUF1 (N9049, N9048);
nor NOR4 (N9050, N9034, N7955, N3157, N376);
nor NOR4 (N9051, N9031, N2771, N4852, N5877);
buf BUF1 (N9052, N9045);
buf BUF1 (N9053, N9043);
xor XOR2 (N9054, N9041, N4110);
and AND2 (N9055, N9047, N818);
nand NAND4 (N9056, N9050, N8153, N1387, N6147);
nand NAND3 (N9057, N9056, N4865, N4424);
buf BUF1 (N9058, N9051);
and AND3 (N9059, N9044, N8535, N8605);
nand NAND2 (N9060, N9015, N4721);
and AND4 (N9061, N9055, N5901, N7922, N7380);
and AND3 (N9062, N9057, N4585, N660);
not NOT1 (N9063, N9005);
nand NAND3 (N9064, N9058, N2404, N1186);
or OR3 (N9065, N9053, N6386, N7838);
or OR4 (N9066, N9061, N5922, N6404, N4687);
or OR2 (N9067, N9052, N6917);
xor XOR2 (N9068, N9060, N7598);
buf BUF1 (N9069, N9062);
and AND2 (N9070, N9064, N3634);
nor NOR2 (N9071, N9059, N7918);
xor XOR2 (N9072, N9070, N2657);
xor XOR2 (N9073, N9067, N8832);
xor XOR2 (N9074, N9072, N352);
and AND2 (N9075, N9049, N6130);
xor XOR2 (N9076, N9075, N4622);
not NOT1 (N9077, N9069);
or OR4 (N9078, N9065, N1851, N7291, N6176);
and AND4 (N9079, N9077, N8844, N7431, N2920);
or OR4 (N9080, N9073, N4140, N4443, N5739);
and AND2 (N9081, N9071, N8630);
nor NOR2 (N9082, N9081, N942);
not NOT1 (N9083, N9066);
xor XOR2 (N9084, N9079, N6937);
not NOT1 (N9085, N9082);
not NOT1 (N9086, N9078);
or OR2 (N9087, N9074, N4222);
buf BUF1 (N9088, N9080);
xor XOR2 (N9089, N9087, N2385);
nand NAND4 (N9090, N9076, N5423, N6657, N7009);
not NOT1 (N9091, N9086);
nor NOR4 (N9092, N9063, N2230, N401, N1438);
not NOT1 (N9093, N9083);
not NOT1 (N9094, N9085);
nand NAND3 (N9095, N9091, N4687, N6779);
nand NAND3 (N9096, N9068, N726, N6016);
or OR4 (N9097, N9095, N389, N4261, N3516);
and AND4 (N9098, N9097, N1987, N1264, N5276);
nor NOR2 (N9099, N9093, N8651);
nor NOR4 (N9100, N9094, N3636, N8055, N5183);
nand NAND2 (N9101, N9096, N8789);
buf BUF1 (N9102, N9101);
or OR3 (N9103, N9092, N1807, N4828);
nor NOR2 (N9104, N9099, N5860);
nor NOR2 (N9105, N9104, N7620);
nand NAND4 (N9106, N9088, N2055, N5997, N2707);
xor XOR2 (N9107, N9089, N2995);
or OR4 (N9108, N9100, N1863, N5358, N1970);
nor NOR3 (N9109, N9090, N4878, N2071);
and AND3 (N9110, N9109, N371, N2371);
xor XOR2 (N9111, N9108, N810);
nor NOR4 (N9112, N9084, N157, N4121, N3268);
or OR4 (N9113, N9098, N8745, N4766, N7349);
or OR3 (N9114, N9105, N1192, N3764);
buf BUF1 (N9115, N9114);
nor NOR3 (N9116, N9103, N3407, N5107);
not NOT1 (N9117, N9107);
nor NOR2 (N9118, N9115, N4816);
nand NAND2 (N9119, N9113, N7189);
not NOT1 (N9120, N9111);
nand NAND4 (N9121, N9110, N6059, N616, N8890);
nor NOR2 (N9122, N9119, N5151);
buf BUF1 (N9123, N9122);
or OR2 (N9124, N9054, N4506);
buf BUF1 (N9125, N9106);
and AND3 (N9126, N9123, N244, N298);
buf BUF1 (N9127, N9120);
nand NAND4 (N9128, N9102, N1606, N4305, N4464);
not NOT1 (N9129, N9112);
or OR4 (N9130, N9125, N1247, N5626, N2727);
not NOT1 (N9131, N9126);
or OR2 (N9132, N9129, N7170);
nor NOR3 (N9133, N9118, N328, N6563);
and AND3 (N9134, N9127, N588, N6340);
or OR2 (N9135, N9128, N269);
nor NOR3 (N9136, N9131, N2981, N3506);
nand NAND3 (N9137, N9132, N2914, N6605);
buf BUF1 (N9138, N9121);
and AND4 (N9139, N9130, N5436, N6222, N8749);
not NOT1 (N9140, N9135);
xor XOR2 (N9141, N9116, N5457);
and AND3 (N9142, N9139, N189, N7497);
nand NAND4 (N9143, N9138, N6191, N4203, N7658);
nor NOR4 (N9144, N9143, N8022, N1682, N3791);
and AND2 (N9145, N9136, N4447);
xor XOR2 (N9146, N9140, N7706);
or OR3 (N9147, N9134, N8618, N4002);
or OR2 (N9148, N9147, N1268);
buf BUF1 (N9149, N9124);
nand NAND2 (N9150, N9148, N6081);
nand NAND2 (N9151, N9142, N2172);
buf BUF1 (N9152, N9144);
buf BUF1 (N9153, N9137);
not NOT1 (N9154, N9117);
nor NOR2 (N9155, N9150, N6278);
or OR2 (N9156, N9155, N1757);
and AND2 (N9157, N9151, N1208);
nand NAND2 (N9158, N9153, N3429);
nand NAND3 (N9159, N9149, N8308, N371);
buf BUF1 (N9160, N9145);
not NOT1 (N9161, N9158);
nand NAND2 (N9162, N9161, N6647);
and AND4 (N9163, N9160, N3396, N8653, N74);
xor XOR2 (N9164, N9159, N2741);
or OR3 (N9165, N9154, N3158, N2861);
buf BUF1 (N9166, N9152);
nor NOR2 (N9167, N9166, N5473);
nor NOR4 (N9168, N9163, N7476, N8319, N6312);
buf BUF1 (N9169, N9168);
and AND4 (N9170, N9167, N3950, N7228, N3363);
nor NOR4 (N9171, N9169, N8641, N5962, N3867);
nand NAND4 (N9172, N9133, N4969, N1722, N4017);
buf BUF1 (N9173, N9157);
not NOT1 (N9174, N9165);
and AND4 (N9175, N9162, N3461, N1424, N664);
or OR4 (N9176, N9141, N6584, N3406, N8171);
and AND3 (N9177, N9175, N8285, N9064);
xor XOR2 (N9178, N9176, N7804);
nor NOR4 (N9179, N9177, N4994, N8988, N4018);
buf BUF1 (N9180, N9146);
buf BUF1 (N9181, N9174);
not NOT1 (N9182, N9170);
buf BUF1 (N9183, N9172);
buf BUF1 (N9184, N9182);
xor XOR2 (N9185, N9181, N3186);
xor XOR2 (N9186, N9180, N9143);
buf BUF1 (N9187, N9185);
and AND2 (N9188, N9173, N5506);
xor XOR2 (N9189, N9178, N3869);
or OR3 (N9190, N9183, N7228, N6460);
xor XOR2 (N9191, N9188, N2412);
nor NOR4 (N9192, N9191, N8433, N7721, N414);
or OR2 (N9193, N9192, N5660);
and AND4 (N9194, N9164, N8485, N4856, N7800);
buf BUF1 (N9195, N9189);
xor XOR2 (N9196, N9171, N8045);
nand NAND2 (N9197, N9184, N1878);
buf BUF1 (N9198, N9196);
nand NAND4 (N9199, N9186, N8340, N5797, N6521);
nand NAND2 (N9200, N9190, N1703);
xor XOR2 (N9201, N9187, N8703);
not NOT1 (N9202, N9197);
nand NAND2 (N9203, N9200, N1092);
not NOT1 (N9204, N9156);
or OR2 (N9205, N9204, N3387);
or OR2 (N9206, N9199, N4378);
not NOT1 (N9207, N9201);
or OR3 (N9208, N9195, N8696, N7641);
nor NOR2 (N9209, N9193, N3322);
nand NAND2 (N9210, N9194, N7525);
xor XOR2 (N9211, N9208, N7334);
not NOT1 (N9212, N9203);
or OR3 (N9213, N9206, N8432, N4353);
or OR3 (N9214, N9179, N4340, N4364);
not NOT1 (N9215, N9212);
xor XOR2 (N9216, N9210, N1517);
xor XOR2 (N9217, N9209, N5313);
buf BUF1 (N9218, N9207);
nor NOR3 (N9219, N9216, N5584, N6618);
not NOT1 (N9220, N9215);
or OR2 (N9221, N9198, N5071);
not NOT1 (N9222, N9217);
xor XOR2 (N9223, N9211, N5425);
and AND2 (N9224, N9213, N5378);
nand NAND3 (N9225, N9221, N2985, N1496);
buf BUF1 (N9226, N9202);
buf BUF1 (N9227, N9205);
nor NOR3 (N9228, N9225, N8332, N1117);
and AND3 (N9229, N9214, N7671, N2645);
xor XOR2 (N9230, N9220, N2066);
or OR4 (N9231, N9224, N4686, N5256, N918);
buf BUF1 (N9232, N9219);
buf BUF1 (N9233, N9230);
xor XOR2 (N9234, N9231, N1544);
not NOT1 (N9235, N9228);
nand NAND2 (N9236, N9223, N5989);
buf BUF1 (N9237, N9222);
nor NOR3 (N9238, N9232, N5844, N3405);
nor NOR3 (N9239, N9237, N2187, N7277);
or OR2 (N9240, N9218, N5596);
nor NOR4 (N9241, N9238, N2949, N481, N6928);
buf BUF1 (N9242, N9226);
nor NOR2 (N9243, N9236, N7255);
nand NAND4 (N9244, N9227, N6683, N6843, N2018);
or OR3 (N9245, N9235, N6603, N3938);
and AND3 (N9246, N9234, N2091, N1128);
or OR3 (N9247, N9246, N7821, N4928);
or OR3 (N9248, N9239, N268, N4490);
nor NOR3 (N9249, N9243, N493, N4609);
and AND4 (N9250, N9245, N7544, N4660, N5316);
xor XOR2 (N9251, N9248, N1723);
or OR2 (N9252, N9244, N3221);
nor NOR4 (N9253, N9249, N7030, N5380, N7586);
xor XOR2 (N9254, N9240, N5194);
nand NAND3 (N9255, N9251, N8061, N3240);
xor XOR2 (N9256, N9252, N1352);
nor NOR3 (N9257, N9242, N3044, N3827);
xor XOR2 (N9258, N9250, N885);
nand NAND4 (N9259, N9256, N6836, N2291, N8133);
xor XOR2 (N9260, N9247, N2676);
not NOT1 (N9261, N9233);
xor XOR2 (N9262, N9255, N8595);
buf BUF1 (N9263, N9260);
not NOT1 (N9264, N9257);
buf BUF1 (N9265, N9241);
buf BUF1 (N9266, N9262);
or OR4 (N9267, N9229, N6010, N7579, N5593);
and AND2 (N9268, N9261, N3463);
and AND4 (N9269, N9268, N1538, N784, N5671);
or OR3 (N9270, N9266, N5168, N2226);
or OR2 (N9271, N9265, N1324);
not NOT1 (N9272, N9267);
and AND2 (N9273, N9269, N8062);
and AND2 (N9274, N9258, N5646);
nand NAND2 (N9275, N9259, N8397);
xor XOR2 (N9276, N9264, N1892);
or OR4 (N9277, N9270, N7287, N6495, N5827);
or OR3 (N9278, N9271, N4356, N4823);
nor NOR4 (N9279, N9274, N4868, N2922, N2820);
xor XOR2 (N9280, N9254, N6315);
and AND3 (N9281, N9263, N3830, N2501);
buf BUF1 (N9282, N9280);
not NOT1 (N9283, N9275);
buf BUF1 (N9284, N9277);
nand NAND3 (N9285, N9281, N1324, N533);
not NOT1 (N9286, N9279);
nor NOR3 (N9287, N9278, N823, N3706);
nor NOR2 (N9288, N9272, N4804);
nand NAND2 (N9289, N9253, N1492);
not NOT1 (N9290, N9283);
nor NOR2 (N9291, N9287, N8786);
or OR3 (N9292, N9288, N8530, N2593);
or OR2 (N9293, N9285, N3342);
xor XOR2 (N9294, N9290, N5475);
xor XOR2 (N9295, N9282, N7056);
and AND3 (N9296, N9286, N182, N4494);
or OR2 (N9297, N9291, N5720);
or OR4 (N9298, N9294, N5440, N4577, N5620);
nor NOR3 (N9299, N9297, N1160, N5230);
or OR4 (N9300, N9298, N6952, N7968, N5371);
and AND2 (N9301, N9273, N6515);
and AND4 (N9302, N9301, N6653, N4446, N5936);
or OR4 (N9303, N9299, N3869, N6296, N5077);
not NOT1 (N9304, N9289);
nand NAND2 (N9305, N9295, N4737);
nand NAND3 (N9306, N9303, N947, N6972);
buf BUF1 (N9307, N9305);
or OR4 (N9308, N9302, N4731, N5259, N694);
buf BUF1 (N9309, N9307);
xor XOR2 (N9310, N9292, N5560);
buf BUF1 (N9311, N9276);
nand NAND3 (N9312, N9296, N6295, N4799);
not NOT1 (N9313, N9304);
not NOT1 (N9314, N9311);
nor NOR3 (N9315, N9300, N8126, N5032);
nor NOR3 (N9316, N9306, N2389, N5356);
xor XOR2 (N9317, N9284, N5345);
buf BUF1 (N9318, N9293);
nor NOR3 (N9319, N9308, N5319, N6141);
not NOT1 (N9320, N9317);
xor XOR2 (N9321, N9315, N2538);
and AND2 (N9322, N9313, N8798);
xor XOR2 (N9323, N9322, N6296);
or OR4 (N9324, N9323, N7775, N8343, N5291);
or OR4 (N9325, N9312, N9011, N6189, N9151);
nand NAND2 (N9326, N9320, N5860);
and AND2 (N9327, N9319, N1888);
nand NAND3 (N9328, N9309, N9308, N96);
not NOT1 (N9329, N9318);
buf BUF1 (N9330, N9325);
or OR2 (N9331, N9314, N7974);
nand NAND2 (N9332, N9331, N6769);
buf BUF1 (N9333, N9328);
nor NOR2 (N9334, N9321, N4654);
not NOT1 (N9335, N9310);
xor XOR2 (N9336, N9335, N7636);
or OR3 (N9337, N9327, N7228, N5356);
xor XOR2 (N9338, N9333, N4990);
and AND4 (N9339, N9338, N2020, N8005, N5820);
and AND4 (N9340, N9329, N2894, N416, N8376);
buf BUF1 (N9341, N9316);
buf BUF1 (N9342, N9341);
not NOT1 (N9343, N9326);
xor XOR2 (N9344, N9343, N8928);
nor NOR3 (N9345, N9336, N7691, N2391);
buf BUF1 (N9346, N9324);
nand NAND2 (N9347, N9345, N7706);
nor NOR2 (N9348, N9346, N8179);
buf BUF1 (N9349, N9342);
nand NAND2 (N9350, N9340, N8051);
nand NAND3 (N9351, N9330, N549, N6696);
buf BUF1 (N9352, N9334);
buf BUF1 (N9353, N9347);
or OR3 (N9354, N9332, N6633, N4290);
nand NAND4 (N9355, N9348, N5328, N4340, N9274);
or OR2 (N9356, N9339, N7907);
or OR2 (N9357, N9354, N205);
buf BUF1 (N9358, N9350);
xor XOR2 (N9359, N9349, N7377);
buf BUF1 (N9360, N9353);
nor NOR4 (N9361, N9357, N2238, N2510, N2488);
and AND3 (N9362, N9356, N3246, N2683);
nor NOR3 (N9363, N9360, N6796, N912);
not NOT1 (N9364, N9351);
xor XOR2 (N9365, N9359, N3144);
xor XOR2 (N9366, N9362, N1226);
nand NAND3 (N9367, N9358, N8501, N4437);
buf BUF1 (N9368, N9366);
and AND2 (N9369, N9352, N6093);
xor XOR2 (N9370, N9364, N2021);
xor XOR2 (N9371, N9370, N864);
xor XOR2 (N9372, N9344, N4761);
nand NAND3 (N9373, N9365, N8011, N1193);
not NOT1 (N9374, N9361);
or OR3 (N9375, N9369, N2681, N6748);
or OR2 (N9376, N9373, N2298);
nand NAND3 (N9377, N9355, N654, N1055);
or OR4 (N9378, N9367, N1243, N8989, N2828);
nor NOR3 (N9379, N9371, N8144, N5878);
nand NAND2 (N9380, N9377, N790);
buf BUF1 (N9381, N9337);
nor NOR4 (N9382, N9372, N8009, N4013, N8904);
nor NOR4 (N9383, N9374, N170, N8970, N7469);
xor XOR2 (N9384, N9380, N2108);
not NOT1 (N9385, N9368);
and AND3 (N9386, N9379, N4796, N6325);
nor NOR3 (N9387, N9385, N9155, N6666);
or OR4 (N9388, N9387, N744, N5032, N5714);
not NOT1 (N9389, N9376);
buf BUF1 (N9390, N9383);
xor XOR2 (N9391, N9388, N1296);
or OR4 (N9392, N9382, N2167, N4802, N2900);
buf BUF1 (N9393, N9363);
nor NOR2 (N9394, N9378, N3884);
nand NAND4 (N9395, N9390, N4028, N2467, N2956);
buf BUF1 (N9396, N9381);
buf BUF1 (N9397, N9391);
not NOT1 (N9398, N9393);
nor NOR2 (N9399, N9397, N3095);
buf BUF1 (N9400, N9384);
buf BUF1 (N9401, N9395);
not NOT1 (N9402, N9392);
xor XOR2 (N9403, N9394, N4673);
nor NOR2 (N9404, N9401, N7154);
xor XOR2 (N9405, N9403, N6224);
or OR3 (N9406, N9400, N2778, N5064);
not NOT1 (N9407, N9396);
not NOT1 (N9408, N9386);
xor XOR2 (N9409, N9405, N7559);
nor NOR4 (N9410, N9402, N7729, N2787, N8142);
nor NOR3 (N9411, N9406, N5608, N1059);
and AND3 (N9412, N9399, N8619, N9343);
and AND4 (N9413, N9408, N6685, N7041, N1655);
or OR2 (N9414, N9409, N7225);
xor XOR2 (N9415, N9407, N4858);
buf BUF1 (N9416, N9411);
xor XOR2 (N9417, N9414, N6612);
nand NAND2 (N9418, N9413, N6761);
not NOT1 (N9419, N9415);
not NOT1 (N9420, N9375);
not NOT1 (N9421, N9404);
buf BUF1 (N9422, N9419);
buf BUF1 (N9423, N9417);
and AND3 (N9424, N9421, N2839, N5878);
or OR2 (N9425, N9424, N1136);
buf BUF1 (N9426, N9389);
and AND3 (N9427, N9425, N4908, N2690);
buf BUF1 (N9428, N9423);
and AND2 (N9429, N9422, N3695);
nand NAND3 (N9430, N9416, N8080, N8708);
nor NOR2 (N9431, N9427, N6837);
buf BUF1 (N9432, N9420);
nand NAND4 (N9433, N9418, N2128, N7434, N1049);
and AND3 (N9434, N9412, N481, N3602);
xor XOR2 (N9435, N9429, N6382);
xor XOR2 (N9436, N9410, N4327);
nand NAND4 (N9437, N9432, N1201, N2177, N1141);
or OR4 (N9438, N9433, N169, N1021, N2667);
nand NAND4 (N9439, N9437, N9103, N3337, N6934);
nor NOR4 (N9440, N9439, N4621, N3045, N7165);
not NOT1 (N9441, N9428);
buf BUF1 (N9442, N9430);
nand NAND4 (N9443, N9442, N7872, N2483, N531);
nand NAND3 (N9444, N9426, N3652, N7988);
buf BUF1 (N9445, N9398);
nor NOR2 (N9446, N9434, N5718);
nor NOR2 (N9447, N9443, N507);
nand NAND4 (N9448, N9444, N7729, N4656, N4105);
buf BUF1 (N9449, N9447);
nor NOR2 (N9450, N9440, N6692);
and AND3 (N9451, N9449, N655, N66);
buf BUF1 (N9452, N9448);
buf BUF1 (N9453, N9431);
nor NOR2 (N9454, N9445, N8807);
nor NOR4 (N9455, N9451, N2237, N8709, N8642);
nand NAND3 (N9456, N9454, N5171, N7293);
nor NOR3 (N9457, N9455, N960, N5978);
nor NOR3 (N9458, N9441, N82, N2570);
and AND3 (N9459, N9453, N6108, N6187);
buf BUF1 (N9460, N9436);
or OR3 (N9461, N9446, N5073, N1073);
and AND4 (N9462, N9459, N3775, N4702, N5400);
nor NOR4 (N9463, N9435, N6217, N136, N8938);
or OR3 (N9464, N9462, N8433, N6028);
not NOT1 (N9465, N9438);
or OR4 (N9466, N9458, N7555, N2693, N1816);
buf BUF1 (N9467, N9464);
and AND3 (N9468, N9452, N4303, N7190);
or OR4 (N9469, N9456, N2894, N5722, N1647);
not NOT1 (N9470, N9468);
nand NAND3 (N9471, N9469, N2515, N5888);
and AND3 (N9472, N9457, N3023, N4191);
nor NOR4 (N9473, N9450, N7794, N8283, N4822);
or OR2 (N9474, N9460, N2899);
nand NAND4 (N9475, N9470, N6544, N4814, N1623);
not NOT1 (N9476, N9472);
not NOT1 (N9477, N9465);
not NOT1 (N9478, N9467);
and AND3 (N9479, N9463, N241, N6307);
not NOT1 (N9480, N9478);
not NOT1 (N9481, N9471);
nor NOR4 (N9482, N9476, N4358, N6854, N9365);
or OR4 (N9483, N9461, N8080, N8234, N3214);
or OR3 (N9484, N9474, N3337, N1473);
not NOT1 (N9485, N9473);
nor NOR2 (N9486, N9479, N4177);
nand NAND3 (N9487, N9483, N6873, N4571);
nand NAND2 (N9488, N9485, N3426);
nor NOR2 (N9489, N9477, N9022);
nor NOR2 (N9490, N9484, N5136);
xor XOR2 (N9491, N9466, N6147);
and AND3 (N9492, N9488, N5140, N9341);
nand NAND4 (N9493, N9492, N7769, N7620, N6703);
not NOT1 (N9494, N9490);
and AND2 (N9495, N9475, N2092);
not NOT1 (N9496, N9480);
buf BUF1 (N9497, N9489);
nand NAND4 (N9498, N9496, N7248, N5446, N5615);
not NOT1 (N9499, N9481);
nand NAND3 (N9500, N9498, N2992, N6788);
or OR2 (N9501, N9494, N4915);
buf BUF1 (N9502, N9486);
nand NAND2 (N9503, N9501, N7714);
nand NAND2 (N9504, N9500, N4507);
not NOT1 (N9505, N9482);
nand NAND3 (N9506, N9487, N2889, N5189);
or OR3 (N9507, N9491, N7677, N2010);
buf BUF1 (N9508, N9504);
nor NOR3 (N9509, N9505, N833, N8409);
and AND3 (N9510, N9503, N3410, N7777);
not NOT1 (N9511, N9495);
xor XOR2 (N9512, N9493, N9441);
nor NOR2 (N9513, N9502, N9443);
or OR3 (N9514, N9509, N8568, N8166);
or OR3 (N9515, N9511, N339, N9372);
xor XOR2 (N9516, N9497, N1711);
buf BUF1 (N9517, N9512);
and AND4 (N9518, N9513, N2403, N1050, N6821);
nand NAND4 (N9519, N9518, N5990, N5646, N7323);
nor NOR2 (N9520, N9510, N5345);
nor NOR2 (N9521, N9499, N5496);
buf BUF1 (N9522, N9507);
or OR2 (N9523, N9506, N402);
or OR2 (N9524, N9517, N9113);
not NOT1 (N9525, N9514);
nor NOR3 (N9526, N9520, N2991, N3309);
not NOT1 (N9527, N9524);
or OR2 (N9528, N9525, N2821);
not NOT1 (N9529, N9523);
nand NAND4 (N9530, N9526, N1195, N6019, N7075);
xor XOR2 (N9531, N9516, N3161);
xor XOR2 (N9532, N9527, N394);
xor XOR2 (N9533, N9508, N8133);
and AND4 (N9534, N9532, N2048, N141, N8227);
buf BUF1 (N9535, N9515);
nand NAND2 (N9536, N9522, N7371);
not NOT1 (N9537, N9536);
not NOT1 (N9538, N9534);
or OR3 (N9539, N9519, N5141, N2587);
or OR2 (N9540, N9521, N27);
nand NAND4 (N9541, N9528, N6046, N8758, N912);
xor XOR2 (N9542, N9541, N3181);
and AND3 (N9543, N9529, N5150, N3389);
nor NOR3 (N9544, N9543, N1671, N1855);
xor XOR2 (N9545, N9539, N904);
nor NOR3 (N9546, N9530, N8980, N3601);
not NOT1 (N9547, N9538);
buf BUF1 (N9548, N9531);
or OR4 (N9549, N9540, N7463, N7364, N5313);
nor NOR4 (N9550, N9549, N1397, N3891, N821);
buf BUF1 (N9551, N9533);
not NOT1 (N9552, N9546);
nor NOR3 (N9553, N9550, N7507, N9028);
xor XOR2 (N9554, N9545, N8957);
nand NAND2 (N9555, N9551, N793);
or OR2 (N9556, N9554, N8459);
nand NAND4 (N9557, N9553, N6838, N5904, N6998);
buf BUF1 (N9558, N9544);
xor XOR2 (N9559, N9535, N1740);
xor XOR2 (N9560, N9552, N1464);
and AND3 (N9561, N9542, N4281, N4917);
nand NAND2 (N9562, N9556, N4628);
nand NAND4 (N9563, N9555, N4282, N6222, N4680);
nand NAND4 (N9564, N9561, N179, N243, N8888);
xor XOR2 (N9565, N9560, N2821);
xor XOR2 (N9566, N9557, N6952);
or OR2 (N9567, N9548, N7248);
not NOT1 (N9568, N9562);
xor XOR2 (N9569, N9564, N3437);
and AND3 (N9570, N9559, N7562, N3710);
xor XOR2 (N9571, N9566, N7125);
and AND2 (N9572, N9567, N5280);
not NOT1 (N9573, N9565);
xor XOR2 (N9574, N9572, N3353);
xor XOR2 (N9575, N9573, N7726);
not NOT1 (N9576, N9574);
and AND2 (N9577, N9537, N6877);
or OR2 (N9578, N9558, N7461);
buf BUF1 (N9579, N9577);
nor NOR2 (N9580, N9578, N1248);
or OR3 (N9581, N9568, N694, N8050);
nor NOR3 (N9582, N9579, N3475, N6095);
nand NAND2 (N9583, N9571, N928);
and AND2 (N9584, N9580, N1075);
xor XOR2 (N9585, N9547, N7810);
and AND2 (N9586, N9581, N2058);
and AND4 (N9587, N9583, N2813, N9111, N9378);
nand NAND3 (N9588, N9563, N3087, N1877);
buf BUF1 (N9589, N9569);
nand NAND4 (N9590, N9586, N3461, N1796, N6852);
not NOT1 (N9591, N9588);
xor XOR2 (N9592, N9584, N2669);
nand NAND2 (N9593, N9585, N5657);
buf BUF1 (N9594, N9575);
or OR2 (N9595, N9589, N5348);
and AND3 (N9596, N9576, N6523, N5528);
xor XOR2 (N9597, N9595, N7155);
not NOT1 (N9598, N9597);
not NOT1 (N9599, N9591);
not NOT1 (N9600, N9593);
not NOT1 (N9601, N9598);
or OR2 (N9602, N9601, N1782);
and AND3 (N9603, N9599, N1840, N3273);
buf BUF1 (N9604, N9587);
and AND2 (N9605, N9590, N2694);
not NOT1 (N9606, N9592);
xor XOR2 (N9607, N9602, N7807);
and AND4 (N9608, N9600, N8931, N3418, N3767);
buf BUF1 (N9609, N9570);
buf BUF1 (N9610, N9609);
nor NOR2 (N9611, N9605, N4590);
or OR4 (N9612, N9582, N6073, N4350, N7869);
or OR2 (N9613, N9603, N9332);
or OR3 (N9614, N9613, N8459, N2408);
not NOT1 (N9615, N9604);
or OR2 (N9616, N9614, N3859);
nand NAND3 (N9617, N9615, N7888, N8570);
or OR3 (N9618, N9610, N5441, N3436);
buf BUF1 (N9619, N9617);
nor NOR2 (N9620, N9606, N7048);
not NOT1 (N9621, N9608);
and AND2 (N9622, N9607, N8154);
not NOT1 (N9623, N9620);
xor XOR2 (N9624, N9594, N3898);
not NOT1 (N9625, N9622);
buf BUF1 (N9626, N9618);
nand NAND2 (N9627, N9616, N6853);
xor XOR2 (N9628, N9621, N9143);
and AND2 (N9629, N9612, N5695);
or OR4 (N9630, N9596, N6941, N5624, N5185);
xor XOR2 (N9631, N9630, N8652);
and AND3 (N9632, N9625, N7573, N3610);
and AND3 (N9633, N9624, N4399, N6081);
and AND2 (N9634, N9623, N7936);
xor XOR2 (N9635, N9627, N1584);
xor XOR2 (N9636, N9631, N1635);
or OR3 (N9637, N9629, N5478, N3558);
and AND2 (N9638, N9632, N8093);
nand NAND4 (N9639, N9636, N1715, N2060, N3323);
or OR4 (N9640, N9633, N2419, N9150, N5461);
or OR4 (N9641, N9637, N4625, N2853, N6515);
not NOT1 (N9642, N9634);
not NOT1 (N9643, N9640);
or OR4 (N9644, N9642, N177, N378, N6405);
nor NOR3 (N9645, N9644, N6491, N1905);
xor XOR2 (N9646, N9645, N2877);
not NOT1 (N9647, N9626);
or OR3 (N9648, N9628, N4210, N2025);
not NOT1 (N9649, N9646);
xor XOR2 (N9650, N9648, N3421);
or OR2 (N9651, N9641, N4887);
and AND3 (N9652, N9643, N3180, N6080);
and AND3 (N9653, N9638, N6668, N81);
not NOT1 (N9654, N9647);
xor XOR2 (N9655, N9635, N1127);
nor NOR2 (N9656, N9651, N9501);
or OR4 (N9657, N9655, N2705, N8413, N1294);
nor NOR2 (N9658, N9639, N8788);
not NOT1 (N9659, N9652);
nand NAND2 (N9660, N9653, N7578);
buf BUF1 (N9661, N9619);
nand NAND4 (N9662, N9657, N3248, N340, N3340);
nand NAND2 (N9663, N9660, N4816);
xor XOR2 (N9664, N9649, N2957);
buf BUF1 (N9665, N9663);
or OR4 (N9666, N9661, N3587, N5447, N5567);
or OR4 (N9667, N9654, N8278, N7360, N7781);
buf BUF1 (N9668, N9666);
nor NOR3 (N9669, N9650, N4524, N2571);
or OR2 (N9670, N9667, N7528);
and AND2 (N9671, N9670, N3472);
and AND4 (N9672, N9664, N7020, N7675, N8996);
nor NOR2 (N9673, N9662, N5302);
buf BUF1 (N9674, N9656);
or OR2 (N9675, N9659, N2859);
not NOT1 (N9676, N9669);
xor XOR2 (N9677, N9676, N1300);
nor NOR2 (N9678, N9668, N824);
xor XOR2 (N9679, N9672, N9303);
and AND2 (N9680, N9679, N5960);
nor NOR4 (N9681, N9671, N5192, N2671, N3129);
xor XOR2 (N9682, N9677, N2457);
buf BUF1 (N9683, N9675);
xor XOR2 (N9684, N9665, N6320);
and AND3 (N9685, N9680, N137, N5782);
not NOT1 (N9686, N9685);
buf BUF1 (N9687, N9658);
buf BUF1 (N9688, N9674);
xor XOR2 (N9689, N9688, N3569);
nand NAND4 (N9690, N9687, N1678, N642, N3985);
or OR2 (N9691, N9689, N7742);
nor NOR3 (N9692, N9681, N4334, N11);
nor NOR2 (N9693, N9690, N3947);
nand NAND4 (N9694, N9678, N3879, N8811, N639);
nand NAND3 (N9695, N9692, N2573, N1534);
and AND4 (N9696, N9693, N7706, N6156, N8417);
not NOT1 (N9697, N9683);
and AND3 (N9698, N9691, N1862, N5095);
xor XOR2 (N9699, N9694, N3573);
xor XOR2 (N9700, N9698, N9515);
buf BUF1 (N9701, N9695);
nand NAND4 (N9702, N9696, N7494, N8378, N9435);
nand NAND3 (N9703, N9611, N1875, N507);
nand NAND3 (N9704, N9697, N1468, N595);
xor XOR2 (N9705, N9703, N3915);
nand NAND3 (N9706, N9702, N1978, N3899);
and AND2 (N9707, N9706, N6859);
xor XOR2 (N9708, N9701, N183);
buf BUF1 (N9709, N9682);
nand NAND3 (N9710, N9705, N7897, N682);
nor NOR3 (N9711, N9707, N2870, N2039);
or OR3 (N9712, N9673, N9689, N9244);
not NOT1 (N9713, N9710);
not NOT1 (N9714, N9712);
not NOT1 (N9715, N9699);
xor XOR2 (N9716, N9704, N9154);
buf BUF1 (N9717, N9686);
not NOT1 (N9718, N9714);
or OR4 (N9719, N9684, N7227, N8544, N5522);
not NOT1 (N9720, N9708);
nor NOR2 (N9721, N9713, N6730);
not NOT1 (N9722, N9711);
xor XOR2 (N9723, N9716, N7252);
xor XOR2 (N9724, N9718, N2017);
nor NOR4 (N9725, N9709, N9720, N5843, N1706);
and AND2 (N9726, N5323, N8803);
and AND3 (N9727, N9722, N8192, N7302);
xor XOR2 (N9728, N9726, N584);
nor NOR4 (N9729, N9721, N7033, N8024, N5460);
buf BUF1 (N9730, N9723);
buf BUF1 (N9731, N9700);
buf BUF1 (N9732, N9725);
buf BUF1 (N9733, N9732);
not NOT1 (N9734, N9733);
nand NAND4 (N9735, N9724, N7002, N7656, N6181);
nor NOR2 (N9736, N9734, N6969);
xor XOR2 (N9737, N9717, N3643);
nor NOR4 (N9738, N9735, N2004, N1185, N4312);
or OR3 (N9739, N9715, N8418, N2896);
xor XOR2 (N9740, N9728, N7964);
buf BUF1 (N9741, N9737);
nand NAND3 (N9742, N9729, N4014, N7833);
nor NOR2 (N9743, N9719, N2867);
nor NOR2 (N9744, N9739, N9371);
or OR4 (N9745, N9741, N1923, N9665, N3057);
or OR2 (N9746, N9727, N3531);
and AND4 (N9747, N9730, N5578, N2421, N8668);
xor XOR2 (N9748, N9731, N9301);
nor NOR3 (N9749, N9736, N7556, N1187);
nor NOR3 (N9750, N9744, N5049, N1172);
nor NOR3 (N9751, N9740, N6281, N1290);
xor XOR2 (N9752, N9746, N8866);
xor XOR2 (N9753, N9747, N5587);
or OR4 (N9754, N9752, N3753, N8401, N9309);
nand NAND3 (N9755, N9745, N2521, N8127);
and AND3 (N9756, N9738, N8884, N4376);
and AND4 (N9757, N9742, N6676, N8517, N6040);
nor NOR4 (N9758, N9748, N79, N8241, N8073);
nor NOR3 (N9759, N9757, N8115, N7579);
xor XOR2 (N9760, N9758, N7453);
buf BUF1 (N9761, N9743);
nand NAND3 (N9762, N9751, N2435, N1809);
not NOT1 (N9763, N9750);
xor XOR2 (N9764, N9749, N692);
buf BUF1 (N9765, N9754);
xor XOR2 (N9766, N9761, N9156);
nor NOR4 (N9767, N9766, N4942, N1354, N1342);
xor XOR2 (N9768, N9755, N5966);
and AND4 (N9769, N9767, N5360, N2939, N9170);
nand NAND2 (N9770, N9769, N3377);
nor NOR3 (N9771, N9759, N8768, N1896);
xor XOR2 (N9772, N9770, N9621);
not NOT1 (N9773, N9771);
or OR3 (N9774, N9772, N4440, N2159);
not NOT1 (N9775, N9763);
and AND3 (N9776, N9764, N6093, N9607);
and AND4 (N9777, N9774, N2, N5504, N2203);
and AND3 (N9778, N9777, N7896, N6860);
buf BUF1 (N9779, N9765);
xor XOR2 (N9780, N9775, N400);
or OR2 (N9781, N9756, N6303);
nand NAND2 (N9782, N9776, N9763);
or OR3 (N9783, N9773, N3754, N543);
not NOT1 (N9784, N9768);
and AND2 (N9785, N9762, N8845);
not NOT1 (N9786, N9779);
and AND2 (N9787, N9778, N8335);
not NOT1 (N9788, N9780);
buf BUF1 (N9789, N9785);
nor NOR3 (N9790, N9789, N7889, N9738);
nor NOR4 (N9791, N9760, N6622, N558, N6958);
and AND4 (N9792, N9788, N5226, N3678, N2033);
nand NAND2 (N9793, N9786, N5907);
nor NOR3 (N9794, N9793, N1581, N5444);
not NOT1 (N9795, N9794);
nor NOR3 (N9796, N9781, N8544, N3815);
nor NOR4 (N9797, N9790, N6692, N4434, N8538);
buf BUF1 (N9798, N9796);
buf BUF1 (N9799, N9798);
and AND3 (N9800, N9791, N9757, N7604);
nor NOR4 (N9801, N9792, N9393, N7419, N4080);
nand NAND2 (N9802, N9797, N2846);
buf BUF1 (N9803, N9787);
or OR4 (N9804, N9802, N513, N3609, N5129);
xor XOR2 (N9805, N9753, N1453);
nand NAND3 (N9806, N9803, N3520, N5820);
xor XOR2 (N9807, N9805, N5608);
or OR2 (N9808, N9806, N3247);
not NOT1 (N9809, N9808);
nand NAND4 (N9810, N9783, N7739, N8154, N5571);
xor XOR2 (N9811, N9784, N5345);
or OR4 (N9812, N9800, N4899, N1937, N8989);
nor NOR4 (N9813, N9809, N7193, N597, N4256);
nand NAND3 (N9814, N9795, N505, N4248);
or OR2 (N9815, N9782, N997);
or OR3 (N9816, N9807, N610, N8437);
xor XOR2 (N9817, N9804, N6184);
or OR2 (N9818, N9814, N2921);
xor XOR2 (N9819, N9815, N2790);
nor NOR4 (N9820, N9810, N9392, N4620, N3219);
nor NOR2 (N9821, N9819, N7924);
nor NOR4 (N9822, N9817, N4981, N9281, N2704);
buf BUF1 (N9823, N9811);
nor NOR4 (N9824, N9812, N7300, N4410, N3555);
nand NAND4 (N9825, N9799, N2285, N5357, N9090);
not NOT1 (N9826, N9822);
nor NOR3 (N9827, N9820, N5512, N2475);
buf BUF1 (N9828, N9821);
xor XOR2 (N9829, N9801, N5363);
not NOT1 (N9830, N9828);
xor XOR2 (N9831, N9824, N3921);
nor NOR3 (N9832, N9829, N8803, N2733);
or OR4 (N9833, N9825, N2666, N9220, N7403);
and AND2 (N9834, N9831, N1507);
and AND2 (N9835, N9833, N1378);
buf BUF1 (N9836, N9830);
and AND4 (N9837, N9827, N7608, N8482, N9697);
xor XOR2 (N9838, N9834, N4170);
xor XOR2 (N9839, N9816, N2124);
not NOT1 (N9840, N9838);
buf BUF1 (N9841, N9837);
not NOT1 (N9842, N9826);
nor NOR2 (N9843, N9839, N403);
and AND2 (N9844, N9832, N1454);
and AND4 (N9845, N9844, N3647, N8172, N5095);
nand NAND2 (N9846, N9813, N7492);
xor XOR2 (N9847, N9841, N7083);
or OR3 (N9848, N9843, N628, N1993);
nor NOR3 (N9849, N9840, N3301, N6711);
nand NAND2 (N9850, N9835, N848);
nand NAND2 (N9851, N9818, N4661);
buf BUF1 (N9852, N9823);
buf BUF1 (N9853, N9850);
nor NOR4 (N9854, N9847, N6675, N2387, N5704);
nor NOR2 (N9855, N9851, N7687);
or OR3 (N9856, N9854, N9764, N8110);
or OR2 (N9857, N9845, N8016);
buf BUF1 (N9858, N9855);
xor XOR2 (N9859, N9856, N3773);
or OR2 (N9860, N9857, N8774);
nor NOR3 (N9861, N9853, N3091, N3917);
or OR2 (N9862, N9842, N486);
xor XOR2 (N9863, N9861, N997);
buf BUF1 (N9864, N9846);
or OR4 (N9865, N9860, N3064, N5040, N4603);
not NOT1 (N9866, N9864);
nand NAND2 (N9867, N9863, N4612);
buf BUF1 (N9868, N9858);
and AND2 (N9869, N9852, N6221);
buf BUF1 (N9870, N9859);
and AND3 (N9871, N9836, N7132, N8421);
or OR4 (N9872, N9870, N1244, N4253, N3702);
not NOT1 (N9873, N9868);
nor NOR2 (N9874, N9869, N69);
not NOT1 (N9875, N9862);
buf BUF1 (N9876, N9865);
xor XOR2 (N9877, N9876, N6884);
nor NOR4 (N9878, N9873, N3279, N5723, N1237);
not NOT1 (N9879, N9866);
xor XOR2 (N9880, N9879, N1405);
and AND3 (N9881, N9872, N2669, N2507);
buf BUF1 (N9882, N9881);
xor XOR2 (N9883, N9882, N7893);
nand NAND2 (N9884, N9877, N7149);
buf BUF1 (N9885, N9871);
nor NOR3 (N9886, N9880, N2172, N7754);
and AND3 (N9887, N9867, N7734, N1679);
nor NOR4 (N9888, N9885, N5637, N1079, N4789);
nor NOR4 (N9889, N9883, N6500, N3741, N8085);
and AND2 (N9890, N9886, N9084);
nand NAND4 (N9891, N9874, N4324, N5353, N3732);
not NOT1 (N9892, N9848);
not NOT1 (N9893, N9887);
nand NAND2 (N9894, N9884, N6840);
not NOT1 (N9895, N9890);
and AND4 (N9896, N9878, N8157, N4498, N2140);
not NOT1 (N9897, N9896);
or OR2 (N9898, N9849, N4363);
nor NOR2 (N9899, N9893, N2889);
or OR2 (N9900, N9897, N4637);
buf BUF1 (N9901, N9891);
nand NAND4 (N9902, N9889, N5774, N8777, N6584);
or OR2 (N9903, N9892, N8388);
and AND3 (N9904, N9902, N4305, N1337);
nand NAND2 (N9905, N9894, N7129);
not NOT1 (N9906, N9903);
nor NOR2 (N9907, N9901, N1509);
nor NOR2 (N9908, N9905, N847);
nor NOR3 (N9909, N9899, N255, N4388);
nor NOR4 (N9910, N9904, N3340, N7334, N6352);
not NOT1 (N9911, N9909);
buf BUF1 (N9912, N9908);
xor XOR2 (N9913, N9900, N6421);
xor XOR2 (N9914, N9898, N2205);
nor NOR2 (N9915, N9912, N5973);
or OR4 (N9916, N9888, N9633, N3547, N7830);
or OR4 (N9917, N9875, N358, N7428, N2758);
nand NAND4 (N9918, N9911, N5919, N6763, N2440);
or OR2 (N9919, N9913, N360);
not NOT1 (N9920, N9916);
not NOT1 (N9921, N9895);
and AND2 (N9922, N9906, N3476);
or OR4 (N9923, N9920, N9838, N5822, N2403);
not NOT1 (N9924, N9910);
not NOT1 (N9925, N9914);
nand NAND4 (N9926, N9922, N3068, N3498, N756);
nor NOR2 (N9927, N9923, N8633);
xor XOR2 (N9928, N9907, N6130);
buf BUF1 (N9929, N9928);
and AND3 (N9930, N9927, N6390, N9687);
buf BUF1 (N9931, N9926);
nor NOR4 (N9932, N9918, N65, N7813, N4449);
nor NOR3 (N9933, N9930, N9649, N3540);
or OR3 (N9934, N9931, N4237, N982);
nor NOR4 (N9935, N9932, N522, N1580, N1899);
nor NOR2 (N9936, N9933, N1396);
nand NAND3 (N9937, N9936, N3755, N7917);
and AND4 (N9938, N9937, N4692, N3598, N2518);
or OR2 (N9939, N9929, N5646);
xor XOR2 (N9940, N9915, N5720);
nand NAND4 (N9941, N9917, N7635, N9882, N1845);
nand NAND4 (N9942, N9935, N1868, N6756, N4862);
xor XOR2 (N9943, N9938, N3977);
and AND4 (N9944, N9940, N5465, N2056, N2419);
buf BUF1 (N9945, N9934);
nand NAND4 (N9946, N9919, N9879, N3332, N8087);
or OR4 (N9947, N9939, N1866, N2287, N5581);
or OR2 (N9948, N9942, N5883);
not NOT1 (N9949, N9925);
and AND4 (N9950, N9941, N2425, N7231, N7645);
buf BUF1 (N9951, N9924);
not NOT1 (N9952, N9946);
and AND4 (N9953, N9943, N2279, N1035, N7854);
xor XOR2 (N9954, N9948, N5906);
or OR4 (N9955, N9953, N5666, N5628, N4435);
nor NOR4 (N9956, N9952, N4379, N2529, N1814);
not NOT1 (N9957, N9956);
not NOT1 (N9958, N9947);
or OR4 (N9959, N9957, N5483, N4689, N541);
nand NAND4 (N9960, N9949, N5005, N801, N4450);
and AND3 (N9961, N9950, N9115, N1631);
buf BUF1 (N9962, N9945);
or OR3 (N9963, N9958, N8645, N6009);
or OR3 (N9964, N9921, N2956, N7170);
or OR3 (N9965, N9951, N845, N1680);
xor XOR2 (N9966, N9964, N3891);
not NOT1 (N9967, N9954);
and AND2 (N9968, N9944, N7004);
buf BUF1 (N9969, N9966);
not NOT1 (N9970, N9969);
or OR2 (N9971, N9963, N6783);
xor XOR2 (N9972, N9968, N5510);
and AND2 (N9973, N9967, N9477);
xor XOR2 (N9974, N9955, N347);
not NOT1 (N9975, N9972);
not NOT1 (N9976, N9962);
or OR2 (N9977, N9975, N3698);
nor NOR2 (N9978, N9960, N6102);
nor NOR2 (N9979, N9965, N3915);
buf BUF1 (N9980, N9970);
nand NAND2 (N9981, N9961, N9887);
not NOT1 (N9982, N9977);
xor XOR2 (N9983, N9980, N3712);
nor NOR2 (N9984, N9974, N9213);
xor XOR2 (N9985, N9982, N6629);
and AND4 (N9986, N9979, N2498, N7071, N7309);
nor NOR3 (N9987, N9985, N9959, N9752);
or OR3 (N9988, N1793, N5645, N5721);
buf BUF1 (N9989, N9981);
and AND2 (N9990, N9984, N4359);
not NOT1 (N9991, N9986);
nor NOR4 (N9992, N9989, N8647, N3113, N3648);
or OR3 (N9993, N9988, N9431, N268);
nor NOR4 (N9994, N9971, N9628, N8326, N6306);
and AND2 (N9995, N9994, N2188);
nand NAND2 (N9996, N9990, N7338);
and AND2 (N9997, N9996, N3795);
and AND3 (N9998, N9983, N6672, N627);
or OR2 (N9999, N9987, N7511);
nand NAND4 (N10000, N9997, N3053, N6028, N8665);
buf BUF1 (N10001, N9993);
buf BUF1 (N10002, N9978);
or OR3 (N10003, N9973, N6757, N2401);
xor XOR2 (N10004, N10002, N1226);
nor NOR3 (N10005, N10004, N4887, N1811);
xor XOR2 (N10006, N9976, N9565);
not NOT1 (N10007, N10001);
xor XOR2 (N10008, N9998, N9099);
not NOT1 (N10009, N9999);
and AND3 (N10010, N10006, N7852, N3212);
nor NOR4 (N10011, N10010, N7829, N6939, N3274);
nor NOR3 (N10012, N10011, N6903, N2557);
xor XOR2 (N10013, N10005, N8202);
not NOT1 (N10014, N10007);
and AND3 (N10015, N10000, N5190, N3114);
xor XOR2 (N10016, N10015, N3467);
nor NOR2 (N10017, N10008, N5992);
nor NOR4 (N10018, N10016, N9618, N6784, N2743);
not NOT1 (N10019, N10014);
or OR4 (N10020, N10013, N7272, N8467, N3257);
and AND2 (N10021, N10012, N1958);
buf BUF1 (N10022, N10021);
not NOT1 (N10023, N10022);
nor NOR2 (N10024, N10023, N4573);
nor NOR2 (N10025, N10009, N6491);
xor XOR2 (N10026, N10024, N4295);
or OR2 (N10027, N9991, N3222);
buf BUF1 (N10028, N9992);
xor XOR2 (N10029, N10025, N4193);
nand NAND3 (N10030, N10027, N8743, N9193);
xor XOR2 (N10031, N10026, N7304);
buf BUF1 (N10032, N10031);
not NOT1 (N10033, N10003);
nand NAND3 (N10034, N10020, N861, N116);
not NOT1 (N10035, N10032);
buf BUF1 (N10036, N10034);
or OR2 (N10037, N10019, N1459);
and AND4 (N10038, N10017, N5756, N356, N6533);
buf BUF1 (N10039, N10035);
nand NAND2 (N10040, N10030, N7689);
buf BUF1 (N10041, N10039);
and AND2 (N10042, N10041, N5937);
nand NAND4 (N10043, N10038, N4205, N7165, N9096);
buf BUF1 (N10044, N10029);
and AND4 (N10045, N10042, N5896, N533, N6869);
nand NAND2 (N10046, N10044, N4396);
nor NOR3 (N10047, N10040, N3288, N7499);
buf BUF1 (N10048, N10018);
or OR4 (N10049, N10036, N4611, N9619, N6252);
buf BUF1 (N10050, N10028);
nor NOR3 (N10051, N10047, N8855, N1695);
nand NAND2 (N10052, N10045, N7181);
nor NOR3 (N10053, N10051, N3280, N772);
nor NOR3 (N10054, N10033, N3009, N8147);
not NOT1 (N10055, N10053);
buf BUF1 (N10056, N10054);
xor XOR2 (N10057, N10049, N9500);
not NOT1 (N10058, N10037);
nand NAND3 (N10059, N10056, N1411, N4170);
nor NOR3 (N10060, N10058, N9802, N115);
not NOT1 (N10061, N10057);
nor NOR4 (N10062, N10055, N4528, N5717, N1960);
not NOT1 (N10063, N10059);
nor NOR3 (N10064, N10052, N9839, N2099);
nand NAND3 (N10065, N10060, N5944, N1100);
or OR4 (N10066, N10043, N6986, N5868, N2687);
and AND4 (N10067, N10066, N468, N7942, N2607);
xor XOR2 (N10068, N10050, N1737);
nor NOR3 (N10069, N10062, N884, N8363);
buf BUF1 (N10070, N10064);
not NOT1 (N10071, N10070);
not NOT1 (N10072, N10061);
nor NOR2 (N10073, N10069, N6968);
nand NAND3 (N10074, N10046, N4716, N7704);
or OR3 (N10075, N9995, N3231, N5530);
nand NAND4 (N10076, N10048, N7450, N6886, N9348);
not NOT1 (N10077, N10068);
buf BUF1 (N10078, N10073);
nor NOR2 (N10079, N10067, N162);
and AND4 (N10080, N10077, N8291, N1888, N962);
or OR2 (N10081, N10072, N8675);
or OR4 (N10082, N10081, N9327, N5812, N7737);
not NOT1 (N10083, N10079);
and AND4 (N10084, N10063, N849, N2749, N6790);
and AND4 (N10085, N10080, N3565, N902, N453);
buf BUF1 (N10086, N10071);
not NOT1 (N10087, N10086);
xor XOR2 (N10088, N10085, N6630);
buf BUF1 (N10089, N10065);
buf BUF1 (N10090, N10075);
nand NAND3 (N10091, N10078, N4979, N1640);
not NOT1 (N10092, N10082);
nand NAND2 (N10093, N10092, N3693);
nand NAND4 (N10094, N10091, N6832, N8810, N4185);
buf BUF1 (N10095, N10093);
nand NAND2 (N10096, N10089, N1298);
nand NAND4 (N10097, N10096, N2920, N8723, N216);
and AND4 (N10098, N10074, N4157, N4679, N932);
buf BUF1 (N10099, N10097);
xor XOR2 (N10100, N10094, N1109);
nand NAND4 (N10101, N10099, N6395, N2397, N8577);
not NOT1 (N10102, N10084);
not NOT1 (N10103, N10087);
buf BUF1 (N10104, N10098);
and AND4 (N10105, N10102, N7460, N369, N3209);
or OR2 (N10106, N10101, N1769);
nand NAND3 (N10107, N10103, N645, N9600);
nand NAND2 (N10108, N10100, N5287);
not NOT1 (N10109, N10083);
or OR4 (N10110, N10109, N1021, N3791, N7325);
buf BUF1 (N10111, N10106);
not NOT1 (N10112, N10111);
and AND4 (N10113, N10088, N9517, N4003, N2214);
and AND3 (N10114, N10110, N7103, N6147);
nand NAND2 (N10115, N10108, N6529);
or OR3 (N10116, N10113, N8159, N5879);
nand NAND2 (N10117, N10114, N8205);
nand NAND3 (N10118, N10112, N7694, N4127);
nand NAND4 (N10119, N10095, N3039, N8042, N8395);
and AND4 (N10120, N10076, N1406, N6705, N6710);
xor XOR2 (N10121, N10118, N9341);
and AND2 (N10122, N10120, N9848);
nand NAND2 (N10123, N10122, N1448);
buf BUF1 (N10124, N10119);
nor NOR4 (N10125, N10104, N3708, N2582, N3894);
and AND2 (N10126, N10116, N6266);
xor XOR2 (N10127, N10125, N5079);
nand NAND4 (N10128, N10124, N1424, N7683, N7531);
and AND2 (N10129, N10090, N349);
or OR3 (N10130, N10107, N3139, N2092);
not NOT1 (N10131, N10128);
not NOT1 (N10132, N10121);
nand NAND3 (N10133, N10129, N4032, N2155);
not NOT1 (N10134, N10126);
buf BUF1 (N10135, N10105);
nor NOR2 (N10136, N10131, N7133);
not NOT1 (N10137, N10136);
xor XOR2 (N10138, N10135, N4085);
buf BUF1 (N10139, N10117);
and AND3 (N10140, N10132, N9323, N9629);
not NOT1 (N10141, N10123);
nor NOR3 (N10142, N10127, N4932, N5644);
not NOT1 (N10143, N10130);
buf BUF1 (N10144, N10133);
nor NOR3 (N10145, N10144, N1899, N7213);
not NOT1 (N10146, N10145);
not NOT1 (N10147, N10146);
nor NOR4 (N10148, N10138, N3387, N1340, N4682);
xor XOR2 (N10149, N10115, N2834);
buf BUF1 (N10150, N10143);
or OR3 (N10151, N10148, N9581, N2633);
and AND4 (N10152, N10142, N6078, N9529, N1218);
or OR2 (N10153, N10150, N420);
nor NOR4 (N10154, N10153, N3764, N5133, N3084);
or OR3 (N10155, N10152, N7308, N3203);
not NOT1 (N10156, N10140);
nand NAND3 (N10157, N10149, N9294, N7428);
and AND4 (N10158, N10157, N5359, N1225, N3456);
xor XOR2 (N10159, N10156, N4523);
xor XOR2 (N10160, N10154, N4632);
nor NOR4 (N10161, N10159, N4754, N9170, N1352);
nor NOR3 (N10162, N10151, N1366, N3916);
not NOT1 (N10163, N10141);
or OR4 (N10164, N10160, N8784, N1901, N1607);
xor XOR2 (N10165, N10147, N8694);
nand NAND3 (N10166, N10134, N8745, N7265);
not NOT1 (N10167, N10162);
not NOT1 (N10168, N10161);
xor XOR2 (N10169, N10155, N2919);
and AND3 (N10170, N10167, N88, N4042);
buf BUF1 (N10171, N10169);
not NOT1 (N10172, N10163);
or OR4 (N10173, N10166, N2721, N5533, N3258);
or OR2 (N10174, N10139, N8841);
xor XOR2 (N10175, N10164, N1610);
xor XOR2 (N10176, N10172, N5749);
and AND2 (N10177, N10176, N5362);
and AND3 (N10178, N10170, N7662, N751);
nor NOR4 (N10179, N10178, N5732, N653, N1172);
buf BUF1 (N10180, N10175);
buf BUF1 (N10181, N10177);
nand NAND2 (N10182, N10174, N4204);
xor XOR2 (N10183, N10180, N4970);
or OR2 (N10184, N10179, N5528);
or OR3 (N10185, N10158, N9705, N6137);
nor NOR2 (N10186, N10165, N3525);
and AND4 (N10187, N10137, N9679, N7620, N2525);
xor XOR2 (N10188, N10186, N8274);
nand NAND2 (N10189, N10173, N6219);
or OR3 (N10190, N10171, N2632, N6110);
nand NAND4 (N10191, N10189, N81, N9998, N4398);
not NOT1 (N10192, N10183);
and AND3 (N10193, N10188, N4461, N7102);
xor XOR2 (N10194, N10184, N6742);
xor XOR2 (N10195, N10182, N6157);
nor NOR3 (N10196, N10185, N171, N1480);
not NOT1 (N10197, N10190);
nor NOR2 (N10198, N10187, N1307);
buf BUF1 (N10199, N10181);
and AND2 (N10200, N10168, N7850);
and AND3 (N10201, N10200, N4263, N3166);
nand NAND3 (N10202, N10198, N5995, N2378);
nor NOR3 (N10203, N10197, N3915, N8186);
or OR2 (N10204, N10191, N5402);
or OR3 (N10205, N10196, N9725, N4203);
nand NAND3 (N10206, N10193, N9002, N3839);
or OR2 (N10207, N10194, N3161);
nand NAND2 (N10208, N10195, N312);
nor NOR3 (N10209, N10201, N3950, N9923);
nand NAND4 (N10210, N10207, N10040, N7117, N2009);
nand NAND4 (N10211, N10209, N5114, N97, N2296);
xor XOR2 (N10212, N10208, N9882);
buf BUF1 (N10213, N10205);
buf BUF1 (N10214, N10204);
xor XOR2 (N10215, N10210, N3107);
and AND2 (N10216, N10215, N6482);
or OR2 (N10217, N10212, N638);
and AND3 (N10218, N10213, N2134, N580);
buf BUF1 (N10219, N10202);
and AND2 (N10220, N10214, N4872);
or OR2 (N10221, N10211, N3224);
not NOT1 (N10222, N10199);
nor NOR2 (N10223, N10203, N4958);
and AND2 (N10224, N10218, N5364);
buf BUF1 (N10225, N10219);
or OR4 (N10226, N10221, N5624, N155, N5579);
and AND4 (N10227, N10192, N3549, N3857, N6700);
nand NAND3 (N10228, N10216, N8280, N1115);
nand NAND2 (N10229, N10227, N7488);
xor XOR2 (N10230, N10228, N3300);
buf BUF1 (N10231, N10229);
or OR4 (N10232, N10217, N8750, N1201, N2648);
xor XOR2 (N10233, N10232, N8875);
and AND2 (N10234, N10224, N5857);
nand NAND4 (N10235, N10220, N9328, N9164, N2734);
and AND2 (N10236, N10234, N2876);
nand NAND2 (N10237, N10206, N5695);
buf BUF1 (N10238, N10233);
not NOT1 (N10239, N10222);
not NOT1 (N10240, N10223);
xor XOR2 (N10241, N10236, N9335);
or OR3 (N10242, N10241, N5134, N348);
nor NOR2 (N10243, N10226, N3388);
buf BUF1 (N10244, N10225);
not NOT1 (N10245, N10243);
nor NOR4 (N10246, N10245, N4729, N4646, N2661);
nand NAND3 (N10247, N10239, N5816, N7730);
nand NAND4 (N10248, N10240, N4688, N7643, N10084);
nand NAND4 (N10249, N10231, N7937, N6936, N162);
or OR3 (N10250, N10238, N4179, N276);
xor XOR2 (N10251, N10249, N780);
nor NOR3 (N10252, N10247, N652, N3766);
and AND3 (N10253, N10242, N3521, N3533);
nor NOR2 (N10254, N10230, N3125);
buf BUF1 (N10255, N10235);
nand NAND2 (N10256, N10253, N9076);
not NOT1 (N10257, N10246);
nand NAND4 (N10258, N10251, N2145, N3436, N1041);
xor XOR2 (N10259, N10254, N9314);
not NOT1 (N10260, N10250);
nand NAND4 (N10261, N10260, N2219, N4365, N3378);
and AND4 (N10262, N10237, N1070, N9203, N5474);
or OR2 (N10263, N10248, N300);
buf BUF1 (N10264, N10252);
nor NOR2 (N10265, N10262, N977);
and AND4 (N10266, N10256, N2143, N230, N6072);
and AND2 (N10267, N10255, N8263);
nand NAND3 (N10268, N10259, N1455, N377);
and AND4 (N10269, N10265, N8391, N2534, N8165);
and AND4 (N10270, N10268, N2434, N9823, N7467);
nor NOR3 (N10271, N10258, N3750, N529);
not NOT1 (N10272, N10261);
buf BUF1 (N10273, N10270);
xor XOR2 (N10274, N10264, N5152);
or OR4 (N10275, N10272, N1687, N10096, N2503);
not NOT1 (N10276, N10244);
buf BUF1 (N10277, N10266);
nor NOR4 (N10278, N10277, N6680, N5697, N153);
not NOT1 (N10279, N10271);
buf BUF1 (N10280, N10267);
xor XOR2 (N10281, N10278, N9015);
or OR3 (N10282, N10276, N6301, N8911);
and AND3 (N10283, N10273, N2351, N1539);
and AND4 (N10284, N10269, N52, N6013, N2985);
xor XOR2 (N10285, N10279, N549);
and AND4 (N10286, N10275, N1537, N1169, N1619);
and AND4 (N10287, N10285, N7823, N473, N1781);
not NOT1 (N10288, N10283);
and AND4 (N10289, N10288, N6512, N8578, N2386);
buf BUF1 (N10290, N10281);
nor NOR4 (N10291, N10284, N1082, N9757, N1082);
nand NAND3 (N10292, N10282, N5688, N3396);
nor NOR4 (N10293, N10257, N968, N2662, N6395);
nor NOR2 (N10294, N10292, N6531);
buf BUF1 (N10295, N10263);
or OR2 (N10296, N10291, N3633);
nor NOR2 (N10297, N10274, N1090);
xor XOR2 (N10298, N10286, N975);
not NOT1 (N10299, N10289);
nor NOR4 (N10300, N10293, N8788, N5048, N3963);
nand NAND4 (N10301, N10290, N10258, N8777, N4643);
not NOT1 (N10302, N10297);
buf BUF1 (N10303, N10302);
or OR4 (N10304, N10287, N722, N10215, N4926);
and AND2 (N10305, N10299, N2750);
nor NOR3 (N10306, N10300, N1977, N2368);
xor XOR2 (N10307, N10301, N7398);
and AND2 (N10308, N10294, N2527);
xor XOR2 (N10309, N10306, N5847);
buf BUF1 (N10310, N10280);
not NOT1 (N10311, N10307);
or OR2 (N10312, N10296, N2933);
buf BUF1 (N10313, N10308);
and AND2 (N10314, N10304, N8054);
nor NOR3 (N10315, N10314, N4644, N3385);
xor XOR2 (N10316, N10303, N3495);
buf BUF1 (N10317, N10313);
and AND2 (N10318, N10298, N3624);
nor NOR4 (N10319, N10312, N3900, N5618, N8236);
nand NAND4 (N10320, N10317, N5915, N9280, N2215);
nand NAND3 (N10321, N10311, N8698, N5298);
or OR4 (N10322, N10318, N5204, N8704, N2987);
and AND4 (N10323, N10322, N5465, N4617, N166);
not NOT1 (N10324, N10305);
not NOT1 (N10325, N10321);
buf BUF1 (N10326, N10323);
or OR3 (N10327, N10320, N629, N7723);
and AND4 (N10328, N10309, N2267, N7730, N1386);
nor NOR3 (N10329, N10295, N8214, N5098);
buf BUF1 (N10330, N10328);
and AND3 (N10331, N10326, N1814, N591);
xor XOR2 (N10332, N10310, N9205);
and AND2 (N10333, N10327, N8704);
or OR2 (N10334, N10324, N4416);
nor NOR2 (N10335, N10319, N9759);
nand NAND4 (N10336, N10331, N4046, N6656, N7809);
and AND3 (N10337, N10316, N9974, N8280);
nand NAND3 (N10338, N10336, N8089, N2728);
xor XOR2 (N10339, N10330, N9398);
or OR2 (N10340, N10332, N9008);
xor XOR2 (N10341, N10325, N8519);
xor XOR2 (N10342, N10335, N3466);
and AND3 (N10343, N10333, N1716, N7940);
xor XOR2 (N10344, N10343, N3740);
xor XOR2 (N10345, N10339, N4819);
or OR2 (N10346, N10338, N8527);
nor NOR2 (N10347, N10337, N1230);
not NOT1 (N10348, N10329);
xor XOR2 (N10349, N10346, N7877);
and AND3 (N10350, N10341, N5840, N7689);
nand NAND2 (N10351, N10349, N4740);
nand NAND3 (N10352, N10342, N3966, N781);
nor NOR4 (N10353, N10334, N6600, N7212, N1757);
nand NAND2 (N10354, N10348, N271);
or OR2 (N10355, N10352, N5783);
xor XOR2 (N10356, N10355, N5671);
nand NAND4 (N10357, N10347, N6979, N6955, N9776);
and AND3 (N10358, N10340, N6855, N6469);
nand NAND4 (N10359, N10357, N710, N7101, N3399);
xor XOR2 (N10360, N10344, N1448);
nor NOR3 (N10361, N10356, N1358, N8641);
nor NOR4 (N10362, N10358, N3794, N7274, N6009);
and AND3 (N10363, N10361, N9082, N130);
nor NOR2 (N10364, N10362, N8563);
buf BUF1 (N10365, N10354);
nor NOR4 (N10366, N10360, N5532, N7959, N8933);
not NOT1 (N10367, N10364);
and AND2 (N10368, N10367, N3376);
nor NOR3 (N10369, N10366, N7377, N7379);
nor NOR4 (N10370, N10350, N363, N2522, N7093);
xor XOR2 (N10371, N10368, N4209);
not NOT1 (N10372, N10351);
nand NAND2 (N10373, N10345, N4292);
not NOT1 (N10374, N10363);
buf BUF1 (N10375, N10374);
not NOT1 (N10376, N10369);
or OR4 (N10377, N10376, N2305, N1190, N8143);
not NOT1 (N10378, N10370);
nor NOR3 (N10379, N10365, N3945, N7027);
not NOT1 (N10380, N10353);
and AND2 (N10381, N10375, N2686);
nand NAND2 (N10382, N10373, N3592);
or OR4 (N10383, N10380, N9819, N7749, N6002);
not NOT1 (N10384, N10381);
and AND2 (N10385, N10372, N523);
and AND3 (N10386, N10378, N10112, N6516);
nand NAND3 (N10387, N10359, N6023, N2262);
xor XOR2 (N10388, N10384, N3072);
nor NOR4 (N10389, N10371, N5059, N2202, N4239);
xor XOR2 (N10390, N10387, N4892);
nand NAND2 (N10391, N10382, N2419);
and AND3 (N10392, N10379, N3481, N5332);
and AND4 (N10393, N10389, N9951, N7821, N7740);
nor NOR2 (N10394, N10386, N6258);
xor XOR2 (N10395, N10390, N3011);
or OR2 (N10396, N10393, N7135);
nor NOR2 (N10397, N10383, N7030);
or OR3 (N10398, N10392, N242, N9459);
xor XOR2 (N10399, N10377, N4455);
and AND3 (N10400, N10398, N331, N3487);
nor NOR3 (N10401, N10388, N5158, N1006);
buf BUF1 (N10402, N10315);
not NOT1 (N10403, N10391);
nor NOR4 (N10404, N10399, N2192, N326, N9714);
not NOT1 (N10405, N10400);
nand NAND4 (N10406, N10405, N6323, N8896, N10107);
buf BUF1 (N10407, N10404);
nand NAND2 (N10408, N10396, N984);
buf BUF1 (N10409, N10408);
nor NOR2 (N10410, N10395, N4090);
nor NOR2 (N10411, N10385, N6661);
nor NOR4 (N10412, N10406, N10163, N7014, N5922);
or OR2 (N10413, N10394, N10234);
nor NOR3 (N10414, N10402, N4659, N7235);
and AND3 (N10415, N10401, N1054, N7923);
nor NOR4 (N10416, N10397, N4928, N1963, N7336);
buf BUF1 (N10417, N10403);
and AND2 (N10418, N10411, N3483);
nand NAND4 (N10419, N10410, N3033, N8543, N156);
nand NAND2 (N10420, N10417, N3956);
nor NOR2 (N10421, N10419, N2896);
nor NOR3 (N10422, N10418, N7918, N5296);
nor NOR2 (N10423, N10414, N6766);
or OR2 (N10424, N10415, N10349);
or OR3 (N10425, N10423, N174, N2644);
nand NAND3 (N10426, N10412, N2418, N2840);
xor XOR2 (N10427, N10424, N9745);
nor NOR2 (N10428, N10425, N3419);
buf BUF1 (N10429, N10407);
buf BUF1 (N10430, N10428);
nand NAND2 (N10431, N10429, N5530);
buf BUF1 (N10432, N10426);
xor XOR2 (N10433, N10416, N3055);
buf BUF1 (N10434, N10409);
buf BUF1 (N10435, N10434);
not NOT1 (N10436, N10420);
xor XOR2 (N10437, N10436, N6702);
nor NOR3 (N10438, N10431, N6061, N8609);
and AND2 (N10439, N10438, N7659);
or OR4 (N10440, N10435, N1077, N8197, N8799);
buf BUF1 (N10441, N10430);
buf BUF1 (N10442, N10440);
nor NOR3 (N10443, N10422, N7059, N1591);
or OR4 (N10444, N10427, N9673, N5241, N4759);
not NOT1 (N10445, N10432);
or OR4 (N10446, N10445, N3237, N8569, N9172);
buf BUF1 (N10447, N10439);
nand NAND3 (N10448, N10433, N9245, N6266);
xor XOR2 (N10449, N10444, N9152);
and AND3 (N10450, N10443, N3963, N3943);
not NOT1 (N10451, N10450);
nand NAND4 (N10452, N10437, N6657, N2890, N6959);
nor NOR4 (N10453, N10442, N3792, N7139, N6703);
and AND3 (N10454, N10413, N4033, N10054);
and AND2 (N10455, N10447, N4398);
or OR2 (N10456, N10446, N3567);
nand NAND2 (N10457, N10455, N9849);
and AND4 (N10458, N10449, N4896, N3786, N2565);
nand NAND2 (N10459, N10454, N3574);
nand NAND3 (N10460, N10453, N6577, N8785);
xor XOR2 (N10461, N10421, N9581);
nand NAND4 (N10462, N10457, N901, N2831, N989);
buf BUF1 (N10463, N10460);
or OR2 (N10464, N10456, N8161);
or OR2 (N10465, N10448, N4488);
nand NAND4 (N10466, N10463, N8103, N8454, N721);
nand NAND2 (N10467, N10466, N1627);
nand NAND2 (N10468, N10441, N10357);
or OR2 (N10469, N10459, N7730);
and AND3 (N10470, N10462, N1638, N5593);
nand NAND4 (N10471, N10458, N801, N5522, N7384);
xor XOR2 (N10472, N10451, N9351);
buf BUF1 (N10473, N10471);
buf BUF1 (N10474, N10464);
nor NOR2 (N10475, N10465, N3821);
and AND3 (N10476, N10452, N762, N3412);
buf BUF1 (N10477, N10470);
and AND3 (N10478, N10461, N6494, N7993);
and AND3 (N10479, N10474, N7754, N9178);
buf BUF1 (N10480, N10468);
xor XOR2 (N10481, N10479, N6331);
xor XOR2 (N10482, N10476, N1809);
not NOT1 (N10483, N10482);
nand NAND4 (N10484, N10469, N8529, N6499, N10037);
not NOT1 (N10485, N10467);
and AND2 (N10486, N10481, N9195);
not NOT1 (N10487, N10478);
nand NAND4 (N10488, N10486, N3607, N4258, N5568);
or OR4 (N10489, N10480, N5452, N782, N9811);
nor NOR4 (N10490, N10488, N2001, N1882, N8834);
xor XOR2 (N10491, N10475, N1046);
not NOT1 (N10492, N10487);
nand NAND2 (N10493, N10483, N1247);
nor NOR4 (N10494, N10492, N5216, N3609, N6291);
and AND2 (N10495, N10490, N7718);
and AND2 (N10496, N10472, N3613);
not NOT1 (N10497, N10495);
and AND3 (N10498, N10489, N4916, N9312);
buf BUF1 (N10499, N10484);
or OR2 (N10500, N10494, N5021);
buf BUF1 (N10501, N10498);
not NOT1 (N10502, N10496);
not NOT1 (N10503, N10473);
buf BUF1 (N10504, N10485);
not NOT1 (N10505, N10491);
buf BUF1 (N10506, N10499);
not NOT1 (N10507, N10502);
buf BUF1 (N10508, N10501);
xor XOR2 (N10509, N10477, N7699);
nor NOR3 (N10510, N10500, N3418, N3013);
buf BUF1 (N10511, N10503);
nand NAND3 (N10512, N10507, N3097, N9772);
or OR4 (N10513, N10493, N2064, N212, N3344);
xor XOR2 (N10514, N10512, N7742);
or OR4 (N10515, N10505, N6132, N10285, N6172);
xor XOR2 (N10516, N10515, N9774);
buf BUF1 (N10517, N10511);
nand NAND3 (N10518, N10517, N8669, N8414);
xor XOR2 (N10519, N10506, N7334);
xor XOR2 (N10520, N10508, N3889);
nor NOR3 (N10521, N10518, N7970, N10346);
xor XOR2 (N10522, N10497, N5290);
and AND2 (N10523, N10519, N4474);
not NOT1 (N10524, N10510);
not NOT1 (N10525, N10513);
buf BUF1 (N10526, N10524);
and AND3 (N10527, N10526, N918, N7972);
nand NAND4 (N10528, N10522, N5954, N1514, N6880);
or OR3 (N10529, N10523, N3765, N74);
or OR2 (N10530, N10528, N8650);
or OR3 (N10531, N10527, N2682, N10265);
nor NOR3 (N10532, N10514, N7794, N1525);
nand NAND2 (N10533, N10521, N5225);
nor NOR3 (N10534, N10533, N71, N1108);
not NOT1 (N10535, N10532);
nor NOR4 (N10536, N10529, N3093, N4784, N3860);
and AND4 (N10537, N10535, N8568, N3710, N3863);
nand NAND2 (N10538, N10520, N2819);
nand NAND3 (N10539, N10516, N3214, N3994);
buf BUF1 (N10540, N10531);
not NOT1 (N10541, N10536);
xor XOR2 (N10542, N10525, N5148);
buf BUF1 (N10543, N10539);
buf BUF1 (N10544, N10509);
nand NAND2 (N10545, N10541, N1197);
or OR4 (N10546, N10534, N3504, N7941, N5118);
xor XOR2 (N10547, N10545, N1385);
not NOT1 (N10548, N10530);
and AND4 (N10549, N10548, N938, N9871, N7322);
nor NOR2 (N10550, N10546, N3414);
nand NAND3 (N10551, N10540, N313, N9125);
nor NOR4 (N10552, N10544, N2452, N243, N9851);
nand NAND3 (N10553, N10537, N1487, N7039);
buf BUF1 (N10554, N10553);
nand NAND4 (N10555, N10549, N7907, N7586, N1661);
nand NAND4 (N10556, N10538, N5060, N8767, N5044);
nor NOR3 (N10557, N10554, N4563, N10373);
nor NOR3 (N10558, N10555, N1237, N7813);
not NOT1 (N10559, N10557);
nand NAND4 (N10560, N10551, N9478, N9994, N3857);
nand NAND2 (N10561, N10550, N2677);
nor NOR4 (N10562, N10547, N8631, N6312, N2674);
and AND2 (N10563, N10543, N3012);
nor NOR3 (N10564, N10542, N3707, N3999);
or OR3 (N10565, N10561, N2098, N8212);
xor XOR2 (N10566, N10563, N2883);
buf BUF1 (N10567, N10565);
nor NOR4 (N10568, N10567, N9595, N9561, N6389);
xor XOR2 (N10569, N10558, N3940);
and AND4 (N10570, N10566, N2199, N79, N6398);
nor NOR2 (N10571, N10560, N472);
buf BUF1 (N10572, N10559);
and AND3 (N10573, N10564, N10145, N9098);
nor NOR4 (N10574, N10573, N9712, N5009, N6499);
nor NOR3 (N10575, N10552, N4803, N2279);
and AND3 (N10576, N10556, N4634, N6998);
nor NOR4 (N10577, N10504, N5815, N4358, N7179);
or OR3 (N10578, N10571, N298, N9290);
buf BUF1 (N10579, N10574);
xor XOR2 (N10580, N10572, N8358);
not NOT1 (N10581, N10576);
nor NOR3 (N10582, N10577, N5746, N1468);
not NOT1 (N10583, N10575);
and AND4 (N10584, N10583, N5586, N10378, N1215);
not NOT1 (N10585, N10582);
not NOT1 (N10586, N10581);
xor XOR2 (N10587, N10585, N7942);
xor XOR2 (N10588, N10587, N2475);
buf BUF1 (N10589, N10579);
and AND3 (N10590, N10568, N9056, N6106);
nand NAND2 (N10591, N10584, N8670);
nand NAND2 (N10592, N10588, N5655);
nand NAND4 (N10593, N10589, N504, N6436, N3259);
not NOT1 (N10594, N10580);
nand NAND3 (N10595, N10562, N9451, N3818);
nand NAND4 (N10596, N10590, N4018, N8193, N6895);
and AND2 (N10597, N10596, N9096);
or OR4 (N10598, N10592, N9474, N7692, N2876);
xor XOR2 (N10599, N10578, N9736);
and AND4 (N10600, N10586, N6946, N6307, N10499);
nor NOR2 (N10601, N10595, N452);
or OR4 (N10602, N10599, N1042, N9053, N9196);
or OR4 (N10603, N10591, N9861, N6062, N1695);
and AND3 (N10604, N10601, N8615, N8987);
not NOT1 (N10605, N10603);
and AND4 (N10606, N10597, N3635, N9909, N2876);
or OR2 (N10607, N10594, N9825);
or OR2 (N10608, N10593, N7999);
xor XOR2 (N10609, N10602, N2540);
buf BUF1 (N10610, N10569);
buf BUF1 (N10611, N10610);
xor XOR2 (N10612, N10605, N2495);
or OR4 (N10613, N10609, N9180, N8350, N9366);
nand NAND2 (N10614, N10600, N4675);
or OR4 (N10615, N10614, N4053, N9305, N8218);
nor NOR4 (N10616, N10615, N1159, N8119, N4509);
not NOT1 (N10617, N10612);
and AND2 (N10618, N10606, N9555);
not NOT1 (N10619, N10611);
not NOT1 (N10620, N10613);
nand NAND4 (N10621, N10608, N4420, N10095, N1127);
and AND2 (N10622, N10616, N5360);
buf BUF1 (N10623, N10621);
nand NAND4 (N10624, N10607, N4621, N4628, N7922);
xor XOR2 (N10625, N10623, N3102);
nor NOR2 (N10626, N10625, N6201);
or OR4 (N10627, N10604, N999, N6423, N9174);
nor NOR4 (N10628, N10619, N1155, N7922, N8420);
not NOT1 (N10629, N10598);
and AND4 (N10630, N10629, N745, N5752, N9297);
xor XOR2 (N10631, N10630, N9252);
xor XOR2 (N10632, N10617, N4196);
or OR3 (N10633, N10570, N5745, N10539);
xor XOR2 (N10634, N10620, N6183);
nor NOR2 (N10635, N10618, N10212);
or OR3 (N10636, N10628, N9345, N9503);
xor XOR2 (N10637, N10632, N8000);
not NOT1 (N10638, N10631);
buf BUF1 (N10639, N10633);
not NOT1 (N10640, N10635);
nor NOR3 (N10641, N10624, N5766, N618);
buf BUF1 (N10642, N10639);
nand NAND2 (N10643, N10641, N2490);
buf BUF1 (N10644, N10622);
not NOT1 (N10645, N10634);
nor NOR4 (N10646, N10644, N5286, N1661, N10119);
nor NOR4 (N10647, N10627, N2957, N9402, N6295);
and AND3 (N10648, N10637, N10457, N1889);
buf BUF1 (N10649, N10636);
nand NAND4 (N10650, N10645, N8214, N3973, N4783);
or OR4 (N10651, N10643, N232, N1399, N9466);
xor XOR2 (N10652, N10642, N1304);
or OR2 (N10653, N10647, N8987);
not NOT1 (N10654, N10649);
and AND2 (N10655, N10648, N10407);
nand NAND2 (N10656, N10654, N10626);
not NOT1 (N10657, N4215);
not NOT1 (N10658, N10646);
and AND2 (N10659, N10653, N9458);
nand NAND4 (N10660, N10656, N8109, N6541, N6356);
nor NOR2 (N10661, N10657, N2300);
nor NOR3 (N10662, N10652, N7122, N2057);
buf BUF1 (N10663, N10662);
or OR4 (N10664, N10659, N8512, N848, N7572);
not NOT1 (N10665, N10658);
or OR2 (N10666, N10665, N8433);
xor XOR2 (N10667, N10651, N194);
not NOT1 (N10668, N10664);
xor XOR2 (N10669, N10638, N628);
buf BUF1 (N10670, N10661);
not NOT1 (N10671, N10655);
nand NAND2 (N10672, N10660, N10048);
nor NOR4 (N10673, N10671, N5384, N5342, N3739);
nor NOR3 (N10674, N10670, N4119, N1464);
and AND3 (N10675, N10669, N688, N8276);
buf BUF1 (N10676, N10675);
buf BUF1 (N10677, N10666);
not NOT1 (N10678, N10673);
xor XOR2 (N10679, N10650, N1716);
and AND2 (N10680, N10676, N1350);
not NOT1 (N10681, N10640);
and AND4 (N10682, N10678, N6891, N6653, N1381);
xor XOR2 (N10683, N10679, N2596);
xor XOR2 (N10684, N10677, N6422);
xor XOR2 (N10685, N10682, N10229);
nand NAND3 (N10686, N10685, N5833, N7937);
nor NOR3 (N10687, N10686, N7831, N19);
nand NAND4 (N10688, N10681, N3648, N8096, N6386);
xor XOR2 (N10689, N10663, N5354);
xor XOR2 (N10690, N10683, N7167);
xor XOR2 (N10691, N10680, N6919);
buf BUF1 (N10692, N10674);
nor NOR2 (N10693, N10692, N7909);
buf BUF1 (N10694, N10687);
nand NAND4 (N10695, N10688, N5262, N6457, N9475);
not NOT1 (N10696, N10693);
nor NOR2 (N10697, N10690, N7259);
nand NAND4 (N10698, N10696, N7180, N1472, N7073);
buf BUF1 (N10699, N10684);
or OR2 (N10700, N10667, N3260);
nor NOR2 (N10701, N10697, N6437);
nor NOR4 (N10702, N10689, N9051, N10524, N9320);
xor XOR2 (N10703, N10701, N3984);
not NOT1 (N10704, N10695);
nor NOR3 (N10705, N10694, N8868, N6822);
buf BUF1 (N10706, N10703);
nand NAND4 (N10707, N10698, N5440, N9546, N3117);
nor NOR3 (N10708, N10707, N10012, N3795);
nand NAND3 (N10709, N10708, N3615, N10278);
or OR2 (N10710, N10702, N5573);
or OR2 (N10711, N10705, N4581);
nor NOR2 (N10712, N10709, N641);
nor NOR2 (N10713, N10706, N4643);
nor NOR4 (N10714, N10699, N7081, N5995, N9695);
nor NOR4 (N10715, N10711, N3875, N3470, N7809);
and AND2 (N10716, N10672, N5871);
buf BUF1 (N10717, N10668);
not NOT1 (N10718, N10704);
and AND4 (N10719, N10714, N1986, N6870, N179);
not NOT1 (N10720, N10700);
and AND2 (N10721, N10720, N10011);
nor NOR3 (N10722, N10718, N1250, N9661);
buf BUF1 (N10723, N10717);
or OR3 (N10724, N10723, N4971, N2492);
not NOT1 (N10725, N10724);
buf BUF1 (N10726, N10721);
not NOT1 (N10727, N10713);
xor XOR2 (N10728, N10725, N6668);
nand NAND2 (N10729, N10722, N10617);
buf BUF1 (N10730, N10715);
xor XOR2 (N10731, N10719, N631);
not NOT1 (N10732, N10726);
or OR3 (N10733, N10732, N9683, N5266);
buf BUF1 (N10734, N10710);
not NOT1 (N10735, N10716);
and AND4 (N10736, N10691, N6797, N6311, N1664);
xor XOR2 (N10737, N10727, N6369);
buf BUF1 (N10738, N10712);
buf BUF1 (N10739, N10728);
xor XOR2 (N10740, N10739, N3332);
not NOT1 (N10741, N10731);
buf BUF1 (N10742, N10738);
nand NAND3 (N10743, N10740, N8405, N4504);
xor XOR2 (N10744, N10729, N4494);
buf BUF1 (N10745, N10730);
nand NAND2 (N10746, N10743, N6482);
or OR3 (N10747, N10735, N7540, N3278);
xor XOR2 (N10748, N10747, N4432);
or OR3 (N10749, N10748, N6785, N8691);
or OR4 (N10750, N10741, N9493, N4439, N4838);
buf BUF1 (N10751, N10734);
nand NAND2 (N10752, N10751, N10327);
xor XOR2 (N10753, N10733, N5450);
not NOT1 (N10754, N10744);
not NOT1 (N10755, N10737);
and AND2 (N10756, N10749, N2922);
nor NOR4 (N10757, N10746, N9784, N2940, N5977);
nor NOR2 (N10758, N10753, N2679);
or OR3 (N10759, N10756, N6254, N3242);
or OR4 (N10760, N10750, N1047, N5517, N9134);
not NOT1 (N10761, N10757);
nor NOR4 (N10762, N10752, N6675, N4661, N3992);
nand NAND4 (N10763, N10759, N8518, N2448, N1893);
and AND4 (N10764, N10736, N4130, N1312, N10457);
buf BUF1 (N10765, N10754);
nor NOR3 (N10766, N10760, N1117, N3310);
nor NOR3 (N10767, N10762, N2512, N9715);
or OR4 (N10768, N10763, N5192, N441, N6568);
nor NOR4 (N10769, N10761, N6643, N3327, N2282);
not NOT1 (N10770, N10755);
and AND2 (N10771, N10745, N8943);
nor NOR3 (N10772, N10769, N4248, N8581);
or OR2 (N10773, N10766, N6326);
xor XOR2 (N10774, N10758, N4154);
xor XOR2 (N10775, N10774, N9700);
or OR4 (N10776, N10765, N736, N823, N8534);
nand NAND3 (N10777, N10768, N8405, N7252);
and AND4 (N10778, N10773, N2009, N7977, N7076);
xor XOR2 (N10779, N10776, N5363);
xor XOR2 (N10780, N10778, N8864);
not NOT1 (N10781, N10742);
xor XOR2 (N10782, N10779, N5873);
buf BUF1 (N10783, N10782);
nand NAND3 (N10784, N10777, N6115, N9418);
buf BUF1 (N10785, N10767);
nand NAND2 (N10786, N10771, N549);
not NOT1 (N10787, N10775);
nand NAND2 (N10788, N10785, N10142);
or OR4 (N10789, N10780, N1983, N2562, N118);
nand NAND4 (N10790, N10772, N1264, N1690, N7946);
not NOT1 (N10791, N10788);
xor XOR2 (N10792, N10764, N251);
buf BUF1 (N10793, N10792);
buf BUF1 (N10794, N10787);
or OR2 (N10795, N10789, N9986);
nand NAND2 (N10796, N10794, N896);
or OR4 (N10797, N10790, N9121, N4885, N9867);
or OR3 (N10798, N10796, N7207, N8200);
buf BUF1 (N10799, N10798);
and AND2 (N10800, N10784, N7322);
xor XOR2 (N10801, N10799, N6651);
nor NOR4 (N10802, N10797, N1103, N3408, N3171);
buf BUF1 (N10803, N10795);
or OR2 (N10804, N10802, N3471);
not NOT1 (N10805, N10804);
not NOT1 (N10806, N10793);
nand NAND4 (N10807, N10791, N2629, N7434, N4240);
nor NOR3 (N10808, N10806, N2035, N9383);
nand NAND4 (N10809, N10770, N2479, N2015, N1129);
nor NOR4 (N10810, N10803, N10600, N6247, N5936);
nor NOR2 (N10811, N10810, N3106);
or OR4 (N10812, N10783, N5920, N10364, N7524);
or OR3 (N10813, N10811, N5452, N7113);
not NOT1 (N10814, N10801);
or OR4 (N10815, N10807, N10046, N4273, N7098);
nand NAND2 (N10816, N10809, N10177);
and AND4 (N10817, N10805, N3137, N3305, N9515);
xor XOR2 (N10818, N10781, N9374);
nor NOR2 (N10819, N10817, N2651);
not NOT1 (N10820, N10819);
buf BUF1 (N10821, N10786);
xor XOR2 (N10822, N10800, N9770);
or OR4 (N10823, N10815, N7757, N7889, N4823);
nor NOR4 (N10824, N10814, N7001, N508, N6652);
or OR3 (N10825, N10823, N1423, N8222);
buf BUF1 (N10826, N10808);
and AND4 (N10827, N10822, N4268, N3695, N3058);
and AND3 (N10828, N10816, N2603, N2258);
or OR4 (N10829, N10820, N5808, N2592, N1873);
or OR3 (N10830, N10824, N9971, N687);
or OR3 (N10831, N10828, N6154, N2746);
buf BUF1 (N10832, N10830);
nor NOR2 (N10833, N10812, N1448);
buf BUF1 (N10834, N10825);
and AND4 (N10835, N10821, N9241, N9430, N5591);
nand NAND3 (N10836, N10827, N6996, N5445);
and AND4 (N10837, N10836, N10138, N3724, N2203);
xor XOR2 (N10838, N10818, N3125);
xor XOR2 (N10839, N10829, N7442);
nor NOR3 (N10840, N10834, N3038, N527);
buf BUF1 (N10841, N10833);
not NOT1 (N10842, N10840);
xor XOR2 (N10843, N10841, N5204);
xor XOR2 (N10844, N10839, N5065);
buf BUF1 (N10845, N10835);
or OR4 (N10846, N10838, N3456, N672, N556);
nor NOR2 (N10847, N10826, N8736);
xor XOR2 (N10848, N10847, N1693);
nand NAND4 (N10849, N10844, N6916, N230, N3827);
and AND3 (N10850, N10813, N625, N7753);
nand NAND2 (N10851, N10837, N5525);
not NOT1 (N10852, N10851);
and AND3 (N10853, N10848, N9444, N9120);
nor NOR2 (N10854, N10852, N9032);
not NOT1 (N10855, N10842);
buf BUF1 (N10856, N10849);
not NOT1 (N10857, N10853);
nand NAND3 (N10858, N10831, N5808, N8569);
or OR3 (N10859, N10858, N78, N7848);
not NOT1 (N10860, N10843);
buf BUF1 (N10861, N10856);
not NOT1 (N10862, N10850);
buf BUF1 (N10863, N10854);
and AND4 (N10864, N10832, N5476, N6329, N8823);
xor XOR2 (N10865, N10857, N1741);
nand NAND4 (N10866, N10863, N4586, N1456, N790);
or OR3 (N10867, N10855, N1847, N3526);
or OR3 (N10868, N10860, N2017, N10182);
or OR3 (N10869, N10866, N9747, N7537);
xor XOR2 (N10870, N10862, N875);
buf BUF1 (N10871, N10870);
xor XOR2 (N10872, N10861, N2577);
xor XOR2 (N10873, N10869, N3620);
nor NOR4 (N10874, N10864, N139, N3073, N6845);
not NOT1 (N10875, N10845);
not NOT1 (N10876, N10846);
xor XOR2 (N10877, N10876, N3191);
nor NOR2 (N10878, N10867, N5575);
buf BUF1 (N10879, N10865);
xor XOR2 (N10880, N10871, N10267);
and AND2 (N10881, N10878, N8846);
nor NOR3 (N10882, N10875, N1050, N5674);
nand NAND3 (N10883, N10880, N2632, N3509);
xor XOR2 (N10884, N10877, N3090);
and AND2 (N10885, N10881, N7511);
or OR3 (N10886, N10874, N1112, N7286);
not NOT1 (N10887, N10884);
and AND2 (N10888, N10883, N2816);
nor NOR2 (N10889, N10872, N4576);
xor XOR2 (N10890, N10886, N5631);
nor NOR2 (N10891, N10882, N2467);
nand NAND2 (N10892, N10859, N6089);
nand NAND3 (N10893, N10885, N1464, N7195);
not NOT1 (N10894, N10879);
buf BUF1 (N10895, N10890);
not NOT1 (N10896, N10887);
nor NOR3 (N10897, N10894, N7811, N10419);
xor XOR2 (N10898, N10895, N6909);
nor NOR2 (N10899, N10873, N8386);
nand NAND3 (N10900, N10898, N8937, N1156);
buf BUF1 (N10901, N10891);
nor NOR3 (N10902, N10899, N10819, N3188);
or OR2 (N10903, N10888, N5489);
nor NOR2 (N10904, N10902, N3496);
not NOT1 (N10905, N10896);
or OR3 (N10906, N10892, N6154, N655);
or OR2 (N10907, N10897, N8701);
not NOT1 (N10908, N10893);
not NOT1 (N10909, N10900);
nand NAND4 (N10910, N10889, N2102, N7192, N2599);
buf BUF1 (N10911, N10909);
not NOT1 (N10912, N10903);
or OR2 (N10913, N10912, N3057);
nor NOR3 (N10914, N10906, N2301, N231);
nand NAND4 (N10915, N10914, N1616, N6974, N5072);
and AND3 (N10916, N10868, N8876, N10254);
not NOT1 (N10917, N10913);
nand NAND4 (N10918, N10910, N10550, N6889, N8960);
buf BUF1 (N10919, N10908);
buf BUF1 (N10920, N10907);
nand NAND2 (N10921, N10901, N3067);
nand NAND3 (N10922, N10920, N1924, N7921);
nand NAND3 (N10923, N10905, N3909, N10098);
not NOT1 (N10924, N10923);
nor NOR3 (N10925, N10922, N6252, N9048);
and AND4 (N10926, N10924, N6539, N1545, N5367);
or OR2 (N10927, N10904, N1322);
nand NAND3 (N10928, N10926, N433, N8222);
and AND2 (N10929, N10921, N6715);
not NOT1 (N10930, N10919);
not NOT1 (N10931, N10930);
xor XOR2 (N10932, N10917, N6514);
not NOT1 (N10933, N10918);
xor XOR2 (N10934, N10927, N3974);
buf BUF1 (N10935, N10925);
buf BUF1 (N10936, N10929);
nor NOR3 (N10937, N10915, N2287, N4642);
or OR2 (N10938, N10916, N5687);
xor XOR2 (N10939, N10936, N8935);
nor NOR4 (N10940, N10939, N9761, N5250, N218);
buf BUF1 (N10941, N10937);
nand NAND2 (N10942, N10935, N8423);
nand NAND4 (N10943, N10940, N1979, N6505, N7699);
not NOT1 (N10944, N10934);
nor NOR2 (N10945, N10911, N5633);
nand NAND4 (N10946, N10938, N10117, N1967, N9761);
buf BUF1 (N10947, N10944);
not NOT1 (N10948, N10943);
buf BUF1 (N10949, N10931);
and AND4 (N10950, N10941, N3686, N9382, N10475);
buf BUF1 (N10951, N10950);
buf BUF1 (N10952, N10948);
buf BUF1 (N10953, N10947);
or OR3 (N10954, N10945, N8765, N4124);
nand NAND2 (N10955, N10932, N2804);
and AND3 (N10956, N10953, N9830, N3506);
xor XOR2 (N10957, N10933, N8333);
nor NOR2 (N10958, N10949, N5345);
nor NOR4 (N10959, N10928, N8597, N4214, N9118);
or OR4 (N10960, N10957, N662, N4733, N2337);
not NOT1 (N10961, N10958);
buf BUF1 (N10962, N10955);
not NOT1 (N10963, N10956);
not NOT1 (N10964, N10952);
not NOT1 (N10965, N10946);
not NOT1 (N10966, N10954);
or OR3 (N10967, N10964, N7790, N10432);
and AND3 (N10968, N10966, N5806, N3526);
xor XOR2 (N10969, N10962, N10213);
buf BUF1 (N10970, N10961);
and AND4 (N10971, N10960, N10541, N488, N7628);
or OR4 (N10972, N10970, N590, N8474, N4469);
not NOT1 (N10973, N10942);
xor XOR2 (N10974, N10968, N2925);
xor XOR2 (N10975, N10967, N1272);
xor XOR2 (N10976, N10951, N4346);
or OR2 (N10977, N10971, N10117);
nor NOR4 (N10978, N10963, N7078, N2497, N2352);
xor XOR2 (N10979, N10977, N4750);
buf BUF1 (N10980, N10979);
buf BUF1 (N10981, N10975);
not NOT1 (N10982, N10976);
nand NAND3 (N10983, N10965, N6970, N5747);
buf BUF1 (N10984, N10969);
or OR2 (N10985, N10978, N10893);
nand NAND2 (N10986, N10985, N2516);
and AND2 (N10987, N10981, N9169);
xor XOR2 (N10988, N10959, N5218);
not NOT1 (N10989, N10984);
nand NAND2 (N10990, N10987, N10703);
or OR2 (N10991, N10988, N9707);
or OR3 (N10992, N10973, N3317, N9962);
or OR4 (N10993, N10974, N9805, N1353, N4061);
nand NAND4 (N10994, N10982, N1373, N6414, N9699);
and AND3 (N10995, N10992, N5972, N7946);
not NOT1 (N10996, N10993);
or OR3 (N10997, N10991, N6033, N922);
not NOT1 (N10998, N10980);
xor XOR2 (N10999, N10990, N10254);
nand NAND4 (N11000, N10995, N3730, N5767, N2900);
nand NAND2 (N11001, N10994, N4624);
buf BUF1 (N11002, N10983);
and AND3 (N11003, N10998, N945, N1946);
xor XOR2 (N11004, N11002, N3311);
or OR3 (N11005, N10999, N5623, N9932);
xor XOR2 (N11006, N11003, N7615);
nor NOR2 (N11007, N10986, N2530);
nand NAND2 (N11008, N10997, N3801);
nand NAND3 (N11009, N10972, N5037, N4834);
and AND3 (N11010, N11000, N4444, N3050);
nor NOR4 (N11011, N10996, N2259, N4485, N2887);
or OR4 (N11012, N10989, N4131, N10276, N3072);
xor XOR2 (N11013, N11010, N4909);
nand NAND4 (N11014, N11001, N4928, N5279, N7474);
nand NAND4 (N11015, N11012, N10016, N1733, N2566);
nor NOR2 (N11016, N11013, N6039);
xor XOR2 (N11017, N11008, N3877);
nand NAND3 (N11018, N11005, N3483, N4186);
xor XOR2 (N11019, N11004, N8270);
and AND2 (N11020, N11016, N5017);
nand NAND3 (N11021, N11019, N3425, N5184);
or OR4 (N11022, N11018, N4106, N6128, N6776);
nand NAND3 (N11023, N11021, N3169, N4695);
nor NOR4 (N11024, N11015, N9347, N2857, N1805);
nor NOR3 (N11025, N11023, N5212, N6338);
buf BUF1 (N11026, N11009);
and AND3 (N11027, N11026, N7793, N10217);
or OR2 (N11028, N11006, N10501);
or OR2 (N11029, N11022, N1267);
and AND3 (N11030, N11017, N2219, N4181);
nand NAND3 (N11031, N11029, N9586, N4827);
not NOT1 (N11032, N11031);
nor NOR4 (N11033, N11024, N746, N7438, N4750);
or OR4 (N11034, N11028, N4281, N9334, N2690);
nand NAND4 (N11035, N11014, N6655, N8739, N4809);
or OR3 (N11036, N11025, N200, N4550);
or OR2 (N11037, N11030, N4022);
nand NAND3 (N11038, N11033, N3703, N6548);
nor NOR2 (N11039, N11034, N6327);
and AND4 (N11040, N11035, N8731, N6271, N6920);
nand NAND2 (N11041, N11036, N5697);
not NOT1 (N11042, N11020);
or OR2 (N11043, N11037, N9085);
nand NAND4 (N11044, N11032, N9059, N1761, N6906);
nor NOR3 (N11045, N11007, N2030, N23);
nor NOR2 (N11046, N11038, N7492);
nand NAND3 (N11047, N11027, N8547, N1572);
not NOT1 (N11048, N11042);
and AND2 (N11049, N11047, N7306);
or OR4 (N11050, N11045, N5882, N10227, N543);
xor XOR2 (N11051, N11046, N3828);
or OR3 (N11052, N11039, N1401, N9713);
xor XOR2 (N11053, N11049, N3491);
xor XOR2 (N11054, N11040, N9407);
nand NAND2 (N11055, N11051, N4437);
buf BUF1 (N11056, N11055);
nor NOR3 (N11057, N11056, N480, N5722);
nor NOR2 (N11058, N11050, N7576);
or OR4 (N11059, N11058, N9233, N5898, N5923);
nand NAND2 (N11060, N11011, N3301);
or OR3 (N11061, N11044, N10767, N3700);
xor XOR2 (N11062, N11052, N10024);
xor XOR2 (N11063, N11059, N9025);
and AND4 (N11064, N11041, N2864, N5873, N6375);
buf BUF1 (N11065, N11064);
buf BUF1 (N11066, N11060);
nor NOR4 (N11067, N11062, N7836, N8717, N5149);
and AND3 (N11068, N11063, N259, N10814);
nor NOR3 (N11069, N11067, N9453, N10858);
or OR3 (N11070, N11068, N4993, N6773);
xor XOR2 (N11071, N11069, N6362);
xor XOR2 (N11072, N11071, N787);
not NOT1 (N11073, N11070);
buf BUF1 (N11074, N11065);
nor NOR3 (N11075, N11054, N1366, N5727);
and AND2 (N11076, N11066, N2437);
or OR4 (N11077, N11075, N1146, N4500, N1753);
not NOT1 (N11078, N11053);
xor XOR2 (N11079, N11043, N3503);
nor NOR3 (N11080, N11078, N3668, N4623);
not NOT1 (N11081, N11073);
and AND2 (N11082, N11079, N1121);
nor NOR2 (N11083, N11072, N5465);
or OR4 (N11084, N11048, N4610, N390, N6269);
and AND4 (N11085, N11084, N709, N9312, N9670);
xor XOR2 (N11086, N11082, N9690);
nand NAND3 (N11087, N11086, N6850, N8910);
not NOT1 (N11088, N11081);
not NOT1 (N11089, N11080);
not NOT1 (N11090, N11057);
nand NAND4 (N11091, N11089, N2048, N4273, N7421);
buf BUF1 (N11092, N11088);
buf BUF1 (N11093, N11074);
xor XOR2 (N11094, N11076, N7277);
or OR2 (N11095, N11077, N2001);
and AND3 (N11096, N11085, N7107, N6818);
nor NOR2 (N11097, N11095, N6915);
nor NOR2 (N11098, N11096, N3581);
nand NAND3 (N11099, N11092, N4376, N2282);
xor XOR2 (N11100, N11083, N6761);
xor XOR2 (N11101, N11098, N4);
nand NAND2 (N11102, N11091, N3765);
nor NOR3 (N11103, N11101, N2092, N7316);
or OR4 (N11104, N11087, N9077, N6353, N7486);
nand NAND3 (N11105, N11102, N39, N4240);
buf BUF1 (N11106, N11103);
and AND2 (N11107, N11100, N3008);
nand NAND4 (N11108, N11097, N3571, N7677, N3263);
or OR3 (N11109, N11108, N6722, N8350);
buf BUF1 (N11110, N11061);
nor NOR4 (N11111, N11107, N10189, N6740, N7749);
and AND4 (N11112, N11105, N9033, N10105, N4747);
nand NAND4 (N11113, N11090, N9700, N3636, N5035);
and AND2 (N11114, N11111, N999);
nor NOR4 (N11115, N11112, N3581, N2059, N2065);
nand NAND2 (N11116, N11106, N5339);
nor NOR3 (N11117, N11116, N1394, N777);
buf BUF1 (N11118, N11114);
not NOT1 (N11119, N11109);
nand NAND2 (N11120, N11104, N4745);
or OR3 (N11121, N11118, N6223, N7659);
and AND3 (N11122, N11120, N10702, N988);
nor NOR3 (N11123, N11093, N5782, N2407);
nand NAND4 (N11124, N11121, N1692, N6877, N7294);
xor XOR2 (N11125, N11119, N10614);
and AND3 (N11126, N11117, N9467, N10616);
and AND4 (N11127, N11123, N6532, N10120, N3922);
xor XOR2 (N11128, N11124, N8797);
nor NOR3 (N11129, N11126, N3900, N11010);
not NOT1 (N11130, N11122);
not NOT1 (N11131, N11094);
or OR3 (N11132, N11129, N5338, N7005);
and AND2 (N11133, N11113, N9610);
nand NAND2 (N11134, N11132, N1596);
and AND4 (N11135, N11131, N2341, N318, N10894);
not NOT1 (N11136, N11128);
and AND3 (N11137, N11110, N7854, N6911);
nand NAND2 (N11138, N11127, N5604);
nand NAND3 (N11139, N11115, N5368, N521);
xor XOR2 (N11140, N11099, N10783);
or OR4 (N11141, N11136, N4059, N6009, N1549);
xor XOR2 (N11142, N11140, N2576);
xor XOR2 (N11143, N11138, N7451);
and AND4 (N11144, N11125, N10502, N5132, N3623);
and AND4 (N11145, N11134, N2356, N8466, N3335);
and AND2 (N11146, N11142, N3877);
not NOT1 (N11147, N11144);
nor NOR2 (N11148, N11146, N9831);
nor NOR4 (N11149, N11133, N8428, N10237, N3578);
or OR2 (N11150, N11130, N9947);
xor XOR2 (N11151, N11137, N3008);
or OR4 (N11152, N11149, N7994, N7786, N3701);
xor XOR2 (N11153, N11147, N158);
xor XOR2 (N11154, N11143, N1547);
and AND4 (N11155, N11135, N3202, N2429, N10731);
nor NOR2 (N11156, N11151, N8290);
nor NOR2 (N11157, N11139, N9308);
nand NAND3 (N11158, N11145, N6821, N874);
nand NAND2 (N11159, N11156, N6361);
nor NOR4 (N11160, N11148, N10910, N1169, N4812);
not NOT1 (N11161, N11158);
nand NAND3 (N11162, N11153, N5196, N3376);
or OR2 (N11163, N11150, N10800);
buf BUF1 (N11164, N11157);
and AND3 (N11165, N11154, N6469, N9662);
nor NOR2 (N11166, N11159, N3627);
not NOT1 (N11167, N11152);
not NOT1 (N11168, N11166);
nor NOR2 (N11169, N11163, N3302);
xor XOR2 (N11170, N11168, N1387);
buf BUF1 (N11171, N11167);
nand NAND4 (N11172, N11160, N6301, N6434, N3674);
nor NOR4 (N11173, N11141, N5814, N5974, N6327);
not NOT1 (N11174, N11169);
and AND3 (N11175, N11161, N8623, N7990);
or OR3 (N11176, N11162, N5065, N1946);
buf BUF1 (N11177, N11174);
xor XOR2 (N11178, N11173, N9082);
and AND3 (N11179, N11175, N5176, N5705);
and AND3 (N11180, N11176, N9021, N327);
nand NAND3 (N11181, N11155, N11150, N6804);
or OR2 (N11182, N11178, N2222);
and AND3 (N11183, N11165, N10597, N4107);
or OR2 (N11184, N11182, N2260);
buf BUF1 (N11185, N11184);
and AND2 (N11186, N11172, N5039);
nor NOR2 (N11187, N11177, N9502);
buf BUF1 (N11188, N11186);
xor XOR2 (N11189, N11185, N6258);
buf BUF1 (N11190, N11181);
and AND4 (N11191, N11187, N10674, N77, N5139);
or OR3 (N11192, N11191, N1798, N676);
and AND3 (N11193, N11192, N3953, N4640);
nor NOR4 (N11194, N11179, N8517, N53, N10997);
or OR3 (N11195, N11180, N5606, N1270);
and AND3 (N11196, N11188, N7660, N10924);
buf BUF1 (N11197, N11183);
and AND4 (N11198, N11171, N3056, N6213, N7125);
buf BUF1 (N11199, N11198);
and AND4 (N11200, N11193, N6588, N7534, N4404);
buf BUF1 (N11201, N11164);
not NOT1 (N11202, N11194);
buf BUF1 (N11203, N11197);
not NOT1 (N11204, N11201);
nand NAND3 (N11205, N11196, N6445, N6431);
xor XOR2 (N11206, N11199, N6019);
nand NAND2 (N11207, N11204, N2993);
xor XOR2 (N11208, N11200, N2045);
buf BUF1 (N11209, N11189);
buf BUF1 (N11210, N11203);
buf BUF1 (N11211, N11208);
nor NOR3 (N11212, N11207, N2900, N5094);
and AND2 (N11213, N11212, N2402);
or OR2 (N11214, N11213, N7401);
xor XOR2 (N11215, N11205, N9453);
nand NAND3 (N11216, N11209, N5125, N668);
xor XOR2 (N11217, N11170, N3908);
buf BUF1 (N11218, N11202);
buf BUF1 (N11219, N11190);
or OR4 (N11220, N11211, N8013, N1471, N4427);
or OR4 (N11221, N11206, N134, N2423, N4292);
and AND3 (N11222, N11195, N2882, N10755);
not NOT1 (N11223, N11214);
nand NAND3 (N11224, N11221, N5649, N11208);
not NOT1 (N11225, N11218);
buf BUF1 (N11226, N11219);
nor NOR2 (N11227, N11217, N1351);
nand NAND4 (N11228, N11225, N4256, N1585, N4809);
nor NOR2 (N11229, N11215, N8593);
xor XOR2 (N11230, N11229, N2734);
not NOT1 (N11231, N11224);
xor XOR2 (N11232, N11222, N8503);
nor NOR2 (N11233, N11216, N3294);
nor NOR4 (N11234, N11226, N8266, N10060, N1162);
or OR4 (N11235, N11228, N676, N10770, N10164);
nand NAND3 (N11236, N11233, N10708, N9099);
or OR2 (N11237, N11231, N4308);
not NOT1 (N11238, N11236);
xor XOR2 (N11239, N11223, N10983);
xor XOR2 (N11240, N11235, N322);
nand NAND3 (N11241, N11240, N620, N1473);
or OR2 (N11242, N11239, N1272);
or OR2 (N11243, N11242, N1506);
and AND2 (N11244, N11232, N3565);
or OR3 (N11245, N11220, N4241, N5935);
and AND4 (N11246, N11230, N9232, N9537, N1609);
or OR4 (N11247, N11234, N10516, N4703, N1234);
xor XOR2 (N11248, N11247, N753);
xor XOR2 (N11249, N11238, N3307);
and AND3 (N11250, N11210, N3456, N3789);
buf BUF1 (N11251, N11243);
nor NOR2 (N11252, N11249, N6762);
not NOT1 (N11253, N11237);
nor NOR4 (N11254, N11241, N3594, N5676, N9811);
xor XOR2 (N11255, N11244, N9517);
xor XOR2 (N11256, N11227, N5213);
nor NOR4 (N11257, N11253, N2136, N5662, N9995);
and AND2 (N11258, N11246, N11212);
or OR4 (N11259, N11252, N7537, N1652, N7998);
not NOT1 (N11260, N11254);
and AND2 (N11261, N11256, N1638);
xor XOR2 (N11262, N11245, N10741);
xor XOR2 (N11263, N11262, N3093);
nor NOR4 (N11264, N11259, N4320, N8105, N9736);
or OR4 (N11265, N11258, N5839, N10188, N6637);
xor XOR2 (N11266, N11260, N9589);
xor XOR2 (N11267, N11261, N10372);
buf BUF1 (N11268, N11267);
xor XOR2 (N11269, N11257, N10503);
and AND3 (N11270, N11268, N10746, N8175);
nand NAND2 (N11271, N11265, N5093);
not NOT1 (N11272, N11263);
nor NOR3 (N11273, N11264, N5875, N8725);
xor XOR2 (N11274, N11250, N2839);
nor NOR2 (N11275, N11255, N10915);
nor NOR4 (N11276, N11266, N3140, N7165, N4684);
or OR3 (N11277, N11271, N984, N9753);
buf BUF1 (N11278, N11270);
or OR4 (N11279, N11278, N8239, N9841, N2121);
not NOT1 (N11280, N11277);
buf BUF1 (N11281, N11269);
or OR4 (N11282, N11248, N10806, N1866, N4439);
nand NAND4 (N11283, N11275, N1338, N10234, N7256);
or OR3 (N11284, N11274, N7249, N4335);
nor NOR4 (N11285, N11272, N2696, N2773, N10008);
or OR3 (N11286, N11281, N3444, N8412);
and AND4 (N11287, N11251, N1985, N6955, N3011);
nor NOR2 (N11288, N11287, N4102);
xor XOR2 (N11289, N11288, N4760);
buf BUF1 (N11290, N11280);
nand NAND3 (N11291, N11273, N6971, N3517);
or OR3 (N11292, N11290, N6688, N9545);
or OR4 (N11293, N11289, N7745, N11139, N7557);
nand NAND3 (N11294, N11283, N11201, N3481);
or OR3 (N11295, N11276, N4791, N6732);
nor NOR3 (N11296, N11282, N8752, N9500);
xor XOR2 (N11297, N11284, N5954);
or OR4 (N11298, N11295, N7232, N9451, N749);
nand NAND3 (N11299, N11298, N300, N5088);
not NOT1 (N11300, N11296);
nand NAND3 (N11301, N11279, N9535, N7030);
nor NOR4 (N11302, N11301, N3817, N6225, N5298);
xor XOR2 (N11303, N11294, N10990);
not NOT1 (N11304, N11285);
xor XOR2 (N11305, N11304, N8923);
not NOT1 (N11306, N11291);
buf BUF1 (N11307, N11300);
nor NOR2 (N11308, N11286, N7567);
nand NAND3 (N11309, N11302, N8095, N5628);
xor XOR2 (N11310, N11306, N4713);
nor NOR4 (N11311, N11305, N6801, N545, N3050);
not NOT1 (N11312, N11292);
nor NOR2 (N11313, N11311, N6939);
nand NAND3 (N11314, N11310, N8428, N9747);
buf BUF1 (N11315, N11313);
and AND3 (N11316, N11307, N1862, N8922);
nor NOR2 (N11317, N11316, N4049);
not NOT1 (N11318, N11297);
not NOT1 (N11319, N11303);
xor XOR2 (N11320, N11299, N7106);
buf BUF1 (N11321, N11317);
not NOT1 (N11322, N11314);
nor NOR4 (N11323, N11322, N9598, N5178, N6478);
or OR3 (N11324, N11315, N8306, N10038);
xor XOR2 (N11325, N11309, N5027);
nor NOR4 (N11326, N11308, N1845, N10706, N6154);
not NOT1 (N11327, N11323);
buf BUF1 (N11328, N11319);
nand NAND2 (N11329, N11328, N8611);
xor XOR2 (N11330, N11312, N9303);
buf BUF1 (N11331, N11321);
nand NAND2 (N11332, N11324, N6459);
or OR3 (N11333, N11325, N1836, N3922);
nor NOR2 (N11334, N11333, N655);
nand NAND4 (N11335, N11326, N2657, N716, N9705);
and AND3 (N11336, N11332, N10110, N10838);
buf BUF1 (N11337, N11330);
xor XOR2 (N11338, N11334, N7245);
and AND4 (N11339, N11331, N2307, N7327, N844);
or OR4 (N11340, N11339, N6892, N7381, N6456);
not NOT1 (N11341, N11337);
xor XOR2 (N11342, N11327, N6986);
nand NAND3 (N11343, N11341, N3357, N10902);
buf BUF1 (N11344, N11340);
or OR2 (N11345, N11343, N9371);
xor XOR2 (N11346, N11329, N4905);
xor XOR2 (N11347, N11346, N1228);
nor NOR3 (N11348, N11342, N1852, N7487);
or OR2 (N11349, N11336, N11216);
and AND4 (N11350, N11344, N11035, N1495, N9948);
or OR2 (N11351, N11345, N360);
nand NAND3 (N11352, N11293, N9646, N7462);
buf BUF1 (N11353, N11338);
not NOT1 (N11354, N11350);
xor XOR2 (N11355, N11318, N3114);
or OR2 (N11356, N11352, N3237);
xor XOR2 (N11357, N11351, N6260);
and AND3 (N11358, N11348, N3411, N5702);
or OR2 (N11359, N11320, N4717);
not NOT1 (N11360, N11358);
not NOT1 (N11361, N11356);
buf BUF1 (N11362, N11355);
and AND3 (N11363, N11354, N2192, N11014);
xor XOR2 (N11364, N11349, N7093);
nand NAND3 (N11365, N11364, N10049, N10650);
nand NAND3 (N11366, N11360, N2520, N2948);
and AND4 (N11367, N11365, N107, N4294, N3399);
xor XOR2 (N11368, N11366, N7670);
or OR3 (N11369, N11362, N8909, N10645);
or OR3 (N11370, N11353, N10875, N3449);
not NOT1 (N11371, N11361);
xor XOR2 (N11372, N11357, N8419);
or OR4 (N11373, N11367, N10080, N9572, N6053);
or OR2 (N11374, N11372, N5691);
nor NOR3 (N11375, N11373, N3390, N10863);
nand NAND3 (N11376, N11371, N2413, N10106);
nor NOR3 (N11377, N11370, N7214, N8248);
nor NOR3 (N11378, N11374, N6469, N5340);
nand NAND2 (N11379, N11376, N2969);
buf BUF1 (N11380, N11368);
nor NOR2 (N11381, N11380, N2584);
not NOT1 (N11382, N11381);
not NOT1 (N11383, N11369);
xor XOR2 (N11384, N11359, N11289);
or OR2 (N11385, N11335, N4428);
nand NAND3 (N11386, N11375, N11228, N1029);
or OR4 (N11387, N11363, N5407, N9041, N11028);
not NOT1 (N11388, N11378);
xor XOR2 (N11389, N11384, N5413);
or OR4 (N11390, N11388, N5050, N4325, N8343);
xor XOR2 (N11391, N11389, N694);
and AND2 (N11392, N11379, N453);
nand NAND3 (N11393, N11383, N8111, N5527);
and AND4 (N11394, N11385, N1534, N3044, N4031);
or OR2 (N11395, N11386, N1183);
xor XOR2 (N11396, N11347, N4376);
xor XOR2 (N11397, N11392, N9657);
xor XOR2 (N11398, N11390, N8955);
buf BUF1 (N11399, N11398);
buf BUF1 (N11400, N11377);
or OR4 (N11401, N11396, N9969, N5379, N2038);
xor XOR2 (N11402, N11397, N7326);
nand NAND4 (N11403, N11391, N257, N5163, N4002);
xor XOR2 (N11404, N11394, N2581);
not NOT1 (N11405, N11395);
nand NAND4 (N11406, N11382, N10098, N7542, N9421);
xor XOR2 (N11407, N11401, N2567);
nand NAND4 (N11408, N11393, N8161, N7444, N1518);
and AND2 (N11409, N11400, N3140);
buf BUF1 (N11410, N11402);
nor NOR4 (N11411, N11408, N277, N5969, N4669);
xor XOR2 (N11412, N11387, N6194);
and AND4 (N11413, N11403, N10527, N579, N1450);
xor XOR2 (N11414, N11406, N5342);
or OR2 (N11415, N11410, N10887);
or OR2 (N11416, N11399, N5018);
nor NOR2 (N11417, N11416, N10149);
nand NAND4 (N11418, N11415, N8132, N3420, N6399);
or OR4 (N11419, N11409, N5917, N4302, N2829);
and AND4 (N11420, N11414, N9596, N2476, N10551);
or OR2 (N11421, N11417, N3085);
nand NAND2 (N11422, N11419, N546);
xor XOR2 (N11423, N11421, N9542);
not NOT1 (N11424, N11423);
nand NAND4 (N11425, N11420, N5660, N4379, N6168);
and AND2 (N11426, N11404, N1694);
and AND2 (N11427, N11405, N4546);
or OR4 (N11428, N11424, N5416, N9280, N10895);
nor NOR3 (N11429, N11426, N8596, N7941);
nand NAND4 (N11430, N11429, N9052, N2388, N3906);
xor XOR2 (N11431, N11428, N4899);
or OR4 (N11432, N11413, N7436, N3754, N9979);
buf BUF1 (N11433, N11418);
xor XOR2 (N11434, N11425, N1608);
nor NOR4 (N11435, N11433, N7492, N5992, N569);
buf BUF1 (N11436, N11431);
not NOT1 (N11437, N11422);
nand NAND4 (N11438, N11434, N653, N553, N7223);
not NOT1 (N11439, N11407);
xor XOR2 (N11440, N11438, N3436);
not NOT1 (N11441, N11432);
nor NOR2 (N11442, N11441, N9313);
and AND4 (N11443, N11412, N3998, N3869, N7393);
not NOT1 (N11444, N11436);
and AND3 (N11445, N11440, N9354, N5617);
nand NAND2 (N11446, N11445, N7445);
nand NAND4 (N11447, N11443, N8495, N3333, N10811);
xor XOR2 (N11448, N11430, N3417);
buf BUF1 (N11449, N11427);
nand NAND4 (N11450, N11435, N5870, N10408, N5981);
nor NOR4 (N11451, N11442, N10635, N8643, N2290);
nand NAND4 (N11452, N11450, N6881, N5166, N847);
xor XOR2 (N11453, N11437, N8860);
nand NAND2 (N11454, N11446, N7762);
not NOT1 (N11455, N11447);
buf BUF1 (N11456, N11449);
or OR2 (N11457, N11456, N10047);
or OR2 (N11458, N11411, N425);
and AND4 (N11459, N11454, N3555, N7850, N1878);
not NOT1 (N11460, N11451);
xor XOR2 (N11461, N11458, N11080);
or OR2 (N11462, N11452, N3411);
not NOT1 (N11463, N11455);
or OR4 (N11464, N11459, N3355, N7937, N2250);
nor NOR2 (N11465, N11463, N3597);
buf BUF1 (N11466, N11439);
buf BUF1 (N11467, N11464);
xor XOR2 (N11468, N11444, N3950);
or OR2 (N11469, N11462, N11268);
not NOT1 (N11470, N11453);
xor XOR2 (N11471, N11466, N3964);
nor NOR3 (N11472, N11448, N3067, N684);
and AND2 (N11473, N11460, N6231);
buf BUF1 (N11474, N11457);
buf BUF1 (N11475, N11472);
not NOT1 (N11476, N11474);
nor NOR3 (N11477, N11469, N1749, N9778);
xor XOR2 (N11478, N11465, N3099);
not NOT1 (N11479, N11461);
not NOT1 (N11480, N11471);
nand NAND2 (N11481, N11479, N9298);
nand NAND2 (N11482, N11477, N10563);
and AND3 (N11483, N11476, N852, N7180);
nor NOR3 (N11484, N11480, N2985, N6023);
nor NOR4 (N11485, N11483, N6127, N7655, N7289);
buf BUF1 (N11486, N11485);
buf BUF1 (N11487, N11478);
and AND4 (N11488, N11484, N3787, N2651, N8413);
and AND3 (N11489, N11475, N10843, N10151);
xor XOR2 (N11490, N11488, N7580);
nand NAND4 (N11491, N11490, N3924, N7474, N11121);
or OR4 (N11492, N11489, N4036, N10694, N4241);
nor NOR3 (N11493, N11482, N9300, N7962);
or OR4 (N11494, N11487, N8112, N2556, N4266);
and AND3 (N11495, N11491, N6779, N8546);
nor NOR4 (N11496, N11493, N8481, N2825, N424);
xor XOR2 (N11497, N11473, N9319);
xor XOR2 (N11498, N11481, N7199);
or OR3 (N11499, N11467, N7237, N3133);
nor NOR4 (N11500, N11494, N7679, N6723, N3809);
nor NOR3 (N11501, N11492, N1228, N8346);
or OR2 (N11502, N11468, N11049);
and AND3 (N11503, N11486, N9582, N6053);
buf BUF1 (N11504, N11498);
buf BUF1 (N11505, N11504);
xor XOR2 (N11506, N11502, N8937);
or OR4 (N11507, N11499, N6548, N11026, N7094);
nor NOR4 (N11508, N11507, N667, N7210, N3308);
buf BUF1 (N11509, N11470);
xor XOR2 (N11510, N11506, N2846);
not NOT1 (N11511, N11510);
or OR2 (N11512, N11497, N1945);
nor NOR2 (N11513, N11500, N9451);
or OR4 (N11514, N11505, N10178, N7593, N6450);
nand NAND2 (N11515, N11508, N2097);
and AND2 (N11516, N11515, N2413);
nor NOR3 (N11517, N11503, N10354, N11269);
nor NOR3 (N11518, N11513, N6515, N10024);
xor XOR2 (N11519, N11518, N3847);
not NOT1 (N11520, N11511);
nand NAND4 (N11521, N11512, N1697, N9428, N100);
or OR3 (N11522, N11496, N2240, N3358);
and AND3 (N11523, N11501, N11494, N9698);
or OR2 (N11524, N11520, N1464);
not NOT1 (N11525, N11524);
buf BUF1 (N11526, N11517);
and AND3 (N11527, N11521, N12, N7249);
or OR3 (N11528, N11514, N6613, N316);
xor XOR2 (N11529, N11519, N4240);
buf BUF1 (N11530, N11528);
and AND2 (N11531, N11526, N8775);
or OR4 (N11532, N11509, N5680, N5433, N545);
and AND2 (N11533, N11525, N1228);
not NOT1 (N11534, N11522);
xor XOR2 (N11535, N11527, N10384);
not NOT1 (N11536, N11533);
not NOT1 (N11537, N11536);
nand NAND3 (N11538, N11534, N2923, N10158);
nand NAND3 (N11539, N11538, N7191, N4415);
nor NOR2 (N11540, N11539, N1926);
xor XOR2 (N11541, N11529, N7074);
and AND2 (N11542, N11535, N2183);
xor XOR2 (N11543, N11495, N6939);
buf BUF1 (N11544, N11516);
not NOT1 (N11545, N11544);
buf BUF1 (N11546, N11541);
xor XOR2 (N11547, N11530, N543);
xor XOR2 (N11548, N11523, N5289);
nand NAND3 (N11549, N11542, N4148, N9409);
not NOT1 (N11550, N11546);
not NOT1 (N11551, N11548);
xor XOR2 (N11552, N11531, N5435);
and AND3 (N11553, N11532, N4120, N8497);
or OR4 (N11554, N11543, N9708, N7688, N11359);
xor XOR2 (N11555, N11547, N1039);
and AND2 (N11556, N11554, N957);
nor NOR3 (N11557, N11540, N7027, N10072);
nor NOR3 (N11558, N11552, N8318, N5344);
or OR2 (N11559, N11558, N6012);
or OR4 (N11560, N11559, N2359, N8315, N10732);
buf BUF1 (N11561, N11551);
or OR4 (N11562, N11557, N975, N1510, N10921);
buf BUF1 (N11563, N11560);
or OR2 (N11564, N11563, N7625);
not NOT1 (N11565, N11564);
nand NAND2 (N11566, N11537, N95);
or OR3 (N11567, N11566, N8927, N683);
and AND4 (N11568, N11561, N3959, N3649, N2456);
and AND3 (N11569, N11553, N8134, N2504);
nor NOR2 (N11570, N11568, N9006);
or OR3 (N11571, N11569, N2278, N5317);
xor XOR2 (N11572, N11555, N8918);
and AND4 (N11573, N11565, N9152, N9648, N6771);
and AND3 (N11574, N11562, N7447, N1436);
nand NAND2 (N11575, N11573, N4106);
nor NOR3 (N11576, N11571, N10551, N7803);
xor XOR2 (N11577, N11570, N2920);
xor XOR2 (N11578, N11549, N9598);
xor XOR2 (N11579, N11556, N4184);
or OR2 (N11580, N11576, N2067);
nor NOR2 (N11581, N11579, N10976);
or OR4 (N11582, N11572, N4332, N11254, N1623);
nand NAND4 (N11583, N11581, N10094, N6841, N9832);
not NOT1 (N11584, N11580);
nor NOR3 (N11585, N11574, N11581, N10833);
and AND3 (N11586, N11578, N5549, N8778);
or OR4 (N11587, N11583, N6313, N1820, N8057);
or OR3 (N11588, N11586, N11513, N4216);
xor XOR2 (N11589, N11567, N8939);
and AND4 (N11590, N11575, N10965, N8900, N555);
nor NOR2 (N11591, N11550, N8450);
not NOT1 (N11592, N11584);
not NOT1 (N11593, N11588);
nor NOR4 (N11594, N11591, N3241, N1684, N8713);
nor NOR3 (N11595, N11593, N5261, N9707);
buf BUF1 (N11596, N11589);
nand NAND4 (N11597, N11545, N5333, N8270, N7684);
nor NOR2 (N11598, N11587, N4365);
nand NAND4 (N11599, N11577, N4276, N8617, N8850);
not NOT1 (N11600, N11590);
not NOT1 (N11601, N11596);
xor XOR2 (N11602, N11598, N4215);
nand NAND4 (N11603, N11602, N10040, N8458, N7357);
or OR2 (N11604, N11599, N9777);
nor NOR3 (N11605, N11603, N4197, N2295);
and AND3 (N11606, N11595, N9039, N7951);
nor NOR4 (N11607, N11592, N9814, N2265, N6511);
and AND2 (N11608, N11582, N2725);
and AND2 (N11609, N11601, N3169);
xor XOR2 (N11610, N11609, N405);
not NOT1 (N11611, N11610);
or OR4 (N11612, N11585, N8492, N4451, N1430);
and AND3 (N11613, N11604, N7100, N9595);
xor XOR2 (N11614, N11600, N4666);
or OR3 (N11615, N11611, N9771, N10327);
not NOT1 (N11616, N11613);
not NOT1 (N11617, N11607);
not NOT1 (N11618, N11612);
xor XOR2 (N11619, N11606, N2565);
xor XOR2 (N11620, N11597, N10351);
nor NOR3 (N11621, N11618, N9634, N8215);
or OR3 (N11622, N11615, N5467, N7415);
nor NOR4 (N11623, N11614, N4034, N442, N5984);
not NOT1 (N11624, N11617);
nand NAND4 (N11625, N11620, N921, N2316, N3416);
xor XOR2 (N11626, N11621, N5986);
nor NOR2 (N11627, N11605, N8349);
buf BUF1 (N11628, N11625);
buf BUF1 (N11629, N11619);
or OR3 (N11630, N11627, N3563, N2933);
xor XOR2 (N11631, N11624, N5848);
buf BUF1 (N11632, N11622);
nor NOR2 (N11633, N11623, N10082);
nand NAND4 (N11634, N11628, N9336, N5420, N6085);
and AND3 (N11635, N11629, N1492, N5872);
not NOT1 (N11636, N11594);
buf BUF1 (N11637, N11633);
nor NOR3 (N11638, N11634, N4268, N10051);
buf BUF1 (N11639, N11636);
xor XOR2 (N11640, N11608, N7887);
nand NAND4 (N11641, N11635, N6180, N6990, N4034);
not NOT1 (N11642, N11632);
or OR4 (N11643, N11626, N3448, N4294, N5106);
nand NAND4 (N11644, N11638, N2888, N4714, N9998);
nor NOR3 (N11645, N11637, N6166, N5824);
and AND3 (N11646, N11631, N536, N382);
and AND4 (N11647, N11630, N11281, N6356, N2292);
buf BUF1 (N11648, N11641);
nand NAND3 (N11649, N11648, N6422, N7103);
and AND3 (N11650, N11642, N9506, N1962);
not NOT1 (N11651, N11646);
or OR4 (N11652, N11650, N9574, N4218, N753);
buf BUF1 (N11653, N11643);
nand NAND2 (N11654, N11653, N9230);
nor NOR2 (N11655, N11640, N1373);
buf BUF1 (N11656, N11649);
or OR4 (N11657, N11655, N9746, N10077, N428);
not NOT1 (N11658, N11645);
not NOT1 (N11659, N11639);
not NOT1 (N11660, N11644);
xor XOR2 (N11661, N11659, N99);
nand NAND4 (N11662, N11651, N5934, N4853, N2060);
or OR2 (N11663, N11657, N5270);
nor NOR2 (N11664, N11658, N3436);
and AND3 (N11665, N11647, N4471, N9947);
not NOT1 (N11666, N11616);
and AND3 (N11667, N11661, N745, N11635);
nand NAND4 (N11668, N11662, N6996, N5250, N5459);
xor XOR2 (N11669, N11656, N7641);
nor NOR3 (N11670, N11652, N5344, N8333);
xor XOR2 (N11671, N11668, N9408);
buf BUF1 (N11672, N11654);
xor XOR2 (N11673, N11666, N4709);
nor NOR2 (N11674, N11669, N618);
nor NOR2 (N11675, N11665, N280);
nand NAND4 (N11676, N11670, N10226, N9627, N1744);
nand NAND2 (N11677, N11676, N2276);
and AND2 (N11678, N11667, N6889);
or OR4 (N11679, N11678, N8443, N260, N10420);
and AND4 (N11680, N11674, N1105, N3610, N5957);
and AND3 (N11681, N11672, N10701, N10183);
not NOT1 (N11682, N11664);
not NOT1 (N11683, N11680);
or OR2 (N11684, N11675, N3807);
and AND4 (N11685, N11671, N10111, N5738, N10099);
buf BUF1 (N11686, N11684);
or OR4 (N11687, N11677, N9431, N10902, N4111);
xor XOR2 (N11688, N11660, N3434);
xor XOR2 (N11689, N11683, N233);
xor XOR2 (N11690, N11663, N11098);
buf BUF1 (N11691, N11673);
xor XOR2 (N11692, N11690, N6381);
or OR2 (N11693, N11689, N11444);
not NOT1 (N11694, N11686);
not NOT1 (N11695, N11679);
not NOT1 (N11696, N11694);
nor NOR3 (N11697, N11681, N6938, N549);
and AND4 (N11698, N11682, N5034, N5205, N2357);
nor NOR2 (N11699, N11691, N3672);
and AND3 (N11700, N11685, N9622, N7769);
not NOT1 (N11701, N11688);
and AND3 (N11702, N11696, N3608, N11312);
and AND4 (N11703, N11700, N5778, N5109, N4978);
or OR2 (N11704, N11695, N101);
and AND3 (N11705, N11704, N2872, N7159);
xor XOR2 (N11706, N11705, N5696);
nor NOR2 (N11707, N11687, N11496);
not NOT1 (N11708, N11699);
xor XOR2 (N11709, N11698, N5839);
or OR2 (N11710, N11692, N8474);
or OR4 (N11711, N11707, N1096, N5402, N10753);
not NOT1 (N11712, N11711);
buf BUF1 (N11713, N11693);
or OR4 (N11714, N11709, N4173, N1832, N4148);
and AND3 (N11715, N11706, N61, N11521);
nand NAND2 (N11716, N11713, N7353);
nor NOR3 (N11717, N11697, N3240, N10691);
not NOT1 (N11718, N11702);
nand NAND4 (N11719, N11701, N527, N6535, N10742);
nor NOR2 (N11720, N11718, N11082);
nor NOR4 (N11721, N11708, N353, N9686, N7107);
or OR4 (N11722, N11714, N617, N4377, N5800);
nor NOR4 (N11723, N11716, N9750, N8764, N8990);
and AND4 (N11724, N11717, N1297, N6929, N3148);
xor XOR2 (N11725, N11724, N4222);
xor XOR2 (N11726, N11725, N3455);
buf BUF1 (N11727, N11710);
nand NAND3 (N11728, N11720, N4191, N2396);
or OR2 (N11729, N11715, N1327);
xor XOR2 (N11730, N11729, N3712);
nor NOR2 (N11731, N11721, N5554);
nand NAND3 (N11732, N11730, N6897, N7839);
buf BUF1 (N11733, N11719);
nand NAND4 (N11734, N11733, N4305, N7254, N1996);
not NOT1 (N11735, N11734);
nor NOR3 (N11736, N11735, N69, N7430);
not NOT1 (N11737, N11727);
xor XOR2 (N11738, N11723, N8157);
not NOT1 (N11739, N11731);
nor NOR2 (N11740, N11739, N1492);
nor NOR3 (N11741, N11736, N5271, N8164);
nand NAND4 (N11742, N11740, N5794, N8372, N9056);
not NOT1 (N11743, N11712);
not NOT1 (N11744, N11743);
or OR3 (N11745, N11742, N6400, N6238);
buf BUF1 (N11746, N11722);
or OR3 (N11747, N11737, N3607, N6134);
buf BUF1 (N11748, N11741);
and AND2 (N11749, N11744, N10233);
xor XOR2 (N11750, N11738, N3525);
buf BUF1 (N11751, N11747);
nand NAND2 (N11752, N11732, N8162);
not NOT1 (N11753, N11745);
and AND4 (N11754, N11750, N680, N1, N4125);
nor NOR4 (N11755, N11752, N1689, N7565, N7528);
or OR3 (N11756, N11703, N6519, N83);
or OR2 (N11757, N11751, N1911);
xor XOR2 (N11758, N11748, N7980);
and AND2 (N11759, N11726, N5817);
and AND4 (N11760, N11757, N11172, N6530, N1881);
xor XOR2 (N11761, N11749, N4332);
nor NOR2 (N11762, N11758, N8600);
and AND4 (N11763, N11755, N799, N7412, N1649);
nor NOR3 (N11764, N11753, N2819, N11202);
buf BUF1 (N11765, N11761);
buf BUF1 (N11766, N11728);
xor XOR2 (N11767, N11765, N6961);
nand NAND3 (N11768, N11759, N10769, N1281);
buf BUF1 (N11769, N11760);
nand NAND4 (N11770, N11769, N6776, N3184, N341);
nor NOR3 (N11771, N11756, N3931, N7249);
not NOT1 (N11772, N11766);
nor NOR4 (N11773, N11772, N8313, N4025, N432);
nand NAND2 (N11774, N11754, N598);
nand NAND4 (N11775, N11771, N6059, N4890, N1225);
or OR4 (N11776, N11773, N4843, N11712, N155);
and AND4 (N11777, N11776, N10379, N84, N9401);
and AND2 (N11778, N11764, N7622);
not NOT1 (N11779, N11763);
xor XOR2 (N11780, N11778, N8963);
and AND3 (N11781, N11779, N6602, N5568);
not NOT1 (N11782, N11770);
xor XOR2 (N11783, N11767, N4368);
nand NAND4 (N11784, N11768, N4969, N4173, N3743);
nor NOR4 (N11785, N11783, N7696, N9346, N11569);
nor NOR3 (N11786, N11781, N6621, N6837);
buf BUF1 (N11787, N11780);
nor NOR3 (N11788, N11787, N6693, N280);
buf BUF1 (N11789, N11788);
or OR2 (N11790, N11746, N1906);
nand NAND3 (N11791, N11790, N10098, N1114);
nand NAND4 (N11792, N11762, N673, N10387, N9201);
or OR4 (N11793, N11786, N4360, N6132, N1591);
and AND3 (N11794, N11792, N737, N980);
and AND4 (N11795, N11775, N10260, N3393, N7728);
xor XOR2 (N11796, N11795, N3666);
nand NAND4 (N11797, N11793, N10180, N628, N187);
xor XOR2 (N11798, N11797, N4286);
not NOT1 (N11799, N11784);
buf BUF1 (N11800, N11799);
not NOT1 (N11801, N11794);
buf BUF1 (N11802, N11785);
xor XOR2 (N11803, N11801, N4520);
xor XOR2 (N11804, N11791, N9254);
not NOT1 (N11805, N11774);
xor XOR2 (N11806, N11789, N4099);
xor XOR2 (N11807, N11796, N1716);
nand NAND2 (N11808, N11798, N7703);
xor XOR2 (N11809, N11804, N3125);
buf BUF1 (N11810, N11808);
nor NOR4 (N11811, N11800, N4147, N8010, N11758);
xor XOR2 (N11812, N11806, N8087);
xor XOR2 (N11813, N11812, N620);
xor XOR2 (N11814, N11810, N11166);
nand NAND4 (N11815, N11782, N5879, N416, N9771);
not NOT1 (N11816, N11813);
and AND4 (N11817, N11803, N9684, N906, N10477);
xor XOR2 (N11818, N11777, N7737);
nor NOR3 (N11819, N11811, N5555, N11653);
nand NAND3 (N11820, N11802, N8206, N9829);
nor NOR2 (N11821, N11819, N10498);
nor NOR4 (N11822, N11818, N224, N6091, N7131);
nor NOR2 (N11823, N11822, N9558);
and AND2 (N11824, N11817, N9296);
buf BUF1 (N11825, N11824);
xor XOR2 (N11826, N11820, N11679);
xor XOR2 (N11827, N11805, N5455);
buf BUF1 (N11828, N11821);
or OR3 (N11829, N11823, N100, N8326);
not NOT1 (N11830, N11816);
nand NAND2 (N11831, N11807, N4252);
buf BUF1 (N11832, N11814);
or OR3 (N11833, N11809, N96, N622);
xor XOR2 (N11834, N11815, N590);
nand NAND2 (N11835, N11826, N898);
or OR4 (N11836, N11828, N1275, N4736, N7199);
nand NAND2 (N11837, N11827, N2927);
buf BUF1 (N11838, N11834);
xor XOR2 (N11839, N11831, N9029);
nand NAND2 (N11840, N11838, N996);
nand NAND3 (N11841, N11832, N3608, N10142);
nor NOR4 (N11842, N11836, N1726, N10116, N9047);
and AND4 (N11843, N11825, N3882, N3771, N4026);
xor XOR2 (N11844, N11830, N5139);
not NOT1 (N11845, N11840);
and AND2 (N11846, N11845, N4924);
buf BUF1 (N11847, N11833);
xor XOR2 (N11848, N11847, N3457);
xor XOR2 (N11849, N11837, N2613);
and AND4 (N11850, N11844, N6121, N9351, N7382);
and AND4 (N11851, N11846, N1992, N8693, N7995);
or OR3 (N11852, N11843, N1530, N6226);
not NOT1 (N11853, N11829);
not NOT1 (N11854, N11842);
xor XOR2 (N11855, N11849, N11731);
or OR3 (N11856, N11839, N3496, N7084);
xor XOR2 (N11857, N11854, N3423);
xor XOR2 (N11858, N11855, N1302);
xor XOR2 (N11859, N11857, N6449);
and AND4 (N11860, N11859, N663, N11690, N6386);
nand NAND4 (N11861, N11835, N3377, N3594, N11611);
not NOT1 (N11862, N11848);
nand NAND2 (N11863, N11858, N7097);
xor XOR2 (N11864, N11841, N8433);
and AND4 (N11865, N11864, N4812, N5938, N5041);
and AND3 (N11866, N11851, N1463, N893);
nor NOR2 (N11867, N11863, N7669);
xor XOR2 (N11868, N11866, N2037);
or OR2 (N11869, N11856, N8812);
not NOT1 (N11870, N11865);
not NOT1 (N11871, N11861);
buf BUF1 (N11872, N11850);
and AND2 (N11873, N11852, N8084);
and AND4 (N11874, N11871, N10704, N833, N6935);
nand NAND2 (N11875, N11874, N7469);
buf BUF1 (N11876, N11873);
nor NOR3 (N11877, N11870, N10330, N9421);
xor XOR2 (N11878, N11876, N3698);
nor NOR2 (N11879, N11868, N4542);
or OR2 (N11880, N11862, N11274);
not NOT1 (N11881, N11879);
or OR4 (N11882, N11880, N6276, N9941, N11804);
and AND4 (N11883, N11877, N3604, N7258, N17);
not NOT1 (N11884, N11872);
xor XOR2 (N11885, N11875, N6007);
buf BUF1 (N11886, N11884);
xor XOR2 (N11887, N11867, N1328);
nor NOR4 (N11888, N11885, N334, N9287, N6059);
xor XOR2 (N11889, N11860, N11405);
xor XOR2 (N11890, N11886, N3944);
xor XOR2 (N11891, N11881, N11457);
not NOT1 (N11892, N11890);
or OR3 (N11893, N11878, N6909, N3115);
not NOT1 (N11894, N11883);
nand NAND2 (N11895, N11869, N4668);
xor XOR2 (N11896, N11889, N11229);
buf BUF1 (N11897, N11887);
xor XOR2 (N11898, N11893, N10452);
buf BUF1 (N11899, N11894);
not NOT1 (N11900, N11882);
not NOT1 (N11901, N11897);
or OR3 (N11902, N11853, N3236, N5787);
buf BUF1 (N11903, N11896);
nand NAND4 (N11904, N11899, N6803, N3968, N2559);
buf BUF1 (N11905, N11892);
xor XOR2 (N11906, N11904, N5239);
xor XOR2 (N11907, N11903, N1102);
not NOT1 (N11908, N11901);
or OR3 (N11909, N11900, N2168, N1175);
buf BUF1 (N11910, N11891);
xor XOR2 (N11911, N11895, N1191);
nand NAND3 (N11912, N11898, N11192, N10113);
buf BUF1 (N11913, N11912);
and AND4 (N11914, N11913, N947, N11729, N295);
nor NOR4 (N11915, N11907, N5390, N3081, N7133);
and AND3 (N11916, N11915, N1214, N747);
or OR2 (N11917, N11914, N897);
not NOT1 (N11918, N11909);
nor NOR3 (N11919, N11905, N7536, N318);
and AND2 (N11920, N11910, N9807);
buf BUF1 (N11921, N11911);
and AND3 (N11922, N11902, N9276, N11533);
nor NOR3 (N11923, N11921, N1101, N3657);
or OR3 (N11924, N11919, N4667, N9491);
nand NAND4 (N11925, N11906, N11307, N5634, N5954);
xor XOR2 (N11926, N11908, N8449);
not NOT1 (N11927, N11925);
not NOT1 (N11928, N11888);
xor XOR2 (N11929, N11924, N5632);
buf BUF1 (N11930, N11917);
not NOT1 (N11931, N11927);
nor NOR4 (N11932, N11922, N9406, N2978, N10839);
nand NAND3 (N11933, N11916, N814, N478);
nand NAND4 (N11934, N11930, N948, N11234, N8225);
buf BUF1 (N11935, N11931);
and AND3 (N11936, N11929, N4013, N5687);
not NOT1 (N11937, N11936);
xor XOR2 (N11938, N11918, N5283);
and AND4 (N11939, N11934, N9380, N2892, N4040);
xor XOR2 (N11940, N11926, N1832);
nand NAND4 (N11941, N11932, N627, N8307, N4847);
and AND3 (N11942, N11933, N107, N4373);
nand NAND2 (N11943, N11942, N2755);
nand NAND3 (N11944, N11940, N7113, N9212);
nand NAND3 (N11945, N11920, N6701, N8096);
buf BUF1 (N11946, N11944);
buf BUF1 (N11947, N11928);
not NOT1 (N11948, N11943);
nand NAND4 (N11949, N11941, N9478, N6270, N9795);
and AND4 (N11950, N11937, N8590, N4874, N5418);
or OR2 (N11951, N11949, N1963);
nand NAND3 (N11952, N11939, N495, N7316);
buf BUF1 (N11953, N11946);
or OR2 (N11954, N11951, N4390);
or OR2 (N11955, N11938, N7115);
or OR4 (N11956, N11935, N10394, N4157, N10740);
and AND3 (N11957, N11953, N1444, N5087);
or OR3 (N11958, N11947, N3857, N5290);
not NOT1 (N11959, N11957);
nand NAND2 (N11960, N11952, N9808);
and AND3 (N11961, N11960, N6340, N6049);
xor XOR2 (N11962, N11961, N3260);
xor XOR2 (N11963, N11950, N10979);
not NOT1 (N11964, N11923);
and AND2 (N11965, N11963, N10426);
or OR3 (N11966, N11959, N4846, N3845);
xor XOR2 (N11967, N11945, N1479);
or OR2 (N11968, N11954, N9821);
nand NAND2 (N11969, N11948, N7238);
buf BUF1 (N11970, N11967);
not NOT1 (N11971, N11970);
buf BUF1 (N11972, N11958);
nor NOR2 (N11973, N11966, N2690);
nor NOR3 (N11974, N11972, N2816, N1092);
or OR2 (N11975, N11974, N9294);
buf BUF1 (N11976, N11971);
nand NAND2 (N11977, N11973, N10055);
and AND2 (N11978, N11969, N7465);
nor NOR4 (N11979, N11955, N10542, N5215, N3748);
and AND4 (N11980, N11964, N4568, N10171, N10102);
not NOT1 (N11981, N11965);
not NOT1 (N11982, N11979);
not NOT1 (N11983, N11981);
buf BUF1 (N11984, N11962);
nor NOR2 (N11985, N11983, N393);
xor XOR2 (N11986, N11975, N10836);
nand NAND2 (N11987, N11968, N3544);
and AND4 (N11988, N11987, N9694, N4991, N1223);
nor NOR4 (N11989, N11986, N176, N11927, N7908);
xor XOR2 (N11990, N11956, N9125);
or OR3 (N11991, N11984, N11538, N2772);
xor XOR2 (N11992, N11982, N6054);
xor XOR2 (N11993, N11980, N4437);
xor XOR2 (N11994, N11992, N9696);
or OR3 (N11995, N11988, N744, N2830);
nor NOR2 (N11996, N11993, N10073);
buf BUF1 (N11997, N11990);
nor NOR3 (N11998, N11985, N6645, N4255);
nand NAND2 (N11999, N11977, N9019);
and AND2 (N12000, N11995, N9869);
xor XOR2 (N12001, N11999, N4970);
xor XOR2 (N12002, N12000, N9902);
and AND2 (N12003, N11976, N11211);
nand NAND2 (N12004, N11996, N7236);
nand NAND2 (N12005, N12002, N11893);
not NOT1 (N12006, N12003);
xor XOR2 (N12007, N12005, N6302);
or OR2 (N12008, N12004, N6812);
and AND4 (N12009, N12001, N597, N6951, N2816);
and AND4 (N12010, N11997, N4424, N6625, N5627);
buf BUF1 (N12011, N11991);
or OR4 (N12012, N11989, N8173, N3514, N1906);
nand NAND2 (N12013, N12008, N4687);
not NOT1 (N12014, N12011);
and AND3 (N12015, N12013, N7684, N8911);
or OR3 (N12016, N12010, N3002, N7164);
and AND3 (N12017, N11998, N5405, N7983);
buf BUF1 (N12018, N12006);
or OR2 (N12019, N12007, N627);
buf BUF1 (N12020, N12018);
nor NOR4 (N12021, N12020, N10431, N699, N11220);
xor XOR2 (N12022, N11978, N2702);
xor XOR2 (N12023, N12022, N7379);
not NOT1 (N12024, N12017);
nand NAND4 (N12025, N12023, N9744, N11426, N11298);
nor NOR3 (N12026, N12025, N4631, N4717);
nand NAND3 (N12027, N12026, N7321, N5843);
xor XOR2 (N12028, N11994, N4360);
nor NOR4 (N12029, N12028, N9489, N11482, N9645);
and AND3 (N12030, N12021, N9909, N11809);
nor NOR3 (N12031, N12027, N11528, N11177);
buf BUF1 (N12032, N12030);
xor XOR2 (N12033, N12029, N6035);
nand NAND4 (N12034, N12019, N6561, N2370, N4924);
nor NOR4 (N12035, N12031, N9384, N5970, N10775);
xor XOR2 (N12036, N12035, N7052);
and AND3 (N12037, N12036, N10081, N10746);
or OR4 (N12038, N12012, N7220, N2687, N7992);
buf BUF1 (N12039, N12024);
xor XOR2 (N12040, N12038, N3504);
not NOT1 (N12041, N12033);
or OR3 (N12042, N12032, N10969, N7880);
nand NAND2 (N12043, N12034, N10131);
and AND2 (N12044, N12043, N7864);
and AND4 (N12045, N12014, N4257, N4603, N9468);
xor XOR2 (N12046, N12009, N2479);
nand NAND4 (N12047, N12015, N7671, N4897, N9313);
nor NOR2 (N12048, N12040, N7794);
buf BUF1 (N12049, N12041);
or OR3 (N12050, N12045, N6399, N7582);
not NOT1 (N12051, N12044);
and AND3 (N12052, N12042, N4937, N8290);
buf BUF1 (N12053, N12016);
and AND3 (N12054, N12037, N8359, N10249);
not NOT1 (N12055, N12047);
nor NOR4 (N12056, N12054, N5151, N5912, N2595);
xor XOR2 (N12057, N12048, N27);
xor XOR2 (N12058, N12057, N6319);
or OR3 (N12059, N12039, N6703, N5549);
not NOT1 (N12060, N12058);
buf BUF1 (N12061, N12050);
nand NAND3 (N12062, N12051, N3805, N4784);
and AND3 (N12063, N12062, N4395, N9646);
and AND3 (N12064, N12060, N479, N1176);
nand NAND3 (N12065, N12061, N4210, N11278);
xor XOR2 (N12066, N12052, N8479);
nand NAND4 (N12067, N12063, N1318, N982, N3877);
buf BUF1 (N12068, N12065);
buf BUF1 (N12069, N12055);
not NOT1 (N12070, N12059);
nand NAND2 (N12071, N12070, N7976);
buf BUF1 (N12072, N12053);
nand NAND2 (N12073, N12068, N3573);
buf BUF1 (N12074, N12056);
or OR4 (N12075, N12066, N8675, N4180, N11800);
not NOT1 (N12076, N12073);
buf BUF1 (N12077, N12049);
buf BUF1 (N12078, N12067);
nand NAND2 (N12079, N12077, N1627);
nand NAND4 (N12080, N12075, N9178, N3665, N5108);
buf BUF1 (N12081, N12064);
nand NAND2 (N12082, N12078, N924);
buf BUF1 (N12083, N12076);
nand NAND3 (N12084, N12069, N3000, N9465);
nand NAND4 (N12085, N12083, N5763, N5106, N3024);
nand NAND2 (N12086, N12084, N6360);
buf BUF1 (N12087, N12046);
nor NOR3 (N12088, N12072, N5636, N5087);
buf BUF1 (N12089, N12086);
xor XOR2 (N12090, N12080, N3203);
xor XOR2 (N12091, N12081, N3170);
xor XOR2 (N12092, N12089, N2807);
nor NOR2 (N12093, N12071, N1851);
nor NOR4 (N12094, N12090, N410, N9119, N2606);
not NOT1 (N12095, N12074);
buf BUF1 (N12096, N12085);
nor NOR2 (N12097, N12088, N11284);
and AND4 (N12098, N12096, N4433, N4996, N1212);
nor NOR2 (N12099, N12082, N11468);
nor NOR4 (N12100, N12079, N1526, N8151, N9055);
nand NAND3 (N12101, N12100, N6092, N3925);
and AND4 (N12102, N12091, N3912, N320, N8121);
nand NAND2 (N12103, N12093, N22);
buf BUF1 (N12104, N12102);
or OR4 (N12105, N12092, N3321, N9077, N3865);
nor NOR3 (N12106, N12095, N7077, N1144);
nand NAND4 (N12107, N12105, N163, N3789, N3843);
nand NAND3 (N12108, N12099, N9179, N450);
or OR3 (N12109, N12103, N7208, N8538);
or OR3 (N12110, N12098, N11660, N5128);
buf BUF1 (N12111, N12110);
nand NAND3 (N12112, N12108, N5781, N5624);
nor NOR3 (N12113, N12094, N1764, N2332);
xor XOR2 (N12114, N12087, N6897);
nor NOR3 (N12115, N12107, N11241, N3179);
nor NOR4 (N12116, N12101, N10878, N104, N3958);
and AND4 (N12117, N12114, N8120, N1389, N10620);
buf BUF1 (N12118, N12116);
nor NOR2 (N12119, N12112, N5812);
not NOT1 (N12120, N12113);
and AND3 (N12121, N12117, N10802, N1163);
xor XOR2 (N12122, N12118, N2832);
not NOT1 (N12123, N12119);
buf BUF1 (N12124, N12104);
nand NAND2 (N12125, N12109, N1098);
or OR4 (N12126, N12121, N868, N11836, N6631);
nand NAND4 (N12127, N12122, N3565, N10713, N608);
and AND3 (N12128, N12106, N4640, N8413);
or OR4 (N12129, N12127, N7871, N9372, N2963);
nor NOR2 (N12130, N12111, N11717);
or OR3 (N12131, N12126, N3435, N2367);
nor NOR3 (N12132, N12130, N10382, N9473);
or OR3 (N12133, N12124, N9297, N5790);
xor XOR2 (N12134, N12132, N10545);
buf BUF1 (N12135, N12123);
nor NOR2 (N12136, N12097, N706);
or OR2 (N12137, N12115, N2095);
or OR4 (N12138, N12128, N4493, N9020, N1215);
or OR4 (N12139, N12135, N80, N2960, N3823);
nor NOR3 (N12140, N12131, N9015, N7545);
xor XOR2 (N12141, N12133, N5246);
nand NAND4 (N12142, N12120, N7126, N2712, N2631);
buf BUF1 (N12143, N12142);
not NOT1 (N12144, N12125);
xor XOR2 (N12145, N12137, N7579);
nor NOR4 (N12146, N12139, N5877, N7995, N5561);
nand NAND3 (N12147, N12144, N2279, N7931);
and AND2 (N12148, N12129, N6798);
nand NAND2 (N12149, N12138, N10753);
not NOT1 (N12150, N12146);
xor XOR2 (N12151, N12134, N10089);
buf BUF1 (N12152, N12148);
buf BUF1 (N12153, N12141);
and AND3 (N12154, N12136, N6881, N9253);
or OR2 (N12155, N12147, N5061);
nand NAND2 (N12156, N12154, N11031);
buf BUF1 (N12157, N12155);
and AND2 (N12158, N12145, N3690);
or OR3 (N12159, N12157, N9398, N1227);
or OR2 (N12160, N12150, N2632);
xor XOR2 (N12161, N12159, N2801);
or OR4 (N12162, N12153, N3868, N1165, N3093);
xor XOR2 (N12163, N12143, N11545);
xor XOR2 (N12164, N12151, N9906);
or OR2 (N12165, N12140, N10790);
buf BUF1 (N12166, N12161);
buf BUF1 (N12167, N12165);
buf BUF1 (N12168, N12152);
nand NAND3 (N12169, N12167, N11847, N6943);
and AND2 (N12170, N12164, N4166);
xor XOR2 (N12171, N12156, N3782);
not NOT1 (N12172, N12162);
xor XOR2 (N12173, N12163, N10393);
or OR4 (N12174, N12173, N3184, N9465, N934);
xor XOR2 (N12175, N12166, N11743);
xor XOR2 (N12176, N12160, N5467);
nor NOR4 (N12177, N12158, N230, N7761, N11414);
nor NOR4 (N12178, N12175, N11947, N4818, N8917);
not NOT1 (N12179, N12171);
not NOT1 (N12180, N12176);
or OR3 (N12181, N12168, N6904, N2533);
nand NAND3 (N12182, N12180, N11991, N6577);
nor NOR4 (N12183, N12179, N11333, N5690, N2945);
not NOT1 (N12184, N12177);
not NOT1 (N12185, N12183);
nor NOR4 (N12186, N12170, N6448, N3248, N10519);
buf BUF1 (N12187, N12174);
nor NOR3 (N12188, N12187, N2934, N11799);
or OR4 (N12189, N12182, N4358, N7782, N1360);
buf BUF1 (N12190, N12149);
buf BUF1 (N12191, N12184);
nor NOR2 (N12192, N12178, N11452);
xor XOR2 (N12193, N12190, N4069);
or OR2 (N12194, N12181, N4323);
and AND3 (N12195, N12169, N4965, N6114);
or OR2 (N12196, N12172, N3068);
buf BUF1 (N12197, N12189);
and AND2 (N12198, N12197, N3578);
and AND4 (N12199, N12198, N12118, N1000, N9272);
xor XOR2 (N12200, N12186, N4565);
and AND2 (N12201, N12196, N395);
or OR2 (N12202, N12195, N10955);
not NOT1 (N12203, N12199);
and AND3 (N12204, N12200, N8677, N12157);
nand NAND4 (N12205, N12194, N11758, N10608, N863);
not NOT1 (N12206, N12188);
xor XOR2 (N12207, N12205, N3407);
and AND2 (N12208, N12207, N2391);
buf BUF1 (N12209, N12193);
buf BUF1 (N12210, N12209);
buf BUF1 (N12211, N12202);
buf BUF1 (N12212, N12210);
xor XOR2 (N12213, N12212, N8370);
nand NAND3 (N12214, N12208, N6913, N428);
buf BUF1 (N12215, N12201);
xor XOR2 (N12216, N12192, N7958);
nor NOR4 (N12217, N12211, N9857, N11128, N3241);
or OR3 (N12218, N12216, N11817, N2459);
nand NAND3 (N12219, N12217, N3137, N12024);
xor XOR2 (N12220, N12218, N8995);
buf BUF1 (N12221, N12204);
not NOT1 (N12222, N12215);
nand NAND3 (N12223, N12185, N10946, N1608);
nor NOR4 (N12224, N12221, N5559, N4151, N3653);
nand NAND3 (N12225, N12191, N3029, N9669);
or OR4 (N12226, N12224, N9766, N3840, N7352);
or OR4 (N12227, N12225, N6938, N4509, N8647);
and AND3 (N12228, N12203, N9212, N492);
nor NOR2 (N12229, N12214, N8256);
and AND3 (N12230, N12226, N7725, N4109);
buf BUF1 (N12231, N12219);
not NOT1 (N12232, N12223);
nor NOR2 (N12233, N12222, N7069);
nor NOR2 (N12234, N12220, N1025);
or OR2 (N12235, N12213, N5518);
nand NAND2 (N12236, N12232, N2359);
or OR4 (N12237, N12228, N2973, N7557, N12140);
xor XOR2 (N12238, N12233, N5694);
nand NAND4 (N12239, N12234, N3007, N7137, N313);
buf BUF1 (N12240, N12235);
not NOT1 (N12241, N12236);
xor XOR2 (N12242, N12238, N53);
not NOT1 (N12243, N12242);
nor NOR3 (N12244, N12237, N9759, N10997);
not NOT1 (N12245, N12243);
or OR4 (N12246, N12227, N2283, N6991, N8067);
not NOT1 (N12247, N12241);
xor XOR2 (N12248, N12230, N11754);
and AND4 (N12249, N12246, N5610, N2429, N4565);
buf BUF1 (N12250, N12244);
buf BUF1 (N12251, N12247);
nand NAND2 (N12252, N12251, N8807);
nor NOR2 (N12253, N12249, N1721);
xor XOR2 (N12254, N12231, N1339);
xor XOR2 (N12255, N12206, N5134);
nor NOR2 (N12256, N12253, N6953);
nand NAND3 (N12257, N12252, N3768, N2822);
not NOT1 (N12258, N12254);
and AND4 (N12259, N12255, N7076, N8434, N5723);
or OR3 (N12260, N12240, N1103, N5598);
buf BUF1 (N12261, N12258);
xor XOR2 (N12262, N12239, N9873);
buf BUF1 (N12263, N12256);
nor NOR3 (N12264, N12248, N10871, N1838);
and AND3 (N12265, N12245, N8432, N5719);
nor NOR3 (N12266, N12257, N6699, N13);
or OR3 (N12267, N12265, N2454, N5315);
and AND2 (N12268, N12267, N2388);
nor NOR3 (N12269, N12260, N2925, N6182);
not NOT1 (N12270, N12250);
and AND3 (N12271, N12229, N12123, N1483);
or OR4 (N12272, N12268, N9857, N3479, N836);
nor NOR2 (N12273, N12270, N5391);
xor XOR2 (N12274, N12272, N8110);
or OR4 (N12275, N12263, N9207, N2811, N5133);
nand NAND4 (N12276, N12275, N5559, N7012, N8813);
xor XOR2 (N12277, N12274, N6290);
xor XOR2 (N12278, N12273, N8133);
and AND3 (N12279, N12262, N10844, N2162);
or OR3 (N12280, N12259, N11021, N193);
nand NAND3 (N12281, N12276, N2840, N1056);
xor XOR2 (N12282, N12279, N3793);
xor XOR2 (N12283, N12278, N5747);
not NOT1 (N12284, N12261);
nor NOR3 (N12285, N12284, N8359, N10781);
and AND4 (N12286, N12269, N3954, N11505, N3749);
nand NAND2 (N12287, N12280, N820);
nand NAND4 (N12288, N12277, N39, N4348, N6973);
nor NOR3 (N12289, N12281, N11044, N10153);
xor XOR2 (N12290, N12283, N6562);
not NOT1 (N12291, N12282);
and AND4 (N12292, N12289, N11848, N1094, N360);
not NOT1 (N12293, N12291);
or OR4 (N12294, N12288, N3357, N10205, N12002);
not NOT1 (N12295, N12286);
nor NOR2 (N12296, N12292, N7846);
nor NOR2 (N12297, N12294, N6039);
nor NOR2 (N12298, N12296, N8283);
not NOT1 (N12299, N12293);
and AND2 (N12300, N12299, N483);
buf BUF1 (N12301, N12297);
not NOT1 (N12302, N12301);
xor XOR2 (N12303, N12285, N6299);
buf BUF1 (N12304, N12290);
buf BUF1 (N12305, N12264);
nor NOR3 (N12306, N12266, N7871, N8171);
not NOT1 (N12307, N12304);
and AND3 (N12308, N12287, N11928, N5591);
nand NAND2 (N12309, N12295, N8829);
buf BUF1 (N12310, N12306);
nor NOR3 (N12311, N12305, N10189, N7807);
nor NOR3 (N12312, N12302, N11918, N3777);
buf BUF1 (N12313, N12271);
nand NAND4 (N12314, N12311, N3984, N3378, N9419);
or OR2 (N12315, N12308, N604);
buf BUF1 (N12316, N12312);
and AND3 (N12317, N12316, N11781, N11871);
and AND4 (N12318, N12313, N2906, N9755, N9987);
xor XOR2 (N12319, N12310, N2802);
nand NAND4 (N12320, N12319, N1413, N551, N7883);
nand NAND3 (N12321, N12300, N4390, N5391);
and AND4 (N12322, N12320, N9273, N8768, N11514);
nand NAND2 (N12323, N12298, N6330);
not NOT1 (N12324, N12314);
xor XOR2 (N12325, N12324, N8338);
nor NOR4 (N12326, N12321, N11481, N11701, N10515);
not NOT1 (N12327, N12325);
or OR3 (N12328, N12307, N9711, N2953);
nor NOR3 (N12329, N12309, N5957, N2109);
or OR2 (N12330, N12328, N4734);
and AND4 (N12331, N12323, N10842, N4812, N10174);
nor NOR3 (N12332, N12329, N11247, N3070);
nor NOR4 (N12333, N12317, N7684, N7053, N10653);
buf BUF1 (N12334, N12326);
and AND2 (N12335, N12330, N6453);
not NOT1 (N12336, N12318);
nand NAND3 (N12337, N12303, N9050, N2699);
nand NAND4 (N12338, N12322, N6860, N10108, N134);
nor NOR3 (N12339, N12335, N7379, N8594);
and AND3 (N12340, N12327, N7974, N4422);
not NOT1 (N12341, N12339);
and AND3 (N12342, N12336, N10938, N6766);
nand NAND3 (N12343, N12332, N10405, N10654);
not NOT1 (N12344, N12343);
buf BUF1 (N12345, N12331);
not NOT1 (N12346, N12345);
nand NAND3 (N12347, N12342, N2347, N2154);
nor NOR4 (N12348, N12344, N10186, N5095, N951);
buf BUF1 (N12349, N12334);
nor NOR4 (N12350, N12337, N6758, N9817, N10792);
nor NOR4 (N12351, N12348, N2663, N11086, N5607);
buf BUF1 (N12352, N12338);
and AND3 (N12353, N12346, N11713, N11055);
nand NAND2 (N12354, N12341, N11803);
xor XOR2 (N12355, N12351, N10767);
and AND2 (N12356, N12354, N6562);
or OR4 (N12357, N12349, N4068, N2818, N7664);
buf BUF1 (N12358, N12333);
and AND4 (N12359, N12347, N12112, N5534, N5077);
not NOT1 (N12360, N12357);
nand NAND2 (N12361, N12355, N4078);
or OR4 (N12362, N12356, N4962, N1992, N6189);
xor XOR2 (N12363, N12350, N6838);
and AND4 (N12364, N12352, N8715, N5163, N3322);
nand NAND4 (N12365, N12353, N1498, N9721, N5625);
not NOT1 (N12366, N12365);
nor NOR2 (N12367, N12360, N1430);
xor XOR2 (N12368, N12367, N2305);
xor XOR2 (N12369, N12361, N10254);
nor NOR4 (N12370, N12366, N3191, N989, N2024);
buf BUF1 (N12371, N12363);
and AND2 (N12372, N12370, N7623);
or OR2 (N12373, N12372, N44);
nor NOR2 (N12374, N12362, N2850);
nand NAND3 (N12375, N12369, N1483, N1775);
or OR2 (N12376, N12359, N5951);
buf BUF1 (N12377, N12364);
nand NAND4 (N12378, N12315, N5239, N8252, N1725);
buf BUF1 (N12379, N12376);
and AND3 (N12380, N12377, N11336, N5891);
and AND3 (N12381, N12373, N1046, N11387);
nand NAND2 (N12382, N12380, N6755);
nand NAND3 (N12383, N12382, N2513, N8619);
or OR2 (N12384, N12381, N6282);
nor NOR4 (N12385, N12379, N9685, N2938, N2924);
nor NOR3 (N12386, N12375, N8141, N5754);
or OR4 (N12387, N12368, N4881, N8044, N2905);
or OR3 (N12388, N12383, N6806, N2971);
and AND4 (N12389, N12384, N2548, N10550, N5222);
xor XOR2 (N12390, N12358, N194);
and AND2 (N12391, N12385, N10976);
buf BUF1 (N12392, N12389);
buf BUF1 (N12393, N12391);
and AND4 (N12394, N12378, N10072, N6146, N11597);
xor XOR2 (N12395, N12371, N2235);
nor NOR3 (N12396, N12392, N1734, N2073);
buf BUF1 (N12397, N12394);
not NOT1 (N12398, N12387);
or OR3 (N12399, N12395, N1691, N10825);
not NOT1 (N12400, N12398);
xor XOR2 (N12401, N12388, N9477);
buf BUF1 (N12402, N12396);
and AND4 (N12403, N12393, N9787, N5882, N9678);
not NOT1 (N12404, N12397);
and AND2 (N12405, N12386, N1066);
not NOT1 (N12406, N12403);
xor XOR2 (N12407, N12402, N1282);
not NOT1 (N12408, N12400);
buf BUF1 (N12409, N12401);
buf BUF1 (N12410, N12406);
nand NAND4 (N12411, N12399, N154, N6086, N11319);
buf BUF1 (N12412, N12408);
not NOT1 (N12413, N12340);
xor XOR2 (N12414, N12413, N8619);
nand NAND3 (N12415, N12407, N635, N7642);
and AND2 (N12416, N12405, N5476);
xor XOR2 (N12417, N12410, N10621);
buf BUF1 (N12418, N12417);
xor XOR2 (N12419, N12411, N3697);
nand NAND3 (N12420, N12412, N11595, N867);
not NOT1 (N12421, N12415);
and AND2 (N12422, N12409, N10799);
nand NAND4 (N12423, N12414, N3756, N2162, N2527);
nand NAND4 (N12424, N12404, N1966, N3831, N287);
nor NOR2 (N12425, N12423, N3287);
xor XOR2 (N12426, N12418, N8408);
xor XOR2 (N12427, N12419, N1071);
nand NAND3 (N12428, N12427, N3712, N5902);
buf BUF1 (N12429, N12422);
xor XOR2 (N12430, N12374, N6340);
or OR3 (N12431, N12421, N12238, N5980);
nand NAND4 (N12432, N12420, N7958, N7548, N6818);
buf BUF1 (N12433, N12428);
or OR2 (N12434, N12431, N6832);
or OR2 (N12435, N12429, N2542);
nand NAND3 (N12436, N12433, N1303, N2291);
nand NAND2 (N12437, N12436, N6030);
nor NOR3 (N12438, N12434, N1912, N5944);
nand NAND2 (N12439, N12424, N9755);
and AND3 (N12440, N12425, N8933, N11752);
xor XOR2 (N12441, N12439, N11319);
and AND4 (N12442, N12435, N1334, N11561, N439);
buf BUF1 (N12443, N12442);
buf BUF1 (N12444, N12426);
and AND2 (N12445, N12430, N3218);
xor XOR2 (N12446, N12416, N2061);
nor NOR2 (N12447, N12432, N2889);
xor XOR2 (N12448, N12440, N5205);
buf BUF1 (N12449, N12448);
and AND2 (N12450, N12441, N4646);
not NOT1 (N12451, N12445);
and AND3 (N12452, N12449, N7232, N6895);
nor NOR4 (N12453, N12446, N1988, N11680, N4496);
nand NAND4 (N12454, N12444, N5384, N10474, N9048);
and AND3 (N12455, N12390, N11434, N7332);
buf BUF1 (N12456, N12450);
or OR4 (N12457, N12454, N10490, N10924, N7854);
nand NAND4 (N12458, N12456, N1627, N406, N3562);
xor XOR2 (N12459, N12437, N11758);
and AND3 (N12460, N12443, N10826, N10437);
or OR2 (N12461, N12451, N11552);
or OR4 (N12462, N12455, N1256, N5081, N4808);
xor XOR2 (N12463, N12453, N8666);
or OR4 (N12464, N12463, N12295, N4027, N234);
buf BUF1 (N12465, N12457);
nand NAND2 (N12466, N12438, N1378);
and AND3 (N12467, N12458, N11537, N10933);
and AND4 (N12468, N12462, N5536, N6597, N3667);
or OR4 (N12469, N12459, N241, N2946, N8542);
not NOT1 (N12470, N12461);
not NOT1 (N12471, N12467);
or OR2 (N12472, N12471, N9976);
buf BUF1 (N12473, N12469);
not NOT1 (N12474, N12468);
xor XOR2 (N12475, N12464, N6993);
and AND2 (N12476, N12475, N299);
not NOT1 (N12477, N12472);
or OR2 (N12478, N12452, N10699);
or OR2 (N12479, N12466, N8370);
nand NAND2 (N12480, N12476, N3528);
buf BUF1 (N12481, N12465);
nor NOR3 (N12482, N12473, N7940, N11299);
or OR2 (N12483, N12470, N4438);
xor XOR2 (N12484, N12478, N9980);
xor XOR2 (N12485, N12477, N5187);
or OR4 (N12486, N12479, N5751, N9749, N3301);
or OR4 (N12487, N12482, N4997, N10123, N8476);
or OR3 (N12488, N12481, N461, N8462);
or OR2 (N12489, N12485, N2811);
not NOT1 (N12490, N12460);
nor NOR3 (N12491, N12486, N4972, N10316);
not NOT1 (N12492, N12484);
nand NAND3 (N12493, N12487, N5885, N6610);
buf BUF1 (N12494, N12492);
not NOT1 (N12495, N12447);
nor NOR2 (N12496, N12491, N8743);
not NOT1 (N12497, N12490);
buf BUF1 (N12498, N12480);
xor XOR2 (N12499, N12474, N3433);
nor NOR3 (N12500, N12496, N4163, N673);
nand NAND2 (N12501, N12499, N8392);
xor XOR2 (N12502, N12495, N1754);
not NOT1 (N12503, N12494);
nand NAND4 (N12504, N12502, N1802, N9326, N1802);
not NOT1 (N12505, N12498);
or OR3 (N12506, N12497, N297, N1960);
buf BUF1 (N12507, N12483);
not NOT1 (N12508, N12500);
buf BUF1 (N12509, N12505);
and AND2 (N12510, N12501, N2233);
buf BUF1 (N12511, N12504);
and AND4 (N12512, N12493, N1675, N4023, N6828);
xor XOR2 (N12513, N12509, N1662);
nor NOR4 (N12514, N12511, N8101, N6743, N7408);
nor NOR2 (N12515, N12512, N8209);
nand NAND4 (N12516, N12507, N2262, N8765, N7529);
nand NAND4 (N12517, N12508, N7572, N7398, N4306);
nor NOR3 (N12518, N12513, N10127, N5741);
nand NAND4 (N12519, N12516, N4575, N3956, N3839);
buf BUF1 (N12520, N12489);
buf BUF1 (N12521, N12506);
nand NAND4 (N12522, N12510, N2438, N2863, N10977);
buf BUF1 (N12523, N12514);
or OR4 (N12524, N12519, N11156, N9380, N3260);
and AND3 (N12525, N12521, N2034, N8111);
nor NOR2 (N12526, N12518, N8652);
nand NAND4 (N12527, N12525, N4457, N8871, N10755);
and AND4 (N12528, N12515, N3711, N7772, N7120);
not NOT1 (N12529, N12517);
not NOT1 (N12530, N12526);
xor XOR2 (N12531, N12530, N3727);
nor NOR2 (N12532, N12531, N11785);
and AND2 (N12533, N12523, N9014);
xor XOR2 (N12534, N12532, N6773);
nor NOR4 (N12535, N12534, N2961, N10248, N6260);
buf BUF1 (N12536, N12533);
xor XOR2 (N12537, N12522, N9246);
xor XOR2 (N12538, N12536, N4600);
xor XOR2 (N12539, N12488, N8642);
xor XOR2 (N12540, N12538, N11166);
nor NOR3 (N12541, N12503, N3135, N8139);
or OR4 (N12542, N12524, N8800, N12287, N7537);
and AND3 (N12543, N12540, N5527, N6667);
nand NAND4 (N12544, N12541, N8257, N3135, N4412);
and AND4 (N12545, N12542, N4873, N2020, N9087);
buf BUF1 (N12546, N12528);
nor NOR3 (N12547, N12537, N697, N8357);
buf BUF1 (N12548, N12547);
and AND4 (N12549, N12520, N7332, N4180, N8225);
and AND4 (N12550, N12535, N3374, N12288, N5997);
and AND3 (N12551, N12539, N4911, N1869);
xor XOR2 (N12552, N12544, N8372);
not NOT1 (N12553, N12543);
xor XOR2 (N12554, N12529, N2946);
not NOT1 (N12555, N12549);
and AND3 (N12556, N12552, N7323, N8634);
nor NOR4 (N12557, N12553, N6096, N8320, N8489);
xor XOR2 (N12558, N12551, N5492);
and AND2 (N12559, N12558, N1895);
xor XOR2 (N12560, N12556, N8978);
xor XOR2 (N12561, N12545, N11657);
nand NAND2 (N12562, N12559, N9795);
nand NAND4 (N12563, N12550, N4122, N9438, N6356);
not NOT1 (N12564, N12546);
nand NAND4 (N12565, N12560, N7361, N1143, N3141);
nor NOR3 (N12566, N12564, N9338, N2620);
or OR4 (N12567, N12557, N1900, N7693, N6280);
buf BUF1 (N12568, N12555);
nor NOR3 (N12569, N12565, N12023, N8894);
or OR2 (N12570, N12566, N9213);
nand NAND2 (N12571, N12570, N9991);
nand NAND3 (N12572, N12567, N2782, N6307);
not NOT1 (N12573, N12527);
xor XOR2 (N12574, N12554, N3165);
buf BUF1 (N12575, N12561);
xor XOR2 (N12576, N12572, N11233);
xor XOR2 (N12577, N12548, N704);
or OR4 (N12578, N12568, N7739, N11852, N8849);
or OR3 (N12579, N12578, N11073, N11245);
buf BUF1 (N12580, N12575);
or OR4 (N12581, N12573, N8387, N9674, N304);
buf BUF1 (N12582, N12562);
xor XOR2 (N12583, N12579, N5006);
not NOT1 (N12584, N12569);
xor XOR2 (N12585, N12583, N9439);
or OR3 (N12586, N12584, N3171, N12550);
nor NOR2 (N12587, N12582, N4405);
nand NAND4 (N12588, N12585, N12318, N6761, N4769);
or OR4 (N12589, N12587, N12105, N3652, N9394);
nand NAND3 (N12590, N12563, N8473, N12031);
nor NOR4 (N12591, N12581, N5067, N10064, N2960);
or OR3 (N12592, N12586, N1663, N9224);
nand NAND4 (N12593, N12589, N8941, N7693, N7635);
nand NAND3 (N12594, N12588, N6163, N4658);
nor NOR2 (N12595, N12594, N3440);
or OR3 (N12596, N12576, N7828, N2704);
xor XOR2 (N12597, N12577, N11245);
nand NAND4 (N12598, N12592, N4762, N6844, N3809);
or OR4 (N12599, N12580, N2201, N297, N11587);
buf BUF1 (N12600, N12574);
nand NAND2 (N12601, N12597, N2912);
nand NAND2 (N12602, N12600, N7303);
nand NAND2 (N12603, N12591, N8383);
buf BUF1 (N12604, N12596);
or OR2 (N12605, N12593, N2431);
and AND2 (N12606, N12571, N6538);
buf BUF1 (N12607, N12601);
or OR4 (N12608, N12599, N11070, N1266, N10624);
nand NAND4 (N12609, N12607, N7777, N8337, N7068);
not NOT1 (N12610, N12603);
buf BUF1 (N12611, N12598);
nand NAND3 (N12612, N12605, N5582, N4040);
not NOT1 (N12613, N12590);
or OR4 (N12614, N12595, N10998, N6957, N2922);
xor XOR2 (N12615, N12611, N6270);
buf BUF1 (N12616, N12610);
nor NOR4 (N12617, N12606, N12418, N12265, N3294);
and AND2 (N12618, N12604, N10036);
xor XOR2 (N12619, N12602, N131);
and AND2 (N12620, N12615, N8479);
nor NOR4 (N12621, N12616, N260, N1001, N5386);
or OR2 (N12622, N12609, N4060);
buf BUF1 (N12623, N12612);
and AND3 (N12624, N12620, N7329, N5034);
buf BUF1 (N12625, N12617);
nor NOR4 (N12626, N12622, N977, N7403, N5852);
not NOT1 (N12627, N12613);
buf BUF1 (N12628, N12624);
not NOT1 (N12629, N12627);
nand NAND4 (N12630, N12608, N5232, N9249, N9936);
xor XOR2 (N12631, N12628, N5079);
xor XOR2 (N12632, N12621, N3819);
buf BUF1 (N12633, N12631);
nand NAND3 (N12634, N12623, N6458, N10551);
and AND4 (N12635, N12619, N12554, N1574, N6022);
and AND4 (N12636, N12635, N1521, N4734, N9718);
buf BUF1 (N12637, N12614);
buf BUF1 (N12638, N12625);
buf BUF1 (N12639, N12629);
xor XOR2 (N12640, N12638, N3062);
buf BUF1 (N12641, N12636);
nor NOR4 (N12642, N12634, N12219, N6097, N8690);
and AND4 (N12643, N12641, N7774, N6758, N9860);
nand NAND3 (N12644, N12642, N972, N7826);
buf BUF1 (N12645, N12633);
and AND4 (N12646, N12643, N10001, N2894, N7098);
xor XOR2 (N12647, N12639, N10961);
buf BUF1 (N12648, N12645);
nor NOR4 (N12649, N12646, N9837, N8238, N10846);
xor XOR2 (N12650, N12647, N5375);
not NOT1 (N12651, N12644);
xor XOR2 (N12652, N12632, N5569);
xor XOR2 (N12653, N12640, N9354);
xor XOR2 (N12654, N12618, N71);
and AND3 (N12655, N12648, N9251, N11771);
and AND2 (N12656, N12626, N5671);
nor NOR3 (N12657, N12656, N9170, N10086);
and AND2 (N12658, N12650, N5288);
not NOT1 (N12659, N12654);
not NOT1 (N12660, N12652);
not NOT1 (N12661, N12660);
not NOT1 (N12662, N12661);
xor XOR2 (N12663, N12649, N9061);
xor XOR2 (N12664, N12655, N6063);
buf BUF1 (N12665, N12653);
or OR3 (N12666, N12630, N2681, N566);
xor XOR2 (N12667, N12666, N11150);
nand NAND4 (N12668, N12659, N7390, N12629, N5893);
xor XOR2 (N12669, N12664, N10794);
not NOT1 (N12670, N12665);
and AND4 (N12671, N12667, N3374, N328, N2749);
not NOT1 (N12672, N12669);
nor NOR3 (N12673, N12670, N6374, N7666);
nor NOR4 (N12674, N12663, N9160, N7218, N3828);
nor NOR3 (N12675, N12637, N4102, N12333);
not NOT1 (N12676, N12651);
nand NAND3 (N12677, N12676, N10533, N7772);
buf BUF1 (N12678, N12658);
or OR2 (N12679, N12674, N9094);
xor XOR2 (N12680, N12677, N2478);
xor XOR2 (N12681, N12668, N8981);
buf BUF1 (N12682, N12662);
nor NOR4 (N12683, N12673, N11548, N10566, N7217);
nand NAND3 (N12684, N12678, N2499, N12563);
or OR4 (N12685, N12681, N7701, N2600, N3273);
nand NAND4 (N12686, N12683, N5470, N8167, N5576);
xor XOR2 (N12687, N12671, N3838);
xor XOR2 (N12688, N12685, N4948);
nand NAND3 (N12689, N12688, N3939, N11513);
buf BUF1 (N12690, N12686);
buf BUF1 (N12691, N12672);
xor XOR2 (N12692, N12679, N9988);
buf BUF1 (N12693, N12680);
not NOT1 (N12694, N12691);
nor NOR2 (N12695, N12692, N8869);
not NOT1 (N12696, N12684);
buf BUF1 (N12697, N12682);
nand NAND2 (N12698, N12687, N2039);
or OR3 (N12699, N12697, N4899, N12530);
buf BUF1 (N12700, N12695);
xor XOR2 (N12701, N12694, N7387);
nor NOR4 (N12702, N12693, N11457, N9314, N4839);
nand NAND2 (N12703, N12700, N11286);
or OR3 (N12704, N12698, N11747, N9421);
nand NAND3 (N12705, N12689, N8681, N9069);
nand NAND4 (N12706, N12690, N9885, N1011, N7501);
or OR4 (N12707, N12702, N4508, N7026, N9160);
and AND2 (N12708, N12696, N1187);
nand NAND4 (N12709, N12706, N5392, N9402, N6016);
or OR2 (N12710, N12708, N8458);
buf BUF1 (N12711, N12699);
nand NAND2 (N12712, N12675, N5660);
nand NAND4 (N12713, N12710, N926, N230, N12597);
buf BUF1 (N12714, N12705);
not NOT1 (N12715, N12712);
buf BUF1 (N12716, N12701);
buf BUF1 (N12717, N12709);
and AND2 (N12718, N12713, N4759);
or OR2 (N12719, N12711, N11068);
nor NOR2 (N12720, N12715, N11789);
buf BUF1 (N12721, N12704);
xor XOR2 (N12722, N12657, N1237);
and AND3 (N12723, N12716, N2452, N2084);
nand NAND3 (N12724, N12720, N7014, N1357);
buf BUF1 (N12725, N12707);
and AND3 (N12726, N12703, N11898, N3390);
nor NOR4 (N12727, N12714, N3296, N9850, N1914);
nand NAND4 (N12728, N12722, N3168, N6064, N7989);
xor XOR2 (N12729, N12724, N7836);
nor NOR3 (N12730, N12728, N5858, N1743);
not NOT1 (N12731, N12729);
or OR2 (N12732, N12719, N5940);
or OR4 (N12733, N12723, N6430, N12170, N3382);
buf BUF1 (N12734, N12733);
or OR4 (N12735, N12721, N12465, N3255, N11402);
and AND3 (N12736, N12718, N8262, N6324);
nand NAND4 (N12737, N12727, N3017, N11133, N3272);
nand NAND2 (N12738, N12725, N6000);
not NOT1 (N12739, N12738);
not NOT1 (N12740, N12736);
xor XOR2 (N12741, N12740, N10705);
xor XOR2 (N12742, N12732, N6515);
buf BUF1 (N12743, N12739);
or OR4 (N12744, N12742, N3300, N7381, N10856);
and AND3 (N12745, N12731, N5577, N8320);
buf BUF1 (N12746, N12737);
xor XOR2 (N12747, N12744, N12681);
or OR3 (N12748, N12734, N9838, N6520);
or OR2 (N12749, N12745, N11980);
xor XOR2 (N12750, N12746, N10925);
and AND2 (N12751, N12743, N8642);
xor XOR2 (N12752, N12748, N10558);
nor NOR2 (N12753, N12735, N12194);
xor XOR2 (N12754, N12747, N11233);
not NOT1 (N12755, N12726);
xor XOR2 (N12756, N12755, N6442);
xor XOR2 (N12757, N12751, N1492);
not NOT1 (N12758, N12741);
xor XOR2 (N12759, N12758, N2479);
not NOT1 (N12760, N12717);
nand NAND3 (N12761, N12750, N8611, N10063);
or OR4 (N12762, N12760, N11295, N4929, N9011);
nor NOR2 (N12763, N12753, N1982);
xor XOR2 (N12764, N12759, N6964);
buf BUF1 (N12765, N12754);
not NOT1 (N12766, N12752);
buf BUF1 (N12767, N12763);
nor NOR3 (N12768, N12756, N12610, N9798);
nand NAND3 (N12769, N12757, N3398, N11308);
not NOT1 (N12770, N12749);
and AND4 (N12771, N12768, N3236, N1629, N4339);
nor NOR4 (N12772, N12770, N9731, N2363, N1925);
buf BUF1 (N12773, N12769);
xor XOR2 (N12774, N12772, N4350);
or OR4 (N12775, N12730, N5839, N9475, N3948);
and AND3 (N12776, N12764, N3241, N7049);
or OR3 (N12777, N12771, N9927, N10605);
nand NAND2 (N12778, N12762, N8936);
nand NAND3 (N12779, N12766, N12110, N12150);
not NOT1 (N12780, N12774);
not NOT1 (N12781, N12761);
and AND2 (N12782, N12773, N3773);
nand NAND4 (N12783, N12775, N7393, N9786, N927);
not NOT1 (N12784, N12783);
buf BUF1 (N12785, N12765);
nand NAND3 (N12786, N12780, N8370, N1638);
not NOT1 (N12787, N12778);
buf BUF1 (N12788, N12779);
buf BUF1 (N12789, N12786);
xor XOR2 (N12790, N12789, N12739);
nand NAND3 (N12791, N12790, N8039, N6083);
or OR3 (N12792, N12784, N6149, N128);
not NOT1 (N12793, N12791);
buf BUF1 (N12794, N12782);
nand NAND2 (N12795, N12767, N919);
and AND4 (N12796, N12776, N1563, N9486, N4560);
nor NOR4 (N12797, N12785, N5055, N3, N6866);
not NOT1 (N12798, N12793);
nor NOR3 (N12799, N12797, N4968, N4975);
or OR2 (N12800, N12781, N3260);
xor XOR2 (N12801, N12777, N11730);
or OR2 (N12802, N12800, N4579);
buf BUF1 (N12803, N12796);
nand NAND4 (N12804, N12787, N2527, N8443, N1619);
nand NAND2 (N12805, N12802, N9858);
nand NAND2 (N12806, N12788, N4835);
nor NOR4 (N12807, N12801, N856, N12623, N9624);
and AND3 (N12808, N12799, N649, N1508);
and AND3 (N12809, N12805, N8490, N1989);
not NOT1 (N12810, N12803);
xor XOR2 (N12811, N12808, N1370);
not NOT1 (N12812, N12804);
or OR3 (N12813, N12806, N1823, N12204);
buf BUF1 (N12814, N12809);
nand NAND3 (N12815, N12794, N9343, N12061);
and AND2 (N12816, N12807, N6686);
nor NOR3 (N12817, N12811, N10384, N8378);
nor NOR2 (N12818, N12815, N3701);
not NOT1 (N12819, N12798);
nand NAND2 (N12820, N12795, N11692);
nor NOR2 (N12821, N12818, N12745);
nand NAND4 (N12822, N12816, N1668, N832, N9772);
not NOT1 (N12823, N12814);
nor NOR2 (N12824, N12820, N4885);
or OR2 (N12825, N12810, N646);
buf BUF1 (N12826, N12792);
nor NOR4 (N12827, N12822, N9212, N10989, N5234);
xor XOR2 (N12828, N12827, N10013);
xor XOR2 (N12829, N12826, N4190);
nand NAND2 (N12830, N12823, N8606);
nand NAND4 (N12831, N12829, N11613, N129, N1502);
or OR4 (N12832, N12817, N7210, N11751, N10164);
or OR4 (N12833, N12825, N12110, N12376, N11456);
and AND3 (N12834, N12830, N5809, N7977);
nand NAND3 (N12835, N12813, N11564, N2691);
and AND3 (N12836, N12821, N8245, N4212);
not NOT1 (N12837, N12836);
nand NAND4 (N12838, N12831, N1578, N2602, N12267);
and AND3 (N12839, N12832, N6166, N9324);
buf BUF1 (N12840, N12838);
or OR2 (N12841, N12840, N11244);
and AND2 (N12842, N12839, N9509);
not NOT1 (N12843, N12833);
xor XOR2 (N12844, N12837, N2358);
or OR4 (N12845, N12812, N10170, N11330, N9102);
nand NAND3 (N12846, N12835, N11424, N12401);
nand NAND2 (N12847, N12843, N3875);
buf BUF1 (N12848, N12842);
nand NAND2 (N12849, N12847, N6695);
not NOT1 (N12850, N12824);
nand NAND4 (N12851, N12841, N955, N9334, N7313);
not NOT1 (N12852, N12846);
and AND2 (N12853, N12852, N2858);
nor NOR4 (N12854, N12849, N8980, N6219, N9068);
xor XOR2 (N12855, N12834, N4841);
and AND3 (N12856, N12851, N12523, N6948);
or OR4 (N12857, N12844, N531, N10674, N4686);
nand NAND3 (N12858, N12856, N1214, N10784);
not NOT1 (N12859, N12850);
xor XOR2 (N12860, N12855, N5783);
and AND2 (N12861, N12858, N4496);
and AND3 (N12862, N12828, N7335, N6719);
xor XOR2 (N12863, N12819, N10625);
not NOT1 (N12864, N12853);
nand NAND3 (N12865, N12861, N9571, N9666);
buf BUF1 (N12866, N12860);
and AND3 (N12867, N12864, N5105, N3841);
xor XOR2 (N12868, N12866, N10819);
buf BUF1 (N12869, N12859);
nand NAND4 (N12870, N12854, N9592, N2080, N4915);
or OR2 (N12871, N12845, N4242);
nor NOR2 (N12872, N12870, N4436);
and AND2 (N12873, N12868, N1153);
or OR4 (N12874, N12867, N2124, N1140, N3001);
xor XOR2 (N12875, N12874, N10584);
not NOT1 (N12876, N12863);
or OR4 (N12877, N12862, N3493, N10000, N11389);
or OR4 (N12878, N12875, N12815, N10637, N10512);
buf BUF1 (N12879, N12878);
buf BUF1 (N12880, N12865);
or OR2 (N12881, N12848, N6128);
not NOT1 (N12882, N12876);
buf BUF1 (N12883, N12879);
or OR3 (N12884, N12882, N3803, N2143);
and AND4 (N12885, N12872, N474, N9971, N7057);
or OR3 (N12886, N12873, N2017, N3565);
nor NOR4 (N12887, N12869, N1292, N11643, N10208);
nand NAND4 (N12888, N12884, N1414, N4516, N4462);
or OR3 (N12889, N12877, N11898, N5859);
xor XOR2 (N12890, N12888, N4587);
and AND4 (N12891, N12890, N3691, N8890, N7683);
or OR3 (N12892, N12883, N5248, N602);
nand NAND4 (N12893, N12891, N2185, N11451, N7972);
not NOT1 (N12894, N12880);
nor NOR3 (N12895, N12886, N6876, N5108);
buf BUF1 (N12896, N12892);
nand NAND2 (N12897, N12871, N10309);
nor NOR2 (N12898, N12857, N2965);
nor NOR2 (N12899, N12896, N4688);
nor NOR3 (N12900, N12881, N8690, N1739);
buf BUF1 (N12901, N12899);
and AND4 (N12902, N12893, N11533, N2136, N8346);
buf BUF1 (N12903, N12889);
and AND4 (N12904, N12894, N12635, N10329, N4914);
or OR2 (N12905, N12902, N1390);
nand NAND2 (N12906, N12898, N2654);
nor NOR4 (N12907, N12901, N9450, N2984, N6247);
xor XOR2 (N12908, N12906, N5704);
and AND3 (N12909, N12897, N1595, N3431);
or OR4 (N12910, N12895, N12767, N2387, N10755);
nor NOR4 (N12911, N12887, N4794, N672, N8087);
xor XOR2 (N12912, N12905, N5395);
or OR4 (N12913, N12907, N3287, N10247, N8963);
nand NAND2 (N12914, N12908, N5305);
not NOT1 (N12915, N12911);
not NOT1 (N12916, N12915);
nor NOR3 (N12917, N12910, N6860, N11343);
or OR4 (N12918, N12900, N3744, N4612, N11208);
nor NOR3 (N12919, N12904, N8893, N198);
nand NAND3 (N12920, N12918, N1756, N11310);
not NOT1 (N12921, N12919);
nor NOR4 (N12922, N12916, N4822, N10014, N7343);
xor XOR2 (N12923, N12917, N251);
and AND3 (N12924, N12914, N1330, N4105);
xor XOR2 (N12925, N12923, N8305);
buf BUF1 (N12926, N12913);
and AND4 (N12927, N12924, N8492, N4620, N7609);
buf BUF1 (N12928, N12885);
and AND2 (N12929, N12921, N7444);
xor XOR2 (N12930, N12903, N9157);
nand NAND3 (N12931, N12927, N4490, N12886);
or OR2 (N12932, N12912, N9742);
xor XOR2 (N12933, N12920, N2374);
not NOT1 (N12934, N12930);
buf BUF1 (N12935, N12928);
nand NAND2 (N12936, N12932, N7048);
xor XOR2 (N12937, N12909, N5476);
nand NAND3 (N12938, N12931, N8544, N1991);
nand NAND3 (N12939, N12925, N3343, N10032);
nor NOR3 (N12940, N12933, N4274, N5470);
xor XOR2 (N12941, N12938, N11633);
buf BUF1 (N12942, N12934);
not NOT1 (N12943, N12936);
not NOT1 (N12944, N12940);
and AND3 (N12945, N12944, N2562, N12537);
or OR3 (N12946, N12926, N11185, N12663);
nand NAND2 (N12947, N12937, N3904);
and AND3 (N12948, N12947, N10424, N2483);
xor XOR2 (N12949, N12945, N5835);
and AND4 (N12950, N12946, N3999, N10019, N6644);
buf BUF1 (N12951, N12948);
buf BUF1 (N12952, N12929);
and AND3 (N12953, N12950, N4744, N5651);
not NOT1 (N12954, N12941);
not NOT1 (N12955, N12951);
nor NOR2 (N12956, N12922, N1202);
and AND3 (N12957, N12952, N10784, N6926);
nor NOR4 (N12958, N12935, N11229, N6419, N10953);
not NOT1 (N12959, N12954);
xor XOR2 (N12960, N12955, N6118);
nor NOR3 (N12961, N12949, N7086, N3997);
or OR2 (N12962, N12958, N9727);
nand NAND3 (N12963, N12953, N12587, N8353);
xor XOR2 (N12964, N12956, N11195);
not NOT1 (N12965, N12939);
and AND2 (N12966, N12961, N6149);
xor XOR2 (N12967, N12962, N2411);
nand NAND4 (N12968, N12965, N7376, N6131, N11371);
or OR3 (N12969, N12963, N10456, N6264);
or OR3 (N12970, N12969, N7190, N8416);
not NOT1 (N12971, N12967);
not NOT1 (N12972, N12968);
nor NOR2 (N12973, N12966, N182);
nor NOR2 (N12974, N12957, N3645);
or OR3 (N12975, N12942, N3632, N404);
and AND4 (N12976, N12972, N492, N12164, N322);
nand NAND2 (N12977, N12975, N9153);
xor XOR2 (N12978, N12976, N12227);
xor XOR2 (N12979, N12971, N3047);
nand NAND3 (N12980, N12973, N485, N12179);
nand NAND3 (N12981, N12964, N2902, N7736);
nor NOR2 (N12982, N12981, N8843);
and AND2 (N12983, N12978, N12224);
nor NOR2 (N12984, N12943, N853);
buf BUF1 (N12985, N12959);
or OR3 (N12986, N12979, N1267, N8583);
or OR2 (N12987, N12977, N12280);
not NOT1 (N12988, N12970);
and AND2 (N12989, N12960, N3781);
buf BUF1 (N12990, N12974);
and AND4 (N12991, N12982, N8059, N258, N8680);
and AND2 (N12992, N12980, N3148);
not NOT1 (N12993, N12992);
xor XOR2 (N12994, N12985, N5534);
not NOT1 (N12995, N12988);
nor NOR2 (N12996, N12986, N5566);
not NOT1 (N12997, N12994);
and AND2 (N12998, N12996, N660);
nand NAND2 (N12999, N12989, N8265);
xor XOR2 (N13000, N12990, N9142);
nand NAND4 (N13001, N12987, N7257, N8259, N2419);
not NOT1 (N13002, N12991);
and AND3 (N13003, N12999, N4062, N1962);
buf BUF1 (N13004, N13002);
xor XOR2 (N13005, N12995, N10130);
buf BUF1 (N13006, N13000);
nor NOR4 (N13007, N12997, N5218, N11728, N9996);
or OR3 (N13008, N13001, N9699, N4692);
nor NOR4 (N13009, N13004, N10, N12775, N9879);
nand NAND4 (N13010, N12998, N872, N12676, N7366);
nor NOR3 (N13011, N13006, N4994, N6888);
or OR3 (N13012, N12984, N3754, N1195);
xor XOR2 (N13013, N13007, N10192);
not NOT1 (N13014, N13005);
xor XOR2 (N13015, N13010, N8314);
or OR2 (N13016, N13013, N8180);
xor XOR2 (N13017, N13012, N10271);
xor XOR2 (N13018, N13014, N5664);
nor NOR2 (N13019, N13018, N3421);
nor NOR3 (N13020, N13008, N1125, N10681);
and AND3 (N13021, N13009, N4776, N12660);
nor NOR4 (N13022, N13015, N6422, N9249, N11024);
and AND2 (N13023, N12993, N12050);
nor NOR2 (N13024, N12983, N5191);
buf BUF1 (N13025, N13019);
not NOT1 (N13026, N13020);
nand NAND2 (N13027, N13003, N2764);
or OR3 (N13028, N13016, N3152, N413);
not NOT1 (N13029, N13017);
and AND3 (N13030, N13021, N8520, N3888);
xor XOR2 (N13031, N13028, N7445);
buf BUF1 (N13032, N13027);
or OR4 (N13033, N13011, N1660, N2444, N11307);
nor NOR3 (N13034, N13024, N4303, N8342);
nor NOR4 (N13035, N13030, N1066, N8196, N12031);
buf BUF1 (N13036, N13035);
not NOT1 (N13037, N13032);
or OR3 (N13038, N13029, N9412, N7691);
xor XOR2 (N13039, N13031, N298);
xor XOR2 (N13040, N13023, N5236);
xor XOR2 (N13041, N13034, N1182);
buf BUF1 (N13042, N13039);
xor XOR2 (N13043, N13040, N12420);
nand NAND3 (N13044, N13038, N9418, N8033);
nor NOR4 (N13045, N13044, N590, N4596, N342);
buf BUF1 (N13046, N13041);
not NOT1 (N13047, N13025);
nor NOR2 (N13048, N13046, N8773);
xor XOR2 (N13049, N13022, N5091);
not NOT1 (N13050, N13047);
nand NAND3 (N13051, N13033, N10956, N1013);
or OR3 (N13052, N13026, N4823, N3894);
buf BUF1 (N13053, N13049);
xor XOR2 (N13054, N13036, N2002);
buf BUF1 (N13055, N13042);
and AND2 (N13056, N13055, N11942);
buf BUF1 (N13057, N13050);
buf BUF1 (N13058, N13037);
buf BUF1 (N13059, N13053);
or OR3 (N13060, N13048, N10975, N12168);
or OR4 (N13061, N13060, N9196, N6663, N1623);
nand NAND3 (N13062, N13051, N3378, N5825);
and AND2 (N13063, N13062, N9982);
not NOT1 (N13064, N13052);
nand NAND4 (N13065, N13061, N2342, N1256, N7391);
or OR3 (N13066, N13054, N12221, N11348);
or OR4 (N13067, N13056, N3565, N9158, N10729);
or OR4 (N13068, N13059, N8686, N11728, N3855);
buf BUF1 (N13069, N13065);
and AND3 (N13070, N13057, N11439, N6922);
not NOT1 (N13071, N13069);
xor XOR2 (N13072, N13064, N1594);
xor XOR2 (N13073, N13045, N10664);
or OR3 (N13074, N13058, N9635, N5253);
or OR4 (N13075, N13073, N2899, N6327, N9770);
nand NAND2 (N13076, N13071, N11711);
nand NAND3 (N13077, N13070, N9367, N3264);
nand NAND3 (N13078, N13063, N9157, N5469);
nand NAND3 (N13079, N13067, N2260, N4009);
or OR3 (N13080, N13072, N1293, N2360);
nand NAND2 (N13081, N13075, N5273);
not NOT1 (N13082, N13043);
buf BUF1 (N13083, N13068);
nand NAND3 (N13084, N13076, N1759, N2342);
nand NAND2 (N13085, N13077, N10014);
not NOT1 (N13086, N13084);
nand NAND4 (N13087, N13085, N3688, N3902, N21);
not NOT1 (N13088, N13081);
or OR4 (N13089, N13074, N3991, N9012, N9891);
nor NOR3 (N13090, N13089, N6785, N12340);
nand NAND4 (N13091, N13090, N4221, N2766, N4912);
nor NOR4 (N13092, N13083, N6430, N9265, N7699);
not NOT1 (N13093, N13080);
and AND2 (N13094, N13093, N12486);
and AND4 (N13095, N13066, N12495, N10951, N11658);
not NOT1 (N13096, N13092);
buf BUF1 (N13097, N13091);
and AND4 (N13098, N13096, N12521, N8878, N4972);
or OR3 (N13099, N13094, N162, N6112);
xor XOR2 (N13100, N13078, N5277);
or OR4 (N13101, N13095, N6273, N4463, N6766);
buf BUF1 (N13102, N13099);
nand NAND4 (N13103, N13082, N1146, N1928, N8542);
xor XOR2 (N13104, N13087, N963);
not NOT1 (N13105, N13079);
nand NAND3 (N13106, N13100, N12653, N8469);
and AND3 (N13107, N13086, N121, N4504);
buf BUF1 (N13108, N13103);
nor NOR4 (N13109, N13088, N10827, N9819, N4425);
and AND2 (N13110, N13097, N2543);
not NOT1 (N13111, N13108);
buf BUF1 (N13112, N13098);
nand NAND4 (N13113, N13106, N868, N12220, N197);
xor XOR2 (N13114, N13104, N2302);
nor NOR3 (N13115, N13107, N12982, N6654);
nand NAND4 (N13116, N13113, N7230, N290, N8325);
nor NOR2 (N13117, N13115, N1485);
xor XOR2 (N13118, N13112, N10966);
xor XOR2 (N13119, N13118, N7718);
or OR4 (N13120, N13116, N4057, N7293, N9373);
nand NAND4 (N13121, N13120, N4072, N11031, N3621);
and AND2 (N13122, N13109, N5901);
nand NAND2 (N13123, N13122, N6808);
and AND3 (N13124, N13102, N6557, N1443);
or OR2 (N13125, N13114, N4704);
buf BUF1 (N13126, N13117);
xor XOR2 (N13127, N13125, N1277);
nand NAND3 (N13128, N13111, N9022, N3705);
nand NAND2 (N13129, N13123, N12324);
nor NOR3 (N13130, N13124, N4218, N1501);
and AND3 (N13131, N13126, N3773, N12678);
buf BUF1 (N13132, N13119);
or OR4 (N13133, N13101, N7770, N5211, N669);
buf BUF1 (N13134, N13129);
nand NAND4 (N13135, N13110, N11898, N925, N3594);
nor NOR3 (N13136, N13131, N11987, N1737);
nor NOR4 (N13137, N13130, N10582, N4357, N5758);
xor XOR2 (N13138, N13136, N2811);
nor NOR3 (N13139, N13134, N12161, N12775);
buf BUF1 (N13140, N13138);
not NOT1 (N13141, N13105);
xor XOR2 (N13142, N13133, N11475);
and AND2 (N13143, N13121, N12106);
xor XOR2 (N13144, N13141, N4946);
buf BUF1 (N13145, N13135);
xor XOR2 (N13146, N13145, N9879);
not NOT1 (N13147, N13128);
not NOT1 (N13148, N13143);
not NOT1 (N13149, N13132);
xor XOR2 (N13150, N13139, N6607);
not NOT1 (N13151, N13148);
nand NAND2 (N13152, N13144, N5520);
xor XOR2 (N13153, N13127, N12367);
nor NOR2 (N13154, N13150, N621);
buf BUF1 (N13155, N13146);
nand NAND3 (N13156, N13152, N8815, N12272);
nor NOR4 (N13157, N13140, N10942, N5876, N3895);
not NOT1 (N13158, N13153);
nor NOR3 (N13159, N13156, N2764, N8252);
xor XOR2 (N13160, N13159, N6266);
buf BUF1 (N13161, N13157);
xor XOR2 (N13162, N13158, N4174);
or OR4 (N13163, N13154, N12850, N1388, N3162);
nand NAND3 (N13164, N13142, N711, N281);
not NOT1 (N13165, N13151);
and AND2 (N13166, N13155, N4570);
not NOT1 (N13167, N13164);
and AND4 (N13168, N13149, N4750, N8580, N12602);
and AND4 (N13169, N13166, N6514, N856, N5359);
not NOT1 (N13170, N13167);
nor NOR4 (N13171, N13162, N2956, N9911, N4081);
xor XOR2 (N13172, N13160, N7649);
or OR3 (N13173, N13137, N1444, N11351);
xor XOR2 (N13174, N13161, N1006);
nor NOR3 (N13175, N13147, N8269, N4625);
xor XOR2 (N13176, N13169, N2523);
nand NAND3 (N13177, N13171, N5509, N5455);
or OR4 (N13178, N13173, N6557, N1047, N2387);
xor XOR2 (N13179, N13176, N1282);
and AND4 (N13180, N13163, N3429, N29, N5565);
xor XOR2 (N13181, N13180, N12467);
or OR4 (N13182, N13174, N11515, N10335, N6623);
nor NOR4 (N13183, N13168, N4899, N3587, N9456);
nand NAND4 (N13184, N13172, N3447, N12619, N7817);
buf BUF1 (N13185, N13184);
xor XOR2 (N13186, N13183, N10376);
nand NAND4 (N13187, N13175, N8729, N12216, N9049);
and AND3 (N13188, N13185, N4886, N10907);
nor NOR2 (N13189, N13177, N2792);
buf BUF1 (N13190, N13188);
not NOT1 (N13191, N13165);
nand NAND2 (N13192, N13187, N5382);
or OR3 (N13193, N13170, N8110, N12348);
nor NOR2 (N13194, N13190, N12967);
not NOT1 (N13195, N13181);
xor XOR2 (N13196, N13194, N13028);
nor NOR2 (N13197, N13195, N4268);
nand NAND2 (N13198, N13191, N1563);
and AND4 (N13199, N13186, N4147, N7807, N10874);
xor XOR2 (N13200, N13193, N9194);
xor XOR2 (N13201, N13199, N9031);
nand NAND2 (N13202, N13179, N13039);
and AND4 (N13203, N13189, N12994, N3145, N7664);
nand NAND4 (N13204, N13197, N6077, N10649, N3203);
not NOT1 (N13205, N13178);
and AND2 (N13206, N13196, N8686);
buf BUF1 (N13207, N13205);
or OR2 (N13208, N13203, N12919);
xor XOR2 (N13209, N13207, N2228);
or OR4 (N13210, N13209, N7042, N11010, N2274);
nand NAND4 (N13211, N13200, N1229, N5624, N5535);
or OR2 (N13212, N13211, N7510);
and AND3 (N13213, N13206, N10416, N9438);
buf BUF1 (N13214, N13208);
or OR4 (N13215, N13202, N6078, N11548, N4915);
and AND4 (N13216, N13212, N7433, N3669, N2641);
and AND4 (N13217, N13198, N2465, N12905, N10952);
nand NAND4 (N13218, N13214, N3168, N7453, N8651);
not NOT1 (N13219, N13217);
buf BUF1 (N13220, N13213);
nor NOR4 (N13221, N13218, N10401, N12577, N8549);
or OR2 (N13222, N13192, N4458);
and AND2 (N13223, N13221, N2365);
and AND4 (N13224, N13220, N6021, N3857, N7802);
nand NAND2 (N13225, N13210, N3653);
buf BUF1 (N13226, N13224);
or OR4 (N13227, N13226, N12209, N11871, N10465);
not NOT1 (N13228, N13182);
and AND2 (N13229, N13219, N10581);
not NOT1 (N13230, N13227);
nand NAND4 (N13231, N13228, N10873, N1386, N4036);
buf BUF1 (N13232, N13230);
not NOT1 (N13233, N13204);
and AND4 (N13234, N13233, N6120, N9772, N12125);
nor NOR2 (N13235, N13229, N8105);
not NOT1 (N13236, N13232);
nor NOR4 (N13237, N13215, N3736, N4068, N12871);
not NOT1 (N13238, N13201);
not NOT1 (N13239, N13216);
not NOT1 (N13240, N13237);
nand NAND2 (N13241, N13231, N11545);
xor XOR2 (N13242, N13241, N2702);
buf BUF1 (N13243, N13225);
and AND3 (N13244, N13242, N3455, N12540);
buf BUF1 (N13245, N13243);
or OR4 (N13246, N13239, N8514, N765, N5938);
xor XOR2 (N13247, N13245, N11964);
buf BUF1 (N13248, N13234);
buf BUF1 (N13249, N13246);
nand NAND4 (N13250, N13244, N2530, N2619, N6288);
nor NOR3 (N13251, N13238, N11649, N9350);
buf BUF1 (N13252, N13223);
or OR4 (N13253, N13251, N7160, N7255, N11158);
buf BUF1 (N13254, N13240);
nand NAND2 (N13255, N13236, N12115);
and AND3 (N13256, N13249, N7602, N8638);
xor XOR2 (N13257, N13252, N7999);
buf BUF1 (N13258, N13248);
nor NOR2 (N13259, N13250, N562);
or OR2 (N13260, N13235, N1649);
or OR3 (N13261, N13253, N5277, N8616);
or OR3 (N13262, N13254, N12822, N4574);
buf BUF1 (N13263, N13257);
or OR4 (N13264, N13247, N11483, N4044, N13159);
nand NAND3 (N13265, N13222, N2970, N10297);
nor NOR2 (N13266, N13265, N12097);
and AND4 (N13267, N13255, N1102, N8956, N4818);
nor NOR4 (N13268, N13258, N4512, N2450, N12757);
nor NOR3 (N13269, N13263, N3797, N226);
buf BUF1 (N13270, N13268);
nor NOR3 (N13271, N13256, N11655, N12510);
buf BUF1 (N13272, N13270);
nand NAND2 (N13273, N13259, N2885);
not NOT1 (N13274, N13272);
nor NOR2 (N13275, N13274, N12887);
xor XOR2 (N13276, N13264, N10386);
xor XOR2 (N13277, N13269, N11641);
or OR3 (N13278, N13271, N8565, N11739);
nand NAND2 (N13279, N13273, N7351);
xor XOR2 (N13280, N13279, N3866);
nor NOR2 (N13281, N13262, N13260);
buf BUF1 (N13282, N7809);
and AND2 (N13283, N13267, N4797);
buf BUF1 (N13284, N13280);
nand NAND2 (N13285, N13284, N4564);
buf BUF1 (N13286, N13275);
nor NOR4 (N13287, N13281, N3362, N12271, N8372);
and AND2 (N13288, N13261, N9589);
xor XOR2 (N13289, N13277, N711);
nor NOR2 (N13290, N13283, N1182);
nand NAND2 (N13291, N13278, N7997);
xor XOR2 (N13292, N13290, N4334);
not NOT1 (N13293, N13282);
and AND4 (N13294, N13289, N12570, N6433, N4672);
or OR3 (N13295, N13294, N688, N4203);
nand NAND4 (N13296, N13285, N8575, N3663, N7180);
nor NOR4 (N13297, N13292, N8165, N2584, N4615);
nand NAND4 (N13298, N13297, N423, N2681, N1781);
buf BUF1 (N13299, N13291);
nor NOR2 (N13300, N13266, N13259);
nand NAND2 (N13301, N13276, N4530);
and AND4 (N13302, N13293, N4524, N7680, N4453);
not NOT1 (N13303, N13295);
xor XOR2 (N13304, N13296, N13041);
nor NOR3 (N13305, N13298, N9293, N9420);
nand NAND3 (N13306, N13301, N11152, N12314);
nand NAND4 (N13307, N13302, N11365, N5572, N4840);
not NOT1 (N13308, N13300);
nor NOR2 (N13309, N13287, N6495);
not NOT1 (N13310, N13306);
or OR3 (N13311, N13307, N6247, N4387);
nand NAND2 (N13312, N13304, N10192);
nand NAND3 (N13313, N13305, N4183, N2992);
nand NAND3 (N13314, N13286, N9778, N952);
xor XOR2 (N13315, N13288, N9019);
and AND2 (N13316, N13315, N7852);
nand NAND3 (N13317, N13311, N4374, N3033);
nor NOR3 (N13318, N13303, N7611, N12828);
nor NOR4 (N13319, N13309, N9880, N7937, N9555);
buf BUF1 (N13320, N13312);
and AND4 (N13321, N13318, N1418, N11051, N13150);
xor XOR2 (N13322, N13319, N1822);
xor XOR2 (N13323, N13316, N11052);
nor NOR4 (N13324, N13299, N3290, N7140, N4083);
or OR3 (N13325, N13313, N190, N9004);
nor NOR2 (N13326, N13321, N5013);
and AND2 (N13327, N13310, N8180);
xor XOR2 (N13328, N13327, N6444);
buf BUF1 (N13329, N13324);
nor NOR4 (N13330, N13308, N6664, N12591, N12702);
not NOT1 (N13331, N13329);
xor XOR2 (N13332, N13331, N12994);
nor NOR2 (N13333, N13328, N9418);
or OR3 (N13334, N13317, N8064, N203);
nand NAND3 (N13335, N13323, N2872, N4359);
nor NOR4 (N13336, N13325, N2068, N9264, N1958);
buf BUF1 (N13337, N13336);
nor NOR4 (N13338, N13333, N1193, N8236, N3304);
buf BUF1 (N13339, N13335);
not NOT1 (N13340, N13332);
not NOT1 (N13341, N13340);
not NOT1 (N13342, N13339);
or OR3 (N13343, N13338, N380, N8238);
xor XOR2 (N13344, N13342, N12586);
or OR3 (N13345, N13322, N3669, N6957);
not NOT1 (N13346, N13341);
and AND4 (N13347, N13326, N9135, N6029, N3632);
or OR4 (N13348, N13347, N9842, N1477, N1327);
nor NOR3 (N13349, N13346, N10836, N6550);
nor NOR3 (N13350, N13314, N2269, N8867);
nor NOR3 (N13351, N13337, N11019, N2017);
nor NOR2 (N13352, N13351, N11352);
nor NOR4 (N13353, N13330, N5340, N4614, N3469);
buf BUF1 (N13354, N13320);
nor NOR4 (N13355, N13354, N11382, N5248, N182);
nor NOR4 (N13356, N13345, N6574, N12104, N12973);
and AND4 (N13357, N13343, N8094, N2183, N7741);
or OR3 (N13358, N13334, N923, N12836);
nand NAND2 (N13359, N13356, N9115);
xor XOR2 (N13360, N13357, N11140);
not NOT1 (N13361, N13352);
nand NAND4 (N13362, N13344, N12670, N1734, N6482);
nor NOR3 (N13363, N13358, N3591, N3479);
buf BUF1 (N13364, N13359);
or OR2 (N13365, N13361, N11753);
and AND3 (N13366, N13365, N6816, N7501);
xor XOR2 (N13367, N13353, N3937);
nor NOR3 (N13368, N13362, N7637, N9018);
buf BUF1 (N13369, N13368);
nor NOR3 (N13370, N13364, N4989, N12919);
and AND2 (N13371, N13355, N8742);
buf BUF1 (N13372, N13370);
and AND4 (N13373, N13371, N199, N1921, N4030);
xor XOR2 (N13374, N13348, N12669);
buf BUF1 (N13375, N13350);
and AND4 (N13376, N13373, N128, N7961, N556);
not NOT1 (N13377, N13376);
not NOT1 (N13378, N13363);
or OR3 (N13379, N13372, N274, N4845);
buf BUF1 (N13380, N13360);
buf BUF1 (N13381, N13380);
xor XOR2 (N13382, N13378, N1536);
nand NAND3 (N13383, N13349, N5656, N10342);
nand NAND2 (N13384, N13377, N9547);
or OR4 (N13385, N13384, N3055, N1335, N11458);
or OR4 (N13386, N13367, N10048, N6823, N8662);
nand NAND4 (N13387, N13385, N4016, N10643, N8663);
and AND2 (N13388, N13386, N4988);
or OR3 (N13389, N13375, N5736, N8923);
or OR3 (N13390, N13389, N1610, N9942);
xor XOR2 (N13391, N13379, N2344);
buf BUF1 (N13392, N13382);
not NOT1 (N13393, N13369);
or OR2 (N13394, N13387, N11845);
and AND3 (N13395, N13388, N12141, N9406);
nand NAND2 (N13396, N13395, N10868);
nor NOR3 (N13397, N13374, N4475, N7211);
xor XOR2 (N13398, N13394, N11724);
and AND3 (N13399, N13396, N11487, N10896);
nand NAND3 (N13400, N13391, N3027, N8064);
buf BUF1 (N13401, N13366);
or OR3 (N13402, N13393, N7701, N7852);
nor NOR2 (N13403, N13401, N8739);
nor NOR4 (N13404, N13403, N5054, N1726, N3256);
or OR2 (N13405, N13397, N11686);
buf BUF1 (N13406, N13399);
buf BUF1 (N13407, N13404);
xor XOR2 (N13408, N13406, N9809);
or OR2 (N13409, N13392, N12444);
and AND2 (N13410, N13383, N6077);
nand NAND4 (N13411, N13405, N7342, N12184, N6218);
xor XOR2 (N13412, N13390, N6095);
and AND4 (N13413, N13409, N13230, N8947, N970);
or OR4 (N13414, N13400, N10639, N2079, N348);
nor NOR4 (N13415, N13408, N1231, N2829, N3664);
buf BUF1 (N13416, N13410);
nand NAND2 (N13417, N13414, N2434);
nor NOR4 (N13418, N13417, N11981, N1473, N9115);
nand NAND3 (N13419, N13411, N8423, N5106);
nor NOR2 (N13420, N13415, N1237);
or OR3 (N13421, N13412, N5994, N1670);
nor NOR4 (N13422, N13421, N2621, N3888, N6749);
xor XOR2 (N13423, N13402, N1134);
nand NAND4 (N13424, N13381, N129, N13123, N9980);
nor NOR4 (N13425, N13419, N1318, N3052, N1899);
or OR4 (N13426, N13413, N7061, N4322, N10813);
and AND3 (N13427, N13420, N12730, N387);
or OR4 (N13428, N13425, N13317, N9752, N5733);
not NOT1 (N13429, N13428);
or OR4 (N13430, N13416, N11203, N10127, N5592);
or OR3 (N13431, N13430, N2100, N7776);
or OR2 (N13432, N13427, N2056);
xor XOR2 (N13433, N13424, N3249);
nand NAND4 (N13434, N13418, N5646, N10051, N7238);
xor XOR2 (N13435, N13426, N6050);
xor XOR2 (N13436, N13431, N10506);
and AND4 (N13437, N13434, N2783, N7991, N12920);
not NOT1 (N13438, N13436);
nor NOR2 (N13439, N13429, N321);
and AND2 (N13440, N13438, N7738);
or OR3 (N13441, N13440, N3626, N6686);
nor NOR3 (N13442, N13435, N1519, N8816);
nand NAND2 (N13443, N13439, N395);
and AND3 (N13444, N13443, N7171, N5939);
not NOT1 (N13445, N13441);
nor NOR3 (N13446, N13423, N11249, N9860);
buf BUF1 (N13447, N13432);
or OR2 (N13448, N13422, N10087);
buf BUF1 (N13449, N13444);
and AND4 (N13450, N13437, N7970, N3420, N5591);
or OR3 (N13451, N13448, N2214, N6395);
or OR4 (N13452, N13446, N7428, N5223, N6393);
buf BUF1 (N13453, N13449);
nor NOR2 (N13454, N13398, N12180);
buf BUF1 (N13455, N13445);
or OR3 (N13456, N13451, N12364, N306);
buf BUF1 (N13457, N13452);
nand NAND2 (N13458, N13433, N5755);
xor XOR2 (N13459, N13453, N11390);
buf BUF1 (N13460, N13454);
buf BUF1 (N13461, N13455);
and AND4 (N13462, N13458, N6812, N130, N2356);
xor XOR2 (N13463, N13442, N1123);
or OR4 (N13464, N13459, N2642, N4401, N1855);
xor XOR2 (N13465, N13407, N7598);
or OR2 (N13466, N13450, N8318);
and AND3 (N13467, N13462, N6238, N8533);
and AND3 (N13468, N13465, N410, N9170);
and AND3 (N13469, N13464, N9752, N13333);
and AND4 (N13470, N13466, N6829, N7208, N1829);
or OR3 (N13471, N13463, N8267, N12767);
xor XOR2 (N13472, N13467, N4643);
xor XOR2 (N13473, N13468, N6488);
and AND4 (N13474, N13461, N10948, N13159, N11299);
or OR3 (N13475, N13460, N3349, N4595);
and AND3 (N13476, N13447, N6687, N7526);
not NOT1 (N13477, N13469);
nand NAND3 (N13478, N13470, N1619, N11606);
xor XOR2 (N13479, N13477, N11388);
or OR4 (N13480, N13473, N7868, N8963, N37);
nand NAND4 (N13481, N13475, N5437, N8756, N9553);
or OR3 (N13482, N13472, N3323, N10068);
nor NOR3 (N13483, N13482, N10780, N8816);
or OR3 (N13484, N13456, N4546, N12037);
xor XOR2 (N13485, N13483, N2072);
nor NOR2 (N13486, N13457, N1186);
or OR3 (N13487, N13471, N2856, N11323);
nor NOR2 (N13488, N13487, N5036);
or OR3 (N13489, N13480, N8621, N7596);
or OR2 (N13490, N13479, N4799);
nand NAND3 (N13491, N13484, N12518, N5457);
nor NOR2 (N13492, N13476, N730);
and AND3 (N13493, N13486, N8247, N13308);
or OR4 (N13494, N13492, N6414, N2782, N10978);
and AND4 (N13495, N13481, N737, N782, N7150);
nor NOR4 (N13496, N13485, N2919, N5916, N1509);
buf BUF1 (N13497, N13490);
not NOT1 (N13498, N13478);
and AND3 (N13499, N13488, N125, N3327);
and AND3 (N13500, N13496, N12792, N5090);
buf BUF1 (N13501, N13497);
buf BUF1 (N13502, N13489);
xor XOR2 (N13503, N13474, N6459);
and AND3 (N13504, N13501, N5279, N4821);
and AND4 (N13505, N13502, N6264, N3073, N1889);
nand NAND2 (N13506, N13493, N326);
and AND3 (N13507, N13491, N4093, N2318);
xor XOR2 (N13508, N13495, N5563);
buf BUF1 (N13509, N13494);
nor NOR3 (N13510, N13500, N719, N12274);
or OR3 (N13511, N13504, N11875, N10374);
nor NOR4 (N13512, N13509, N10967, N1208, N10788);
or OR4 (N13513, N13499, N10453, N7919, N9962);
buf BUF1 (N13514, N13507);
nor NOR4 (N13515, N13503, N4795, N8282, N2279);
buf BUF1 (N13516, N13508);
and AND2 (N13517, N13506, N7449);
buf BUF1 (N13518, N13517);
nand NAND3 (N13519, N13498, N6614, N727);
not NOT1 (N13520, N13511);
not NOT1 (N13521, N13516);
buf BUF1 (N13522, N13505);
xor XOR2 (N13523, N13522, N5369);
nor NOR2 (N13524, N13513, N6720);
buf BUF1 (N13525, N13514);
xor XOR2 (N13526, N13523, N1115);
nand NAND2 (N13527, N13515, N9202);
xor XOR2 (N13528, N13524, N11895);
buf BUF1 (N13529, N13526);
or OR3 (N13530, N13518, N255, N11549);
and AND4 (N13531, N13528, N3466, N1097, N13248);
buf BUF1 (N13532, N13525);
xor XOR2 (N13533, N13512, N5705);
and AND4 (N13534, N13520, N5181, N9776, N11171);
or OR3 (N13535, N13533, N7571, N8663);
xor XOR2 (N13536, N13521, N9212);
buf BUF1 (N13537, N13536);
buf BUF1 (N13538, N13537);
nand NAND4 (N13539, N13527, N8790, N5833, N11363);
nor NOR4 (N13540, N13530, N9704, N12640, N2859);
not NOT1 (N13541, N13539);
not NOT1 (N13542, N13510);
and AND4 (N13543, N13542, N4328, N6610, N11842);
not NOT1 (N13544, N13538);
or OR3 (N13545, N13540, N2906, N4088);
not NOT1 (N13546, N13535);
or OR3 (N13547, N13544, N3773, N11685);
buf BUF1 (N13548, N13545);
buf BUF1 (N13549, N13541);
or OR2 (N13550, N13529, N8317);
and AND3 (N13551, N13546, N4172, N5287);
and AND2 (N13552, N13519, N5122);
xor XOR2 (N13553, N13543, N932);
buf BUF1 (N13554, N13553);
xor XOR2 (N13555, N13531, N3142);
nor NOR4 (N13556, N13532, N11976, N5944, N6503);
not NOT1 (N13557, N13556);
nor NOR3 (N13558, N13548, N8230, N9240);
xor XOR2 (N13559, N13555, N11497);
and AND4 (N13560, N13534, N7100, N1762, N13419);
xor XOR2 (N13561, N13560, N10777);
nor NOR4 (N13562, N13552, N12882, N1703, N4182);
buf BUF1 (N13563, N13559);
nor NOR3 (N13564, N13547, N5661, N11971);
or OR2 (N13565, N13562, N1230);
nor NOR2 (N13566, N13550, N577);
xor XOR2 (N13567, N13554, N2611);
nand NAND2 (N13568, N13565, N11090);
or OR2 (N13569, N13561, N1030);
buf BUF1 (N13570, N13567);
buf BUF1 (N13571, N13557);
not NOT1 (N13572, N13563);
and AND3 (N13573, N13570, N7423, N2950);
buf BUF1 (N13574, N13572);
xor XOR2 (N13575, N13569, N3423);
and AND3 (N13576, N13574, N5849, N10125);
nor NOR3 (N13577, N13568, N1822, N5284);
buf BUF1 (N13578, N13551);
nor NOR3 (N13579, N13566, N2871, N8819);
xor XOR2 (N13580, N13577, N9274);
nor NOR2 (N13581, N13564, N2385);
not NOT1 (N13582, N13581);
nand NAND4 (N13583, N13573, N3418, N2137, N10100);
nand NAND3 (N13584, N13582, N2613, N5592);
not NOT1 (N13585, N13558);
buf BUF1 (N13586, N13579);
and AND2 (N13587, N13549, N10515);
nor NOR4 (N13588, N13571, N6037, N13042, N2337);
nand NAND2 (N13589, N13584, N7828);
xor XOR2 (N13590, N13583, N2501);
or OR3 (N13591, N13575, N12506, N100);
and AND3 (N13592, N13578, N951, N190);
nand NAND3 (N13593, N13589, N1692, N12353);
or OR4 (N13594, N13588, N2480, N8711, N7206);
and AND2 (N13595, N13587, N9400);
or OR4 (N13596, N13576, N6937, N2470, N3566);
nand NAND4 (N13597, N13592, N6690, N3239, N11356);
xor XOR2 (N13598, N13597, N3193);
buf BUF1 (N13599, N13590);
nand NAND3 (N13600, N13598, N5940, N5085);
and AND2 (N13601, N13586, N2030);
and AND4 (N13602, N13580, N12385, N6964, N7023);
buf BUF1 (N13603, N13593);
and AND2 (N13604, N13601, N11363);
not NOT1 (N13605, N13604);
xor XOR2 (N13606, N13596, N11231);
buf BUF1 (N13607, N13602);
or OR4 (N13608, N13606, N9517, N8374, N4371);
and AND4 (N13609, N13607, N6939, N2863, N1228);
nand NAND2 (N13610, N13603, N11799);
nand NAND4 (N13611, N13599, N3286, N9197, N2437);
not NOT1 (N13612, N13610);
nand NAND4 (N13613, N13605, N13166, N5663, N13068);
and AND3 (N13614, N13609, N11983, N359);
xor XOR2 (N13615, N13595, N9245);
not NOT1 (N13616, N13611);
or OR4 (N13617, N13594, N2359, N4459, N3839);
nand NAND2 (N13618, N13600, N5352);
xor XOR2 (N13619, N13617, N3723);
xor XOR2 (N13620, N13619, N5617);
nor NOR3 (N13621, N13585, N13614, N13273);
buf BUF1 (N13622, N7494);
or OR4 (N13623, N13591, N10443, N11623, N10418);
nand NAND4 (N13624, N13623, N4199, N1738, N6084);
nand NAND2 (N13625, N13615, N9451);
or OR2 (N13626, N13616, N1894);
buf BUF1 (N13627, N13608);
nand NAND2 (N13628, N13622, N11347);
nor NOR2 (N13629, N13613, N473);
nor NOR4 (N13630, N13626, N7083, N6201, N9069);
or OR4 (N13631, N13620, N6371, N1584, N6542);
xor XOR2 (N13632, N13627, N6217);
xor XOR2 (N13633, N13612, N6482);
or OR4 (N13634, N13632, N6801, N10820, N11605);
nand NAND2 (N13635, N13633, N6916);
or OR3 (N13636, N13631, N9716, N12379);
nand NAND2 (N13637, N13618, N10474);
or OR4 (N13638, N13621, N10339, N4798, N2515);
xor XOR2 (N13639, N13630, N2181);
nor NOR4 (N13640, N13637, N5570, N11090, N2323);
not NOT1 (N13641, N13635);
buf BUF1 (N13642, N13629);
nand NAND4 (N13643, N13636, N2397, N2648, N5143);
nand NAND3 (N13644, N13641, N12498, N305);
nand NAND3 (N13645, N13644, N11698, N9277);
or OR2 (N13646, N13642, N13194);
xor XOR2 (N13647, N13639, N11991);
xor XOR2 (N13648, N13624, N13630);
xor XOR2 (N13649, N13643, N2995);
and AND4 (N13650, N13646, N3421, N12046, N2468);
nand NAND2 (N13651, N13647, N3254);
xor XOR2 (N13652, N13634, N2174);
or OR4 (N13653, N13645, N9511, N7812, N8783);
xor XOR2 (N13654, N13653, N5416);
or OR4 (N13655, N13640, N10488, N8051, N7016);
nand NAND4 (N13656, N13652, N7513, N10271, N13054);
or OR3 (N13657, N13654, N987, N13090);
buf BUF1 (N13658, N13628);
nand NAND4 (N13659, N13657, N7522, N6744, N8173);
xor XOR2 (N13660, N13658, N7602);
not NOT1 (N13661, N13655);
or OR2 (N13662, N13660, N6809);
nor NOR3 (N13663, N13656, N9901, N10436);
buf BUF1 (N13664, N13661);
and AND4 (N13665, N13648, N11183, N9714, N13578);
nand NAND4 (N13666, N13659, N10986, N11313, N9177);
nor NOR4 (N13667, N13663, N12362, N11769, N13075);
or OR2 (N13668, N13638, N1942);
or OR4 (N13669, N13665, N13159, N1110, N12383);
and AND2 (N13670, N13669, N13103);
xor XOR2 (N13671, N13666, N417);
xor XOR2 (N13672, N13651, N2761);
not NOT1 (N13673, N13672);
not NOT1 (N13674, N13662);
and AND3 (N13675, N13674, N4521, N10461);
xor XOR2 (N13676, N13671, N4018);
buf BUF1 (N13677, N13676);
and AND3 (N13678, N13650, N1678, N1905);
not NOT1 (N13679, N13649);
not NOT1 (N13680, N13664);
not NOT1 (N13681, N13670);
nand NAND4 (N13682, N13678, N7928, N5513, N11984);
nor NOR2 (N13683, N13667, N10838);
or OR3 (N13684, N13681, N8868, N732);
not NOT1 (N13685, N13668);
not NOT1 (N13686, N13673);
or OR3 (N13687, N13682, N11290, N4003);
xor XOR2 (N13688, N13679, N10280);
buf BUF1 (N13689, N13675);
and AND4 (N13690, N13625, N7357, N6281, N6572);
nand NAND3 (N13691, N13684, N1050, N1892);
not NOT1 (N13692, N13691);
or OR3 (N13693, N13688, N3421, N9750);
nand NAND3 (N13694, N13690, N13332, N1690);
nor NOR2 (N13695, N13694, N13199);
and AND2 (N13696, N13677, N5543);
not NOT1 (N13697, N13680);
buf BUF1 (N13698, N13685);
and AND2 (N13699, N13692, N11896);
and AND3 (N13700, N13695, N2231, N11213);
nor NOR2 (N13701, N13698, N9121);
buf BUF1 (N13702, N13697);
not NOT1 (N13703, N13683);
and AND2 (N13704, N13701, N12159);
and AND3 (N13705, N13689, N9926, N8971);
nor NOR2 (N13706, N13696, N2371);
buf BUF1 (N13707, N13687);
buf BUF1 (N13708, N13705);
not NOT1 (N13709, N13706);
and AND3 (N13710, N13707, N10746, N6261);
buf BUF1 (N13711, N13686);
not NOT1 (N13712, N13711);
nor NOR4 (N13713, N13709, N4200, N6265, N6528);
nor NOR3 (N13714, N13699, N11220, N10663);
and AND3 (N13715, N13713, N11698, N13307);
and AND4 (N13716, N13712, N9032, N12114, N7077);
and AND3 (N13717, N13700, N10085, N9588);
nor NOR4 (N13718, N13710, N2444, N4309, N5584);
and AND4 (N13719, N13703, N2852, N1388, N4150);
nor NOR3 (N13720, N13714, N5185, N6463);
nand NAND3 (N13721, N13720, N29, N481);
nor NOR4 (N13722, N13702, N1171, N13192, N2700);
not NOT1 (N13723, N13704);
xor XOR2 (N13724, N13693, N10767);
and AND4 (N13725, N13715, N7075, N3215, N6637);
or OR4 (N13726, N13718, N10751, N1831, N4017);
xor XOR2 (N13727, N13721, N13326);
and AND4 (N13728, N13724, N12334, N4454, N9050);
or OR4 (N13729, N13719, N2727, N13440, N11882);
nor NOR2 (N13730, N13722, N8316);
nor NOR2 (N13731, N13727, N10595);
nand NAND2 (N13732, N13731, N5332);
buf BUF1 (N13733, N13728);
not NOT1 (N13734, N13708);
or OR2 (N13735, N13726, N1208);
not NOT1 (N13736, N13732);
not NOT1 (N13737, N13735);
nand NAND2 (N13738, N13734, N2190);
xor XOR2 (N13739, N13736, N10510);
or OR4 (N13740, N13716, N10654, N5447, N1763);
or OR4 (N13741, N13730, N10207, N5087, N12116);
xor XOR2 (N13742, N13729, N9257);
not NOT1 (N13743, N13740);
or OR3 (N13744, N13741, N782, N845);
buf BUF1 (N13745, N13738);
nand NAND2 (N13746, N13744, N1306);
or OR2 (N13747, N13746, N6222);
xor XOR2 (N13748, N13733, N2817);
and AND4 (N13749, N13737, N8602, N1734, N13732);
buf BUF1 (N13750, N13725);
not NOT1 (N13751, N13717);
nor NOR2 (N13752, N13742, N9101);
and AND2 (N13753, N13723, N6217);
xor XOR2 (N13754, N13745, N5245);
or OR4 (N13755, N13739, N4150, N1931, N8358);
nor NOR2 (N13756, N13749, N892);
nand NAND4 (N13757, N13750, N2959, N996, N10886);
not NOT1 (N13758, N13755);
xor XOR2 (N13759, N13758, N2226);
and AND4 (N13760, N13753, N2312, N2779, N719);
or OR2 (N13761, N13757, N1611);
buf BUF1 (N13762, N13760);
xor XOR2 (N13763, N13756, N6128);
xor XOR2 (N13764, N13759, N2533);
not NOT1 (N13765, N13751);
or OR4 (N13766, N13763, N11076, N10557, N10081);
nor NOR2 (N13767, N13765, N4430);
or OR2 (N13768, N13752, N8057);
xor XOR2 (N13769, N13754, N5010);
and AND2 (N13770, N13762, N8949);
xor XOR2 (N13771, N13768, N12247);
buf BUF1 (N13772, N13769);
buf BUF1 (N13773, N13764);
buf BUF1 (N13774, N13743);
nand NAND3 (N13775, N13761, N3723, N49);
not NOT1 (N13776, N13770);
xor XOR2 (N13777, N13775, N9073);
not NOT1 (N13778, N13776);
xor XOR2 (N13779, N13767, N9159);
and AND3 (N13780, N13747, N9405, N2854);
buf BUF1 (N13781, N13778);
or OR3 (N13782, N13773, N9374, N12910);
buf BUF1 (N13783, N13777);
not NOT1 (N13784, N13766);
and AND4 (N13785, N13784, N1504, N11172, N12814);
nand NAND3 (N13786, N13782, N7268, N3336);
nor NOR4 (N13787, N13771, N2576, N9888, N11369);
and AND4 (N13788, N13785, N4715, N1711, N10421);
buf BUF1 (N13789, N13774);
not NOT1 (N13790, N13789);
or OR4 (N13791, N13786, N3744, N1867, N3832);
nand NAND3 (N13792, N13787, N8519, N6667);
or OR2 (N13793, N13779, N3655);
not NOT1 (N13794, N13792);
nor NOR2 (N13795, N13788, N3620);
nor NOR4 (N13796, N13791, N12491, N13593, N6950);
buf BUF1 (N13797, N13783);
nor NOR4 (N13798, N13797, N7126, N11631, N10177);
nand NAND2 (N13799, N13794, N8430);
xor XOR2 (N13800, N13795, N2776);
nor NOR4 (N13801, N13793, N10092, N4350, N6623);
or OR4 (N13802, N13780, N2943, N10177, N163);
or OR3 (N13803, N13790, N12825, N13685);
and AND4 (N13804, N13772, N9199, N515, N5709);
not NOT1 (N13805, N13803);
xor XOR2 (N13806, N13781, N12643);
nand NAND3 (N13807, N13796, N8741, N9952);
and AND2 (N13808, N13798, N9790);
buf BUF1 (N13809, N13799);
nor NOR4 (N13810, N13805, N12263, N3777, N13743);
and AND2 (N13811, N13800, N6438);
xor XOR2 (N13812, N13802, N7227);
buf BUF1 (N13813, N13806);
buf BUF1 (N13814, N13801);
buf BUF1 (N13815, N13748);
nor NOR3 (N13816, N13813, N4798, N7558);
or OR2 (N13817, N13807, N10016);
nor NOR2 (N13818, N13809, N4511);
nor NOR2 (N13819, N13810, N7350);
xor XOR2 (N13820, N13811, N4848);
xor XOR2 (N13821, N13804, N5951);
buf BUF1 (N13822, N13821);
not NOT1 (N13823, N13814);
nand NAND4 (N13824, N13819, N9916, N8444, N13250);
buf BUF1 (N13825, N13824);
not NOT1 (N13826, N13825);
buf BUF1 (N13827, N13818);
xor XOR2 (N13828, N13827, N610);
not NOT1 (N13829, N13828);
nor NOR2 (N13830, N13829, N902);
not NOT1 (N13831, N13812);
xor XOR2 (N13832, N13815, N10712);
buf BUF1 (N13833, N13822);
and AND4 (N13834, N13832, N5058, N8955, N8471);
or OR2 (N13835, N13831, N3621);
xor XOR2 (N13836, N13830, N9501);
nor NOR4 (N13837, N13823, N9457, N3595, N10478);
not NOT1 (N13838, N13820);
xor XOR2 (N13839, N13833, N8850);
not NOT1 (N13840, N13817);
and AND3 (N13841, N13816, N1523, N4633);
xor XOR2 (N13842, N13808, N13796);
and AND3 (N13843, N13834, N90, N10466);
buf BUF1 (N13844, N13826);
and AND4 (N13845, N13839, N845, N10400, N11552);
nand NAND2 (N13846, N13841, N8182);
nor NOR2 (N13847, N13846, N11728);
nor NOR4 (N13848, N13844, N6379, N12569, N1838);
xor XOR2 (N13849, N13838, N5599);
nor NOR4 (N13850, N13845, N4087, N11781, N3006);
not NOT1 (N13851, N13842);
nor NOR2 (N13852, N13851, N13380);
xor XOR2 (N13853, N13835, N8099);
not NOT1 (N13854, N13848);
and AND4 (N13855, N13843, N4594, N5410, N1160);
and AND2 (N13856, N13852, N4862);
nand NAND3 (N13857, N13850, N13289, N13401);
or OR3 (N13858, N13856, N5820, N7650);
buf BUF1 (N13859, N13858);
or OR4 (N13860, N13855, N3529, N9609, N13433);
nor NOR3 (N13861, N13840, N13145, N69);
not NOT1 (N13862, N13849);
nor NOR2 (N13863, N13857, N9838);
and AND2 (N13864, N13859, N3567);
and AND3 (N13865, N13861, N2296, N12658);
and AND2 (N13866, N13853, N2271);
xor XOR2 (N13867, N13837, N8248);
and AND3 (N13868, N13854, N13073, N9596);
not NOT1 (N13869, N13864);
buf BUF1 (N13870, N13862);
nand NAND3 (N13871, N13866, N7727, N11088);
nor NOR2 (N13872, N13863, N2532);
buf BUF1 (N13873, N13836);
or OR3 (N13874, N13868, N1806, N6531);
and AND2 (N13875, N13872, N13851);
xor XOR2 (N13876, N13875, N12418);
not NOT1 (N13877, N13869);
or OR3 (N13878, N13865, N4790, N3375);
nor NOR3 (N13879, N13876, N6162, N9942);
nor NOR4 (N13880, N13860, N10685, N1021, N10701);
nand NAND2 (N13881, N13870, N11886);
and AND2 (N13882, N13878, N13260);
or OR3 (N13883, N13871, N9134, N12801);
nand NAND4 (N13884, N13847, N2905, N6382, N10631);
and AND4 (N13885, N13877, N932, N6818, N5385);
buf BUF1 (N13886, N13882);
xor XOR2 (N13887, N13873, N7863);
nand NAND3 (N13888, N13881, N10050, N8105);
nand NAND2 (N13889, N13879, N9323);
buf BUF1 (N13890, N13889);
not NOT1 (N13891, N13890);
not NOT1 (N13892, N13886);
nor NOR4 (N13893, N13891, N1465, N7968, N2049);
xor XOR2 (N13894, N13867, N13661);
nor NOR3 (N13895, N13887, N4493, N11092);
not NOT1 (N13896, N13893);
xor XOR2 (N13897, N13892, N7618);
or OR4 (N13898, N13895, N996, N3202, N4813);
xor XOR2 (N13899, N13897, N8804);
buf BUF1 (N13900, N13894);
or OR4 (N13901, N13880, N9489, N13740, N12624);
and AND3 (N13902, N13899, N12441, N13519);
buf BUF1 (N13903, N13900);
not NOT1 (N13904, N13898);
xor XOR2 (N13905, N13903, N3534);
or OR3 (N13906, N13902, N10490, N5054);
nand NAND3 (N13907, N13901, N7889, N987);
buf BUF1 (N13908, N13905);
or OR4 (N13909, N13904, N13514, N7017, N2261);
nor NOR2 (N13910, N13885, N8991);
nand NAND3 (N13911, N13888, N340, N7616);
xor XOR2 (N13912, N13896, N6867);
buf BUF1 (N13913, N13912);
and AND4 (N13914, N13909, N10863, N3867, N4735);
and AND3 (N13915, N13914, N2570, N7455);
and AND2 (N13916, N13913, N12123);
and AND3 (N13917, N13884, N6108, N7545);
or OR2 (N13918, N13911, N6718);
buf BUF1 (N13919, N13883);
or OR3 (N13920, N13910, N13513, N9187);
or OR3 (N13921, N13915, N6659, N674);
xor XOR2 (N13922, N13907, N3367);
xor XOR2 (N13923, N13922, N11713);
buf BUF1 (N13924, N13908);
buf BUF1 (N13925, N13923);
nand NAND2 (N13926, N13919, N6642);
buf BUF1 (N13927, N13874);
nand NAND3 (N13928, N13917, N8359, N5983);
nand NAND3 (N13929, N13916, N7939, N7570);
nor NOR3 (N13930, N13925, N9407, N8521);
and AND3 (N13931, N13920, N9626, N8651);
nand NAND3 (N13932, N13906, N9546, N3429);
buf BUF1 (N13933, N13928);
not NOT1 (N13934, N13933);
nand NAND3 (N13935, N13930, N7378, N11079);
or OR2 (N13936, N13927, N6488);
not NOT1 (N13937, N13935);
buf BUF1 (N13938, N13934);
not NOT1 (N13939, N13921);
and AND2 (N13940, N13918, N6654);
or OR3 (N13941, N13929, N1367, N7614);
xor XOR2 (N13942, N13931, N2034);
and AND2 (N13943, N13939, N9127);
buf BUF1 (N13944, N13924);
not NOT1 (N13945, N13932);
and AND3 (N13946, N13942, N2455, N1109);
nand NAND3 (N13947, N13940, N5982, N1805);
nand NAND4 (N13948, N13947, N5889, N3771, N3900);
xor XOR2 (N13949, N13936, N11936);
nor NOR4 (N13950, N13943, N10688, N8362, N9073);
not NOT1 (N13951, N13948);
nor NOR2 (N13952, N13938, N5266);
nand NAND3 (N13953, N13944, N10497, N3359);
and AND3 (N13954, N13926, N3816, N4473);
buf BUF1 (N13955, N13937);
xor XOR2 (N13956, N13941, N1985);
xor XOR2 (N13957, N13952, N376);
nor NOR4 (N13958, N13946, N12822, N2911, N4385);
nand NAND4 (N13959, N13957, N10949, N4717, N5461);
xor XOR2 (N13960, N13958, N1435);
buf BUF1 (N13961, N13945);
xor XOR2 (N13962, N13953, N8579);
and AND2 (N13963, N13949, N11942);
and AND2 (N13964, N13950, N7102);
or OR3 (N13965, N13955, N11724, N8898);
and AND2 (N13966, N13960, N6997);
buf BUF1 (N13967, N13965);
buf BUF1 (N13968, N13963);
not NOT1 (N13969, N13959);
nor NOR4 (N13970, N13951, N10910, N8709, N13582);
or OR4 (N13971, N13961, N5307, N2388, N5093);
or OR3 (N13972, N13969, N1354, N13356);
not NOT1 (N13973, N13964);
not NOT1 (N13974, N13966);
and AND3 (N13975, N13973, N10632, N2796);
nor NOR3 (N13976, N13971, N9302, N6264);
nor NOR4 (N13977, N13972, N6968, N1335, N8556);
buf BUF1 (N13978, N13976);
nand NAND4 (N13979, N13974, N6972, N8928, N8534);
buf BUF1 (N13980, N13956);
not NOT1 (N13981, N13980);
nor NOR2 (N13982, N13978, N5706);
and AND3 (N13983, N13968, N8510, N7375);
and AND2 (N13984, N13983, N11988);
nand NAND3 (N13985, N13967, N9576, N8680);
xor XOR2 (N13986, N13985, N7943);
and AND4 (N13987, N13954, N7306, N13150, N12861);
and AND4 (N13988, N13962, N9269, N10020, N9721);
and AND4 (N13989, N13982, N2091, N8756, N11707);
nand NAND2 (N13990, N13970, N4876);
nor NOR2 (N13991, N13984, N10375);
xor XOR2 (N13992, N13990, N1346);
or OR3 (N13993, N13991, N3489, N3047);
buf BUF1 (N13994, N13989);
not NOT1 (N13995, N13993);
nor NOR3 (N13996, N13979, N4037, N561);
nor NOR3 (N13997, N13996, N5789, N9931);
buf BUF1 (N13998, N13988);
and AND2 (N13999, N13997, N3289);
nand NAND3 (N14000, N13987, N10911, N11906);
xor XOR2 (N14001, N13975, N10310);
nand NAND2 (N14002, N13981, N10093);
not NOT1 (N14003, N13999);
buf BUF1 (N14004, N14003);
nor NOR4 (N14005, N13994, N9039, N1882, N3861);
or OR4 (N14006, N14000, N13956, N7004, N10334);
and AND2 (N14007, N14001, N3500);
xor XOR2 (N14008, N14002, N4154);
or OR3 (N14009, N13995, N8446, N11253);
nand NAND2 (N14010, N14005, N7965);
nor NOR2 (N14011, N13986, N13338);
nand NAND4 (N14012, N13977, N7624, N5626, N8249);
xor XOR2 (N14013, N13998, N13165);
or OR3 (N14014, N14006, N11760, N5585);
xor XOR2 (N14015, N13992, N1405);
nor NOR3 (N14016, N14009, N5591, N5022);
nand NAND4 (N14017, N14011, N3267, N5787, N10567);
buf BUF1 (N14018, N14010);
or OR4 (N14019, N14004, N8812, N5245, N5033);
nor NOR2 (N14020, N14018, N5018);
nor NOR3 (N14021, N14007, N847, N3535);
or OR2 (N14022, N14014, N11492);
or OR4 (N14023, N14019, N9192, N6711, N12563);
nand NAND2 (N14024, N14008, N11857);
xor XOR2 (N14025, N14021, N8111);
and AND2 (N14026, N14023, N6878);
xor XOR2 (N14027, N14022, N12576);
xor XOR2 (N14028, N14013, N6079);
nor NOR3 (N14029, N14026, N1552, N7954);
buf BUF1 (N14030, N14025);
not NOT1 (N14031, N14028);
nor NOR3 (N14032, N14016, N4442, N866);
nand NAND3 (N14033, N14015, N12489, N9998);
nand NAND3 (N14034, N14029, N7244, N11140);
or OR3 (N14035, N14024, N10436, N10780);
not NOT1 (N14036, N14034);
nand NAND2 (N14037, N14020, N11028);
or OR4 (N14038, N14032, N12623, N6259, N13699);
xor XOR2 (N14039, N14037, N9062);
nor NOR3 (N14040, N14036, N11270, N19);
xor XOR2 (N14041, N14031, N7140);
or OR3 (N14042, N14027, N3392, N10458);
nor NOR2 (N14043, N14041, N470);
or OR2 (N14044, N14035, N12172);
nand NAND4 (N14045, N14012, N12949, N5337, N4595);
xor XOR2 (N14046, N14039, N7152);
xor XOR2 (N14047, N14033, N4280);
nand NAND4 (N14048, N14038, N508, N3007, N2754);
nand NAND3 (N14049, N14030, N6658, N11236);
nor NOR4 (N14050, N14043, N6546, N9557, N6985);
buf BUF1 (N14051, N14042);
and AND4 (N14052, N14044, N121, N11220, N1088);
xor XOR2 (N14053, N14017, N8328);
nor NOR4 (N14054, N14049, N7474, N11213, N10019);
not NOT1 (N14055, N14045);
nor NOR4 (N14056, N14051, N5029, N2116, N4902);
or OR4 (N14057, N14047, N7704, N9358, N12296);
nor NOR4 (N14058, N14053, N10067, N8679, N1043);
xor XOR2 (N14059, N14050, N8564);
and AND3 (N14060, N14048, N7259, N4125);
not NOT1 (N14061, N14052);
nand NAND4 (N14062, N14056, N8021, N8043, N6592);
xor XOR2 (N14063, N14054, N4916);
and AND2 (N14064, N14063, N8030);
not NOT1 (N14065, N14059);
not NOT1 (N14066, N14062);
or OR3 (N14067, N14060, N12728, N10628);
buf BUF1 (N14068, N14055);
xor XOR2 (N14069, N14046, N7372);
xor XOR2 (N14070, N14057, N11069);
not NOT1 (N14071, N14068);
not NOT1 (N14072, N14066);
nor NOR4 (N14073, N14040, N6599, N4023, N10314);
nor NOR3 (N14074, N14065, N12253, N10078);
xor XOR2 (N14075, N14070, N13961);
buf BUF1 (N14076, N14064);
or OR2 (N14077, N14061, N1537);
not NOT1 (N14078, N14074);
buf BUF1 (N14079, N14078);
or OR2 (N14080, N14069, N61);
or OR3 (N14081, N14073, N7282, N13597);
nand NAND2 (N14082, N14071, N8316);
xor XOR2 (N14083, N14079, N11508);
not NOT1 (N14084, N14075);
nor NOR2 (N14085, N14072, N13741);
nand NAND2 (N14086, N14083, N3610);
or OR3 (N14087, N14085, N11968, N5534);
xor XOR2 (N14088, N14058, N12096);
or OR2 (N14089, N14080, N3301);
or OR2 (N14090, N14076, N6755);
and AND3 (N14091, N14084, N6727, N7766);
and AND4 (N14092, N14067, N4391, N5952, N3904);
nand NAND4 (N14093, N14090, N10292, N6104, N9176);
buf BUF1 (N14094, N14092);
buf BUF1 (N14095, N14094);
buf BUF1 (N14096, N14088);
xor XOR2 (N14097, N14087, N5744);
buf BUF1 (N14098, N14081);
xor XOR2 (N14099, N14095, N3647);
and AND3 (N14100, N14093, N13377, N953);
xor XOR2 (N14101, N14082, N13762);
not NOT1 (N14102, N14077);
not NOT1 (N14103, N14099);
or OR3 (N14104, N14086, N10456, N12801);
or OR2 (N14105, N14100, N8891);
nor NOR4 (N14106, N14103, N4962, N4755, N7435);
not NOT1 (N14107, N14104);
buf BUF1 (N14108, N14096);
nor NOR2 (N14109, N14091, N8266);
xor XOR2 (N14110, N14108, N5935);
buf BUF1 (N14111, N14107);
buf BUF1 (N14112, N14089);
nor NOR2 (N14113, N14111, N5645);
nor NOR3 (N14114, N14106, N13154, N11883);
or OR3 (N14115, N14105, N1616, N2457);
and AND4 (N14116, N14112, N1394, N7971, N9986);
nand NAND3 (N14117, N14110, N1576, N10079);
buf BUF1 (N14118, N14115);
xor XOR2 (N14119, N14118, N3505);
buf BUF1 (N14120, N14101);
nor NOR2 (N14121, N14113, N1275);
buf BUF1 (N14122, N14109);
xor XOR2 (N14123, N14122, N762);
and AND3 (N14124, N14098, N10077, N7939);
or OR4 (N14125, N14114, N7188, N11631, N1681);
nand NAND2 (N14126, N14123, N4373);
nor NOR2 (N14127, N14117, N8429);
nand NAND4 (N14128, N14125, N13780, N3134, N1596);
and AND4 (N14129, N14128, N7798, N8442, N8158);
buf BUF1 (N14130, N14129);
not NOT1 (N14131, N14097);
not NOT1 (N14132, N14131);
nor NOR4 (N14133, N14102, N623, N9932, N8928);
nor NOR3 (N14134, N14119, N2533, N1345);
xor XOR2 (N14135, N14130, N11765);
xor XOR2 (N14136, N14127, N8279);
not NOT1 (N14137, N14133);
buf BUF1 (N14138, N14116);
nand NAND4 (N14139, N14121, N5083, N5398, N12722);
buf BUF1 (N14140, N14120);
buf BUF1 (N14141, N14140);
and AND2 (N14142, N14132, N1619);
buf BUF1 (N14143, N14134);
or OR2 (N14144, N14137, N14055);
xor XOR2 (N14145, N14135, N6094);
nand NAND3 (N14146, N14139, N3954, N2779);
nand NAND2 (N14147, N14141, N12872);
not NOT1 (N14148, N14136);
not NOT1 (N14149, N14138);
not NOT1 (N14150, N14149);
buf BUF1 (N14151, N14142);
or OR3 (N14152, N14144, N3931, N372);
xor XOR2 (N14153, N14145, N1199);
nor NOR4 (N14154, N14148, N5238, N2336, N12001);
nand NAND3 (N14155, N14126, N5783, N1742);
and AND3 (N14156, N14147, N4344, N12533);
nand NAND2 (N14157, N14151, N5509);
buf BUF1 (N14158, N14157);
and AND2 (N14159, N14146, N3028);
xor XOR2 (N14160, N14150, N5010);
and AND4 (N14161, N14152, N8260, N12053, N13154);
nand NAND3 (N14162, N14143, N9512, N2755);
nand NAND2 (N14163, N14156, N1484);
nand NAND2 (N14164, N14155, N2329);
or OR4 (N14165, N14160, N9568, N12424, N2);
nor NOR3 (N14166, N14164, N4200, N1086);
buf BUF1 (N14167, N14153);
nor NOR4 (N14168, N14167, N565, N4968, N5696);
xor XOR2 (N14169, N14154, N2893);
or OR3 (N14170, N14161, N334, N12940);
buf BUF1 (N14171, N14159);
nor NOR3 (N14172, N14158, N8661, N9008);
xor XOR2 (N14173, N14162, N2571);
or OR3 (N14174, N14165, N3269, N10349);
not NOT1 (N14175, N14169);
or OR4 (N14176, N14166, N9315, N11451, N12746);
and AND2 (N14177, N14171, N7681);
nand NAND3 (N14178, N14163, N3745, N9129);
or OR2 (N14179, N14124, N4054);
nand NAND4 (N14180, N14179, N9398, N5861, N1139);
and AND4 (N14181, N14180, N9785, N9002, N2012);
and AND2 (N14182, N14181, N3679);
xor XOR2 (N14183, N14182, N10250);
nor NOR2 (N14184, N14175, N7709);
nor NOR3 (N14185, N14184, N13450, N7767);
not NOT1 (N14186, N14183);
or OR3 (N14187, N14173, N172, N9370);
nor NOR4 (N14188, N14172, N5098, N8387, N9012);
nand NAND4 (N14189, N14174, N5599, N2305, N4255);
xor XOR2 (N14190, N14168, N9492);
xor XOR2 (N14191, N14190, N4313);
nor NOR4 (N14192, N14176, N3896, N453, N11106);
nand NAND2 (N14193, N14187, N1974);
nor NOR4 (N14194, N14178, N10886, N885, N3432);
nor NOR4 (N14195, N14188, N11256, N7357, N11960);
nand NAND2 (N14196, N14193, N9204);
buf BUF1 (N14197, N14177);
xor XOR2 (N14198, N14194, N1123);
nor NOR2 (N14199, N14189, N10132);
xor XOR2 (N14200, N14196, N2269);
buf BUF1 (N14201, N14200);
nand NAND2 (N14202, N14195, N13198);
or OR3 (N14203, N14197, N7260, N2730);
xor XOR2 (N14204, N14199, N12183);
nor NOR3 (N14205, N14191, N8754, N13481);
or OR2 (N14206, N14186, N5624);
or OR3 (N14207, N14192, N5859, N4161);
and AND3 (N14208, N14205, N3280, N11630);
nor NOR4 (N14209, N14207, N7895, N9063, N10519);
xor XOR2 (N14210, N14204, N8264);
nand NAND4 (N14211, N14201, N1588, N13845, N7414);
or OR3 (N14212, N14170, N12513, N4451);
nand NAND2 (N14213, N14198, N145);
nor NOR4 (N14214, N14203, N33, N9306, N10317);
or OR4 (N14215, N14210, N9427, N11981, N6586);
or OR3 (N14216, N14215, N10398, N1931);
nor NOR4 (N14217, N14212, N6400, N13434, N3812);
xor XOR2 (N14218, N14217, N4284);
buf BUF1 (N14219, N14211);
nand NAND4 (N14220, N14208, N1028, N744, N3180);
or OR4 (N14221, N14216, N7510, N511, N2139);
nand NAND3 (N14222, N14218, N6117, N3102);
nor NOR3 (N14223, N14219, N1336, N5259);
buf BUF1 (N14224, N14209);
xor XOR2 (N14225, N14185, N4963);
nor NOR4 (N14226, N14222, N6850, N4598, N4483);
nand NAND4 (N14227, N14225, N2474, N9452, N7556);
and AND3 (N14228, N14221, N5002, N9900);
or OR3 (N14229, N14228, N12648, N4614);
nor NOR2 (N14230, N14213, N10914);
nor NOR4 (N14231, N14224, N861, N10073, N10920);
and AND3 (N14232, N14202, N10226, N14022);
not NOT1 (N14233, N14232);
or OR4 (N14234, N14214, N7194, N4867, N3249);
nand NAND4 (N14235, N14231, N5526, N13841, N2949);
not NOT1 (N14236, N14234);
nor NOR2 (N14237, N14229, N7434);
buf BUF1 (N14238, N14223);
xor XOR2 (N14239, N14206, N11581);
nand NAND2 (N14240, N14220, N12946);
buf BUF1 (N14241, N14239);
buf BUF1 (N14242, N14241);
buf BUF1 (N14243, N14236);
buf BUF1 (N14244, N14235);
and AND3 (N14245, N14244, N13483, N2083);
xor XOR2 (N14246, N14242, N4585);
xor XOR2 (N14247, N14227, N12386);
xor XOR2 (N14248, N14237, N6496);
nor NOR2 (N14249, N14238, N11763);
and AND3 (N14250, N14249, N10093, N7749);
nor NOR4 (N14251, N14247, N7710, N6395, N5307);
not NOT1 (N14252, N14246);
or OR4 (N14253, N14245, N2216, N3239, N13770);
not NOT1 (N14254, N14253);
and AND4 (N14255, N14240, N9400, N13807, N11350);
nor NOR3 (N14256, N14252, N1809, N9611);
or OR4 (N14257, N14243, N10000, N12428, N5040);
not NOT1 (N14258, N14256);
nand NAND4 (N14259, N14254, N319, N6707, N11826);
and AND4 (N14260, N14233, N656, N13146, N4037);
or OR4 (N14261, N14230, N1675, N4433, N9671);
or OR2 (N14262, N14257, N7295);
nor NOR2 (N14263, N14258, N5836);
nor NOR4 (N14264, N14255, N7246, N5007, N10499);
buf BUF1 (N14265, N14250);
not NOT1 (N14266, N14251);
and AND4 (N14267, N14226, N5098, N13523, N7685);
and AND4 (N14268, N14261, N380, N6655, N8536);
and AND4 (N14269, N14266, N3368, N11401, N2641);
xor XOR2 (N14270, N14260, N10581);
and AND2 (N14271, N14263, N1907);
and AND2 (N14272, N14271, N6876);
nor NOR3 (N14273, N14269, N1400, N7872);
or OR4 (N14274, N14270, N1149, N1917, N3578);
not NOT1 (N14275, N14264);
nor NOR3 (N14276, N14267, N2928, N10640);
not NOT1 (N14277, N14273);
buf BUF1 (N14278, N14259);
buf BUF1 (N14279, N14265);
or OR2 (N14280, N14262, N5403);
nor NOR2 (N14281, N14248, N13251);
and AND2 (N14282, N14276, N10246);
xor XOR2 (N14283, N14277, N10881);
nor NOR2 (N14284, N14268, N5247);
not NOT1 (N14285, N14274);
xor XOR2 (N14286, N14278, N3469);
buf BUF1 (N14287, N14284);
not NOT1 (N14288, N14281);
nand NAND2 (N14289, N14272, N2402);
nor NOR4 (N14290, N14279, N6268, N395, N6849);
buf BUF1 (N14291, N14288);
buf BUF1 (N14292, N14291);
buf BUF1 (N14293, N14275);
buf BUF1 (N14294, N14282);
buf BUF1 (N14295, N14280);
not NOT1 (N14296, N14293);
xor XOR2 (N14297, N14283, N12988);
buf BUF1 (N14298, N14297);
and AND4 (N14299, N14298, N4225, N4463, N7172);
buf BUF1 (N14300, N14286);
nand NAND2 (N14301, N14289, N2714);
nand NAND3 (N14302, N14300, N7849, N10216);
xor XOR2 (N14303, N14299, N3685);
not NOT1 (N14304, N14294);
buf BUF1 (N14305, N14302);
and AND3 (N14306, N14296, N888, N2247);
not NOT1 (N14307, N14292);
and AND4 (N14308, N14301, N8952, N7153, N12125);
nor NOR3 (N14309, N14295, N13100, N9315);
and AND4 (N14310, N14307, N7329, N3522, N13296);
xor XOR2 (N14311, N14303, N10530);
or OR2 (N14312, N14285, N5124);
buf BUF1 (N14313, N14312);
nand NAND3 (N14314, N14287, N11301, N7408);
not NOT1 (N14315, N14309);
not NOT1 (N14316, N14306);
nand NAND2 (N14317, N14313, N7306);
buf BUF1 (N14318, N14308);
and AND4 (N14319, N14314, N1069, N10618, N13289);
xor XOR2 (N14320, N14317, N13508);
xor XOR2 (N14321, N14304, N4279);
and AND4 (N14322, N14320, N4626, N2551, N911);
and AND4 (N14323, N14311, N13019, N13670, N5191);
nand NAND3 (N14324, N14318, N335, N11928);
xor XOR2 (N14325, N14316, N13310);
and AND2 (N14326, N14315, N9130);
nand NAND3 (N14327, N14326, N10113, N3108);
nand NAND3 (N14328, N14305, N1634, N6673);
and AND3 (N14329, N14310, N7787, N3846);
and AND3 (N14330, N14328, N9394, N10298);
nor NOR3 (N14331, N14327, N12266, N9009);
or OR4 (N14332, N14323, N8736, N7367, N7886);
buf BUF1 (N14333, N14331);
nor NOR3 (N14334, N14324, N2023, N7255);
and AND2 (N14335, N14290, N8533);
xor XOR2 (N14336, N14319, N2193);
not NOT1 (N14337, N14332);
xor XOR2 (N14338, N14333, N1439);
xor XOR2 (N14339, N14338, N1540);
buf BUF1 (N14340, N14339);
or OR2 (N14341, N14330, N6566);
or OR4 (N14342, N14329, N13384, N11423, N2744);
xor XOR2 (N14343, N14334, N2717);
not NOT1 (N14344, N14335);
or OR3 (N14345, N14325, N11857, N3469);
and AND3 (N14346, N14345, N2222, N9344);
and AND2 (N14347, N14342, N785);
and AND3 (N14348, N14347, N12830, N141);
xor XOR2 (N14349, N14341, N10333);
not NOT1 (N14350, N14346);
xor XOR2 (N14351, N14343, N12230);
not NOT1 (N14352, N14344);
nor NOR2 (N14353, N14351, N8242);
or OR2 (N14354, N14350, N5199);
nor NOR4 (N14355, N14348, N8126, N11536, N2276);
xor XOR2 (N14356, N14354, N13525);
not NOT1 (N14357, N14336);
and AND4 (N14358, N14349, N5031, N8176, N3884);
xor XOR2 (N14359, N14353, N12294);
and AND2 (N14360, N14357, N7744);
buf BUF1 (N14361, N14352);
nand NAND3 (N14362, N14321, N10577, N11375);
not NOT1 (N14363, N14359);
and AND3 (N14364, N14337, N10401, N1233);
and AND2 (N14365, N14364, N7890);
and AND3 (N14366, N14322, N13843, N9981);
nor NOR2 (N14367, N14361, N5093);
nand NAND3 (N14368, N14340, N1894, N7651);
xor XOR2 (N14369, N14363, N5131);
not NOT1 (N14370, N14368);
not NOT1 (N14371, N14369);
nor NOR2 (N14372, N14358, N600);
and AND4 (N14373, N14367, N2739, N9499, N1731);
nand NAND4 (N14374, N14356, N13950, N12362, N13731);
and AND2 (N14375, N14365, N9169);
nand NAND2 (N14376, N14374, N6000);
xor XOR2 (N14377, N14362, N12166);
and AND4 (N14378, N14355, N13695, N1238, N840);
nor NOR3 (N14379, N14366, N10867, N5520);
not NOT1 (N14380, N14371);
xor XOR2 (N14381, N14370, N7969);
nand NAND3 (N14382, N14378, N3101, N1842);
buf BUF1 (N14383, N14375);
not NOT1 (N14384, N14380);
nand NAND2 (N14385, N14384, N13932);
xor XOR2 (N14386, N14376, N2782);
xor XOR2 (N14387, N14360, N11609);
nand NAND4 (N14388, N14379, N11735, N5473, N12264);
xor XOR2 (N14389, N14385, N9762);
buf BUF1 (N14390, N14372);
and AND4 (N14391, N14388, N11999, N11318, N9054);
nand NAND3 (N14392, N14383, N4342, N800);
nor NOR3 (N14393, N14381, N2178, N12526);
buf BUF1 (N14394, N14382);
buf BUF1 (N14395, N14389);
and AND3 (N14396, N14394, N12027, N13666);
not NOT1 (N14397, N14387);
and AND3 (N14398, N14390, N4837, N1552);
or OR3 (N14399, N14392, N3135, N12080);
and AND2 (N14400, N14393, N13670);
nor NOR2 (N14401, N14396, N2698);
not NOT1 (N14402, N14398);
xor XOR2 (N14403, N14386, N8919);
buf BUF1 (N14404, N14377);
xor XOR2 (N14405, N14397, N6796);
nand NAND3 (N14406, N14403, N6052, N1723);
not NOT1 (N14407, N14404);
and AND3 (N14408, N14400, N12947, N2091);
buf BUF1 (N14409, N14391);
buf BUF1 (N14410, N14407);
not NOT1 (N14411, N14409);
xor XOR2 (N14412, N14399, N4673);
nor NOR4 (N14413, N14402, N3174, N2151, N4220);
or OR3 (N14414, N14401, N12013, N1833);
nand NAND3 (N14415, N14414, N6087, N92);
xor XOR2 (N14416, N14408, N7493);
nor NOR4 (N14417, N14415, N8831, N13490, N10307);
nand NAND3 (N14418, N14410, N8433, N619);
xor XOR2 (N14419, N14406, N7753);
nand NAND4 (N14420, N14405, N852, N7773, N5350);
buf BUF1 (N14421, N14412);
and AND3 (N14422, N14421, N3598, N5034);
not NOT1 (N14423, N14416);
and AND3 (N14424, N14422, N7698, N9765);
and AND4 (N14425, N14411, N7234, N5240, N13331);
nand NAND2 (N14426, N14418, N2070);
nor NOR2 (N14427, N14426, N13036);
nand NAND4 (N14428, N14413, N1135, N3668, N2741);
buf BUF1 (N14429, N14424);
and AND2 (N14430, N14423, N200);
and AND4 (N14431, N14373, N8952, N3431, N5771);
not NOT1 (N14432, N14395);
nor NOR2 (N14433, N14420, N4545);
xor XOR2 (N14434, N14431, N6284);
nor NOR3 (N14435, N14429, N12150, N2691);
buf BUF1 (N14436, N14428);
and AND2 (N14437, N14433, N9659);
nand NAND4 (N14438, N14436, N10856, N12774, N9264);
and AND4 (N14439, N14438, N2491, N10001, N3141);
xor XOR2 (N14440, N14432, N3768);
not NOT1 (N14441, N14419);
nand NAND4 (N14442, N14439, N3650, N11096, N1999);
or OR2 (N14443, N14425, N10946);
and AND3 (N14444, N14427, N4812, N12393);
nand NAND4 (N14445, N14444, N12926, N1117, N2598);
and AND4 (N14446, N14443, N13574, N12779, N11239);
nand NAND3 (N14447, N14437, N1081, N12693);
not NOT1 (N14448, N14417);
nor NOR3 (N14449, N14435, N9244, N5515);
nand NAND3 (N14450, N14440, N3723, N2301);
and AND3 (N14451, N14450, N5667, N11489);
and AND3 (N14452, N14434, N14163, N11249);
or OR2 (N14453, N14447, N3743);
and AND4 (N14454, N14452, N3254, N5922, N623);
buf BUF1 (N14455, N14453);
xor XOR2 (N14456, N14448, N11186);
xor XOR2 (N14457, N14449, N11205);
not NOT1 (N14458, N14446);
nand NAND4 (N14459, N14441, N3895, N7612, N11525);
or OR3 (N14460, N14451, N4873, N8295);
buf BUF1 (N14461, N14456);
buf BUF1 (N14462, N14460);
and AND2 (N14463, N14457, N4191);
and AND2 (N14464, N14445, N5961);
buf BUF1 (N14465, N14464);
xor XOR2 (N14466, N14455, N4387);
buf BUF1 (N14467, N14442);
not NOT1 (N14468, N14467);
nor NOR2 (N14469, N14461, N7182);
nand NAND3 (N14470, N14459, N5311, N457);
not NOT1 (N14471, N14465);
nand NAND2 (N14472, N14430, N8359);
nor NOR4 (N14473, N14463, N7440, N4493, N8376);
and AND3 (N14474, N14468, N11160, N6604);
buf BUF1 (N14475, N14469);
not NOT1 (N14476, N14473);
nor NOR2 (N14477, N14476, N4024);
and AND4 (N14478, N14474, N6375, N1015, N7494);
nand NAND4 (N14479, N14470, N11324, N11127, N2321);
xor XOR2 (N14480, N14479, N9139);
or OR4 (N14481, N14458, N5528, N9540, N9102);
not NOT1 (N14482, N14471);
nor NOR4 (N14483, N14482, N5134, N4839, N11450);
or OR3 (N14484, N14483, N1387, N3075);
not NOT1 (N14485, N14480);
xor XOR2 (N14486, N14478, N6288);
nand NAND4 (N14487, N14477, N13904, N12088, N10008);
buf BUF1 (N14488, N14462);
buf BUF1 (N14489, N14475);
buf BUF1 (N14490, N14484);
buf BUF1 (N14491, N14490);
buf BUF1 (N14492, N14488);
buf BUF1 (N14493, N14489);
or OR2 (N14494, N14491, N8344);
not NOT1 (N14495, N14454);
or OR2 (N14496, N14486, N1877);
buf BUF1 (N14497, N14492);
buf BUF1 (N14498, N14481);
nand NAND4 (N14499, N14487, N9566, N11915, N2766);
nor NOR2 (N14500, N14466, N10456);
nand NAND3 (N14501, N14497, N3568, N11333);
and AND2 (N14502, N14496, N10400);
and AND4 (N14503, N14501, N12157, N2357, N4188);
nor NOR4 (N14504, N14503, N6610, N8977, N966);
or OR4 (N14505, N14499, N9276, N1389, N14249);
buf BUF1 (N14506, N14495);
xor XOR2 (N14507, N14500, N10696);
or OR3 (N14508, N14504, N11643, N4809);
nor NOR2 (N14509, N14498, N8537);
buf BUF1 (N14510, N14506);
and AND3 (N14511, N14510, N2209, N12198);
buf BUF1 (N14512, N14505);
nand NAND2 (N14513, N14507, N578);
xor XOR2 (N14514, N14511, N3745);
or OR4 (N14515, N14494, N11956, N7479, N8726);
nand NAND2 (N14516, N14485, N610);
xor XOR2 (N14517, N14493, N10880);
xor XOR2 (N14518, N14514, N3267);
and AND3 (N14519, N14513, N9842, N12328);
and AND2 (N14520, N14517, N6494);
nand NAND3 (N14521, N14518, N10219, N6191);
and AND2 (N14522, N14512, N7067);
and AND2 (N14523, N14520, N8224);
or OR4 (N14524, N14516, N3275, N2596, N2133);
and AND3 (N14525, N14502, N14313, N12264);
nand NAND3 (N14526, N14521, N10641, N1951);
nor NOR2 (N14527, N14522, N7635);
or OR3 (N14528, N14509, N11240, N301);
nor NOR3 (N14529, N14528, N5642, N5356);
not NOT1 (N14530, N14472);
and AND2 (N14531, N14530, N13238);
and AND3 (N14532, N14524, N7951, N2255);
and AND2 (N14533, N14515, N9937);
and AND4 (N14534, N14525, N682, N7223, N8087);
nand NAND3 (N14535, N14529, N6948, N6372);
nor NOR3 (N14536, N14523, N8587, N11999);
not NOT1 (N14537, N14519);
nor NOR4 (N14538, N14535, N7498, N5838, N12862);
buf BUF1 (N14539, N14534);
buf BUF1 (N14540, N14538);
and AND4 (N14541, N14508, N1373, N8917, N5297);
nor NOR2 (N14542, N14532, N11096);
nor NOR2 (N14543, N14533, N4814);
and AND2 (N14544, N14536, N11083);
xor XOR2 (N14545, N14527, N13415);
and AND4 (N14546, N14544, N7950, N4464, N4682);
nor NOR2 (N14547, N14531, N3598);
xor XOR2 (N14548, N14540, N745);
nor NOR3 (N14549, N14542, N13514, N3700);
buf BUF1 (N14550, N14543);
xor XOR2 (N14551, N14549, N13874);
or OR3 (N14552, N14537, N4072, N11516);
or OR2 (N14553, N14552, N10817);
or OR2 (N14554, N14550, N11411);
or OR4 (N14555, N14546, N4171, N210, N10434);
xor XOR2 (N14556, N14539, N3482);
nand NAND2 (N14557, N14541, N2863);
or OR3 (N14558, N14553, N8324, N14383);
nand NAND3 (N14559, N14526, N9872, N5167);
xor XOR2 (N14560, N14548, N8269);
nand NAND2 (N14561, N14557, N10493);
nor NOR4 (N14562, N14554, N13857, N6025, N10643);
nor NOR2 (N14563, N14555, N11592);
buf BUF1 (N14564, N14556);
and AND2 (N14565, N14561, N12195);
not NOT1 (N14566, N14559);
not NOT1 (N14567, N14551);
nand NAND4 (N14568, N14567, N13492, N8704, N2551);
xor XOR2 (N14569, N14558, N14169);
xor XOR2 (N14570, N14566, N631);
and AND2 (N14571, N14545, N7715);
buf BUF1 (N14572, N14562);
xor XOR2 (N14573, N14569, N2258);
xor XOR2 (N14574, N14573, N6097);
and AND3 (N14575, N14564, N8611, N6275);
not NOT1 (N14576, N14570);
buf BUF1 (N14577, N14575);
and AND4 (N14578, N14547, N8877, N13623, N6251);
buf BUF1 (N14579, N14568);
or OR4 (N14580, N14560, N11664, N4677, N14184);
not NOT1 (N14581, N14571);
and AND3 (N14582, N14577, N11996, N13296);
xor XOR2 (N14583, N14582, N3324);
nand NAND3 (N14584, N14581, N8739, N5404);
nand NAND2 (N14585, N14576, N13931);
buf BUF1 (N14586, N14574);
nand NAND3 (N14587, N14580, N11740, N6909);
and AND2 (N14588, N14583, N1086);
buf BUF1 (N14589, N14588);
or OR3 (N14590, N14565, N7546, N10958);
or OR2 (N14591, N14590, N7820);
nand NAND3 (N14592, N14572, N9000, N11577);
nor NOR2 (N14593, N14584, N5913);
nand NAND2 (N14594, N14585, N6994);
or OR3 (N14595, N14587, N12888, N406);
buf BUF1 (N14596, N14578);
nand NAND4 (N14597, N14594, N7782, N7866, N7433);
nand NAND4 (N14598, N14593, N4248, N7090, N6367);
or OR3 (N14599, N14591, N2739, N2779);
nor NOR3 (N14600, N14595, N2922, N13077);
nor NOR4 (N14601, N14586, N4762, N1588, N205);
and AND2 (N14602, N14598, N5327);
not NOT1 (N14603, N14599);
and AND4 (N14604, N14579, N8969, N13677, N8223);
xor XOR2 (N14605, N14603, N12598);
or OR2 (N14606, N14602, N3658);
or OR2 (N14607, N14600, N6015);
and AND3 (N14608, N14604, N2593, N10097);
and AND3 (N14609, N14592, N1083, N1129);
buf BUF1 (N14610, N14605);
not NOT1 (N14611, N14609);
or OR3 (N14612, N14597, N3528, N4841);
nand NAND2 (N14613, N14601, N12197);
nor NOR2 (N14614, N14613, N13141);
and AND4 (N14615, N14611, N12288, N11227, N3740);
nor NOR3 (N14616, N14563, N8454, N2664);
buf BUF1 (N14617, N14612);
and AND3 (N14618, N14596, N12285, N1173);
nor NOR3 (N14619, N14616, N7301, N7527);
nor NOR2 (N14620, N14618, N3871);
or OR4 (N14621, N14606, N13817, N8839, N4934);
buf BUF1 (N14622, N14614);
and AND3 (N14623, N14622, N13210, N14618);
nand NAND3 (N14624, N14620, N3360, N4893);
or OR3 (N14625, N14619, N5922, N4546);
and AND3 (N14626, N14610, N14470, N5649);
nand NAND3 (N14627, N14589, N2549, N1056);
and AND2 (N14628, N14623, N8525);
buf BUF1 (N14629, N14628);
and AND2 (N14630, N14626, N6161);
nor NOR4 (N14631, N14625, N10266, N7851, N11217);
not NOT1 (N14632, N14617);
or OR2 (N14633, N14615, N12647);
and AND2 (N14634, N14624, N12283);
and AND2 (N14635, N14607, N7804);
buf BUF1 (N14636, N14632);
buf BUF1 (N14637, N14634);
xor XOR2 (N14638, N14636, N7277);
or OR2 (N14639, N14633, N5176);
buf BUF1 (N14640, N14637);
nor NOR2 (N14641, N14627, N5826);
not NOT1 (N14642, N14629);
not NOT1 (N14643, N14641);
buf BUF1 (N14644, N14640);
buf BUF1 (N14645, N14630);
nand NAND3 (N14646, N14638, N9131, N5014);
nor NOR3 (N14647, N14642, N80, N11991);
nor NOR4 (N14648, N14644, N5795, N2787, N6493);
and AND2 (N14649, N14647, N11859);
and AND3 (N14650, N14621, N7905, N6743);
or OR4 (N14651, N14650, N6728, N13121, N10938);
and AND2 (N14652, N14651, N9693);
or OR4 (N14653, N14608, N7762, N323, N1395);
xor XOR2 (N14654, N14649, N7127);
not NOT1 (N14655, N14635);
or OR2 (N14656, N14654, N11701);
buf BUF1 (N14657, N14639);
buf BUF1 (N14658, N14655);
nor NOR3 (N14659, N14648, N13745, N121);
nand NAND4 (N14660, N14645, N1102, N9815, N1011);
buf BUF1 (N14661, N14646);
buf BUF1 (N14662, N14643);
nor NOR4 (N14663, N14659, N5639, N5713, N4289);
nor NOR3 (N14664, N14661, N11206, N6740);
nand NAND2 (N14665, N14662, N6084);
xor XOR2 (N14666, N14664, N11937);
nor NOR4 (N14667, N14652, N14124, N9599, N9254);
and AND4 (N14668, N14666, N281, N9441, N4152);
buf BUF1 (N14669, N14660);
xor XOR2 (N14670, N14631, N7179);
and AND2 (N14671, N14665, N13917);
not NOT1 (N14672, N14658);
not NOT1 (N14673, N14663);
or OR2 (N14674, N14653, N5385);
buf BUF1 (N14675, N14670);
buf BUF1 (N14676, N14656);
xor XOR2 (N14677, N14667, N11441);
nor NOR3 (N14678, N14669, N857, N11151);
not NOT1 (N14679, N14677);
or OR3 (N14680, N14671, N9132, N5655);
not NOT1 (N14681, N14673);
nand NAND2 (N14682, N14672, N283);
nand NAND4 (N14683, N14668, N11588, N7062, N10622);
nand NAND4 (N14684, N14681, N12546, N8263, N11785);
buf BUF1 (N14685, N14657);
nor NOR3 (N14686, N14680, N11561, N131);
xor XOR2 (N14687, N14682, N617);
buf BUF1 (N14688, N14687);
nand NAND3 (N14689, N14679, N11019, N10669);
not NOT1 (N14690, N14674);
or OR4 (N14691, N14675, N4364, N9251, N9593);
xor XOR2 (N14692, N14691, N13503);
not NOT1 (N14693, N14688);
nand NAND3 (N14694, N14689, N14398, N3946);
xor XOR2 (N14695, N14685, N1979);
xor XOR2 (N14696, N14694, N12344);
buf BUF1 (N14697, N14683);
nor NOR2 (N14698, N14686, N9461);
and AND2 (N14699, N14698, N5545);
or OR2 (N14700, N14676, N1248);
nor NOR3 (N14701, N14695, N9358, N1109);
nand NAND4 (N14702, N14690, N6888, N7705, N14673);
buf BUF1 (N14703, N14692);
nand NAND3 (N14704, N14701, N9490, N11364);
nand NAND2 (N14705, N14703, N3964);
xor XOR2 (N14706, N14704, N9768);
nand NAND4 (N14707, N14697, N5010, N4256, N13579);
not NOT1 (N14708, N14707);
buf BUF1 (N14709, N14684);
xor XOR2 (N14710, N14693, N1236);
and AND4 (N14711, N14678, N11409, N11907, N8317);
not NOT1 (N14712, N14706);
nor NOR3 (N14713, N14711, N2968, N34);
and AND3 (N14714, N14696, N12717, N3491);
not NOT1 (N14715, N14709);
or OR2 (N14716, N14710, N3902);
buf BUF1 (N14717, N14713);
nor NOR2 (N14718, N14714, N4311);
or OR4 (N14719, N14700, N5781, N14090, N13242);
buf BUF1 (N14720, N14717);
nand NAND3 (N14721, N14719, N176, N1581);
nand NAND4 (N14722, N14712, N1347, N11953, N13621);
nand NAND4 (N14723, N14699, N11796, N7236, N12109);
or OR2 (N14724, N14721, N12181);
or OR4 (N14725, N14702, N1270, N13338, N12158);
buf BUF1 (N14726, N14724);
nand NAND3 (N14727, N14722, N11037, N3673);
buf BUF1 (N14728, N14715);
not NOT1 (N14729, N14727);
or OR2 (N14730, N14708, N627);
or OR3 (N14731, N14716, N10169, N12637);
xor XOR2 (N14732, N14730, N12655);
and AND3 (N14733, N14720, N1928, N13549);
or OR3 (N14734, N14733, N3372, N13173);
buf BUF1 (N14735, N14732);
buf BUF1 (N14736, N14734);
buf BUF1 (N14737, N14728);
nor NOR2 (N14738, N14725, N8381);
xor XOR2 (N14739, N14705, N4655);
buf BUF1 (N14740, N14726);
and AND2 (N14741, N14738, N1680);
nand NAND3 (N14742, N14718, N8080, N11282);
buf BUF1 (N14743, N14731);
and AND2 (N14744, N14739, N2082);
buf BUF1 (N14745, N14743);
xor XOR2 (N14746, N14723, N13400);
and AND3 (N14747, N14746, N3385, N1499);
and AND2 (N14748, N14744, N2114);
not NOT1 (N14749, N14736);
or OR4 (N14750, N14737, N13134, N4543, N11539);
xor XOR2 (N14751, N14742, N8254);
xor XOR2 (N14752, N14751, N11430);
and AND4 (N14753, N14735, N3570, N10925, N2825);
and AND2 (N14754, N14740, N5630);
and AND2 (N14755, N14745, N12027);
or OR4 (N14756, N14752, N6285, N3229, N12901);
nor NOR2 (N14757, N14741, N14427);
nand NAND3 (N14758, N14749, N8591, N6058);
not NOT1 (N14759, N14758);
and AND2 (N14760, N14759, N10048);
buf BUF1 (N14761, N14757);
xor XOR2 (N14762, N14755, N9824);
buf BUF1 (N14763, N14747);
and AND3 (N14764, N14762, N2638, N5829);
nor NOR3 (N14765, N14756, N3027, N886);
not NOT1 (N14766, N14753);
nand NAND2 (N14767, N14765, N13623);
or OR4 (N14768, N14764, N12436, N11876, N14683);
and AND2 (N14769, N14760, N7925);
xor XOR2 (N14770, N14761, N3261);
not NOT1 (N14771, N14754);
nor NOR4 (N14772, N14750, N10220, N4458, N11616);
and AND4 (N14773, N14769, N2405, N3890, N7336);
not NOT1 (N14774, N14773);
or OR4 (N14775, N14768, N143, N9937, N10378);
buf BUF1 (N14776, N14774);
not NOT1 (N14777, N14766);
buf BUF1 (N14778, N14771);
buf BUF1 (N14779, N14772);
nand NAND2 (N14780, N14778, N8424);
buf BUF1 (N14781, N14767);
buf BUF1 (N14782, N14776);
xor XOR2 (N14783, N14770, N5842);
nand NAND3 (N14784, N14783, N11712, N3781);
or OR3 (N14785, N14781, N9298, N1606);
and AND3 (N14786, N14763, N2058, N7990);
buf BUF1 (N14787, N14780);
nor NOR4 (N14788, N14785, N2336, N6828, N8211);
xor XOR2 (N14789, N14787, N8280);
not NOT1 (N14790, N14779);
or OR3 (N14791, N14786, N14776, N13565);
nor NOR3 (N14792, N14775, N9476, N12073);
nor NOR4 (N14793, N14748, N2497, N14069, N5924);
xor XOR2 (N14794, N14777, N7963);
and AND2 (N14795, N14792, N5427);
or OR4 (N14796, N14791, N1012, N13541, N5545);
xor XOR2 (N14797, N14789, N673);
and AND3 (N14798, N14729, N9240, N1233);
nand NAND4 (N14799, N14784, N8541, N2049, N8642);
or OR3 (N14800, N14797, N4493, N6614);
nor NOR2 (N14801, N14782, N9690);
nand NAND3 (N14802, N14801, N7657, N1506);
not NOT1 (N14803, N14798);
or OR2 (N14804, N14802, N4083);
nor NOR3 (N14805, N14793, N13839, N2029);
and AND4 (N14806, N14799, N4361, N7971, N10872);
not NOT1 (N14807, N14788);
nand NAND2 (N14808, N14804, N12334);
nor NOR3 (N14809, N14794, N6780, N6155);
not NOT1 (N14810, N14805);
or OR3 (N14811, N14808, N11926, N6562);
xor XOR2 (N14812, N14807, N8026);
nand NAND3 (N14813, N14803, N2668, N14578);
or OR3 (N14814, N14800, N3147, N13022);
xor XOR2 (N14815, N14814, N6016);
and AND3 (N14816, N14812, N6070, N7842);
and AND3 (N14817, N14813, N3679, N2139);
buf BUF1 (N14818, N14806);
nand NAND2 (N14819, N14796, N5830);
xor XOR2 (N14820, N14815, N7291);
xor XOR2 (N14821, N14790, N523);
xor XOR2 (N14822, N14821, N12759);
buf BUF1 (N14823, N14820);
or OR2 (N14824, N14817, N11655);
nand NAND4 (N14825, N14795, N7257, N1286, N12792);
nand NAND3 (N14826, N14818, N3836, N495);
or OR4 (N14827, N14822, N13749, N4965, N2940);
or OR2 (N14828, N14825, N4077);
xor XOR2 (N14829, N14823, N93);
xor XOR2 (N14830, N14819, N12966);
not NOT1 (N14831, N14826);
buf BUF1 (N14832, N14811);
nor NOR2 (N14833, N14829, N2950);
or OR2 (N14834, N14831, N4275);
not NOT1 (N14835, N14809);
nor NOR3 (N14836, N14833, N1145, N9863);
or OR2 (N14837, N14810, N13214);
nand NAND2 (N14838, N14827, N14351);
buf BUF1 (N14839, N14816);
or OR3 (N14840, N14838, N11594, N6890);
xor XOR2 (N14841, N14836, N3845);
nand NAND2 (N14842, N14837, N12806);
not NOT1 (N14843, N14834);
xor XOR2 (N14844, N14842, N990);
and AND4 (N14845, N14828, N4033, N5103, N10180);
nand NAND2 (N14846, N14824, N8811);
or OR2 (N14847, N14845, N8697);
buf BUF1 (N14848, N14835);
not NOT1 (N14849, N14846);
xor XOR2 (N14850, N14847, N10969);
or OR4 (N14851, N14840, N14206, N7985, N12169);
not NOT1 (N14852, N14849);
and AND3 (N14853, N14843, N11520, N10331);
and AND2 (N14854, N14844, N475);
and AND2 (N14855, N14851, N30);
buf BUF1 (N14856, N14852);
buf BUF1 (N14857, N14850);
not NOT1 (N14858, N14830);
nor NOR2 (N14859, N14856, N13997);
nand NAND3 (N14860, N14853, N3953, N10577);
and AND2 (N14861, N14854, N2286);
xor XOR2 (N14862, N14855, N3977);
nor NOR4 (N14863, N14841, N14226, N3499, N14622);
nor NOR4 (N14864, N14861, N12069, N488, N6000);
nor NOR3 (N14865, N14832, N13870, N5974);
not NOT1 (N14866, N14865);
buf BUF1 (N14867, N14839);
nand NAND3 (N14868, N14857, N7583, N4830);
and AND4 (N14869, N14864, N5771, N11099, N10059);
or OR2 (N14870, N14867, N8066);
xor XOR2 (N14871, N14863, N3669);
buf BUF1 (N14872, N14848);
nor NOR4 (N14873, N14859, N6123, N10548, N6159);
and AND3 (N14874, N14870, N6093, N1571);
xor XOR2 (N14875, N14871, N3894);
nor NOR3 (N14876, N14868, N9646, N6706);
not NOT1 (N14877, N14866);
not NOT1 (N14878, N14858);
not NOT1 (N14879, N14862);
buf BUF1 (N14880, N14872);
xor XOR2 (N14881, N14869, N6259);
xor XOR2 (N14882, N14876, N10598);
not NOT1 (N14883, N14878);
xor XOR2 (N14884, N14879, N8721);
or OR4 (N14885, N14877, N8368, N3737, N949);
nand NAND2 (N14886, N14883, N12905);
nand NAND2 (N14887, N14860, N131);
xor XOR2 (N14888, N14873, N8269);
nand NAND3 (N14889, N14875, N4782, N2173);
not NOT1 (N14890, N14885);
buf BUF1 (N14891, N14881);
xor XOR2 (N14892, N14888, N873);
buf BUF1 (N14893, N14882);
nand NAND4 (N14894, N14884, N5441, N12634, N9182);
buf BUF1 (N14895, N14887);
nor NOR2 (N14896, N14895, N3979);
buf BUF1 (N14897, N14890);
buf BUF1 (N14898, N14874);
and AND3 (N14899, N14894, N1474, N5897);
nand NAND4 (N14900, N14893, N9478, N2515, N12491);
buf BUF1 (N14901, N14896);
not NOT1 (N14902, N14886);
not NOT1 (N14903, N14892);
not NOT1 (N14904, N14889);
xor XOR2 (N14905, N14897, N12386);
nand NAND2 (N14906, N14899, N11004);
or OR4 (N14907, N14880, N11953, N13866, N11469);
nand NAND4 (N14908, N14901, N1684, N12295, N11144);
xor XOR2 (N14909, N14905, N6645);
or OR4 (N14910, N14900, N7096, N10589, N6935);
buf BUF1 (N14911, N14910);
buf BUF1 (N14912, N14911);
xor XOR2 (N14913, N14912, N6495);
and AND4 (N14914, N14906, N8141, N3033, N7846);
not NOT1 (N14915, N14908);
nand NAND3 (N14916, N14913, N2823, N1737);
or OR2 (N14917, N14902, N8714);
and AND4 (N14918, N14904, N1531, N14229, N1710);
nand NAND3 (N14919, N14909, N11145, N33);
not NOT1 (N14920, N14915);
nor NOR4 (N14921, N14891, N2915, N11991, N9984);
not NOT1 (N14922, N14921);
nor NOR2 (N14923, N14916, N6531);
nand NAND4 (N14924, N14918, N8000, N5261, N3597);
and AND4 (N14925, N14924, N9418, N1704, N864);
nand NAND2 (N14926, N14923, N1134);
nand NAND2 (N14927, N14917, N34);
buf BUF1 (N14928, N14903);
or OR3 (N14929, N14925, N8641, N9604);
nand NAND4 (N14930, N14928, N1730, N7586, N5283);
not NOT1 (N14931, N14920);
or OR3 (N14932, N14922, N9011, N13865);
and AND3 (N14933, N14926, N8754, N12254);
not NOT1 (N14934, N14927);
or OR3 (N14935, N14933, N12763, N2478);
nand NAND4 (N14936, N14929, N10808, N14349, N11658);
xor XOR2 (N14937, N14930, N6330);
buf BUF1 (N14938, N14935);
xor XOR2 (N14939, N14936, N10688);
xor XOR2 (N14940, N14932, N9359);
buf BUF1 (N14941, N14940);
and AND3 (N14942, N14898, N4606, N14497);
nor NOR3 (N14943, N14907, N14500, N5148);
or OR2 (N14944, N14937, N2765);
nor NOR4 (N14945, N14919, N6506, N2351, N3352);
xor XOR2 (N14946, N14943, N4985);
not NOT1 (N14947, N14942);
not NOT1 (N14948, N14934);
or OR3 (N14949, N14941, N8005, N7624);
buf BUF1 (N14950, N14947);
nor NOR2 (N14951, N14946, N2917);
not NOT1 (N14952, N14944);
not NOT1 (N14953, N14914);
not NOT1 (N14954, N14953);
or OR3 (N14955, N14938, N11005, N14570);
xor XOR2 (N14956, N14948, N12846);
and AND2 (N14957, N14956, N11221);
and AND2 (N14958, N14939, N13332);
xor XOR2 (N14959, N14950, N3862);
xor XOR2 (N14960, N14954, N5193);
buf BUF1 (N14961, N14949);
nor NOR2 (N14962, N14931, N4468);
nand NAND2 (N14963, N14958, N13928);
nor NOR4 (N14964, N14945, N5200, N8293, N7058);
and AND2 (N14965, N14952, N4365);
or OR3 (N14966, N14961, N4723, N10547);
xor XOR2 (N14967, N14965, N14388);
xor XOR2 (N14968, N14957, N12362);
and AND2 (N14969, N14964, N100);
not NOT1 (N14970, N14959);
and AND4 (N14971, N14966, N2018, N11285, N2881);
or OR4 (N14972, N14962, N11773, N4442, N12910);
xor XOR2 (N14973, N14955, N6794);
nand NAND2 (N14974, N14969, N670);
xor XOR2 (N14975, N14970, N10731);
buf BUF1 (N14976, N14968);
nor NOR2 (N14977, N14963, N14963);
and AND2 (N14978, N14975, N1645);
buf BUF1 (N14979, N14971);
buf BUF1 (N14980, N14978);
nand NAND3 (N14981, N14967, N170, N4174);
nor NOR2 (N14982, N14974, N12541);
and AND4 (N14983, N14972, N1064, N8249, N11922);
not NOT1 (N14984, N14960);
buf BUF1 (N14985, N14984);
nor NOR3 (N14986, N14983, N7506, N2415);
buf BUF1 (N14987, N14976);
or OR4 (N14988, N14985, N5810, N12357, N9388);
buf BUF1 (N14989, N14951);
nand NAND4 (N14990, N14986, N8337, N112, N2458);
xor XOR2 (N14991, N14980, N9942);
nand NAND4 (N14992, N14990, N12895, N10983, N6995);
not NOT1 (N14993, N14992);
not NOT1 (N14994, N14977);
nor NOR4 (N14995, N14993, N9843, N9732, N7179);
or OR2 (N14996, N14973, N13089);
nand NAND4 (N14997, N14996, N8286, N8852, N14473);
not NOT1 (N14998, N14997);
and AND3 (N14999, N14995, N9299, N11729);
buf BUF1 (N15000, N14989);
not NOT1 (N15001, N14988);
buf BUF1 (N15002, N14987);
not NOT1 (N15003, N15002);
or OR4 (N15004, N14998, N44, N9715, N9123);
xor XOR2 (N15005, N15000, N3684);
nand NAND3 (N15006, N15001, N3213, N10751);
buf BUF1 (N15007, N15005);
xor XOR2 (N15008, N14981, N7914);
xor XOR2 (N15009, N15008, N3425);
xor XOR2 (N15010, N15007, N6222);
and AND2 (N15011, N15006, N10961);
nand NAND2 (N15012, N14994, N11167);
or OR2 (N15013, N15010, N9246);
and AND4 (N15014, N15003, N13315, N7802, N7059);
nand NAND4 (N15015, N14991, N6688, N7812, N12161);
nand NAND2 (N15016, N14982, N9962);
or OR4 (N15017, N14999, N12833, N8986, N12839);
buf BUF1 (N15018, N14979);
xor XOR2 (N15019, N15009, N8453);
buf BUF1 (N15020, N15011);
and AND4 (N15021, N15017, N2438, N6461, N1059);
not NOT1 (N15022, N15015);
nor NOR3 (N15023, N15004, N3381, N6075);
nor NOR4 (N15024, N15018, N5619, N8918, N898);
xor XOR2 (N15025, N15014, N9420);
nor NOR3 (N15026, N15025, N6114, N13275);
or OR3 (N15027, N15013, N14295, N8562);
nand NAND3 (N15028, N15024, N13872, N3235);
and AND3 (N15029, N15020, N7726, N5151);
xor XOR2 (N15030, N15021, N6429);
or OR3 (N15031, N15029, N5558, N13675);
or OR2 (N15032, N15023, N10794);
xor XOR2 (N15033, N15027, N4641);
nor NOR2 (N15034, N15030, N5948);
xor XOR2 (N15035, N15033, N13713);
or OR3 (N15036, N15019, N6849, N5461);
buf BUF1 (N15037, N15034);
nor NOR4 (N15038, N15028, N148, N8223, N2708);
buf BUF1 (N15039, N15016);
not NOT1 (N15040, N15031);
nand NAND3 (N15041, N15037, N12763, N13437);
and AND4 (N15042, N15012, N8454, N6413, N6740);
nand NAND3 (N15043, N15041, N858, N9896);
buf BUF1 (N15044, N15042);
nor NOR2 (N15045, N15038, N8707);
nor NOR4 (N15046, N15040, N1770, N2908, N8599);
not NOT1 (N15047, N15026);
buf BUF1 (N15048, N15044);
or OR3 (N15049, N15047, N3067, N739);
or OR3 (N15050, N15045, N11974, N8282);
and AND4 (N15051, N15050, N8693, N8418, N3900);
and AND4 (N15052, N15051, N12738, N8583, N473);
or OR4 (N15053, N15032, N10097, N9497, N11096);
xor XOR2 (N15054, N15043, N300);
buf BUF1 (N15055, N15046);
and AND2 (N15056, N15039, N2417);
not NOT1 (N15057, N15048);
and AND2 (N15058, N15053, N6514);
or OR3 (N15059, N15058, N4913, N1448);
nand NAND4 (N15060, N15057, N3342, N5604, N9716);
buf BUF1 (N15061, N15036);
or OR4 (N15062, N15049, N7447, N3746, N3750);
nor NOR3 (N15063, N15062, N4591, N2167);
nand NAND2 (N15064, N15056, N2996);
xor XOR2 (N15065, N15054, N3443);
and AND3 (N15066, N15061, N5436, N11925);
buf BUF1 (N15067, N15052);
not NOT1 (N15068, N15035);
nor NOR2 (N15069, N15065, N11474);
not NOT1 (N15070, N15064);
and AND2 (N15071, N15063, N9033);
xor XOR2 (N15072, N15070, N13429);
nor NOR3 (N15073, N15072, N13166, N10730);
buf BUF1 (N15074, N15059);
nand NAND3 (N15075, N15067, N2436, N3025);
or OR2 (N15076, N15069, N13635);
or OR3 (N15077, N15075, N328, N854);
nand NAND3 (N15078, N15073, N9655, N8019);
xor XOR2 (N15079, N15060, N12016);
and AND2 (N15080, N15022, N13697);
or OR3 (N15081, N15055, N10349, N180);
buf BUF1 (N15082, N15080);
or OR3 (N15083, N15071, N3851, N7667);
buf BUF1 (N15084, N15076);
xor XOR2 (N15085, N15079, N10879);
xor XOR2 (N15086, N15084, N6030);
or OR4 (N15087, N15068, N7348, N5849, N9475);
nand NAND4 (N15088, N15077, N3096, N858, N5080);
buf BUF1 (N15089, N15082);
xor XOR2 (N15090, N15074, N3872);
nand NAND4 (N15091, N15081, N5579, N718, N9076);
xor XOR2 (N15092, N15066, N220);
and AND2 (N15093, N15089, N1366);
nand NAND4 (N15094, N15086, N13705, N2971, N8493);
nor NOR4 (N15095, N15087, N4857, N4688, N13736);
nand NAND3 (N15096, N15094, N4380, N13402);
or OR4 (N15097, N15093, N468, N9340, N3046);
not NOT1 (N15098, N15095);
not NOT1 (N15099, N15098);
not NOT1 (N15100, N15088);
nand NAND3 (N15101, N15085, N12760, N9589);
or OR2 (N15102, N15092, N4232);
nor NOR3 (N15103, N15091, N1446, N14698);
buf BUF1 (N15104, N15078);
buf BUF1 (N15105, N15099);
xor XOR2 (N15106, N15105, N8405);
and AND3 (N15107, N15101, N7815, N2773);
or OR3 (N15108, N15097, N3034, N6095);
or OR4 (N15109, N15102, N8827, N13507, N2652);
or OR3 (N15110, N15096, N5743, N8306);
buf BUF1 (N15111, N15110);
xor XOR2 (N15112, N15106, N9075);
buf BUF1 (N15113, N15109);
nor NOR2 (N15114, N15083, N4690);
and AND3 (N15115, N15108, N358, N12848);
not NOT1 (N15116, N15104);
not NOT1 (N15117, N15111);
and AND2 (N15118, N15116, N12306);
nor NOR4 (N15119, N15090, N13322, N4767, N1608);
not NOT1 (N15120, N15100);
and AND4 (N15121, N15118, N13572, N11580, N1192);
nor NOR4 (N15122, N15117, N2950, N10127, N14889);
xor XOR2 (N15123, N15121, N12171);
or OR3 (N15124, N15103, N6657, N2393);
or OR2 (N15125, N15112, N2358);
and AND2 (N15126, N15124, N9889);
nand NAND4 (N15127, N15114, N13664, N11757, N4982);
and AND2 (N15128, N15113, N7960);
or OR3 (N15129, N15115, N4621, N9346);
nand NAND4 (N15130, N15127, N2847, N307, N8867);
not NOT1 (N15131, N15128);
xor XOR2 (N15132, N15122, N13476);
and AND3 (N15133, N15132, N3386, N14436);
xor XOR2 (N15134, N15130, N11021);
and AND4 (N15135, N15125, N11912, N4217, N9678);
xor XOR2 (N15136, N15107, N6239);
not NOT1 (N15137, N15120);
nor NOR3 (N15138, N15119, N14165, N5780);
or OR3 (N15139, N15123, N14779, N6382);
not NOT1 (N15140, N15137);
not NOT1 (N15141, N15139);
nor NOR4 (N15142, N15136, N11241, N2637, N7831);
and AND3 (N15143, N15129, N10646, N1478);
not NOT1 (N15144, N15126);
not NOT1 (N15145, N15135);
or OR3 (N15146, N15138, N729, N3790);
or OR3 (N15147, N15140, N1354, N5778);
buf BUF1 (N15148, N15131);
and AND4 (N15149, N15147, N4187, N1946, N8517);
xor XOR2 (N15150, N15143, N12955);
or OR2 (N15151, N15146, N12123);
nand NAND4 (N15152, N15149, N5676, N13729, N1373);
buf BUF1 (N15153, N15151);
or OR2 (N15154, N15148, N6087);
xor XOR2 (N15155, N15133, N1188);
and AND4 (N15156, N15152, N3674, N7254, N5302);
xor XOR2 (N15157, N15154, N11750);
nand NAND4 (N15158, N15157, N2146, N12733, N13953);
nor NOR2 (N15159, N15158, N5929);
nand NAND4 (N15160, N15141, N11341, N1342, N13271);
not NOT1 (N15161, N15155);
nor NOR4 (N15162, N15153, N9484, N10791, N12690);
not NOT1 (N15163, N15142);
and AND2 (N15164, N15161, N13138);
or OR4 (N15165, N15134, N1791, N9885, N12113);
xor XOR2 (N15166, N15159, N709);
nor NOR4 (N15167, N15150, N4534, N11154, N1432);
and AND2 (N15168, N15156, N4369);
or OR2 (N15169, N15145, N13452);
nand NAND4 (N15170, N15144, N3112, N12562, N13398);
buf BUF1 (N15171, N15160);
xor XOR2 (N15172, N15170, N3743);
or OR2 (N15173, N15163, N38);
and AND2 (N15174, N15168, N14872);
or OR4 (N15175, N15172, N13351, N2962, N4693);
or OR4 (N15176, N15164, N3637, N14450, N5432);
not NOT1 (N15177, N15169);
not NOT1 (N15178, N15171);
nand NAND2 (N15179, N15165, N14754);
xor XOR2 (N15180, N15167, N1973);
not NOT1 (N15181, N15174);
buf BUF1 (N15182, N15176);
xor XOR2 (N15183, N15162, N9629);
nand NAND2 (N15184, N15181, N8384);
nand NAND3 (N15185, N15184, N8392, N10734);
nor NOR4 (N15186, N15185, N5629, N4159, N4867);
and AND4 (N15187, N15179, N14823, N437, N1986);
and AND2 (N15188, N15166, N8567);
or OR4 (N15189, N15173, N13061, N11226, N10495);
xor XOR2 (N15190, N15187, N1234);
and AND3 (N15191, N15182, N8823, N2058);
buf BUF1 (N15192, N15188);
not NOT1 (N15193, N15177);
xor XOR2 (N15194, N15193, N5210);
nand NAND2 (N15195, N15180, N2635);
nor NOR3 (N15196, N15192, N1768, N10105);
xor XOR2 (N15197, N15189, N5036);
not NOT1 (N15198, N15175);
nand NAND3 (N15199, N15194, N4919, N547);
not NOT1 (N15200, N15183);
buf BUF1 (N15201, N15190);
not NOT1 (N15202, N15197);
not NOT1 (N15203, N15202);
and AND4 (N15204, N15200, N7901, N14314, N5949);
and AND4 (N15205, N15178, N4948, N8246, N10947);
not NOT1 (N15206, N15198);
xor XOR2 (N15207, N15203, N3383);
or OR3 (N15208, N15199, N7635, N6648);
and AND3 (N15209, N15201, N4912, N8283);
xor XOR2 (N15210, N15204, N12374);
nand NAND2 (N15211, N15195, N10283);
nand NAND3 (N15212, N15191, N13183, N5745);
nor NOR3 (N15213, N15211, N7040, N953);
xor XOR2 (N15214, N15207, N582);
nor NOR3 (N15215, N15212, N11458, N2531);
xor XOR2 (N15216, N15196, N2993);
buf BUF1 (N15217, N15206);
xor XOR2 (N15218, N15186, N7578);
nand NAND4 (N15219, N15218, N11044, N3829, N11039);
buf BUF1 (N15220, N15209);
nand NAND4 (N15221, N15213, N8523, N12670, N7578);
nand NAND3 (N15222, N15214, N4547, N10229);
and AND4 (N15223, N15219, N14068, N10744, N8566);
xor XOR2 (N15224, N15215, N613);
not NOT1 (N15225, N15223);
or OR2 (N15226, N15208, N11527);
not NOT1 (N15227, N15224);
nand NAND4 (N15228, N15220, N3482, N14086, N13303);
xor XOR2 (N15229, N15228, N3804);
xor XOR2 (N15230, N15221, N3757);
and AND2 (N15231, N15229, N6411);
xor XOR2 (N15232, N15225, N14728);
xor XOR2 (N15233, N15230, N7733);
or OR2 (N15234, N15233, N6763);
buf BUF1 (N15235, N15217);
buf BUF1 (N15236, N15226);
buf BUF1 (N15237, N15210);
not NOT1 (N15238, N15237);
or OR2 (N15239, N15205, N10248);
nor NOR4 (N15240, N15238, N2558, N11142, N11269);
and AND2 (N15241, N15232, N11643);
nor NOR3 (N15242, N15216, N9466, N7318);
nand NAND3 (N15243, N15236, N2571, N6409);
nand NAND3 (N15244, N15227, N1179, N2055);
nor NOR4 (N15245, N15242, N13826, N13233, N5900);
nand NAND3 (N15246, N15244, N6362, N972);
or OR4 (N15247, N15245, N13944, N7313, N10708);
nor NOR2 (N15248, N15241, N4828);
nor NOR2 (N15249, N15246, N7542);
xor XOR2 (N15250, N15234, N6592);
nor NOR2 (N15251, N15240, N6274);
nor NOR3 (N15252, N15231, N14665, N1107);
not NOT1 (N15253, N15247);
not NOT1 (N15254, N15252);
not NOT1 (N15255, N15250);
not NOT1 (N15256, N15248);
buf BUF1 (N15257, N15249);
nor NOR4 (N15258, N15254, N5123, N2051, N5530);
and AND4 (N15259, N15258, N7754, N3554, N8672);
nor NOR3 (N15260, N15235, N5735, N7664);
nand NAND2 (N15261, N15255, N6658);
buf BUF1 (N15262, N15260);
nand NAND3 (N15263, N15251, N4466, N7206);
or OR4 (N15264, N15256, N13787, N7258, N260);
nand NAND3 (N15265, N15264, N5674, N7143);
xor XOR2 (N15266, N15262, N14452);
and AND3 (N15267, N15222, N11145, N14814);
or OR2 (N15268, N15243, N5463);
not NOT1 (N15269, N15268);
xor XOR2 (N15270, N15263, N12294);
xor XOR2 (N15271, N15257, N2583);
and AND4 (N15272, N15259, N4961, N5827, N5878);
nand NAND2 (N15273, N15271, N6089);
nand NAND2 (N15274, N15253, N15206);
nor NOR3 (N15275, N15270, N14234, N10116);
nor NOR3 (N15276, N15272, N3625, N7446);
xor XOR2 (N15277, N15276, N8559);
and AND3 (N15278, N15261, N11193, N9581);
or OR2 (N15279, N15266, N789);
xor XOR2 (N15280, N15269, N14734);
xor XOR2 (N15281, N15279, N6151);
nor NOR3 (N15282, N15265, N4611, N10706);
or OR3 (N15283, N15273, N2174, N12308);
not NOT1 (N15284, N15283);
nor NOR3 (N15285, N15267, N14271, N10967);
and AND4 (N15286, N15274, N289, N4594, N7825);
xor XOR2 (N15287, N15282, N11772);
buf BUF1 (N15288, N15286);
not NOT1 (N15289, N15281);
or OR3 (N15290, N15289, N11981, N4313);
or OR3 (N15291, N15290, N9501, N2757);
xor XOR2 (N15292, N15285, N11962);
nor NOR2 (N15293, N15284, N6485);
buf BUF1 (N15294, N15287);
buf BUF1 (N15295, N15275);
or OR2 (N15296, N15288, N1941);
not NOT1 (N15297, N15293);
and AND4 (N15298, N15291, N1846, N4418, N14545);
xor XOR2 (N15299, N15277, N7626);
and AND2 (N15300, N15292, N9794);
and AND3 (N15301, N15239, N10904, N3282);
and AND2 (N15302, N15294, N11065);
buf BUF1 (N15303, N15300);
xor XOR2 (N15304, N15296, N11266);
nor NOR4 (N15305, N15297, N5398, N12564, N14751);
nand NAND4 (N15306, N15302, N11628, N13634, N3416);
buf BUF1 (N15307, N15278);
not NOT1 (N15308, N15306);
xor XOR2 (N15309, N15298, N5204);
nand NAND4 (N15310, N15307, N4656, N8323, N12546);
xor XOR2 (N15311, N15295, N13054);
nand NAND2 (N15312, N15311, N7432);
nand NAND2 (N15313, N15310, N6294);
xor XOR2 (N15314, N15304, N14887);
not NOT1 (N15315, N15308);
nand NAND2 (N15316, N15280, N5499);
not NOT1 (N15317, N15305);
xor XOR2 (N15318, N15301, N5591);
or OR3 (N15319, N15315, N634, N5455);
buf BUF1 (N15320, N15299);
nor NOR3 (N15321, N15320, N9534, N9957);
buf BUF1 (N15322, N15313);
buf BUF1 (N15323, N15319);
nor NOR3 (N15324, N15321, N2644, N11100);
nand NAND3 (N15325, N15323, N2721, N6411);
buf BUF1 (N15326, N15309);
or OR3 (N15327, N15324, N9958, N3295);
and AND3 (N15328, N15314, N657, N8088);
nand NAND4 (N15329, N15303, N11460, N9957, N3635);
nor NOR2 (N15330, N15326, N3838);
or OR3 (N15331, N15325, N11034, N15013);
nor NOR4 (N15332, N15317, N3918, N4543, N12317);
nand NAND3 (N15333, N15329, N15084, N3309);
nand NAND3 (N15334, N15318, N7278, N7671);
or OR3 (N15335, N15328, N10568, N11912);
nand NAND2 (N15336, N15333, N12821);
not NOT1 (N15337, N15322);
nand NAND2 (N15338, N15335, N8155);
or OR3 (N15339, N15334, N9167, N11426);
nor NOR4 (N15340, N15316, N8291, N11642, N7783);
and AND2 (N15341, N15312, N5417);
nand NAND3 (N15342, N15330, N1800, N6718);
buf BUF1 (N15343, N15342);
or OR3 (N15344, N15340, N12428, N2571);
nand NAND2 (N15345, N15337, N1670);
xor XOR2 (N15346, N15331, N6533);
buf BUF1 (N15347, N15338);
not NOT1 (N15348, N15344);
or OR3 (N15349, N15343, N14633, N6521);
buf BUF1 (N15350, N15332);
and AND4 (N15351, N15350, N11455, N5287, N8452);
nand NAND4 (N15352, N15346, N4492, N2713, N14283);
nor NOR3 (N15353, N15327, N1655, N1733);
not NOT1 (N15354, N15341);
nand NAND3 (N15355, N15353, N11511, N13844);
xor XOR2 (N15356, N15349, N7073);
nor NOR3 (N15357, N15352, N11922, N10383);
or OR4 (N15358, N15336, N10951, N8222, N8764);
or OR4 (N15359, N15355, N11940, N12637, N1989);
or OR2 (N15360, N15358, N6050);
nand NAND2 (N15361, N15348, N6612);
not NOT1 (N15362, N15357);
or OR3 (N15363, N15351, N1276, N6037);
and AND3 (N15364, N15347, N4649, N12553);
xor XOR2 (N15365, N15356, N12040);
or OR2 (N15366, N15365, N6153);
nand NAND3 (N15367, N15360, N6967, N10197);
or OR3 (N15368, N15362, N8513, N5195);
not NOT1 (N15369, N15364);
not NOT1 (N15370, N15345);
or OR3 (N15371, N15359, N9572, N1495);
nor NOR2 (N15372, N15354, N7981);
nor NOR2 (N15373, N15370, N14540);
or OR2 (N15374, N15363, N13619);
nand NAND2 (N15375, N15372, N141);
xor XOR2 (N15376, N15367, N7775);
or OR2 (N15377, N15375, N1474);
not NOT1 (N15378, N15339);
xor XOR2 (N15379, N15371, N13381);
not NOT1 (N15380, N15368);
nand NAND3 (N15381, N15378, N3325, N11282);
and AND3 (N15382, N15369, N9695, N13104);
or OR2 (N15383, N15374, N11691);
not NOT1 (N15384, N15380);
xor XOR2 (N15385, N15382, N1652);
buf BUF1 (N15386, N15377);
buf BUF1 (N15387, N15379);
buf BUF1 (N15388, N15383);
or OR3 (N15389, N15385, N14503, N8114);
xor XOR2 (N15390, N15386, N2400);
buf BUF1 (N15391, N15384);
or OR3 (N15392, N15381, N11616, N13518);
nor NOR3 (N15393, N15392, N10853, N4504);
xor XOR2 (N15394, N15391, N6462);
or OR4 (N15395, N15388, N7484, N7495, N737);
not NOT1 (N15396, N15393);
nand NAND2 (N15397, N15376, N9454);
nand NAND4 (N15398, N15397, N15159, N13572, N10998);
and AND2 (N15399, N15361, N1420);
and AND2 (N15400, N15366, N11301);
xor XOR2 (N15401, N15394, N12936);
nand NAND4 (N15402, N15400, N8279, N6965, N8176);
buf BUF1 (N15403, N15373);
or OR3 (N15404, N15398, N12234, N13658);
nand NAND3 (N15405, N15402, N11035, N14609);
or OR2 (N15406, N15389, N14001);
xor XOR2 (N15407, N15406, N11329);
nand NAND2 (N15408, N15403, N14619);
xor XOR2 (N15409, N15396, N14536);
or OR3 (N15410, N15387, N1096, N9184);
or OR3 (N15411, N15407, N3970, N1464);
xor XOR2 (N15412, N15404, N9008);
xor XOR2 (N15413, N15395, N7069);
or OR2 (N15414, N15405, N11398);
and AND2 (N15415, N15414, N8702);
nor NOR2 (N15416, N15399, N7017);
buf BUF1 (N15417, N15412);
buf BUF1 (N15418, N15401);
nor NOR2 (N15419, N15417, N6863);
not NOT1 (N15420, N15409);
nand NAND4 (N15421, N15418, N8966, N3551, N4946);
and AND3 (N15422, N15419, N6604, N12524);
buf BUF1 (N15423, N15422);
buf BUF1 (N15424, N15421);
or OR3 (N15425, N15413, N13907, N15029);
nor NOR4 (N15426, N15408, N9113, N13141, N69);
nand NAND2 (N15427, N15416, N5948);
not NOT1 (N15428, N15390);
nand NAND2 (N15429, N15423, N9521);
and AND4 (N15430, N15420, N6309, N3777, N4232);
and AND4 (N15431, N15425, N13420, N11700, N194);
xor XOR2 (N15432, N15428, N14900);
nor NOR2 (N15433, N15424, N13267);
xor XOR2 (N15434, N15426, N235);
and AND4 (N15435, N15427, N7935, N13163, N6226);
buf BUF1 (N15436, N15429);
nand NAND2 (N15437, N15432, N412);
not NOT1 (N15438, N15431);
nor NOR2 (N15439, N15434, N8194);
and AND3 (N15440, N15430, N526, N12115);
buf BUF1 (N15441, N15437);
not NOT1 (N15442, N15441);
or OR3 (N15443, N15411, N3782, N5508);
or OR4 (N15444, N15435, N6760, N4088, N2960);
not NOT1 (N15445, N15439);
buf BUF1 (N15446, N15445);
buf BUF1 (N15447, N15436);
or OR3 (N15448, N15446, N8332, N6535);
nor NOR4 (N15449, N15447, N9030, N7868, N14891);
not NOT1 (N15450, N15449);
and AND3 (N15451, N15433, N14592, N1377);
xor XOR2 (N15452, N15450, N8131);
xor XOR2 (N15453, N15440, N6235);
nand NAND4 (N15454, N15443, N5823, N10410, N11943);
not NOT1 (N15455, N15438);
nand NAND2 (N15456, N15444, N6184);
nand NAND3 (N15457, N15451, N5941, N2241);
nor NOR3 (N15458, N15455, N11890, N8356);
nand NAND2 (N15459, N15456, N8344);
nor NOR3 (N15460, N15454, N6833, N1163);
not NOT1 (N15461, N15410);
or OR2 (N15462, N15453, N10269);
not NOT1 (N15463, N15460);
and AND3 (N15464, N15459, N3123, N905);
buf BUF1 (N15465, N15462);
or OR3 (N15466, N15457, N6395, N6186);
or OR3 (N15467, N15458, N8520, N10387);
and AND2 (N15468, N15467, N12982);
and AND4 (N15469, N15452, N1735, N1902, N6189);
or OR2 (N15470, N15466, N1948);
or OR2 (N15471, N15469, N9884);
nor NOR2 (N15472, N15470, N1866);
and AND3 (N15473, N15463, N2201, N7088);
or OR4 (N15474, N15471, N11424, N11825, N12177);
nor NOR4 (N15475, N15472, N14197, N1019, N7799);
nor NOR3 (N15476, N15442, N13362, N4732);
nor NOR3 (N15477, N15448, N6265, N13079);
buf BUF1 (N15478, N15415);
nand NAND4 (N15479, N15476, N12467, N4423, N3297);
xor XOR2 (N15480, N15478, N305);
buf BUF1 (N15481, N15479);
nor NOR4 (N15482, N15481, N10775, N1467, N10411);
xor XOR2 (N15483, N15464, N817);
or OR3 (N15484, N15477, N8294, N14872);
buf BUF1 (N15485, N15474);
and AND2 (N15486, N15461, N13154);
nor NOR2 (N15487, N15484, N2533);
not NOT1 (N15488, N15483);
buf BUF1 (N15489, N15473);
or OR4 (N15490, N15482, N10925, N1377, N1101);
and AND2 (N15491, N15480, N5220);
xor XOR2 (N15492, N15491, N15323);
not NOT1 (N15493, N15492);
and AND2 (N15494, N15465, N15321);
not NOT1 (N15495, N15489);
nand NAND2 (N15496, N15486, N14044);
nand NAND2 (N15497, N15488, N13481);
or OR2 (N15498, N15475, N13310);
not NOT1 (N15499, N15495);
nor NOR2 (N15500, N15498, N8182);
not NOT1 (N15501, N15468);
not NOT1 (N15502, N15500);
nor NOR3 (N15503, N15485, N11989, N995);
nor NOR3 (N15504, N15497, N939, N6685);
nand NAND4 (N15505, N15496, N12, N9796, N12043);
nor NOR4 (N15506, N15501, N4, N7121, N7419);
nand NAND4 (N15507, N15504, N2854, N6528, N9376);
not NOT1 (N15508, N15494);
nand NAND2 (N15509, N15487, N7417);
buf BUF1 (N15510, N15507);
nand NAND2 (N15511, N15508, N12896);
nor NOR4 (N15512, N15509, N4786, N10042, N4588);
or OR3 (N15513, N15511, N2684, N4993);
nor NOR2 (N15514, N15493, N12384);
or OR4 (N15515, N15505, N12433, N3009, N5872);
nor NOR3 (N15516, N15490, N165, N1615);
nand NAND4 (N15517, N15515, N11268, N2222, N3411);
nand NAND3 (N15518, N15513, N6057, N3562);
and AND3 (N15519, N15518, N5466, N7842);
or OR2 (N15520, N15510, N11454);
or OR3 (N15521, N15506, N5855, N5238);
not NOT1 (N15522, N15503);
nor NOR2 (N15523, N15521, N6926);
or OR3 (N15524, N15517, N4259, N15477);
not NOT1 (N15525, N15512);
and AND2 (N15526, N15525, N9182);
or OR2 (N15527, N15502, N8008);
not NOT1 (N15528, N15522);
or OR3 (N15529, N15526, N2227, N2992);
nand NAND2 (N15530, N15514, N12483);
not NOT1 (N15531, N15516);
xor XOR2 (N15532, N15519, N3593);
and AND3 (N15533, N15499, N11266, N13038);
and AND3 (N15534, N15533, N13284, N9889);
xor XOR2 (N15535, N15531, N7908);
buf BUF1 (N15536, N15527);
xor XOR2 (N15537, N15528, N6998);
xor XOR2 (N15538, N15523, N11822);
xor XOR2 (N15539, N15538, N9138);
buf BUF1 (N15540, N15534);
nor NOR2 (N15541, N15535, N3365);
nor NOR4 (N15542, N15539, N8057, N7902, N14854);
nand NAND2 (N15543, N15532, N5825);
nand NAND3 (N15544, N15541, N11004, N14499);
and AND4 (N15545, N15542, N2263, N12696, N9126);
nand NAND3 (N15546, N15524, N3751, N3932);
buf BUF1 (N15547, N15543);
nor NOR3 (N15548, N15537, N13035, N8776);
and AND2 (N15549, N15529, N3680);
buf BUF1 (N15550, N15545);
nor NOR4 (N15551, N15540, N10800, N765, N4307);
not NOT1 (N15552, N15548);
not NOT1 (N15553, N15550);
not NOT1 (N15554, N15530);
nand NAND4 (N15555, N15546, N6840, N14069, N3152);
nand NAND2 (N15556, N15536, N14164);
nor NOR3 (N15557, N15520, N8041, N13831);
and AND2 (N15558, N15554, N5283);
xor XOR2 (N15559, N15557, N2341);
nand NAND4 (N15560, N15551, N3844, N14597, N13015);
xor XOR2 (N15561, N15556, N7009);
buf BUF1 (N15562, N15560);
and AND2 (N15563, N15553, N3615);
not NOT1 (N15564, N15559);
and AND4 (N15565, N15558, N12575, N2471, N4975);
not NOT1 (N15566, N15562);
and AND3 (N15567, N15564, N11220, N4240);
or OR3 (N15568, N15549, N10697, N6049);
or OR2 (N15569, N15561, N3202);
nand NAND4 (N15570, N15568, N2949, N14093, N8304);
xor XOR2 (N15571, N15552, N7414);
xor XOR2 (N15572, N15567, N1733);
not NOT1 (N15573, N15565);
nor NOR3 (N15574, N15571, N3635, N2926);
buf BUF1 (N15575, N15573);
and AND3 (N15576, N15572, N4728, N3744);
xor XOR2 (N15577, N15566, N9276);
and AND2 (N15578, N15575, N74);
nor NOR4 (N15579, N15576, N14199, N9319, N9562);
buf BUF1 (N15580, N15563);
not NOT1 (N15581, N15570);
or OR3 (N15582, N15544, N3963, N13378);
xor XOR2 (N15583, N15547, N11397);
or OR2 (N15584, N15579, N14320);
buf BUF1 (N15585, N15580);
xor XOR2 (N15586, N15582, N4968);
or OR4 (N15587, N15581, N8662, N8667, N7661);
nor NOR3 (N15588, N15583, N5585, N11902);
nand NAND4 (N15589, N15578, N5246, N9306, N8336);
nand NAND4 (N15590, N15589, N6260, N1405, N2683);
buf BUF1 (N15591, N15588);
or OR2 (N15592, N15577, N14663);
and AND2 (N15593, N15587, N4631);
nor NOR3 (N15594, N15585, N11657, N14252);
nand NAND3 (N15595, N15555, N3549, N8912);
and AND2 (N15596, N15586, N14514);
not NOT1 (N15597, N15574);
nand NAND3 (N15598, N15592, N7741, N8706);
nand NAND4 (N15599, N15595, N4560, N12985, N3662);
nor NOR3 (N15600, N15594, N9536, N2811);
nor NOR3 (N15601, N15593, N13449, N2754);
or OR4 (N15602, N15591, N6714, N987, N15145);
xor XOR2 (N15603, N15590, N3133);
not NOT1 (N15604, N15600);
and AND2 (N15605, N15598, N754);
nor NOR3 (N15606, N15601, N15374, N13954);
and AND2 (N15607, N15606, N1773);
nand NAND2 (N15608, N15584, N8942);
and AND2 (N15609, N15605, N5739);
xor XOR2 (N15610, N15609, N6896);
or OR3 (N15611, N15599, N846, N6273);
and AND3 (N15612, N15611, N4354, N8177);
nand NAND3 (N15613, N15603, N8296, N7698);
xor XOR2 (N15614, N15613, N609);
buf BUF1 (N15615, N15608);
not NOT1 (N15616, N15607);
and AND2 (N15617, N15612, N13837);
xor XOR2 (N15618, N15617, N9603);
nand NAND3 (N15619, N15618, N14246, N587);
or OR4 (N15620, N15610, N13118, N3001, N12132);
or OR4 (N15621, N15614, N14120, N5502, N12012);
or OR4 (N15622, N15597, N7533, N9249, N10057);
xor XOR2 (N15623, N15619, N10000);
and AND3 (N15624, N15621, N1585, N11386);
or OR2 (N15625, N15616, N6620);
not NOT1 (N15626, N15624);
nand NAND3 (N15627, N15615, N6148, N9529);
nand NAND3 (N15628, N15569, N1858, N6494);
buf BUF1 (N15629, N15622);
buf BUF1 (N15630, N15627);
not NOT1 (N15631, N15625);
nand NAND2 (N15632, N15602, N4264);
or OR3 (N15633, N15620, N651, N14090);
and AND3 (N15634, N15629, N6946, N9740);
nor NOR2 (N15635, N15596, N12577);
nand NAND2 (N15636, N15631, N10482);
and AND2 (N15637, N15630, N7260);
buf BUF1 (N15638, N15633);
xor XOR2 (N15639, N15637, N9799);
nand NAND4 (N15640, N15636, N8809, N6576, N11687);
or OR2 (N15641, N15628, N7782);
xor XOR2 (N15642, N15626, N5678);
and AND4 (N15643, N15641, N3610, N763, N7311);
buf BUF1 (N15644, N15623);
nor NOR3 (N15645, N15604, N12324, N13403);
or OR3 (N15646, N15635, N2895, N10826);
xor XOR2 (N15647, N15632, N4577);
xor XOR2 (N15648, N15639, N6866);
xor XOR2 (N15649, N15634, N8409);
nand NAND2 (N15650, N15638, N14171);
buf BUF1 (N15651, N15644);
or OR3 (N15652, N15645, N2192, N1325);
nand NAND3 (N15653, N15650, N9898, N14472);
and AND2 (N15654, N15649, N114);
buf BUF1 (N15655, N15647);
and AND4 (N15656, N15651, N1848, N14289, N6607);
nand NAND2 (N15657, N15648, N14836);
buf BUF1 (N15658, N15653);
not NOT1 (N15659, N15656);
xor XOR2 (N15660, N15642, N766);
buf BUF1 (N15661, N15660);
not NOT1 (N15662, N15646);
and AND4 (N15663, N15655, N9249, N15399, N9611);
nor NOR2 (N15664, N15657, N6896);
buf BUF1 (N15665, N15662);
xor XOR2 (N15666, N15661, N8886);
buf BUF1 (N15667, N15643);
xor XOR2 (N15668, N15664, N9202);
buf BUF1 (N15669, N15666);
buf BUF1 (N15670, N15654);
nor NOR3 (N15671, N15667, N10060, N5841);
nor NOR2 (N15672, N15663, N14767);
nor NOR3 (N15673, N15668, N8953, N147);
nand NAND4 (N15674, N15672, N121, N3505, N14738);
not NOT1 (N15675, N15671);
not NOT1 (N15676, N15673);
xor XOR2 (N15677, N15669, N4414);
not NOT1 (N15678, N15676);
nor NOR2 (N15679, N15675, N7944);
xor XOR2 (N15680, N15670, N7287);
nor NOR2 (N15681, N15652, N11938);
nor NOR4 (N15682, N15679, N14459, N5310, N6391);
or OR4 (N15683, N15682, N9836, N9903, N2847);
not NOT1 (N15684, N15658);
xor XOR2 (N15685, N15683, N4153);
nand NAND3 (N15686, N15659, N14074, N12993);
nor NOR3 (N15687, N15680, N15164, N1547);
nand NAND2 (N15688, N15686, N13056);
nor NOR3 (N15689, N15685, N12842, N15264);
or OR4 (N15690, N15681, N12546, N13887, N3235);
buf BUF1 (N15691, N15674);
not NOT1 (N15692, N15688);
not NOT1 (N15693, N15687);
buf BUF1 (N15694, N15693);
and AND3 (N15695, N15690, N11199, N9353);
and AND3 (N15696, N15692, N1301, N15110);
and AND4 (N15697, N15677, N8302, N5689, N5800);
nand NAND4 (N15698, N15684, N859, N11265, N4420);
not NOT1 (N15699, N15696);
buf BUF1 (N15700, N15665);
not NOT1 (N15701, N15698);
not NOT1 (N15702, N15700);
nor NOR2 (N15703, N15678, N6944);
or OR3 (N15704, N15689, N1106, N2050);
xor XOR2 (N15705, N15704, N4421);
or OR2 (N15706, N15640, N9364);
or OR4 (N15707, N15701, N3150, N9121, N7941);
or OR4 (N15708, N15695, N9818, N6429, N9530);
nand NAND4 (N15709, N15705, N14832, N11619, N12905);
buf BUF1 (N15710, N15697);
and AND3 (N15711, N15699, N1341, N5236);
buf BUF1 (N15712, N15710);
nand NAND3 (N15713, N15706, N11894, N11935);
buf BUF1 (N15714, N15691);
buf BUF1 (N15715, N15707);
xor XOR2 (N15716, N15713, N11978);
nor NOR4 (N15717, N15714, N8969, N9818, N2936);
buf BUF1 (N15718, N15702);
or OR4 (N15719, N15712, N10600, N1357, N5831);
xor XOR2 (N15720, N15719, N10890);
buf BUF1 (N15721, N15711);
buf BUF1 (N15722, N15716);
xor XOR2 (N15723, N15718, N5376);
or OR2 (N15724, N15717, N3431);
nand NAND4 (N15725, N15724, N12473, N10955, N2189);
not NOT1 (N15726, N15722);
nand NAND2 (N15727, N15708, N9300);
nor NOR3 (N15728, N15726, N1781, N1500);
nor NOR4 (N15729, N15720, N7619, N14663, N12994);
and AND3 (N15730, N15723, N7668, N10960);
and AND3 (N15731, N15727, N9420, N13467);
and AND3 (N15732, N15731, N14971, N4806);
nand NAND2 (N15733, N15703, N824);
and AND2 (N15734, N15728, N1402);
nand NAND4 (N15735, N15694, N6460, N1309, N7751);
buf BUF1 (N15736, N15709);
or OR3 (N15737, N15721, N5465, N4201);
nor NOR3 (N15738, N15737, N13800, N6235);
and AND2 (N15739, N15729, N4592);
not NOT1 (N15740, N15725);
buf BUF1 (N15741, N15730);
nand NAND4 (N15742, N15733, N4022, N7964, N9234);
nor NOR3 (N15743, N15732, N15005, N4142);
nand NAND4 (N15744, N15736, N469, N2651, N7676);
nand NAND4 (N15745, N15735, N4323, N9243, N2117);
nand NAND2 (N15746, N15741, N2270);
and AND2 (N15747, N15743, N11320);
nor NOR3 (N15748, N15739, N1250, N14585);
or OR2 (N15749, N15748, N13053);
not NOT1 (N15750, N15744);
and AND3 (N15751, N15746, N7828, N5682);
not NOT1 (N15752, N15715);
or OR4 (N15753, N15745, N7394, N112, N15329);
xor XOR2 (N15754, N15747, N6596);
xor XOR2 (N15755, N15749, N6274);
nor NOR4 (N15756, N15754, N5640, N10093, N11908);
nand NAND3 (N15757, N15755, N707, N817);
xor XOR2 (N15758, N15751, N14400);
buf BUF1 (N15759, N15742);
xor XOR2 (N15760, N15759, N9349);
nand NAND4 (N15761, N15752, N11812, N4295, N7943);
and AND4 (N15762, N15761, N1584, N6100, N8030);
or OR2 (N15763, N15758, N4864);
buf BUF1 (N15764, N15756);
nand NAND3 (N15765, N15760, N5999, N15340);
not NOT1 (N15766, N15757);
nor NOR3 (N15767, N15765, N14290, N9886);
nand NAND3 (N15768, N15753, N7647, N3451);
and AND2 (N15769, N15740, N12335);
xor XOR2 (N15770, N15734, N1307);
xor XOR2 (N15771, N15768, N3502);
or OR3 (N15772, N15769, N10692, N5017);
and AND4 (N15773, N15766, N5071, N1606, N10565);
nor NOR2 (N15774, N15772, N9861);
nor NOR4 (N15775, N15767, N10817, N844, N11785);
not NOT1 (N15776, N15762);
not NOT1 (N15777, N15771);
not NOT1 (N15778, N15750);
xor XOR2 (N15779, N15763, N1719);
not NOT1 (N15780, N15779);
buf BUF1 (N15781, N15738);
xor XOR2 (N15782, N15777, N4087);
and AND3 (N15783, N15780, N10730, N4208);
xor XOR2 (N15784, N15775, N7815);
nand NAND2 (N15785, N15782, N9164);
nor NOR3 (N15786, N15774, N1615, N1603);
and AND3 (N15787, N15770, N3077, N15344);
nor NOR4 (N15788, N15773, N8928, N4265, N8058);
or OR4 (N15789, N15781, N7816, N5443, N637);
and AND4 (N15790, N15776, N9003, N13488, N11526);
and AND3 (N15791, N15788, N2950, N4965);
or OR3 (N15792, N15786, N7212, N7255);
or OR3 (N15793, N15789, N10256, N9077);
xor XOR2 (N15794, N15764, N11890);
and AND4 (N15795, N15784, N6141, N12149, N13154);
not NOT1 (N15796, N15787);
xor XOR2 (N15797, N15785, N2734);
xor XOR2 (N15798, N15797, N8257);
xor XOR2 (N15799, N15783, N14305);
nor NOR2 (N15800, N15796, N9761);
xor XOR2 (N15801, N15790, N8412);
not NOT1 (N15802, N15778);
or OR4 (N15803, N15799, N1239, N14863, N10645);
nand NAND3 (N15804, N15793, N6918, N15198);
and AND3 (N15805, N15794, N3084, N1245);
nand NAND4 (N15806, N15791, N431, N9742, N3030);
not NOT1 (N15807, N15805);
not NOT1 (N15808, N15800);
or OR2 (N15809, N15792, N2729);
not NOT1 (N15810, N15795);
not NOT1 (N15811, N15798);
buf BUF1 (N15812, N15804);
nand NAND3 (N15813, N15802, N4535, N15673);
buf BUF1 (N15814, N15813);
or OR2 (N15815, N15811, N4810);
buf BUF1 (N15816, N15814);
nand NAND3 (N15817, N15806, N9464, N7098);
nand NAND4 (N15818, N15817, N6058, N1926, N4665);
buf BUF1 (N15819, N15809);
xor XOR2 (N15820, N15808, N594);
and AND2 (N15821, N15803, N15036);
xor XOR2 (N15822, N15820, N9643);
and AND2 (N15823, N15807, N3106);
nor NOR4 (N15824, N15822, N4980, N2195, N11925);
buf BUF1 (N15825, N15818);
not NOT1 (N15826, N15812);
xor XOR2 (N15827, N15824, N5107);
not NOT1 (N15828, N15815);
nand NAND3 (N15829, N15821, N7980, N678);
buf BUF1 (N15830, N15827);
xor XOR2 (N15831, N15823, N2712);
or OR4 (N15832, N15831, N14949, N7368, N11099);
nor NOR3 (N15833, N15832, N924, N6330);
xor XOR2 (N15834, N15830, N9938);
buf BUF1 (N15835, N15825);
buf BUF1 (N15836, N15816);
not NOT1 (N15837, N15801);
not NOT1 (N15838, N15833);
and AND2 (N15839, N15834, N6205);
or OR3 (N15840, N15836, N14110, N114);
nand NAND4 (N15841, N15826, N8953, N13748, N1059);
xor XOR2 (N15842, N15829, N3061);
and AND3 (N15843, N15828, N307, N8298);
not NOT1 (N15844, N15838);
xor XOR2 (N15845, N15842, N486);
nor NOR2 (N15846, N15837, N5667);
xor XOR2 (N15847, N15810, N242);
buf BUF1 (N15848, N15845);
buf BUF1 (N15849, N15847);
nor NOR3 (N15850, N15844, N6838, N14739);
xor XOR2 (N15851, N15839, N13601);
or OR4 (N15852, N15846, N3109, N342, N1108);
not NOT1 (N15853, N15850);
not NOT1 (N15854, N15852);
not NOT1 (N15855, N15849);
nand NAND2 (N15856, N15843, N810);
not NOT1 (N15857, N15848);
or OR2 (N15858, N15851, N9830);
buf BUF1 (N15859, N15856);
xor XOR2 (N15860, N15841, N11965);
nor NOR2 (N15861, N15840, N11910);
not NOT1 (N15862, N15858);
or OR3 (N15863, N15860, N11997, N1787);
nand NAND3 (N15864, N15835, N15494, N6783);
buf BUF1 (N15865, N15857);
xor XOR2 (N15866, N15859, N6817);
buf BUF1 (N15867, N15853);
nor NOR3 (N15868, N15865, N1727, N15469);
buf BUF1 (N15869, N15861);
or OR3 (N15870, N15868, N3976, N12164);
buf BUF1 (N15871, N15855);
buf BUF1 (N15872, N15854);
nor NOR3 (N15873, N15863, N15255, N4780);
or OR4 (N15874, N15864, N15536, N3449, N1386);
buf BUF1 (N15875, N15862);
nand NAND2 (N15876, N15869, N12119);
and AND2 (N15877, N15866, N4367);
and AND2 (N15878, N15871, N7834);
or OR2 (N15879, N15872, N5554);
or OR2 (N15880, N15819, N8981);
nand NAND2 (N15881, N15874, N8007);
nor NOR3 (N15882, N15879, N12240, N12515);
or OR2 (N15883, N15880, N1769);
not NOT1 (N15884, N15873);
nor NOR3 (N15885, N15876, N10926, N12113);
nor NOR3 (N15886, N15878, N2735, N8429);
or OR4 (N15887, N15882, N1316, N9987, N11308);
and AND3 (N15888, N15886, N2676, N332);
buf BUF1 (N15889, N15881);
not NOT1 (N15890, N15883);
nor NOR2 (N15891, N15884, N295);
or OR4 (N15892, N15887, N5834, N2427, N4508);
or OR4 (N15893, N15885, N1696, N2453, N8702);
nor NOR2 (N15894, N15877, N4365);
not NOT1 (N15895, N15892);
nand NAND3 (N15896, N15888, N158, N8477);
not NOT1 (N15897, N15895);
nand NAND4 (N15898, N15867, N13136, N4001, N11);
not NOT1 (N15899, N15898);
nand NAND3 (N15900, N15889, N14319, N15109);
nor NOR3 (N15901, N15893, N10706, N1524);
buf BUF1 (N15902, N15875);
xor XOR2 (N15903, N15900, N13242);
and AND4 (N15904, N15901, N2720, N13349, N12543);
nor NOR2 (N15905, N15894, N13011);
xor XOR2 (N15906, N15896, N2028);
nand NAND4 (N15907, N15870, N6948, N12077, N15622);
not NOT1 (N15908, N15905);
not NOT1 (N15909, N15906);
nor NOR2 (N15910, N15899, N9480);
nand NAND2 (N15911, N15897, N2203);
and AND3 (N15912, N15902, N12395, N3147);
not NOT1 (N15913, N15910);
and AND2 (N15914, N15911, N8906);
not NOT1 (N15915, N15908);
xor XOR2 (N15916, N15904, N654);
buf BUF1 (N15917, N15912);
nand NAND4 (N15918, N15909, N15472, N3151, N1426);
buf BUF1 (N15919, N15913);
nand NAND3 (N15920, N15914, N15286, N99);
xor XOR2 (N15921, N15918, N1900);
or OR4 (N15922, N15915, N12096, N7588, N14881);
xor XOR2 (N15923, N15920, N13288);
buf BUF1 (N15924, N15917);
nand NAND2 (N15925, N15916, N14444);
and AND4 (N15926, N15924, N13586, N3554, N3751);
xor XOR2 (N15927, N15891, N11944);
or OR3 (N15928, N15890, N12955, N12040);
xor XOR2 (N15929, N15907, N10355);
nand NAND4 (N15930, N15929, N8785, N1818, N295);
or OR4 (N15931, N15923, N12098, N3351, N4059);
or OR4 (N15932, N15927, N3523, N11161, N15599);
not NOT1 (N15933, N15928);
buf BUF1 (N15934, N15919);
buf BUF1 (N15935, N15932);
buf BUF1 (N15936, N15933);
buf BUF1 (N15937, N15903);
xor XOR2 (N15938, N15936, N4149);
or OR3 (N15939, N15938, N14151, N8773);
xor XOR2 (N15940, N15937, N8907);
nand NAND3 (N15941, N15940, N9038, N3502);
nand NAND2 (N15942, N15934, N13100);
nand NAND2 (N15943, N15941, N2913);
nand NAND2 (N15944, N15921, N8362);
and AND3 (N15945, N15942, N4925, N3229);
nor NOR2 (N15946, N15935, N9936);
buf BUF1 (N15947, N15926);
or OR2 (N15948, N15931, N10319);
or OR2 (N15949, N15922, N13323);
buf BUF1 (N15950, N15939);
or OR4 (N15951, N15944, N7481, N5347, N12151);
nand NAND2 (N15952, N15943, N1944);
or OR2 (N15953, N15950, N12825);
buf BUF1 (N15954, N15948);
or OR3 (N15955, N15930, N1268, N15637);
not NOT1 (N15956, N15947);
or OR4 (N15957, N15946, N11781, N2801, N247);
not NOT1 (N15958, N15953);
xor XOR2 (N15959, N15925, N5237);
nand NAND3 (N15960, N15959, N13973, N5121);
nand NAND3 (N15961, N15958, N5321, N10633);
buf BUF1 (N15962, N15955);
xor XOR2 (N15963, N15951, N2178);
buf BUF1 (N15964, N15949);
xor XOR2 (N15965, N15963, N5680);
xor XOR2 (N15966, N15965, N1044);
nor NOR3 (N15967, N15964, N4048, N15733);
nand NAND3 (N15968, N15966, N6796, N6880);
not NOT1 (N15969, N15945);
buf BUF1 (N15970, N15967);
xor XOR2 (N15971, N15968, N3673);
nand NAND2 (N15972, N15952, N516);
and AND2 (N15973, N15962, N1691);
not NOT1 (N15974, N15957);
nand NAND3 (N15975, N15961, N2232, N4956);
nand NAND4 (N15976, N15973, N6700, N15134, N2784);
not NOT1 (N15977, N15960);
and AND2 (N15978, N15977, N7271);
not NOT1 (N15979, N15972);
or OR3 (N15980, N15956, N10113, N9510);
nand NAND4 (N15981, N15969, N7667, N13508, N599);
buf BUF1 (N15982, N15979);
xor XOR2 (N15983, N15971, N6227);
nand NAND4 (N15984, N15974, N14084, N10762, N2468);
xor XOR2 (N15985, N15975, N10196);
nand NAND4 (N15986, N15980, N2507, N10024, N12909);
not NOT1 (N15987, N15976);
or OR4 (N15988, N15978, N23, N10518, N12383);
nand NAND2 (N15989, N15987, N11684);
nand NAND3 (N15990, N15970, N10171, N9647);
and AND4 (N15991, N15988, N2997, N5516, N7005);
buf BUF1 (N15992, N15985);
xor XOR2 (N15993, N15990, N10106);
buf BUF1 (N15994, N15981);
buf BUF1 (N15995, N15984);
nor NOR3 (N15996, N15994, N7191, N8331);
xor XOR2 (N15997, N15983, N6744);
and AND2 (N15998, N15989, N7470);
xor XOR2 (N15999, N15954, N2516);
nor NOR4 (N16000, N15995, N1714, N1936, N15248);
not NOT1 (N16001, N15992);
nand NAND3 (N16002, N15998, N3085, N14424);
xor XOR2 (N16003, N15997, N2462);
xor XOR2 (N16004, N15999, N6423);
buf BUF1 (N16005, N15991);
and AND2 (N16006, N15986, N2657);
buf BUF1 (N16007, N15993);
nor NOR4 (N16008, N16000, N8469, N8045, N11445);
or OR4 (N16009, N15982, N8476, N13778, N13901);
nor NOR4 (N16010, N16007, N14636, N11673, N2807);
and AND2 (N16011, N16005, N5713);
or OR2 (N16012, N16004, N10622);
nor NOR2 (N16013, N15996, N8911);
not NOT1 (N16014, N16008);
and AND2 (N16015, N16001, N13236);
buf BUF1 (N16016, N16015);
or OR2 (N16017, N16012, N3637);
buf BUF1 (N16018, N16006);
not NOT1 (N16019, N16016);
nand NAND3 (N16020, N16002, N14552, N7649);
not NOT1 (N16021, N16017);
and AND3 (N16022, N16011, N13260, N2270);
or OR2 (N16023, N16010, N11497);
buf BUF1 (N16024, N16003);
nand NAND3 (N16025, N16018, N7142, N667);
nor NOR4 (N16026, N16009, N11121, N7519, N12800);
buf BUF1 (N16027, N16020);
xor XOR2 (N16028, N16014, N2104);
nor NOR4 (N16029, N16025, N1726, N5846, N972);
and AND3 (N16030, N16027, N7401, N486);
and AND2 (N16031, N16021, N2235);
nor NOR3 (N16032, N16024, N8363, N287);
nand NAND3 (N16033, N16026, N14954, N5452);
nand NAND3 (N16034, N16029, N14629, N7711);
xor XOR2 (N16035, N16032, N7377);
or OR3 (N16036, N16023, N8610, N7266);
and AND2 (N16037, N16013, N1816);
not NOT1 (N16038, N16019);
and AND4 (N16039, N16035, N9063, N2105, N2697);
and AND2 (N16040, N16034, N10036);
and AND2 (N16041, N16028, N1609);
and AND2 (N16042, N16039, N2259);
xor XOR2 (N16043, N16031, N12156);
buf BUF1 (N16044, N16037);
buf BUF1 (N16045, N16036);
nor NOR3 (N16046, N16022, N5051, N13788);
not NOT1 (N16047, N16038);
nor NOR3 (N16048, N16030, N9818, N6280);
not NOT1 (N16049, N16042);
not NOT1 (N16050, N16046);
buf BUF1 (N16051, N16040);
xor XOR2 (N16052, N16033, N6074);
not NOT1 (N16053, N16048);
nand NAND4 (N16054, N16050, N13572, N8444, N277);
nand NAND4 (N16055, N16051, N3787, N2811, N5005);
not NOT1 (N16056, N16044);
or OR4 (N16057, N16052, N2913, N13130, N6069);
or OR3 (N16058, N16056, N7590, N1998);
buf BUF1 (N16059, N16049);
or OR4 (N16060, N16047, N15710, N2164, N3580);
or OR4 (N16061, N16053, N14735, N5067, N9181);
not NOT1 (N16062, N16061);
not NOT1 (N16063, N16060);
and AND2 (N16064, N16043, N7965);
xor XOR2 (N16065, N16064, N5497);
and AND2 (N16066, N16065, N12768);
xor XOR2 (N16067, N16063, N3953);
nand NAND2 (N16068, N16066, N14077);
or OR2 (N16069, N16045, N3204);
xor XOR2 (N16070, N16062, N3744);
not NOT1 (N16071, N16058);
xor XOR2 (N16072, N16068, N2680);
nand NAND3 (N16073, N16071, N6635, N4999);
and AND3 (N16074, N16059, N2160, N8127);
buf BUF1 (N16075, N16041);
nand NAND4 (N16076, N16075, N7868, N1373, N10515);
nor NOR2 (N16077, N16072, N11631);
not NOT1 (N16078, N16054);
nand NAND4 (N16079, N16069, N7215, N13109, N1536);
nand NAND3 (N16080, N16067, N9554, N1903);
and AND2 (N16081, N16076, N10775);
and AND3 (N16082, N16081, N15823, N5868);
xor XOR2 (N16083, N16074, N12541);
buf BUF1 (N16084, N16083);
nand NAND4 (N16085, N16084, N4366, N2737, N12673);
xor XOR2 (N16086, N16055, N4544);
nor NOR4 (N16087, N16057, N8179, N13370, N16019);
nand NAND3 (N16088, N16087, N4165, N7002);
buf BUF1 (N16089, N16080);
nor NOR3 (N16090, N16089, N16029, N4798);
nand NAND2 (N16091, N16085, N10201);
not NOT1 (N16092, N16070);
not NOT1 (N16093, N16073);
buf BUF1 (N16094, N16093);
nor NOR2 (N16095, N16078, N1443);
nand NAND4 (N16096, N16090, N12904, N8800, N1470);
nand NAND4 (N16097, N16077, N14946, N7164, N12721);
or OR4 (N16098, N16091, N12980, N1999, N7609);
nor NOR3 (N16099, N16092, N3793, N8744);
nand NAND4 (N16100, N16082, N9192, N15722, N14816);
or OR3 (N16101, N16086, N11821, N1178);
and AND4 (N16102, N16094, N11737, N11049, N11016);
and AND3 (N16103, N16088, N9176, N12007);
and AND4 (N16104, N16102, N12451, N6386, N5291);
xor XOR2 (N16105, N16101, N7875);
nand NAND3 (N16106, N16098, N1823, N7214);
or OR2 (N16107, N16106, N12791);
nor NOR4 (N16108, N16100, N13766, N4872, N13164);
or OR2 (N16109, N16108, N3826);
and AND3 (N16110, N16105, N7035, N4317);
nor NOR2 (N16111, N16104, N9996);
not NOT1 (N16112, N16099);
xor XOR2 (N16113, N16079, N1552);
xor XOR2 (N16114, N16109, N15636);
nand NAND3 (N16115, N16097, N15690, N11927);
and AND2 (N16116, N16110, N10721);
xor XOR2 (N16117, N16116, N4375);
nand NAND2 (N16118, N16111, N9574);
nor NOR2 (N16119, N16113, N9518);
nand NAND2 (N16120, N16112, N390);
nand NAND4 (N16121, N16103, N10243, N16001, N9578);
buf BUF1 (N16122, N16117);
nand NAND2 (N16123, N16118, N11481);
nor NOR4 (N16124, N16095, N10297, N15654, N6791);
xor XOR2 (N16125, N16107, N14651);
or OR3 (N16126, N16123, N2558, N3646);
or OR4 (N16127, N16096, N1808, N10064, N5525);
not NOT1 (N16128, N16127);
or OR3 (N16129, N16125, N9146, N8788);
xor XOR2 (N16130, N16128, N3099);
nor NOR3 (N16131, N16120, N3559, N4957);
buf BUF1 (N16132, N16119);
xor XOR2 (N16133, N16130, N8151);
xor XOR2 (N16134, N16121, N14182);
nand NAND4 (N16135, N16126, N4923, N14932, N6286);
or OR3 (N16136, N16129, N12701, N3947);
nand NAND4 (N16137, N16136, N8948, N13005, N2700);
nor NOR3 (N16138, N16131, N14423, N4696);
nor NOR4 (N16139, N16135, N13547, N13836, N3636);
nor NOR4 (N16140, N16124, N12480, N13636, N10816);
or OR3 (N16141, N16137, N6405, N4049);
buf BUF1 (N16142, N16114);
nor NOR2 (N16143, N16138, N6827);
buf BUF1 (N16144, N16133);
or OR3 (N16145, N16141, N13810, N3098);
buf BUF1 (N16146, N16145);
xor XOR2 (N16147, N16143, N7288);
nand NAND4 (N16148, N16146, N5309, N6410, N8076);
xor XOR2 (N16149, N16115, N11475);
and AND3 (N16150, N16132, N13971, N14952);
nand NAND3 (N16151, N16148, N12853, N14380);
nand NAND2 (N16152, N16147, N9101);
not NOT1 (N16153, N16142);
nor NOR3 (N16154, N16140, N3972, N2961);
nor NOR2 (N16155, N16151, N10289);
and AND3 (N16156, N16154, N4552, N9268);
xor XOR2 (N16157, N16155, N14278);
not NOT1 (N16158, N16150);
and AND3 (N16159, N16122, N6602, N642);
and AND3 (N16160, N16156, N9912, N15241);
or OR2 (N16161, N16134, N13476);
or OR3 (N16162, N16157, N6109, N6271);
or OR4 (N16163, N16139, N2201, N11208, N2001);
xor XOR2 (N16164, N16159, N15822);
buf BUF1 (N16165, N16153);
nand NAND3 (N16166, N16161, N10483, N5041);
not NOT1 (N16167, N16152);
xor XOR2 (N16168, N16160, N11454);
buf BUF1 (N16169, N16144);
buf BUF1 (N16170, N16158);
not NOT1 (N16171, N16165);
xor XOR2 (N16172, N16166, N6467);
buf BUF1 (N16173, N16167);
nor NOR2 (N16174, N16173, N9106);
nor NOR2 (N16175, N16163, N9812);
or OR2 (N16176, N16169, N11624);
nor NOR4 (N16177, N16168, N6908, N7444, N13922);
nor NOR4 (N16178, N16162, N13298, N12784, N3770);
xor XOR2 (N16179, N16177, N1487);
nand NAND3 (N16180, N16176, N11875, N7410);
xor XOR2 (N16181, N16180, N266);
nand NAND2 (N16182, N16174, N9509);
xor XOR2 (N16183, N16171, N16074);
nand NAND4 (N16184, N16183, N5840, N12049, N5264);
and AND2 (N16185, N16170, N11389);
and AND4 (N16186, N16184, N3794, N11172, N8004);
nand NAND2 (N16187, N16149, N12781);
xor XOR2 (N16188, N16179, N15709);
and AND2 (N16189, N16164, N11235);
or OR3 (N16190, N16175, N3211, N1470);
or OR2 (N16191, N16190, N16014);
not NOT1 (N16192, N16181);
nor NOR4 (N16193, N16185, N9900, N618, N8672);
not NOT1 (N16194, N16182);
or OR2 (N16195, N16189, N4770);
buf BUF1 (N16196, N16187);
xor XOR2 (N16197, N16193, N13241);
nand NAND4 (N16198, N16188, N8935, N1105, N651);
nor NOR2 (N16199, N16178, N13462);
nor NOR3 (N16200, N16196, N9179, N9187);
and AND4 (N16201, N16186, N304, N9369, N10566);
and AND4 (N16202, N16191, N9934, N12045, N5057);
xor XOR2 (N16203, N16195, N8399);
or OR4 (N16204, N16194, N3939, N1529, N14198);
and AND4 (N16205, N16204, N15275, N6228, N288);
buf BUF1 (N16206, N16192);
not NOT1 (N16207, N16198);
buf BUF1 (N16208, N16202);
or OR3 (N16209, N16206, N13295, N15616);
and AND3 (N16210, N16199, N5761, N10519);
and AND2 (N16211, N16201, N14129);
or OR4 (N16212, N16200, N1725, N1100, N8053);
and AND2 (N16213, N16210, N441);
xor XOR2 (N16214, N16203, N2620);
nand NAND3 (N16215, N16211, N5794, N12957);
nand NAND3 (N16216, N16213, N1161, N4855);
nor NOR4 (N16217, N16216, N15529, N9206, N12946);
nand NAND3 (N16218, N16197, N11666, N956);
and AND3 (N16219, N16209, N7843, N547);
nor NOR2 (N16220, N16207, N1757);
and AND2 (N16221, N16172, N5074);
not NOT1 (N16222, N16221);
nand NAND3 (N16223, N16215, N7022, N543);
not NOT1 (N16224, N16214);
or OR2 (N16225, N16205, N5627);
nand NAND4 (N16226, N16217, N12751, N14441, N1777);
and AND3 (N16227, N16219, N6035, N7132);
nand NAND3 (N16228, N16223, N5843, N2680);
buf BUF1 (N16229, N16224);
buf BUF1 (N16230, N16208);
nand NAND3 (N16231, N16225, N11376, N2423);
buf BUF1 (N16232, N16220);
nand NAND2 (N16233, N16222, N5902);
buf BUF1 (N16234, N16226);
buf BUF1 (N16235, N16231);
and AND2 (N16236, N16228, N7158);
buf BUF1 (N16237, N16236);
buf BUF1 (N16238, N16237);
nand NAND4 (N16239, N16238, N876, N3734, N2057);
nor NOR3 (N16240, N16227, N2318, N11673);
buf BUF1 (N16241, N16218);
or OR2 (N16242, N16239, N7018);
nand NAND3 (N16243, N16230, N11105, N1761);
nor NOR2 (N16244, N16232, N9176);
and AND3 (N16245, N16242, N5251, N14143);
and AND4 (N16246, N16235, N8785, N7238, N51);
xor XOR2 (N16247, N16246, N6412);
and AND3 (N16248, N16245, N14619, N6727);
nor NOR4 (N16249, N16247, N9096, N11691, N11260);
nand NAND4 (N16250, N16244, N315, N1083, N4872);
buf BUF1 (N16251, N16233);
not NOT1 (N16252, N16250);
or OR2 (N16253, N16241, N9071);
or OR4 (N16254, N16243, N14788, N7507, N13970);
nand NAND3 (N16255, N16240, N1901, N11187);
and AND3 (N16256, N16249, N11273, N3920);
xor XOR2 (N16257, N16254, N2302);
or OR2 (N16258, N16255, N2672);
xor XOR2 (N16259, N16257, N6590);
nor NOR3 (N16260, N16252, N11670, N4179);
and AND2 (N16261, N16253, N3139);
buf BUF1 (N16262, N16251);
and AND2 (N16263, N16256, N2917);
nand NAND3 (N16264, N16262, N10615, N1255);
buf BUF1 (N16265, N16258);
xor XOR2 (N16266, N16259, N1950);
and AND3 (N16267, N16260, N7903, N3842);
or OR2 (N16268, N16212, N6395);
nor NOR3 (N16269, N16234, N13834, N3895);
nand NAND2 (N16270, N16265, N9026);
nand NAND4 (N16271, N16268, N11290, N7279, N12250);
nand NAND4 (N16272, N16261, N4071, N14951, N3248);
nor NOR2 (N16273, N16263, N172);
buf BUF1 (N16274, N16272);
buf BUF1 (N16275, N16270);
nor NOR3 (N16276, N16274, N3942, N8705);
or OR3 (N16277, N16271, N2070, N4081);
xor XOR2 (N16278, N16276, N4305);
nand NAND4 (N16279, N16269, N16092, N12498, N2060);
nor NOR2 (N16280, N16273, N4708);
and AND2 (N16281, N16278, N13372);
not NOT1 (N16282, N16281);
xor XOR2 (N16283, N16279, N3052);
nor NOR3 (N16284, N16283, N14422, N13777);
not NOT1 (N16285, N16248);
and AND2 (N16286, N16275, N1214);
buf BUF1 (N16287, N16285);
or OR2 (N16288, N16266, N6540);
nand NAND3 (N16289, N16280, N15366, N9577);
xor XOR2 (N16290, N16286, N10689);
not NOT1 (N16291, N16288);
and AND2 (N16292, N16284, N2101);
not NOT1 (N16293, N16277);
not NOT1 (N16294, N16229);
nor NOR4 (N16295, N16267, N868, N8258, N9094);
and AND3 (N16296, N16291, N6388, N10381);
xor XOR2 (N16297, N16294, N1334);
not NOT1 (N16298, N16287);
buf BUF1 (N16299, N16296);
and AND2 (N16300, N16264, N12088);
not NOT1 (N16301, N16300);
or OR4 (N16302, N16282, N6783, N9681, N15667);
not NOT1 (N16303, N16299);
buf BUF1 (N16304, N16289);
nor NOR3 (N16305, N16292, N4866, N12646);
nor NOR2 (N16306, N16304, N11780);
not NOT1 (N16307, N16303);
nor NOR4 (N16308, N16307, N2427, N10090, N6018);
xor XOR2 (N16309, N16301, N4155);
nand NAND2 (N16310, N16297, N11145);
buf BUF1 (N16311, N16293);
and AND4 (N16312, N16309, N13719, N9773, N5457);
and AND4 (N16313, N16295, N7049, N99, N5943);
nor NOR3 (N16314, N16298, N3648, N2407);
xor XOR2 (N16315, N16312, N9692);
or OR3 (N16316, N16302, N9070, N11577);
nand NAND3 (N16317, N16313, N14499, N1701);
buf BUF1 (N16318, N16316);
nor NOR3 (N16319, N16317, N3394, N8300);
not NOT1 (N16320, N16311);
nor NOR2 (N16321, N16310, N14605);
buf BUF1 (N16322, N16308);
buf BUF1 (N16323, N16290);
not NOT1 (N16324, N16315);
nand NAND2 (N16325, N16314, N10731);
nand NAND4 (N16326, N16324, N8890, N92, N6775);
nand NAND2 (N16327, N16321, N6255);
nand NAND2 (N16328, N16305, N14745);
not NOT1 (N16329, N16325);
and AND4 (N16330, N16328, N10977, N5449, N9932);
not NOT1 (N16331, N16306);
or OR4 (N16332, N16330, N7927, N14604, N14872);
not NOT1 (N16333, N16327);
nand NAND3 (N16334, N16320, N2190, N11705);
xor XOR2 (N16335, N16331, N14532);
nor NOR4 (N16336, N16318, N14353, N13145, N13916);
nand NAND2 (N16337, N16332, N266);
or OR2 (N16338, N16334, N8451);
not NOT1 (N16339, N16336);
buf BUF1 (N16340, N16323);
or OR4 (N16341, N16319, N11310, N10385, N16323);
and AND2 (N16342, N16333, N14299);
and AND3 (N16343, N16322, N4834, N14801);
nor NOR4 (N16344, N16339, N12904, N6311, N7331);
buf BUF1 (N16345, N16341);
nand NAND3 (N16346, N16342, N11363, N13892);
or OR3 (N16347, N16335, N13787, N2341);
buf BUF1 (N16348, N16329);
and AND3 (N16349, N16338, N69, N15803);
buf BUF1 (N16350, N16346);
not NOT1 (N16351, N16326);
or OR4 (N16352, N16343, N3717, N448, N42);
nor NOR3 (N16353, N16352, N198, N7648);
nor NOR3 (N16354, N16340, N4758, N2582);
xor XOR2 (N16355, N16337, N15873);
and AND4 (N16356, N16345, N13373, N7895, N15909);
or OR2 (N16357, N16355, N3175);
xor XOR2 (N16358, N16353, N4709);
or OR3 (N16359, N16357, N14965, N1566);
nor NOR4 (N16360, N16351, N5642, N10697, N5260);
and AND3 (N16361, N16356, N820, N5560);
not NOT1 (N16362, N16348);
or OR3 (N16363, N16344, N11476, N13713);
and AND4 (N16364, N16354, N5373, N8620, N6386);
xor XOR2 (N16365, N16358, N11193);
nor NOR2 (N16366, N16349, N2485);
xor XOR2 (N16367, N16360, N15236);
or OR3 (N16368, N16359, N1693, N13743);
or OR4 (N16369, N16362, N14136, N9069, N142);
buf BUF1 (N16370, N16365);
nor NOR2 (N16371, N16364, N9218);
or OR4 (N16372, N16363, N14031, N8095, N11436);
nor NOR3 (N16373, N16369, N16034, N312);
buf BUF1 (N16374, N16370);
not NOT1 (N16375, N16350);
xor XOR2 (N16376, N16373, N849);
buf BUF1 (N16377, N16371);
not NOT1 (N16378, N16372);
nand NAND2 (N16379, N16361, N6257);
nand NAND4 (N16380, N16367, N15888, N5687, N11890);
buf BUF1 (N16381, N16379);
nand NAND2 (N16382, N16381, N1753);
xor XOR2 (N16383, N16368, N11366);
xor XOR2 (N16384, N16383, N10988);
or OR4 (N16385, N16376, N8509, N10089, N3396);
not NOT1 (N16386, N16375);
xor XOR2 (N16387, N16347, N7121);
xor XOR2 (N16388, N16387, N1403);
buf BUF1 (N16389, N16384);
buf BUF1 (N16390, N16380);
not NOT1 (N16391, N16389);
buf BUF1 (N16392, N16386);
and AND3 (N16393, N16374, N15650, N1601);
buf BUF1 (N16394, N16391);
nand NAND2 (N16395, N16388, N12970);
buf BUF1 (N16396, N16382);
not NOT1 (N16397, N16395);
not NOT1 (N16398, N16378);
buf BUF1 (N16399, N16377);
or OR2 (N16400, N16394, N6169);
and AND2 (N16401, N16392, N11459);
nand NAND3 (N16402, N16366, N16241, N4254);
and AND3 (N16403, N16385, N15973, N8067);
nand NAND3 (N16404, N16393, N10076, N822);
and AND2 (N16405, N16401, N6343);
xor XOR2 (N16406, N16402, N10366);
xor XOR2 (N16407, N16406, N14128);
and AND3 (N16408, N16397, N12966, N6070);
buf BUF1 (N16409, N16403);
buf BUF1 (N16410, N16405);
nand NAND2 (N16411, N16390, N44);
nand NAND2 (N16412, N16400, N6311);
xor XOR2 (N16413, N16408, N3633);
or OR2 (N16414, N16407, N104);
and AND2 (N16415, N16404, N13366);
nor NOR3 (N16416, N16409, N8494, N7994);
or OR3 (N16417, N16396, N10432, N6884);
xor XOR2 (N16418, N16411, N10619);
and AND2 (N16419, N16418, N11759);
and AND4 (N16420, N16413, N6172, N10396, N1195);
and AND2 (N16421, N16398, N16379);
nor NOR2 (N16422, N16399, N10383);
or OR3 (N16423, N16412, N13322, N5908);
or OR4 (N16424, N16420, N12782, N3772, N12883);
not NOT1 (N16425, N16410);
nand NAND2 (N16426, N16419, N2584);
or OR2 (N16427, N16422, N9424);
not NOT1 (N16428, N16416);
and AND3 (N16429, N16414, N1763, N2352);
nand NAND2 (N16430, N16424, N5685);
xor XOR2 (N16431, N16429, N11026);
and AND3 (N16432, N16425, N9469, N4225);
nand NAND2 (N16433, N16430, N3475);
nor NOR2 (N16434, N16426, N13098);
not NOT1 (N16435, N16417);
or OR2 (N16436, N16415, N7058);
nor NOR4 (N16437, N16423, N160, N15038, N3251);
and AND4 (N16438, N16428, N2891, N3209, N4880);
nand NAND2 (N16439, N16431, N6058);
nand NAND3 (N16440, N16432, N6665, N14008);
nor NOR3 (N16441, N16436, N7315, N4384);
and AND2 (N16442, N16439, N8907);
nand NAND2 (N16443, N16434, N9319);
or OR4 (N16444, N16421, N7697, N16395, N7157);
nor NOR2 (N16445, N16444, N12713);
and AND4 (N16446, N16441, N7012, N7240, N7019);
or OR3 (N16447, N16440, N12428, N8);
or OR2 (N16448, N16435, N14588);
nor NOR2 (N16449, N16448, N11369);
or OR4 (N16450, N16427, N8449, N4442, N585);
xor XOR2 (N16451, N16433, N540);
or OR2 (N16452, N16447, N5777);
and AND3 (N16453, N16449, N15656, N11703);
and AND3 (N16454, N16446, N2408, N473);
nand NAND4 (N16455, N16452, N451, N12670, N997);
xor XOR2 (N16456, N16437, N12420);
nor NOR2 (N16457, N16451, N14915);
not NOT1 (N16458, N16453);
not NOT1 (N16459, N16458);
nor NOR3 (N16460, N16442, N2770, N14477);
or OR3 (N16461, N16455, N10022, N7819);
nand NAND3 (N16462, N16459, N3853, N4727);
or OR4 (N16463, N16462, N13505, N12983, N12513);
buf BUF1 (N16464, N16438);
nor NOR2 (N16465, N16443, N5774);
xor XOR2 (N16466, N16457, N14187);
buf BUF1 (N16467, N16445);
buf BUF1 (N16468, N16465);
not NOT1 (N16469, N16466);
not NOT1 (N16470, N16467);
and AND4 (N16471, N16463, N2749, N15968, N5215);
nor NOR2 (N16472, N16470, N993);
buf BUF1 (N16473, N16469);
buf BUF1 (N16474, N16472);
nor NOR2 (N16475, N16473, N9991);
and AND3 (N16476, N16456, N14901, N6792);
buf BUF1 (N16477, N16460);
or OR2 (N16478, N16475, N3516);
not NOT1 (N16479, N16461);
or OR2 (N16480, N16464, N8799);
nor NOR3 (N16481, N16450, N9462, N3957);
and AND2 (N16482, N16454, N370);
xor XOR2 (N16483, N16481, N8536);
or OR2 (N16484, N16468, N1857);
xor XOR2 (N16485, N16477, N8278);
buf BUF1 (N16486, N16480);
nor NOR4 (N16487, N16471, N6391, N6194, N7256);
and AND3 (N16488, N16479, N13347, N14644);
xor XOR2 (N16489, N16486, N1693);
not NOT1 (N16490, N16488);
not NOT1 (N16491, N16474);
nand NAND2 (N16492, N16485, N4734);
nor NOR2 (N16493, N16492, N3377);
nand NAND4 (N16494, N16490, N3504, N14924, N3171);
buf BUF1 (N16495, N16478);
and AND3 (N16496, N16484, N1996, N16265);
buf BUF1 (N16497, N16489);
or OR4 (N16498, N16493, N9957, N3007, N12376);
and AND2 (N16499, N16483, N9128);
or OR2 (N16500, N16499, N1015);
xor XOR2 (N16501, N16491, N8712);
nor NOR3 (N16502, N16496, N8653, N14690);
or OR4 (N16503, N16498, N13417, N4999, N7980);
xor XOR2 (N16504, N16494, N5733);
nor NOR4 (N16505, N16503, N7086, N13025, N10232);
nor NOR3 (N16506, N16482, N2366, N15834);
or OR2 (N16507, N16502, N9651);
not NOT1 (N16508, N16501);
nor NOR3 (N16509, N16500, N1562, N5645);
not NOT1 (N16510, N16508);
nand NAND3 (N16511, N16509, N4702, N4780);
nor NOR4 (N16512, N16510, N9417, N12100, N2244);
xor XOR2 (N16513, N16495, N14744);
nand NAND4 (N16514, N16507, N309, N9831, N13525);
buf BUF1 (N16515, N16505);
not NOT1 (N16516, N16506);
buf BUF1 (N16517, N16487);
buf BUF1 (N16518, N16514);
nand NAND4 (N16519, N16518, N6591, N13920, N2395);
nand NAND4 (N16520, N16513, N15994, N2344, N3985);
nand NAND4 (N16521, N16519, N10923, N8398, N364);
and AND2 (N16522, N16516, N11043);
xor XOR2 (N16523, N16512, N9031);
nand NAND2 (N16524, N16504, N11887);
xor XOR2 (N16525, N16517, N7932);
nor NOR3 (N16526, N16524, N10534, N8939);
and AND2 (N16527, N16520, N14934);
not NOT1 (N16528, N16526);
nor NOR3 (N16529, N16515, N5209, N14407);
or OR2 (N16530, N16525, N5715);
buf BUF1 (N16531, N16497);
nand NAND2 (N16532, N16531, N10108);
buf BUF1 (N16533, N16522);
nand NAND2 (N16534, N16523, N5878);
or OR4 (N16535, N16521, N3891, N10920, N16036);
or OR2 (N16536, N16528, N3850);
buf BUF1 (N16537, N16534);
or OR3 (N16538, N16535, N8374, N5023);
xor XOR2 (N16539, N16527, N5986);
xor XOR2 (N16540, N16533, N12022);
or OR4 (N16541, N16536, N13863, N8542, N12855);
nor NOR3 (N16542, N16476, N3039, N9478);
buf BUF1 (N16543, N16541);
or OR3 (N16544, N16537, N4227, N2614);
nand NAND2 (N16545, N16543, N2322);
not NOT1 (N16546, N16529);
xor XOR2 (N16547, N16540, N6881);
nand NAND2 (N16548, N16538, N6063);
and AND2 (N16549, N16546, N13265);
xor XOR2 (N16550, N16545, N4195);
or OR2 (N16551, N16532, N1571);
nand NAND2 (N16552, N16530, N2244);
xor XOR2 (N16553, N16551, N473);
and AND2 (N16554, N16553, N257);
nand NAND2 (N16555, N16552, N15905);
not NOT1 (N16556, N16544);
or OR3 (N16557, N16550, N11938, N14553);
not NOT1 (N16558, N16542);
buf BUF1 (N16559, N16555);
not NOT1 (N16560, N16547);
and AND2 (N16561, N16511, N7105);
nand NAND3 (N16562, N16557, N9037, N11574);
and AND3 (N16563, N16558, N3664, N11463);
and AND4 (N16564, N16559, N7457, N5095, N3907);
nor NOR4 (N16565, N16560, N2207, N12818, N5806);
buf BUF1 (N16566, N16561);
and AND3 (N16567, N16563, N9097, N15427);
and AND4 (N16568, N16556, N15355, N4578, N16135);
buf BUF1 (N16569, N16567);
nor NOR3 (N16570, N16566, N2915, N13010);
nand NAND2 (N16571, N16548, N2392);
xor XOR2 (N16572, N16554, N387);
buf BUF1 (N16573, N16569);
and AND2 (N16574, N16570, N14187);
nand NAND3 (N16575, N16565, N9549, N5504);
or OR3 (N16576, N16568, N2784, N1111);
and AND3 (N16577, N16562, N14085, N14958);
xor XOR2 (N16578, N16575, N9825);
and AND2 (N16579, N16571, N6387);
not NOT1 (N16580, N16579);
not NOT1 (N16581, N16564);
xor XOR2 (N16582, N16573, N13131);
xor XOR2 (N16583, N16539, N9134);
not NOT1 (N16584, N16549);
nand NAND4 (N16585, N16584, N15153, N9703, N10280);
nand NAND4 (N16586, N16583, N14034, N9852, N14263);
nand NAND2 (N16587, N16580, N15179);
buf BUF1 (N16588, N16578);
or OR3 (N16589, N16588, N1217, N8813);
buf BUF1 (N16590, N16581);
and AND4 (N16591, N16589, N16129, N747, N14051);
and AND2 (N16592, N16574, N6019);
or OR2 (N16593, N16592, N6060);
xor XOR2 (N16594, N16590, N3243);
and AND3 (N16595, N16586, N6524, N4307);
nand NAND4 (N16596, N16585, N10297, N6969, N2946);
not NOT1 (N16597, N16587);
buf BUF1 (N16598, N16572);
buf BUF1 (N16599, N16577);
and AND4 (N16600, N16576, N7999, N8400, N9180);
nor NOR3 (N16601, N16594, N4198, N1057);
buf BUF1 (N16602, N16596);
nand NAND2 (N16603, N16601, N9738);
and AND2 (N16604, N16598, N3549);
not NOT1 (N16605, N16593);
nand NAND4 (N16606, N16599, N9731, N15615, N6007);
or OR4 (N16607, N16597, N3469, N10578, N15054);
xor XOR2 (N16608, N16605, N16304);
not NOT1 (N16609, N16604);
or OR3 (N16610, N16602, N1557, N5130);
and AND3 (N16611, N16582, N13097, N5194);
and AND2 (N16612, N16609, N8197);
and AND3 (N16613, N16591, N15524, N11514);
nor NOR2 (N16614, N16603, N14387);
nand NAND3 (N16615, N16595, N3907, N2421);
nand NAND3 (N16616, N16615, N12363, N3313);
xor XOR2 (N16617, N16614, N12942);
or OR3 (N16618, N16612, N6588, N16294);
not NOT1 (N16619, N16607);
xor XOR2 (N16620, N16618, N4406);
nor NOR4 (N16621, N16600, N13562, N15702, N13611);
buf BUF1 (N16622, N16616);
or OR4 (N16623, N16606, N5435, N3364, N15564);
not NOT1 (N16624, N16619);
or OR4 (N16625, N16617, N1461, N2587, N10183);
nand NAND4 (N16626, N16610, N10405, N7100, N13325);
xor XOR2 (N16627, N16622, N15125);
xor XOR2 (N16628, N16621, N15967);
buf BUF1 (N16629, N16608);
and AND3 (N16630, N16625, N9021, N1947);
buf BUF1 (N16631, N16623);
or OR2 (N16632, N16620, N4367);
nand NAND2 (N16633, N16628, N4873);
nand NAND3 (N16634, N16632, N9994, N11444);
not NOT1 (N16635, N16634);
buf BUF1 (N16636, N16626);
or OR2 (N16637, N16635, N188);
and AND2 (N16638, N16636, N16197);
buf BUF1 (N16639, N16611);
xor XOR2 (N16640, N16639, N5116);
and AND2 (N16641, N16630, N547);
nand NAND3 (N16642, N16631, N15033, N178);
or OR4 (N16643, N16613, N3035, N15385, N15101);
nand NAND4 (N16644, N16629, N8682, N5596, N2559);
xor XOR2 (N16645, N16638, N1978);
nand NAND3 (N16646, N16627, N7860, N5225);
not NOT1 (N16647, N16646);
or OR4 (N16648, N16641, N13768, N14858, N3911);
and AND4 (N16649, N16647, N11071, N13091, N1823);
not NOT1 (N16650, N16644);
or OR4 (N16651, N16637, N13154, N5717, N7916);
or OR3 (N16652, N16648, N2009, N12043);
nand NAND3 (N16653, N16649, N13316, N6115);
or OR4 (N16654, N16652, N2767, N11640, N12372);
and AND2 (N16655, N16642, N6069);
not NOT1 (N16656, N16654);
buf BUF1 (N16657, N16633);
buf BUF1 (N16658, N16645);
not NOT1 (N16659, N16656);
buf BUF1 (N16660, N16659);
not NOT1 (N16661, N16657);
nand NAND3 (N16662, N16640, N1686, N1114);
and AND2 (N16663, N16653, N11251);
xor XOR2 (N16664, N16661, N4927);
or OR4 (N16665, N16660, N8772, N3998, N2199);
not NOT1 (N16666, N16658);
or OR2 (N16667, N16650, N15012);
or OR4 (N16668, N16665, N14930, N9797, N4572);
xor XOR2 (N16669, N16668, N9141);
or OR2 (N16670, N16663, N14637);
or OR4 (N16671, N16669, N8711, N14452, N489);
or OR4 (N16672, N16651, N4802, N3339, N9836);
not NOT1 (N16673, N16672);
buf BUF1 (N16674, N16643);
buf BUF1 (N16675, N16674);
nor NOR2 (N16676, N16666, N7847);
nor NOR4 (N16677, N16662, N540, N3022, N8275);
buf BUF1 (N16678, N16624);
buf BUF1 (N16679, N16673);
xor XOR2 (N16680, N16675, N6503);
nand NAND2 (N16681, N16671, N998);
xor XOR2 (N16682, N16667, N9822);
or OR4 (N16683, N16664, N12730, N12980, N1324);
nand NAND3 (N16684, N16683, N14219, N14605);
nor NOR3 (N16685, N16670, N13123, N10849);
buf BUF1 (N16686, N16681);
buf BUF1 (N16687, N16680);
not NOT1 (N16688, N16682);
or OR2 (N16689, N16686, N4054);
and AND2 (N16690, N16685, N16520);
nand NAND4 (N16691, N16690, N16215, N14080, N10692);
xor XOR2 (N16692, N16679, N11336);
buf BUF1 (N16693, N16678);
or OR2 (N16694, N16687, N14510);
not NOT1 (N16695, N16694);
nand NAND3 (N16696, N16692, N14416, N7665);
and AND2 (N16697, N16688, N7211);
and AND3 (N16698, N16689, N14479, N4261);
buf BUF1 (N16699, N16677);
nand NAND3 (N16700, N16691, N2592, N55);
xor XOR2 (N16701, N16655, N5011);
not NOT1 (N16702, N16693);
buf BUF1 (N16703, N16700);
and AND2 (N16704, N16684, N11257);
or OR3 (N16705, N16699, N8397, N11959);
and AND3 (N16706, N16697, N8610, N5915);
and AND2 (N16707, N16705, N13635);
buf BUF1 (N16708, N16702);
not NOT1 (N16709, N16698);
and AND4 (N16710, N16707, N11450, N6642, N7464);
or OR3 (N16711, N16706, N8040, N7130);
and AND2 (N16712, N16676, N16692);
nor NOR4 (N16713, N16711, N202, N4667, N11198);
nor NOR2 (N16714, N16703, N1918);
not NOT1 (N16715, N16708);
and AND4 (N16716, N16715, N3649, N3063, N12339);
not NOT1 (N16717, N16716);
nand NAND3 (N16718, N16717, N5594, N4002);
buf BUF1 (N16719, N16696);
nand NAND4 (N16720, N16713, N14012, N9081, N4769);
nor NOR2 (N16721, N16709, N3888);
buf BUF1 (N16722, N16710);
nand NAND3 (N16723, N16695, N10688, N9257);
not NOT1 (N16724, N16723);
or OR3 (N16725, N16721, N1942, N2045);
not NOT1 (N16726, N16719);
nand NAND3 (N16727, N16720, N12236, N3522);
nor NOR2 (N16728, N16718, N4420);
not NOT1 (N16729, N16726);
not NOT1 (N16730, N16729);
not NOT1 (N16731, N16724);
nor NOR3 (N16732, N16728, N15669, N4547);
xor XOR2 (N16733, N16714, N13203);
buf BUF1 (N16734, N16733);
nor NOR2 (N16735, N16722, N9691);
nor NOR3 (N16736, N16725, N13174, N5578);
and AND2 (N16737, N16732, N5937);
nand NAND3 (N16738, N16736, N8160, N9854);
nor NOR2 (N16739, N16730, N14437);
buf BUF1 (N16740, N16734);
nand NAND4 (N16741, N16735, N10329, N12747, N16149);
xor XOR2 (N16742, N16740, N2556);
nor NOR3 (N16743, N16738, N4930, N134);
xor XOR2 (N16744, N16742, N15067);
nor NOR3 (N16745, N16739, N5612, N14019);
buf BUF1 (N16746, N16727);
xor XOR2 (N16747, N16704, N3561);
not NOT1 (N16748, N16747);
nand NAND4 (N16749, N16712, N10516, N7211, N12824);
and AND4 (N16750, N16743, N3220, N14885, N7257);
nand NAND3 (N16751, N16701, N8841, N16435);
not NOT1 (N16752, N16737);
or OR4 (N16753, N16752, N12077, N13124, N11618);
buf BUF1 (N16754, N16745);
or OR3 (N16755, N16746, N15010, N10272);
nand NAND2 (N16756, N16741, N9786);
or OR3 (N16757, N16750, N8754, N2198);
not NOT1 (N16758, N16748);
and AND3 (N16759, N16754, N134, N10432);
and AND3 (N16760, N16751, N3564, N5628);
xor XOR2 (N16761, N16753, N14655);
nor NOR4 (N16762, N16761, N4672, N1280, N4614);
buf BUF1 (N16763, N16757);
or OR2 (N16764, N16731, N12371);
xor XOR2 (N16765, N16762, N12650);
and AND3 (N16766, N16755, N8806, N5276);
xor XOR2 (N16767, N16758, N12742);
buf BUF1 (N16768, N16766);
and AND2 (N16769, N16760, N5836);
nand NAND3 (N16770, N16756, N7520, N7898);
not NOT1 (N16771, N16763);
or OR2 (N16772, N16744, N11299);
or OR3 (N16773, N16767, N4577, N7217);
buf BUF1 (N16774, N16749);
nor NOR2 (N16775, N16769, N16162);
buf BUF1 (N16776, N16774);
buf BUF1 (N16777, N16772);
not NOT1 (N16778, N16773);
and AND3 (N16779, N16770, N13328, N12580);
xor XOR2 (N16780, N16779, N3090);
xor XOR2 (N16781, N16765, N4610);
and AND2 (N16782, N16780, N160);
nand NAND4 (N16783, N16781, N8676, N11670, N8117);
nand NAND3 (N16784, N16776, N9955, N14961);
nand NAND2 (N16785, N16783, N10103);
and AND4 (N16786, N16759, N9743, N13179, N9351);
not NOT1 (N16787, N16784);
not NOT1 (N16788, N16764);
and AND3 (N16789, N16777, N13718, N16193);
or OR2 (N16790, N16775, N2527);
nor NOR3 (N16791, N16768, N7392, N10667);
not NOT1 (N16792, N16786);
buf BUF1 (N16793, N16787);
not NOT1 (N16794, N16790);
or OR2 (N16795, N16771, N12229);
nor NOR4 (N16796, N16782, N5940, N7164, N6891);
buf BUF1 (N16797, N16794);
nor NOR3 (N16798, N16797, N13303, N14439);
and AND4 (N16799, N16796, N3459, N16742, N11997);
or OR2 (N16800, N16788, N15481);
buf BUF1 (N16801, N16778);
or OR4 (N16802, N16798, N618, N8696, N7590);
nand NAND3 (N16803, N16793, N14864, N14613);
xor XOR2 (N16804, N16791, N9531);
nand NAND2 (N16805, N16800, N2250);
and AND4 (N16806, N16803, N678, N10016, N484);
and AND3 (N16807, N16799, N6411, N76);
nand NAND4 (N16808, N16789, N9720, N8083, N10705);
nand NAND4 (N16809, N16792, N1351, N7425, N9361);
nor NOR3 (N16810, N16785, N9532, N14934);
nand NAND4 (N16811, N16808, N11808, N4014, N1208);
nand NAND3 (N16812, N16795, N16374, N7158);
or OR4 (N16813, N16801, N3827, N14764, N16617);
not NOT1 (N16814, N16805);
and AND3 (N16815, N16804, N7989, N4372);
buf BUF1 (N16816, N16809);
nor NOR2 (N16817, N16806, N3390);
and AND4 (N16818, N16807, N4825, N13944, N14158);
buf BUF1 (N16819, N16813);
xor XOR2 (N16820, N16812, N4682);
buf BUF1 (N16821, N16811);
and AND3 (N16822, N16810, N6979, N9263);
and AND3 (N16823, N16820, N6685, N2661);
buf BUF1 (N16824, N16816);
nor NOR4 (N16825, N16815, N11601, N6115, N8131);
or OR3 (N16826, N16817, N4582, N15685);
nor NOR4 (N16827, N16826, N6825, N1853, N3703);
buf BUF1 (N16828, N16823);
nor NOR3 (N16829, N16814, N14919, N4601);
nand NAND3 (N16830, N16822, N12885, N3042);
not NOT1 (N16831, N16825);
nor NOR2 (N16832, N16830, N2544);
and AND4 (N16833, N16824, N1346, N2468, N3047);
nor NOR4 (N16834, N16829, N6054, N11889, N8407);
not NOT1 (N16835, N16821);
not NOT1 (N16836, N16832);
and AND3 (N16837, N16835, N9026, N8671);
buf BUF1 (N16838, N16827);
and AND4 (N16839, N16836, N4785, N7214, N14680);
not NOT1 (N16840, N16834);
and AND4 (N16841, N16839, N13235, N4937, N14059);
buf BUF1 (N16842, N16828);
buf BUF1 (N16843, N16841);
nand NAND3 (N16844, N16802, N5544, N10882);
xor XOR2 (N16845, N16838, N12839);
or OR3 (N16846, N16845, N5582, N7453);
not NOT1 (N16847, N16837);
nor NOR3 (N16848, N16847, N8075, N2392);
nor NOR2 (N16849, N16848, N14052);
xor XOR2 (N16850, N16819, N10189);
nor NOR2 (N16851, N16843, N1422);
xor XOR2 (N16852, N16844, N14021);
buf BUF1 (N16853, N16842);
buf BUF1 (N16854, N16818);
xor XOR2 (N16855, N16852, N6578);
and AND4 (N16856, N16854, N15615, N9016, N16548);
nor NOR2 (N16857, N16850, N15217);
or OR3 (N16858, N16855, N8365, N2082);
buf BUF1 (N16859, N16851);
not NOT1 (N16860, N16858);
nor NOR2 (N16861, N16853, N3346);
or OR3 (N16862, N16860, N14148, N6105);
buf BUF1 (N16863, N16840);
xor XOR2 (N16864, N16846, N10678);
xor XOR2 (N16865, N16857, N9036);
nor NOR4 (N16866, N16863, N8314, N2703, N13345);
buf BUF1 (N16867, N16861);
xor XOR2 (N16868, N16867, N15913);
or OR2 (N16869, N16862, N11528);
or OR3 (N16870, N16859, N5139, N10434);
nand NAND4 (N16871, N16865, N11975, N12009, N3102);
nand NAND2 (N16872, N16833, N1493);
and AND4 (N16873, N16869, N11047, N5484, N2271);
or OR2 (N16874, N16864, N5269);
nand NAND3 (N16875, N16871, N6225, N10632);
xor XOR2 (N16876, N16868, N15799);
not NOT1 (N16877, N16874);
not NOT1 (N16878, N16873);
not NOT1 (N16879, N16872);
and AND4 (N16880, N16878, N14742, N10738, N13553);
and AND2 (N16881, N16870, N865);
or OR2 (N16882, N16879, N7272);
nor NOR4 (N16883, N16881, N9486, N1490, N1363);
and AND2 (N16884, N16849, N16421);
and AND4 (N16885, N16856, N13843, N4021, N7607);
xor XOR2 (N16886, N16875, N2557);
xor XOR2 (N16887, N16882, N229);
nor NOR2 (N16888, N16884, N14860);
nor NOR3 (N16889, N16866, N14637, N6451);
not NOT1 (N16890, N16880);
or OR4 (N16891, N16890, N777, N3723, N586);
and AND2 (N16892, N16891, N10275);
nor NOR4 (N16893, N16886, N6983, N5460, N5137);
not NOT1 (N16894, N16883);
and AND4 (N16895, N16889, N2241, N1921, N6226);
or OR3 (N16896, N16895, N2872, N16699);
nand NAND4 (N16897, N16896, N15571, N1699, N10131);
and AND4 (N16898, N16897, N789, N1502, N11786);
xor XOR2 (N16899, N16831, N1409);
nor NOR4 (N16900, N16893, N2884, N9183, N5246);
and AND2 (N16901, N16900, N16873);
not NOT1 (N16902, N16887);
and AND2 (N16903, N16892, N2283);
not NOT1 (N16904, N16885);
and AND3 (N16905, N16888, N12048, N9272);
nor NOR2 (N16906, N16902, N10913);
not NOT1 (N16907, N16903);
or OR3 (N16908, N16899, N9975, N3382);
xor XOR2 (N16909, N16901, N3147);
not NOT1 (N16910, N16898);
or OR2 (N16911, N16894, N9318);
and AND4 (N16912, N16911, N15984, N7131, N6456);
or OR4 (N16913, N16907, N13104, N1858, N12235);
xor XOR2 (N16914, N16904, N2736);
nand NAND3 (N16915, N16876, N5934, N2807);
and AND3 (N16916, N16912, N10893, N11408);
and AND3 (N16917, N16913, N34, N13100);
and AND4 (N16918, N16910, N16534, N7585, N11409);
or OR3 (N16919, N16918, N10578, N4891);
and AND3 (N16920, N16908, N1232, N15646);
xor XOR2 (N16921, N16905, N2821);
xor XOR2 (N16922, N16919, N12280);
and AND4 (N16923, N16915, N11255, N9116, N2724);
nand NAND4 (N16924, N16906, N14228, N7304, N6227);
buf BUF1 (N16925, N16923);
buf BUF1 (N16926, N16916);
nand NAND4 (N16927, N16924, N12719, N1672, N12378);
nor NOR4 (N16928, N16917, N14907, N6882, N16112);
nand NAND4 (N16929, N16920, N886, N15397, N12198);
not NOT1 (N16930, N16929);
xor XOR2 (N16931, N16921, N5709);
xor XOR2 (N16932, N16877, N373);
nand NAND4 (N16933, N16932, N4985, N64, N1756);
not NOT1 (N16934, N16930);
not NOT1 (N16935, N16931);
and AND4 (N16936, N16925, N12481, N9490, N1292);
and AND3 (N16937, N16935, N15686, N14163);
not NOT1 (N16938, N16914);
buf BUF1 (N16939, N16933);
nor NOR4 (N16940, N16939, N9905, N16037, N12213);
xor XOR2 (N16941, N16937, N16065);
or OR4 (N16942, N16940, N6691, N1104, N7495);
and AND3 (N16943, N16941, N15190, N10428);
xor XOR2 (N16944, N16936, N9124);
and AND4 (N16945, N16926, N11714, N14953, N16202);
or OR3 (N16946, N16943, N11104, N16704);
not NOT1 (N16947, N16946);
xor XOR2 (N16948, N16942, N3240);
nor NOR3 (N16949, N16928, N13504, N11762);
nor NOR4 (N16950, N16922, N2227, N13298, N4724);
nand NAND4 (N16951, N16945, N9456, N12385, N7403);
and AND3 (N16952, N16927, N10702, N16939);
or OR3 (N16953, N16949, N5399, N13271);
nand NAND2 (N16954, N16951, N1896);
buf BUF1 (N16955, N16944);
buf BUF1 (N16956, N16947);
nand NAND2 (N16957, N16948, N7111);
nand NAND4 (N16958, N16955, N365, N7677, N12227);
buf BUF1 (N16959, N16953);
not NOT1 (N16960, N16950);
buf BUF1 (N16961, N16954);
nand NAND4 (N16962, N16958, N12597, N11046, N9138);
buf BUF1 (N16963, N16960);
buf BUF1 (N16964, N16959);
nand NAND4 (N16965, N16962, N16225, N4149, N13745);
nand NAND3 (N16966, N16964, N11213, N4480);
xor XOR2 (N16967, N16956, N15341);
nand NAND3 (N16968, N16957, N2821, N16758);
not NOT1 (N16969, N16934);
or OR2 (N16970, N16966, N6278);
and AND4 (N16971, N16969, N12685, N2681, N2158);
or OR2 (N16972, N16938, N16006);
nor NOR4 (N16973, N16970, N8786, N12512, N14770);
not NOT1 (N16974, N16961);
buf BUF1 (N16975, N16968);
not NOT1 (N16976, N16973);
xor XOR2 (N16977, N16963, N13585);
buf BUF1 (N16978, N16971);
or OR3 (N16979, N16972, N5505, N591);
or OR4 (N16980, N16975, N12143, N11589, N1541);
not NOT1 (N16981, N16977);
nor NOR4 (N16982, N16980, N14215, N8050, N4515);
not NOT1 (N16983, N16979);
not NOT1 (N16984, N16981);
buf BUF1 (N16985, N16978);
or OR4 (N16986, N16982, N12135, N13877, N16185);
nor NOR3 (N16987, N16965, N15855, N3552);
not NOT1 (N16988, N16983);
xor XOR2 (N16989, N16986, N2325);
nor NOR3 (N16990, N16984, N12610, N6615);
nand NAND2 (N16991, N16967, N8228);
nand NAND2 (N16992, N16987, N7616);
not NOT1 (N16993, N16985);
or OR3 (N16994, N16988, N15377, N1722);
nor NOR4 (N16995, N16991, N655, N13534, N3029);
or OR3 (N16996, N16976, N13598, N16312);
nor NOR3 (N16997, N16996, N3520, N13834);
nand NAND3 (N16998, N16992, N3757, N7372);
nand NAND3 (N16999, N16993, N15014, N11963);
or OR2 (N17000, N16974, N14837);
buf BUF1 (N17001, N16909);
and AND2 (N17002, N16952, N16637);
nand NAND4 (N17003, N16997, N13750, N1926, N5429);
buf BUF1 (N17004, N16989);
and AND4 (N17005, N16990, N15172, N2785, N13861);
nor NOR2 (N17006, N17000, N15865);
nor NOR4 (N17007, N17002, N3304, N8143, N1867);
and AND4 (N17008, N16999, N3662, N6272, N9031);
nand NAND2 (N17009, N17004, N13769);
and AND3 (N17010, N17009, N9185, N10086);
xor XOR2 (N17011, N17007, N14496);
and AND4 (N17012, N17006, N12202, N5480, N2773);
not NOT1 (N17013, N17012);
or OR3 (N17014, N16995, N2758, N5966);
and AND4 (N17015, N17011, N2495, N8722, N14216);
buf BUF1 (N17016, N16994);
nand NAND3 (N17017, N17003, N9637, N12337);
nand NAND4 (N17018, N17014, N9479, N14707, N9206);
nor NOR2 (N17019, N17018, N14122);
or OR3 (N17020, N16998, N8918, N12527);
buf BUF1 (N17021, N17001);
or OR3 (N17022, N17008, N15748, N1328);
nor NOR2 (N17023, N17021, N7698);
and AND3 (N17024, N17022, N5610, N1653);
xor XOR2 (N17025, N17015, N9095);
buf BUF1 (N17026, N17013);
buf BUF1 (N17027, N17020);
buf BUF1 (N17028, N17010);
not NOT1 (N17029, N17028);
and AND4 (N17030, N17019, N3184, N6718, N11657);
nor NOR3 (N17031, N17025, N15417, N9795);
nor NOR3 (N17032, N17016, N11209, N589);
not NOT1 (N17033, N17024);
nor NOR4 (N17034, N17026, N10257, N14317, N10597);
not NOT1 (N17035, N17033);
nand NAND2 (N17036, N17031, N2220);
xor XOR2 (N17037, N17027, N6668);
not NOT1 (N17038, N17037);
xor XOR2 (N17039, N17005, N7590);
nand NAND3 (N17040, N17038, N16339, N9002);
buf BUF1 (N17041, N17040);
nor NOR4 (N17042, N17034, N4433, N5316, N921);
not NOT1 (N17043, N17036);
nand NAND3 (N17044, N17042, N79, N6199);
nand NAND2 (N17045, N17017, N9010);
nand NAND4 (N17046, N17045, N12939, N7779, N1559);
buf BUF1 (N17047, N17030);
nand NAND3 (N17048, N17041, N2967, N2359);
nor NOR4 (N17049, N17047, N12921, N6683, N6954);
nor NOR3 (N17050, N17048, N6413, N6263);
and AND2 (N17051, N17050, N16604);
nand NAND3 (N17052, N17044, N12348, N7657);
buf BUF1 (N17053, N17029);
or OR2 (N17054, N17052, N13885);
xor XOR2 (N17055, N17039, N4128);
not NOT1 (N17056, N17055);
nand NAND4 (N17057, N17043, N11171, N15786, N2271);
nand NAND3 (N17058, N17049, N3754, N6980);
nand NAND4 (N17059, N17053, N9140, N3418, N4368);
not NOT1 (N17060, N17035);
nor NOR2 (N17061, N17051, N9194);
xor XOR2 (N17062, N17058, N16902);
and AND4 (N17063, N17057, N8007, N7775, N912);
nor NOR2 (N17064, N17061, N10925);
or OR3 (N17065, N17063, N14307, N2809);
nor NOR3 (N17066, N17060, N924, N3363);
or OR4 (N17067, N17064, N2099, N9524, N15134);
not NOT1 (N17068, N17046);
or OR3 (N17069, N17032, N463, N10192);
buf BUF1 (N17070, N17056);
nor NOR2 (N17071, N17023, N16983);
nor NOR2 (N17072, N17070, N10394);
nand NAND2 (N17073, N17071, N10295);
not NOT1 (N17074, N17069);
and AND3 (N17075, N17068, N2760, N713);
or OR3 (N17076, N17075, N8738, N3740);
xor XOR2 (N17077, N17076, N14172);
xor XOR2 (N17078, N17077, N524);
and AND4 (N17079, N17074, N13429, N13770, N14292);
not NOT1 (N17080, N17054);
xor XOR2 (N17081, N17073, N5424);
nand NAND2 (N17082, N17059, N6761);
not NOT1 (N17083, N17079);
nand NAND3 (N17084, N17072, N8723, N1242);
buf BUF1 (N17085, N17084);
and AND3 (N17086, N17083, N3813, N3764);
or OR4 (N17087, N17082, N4172, N5807, N4801);
xor XOR2 (N17088, N17080, N15027);
xor XOR2 (N17089, N17085, N9273);
nand NAND4 (N17090, N17087, N6866, N2055, N1747);
and AND3 (N17091, N17081, N7653, N14121);
and AND3 (N17092, N17066, N12553, N5350);
buf BUF1 (N17093, N17078);
or OR3 (N17094, N17090, N10527, N973);
nor NOR3 (N17095, N17086, N7752, N6140);
buf BUF1 (N17096, N17095);
buf BUF1 (N17097, N17094);
or OR2 (N17098, N17093, N3813);
buf BUF1 (N17099, N17098);
xor XOR2 (N17100, N17097, N8945);
nand NAND3 (N17101, N17065, N12748, N3038);
xor XOR2 (N17102, N17089, N164);
not NOT1 (N17103, N17092);
and AND4 (N17104, N17088, N15820, N14849, N2628);
nor NOR2 (N17105, N17091, N13983);
nand NAND3 (N17106, N17104, N11019, N10959);
buf BUF1 (N17107, N17099);
buf BUF1 (N17108, N17103);
xor XOR2 (N17109, N17102, N13679);
xor XOR2 (N17110, N17062, N258);
nor NOR2 (N17111, N17100, N14972);
and AND2 (N17112, N17106, N3542);
xor XOR2 (N17113, N17110, N9465);
xor XOR2 (N17114, N17109, N7335);
xor XOR2 (N17115, N17096, N2744);
nand NAND3 (N17116, N17111, N8419, N16566);
or OR2 (N17117, N17108, N12639);
nor NOR2 (N17118, N17107, N12811);
and AND2 (N17119, N17115, N9590);
not NOT1 (N17120, N17113);
nor NOR3 (N17121, N17116, N521, N2341);
buf BUF1 (N17122, N17117);
and AND4 (N17123, N17105, N1714, N1086, N8075);
nor NOR3 (N17124, N17122, N13964, N6241);
xor XOR2 (N17125, N17121, N12818);
nand NAND4 (N17126, N17118, N7191, N1841, N15884);
xor XOR2 (N17127, N17119, N14982);
nor NOR3 (N17128, N17123, N7876, N12115);
nor NOR2 (N17129, N17128, N13471);
or OR4 (N17130, N17114, N6596, N10533, N8122);
and AND4 (N17131, N17067, N8850, N14329, N4474);
and AND4 (N17132, N17124, N8404, N9407, N13764);
nand NAND3 (N17133, N17112, N17002, N15169);
xor XOR2 (N17134, N17130, N1669);
xor XOR2 (N17135, N17134, N11037);
xor XOR2 (N17136, N17129, N32);
nand NAND4 (N17137, N17133, N13141, N14426, N11194);
nor NOR2 (N17138, N17132, N2840);
nand NAND2 (N17139, N17127, N10854);
not NOT1 (N17140, N17101);
xor XOR2 (N17141, N17139, N3817);
xor XOR2 (N17142, N17131, N5185);
buf BUF1 (N17143, N17141);
and AND4 (N17144, N17142, N4432, N17061, N15499);
or OR3 (N17145, N17126, N9170, N15023);
buf BUF1 (N17146, N17143);
not NOT1 (N17147, N17140);
nor NOR2 (N17148, N17138, N10814);
not NOT1 (N17149, N17147);
buf BUF1 (N17150, N17148);
not NOT1 (N17151, N17150);
and AND2 (N17152, N17136, N13104);
and AND2 (N17153, N17135, N11018);
not NOT1 (N17154, N17137);
not NOT1 (N17155, N17125);
nand NAND4 (N17156, N17151, N8094, N1111, N19);
xor XOR2 (N17157, N17146, N9432);
not NOT1 (N17158, N17155);
nand NAND3 (N17159, N17158, N1754, N8041);
buf BUF1 (N17160, N17159);
or OR4 (N17161, N17160, N10509, N8715, N5346);
xor XOR2 (N17162, N17156, N11020);
nor NOR2 (N17163, N17145, N3406);
xor XOR2 (N17164, N17153, N11159);
or OR3 (N17165, N17163, N4526, N11190);
nand NAND2 (N17166, N17157, N5059);
and AND2 (N17167, N17144, N1414);
buf BUF1 (N17168, N17167);
not NOT1 (N17169, N17161);
nor NOR2 (N17170, N17165, N14712);
and AND2 (N17171, N17120, N13758);
xor XOR2 (N17172, N17171, N7621);
not NOT1 (N17173, N17152);
buf BUF1 (N17174, N17168);
buf BUF1 (N17175, N17169);
or OR3 (N17176, N17149, N16043, N144);
and AND2 (N17177, N17154, N4445);
and AND3 (N17178, N17177, N2920, N13019);
buf BUF1 (N17179, N17170);
nor NOR4 (N17180, N17176, N7520, N2484, N3464);
or OR3 (N17181, N17175, N5870, N7173);
buf BUF1 (N17182, N17172);
nand NAND2 (N17183, N17174, N14479);
nor NOR4 (N17184, N17182, N6850, N6868, N807);
xor XOR2 (N17185, N17166, N16449);
or OR2 (N17186, N17164, N6606);
buf BUF1 (N17187, N17186);
buf BUF1 (N17188, N17173);
buf BUF1 (N17189, N17183);
nand NAND3 (N17190, N17180, N13432, N15256);
not NOT1 (N17191, N17181);
xor XOR2 (N17192, N17188, N10661);
xor XOR2 (N17193, N17179, N3122);
xor XOR2 (N17194, N17192, N7557);
or OR4 (N17195, N17193, N17177, N15884, N2320);
not NOT1 (N17196, N17191);
buf BUF1 (N17197, N17185);
buf BUF1 (N17198, N17184);
buf BUF1 (N17199, N17198);
not NOT1 (N17200, N17178);
nand NAND4 (N17201, N17200, N5983, N5897, N2644);
nor NOR2 (N17202, N17190, N4597);
or OR4 (N17203, N17189, N13958, N295, N6839);
and AND2 (N17204, N17187, N2517);
xor XOR2 (N17205, N17202, N14367);
nand NAND2 (N17206, N17201, N8944);
nor NOR4 (N17207, N17194, N14838, N2098, N3505);
not NOT1 (N17208, N17197);
buf BUF1 (N17209, N17206);
and AND2 (N17210, N17208, N4314);
xor XOR2 (N17211, N17196, N3945);
nand NAND4 (N17212, N17195, N11196, N312, N3961);
nor NOR4 (N17213, N17209, N15864, N1338, N3593);
buf BUF1 (N17214, N17212);
not NOT1 (N17215, N17203);
not NOT1 (N17216, N17211);
buf BUF1 (N17217, N17205);
or OR2 (N17218, N17204, N1153);
xor XOR2 (N17219, N17199, N4582);
xor XOR2 (N17220, N17162, N15019);
and AND2 (N17221, N17216, N6139);
nor NOR3 (N17222, N17219, N7288, N15842);
xor XOR2 (N17223, N17213, N4407);
or OR4 (N17224, N17223, N10024, N11644, N7551);
nor NOR4 (N17225, N17222, N3092, N4923, N1140);
and AND2 (N17226, N17210, N10496);
nand NAND3 (N17227, N17225, N4988, N6993);
nor NOR4 (N17228, N17221, N11915, N5678, N6201);
and AND2 (N17229, N17215, N15503);
or OR2 (N17230, N17226, N15917);
nor NOR2 (N17231, N17229, N10712);
xor XOR2 (N17232, N17228, N10731);
buf BUF1 (N17233, N17207);
xor XOR2 (N17234, N17220, N8132);
nand NAND4 (N17235, N17214, N15460, N7372, N5564);
buf BUF1 (N17236, N17230);
not NOT1 (N17237, N17217);
nor NOR4 (N17238, N17227, N11968, N4122, N6837);
buf BUF1 (N17239, N17234);
and AND2 (N17240, N17231, N10367);
buf BUF1 (N17241, N17239);
not NOT1 (N17242, N17236);
not NOT1 (N17243, N17238);
buf BUF1 (N17244, N17242);
or OR3 (N17245, N17224, N11734, N1313);
xor XOR2 (N17246, N17245, N4018);
nand NAND2 (N17247, N17241, N12916);
xor XOR2 (N17248, N17218, N6277);
buf BUF1 (N17249, N17243);
buf BUF1 (N17250, N17237);
or OR3 (N17251, N17235, N7635, N602);
buf BUF1 (N17252, N17251);
nand NAND2 (N17253, N17247, N3219);
buf BUF1 (N17254, N17250);
xor XOR2 (N17255, N17240, N1715);
nor NOR2 (N17256, N17253, N6151);
buf BUF1 (N17257, N17244);
buf BUF1 (N17258, N17254);
nor NOR2 (N17259, N17246, N14855);
and AND2 (N17260, N17233, N15358);
nor NOR3 (N17261, N17252, N7063, N10525);
or OR4 (N17262, N17259, N11763, N6734, N13194);
nor NOR4 (N17263, N17257, N8345, N6030, N297);
buf BUF1 (N17264, N17260);
nand NAND4 (N17265, N17255, N11214, N7851, N6958);
nand NAND4 (N17266, N17263, N16248, N13433, N13928);
xor XOR2 (N17267, N17266, N12788);
nand NAND3 (N17268, N17264, N6446, N13276);
nor NOR4 (N17269, N17261, N16648, N7272, N9119);
and AND2 (N17270, N17232, N15997);
buf BUF1 (N17271, N17249);
and AND2 (N17272, N17258, N3879);
nand NAND2 (N17273, N17267, N11750);
and AND3 (N17274, N17269, N361, N13338);
nand NAND4 (N17275, N17271, N7942, N9331, N1161);
not NOT1 (N17276, N17268);
buf BUF1 (N17277, N17272);
or OR4 (N17278, N17274, N2697, N6092, N15895);
not NOT1 (N17279, N17276);
not NOT1 (N17280, N17270);
and AND3 (N17281, N17279, N9675, N843);
nor NOR4 (N17282, N17265, N2098, N843, N2491);
and AND4 (N17283, N17262, N9507, N10264, N4199);
nand NAND4 (N17284, N17283, N12899, N11502, N10487);
buf BUF1 (N17285, N17273);
xor XOR2 (N17286, N17278, N1139);
xor XOR2 (N17287, N17256, N6901);
nor NOR4 (N17288, N17284, N6018, N7519, N15693);
nor NOR4 (N17289, N17286, N11473, N5753, N9012);
and AND2 (N17290, N17277, N7619);
buf BUF1 (N17291, N17248);
xor XOR2 (N17292, N17287, N17073);
xor XOR2 (N17293, N17282, N5174);
nor NOR3 (N17294, N17293, N15204, N1754);
or OR3 (N17295, N17288, N10722, N1377);
or OR2 (N17296, N17291, N12937);
or OR2 (N17297, N17290, N8184);
nand NAND2 (N17298, N17292, N5013);
or OR2 (N17299, N17289, N7502);
nand NAND3 (N17300, N17294, N2115, N16844);
xor XOR2 (N17301, N17300, N1962);
buf BUF1 (N17302, N17301);
not NOT1 (N17303, N17280);
nor NOR2 (N17304, N17302, N14706);
or OR4 (N17305, N17281, N461, N13906, N850);
not NOT1 (N17306, N17298);
not NOT1 (N17307, N17305);
and AND4 (N17308, N17297, N12658, N10860, N10219);
buf BUF1 (N17309, N17308);
buf BUF1 (N17310, N17309);
and AND4 (N17311, N17310, N699, N2037, N4128);
nor NOR2 (N17312, N17299, N12493);
or OR4 (N17313, N17312, N3853, N8298, N14722);
buf BUF1 (N17314, N17304);
buf BUF1 (N17315, N17314);
not NOT1 (N17316, N17313);
buf BUF1 (N17317, N17311);
and AND2 (N17318, N17315, N14621);
buf BUF1 (N17319, N17296);
nor NOR4 (N17320, N17275, N2976, N9316, N12990);
nand NAND4 (N17321, N17319, N3699, N8705, N647);
xor XOR2 (N17322, N17303, N15074);
or OR3 (N17323, N17316, N16962, N2855);
or OR4 (N17324, N17317, N633, N9085, N14441);
buf BUF1 (N17325, N17318);
xor XOR2 (N17326, N17322, N16488);
or OR4 (N17327, N17324, N9666, N15665, N5291);
or OR2 (N17328, N17320, N12986);
nand NAND3 (N17329, N17323, N12049, N8840);
nor NOR3 (N17330, N17325, N4544, N2124);
not NOT1 (N17331, N17321);
and AND4 (N17332, N17327, N14592, N3794, N13343);
or OR4 (N17333, N17326, N14302, N12756, N9115);
nand NAND2 (N17334, N17295, N583);
buf BUF1 (N17335, N17331);
or OR3 (N17336, N17332, N7797, N6522);
or OR2 (N17337, N17328, N1508);
xor XOR2 (N17338, N17306, N5018);
not NOT1 (N17339, N17337);
buf BUF1 (N17340, N17329);
buf BUF1 (N17341, N17330);
buf BUF1 (N17342, N17336);
and AND3 (N17343, N17338, N174, N9312);
nand NAND4 (N17344, N17341, N390, N8996, N10474);
nand NAND2 (N17345, N17334, N4118);
buf BUF1 (N17346, N17344);
nor NOR3 (N17347, N17285, N2001, N13900);
xor XOR2 (N17348, N17343, N4724);
xor XOR2 (N17349, N17346, N10205);
or OR2 (N17350, N17340, N11230);
not NOT1 (N17351, N17335);
nor NOR2 (N17352, N17307, N7196);
or OR3 (N17353, N17349, N13784, N11981);
xor XOR2 (N17354, N17353, N5925);
or OR3 (N17355, N17339, N3599, N12574);
not NOT1 (N17356, N17345);
xor XOR2 (N17357, N17347, N15320);
not NOT1 (N17358, N17348);
nor NOR4 (N17359, N17357, N10478, N3521, N9925);
buf BUF1 (N17360, N17356);
or OR4 (N17361, N17351, N6516, N6022, N522);
nand NAND3 (N17362, N17342, N15392, N2119);
not NOT1 (N17363, N17352);
xor XOR2 (N17364, N17358, N2129);
nor NOR4 (N17365, N17362, N12375, N7852, N13589);
xor XOR2 (N17366, N17360, N3666);
buf BUF1 (N17367, N17355);
not NOT1 (N17368, N17367);
nand NAND3 (N17369, N17359, N4747, N12679);
xor XOR2 (N17370, N17365, N15);
not NOT1 (N17371, N17354);
and AND2 (N17372, N17363, N14657);
not NOT1 (N17373, N17372);
nand NAND2 (N17374, N17368, N15723);
nor NOR4 (N17375, N17364, N10581, N14645, N9585);
or OR2 (N17376, N17371, N13355);
xor XOR2 (N17377, N17350, N3313);
nand NAND3 (N17378, N17369, N13645, N12951);
nor NOR4 (N17379, N17361, N11516, N1477, N8446);
nor NOR2 (N17380, N17376, N10794);
nand NAND4 (N17381, N17333, N16104, N4959, N11530);
or OR4 (N17382, N17373, N7720, N6940, N13250);
buf BUF1 (N17383, N17381);
xor XOR2 (N17384, N17380, N1823);
xor XOR2 (N17385, N17382, N15892);
or OR3 (N17386, N17375, N14792, N11145);
nand NAND4 (N17387, N17378, N16764, N1572, N8942);
not NOT1 (N17388, N17383);
and AND3 (N17389, N17384, N5771, N5685);
or OR2 (N17390, N17387, N3078);
nor NOR2 (N17391, N17370, N25);
not NOT1 (N17392, N17379);
and AND4 (N17393, N17389, N15509, N17303, N3973);
xor XOR2 (N17394, N17377, N10079);
nor NOR2 (N17395, N17393, N1246);
nand NAND4 (N17396, N17392, N10603, N6265, N13822);
not NOT1 (N17397, N17374);
buf BUF1 (N17398, N17391);
xor XOR2 (N17399, N17397, N12088);
or OR2 (N17400, N17395, N15230);
buf BUF1 (N17401, N17399);
or OR4 (N17402, N17385, N3653, N7217, N2128);
and AND4 (N17403, N17396, N11221, N6954, N8087);
buf BUF1 (N17404, N17403);
nor NOR2 (N17405, N17400, N8802);
xor XOR2 (N17406, N17386, N6729);
nor NOR2 (N17407, N17388, N12873);
not NOT1 (N17408, N17398);
nor NOR2 (N17409, N17401, N3712);
xor XOR2 (N17410, N17366, N9394);
not NOT1 (N17411, N17394);
buf BUF1 (N17412, N17390);
nand NAND4 (N17413, N17412, N14231, N17371, N6312);
buf BUF1 (N17414, N17404);
nor NOR2 (N17415, N17405, N5732);
nand NAND4 (N17416, N17415, N12540, N17242, N2182);
nor NOR2 (N17417, N17407, N6830);
or OR4 (N17418, N17410, N11537, N2895, N10557);
xor XOR2 (N17419, N17406, N9524);
or OR2 (N17420, N17408, N16197);
and AND4 (N17421, N17413, N4986, N13259, N10872);
nand NAND4 (N17422, N17411, N3827, N16870, N11520);
and AND2 (N17423, N17414, N9498);
or OR3 (N17424, N17418, N584, N1604);
and AND2 (N17425, N17420, N8776);
not NOT1 (N17426, N17424);
xor XOR2 (N17427, N17422, N13884);
nand NAND2 (N17428, N17416, N10335);
or OR3 (N17429, N17419, N4333, N794);
nand NAND3 (N17430, N17417, N15460, N16121);
and AND3 (N17431, N17402, N5243, N14589);
and AND4 (N17432, N17431, N6570, N16524, N9595);
xor XOR2 (N17433, N17409, N7396);
not NOT1 (N17434, N17433);
not NOT1 (N17435, N17429);
not NOT1 (N17436, N17432);
nand NAND2 (N17437, N17428, N11568);
xor XOR2 (N17438, N17434, N15647);
nor NOR3 (N17439, N17438, N10062, N3934);
or OR2 (N17440, N17437, N11414);
xor XOR2 (N17441, N17436, N3368);
nand NAND3 (N17442, N17440, N11122, N10257);
xor XOR2 (N17443, N17427, N10320);
nand NAND3 (N17444, N17425, N1227, N12915);
and AND2 (N17445, N17426, N16429);
xor XOR2 (N17446, N17423, N14027);
nand NAND2 (N17447, N17442, N13622);
xor XOR2 (N17448, N17446, N14691);
buf BUF1 (N17449, N17421);
or OR3 (N17450, N17447, N13815, N3931);
not NOT1 (N17451, N17445);
nor NOR2 (N17452, N17448, N7052);
and AND4 (N17453, N17443, N7385, N17065, N1560);
not NOT1 (N17454, N17451);
nor NOR2 (N17455, N17430, N13970);
nor NOR4 (N17456, N17453, N16355, N3747, N8536);
or OR2 (N17457, N17452, N13841);
not NOT1 (N17458, N17454);
buf BUF1 (N17459, N17458);
nor NOR3 (N17460, N17439, N4956, N15710);
buf BUF1 (N17461, N17444);
nand NAND3 (N17462, N17435, N5820, N14268);
nand NAND4 (N17463, N17459, N8678, N6191, N8380);
nor NOR3 (N17464, N17462, N2323, N4825);
nand NAND2 (N17465, N17460, N14914);
not NOT1 (N17466, N17456);
buf BUF1 (N17467, N17441);
and AND2 (N17468, N17461, N1171);
nand NAND2 (N17469, N17455, N4826);
and AND4 (N17470, N17457, N15210, N14400, N9485);
xor XOR2 (N17471, N17463, N5242);
nor NOR3 (N17472, N17470, N9118, N2999);
buf BUF1 (N17473, N17472);
nand NAND4 (N17474, N17468, N2988, N1102, N7942);
and AND3 (N17475, N17450, N14896, N8550);
nand NAND3 (N17476, N17471, N10469, N10108);
nand NAND3 (N17477, N17474, N8505, N11885);
nand NAND2 (N17478, N17476, N10958);
and AND4 (N17479, N17464, N10952, N13688, N11609);
not NOT1 (N17480, N17467);
xor XOR2 (N17481, N17478, N16697);
or OR2 (N17482, N17480, N708);
and AND3 (N17483, N17466, N3593, N15558);
nor NOR3 (N17484, N17477, N6037, N12034);
xor XOR2 (N17485, N17482, N16415);
nor NOR2 (N17486, N17484, N16845);
or OR2 (N17487, N17465, N12272);
nand NAND2 (N17488, N17479, N17141);
nand NAND3 (N17489, N17487, N12846, N10793);
nand NAND3 (N17490, N17485, N6399, N3678);
or OR2 (N17491, N17490, N11489);
or OR3 (N17492, N17473, N5247, N11442);
nand NAND4 (N17493, N17489, N6758, N11808, N4304);
xor XOR2 (N17494, N17475, N16946);
nand NAND4 (N17495, N17491, N12713, N12947, N1158);
and AND2 (N17496, N17495, N16362);
and AND3 (N17497, N17488, N12326, N16634);
not NOT1 (N17498, N17483);
buf BUF1 (N17499, N17493);
not NOT1 (N17500, N17481);
buf BUF1 (N17501, N17486);
not NOT1 (N17502, N17500);
and AND3 (N17503, N17469, N2142, N17249);
xor XOR2 (N17504, N17503, N3687);
nor NOR4 (N17505, N17492, N9426, N13044, N4110);
xor XOR2 (N17506, N17498, N14875);
nand NAND3 (N17507, N17505, N4767, N1237);
not NOT1 (N17508, N17502);
xor XOR2 (N17509, N17508, N1310);
or OR2 (N17510, N17501, N14287);
and AND3 (N17511, N17496, N3509, N6221);
not NOT1 (N17512, N17509);
xor XOR2 (N17513, N17510, N12573);
nor NOR4 (N17514, N17494, N4248, N4701, N244);
buf BUF1 (N17515, N17449);
or OR2 (N17516, N17511, N13485);
and AND3 (N17517, N17513, N2452, N12295);
xor XOR2 (N17518, N17506, N15707);
nor NOR4 (N17519, N17517, N14895, N2132, N12003);
nor NOR4 (N17520, N17516, N4513, N624, N3078);
and AND4 (N17521, N17504, N10688, N3647, N1459);
or OR4 (N17522, N17518, N14325, N9305, N16381);
nand NAND4 (N17523, N17515, N9200, N2518, N11251);
buf BUF1 (N17524, N17507);
and AND3 (N17525, N17521, N12574, N1994);
and AND4 (N17526, N17524, N5713, N14025, N11448);
not NOT1 (N17527, N17514);
nand NAND2 (N17528, N17523, N4178);
nor NOR4 (N17529, N17528, N7392, N11747, N8192);
or OR3 (N17530, N17497, N6512, N14502);
buf BUF1 (N17531, N17527);
nor NOR4 (N17532, N17529, N2246, N1380, N17314);
not NOT1 (N17533, N17522);
or OR4 (N17534, N17532, N674, N12346, N2615);
not NOT1 (N17535, N17525);
nand NAND3 (N17536, N17531, N8803, N5467);
nor NOR2 (N17537, N17512, N14181);
nand NAND2 (N17538, N17536, N12104);
nand NAND4 (N17539, N17526, N13351, N644, N11598);
buf BUF1 (N17540, N17539);
and AND3 (N17541, N17534, N10551, N9531);
xor XOR2 (N17542, N17535, N259);
and AND3 (N17543, N17538, N4255, N9400);
or OR2 (N17544, N17530, N780);
nand NAND2 (N17545, N17537, N3767);
xor XOR2 (N17546, N17540, N7848);
nor NOR3 (N17547, N17541, N2441, N7245);
or OR2 (N17548, N17520, N10802);
xor XOR2 (N17549, N17548, N7567);
nor NOR3 (N17550, N17546, N7525, N13685);
nor NOR2 (N17551, N17549, N14136);
nand NAND3 (N17552, N17551, N12850, N16521);
buf BUF1 (N17553, N17519);
or OR4 (N17554, N17533, N11180, N9968, N1540);
nand NAND3 (N17555, N17542, N1362, N4684);
not NOT1 (N17556, N17544);
nand NAND3 (N17557, N17543, N5954, N4515);
buf BUF1 (N17558, N17554);
nor NOR3 (N17559, N17550, N8519, N957);
nor NOR3 (N17560, N17547, N7457, N6570);
or OR2 (N17561, N17560, N13067);
and AND2 (N17562, N17552, N11121);
and AND3 (N17563, N17545, N12187, N9267);
nor NOR3 (N17564, N17556, N11092, N5290);
nor NOR4 (N17565, N17559, N10001, N5320, N5516);
xor XOR2 (N17566, N17563, N16070);
buf BUF1 (N17567, N17562);
or OR3 (N17568, N17499, N593, N13123);
nand NAND3 (N17569, N17557, N2203, N14572);
and AND4 (N17570, N17569, N10335, N4057, N2164);
buf BUF1 (N17571, N17568);
or OR4 (N17572, N17558, N1124, N9506, N17283);
nand NAND3 (N17573, N17564, N16631, N12756);
nand NAND4 (N17574, N17553, N15495, N11371, N12727);
nand NAND2 (N17575, N17574, N892);
nand NAND3 (N17576, N17566, N10772, N12942);
or OR2 (N17577, N17570, N9104);
nor NOR4 (N17578, N17575, N6960, N7079, N13592);
xor XOR2 (N17579, N17578, N9345);
nand NAND2 (N17580, N17567, N12220);
xor XOR2 (N17581, N17561, N12677);
not NOT1 (N17582, N17577);
or OR3 (N17583, N17573, N14745, N12514);
or OR3 (N17584, N17565, N11347, N7168);
or OR4 (N17585, N17572, N13906, N1949, N6820);
nand NAND3 (N17586, N17571, N2730, N9564);
buf BUF1 (N17587, N17579);
xor XOR2 (N17588, N17581, N8946);
xor XOR2 (N17589, N17586, N4990);
nor NOR4 (N17590, N17589, N15833, N14109, N1042);
or OR3 (N17591, N17585, N11076, N4869);
or OR2 (N17592, N17576, N1182);
xor XOR2 (N17593, N17591, N5110);
xor XOR2 (N17594, N17587, N16292);
not NOT1 (N17595, N17592);
nor NOR3 (N17596, N17555, N8382, N12529);
not NOT1 (N17597, N17582);
xor XOR2 (N17598, N17590, N14010);
and AND4 (N17599, N17596, N446, N17216, N17301);
and AND2 (N17600, N17588, N404);
buf BUF1 (N17601, N17597);
or OR2 (N17602, N17580, N7689);
and AND2 (N17603, N17599, N14001);
buf BUF1 (N17604, N17593);
buf BUF1 (N17605, N17604);
and AND3 (N17606, N17602, N5637, N6534);
buf BUF1 (N17607, N17603);
xor XOR2 (N17608, N17607, N265);
nor NOR4 (N17609, N17605, N7180, N1830, N2702);
buf BUF1 (N17610, N17594);
and AND2 (N17611, N17584, N4549);
nor NOR2 (N17612, N17601, N7629);
nor NOR4 (N17613, N17600, N7573, N169, N12470);
and AND4 (N17614, N17606, N13055, N1706, N7009);
or OR4 (N17615, N17608, N9729, N5705, N4814);
and AND3 (N17616, N17614, N9964, N2424);
nand NAND3 (N17617, N17611, N13707, N4242);
nor NOR4 (N17618, N17612, N12597, N201, N2822);
not NOT1 (N17619, N17598);
and AND4 (N17620, N17619, N6339, N2205, N6231);
not NOT1 (N17621, N17613);
and AND3 (N17622, N17620, N12219, N12036);
and AND4 (N17623, N17610, N9025, N9182, N14165);
not NOT1 (N17624, N17617);
xor XOR2 (N17625, N17622, N16159);
nand NAND2 (N17626, N17609, N5421);
nor NOR2 (N17627, N17615, N2898);
or OR3 (N17628, N17625, N5207, N9952);
nor NOR4 (N17629, N17595, N15163, N16867, N1841);
or OR4 (N17630, N17618, N4470, N15596, N126);
or OR4 (N17631, N17616, N2957, N3935, N842);
nand NAND3 (N17632, N17631, N15659, N1943);
buf BUF1 (N17633, N17628);
nor NOR4 (N17634, N17633, N5152, N3557, N3770);
and AND4 (N17635, N17629, N11751, N15376, N16978);
and AND4 (N17636, N17624, N5759, N9351, N9483);
nor NOR4 (N17637, N17630, N9658, N14844, N974);
or OR3 (N17638, N17634, N8494, N17424);
and AND2 (N17639, N17632, N429);
or OR3 (N17640, N17626, N5375, N17305);
not NOT1 (N17641, N17635);
and AND3 (N17642, N17636, N1663, N7368);
not NOT1 (N17643, N17641);
not NOT1 (N17644, N17623);
xor XOR2 (N17645, N17642, N1232);
and AND3 (N17646, N17645, N4018, N5853);
buf BUF1 (N17647, N17627);
nor NOR3 (N17648, N17621, N8083, N3491);
and AND4 (N17649, N17583, N7260, N5546, N3899);
or OR2 (N17650, N17637, N7500);
nor NOR2 (N17651, N17649, N16907);
nand NAND3 (N17652, N17644, N12817, N8363);
and AND3 (N17653, N17652, N14574, N11906);
and AND2 (N17654, N17638, N5242);
nand NAND4 (N17655, N17654, N2159, N15903, N13341);
nand NAND4 (N17656, N17655, N11939, N5568, N7965);
and AND2 (N17657, N17646, N14536);
not NOT1 (N17658, N17643);
buf BUF1 (N17659, N17648);
xor XOR2 (N17660, N17647, N8413);
nand NAND2 (N17661, N17640, N13135);
nand NAND4 (N17662, N17653, N4749, N2082, N9102);
and AND2 (N17663, N17661, N10615);
and AND4 (N17664, N17650, N769, N2825, N10269);
not NOT1 (N17665, N17656);
nor NOR4 (N17666, N17651, N8118, N7370, N2025);
nor NOR3 (N17667, N17663, N2906, N9750);
buf BUF1 (N17668, N17658);
or OR4 (N17669, N17662, N10826, N6436, N357);
xor XOR2 (N17670, N17667, N744);
not NOT1 (N17671, N17660);
nand NAND4 (N17672, N17657, N17051, N16044, N3569);
xor XOR2 (N17673, N17659, N16983);
xor XOR2 (N17674, N17672, N1097);
nand NAND3 (N17675, N17673, N4062, N4311);
not NOT1 (N17676, N17674);
or OR3 (N17677, N17669, N14123, N16654);
not NOT1 (N17678, N17675);
or OR2 (N17679, N17668, N4458);
or OR2 (N17680, N17671, N15651);
nor NOR3 (N17681, N17639, N13668, N11371);
xor XOR2 (N17682, N17680, N10239);
not NOT1 (N17683, N17664);
nand NAND4 (N17684, N17682, N8342, N2926, N5001);
nand NAND3 (N17685, N17681, N4314, N17144);
and AND3 (N17686, N17666, N9390, N14496);
and AND4 (N17687, N17685, N17491, N10413, N7635);
and AND3 (N17688, N17676, N8995, N16151);
and AND4 (N17689, N17665, N15736, N16408, N11093);
not NOT1 (N17690, N17683);
or OR3 (N17691, N17677, N17319, N997);
or OR3 (N17692, N17689, N14308, N1140);
buf BUF1 (N17693, N17678);
buf BUF1 (N17694, N17691);
xor XOR2 (N17695, N17684, N895);
not NOT1 (N17696, N17692);
not NOT1 (N17697, N17695);
or OR4 (N17698, N17688, N7475, N9865, N102);
nand NAND2 (N17699, N17693, N15671);
xor XOR2 (N17700, N17679, N9941);
not NOT1 (N17701, N17694);
xor XOR2 (N17702, N17700, N13360);
buf BUF1 (N17703, N17696);
not NOT1 (N17704, N17702);
and AND4 (N17705, N17699, N14548, N8278, N17631);
nor NOR3 (N17706, N17670, N12255, N949);
nand NAND2 (N17707, N17704, N17235);
nor NOR2 (N17708, N17705, N13537);
nand NAND2 (N17709, N17686, N4237);
buf BUF1 (N17710, N17698);
nand NAND4 (N17711, N17707, N12218, N2790, N15297);
or OR3 (N17712, N17703, N6283, N16276);
and AND2 (N17713, N17708, N4255);
xor XOR2 (N17714, N17701, N15138);
xor XOR2 (N17715, N17697, N4152);
buf BUF1 (N17716, N17690);
nand NAND4 (N17717, N17687, N6237, N6477, N17155);
not NOT1 (N17718, N17717);
nand NAND2 (N17719, N17718, N1238);
not NOT1 (N17720, N17712);
nor NOR3 (N17721, N17715, N13169, N6713);
or OR4 (N17722, N17721, N14657, N17237, N4493);
or OR2 (N17723, N17716, N14499);
nand NAND2 (N17724, N17709, N1964);
xor XOR2 (N17725, N17719, N3480);
buf BUF1 (N17726, N17706);
or OR2 (N17727, N17713, N10576);
xor XOR2 (N17728, N17723, N8884);
nor NOR4 (N17729, N17720, N5865, N6320, N10498);
or OR3 (N17730, N17711, N11307, N7406);
and AND3 (N17731, N17729, N3919, N4686);
not NOT1 (N17732, N17710);
and AND2 (N17733, N17726, N8702);
nand NAND3 (N17734, N17727, N1045, N10591);
nor NOR4 (N17735, N17733, N9848, N5485, N9532);
xor XOR2 (N17736, N17725, N2918);
and AND2 (N17737, N17722, N3297);
nor NOR2 (N17738, N17731, N47);
nor NOR2 (N17739, N17724, N16645);
not NOT1 (N17740, N17736);
not NOT1 (N17741, N17728);
not NOT1 (N17742, N17741);
and AND2 (N17743, N17737, N5460);
not NOT1 (N17744, N17740);
xor XOR2 (N17745, N17739, N14703);
nand NAND3 (N17746, N17734, N1557, N7542);
and AND3 (N17747, N17735, N10468, N2251);
not NOT1 (N17748, N17738);
nor NOR3 (N17749, N17746, N13754, N13387);
nor NOR4 (N17750, N17714, N5755, N12674, N13323);
buf BUF1 (N17751, N17745);
xor XOR2 (N17752, N17730, N6395);
nor NOR2 (N17753, N17750, N195);
xor XOR2 (N17754, N17748, N8261);
or OR3 (N17755, N17749, N5610, N2217);
nand NAND4 (N17756, N17747, N283, N1790, N8262);
not NOT1 (N17757, N17756);
and AND4 (N17758, N17754, N17732, N9317, N8231);
xor XOR2 (N17759, N8605, N14835);
and AND4 (N17760, N17752, N8723, N9972, N8383);
or OR3 (N17761, N17751, N7771, N12108);
buf BUF1 (N17762, N17759);
nor NOR3 (N17763, N17761, N4137, N11338);
and AND2 (N17764, N17762, N10025);
and AND4 (N17765, N17763, N11992, N8064, N4468);
xor XOR2 (N17766, N17743, N11637);
nor NOR2 (N17767, N17760, N15094);
xor XOR2 (N17768, N17767, N3730);
xor XOR2 (N17769, N17755, N3580);
xor XOR2 (N17770, N17753, N13742);
and AND3 (N17771, N17769, N15568, N2931);
not NOT1 (N17772, N17770);
not NOT1 (N17773, N17766);
or OR4 (N17774, N17757, N2054, N11323, N1557);
nand NAND4 (N17775, N17768, N13618, N5029, N13421);
and AND3 (N17776, N17773, N9771, N10707);
buf BUF1 (N17777, N17764);
and AND4 (N17778, N17774, N3657, N7668, N15267);
xor XOR2 (N17779, N17758, N4888);
nor NOR3 (N17780, N17776, N11311, N633);
or OR3 (N17781, N17765, N8083, N3678);
xor XOR2 (N17782, N17742, N2307);
nor NOR4 (N17783, N17781, N7655, N9963, N4095);
buf BUF1 (N17784, N17771);
or OR2 (N17785, N17744, N3555);
or OR4 (N17786, N17779, N1314, N1750, N2896);
xor XOR2 (N17787, N17785, N12409);
and AND2 (N17788, N17782, N16522);
and AND4 (N17789, N17780, N9923, N7656, N16537);
nor NOR2 (N17790, N17783, N9629);
nor NOR4 (N17791, N17787, N7099, N9339, N2310);
nand NAND2 (N17792, N17775, N4403);
not NOT1 (N17793, N17790);
nor NOR3 (N17794, N17792, N14187, N2583);
and AND4 (N17795, N17794, N1482, N13360, N6055);
buf BUF1 (N17796, N17777);
nand NAND2 (N17797, N17788, N12455);
nor NOR3 (N17798, N17778, N3698, N424);
not NOT1 (N17799, N17796);
and AND2 (N17800, N17784, N11943);
or OR4 (N17801, N17797, N4627, N8831, N1244);
xor XOR2 (N17802, N17801, N7593);
and AND2 (N17803, N17800, N12436);
nand NAND4 (N17804, N17772, N14821, N4448, N17086);
or OR2 (N17805, N17798, N15513);
xor XOR2 (N17806, N17805, N9866);
nand NAND4 (N17807, N17789, N4491, N5891, N14985);
nor NOR3 (N17808, N17803, N3929, N14091);
not NOT1 (N17809, N17802);
xor XOR2 (N17810, N17807, N4631);
and AND3 (N17811, N17793, N10349, N1531);
not NOT1 (N17812, N17810);
and AND4 (N17813, N17808, N7172, N3802, N3166);
nand NAND4 (N17814, N17812, N9005, N11194, N10791);
xor XOR2 (N17815, N17791, N2505);
xor XOR2 (N17816, N17813, N1399);
nor NOR4 (N17817, N17814, N5917, N15993, N11895);
nor NOR4 (N17818, N17795, N8018, N13505, N7388);
buf BUF1 (N17819, N17786);
not NOT1 (N17820, N17811);
or OR2 (N17821, N17804, N761);
xor XOR2 (N17822, N17821, N11757);
nand NAND4 (N17823, N17822, N14337, N3307, N14014);
buf BUF1 (N17824, N17806);
nand NAND3 (N17825, N17824, N14045, N7572);
buf BUF1 (N17826, N17818);
or OR4 (N17827, N17823, N14149, N4875, N2726);
not NOT1 (N17828, N17809);
xor XOR2 (N17829, N17819, N13105);
buf BUF1 (N17830, N17826);
and AND3 (N17831, N17829, N9734, N5493);
xor XOR2 (N17832, N17820, N15686);
buf BUF1 (N17833, N17799);
nor NOR2 (N17834, N17816, N6556);
nand NAND3 (N17835, N17833, N1333, N9214);
or OR2 (N17836, N17830, N6742);
nor NOR4 (N17837, N17827, N8321, N13987, N2242);
nor NOR3 (N17838, N17828, N6488, N3658);
buf BUF1 (N17839, N17836);
xor XOR2 (N17840, N17815, N1037);
or OR4 (N17841, N17840, N16821, N5228, N8667);
buf BUF1 (N17842, N17835);
nand NAND2 (N17843, N17832, N6124);
or OR4 (N17844, N17831, N12906, N1522, N14996);
nand NAND2 (N17845, N17838, N6411);
xor XOR2 (N17846, N17834, N17138);
nor NOR2 (N17847, N17825, N14973);
and AND3 (N17848, N17817, N6676, N664);
nor NOR3 (N17849, N17844, N2350, N16823);
not NOT1 (N17850, N17846);
and AND2 (N17851, N17842, N13337);
and AND2 (N17852, N17847, N2378);
nand NAND3 (N17853, N17837, N8429, N6611);
nand NAND4 (N17854, N17839, N17139, N16046, N6956);
not NOT1 (N17855, N17851);
not NOT1 (N17856, N17854);
buf BUF1 (N17857, N17848);
buf BUF1 (N17858, N17856);
not NOT1 (N17859, N17858);
and AND4 (N17860, N17850, N3235, N10090, N10234);
or OR3 (N17861, N17845, N6058, N14630);
nor NOR3 (N17862, N17852, N1438, N17748);
and AND4 (N17863, N17859, N16006, N17462, N11160);
and AND3 (N17864, N17843, N10032, N13182);
xor XOR2 (N17865, N17864, N3836);
and AND2 (N17866, N17841, N13566);
or OR4 (N17867, N17861, N8382, N8489, N15647);
nand NAND4 (N17868, N17855, N7936, N10987, N17406);
nor NOR4 (N17869, N17849, N762, N8303, N12147);
buf BUF1 (N17870, N17857);
or OR4 (N17871, N17869, N11775, N1392, N336);
buf BUF1 (N17872, N17862);
nand NAND4 (N17873, N17872, N16223, N3325, N10310);
buf BUF1 (N17874, N17853);
nand NAND2 (N17875, N17866, N2625);
and AND2 (N17876, N17868, N5835);
nand NAND3 (N17877, N17865, N16860, N5448);
xor XOR2 (N17878, N17860, N7982);
buf BUF1 (N17879, N17878);
xor XOR2 (N17880, N17871, N11434);
or OR3 (N17881, N17877, N8199, N9368);
nand NAND4 (N17882, N17874, N4370, N16272, N9445);
and AND2 (N17883, N17873, N4542);
or OR2 (N17884, N17863, N12397);
not NOT1 (N17885, N17876);
or OR2 (N17886, N17879, N3686);
or OR3 (N17887, N17886, N5738, N13930);
not NOT1 (N17888, N17870);
buf BUF1 (N17889, N17875);
xor XOR2 (N17890, N17888, N11985);
nand NAND4 (N17891, N17885, N8219, N7780, N2640);
xor XOR2 (N17892, N17883, N1313);
nand NAND4 (N17893, N17892, N17284, N8501, N504);
not NOT1 (N17894, N17867);
nor NOR3 (N17895, N17880, N622, N9629);
not NOT1 (N17896, N17890);
nand NAND3 (N17897, N17896, N7694, N4847);
xor XOR2 (N17898, N17895, N11634);
xor XOR2 (N17899, N17882, N13130);
or OR3 (N17900, N17897, N9415, N9355);
nand NAND3 (N17901, N17891, N10981, N12496);
not NOT1 (N17902, N17893);
xor XOR2 (N17903, N17901, N379);
or OR4 (N17904, N17899, N8232, N16187, N14657);
buf BUF1 (N17905, N17894);
nand NAND2 (N17906, N17884, N10875);
or OR3 (N17907, N17889, N5253, N5614);
nand NAND4 (N17908, N17906, N2934, N5684, N8135);
nor NOR4 (N17909, N17908, N10475, N5936, N7813);
or OR3 (N17910, N17902, N1944, N12780);
and AND3 (N17911, N17887, N12499, N15598);
buf BUF1 (N17912, N17898);
xor XOR2 (N17913, N17881, N10279);
nand NAND2 (N17914, N17911, N307);
not NOT1 (N17915, N17907);
nand NAND2 (N17916, N17904, N131);
nand NAND3 (N17917, N17915, N13883, N14957);
buf BUF1 (N17918, N17903);
nand NAND3 (N17919, N17917, N10156, N9078);
nand NAND2 (N17920, N17910, N9030);
nor NOR3 (N17921, N17913, N3866, N16218);
buf BUF1 (N17922, N17900);
nor NOR2 (N17923, N17909, N11086);
nor NOR2 (N17924, N17905, N1436);
and AND4 (N17925, N17920, N2750, N6384, N5190);
buf BUF1 (N17926, N17921);
nor NOR2 (N17927, N17914, N10448);
not NOT1 (N17928, N17923);
buf BUF1 (N17929, N17918);
and AND4 (N17930, N17924, N13454, N5859, N12651);
nand NAND4 (N17931, N17919, N6987, N5796, N9632);
buf BUF1 (N17932, N17925);
xor XOR2 (N17933, N17922, N8825);
nand NAND4 (N17934, N17931, N11284, N10850, N9793);
nand NAND4 (N17935, N17930, N1089, N7992, N2323);
nand NAND2 (N17936, N17933, N13364);
nand NAND4 (N17937, N17935, N13458, N3417, N9401);
buf BUF1 (N17938, N17928);
not NOT1 (N17939, N17934);
nand NAND4 (N17940, N17937, N8221, N6712, N2474);
and AND4 (N17941, N17940, N8531, N9623, N1415);
or OR3 (N17942, N17926, N15589, N1513);
or OR2 (N17943, N17938, N16728);
not NOT1 (N17944, N17943);
buf BUF1 (N17945, N17929);
nor NOR2 (N17946, N17939, N11985);
nor NOR3 (N17947, N17936, N15726, N9751);
buf BUF1 (N17948, N17927);
not NOT1 (N17949, N17941);
or OR3 (N17950, N17949, N17821, N15391);
nor NOR4 (N17951, N17947, N2332, N17311, N16594);
nand NAND4 (N17952, N17912, N9182, N5181, N4299);
not NOT1 (N17953, N17945);
buf BUF1 (N17954, N17951);
xor XOR2 (N17955, N17950, N4254);
buf BUF1 (N17956, N17944);
not NOT1 (N17957, N17953);
nand NAND4 (N17958, N17956, N10393, N5858, N12497);
nor NOR4 (N17959, N17916, N4783, N10053, N14664);
and AND4 (N17960, N17959, N10728, N15490, N5072);
not NOT1 (N17961, N17957);
and AND3 (N17962, N17948, N1405, N16788);
and AND2 (N17963, N17960, N6481);
buf BUF1 (N17964, N17954);
or OR2 (N17965, N17962, N8166);
or OR4 (N17966, N17955, N3874, N15456, N50);
nand NAND4 (N17967, N17965, N12333, N5125, N11528);
not NOT1 (N17968, N17952);
not NOT1 (N17969, N17946);
nand NAND4 (N17970, N17958, N9737, N14973, N9135);
xor XOR2 (N17971, N17969, N17590);
buf BUF1 (N17972, N17970);
nand NAND3 (N17973, N17966, N17187, N13477);
nand NAND2 (N17974, N17967, N16339);
not NOT1 (N17975, N17973);
or OR4 (N17976, N17974, N10282, N16463, N8401);
and AND3 (N17977, N17972, N13642, N471);
xor XOR2 (N17978, N17942, N8681);
buf BUF1 (N17979, N17976);
xor XOR2 (N17980, N17977, N10925);
and AND2 (N17981, N17975, N10642);
and AND4 (N17982, N17971, N14797, N14410, N5340);
not NOT1 (N17983, N17979);
xor XOR2 (N17984, N17980, N11377);
xor XOR2 (N17985, N17982, N8598);
not NOT1 (N17986, N17932);
nand NAND3 (N17987, N17981, N12955, N14068);
nor NOR3 (N17988, N17987, N4707, N10464);
not NOT1 (N17989, N17964);
nand NAND2 (N17990, N17986, N14314);
buf BUF1 (N17991, N17985);
buf BUF1 (N17992, N17989);
buf BUF1 (N17993, N17990);
and AND4 (N17994, N17993, N12466, N14725, N2257);
nand NAND2 (N17995, N17988, N6196);
nand NAND4 (N17996, N17983, N12195, N3788, N4174);
xor XOR2 (N17997, N17978, N17478);
nand NAND3 (N17998, N17968, N8797, N2458);
or OR2 (N17999, N17961, N17079);
or OR4 (N18000, N17984, N7958, N6076, N7133);
not NOT1 (N18001, N17992);
nor NOR2 (N18002, N17991, N6198);
and AND3 (N18003, N17994, N1402, N539);
buf BUF1 (N18004, N18001);
or OR4 (N18005, N17996, N8051, N7573, N1100);
and AND4 (N18006, N18005, N11981, N15875, N5003);
nand NAND4 (N18007, N18000, N2778, N15275, N11520);
nor NOR3 (N18008, N17999, N13141, N2778);
not NOT1 (N18009, N17995);
and AND2 (N18010, N17998, N8373);
or OR4 (N18011, N18002, N7887, N11952, N5074);
buf BUF1 (N18012, N18010);
nor NOR3 (N18013, N18008, N4433, N17469);
xor XOR2 (N18014, N18011, N14176);
nor NOR4 (N18015, N18004, N11838, N16991, N15331);
nand NAND3 (N18016, N18013, N3285, N16486);
buf BUF1 (N18017, N18015);
buf BUF1 (N18018, N18016);
nand NAND4 (N18019, N18007, N15091, N10544, N4350);
buf BUF1 (N18020, N18019);
nor NOR2 (N18021, N18017, N723);
buf BUF1 (N18022, N18012);
or OR4 (N18023, N18009, N4541, N16597, N6188);
nor NOR2 (N18024, N18018, N325);
nor NOR4 (N18025, N18023, N16031, N12736, N6625);
nor NOR2 (N18026, N17997, N8229);
nor NOR3 (N18027, N18021, N2623, N14535);
or OR3 (N18028, N18022, N7548, N9291);
nor NOR2 (N18029, N18027, N10481);
nor NOR2 (N18030, N18026, N2116);
buf BUF1 (N18031, N17963);
and AND3 (N18032, N18020, N4447, N4124);
buf BUF1 (N18033, N18014);
xor XOR2 (N18034, N18029, N14113);
xor XOR2 (N18035, N18031, N5228);
nor NOR3 (N18036, N18028, N11457, N6543);
xor XOR2 (N18037, N18006, N4456);
nand NAND2 (N18038, N18024, N6724);
buf BUF1 (N18039, N18037);
or OR4 (N18040, N18035, N4121, N612, N14515);
xor XOR2 (N18041, N18033, N2917);
and AND3 (N18042, N18032, N3660, N5717);
and AND4 (N18043, N18039, N9388, N11284, N8275);
or OR4 (N18044, N18041, N13806, N3893, N17685);
and AND3 (N18045, N18040, N8222, N8292);
nor NOR4 (N18046, N18036, N2696, N7532, N4853);
and AND4 (N18047, N18042, N1830, N3605, N3845);
nand NAND3 (N18048, N18047, N16772, N10629);
and AND4 (N18049, N18043, N8138, N2897, N7599);
buf BUF1 (N18050, N18030);
not NOT1 (N18051, N18025);
nand NAND3 (N18052, N18046, N4221, N14846);
and AND4 (N18053, N18052, N13035, N17818, N187);
not NOT1 (N18054, N18038);
nor NOR2 (N18055, N18049, N11530);
nor NOR4 (N18056, N18048, N8066, N2966, N3421);
or OR2 (N18057, N18054, N3086);
not NOT1 (N18058, N18056);
or OR4 (N18059, N18055, N10345, N2735, N9110);
not NOT1 (N18060, N18053);
xor XOR2 (N18061, N18060, N9774);
nand NAND4 (N18062, N18034, N18052, N13799, N3419);
xor XOR2 (N18063, N18057, N8812);
or OR2 (N18064, N18044, N8803);
not NOT1 (N18065, N18050);
nand NAND2 (N18066, N18051, N16988);
buf BUF1 (N18067, N18061);
and AND3 (N18068, N18064, N8920, N10878);
buf BUF1 (N18069, N18068);
nand NAND2 (N18070, N18067, N4559);
nand NAND3 (N18071, N18065, N12491, N14059);
xor XOR2 (N18072, N18003, N13716);
nand NAND3 (N18073, N18066, N7612, N3066);
nor NOR2 (N18074, N18058, N4212);
or OR4 (N18075, N18074, N6011, N747, N14749);
nand NAND3 (N18076, N18071, N15360, N3829);
and AND4 (N18077, N18069, N2740, N13201, N544);
buf BUF1 (N18078, N18062);
xor XOR2 (N18079, N18076, N6365);
buf BUF1 (N18080, N18073);
xor XOR2 (N18081, N18079, N7187);
nor NOR2 (N18082, N18059, N8875);
and AND3 (N18083, N18082, N17360, N8757);
nand NAND2 (N18084, N18063, N4425);
not NOT1 (N18085, N18080);
xor XOR2 (N18086, N18084, N6740);
buf BUF1 (N18087, N18078);
or OR4 (N18088, N18087, N69, N3302, N14935);
buf BUF1 (N18089, N18072);
nand NAND3 (N18090, N18086, N6420, N917);
not NOT1 (N18091, N18075);
buf BUF1 (N18092, N18088);
or OR4 (N18093, N18092, N16803, N8750, N945);
buf BUF1 (N18094, N18089);
not NOT1 (N18095, N18091);
or OR3 (N18096, N18094, N8682, N7422);
nand NAND4 (N18097, N18090, N3971, N5265, N15340);
and AND4 (N18098, N18096, N14747, N16395, N15167);
nand NAND2 (N18099, N18083, N12602);
or OR2 (N18100, N18098, N7689);
nand NAND2 (N18101, N18045, N6574);
nand NAND4 (N18102, N18101, N5274, N16561, N13287);
buf BUF1 (N18103, N18097);
buf BUF1 (N18104, N18103);
nand NAND4 (N18105, N18104, N9102, N17693, N12372);
and AND2 (N18106, N18102, N8088);
nor NOR2 (N18107, N18085, N1659);
nor NOR3 (N18108, N18093, N11471, N3374);
buf BUF1 (N18109, N18070);
nand NAND3 (N18110, N18077, N6441, N6480);
nor NOR2 (N18111, N18099, N4229);
not NOT1 (N18112, N18110);
nor NOR2 (N18113, N18095, N5543);
or OR4 (N18114, N18113, N8903, N10883, N7654);
and AND4 (N18115, N18105, N3042, N9813, N4795);
nand NAND4 (N18116, N18115, N2400, N299, N15758);
not NOT1 (N18117, N18109);
xor XOR2 (N18118, N18108, N13686);
or OR4 (N18119, N18116, N15169, N14616, N9961);
nand NAND4 (N18120, N18081, N13624, N12769, N10370);
not NOT1 (N18121, N18100);
or OR3 (N18122, N18107, N3197, N5899);
xor XOR2 (N18123, N18118, N9313);
not NOT1 (N18124, N18112);
and AND2 (N18125, N18117, N17759);
not NOT1 (N18126, N18111);
not NOT1 (N18127, N18106);
nand NAND2 (N18128, N18119, N9095);
or OR3 (N18129, N18123, N2135, N4558);
xor XOR2 (N18130, N18127, N1888);
not NOT1 (N18131, N18121);
xor XOR2 (N18132, N18120, N10276);
xor XOR2 (N18133, N18129, N15777);
buf BUF1 (N18134, N18131);
and AND4 (N18135, N18133, N1562, N5535, N11465);
not NOT1 (N18136, N18122);
nor NOR2 (N18137, N18132, N7292);
buf BUF1 (N18138, N18136);
xor XOR2 (N18139, N18126, N12859);
nor NOR4 (N18140, N18137, N2228, N11923, N7858);
and AND2 (N18141, N18135, N10508);
nor NOR2 (N18142, N18128, N14370);
and AND4 (N18143, N18140, N1503, N12586, N2143);
nor NOR2 (N18144, N18124, N6763);
nor NOR2 (N18145, N18144, N13574);
or OR3 (N18146, N18125, N11952, N8121);
xor XOR2 (N18147, N18139, N16587);
not NOT1 (N18148, N18114);
xor XOR2 (N18149, N18143, N3251);
xor XOR2 (N18150, N18134, N14762);
nor NOR4 (N18151, N18138, N10942, N16756, N259);
buf BUF1 (N18152, N18151);
nor NOR2 (N18153, N18142, N7550);
nor NOR4 (N18154, N18130, N4656, N4163, N9413);
not NOT1 (N18155, N18148);
and AND3 (N18156, N18154, N2605, N12722);
buf BUF1 (N18157, N18141);
buf BUF1 (N18158, N18147);
nor NOR3 (N18159, N18155, N17541, N17597);
not NOT1 (N18160, N18150);
nand NAND3 (N18161, N18158, N5048, N8874);
or OR4 (N18162, N18145, N17191, N10903, N1019);
buf BUF1 (N18163, N18159);
or OR4 (N18164, N18161, N9778, N9170, N14780);
nor NOR3 (N18165, N18164, N6825, N9433);
not NOT1 (N18166, N18156);
nand NAND4 (N18167, N18160, N6766, N14903, N1052);
not NOT1 (N18168, N18162);
nor NOR4 (N18169, N18165, N15013, N9228, N2007);
xor XOR2 (N18170, N18157, N10562);
xor XOR2 (N18171, N18170, N8312);
nor NOR4 (N18172, N18146, N2467, N8996, N12422);
xor XOR2 (N18173, N18168, N7475);
nor NOR3 (N18174, N18172, N267, N15762);
nor NOR4 (N18175, N18167, N98, N11967, N12649);
buf BUF1 (N18176, N18166);
not NOT1 (N18177, N18175);
buf BUF1 (N18178, N18173);
or OR4 (N18179, N18163, N7880, N12349, N15865);
buf BUF1 (N18180, N18176);
and AND4 (N18181, N18169, N12839, N11737, N2323);
not NOT1 (N18182, N18179);
or OR2 (N18183, N18178, N10886);
buf BUF1 (N18184, N18152);
and AND2 (N18185, N18183, N16559);
or OR2 (N18186, N18153, N13887);
and AND3 (N18187, N18177, N15741, N2287);
and AND2 (N18188, N18184, N16395);
nand NAND3 (N18189, N18174, N5003, N2451);
nor NOR4 (N18190, N18149, N11378, N7139, N12000);
not NOT1 (N18191, N18182);
not NOT1 (N18192, N18186);
or OR4 (N18193, N18171, N5348, N745, N11520);
xor XOR2 (N18194, N18185, N16113);
or OR3 (N18195, N18188, N10273, N2837);
nand NAND4 (N18196, N18181, N16859, N897, N16550);
or OR2 (N18197, N18191, N1248);
xor XOR2 (N18198, N18197, N7136);
or OR3 (N18199, N18187, N17189, N3829);
buf BUF1 (N18200, N18195);
not NOT1 (N18201, N18198);
or OR4 (N18202, N18201, N16553, N17185, N16693);
and AND4 (N18203, N18200, N9891, N11104, N8913);
nor NOR2 (N18204, N18199, N14275);
and AND3 (N18205, N18202, N15325, N10597);
nand NAND3 (N18206, N18196, N10971, N11725);
or OR2 (N18207, N18206, N10427);
nor NOR2 (N18208, N18205, N4089);
not NOT1 (N18209, N18208);
xor XOR2 (N18210, N18203, N3936);
or OR2 (N18211, N18194, N15528);
not NOT1 (N18212, N18210);
not NOT1 (N18213, N18180);
nor NOR4 (N18214, N18190, N11871, N11979, N13046);
and AND4 (N18215, N18214, N15177, N7199, N1291);
xor XOR2 (N18216, N18192, N9364);
not NOT1 (N18217, N18204);
or OR4 (N18218, N18193, N3608, N9422, N7680);
buf BUF1 (N18219, N18211);
or OR4 (N18220, N18215, N16655, N11174, N13907);
nor NOR4 (N18221, N18207, N14466, N18010, N3902);
xor XOR2 (N18222, N18212, N13152);
buf BUF1 (N18223, N18222);
buf BUF1 (N18224, N18217);
not NOT1 (N18225, N18223);
or OR4 (N18226, N18218, N9121, N17120, N18046);
or OR4 (N18227, N18225, N14973, N13625, N7604);
xor XOR2 (N18228, N18224, N4041);
or OR4 (N18229, N18221, N7921, N4261, N12168);
buf BUF1 (N18230, N18209);
xor XOR2 (N18231, N18189, N4189);
and AND3 (N18232, N18219, N7478, N17247);
buf BUF1 (N18233, N18228);
nor NOR4 (N18234, N18227, N6144, N13870, N16339);
and AND2 (N18235, N18233, N7417);
or OR2 (N18236, N18232, N5339);
xor XOR2 (N18237, N18229, N16483);
xor XOR2 (N18238, N18235, N2669);
or OR3 (N18239, N18226, N1994, N15687);
buf BUF1 (N18240, N18220);
not NOT1 (N18241, N18231);
nor NOR3 (N18242, N18241, N9178, N16466);
xor XOR2 (N18243, N18242, N11204);
not NOT1 (N18244, N18237);
nor NOR2 (N18245, N18236, N12090);
nor NOR3 (N18246, N18239, N6823, N12934);
xor XOR2 (N18247, N18240, N17305);
xor XOR2 (N18248, N18244, N1124);
or OR3 (N18249, N18230, N200, N3816);
nor NOR4 (N18250, N18247, N5561, N11592, N12461);
and AND4 (N18251, N18248, N12962, N14016, N17398);
or OR2 (N18252, N18234, N17052);
nand NAND4 (N18253, N18252, N17797, N942, N13678);
and AND3 (N18254, N18250, N7753, N17096);
and AND3 (N18255, N18213, N2033, N7843);
or OR2 (N18256, N18238, N16593);
or OR3 (N18257, N18216, N11233, N9060);
xor XOR2 (N18258, N18245, N2603);
xor XOR2 (N18259, N18246, N5405);
or OR4 (N18260, N18255, N9242, N17864, N9891);
nor NOR4 (N18261, N18243, N12774, N17884, N17612);
xor XOR2 (N18262, N18254, N5738);
xor XOR2 (N18263, N18261, N10867);
not NOT1 (N18264, N18257);
or OR2 (N18265, N18253, N324);
xor XOR2 (N18266, N18256, N3995);
nand NAND2 (N18267, N18265, N10744);
nor NOR2 (N18268, N18266, N2772);
and AND3 (N18269, N18268, N14022, N13521);
nand NAND3 (N18270, N18263, N9450, N13718);
xor XOR2 (N18271, N18264, N6879);
or OR2 (N18272, N18249, N14407);
nand NAND4 (N18273, N18270, N874, N5513, N10459);
and AND2 (N18274, N18260, N15777);
buf BUF1 (N18275, N18273);
xor XOR2 (N18276, N18267, N8118);
nand NAND4 (N18277, N18271, N8057, N11698, N14468);
or OR3 (N18278, N18276, N3639, N7274);
xor XOR2 (N18279, N18278, N1868);
nand NAND4 (N18280, N18258, N6981, N4589, N17801);
xor XOR2 (N18281, N18269, N11682);
or OR4 (N18282, N18275, N7560, N5964, N8345);
and AND2 (N18283, N18262, N3761);
xor XOR2 (N18284, N18274, N17878);
buf BUF1 (N18285, N18280);
nand NAND4 (N18286, N18281, N6402, N12242, N14890);
or OR4 (N18287, N18282, N11728, N8275, N10624);
and AND4 (N18288, N18251, N5608, N4012, N3983);
xor XOR2 (N18289, N18288, N8285);
nor NOR3 (N18290, N18283, N16429, N7038);
not NOT1 (N18291, N18289);
nor NOR3 (N18292, N18272, N4898, N8066);
nand NAND3 (N18293, N18286, N7580, N15847);
or OR2 (N18294, N18285, N2445);
not NOT1 (N18295, N18292);
and AND3 (N18296, N18277, N12757, N7842);
xor XOR2 (N18297, N18293, N13338);
or OR3 (N18298, N18297, N9357, N3478);
and AND2 (N18299, N18290, N2730);
or OR2 (N18300, N18284, N1732);
and AND4 (N18301, N18300, N6752, N9157, N17533);
xor XOR2 (N18302, N18296, N11782);
not NOT1 (N18303, N18291);
xor XOR2 (N18304, N18299, N14677);
or OR4 (N18305, N18298, N4836, N354, N1176);
nor NOR4 (N18306, N18295, N3953, N6721, N1134);
nand NAND2 (N18307, N18294, N9880);
nor NOR2 (N18308, N18304, N10294);
and AND4 (N18309, N18303, N7981, N11881, N4760);
nor NOR2 (N18310, N18279, N1098);
nand NAND3 (N18311, N18308, N12867, N17703);
xor XOR2 (N18312, N18309, N9534);
not NOT1 (N18313, N18302);
buf BUF1 (N18314, N18312);
xor XOR2 (N18315, N18306, N7224);
buf BUF1 (N18316, N18259);
nor NOR2 (N18317, N18305, N9239);
buf BUF1 (N18318, N18301);
or OR4 (N18319, N18317, N3821, N199, N6770);
nor NOR3 (N18320, N18316, N11191, N1631);
buf BUF1 (N18321, N18313);
xor XOR2 (N18322, N18319, N1292);
xor XOR2 (N18323, N18315, N6980);
xor XOR2 (N18324, N18321, N13541);
buf BUF1 (N18325, N18287);
not NOT1 (N18326, N18323);
xor XOR2 (N18327, N18310, N5011);
nor NOR3 (N18328, N18322, N6969, N8239);
xor XOR2 (N18329, N18328, N14692);
xor XOR2 (N18330, N18326, N1665);
and AND2 (N18331, N18325, N14423);
nand NAND3 (N18332, N18320, N3446, N4073);
or OR4 (N18333, N18307, N16277, N4908, N12513);
and AND3 (N18334, N18329, N1731, N1860);
or OR2 (N18335, N18311, N4786);
or OR3 (N18336, N18332, N6719, N18323);
not NOT1 (N18337, N18336);
nor NOR4 (N18338, N18314, N10317, N17647, N15949);
or OR2 (N18339, N18333, N2136);
buf BUF1 (N18340, N18324);
nand NAND3 (N18341, N18335, N6733, N12529);
nor NOR4 (N18342, N18327, N2497, N11999, N4612);
xor XOR2 (N18343, N18318, N13346);
nor NOR4 (N18344, N18334, N15868, N4651, N6951);
nand NAND2 (N18345, N18341, N9959);
not NOT1 (N18346, N18344);
nand NAND4 (N18347, N18345, N3258, N12908, N12354);
and AND3 (N18348, N18337, N2185, N10952);
not NOT1 (N18349, N18340);
nor NOR4 (N18350, N18330, N14834, N16759, N3862);
not NOT1 (N18351, N18349);
or OR4 (N18352, N18348, N1663, N11566, N3998);
and AND3 (N18353, N18338, N1413, N16975);
xor XOR2 (N18354, N18350, N17536);
xor XOR2 (N18355, N18339, N7641);
or OR2 (N18356, N18347, N16195);
nor NOR4 (N18357, N18342, N6832, N1597, N9628);
buf BUF1 (N18358, N18346);
or OR4 (N18359, N18352, N17514, N18327, N15800);
not NOT1 (N18360, N18331);
and AND2 (N18361, N18357, N16901);
buf BUF1 (N18362, N18355);
not NOT1 (N18363, N18356);
not NOT1 (N18364, N18353);
and AND3 (N18365, N18364, N5983, N4370);
nor NOR3 (N18366, N18363, N15904, N9970);
or OR4 (N18367, N18362, N1120, N4124, N2320);
not NOT1 (N18368, N18367);
and AND2 (N18369, N18343, N12350);
buf BUF1 (N18370, N18365);
not NOT1 (N18371, N18360);
not NOT1 (N18372, N18361);
and AND4 (N18373, N18369, N12850, N3204, N13103);
buf BUF1 (N18374, N18370);
nand NAND4 (N18375, N18372, N4494, N276, N12906);
buf BUF1 (N18376, N18375);
not NOT1 (N18377, N18358);
and AND4 (N18378, N18373, N10139, N16371, N14003);
not NOT1 (N18379, N18351);
or OR3 (N18380, N18378, N13133, N6130);
xor XOR2 (N18381, N18354, N15070);
not NOT1 (N18382, N18379);
and AND4 (N18383, N18374, N13559, N3497, N15348);
nand NAND4 (N18384, N18381, N6574, N6603, N15472);
nand NAND2 (N18385, N18359, N15145);
nor NOR3 (N18386, N18377, N2074, N9480);
nand NAND3 (N18387, N18368, N14458, N8420);
nor NOR3 (N18388, N18386, N11461, N17490);
xor XOR2 (N18389, N18388, N7605);
and AND3 (N18390, N18385, N14141, N8186);
or OR4 (N18391, N18383, N16724, N212, N15818);
xor XOR2 (N18392, N18387, N10080);
xor XOR2 (N18393, N18371, N4572);
nor NOR3 (N18394, N18391, N7832, N14970);
and AND3 (N18395, N18380, N15794, N12825);
buf BUF1 (N18396, N18384);
nand NAND3 (N18397, N18390, N17626, N12597);
nor NOR2 (N18398, N18389, N7509);
nor NOR2 (N18399, N18366, N3903);
xor XOR2 (N18400, N18393, N3712);
nor NOR2 (N18401, N18392, N10533);
nor NOR2 (N18402, N18397, N17522);
xor XOR2 (N18403, N18402, N17319);
xor XOR2 (N18404, N18400, N12234);
nor NOR4 (N18405, N18376, N1571, N5641, N17079);
xor XOR2 (N18406, N18405, N15232);
nor NOR2 (N18407, N18403, N2487);
xor XOR2 (N18408, N18396, N234);
or OR3 (N18409, N18404, N3695, N1477);
nor NOR2 (N18410, N18382, N4573);
xor XOR2 (N18411, N18409, N14788);
nand NAND2 (N18412, N18394, N8455);
not NOT1 (N18413, N18412);
xor XOR2 (N18414, N18406, N8850);
and AND2 (N18415, N18399, N11939);
nand NAND3 (N18416, N18395, N10485, N11591);
and AND2 (N18417, N18414, N9498);
or OR3 (N18418, N18398, N1575, N393);
xor XOR2 (N18419, N18418, N16047);
nand NAND2 (N18420, N18407, N9127);
xor XOR2 (N18421, N18408, N4623);
buf BUF1 (N18422, N18411);
xor XOR2 (N18423, N18417, N13228);
nand NAND4 (N18424, N18416, N9214, N16122, N7958);
buf BUF1 (N18425, N18401);
xor XOR2 (N18426, N18425, N6242);
or OR3 (N18427, N18426, N10552, N9427);
nand NAND2 (N18428, N18410, N1901);
buf BUF1 (N18429, N18423);
nor NOR2 (N18430, N18413, N8307);
nor NOR2 (N18431, N18428, N16501);
nand NAND3 (N18432, N18427, N11081, N8429);
nor NOR2 (N18433, N18431, N1438);
and AND3 (N18434, N18419, N15695, N13394);
nand NAND2 (N18435, N18424, N16745);
or OR2 (N18436, N18433, N3483);
not NOT1 (N18437, N18434);
buf BUF1 (N18438, N18435);
nand NAND3 (N18439, N18436, N660, N11865);
xor XOR2 (N18440, N18439, N5923);
xor XOR2 (N18441, N18438, N14267);
buf BUF1 (N18442, N18421);
or OR2 (N18443, N18442, N3591);
nor NOR3 (N18444, N18420, N6931, N9791);
buf BUF1 (N18445, N18444);
nand NAND3 (N18446, N18430, N4594, N10301);
xor XOR2 (N18447, N18429, N11372);
not NOT1 (N18448, N18415);
xor XOR2 (N18449, N18446, N4428);
not NOT1 (N18450, N18422);
buf BUF1 (N18451, N18450);
nor NOR2 (N18452, N18448, N7188);
and AND4 (N18453, N18451, N4714, N16148, N13331);
not NOT1 (N18454, N18437);
nor NOR2 (N18455, N18440, N8414);
not NOT1 (N18456, N18443);
or OR3 (N18457, N18452, N11916, N15480);
buf BUF1 (N18458, N18455);
nor NOR2 (N18459, N18453, N12634);
or OR4 (N18460, N18441, N8636, N14930, N4957);
nor NOR3 (N18461, N18458, N5642, N15056);
xor XOR2 (N18462, N18447, N9949);
nor NOR3 (N18463, N18454, N5665, N12237);
and AND4 (N18464, N18449, N6153, N5162, N11707);
or OR3 (N18465, N18456, N11094, N2900);
and AND4 (N18466, N18464, N11710, N8849, N9864);
and AND2 (N18467, N18445, N15475);
and AND3 (N18468, N18432, N4700, N3544);
and AND2 (N18469, N18460, N5484);
buf BUF1 (N18470, N18465);
xor XOR2 (N18471, N18468, N13682);
nand NAND2 (N18472, N18459, N907);
nor NOR3 (N18473, N18471, N5816, N7162);
not NOT1 (N18474, N18461);
nand NAND2 (N18475, N18462, N17671);
and AND3 (N18476, N18474, N14416, N15746);
buf BUF1 (N18477, N18463);
nor NOR3 (N18478, N18467, N3259, N3489);
nor NOR2 (N18479, N18457, N6439);
nor NOR4 (N18480, N18477, N6790, N13946, N16321);
and AND3 (N18481, N18480, N5486, N781);
buf BUF1 (N18482, N18470);
nor NOR4 (N18483, N18476, N9220, N2501, N13744);
not NOT1 (N18484, N18483);
xor XOR2 (N18485, N18472, N16994);
buf BUF1 (N18486, N18469);
nor NOR3 (N18487, N18475, N3105, N10401);
xor XOR2 (N18488, N18487, N1386);
not NOT1 (N18489, N18488);
and AND2 (N18490, N18473, N4158);
nand NAND3 (N18491, N18484, N2955, N12571);
nor NOR3 (N18492, N18482, N9574, N5450);
xor XOR2 (N18493, N18485, N9832);
and AND2 (N18494, N18466, N14988);
buf BUF1 (N18495, N18491);
not NOT1 (N18496, N18493);
nor NOR4 (N18497, N18496, N6247, N1066, N2475);
or OR3 (N18498, N18497, N3415, N15217);
and AND2 (N18499, N18489, N5803);
not NOT1 (N18500, N18498);
nand NAND3 (N18501, N18494, N16771, N11386);
and AND2 (N18502, N18490, N10105);
nor NOR2 (N18503, N18502, N11038);
nand NAND4 (N18504, N18503, N16220, N17114, N403);
and AND3 (N18505, N18486, N1565, N4838);
and AND2 (N18506, N18504, N1653);
xor XOR2 (N18507, N18479, N4512);
not NOT1 (N18508, N18507);
not NOT1 (N18509, N18500);
and AND3 (N18510, N18481, N4525, N7899);
not NOT1 (N18511, N18499);
and AND4 (N18512, N18505, N14852, N236, N16642);
xor XOR2 (N18513, N18495, N12499);
or OR2 (N18514, N18506, N16919);
and AND2 (N18515, N18513, N8453);
nand NAND4 (N18516, N18509, N9020, N3523, N9235);
or OR2 (N18517, N18508, N11430);
and AND4 (N18518, N18501, N3871, N16125, N9244);
nand NAND3 (N18519, N18516, N2200, N10486);
not NOT1 (N18520, N18512);
xor XOR2 (N18521, N18514, N5319);
nor NOR4 (N18522, N18515, N6525, N5663, N18450);
xor XOR2 (N18523, N18521, N15160);
buf BUF1 (N18524, N18523);
not NOT1 (N18525, N18478);
and AND4 (N18526, N18522, N5102, N5975, N13170);
not NOT1 (N18527, N18517);
or OR3 (N18528, N18518, N8321, N9527);
buf BUF1 (N18529, N18526);
buf BUF1 (N18530, N18527);
and AND2 (N18531, N18510, N1172);
and AND4 (N18532, N18520, N2144, N6200, N4868);
buf BUF1 (N18533, N18511);
xor XOR2 (N18534, N18530, N3120);
xor XOR2 (N18535, N18528, N13382);
nand NAND2 (N18536, N18519, N10448);
not NOT1 (N18537, N18492);
buf BUF1 (N18538, N18535);
and AND2 (N18539, N18538, N17776);
xor XOR2 (N18540, N18532, N3506);
xor XOR2 (N18541, N18525, N2831);
nor NOR2 (N18542, N18533, N12629);
nand NAND4 (N18543, N18542, N7083, N8492, N11536);
nand NAND2 (N18544, N18534, N14636);
and AND4 (N18545, N18541, N15003, N16293, N1300);
or OR2 (N18546, N18545, N10542);
xor XOR2 (N18547, N18539, N2277);
or OR2 (N18548, N18543, N1892);
and AND3 (N18549, N18544, N6876, N6700);
or OR2 (N18550, N18537, N12256);
and AND3 (N18551, N18540, N13436, N1079);
not NOT1 (N18552, N18551);
buf BUF1 (N18553, N18548);
nor NOR4 (N18554, N18547, N4686, N12822, N9701);
nand NAND3 (N18555, N18552, N11576, N1153);
xor XOR2 (N18556, N18536, N16163);
buf BUF1 (N18557, N18549);
and AND4 (N18558, N18524, N18301, N12900, N9159);
xor XOR2 (N18559, N18555, N2953);
nand NAND2 (N18560, N18554, N5890);
and AND4 (N18561, N18531, N18142, N4004, N15742);
xor XOR2 (N18562, N18529, N18366);
not NOT1 (N18563, N18557);
nand NAND3 (N18564, N18563, N15608, N11070);
xor XOR2 (N18565, N18559, N2894);
or OR2 (N18566, N18556, N6191);
and AND2 (N18567, N18564, N8079);
xor XOR2 (N18568, N18550, N5057);
nand NAND4 (N18569, N18568, N1564, N15684, N7689);
xor XOR2 (N18570, N18562, N9693);
nor NOR3 (N18571, N18569, N11329, N17105);
nand NAND4 (N18572, N18565, N4300, N2689, N10216);
or OR2 (N18573, N18546, N17171);
buf BUF1 (N18574, N18571);
xor XOR2 (N18575, N18567, N12761);
or OR2 (N18576, N18560, N8808);
and AND3 (N18577, N18561, N2954, N12638);
nor NOR4 (N18578, N18566, N17207, N2543, N1334);
nor NOR2 (N18579, N18575, N20);
xor XOR2 (N18580, N18577, N16279);
or OR2 (N18581, N18580, N11495);
or OR4 (N18582, N18576, N16359, N10187, N7195);
not NOT1 (N18583, N18572);
nor NOR4 (N18584, N18578, N14536, N16967, N3042);
buf BUF1 (N18585, N18579);
and AND4 (N18586, N18573, N10476, N11164, N17862);
nand NAND4 (N18587, N18574, N16666, N1624, N5217);
and AND4 (N18588, N18558, N2473, N9058, N12798);
buf BUF1 (N18589, N18585);
buf BUF1 (N18590, N18570);
buf BUF1 (N18591, N18553);
nand NAND4 (N18592, N18582, N3047, N5096, N5761);
nor NOR2 (N18593, N18592, N4095);
and AND4 (N18594, N18590, N16365, N2044, N836);
xor XOR2 (N18595, N18581, N2370);
or OR3 (N18596, N18589, N15431, N14234);
xor XOR2 (N18597, N18593, N3953);
nand NAND3 (N18598, N18586, N11878, N11593);
and AND4 (N18599, N18591, N17186, N16561, N10458);
buf BUF1 (N18600, N18588);
nand NAND3 (N18601, N18599, N7688, N9280);
not NOT1 (N18602, N18596);
nor NOR2 (N18603, N18602, N4809);
not NOT1 (N18604, N18584);
nor NOR4 (N18605, N18597, N9868, N9835, N8066);
or OR3 (N18606, N18601, N13229, N14284);
nor NOR2 (N18607, N18587, N8089);
not NOT1 (N18608, N18594);
buf BUF1 (N18609, N18603);
nor NOR4 (N18610, N18608, N12716, N12352, N8873);
nor NOR2 (N18611, N18610, N11582);
or OR2 (N18612, N18604, N2847);
nand NAND2 (N18613, N18607, N10870);
or OR2 (N18614, N18612, N12793);
and AND2 (N18615, N18598, N4347);
nor NOR2 (N18616, N18583, N6472);
nor NOR4 (N18617, N18613, N18429, N2915, N10913);
or OR2 (N18618, N18614, N13959);
or OR4 (N18619, N18615, N3596, N14725, N1731);
and AND2 (N18620, N18617, N10267);
not NOT1 (N18621, N18606);
not NOT1 (N18622, N18620);
and AND3 (N18623, N18616, N17666, N8169);
nor NOR4 (N18624, N18623, N4221, N8254, N9469);
nand NAND4 (N18625, N18619, N6220, N17027, N7660);
or OR4 (N18626, N18600, N6485, N15522, N9402);
buf BUF1 (N18627, N18625);
not NOT1 (N18628, N18595);
or OR4 (N18629, N18626, N3557, N7097, N62);
nand NAND3 (N18630, N18611, N620, N17293);
buf BUF1 (N18631, N18621);
and AND4 (N18632, N18618, N12450, N2568, N3334);
or OR4 (N18633, N18630, N13530, N17130, N3076);
and AND2 (N18634, N18627, N13091);
xor XOR2 (N18635, N18628, N12333);
xor XOR2 (N18636, N18622, N8197);
or OR4 (N18637, N18636, N3308, N3121, N16157);
and AND4 (N18638, N18631, N14598, N12354, N13597);
nor NOR3 (N18639, N18629, N603, N10421);
buf BUF1 (N18640, N18638);
buf BUF1 (N18641, N18634);
buf BUF1 (N18642, N18633);
xor XOR2 (N18643, N18640, N14279);
xor XOR2 (N18644, N18632, N6007);
and AND2 (N18645, N18637, N17600);
and AND3 (N18646, N18642, N11221, N8556);
and AND2 (N18647, N18644, N5415);
buf BUF1 (N18648, N18639);
xor XOR2 (N18649, N18624, N918);
nor NOR3 (N18650, N18605, N8408, N6211);
nand NAND4 (N18651, N18648, N12995, N3442, N5407);
buf BUF1 (N18652, N18641);
xor XOR2 (N18653, N18651, N491);
xor XOR2 (N18654, N18635, N12700);
buf BUF1 (N18655, N18647);
xor XOR2 (N18656, N18650, N5194);
and AND2 (N18657, N18609, N14606);
nor NOR2 (N18658, N18657, N1833);
or OR3 (N18659, N18649, N14703, N1217);
not NOT1 (N18660, N18653);
nand NAND3 (N18661, N18660, N5763, N4496);
and AND4 (N18662, N18655, N9740, N9555, N11091);
xor XOR2 (N18663, N18646, N16859);
or OR2 (N18664, N18661, N3828);
and AND4 (N18665, N18662, N16172, N286, N1101);
buf BUF1 (N18666, N18665);
not NOT1 (N18667, N18645);
not NOT1 (N18668, N18643);
not NOT1 (N18669, N18656);
xor XOR2 (N18670, N18658, N539);
buf BUF1 (N18671, N18654);
nor NOR2 (N18672, N18659, N9607);
buf BUF1 (N18673, N18672);
nand NAND3 (N18674, N18663, N2233, N9373);
and AND3 (N18675, N18667, N7848, N9652);
nand NAND2 (N18676, N18668, N14776);
nand NAND3 (N18677, N18675, N17022, N8473);
xor XOR2 (N18678, N18674, N16257);
not NOT1 (N18679, N18652);
nand NAND3 (N18680, N18678, N6747, N3627);
buf BUF1 (N18681, N18664);
or OR4 (N18682, N18669, N4852, N16507, N18058);
nor NOR2 (N18683, N18681, N5269);
nor NOR4 (N18684, N18677, N13886, N5127, N8243);
nand NAND2 (N18685, N18684, N16430);
xor XOR2 (N18686, N18671, N8854);
nor NOR2 (N18687, N18680, N698);
xor XOR2 (N18688, N18670, N15820);
nor NOR4 (N18689, N18673, N16334, N9318, N10229);
and AND3 (N18690, N18679, N14694, N3482);
buf BUF1 (N18691, N18690);
or OR2 (N18692, N18683, N10131);
nor NOR4 (N18693, N18691, N2169, N8412, N17314);
nor NOR4 (N18694, N18676, N1001, N17080, N493);
buf BUF1 (N18695, N18666);
not NOT1 (N18696, N18687);
buf BUF1 (N18697, N18696);
nor NOR4 (N18698, N18697, N589, N8077, N4800);
and AND4 (N18699, N18689, N16787, N629, N15288);
and AND3 (N18700, N18699, N16610, N4108);
and AND4 (N18701, N18685, N8257, N15490, N5607);
nand NAND4 (N18702, N18693, N11657, N16403, N1222);
nand NAND4 (N18703, N18692, N8630, N13281, N10792);
not NOT1 (N18704, N18688);
buf BUF1 (N18705, N18695);
xor XOR2 (N18706, N18698, N4486);
xor XOR2 (N18707, N18682, N9687);
not NOT1 (N18708, N18694);
buf BUF1 (N18709, N18701);
nand NAND3 (N18710, N18707, N10828, N9553);
or OR3 (N18711, N18710, N2333, N4648);
nor NOR3 (N18712, N18704, N2228, N18159);
xor XOR2 (N18713, N18706, N15352);
not NOT1 (N18714, N18702);
or OR3 (N18715, N18708, N14402, N4513);
not NOT1 (N18716, N18686);
and AND2 (N18717, N18700, N14859);
xor XOR2 (N18718, N18715, N9113);
and AND2 (N18719, N18712, N12291);
not NOT1 (N18720, N18709);
xor XOR2 (N18721, N18719, N18110);
xor XOR2 (N18722, N18718, N8983);
buf BUF1 (N18723, N18713);
not NOT1 (N18724, N18717);
and AND4 (N18725, N18724, N2295, N7970, N12578);
nor NOR2 (N18726, N18716, N692);
xor XOR2 (N18727, N18725, N7947);
buf BUF1 (N18728, N18726);
buf BUF1 (N18729, N18714);
buf BUF1 (N18730, N18722);
not NOT1 (N18731, N18711);
nor NOR2 (N18732, N18723, N14850);
not NOT1 (N18733, N18703);
nand NAND4 (N18734, N18727, N7005, N17179, N16724);
buf BUF1 (N18735, N18731);
or OR4 (N18736, N18721, N2864, N13761, N7547);
and AND2 (N18737, N18728, N6281);
and AND4 (N18738, N18735, N1842, N17481, N12877);
or OR2 (N18739, N18729, N7199);
and AND2 (N18740, N18730, N5765);
not NOT1 (N18741, N18733);
nor NOR2 (N18742, N18738, N5727);
xor XOR2 (N18743, N18742, N12374);
nor NOR2 (N18744, N18740, N18020);
xor XOR2 (N18745, N18705, N1287);
not NOT1 (N18746, N18741);
or OR2 (N18747, N18744, N11153);
xor XOR2 (N18748, N18746, N4317);
or OR3 (N18749, N18739, N7351, N7534);
not NOT1 (N18750, N18748);
and AND3 (N18751, N18720, N4232, N11055);
and AND4 (N18752, N18745, N918, N8476, N7350);
or OR4 (N18753, N18751, N4235, N10683, N3568);
xor XOR2 (N18754, N18736, N1325);
and AND3 (N18755, N18749, N4296, N4148);
not NOT1 (N18756, N18734);
buf BUF1 (N18757, N18737);
not NOT1 (N18758, N18753);
nor NOR2 (N18759, N18754, N5395);
and AND4 (N18760, N18752, N12950, N8803, N7857);
not NOT1 (N18761, N18758);
nor NOR4 (N18762, N18750, N4878, N5192, N6408);
or OR4 (N18763, N18759, N4410, N8367, N2339);
nand NAND4 (N18764, N18757, N10761, N6439, N2577);
nand NAND2 (N18765, N18761, N10627);
nand NAND2 (N18766, N18755, N14127);
and AND4 (N18767, N18760, N14629, N11432, N10418);
buf BUF1 (N18768, N18762);
and AND3 (N18769, N18766, N17484, N8196);
not NOT1 (N18770, N18768);
nand NAND4 (N18771, N18765, N4878, N4056, N5513);
or OR3 (N18772, N18732, N17683, N9751);
nor NOR3 (N18773, N18756, N16934, N6600);
nand NAND2 (N18774, N18767, N15101);
buf BUF1 (N18775, N18770);
xor XOR2 (N18776, N18763, N11327);
xor XOR2 (N18777, N18773, N17527);
xor XOR2 (N18778, N18771, N202);
and AND2 (N18779, N18776, N3680);
not NOT1 (N18780, N18777);
nor NOR4 (N18781, N18747, N13440, N5031, N1245);
not NOT1 (N18782, N18769);
buf BUF1 (N18783, N18774);
nor NOR3 (N18784, N18764, N4006, N2773);
xor XOR2 (N18785, N18743, N2771);
or OR4 (N18786, N18778, N8402, N4124, N14616);
and AND3 (N18787, N18786, N878, N5333);
or OR3 (N18788, N18781, N15679, N13669);
and AND4 (N18789, N18783, N4436, N18098, N4150);
not NOT1 (N18790, N18785);
or OR3 (N18791, N18790, N5916, N6993);
and AND3 (N18792, N18772, N10108, N168);
xor XOR2 (N18793, N18789, N6528);
nor NOR4 (N18794, N18787, N7347, N7145, N6536);
nand NAND2 (N18795, N18792, N9273);
nor NOR4 (N18796, N18780, N10171, N10053, N15900);
or OR4 (N18797, N18796, N17516, N8381, N9363);
and AND3 (N18798, N18794, N15667, N14646);
nand NAND2 (N18799, N18795, N12894);
nor NOR4 (N18800, N18775, N13323, N1695, N2116);
not NOT1 (N18801, N18788);
buf BUF1 (N18802, N18801);
and AND3 (N18803, N18782, N15688, N3538);
or OR4 (N18804, N18779, N8320, N6762, N7830);
xor XOR2 (N18805, N18802, N7545);
nand NAND3 (N18806, N18799, N5506, N12630);
not NOT1 (N18807, N18793);
nand NAND3 (N18808, N18803, N10499, N18801);
xor XOR2 (N18809, N18808, N15595);
or OR4 (N18810, N18800, N14922, N14867, N805);
nor NOR4 (N18811, N18784, N970, N6360, N18376);
buf BUF1 (N18812, N18809);
not NOT1 (N18813, N18812);
buf BUF1 (N18814, N18807);
nand NAND2 (N18815, N18810, N389);
and AND3 (N18816, N18804, N3435, N17708);
not NOT1 (N18817, N18798);
nor NOR2 (N18818, N18815, N1248);
and AND2 (N18819, N18811, N2932);
buf BUF1 (N18820, N18813);
nand NAND2 (N18821, N18820, N6148);
nor NOR4 (N18822, N18805, N14007, N1987, N18569);
buf BUF1 (N18823, N18817);
or OR3 (N18824, N18822, N7677, N13210);
nor NOR4 (N18825, N18821, N8278, N5530, N11984);
and AND4 (N18826, N18818, N879, N536, N3786);
not NOT1 (N18827, N18797);
or OR3 (N18828, N18816, N14684, N14314);
not NOT1 (N18829, N18825);
nor NOR3 (N18830, N18806, N16164, N15972);
xor XOR2 (N18831, N18823, N17842);
and AND4 (N18832, N18827, N5822, N10190, N10492);
xor XOR2 (N18833, N18791, N17531);
xor XOR2 (N18834, N18830, N2992);
buf BUF1 (N18835, N18826);
buf BUF1 (N18836, N18832);
xor XOR2 (N18837, N18819, N1539);
or OR2 (N18838, N18837, N7131);
or OR2 (N18839, N18836, N11851);
nor NOR3 (N18840, N18828, N10256, N1356);
buf BUF1 (N18841, N18829);
xor XOR2 (N18842, N18839, N15680);
xor XOR2 (N18843, N18814, N956);
not NOT1 (N18844, N18824);
and AND4 (N18845, N18833, N5111, N8747, N1518);
or OR4 (N18846, N18845, N15388, N15602, N16614);
xor XOR2 (N18847, N18842, N9930);
not NOT1 (N18848, N18831);
buf BUF1 (N18849, N18834);
not NOT1 (N18850, N18848);
and AND2 (N18851, N18841, N15173);
or OR2 (N18852, N18847, N9124);
nand NAND3 (N18853, N18844, N3824, N3850);
not NOT1 (N18854, N18838);
or OR4 (N18855, N18849, N18470, N16848, N5694);
buf BUF1 (N18856, N18855);
or OR3 (N18857, N18853, N2947, N16018);
nor NOR2 (N18858, N18857, N6260);
xor XOR2 (N18859, N18851, N13564);
xor XOR2 (N18860, N18856, N1198);
or OR4 (N18861, N18850, N11323, N11368, N6932);
nor NOR2 (N18862, N18861, N5013);
and AND4 (N18863, N18840, N4757, N7456, N12032);
nor NOR3 (N18864, N18852, N17913, N4259);
xor XOR2 (N18865, N18862, N2396);
not NOT1 (N18866, N18854);
xor XOR2 (N18867, N18846, N15246);
or OR3 (N18868, N18865, N11062, N11906);
xor XOR2 (N18869, N18867, N10500);
buf BUF1 (N18870, N18868);
nor NOR2 (N18871, N18864, N18441);
nor NOR2 (N18872, N18869, N7113);
not NOT1 (N18873, N18866);
not NOT1 (N18874, N18843);
nor NOR3 (N18875, N18870, N13332, N1528);
xor XOR2 (N18876, N18835, N12415);
and AND2 (N18877, N18871, N13838);
buf BUF1 (N18878, N18875);
nor NOR4 (N18879, N18863, N16164, N11532, N10049);
and AND3 (N18880, N18878, N302, N6996);
nor NOR4 (N18881, N18879, N8491, N13542, N2826);
xor XOR2 (N18882, N18880, N3027);
not NOT1 (N18883, N18881);
xor XOR2 (N18884, N18883, N18858);
xor XOR2 (N18885, N18385, N16854);
nand NAND4 (N18886, N18859, N13595, N6101, N6776);
xor XOR2 (N18887, N18882, N8489);
or OR2 (N18888, N18885, N15760);
xor XOR2 (N18889, N18884, N14379);
nor NOR3 (N18890, N18873, N5068, N4922);
buf BUF1 (N18891, N18874);
buf BUF1 (N18892, N18890);
buf BUF1 (N18893, N18892);
buf BUF1 (N18894, N18886);
buf BUF1 (N18895, N18891);
xor XOR2 (N18896, N18860, N11494);
not NOT1 (N18897, N18896);
or OR3 (N18898, N18876, N17883, N2507);
nor NOR2 (N18899, N18895, N7406);
nor NOR2 (N18900, N18887, N1507);
or OR4 (N18901, N18900, N8456, N15367, N6574);
buf BUF1 (N18902, N18872);
nor NOR3 (N18903, N18894, N55, N18400);
xor XOR2 (N18904, N18889, N12271);
buf BUF1 (N18905, N18904);
xor XOR2 (N18906, N18898, N18551);
xor XOR2 (N18907, N18897, N13898);
buf BUF1 (N18908, N18906);
nor NOR3 (N18909, N18888, N15695, N8570);
nor NOR2 (N18910, N18908, N8452);
nand NAND3 (N18911, N18893, N7082, N15808);
or OR3 (N18912, N18910, N1026, N11151);
nor NOR4 (N18913, N18899, N5110, N13483, N9513);
buf BUF1 (N18914, N18901);
buf BUF1 (N18915, N18914);
nor NOR2 (N18916, N18907, N3528);
or OR3 (N18917, N18909, N7835, N12729);
or OR2 (N18918, N18916, N6119);
nand NAND2 (N18919, N18915, N15175);
nand NAND3 (N18920, N18918, N1736, N10368);
not NOT1 (N18921, N18911);
buf BUF1 (N18922, N18912);
nand NAND3 (N18923, N18920, N11327, N13187);
nor NOR4 (N18924, N18919, N7460, N13155, N12023);
nand NAND3 (N18925, N18917, N12417, N1529);
nor NOR2 (N18926, N18913, N17248);
not NOT1 (N18927, N18924);
and AND2 (N18928, N18927, N15896);
or OR4 (N18929, N18928, N7731, N4002, N16788);
buf BUF1 (N18930, N18929);
xor XOR2 (N18931, N18930, N6318);
and AND4 (N18932, N18902, N10877, N16741, N5995);
xor XOR2 (N18933, N18925, N15339);
not NOT1 (N18934, N18931);
and AND4 (N18935, N18923, N18387, N1021, N7498);
nor NOR2 (N18936, N18926, N10052);
nand NAND4 (N18937, N18935, N17112, N6856, N8300);
xor XOR2 (N18938, N18905, N1826);
nor NOR3 (N18939, N18903, N36, N8014);
xor XOR2 (N18940, N18932, N544);
and AND4 (N18941, N18934, N15019, N9958, N3923);
xor XOR2 (N18942, N18938, N11213);
not NOT1 (N18943, N18933);
buf BUF1 (N18944, N18941);
xor XOR2 (N18945, N18944, N9209);
or OR4 (N18946, N18921, N1178, N7963, N11813);
nor NOR3 (N18947, N18936, N4998, N2398);
xor XOR2 (N18948, N18943, N10153);
nor NOR2 (N18949, N18947, N13264);
or OR2 (N18950, N18922, N9571);
nand NAND3 (N18951, N18946, N17412, N17076);
xor XOR2 (N18952, N18940, N8433);
or OR2 (N18953, N18937, N7311);
not NOT1 (N18954, N18953);
nor NOR2 (N18955, N18954, N4531);
buf BUF1 (N18956, N18955);
not NOT1 (N18957, N18956);
and AND2 (N18958, N18957, N18361);
nand NAND3 (N18959, N18942, N5971, N7466);
and AND2 (N18960, N18939, N6221);
and AND3 (N18961, N18877, N13711, N17179);
not NOT1 (N18962, N18949);
and AND3 (N18963, N18959, N18497, N14515);
nor NOR2 (N18964, N18945, N8755);
or OR2 (N18965, N18962, N11812);
nand NAND4 (N18966, N18961, N4240, N222, N6875);
nor NOR4 (N18967, N18965, N1666, N4616, N4663);
not NOT1 (N18968, N18948);
buf BUF1 (N18969, N18951);
and AND2 (N18970, N18960, N751);
or OR2 (N18971, N18968, N7067);
not NOT1 (N18972, N18970);
buf BUF1 (N18973, N18967);
nand NAND4 (N18974, N18966, N10257, N7153, N1439);
buf BUF1 (N18975, N18972);
xor XOR2 (N18976, N18952, N4582);
not NOT1 (N18977, N18958);
nand NAND2 (N18978, N18971, N18871);
xor XOR2 (N18979, N18977, N2014);
xor XOR2 (N18980, N18976, N7344);
and AND2 (N18981, N18975, N10782);
not NOT1 (N18982, N18978);
or OR3 (N18983, N18981, N16821, N4227);
nor NOR2 (N18984, N18983, N17340);
nand NAND3 (N18985, N18950, N8216, N12178);
not NOT1 (N18986, N18979);
nor NOR4 (N18987, N18985, N14966, N14112, N9975);
not NOT1 (N18988, N18980);
or OR4 (N18989, N18988, N11974, N4709, N18492);
nor NOR3 (N18990, N18989, N4573, N2016);
nor NOR2 (N18991, N18969, N816);
xor XOR2 (N18992, N18964, N15317);
nor NOR3 (N18993, N18986, N9881, N18312);
or OR3 (N18994, N18974, N5053, N11236);
not NOT1 (N18995, N18973);
nor NOR2 (N18996, N18984, N18537);
nand NAND3 (N18997, N18994, N12589, N3420);
nand NAND4 (N18998, N18991, N13630, N848, N14617);
nand NAND3 (N18999, N18995, N1966, N1557);
nand NAND2 (N19000, N18999, N21);
nor NOR4 (N19001, N18998, N3342, N6344, N4626);
nor NOR3 (N19002, N18982, N14766, N11061);
or OR4 (N19003, N18993, N14811, N3065, N17867);
nand NAND4 (N19004, N18990, N10810, N15748, N9071);
not NOT1 (N19005, N18992);
or OR4 (N19006, N19004, N7724, N16677, N7412);
and AND3 (N19007, N19005, N14307, N12596);
and AND2 (N19008, N18963, N5772);
nor NOR4 (N19009, N19003, N15495, N16881, N5894);
nor NOR4 (N19010, N19008, N2514, N2450, N654);
not NOT1 (N19011, N19001);
and AND2 (N19012, N19011, N13867);
and AND4 (N19013, N19010, N1426, N8612, N6216);
nor NOR4 (N19014, N19007, N18662, N3428, N17151);
nor NOR3 (N19015, N19000, N11115, N14607);
nand NAND3 (N19016, N19006, N11586, N11381);
and AND2 (N19017, N19016, N13772);
or OR4 (N19018, N18987, N7274, N1338, N13880);
nand NAND4 (N19019, N19014, N16491, N1546, N4161);
nor NOR2 (N19020, N19012, N3559);
nor NOR4 (N19021, N19018, N10407, N6984, N3504);
xor XOR2 (N19022, N19021, N13380);
or OR3 (N19023, N18996, N12191, N15010);
nand NAND4 (N19024, N18997, N13307, N6939, N2240);
or OR4 (N19025, N19024, N10979, N16215, N13873);
buf BUF1 (N19026, N19002);
xor XOR2 (N19027, N19022, N15625);
or OR4 (N19028, N19017, N12383, N85, N16093);
nand NAND4 (N19029, N19009, N7259, N17521, N15096);
nand NAND2 (N19030, N19029, N6599);
and AND3 (N19031, N19026, N12561, N18709);
or OR2 (N19032, N19027, N15707);
or OR3 (N19033, N19019, N8, N15821);
not NOT1 (N19034, N19015);
buf BUF1 (N19035, N19033);
nor NOR3 (N19036, N19035, N12279, N7712);
and AND3 (N19037, N19023, N3733, N2234);
or OR4 (N19038, N19031, N10370, N17887, N1257);
buf BUF1 (N19039, N19036);
not NOT1 (N19040, N19013);
or OR3 (N19041, N19030, N6580, N1175);
not NOT1 (N19042, N19041);
nor NOR4 (N19043, N19032, N9687, N10501, N10097);
nand NAND2 (N19044, N19020, N262);
not NOT1 (N19045, N19037);
xor XOR2 (N19046, N19039, N3146);
nor NOR2 (N19047, N19046, N14205);
not NOT1 (N19048, N19040);
or OR4 (N19049, N19042, N17274, N14361, N18737);
buf BUF1 (N19050, N19049);
not NOT1 (N19051, N19028);
nor NOR4 (N19052, N19045, N15888, N15915, N13880);
buf BUF1 (N19053, N19043);
nor NOR3 (N19054, N19051, N14457, N6522);
buf BUF1 (N19055, N19052);
or OR2 (N19056, N19038, N18540);
nor NOR4 (N19057, N19044, N18149, N7893, N3721);
buf BUF1 (N19058, N19055);
not NOT1 (N19059, N19056);
nand NAND3 (N19060, N19047, N18923, N4013);
and AND3 (N19061, N19058, N5411, N2241);
nor NOR3 (N19062, N19034, N14818, N767);
not NOT1 (N19063, N19054);
and AND3 (N19064, N19063, N11755, N10991);
or OR3 (N19065, N19061, N18770, N8029);
buf BUF1 (N19066, N19060);
nor NOR3 (N19067, N19025, N14131, N18132);
and AND4 (N19068, N19057, N10207, N9759, N15906);
or OR3 (N19069, N19064, N13141, N1403);
not NOT1 (N19070, N19050);
xor XOR2 (N19071, N19059, N6900);
buf BUF1 (N19072, N19048);
or OR3 (N19073, N19070, N8071, N5955);
buf BUF1 (N19074, N19067);
xor XOR2 (N19075, N19074, N11534);
not NOT1 (N19076, N19065);
or OR3 (N19077, N19068, N1165, N6993);
xor XOR2 (N19078, N19053, N11555);
and AND4 (N19079, N19076, N16370, N4861, N1315);
nor NOR3 (N19080, N19073, N12020, N1401);
or OR3 (N19081, N19062, N4417, N4119);
and AND3 (N19082, N19080, N11857, N16133);
or OR4 (N19083, N19066, N3467, N14110, N320);
nor NOR2 (N19084, N19069, N12274);
xor XOR2 (N19085, N19075, N2589);
not NOT1 (N19086, N19071);
or OR2 (N19087, N19077, N10542);
nand NAND2 (N19088, N19083, N10513);
not NOT1 (N19089, N19078);
buf BUF1 (N19090, N19089);
nand NAND2 (N19091, N19082, N17950);
buf BUF1 (N19092, N19079);
nand NAND4 (N19093, N19086, N17373, N3028, N3656);
xor XOR2 (N19094, N19084, N2103);
or OR3 (N19095, N19090, N16887, N12710);
and AND2 (N19096, N19094, N6176);
buf BUF1 (N19097, N19081);
and AND3 (N19098, N19087, N5060, N13445);
nor NOR3 (N19099, N19096, N6838, N13090);
and AND3 (N19100, N19098, N467, N11411);
and AND2 (N19101, N19093, N16358);
and AND3 (N19102, N19088, N18875, N17908);
or OR4 (N19103, N19097, N9358, N18655, N17784);
and AND3 (N19104, N19095, N16103, N10553);
nor NOR3 (N19105, N19103, N13054, N2109);
nand NAND4 (N19106, N19100, N11275, N2774, N14456);
or OR2 (N19107, N19099, N7392);
xor XOR2 (N19108, N19104, N9877);
nor NOR3 (N19109, N19105, N17602, N11027);
and AND3 (N19110, N19109, N13842, N2213);
nor NOR4 (N19111, N19092, N17864, N9289, N17913);
and AND2 (N19112, N19102, N6902);
nand NAND3 (N19113, N19085, N1780, N17157);
nor NOR4 (N19114, N19091, N476, N7430, N16873);
nor NOR4 (N19115, N19111, N19006, N7249, N6664);
not NOT1 (N19116, N19072);
xor XOR2 (N19117, N19112, N9676);
not NOT1 (N19118, N19114);
xor XOR2 (N19119, N19113, N6914);
nand NAND4 (N19120, N19117, N18949, N8166, N18360);
or OR2 (N19121, N19119, N619);
and AND4 (N19122, N19110, N13753, N10702, N4234);
nor NOR4 (N19123, N19121, N8492, N16138, N14185);
and AND2 (N19124, N19118, N15185);
xor XOR2 (N19125, N19124, N15515);
and AND2 (N19126, N19106, N16959);
not NOT1 (N19127, N19108);
not NOT1 (N19128, N19101);
or OR4 (N19129, N19116, N11163, N9651, N15268);
nor NOR4 (N19130, N19123, N2646, N16197, N18127);
buf BUF1 (N19131, N19122);
or OR2 (N19132, N19125, N3696);
buf BUF1 (N19133, N19115);
xor XOR2 (N19134, N19133, N16574);
nand NAND3 (N19135, N19131, N19065, N4102);
xor XOR2 (N19136, N19132, N1160);
or OR3 (N19137, N19130, N2200, N1064);
and AND3 (N19138, N19137, N1962, N7695);
xor XOR2 (N19139, N19126, N7027);
nor NOR2 (N19140, N19129, N5709);
nand NAND2 (N19141, N19128, N2713);
buf BUF1 (N19142, N19134);
nor NOR2 (N19143, N19142, N2341);
and AND3 (N19144, N19138, N2234, N11140);
or OR2 (N19145, N19144, N2927);
buf BUF1 (N19146, N19143);
nor NOR2 (N19147, N19139, N1899);
buf BUF1 (N19148, N19135);
nor NOR4 (N19149, N19140, N9489, N6397, N5142);
not NOT1 (N19150, N19145);
not NOT1 (N19151, N19127);
nand NAND4 (N19152, N19146, N4715, N364, N7968);
or OR4 (N19153, N19107, N16679, N6073, N17691);
not NOT1 (N19154, N19136);
xor XOR2 (N19155, N19147, N4176);
or OR4 (N19156, N19120, N4835, N4920, N10895);
nor NOR2 (N19157, N19152, N18103);
and AND2 (N19158, N19154, N15448);
and AND3 (N19159, N19151, N15393, N6180);
xor XOR2 (N19160, N19148, N8640);
or OR4 (N19161, N19157, N18688, N6424, N4249);
and AND3 (N19162, N19149, N4608, N13576);
xor XOR2 (N19163, N19141, N13579);
and AND2 (N19164, N19158, N764);
and AND3 (N19165, N19163, N13825, N12937);
nand NAND4 (N19166, N19156, N13290, N10856, N6738);
not NOT1 (N19167, N19150);
nand NAND2 (N19168, N19164, N8063);
nor NOR4 (N19169, N19155, N1301, N11653, N2356);
or OR4 (N19170, N19161, N3531, N6267, N3959);
buf BUF1 (N19171, N19165);
nor NOR3 (N19172, N19167, N14022, N12489);
and AND3 (N19173, N19153, N18881, N180);
or OR4 (N19174, N19170, N7860, N15172, N17203);
nand NAND2 (N19175, N19169, N11151);
xor XOR2 (N19176, N19159, N8193);
and AND3 (N19177, N19166, N9062, N15078);
xor XOR2 (N19178, N19162, N10313);
nand NAND2 (N19179, N19175, N7262);
or OR3 (N19180, N19171, N16180, N18691);
nor NOR3 (N19181, N19176, N4389, N6245);
and AND3 (N19182, N19180, N6076, N6192);
xor XOR2 (N19183, N19181, N14906);
xor XOR2 (N19184, N19172, N3496);
not NOT1 (N19185, N19184);
not NOT1 (N19186, N19168);
xor XOR2 (N19187, N19173, N11535);
xor XOR2 (N19188, N19186, N2234);
xor XOR2 (N19189, N19185, N2382);
nor NOR4 (N19190, N19179, N15794, N6901, N15166);
or OR2 (N19191, N19188, N4568);
xor XOR2 (N19192, N19160, N14496);
buf BUF1 (N19193, N19174);
not NOT1 (N19194, N19182);
and AND4 (N19195, N19193, N17299, N706, N14637);
and AND2 (N19196, N19192, N13178);
xor XOR2 (N19197, N19194, N3593);
not NOT1 (N19198, N19177);
and AND3 (N19199, N19187, N12764, N5749);
buf BUF1 (N19200, N19191);
not NOT1 (N19201, N19199);
not NOT1 (N19202, N19195);
nor NOR3 (N19203, N19197, N10990, N17585);
and AND2 (N19204, N19200, N8659);
xor XOR2 (N19205, N19190, N7397);
nor NOR2 (N19206, N19203, N13836);
xor XOR2 (N19207, N19201, N6135);
not NOT1 (N19208, N19207);
and AND2 (N19209, N19205, N870);
not NOT1 (N19210, N19204);
not NOT1 (N19211, N19178);
nand NAND2 (N19212, N19189, N2360);
xor XOR2 (N19213, N19209, N5123);
and AND3 (N19214, N19196, N15936, N6702);
nand NAND2 (N19215, N19202, N2316);
buf BUF1 (N19216, N19211);
or OR4 (N19217, N19206, N5868, N17019, N18543);
nand NAND4 (N19218, N19214, N16948, N11952, N8033);
and AND2 (N19219, N19216, N899);
xor XOR2 (N19220, N19210, N17919);
xor XOR2 (N19221, N19213, N3358);
and AND3 (N19222, N19219, N12284, N341);
xor XOR2 (N19223, N19208, N578);
nor NOR3 (N19224, N19222, N14589, N4961);
buf BUF1 (N19225, N19183);
nand NAND3 (N19226, N19224, N4596, N17501);
xor XOR2 (N19227, N19217, N5610);
not NOT1 (N19228, N19218);
xor XOR2 (N19229, N19212, N5324);
or OR3 (N19230, N19223, N18122, N9944);
nor NOR4 (N19231, N19198, N5027, N14164, N235);
and AND2 (N19232, N19220, N16627);
xor XOR2 (N19233, N19226, N8795);
nand NAND3 (N19234, N19229, N12307, N5303);
or OR2 (N19235, N19221, N2942);
xor XOR2 (N19236, N19233, N16107);
not NOT1 (N19237, N19228);
and AND2 (N19238, N19237, N5744);
and AND3 (N19239, N19236, N14094, N13949);
nand NAND3 (N19240, N19225, N15956, N1926);
buf BUF1 (N19241, N19215);
buf BUF1 (N19242, N19230);
not NOT1 (N19243, N19238);
xor XOR2 (N19244, N19235, N6823);
and AND3 (N19245, N19240, N17518, N1638);
nor NOR2 (N19246, N19239, N1049);
and AND4 (N19247, N19227, N4114, N12017, N15141);
and AND2 (N19248, N19231, N10475);
or OR2 (N19249, N19246, N7456);
buf BUF1 (N19250, N19234);
nand NAND2 (N19251, N19244, N2585);
buf BUF1 (N19252, N19250);
nor NOR2 (N19253, N19241, N2746);
nand NAND3 (N19254, N19243, N3270, N3084);
or OR4 (N19255, N19232, N13976, N16404, N5525);
and AND3 (N19256, N19248, N6039, N5311);
buf BUF1 (N19257, N19255);
not NOT1 (N19258, N19242);
xor XOR2 (N19259, N19258, N5545);
or OR2 (N19260, N19253, N1641);
nor NOR4 (N19261, N19247, N1636, N15950, N4548);
and AND4 (N19262, N19245, N16130, N11229, N11728);
nand NAND4 (N19263, N19259, N2543, N15298, N12658);
nor NOR4 (N19264, N19252, N12015, N15934, N6707);
nor NOR2 (N19265, N19257, N8641);
nor NOR3 (N19266, N19265, N981, N8163);
buf BUF1 (N19267, N19256);
not NOT1 (N19268, N19266);
xor XOR2 (N19269, N19261, N3140);
nand NAND2 (N19270, N19254, N4387);
and AND3 (N19271, N19264, N1334, N2567);
and AND2 (N19272, N19270, N4127);
nand NAND3 (N19273, N19262, N12540, N2065);
nand NAND4 (N19274, N19249, N17492, N16712, N12657);
or OR2 (N19275, N19263, N16689);
not NOT1 (N19276, N19267);
and AND4 (N19277, N19275, N5299, N16215, N10862);
and AND2 (N19278, N19273, N11828);
or OR4 (N19279, N19272, N15538, N5250, N17970);
buf BUF1 (N19280, N19268);
and AND2 (N19281, N19274, N14556);
buf BUF1 (N19282, N19281);
or OR3 (N19283, N19276, N3681, N9590);
xor XOR2 (N19284, N19282, N3851);
xor XOR2 (N19285, N19279, N9723);
not NOT1 (N19286, N19278);
or OR2 (N19287, N19286, N6788);
nor NOR3 (N19288, N19277, N16555, N1262);
nand NAND3 (N19289, N19271, N3739, N1366);
nor NOR3 (N19290, N19269, N16680, N11599);
or OR3 (N19291, N19284, N3092, N830);
nor NOR2 (N19292, N19283, N9502);
or OR4 (N19293, N19251, N14265, N10247, N2298);
nor NOR4 (N19294, N19290, N15163, N11384, N8704);
buf BUF1 (N19295, N19292);
and AND3 (N19296, N19289, N6347, N16033);
nor NOR4 (N19297, N19293, N18178, N14464, N15361);
nand NAND2 (N19298, N19295, N2168);
buf BUF1 (N19299, N19285);
buf BUF1 (N19300, N19298);
nand NAND3 (N19301, N19299, N8349, N6684);
nand NAND4 (N19302, N19300, N5184, N14347, N9607);
nor NOR4 (N19303, N19302, N12122, N17099, N4949);
buf BUF1 (N19304, N19294);
nor NOR2 (N19305, N19301, N12959);
nand NAND2 (N19306, N19304, N16925);
not NOT1 (N19307, N19287);
nand NAND3 (N19308, N19296, N14056, N7236);
nand NAND3 (N19309, N19260, N17001, N8942);
buf BUF1 (N19310, N19291);
or OR4 (N19311, N19306, N8912, N6327, N17608);
or OR4 (N19312, N19280, N5332, N4834, N8808);
and AND3 (N19313, N19288, N15319, N12371);
not NOT1 (N19314, N19311);
xor XOR2 (N19315, N19312, N8567);
and AND2 (N19316, N19309, N4109);
nor NOR4 (N19317, N19316, N5384, N243, N12986);
xor XOR2 (N19318, N19313, N12210);
and AND3 (N19319, N19308, N2145, N13766);
nor NOR4 (N19320, N19319, N10460, N3971, N9222);
xor XOR2 (N19321, N19315, N7996);
and AND4 (N19322, N19307, N17274, N16274, N13612);
nor NOR2 (N19323, N19314, N16965);
nand NAND3 (N19324, N19320, N14565, N5695);
buf BUF1 (N19325, N19317);
nor NOR4 (N19326, N19318, N1977, N8477, N15382);
nor NOR3 (N19327, N19303, N18957, N12488);
not NOT1 (N19328, N19321);
nor NOR3 (N19329, N19297, N10000, N14334);
or OR2 (N19330, N19324, N13527);
nand NAND3 (N19331, N19325, N10802, N15210);
buf BUF1 (N19332, N19323);
not NOT1 (N19333, N19326);
or OR2 (N19334, N19329, N5555);
nand NAND2 (N19335, N19305, N15020);
nor NOR4 (N19336, N19328, N15377, N14061, N544);
nor NOR2 (N19337, N19330, N15255);
and AND4 (N19338, N19327, N11554, N6608, N2026);
and AND2 (N19339, N19331, N4305);
or OR4 (N19340, N19334, N3216, N4156, N15340);
xor XOR2 (N19341, N19332, N11513);
buf BUF1 (N19342, N19338);
nand NAND3 (N19343, N19333, N13929, N4481);
not NOT1 (N19344, N19322);
xor XOR2 (N19345, N19340, N4508);
buf BUF1 (N19346, N19336);
buf BUF1 (N19347, N19337);
nor NOR4 (N19348, N19344, N18657, N9879, N8383);
buf BUF1 (N19349, N19345);
and AND3 (N19350, N19346, N4670, N8811);
nor NOR2 (N19351, N19348, N9373);
nor NOR2 (N19352, N19339, N15069);
buf BUF1 (N19353, N19352);
not NOT1 (N19354, N19351);
nor NOR2 (N19355, N19353, N16200);
nor NOR4 (N19356, N19342, N7716, N833, N941);
not NOT1 (N19357, N19356);
nand NAND4 (N19358, N19335, N17649, N6628, N12268);
xor XOR2 (N19359, N19310, N9423);
buf BUF1 (N19360, N19355);
xor XOR2 (N19361, N19358, N17630);
buf BUF1 (N19362, N19361);
nor NOR4 (N19363, N19359, N16210, N15945, N4141);
and AND2 (N19364, N19360, N18411);
buf BUF1 (N19365, N19357);
or OR2 (N19366, N19350, N9869);
not NOT1 (N19367, N19349);
nand NAND4 (N19368, N19365, N13600, N941, N1366);
buf BUF1 (N19369, N19364);
or OR3 (N19370, N19354, N6086, N7345);
or OR3 (N19371, N19363, N9914, N1555);
nor NOR2 (N19372, N19347, N14400);
not NOT1 (N19373, N19367);
not NOT1 (N19374, N19341);
nand NAND2 (N19375, N19372, N18625);
xor XOR2 (N19376, N19368, N6149);
nor NOR2 (N19377, N19370, N18066);
buf BUF1 (N19378, N19371);
not NOT1 (N19379, N19362);
nor NOR3 (N19380, N19379, N7044, N14215);
not NOT1 (N19381, N19373);
xor XOR2 (N19382, N19378, N16923);
nand NAND3 (N19383, N19375, N19067, N1066);
nand NAND2 (N19384, N19377, N17201);
or OR2 (N19385, N19376, N16587);
and AND2 (N19386, N19366, N15826);
nand NAND3 (N19387, N19343, N5029, N18782);
nand NAND3 (N19388, N19374, N17815, N11343);
and AND2 (N19389, N19386, N13755);
buf BUF1 (N19390, N19387);
nand NAND3 (N19391, N19383, N6023, N18031);
not NOT1 (N19392, N19384);
or OR2 (N19393, N19389, N1788);
not NOT1 (N19394, N19381);
or OR3 (N19395, N19392, N7311, N8362);
xor XOR2 (N19396, N19391, N14532);
or OR4 (N19397, N19390, N16562, N667, N12971);
buf BUF1 (N19398, N19380);
and AND2 (N19399, N19394, N4260);
buf BUF1 (N19400, N19397);
buf BUF1 (N19401, N19398);
and AND4 (N19402, N19369, N13241, N838, N15651);
buf BUF1 (N19403, N19401);
not NOT1 (N19404, N19396);
or OR4 (N19405, N19395, N12045, N15758, N12720);
xor XOR2 (N19406, N19393, N6255);
nand NAND3 (N19407, N19382, N1249, N4645);
and AND4 (N19408, N19402, N11961, N18898, N2335);
or OR3 (N19409, N19408, N17102, N6553);
or OR3 (N19410, N19404, N17458, N4342);
nand NAND2 (N19411, N19406, N8633);
buf BUF1 (N19412, N19400);
not NOT1 (N19413, N19399);
nor NOR2 (N19414, N19407, N16861);
nor NOR4 (N19415, N19413, N5642, N7748, N14414);
xor XOR2 (N19416, N19403, N3691);
xor XOR2 (N19417, N19409, N1899);
buf BUF1 (N19418, N19415);
xor XOR2 (N19419, N19411, N16516);
or OR2 (N19420, N19419, N17384);
nand NAND2 (N19421, N19417, N13030);
or OR3 (N19422, N19420, N6419, N11132);
buf BUF1 (N19423, N19412);
nor NOR2 (N19424, N19388, N1381);
buf BUF1 (N19425, N19410);
nand NAND2 (N19426, N19385, N4640);
xor XOR2 (N19427, N19421, N6197);
xor XOR2 (N19428, N19422, N11242);
nor NOR3 (N19429, N19414, N5918, N17996);
or OR2 (N19430, N19423, N19130);
not NOT1 (N19431, N19424);
nand NAND3 (N19432, N19430, N13718, N4192);
buf BUF1 (N19433, N19416);
not NOT1 (N19434, N19426);
and AND2 (N19435, N19425, N16717);
nand NAND4 (N19436, N19435, N850, N7648, N6119);
or OR4 (N19437, N19431, N15268, N12181, N4817);
or OR2 (N19438, N19428, N11525);
nor NOR4 (N19439, N19432, N18616, N6369, N1708);
buf BUF1 (N19440, N19433);
or OR2 (N19441, N19436, N431);
nand NAND4 (N19442, N19405, N6562, N16268, N17154);
not NOT1 (N19443, N19440);
buf BUF1 (N19444, N19418);
xor XOR2 (N19445, N19438, N188);
nor NOR3 (N19446, N19442, N4206, N4032);
not NOT1 (N19447, N19427);
xor XOR2 (N19448, N19429, N13190);
buf BUF1 (N19449, N19446);
or OR2 (N19450, N19443, N8042);
nor NOR2 (N19451, N19445, N12500);
or OR2 (N19452, N19448, N5741);
buf BUF1 (N19453, N19439);
xor XOR2 (N19454, N19441, N1715);
not NOT1 (N19455, N19454);
and AND3 (N19456, N19437, N11319, N3663);
or OR4 (N19457, N19450, N7786, N11241, N6801);
nand NAND4 (N19458, N19449, N17581, N2961, N10611);
not NOT1 (N19459, N19451);
or OR2 (N19460, N19455, N18297);
nand NAND4 (N19461, N19453, N12421, N9715, N2705);
xor XOR2 (N19462, N19461, N16935);
buf BUF1 (N19463, N19447);
nor NOR3 (N19464, N19459, N4507, N7998);
nand NAND4 (N19465, N19452, N101, N11610, N18333);
and AND2 (N19466, N19434, N7646);
buf BUF1 (N19467, N19464);
xor XOR2 (N19468, N19462, N14212);
nand NAND4 (N19469, N19467, N3000, N15234, N18815);
or OR3 (N19470, N19468, N19274, N13021);
not NOT1 (N19471, N19457);
buf BUF1 (N19472, N19471);
or OR3 (N19473, N19469, N12351, N543);
and AND3 (N19474, N19458, N9513, N14979);
buf BUF1 (N19475, N19444);
buf BUF1 (N19476, N19463);
nor NOR2 (N19477, N19465, N4220);
not NOT1 (N19478, N19473);
buf BUF1 (N19479, N19477);
buf BUF1 (N19480, N19478);
and AND4 (N19481, N19466, N5622, N16949, N7199);
or OR2 (N19482, N19480, N2605);
xor XOR2 (N19483, N19475, N9675);
not NOT1 (N19484, N19476);
buf BUF1 (N19485, N19483);
nand NAND3 (N19486, N19482, N12379, N12538);
not NOT1 (N19487, N19460);
xor XOR2 (N19488, N19479, N12988);
nor NOR3 (N19489, N19470, N4215, N16352);
and AND2 (N19490, N19486, N18751);
buf BUF1 (N19491, N19488);
nor NOR2 (N19492, N19485, N5701);
and AND4 (N19493, N19492, N2221, N18319, N19168);
xor XOR2 (N19494, N19490, N9397);
and AND2 (N19495, N19484, N14877);
buf BUF1 (N19496, N19472);
xor XOR2 (N19497, N19493, N2925);
not NOT1 (N19498, N19496);
buf BUF1 (N19499, N19495);
or OR2 (N19500, N19499, N11544);
nor NOR3 (N19501, N19498, N3582, N17234);
buf BUF1 (N19502, N19501);
xor XOR2 (N19503, N19502, N3501);
nor NOR3 (N19504, N19494, N16387, N11199);
or OR3 (N19505, N19497, N15094, N7216);
and AND3 (N19506, N19503, N5525, N5067);
not NOT1 (N19507, N19487);
xor XOR2 (N19508, N19500, N4130);
xor XOR2 (N19509, N19481, N9381);
and AND3 (N19510, N19508, N11237, N12134);
or OR3 (N19511, N19504, N7531, N12388);
nor NOR2 (N19512, N19506, N16867);
not NOT1 (N19513, N19474);
buf BUF1 (N19514, N19456);
nor NOR3 (N19515, N19507, N4457, N4250);
nor NOR3 (N19516, N19489, N17894, N11819);
nand NAND3 (N19517, N19509, N16032, N1122);
and AND4 (N19518, N19514, N2141, N3840, N15988);
or OR2 (N19519, N19510, N14339);
buf BUF1 (N19520, N19511);
buf BUF1 (N19521, N19512);
nand NAND2 (N19522, N19491, N5082);
nor NOR2 (N19523, N19517, N2960);
or OR2 (N19524, N19519, N4298);
and AND3 (N19525, N19521, N17743, N6009);
and AND4 (N19526, N19525, N5500, N14097, N8701);
buf BUF1 (N19527, N19513);
not NOT1 (N19528, N19526);
xor XOR2 (N19529, N19528, N10826);
and AND4 (N19530, N19520, N15622, N9445, N12664);
nand NAND3 (N19531, N19518, N2433, N3384);
nand NAND2 (N19532, N19530, N16088);
or OR4 (N19533, N19516, N15509, N3081, N8038);
xor XOR2 (N19534, N19533, N11685);
xor XOR2 (N19535, N19522, N7947);
nand NAND4 (N19536, N19515, N13932, N16234, N11931);
not NOT1 (N19537, N19535);
buf BUF1 (N19538, N19534);
buf BUF1 (N19539, N19524);
not NOT1 (N19540, N19505);
nor NOR4 (N19541, N19527, N5554, N17536, N10536);
xor XOR2 (N19542, N19540, N10656);
or OR2 (N19543, N19537, N17988);
nor NOR2 (N19544, N19538, N18198);
or OR3 (N19545, N19523, N3833, N1107);
nor NOR3 (N19546, N19539, N2568, N9385);
xor XOR2 (N19547, N19529, N11923);
nand NAND4 (N19548, N19547, N14639, N8751, N1333);
buf BUF1 (N19549, N19532);
nand NAND4 (N19550, N19543, N15979, N6309, N6941);
not NOT1 (N19551, N19536);
or OR2 (N19552, N19549, N17970);
or OR4 (N19553, N19544, N14223, N693, N4602);
buf BUF1 (N19554, N19551);
buf BUF1 (N19555, N19550);
nand NAND3 (N19556, N19542, N9190, N10904);
nand NAND3 (N19557, N19548, N1718, N15077);
and AND2 (N19558, N19557, N10925);
not NOT1 (N19559, N19541);
not NOT1 (N19560, N19531);
nor NOR3 (N19561, N19554, N19436, N850);
nand NAND3 (N19562, N19546, N5554, N6137);
or OR2 (N19563, N19552, N8487);
nor NOR3 (N19564, N19553, N8267, N12689);
or OR2 (N19565, N19563, N16288);
xor XOR2 (N19566, N19545, N4148);
and AND2 (N19567, N19561, N4792);
nor NOR3 (N19568, N19555, N18202, N12161);
not NOT1 (N19569, N19556);
not NOT1 (N19570, N19558);
buf BUF1 (N19571, N19559);
or OR2 (N19572, N19562, N1269);
nand NAND3 (N19573, N19568, N12954, N5624);
xor XOR2 (N19574, N19560, N13004);
not NOT1 (N19575, N19564);
not NOT1 (N19576, N19573);
nand NAND2 (N19577, N19565, N19503);
not NOT1 (N19578, N19576);
not NOT1 (N19579, N19572);
nand NAND3 (N19580, N19578, N12405, N18103);
xor XOR2 (N19581, N19574, N11996);
nor NOR2 (N19582, N19577, N8056);
xor XOR2 (N19583, N19575, N8339);
nand NAND3 (N19584, N19579, N12977, N11910);
buf BUF1 (N19585, N19571);
xor XOR2 (N19586, N19583, N17596);
nor NOR2 (N19587, N19570, N13753);
buf BUF1 (N19588, N19584);
and AND2 (N19589, N19569, N13870);
nand NAND4 (N19590, N19587, N14370, N16388, N14394);
nand NAND4 (N19591, N19580, N15956, N8857, N15539);
buf BUF1 (N19592, N19588);
and AND3 (N19593, N19591, N7891, N15340);
nand NAND4 (N19594, N19567, N7801, N1708, N16705);
nand NAND3 (N19595, N19585, N7100, N5108);
nor NOR4 (N19596, N19586, N2612, N17116, N5586);
or OR4 (N19597, N19593, N6798, N11094, N14656);
nor NOR2 (N19598, N19594, N6733);
and AND2 (N19599, N19596, N5289);
buf BUF1 (N19600, N19590);
nand NAND2 (N19601, N19598, N8515);
nor NOR3 (N19602, N19600, N17044, N16453);
xor XOR2 (N19603, N19582, N15838);
xor XOR2 (N19604, N19592, N4100);
and AND2 (N19605, N19602, N811);
and AND3 (N19606, N19581, N3152, N5369);
and AND3 (N19607, N19604, N12101, N18884);
and AND2 (N19608, N19597, N2678);
nor NOR2 (N19609, N19566, N19580);
xor XOR2 (N19610, N19607, N14239);
xor XOR2 (N19611, N19599, N850);
xor XOR2 (N19612, N19611, N6381);
nand NAND3 (N19613, N19612, N1514, N1374);
nor NOR4 (N19614, N19589, N398, N10752, N18759);
xor XOR2 (N19615, N19603, N3713);
nor NOR2 (N19616, N19610, N2701);
or OR4 (N19617, N19606, N19583, N10014, N16942);
nor NOR4 (N19618, N19608, N12184, N1713, N18763);
or OR2 (N19619, N19614, N6631);
xor XOR2 (N19620, N19609, N2134);
or OR4 (N19621, N19613, N11626, N207, N6790);
or OR4 (N19622, N19617, N112, N18125, N1483);
or OR2 (N19623, N19601, N8268);
nor NOR3 (N19624, N19618, N1470, N5103);
and AND4 (N19625, N19620, N16866, N12616, N1392);
and AND2 (N19626, N19595, N16966);
or OR3 (N19627, N19623, N19624, N7450);
or OR3 (N19628, N11621, N3404, N5838);
and AND4 (N19629, N19615, N5158, N3464, N2806);
nor NOR4 (N19630, N19621, N7673, N19142, N13316);
or OR4 (N19631, N19627, N2517, N13111, N1976);
or OR3 (N19632, N19605, N318, N12422);
xor XOR2 (N19633, N19625, N14719);
buf BUF1 (N19634, N19616);
not NOT1 (N19635, N19632);
nand NAND3 (N19636, N19626, N12477, N7805);
buf BUF1 (N19637, N19628);
buf BUF1 (N19638, N19636);
xor XOR2 (N19639, N19638, N4130);
nand NAND3 (N19640, N19635, N6922, N3319);
xor XOR2 (N19641, N19630, N2425);
not NOT1 (N19642, N19629);
buf BUF1 (N19643, N19633);
or OR2 (N19644, N19631, N10346);
and AND2 (N19645, N19622, N8306);
nand NAND4 (N19646, N19644, N17874, N2698, N636);
xor XOR2 (N19647, N19641, N19016);
buf BUF1 (N19648, N19637);
not NOT1 (N19649, N19619);
not NOT1 (N19650, N19647);
xor XOR2 (N19651, N19642, N7680);
or OR2 (N19652, N19639, N11667);
nor NOR2 (N19653, N19651, N7137);
xor XOR2 (N19654, N19648, N10482);
nand NAND3 (N19655, N19650, N4928, N13597);
nor NOR2 (N19656, N19652, N18747);
xor XOR2 (N19657, N19643, N11158);
xor XOR2 (N19658, N19656, N13659);
nor NOR2 (N19659, N19655, N14747);
and AND3 (N19660, N19640, N447, N4976);
and AND4 (N19661, N19653, N6872, N818, N18173);
buf BUF1 (N19662, N19658);
buf BUF1 (N19663, N19659);
nor NOR3 (N19664, N19646, N19097, N13503);
nor NOR4 (N19665, N19634, N15034, N3557, N18135);
nor NOR3 (N19666, N19663, N17528, N7165);
or OR4 (N19667, N19661, N5903, N14070, N6039);
or OR4 (N19668, N19664, N14532, N10278, N8680);
xor XOR2 (N19669, N19668, N3355);
or OR2 (N19670, N19657, N10378);
nor NOR4 (N19671, N19666, N18274, N14883, N16777);
nand NAND4 (N19672, N19649, N11946, N2913, N13875);
not NOT1 (N19673, N19671);
or OR4 (N19674, N19662, N14390, N3919, N6128);
and AND3 (N19675, N19669, N5102, N16243);
xor XOR2 (N19676, N19670, N13227);
or OR2 (N19677, N19672, N524);
nand NAND2 (N19678, N19667, N15991);
xor XOR2 (N19679, N19675, N18122);
buf BUF1 (N19680, N19674);
nand NAND4 (N19681, N19677, N18117, N2384, N6554);
buf BUF1 (N19682, N19654);
and AND2 (N19683, N19680, N15393);
nand NAND2 (N19684, N19665, N10058);
xor XOR2 (N19685, N19676, N9108);
and AND4 (N19686, N19660, N18941, N17327, N2734);
xor XOR2 (N19687, N19678, N11533);
xor XOR2 (N19688, N19679, N833);
not NOT1 (N19689, N19685);
nor NOR3 (N19690, N19687, N1038, N14247);
not NOT1 (N19691, N19681);
or OR3 (N19692, N19682, N15853, N10335);
buf BUF1 (N19693, N19690);
nand NAND3 (N19694, N19686, N10358, N15107);
nor NOR3 (N19695, N19691, N361, N4724);
nor NOR2 (N19696, N19689, N3157);
nand NAND2 (N19697, N19645, N19142);
nor NOR4 (N19698, N19688, N16581, N15543, N14086);
buf BUF1 (N19699, N19696);
buf BUF1 (N19700, N19695);
and AND3 (N19701, N19699, N7066, N9977);
and AND2 (N19702, N19697, N9721);
buf BUF1 (N19703, N19692);
not NOT1 (N19704, N19703);
and AND2 (N19705, N19701, N19026);
nor NOR2 (N19706, N19702, N14989);
xor XOR2 (N19707, N19673, N15155);
xor XOR2 (N19708, N19704, N1629);
nor NOR2 (N19709, N19708, N4028);
buf BUF1 (N19710, N19698);
and AND4 (N19711, N19705, N14040, N14949, N14907);
or OR2 (N19712, N19700, N17068);
and AND4 (N19713, N19683, N2544, N8346, N19398);
or OR3 (N19714, N19709, N15499, N16440);
buf BUF1 (N19715, N19706);
buf BUF1 (N19716, N19707);
nand NAND2 (N19717, N19714, N7974);
not NOT1 (N19718, N19710);
not NOT1 (N19719, N19711);
buf BUF1 (N19720, N19684);
nor NOR3 (N19721, N19720, N9484, N11347);
and AND3 (N19722, N19717, N1313, N14376);
buf BUF1 (N19723, N19693);
or OR3 (N19724, N19712, N7496, N900);
xor XOR2 (N19725, N19721, N8780);
buf BUF1 (N19726, N19722);
not NOT1 (N19727, N19724);
nand NAND3 (N19728, N19726, N10430, N1220);
nor NOR2 (N19729, N19715, N15379);
nand NAND2 (N19730, N19718, N16090);
nand NAND4 (N19731, N19727, N3217, N3479, N508);
nor NOR4 (N19732, N19728, N10877, N13949, N15027);
and AND3 (N19733, N19730, N14762, N19053);
nor NOR4 (N19734, N19733, N8236, N9123, N11128);
buf BUF1 (N19735, N19734);
xor XOR2 (N19736, N19694, N10874);
or OR2 (N19737, N19723, N15410);
xor XOR2 (N19738, N19732, N6770);
not NOT1 (N19739, N19716);
not NOT1 (N19740, N19719);
xor XOR2 (N19741, N19735, N2961);
and AND3 (N19742, N19738, N6634, N18121);
not NOT1 (N19743, N19736);
not NOT1 (N19744, N19737);
buf BUF1 (N19745, N19744);
xor XOR2 (N19746, N19742, N18908);
nor NOR3 (N19747, N19725, N4575, N16320);
not NOT1 (N19748, N19740);
or OR2 (N19749, N19739, N12215);
and AND2 (N19750, N19741, N17106);
and AND2 (N19751, N19750, N14637);
or OR4 (N19752, N19745, N19302, N19589, N17057);
nand NAND2 (N19753, N19751, N634);
nand NAND3 (N19754, N19746, N18545, N8052);
nand NAND4 (N19755, N19743, N10564, N8188, N17027);
xor XOR2 (N19756, N19747, N8516);
xor XOR2 (N19757, N19754, N8425);
and AND4 (N19758, N19713, N18284, N5309, N8390);
not NOT1 (N19759, N19758);
xor XOR2 (N19760, N19752, N19611);
xor XOR2 (N19761, N19757, N8796);
xor XOR2 (N19762, N19731, N15026);
nor NOR4 (N19763, N19761, N19577, N3580, N15673);
xor XOR2 (N19764, N19760, N14419);
not NOT1 (N19765, N19763);
nor NOR3 (N19766, N19753, N5200, N14431);
buf BUF1 (N19767, N19764);
or OR4 (N19768, N19729, N12271, N5932, N18089);
xor XOR2 (N19769, N19765, N16908);
and AND3 (N19770, N19756, N9677, N2905);
and AND2 (N19771, N19768, N16566);
or OR4 (N19772, N19749, N11487, N4557, N5892);
not NOT1 (N19773, N19766);
or OR3 (N19774, N19767, N8428, N13226);
nor NOR4 (N19775, N19762, N9939, N7753, N10079);
xor XOR2 (N19776, N19759, N13764);
not NOT1 (N19777, N19774);
and AND4 (N19778, N19769, N8401, N66, N2047);
nor NOR2 (N19779, N19770, N3895);
and AND3 (N19780, N19775, N12099, N9104);
xor XOR2 (N19781, N19773, N14986);
or OR3 (N19782, N19780, N9976, N6281);
not NOT1 (N19783, N19772);
nand NAND2 (N19784, N19781, N6916);
buf BUF1 (N19785, N19777);
nor NOR3 (N19786, N19755, N11393, N11932);
and AND4 (N19787, N19782, N11023, N10210, N19725);
and AND2 (N19788, N19776, N19711);
or OR3 (N19789, N19784, N8900, N10747);
nor NOR2 (N19790, N19788, N7492);
buf BUF1 (N19791, N19786);
nor NOR3 (N19792, N19787, N6787, N15331);
nand NAND3 (N19793, N19783, N19267, N1469);
buf BUF1 (N19794, N19771);
xor XOR2 (N19795, N19794, N14065);
not NOT1 (N19796, N19785);
buf BUF1 (N19797, N19793);
and AND2 (N19798, N19791, N11976);
buf BUF1 (N19799, N19748);
xor XOR2 (N19800, N19796, N17602);
buf BUF1 (N19801, N19797);
and AND4 (N19802, N19800, N12522, N12200, N10289);
or OR3 (N19803, N19792, N8262, N1756);
nand NAND3 (N19804, N19789, N18475, N17096);
or OR3 (N19805, N19779, N17448, N1750);
not NOT1 (N19806, N19798);
and AND4 (N19807, N19806, N7734, N11438, N16993);
not NOT1 (N19808, N19807);
and AND3 (N19809, N19795, N8864, N12285);
or OR2 (N19810, N19778, N16897);
nand NAND3 (N19811, N19801, N10066, N14914);
and AND2 (N19812, N19808, N12216);
or OR4 (N19813, N19811, N19658, N219, N17452);
buf BUF1 (N19814, N19790);
nand NAND2 (N19815, N19810, N5102);
nor NOR4 (N19816, N19809, N11956, N18775, N3753);
xor XOR2 (N19817, N19803, N16956);
and AND4 (N19818, N19804, N1358, N16667, N12385);
xor XOR2 (N19819, N19805, N18976);
buf BUF1 (N19820, N19817);
xor XOR2 (N19821, N19818, N4652);
nor NOR2 (N19822, N19802, N8608);
not NOT1 (N19823, N19814);
not NOT1 (N19824, N19820);
or OR3 (N19825, N19824, N14671, N10593);
and AND3 (N19826, N19821, N1836, N3237);
nand NAND4 (N19827, N19826, N9312, N3088, N5100);
xor XOR2 (N19828, N19819, N13590);
buf BUF1 (N19829, N19825);
and AND3 (N19830, N19827, N11847, N11422);
buf BUF1 (N19831, N19828);
nor NOR3 (N19832, N19813, N3565, N1666);
buf BUF1 (N19833, N19823);
and AND2 (N19834, N19799, N19447);
nand NAND4 (N19835, N19834, N1111, N8102, N6146);
or OR2 (N19836, N19822, N4204);
and AND3 (N19837, N19816, N11102, N3085);
and AND3 (N19838, N19833, N11857, N12328);
buf BUF1 (N19839, N19830);
buf BUF1 (N19840, N19829);
nor NOR3 (N19841, N19839, N3889, N6322);
xor XOR2 (N19842, N19836, N16921);
and AND4 (N19843, N19838, N4433, N12535, N11893);
or OR4 (N19844, N19837, N15238, N2197, N19078);
xor XOR2 (N19845, N19831, N12360);
or OR3 (N19846, N19812, N6084, N9275);
nand NAND4 (N19847, N19845, N982, N13964, N15907);
or OR2 (N19848, N19840, N3976);
and AND3 (N19849, N19841, N13185, N7508);
nor NOR4 (N19850, N19849, N17500, N16581, N18709);
nor NOR4 (N19851, N19843, N14783, N8649, N12093);
nor NOR2 (N19852, N19847, N10657);
xor XOR2 (N19853, N19851, N7916);
or OR2 (N19854, N19848, N8343);
or OR2 (N19855, N19853, N4551);
not NOT1 (N19856, N19854);
buf BUF1 (N19857, N19842);
buf BUF1 (N19858, N19832);
buf BUF1 (N19859, N19858);
not NOT1 (N19860, N19844);
xor XOR2 (N19861, N19857, N5134);
nor NOR2 (N19862, N19861, N363);
xor XOR2 (N19863, N19856, N5725);
buf BUF1 (N19864, N19855);
or OR3 (N19865, N19835, N8195, N116);
buf BUF1 (N19866, N19862);
or OR3 (N19867, N19860, N3923, N17827);
nor NOR2 (N19868, N19852, N330);
and AND3 (N19869, N19850, N14545, N18893);
nor NOR3 (N19870, N19866, N1013, N11747);
buf BUF1 (N19871, N19859);
buf BUF1 (N19872, N19871);
and AND4 (N19873, N19846, N15827, N11504, N18966);
nand NAND2 (N19874, N19864, N17306);
xor XOR2 (N19875, N19872, N7718);
or OR3 (N19876, N19870, N18430, N18610);
buf BUF1 (N19877, N19873);
and AND4 (N19878, N19869, N1703, N6109, N12101);
or OR3 (N19879, N19867, N4565, N13728);
nor NOR3 (N19880, N19879, N18240, N17657);
not NOT1 (N19881, N19874);
or OR2 (N19882, N19863, N1547);
not NOT1 (N19883, N19880);
xor XOR2 (N19884, N19881, N5820);
not NOT1 (N19885, N19865);
xor XOR2 (N19886, N19885, N9363);
or OR4 (N19887, N19815, N7805, N13689, N2715);
and AND4 (N19888, N19887, N19072, N19274, N2817);
or OR4 (N19889, N19876, N4009, N19085, N16564);
not NOT1 (N19890, N19886);
nand NAND3 (N19891, N19882, N11156, N16815);
nand NAND3 (N19892, N19889, N8612, N14869);
not NOT1 (N19893, N19892);
and AND3 (N19894, N19877, N6014, N14654);
nor NOR4 (N19895, N19890, N17129, N3213, N2767);
nor NOR4 (N19896, N19894, N9171, N15574, N14703);
xor XOR2 (N19897, N19884, N7454);
and AND2 (N19898, N19893, N16571);
or OR4 (N19899, N19875, N12801, N12777, N8264);
nor NOR4 (N19900, N19891, N13304, N2044, N15501);
and AND2 (N19901, N19896, N16336);
buf BUF1 (N19902, N19898);
nor NOR3 (N19903, N19902, N16265, N6444);
nor NOR2 (N19904, N19903, N6400);
nand NAND3 (N19905, N19897, N8063, N15009);
nor NOR4 (N19906, N19900, N17495, N17733, N1866);
nor NOR4 (N19907, N19868, N9098, N18803, N2373);
or OR4 (N19908, N19899, N5175, N12356, N17433);
xor XOR2 (N19909, N19888, N9266);
nand NAND4 (N19910, N19905, N7861, N3270, N7755);
and AND3 (N19911, N19901, N15841, N16667);
not NOT1 (N19912, N19907);
buf BUF1 (N19913, N19883);
nor NOR2 (N19914, N19909, N12291);
or OR4 (N19915, N19895, N191, N16726, N16702);
nand NAND3 (N19916, N19915, N556, N5719);
buf BUF1 (N19917, N19913);
not NOT1 (N19918, N19917);
not NOT1 (N19919, N19904);
and AND4 (N19920, N19916, N6047, N18910, N16006);
not NOT1 (N19921, N19908);
or OR3 (N19922, N19910, N308, N17923);
and AND4 (N19923, N19878, N12238, N4555, N15537);
nand NAND3 (N19924, N19912, N10463, N18017);
nor NOR2 (N19925, N19922, N2566);
or OR4 (N19926, N19925, N3347, N11899, N1115);
not NOT1 (N19927, N19926);
buf BUF1 (N19928, N19923);
and AND3 (N19929, N19918, N12121, N14908);
xor XOR2 (N19930, N19928, N12485);
nor NOR2 (N19931, N19924, N18479);
nand NAND4 (N19932, N19929, N16797, N7708, N2437);
and AND2 (N19933, N19914, N5302);
nand NAND4 (N19934, N19932, N4909, N14131, N4980);
buf BUF1 (N19935, N19927);
and AND3 (N19936, N19911, N14000, N1790);
xor XOR2 (N19937, N19906, N17085);
nand NAND2 (N19938, N19931, N3179);
xor XOR2 (N19939, N19921, N11567);
nand NAND2 (N19940, N19919, N558);
or OR4 (N19941, N19939, N4153, N8030, N8066);
xor XOR2 (N19942, N19937, N19304);
buf BUF1 (N19943, N19935);
and AND3 (N19944, N19920, N9165, N9462);
buf BUF1 (N19945, N19940);
not NOT1 (N19946, N19943);
not NOT1 (N19947, N19936);
buf BUF1 (N19948, N19945);
not NOT1 (N19949, N19942);
xor XOR2 (N19950, N19947, N19358);
and AND4 (N19951, N19938, N15726, N3512, N4529);
nor NOR3 (N19952, N19934, N14639, N15914);
or OR4 (N19953, N19946, N18488, N8722, N17969);
buf BUF1 (N19954, N19952);
not NOT1 (N19955, N19933);
or OR2 (N19956, N19949, N16624);
or OR3 (N19957, N19954, N5217, N2572);
buf BUF1 (N19958, N19941);
not NOT1 (N19959, N19951);
not NOT1 (N19960, N19958);
xor XOR2 (N19961, N19956, N10890);
buf BUF1 (N19962, N19944);
buf BUF1 (N19963, N19960);
nor NOR4 (N19964, N19962, N12213, N12755, N8496);
not NOT1 (N19965, N19963);
and AND2 (N19966, N19950, N6587);
not NOT1 (N19967, N19953);
buf BUF1 (N19968, N19967);
buf BUF1 (N19969, N19948);
buf BUF1 (N19970, N19930);
buf BUF1 (N19971, N19961);
and AND4 (N19972, N19966, N2964, N5036, N18058);
or OR4 (N19973, N19971, N729, N5167, N172);
nor NOR4 (N19974, N19968, N10910, N13611, N3804);
not NOT1 (N19975, N19964);
and AND2 (N19976, N19959, N10681);
not NOT1 (N19977, N19970);
nor NOR2 (N19978, N19975, N6005);
and AND4 (N19979, N19957, N16409, N13376, N18335);
and AND3 (N19980, N19976, N3221, N7373);
and AND2 (N19981, N19972, N12106);
buf BUF1 (N19982, N19973);
nor NOR4 (N19983, N19979, N14037, N4501, N4848);
and AND3 (N19984, N19955, N2559, N15221);
nor NOR3 (N19985, N19983, N1003, N18620);
or OR2 (N19986, N19974, N318);
or OR3 (N19987, N19965, N2568, N15097);
nand NAND3 (N19988, N19978, N11574, N18198);
not NOT1 (N19989, N19986);
and AND3 (N19990, N19977, N8793, N5210);
and AND3 (N19991, N19980, N15089, N12939);
and AND4 (N19992, N19987, N6160, N15080, N6465);
buf BUF1 (N19993, N19990);
nor NOR3 (N19994, N19992, N3949, N2384);
nand NAND3 (N19995, N19993, N4247, N15571);
or OR3 (N19996, N19995, N5477, N308);
nand NAND2 (N19997, N19982, N9747);
xor XOR2 (N19998, N19988, N5854);
and AND4 (N19999, N19989, N7092, N14740, N8109);
buf BUF1 (N20000, N19998);
or OR3 (N20001, N20000, N11412, N12337);
nor NOR4 (N20002, N19984, N14418, N18696, N3931);
xor XOR2 (N20003, N19969, N14215);
or OR4 (N20004, N19985, N4919, N3989, N13619);
nand NAND4 (N20005, N19997, N10179, N12295, N1242);
not NOT1 (N20006, N19999);
nand NAND3 (N20007, N19994, N7327, N13797);
xor XOR2 (N20008, N20003, N11745);
not NOT1 (N20009, N20007);
xor XOR2 (N20010, N20005, N5961);
or OR3 (N20011, N20010, N9701, N11674);
nand NAND3 (N20012, N19991, N18328, N11455);
xor XOR2 (N20013, N20002, N15526);
buf BUF1 (N20014, N20013);
and AND4 (N20015, N20011, N19471, N13207, N18366);
or OR4 (N20016, N20015, N11069, N16587, N14501);
buf BUF1 (N20017, N20006);
nor NOR4 (N20018, N20009, N11062, N15188, N1048);
and AND4 (N20019, N20017, N15605, N11317, N30);
nor NOR2 (N20020, N20016, N19385);
or OR2 (N20021, N19996, N17291);
and AND4 (N20022, N20019, N1787, N8977, N17151);
nor NOR4 (N20023, N20014, N7090, N4599, N17300);
or OR2 (N20024, N20012, N9409);
and AND4 (N20025, N20021, N1566, N8444, N5261);
buf BUF1 (N20026, N20018);
nor NOR3 (N20027, N19981, N14114, N4201);
not NOT1 (N20028, N20020);
not NOT1 (N20029, N20024);
and AND3 (N20030, N20022, N10618, N15570);
nand NAND2 (N20031, N20023, N10095);
xor XOR2 (N20032, N20004, N3805);
or OR2 (N20033, N20031, N1853);
not NOT1 (N20034, N20001);
xor XOR2 (N20035, N20027, N7975);
buf BUF1 (N20036, N20033);
and AND4 (N20037, N20026, N8421, N1788, N11592);
and AND3 (N20038, N20035, N14469, N499);
not NOT1 (N20039, N20032);
and AND4 (N20040, N20039, N4451, N18966, N9109);
and AND3 (N20041, N20008, N10305, N680);
nor NOR3 (N20042, N20028, N10367, N15707);
xor XOR2 (N20043, N20042, N12138);
nand NAND3 (N20044, N20030, N5147, N6815);
and AND3 (N20045, N20040, N9018, N481);
xor XOR2 (N20046, N20034, N10126);
and AND4 (N20047, N20043, N15568, N11601, N9231);
xor XOR2 (N20048, N20041, N10645);
or OR4 (N20049, N20037, N8314, N5092, N1427);
and AND3 (N20050, N20044, N2951, N18381);
nand NAND2 (N20051, N20025, N14708);
buf BUF1 (N20052, N20045);
and AND2 (N20053, N20029, N13373);
nor NOR2 (N20054, N20051, N19510);
nor NOR2 (N20055, N20038, N18253);
not NOT1 (N20056, N20036);
not NOT1 (N20057, N20048);
and AND4 (N20058, N20047, N637, N4859, N11670);
or OR3 (N20059, N20053, N17143, N5232);
or OR3 (N20060, N20057, N18583, N9225);
nand NAND3 (N20061, N20059, N6322, N1479);
and AND3 (N20062, N20060, N11035, N16840);
not NOT1 (N20063, N20050);
and AND2 (N20064, N20062, N6063);
buf BUF1 (N20065, N20061);
or OR3 (N20066, N20052, N5913, N17773);
xor XOR2 (N20067, N20055, N7137);
not NOT1 (N20068, N20065);
buf BUF1 (N20069, N20054);
xor XOR2 (N20070, N20049, N10643);
buf BUF1 (N20071, N20066);
or OR4 (N20072, N20056, N2675, N999, N176);
not NOT1 (N20073, N20046);
nand NAND2 (N20074, N20067, N14296);
nor NOR2 (N20075, N20068, N5745);
and AND4 (N20076, N20075, N17209, N13025, N3231);
not NOT1 (N20077, N20069);
and AND2 (N20078, N20077, N1108);
nand NAND4 (N20079, N20076, N12869, N1126, N7203);
nor NOR2 (N20080, N20072, N10732);
or OR2 (N20081, N20070, N18219);
not NOT1 (N20082, N20080);
or OR2 (N20083, N20081, N2168);
xor XOR2 (N20084, N20083, N18662);
xor XOR2 (N20085, N20063, N19487);
nand NAND3 (N20086, N20084, N13808, N926);
xor XOR2 (N20087, N20086, N13513);
xor XOR2 (N20088, N20087, N14482);
or OR3 (N20089, N20074, N10692, N13941);
or OR4 (N20090, N20082, N14964, N11336, N9160);
nor NOR3 (N20091, N20071, N17995, N3574);
or OR3 (N20092, N20064, N17479, N13209);
or OR2 (N20093, N20091, N2072);
xor XOR2 (N20094, N20092, N8075);
nor NOR2 (N20095, N20089, N4880);
xor XOR2 (N20096, N20095, N18149);
or OR3 (N20097, N20096, N17926, N719);
xor XOR2 (N20098, N20097, N1477);
and AND4 (N20099, N20058, N16281, N4247, N15155);
not NOT1 (N20100, N20079);
xor XOR2 (N20101, N20085, N15412);
nor NOR2 (N20102, N20090, N9909);
nand NAND2 (N20103, N20102, N3447);
xor XOR2 (N20104, N20094, N2700);
nand NAND4 (N20105, N20099, N5926, N10115, N18466);
xor XOR2 (N20106, N20073, N9880);
buf BUF1 (N20107, N20088);
not NOT1 (N20108, N20100);
buf BUF1 (N20109, N20101);
xor XOR2 (N20110, N20093, N16066);
not NOT1 (N20111, N20078);
or OR2 (N20112, N20107, N6311);
and AND2 (N20113, N20103, N16541);
xor XOR2 (N20114, N20098, N8416);
nand NAND2 (N20115, N20110, N10324);
nand NAND3 (N20116, N20112, N19051, N1380);
buf BUF1 (N20117, N20108);
xor XOR2 (N20118, N20111, N4838);
or OR4 (N20119, N20116, N15298, N112, N11134);
xor XOR2 (N20120, N20105, N6597);
and AND3 (N20121, N20106, N1667, N15304);
buf BUF1 (N20122, N20117);
not NOT1 (N20123, N20118);
not NOT1 (N20124, N20113);
and AND3 (N20125, N20114, N7568, N3021);
nor NOR2 (N20126, N20115, N1917);
xor XOR2 (N20127, N20121, N17940);
or OR3 (N20128, N20123, N15371, N11546);
nand NAND2 (N20129, N20109, N1520);
and AND3 (N20130, N20104, N16066, N16957);
nand NAND3 (N20131, N20124, N257, N16988);
or OR2 (N20132, N20128, N5959);
or OR4 (N20133, N20132, N8153, N17524, N826);
xor XOR2 (N20134, N20119, N8663);
and AND4 (N20135, N20131, N9738, N11636, N1354);
buf BUF1 (N20136, N20122);
or OR3 (N20137, N20129, N6064, N11441);
buf BUF1 (N20138, N20130);
and AND4 (N20139, N20133, N100, N8976, N13097);
and AND2 (N20140, N20125, N9808);
buf BUF1 (N20141, N20134);
buf BUF1 (N20142, N20140);
or OR3 (N20143, N20126, N8484, N7179);
nand NAND3 (N20144, N20120, N13698, N13310);
nand NAND3 (N20145, N20135, N8210, N11068);
buf BUF1 (N20146, N20142);
nand NAND2 (N20147, N20143, N2233);
and AND4 (N20148, N20138, N2037, N3030, N3729);
and AND2 (N20149, N20139, N18689);
and AND3 (N20150, N20149, N17345, N5018);
xor XOR2 (N20151, N20146, N13634);
nor NOR2 (N20152, N20148, N13660);
nor NOR4 (N20153, N20152, N4132, N714, N16454);
and AND2 (N20154, N20153, N10700);
or OR4 (N20155, N20154, N8505, N11871, N15207);
not NOT1 (N20156, N20141);
nand NAND2 (N20157, N20151, N16431);
or OR3 (N20158, N20155, N16625, N2672);
buf BUF1 (N20159, N20150);
and AND3 (N20160, N20158, N5413, N16529);
and AND2 (N20161, N20157, N17720);
and AND2 (N20162, N20145, N16392);
nand NAND3 (N20163, N20136, N19849, N18025);
or OR2 (N20164, N20156, N18265);
and AND4 (N20165, N20137, N6084, N11958, N2224);
not NOT1 (N20166, N20165);
or OR4 (N20167, N20161, N7376, N12929, N19474);
or OR2 (N20168, N20166, N13280);
nor NOR4 (N20169, N20167, N5078, N720, N8244);
and AND3 (N20170, N20160, N8500, N11861);
nand NAND4 (N20171, N20159, N5582, N9436, N716);
xor XOR2 (N20172, N20168, N5355);
xor XOR2 (N20173, N20170, N13380);
not NOT1 (N20174, N20173);
or OR3 (N20175, N20172, N8239, N3378);
nand NAND3 (N20176, N20144, N3868, N3383);
not NOT1 (N20177, N20162);
buf BUF1 (N20178, N20175);
nor NOR3 (N20179, N20164, N12244, N15734);
and AND3 (N20180, N20163, N4966, N9220);
nor NOR4 (N20181, N20179, N4106, N1968, N19198);
nand NAND3 (N20182, N20181, N8718, N14770);
not NOT1 (N20183, N20147);
xor XOR2 (N20184, N20176, N19397);
not NOT1 (N20185, N20180);
and AND2 (N20186, N20174, N12370);
nor NOR2 (N20187, N20177, N13476);
or OR3 (N20188, N20127, N16208, N4936);
xor XOR2 (N20189, N20185, N6069);
nor NOR2 (N20190, N20182, N16882);
and AND4 (N20191, N20184, N14362, N1904, N15117);
or OR3 (N20192, N20169, N5318, N15475);
buf BUF1 (N20193, N20187);
buf BUF1 (N20194, N20186);
and AND2 (N20195, N20192, N7482);
and AND3 (N20196, N20195, N9523, N14865);
buf BUF1 (N20197, N20196);
and AND4 (N20198, N20183, N9601, N10340, N13013);
buf BUF1 (N20199, N20198);
and AND4 (N20200, N20199, N9096, N16729, N4706);
nor NOR3 (N20201, N20191, N7387, N1446);
buf BUF1 (N20202, N20193);
not NOT1 (N20203, N20197);
and AND4 (N20204, N20201, N18874, N13629, N8542);
and AND2 (N20205, N20189, N13068);
or OR3 (N20206, N20200, N9504, N2987);
buf BUF1 (N20207, N20190);
and AND3 (N20208, N20188, N1580, N18567);
nor NOR4 (N20209, N20171, N19590, N17636, N18358);
xor XOR2 (N20210, N20202, N6326);
buf BUF1 (N20211, N20208);
buf BUF1 (N20212, N20207);
not NOT1 (N20213, N20194);
xor XOR2 (N20214, N20206, N19641);
nand NAND2 (N20215, N20203, N10552);
buf BUF1 (N20216, N20204);
nand NAND2 (N20217, N20178, N10655);
xor XOR2 (N20218, N20215, N7840);
nor NOR4 (N20219, N20210, N18528, N9758, N2475);
or OR2 (N20220, N20209, N9235);
nor NOR4 (N20221, N20214, N9040, N4780, N7189);
buf BUF1 (N20222, N20217);
or OR4 (N20223, N20219, N7194, N8732, N13758);
nand NAND4 (N20224, N20221, N4316, N12069, N10668);
not NOT1 (N20225, N20222);
not NOT1 (N20226, N20205);
nand NAND2 (N20227, N20211, N16958);
and AND2 (N20228, N20227, N11559);
nand NAND4 (N20229, N20212, N18578, N11958, N10168);
buf BUF1 (N20230, N20228);
or OR3 (N20231, N20218, N7823, N1067);
xor XOR2 (N20232, N20220, N3997);
nor NOR4 (N20233, N20224, N16863, N17882, N4710);
xor XOR2 (N20234, N20233, N11403);
nand NAND2 (N20235, N20223, N1677);
or OR3 (N20236, N20226, N5446, N7257);
not NOT1 (N20237, N20235);
or OR4 (N20238, N20232, N6163, N10132, N371);
and AND4 (N20239, N20236, N11455, N3343, N11498);
nor NOR2 (N20240, N20237, N12499);
xor XOR2 (N20241, N20229, N19999);
xor XOR2 (N20242, N20225, N15870);
or OR2 (N20243, N20238, N13923);
and AND4 (N20244, N20216, N844, N1802, N4671);
buf BUF1 (N20245, N20241);
not NOT1 (N20246, N20213);
or OR2 (N20247, N20231, N12613);
or OR3 (N20248, N20239, N13815, N18917);
nand NAND2 (N20249, N20244, N13920);
buf BUF1 (N20250, N20240);
nor NOR4 (N20251, N20245, N13892, N6884, N7292);
and AND4 (N20252, N20243, N10853, N7731, N15007);
and AND2 (N20253, N20234, N1488);
xor XOR2 (N20254, N20246, N9195);
buf BUF1 (N20255, N20230);
nand NAND3 (N20256, N20254, N18064, N3428);
not NOT1 (N20257, N20255);
nor NOR3 (N20258, N20256, N15976, N3788);
xor XOR2 (N20259, N20250, N3903);
or OR3 (N20260, N20251, N17690, N18533);
and AND4 (N20261, N20257, N1977, N5607, N15423);
not NOT1 (N20262, N20248);
xor XOR2 (N20263, N20253, N12593);
and AND3 (N20264, N20260, N3519, N7256);
and AND4 (N20265, N20262, N16329, N20190, N18700);
not NOT1 (N20266, N20242);
not NOT1 (N20267, N20266);
buf BUF1 (N20268, N20252);
not NOT1 (N20269, N20261);
buf BUF1 (N20270, N20259);
buf BUF1 (N20271, N20270);
buf BUF1 (N20272, N20271);
xor XOR2 (N20273, N20247, N7744);
xor XOR2 (N20274, N20263, N13943);
or OR4 (N20275, N20269, N15499, N19908, N7119);
not NOT1 (N20276, N20267);
xor XOR2 (N20277, N20249, N7536);
xor XOR2 (N20278, N20268, N3120);
or OR3 (N20279, N20277, N9930, N15422);
not NOT1 (N20280, N20279);
xor XOR2 (N20281, N20276, N17875);
not NOT1 (N20282, N20258);
not NOT1 (N20283, N20273);
nor NOR2 (N20284, N20280, N14010);
and AND3 (N20285, N20264, N6982, N11093);
and AND3 (N20286, N20274, N16801, N10238);
xor XOR2 (N20287, N20272, N11527);
buf BUF1 (N20288, N20281);
nand NAND3 (N20289, N20285, N15551, N4675);
buf BUF1 (N20290, N20286);
buf BUF1 (N20291, N20287);
or OR4 (N20292, N20275, N3344, N4240, N19399);
or OR4 (N20293, N20290, N3526, N4914, N10230);
buf BUF1 (N20294, N20289);
not NOT1 (N20295, N20284);
nand NAND4 (N20296, N20283, N4621, N10897, N15507);
buf BUF1 (N20297, N20265);
or OR4 (N20298, N20291, N6739, N6294, N12072);
not NOT1 (N20299, N20288);
nand NAND2 (N20300, N20292, N6409);
xor XOR2 (N20301, N20295, N10177);
buf BUF1 (N20302, N20278);
xor XOR2 (N20303, N20299, N4382);
nand NAND3 (N20304, N20296, N12403, N7203);
xor XOR2 (N20305, N20297, N13396);
buf BUF1 (N20306, N20293);
buf BUF1 (N20307, N20306);
xor XOR2 (N20308, N20304, N11517);
xor XOR2 (N20309, N20298, N20036);
and AND4 (N20310, N20305, N7854, N16025, N16919);
and AND4 (N20311, N20302, N3578, N6168, N9915);
xor XOR2 (N20312, N20307, N16526);
nand NAND3 (N20313, N20308, N3718, N5277);
not NOT1 (N20314, N20282);
not NOT1 (N20315, N20311);
buf BUF1 (N20316, N20303);
nor NOR4 (N20317, N20314, N14571, N101, N12054);
nand NAND4 (N20318, N20316, N13213, N8976, N2668);
not NOT1 (N20319, N20300);
not NOT1 (N20320, N20313);
and AND3 (N20321, N20312, N8240, N16725);
buf BUF1 (N20322, N20319);
or OR4 (N20323, N20322, N5201, N14027, N17145);
and AND3 (N20324, N20309, N14911, N15781);
nor NOR3 (N20325, N20315, N13448, N13799);
not NOT1 (N20326, N20321);
buf BUF1 (N20327, N20301);
buf BUF1 (N20328, N20324);
nand NAND2 (N20329, N20294, N17180);
and AND3 (N20330, N20325, N4916, N3313);
nand NAND4 (N20331, N20323, N20176, N12818, N7920);
buf BUF1 (N20332, N20320);
xor XOR2 (N20333, N20326, N7979);
xor XOR2 (N20334, N20330, N12422);
nand NAND4 (N20335, N20317, N17524, N17324, N15521);
and AND3 (N20336, N20334, N15185, N18960);
or OR4 (N20337, N20328, N19852, N9729, N7724);
buf BUF1 (N20338, N20333);
and AND2 (N20339, N20337, N5673);
or OR2 (N20340, N20336, N4920);
buf BUF1 (N20341, N20338);
or OR3 (N20342, N20327, N10410, N53);
not NOT1 (N20343, N20331);
buf BUF1 (N20344, N20329);
not NOT1 (N20345, N20310);
xor XOR2 (N20346, N20344, N12585);
buf BUF1 (N20347, N20318);
not NOT1 (N20348, N20332);
not NOT1 (N20349, N20339);
nand NAND4 (N20350, N20342, N5015, N13324, N3474);
and AND4 (N20351, N20335, N10682, N5734, N10263);
and AND3 (N20352, N20341, N7717, N6917);
nand NAND2 (N20353, N20349, N6435);
not NOT1 (N20354, N20340);
nor NOR3 (N20355, N20343, N19058, N15418);
nand NAND4 (N20356, N20350, N8940, N11101, N8354);
nand NAND3 (N20357, N20354, N1259, N16051);
and AND3 (N20358, N20351, N19105, N13818);
or OR4 (N20359, N20347, N15242, N10204, N7101);
nand NAND3 (N20360, N20346, N7348, N4217);
or OR2 (N20361, N20353, N3826);
or OR2 (N20362, N20348, N7187);
nor NOR2 (N20363, N20359, N9953);
nor NOR4 (N20364, N20355, N3291, N701, N909);
not NOT1 (N20365, N20362);
buf BUF1 (N20366, N20345);
not NOT1 (N20367, N20361);
not NOT1 (N20368, N20367);
not NOT1 (N20369, N20358);
or OR3 (N20370, N20360, N19380, N13843);
nor NOR2 (N20371, N20364, N10500);
or OR4 (N20372, N20366, N20028, N4980, N13213);
nor NOR2 (N20373, N20372, N11529);
not NOT1 (N20374, N20370);
nor NOR3 (N20375, N20368, N64, N485);
xor XOR2 (N20376, N20371, N2689);
or OR4 (N20377, N20356, N5720, N6770, N284);
buf BUF1 (N20378, N20376);
buf BUF1 (N20379, N20373);
buf BUF1 (N20380, N20357);
or OR3 (N20381, N20378, N14723, N16501);
xor XOR2 (N20382, N20380, N7281);
buf BUF1 (N20383, N20377);
buf BUF1 (N20384, N20375);
not NOT1 (N20385, N20365);
not NOT1 (N20386, N20363);
and AND4 (N20387, N20352, N15431, N7711, N14878);
xor XOR2 (N20388, N20374, N5402);
xor XOR2 (N20389, N20385, N7345);
and AND4 (N20390, N20381, N20064, N14852, N18951);
buf BUF1 (N20391, N20379);
not NOT1 (N20392, N20388);
nor NOR3 (N20393, N20386, N14766, N16910);
and AND2 (N20394, N20383, N9163);
not NOT1 (N20395, N20392);
buf BUF1 (N20396, N20387);
or OR2 (N20397, N20395, N6379);
xor XOR2 (N20398, N20397, N14071);
or OR4 (N20399, N20393, N2574, N8222, N16958);
nand NAND3 (N20400, N20391, N76, N10028);
nand NAND3 (N20401, N20396, N8331, N9764);
buf BUF1 (N20402, N20389);
xor XOR2 (N20403, N20398, N14521);
not NOT1 (N20404, N20401);
or OR3 (N20405, N20399, N3995, N14929);
buf BUF1 (N20406, N20400);
nand NAND4 (N20407, N20403, N6616, N19438, N7097);
and AND4 (N20408, N20394, N16359, N4717, N8875);
nand NAND4 (N20409, N20402, N12817, N7263, N9145);
or OR4 (N20410, N20382, N5322, N10076, N8238);
nand NAND2 (N20411, N20410, N8062);
and AND2 (N20412, N20390, N15123);
or OR2 (N20413, N20412, N1311);
nand NAND3 (N20414, N20409, N4061, N16247);
buf BUF1 (N20415, N20407);
buf BUF1 (N20416, N20404);
xor XOR2 (N20417, N20415, N10494);
not NOT1 (N20418, N20369);
xor XOR2 (N20419, N20417, N14237);
and AND2 (N20420, N20418, N3075);
xor XOR2 (N20421, N20413, N13650);
or OR2 (N20422, N20405, N5785);
not NOT1 (N20423, N20384);
xor XOR2 (N20424, N20416, N4684);
not NOT1 (N20425, N20424);
nor NOR2 (N20426, N20419, N1217);
not NOT1 (N20427, N20425);
nand NAND3 (N20428, N20423, N9253, N2655);
and AND2 (N20429, N20411, N1156);
buf BUF1 (N20430, N20427);
nor NOR2 (N20431, N20429, N4514);
and AND4 (N20432, N20430, N17235, N8324, N12175);
and AND4 (N20433, N20431, N7715, N19874, N13039);
buf BUF1 (N20434, N20422);
or OR3 (N20435, N20434, N9411, N19655);
nor NOR4 (N20436, N20406, N15597, N7680, N11828);
nor NOR4 (N20437, N20436, N1812, N7661, N13690);
not NOT1 (N20438, N20432);
xor XOR2 (N20439, N20437, N13759);
buf BUF1 (N20440, N20421);
not NOT1 (N20441, N20438);
or OR2 (N20442, N20435, N6357);
or OR2 (N20443, N20426, N3767);
not NOT1 (N20444, N20414);
xor XOR2 (N20445, N20440, N4206);
xor XOR2 (N20446, N20444, N9096);
nor NOR2 (N20447, N20428, N20361);
nand NAND3 (N20448, N20433, N7618, N18928);
nor NOR2 (N20449, N20448, N18823);
and AND3 (N20450, N20443, N3791, N13877);
not NOT1 (N20451, N20446);
xor XOR2 (N20452, N20450, N17995);
or OR2 (N20453, N20441, N17924);
and AND3 (N20454, N20453, N1701, N14249);
or OR2 (N20455, N20408, N9426);
and AND2 (N20456, N20445, N4741);
or OR2 (N20457, N20439, N9887);
not NOT1 (N20458, N20449);
not NOT1 (N20459, N20456);
nand NAND4 (N20460, N20451, N20398, N11131, N7391);
or OR4 (N20461, N20442, N16044, N8177, N3396);
nand NAND3 (N20462, N20459, N2745, N13167);
nand NAND4 (N20463, N20454, N8468, N17272, N9477);
xor XOR2 (N20464, N20458, N17368);
and AND4 (N20465, N20457, N16012, N8992, N9583);
xor XOR2 (N20466, N20447, N11173);
not NOT1 (N20467, N20460);
or OR3 (N20468, N20420, N8058, N9977);
buf BUF1 (N20469, N20452);
xor XOR2 (N20470, N20465, N20153);
xor XOR2 (N20471, N20463, N14982);
nand NAND4 (N20472, N20469, N13712, N5764, N1188);
xor XOR2 (N20473, N20471, N11448);
xor XOR2 (N20474, N20467, N19006);
and AND3 (N20475, N20464, N12624, N1763);
nor NOR2 (N20476, N20461, N9414);
xor XOR2 (N20477, N20476, N3511);
xor XOR2 (N20478, N20477, N4869);
nand NAND4 (N20479, N20468, N2710, N4919, N10759);
xor XOR2 (N20480, N20466, N15622);
and AND3 (N20481, N20462, N13991, N14999);
and AND2 (N20482, N20474, N3987);
xor XOR2 (N20483, N20455, N14322);
buf BUF1 (N20484, N20472);
xor XOR2 (N20485, N20482, N16445);
and AND2 (N20486, N20484, N7370);
and AND3 (N20487, N20475, N10280, N20129);
xor XOR2 (N20488, N20478, N8359);
nand NAND4 (N20489, N20473, N11473, N18155, N9357);
not NOT1 (N20490, N20487);
buf BUF1 (N20491, N20481);
buf BUF1 (N20492, N20489);
buf BUF1 (N20493, N20491);
nor NOR3 (N20494, N20479, N4911, N118);
and AND3 (N20495, N20486, N19284, N5134);
and AND2 (N20496, N20470, N10947);
not NOT1 (N20497, N20488);
or OR3 (N20498, N20497, N3105, N20381);
and AND2 (N20499, N20485, N12845);
or OR3 (N20500, N20498, N849, N4984);
nand NAND4 (N20501, N20495, N14435, N15480, N20428);
and AND4 (N20502, N20493, N1074, N11212, N17120);
nand NAND3 (N20503, N20483, N19208, N3562);
buf BUF1 (N20504, N20490);
nand NAND4 (N20505, N20502, N2981, N2878, N18161);
buf BUF1 (N20506, N20494);
not NOT1 (N20507, N20499);
and AND3 (N20508, N20505, N2489, N2528);
nor NOR4 (N20509, N20506, N5994, N2815, N13851);
buf BUF1 (N20510, N20500);
nor NOR3 (N20511, N20509, N12996, N5443);
nor NOR4 (N20512, N20504, N6852, N18658, N2873);
and AND4 (N20513, N20512, N12350, N2344, N6431);
and AND2 (N20514, N20480, N4142);
xor XOR2 (N20515, N20511, N15764);
nand NAND4 (N20516, N20492, N8675, N2878, N5833);
xor XOR2 (N20517, N20508, N17276);
nand NAND2 (N20518, N20501, N405);
xor XOR2 (N20519, N20514, N9294);
not NOT1 (N20520, N20507);
xor XOR2 (N20521, N20503, N18600);
nand NAND4 (N20522, N20516, N8322, N16779, N1227);
nand NAND2 (N20523, N20521, N8713);
nand NAND4 (N20524, N20517, N19058, N18671, N8223);
and AND4 (N20525, N20524, N18245, N3066, N11049);
or OR3 (N20526, N20496, N14683, N3912);
not NOT1 (N20527, N20523);
buf BUF1 (N20528, N20513);
xor XOR2 (N20529, N20527, N14038);
nor NOR2 (N20530, N20528, N8396);
nor NOR4 (N20531, N20522, N6444, N18923, N14916);
and AND3 (N20532, N20526, N561, N12776);
and AND2 (N20533, N20530, N3431);
and AND4 (N20534, N20519, N9919, N1477, N18288);
or OR2 (N20535, N20533, N19503);
nand NAND4 (N20536, N20531, N2138, N11112, N14831);
not NOT1 (N20537, N20529);
nor NOR2 (N20538, N20515, N6333);
not NOT1 (N20539, N20536);
buf BUF1 (N20540, N20539);
buf BUF1 (N20541, N20535);
nand NAND3 (N20542, N20510, N1452, N5734);
buf BUF1 (N20543, N20518);
xor XOR2 (N20544, N20525, N18255);
and AND4 (N20545, N20541, N259, N1057, N9752);
not NOT1 (N20546, N20542);
buf BUF1 (N20547, N20540);
and AND3 (N20548, N20546, N13323, N10893);
buf BUF1 (N20549, N20544);
xor XOR2 (N20550, N20543, N17500);
xor XOR2 (N20551, N20537, N10262);
nand NAND4 (N20552, N20549, N10869, N10405, N19976);
and AND3 (N20553, N20545, N9209, N15366);
buf BUF1 (N20554, N20550);
nor NOR3 (N20555, N20534, N4146, N12960);
buf BUF1 (N20556, N20548);
xor XOR2 (N20557, N20555, N5471);
buf BUF1 (N20558, N20557);
buf BUF1 (N20559, N20538);
xor XOR2 (N20560, N20553, N8111);
and AND4 (N20561, N20532, N11845, N8665, N12824);
not NOT1 (N20562, N20554);
buf BUF1 (N20563, N20560);
nor NOR2 (N20564, N20559, N3425);
or OR3 (N20565, N20561, N2480, N14497);
and AND3 (N20566, N20562, N14846, N10371);
or OR2 (N20567, N20566, N19232);
xor XOR2 (N20568, N20552, N19509);
nand NAND3 (N20569, N20567, N10836, N19316);
nand NAND2 (N20570, N20556, N5554);
buf BUF1 (N20571, N20551);
buf BUF1 (N20572, N20569);
nand NAND3 (N20573, N20568, N17012, N9979);
xor XOR2 (N20574, N20570, N16463);
not NOT1 (N20575, N20563);
and AND3 (N20576, N20520, N16867, N19974);
and AND2 (N20577, N20547, N16468);
xor XOR2 (N20578, N20577, N8050);
not NOT1 (N20579, N20578);
not NOT1 (N20580, N20576);
or OR2 (N20581, N20571, N5466);
buf BUF1 (N20582, N20581);
buf BUF1 (N20583, N20572);
xor XOR2 (N20584, N20579, N5353);
nor NOR2 (N20585, N20580, N6214);
nor NOR4 (N20586, N20565, N19009, N13008, N6548);
nor NOR3 (N20587, N20584, N10877, N13978);
nor NOR4 (N20588, N20558, N46, N15864, N12869);
or OR4 (N20589, N20564, N1287, N15702, N16857);
buf BUF1 (N20590, N20587);
not NOT1 (N20591, N20574);
nand NAND3 (N20592, N20590, N2753, N9485);
xor XOR2 (N20593, N20586, N8463);
buf BUF1 (N20594, N20582);
or OR2 (N20595, N20593, N2039);
not NOT1 (N20596, N20591);
or OR4 (N20597, N20596, N15993, N7124, N6316);
xor XOR2 (N20598, N20588, N4177);
and AND4 (N20599, N20597, N12069, N7410, N11693);
xor XOR2 (N20600, N20575, N6602);
buf BUF1 (N20601, N20592);
or OR3 (N20602, N20595, N18003, N2678);
nor NOR3 (N20603, N20598, N3474, N214);
buf BUF1 (N20604, N20573);
nand NAND4 (N20605, N20599, N3107, N15025, N887);
xor XOR2 (N20606, N20583, N3865);
or OR2 (N20607, N20585, N16492);
and AND2 (N20608, N20589, N5819);
nor NOR4 (N20609, N20606, N16410, N5939, N3583);
buf BUF1 (N20610, N20602);
xor XOR2 (N20611, N20609, N8105);
xor XOR2 (N20612, N20603, N2781);
buf BUF1 (N20613, N20605);
nor NOR3 (N20614, N20601, N14272, N9050);
nor NOR2 (N20615, N20608, N19569);
xor XOR2 (N20616, N20604, N7045);
not NOT1 (N20617, N20607);
nor NOR4 (N20618, N20610, N9416, N9511, N5862);
or OR3 (N20619, N20600, N20060, N6607);
buf BUF1 (N20620, N20615);
not NOT1 (N20621, N20618);
buf BUF1 (N20622, N20621);
buf BUF1 (N20623, N20617);
nand NAND2 (N20624, N20623, N3851);
and AND3 (N20625, N20619, N9478, N8436);
not NOT1 (N20626, N20613);
nor NOR3 (N20627, N20626, N20377, N18002);
nand NAND4 (N20628, N20616, N18449, N7909, N6991);
buf BUF1 (N20629, N20624);
and AND3 (N20630, N20628, N8847, N5316);
buf BUF1 (N20631, N20612);
xor XOR2 (N20632, N20614, N8644);
xor XOR2 (N20633, N20632, N2199);
not NOT1 (N20634, N20630);
nand NAND3 (N20635, N20634, N18694, N17553);
nor NOR2 (N20636, N20625, N5981);
or OR2 (N20637, N20636, N11143);
and AND3 (N20638, N20622, N67, N5273);
xor XOR2 (N20639, N20594, N17772);
buf BUF1 (N20640, N20631);
and AND4 (N20641, N20629, N8444, N11957, N2446);
buf BUF1 (N20642, N20627);
buf BUF1 (N20643, N20638);
buf BUF1 (N20644, N20637);
or OR4 (N20645, N20642, N18694, N8039, N12637);
nor NOR4 (N20646, N20644, N12291, N4333, N6091);
nor NOR2 (N20647, N20639, N5643);
xor XOR2 (N20648, N20611, N798);
nand NAND4 (N20649, N20647, N5175, N6803, N16797);
or OR2 (N20650, N20620, N7976);
buf BUF1 (N20651, N20646);
nor NOR4 (N20652, N20645, N599, N18013, N14774);
nand NAND2 (N20653, N20635, N6229);
xor XOR2 (N20654, N20650, N13659);
not NOT1 (N20655, N20649);
not NOT1 (N20656, N20653);
nand NAND3 (N20657, N20656, N16005, N6127);
buf BUF1 (N20658, N20651);
not NOT1 (N20659, N20641);
xor XOR2 (N20660, N20655, N13628);
nor NOR3 (N20661, N20633, N947, N10649);
nor NOR4 (N20662, N20652, N3589, N17704, N17109);
not NOT1 (N20663, N20662);
or OR4 (N20664, N20663, N8727, N16983, N10503);
not NOT1 (N20665, N20660);
not NOT1 (N20666, N20659);
nand NAND2 (N20667, N20658, N6077);
and AND3 (N20668, N20667, N9986, N9864);
not NOT1 (N20669, N20664);
buf BUF1 (N20670, N20668);
not NOT1 (N20671, N20666);
nor NOR3 (N20672, N20648, N5494, N18482);
xor XOR2 (N20673, N20672, N6134);
nor NOR3 (N20674, N20643, N5931, N10541);
nand NAND2 (N20675, N20669, N17131);
xor XOR2 (N20676, N20670, N13633);
buf BUF1 (N20677, N20640);
or OR2 (N20678, N20673, N2312);
and AND3 (N20679, N20677, N17310, N19099);
or OR4 (N20680, N20676, N18394, N8251, N1232);
and AND3 (N20681, N20679, N13174, N17386);
xor XOR2 (N20682, N20657, N7911);
xor XOR2 (N20683, N20680, N17295);
buf BUF1 (N20684, N20678);
xor XOR2 (N20685, N20681, N13841);
or OR2 (N20686, N20661, N20276);
buf BUF1 (N20687, N20674);
and AND2 (N20688, N20665, N11892);
or OR4 (N20689, N20654, N7808, N6257, N7936);
and AND2 (N20690, N20671, N6368);
buf BUF1 (N20691, N20689);
or OR4 (N20692, N20675, N12386, N5581, N9507);
or OR2 (N20693, N20691, N7638);
and AND4 (N20694, N20682, N2456, N16045, N4921);
or OR4 (N20695, N20693, N8781, N14324, N9852);
nand NAND4 (N20696, N20685, N459, N12658, N16090);
not NOT1 (N20697, N20694);
nor NOR4 (N20698, N20690, N17593, N5394, N18605);
xor XOR2 (N20699, N20695, N10909);
and AND4 (N20700, N20686, N12494, N14817, N8060);
buf BUF1 (N20701, N20700);
and AND3 (N20702, N20696, N13459, N18343);
xor XOR2 (N20703, N20688, N7091);
or OR3 (N20704, N20684, N399, N17009);
not NOT1 (N20705, N20687);
not NOT1 (N20706, N20703);
and AND2 (N20707, N20699, N10403);
nand NAND2 (N20708, N20706, N17911);
nor NOR3 (N20709, N20692, N14969, N9691);
nand NAND4 (N20710, N20707, N2830, N13779, N5806);
xor XOR2 (N20711, N20708, N4218);
buf BUF1 (N20712, N20697);
not NOT1 (N20713, N20710);
nor NOR2 (N20714, N20712, N18383);
nand NAND2 (N20715, N20711, N15176);
and AND2 (N20716, N20715, N11465);
and AND2 (N20717, N20713, N13073);
nor NOR2 (N20718, N20683, N4996);
xor XOR2 (N20719, N20716, N5999);
nand NAND3 (N20720, N20704, N3514, N4526);
or OR2 (N20721, N20720, N2767);
nor NOR3 (N20722, N20719, N15874, N3907);
and AND4 (N20723, N20718, N4726, N9951, N16935);
buf BUF1 (N20724, N20722);
and AND3 (N20725, N20723, N2805, N7104);
nor NOR3 (N20726, N20717, N17574, N14618);
and AND4 (N20727, N20701, N7433, N4484, N6997);
nand NAND2 (N20728, N20727, N2104);
not NOT1 (N20729, N20698);
nor NOR4 (N20730, N20728, N5839, N5715, N14182);
nor NOR2 (N20731, N20705, N16912);
xor XOR2 (N20732, N20702, N17579);
xor XOR2 (N20733, N20731, N14307);
nand NAND3 (N20734, N20725, N14934, N11331);
nor NOR3 (N20735, N20709, N9375, N18901);
nand NAND2 (N20736, N20721, N8650);
buf BUF1 (N20737, N20726);
not NOT1 (N20738, N20736);
buf BUF1 (N20739, N20732);
xor XOR2 (N20740, N20735, N17051);
and AND3 (N20741, N20714, N16334, N2638);
nor NOR4 (N20742, N20738, N7315, N762, N15580);
and AND2 (N20743, N20724, N19453);
not NOT1 (N20744, N20741);
not NOT1 (N20745, N20729);
nand NAND2 (N20746, N20739, N20300);
nor NOR3 (N20747, N20740, N16037, N11428);
xor XOR2 (N20748, N20733, N18080);
buf BUF1 (N20749, N20748);
buf BUF1 (N20750, N20734);
and AND4 (N20751, N20742, N14002, N8261, N3019);
xor XOR2 (N20752, N20751, N12225);
nand NAND3 (N20753, N20743, N19979, N16280);
nand NAND2 (N20754, N20753, N16163);
buf BUF1 (N20755, N20730);
xor XOR2 (N20756, N20747, N13614);
nor NOR4 (N20757, N20750, N5074, N1452, N9293);
not NOT1 (N20758, N20744);
not NOT1 (N20759, N20752);
and AND3 (N20760, N20754, N1429, N6507);
nor NOR2 (N20761, N20737, N3635);
and AND3 (N20762, N20756, N10110, N15186);
buf BUF1 (N20763, N20761);
and AND3 (N20764, N20746, N13471, N956);
nor NOR4 (N20765, N20758, N8439, N12078, N8713);
xor XOR2 (N20766, N20757, N10523);
and AND2 (N20767, N20760, N2691);
or OR3 (N20768, N20755, N4267, N6403);
nand NAND3 (N20769, N20768, N6619, N5710);
or OR4 (N20770, N20769, N909, N6826, N500);
not NOT1 (N20771, N20764);
not NOT1 (N20772, N20771);
nand NAND2 (N20773, N20763, N12057);
and AND3 (N20774, N20749, N7745, N2246);
xor XOR2 (N20775, N20774, N13469);
or OR2 (N20776, N20762, N1961);
nand NAND4 (N20777, N20759, N14782, N2903, N15289);
not NOT1 (N20778, N20767);
xor XOR2 (N20779, N20745, N8394);
and AND4 (N20780, N20778, N16642, N1493, N14567);
nor NOR2 (N20781, N20777, N13785);
not NOT1 (N20782, N20765);
nor NOR2 (N20783, N20766, N19329);
nand NAND3 (N20784, N20775, N11009, N13341);
buf BUF1 (N20785, N20780);
buf BUF1 (N20786, N20772);
buf BUF1 (N20787, N20783);
xor XOR2 (N20788, N20786, N13401);
nand NAND2 (N20789, N20788, N13460);
not NOT1 (N20790, N20785);
nand NAND3 (N20791, N20782, N19521, N2138);
or OR4 (N20792, N20770, N1814, N8070, N1074);
not NOT1 (N20793, N20773);
not NOT1 (N20794, N20784);
and AND2 (N20795, N20779, N11576);
not NOT1 (N20796, N20794);
xor XOR2 (N20797, N20787, N5021);
nand NAND3 (N20798, N20789, N19169, N6792);
buf BUF1 (N20799, N20791);
and AND4 (N20800, N20793, N10268, N9460, N9824);
buf BUF1 (N20801, N20797);
not NOT1 (N20802, N20796);
xor XOR2 (N20803, N20801, N7542);
nand NAND4 (N20804, N20781, N9366, N6794, N14663);
nand NAND3 (N20805, N20804, N12684, N7464);
nor NOR4 (N20806, N20776, N5070, N18410, N3409);
buf BUF1 (N20807, N20795);
nor NOR3 (N20808, N20799, N13017, N19736);
xor XOR2 (N20809, N20792, N18908);
xor XOR2 (N20810, N20805, N12193);
or OR2 (N20811, N20809, N14211);
nand NAND3 (N20812, N20807, N15727, N16146);
or OR4 (N20813, N20808, N10579, N7009, N2545);
buf BUF1 (N20814, N20798);
nand NAND2 (N20815, N20812, N2359);
nor NOR4 (N20816, N20803, N17701, N14338, N10557);
not NOT1 (N20817, N20800);
buf BUF1 (N20818, N20814);
or OR3 (N20819, N20806, N7555, N19349);
and AND3 (N20820, N20816, N19383, N13895);
xor XOR2 (N20821, N20790, N4315);
not NOT1 (N20822, N20820);
and AND3 (N20823, N20815, N2990, N3373);
not NOT1 (N20824, N20818);
nor NOR3 (N20825, N20817, N13208, N17815);
nor NOR2 (N20826, N20819, N13584);
nand NAND2 (N20827, N20813, N8316);
or OR4 (N20828, N20825, N4932, N10134, N12080);
and AND4 (N20829, N20802, N16489, N531, N3396);
nor NOR2 (N20830, N20822, N17794);
nor NOR3 (N20831, N20821, N2028, N4947);
nor NOR4 (N20832, N20826, N11531, N11173, N5023);
nor NOR3 (N20833, N20823, N12119, N17777);
and AND2 (N20834, N20810, N15855);
nand NAND4 (N20835, N20811, N10904, N11999, N11797);
and AND4 (N20836, N20835, N10137, N16716, N6059);
or OR2 (N20837, N20832, N15847);
or OR4 (N20838, N20829, N8388, N11513, N4082);
buf BUF1 (N20839, N20827);
buf BUF1 (N20840, N20834);
or OR4 (N20841, N20833, N18933, N4193, N8814);
xor XOR2 (N20842, N20840, N11558);
and AND4 (N20843, N20836, N20637, N5478, N10016);
xor XOR2 (N20844, N20824, N16482);
nor NOR3 (N20845, N20837, N11394, N14474);
and AND3 (N20846, N20839, N13543, N16810);
not NOT1 (N20847, N20846);
xor XOR2 (N20848, N20831, N4799);
buf BUF1 (N20849, N20828);
buf BUF1 (N20850, N20830);
and AND4 (N20851, N20844, N17354, N14037, N15380);
buf BUF1 (N20852, N20851);
or OR3 (N20853, N20841, N3992, N626);
and AND3 (N20854, N20849, N5677, N4171);
or OR2 (N20855, N20843, N4664);
or OR3 (N20856, N20845, N10687, N12236);
and AND4 (N20857, N20847, N3723, N15919, N7644);
nor NOR2 (N20858, N20842, N11232);
or OR4 (N20859, N20856, N3566, N18006, N5208);
or OR3 (N20860, N20859, N20447, N20326);
not NOT1 (N20861, N20853);
or OR3 (N20862, N20857, N5858, N20044);
nor NOR4 (N20863, N20861, N5739, N20725, N10856);
nand NAND3 (N20864, N20838, N5113, N752);
xor XOR2 (N20865, N20848, N19805);
and AND2 (N20866, N20855, N88);
buf BUF1 (N20867, N20850);
nand NAND3 (N20868, N20862, N17060, N9187);
buf BUF1 (N20869, N20852);
and AND3 (N20870, N20869, N10463, N10202);
nand NAND3 (N20871, N20870, N10124, N1293);
nor NOR2 (N20872, N20860, N587);
nor NOR4 (N20873, N20868, N7700, N3891, N7436);
xor XOR2 (N20874, N20864, N8586);
nand NAND3 (N20875, N20871, N2336, N10997);
not NOT1 (N20876, N20867);
or OR2 (N20877, N20873, N14282);
not NOT1 (N20878, N20876);
nand NAND3 (N20879, N20878, N2348, N10838);
nor NOR3 (N20880, N20858, N18856, N291);
xor XOR2 (N20881, N20866, N17851);
xor XOR2 (N20882, N20880, N12648);
and AND3 (N20883, N20854, N8709, N20056);
nand NAND3 (N20884, N20865, N12149, N9192);
buf BUF1 (N20885, N20881);
or OR4 (N20886, N20879, N16595, N17789, N16049);
buf BUF1 (N20887, N20874);
buf BUF1 (N20888, N20883);
not NOT1 (N20889, N20872);
or OR2 (N20890, N20886, N8767);
buf BUF1 (N20891, N20890);
nor NOR4 (N20892, N20891, N10413, N5408, N2174);
buf BUF1 (N20893, N20892);
xor XOR2 (N20894, N20884, N17601);
nand NAND4 (N20895, N20877, N1117, N7950, N1115);
and AND4 (N20896, N20882, N17748, N11819, N3574);
nand NAND2 (N20897, N20863, N16607);
xor XOR2 (N20898, N20893, N14900);
nand NAND2 (N20899, N20889, N16653);
xor XOR2 (N20900, N20885, N19394);
xor XOR2 (N20901, N20897, N7490);
buf BUF1 (N20902, N20896);
xor XOR2 (N20903, N20888, N507);
xor XOR2 (N20904, N20895, N16873);
nand NAND3 (N20905, N20900, N871, N16336);
xor XOR2 (N20906, N20903, N8566);
nor NOR3 (N20907, N20898, N7104, N19980);
xor XOR2 (N20908, N20905, N15948);
or OR3 (N20909, N20902, N13558, N8141);
not NOT1 (N20910, N20875);
nand NAND4 (N20911, N20910, N15896, N17785, N18968);
xor XOR2 (N20912, N20894, N12502);
nor NOR3 (N20913, N20906, N11274, N6884);
xor XOR2 (N20914, N20899, N15252);
not NOT1 (N20915, N20911);
buf BUF1 (N20916, N20915);
not NOT1 (N20917, N20913);
buf BUF1 (N20918, N20907);
xor XOR2 (N20919, N20917, N1569);
not NOT1 (N20920, N20904);
not NOT1 (N20921, N20908);
or OR4 (N20922, N20919, N18885, N20739, N3495);
xor XOR2 (N20923, N20887, N4921);
nand NAND3 (N20924, N20912, N1330, N9003);
buf BUF1 (N20925, N20918);
nor NOR3 (N20926, N20914, N5085, N2057);
nor NOR4 (N20927, N20922, N1582, N4134, N7078);
not NOT1 (N20928, N20923);
not NOT1 (N20929, N20920);
buf BUF1 (N20930, N20921);
xor XOR2 (N20931, N20916, N17670);
buf BUF1 (N20932, N20925);
xor XOR2 (N20933, N20930, N15219);
buf BUF1 (N20934, N20931);
not NOT1 (N20935, N20933);
xor XOR2 (N20936, N20927, N1333);
and AND4 (N20937, N20936, N5531, N15389, N7711);
or OR3 (N20938, N20924, N9381, N3474);
nor NOR3 (N20939, N20901, N14620, N17807);
or OR3 (N20940, N20938, N12340, N7120);
xor XOR2 (N20941, N20935, N13706);
and AND4 (N20942, N20941, N7424, N5345, N13592);
xor XOR2 (N20943, N20909, N8197);
nand NAND4 (N20944, N20934, N9930, N13455, N7513);
not NOT1 (N20945, N20926);
and AND2 (N20946, N20939, N11213);
or OR2 (N20947, N20928, N20694);
buf BUF1 (N20948, N20937);
or OR2 (N20949, N20932, N19276);
buf BUF1 (N20950, N20948);
and AND2 (N20951, N20929, N10801);
and AND3 (N20952, N20945, N9071, N14370);
not NOT1 (N20953, N20951);
xor XOR2 (N20954, N20944, N14824);
buf BUF1 (N20955, N20946);
nand NAND4 (N20956, N20952, N2062, N6316, N20357);
buf BUF1 (N20957, N20947);
buf BUF1 (N20958, N20956);
or OR3 (N20959, N20949, N19039, N3683);
xor XOR2 (N20960, N20942, N15071);
nor NOR2 (N20961, N20958, N5148);
or OR4 (N20962, N20943, N10475, N20825, N2837);
or OR3 (N20963, N20962, N314, N2191);
nor NOR2 (N20964, N20961, N12025);
or OR2 (N20965, N20957, N2314);
nand NAND2 (N20966, N20954, N257);
buf BUF1 (N20967, N20966);
buf BUF1 (N20968, N20967);
nor NOR3 (N20969, N20959, N1855, N17404);
xor XOR2 (N20970, N20965, N5521);
buf BUF1 (N20971, N20955);
or OR4 (N20972, N20968, N19476, N14778, N17930);
nor NOR3 (N20973, N20963, N13911, N15558);
or OR2 (N20974, N20970, N5008);
or OR4 (N20975, N20953, N14068, N17083, N18714);
nand NAND4 (N20976, N20973, N18430, N15517, N758);
xor XOR2 (N20977, N20969, N8824);
not NOT1 (N20978, N20977);
buf BUF1 (N20979, N20971);
xor XOR2 (N20980, N20979, N6240);
nor NOR2 (N20981, N20960, N180);
nor NOR3 (N20982, N20940, N2884, N8457);
nand NAND3 (N20983, N20972, N20617, N18937);
nor NOR3 (N20984, N20978, N8682, N16745);
nand NAND3 (N20985, N20981, N1180, N12618);
and AND2 (N20986, N20974, N3731);
buf BUF1 (N20987, N20975);
nand NAND3 (N20988, N20982, N10826, N2783);
or OR2 (N20989, N20984, N19864);
nand NAND3 (N20990, N20985, N20149, N9677);
nor NOR4 (N20991, N20964, N18726, N16515, N16689);
and AND4 (N20992, N20950, N17520, N14620, N11407);
xor XOR2 (N20993, N20990, N18706);
xor XOR2 (N20994, N20993, N20803);
or OR3 (N20995, N20989, N5013, N20060);
nand NAND3 (N20996, N20994, N2698, N10316);
not NOT1 (N20997, N20986);
nor NOR3 (N20998, N20980, N15438, N8390);
and AND2 (N20999, N20992, N9650);
buf BUF1 (N21000, N20983);
and AND3 (N21001, N20988, N8100, N4893);
not NOT1 (N21002, N20999);
or OR4 (N21003, N21000, N20872, N7285, N20186);
or OR3 (N21004, N20991, N15221, N3414);
nor NOR2 (N21005, N20998, N15273);
buf BUF1 (N21006, N21001);
or OR2 (N21007, N20997, N7478);
and AND3 (N21008, N20996, N10, N12531);
nor NOR2 (N21009, N21005, N4123);
or OR4 (N21010, N21002, N18927, N14468, N8438);
nor NOR4 (N21011, N21007, N7398, N4257, N15126);
nor NOR2 (N21012, N21004, N7966);
not NOT1 (N21013, N20987);
or OR4 (N21014, N20976, N16620, N10747, N5895);
buf BUF1 (N21015, N21003);
xor XOR2 (N21016, N21013, N17963);
buf BUF1 (N21017, N21010);
not NOT1 (N21018, N21017);
nor NOR2 (N21019, N21006, N16605);
and AND4 (N21020, N21016, N12293, N11689, N14193);
nand NAND4 (N21021, N21015, N13405, N10251, N18421);
nor NOR4 (N21022, N21011, N20886, N3343, N3573);
and AND3 (N21023, N20995, N5884, N2440);
not NOT1 (N21024, N21021);
nand NAND2 (N21025, N21023, N15181);
xor XOR2 (N21026, N21024, N8421);
or OR4 (N21027, N21022, N16751, N11239, N7133);
not NOT1 (N21028, N21025);
nor NOR4 (N21029, N21014, N13014, N11433, N3430);
nand NAND3 (N21030, N21026, N11153, N1625);
and AND4 (N21031, N21009, N18502, N19288, N12648);
buf BUF1 (N21032, N21019);
buf BUF1 (N21033, N21032);
nand NAND2 (N21034, N21018, N1074);
not NOT1 (N21035, N21033);
not NOT1 (N21036, N21034);
not NOT1 (N21037, N21035);
nor NOR4 (N21038, N21020, N3156, N3825, N15211);
not NOT1 (N21039, N21012);
and AND2 (N21040, N21037, N11721);
nor NOR2 (N21041, N21028, N19918);
or OR3 (N21042, N21041, N20895, N16325);
not NOT1 (N21043, N21036);
not NOT1 (N21044, N21043);
and AND2 (N21045, N21030, N15457);
nand NAND3 (N21046, N21045, N8847, N8477);
xor XOR2 (N21047, N21029, N12617);
nand NAND4 (N21048, N21008, N16699, N20846, N3049);
not NOT1 (N21049, N21048);
xor XOR2 (N21050, N21047, N20937);
buf BUF1 (N21051, N21046);
buf BUF1 (N21052, N21040);
nand NAND3 (N21053, N21031, N17911, N17602);
xor XOR2 (N21054, N21049, N14327);
nor NOR2 (N21055, N21051, N19797);
nand NAND4 (N21056, N21050, N14196, N4781, N9044);
or OR2 (N21057, N21042, N10830);
nand NAND3 (N21058, N21052, N16296, N18529);
nor NOR4 (N21059, N21054, N15362, N1534, N16883);
not NOT1 (N21060, N21039);
xor XOR2 (N21061, N21060, N531);
and AND3 (N21062, N21061, N6484, N9622);
or OR2 (N21063, N21062, N15197);
and AND4 (N21064, N21057, N19701, N20437, N17805);
buf BUF1 (N21065, N21063);
buf BUF1 (N21066, N21044);
not NOT1 (N21067, N21056);
not NOT1 (N21068, N21059);
nand NAND4 (N21069, N21053, N317, N14755, N12906);
and AND3 (N21070, N21069, N11541, N7258);
and AND4 (N21071, N21065, N16206, N1637, N11590);
or OR4 (N21072, N21038, N768, N15836, N423);
xor XOR2 (N21073, N21068, N6873);
buf BUF1 (N21074, N21027);
or OR3 (N21075, N21071, N12972, N1519);
and AND2 (N21076, N21072, N19287);
not NOT1 (N21077, N21067);
buf BUF1 (N21078, N21058);
not NOT1 (N21079, N21055);
not NOT1 (N21080, N21070);
nand NAND2 (N21081, N21066, N789);
nor NOR4 (N21082, N21081, N16529, N3921, N15966);
and AND2 (N21083, N21080, N5825);
not NOT1 (N21084, N21082);
xor XOR2 (N21085, N21076, N17881);
or OR3 (N21086, N21084, N13552, N10285);
nand NAND4 (N21087, N21074, N20468, N13399, N6934);
buf BUF1 (N21088, N21086);
buf BUF1 (N21089, N21073);
nor NOR3 (N21090, N21078, N6086, N12770);
not NOT1 (N21091, N21087);
not NOT1 (N21092, N21075);
xor XOR2 (N21093, N21091, N20143);
buf BUF1 (N21094, N21083);
xor XOR2 (N21095, N21094, N4944);
not NOT1 (N21096, N21095);
nor NOR2 (N21097, N21079, N20145);
not NOT1 (N21098, N21088);
nand NAND3 (N21099, N21089, N13119, N1200);
xor XOR2 (N21100, N21093, N12313);
nor NOR2 (N21101, N21097, N10591);
and AND4 (N21102, N21101, N725, N13634, N19561);
xor XOR2 (N21103, N21090, N8986);
not NOT1 (N21104, N21099);
or OR2 (N21105, N21102, N15435);
nand NAND4 (N21106, N21098, N12959, N2245, N20374);
xor XOR2 (N21107, N21105, N14498);
xor XOR2 (N21108, N21085, N13449);
nand NAND3 (N21109, N21100, N10143, N15827);
xor XOR2 (N21110, N21104, N5293);
nor NOR4 (N21111, N21077, N3715, N17400, N2664);
or OR4 (N21112, N21103, N10446, N15069, N16461);
nand NAND3 (N21113, N21108, N6097, N2224);
nand NAND4 (N21114, N21110, N1333, N10204, N12863);
nand NAND4 (N21115, N21113, N7138, N7735, N11694);
not NOT1 (N21116, N21092);
not NOT1 (N21117, N21111);
not NOT1 (N21118, N21112);
nand NAND2 (N21119, N21116, N4497);
nor NOR2 (N21120, N21115, N15653);
not NOT1 (N21121, N21120);
nor NOR4 (N21122, N21117, N256, N346, N211);
nor NOR3 (N21123, N21109, N12180, N13792);
xor XOR2 (N21124, N21114, N17133);
nand NAND4 (N21125, N21064, N3371, N14227, N7904);
not NOT1 (N21126, N21122);
xor XOR2 (N21127, N21126, N16814);
xor XOR2 (N21128, N21125, N18734);
xor XOR2 (N21129, N21127, N12420);
nor NOR2 (N21130, N21118, N15638);
and AND2 (N21131, N21106, N16038);
and AND4 (N21132, N21096, N10118, N18346, N13264);
and AND4 (N21133, N21123, N12074, N6620, N19809);
xor XOR2 (N21134, N21124, N18329);
nor NOR4 (N21135, N21121, N19098, N473, N16095);
buf BUF1 (N21136, N21131);
or OR4 (N21137, N21107, N6216, N1757, N6558);
or OR3 (N21138, N21136, N19282, N20261);
xor XOR2 (N21139, N21138, N9115);
nor NOR3 (N21140, N21137, N5123, N3502);
nand NAND3 (N21141, N21139, N18628, N6205);
nand NAND3 (N21142, N21129, N12590, N15346);
nand NAND2 (N21143, N21119, N5277);
nand NAND2 (N21144, N21140, N6451);
buf BUF1 (N21145, N21141);
nor NOR3 (N21146, N21143, N19437, N13525);
and AND2 (N21147, N21145, N9706);
nor NOR4 (N21148, N21135, N11418, N17494, N6799);
and AND4 (N21149, N21148, N17432, N5953, N16125);
and AND3 (N21150, N21128, N9670, N9824);
nor NOR4 (N21151, N21133, N13209, N10198, N14925);
xor XOR2 (N21152, N21142, N17183);
xor XOR2 (N21153, N21130, N9297);
or OR3 (N21154, N21150, N6674, N6599);
or OR2 (N21155, N21151, N8886);
or OR2 (N21156, N21155, N11164);
nor NOR2 (N21157, N21153, N16533);
xor XOR2 (N21158, N21157, N17296);
buf BUF1 (N21159, N21144);
xor XOR2 (N21160, N21134, N2157);
nor NOR2 (N21161, N21156, N16086);
or OR2 (N21162, N21161, N888);
nor NOR4 (N21163, N21149, N1094, N6203, N6426);
or OR4 (N21164, N21158, N13704, N10278, N10027);
nand NAND4 (N21165, N21162, N3865, N4281, N2095);
nor NOR3 (N21166, N21146, N9188, N17260);
and AND4 (N21167, N21152, N11565, N4644, N9425);
nor NOR2 (N21168, N21160, N13416);
or OR4 (N21169, N21165, N10924, N1363, N18057);
nand NAND2 (N21170, N21166, N7647);
or OR2 (N21171, N21168, N4090);
nor NOR2 (N21172, N21163, N20488);
nand NAND4 (N21173, N21171, N14396, N1438, N16705);
buf BUF1 (N21174, N21159);
nor NOR3 (N21175, N21174, N2745, N4403);
not NOT1 (N21176, N21147);
not NOT1 (N21177, N21167);
not NOT1 (N21178, N21175);
buf BUF1 (N21179, N21170);
buf BUF1 (N21180, N21179);
not NOT1 (N21181, N21173);
nand NAND2 (N21182, N21176, N8631);
nand NAND4 (N21183, N21154, N9548, N5108, N8734);
or OR2 (N21184, N21182, N18961);
xor XOR2 (N21185, N21178, N11711);
xor XOR2 (N21186, N21185, N12921);
and AND3 (N21187, N21180, N16724, N3769);
or OR2 (N21188, N21183, N10586);
or OR2 (N21189, N21169, N15442);
and AND2 (N21190, N21164, N9659);
and AND3 (N21191, N21184, N2365, N17942);
buf BUF1 (N21192, N21132);
and AND3 (N21193, N21181, N10966, N6991);
xor XOR2 (N21194, N21191, N5817);
xor XOR2 (N21195, N21188, N16422);
xor XOR2 (N21196, N21172, N224);
xor XOR2 (N21197, N21187, N15164);
or OR2 (N21198, N21197, N20461);
nor NOR4 (N21199, N21177, N18828, N14429, N13311);
nor NOR4 (N21200, N21196, N482, N10550, N15022);
buf BUF1 (N21201, N21193);
buf BUF1 (N21202, N21195);
nand NAND3 (N21203, N21186, N7282, N3340);
and AND4 (N21204, N21190, N18522, N15575, N20566);
xor XOR2 (N21205, N21204, N13957);
nand NAND3 (N21206, N21201, N6910, N19240);
nor NOR4 (N21207, N21206, N19473, N20938, N799);
nand NAND3 (N21208, N21199, N7706, N15628);
nand NAND4 (N21209, N21194, N6635, N11469, N10073);
not NOT1 (N21210, N21203);
and AND3 (N21211, N21210, N16331, N5418);
nor NOR4 (N21212, N21198, N1471, N19128, N12436);
nor NOR2 (N21213, N21209, N14384);
buf BUF1 (N21214, N21207);
not NOT1 (N21215, N21189);
nand NAND4 (N21216, N21202, N11482, N4868, N16070);
not NOT1 (N21217, N21205);
not NOT1 (N21218, N21216);
or OR4 (N21219, N21218, N6024, N2200, N13389);
and AND4 (N21220, N21211, N18226, N16833, N835);
nor NOR3 (N21221, N21217, N15716, N11758);
or OR2 (N21222, N21220, N14429);
and AND4 (N21223, N21214, N17971, N5329, N14698);
nand NAND4 (N21224, N21213, N17924, N20765, N20489);
buf BUF1 (N21225, N21224);
xor XOR2 (N21226, N21212, N1202);
buf BUF1 (N21227, N21221);
buf BUF1 (N21228, N21219);
buf BUF1 (N21229, N21200);
not NOT1 (N21230, N21223);
and AND2 (N21231, N21192, N20008);
nand NAND4 (N21232, N21228, N20246, N9095, N15082);
xor XOR2 (N21233, N21208, N19711);
buf BUF1 (N21234, N21229);
nand NAND4 (N21235, N21225, N20356, N13079, N6666);
and AND2 (N21236, N21232, N12565);
xor XOR2 (N21237, N21236, N14099);
nand NAND4 (N21238, N21235, N711, N44, N7652);
and AND3 (N21239, N21238, N2447, N3141);
not NOT1 (N21240, N21226);
and AND3 (N21241, N21222, N14139, N13449);
and AND3 (N21242, N21237, N13644, N11487);
nand NAND2 (N21243, N21231, N8727);
and AND3 (N21244, N21215, N19467, N5005);
not NOT1 (N21245, N21240);
xor XOR2 (N21246, N21230, N18694);
or OR2 (N21247, N21243, N11151);
nor NOR4 (N21248, N21246, N8038, N15837, N15326);
nor NOR2 (N21249, N21242, N6318);
nand NAND3 (N21250, N21249, N433, N7725);
nand NAND3 (N21251, N21248, N13634, N4198);
nor NOR2 (N21252, N21239, N16431);
nor NOR3 (N21253, N21241, N16079, N17882);
xor XOR2 (N21254, N21244, N13503);
and AND2 (N21255, N21233, N17419);
xor XOR2 (N21256, N21247, N8542);
xor XOR2 (N21257, N21250, N17880);
nand NAND3 (N21258, N21251, N11403, N5034);
not NOT1 (N21259, N21234);
not NOT1 (N21260, N21257);
and AND4 (N21261, N21252, N12579, N4826, N16199);
buf BUF1 (N21262, N21245);
buf BUF1 (N21263, N21256);
or OR2 (N21264, N21254, N3477);
nand NAND3 (N21265, N21259, N6960, N21089);
not NOT1 (N21266, N21255);
or OR2 (N21267, N21261, N14218);
or OR4 (N21268, N21258, N8144, N17605, N8113);
not NOT1 (N21269, N21267);
nand NAND4 (N21270, N21253, N6552, N1567, N10108);
or OR3 (N21271, N21262, N9535, N12318);
nor NOR2 (N21272, N21266, N11338);
or OR2 (N21273, N21270, N1565);
nor NOR3 (N21274, N21263, N19715, N9785);
or OR3 (N21275, N21272, N5283, N1234);
not NOT1 (N21276, N21271);
nor NOR4 (N21277, N21275, N13175, N3802, N4664);
or OR4 (N21278, N21269, N8349, N13766, N16489);
xor XOR2 (N21279, N21276, N1821);
or OR4 (N21280, N21227, N13347, N19533, N18722);
and AND3 (N21281, N21273, N600, N2682);
xor XOR2 (N21282, N21279, N4166);
nand NAND2 (N21283, N21282, N20232);
buf BUF1 (N21284, N21268);
buf BUF1 (N21285, N21283);
and AND4 (N21286, N21264, N10134, N12332, N7505);
xor XOR2 (N21287, N21274, N19487);
and AND3 (N21288, N21286, N20727, N3919);
buf BUF1 (N21289, N21260);
nand NAND2 (N21290, N21280, N4114);
nor NOR3 (N21291, N21288, N8098, N789);
or OR3 (N21292, N21290, N8884, N21208);
or OR3 (N21293, N21285, N15827, N8754);
buf BUF1 (N21294, N21278);
buf BUF1 (N21295, N21284);
nor NOR3 (N21296, N21293, N3906, N7170);
and AND4 (N21297, N21289, N19777, N694, N1205);
nor NOR4 (N21298, N21297, N4451, N17149, N6718);
nand NAND4 (N21299, N21298, N16045, N17671, N9147);
nor NOR3 (N21300, N21291, N21174, N18436);
and AND2 (N21301, N21277, N10933);
not NOT1 (N21302, N21294);
nor NOR2 (N21303, N21299, N16875);
xor XOR2 (N21304, N21292, N10628);
not NOT1 (N21305, N21295);
or OR2 (N21306, N21296, N16803);
or OR4 (N21307, N21301, N495, N5225, N16225);
and AND2 (N21308, N21307, N7295);
nor NOR3 (N21309, N21306, N16181, N4296);
xor XOR2 (N21310, N21308, N13660);
and AND4 (N21311, N21310, N13734, N20932, N16241);
buf BUF1 (N21312, N21302);
not NOT1 (N21313, N21265);
buf BUF1 (N21314, N21313);
buf BUF1 (N21315, N21300);
buf BUF1 (N21316, N21309);
not NOT1 (N21317, N21287);
not NOT1 (N21318, N21315);
nor NOR3 (N21319, N21318, N19506, N3580);
and AND3 (N21320, N21311, N18175, N8649);
not NOT1 (N21321, N21303);
xor XOR2 (N21322, N21312, N7653);
not NOT1 (N21323, N21314);
and AND4 (N21324, N21305, N18296, N14998, N9990);
nand NAND4 (N21325, N21320, N16728, N5700, N17895);
and AND3 (N21326, N21322, N10415, N7799);
and AND3 (N21327, N21316, N12953, N18160);
not NOT1 (N21328, N21281);
not NOT1 (N21329, N21328);
xor XOR2 (N21330, N21304, N3478);
or OR3 (N21331, N21317, N281, N12024);
xor XOR2 (N21332, N21327, N3626);
not NOT1 (N21333, N21321);
not NOT1 (N21334, N21332);
xor XOR2 (N21335, N21325, N1457);
nor NOR4 (N21336, N21323, N1546, N12721, N9230);
or OR4 (N21337, N21331, N8335, N11687, N4989);
not NOT1 (N21338, N21319);
or OR4 (N21339, N21329, N11648, N16747, N9160);
xor XOR2 (N21340, N21326, N6526);
nor NOR3 (N21341, N21340, N9706, N11078);
xor XOR2 (N21342, N21333, N12989);
nor NOR3 (N21343, N21337, N7208, N14594);
and AND3 (N21344, N21341, N11341, N19763);
nor NOR3 (N21345, N21339, N9175, N13980);
buf BUF1 (N21346, N21344);
buf BUF1 (N21347, N21324);
or OR4 (N21348, N21342, N11689, N12279, N623);
not NOT1 (N21349, N21336);
or OR4 (N21350, N21343, N2744, N20655, N15769);
and AND3 (N21351, N21335, N13156, N11289);
buf BUF1 (N21352, N21351);
xor XOR2 (N21353, N21348, N10148);
nor NOR3 (N21354, N21352, N8681, N8119);
buf BUF1 (N21355, N21353);
nor NOR3 (N21356, N21354, N3937, N7811);
nand NAND2 (N21357, N21330, N11458);
not NOT1 (N21358, N21345);
nand NAND3 (N21359, N21334, N19253, N7306);
nor NOR4 (N21360, N21359, N6501, N3895, N20180);
or OR2 (N21361, N21357, N20595);
xor XOR2 (N21362, N21360, N7968);
not NOT1 (N21363, N21358);
buf BUF1 (N21364, N21362);
and AND2 (N21365, N21356, N3190);
xor XOR2 (N21366, N21361, N7789);
not NOT1 (N21367, N21365);
nand NAND3 (N21368, N21363, N3200, N19847);
xor XOR2 (N21369, N21349, N6583);
xor XOR2 (N21370, N21346, N19666);
nor NOR3 (N21371, N21338, N7670, N3533);
xor XOR2 (N21372, N21364, N9947);
or OR2 (N21373, N21366, N20172);
not NOT1 (N21374, N21373);
xor XOR2 (N21375, N21368, N18817);
not NOT1 (N21376, N21374);
nor NOR4 (N21377, N21375, N15343, N18344, N9755);
buf BUF1 (N21378, N21370);
xor XOR2 (N21379, N21372, N1823);
xor XOR2 (N21380, N21369, N19351);
or OR3 (N21381, N21380, N3704, N5005);
or OR4 (N21382, N21377, N4720, N14830, N7757);
or OR2 (N21383, N21379, N10146);
nor NOR2 (N21384, N21381, N5069);
or OR2 (N21385, N21384, N9260);
xor XOR2 (N21386, N21350, N3171);
or OR2 (N21387, N21367, N1715);
nand NAND4 (N21388, N21385, N10967, N17179, N12663);
or OR4 (N21389, N21355, N19125, N6868, N11770);
not NOT1 (N21390, N21382);
buf BUF1 (N21391, N21378);
nand NAND3 (N21392, N21391, N10778, N15278);
not NOT1 (N21393, N21388);
buf BUF1 (N21394, N21387);
nand NAND3 (N21395, N21392, N12845, N13610);
nand NAND2 (N21396, N21371, N4875);
nand NAND4 (N21397, N21395, N8450, N20397, N6058);
buf BUF1 (N21398, N21390);
nor NOR3 (N21399, N21347, N13995, N15943);
or OR3 (N21400, N21376, N19379, N4070);
nor NOR3 (N21401, N21389, N20403, N19820);
or OR4 (N21402, N21397, N19962, N21286, N4762);
nor NOR2 (N21403, N21393, N9428);
nand NAND2 (N21404, N21400, N3743);
and AND2 (N21405, N21404, N19396);
buf BUF1 (N21406, N21399);
or OR2 (N21407, N21402, N3234);
xor XOR2 (N21408, N21398, N15293);
or OR3 (N21409, N21403, N7196, N10972);
or OR3 (N21410, N21394, N8585, N6082);
nor NOR4 (N21411, N21405, N16755, N8241, N17502);
and AND2 (N21412, N21383, N2958);
nand NAND4 (N21413, N21412, N2296, N19256, N12065);
xor XOR2 (N21414, N21401, N10438);
buf BUF1 (N21415, N21410);
or OR2 (N21416, N21406, N16083);
buf BUF1 (N21417, N21416);
and AND2 (N21418, N21414, N7277);
or OR4 (N21419, N21411, N4022, N4528, N6211);
and AND3 (N21420, N21418, N822, N16250);
not NOT1 (N21421, N21419);
nand NAND4 (N21422, N21415, N15646, N11422, N21060);
nor NOR2 (N21423, N21417, N17281);
nor NOR3 (N21424, N21408, N6230, N14136);
and AND4 (N21425, N21396, N20992, N14646, N10921);
not NOT1 (N21426, N21425);
xor XOR2 (N21427, N21424, N14749);
buf BUF1 (N21428, N21421);
or OR4 (N21429, N21386, N11523, N3552, N10265);
and AND3 (N21430, N21429, N14041, N16718);
nand NAND4 (N21431, N21428, N15333, N14439, N18754);
xor XOR2 (N21432, N21413, N506);
xor XOR2 (N21433, N21409, N7175);
or OR3 (N21434, N21422, N11370, N9573);
nor NOR3 (N21435, N21433, N10988, N15191);
buf BUF1 (N21436, N21427);
not NOT1 (N21437, N21420);
nand NAND4 (N21438, N21423, N15700, N6306, N7398);
and AND4 (N21439, N21435, N18977, N399, N3376);
xor XOR2 (N21440, N21439, N9442);
nor NOR4 (N21441, N21440, N19626, N14919, N7302);
buf BUF1 (N21442, N21437);
nand NAND2 (N21443, N21442, N20990);
buf BUF1 (N21444, N21438);
xor XOR2 (N21445, N21432, N17616);
buf BUF1 (N21446, N21407);
buf BUF1 (N21447, N21434);
buf BUF1 (N21448, N21431);
and AND3 (N21449, N21441, N15077, N5781);
or OR4 (N21450, N21426, N17521, N6635, N13608);
or OR3 (N21451, N21443, N13408, N12578);
xor XOR2 (N21452, N21430, N2109);
nand NAND3 (N21453, N21446, N106, N5765);
nor NOR4 (N21454, N21436, N8413, N10211, N11911);
xor XOR2 (N21455, N21448, N12146);
nand NAND4 (N21456, N21451, N11177, N4123, N13173);
and AND4 (N21457, N21450, N1969, N11959, N13202);
xor XOR2 (N21458, N21456, N3658);
not NOT1 (N21459, N21449);
or OR4 (N21460, N21447, N17696, N21221, N6433);
nor NOR3 (N21461, N21459, N4167, N1391);
and AND4 (N21462, N21444, N8108, N6391, N10356);
or OR2 (N21463, N21454, N8186);
and AND2 (N21464, N21455, N9418);
and AND3 (N21465, N21460, N13078, N15078);
not NOT1 (N21466, N21458);
xor XOR2 (N21467, N21465, N5095);
xor XOR2 (N21468, N21461, N4411);
and AND4 (N21469, N21463, N4143, N110, N18775);
nand NAND2 (N21470, N21464, N1201);
xor XOR2 (N21471, N21468, N16959);
and AND3 (N21472, N21471, N21233, N2417);
or OR2 (N21473, N21466, N4386);
nand NAND4 (N21474, N21472, N8300, N13981, N19008);
or OR3 (N21475, N21473, N16551, N15608);
or OR4 (N21476, N21467, N15847, N1263, N17931);
nor NOR2 (N21477, N21474, N5417);
xor XOR2 (N21478, N21470, N4372);
nand NAND3 (N21479, N21469, N14313, N9137);
nand NAND4 (N21480, N21477, N11078, N8618, N15913);
or OR4 (N21481, N21445, N2661, N10671, N14326);
nand NAND4 (N21482, N21457, N9531, N6433, N15215);
xor XOR2 (N21483, N21452, N18819);
not NOT1 (N21484, N21479);
buf BUF1 (N21485, N21484);
nand NAND2 (N21486, N21482, N9277);
and AND3 (N21487, N21485, N5706, N20789);
xor XOR2 (N21488, N21480, N9660);
nor NOR4 (N21489, N21476, N322, N14775, N889);
not NOT1 (N21490, N21475);
xor XOR2 (N21491, N21483, N9048);
nor NOR4 (N21492, N21488, N15233, N3109, N17966);
or OR4 (N21493, N21486, N12148, N13512, N8448);
or OR2 (N21494, N21489, N7971);
nand NAND3 (N21495, N21493, N10452, N15704);
and AND2 (N21496, N21487, N17437);
or OR4 (N21497, N21496, N10974, N9030, N11952);
not NOT1 (N21498, N21492);
and AND2 (N21499, N21498, N10360);
xor XOR2 (N21500, N21494, N18593);
nand NAND3 (N21501, N21478, N16114, N19032);
nand NAND3 (N21502, N21481, N18513, N20937);
buf BUF1 (N21503, N21490);
nand NAND2 (N21504, N21495, N3170);
not NOT1 (N21505, N21500);
or OR2 (N21506, N21505, N5282);
not NOT1 (N21507, N21503);
or OR4 (N21508, N21502, N8556, N14316, N11032);
xor XOR2 (N21509, N21453, N5602);
nand NAND4 (N21510, N21499, N17245, N12569, N10016);
or OR4 (N21511, N21497, N1243, N7038, N8091);
nand NAND3 (N21512, N21507, N12668, N5806);
or OR4 (N21513, N21511, N9168, N14749, N819);
not NOT1 (N21514, N21462);
nand NAND4 (N21515, N21501, N6014, N658, N6275);
nor NOR4 (N21516, N21510, N15932, N14831, N7151);
xor XOR2 (N21517, N21509, N11666);
and AND2 (N21518, N21506, N16290);
xor XOR2 (N21519, N21504, N15638);
not NOT1 (N21520, N21518);
nor NOR2 (N21521, N21508, N8878);
buf BUF1 (N21522, N21515);
nor NOR4 (N21523, N21522, N21208, N18327, N19712);
nor NOR4 (N21524, N21514, N13022, N1367, N17853);
and AND3 (N21525, N21521, N15891, N15585);
or OR3 (N21526, N21517, N18702, N420);
nor NOR3 (N21527, N21524, N12353, N14407);
xor XOR2 (N21528, N21491, N6187);
xor XOR2 (N21529, N21520, N13811);
xor XOR2 (N21530, N21526, N5);
nand NAND2 (N21531, N21529, N13698);
not NOT1 (N21532, N21523);
nand NAND3 (N21533, N21531, N7158, N15057);
and AND4 (N21534, N21528, N13527, N8213, N18137);
xor XOR2 (N21535, N21519, N7317);
or OR3 (N21536, N21516, N2967, N1145);
nand NAND2 (N21537, N21527, N13548);
or OR4 (N21538, N21532, N5840, N18211, N14624);
nand NAND3 (N21539, N21534, N9549, N6387);
or OR3 (N21540, N21533, N17684, N20077);
nand NAND4 (N21541, N21530, N9714, N13840, N1111);
nand NAND4 (N21542, N21537, N17328, N10107, N18732);
not NOT1 (N21543, N21540);
or OR4 (N21544, N21536, N17743, N19147, N5855);
nor NOR4 (N21545, N21512, N21263, N3245, N5316);
and AND4 (N21546, N21535, N5982, N3177, N14204);
xor XOR2 (N21547, N21542, N1657);
buf BUF1 (N21548, N21543);
and AND4 (N21549, N21539, N19799, N1578, N9101);
nor NOR3 (N21550, N21544, N13108, N161);
buf BUF1 (N21551, N21550);
buf BUF1 (N21552, N21513);
nand NAND3 (N21553, N21525, N21177, N17748);
nor NOR2 (N21554, N21538, N4517);
nor NOR3 (N21555, N21541, N1745, N9567);
not NOT1 (N21556, N21545);
and AND2 (N21557, N21552, N8249);
nor NOR4 (N21558, N21551, N18609, N1773, N11546);
and AND4 (N21559, N21553, N13566, N10017, N19564);
or OR4 (N21560, N21558, N17756, N15730, N4214);
buf BUF1 (N21561, N21557);
not NOT1 (N21562, N21547);
xor XOR2 (N21563, N21556, N17694);
nor NOR4 (N21564, N21560, N20644, N8225, N19964);
buf BUF1 (N21565, N21563);
not NOT1 (N21566, N21549);
nand NAND3 (N21567, N21566, N15845, N7937);
or OR4 (N21568, N21546, N21511, N19367, N3636);
and AND4 (N21569, N21562, N15798, N11491, N14062);
buf BUF1 (N21570, N21564);
and AND4 (N21571, N21568, N1296, N16788, N10846);
buf BUF1 (N21572, N21565);
or OR4 (N21573, N21572, N7792, N4548, N6293);
and AND3 (N21574, N21573, N20727, N13529);
nor NOR4 (N21575, N21554, N8883, N1584, N14262);
and AND4 (N21576, N21575, N1091, N6258, N2540);
or OR4 (N21577, N21576, N13779, N14497, N17572);
not NOT1 (N21578, N21548);
nand NAND4 (N21579, N21559, N5505, N5553, N17749);
and AND3 (N21580, N21561, N12301, N3701);
or OR4 (N21581, N21574, N3455, N2721, N4259);
buf BUF1 (N21582, N21577);
buf BUF1 (N21583, N21578);
nor NOR2 (N21584, N21570, N1478);
nor NOR3 (N21585, N21581, N3036, N19912);
buf BUF1 (N21586, N21571);
nand NAND2 (N21587, N21582, N15107);
or OR3 (N21588, N21585, N8378, N18222);
and AND3 (N21589, N21579, N10203, N12158);
xor XOR2 (N21590, N21580, N15448);
buf BUF1 (N21591, N21567);
buf BUF1 (N21592, N21555);
xor XOR2 (N21593, N21587, N442);
xor XOR2 (N21594, N21593, N14231);
and AND4 (N21595, N21588, N13053, N17155, N1423);
nor NOR3 (N21596, N21595, N20116, N19926);
not NOT1 (N21597, N21592);
xor XOR2 (N21598, N21583, N10672);
xor XOR2 (N21599, N21598, N10668);
or OR3 (N21600, N21586, N471, N12149);
buf BUF1 (N21601, N21589);
nand NAND2 (N21602, N21599, N7998);
not NOT1 (N21603, N21584);
and AND2 (N21604, N21596, N12982);
nand NAND2 (N21605, N21569, N6536);
xor XOR2 (N21606, N21601, N7060);
xor XOR2 (N21607, N21597, N4047);
nand NAND3 (N21608, N21602, N8915, N14725);
and AND2 (N21609, N21608, N21535);
or OR4 (N21610, N21594, N7329, N11618, N14279);
or OR4 (N21611, N21607, N16684, N5067, N1298);
and AND3 (N21612, N21609, N15451, N19372);
buf BUF1 (N21613, N21590);
not NOT1 (N21614, N21600);
or OR2 (N21615, N21611, N11940);
not NOT1 (N21616, N21591);
not NOT1 (N21617, N21616);
nor NOR3 (N21618, N21613, N8098, N9154);
or OR3 (N21619, N21612, N19754, N2214);
nor NOR4 (N21620, N21614, N2562, N11781, N7007);
or OR3 (N21621, N21618, N14381, N20810);
nor NOR2 (N21622, N21621, N13220);
and AND2 (N21623, N21606, N6712);
nand NAND2 (N21624, N21604, N9934);
nand NAND3 (N21625, N21603, N1646, N4973);
buf BUF1 (N21626, N21624);
nand NAND3 (N21627, N21623, N5041, N15983);
not NOT1 (N21628, N21619);
nand NAND2 (N21629, N21625, N17358);
nor NOR3 (N21630, N21615, N10324, N1153);
nor NOR4 (N21631, N21617, N15994, N11010, N19496);
xor XOR2 (N21632, N21605, N1270);
nor NOR2 (N21633, N21630, N4628);
buf BUF1 (N21634, N21628);
nor NOR4 (N21635, N21634, N11693, N11977, N7940);
or OR4 (N21636, N21633, N1543, N5841, N1381);
or OR4 (N21637, N21626, N20016, N16951, N16644);
and AND2 (N21638, N21635, N13405);
not NOT1 (N21639, N21632);
not NOT1 (N21640, N21638);
or OR2 (N21641, N21640, N11086);
not NOT1 (N21642, N21610);
xor XOR2 (N21643, N21629, N12974);
xor XOR2 (N21644, N21622, N18577);
xor XOR2 (N21645, N21643, N21253);
buf BUF1 (N21646, N21644);
buf BUF1 (N21647, N21637);
or OR4 (N21648, N21645, N12626, N1267, N18257);
nor NOR3 (N21649, N21636, N4894, N7196);
xor XOR2 (N21650, N21642, N9330);
nand NAND2 (N21651, N21641, N6957);
and AND4 (N21652, N21646, N20570, N1362, N7421);
and AND3 (N21653, N21647, N3320, N1119);
nand NAND2 (N21654, N21639, N13120);
xor XOR2 (N21655, N21620, N1327);
buf BUF1 (N21656, N21650);
buf BUF1 (N21657, N21631);
buf BUF1 (N21658, N21654);
xor XOR2 (N21659, N21653, N10208);
buf BUF1 (N21660, N21657);
xor XOR2 (N21661, N21658, N5965);
nor NOR2 (N21662, N21656, N1234);
or OR2 (N21663, N21627, N5330);
xor XOR2 (N21664, N21655, N8850);
or OR4 (N21665, N21659, N11126, N14035, N20783);
nor NOR3 (N21666, N21660, N15127, N21598);
nand NAND2 (N21667, N21649, N18557);
nand NAND3 (N21668, N21648, N14863, N5835);
or OR2 (N21669, N21665, N1060);
xor XOR2 (N21670, N21652, N8755);
nand NAND2 (N21671, N21664, N19099);
or OR3 (N21672, N21666, N21497, N12493);
nor NOR3 (N21673, N21663, N10624, N12684);
and AND3 (N21674, N21670, N9231, N14455);
buf BUF1 (N21675, N21671);
and AND2 (N21676, N21661, N849);
not NOT1 (N21677, N21669);
or OR4 (N21678, N21676, N8675, N17394, N11605);
nand NAND4 (N21679, N21674, N15766, N9829, N14696);
not NOT1 (N21680, N21677);
not NOT1 (N21681, N21667);
nor NOR2 (N21682, N21681, N5674);
nor NOR2 (N21683, N21673, N14429);
or OR2 (N21684, N21680, N20764);
nor NOR3 (N21685, N21682, N3475, N8125);
buf BUF1 (N21686, N21672);
not NOT1 (N21687, N21651);
buf BUF1 (N21688, N21662);
buf BUF1 (N21689, N21684);
nor NOR4 (N21690, N21688, N2914, N20134, N7834);
buf BUF1 (N21691, N21679);
buf BUF1 (N21692, N21675);
and AND2 (N21693, N21687, N7733);
nor NOR4 (N21694, N21692, N20725, N8276, N14368);
and AND4 (N21695, N21668, N16890, N5934, N8364);
or OR2 (N21696, N21693, N10968);
buf BUF1 (N21697, N21685);
not NOT1 (N21698, N21686);
and AND2 (N21699, N21690, N11412);
buf BUF1 (N21700, N21697);
or OR3 (N21701, N21678, N3075, N5433);
not NOT1 (N21702, N21689);
not NOT1 (N21703, N21694);
nor NOR4 (N21704, N21683, N20714, N15269, N3202);
nor NOR3 (N21705, N21698, N4780, N19270);
nor NOR3 (N21706, N21702, N11886, N2643);
nor NOR3 (N21707, N21705, N311, N12057);
nand NAND3 (N21708, N21707, N1276, N19972);
nor NOR2 (N21709, N21695, N603);
and AND3 (N21710, N21708, N7230, N556);
or OR2 (N21711, N21703, N10429);
or OR2 (N21712, N21701, N16291);
and AND3 (N21713, N21711, N3109, N755);
nor NOR3 (N21714, N21712, N19946, N5780);
or OR4 (N21715, N21713, N7403, N12549, N12843);
not NOT1 (N21716, N21704);
not NOT1 (N21717, N21715);
nor NOR4 (N21718, N21696, N19780, N8253, N19448);
and AND3 (N21719, N21699, N19665, N5450);
buf BUF1 (N21720, N21717);
or OR3 (N21721, N21716, N5997, N8009);
not NOT1 (N21722, N21691);
and AND4 (N21723, N21719, N4558, N14493, N19027);
and AND2 (N21724, N21714, N3873);
not NOT1 (N21725, N21722);
xor XOR2 (N21726, N21700, N11454);
nor NOR4 (N21727, N21724, N14386, N16903, N11846);
or OR4 (N21728, N21706, N8477, N6440, N19499);
not NOT1 (N21729, N21720);
nor NOR2 (N21730, N21725, N6198);
nand NAND3 (N21731, N21728, N10005, N11471);
buf BUF1 (N21732, N21718);
xor XOR2 (N21733, N21731, N13496);
xor XOR2 (N21734, N21727, N5627);
and AND4 (N21735, N21710, N19624, N18811, N9617);
nand NAND3 (N21736, N21733, N6554, N17496);
not NOT1 (N21737, N21734);
or OR2 (N21738, N21736, N21226);
or OR4 (N21739, N21726, N6684, N4431, N8552);
nand NAND4 (N21740, N21735, N17609, N1010, N19143);
xor XOR2 (N21741, N21739, N18629);
and AND4 (N21742, N21740, N9941, N15718, N13701);
buf BUF1 (N21743, N21732);
nor NOR4 (N21744, N21730, N21515, N15357, N4681);
nand NAND2 (N21745, N21723, N14813);
buf BUF1 (N21746, N21745);
nand NAND4 (N21747, N21741, N1016, N12545, N18437);
not NOT1 (N21748, N21747);
or OR4 (N21749, N21744, N19742, N10017, N16580);
and AND2 (N21750, N21746, N10522);
and AND4 (N21751, N21743, N28, N7612, N6210);
nand NAND4 (N21752, N21738, N18854, N19976, N14061);
not NOT1 (N21753, N21749);
or OR4 (N21754, N21753, N9858, N16737, N8175);
xor XOR2 (N21755, N21729, N7665);
not NOT1 (N21756, N21721);
nor NOR2 (N21757, N21752, N16790);
xor XOR2 (N21758, N21748, N19240);
xor XOR2 (N21759, N21756, N1585);
buf BUF1 (N21760, N21709);
xor XOR2 (N21761, N21754, N20853);
buf BUF1 (N21762, N21751);
nor NOR3 (N21763, N21755, N17774, N6429);
nor NOR4 (N21764, N21758, N3695, N15526, N16962);
not NOT1 (N21765, N21742);
nand NAND3 (N21766, N21760, N17272, N2049);
and AND3 (N21767, N21737, N1279, N7824);
and AND4 (N21768, N21762, N14756, N8608, N18743);
and AND4 (N21769, N21763, N13168, N2890, N1130);
nor NOR4 (N21770, N21766, N20418, N2999, N20381);
not NOT1 (N21771, N21770);
buf BUF1 (N21772, N21765);
and AND3 (N21773, N21771, N11528, N3526);
nor NOR4 (N21774, N21769, N16533, N18549, N14268);
xor XOR2 (N21775, N21759, N14276);
nand NAND2 (N21776, N21768, N10600);
nor NOR4 (N21777, N21767, N9364, N6143, N11891);
nor NOR4 (N21778, N21764, N10700, N919, N12491);
and AND2 (N21779, N21774, N19909);
nor NOR3 (N21780, N21761, N8746, N4273);
nor NOR2 (N21781, N21772, N3537);
nor NOR3 (N21782, N21777, N7261, N11036);
and AND2 (N21783, N21775, N5570);
or OR3 (N21784, N21776, N13045, N13324);
nor NOR4 (N21785, N21784, N10860, N6344, N12011);
xor XOR2 (N21786, N21750, N1855);
nand NAND4 (N21787, N21773, N13385, N10896, N13441);
and AND3 (N21788, N21785, N18967, N109);
or OR4 (N21789, N21778, N19806, N12549, N15707);
nand NAND4 (N21790, N21779, N9708, N17718, N21454);
or OR3 (N21791, N21781, N3599, N9437);
nand NAND3 (N21792, N21789, N5185, N4076);
nand NAND4 (N21793, N21791, N18851, N20986, N8559);
not NOT1 (N21794, N21783);
xor XOR2 (N21795, N21782, N6937);
buf BUF1 (N21796, N21786);
or OR2 (N21797, N21788, N6938);
or OR2 (N21798, N21792, N20563);
xor XOR2 (N21799, N21798, N7504);
or OR4 (N21800, N21794, N15292, N19182, N15647);
nor NOR4 (N21801, N21787, N6600, N6917, N16233);
nor NOR2 (N21802, N21801, N5980);
nor NOR4 (N21803, N21796, N15832, N20361, N17380);
and AND4 (N21804, N21803, N18908, N10721, N2444);
or OR4 (N21805, N21757, N20607, N12162, N15862);
buf BUF1 (N21806, N21790);
nand NAND4 (N21807, N21802, N5587, N17681, N11961);
or OR4 (N21808, N21797, N15314, N3462, N1973);
nand NAND4 (N21809, N21793, N3586, N16674, N18733);
nand NAND3 (N21810, N21808, N6265, N18204);
nor NOR4 (N21811, N21809, N20051, N15658, N4129);
xor XOR2 (N21812, N21795, N17666);
nor NOR2 (N21813, N21807, N3824);
nor NOR4 (N21814, N21805, N3634, N13636, N17950);
xor XOR2 (N21815, N21814, N20603);
buf BUF1 (N21816, N21806);
nand NAND4 (N21817, N21800, N17668, N4169, N12179);
nor NOR4 (N21818, N21815, N15984, N18991, N20403);
xor XOR2 (N21819, N21799, N8306);
xor XOR2 (N21820, N21819, N16629);
or OR4 (N21821, N21820, N16256, N3964, N13029);
or OR2 (N21822, N21804, N19010);
buf BUF1 (N21823, N21816);
buf BUF1 (N21824, N21818);
nand NAND3 (N21825, N21821, N8990, N5286);
nor NOR3 (N21826, N21823, N13725, N10495);
and AND3 (N21827, N21817, N1972, N21154);
or OR2 (N21828, N21812, N21527);
or OR2 (N21829, N21822, N7279);
and AND3 (N21830, N21824, N13968, N10208);
xor XOR2 (N21831, N21829, N4021);
nand NAND4 (N21832, N21811, N5681, N4169, N13820);
not NOT1 (N21833, N21827);
buf BUF1 (N21834, N21813);
not NOT1 (N21835, N21825);
not NOT1 (N21836, N21826);
buf BUF1 (N21837, N21830);
nor NOR2 (N21838, N21837, N10912);
xor XOR2 (N21839, N21834, N9664);
or OR3 (N21840, N21838, N2848, N11659);
buf BUF1 (N21841, N21839);
nand NAND2 (N21842, N21836, N18370);
not NOT1 (N21843, N21833);
nand NAND3 (N21844, N21835, N653, N17353);
and AND4 (N21845, N21831, N20837, N15154, N9635);
or OR3 (N21846, N21841, N14314, N10257);
and AND2 (N21847, N21846, N17028);
not NOT1 (N21848, N21842);
nor NOR3 (N21849, N21832, N20771, N4412);
nor NOR4 (N21850, N21844, N18776, N9587, N13558);
nand NAND2 (N21851, N21849, N6016);
xor XOR2 (N21852, N21828, N7435);
buf BUF1 (N21853, N21851);
nor NOR4 (N21854, N21850, N19449, N9849, N11905);
not NOT1 (N21855, N21843);
buf BUF1 (N21856, N21852);
not NOT1 (N21857, N21854);
and AND4 (N21858, N21810, N10068, N5608, N1031);
nor NOR4 (N21859, N21858, N2668, N12398, N21722);
not NOT1 (N21860, N21855);
and AND4 (N21861, N21840, N17980, N3663, N12229);
and AND3 (N21862, N21860, N2283, N2026);
buf BUF1 (N21863, N21848);
or OR3 (N21864, N21856, N19938, N8708);
and AND2 (N21865, N21859, N8819);
and AND2 (N21866, N21863, N2621);
and AND4 (N21867, N21847, N2435, N2760, N9265);
buf BUF1 (N21868, N21864);
xor XOR2 (N21869, N21868, N10020);
xor XOR2 (N21870, N21867, N17921);
not NOT1 (N21871, N21869);
nor NOR2 (N21872, N21865, N21044);
xor XOR2 (N21873, N21853, N14468);
nand NAND3 (N21874, N21870, N9384, N19786);
or OR3 (N21875, N21874, N13592, N18193);
or OR2 (N21876, N21873, N17988);
not NOT1 (N21877, N21875);
nor NOR3 (N21878, N21861, N9902, N11457);
nor NOR2 (N21879, N21878, N1125);
and AND4 (N21880, N21871, N4169, N21072, N4603);
not NOT1 (N21881, N21872);
nor NOR4 (N21882, N21862, N5375, N15138, N9522);
or OR4 (N21883, N21881, N11718, N14109, N6098);
xor XOR2 (N21884, N21857, N20537);
not NOT1 (N21885, N21877);
xor XOR2 (N21886, N21885, N6237);
xor XOR2 (N21887, N21780, N15297);
nor NOR2 (N21888, N21886, N10449);
nor NOR3 (N21889, N21887, N16343, N14079);
not NOT1 (N21890, N21884);
and AND2 (N21891, N21879, N2413);
and AND4 (N21892, N21866, N20045, N5990, N5683);
or OR2 (N21893, N21883, N5789);
or OR4 (N21894, N21889, N477, N18778, N16237);
buf BUF1 (N21895, N21882);
nand NAND2 (N21896, N21895, N13613);
or OR4 (N21897, N21890, N14590, N11984, N12635);
and AND4 (N21898, N21845, N15901, N6921, N14950);
and AND3 (N21899, N21880, N15497, N1831);
or OR3 (N21900, N21891, N4991, N19810);
xor XOR2 (N21901, N21899, N21606);
not NOT1 (N21902, N21893);
xor XOR2 (N21903, N21896, N1121);
or OR4 (N21904, N21901, N11975, N13222, N16181);
and AND4 (N21905, N21894, N9482, N3325, N15109);
buf BUF1 (N21906, N21900);
buf BUF1 (N21907, N21903);
buf BUF1 (N21908, N21898);
buf BUF1 (N21909, N21902);
buf BUF1 (N21910, N21905);
buf BUF1 (N21911, N21907);
buf BUF1 (N21912, N21911);
not NOT1 (N21913, N21912);
and AND3 (N21914, N21910, N9718, N8946);
or OR3 (N21915, N21913, N21616, N21449);
nand NAND4 (N21916, N21904, N16717, N873, N8298);
or OR2 (N21917, N21916, N6183);
or OR4 (N21918, N21908, N13860, N8108, N12732);
xor XOR2 (N21919, N21915, N822);
xor XOR2 (N21920, N21909, N10240);
nand NAND2 (N21921, N21892, N2253);
buf BUF1 (N21922, N21921);
not NOT1 (N21923, N21876);
nor NOR2 (N21924, N21922, N5714);
or OR4 (N21925, N21897, N15348, N17769, N21283);
nor NOR3 (N21926, N21888, N17568, N12687);
not NOT1 (N21927, N21914);
or OR2 (N21928, N21920, N7345);
xor XOR2 (N21929, N21927, N8768);
nand NAND2 (N21930, N21924, N14334);
or OR3 (N21931, N21926, N9307, N13621);
nor NOR3 (N21932, N21929, N9489, N9371);
and AND4 (N21933, N21906, N7949, N12837, N12709);
xor XOR2 (N21934, N21923, N19586);
or OR3 (N21935, N21932, N7278, N11593);
or OR3 (N21936, N21933, N16127, N7809);
and AND3 (N21937, N21934, N16198, N19063);
nor NOR2 (N21938, N21918, N1067);
xor XOR2 (N21939, N21925, N21119);
not NOT1 (N21940, N21930);
xor XOR2 (N21941, N21917, N13619);
or OR3 (N21942, N21928, N249, N4538);
or OR3 (N21943, N21939, N2176, N13966);
not NOT1 (N21944, N21935);
xor XOR2 (N21945, N21936, N14663);
xor XOR2 (N21946, N21937, N2686);
nor NOR2 (N21947, N21941, N8390);
xor XOR2 (N21948, N21940, N9031);
nor NOR4 (N21949, N21944, N16272, N1976, N12035);
not NOT1 (N21950, N21942);
not NOT1 (N21951, N21947);
nand NAND4 (N21952, N21951, N20053, N13049, N372);
nor NOR4 (N21953, N21952, N13229, N1705, N8571);
and AND2 (N21954, N21945, N12117);
nor NOR2 (N21955, N21949, N11381);
nor NOR2 (N21956, N21954, N728);
not NOT1 (N21957, N21943);
not NOT1 (N21958, N21931);
buf BUF1 (N21959, N21956);
nand NAND3 (N21960, N21958, N9765, N13505);
buf BUF1 (N21961, N21960);
buf BUF1 (N21962, N21957);
not NOT1 (N21963, N21950);
not NOT1 (N21964, N21962);
xor XOR2 (N21965, N21938, N10839);
buf BUF1 (N21966, N21955);
not NOT1 (N21967, N21959);
xor XOR2 (N21968, N21946, N14775);
buf BUF1 (N21969, N21964);
and AND4 (N21970, N21968, N10052, N8316, N8535);
nor NOR4 (N21971, N21966, N2302, N9604, N1053);
nand NAND3 (N21972, N21969, N17386, N5783);
or OR3 (N21973, N21971, N18914, N3414);
not NOT1 (N21974, N21967);
or OR2 (N21975, N21948, N20602);
buf BUF1 (N21976, N21972);
xor XOR2 (N21977, N21970, N1148);
xor XOR2 (N21978, N21953, N10004);
buf BUF1 (N21979, N21974);
and AND3 (N21980, N21976, N907, N10076);
buf BUF1 (N21981, N21965);
xor XOR2 (N21982, N21980, N20558);
not NOT1 (N21983, N21978);
or OR2 (N21984, N21975, N17697);
nand NAND3 (N21985, N21977, N13769, N3551);
buf BUF1 (N21986, N21985);
or OR4 (N21987, N21981, N4868, N16435, N20010);
not NOT1 (N21988, N21982);
not NOT1 (N21989, N21973);
not NOT1 (N21990, N21986);
xor XOR2 (N21991, N21983, N332);
buf BUF1 (N21992, N21963);
xor XOR2 (N21993, N21989, N11260);
nor NOR3 (N21994, N21993, N2754, N795);
xor XOR2 (N21995, N21979, N17820);
not NOT1 (N21996, N21990);
nor NOR4 (N21997, N21984, N10807, N6436, N19965);
buf BUF1 (N21998, N21987);
and AND4 (N21999, N21961, N5377, N2334, N10683);
not NOT1 (N22000, N21991);
xor XOR2 (N22001, N21997, N15666);
nand NAND2 (N22002, N21919, N2120);
buf BUF1 (N22003, N21998);
xor XOR2 (N22004, N22002, N7504);
buf BUF1 (N22005, N21994);
or OR3 (N22006, N22003, N17146, N12888);
not NOT1 (N22007, N22006);
or OR3 (N22008, N21999, N5759, N4257);
not NOT1 (N22009, N22000);
buf BUF1 (N22010, N22005);
not NOT1 (N22011, N22008);
buf BUF1 (N22012, N22004);
and AND3 (N22013, N22010, N8503, N5184);
or OR2 (N22014, N21992, N15057);
nor NOR2 (N22015, N22014, N1476);
not NOT1 (N22016, N22009);
buf BUF1 (N22017, N21995);
nor NOR4 (N22018, N21988, N15102, N3527, N5560);
nand NAND3 (N22019, N22018, N4390, N7734);
xor XOR2 (N22020, N22011, N15979);
nor NOR3 (N22021, N22012, N1968, N1810);
nand NAND3 (N22022, N22013, N6551, N15341);
or OR4 (N22023, N22019, N12279, N3673, N4664);
xor XOR2 (N22024, N22016, N17030);
xor XOR2 (N22025, N22001, N3540);
nor NOR4 (N22026, N21996, N11979, N4202, N5645);
nor NOR4 (N22027, N22026, N17249, N4080, N11476);
buf BUF1 (N22028, N22023);
xor XOR2 (N22029, N22024, N17837);
or OR4 (N22030, N22007, N1240, N21350, N3304);
or OR4 (N22031, N22028, N12569, N2949, N9095);
or OR2 (N22032, N22015, N5701);
nor NOR4 (N22033, N22029, N5922, N13882, N3703);
buf BUF1 (N22034, N22030);
or OR3 (N22035, N22022, N18980, N15141);
or OR2 (N22036, N22027, N21910);
not NOT1 (N22037, N22025);
not NOT1 (N22038, N22033);
not NOT1 (N22039, N22021);
not NOT1 (N22040, N22031);
xor XOR2 (N22041, N22038, N4559);
or OR3 (N22042, N22035, N13230, N15357);
nor NOR4 (N22043, N22032, N15201, N10835, N19986);
nor NOR3 (N22044, N22017, N14483, N4383);
nand NAND2 (N22045, N22043, N11165);
or OR3 (N22046, N22041, N10002, N18900);
or OR4 (N22047, N22036, N16268, N21369, N13485);
or OR4 (N22048, N22044, N7375, N14465, N4806);
or OR4 (N22049, N22034, N3239, N16968, N21211);
not NOT1 (N22050, N22048);
nand NAND3 (N22051, N22050, N8466, N5221);
xor XOR2 (N22052, N22051, N19634);
or OR4 (N22053, N22047, N13215, N4613, N7546);
nand NAND4 (N22054, N22042, N7482, N17390, N17806);
not NOT1 (N22055, N22046);
nor NOR4 (N22056, N22045, N18635, N3867, N14336);
and AND3 (N22057, N22037, N1034, N20709);
not NOT1 (N22058, N22049);
not NOT1 (N22059, N22052);
and AND3 (N22060, N22054, N10908, N7626);
xor XOR2 (N22061, N22055, N12101);
nor NOR2 (N22062, N22059, N5248);
nand NAND3 (N22063, N22062, N21057, N17991);
or OR3 (N22064, N22063, N10058, N1538);
nand NAND2 (N22065, N22039, N6171);
and AND3 (N22066, N22060, N16719, N140);
buf BUF1 (N22067, N22058);
not NOT1 (N22068, N22057);
or OR4 (N22069, N22065, N4721, N8327, N9240);
xor XOR2 (N22070, N22069, N15762);
nor NOR2 (N22071, N22070, N834);
not NOT1 (N22072, N22068);
nand NAND3 (N22073, N22071, N10043, N21595);
buf BUF1 (N22074, N22064);
not NOT1 (N22075, N22074);
buf BUF1 (N22076, N22075);
and AND2 (N22077, N22066, N9422);
xor XOR2 (N22078, N22061, N16028);
buf BUF1 (N22079, N22040);
xor XOR2 (N22080, N22073, N13476);
xor XOR2 (N22081, N22056, N17104);
not NOT1 (N22082, N22081);
nor NOR4 (N22083, N22078, N13362, N17696, N8909);
and AND4 (N22084, N22053, N7970, N15066, N19559);
nor NOR3 (N22085, N22083, N1680, N18542);
and AND4 (N22086, N22085, N8672, N5701, N3547);
or OR2 (N22087, N22084, N10481);
nor NOR2 (N22088, N22076, N19229);
xor XOR2 (N22089, N22088, N21054);
and AND4 (N22090, N22087, N762, N8766, N14031);
nand NAND3 (N22091, N22079, N5236, N13031);
nor NOR4 (N22092, N22080, N17452, N703, N19950);
buf BUF1 (N22093, N22020);
not NOT1 (N22094, N22072);
nor NOR4 (N22095, N22082, N637, N13164, N12988);
xor XOR2 (N22096, N22092, N21645);
buf BUF1 (N22097, N22095);
nand NAND4 (N22098, N22090, N10642, N13968, N7353);
and AND3 (N22099, N22091, N5024, N3314);
buf BUF1 (N22100, N22098);
and AND4 (N22101, N22096, N9026, N7101, N17397);
nor NOR2 (N22102, N22086, N13787);
or OR4 (N22103, N22101, N3611, N21850, N7572);
nor NOR2 (N22104, N22102, N18878);
or OR2 (N22105, N22103, N15632);
nor NOR4 (N22106, N22067, N236, N12731, N14270);
not NOT1 (N22107, N22097);
or OR2 (N22108, N22093, N15401);
buf BUF1 (N22109, N22099);
not NOT1 (N22110, N22077);
not NOT1 (N22111, N22104);
or OR4 (N22112, N22106, N382, N12647, N16965);
buf BUF1 (N22113, N22110);
and AND2 (N22114, N22094, N3537);
nand NAND3 (N22115, N22112, N14594, N7565);
buf BUF1 (N22116, N22111);
not NOT1 (N22117, N22089);
buf BUF1 (N22118, N22100);
xor XOR2 (N22119, N22117, N22072);
buf BUF1 (N22120, N22108);
and AND2 (N22121, N22107, N8681);
not NOT1 (N22122, N22109);
or OR2 (N22123, N22114, N19344);
not NOT1 (N22124, N22116);
xor XOR2 (N22125, N22120, N16958);
not NOT1 (N22126, N22119);
or OR2 (N22127, N22118, N3968);
and AND2 (N22128, N22115, N5641);
nor NOR4 (N22129, N22123, N1459, N1567, N529);
and AND4 (N22130, N22126, N14689, N9645, N19844);
or OR2 (N22131, N22105, N17232);
and AND3 (N22132, N22113, N10819, N439);
buf BUF1 (N22133, N22130);
nand NAND2 (N22134, N22125, N9850);
nor NOR3 (N22135, N22133, N8640, N14498);
not NOT1 (N22136, N22124);
and AND2 (N22137, N22127, N18789);
not NOT1 (N22138, N22128);
nand NAND2 (N22139, N22135, N16096);
or OR3 (N22140, N22139, N11692, N15685);
and AND2 (N22141, N22131, N16119);
buf BUF1 (N22142, N22122);
nand NAND4 (N22143, N22129, N16121, N8780, N19977);
buf BUF1 (N22144, N22132);
or OR4 (N22145, N22138, N13815, N4861, N4579);
buf BUF1 (N22146, N22121);
nor NOR3 (N22147, N22146, N8016, N20297);
and AND2 (N22148, N22145, N12084);
nor NOR2 (N22149, N22143, N14143);
and AND4 (N22150, N22148, N3920, N18930, N3297);
nor NOR4 (N22151, N22140, N19222, N9369, N7640);
nand NAND3 (N22152, N22150, N10375, N17639);
nor NOR4 (N22153, N22136, N402, N18002, N2400);
and AND2 (N22154, N22144, N10742);
xor XOR2 (N22155, N22149, N4832);
nor NOR4 (N22156, N22134, N204, N21477, N21628);
xor XOR2 (N22157, N22155, N561);
nand NAND2 (N22158, N22137, N18985);
buf BUF1 (N22159, N22153);
xor XOR2 (N22160, N22154, N7507);
and AND2 (N22161, N22158, N19156);
not NOT1 (N22162, N22147);
buf BUF1 (N22163, N22151);
nand NAND2 (N22164, N22157, N14680);
buf BUF1 (N22165, N22161);
not NOT1 (N22166, N22156);
and AND3 (N22167, N22166, N13379, N17246);
xor XOR2 (N22168, N22165, N2163);
buf BUF1 (N22169, N22164);
xor XOR2 (N22170, N22152, N12121);
nand NAND4 (N22171, N22167, N13107, N19326, N17834);
xor XOR2 (N22172, N22168, N18924);
not NOT1 (N22173, N22160);
or OR3 (N22174, N22141, N16100, N6335);
or OR4 (N22175, N22159, N18703, N6177, N1062);
buf BUF1 (N22176, N22172);
nand NAND4 (N22177, N22170, N4273, N2427, N3979);
not NOT1 (N22178, N22162);
xor XOR2 (N22179, N22177, N5970);
buf BUF1 (N22180, N22179);
nand NAND2 (N22181, N22178, N8441);
xor XOR2 (N22182, N22169, N9779);
buf BUF1 (N22183, N22176);
nand NAND3 (N22184, N22142, N8239, N15208);
nand NAND3 (N22185, N22182, N8591, N17664);
not NOT1 (N22186, N22175);
nand NAND2 (N22187, N22185, N5196);
nor NOR3 (N22188, N22163, N18704, N367);
and AND3 (N22189, N22180, N14672, N6437);
nand NAND4 (N22190, N22181, N1042, N13884, N20150);
xor XOR2 (N22191, N22186, N574);
nor NOR3 (N22192, N22174, N21696, N19170);
not NOT1 (N22193, N22183);
not NOT1 (N22194, N22187);
xor XOR2 (N22195, N22192, N8888);
nand NAND4 (N22196, N22190, N2252, N8653, N18303);
xor XOR2 (N22197, N22194, N5702);
nand NAND3 (N22198, N22184, N20186, N10876);
not NOT1 (N22199, N22195);
not NOT1 (N22200, N22188);
not NOT1 (N22201, N22173);
not NOT1 (N22202, N22171);
nor NOR3 (N22203, N22198, N1981, N6860);
xor XOR2 (N22204, N22201, N6146);
buf BUF1 (N22205, N22199);
nor NOR2 (N22206, N22191, N4122);
not NOT1 (N22207, N22205);
and AND2 (N22208, N22202, N8358);
not NOT1 (N22209, N22189);
or OR3 (N22210, N22200, N7850, N16106);
and AND4 (N22211, N22197, N12507, N6182, N6364);
not NOT1 (N22212, N22193);
and AND3 (N22213, N22204, N17736, N16524);
not NOT1 (N22214, N22206);
buf BUF1 (N22215, N22203);
xor XOR2 (N22216, N22212, N15779);
buf BUF1 (N22217, N22215);
or OR4 (N22218, N22209, N4910, N9084, N10985);
nor NOR4 (N22219, N22210, N9596, N3615, N19256);
not NOT1 (N22220, N22216);
and AND4 (N22221, N22219, N7860, N770, N11263);
nand NAND4 (N22222, N22196, N3222, N7831, N5820);
buf BUF1 (N22223, N22221);
nor NOR3 (N22224, N22220, N20366, N1173);
nor NOR4 (N22225, N22222, N10335, N14253, N20483);
buf BUF1 (N22226, N22207);
or OR4 (N22227, N22214, N7978, N21210, N19163);
buf BUF1 (N22228, N22224);
nor NOR2 (N22229, N22211, N14077);
buf BUF1 (N22230, N22218);
nand NAND4 (N22231, N22225, N11573, N21584, N7386);
nand NAND2 (N22232, N22231, N13057);
nor NOR4 (N22233, N22232, N20100, N2718, N19273);
nor NOR2 (N22234, N22227, N8355);
nand NAND2 (N22235, N22230, N13944);
buf BUF1 (N22236, N22226);
buf BUF1 (N22237, N22233);
nand NAND2 (N22238, N22217, N8986);
and AND3 (N22239, N22229, N402, N902);
not NOT1 (N22240, N22237);
nand NAND4 (N22241, N22238, N19148, N20669, N4514);
nor NOR2 (N22242, N22228, N7504);
nor NOR3 (N22243, N22235, N13078, N642);
or OR4 (N22244, N22243, N12520, N13722, N14920);
xor XOR2 (N22245, N22208, N5515);
or OR3 (N22246, N22241, N15240, N10787);
or OR4 (N22247, N22236, N20469, N9251, N1285);
buf BUF1 (N22248, N22247);
buf BUF1 (N22249, N22246);
not NOT1 (N22250, N22234);
buf BUF1 (N22251, N22239);
not NOT1 (N22252, N22244);
and AND4 (N22253, N22250, N14790, N2826, N2878);
or OR4 (N22254, N22242, N21112, N9274, N461);
and AND3 (N22255, N22252, N17085, N5923);
not NOT1 (N22256, N22254);
nand NAND4 (N22257, N22223, N3888, N6159, N15428);
xor XOR2 (N22258, N22257, N21827);
and AND4 (N22259, N22249, N6049, N17138, N7201);
and AND4 (N22260, N22248, N14793, N14517, N7724);
nand NAND3 (N22261, N22245, N299, N3351);
not NOT1 (N22262, N22255);
not NOT1 (N22263, N22213);
or OR3 (N22264, N22258, N16877, N1832);
xor XOR2 (N22265, N22259, N19818);
xor XOR2 (N22266, N22260, N5907);
not NOT1 (N22267, N22266);
or OR2 (N22268, N22263, N16487);
or OR2 (N22269, N22265, N18701);
nand NAND2 (N22270, N22253, N18446);
buf BUF1 (N22271, N22256);
buf BUF1 (N22272, N22261);
nor NOR2 (N22273, N22271, N15374);
not NOT1 (N22274, N22273);
and AND4 (N22275, N22269, N1445, N22024, N4486);
xor XOR2 (N22276, N22267, N3246);
and AND3 (N22277, N22268, N20851, N20638);
nor NOR3 (N22278, N22264, N10510, N9387);
xor XOR2 (N22279, N22270, N15057);
and AND2 (N22280, N22279, N3375);
xor XOR2 (N22281, N22274, N2575);
nand NAND2 (N22282, N22276, N2627);
or OR4 (N22283, N22275, N13050, N8067, N1613);
nand NAND4 (N22284, N22278, N18757, N3686, N5265);
not NOT1 (N22285, N22283);
not NOT1 (N22286, N22280);
nand NAND4 (N22287, N22281, N21889, N15881, N5564);
xor XOR2 (N22288, N22251, N1308);
or OR2 (N22289, N22286, N6152);
nor NOR3 (N22290, N22287, N2729, N17322);
nand NAND2 (N22291, N22282, N2223);
or OR3 (N22292, N22288, N1375, N13341);
not NOT1 (N22293, N22277);
and AND3 (N22294, N22289, N12857, N4484);
and AND4 (N22295, N22291, N13524, N225, N5467);
and AND4 (N22296, N22293, N14386, N2061, N7984);
and AND3 (N22297, N22296, N11937, N15901);
not NOT1 (N22298, N22272);
or OR3 (N22299, N22262, N6183, N21793);
xor XOR2 (N22300, N22294, N18648);
or OR3 (N22301, N22298, N15745, N18139);
and AND3 (N22302, N22300, N518, N5819);
buf BUF1 (N22303, N22292);
buf BUF1 (N22304, N22240);
not NOT1 (N22305, N22301);
buf BUF1 (N22306, N22302);
buf BUF1 (N22307, N22299);
and AND2 (N22308, N22307, N10466);
xor XOR2 (N22309, N22306, N10597);
and AND2 (N22310, N22297, N8043);
nor NOR2 (N22311, N22308, N7545);
nand NAND2 (N22312, N22305, N15966);
nor NOR3 (N22313, N22310, N15326, N18291);
not NOT1 (N22314, N22309);
xor XOR2 (N22315, N22303, N2504);
nand NAND4 (N22316, N22313, N15354, N5294, N16817);
nand NAND4 (N22317, N22311, N8084, N7196, N16010);
not NOT1 (N22318, N22317);
and AND4 (N22319, N22285, N8614, N10420, N4422);
not NOT1 (N22320, N22312);
xor XOR2 (N22321, N22295, N18553);
and AND2 (N22322, N22290, N8810);
or OR4 (N22323, N22319, N2418, N15416, N19491);
nor NOR2 (N22324, N22323, N4906);
buf BUF1 (N22325, N22318);
nor NOR4 (N22326, N22316, N12752, N11727, N751);
not NOT1 (N22327, N22320);
buf BUF1 (N22328, N22321);
and AND3 (N22329, N22325, N10372, N5461);
nor NOR4 (N22330, N22314, N20179, N21780, N13451);
not NOT1 (N22331, N22324);
not NOT1 (N22332, N22315);
nor NOR3 (N22333, N22330, N3115, N18971);
nand NAND4 (N22334, N22284, N20441, N7103, N3315);
nor NOR4 (N22335, N22329, N19279, N10000, N4767);
nor NOR2 (N22336, N22326, N742);
nand NAND3 (N22337, N22336, N11540, N4577);
and AND3 (N22338, N22334, N268, N20310);
or OR2 (N22339, N22335, N3741);
or OR2 (N22340, N22328, N2905);
or OR3 (N22341, N22340, N12025, N12930);
nor NOR4 (N22342, N22339, N5925, N7893, N15565);
not NOT1 (N22343, N22332);
buf BUF1 (N22344, N22304);
xor XOR2 (N22345, N22331, N2873);
xor XOR2 (N22346, N22344, N11965);
nand NAND2 (N22347, N22337, N2912);
xor XOR2 (N22348, N22322, N1721);
nand NAND4 (N22349, N22333, N18826, N7179, N9118);
and AND3 (N22350, N22348, N1438, N10491);
not NOT1 (N22351, N22342);
or OR4 (N22352, N22341, N8182, N2962, N120);
nand NAND4 (N22353, N22347, N1963, N10560, N4578);
and AND2 (N22354, N22351, N7755);
nor NOR4 (N22355, N22345, N3846, N15192, N1759);
nor NOR2 (N22356, N22350, N6428);
xor XOR2 (N22357, N22355, N3915);
nor NOR3 (N22358, N22357, N9123, N18298);
nand NAND4 (N22359, N22338, N8212, N2709, N14140);
xor XOR2 (N22360, N22359, N3171);
xor XOR2 (N22361, N22353, N18297);
nor NOR3 (N22362, N22327, N18988, N18858);
not NOT1 (N22363, N22354);
not NOT1 (N22364, N22343);
not NOT1 (N22365, N22361);
buf BUF1 (N22366, N22352);
nand NAND2 (N22367, N22366, N20111);
xor XOR2 (N22368, N22365, N797);
xor XOR2 (N22369, N22364, N17128);
nand NAND3 (N22370, N22369, N9301, N12015);
xor XOR2 (N22371, N22346, N8681);
not NOT1 (N22372, N22367);
xor XOR2 (N22373, N22370, N521);
buf BUF1 (N22374, N22358);
nor NOR4 (N22375, N22374, N3281, N21373, N17593);
and AND2 (N22376, N22372, N19546);
xor XOR2 (N22377, N22349, N1713);
buf BUF1 (N22378, N22360);
nand NAND3 (N22379, N22377, N17332, N1861);
xor XOR2 (N22380, N22371, N22330);
or OR4 (N22381, N22375, N15602, N14096, N1605);
and AND3 (N22382, N22376, N6818, N9472);
and AND2 (N22383, N22379, N15408);
not NOT1 (N22384, N22380);
not NOT1 (N22385, N22381);
nand NAND3 (N22386, N22356, N5964, N18594);
xor XOR2 (N22387, N22368, N2412);
nor NOR4 (N22388, N22383, N21003, N16229, N2073);
not NOT1 (N22389, N22378);
nand NAND3 (N22390, N22373, N10385, N15741);
and AND2 (N22391, N22390, N12515);
xor XOR2 (N22392, N22384, N18301);
buf BUF1 (N22393, N22386);
nor NOR3 (N22394, N22362, N5630, N20168);
xor XOR2 (N22395, N22394, N20529);
nand NAND2 (N22396, N22363, N8974);
and AND2 (N22397, N22385, N4199);
nor NOR3 (N22398, N22396, N10311, N13585);
nand NAND3 (N22399, N22393, N8723, N8063);
not NOT1 (N22400, N22387);
xor XOR2 (N22401, N22388, N22386);
nand NAND3 (N22402, N22399, N3323, N1677);
nor NOR3 (N22403, N22400, N6808, N13825);
or OR3 (N22404, N22398, N7649, N14022);
buf BUF1 (N22405, N22404);
nor NOR2 (N22406, N22397, N17654);
xor XOR2 (N22407, N22403, N20256);
nand NAND3 (N22408, N22401, N9304, N2018);
not NOT1 (N22409, N22392);
not NOT1 (N22410, N22406);
or OR2 (N22411, N22405, N22036);
xor XOR2 (N22412, N22389, N3312);
nor NOR3 (N22413, N22402, N3681, N842);
buf BUF1 (N22414, N22412);
nor NOR3 (N22415, N22408, N2874, N19015);
nor NOR2 (N22416, N22413, N18993);
and AND3 (N22417, N22395, N13823, N20835);
or OR3 (N22418, N22416, N4076, N5227);
xor XOR2 (N22419, N22417, N22251);
or OR3 (N22420, N22391, N17089, N9525);
not NOT1 (N22421, N22407);
not NOT1 (N22422, N22409);
not NOT1 (N22423, N22421);
xor XOR2 (N22424, N22419, N6738);
and AND3 (N22425, N22382, N6739, N376);
nor NOR3 (N22426, N22410, N8059, N634);
nor NOR4 (N22427, N22420, N19924, N7668, N2416);
nor NOR4 (N22428, N22423, N14692, N16138, N22024);
nand NAND3 (N22429, N22425, N3467, N2103);
buf BUF1 (N22430, N22427);
xor XOR2 (N22431, N22415, N21792);
buf BUF1 (N22432, N22411);
nand NAND4 (N22433, N22431, N20736, N596, N4717);
nand NAND2 (N22434, N22418, N12859);
buf BUF1 (N22435, N22432);
not NOT1 (N22436, N22428);
nand NAND4 (N22437, N22424, N8265, N11899, N225);
buf BUF1 (N22438, N22437);
nand NAND2 (N22439, N22436, N16614);
not NOT1 (N22440, N22438);
xor XOR2 (N22441, N22414, N13956);
nor NOR4 (N22442, N22430, N5957, N16671, N6682);
nor NOR2 (N22443, N22434, N20002);
nand NAND2 (N22444, N22441, N5993);
xor XOR2 (N22445, N22443, N13723);
and AND3 (N22446, N22422, N10996, N11696);
buf BUF1 (N22447, N22429);
buf BUF1 (N22448, N22447);
not NOT1 (N22449, N22446);
buf BUF1 (N22450, N22435);
xor XOR2 (N22451, N22439, N992);
and AND3 (N22452, N22445, N17212, N12560);
buf BUF1 (N22453, N22451);
not NOT1 (N22454, N22448);
buf BUF1 (N22455, N22453);
nand NAND4 (N22456, N22455, N1544, N1868, N16578);
or OR3 (N22457, N22433, N5851, N9505);
or OR4 (N22458, N22449, N3620, N12528, N13108);
or OR3 (N22459, N22456, N13705, N10197);
xor XOR2 (N22460, N22450, N20806);
and AND3 (N22461, N22457, N14046, N7392);
xor XOR2 (N22462, N22459, N4170);
nor NOR4 (N22463, N22444, N4279, N2363, N17724);
buf BUF1 (N22464, N22426);
buf BUF1 (N22465, N22464);
and AND2 (N22466, N22440, N21118);
or OR4 (N22467, N22461, N11636, N19119, N4839);
buf BUF1 (N22468, N22465);
buf BUF1 (N22469, N22467);
nor NOR2 (N22470, N22454, N651);
or OR3 (N22471, N22452, N2255, N2331);
or OR4 (N22472, N22471, N3257, N6462, N14795);
not NOT1 (N22473, N22463);
and AND3 (N22474, N22472, N7909, N17126);
nand NAND2 (N22475, N22458, N7612);
nor NOR4 (N22476, N22442, N6241, N15841, N7943);
or OR2 (N22477, N22468, N16348);
nand NAND4 (N22478, N22466, N10609, N16727, N1130);
and AND4 (N22479, N22475, N10512, N3808, N19023);
nor NOR2 (N22480, N22469, N6608);
and AND2 (N22481, N22476, N4540);
nor NOR4 (N22482, N22470, N6182, N140, N16545);
xor XOR2 (N22483, N22479, N8250);
or OR4 (N22484, N22480, N4275, N2254, N12191);
and AND3 (N22485, N22483, N12751, N347);
not NOT1 (N22486, N22481);
nand NAND4 (N22487, N22482, N1712, N8835, N18363);
not NOT1 (N22488, N22460);
not NOT1 (N22489, N22484);
buf BUF1 (N22490, N22478);
nor NOR4 (N22491, N22474, N4200, N6416, N14513);
xor XOR2 (N22492, N22491, N8124);
xor XOR2 (N22493, N22489, N20835);
not NOT1 (N22494, N22490);
nor NOR4 (N22495, N22494, N13722, N6026, N8185);
nor NOR4 (N22496, N22493, N18106, N8631, N14649);
nor NOR3 (N22497, N22477, N6971, N15764);
xor XOR2 (N22498, N22486, N3248);
not NOT1 (N22499, N22473);
nand NAND2 (N22500, N22497, N17500);
not NOT1 (N22501, N22496);
buf BUF1 (N22502, N22498);
not NOT1 (N22503, N22501);
or OR3 (N22504, N22462, N8966, N145);
xor XOR2 (N22505, N22495, N21608);
xor XOR2 (N22506, N22485, N15389);
buf BUF1 (N22507, N22505);
not NOT1 (N22508, N22499);
xor XOR2 (N22509, N22500, N18030);
or OR3 (N22510, N22488, N2900, N342);
not NOT1 (N22511, N22503);
and AND3 (N22512, N22507, N11017, N20811);
nor NOR3 (N22513, N22512, N22498, N22406);
or OR2 (N22514, N22504, N11498);
not NOT1 (N22515, N22502);
or OR2 (N22516, N22514, N2027);
xor XOR2 (N22517, N22510, N251);
xor XOR2 (N22518, N22508, N6390);
nand NAND4 (N22519, N22515, N3270, N7090, N8225);
nand NAND3 (N22520, N22519, N8530, N2993);
nand NAND2 (N22521, N22513, N12785);
not NOT1 (N22522, N22521);
not NOT1 (N22523, N22492);
or OR2 (N22524, N22523, N15616);
xor XOR2 (N22525, N22487, N3570);
buf BUF1 (N22526, N22511);
xor XOR2 (N22527, N22525, N2216);
nand NAND3 (N22528, N22506, N18365, N9952);
and AND4 (N22529, N22520, N7649, N18312, N15513);
nand NAND2 (N22530, N22509, N12001);
nor NOR2 (N22531, N22522, N4549);
or OR4 (N22532, N22518, N11013, N22268, N3899);
nor NOR2 (N22533, N22524, N22069);
not NOT1 (N22534, N22528);
nand NAND2 (N22535, N22526, N16636);
nand NAND2 (N22536, N22530, N4403);
and AND4 (N22537, N22536, N20186, N16382, N3805);
and AND4 (N22538, N22529, N3442, N21242, N18086);
nand NAND2 (N22539, N22535, N782);
or OR3 (N22540, N22517, N5538, N17530);
not NOT1 (N22541, N22540);
buf BUF1 (N22542, N22538);
and AND2 (N22543, N22527, N9);
not NOT1 (N22544, N22541);
buf BUF1 (N22545, N22534);
or OR4 (N22546, N22542, N9732, N17570, N679);
xor XOR2 (N22547, N22543, N19647);
or OR2 (N22548, N22539, N4998);
not NOT1 (N22549, N22532);
nor NOR2 (N22550, N22547, N12524);
nand NAND3 (N22551, N22550, N1013, N7833);
or OR2 (N22552, N22533, N17400);
xor XOR2 (N22553, N22549, N15797);
and AND3 (N22554, N22552, N5668, N21699);
xor XOR2 (N22555, N22546, N15873);
buf BUF1 (N22556, N22537);
nor NOR4 (N22557, N22555, N13119, N11310, N7841);
or OR3 (N22558, N22545, N2046, N14299);
xor XOR2 (N22559, N22553, N7772);
and AND2 (N22560, N22548, N4337);
xor XOR2 (N22561, N22559, N11218);
nand NAND2 (N22562, N22557, N9738);
and AND3 (N22563, N22561, N17718, N8827);
not NOT1 (N22564, N22544);
not NOT1 (N22565, N22564);
nand NAND4 (N22566, N22556, N13767, N6549, N2806);
nand NAND4 (N22567, N22560, N19512, N6752, N5494);
or OR3 (N22568, N22563, N19688, N20526);
or OR4 (N22569, N22558, N11592, N18576, N17948);
nand NAND4 (N22570, N22531, N20967, N11365, N4326);
buf BUF1 (N22571, N22569);
nand NAND3 (N22572, N22566, N2610, N2564);
nand NAND3 (N22573, N22565, N5516, N6219);
nor NOR3 (N22574, N22516, N140, N21017);
xor XOR2 (N22575, N22574, N18446);
nor NOR2 (N22576, N22562, N3583);
nor NOR2 (N22577, N22573, N8417);
xor XOR2 (N22578, N22571, N1744);
xor XOR2 (N22579, N22568, N1027);
buf BUF1 (N22580, N22578);
or OR3 (N22581, N22572, N1814, N19861);
buf BUF1 (N22582, N22579);
nor NOR2 (N22583, N22580, N14566);
nor NOR4 (N22584, N22577, N17529, N7814, N16057);
nor NOR2 (N22585, N22554, N9421);
xor XOR2 (N22586, N22575, N12704);
nor NOR4 (N22587, N22581, N1552, N3247, N7568);
buf BUF1 (N22588, N22585);
buf BUF1 (N22589, N22582);
buf BUF1 (N22590, N22589);
and AND4 (N22591, N22586, N21782, N4837, N3471);
xor XOR2 (N22592, N22551, N1906);
xor XOR2 (N22593, N22570, N20913);
xor XOR2 (N22594, N22593, N4081);
not NOT1 (N22595, N22567);
not NOT1 (N22596, N22576);
or OR2 (N22597, N22583, N22396);
nor NOR2 (N22598, N22597, N19573);
buf BUF1 (N22599, N22588);
xor XOR2 (N22600, N22595, N663);
or OR2 (N22601, N22592, N4097);
nor NOR2 (N22602, N22584, N20893);
and AND2 (N22603, N22600, N8329);
buf BUF1 (N22604, N22599);
nand NAND2 (N22605, N22594, N7263);
and AND3 (N22606, N22587, N2043, N2279);
nand NAND4 (N22607, N22604, N17091, N15626, N7880);
nand NAND4 (N22608, N22603, N18336, N1054, N21644);
xor XOR2 (N22609, N22605, N16511);
nor NOR4 (N22610, N22596, N14554, N843, N10563);
xor XOR2 (N22611, N22601, N11447);
xor XOR2 (N22612, N22609, N8836);
nor NOR2 (N22613, N22606, N21237);
nor NOR4 (N22614, N22612, N14964, N207, N2790);
buf BUF1 (N22615, N22611);
and AND2 (N22616, N22613, N4745);
or OR3 (N22617, N22616, N3325, N10689);
xor XOR2 (N22618, N22607, N8750);
not NOT1 (N22619, N22598);
nor NOR3 (N22620, N22619, N8688, N21075);
and AND2 (N22621, N22615, N17492);
nor NOR3 (N22622, N22602, N10136, N19878);
buf BUF1 (N22623, N22590);
buf BUF1 (N22624, N22622);
or OR3 (N22625, N22608, N17020, N698);
buf BUF1 (N22626, N22621);
and AND3 (N22627, N22623, N7381, N14423);
nor NOR4 (N22628, N22614, N20492, N2530, N20636);
buf BUF1 (N22629, N22625);
xor XOR2 (N22630, N22629, N3150);
nand NAND2 (N22631, N22617, N14286);
nand NAND3 (N22632, N22630, N15022, N14320);
or OR3 (N22633, N22591, N426, N16762);
not NOT1 (N22634, N22628);
or OR4 (N22635, N22631, N5708, N5330, N1198);
nor NOR4 (N22636, N22610, N5442, N9881, N15213);
xor XOR2 (N22637, N22624, N5052);
and AND2 (N22638, N22632, N298);
xor XOR2 (N22639, N22626, N3956);
not NOT1 (N22640, N22635);
xor XOR2 (N22641, N22620, N46);
xor XOR2 (N22642, N22633, N4844);
nand NAND4 (N22643, N22618, N12233, N12530, N4500);
and AND2 (N22644, N22640, N18887);
and AND3 (N22645, N22639, N11466, N18555);
nand NAND3 (N22646, N22637, N17272, N20688);
nand NAND3 (N22647, N22627, N15096, N3315);
nor NOR3 (N22648, N22644, N7524, N10268);
nand NAND4 (N22649, N22642, N15264, N564, N4324);
nand NAND4 (N22650, N22634, N17056, N5813, N13809);
nor NOR3 (N22651, N22648, N1921, N13530);
nor NOR3 (N22652, N22636, N2639, N6245);
nor NOR2 (N22653, N22649, N15333);
buf BUF1 (N22654, N22646);
xor XOR2 (N22655, N22653, N9167);
xor XOR2 (N22656, N22643, N20570);
not NOT1 (N22657, N22652);
or OR2 (N22658, N22655, N8392);
and AND3 (N22659, N22647, N12589, N20333);
nor NOR4 (N22660, N22656, N15330, N17499, N2666);
xor XOR2 (N22661, N22638, N20437);
nor NOR4 (N22662, N22661, N9127, N20108, N2126);
buf BUF1 (N22663, N22641);
nand NAND2 (N22664, N22662, N83);
xor XOR2 (N22665, N22663, N17328);
nand NAND4 (N22666, N22659, N17495, N22537, N12239);
or OR2 (N22667, N22665, N613);
not NOT1 (N22668, N22658);
xor XOR2 (N22669, N22650, N16451);
or OR2 (N22670, N22654, N5760);
buf BUF1 (N22671, N22664);
nor NOR2 (N22672, N22667, N6454);
not NOT1 (N22673, N22657);
buf BUF1 (N22674, N22670);
nor NOR4 (N22675, N22668, N13926, N8007, N13608);
or OR2 (N22676, N22669, N14425);
and AND4 (N22677, N22674, N19566, N7149, N18849);
xor XOR2 (N22678, N22645, N17976);
xor XOR2 (N22679, N22671, N18921);
xor XOR2 (N22680, N22675, N12266);
xor XOR2 (N22681, N22673, N21523);
nand NAND2 (N22682, N22672, N8027);
buf BUF1 (N22683, N22681);
not NOT1 (N22684, N22660);
nor NOR4 (N22685, N22677, N12224, N3705, N4306);
or OR4 (N22686, N22651, N19963, N2298, N18089);
nor NOR2 (N22687, N22680, N20142);
not NOT1 (N22688, N22684);
or OR4 (N22689, N22683, N20625, N4522, N11245);
buf BUF1 (N22690, N22666);
xor XOR2 (N22691, N22676, N15037);
or OR3 (N22692, N22687, N3308, N19162);
and AND3 (N22693, N22691, N1631, N11690);
or OR4 (N22694, N22685, N6359, N15376, N22282);
xor XOR2 (N22695, N22689, N4117);
nand NAND4 (N22696, N22682, N6706, N1513, N7234);
not NOT1 (N22697, N22696);
and AND3 (N22698, N22688, N15562, N2844);
and AND2 (N22699, N22697, N14994);
nand NAND2 (N22700, N22678, N1306);
and AND3 (N22701, N22700, N14557, N656);
and AND3 (N22702, N22692, N10806, N10116);
and AND4 (N22703, N22699, N21677, N17862, N19866);
not NOT1 (N22704, N22694);
buf BUF1 (N22705, N22698);
or OR2 (N22706, N22705, N5235);
nor NOR2 (N22707, N22703, N11335);
nand NAND4 (N22708, N22701, N20787, N22271, N8458);
nor NOR2 (N22709, N22708, N20509);
xor XOR2 (N22710, N22686, N11061);
and AND3 (N22711, N22710, N1274, N2558);
and AND4 (N22712, N22709, N21229, N12554, N7198);
nand NAND2 (N22713, N22690, N22550);
buf BUF1 (N22714, N22702);
and AND3 (N22715, N22679, N1961, N7233);
and AND2 (N22716, N22707, N20189);
and AND2 (N22717, N22714, N15986);
not NOT1 (N22718, N22712);
or OR4 (N22719, N22716, N22438, N19595, N8661);
and AND3 (N22720, N22695, N11230, N3640);
nand NAND4 (N22721, N22693, N19081, N5058, N1557);
and AND3 (N22722, N22719, N2528, N17343);
xor XOR2 (N22723, N22704, N14290);
xor XOR2 (N22724, N22713, N10636);
or OR4 (N22725, N22721, N6573, N4631, N4358);
buf BUF1 (N22726, N22715);
nor NOR2 (N22727, N22711, N19899);
nor NOR3 (N22728, N22722, N6056, N21178);
xor XOR2 (N22729, N22727, N14565);
nor NOR4 (N22730, N22729, N6319, N18609, N14968);
xor XOR2 (N22731, N22728, N1202);
and AND2 (N22732, N22720, N14587);
and AND4 (N22733, N22723, N1103, N19193, N16061);
not NOT1 (N22734, N22730);
nor NOR3 (N22735, N22706, N16163, N15823);
or OR2 (N22736, N22726, N17765);
or OR3 (N22737, N22731, N8157, N12738);
buf BUF1 (N22738, N22732);
and AND3 (N22739, N22738, N10988, N14417);
or OR4 (N22740, N22733, N11891, N14213, N6362);
buf BUF1 (N22741, N22718);
or OR3 (N22742, N22735, N19935, N3288);
or OR2 (N22743, N22742, N9556);
xor XOR2 (N22744, N22737, N266);
buf BUF1 (N22745, N22743);
not NOT1 (N22746, N22744);
xor XOR2 (N22747, N22736, N18195);
not NOT1 (N22748, N22725);
nor NOR2 (N22749, N22748, N21098);
buf BUF1 (N22750, N22745);
or OR4 (N22751, N22741, N4300, N18253, N2545);
and AND2 (N22752, N22749, N1927);
xor XOR2 (N22753, N22739, N8393);
not NOT1 (N22754, N22747);
nor NOR2 (N22755, N22740, N1389);
nand NAND4 (N22756, N22753, N6436, N22108, N15616);
or OR2 (N22757, N22756, N12601);
and AND2 (N22758, N22757, N20375);
xor XOR2 (N22759, N22751, N7735);
xor XOR2 (N22760, N22752, N15245);
nor NOR4 (N22761, N22746, N14109, N17818, N15174);
or OR4 (N22762, N22755, N9413, N11964, N16858);
and AND3 (N22763, N22734, N2840, N6769);
nand NAND4 (N22764, N22759, N1365, N15396, N15464);
and AND3 (N22765, N22763, N1930, N16588);
buf BUF1 (N22766, N22760);
and AND4 (N22767, N22758, N11097, N11745, N809);
xor XOR2 (N22768, N22762, N9459);
and AND3 (N22769, N22766, N9337, N14929);
not NOT1 (N22770, N22750);
and AND2 (N22771, N22717, N16798);
nor NOR2 (N22772, N22724, N3417);
buf BUF1 (N22773, N22754);
or OR3 (N22774, N22767, N7151, N21163);
or OR4 (N22775, N22771, N1507, N22506, N3704);
nor NOR3 (N22776, N22764, N1547, N7263);
or OR2 (N22777, N22774, N10109);
nand NAND3 (N22778, N22777, N20770, N7262);
or OR2 (N22779, N22778, N18851);
nand NAND2 (N22780, N22779, N3554);
and AND2 (N22781, N22769, N5512);
xor XOR2 (N22782, N22761, N22366);
xor XOR2 (N22783, N22773, N8559);
xor XOR2 (N22784, N22783, N20356);
buf BUF1 (N22785, N22780);
not NOT1 (N22786, N22781);
nand NAND4 (N22787, N22770, N9438, N9247, N17324);
and AND3 (N22788, N22776, N17052, N14109);
nand NAND2 (N22789, N22784, N14792);
nand NAND3 (N22790, N22765, N8689, N2612);
xor XOR2 (N22791, N22782, N1078);
xor XOR2 (N22792, N22786, N16211);
and AND2 (N22793, N22788, N4381);
buf BUF1 (N22794, N22772);
nand NAND4 (N22795, N22775, N2832, N9175, N5556);
nor NOR2 (N22796, N22787, N17783);
xor XOR2 (N22797, N22790, N11544);
or OR4 (N22798, N22785, N200, N19046, N20904);
not NOT1 (N22799, N22797);
or OR4 (N22800, N22791, N18033, N11704, N19056);
or OR2 (N22801, N22796, N22413);
nand NAND3 (N22802, N22768, N1422, N13826);
or OR4 (N22803, N22802, N154, N15700, N17893);
and AND3 (N22804, N22793, N3019, N18223);
xor XOR2 (N22805, N22798, N16921);
not NOT1 (N22806, N22801);
nand NAND2 (N22807, N22789, N21682);
nor NOR3 (N22808, N22806, N8066, N10571);
nand NAND2 (N22809, N22808, N730);
or OR3 (N22810, N22792, N2174, N18965);
xor XOR2 (N22811, N22794, N7140);
xor XOR2 (N22812, N22805, N21963);
buf BUF1 (N22813, N22810);
buf BUF1 (N22814, N22795);
nand NAND3 (N22815, N22807, N10115, N4224);
nor NOR2 (N22816, N22799, N9605);
xor XOR2 (N22817, N22811, N1224);
buf BUF1 (N22818, N22813);
not NOT1 (N22819, N22816);
nor NOR3 (N22820, N22812, N15089, N12777);
nand NAND2 (N22821, N22800, N14801);
not NOT1 (N22822, N22818);
nor NOR4 (N22823, N22822, N11118, N4803, N4216);
and AND2 (N22824, N22809, N15366);
buf BUF1 (N22825, N22821);
and AND4 (N22826, N22819, N5080, N17968, N22739);
not NOT1 (N22827, N22825);
or OR3 (N22828, N22820, N1450, N3476);
and AND3 (N22829, N22828, N12209, N12112);
and AND4 (N22830, N22829, N20993, N20811, N9551);
nor NOR2 (N22831, N22804, N11618);
nor NOR2 (N22832, N22823, N19442);
nand NAND2 (N22833, N22814, N6630);
buf BUF1 (N22834, N22824);
or OR2 (N22835, N22834, N13214);
and AND2 (N22836, N22835, N16590);
nor NOR4 (N22837, N22826, N16396, N8211, N13187);
not NOT1 (N22838, N22803);
and AND3 (N22839, N22827, N12960, N5269);
or OR2 (N22840, N22817, N13128);
or OR3 (N22841, N22833, N1028, N18404);
and AND3 (N22842, N22831, N6884, N10897);
nand NAND3 (N22843, N22830, N3668, N14373);
xor XOR2 (N22844, N22837, N5714);
buf BUF1 (N22845, N22839);
nor NOR3 (N22846, N22832, N6522, N15674);
buf BUF1 (N22847, N22815);
nand NAND2 (N22848, N22838, N15971);
nor NOR2 (N22849, N22844, N17779);
and AND4 (N22850, N22846, N14563, N2558, N19946);
nor NOR3 (N22851, N22850, N13645, N21936);
or OR4 (N22852, N22849, N3726, N2986, N18660);
nand NAND2 (N22853, N22843, N3519);
nand NAND4 (N22854, N22841, N18127, N17721, N6714);
or OR3 (N22855, N22852, N567, N15579);
or OR4 (N22856, N22851, N5283, N4128, N1718);
xor XOR2 (N22857, N22842, N18006);
nand NAND4 (N22858, N22848, N17859, N19154, N22495);
or OR2 (N22859, N22847, N13767);
nor NOR3 (N22860, N22855, N10115, N11966);
or OR3 (N22861, N22854, N17416, N11375);
xor XOR2 (N22862, N22845, N14482);
nor NOR3 (N22863, N22857, N10435, N7094);
buf BUF1 (N22864, N22858);
nor NOR2 (N22865, N22853, N20818);
nand NAND4 (N22866, N22862, N17185, N14684, N21753);
and AND4 (N22867, N22840, N20244, N6310, N6172);
nand NAND3 (N22868, N22867, N12912, N8992);
not NOT1 (N22869, N22860);
not NOT1 (N22870, N22864);
nand NAND2 (N22871, N22859, N546);
not NOT1 (N22872, N22868);
nand NAND3 (N22873, N22869, N16541, N9845);
or OR2 (N22874, N22866, N7518);
nor NOR2 (N22875, N22871, N4794);
or OR2 (N22876, N22861, N17471);
nor NOR2 (N22877, N22876, N12840);
nor NOR2 (N22878, N22872, N19427);
buf BUF1 (N22879, N22873);
xor XOR2 (N22880, N22879, N1395);
not NOT1 (N22881, N22880);
nor NOR4 (N22882, N22870, N4070, N12354, N3456);
or OR2 (N22883, N22874, N20757);
nand NAND4 (N22884, N22877, N7304, N21411, N17276);
buf BUF1 (N22885, N22865);
xor XOR2 (N22886, N22884, N4029);
buf BUF1 (N22887, N22883);
buf BUF1 (N22888, N22885);
nor NOR3 (N22889, N22875, N11220, N10946);
or OR2 (N22890, N22836, N3235);
or OR4 (N22891, N22878, N7092, N15687, N4674);
nor NOR4 (N22892, N22891, N13414, N6041, N21574);
and AND2 (N22893, N22890, N21478);
nor NOR4 (N22894, N22889, N22142, N17914, N8383);
nor NOR4 (N22895, N22882, N12080, N18223, N8994);
xor XOR2 (N22896, N22863, N18293);
xor XOR2 (N22897, N22888, N12886);
and AND4 (N22898, N22893, N22723, N6971, N9914);
buf BUF1 (N22899, N22886);
nand NAND4 (N22900, N22856, N7954, N15844, N2883);
xor XOR2 (N22901, N22900, N14844);
or OR3 (N22902, N22897, N19240, N17334);
or OR2 (N22903, N22894, N6511);
not NOT1 (N22904, N22881);
or OR4 (N22905, N22887, N13679, N20391, N17570);
and AND2 (N22906, N22905, N23);
or OR2 (N22907, N22898, N19181);
not NOT1 (N22908, N22902);
nand NAND2 (N22909, N22896, N9582);
nand NAND4 (N22910, N22899, N11932, N10154, N6205);
xor XOR2 (N22911, N22910, N21305);
xor XOR2 (N22912, N22906, N18470);
xor XOR2 (N22913, N22903, N11574);
nor NOR3 (N22914, N22901, N6555, N12269);
not NOT1 (N22915, N22904);
xor XOR2 (N22916, N22915, N15931);
and AND3 (N22917, N22911, N10174, N20251);
not NOT1 (N22918, N22914);
nor NOR3 (N22919, N22916, N2361, N20948);
or OR4 (N22920, N22919, N2129, N13552, N11967);
and AND2 (N22921, N22912, N10184);
nor NOR3 (N22922, N22892, N11829, N4829);
nand NAND3 (N22923, N22921, N1659, N9456);
buf BUF1 (N22924, N22917);
nor NOR4 (N22925, N22920, N12495, N6159, N2469);
and AND3 (N22926, N22918, N8752, N5585);
nand NAND2 (N22927, N22909, N5990);
not NOT1 (N22928, N22913);
not NOT1 (N22929, N22895);
and AND4 (N22930, N22927, N2142, N4118, N745);
xor XOR2 (N22931, N22908, N9536);
nor NOR3 (N22932, N22924, N17147, N17786);
xor XOR2 (N22933, N22932, N22695);
or OR3 (N22934, N22926, N13482, N8415);
or OR4 (N22935, N22934, N9901, N20014, N6646);
not NOT1 (N22936, N22933);
nand NAND3 (N22937, N22936, N11767, N10602);
or OR4 (N22938, N22937, N8559, N20344, N21993);
nand NAND3 (N22939, N22922, N12873, N2490);
nor NOR2 (N22940, N22935, N12487);
or OR3 (N22941, N22925, N19304, N18850);
nor NOR2 (N22942, N22931, N9574);
or OR3 (N22943, N22929, N21050, N2056);
not NOT1 (N22944, N22928);
xor XOR2 (N22945, N22938, N9506);
not NOT1 (N22946, N22944);
not NOT1 (N22947, N22923);
xor XOR2 (N22948, N22930, N19968);
xor XOR2 (N22949, N22939, N2134);
nand NAND2 (N22950, N22943, N5097);
and AND2 (N22951, N22945, N16260);
or OR4 (N22952, N22940, N2094, N1177, N22723);
not NOT1 (N22953, N22950);
or OR3 (N22954, N22946, N2022, N17569);
or OR2 (N22955, N22941, N5394);
nor NOR2 (N22956, N22952, N18172);
not NOT1 (N22957, N22949);
nand NAND2 (N22958, N22953, N19208);
xor XOR2 (N22959, N22955, N17141);
not NOT1 (N22960, N22959);
and AND2 (N22961, N22954, N13071);
and AND4 (N22962, N22942, N5343, N597, N19868);
xor XOR2 (N22963, N22951, N3285);
or OR3 (N22964, N22956, N12444, N3307);
and AND3 (N22965, N22960, N17063, N5124);
nand NAND3 (N22966, N22958, N4562, N30);
nor NOR2 (N22967, N22907, N18039);
or OR4 (N22968, N22957, N6976, N14919, N13344);
buf BUF1 (N22969, N22964);
and AND4 (N22970, N22966, N8508, N22441, N8557);
xor XOR2 (N22971, N22948, N22472);
not NOT1 (N22972, N22967);
and AND2 (N22973, N22968, N16327);
buf BUF1 (N22974, N22973);
or OR4 (N22975, N22961, N14810, N1616, N136);
buf BUF1 (N22976, N22962);
or OR3 (N22977, N22975, N5870, N19108);
buf BUF1 (N22978, N22970);
buf BUF1 (N22979, N22974);
xor XOR2 (N22980, N22963, N5296);
and AND2 (N22981, N22978, N1345);
and AND4 (N22982, N22981, N10236, N13547, N5728);
and AND2 (N22983, N22947, N7974);
not NOT1 (N22984, N22965);
buf BUF1 (N22985, N22971);
xor XOR2 (N22986, N22976, N790);
xor XOR2 (N22987, N22977, N21756);
nand NAND2 (N22988, N22984, N19273);
xor XOR2 (N22989, N22988, N7427);
not NOT1 (N22990, N22983);
xor XOR2 (N22991, N22987, N5987);
not NOT1 (N22992, N22991);
or OR3 (N22993, N22986, N17266, N10778);
or OR3 (N22994, N22969, N16406, N9648);
not NOT1 (N22995, N22972);
not NOT1 (N22996, N22992);
buf BUF1 (N22997, N22985);
and AND3 (N22998, N22996, N10162, N8219);
nand NAND3 (N22999, N22997, N13148, N1312);
nor NOR2 (N23000, N22979, N8539);
and AND4 (N23001, N22998, N2270, N2151, N7830);
not NOT1 (N23002, N22980);
nand NAND3 (N23003, N22994, N21694, N7723);
nand NAND3 (N23004, N22989, N892, N16133);
and AND2 (N23005, N23001, N17598);
or OR3 (N23006, N22999, N9653, N4104);
xor XOR2 (N23007, N23004, N10449);
and AND2 (N23008, N23005, N815);
buf BUF1 (N23009, N23000);
xor XOR2 (N23010, N22995, N13896);
buf BUF1 (N23011, N23010);
xor XOR2 (N23012, N23007, N17320);
nor NOR2 (N23013, N22990, N3448);
xor XOR2 (N23014, N22993, N9225);
nor NOR2 (N23015, N23006, N14622);
and AND2 (N23016, N23014, N14601);
xor XOR2 (N23017, N23016, N3553);
and AND2 (N23018, N23017, N9405);
buf BUF1 (N23019, N23002);
nand NAND3 (N23020, N23018, N12379, N8522);
nand NAND4 (N23021, N23012, N14603, N22519, N6168);
and AND3 (N23022, N23008, N1131, N14011);
buf BUF1 (N23023, N23022);
or OR3 (N23024, N23019, N17945, N13081);
or OR4 (N23025, N23013, N8303, N11434, N1435);
xor XOR2 (N23026, N23021, N710);
buf BUF1 (N23027, N22982);
nor NOR4 (N23028, N23024, N18505, N9867, N7119);
nor NOR4 (N23029, N23011, N14807, N19546, N17566);
not NOT1 (N23030, N23020);
not NOT1 (N23031, N23030);
buf BUF1 (N23032, N23028);
buf BUF1 (N23033, N23027);
buf BUF1 (N23034, N23003);
buf BUF1 (N23035, N23033);
buf BUF1 (N23036, N23034);
nand NAND2 (N23037, N23023, N14934);
nand NAND3 (N23038, N23031, N5703, N14222);
or OR2 (N23039, N23029, N21101);
xor XOR2 (N23040, N23035, N11322);
not NOT1 (N23041, N23040);
nor NOR4 (N23042, N23036, N7881, N11963, N6641);
or OR4 (N23043, N23025, N9477, N64, N14628);
buf BUF1 (N23044, N23041);
or OR2 (N23045, N23015, N1497);
and AND4 (N23046, N23009, N1213, N14384, N15869);
not NOT1 (N23047, N23043);
xor XOR2 (N23048, N23039, N12518);
or OR4 (N23049, N23044, N499, N18688, N5248);
buf BUF1 (N23050, N23046);
nor NOR3 (N23051, N23042, N16973, N12130);
and AND3 (N23052, N23037, N19125, N6599);
nand NAND2 (N23053, N23051, N21213);
and AND4 (N23054, N23045, N1637, N7435, N18840);
buf BUF1 (N23055, N23050);
xor XOR2 (N23056, N23047, N3795);
and AND2 (N23057, N23038, N22930);
nor NOR2 (N23058, N23049, N13350);
or OR2 (N23059, N23053, N13360);
buf BUF1 (N23060, N23052);
xor XOR2 (N23061, N23057, N7157);
not NOT1 (N23062, N23048);
not NOT1 (N23063, N23054);
nor NOR2 (N23064, N23059, N19939);
xor XOR2 (N23065, N23058, N768);
or OR4 (N23066, N23056, N18604, N2267, N6984);
nor NOR3 (N23067, N23066, N7304, N19662);
or OR3 (N23068, N23061, N127, N11770);
nand NAND3 (N23069, N23064, N12851, N19873);
nor NOR4 (N23070, N23065, N5844, N2504, N15163);
nor NOR4 (N23071, N23060, N7507, N2088, N12863);
or OR3 (N23072, N23032, N13441, N211);
not NOT1 (N23073, N23062);
nor NOR3 (N23074, N23067, N22936, N17066);
nor NOR3 (N23075, N23070, N20794, N16041);
and AND3 (N23076, N23074, N3573, N22335);
nor NOR4 (N23077, N23055, N12906, N2025, N18790);
or OR2 (N23078, N23071, N18947);
or OR4 (N23079, N23072, N21951, N14370, N21584);
nand NAND2 (N23080, N23076, N2450);
xor XOR2 (N23081, N23078, N6339);
not NOT1 (N23082, N23075);
nand NAND3 (N23083, N23073, N6576, N786);
nor NOR2 (N23084, N23082, N4721);
nor NOR2 (N23085, N23026, N5166);
not NOT1 (N23086, N23080);
or OR2 (N23087, N23085, N11948);
or OR2 (N23088, N23069, N20496);
buf BUF1 (N23089, N23086);
nand NAND4 (N23090, N23081, N19148, N17940, N18126);
nand NAND4 (N23091, N23063, N21787, N11335, N4568);
nand NAND2 (N23092, N23087, N21543);
xor XOR2 (N23093, N23091, N922);
not NOT1 (N23094, N23079);
xor XOR2 (N23095, N23090, N18444);
nand NAND4 (N23096, N23084, N1667, N5965, N11664);
and AND3 (N23097, N23093, N8317, N13402);
nand NAND3 (N23098, N23094, N5256, N13702);
nand NAND2 (N23099, N23088, N11618);
not NOT1 (N23100, N23083);
not NOT1 (N23101, N23095);
xor XOR2 (N23102, N23101, N21431);
and AND3 (N23103, N23092, N19099, N15558);
not NOT1 (N23104, N23096);
buf BUF1 (N23105, N23104);
nand NAND4 (N23106, N23089, N6416, N19497, N5029);
buf BUF1 (N23107, N23105);
and AND2 (N23108, N23077, N1890);
xor XOR2 (N23109, N23097, N16523);
and AND3 (N23110, N23099, N17821, N12407);
nor NOR2 (N23111, N23106, N3687);
nand NAND2 (N23112, N23107, N6897);
xor XOR2 (N23113, N23110, N17739);
nor NOR4 (N23114, N23113, N2921, N2883, N6348);
and AND3 (N23115, N23102, N17175, N4727);
and AND2 (N23116, N23114, N17258);
buf BUF1 (N23117, N23103);
not NOT1 (N23118, N23115);
buf BUF1 (N23119, N23068);
nor NOR3 (N23120, N23117, N514, N9940);
and AND4 (N23121, N23109, N21136, N1151, N9062);
and AND4 (N23122, N23118, N19713, N13422, N6544);
nand NAND4 (N23123, N23098, N1285, N9335, N2346);
and AND4 (N23124, N23112, N22487, N7934, N1449);
or OR3 (N23125, N23116, N3916, N8031);
nor NOR3 (N23126, N23123, N16492, N11542);
or OR2 (N23127, N23120, N14565);
nor NOR4 (N23128, N23119, N6243, N16039, N2768);
buf BUF1 (N23129, N23121);
buf BUF1 (N23130, N23124);
or OR2 (N23131, N23130, N20158);
nor NOR4 (N23132, N23108, N4979, N278, N5882);
nand NAND2 (N23133, N23125, N8998);
xor XOR2 (N23134, N23122, N20807);
and AND3 (N23135, N23133, N6152, N5044);
nand NAND2 (N23136, N23129, N14277);
xor XOR2 (N23137, N23132, N14980);
and AND3 (N23138, N23128, N1287, N175);
buf BUF1 (N23139, N23135);
or OR3 (N23140, N23138, N5578, N12531);
nor NOR4 (N23141, N23111, N19668, N20236, N1624);
nand NAND3 (N23142, N23127, N9240, N22045);
nand NAND3 (N23143, N23131, N8318, N551);
and AND4 (N23144, N23139, N15798, N20454, N19358);
and AND2 (N23145, N23126, N9746);
xor XOR2 (N23146, N23137, N17415);
and AND3 (N23147, N23144, N14256, N18398);
nand NAND2 (N23148, N23146, N22860);
buf BUF1 (N23149, N23143);
nor NOR4 (N23150, N23100, N16035, N822, N3008);
or OR3 (N23151, N23134, N6278, N20205);
buf BUF1 (N23152, N23141);
nand NAND2 (N23153, N23150, N11770);
or OR2 (N23154, N23145, N13576);
or OR4 (N23155, N23152, N8997, N22757, N13322);
nand NAND2 (N23156, N23151, N17297);
nand NAND4 (N23157, N23153, N20917, N8589, N17463);
not NOT1 (N23158, N23147);
not NOT1 (N23159, N23148);
xor XOR2 (N23160, N23155, N585);
nand NAND4 (N23161, N23136, N8378, N11147, N22923);
nor NOR3 (N23162, N23142, N10516, N6195);
nor NOR2 (N23163, N23159, N5925);
not NOT1 (N23164, N23161);
nand NAND2 (N23165, N23160, N7952);
not NOT1 (N23166, N23157);
not NOT1 (N23167, N23140);
or OR2 (N23168, N23156, N15838);
or OR4 (N23169, N23167, N2292, N21754, N845);
nand NAND4 (N23170, N23154, N7895, N17861, N17578);
nor NOR2 (N23171, N23169, N20457);
buf BUF1 (N23172, N23165);
buf BUF1 (N23173, N23162);
not NOT1 (N23174, N23168);
not NOT1 (N23175, N23174);
and AND3 (N23176, N23163, N12207, N14363);
xor XOR2 (N23177, N23171, N19856);
not NOT1 (N23178, N23164);
nand NAND2 (N23179, N23177, N17793);
and AND4 (N23180, N23166, N8921, N16742, N7223);
xor XOR2 (N23181, N23158, N17779);
nand NAND3 (N23182, N23176, N22566, N11575);
buf BUF1 (N23183, N23173);
or OR4 (N23184, N23179, N5262, N19729, N2691);
xor XOR2 (N23185, N23180, N22848);
nor NOR2 (N23186, N23170, N18415);
and AND2 (N23187, N23172, N13033);
not NOT1 (N23188, N23181);
buf BUF1 (N23189, N23178);
not NOT1 (N23190, N23189);
nand NAND3 (N23191, N23149, N10990, N4567);
buf BUF1 (N23192, N23190);
buf BUF1 (N23193, N23182);
buf BUF1 (N23194, N23187);
nor NOR2 (N23195, N23194, N12029);
or OR4 (N23196, N23193, N21530, N14014, N7008);
nand NAND2 (N23197, N23192, N14525);
xor XOR2 (N23198, N23188, N380);
xor XOR2 (N23199, N23184, N2743);
or OR2 (N23200, N23199, N9424);
buf BUF1 (N23201, N23197);
not NOT1 (N23202, N23186);
buf BUF1 (N23203, N23202);
nand NAND4 (N23204, N23185, N20101, N15596, N15919);
nor NOR3 (N23205, N23198, N6156, N15140);
and AND2 (N23206, N23196, N6840);
xor XOR2 (N23207, N23204, N22171);
xor XOR2 (N23208, N23206, N5154);
not NOT1 (N23209, N23203);
nor NOR3 (N23210, N23195, N14576, N5272);
not NOT1 (N23211, N23191);
or OR3 (N23212, N23210, N21456, N21258);
buf BUF1 (N23213, N23209);
or OR4 (N23214, N23175, N352, N9082, N12036);
nand NAND4 (N23215, N23208, N21623, N2442, N20122);
not NOT1 (N23216, N23215);
and AND4 (N23217, N23211, N4704, N14385, N13374);
or OR3 (N23218, N23205, N9790, N5217);
nand NAND2 (N23219, N23200, N5504);
and AND2 (N23220, N23217, N8260);
buf BUF1 (N23221, N23183);
or OR3 (N23222, N23207, N12792, N17121);
xor XOR2 (N23223, N23221, N18154);
buf BUF1 (N23224, N23213);
nor NOR3 (N23225, N23201, N3495, N21612);
nand NAND4 (N23226, N23214, N18257, N22540, N2817);
or OR3 (N23227, N23220, N13820, N17398);
and AND4 (N23228, N23224, N8234, N14872, N14398);
buf BUF1 (N23229, N23218);
not NOT1 (N23230, N23225);
nand NAND4 (N23231, N23223, N1415, N5980, N19302);
not NOT1 (N23232, N23222);
nor NOR4 (N23233, N23228, N19587, N11580, N8488);
not NOT1 (N23234, N23226);
nand NAND4 (N23235, N23230, N19170, N4146, N5605);
buf BUF1 (N23236, N23235);
xor XOR2 (N23237, N23234, N9091);
nand NAND2 (N23238, N23227, N11727);
and AND2 (N23239, N23233, N10907);
not NOT1 (N23240, N23232);
or OR2 (N23241, N23216, N11551);
not NOT1 (N23242, N23237);
xor XOR2 (N23243, N23212, N6031);
nor NOR3 (N23244, N23239, N9409, N20382);
and AND2 (N23245, N23219, N3957);
or OR3 (N23246, N23245, N5498, N19295);
buf BUF1 (N23247, N23240);
buf BUF1 (N23248, N23241);
xor XOR2 (N23249, N23229, N20149);
or OR2 (N23250, N23231, N11668);
not NOT1 (N23251, N23243);
or OR3 (N23252, N23250, N7691, N10354);
xor XOR2 (N23253, N23246, N1710);
not NOT1 (N23254, N23242);
and AND2 (N23255, N23236, N17234);
buf BUF1 (N23256, N23247);
buf BUF1 (N23257, N23238);
buf BUF1 (N23258, N23244);
not NOT1 (N23259, N23253);
or OR2 (N23260, N23249, N13874);
buf BUF1 (N23261, N23256);
and AND3 (N23262, N23257, N15715, N8069);
nor NOR3 (N23263, N23262, N20985, N11196);
not NOT1 (N23264, N23255);
not NOT1 (N23265, N23251);
nand NAND4 (N23266, N23259, N13103, N7343, N622);
nand NAND3 (N23267, N23266, N2648, N21802);
nand NAND3 (N23268, N23248, N11047, N13024);
nand NAND3 (N23269, N23265, N14882, N10320);
buf BUF1 (N23270, N23267);
not NOT1 (N23271, N23254);
xor XOR2 (N23272, N23264, N3281);
and AND2 (N23273, N23269, N6448);
nand NAND4 (N23274, N23272, N2103, N14730, N12930);
not NOT1 (N23275, N23260);
not NOT1 (N23276, N23274);
and AND3 (N23277, N23270, N21113, N18120);
buf BUF1 (N23278, N23263);
nor NOR2 (N23279, N23277, N19155);
nand NAND3 (N23280, N23278, N17016, N11987);
buf BUF1 (N23281, N23271);
xor XOR2 (N23282, N23258, N9701);
not NOT1 (N23283, N23275);
and AND3 (N23284, N23252, N13055, N21148);
nor NOR2 (N23285, N23261, N2039);
and AND3 (N23286, N23284, N14471, N22078);
xor XOR2 (N23287, N23282, N13540);
buf BUF1 (N23288, N23286);
and AND3 (N23289, N23287, N8161, N9436);
xor XOR2 (N23290, N23288, N20862);
not NOT1 (N23291, N23276);
xor XOR2 (N23292, N23291, N10130);
and AND3 (N23293, N23268, N13432, N20766);
or OR3 (N23294, N23279, N9927, N18475);
and AND2 (N23295, N23289, N4193);
nand NAND3 (N23296, N23285, N18980, N16863);
buf BUF1 (N23297, N23296);
nor NOR2 (N23298, N23290, N16103);
or OR4 (N23299, N23280, N13443, N12866, N12227);
not NOT1 (N23300, N23292);
buf BUF1 (N23301, N23300);
xor XOR2 (N23302, N23297, N17796);
buf BUF1 (N23303, N23294);
or OR4 (N23304, N23298, N19377, N12636, N18495);
nor NOR2 (N23305, N23303, N4761);
nor NOR3 (N23306, N23301, N16960, N20808);
or OR3 (N23307, N23305, N14846, N14464);
not NOT1 (N23308, N23302);
buf BUF1 (N23309, N23306);
nand NAND2 (N23310, N23293, N5611);
nand NAND2 (N23311, N23307, N17714);
nand NAND3 (N23312, N23273, N12548, N4685);
or OR3 (N23313, N23283, N18947, N13906);
not NOT1 (N23314, N23308);
and AND3 (N23315, N23312, N12813, N5061);
buf BUF1 (N23316, N23315);
or OR4 (N23317, N23314, N16123, N7751, N5853);
nor NOR2 (N23318, N23310, N21584);
nand NAND3 (N23319, N23311, N23122, N19887);
or OR4 (N23320, N23309, N13083, N1958, N1396);
buf BUF1 (N23321, N23318);
nor NOR4 (N23322, N23281, N3121, N17121, N8239);
buf BUF1 (N23323, N23319);
not NOT1 (N23324, N23313);
and AND3 (N23325, N23321, N20440, N18384);
not NOT1 (N23326, N23322);
or OR4 (N23327, N23316, N7217, N3245, N6027);
or OR4 (N23328, N23326, N4720, N9487, N3489);
not NOT1 (N23329, N23304);
xor XOR2 (N23330, N23295, N7510);
nand NAND4 (N23331, N23328, N8945, N16986, N16981);
nand NAND2 (N23332, N23323, N11253);
or OR4 (N23333, N23324, N15909, N214, N12843);
and AND4 (N23334, N23325, N16937, N17673, N6363);
or OR3 (N23335, N23333, N10848, N513);
and AND2 (N23336, N23331, N11175);
or OR2 (N23337, N23330, N8968);
not NOT1 (N23338, N23335);
nor NOR2 (N23339, N23332, N7905);
nand NAND4 (N23340, N23338, N9335, N13333, N10562);
not NOT1 (N23341, N23334);
or OR2 (N23342, N23299, N5593);
or OR4 (N23343, N23327, N2127, N22592, N17345);
nor NOR3 (N23344, N23320, N13972, N866);
nor NOR2 (N23345, N23339, N18434);
or OR4 (N23346, N23329, N11526, N16533, N20355);
or OR2 (N23347, N23344, N21661);
not NOT1 (N23348, N23341);
and AND2 (N23349, N23346, N3324);
not NOT1 (N23350, N23345);
buf BUF1 (N23351, N23317);
nand NAND4 (N23352, N23342, N19309, N18864, N4762);
not NOT1 (N23353, N23350);
buf BUF1 (N23354, N23343);
xor XOR2 (N23355, N23353, N3862);
nand NAND2 (N23356, N23355, N16105);
xor XOR2 (N23357, N23349, N6719);
nor NOR2 (N23358, N23340, N1515);
or OR4 (N23359, N23356, N18700, N16516, N6204);
not NOT1 (N23360, N23352);
and AND4 (N23361, N23359, N19213, N22392, N13427);
buf BUF1 (N23362, N23357);
and AND4 (N23363, N23362, N19289, N18340, N22654);
and AND3 (N23364, N23336, N14286, N8082);
buf BUF1 (N23365, N23347);
nor NOR4 (N23366, N23365, N648, N21673, N4661);
buf BUF1 (N23367, N23361);
buf BUF1 (N23368, N23358);
buf BUF1 (N23369, N23354);
buf BUF1 (N23370, N23360);
and AND3 (N23371, N23337, N15662, N17288);
nor NOR4 (N23372, N23348, N435, N20282, N1785);
nand NAND2 (N23373, N23363, N16946);
buf BUF1 (N23374, N23369);
and AND3 (N23375, N23374, N16665, N983);
not NOT1 (N23376, N23364);
nand NAND4 (N23377, N23367, N22445, N9546, N20676);
nand NAND4 (N23378, N23373, N17174, N2790, N17603);
buf BUF1 (N23379, N23378);
nor NOR3 (N23380, N23372, N22295, N18473);
xor XOR2 (N23381, N23351, N16511);
xor XOR2 (N23382, N23370, N3854);
buf BUF1 (N23383, N23366);
nand NAND2 (N23384, N23380, N11388);
and AND3 (N23385, N23381, N17103, N16623);
xor XOR2 (N23386, N23383, N2379);
xor XOR2 (N23387, N23371, N4538);
or OR2 (N23388, N23376, N5757);
not NOT1 (N23389, N23382);
and AND3 (N23390, N23384, N2972, N20047);
nor NOR3 (N23391, N23379, N17962, N15148);
and AND3 (N23392, N23368, N2160, N8992);
and AND4 (N23393, N23390, N17870, N12311, N18994);
xor XOR2 (N23394, N23388, N10863);
not NOT1 (N23395, N23377);
not NOT1 (N23396, N23392);
not NOT1 (N23397, N23396);
or OR4 (N23398, N23386, N8869, N18982, N3357);
nand NAND4 (N23399, N23375, N1741, N5528, N1933);
nand NAND2 (N23400, N23399, N2413);
or OR4 (N23401, N23391, N17869, N7569, N17141);
nor NOR4 (N23402, N23400, N21755, N8665, N13724);
or OR4 (N23403, N23387, N17696, N3759, N7917);
and AND2 (N23404, N23403, N9499);
nand NAND2 (N23405, N23398, N19073);
or OR2 (N23406, N23404, N9217);
nand NAND4 (N23407, N23393, N692, N13148, N14499);
and AND3 (N23408, N23397, N19175, N2131);
buf BUF1 (N23409, N23407);
nor NOR4 (N23410, N23394, N6927, N15210, N21778);
nand NAND3 (N23411, N23405, N8936, N8163);
xor XOR2 (N23412, N23410, N2723);
not NOT1 (N23413, N23385);
not NOT1 (N23414, N23402);
not NOT1 (N23415, N23395);
nand NAND3 (N23416, N23411, N11429, N18225);
buf BUF1 (N23417, N23416);
not NOT1 (N23418, N23417);
and AND3 (N23419, N23414, N6765, N2672);
nand NAND2 (N23420, N23401, N22575);
buf BUF1 (N23421, N23419);
buf BUF1 (N23422, N23406);
or OR4 (N23423, N23409, N6114, N20990, N7385);
nor NOR2 (N23424, N23423, N9790);
nor NOR2 (N23425, N23415, N22141);
xor XOR2 (N23426, N23425, N9691);
nand NAND4 (N23427, N23408, N4996, N22764, N2545);
nand NAND3 (N23428, N23424, N5980, N18372);
xor XOR2 (N23429, N23421, N18060);
nor NOR4 (N23430, N23429, N1013, N9266, N13618);
and AND2 (N23431, N23422, N7338);
and AND3 (N23432, N23427, N5912, N6092);
nor NOR2 (N23433, N23432, N14018);
xor XOR2 (N23434, N23420, N7829);
nor NOR3 (N23435, N23433, N2551, N21079);
not NOT1 (N23436, N23428);
or OR4 (N23437, N23413, N5893, N7013, N9727);
nand NAND3 (N23438, N23412, N8322, N633);
not NOT1 (N23439, N23430);
and AND2 (N23440, N23435, N16401);
or OR4 (N23441, N23434, N9106, N14968, N4932);
and AND4 (N23442, N23426, N15022, N14, N10512);
or OR4 (N23443, N23442, N9319, N14489, N23230);
nand NAND2 (N23444, N23441, N12799);
not NOT1 (N23445, N23431);
or OR2 (N23446, N23436, N16561);
xor XOR2 (N23447, N23446, N18380);
nand NAND3 (N23448, N23389, N15972, N11870);
xor XOR2 (N23449, N23438, N21436);
or OR2 (N23450, N23418, N6664);
nor NOR3 (N23451, N23444, N13224, N839);
buf BUF1 (N23452, N23437);
nor NOR3 (N23453, N23451, N21072, N3590);
not NOT1 (N23454, N23449);
not NOT1 (N23455, N23440);
not NOT1 (N23456, N23450);
not NOT1 (N23457, N23439);
not NOT1 (N23458, N23453);
or OR3 (N23459, N23458, N9642, N842);
not NOT1 (N23460, N23455);
not NOT1 (N23461, N23447);
buf BUF1 (N23462, N23456);
and AND2 (N23463, N23452, N22496);
xor XOR2 (N23464, N23445, N11728);
not NOT1 (N23465, N23459);
nor NOR2 (N23466, N23464, N15776);
nor NOR3 (N23467, N23466, N2296, N16375);
or OR2 (N23468, N23465, N1580);
or OR3 (N23469, N23454, N20651, N3758);
nand NAND4 (N23470, N23460, N21350, N11108, N19063);
or OR4 (N23471, N23470, N9315, N18992, N13329);
nor NOR4 (N23472, N23468, N19396, N21711, N2314);
or OR3 (N23473, N23457, N18831, N8612);
nand NAND4 (N23474, N23472, N19647, N14564, N11878);
nor NOR4 (N23475, N23443, N22988, N15609, N17088);
xor XOR2 (N23476, N23473, N22656);
not NOT1 (N23477, N23462);
and AND4 (N23478, N23461, N15686, N16914, N11123);
not NOT1 (N23479, N23474);
or OR2 (N23480, N23475, N15447);
and AND2 (N23481, N23448, N1875);
not NOT1 (N23482, N23469);
buf BUF1 (N23483, N23481);
xor XOR2 (N23484, N23476, N20006);
and AND4 (N23485, N23478, N10698, N7762, N4566);
nor NOR4 (N23486, N23467, N9910, N16082, N16503);
or OR3 (N23487, N23463, N1050, N13503);
or OR4 (N23488, N23484, N1159, N22072, N11095);
nand NAND2 (N23489, N23488, N14500);
buf BUF1 (N23490, N23489);
buf BUF1 (N23491, N23482);
buf BUF1 (N23492, N23487);
nand NAND2 (N23493, N23483, N11266);
nand NAND4 (N23494, N23480, N12918, N3198, N4798);
nand NAND2 (N23495, N23477, N17021);
and AND3 (N23496, N23495, N14138, N12586);
nor NOR4 (N23497, N23479, N13335, N4923, N6349);
and AND3 (N23498, N23485, N7101, N5164);
and AND3 (N23499, N23497, N14287, N13359);
or OR3 (N23500, N23499, N7034, N22467);
xor XOR2 (N23501, N23490, N4460);
buf BUF1 (N23502, N23496);
or OR4 (N23503, N23492, N6378, N4286, N19207);
xor XOR2 (N23504, N23502, N21879);
xor XOR2 (N23505, N23471, N21810);
buf BUF1 (N23506, N23505);
nand NAND2 (N23507, N23503, N20097);
and AND4 (N23508, N23493, N13574, N17110, N18198);
or OR3 (N23509, N23507, N12495, N23427);
xor XOR2 (N23510, N23501, N22925);
nor NOR4 (N23511, N23506, N4019, N2144, N1363);
nand NAND4 (N23512, N23511, N17922, N15502, N1948);
and AND2 (N23513, N23504, N6935);
xor XOR2 (N23514, N23512, N16040);
nor NOR4 (N23515, N23514, N16212, N8674, N19445);
xor XOR2 (N23516, N23510, N12762);
not NOT1 (N23517, N23508);
or OR3 (N23518, N23500, N21765, N20302);
buf BUF1 (N23519, N23517);
xor XOR2 (N23520, N23491, N403);
xor XOR2 (N23521, N23494, N11988);
or OR4 (N23522, N23521, N12786, N22006, N18607);
nand NAND3 (N23523, N23498, N7616, N13724);
not NOT1 (N23524, N23486);
or OR4 (N23525, N23516, N5295, N386, N9136);
nand NAND4 (N23526, N23523, N20732, N17809, N6946);
not NOT1 (N23527, N23515);
nor NOR3 (N23528, N23525, N19583, N1041);
or OR3 (N23529, N23518, N17841, N22917);
nand NAND2 (N23530, N23527, N16237);
buf BUF1 (N23531, N23522);
or OR2 (N23532, N23520, N2629);
nand NAND2 (N23533, N23526, N19120);
not NOT1 (N23534, N23531);
or OR4 (N23535, N23509, N23422, N16640, N22533);
buf BUF1 (N23536, N23513);
or OR4 (N23537, N23536, N19977, N2117, N1953);
or OR4 (N23538, N23537, N20240, N17491, N16249);
nor NOR4 (N23539, N23535, N5033, N21456, N362);
buf BUF1 (N23540, N23533);
and AND2 (N23541, N23528, N10835);
buf BUF1 (N23542, N23539);
or OR2 (N23543, N23529, N23078);
xor XOR2 (N23544, N23519, N14673);
or OR2 (N23545, N23538, N20393);
not NOT1 (N23546, N23545);
nand NAND4 (N23547, N23544, N15369, N9823, N18973);
nor NOR3 (N23548, N23524, N14348, N17043);
xor XOR2 (N23549, N23530, N9103);
nand NAND4 (N23550, N23540, N578, N13461, N21929);
not NOT1 (N23551, N23547);
xor XOR2 (N23552, N23548, N17863);
xor XOR2 (N23553, N23550, N3296);
buf BUF1 (N23554, N23532);
or OR2 (N23555, N23546, N11858);
or OR3 (N23556, N23549, N23090, N13896);
not NOT1 (N23557, N23543);
xor XOR2 (N23558, N23552, N19326);
nand NAND4 (N23559, N23541, N11706, N12395, N12549);
and AND2 (N23560, N23534, N11092);
or OR2 (N23561, N23553, N5575);
nor NOR4 (N23562, N23558, N7227, N76, N2397);
nor NOR3 (N23563, N23542, N21, N15193);
xor XOR2 (N23564, N23560, N7479);
buf BUF1 (N23565, N23554);
and AND3 (N23566, N23563, N22499, N12852);
and AND4 (N23567, N23562, N6074, N10956, N19869);
nand NAND3 (N23568, N23561, N12072, N10438);
buf BUF1 (N23569, N23559);
not NOT1 (N23570, N23565);
and AND3 (N23571, N23567, N11788, N15980);
buf BUF1 (N23572, N23564);
buf BUF1 (N23573, N23551);
and AND2 (N23574, N23566, N5523);
not NOT1 (N23575, N23570);
and AND3 (N23576, N23572, N9904, N21379);
and AND2 (N23577, N23571, N11607);
nor NOR2 (N23578, N23576, N22906);
and AND3 (N23579, N23573, N21518, N8508);
xor XOR2 (N23580, N23568, N23515);
buf BUF1 (N23581, N23580);
buf BUF1 (N23582, N23574);
buf BUF1 (N23583, N23555);
nand NAND3 (N23584, N23556, N2973, N4552);
nor NOR2 (N23585, N23569, N3988);
nor NOR4 (N23586, N23579, N16297, N16269, N16862);
buf BUF1 (N23587, N23581);
nor NOR4 (N23588, N23577, N11521, N19278, N7880);
nor NOR4 (N23589, N23582, N1152, N12515, N13828);
nor NOR2 (N23590, N23586, N17210);
xor XOR2 (N23591, N23585, N17797);
buf BUF1 (N23592, N23575);
and AND3 (N23593, N23557, N18226, N19551);
xor XOR2 (N23594, N23589, N3894);
or OR4 (N23595, N23593, N18836, N8022, N23525);
and AND4 (N23596, N23594, N8609, N727, N2472);
xor XOR2 (N23597, N23596, N3139);
buf BUF1 (N23598, N23591);
not NOT1 (N23599, N23588);
nand NAND4 (N23600, N23599, N15815, N14445, N5776);
not NOT1 (N23601, N23592);
nor NOR4 (N23602, N23601, N22708, N21771, N15424);
nand NAND2 (N23603, N23587, N15006);
nand NAND3 (N23604, N23597, N12525, N11648);
buf BUF1 (N23605, N23578);
and AND3 (N23606, N23584, N18304, N5830);
and AND3 (N23607, N23600, N16724, N22988);
nor NOR4 (N23608, N23603, N6838, N21018, N5422);
xor XOR2 (N23609, N23604, N3237);
or OR2 (N23610, N23598, N5361);
buf BUF1 (N23611, N23595);
nand NAND3 (N23612, N23610, N20726, N12355);
nand NAND2 (N23613, N23590, N21087);
xor XOR2 (N23614, N23613, N6741);
nor NOR2 (N23615, N23605, N12233);
and AND3 (N23616, N23583, N9883, N3994);
nand NAND4 (N23617, N23614, N19216, N9352, N3307);
and AND3 (N23618, N23617, N19229, N15773);
xor XOR2 (N23619, N23616, N13874);
nand NAND3 (N23620, N23612, N490, N13859);
nor NOR4 (N23621, N23607, N9297, N14605, N15259);
not NOT1 (N23622, N23602);
and AND3 (N23623, N23608, N390, N20325);
nor NOR4 (N23624, N23620, N21759, N2861, N20819);
not NOT1 (N23625, N23609);
and AND4 (N23626, N23622, N16278, N10177, N11881);
buf BUF1 (N23627, N23618);
xor XOR2 (N23628, N23606, N16701);
xor XOR2 (N23629, N23619, N18683);
buf BUF1 (N23630, N23628);
nor NOR2 (N23631, N23626, N10834);
buf BUF1 (N23632, N23629);
buf BUF1 (N23633, N23611);
xor XOR2 (N23634, N23633, N8340);
buf BUF1 (N23635, N23627);
xor XOR2 (N23636, N23623, N19192);
xor XOR2 (N23637, N23625, N10110);
nor NOR2 (N23638, N23615, N4592);
and AND4 (N23639, N23635, N14305, N13169, N6170);
nand NAND4 (N23640, N23624, N22042, N18409, N4914);
nand NAND4 (N23641, N23632, N13800, N20130, N16363);
not NOT1 (N23642, N23636);
nand NAND4 (N23643, N23631, N11388, N10629, N10947);
and AND4 (N23644, N23641, N19729, N2045, N9657);
not NOT1 (N23645, N23639);
xor XOR2 (N23646, N23643, N1044);
or OR4 (N23647, N23644, N17067, N6742, N18911);
nand NAND3 (N23648, N23621, N5913, N9339);
nor NOR2 (N23649, N23638, N11801);
buf BUF1 (N23650, N23637);
xor XOR2 (N23651, N23640, N11567);
nand NAND3 (N23652, N23646, N2875, N19698);
xor XOR2 (N23653, N23648, N14186);
xor XOR2 (N23654, N23642, N21170);
buf BUF1 (N23655, N23649);
and AND2 (N23656, N23630, N13979);
xor XOR2 (N23657, N23654, N18944);
nor NOR2 (N23658, N23656, N2830);
nand NAND4 (N23659, N23657, N10080, N7252, N21425);
or OR3 (N23660, N23653, N10857, N20174);
xor XOR2 (N23661, N23650, N1526);
or OR4 (N23662, N23655, N18829, N4136, N18233);
nand NAND2 (N23663, N23658, N5800);
and AND3 (N23664, N23634, N6660, N20499);
nand NAND3 (N23665, N23645, N20717, N14592);
buf BUF1 (N23666, N23663);
and AND4 (N23667, N23665, N23308, N11914, N20151);
buf BUF1 (N23668, N23662);
buf BUF1 (N23669, N23661);
buf BUF1 (N23670, N23666);
xor XOR2 (N23671, N23667, N18119);
buf BUF1 (N23672, N23651);
nor NOR4 (N23673, N23647, N18169, N21661, N17749);
not NOT1 (N23674, N23670);
not NOT1 (N23675, N23672);
xor XOR2 (N23676, N23674, N21870);
or OR2 (N23677, N23660, N22146);
nand NAND3 (N23678, N23652, N7359, N16358);
xor XOR2 (N23679, N23675, N6227);
or OR3 (N23680, N23676, N17509, N14319);
nor NOR3 (N23681, N23673, N1468, N15336);
and AND2 (N23682, N23664, N23001);
xor XOR2 (N23683, N23677, N23148);
nand NAND3 (N23684, N23683, N5999, N17203);
or OR3 (N23685, N23659, N7756, N19157);
not NOT1 (N23686, N23669);
not NOT1 (N23687, N23685);
and AND2 (N23688, N23671, N18713);
not NOT1 (N23689, N23684);
and AND2 (N23690, N23680, N12134);
or OR2 (N23691, N23687, N14797);
and AND4 (N23692, N23668, N1973, N8404, N22090);
nor NOR2 (N23693, N23681, N19267);
nor NOR2 (N23694, N23692, N11722);
not NOT1 (N23695, N23682);
or OR3 (N23696, N23693, N8790, N6287);
and AND2 (N23697, N23690, N17063);
buf BUF1 (N23698, N23697);
buf BUF1 (N23699, N23691);
nor NOR2 (N23700, N23686, N6134);
or OR3 (N23701, N23699, N3105, N11203);
or OR2 (N23702, N23696, N12149);
xor XOR2 (N23703, N23689, N11265);
nand NAND3 (N23704, N23703, N12585, N22607);
and AND2 (N23705, N23679, N9119);
buf BUF1 (N23706, N23704);
and AND3 (N23707, N23698, N23265, N15494);
nor NOR2 (N23708, N23702, N12395);
xor XOR2 (N23709, N23705, N17638);
xor XOR2 (N23710, N23694, N5306);
nor NOR2 (N23711, N23709, N13168);
nor NOR2 (N23712, N23711, N5590);
nand NAND2 (N23713, N23695, N857);
or OR3 (N23714, N23713, N215, N20661);
buf BUF1 (N23715, N23706);
nor NOR4 (N23716, N23714, N19090, N5255, N503);
nand NAND3 (N23717, N23712, N17353, N694);
or OR4 (N23718, N23716, N8100, N15598, N9497);
nand NAND4 (N23719, N23700, N17847, N8234, N10005);
xor XOR2 (N23720, N23678, N3684);
and AND3 (N23721, N23720, N3074, N20713);
or OR2 (N23722, N23715, N22226);
nor NOR2 (N23723, N23718, N3666);
xor XOR2 (N23724, N23701, N736);
nand NAND2 (N23725, N23708, N5113);
nand NAND3 (N23726, N23688, N3517, N1243);
nor NOR4 (N23727, N23719, N23599, N18724, N9966);
and AND4 (N23728, N23710, N20586, N4050, N8467);
nor NOR2 (N23729, N23723, N13713);
or OR4 (N23730, N23725, N3219, N1517, N11266);
xor XOR2 (N23731, N23729, N21325);
nor NOR4 (N23732, N23707, N5398, N17884, N18501);
or OR2 (N23733, N23717, N21833);
buf BUF1 (N23734, N23733);
not NOT1 (N23735, N23734);
and AND4 (N23736, N23731, N134, N15099, N1810);
xor XOR2 (N23737, N23727, N7409);
buf BUF1 (N23738, N23721);
nor NOR2 (N23739, N23738, N18141);
nand NAND3 (N23740, N23728, N520, N20607);
nand NAND2 (N23741, N23739, N14171);
and AND2 (N23742, N23732, N4670);
or OR3 (N23743, N23730, N23545, N8311);
xor XOR2 (N23744, N23742, N16484);
and AND3 (N23745, N23736, N3126, N23723);
and AND2 (N23746, N23735, N6742);
and AND3 (N23747, N23743, N8840, N10054);
not NOT1 (N23748, N23740);
and AND2 (N23749, N23726, N6177);
xor XOR2 (N23750, N23745, N22195);
not NOT1 (N23751, N23749);
not NOT1 (N23752, N23722);
nand NAND2 (N23753, N23748, N8536);
nor NOR4 (N23754, N23751, N19472, N9107, N14230);
nand NAND4 (N23755, N23750, N5160, N1635, N3180);
and AND4 (N23756, N23754, N21323, N17973, N20822);
nor NOR3 (N23757, N23753, N21937, N10607);
nor NOR4 (N23758, N23756, N7582, N20034, N1384);
nand NAND3 (N23759, N23752, N20071, N8016);
xor XOR2 (N23760, N23758, N13521);
nor NOR2 (N23761, N23757, N22239);
and AND4 (N23762, N23746, N4258, N8064, N1514);
buf BUF1 (N23763, N23724);
xor XOR2 (N23764, N23759, N12814);
and AND3 (N23765, N23755, N17939, N4957);
or OR3 (N23766, N23763, N4478, N19058);
not NOT1 (N23767, N23766);
buf BUF1 (N23768, N23764);
nor NOR4 (N23769, N23761, N18194, N17757, N3294);
xor XOR2 (N23770, N23747, N16887);
buf BUF1 (N23771, N23765);
xor XOR2 (N23772, N23737, N5323);
xor XOR2 (N23773, N23744, N1007);
and AND3 (N23774, N23770, N16846, N11924);
or OR3 (N23775, N23767, N21394, N5656);
nor NOR4 (N23776, N23741, N7900, N15667, N22898);
and AND3 (N23777, N23762, N20914, N22960);
xor XOR2 (N23778, N23773, N7184);
nor NOR2 (N23779, N23760, N3897);
buf BUF1 (N23780, N23779);
and AND3 (N23781, N23772, N21683, N18197);
nor NOR3 (N23782, N23769, N18951, N3331);
not NOT1 (N23783, N23774);
nand NAND3 (N23784, N23775, N12480, N9274);
nor NOR2 (N23785, N23784, N10952);
not NOT1 (N23786, N23781);
not NOT1 (N23787, N23768);
not NOT1 (N23788, N23785);
nand NAND3 (N23789, N23783, N6665, N13909);
nor NOR4 (N23790, N23786, N4312, N4819, N23660);
and AND4 (N23791, N23777, N18786, N12367, N22420);
nand NAND3 (N23792, N23778, N7544, N19790);
buf BUF1 (N23793, N23790);
not NOT1 (N23794, N23787);
buf BUF1 (N23795, N23794);
nor NOR4 (N23796, N23792, N8599, N18705, N981);
nand NAND3 (N23797, N23793, N8428, N9597);
xor XOR2 (N23798, N23789, N20607);
nand NAND4 (N23799, N23788, N17628, N9509, N8451);
not NOT1 (N23800, N23799);
not NOT1 (N23801, N23795);
xor XOR2 (N23802, N23797, N340);
buf BUF1 (N23803, N23798);
nand NAND4 (N23804, N23800, N3830, N19665, N20469);
not NOT1 (N23805, N23780);
nand NAND3 (N23806, N23804, N5879, N1464);
nor NOR2 (N23807, N23771, N9614);
nor NOR2 (N23808, N23807, N2981);
buf BUF1 (N23809, N23805);
and AND2 (N23810, N23808, N16238);
and AND4 (N23811, N23810, N16546, N2645, N17521);
nor NOR3 (N23812, N23796, N4549, N12247);
nor NOR4 (N23813, N23782, N22428, N11709, N10243);
nand NAND4 (N23814, N23812, N3874, N509, N4932);
and AND3 (N23815, N23814, N10131, N4671);
or OR4 (N23816, N23803, N9167, N4525, N20581);
and AND4 (N23817, N23816, N20462, N18101, N14450);
and AND3 (N23818, N23801, N13264, N18660);
nor NOR3 (N23819, N23791, N23378, N4511);
and AND3 (N23820, N23802, N17527, N21502);
buf BUF1 (N23821, N23820);
nor NOR2 (N23822, N23806, N18589);
or OR2 (N23823, N23818, N2322);
or OR2 (N23824, N23819, N3882);
nor NOR2 (N23825, N23821, N23781);
buf BUF1 (N23826, N23823);
and AND2 (N23827, N23776, N19284);
or OR3 (N23828, N23815, N7946, N8885);
nor NOR4 (N23829, N23813, N6554, N2026, N23281);
not NOT1 (N23830, N23828);
or OR2 (N23831, N23830, N8113);
xor XOR2 (N23832, N23817, N22820);
nand NAND4 (N23833, N23809, N20852, N1661, N8484);
or OR2 (N23834, N23811, N3653);
and AND4 (N23835, N23829, N18165, N18145, N12988);
buf BUF1 (N23836, N23824);
buf BUF1 (N23837, N23832);
xor XOR2 (N23838, N23837, N21517);
nor NOR2 (N23839, N23834, N18175);
nor NOR2 (N23840, N23831, N15208);
buf BUF1 (N23841, N23839);
nand NAND3 (N23842, N23826, N5051, N95);
xor XOR2 (N23843, N23835, N13707);
xor XOR2 (N23844, N23833, N14800);
nand NAND4 (N23845, N23822, N12698, N10356, N17134);
buf BUF1 (N23846, N23841);
not NOT1 (N23847, N23846);
or OR4 (N23848, N23847, N23357, N18938, N18833);
buf BUF1 (N23849, N23840);
or OR3 (N23850, N23844, N13782, N14766);
xor XOR2 (N23851, N23838, N5500);
xor XOR2 (N23852, N23827, N8238);
and AND3 (N23853, N23845, N17379, N347);
or OR4 (N23854, N23843, N22583, N4673, N12272);
buf BUF1 (N23855, N23825);
nand NAND4 (N23856, N23854, N21101, N7149, N21003);
nand NAND2 (N23857, N23851, N1217);
xor XOR2 (N23858, N23848, N6599);
not NOT1 (N23859, N23856);
or OR3 (N23860, N23859, N12224, N23853);
nor NOR4 (N23861, N11780, N8385, N7856, N14179);
or OR4 (N23862, N23849, N4656, N54, N16727);
xor XOR2 (N23863, N23842, N20488);
nor NOR2 (N23864, N23858, N8637);
buf BUF1 (N23865, N23860);
nand NAND4 (N23866, N23865, N1721, N12662, N23718);
not NOT1 (N23867, N23850);
not NOT1 (N23868, N23862);
not NOT1 (N23869, N23855);
nand NAND3 (N23870, N23861, N7577, N9968);
nor NOR3 (N23871, N23863, N23784, N7439);
nor NOR4 (N23872, N23867, N8112, N12910, N6071);
not NOT1 (N23873, N23866);
nor NOR4 (N23874, N23836, N2352, N7200, N6411);
buf BUF1 (N23875, N23869);
xor XOR2 (N23876, N23875, N2977);
xor XOR2 (N23877, N23868, N289);
nand NAND3 (N23878, N23874, N6161, N6338);
xor XOR2 (N23879, N23876, N1799);
xor XOR2 (N23880, N23877, N7515);
nand NAND3 (N23881, N23852, N11942, N21218);
buf BUF1 (N23882, N23881);
buf BUF1 (N23883, N23870);
or OR4 (N23884, N23882, N22923, N21143, N19179);
nand NAND3 (N23885, N23880, N21910, N18775);
and AND2 (N23886, N23883, N1914);
buf BUF1 (N23887, N23857);
nor NOR2 (N23888, N23871, N344);
and AND2 (N23889, N23879, N8815);
not NOT1 (N23890, N23886);
or OR4 (N23891, N23887, N10706, N8567, N5897);
and AND2 (N23892, N23890, N16895);
buf BUF1 (N23893, N23889);
buf BUF1 (N23894, N23893);
nand NAND4 (N23895, N23864, N19536, N17918, N15);
buf BUF1 (N23896, N23872);
not NOT1 (N23897, N23888);
xor XOR2 (N23898, N23895, N5333);
nor NOR4 (N23899, N23896, N8017, N20605, N2328);
buf BUF1 (N23900, N23878);
xor XOR2 (N23901, N23884, N3638);
nor NOR3 (N23902, N23894, N17637, N5017);
and AND2 (N23903, N23900, N10804);
xor XOR2 (N23904, N23873, N15300);
and AND4 (N23905, N23891, N3089, N13006, N16979);
and AND2 (N23906, N23904, N6768);
not NOT1 (N23907, N23899);
or OR2 (N23908, N23901, N20866);
nor NOR3 (N23909, N23903, N577, N16175);
nor NOR4 (N23910, N23892, N21685, N11676, N2475);
xor XOR2 (N23911, N23902, N583);
nor NOR3 (N23912, N23906, N3937, N15529);
and AND2 (N23913, N23908, N1925);
buf BUF1 (N23914, N23909);
nor NOR4 (N23915, N23897, N11467, N9751, N23709);
not NOT1 (N23916, N23912);
not NOT1 (N23917, N23913);
xor XOR2 (N23918, N23915, N3362);
or OR3 (N23919, N23916, N16549, N14567);
nor NOR4 (N23920, N23898, N11611, N2685, N23850);
not NOT1 (N23921, N23920);
buf BUF1 (N23922, N23914);
buf BUF1 (N23923, N23922);
nor NOR4 (N23924, N23905, N7385, N22429, N22104);
buf BUF1 (N23925, N23921);
not NOT1 (N23926, N23923);
and AND2 (N23927, N23925, N8135);
and AND4 (N23928, N23926, N14324, N14627, N17345);
not NOT1 (N23929, N23917);
nand NAND2 (N23930, N23929, N8228);
or OR3 (N23931, N23907, N17480, N20359);
xor XOR2 (N23932, N23930, N7529);
not NOT1 (N23933, N23885);
and AND3 (N23934, N23928, N13374, N11751);
buf BUF1 (N23935, N23933);
nand NAND4 (N23936, N23910, N1766, N5287, N16063);
nand NAND4 (N23937, N23919, N4817, N21347, N8585);
and AND2 (N23938, N23937, N4607);
or OR4 (N23939, N23935, N12404, N19154, N18504);
buf BUF1 (N23940, N23924);
buf BUF1 (N23941, N23931);
xor XOR2 (N23942, N23940, N22839);
nor NOR2 (N23943, N23941, N4214);
xor XOR2 (N23944, N23942, N14351);
nand NAND3 (N23945, N23939, N20847, N16714);
and AND2 (N23946, N23932, N17150);
nand NAND3 (N23947, N23938, N9704, N23423);
buf BUF1 (N23948, N23927);
xor XOR2 (N23949, N23947, N2659);
or OR3 (N23950, N23945, N801, N2290);
and AND4 (N23951, N23943, N17043, N9773, N5108);
nand NAND3 (N23952, N23934, N20782, N14124);
not NOT1 (N23953, N23911);
nand NAND4 (N23954, N23953, N19629, N10191, N3767);
buf BUF1 (N23955, N23952);
nand NAND3 (N23956, N23955, N7509, N7309);
nor NOR4 (N23957, N23936, N16658, N18745, N19984);
buf BUF1 (N23958, N23949);
buf BUF1 (N23959, N23946);
nand NAND2 (N23960, N23951, N14516);
xor XOR2 (N23961, N23960, N18528);
nor NOR2 (N23962, N23957, N4426);
nand NAND3 (N23963, N23959, N8724, N17548);
or OR2 (N23964, N23944, N9358);
buf BUF1 (N23965, N23958);
buf BUF1 (N23966, N23950);
nor NOR2 (N23967, N23961, N12722);
not NOT1 (N23968, N23954);
not NOT1 (N23969, N23956);
not NOT1 (N23970, N23964);
not NOT1 (N23971, N23962);
xor XOR2 (N23972, N23967, N15921);
or OR3 (N23973, N23918, N13849, N11745);
and AND3 (N23974, N23972, N20597, N17734);
buf BUF1 (N23975, N23965);
not NOT1 (N23976, N23973);
and AND3 (N23977, N23971, N14312, N3336);
not NOT1 (N23978, N23970);
or OR3 (N23979, N23975, N3329, N4243);
not NOT1 (N23980, N23963);
and AND4 (N23981, N23974, N20558, N19752, N11610);
nand NAND2 (N23982, N23969, N4834);
buf BUF1 (N23983, N23979);
not NOT1 (N23984, N23948);
or OR4 (N23985, N23984, N11689, N1467, N19380);
and AND2 (N23986, N23977, N22604);
xor XOR2 (N23987, N23968, N1711);
buf BUF1 (N23988, N23978);
nand NAND3 (N23989, N23985, N22941, N16153);
nor NOR2 (N23990, N23980, N20798);
or OR3 (N23991, N23986, N14757, N6144);
not NOT1 (N23992, N23982);
not NOT1 (N23993, N23976);
nor NOR2 (N23994, N23990, N16262);
or OR4 (N23995, N23981, N15788, N12172, N15995);
buf BUF1 (N23996, N23992);
xor XOR2 (N23997, N23987, N16873);
xor XOR2 (N23998, N23995, N12252);
xor XOR2 (N23999, N23991, N16804);
xor XOR2 (N24000, N23998, N289);
xor XOR2 (N24001, N23988, N16423);
xor XOR2 (N24002, N23989, N19236);
not NOT1 (N24003, N23993);
nor NOR2 (N24004, N23997, N2161);
nand NAND3 (N24005, N24002, N11450, N7163);
buf BUF1 (N24006, N23983);
and AND2 (N24007, N23966, N23913);
and AND4 (N24008, N24001, N7767, N14034, N12444);
not NOT1 (N24009, N24004);
and AND2 (N24010, N23994, N2714);
buf BUF1 (N24011, N24000);
or OR4 (N24012, N24007, N11097, N17982, N21000);
nor NOR4 (N24013, N24010, N23915, N7111, N21433);
or OR4 (N24014, N23999, N4926, N14789, N7934);
not NOT1 (N24015, N24003);
nor NOR4 (N24016, N24009, N14126, N10719, N11736);
buf BUF1 (N24017, N24013);
buf BUF1 (N24018, N24006);
nand NAND4 (N24019, N23996, N9251, N12593, N8501);
or OR4 (N24020, N24012, N18393, N4902, N21951);
or OR4 (N24021, N24016, N2414, N21821, N6138);
and AND2 (N24022, N24014, N15709);
not NOT1 (N24023, N24019);
not NOT1 (N24024, N24021);
not NOT1 (N24025, N24020);
or OR2 (N24026, N24011, N11685);
nand NAND3 (N24027, N24017, N2297, N9603);
not NOT1 (N24028, N24024);
nor NOR2 (N24029, N24018, N5412);
xor XOR2 (N24030, N24026, N2297);
xor XOR2 (N24031, N24030, N20);
and AND4 (N24032, N24015, N7993, N5072, N4565);
or OR2 (N24033, N24027, N5969);
not NOT1 (N24034, N24028);
nand NAND2 (N24035, N24034, N12056);
xor XOR2 (N24036, N24035, N9899);
xor XOR2 (N24037, N24023, N14402);
nand NAND3 (N24038, N24029, N8989, N224);
and AND4 (N24039, N24032, N329, N13269, N22411);
and AND4 (N24040, N24038, N13922, N20379, N2885);
buf BUF1 (N24041, N24040);
nor NOR4 (N24042, N24036, N15235, N14577, N9400);
and AND4 (N24043, N24008, N15280, N13841, N17494);
xor XOR2 (N24044, N24043, N21516);
nand NAND3 (N24045, N24041, N19162, N2262);
buf BUF1 (N24046, N24037);
nor NOR4 (N24047, N24033, N9770, N3162, N6685);
buf BUF1 (N24048, N24044);
buf BUF1 (N24049, N24045);
xor XOR2 (N24050, N24031, N10343);
and AND4 (N24051, N24048, N20473, N22312, N14229);
xor XOR2 (N24052, N24049, N22078);
nor NOR4 (N24053, N24039, N3555, N4980, N11566);
xor XOR2 (N24054, N24042, N1706);
or OR2 (N24055, N24052, N21580);
nor NOR3 (N24056, N24051, N221, N16790);
or OR4 (N24057, N24046, N19923, N19108, N19729);
and AND4 (N24058, N24054, N13506, N12496, N2486);
xor XOR2 (N24059, N24025, N16571);
nand NAND2 (N24060, N24057, N17301);
nor NOR4 (N24061, N24058, N20779, N12969, N19371);
and AND4 (N24062, N24055, N18961, N13850, N8422);
or OR4 (N24063, N24022, N4977, N22216, N1794);
or OR4 (N24064, N24047, N23211, N5637, N8390);
nor NOR3 (N24065, N24050, N17927, N23346);
xor XOR2 (N24066, N24063, N9360);
not NOT1 (N24067, N24005);
nor NOR4 (N24068, N24059, N3580, N23382, N20871);
xor XOR2 (N24069, N24064, N21575);
or OR3 (N24070, N24060, N2731, N4167);
not NOT1 (N24071, N24070);
nand NAND4 (N24072, N24062, N16191, N9209, N18156);
not NOT1 (N24073, N24069);
and AND4 (N24074, N24071, N19509, N23692, N17650);
buf BUF1 (N24075, N24056);
not NOT1 (N24076, N24068);
xor XOR2 (N24077, N24073, N13244);
not NOT1 (N24078, N24076);
nand NAND2 (N24079, N24061, N5100);
and AND4 (N24080, N24075, N16588, N5514, N10595);
xor XOR2 (N24081, N24077, N10897);
nand NAND2 (N24082, N24080, N7472);
and AND2 (N24083, N24066, N16821);
xor XOR2 (N24084, N24082, N23271);
nor NOR2 (N24085, N24084, N8918);
or OR3 (N24086, N24085, N3895, N7885);
nand NAND3 (N24087, N24081, N22764, N18113);
and AND2 (N24088, N24067, N20371);
xor XOR2 (N24089, N24079, N16063);
or OR4 (N24090, N24088, N8757, N10224, N2917);
xor XOR2 (N24091, N24072, N19937);
or OR2 (N24092, N24065, N21513);
not NOT1 (N24093, N24083);
or OR3 (N24094, N24053, N3965, N12385);
or OR2 (N24095, N24087, N19029);
or OR2 (N24096, N24074, N973);
or OR2 (N24097, N24086, N989);
not NOT1 (N24098, N24089);
nand NAND4 (N24099, N24092, N4937, N19437, N855);
buf BUF1 (N24100, N24096);
or OR4 (N24101, N24097, N19965, N19248, N19852);
or OR4 (N24102, N24090, N16826, N24077, N7093);
or OR2 (N24103, N24098, N15527);
nor NOR4 (N24104, N24094, N9216, N5114, N16233);
not NOT1 (N24105, N24104);
nand NAND2 (N24106, N24101, N4135);
or OR2 (N24107, N24105, N5976);
nor NOR2 (N24108, N24102, N21163);
xor XOR2 (N24109, N24099, N5982);
not NOT1 (N24110, N24091);
not NOT1 (N24111, N24106);
xor XOR2 (N24112, N24108, N19653);
buf BUF1 (N24113, N24110);
xor XOR2 (N24114, N24093, N19690);
nor NOR4 (N24115, N24114, N15967, N4203, N6065);
not NOT1 (N24116, N24112);
nand NAND3 (N24117, N24100, N15310, N14264);
not NOT1 (N24118, N24115);
nor NOR3 (N24119, N24095, N9303, N11200);
xor XOR2 (N24120, N24113, N7284);
or OR4 (N24121, N24116, N2719, N19314, N15014);
nor NOR2 (N24122, N24118, N3200);
nand NAND2 (N24123, N24121, N1827);
buf BUF1 (N24124, N24122);
xor XOR2 (N24125, N24124, N22667);
and AND3 (N24126, N24120, N18809, N10270);
nor NOR3 (N24127, N24123, N6869, N10181);
buf BUF1 (N24128, N24103);
or OR4 (N24129, N24109, N15447, N21227, N3800);
or OR4 (N24130, N24117, N18958, N4692, N7918);
not NOT1 (N24131, N24130);
not NOT1 (N24132, N24078);
nand NAND3 (N24133, N24129, N3621, N19345);
xor XOR2 (N24134, N24133, N14882);
xor XOR2 (N24135, N24134, N950);
and AND3 (N24136, N24111, N7138, N11635);
and AND2 (N24137, N24119, N2109);
xor XOR2 (N24138, N24136, N11462);
nor NOR2 (N24139, N24132, N1312);
nor NOR3 (N24140, N24128, N469, N20657);
or OR2 (N24141, N24140, N15794);
nand NAND2 (N24142, N24131, N4022);
xor XOR2 (N24143, N24139, N5120);
nor NOR4 (N24144, N24107, N1703, N11506, N6045);
or OR2 (N24145, N24126, N6856);
nand NAND2 (N24146, N24127, N8789);
not NOT1 (N24147, N24143);
nand NAND3 (N24148, N24135, N23825, N22016);
buf BUF1 (N24149, N24145);
buf BUF1 (N24150, N24138);
not NOT1 (N24151, N24148);
and AND4 (N24152, N24151, N13101, N10769, N8643);
and AND3 (N24153, N24137, N11130, N23050);
not NOT1 (N24154, N24146);
not NOT1 (N24155, N24141);
nor NOR4 (N24156, N24154, N5523, N22345, N4614);
nand NAND4 (N24157, N24144, N16458, N16129, N22659);
nor NOR3 (N24158, N24147, N20658, N4336);
nand NAND3 (N24159, N24142, N19827, N22808);
buf BUF1 (N24160, N24155);
or OR2 (N24161, N24125, N11089);
nand NAND4 (N24162, N24149, N5050, N16377, N22229);
and AND4 (N24163, N24162, N2375, N15961, N13054);
not NOT1 (N24164, N24161);
not NOT1 (N24165, N24152);
nor NOR4 (N24166, N24159, N15563, N16816, N6288);
not NOT1 (N24167, N24153);
xor XOR2 (N24168, N24160, N5501);
buf BUF1 (N24169, N24164);
or OR3 (N24170, N24165, N3257, N23276);
nor NOR4 (N24171, N24170, N19546, N19937, N50);
xor XOR2 (N24172, N24156, N447);
buf BUF1 (N24173, N24167);
not NOT1 (N24174, N24150);
or OR4 (N24175, N24174, N23903, N2745, N12023);
nand NAND2 (N24176, N24158, N14533);
and AND4 (N24177, N24157, N4222, N6577, N14125);
buf BUF1 (N24178, N24172);
nor NOR4 (N24179, N24166, N14798, N787, N9083);
and AND4 (N24180, N24175, N1057, N22178, N15702);
xor XOR2 (N24181, N24171, N15531);
nor NOR3 (N24182, N24180, N11666, N14286);
nor NOR3 (N24183, N24179, N1262, N20057);
and AND4 (N24184, N24176, N8307, N9549, N20537);
not NOT1 (N24185, N24182);
nand NAND4 (N24186, N24181, N8457, N21369, N18111);
xor XOR2 (N24187, N24168, N15731);
nor NOR4 (N24188, N24186, N19043, N18743, N15233);
nand NAND2 (N24189, N24184, N7725);
buf BUF1 (N24190, N24178);
buf BUF1 (N24191, N24189);
not NOT1 (N24192, N24188);
not NOT1 (N24193, N24173);
and AND3 (N24194, N24183, N13305, N12566);
nand NAND2 (N24195, N24163, N22225);
not NOT1 (N24196, N24177);
nor NOR4 (N24197, N24185, N6025, N12019, N4732);
nor NOR2 (N24198, N24195, N18196);
not NOT1 (N24199, N24198);
not NOT1 (N24200, N24193);
nor NOR2 (N24201, N24187, N13915);
or OR4 (N24202, N24190, N20991, N5463, N21299);
and AND4 (N24203, N24202, N22419, N16575, N17599);
or OR3 (N24204, N24192, N15062, N17945);
xor XOR2 (N24205, N24191, N6276);
xor XOR2 (N24206, N24205, N19993);
and AND2 (N24207, N24197, N1680);
not NOT1 (N24208, N24204);
nor NOR2 (N24209, N24169, N10413);
xor XOR2 (N24210, N24201, N7742);
nand NAND4 (N24211, N24194, N10478, N8322, N5444);
xor XOR2 (N24212, N24199, N14800);
nand NAND4 (N24213, N24209, N15339, N1259, N9682);
xor XOR2 (N24214, N24210, N19047);
and AND3 (N24215, N24211, N19372, N22528);
and AND3 (N24216, N24196, N4679, N23019);
buf BUF1 (N24217, N24203);
nor NOR2 (N24218, N24208, N1369);
or OR4 (N24219, N24207, N21184, N1496, N20707);
nor NOR4 (N24220, N24206, N2598, N20477, N2330);
xor XOR2 (N24221, N24215, N24177);
not NOT1 (N24222, N24214);
not NOT1 (N24223, N24216);
and AND2 (N24224, N24223, N19388);
nor NOR4 (N24225, N24221, N23477, N16665, N16900);
and AND2 (N24226, N24217, N7421);
and AND2 (N24227, N24218, N17265);
not NOT1 (N24228, N24212);
and AND3 (N24229, N24228, N13013, N2015);
and AND3 (N24230, N24229, N424, N10428);
not NOT1 (N24231, N24226);
and AND2 (N24232, N24227, N22238);
and AND4 (N24233, N24231, N6044, N22968, N10834);
nor NOR2 (N24234, N24200, N7304);
and AND3 (N24235, N24233, N20151, N2035);
and AND3 (N24236, N24224, N812, N21974);
nand NAND2 (N24237, N24225, N4579);
nor NOR3 (N24238, N24237, N3651, N15863);
not NOT1 (N24239, N24236);
nand NAND2 (N24240, N24232, N13020);
nor NOR4 (N24241, N24219, N6076, N10781, N4976);
xor XOR2 (N24242, N24230, N21411);
and AND3 (N24243, N24242, N15821, N7852);
xor XOR2 (N24244, N24234, N20189);
nor NOR4 (N24245, N24240, N13793, N10346, N1079);
nand NAND4 (N24246, N24239, N2346, N8332, N12534);
nand NAND4 (N24247, N24243, N15136, N8362, N17912);
nor NOR4 (N24248, N24245, N18363, N6949, N6124);
or OR3 (N24249, N24241, N12459, N13357);
or OR3 (N24250, N24235, N1144, N21196);
and AND2 (N24251, N24246, N2990);
nand NAND3 (N24252, N24251, N20711, N22876);
not NOT1 (N24253, N24250);
nand NAND4 (N24254, N24253, N11656, N10912, N2441);
and AND4 (N24255, N24247, N2554, N22154, N6308);
not NOT1 (N24256, N24213);
or OR3 (N24257, N24222, N11268, N4791);
and AND3 (N24258, N24257, N7583, N14479);
buf BUF1 (N24259, N24249);
nor NOR4 (N24260, N24256, N22108, N23693, N612);
not NOT1 (N24261, N24254);
or OR3 (N24262, N24260, N20177, N5137);
nand NAND2 (N24263, N24259, N4023);
not NOT1 (N24264, N24244);
and AND4 (N24265, N24248, N22730, N126, N19389);
not NOT1 (N24266, N24261);
and AND3 (N24267, N24255, N9489, N21980);
not NOT1 (N24268, N24264);
buf BUF1 (N24269, N24252);
xor XOR2 (N24270, N24267, N21355);
or OR3 (N24271, N24263, N20102, N22655);
nor NOR3 (N24272, N24266, N24092, N2187);
buf BUF1 (N24273, N24258);
nor NOR2 (N24274, N24270, N19159);
nand NAND2 (N24275, N24265, N17907);
nand NAND4 (N24276, N24268, N1168, N10006, N16743);
nand NAND2 (N24277, N24274, N5329);
not NOT1 (N24278, N24220);
not NOT1 (N24279, N24275);
xor XOR2 (N24280, N24277, N18825);
nand NAND3 (N24281, N24238, N20259, N3378);
and AND3 (N24282, N24262, N9225, N7334);
xor XOR2 (N24283, N24279, N11931);
buf BUF1 (N24284, N24271);
or OR4 (N24285, N24283, N4508, N10433, N4068);
xor XOR2 (N24286, N24276, N10880);
xor XOR2 (N24287, N24280, N18586);
xor XOR2 (N24288, N24286, N23855);
nand NAND3 (N24289, N24282, N5542, N11395);
nand NAND3 (N24290, N24278, N9896, N20235);
or OR4 (N24291, N24284, N2881, N20337, N3316);
nor NOR3 (N24292, N24281, N15842, N2843);
nand NAND2 (N24293, N24291, N11824);
and AND3 (N24294, N24287, N9204, N2304);
and AND4 (N24295, N24290, N17738, N16096, N5477);
not NOT1 (N24296, N24294);
and AND3 (N24297, N24293, N8851, N22563);
and AND4 (N24298, N24297, N4210, N16998, N19869);
and AND3 (N24299, N24269, N10811, N21635);
nor NOR4 (N24300, N24288, N11649, N22369, N16637);
and AND4 (N24301, N24289, N21624, N5238, N20067);
buf BUF1 (N24302, N24292);
nor NOR4 (N24303, N24272, N6643, N10477, N20608);
and AND3 (N24304, N24298, N6953, N20872);
not NOT1 (N24305, N24302);
nand NAND3 (N24306, N24303, N23886, N5195);
nand NAND4 (N24307, N24299, N7963, N17706, N23593);
nand NAND2 (N24308, N24306, N15989);
or OR2 (N24309, N24295, N7091);
and AND3 (N24310, N24307, N19743, N15260);
nor NOR4 (N24311, N24309, N7872, N15361, N19077);
or OR4 (N24312, N24311, N11221, N83, N8274);
not NOT1 (N24313, N24312);
not NOT1 (N24314, N24304);
nor NOR3 (N24315, N24308, N21791, N6604);
and AND4 (N24316, N24285, N3995, N14613, N8485);
nand NAND3 (N24317, N24296, N380, N9987);
xor XOR2 (N24318, N24313, N23485);
not NOT1 (N24319, N24273);
nand NAND3 (N24320, N24301, N2766, N11635);
xor XOR2 (N24321, N24300, N5568);
nor NOR4 (N24322, N24305, N21117, N12041, N19316);
or OR2 (N24323, N24321, N15112);
nand NAND4 (N24324, N24310, N9790, N2199, N14103);
and AND4 (N24325, N24314, N2514, N21613, N5537);
buf BUF1 (N24326, N24318);
or OR2 (N24327, N24317, N17214);
nand NAND4 (N24328, N24315, N22513, N16704, N10346);
nand NAND2 (N24329, N24323, N305);
or OR3 (N24330, N24326, N6796, N6669);
and AND2 (N24331, N24325, N21823);
not NOT1 (N24332, N24327);
buf BUF1 (N24333, N24329);
not NOT1 (N24334, N24332);
nor NOR4 (N24335, N24334, N23521, N8618, N21784);
and AND4 (N24336, N24333, N4366, N9712, N14115);
xor XOR2 (N24337, N24320, N21767);
buf BUF1 (N24338, N24336);
nor NOR4 (N24339, N24338, N23356, N12724, N19821);
or OR4 (N24340, N24316, N14119, N5714, N21607);
and AND4 (N24341, N24335, N15481, N682, N8569);
nor NOR4 (N24342, N24341, N13414, N4915, N8597);
nand NAND2 (N24343, N24339, N6620);
xor XOR2 (N24344, N24340, N7164);
or OR3 (N24345, N24322, N16612, N12211);
and AND4 (N24346, N24342, N69, N20306, N14445);
xor XOR2 (N24347, N24319, N15202);
not NOT1 (N24348, N24346);
and AND4 (N24349, N24345, N9904, N9542, N7558);
not NOT1 (N24350, N24349);
xor XOR2 (N24351, N24350, N24018);
not NOT1 (N24352, N24347);
nor NOR4 (N24353, N24352, N19807, N17333, N17016);
nand NAND2 (N24354, N24330, N2627);
and AND4 (N24355, N24348, N23492, N20598, N16614);
and AND4 (N24356, N24337, N21191, N23085, N10652);
xor XOR2 (N24357, N24354, N16722);
buf BUF1 (N24358, N24357);
not NOT1 (N24359, N24355);
nand NAND2 (N24360, N24344, N17109);
xor XOR2 (N24361, N24351, N12748);
nor NOR4 (N24362, N24360, N11752, N23533, N13127);
not NOT1 (N24363, N24358);
xor XOR2 (N24364, N24324, N18076);
xor XOR2 (N24365, N24364, N10011);
and AND4 (N24366, N24328, N22726, N2405, N15101);
nor NOR3 (N24367, N24343, N180, N10813);
buf BUF1 (N24368, N24331);
nor NOR3 (N24369, N24356, N11426, N10036);
not NOT1 (N24370, N24362);
or OR3 (N24371, N24367, N9362, N15312);
or OR3 (N24372, N24366, N8262, N6425);
nor NOR3 (N24373, N24369, N5523, N6355);
xor XOR2 (N24374, N24353, N17742);
nor NOR4 (N24375, N24374, N23658, N1275, N16803);
or OR3 (N24376, N24368, N13990, N11827);
xor XOR2 (N24377, N24361, N1394);
nand NAND3 (N24378, N24365, N22028, N20654);
xor XOR2 (N24379, N24370, N5963);
xor XOR2 (N24380, N24363, N16986);
not NOT1 (N24381, N24371);
buf BUF1 (N24382, N24381);
xor XOR2 (N24383, N24382, N4065);
or OR4 (N24384, N24376, N1423, N23851, N5048);
or OR2 (N24385, N24380, N23228);
nor NOR4 (N24386, N24359, N17762, N2383, N14467);
and AND4 (N24387, N24386, N12737, N1906, N19972);
xor XOR2 (N24388, N24372, N4781);
buf BUF1 (N24389, N24387);
or OR3 (N24390, N24379, N18418, N9523);
buf BUF1 (N24391, N24375);
not NOT1 (N24392, N24384);
nand NAND4 (N24393, N24391, N20185, N3491, N114);
and AND3 (N24394, N24378, N17658, N12765);
xor XOR2 (N24395, N24383, N5346);
nand NAND3 (N24396, N24395, N17441, N12876);
not NOT1 (N24397, N24393);
buf BUF1 (N24398, N24385);
not NOT1 (N24399, N24377);
xor XOR2 (N24400, N24396, N23110);
xor XOR2 (N24401, N24394, N1177);
nand NAND3 (N24402, N24398, N16482, N19898);
not NOT1 (N24403, N24373);
xor XOR2 (N24404, N24401, N5011);
nor NOR2 (N24405, N24399, N6330);
and AND3 (N24406, N24389, N10633, N21838);
xor XOR2 (N24407, N24397, N15534);
and AND3 (N24408, N24406, N890, N2485);
nand NAND3 (N24409, N24408, N10115, N15751);
and AND3 (N24410, N24402, N11118, N21906);
nor NOR4 (N24411, N24404, N22266, N12382, N14712);
nand NAND2 (N24412, N24390, N22694);
nor NOR3 (N24413, N24400, N10927, N7773);
nor NOR3 (N24414, N24392, N5164, N325);
nor NOR2 (N24415, N24409, N13539);
and AND2 (N24416, N24413, N18513);
buf BUF1 (N24417, N24407);
buf BUF1 (N24418, N24412);
xor XOR2 (N24419, N24417, N4389);
nor NOR3 (N24420, N24403, N2925, N5202);
nand NAND2 (N24421, N24418, N13079);
nand NAND4 (N24422, N24410, N2189, N573, N4470);
not NOT1 (N24423, N24414);
xor XOR2 (N24424, N24423, N1005);
xor XOR2 (N24425, N24421, N2193);
and AND2 (N24426, N24405, N18321);
nand NAND3 (N24427, N24420, N1085, N7588);
nand NAND2 (N24428, N24415, N18725);
nand NAND3 (N24429, N24428, N16349, N8847);
or OR2 (N24430, N24425, N12337);
buf BUF1 (N24431, N24427);
buf BUF1 (N24432, N24429);
buf BUF1 (N24433, N24426);
xor XOR2 (N24434, N24430, N24059);
buf BUF1 (N24435, N24433);
not NOT1 (N24436, N24388);
and AND2 (N24437, N24424, N19981);
not NOT1 (N24438, N24436);
nor NOR2 (N24439, N24416, N668);
buf BUF1 (N24440, N24422);
nand NAND4 (N24441, N24437, N19614, N5162, N17720);
or OR4 (N24442, N24419, N6975, N15376, N11762);
and AND3 (N24443, N24439, N9209, N1043);
nor NOR3 (N24444, N24432, N23288, N16177);
or OR2 (N24445, N24434, N3228);
buf BUF1 (N24446, N24435);
buf BUF1 (N24447, N24438);
buf BUF1 (N24448, N24446);
nand NAND3 (N24449, N24448, N9717, N19220);
and AND4 (N24450, N24431, N9727, N14612, N21987);
buf BUF1 (N24451, N24450);
not NOT1 (N24452, N24451);
buf BUF1 (N24453, N24449);
nand NAND2 (N24454, N24440, N6376);
or OR4 (N24455, N24447, N649, N14018, N7377);
nor NOR4 (N24456, N24441, N21769, N4678, N4608);
buf BUF1 (N24457, N24443);
buf BUF1 (N24458, N24456);
nand NAND4 (N24459, N24454, N14508, N21485, N5978);
buf BUF1 (N24460, N24458);
and AND2 (N24461, N24444, N12773);
buf BUF1 (N24462, N24461);
nor NOR3 (N24463, N24457, N5413, N11519);
nor NOR3 (N24464, N24462, N372, N20655);
not NOT1 (N24465, N24452);
and AND2 (N24466, N24453, N8903);
xor XOR2 (N24467, N24466, N11099);
xor XOR2 (N24468, N24445, N12339);
not NOT1 (N24469, N24459);
buf BUF1 (N24470, N24455);
nor NOR4 (N24471, N24467, N23790, N12813, N24282);
and AND2 (N24472, N24468, N7249);
not NOT1 (N24473, N24442);
not NOT1 (N24474, N24464);
and AND3 (N24475, N24474, N10789, N6178);
nand NAND3 (N24476, N24465, N13811, N10473);
not NOT1 (N24477, N24475);
or OR4 (N24478, N24471, N19303, N11972, N23477);
or OR3 (N24479, N24476, N7387, N8583);
xor XOR2 (N24480, N24463, N10883);
xor XOR2 (N24481, N24479, N12862);
and AND4 (N24482, N24478, N20198, N3954, N1887);
nor NOR4 (N24483, N24469, N11896, N16859, N12983);
not NOT1 (N24484, N24483);
xor XOR2 (N24485, N24411, N1738);
xor XOR2 (N24486, N24485, N4489);
or OR2 (N24487, N24477, N5729);
nand NAND3 (N24488, N24470, N2530, N428);
nor NOR3 (N24489, N24484, N4806, N14923);
or OR3 (N24490, N24472, N17207, N9085);
nor NOR3 (N24491, N24489, N20396, N21216);
not NOT1 (N24492, N24473);
not NOT1 (N24493, N24492);
not NOT1 (N24494, N24460);
and AND2 (N24495, N24487, N10918);
xor XOR2 (N24496, N24490, N22601);
not NOT1 (N24497, N24486);
nand NAND4 (N24498, N24491, N18022, N3216, N20803);
buf BUF1 (N24499, N24493);
nand NAND4 (N24500, N24480, N17249, N4599, N22288);
and AND4 (N24501, N24482, N5785, N20120, N21754);
or OR4 (N24502, N24500, N21947, N17753, N20274);
buf BUF1 (N24503, N24496);
nor NOR4 (N24504, N24497, N18523, N22248, N23344);
nor NOR3 (N24505, N24498, N2429, N447);
buf BUF1 (N24506, N24495);
nor NOR3 (N24507, N24494, N7810, N8457);
buf BUF1 (N24508, N24488);
buf BUF1 (N24509, N24499);
and AND2 (N24510, N24504, N17981);
nor NOR2 (N24511, N24501, N3922);
buf BUF1 (N24512, N24502);
xor XOR2 (N24513, N24503, N4710);
and AND2 (N24514, N24507, N9692);
nand NAND3 (N24515, N24511, N1685, N4107);
xor XOR2 (N24516, N24508, N9174);
nand NAND4 (N24517, N24506, N11730, N7008, N5294);
xor XOR2 (N24518, N24510, N3843);
not NOT1 (N24519, N24517);
and AND2 (N24520, N24512, N8723);
xor XOR2 (N24521, N24515, N8299);
and AND3 (N24522, N24519, N6746, N19535);
nand NAND3 (N24523, N24505, N4512, N3191);
not NOT1 (N24524, N24516);
xor XOR2 (N24525, N24513, N20150);
and AND3 (N24526, N24521, N11916, N24434);
or OR2 (N24527, N24523, N4886);
nor NOR3 (N24528, N24518, N14441, N7448);
or OR4 (N24529, N24528, N6197, N16390, N2130);
not NOT1 (N24530, N24481);
and AND2 (N24531, N24527, N21044);
not NOT1 (N24532, N24526);
and AND2 (N24533, N24514, N8671);
or OR2 (N24534, N24520, N8993);
nor NOR3 (N24535, N24532, N22752, N22379);
and AND3 (N24536, N24524, N13368, N20990);
and AND2 (N24537, N24533, N5273);
xor XOR2 (N24538, N24509, N12401);
not NOT1 (N24539, N24522);
or OR4 (N24540, N24529, N18565, N11194, N17100);
nand NAND3 (N24541, N24531, N11249, N4275);
or OR4 (N24542, N24525, N4625, N15987, N9672);
or OR4 (N24543, N24535, N8789, N19608, N5626);
xor XOR2 (N24544, N24537, N22012);
xor XOR2 (N24545, N24541, N23984);
and AND2 (N24546, N24536, N4821);
or OR4 (N24547, N24546, N9787, N24476, N12793);
not NOT1 (N24548, N24540);
or OR3 (N24549, N24539, N22292, N23749);
not NOT1 (N24550, N24547);
nor NOR4 (N24551, N24542, N5889, N22671, N8790);
not NOT1 (N24552, N24544);
and AND3 (N24553, N24538, N3914, N8556);
not NOT1 (N24554, N24550);
nor NOR4 (N24555, N24548, N21850, N15222, N15320);
buf BUF1 (N24556, N24543);
buf BUF1 (N24557, N24534);
or OR3 (N24558, N24556, N16150, N3676);
nor NOR2 (N24559, N24530, N1502);
or OR4 (N24560, N24553, N18083, N21706, N3652);
or OR3 (N24561, N24554, N18171, N13528);
or OR3 (N24562, N24557, N13965, N16797);
and AND3 (N24563, N24552, N14863, N9575);
buf BUF1 (N24564, N24562);
nor NOR3 (N24565, N24563, N17777, N5809);
and AND3 (N24566, N24551, N17291, N22918);
not NOT1 (N24567, N24565);
and AND3 (N24568, N24566, N5678, N47);
not NOT1 (N24569, N24555);
buf BUF1 (N24570, N24560);
or OR3 (N24571, N24569, N11684, N22411);
nor NOR4 (N24572, N24558, N1599, N1857, N12936);
not NOT1 (N24573, N24572);
nor NOR2 (N24574, N24561, N3123);
buf BUF1 (N24575, N24545);
and AND4 (N24576, N24571, N16757, N14279, N1592);
nor NOR4 (N24577, N24570, N7933, N2685, N4760);
nand NAND4 (N24578, N24577, N5891, N1344, N1488);
not NOT1 (N24579, N24578);
xor XOR2 (N24580, N24579, N15906);
nand NAND4 (N24581, N24549, N22217, N5738, N10417);
not NOT1 (N24582, N24574);
not NOT1 (N24583, N24575);
nor NOR4 (N24584, N24559, N24252, N9185, N9370);
not NOT1 (N24585, N24568);
and AND3 (N24586, N24580, N18074, N15336);
not NOT1 (N24587, N24581);
not NOT1 (N24588, N24585);
buf BUF1 (N24589, N24582);
and AND4 (N24590, N24588, N12095, N15027, N19148);
and AND4 (N24591, N24583, N4600, N5437, N8213);
buf BUF1 (N24592, N24590);
xor XOR2 (N24593, N24592, N24120);
nor NOR4 (N24594, N24586, N12245, N6378, N16357);
xor XOR2 (N24595, N24593, N20929);
not NOT1 (N24596, N24587);
buf BUF1 (N24597, N24573);
and AND3 (N24598, N24564, N5839, N14958);
nand NAND2 (N24599, N24567, N3392);
nor NOR4 (N24600, N24591, N10208, N3622, N11152);
buf BUF1 (N24601, N24598);
xor XOR2 (N24602, N24601, N13958);
and AND2 (N24603, N24597, N3076);
buf BUF1 (N24604, N24589);
nand NAND4 (N24605, N24576, N2567, N18127, N22371);
buf BUF1 (N24606, N24604);
or OR3 (N24607, N24603, N16229, N19806);
not NOT1 (N24608, N24607);
nand NAND4 (N24609, N24606, N22006, N619, N10285);
buf BUF1 (N24610, N24605);
and AND3 (N24611, N24594, N5026, N383);
not NOT1 (N24612, N24599);
nor NOR4 (N24613, N24608, N16608, N2650, N14365);
nand NAND3 (N24614, N24613, N6926, N14552);
xor XOR2 (N24615, N24600, N8776);
xor XOR2 (N24616, N24596, N18679);
nand NAND3 (N24617, N24584, N11899, N15251);
xor XOR2 (N24618, N24616, N22287);
or OR3 (N24619, N24618, N1850, N9047);
buf BUF1 (N24620, N24602);
nor NOR4 (N24621, N24615, N15404, N13324, N20230);
or OR4 (N24622, N24614, N12282, N10723, N17142);
nand NAND3 (N24623, N24621, N6436, N18691);
nand NAND4 (N24624, N24617, N23789, N8506, N5580);
or OR2 (N24625, N24612, N22758);
or OR4 (N24626, N24623, N18011, N6967, N4650);
and AND4 (N24627, N24595, N19634, N18857, N297);
buf BUF1 (N24628, N24611);
buf BUF1 (N24629, N24626);
nor NOR2 (N24630, N24624, N3786);
xor XOR2 (N24631, N24622, N8651);
or OR4 (N24632, N24631, N6842, N4079, N12947);
xor XOR2 (N24633, N24625, N3928);
or OR2 (N24634, N24610, N8550);
not NOT1 (N24635, N24630);
not NOT1 (N24636, N24629);
buf BUF1 (N24637, N24636);
nor NOR3 (N24638, N24627, N24111, N5576);
or OR2 (N24639, N24637, N16444);
buf BUF1 (N24640, N24628);
nand NAND4 (N24641, N24620, N19860, N517, N23770);
and AND2 (N24642, N24634, N6190);
nor NOR3 (N24643, N24639, N19594, N5459);
nand NAND3 (N24644, N24643, N19667, N13563);
or OR2 (N24645, N24635, N16988);
and AND4 (N24646, N24642, N15144, N11407, N4226);
xor XOR2 (N24647, N24609, N22055);
xor XOR2 (N24648, N24640, N21484);
not NOT1 (N24649, N24638);
xor XOR2 (N24650, N24645, N8527);
nor NOR2 (N24651, N24619, N8781);
nand NAND3 (N24652, N24632, N14946, N21778);
and AND3 (N24653, N24652, N12108, N6648);
nor NOR2 (N24654, N24646, N18541);
not NOT1 (N24655, N24647);
buf BUF1 (N24656, N24648);
not NOT1 (N24657, N24644);
nand NAND3 (N24658, N24654, N24633, N7958);
buf BUF1 (N24659, N1935);
not NOT1 (N24660, N24656);
and AND4 (N24661, N24649, N10632, N6280, N16514);
xor XOR2 (N24662, N24653, N22049);
buf BUF1 (N24663, N24658);
buf BUF1 (N24664, N24660);
buf BUF1 (N24665, N24657);
xor XOR2 (N24666, N24650, N592);
buf BUF1 (N24667, N24666);
not NOT1 (N24668, N24662);
nand NAND2 (N24669, N24655, N3319);
and AND3 (N24670, N24651, N16164, N17167);
nand NAND2 (N24671, N24668, N801);
xor XOR2 (N24672, N24667, N5376);
or OR4 (N24673, N24672, N2475, N17229, N2636);
xor XOR2 (N24674, N24641, N23038);
not NOT1 (N24675, N24670);
and AND2 (N24676, N24673, N17923);
buf BUF1 (N24677, N24663);
xor XOR2 (N24678, N24675, N5445);
or OR3 (N24679, N24671, N16207, N20754);
xor XOR2 (N24680, N24676, N18529);
or OR2 (N24681, N24659, N11583);
nor NOR4 (N24682, N24661, N10894, N386, N7476);
and AND2 (N24683, N24681, N22628);
or OR2 (N24684, N24682, N15619);
buf BUF1 (N24685, N24683);
or OR3 (N24686, N24677, N11026, N10242);
or OR4 (N24687, N24684, N13922, N21533, N17720);
not NOT1 (N24688, N24669);
or OR2 (N24689, N24685, N5410);
and AND3 (N24690, N24664, N16370, N3201);
or OR4 (N24691, N24688, N1926, N2036, N17938);
nand NAND2 (N24692, N24680, N558);
nand NAND4 (N24693, N24687, N1320, N12287, N15153);
and AND3 (N24694, N24686, N24404, N21619);
nor NOR2 (N24695, N24674, N12059);
nand NAND2 (N24696, N24692, N19629);
nand NAND2 (N24697, N24690, N1442);
not NOT1 (N24698, N24693);
nor NOR3 (N24699, N24698, N1803, N4900);
not NOT1 (N24700, N24696);
nand NAND2 (N24701, N24679, N16379);
buf BUF1 (N24702, N24694);
buf BUF1 (N24703, N24689);
or OR4 (N24704, N24678, N15743, N5377, N17679);
buf BUF1 (N24705, N24701);
xor XOR2 (N24706, N24691, N13108);
not NOT1 (N24707, N24700);
nor NOR3 (N24708, N24702, N19433, N6954);
or OR4 (N24709, N24708, N2420, N12195, N16359);
nor NOR4 (N24710, N24704, N21413, N7033, N1459);
nand NAND3 (N24711, N24665, N12437, N9423);
and AND4 (N24712, N24703, N891, N3986, N18730);
or OR4 (N24713, N24699, N17475, N20357, N21371);
or OR3 (N24714, N24705, N1891, N6575);
buf BUF1 (N24715, N24697);
not NOT1 (N24716, N24706);
not NOT1 (N24717, N24714);
or OR4 (N24718, N24695, N15967, N17657, N21728);
nand NAND4 (N24719, N24711, N9253, N10849, N10386);
nor NOR4 (N24720, N24715, N16317, N1891, N21670);
buf BUF1 (N24721, N24720);
buf BUF1 (N24722, N24712);
buf BUF1 (N24723, N24717);
nand NAND4 (N24724, N24713, N5899, N14572, N21987);
or OR4 (N24725, N24707, N1238, N14617, N21384);
xor XOR2 (N24726, N24718, N19319);
buf BUF1 (N24727, N24725);
and AND3 (N24728, N24709, N23495, N5124);
nor NOR2 (N24729, N24727, N22353);
not NOT1 (N24730, N24723);
buf BUF1 (N24731, N24710);
nand NAND2 (N24732, N24731, N19526);
not NOT1 (N24733, N24728);
xor XOR2 (N24734, N24722, N8244);
or OR3 (N24735, N24716, N23164, N17568);
nor NOR4 (N24736, N24733, N19725, N135, N10805);
and AND2 (N24737, N24719, N23895);
nand NAND2 (N24738, N24732, N2156);
buf BUF1 (N24739, N24726);
nand NAND3 (N24740, N24729, N24657, N5189);
and AND3 (N24741, N24721, N22318, N22446);
and AND2 (N24742, N24736, N11167);
buf BUF1 (N24743, N24738);
not NOT1 (N24744, N24730);
buf BUF1 (N24745, N24735);
not NOT1 (N24746, N24743);
xor XOR2 (N24747, N24741, N8906);
nor NOR2 (N24748, N24747, N803);
nand NAND2 (N24749, N24742, N10244);
not NOT1 (N24750, N24739);
nand NAND4 (N24751, N24749, N18743, N23935, N11549);
and AND3 (N24752, N24748, N14395, N13148);
not NOT1 (N24753, N24734);
not NOT1 (N24754, N24740);
or OR4 (N24755, N24737, N11229, N22388, N17858);
nor NOR4 (N24756, N24751, N2932, N22490, N23612);
not NOT1 (N24757, N24754);
xor XOR2 (N24758, N24756, N2975);
not NOT1 (N24759, N24757);
xor XOR2 (N24760, N24758, N6758);
and AND3 (N24761, N24745, N7855, N24403);
not NOT1 (N24762, N24760);
xor XOR2 (N24763, N24762, N9818);
nor NOR2 (N24764, N24759, N23845);
not NOT1 (N24765, N24752);
or OR4 (N24766, N24724, N18663, N962, N8176);
and AND3 (N24767, N24761, N16157, N913);
buf BUF1 (N24768, N24750);
nor NOR3 (N24769, N24753, N16960, N5994);
nand NAND2 (N24770, N24764, N21596);
and AND4 (N24771, N24768, N17066, N19071, N7631);
not NOT1 (N24772, N24755);
nand NAND3 (N24773, N24763, N11338, N2922);
nand NAND2 (N24774, N24769, N3859);
buf BUF1 (N24775, N24774);
or OR3 (N24776, N24765, N10258, N18394);
buf BUF1 (N24777, N24773);
buf BUF1 (N24778, N24770);
not NOT1 (N24779, N24767);
nand NAND4 (N24780, N24771, N468, N20495, N6771);
and AND3 (N24781, N24746, N5667, N15126);
nor NOR2 (N24782, N24780, N1205);
and AND3 (N24783, N24778, N14440, N11871);
nor NOR3 (N24784, N24776, N21164, N11069);
nor NOR4 (N24785, N24772, N8642, N23881, N21776);
or OR2 (N24786, N24766, N9536);
nor NOR4 (N24787, N24783, N938, N15028, N2594);
or OR3 (N24788, N24785, N24335, N24709);
nor NOR2 (N24789, N24781, N3721);
not NOT1 (N24790, N24784);
or OR4 (N24791, N24775, N17630, N14533, N20927);
nor NOR2 (N24792, N24789, N5046);
or OR4 (N24793, N24779, N22317, N9518, N20966);
xor XOR2 (N24794, N24787, N19030);
nand NAND3 (N24795, N24782, N1564, N11417);
and AND2 (N24796, N24777, N20161);
nand NAND3 (N24797, N24790, N12311, N9077);
nor NOR3 (N24798, N24794, N4658, N17861);
xor XOR2 (N24799, N24793, N15136);
and AND4 (N24800, N24744, N2489, N6803, N13691);
or OR3 (N24801, N24786, N2070, N9093);
and AND2 (N24802, N24800, N7110);
and AND4 (N24803, N24801, N13544, N6004, N4352);
buf BUF1 (N24804, N24799);
and AND2 (N24805, N24792, N23735);
nand NAND4 (N24806, N24796, N17921, N9455, N13388);
buf BUF1 (N24807, N24805);
nand NAND2 (N24808, N24804, N6807);
not NOT1 (N24809, N24808);
nand NAND2 (N24810, N24788, N4322);
nor NOR2 (N24811, N24797, N7270);
xor XOR2 (N24812, N24806, N12154);
buf BUF1 (N24813, N24791);
not NOT1 (N24814, N24811);
buf BUF1 (N24815, N24814);
buf BUF1 (N24816, N24812);
or OR3 (N24817, N24809, N22349, N5267);
nor NOR3 (N24818, N24803, N24706, N18204);
or OR3 (N24819, N24815, N11914, N13577);
xor XOR2 (N24820, N24813, N23626);
and AND4 (N24821, N24810, N24357, N11106, N4278);
xor XOR2 (N24822, N24798, N14467);
nor NOR4 (N24823, N24816, N15906, N1748, N4526);
not NOT1 (N24824, N24807);
xor XOR2 (N24825, N24795, N3236);
nand NAND4 (N24826, N24823, N17783, N14567, N18171);
and AND4 (N24827, N24819, N10511, N2848, N22563);
nand NAND4 (N24828, N24824, N1963, N5755, N8811);
xor XOR2 (N24829, N24828, N3890);
xor XOR2 (N24830, N24817, N19892);
xor XOR2 (N24831, N24830, N14323);
not NOT1 (N24832, N24822);
not NOT1 (N24833, N24829);
and AND3 (N24834, N24827, N12324, N15464);
nand NAND3 (N24835, N24820, N14037, N6476);
and AND4 (N24836, N24831, N15648, N278, N2636);
xor XOR2 (N24837, N24834, N24739);
and AND2 (N24838, N24832, N23820);
and AND3 (N24839, N24826, N21594, N9623);
not NOT1 (N24840, N24837);
xor XOR2 (N24841, N24825, N23891);
buf BUF1 (N24842, N24835);
nor NOR4 (N24843, N24821, N5588, N37, N24323);
xor XOR2 (N24844, N24842, N22187);
and AND3 (N24845, N24840, N16645, N17251);
buf BUF1 (N24846, N24845);
nor NOR3 (N24847, N24839, N13836, N21003);
nor NOR2 (N24848, N24844, N4496);
not NOT1 (N24849, N24848);
xor XOR2 (N24850, N24833, N5726);
buf BUF1 (N24851, N24846);
xor XOR2 (N24852, N24841, N21910);
or OR2 (N24853, N24850, N198);
xor XOR2 (N24854, N24852, N11456);
not NOT1 (N24855, N24849);
xor XOR2 (N24856, N24854, N3521);
xor XOR2 (N24857, N24851, N143);
buf BUF1 (N24858, N24838);
xor XOR2 (N24859, N24858, N14434);
buf BUF1 (N24860, N24856);
not NOT1 (N24861, N24855);
buf BUF1 (N24862, N24843);
nand NAND3 (N24863, N24861, N14178, N1377);
nor NOR3 (N24864, N24818, N17032, N19307);
nand NAND4 (N24865, N24859, N21744, N3782, N10756);
nor NOR4 (N24866, N24860, N2857, N1664, N1499);
nor NOR4 (N24867, N24853, N10750, N24348, N21868);
and AND4 (N24868, N24863, N20086, N1095, N21676);
buf BUF1 (N24869, N24865);
and AND3 (N24870, N24857, N2422, N5853);
xor XOR2 (N24871, N24870, N23028);
nand NAND4 (N24872, N24871, N19775, N3910, N1770);
or OR3 (N24873, N24847, N1464, N10164);
not NOT1 (N24874, N24862);
and AND3 (N24875, N24868, N18090, N11082);
buf BUF1 (N24876, N24874);
and AND3 (N24877, N24873, N18586, N23235);
xor XOR2 (N24878, N24867, N21410);
or OR4 (N24879, N24878, N3445, N24059, N7300);
not NOT1 (N24880, N24875);
not NOT1 (N24881, N24836);
or OR4 (N24882, N24877, N15953, N6707, N23927);
not NOT1 (N24883, N24866);
and AND3 (N24884, N24802, N14858, N24538);
not NOT1 (N24885, N24880);
or OR2 (N24886, N24885, N9246);
buf BUF1 (N24887, N24872);
buf BUF1 (N24888, N24869);
nand NAND3 (N24889, N24881, N128, N14663);
nand NAND3 (N24890, N24889, N3712, N7858);
buf BUF1 (N24891, N24890);
xor XOR2 (N24892, N24891, N2150);
and AND3 (N24893, N24884, N12712, N12826);
not NOT1 (N24894, N24864);
buf BUF1 (N24895, N24876);
buf BUF1 (N24896, N24879);
not NOT1 (N24897, N24886);
xor XOR2 (N24898, N24895, N16576);
buf BUF1 (N24899, N24894);
or OR2 (N24900, N24898, N1337);
buf BUF1 (N24901, N24893);
or OR3 (N24902, N24892, N5068, N21176);
buf BUF1 (N24903, N24900);
nand NAND2 (N24904, N24887, N6530);
buf BUF1 (N24905, N24902);
not NOT1 (N24906, N24903);
buf BUF1 (N24907, N24904);
not NOT1 (N24908, N24883);
nand NAND4 (N24909, N24882, N9485, N2859, N12392);
and AND2 (N24910, N24909, N15105);
or OR4 (N24911, N24888, N15965, N21042, N4748);
xor XOR2 (N24912, N24907, N24299);
not NOT1 (N24913, N24912);
nand NAND3 (N24914, N24899, N21150, N13651);
or OR2 (N24915, N24897, N8399);
buf BUF1 (N24916, N24915);
nand NAND3 (N24917, N24896, N13788, N10497);
xor XOR2 (N24918, N24917, N10029);
xor XOR2 (N24919, N24911, N7943);
buf BUF1 (N24920, N24906);
not NOT1 (N24921, N24920);
and AND3 (N24922, N24914, N4768, N10725);
buf BUF1 (N24923, N24913);
nand NAND4 (N24924, N24923, N17051, N6752, N3708);
nor NOR2 (N24925, N24908, N8691);
nor NOR3 (N24926, N24922, N8171, N13730);
xor XOR2 (N24927, N24926, N4698);
nand NAND4 (N24928, N24916, N14491, N14071, N21443);
or OR2 (N24929, N24901, N12588);
buf BUF1 (N24930, N24905);
or OR2 (N24931, N24927, N5072);
and AND3 (N24932, N24921, N15718, N22782);
buf BUF1 (N24933, N24925);
nor NOR2 (N24934, N24932, N4696);
not NOT1 (N24935, N24928);
nor NOR2 (N24936, N24918, N7771);
or OR3 (N24937, N24919, N17565, N4957);
and AND3 (N24938, N24931, N22252, N5471);
nand NAND3 (N24939, N24938, N1572, N1310);
and AND3 (N24940, N24924, N17985, N13236);
and AND3 (N24941, N24934, N20878, N2306);
nand NAND4 (N24942, N24937, N1873, N16126, N10013);
or OR2 (N24943, N24940, N23073);
and AND3 (N24944, N24933, N6293, N15327);
not NOT1 (N24945, N24941);
buf BUF1 (N24946, N24936);
nor NOR2 (N24947, N24929, N9520);
xor XOR2 (N24948, N24943, N13884);
nor NOR2 (N24949, N24942, N15032);
not NOT1 (N24950, N24930);
or OR3 (N24951, N24939, N12017, N3869);
nand NAND3 (N24952, N24946, N12934, N3285);
and AND4 (N24953, N24944, N1446, N17179, N19028);
or OR3 (N24954, N24948, N3625, N7616);
nor NOR2 (N24955, N24951, N12379);
not NOT1 (N24956, N24953);
not NOT1 (N24957, N24954);
buf BUF1 (N24958, N24910);
nand NAND4 (N24959, N24950, N9664, N10555, N18366);
nand NAND2 (N24960, N24947, N18267);
and AND2 (N24961, N24955, N15045);
buf BUF1 (N24962, N24958);
nand NAND2 (N24963, N24962, N14420);
not NOT1 (N24964, N24961);
buf BUF1 (N24965, N24956);
not NOT1 (N24966, N24952);
or OR2 (N24967, N24949, N9863);
nor NOR4 (N24968, N24960, N15989, N22920, N3292);
or OR2 (N24969, N24945, N22960);
not NOT1 (N24970, N24965);
and AND4 (N24971, N24966, N1979, N5611, N16376);
not NOT1 (N24972, N24970);
and AND3 (N24973, N24971, N15731, N11487);
nor NOR2 (N24974, N24968, N22223);
nand NAND3 (N24975, N24972, N20769, N21675);
or OR3 (N24976, N24935, N20214, N12959);
nor NOR2 (N24977, N24974, N20541);
and AND3 (N24978, N24975, N18346, N22509);
not NOT1 (N24979, N24967);
and AND4 (N24980, N24957, N13705, N17793, N21788);
not NOT1 (N24981, N24979);
nand NAND4 (N24982, N24964, N22703, N6216, N9718);
and AND3 (N24983, N24969, N22378, N15311);
nor NOR3 (N24984, N24963, N19983, N6469);
buf BUF1 (N24985, N24980);
xor XOR2 (N24986, N24983, N21127);
not NOT1 (N24987, N24981);
and AND4 (N24988, N24987, N350, N8003, N5114);
nand NAND3 (N24989, N24977, N20946, N2460);
buf BUF1 (N24990, N24985);
nand NAND4 (N24991, N24976, N8998, N11556, N858);
not NOT1 (N24992, N24988);
xor XOR2 (N24993, N24986, N16868);
buf BUF1 (N24994, N24993);
not NOT1 (N24995, N24992);
buf BUF1 (N24996, N24990);
nand NAND4 (N24997, N24973, N21998, N20001, N313);
not NOT1 (N24998, N24991);
not NOT1 (N24999, N24995);
nand NAND2 (N25000, N24998, N15236);
buf BUF1 (N25001, N24984);
nand NAND3 (N25002, N24999, N16370, N18022);
or OR2 (N25003, N24959, N17410);
or OR3 (N25004, N24982, N24398, N18557);
nor NOR4 (N25005, N24978, N21869, N21594, N22933);
xor XOR2 (N25006, N25001, N7411);
or OR2 (N25007, N25004, N18402);
xor XOR2 (N25008, N25006, N11655);
nand NAND3 (N25009, N25002, N3846, N6036);
and AND2 (N25010, N24994, N16460);
not NOT1 (N25011, N24997);
nand NAND3 (N25012, N24996, N23328, N22729);
or OR4 (N25013, N25009, N5585, N18124, N5276);
xor XOR2 (N25014, N25010, N4497);
xor XOR2 (N25015, N25014, N4017);
and AND3 (N25016, N25000, N10602, N20639);
nor NOR4 (N25017, N25012, N6338, N23506, N23716);
and AND2 (N25018, N25015, N4683);
nor NOR4 (N25019, N25013, N12772, N24562, N21843);
nor NOR4 (N25020, N25019, N7580, N6819, N20377);
not NOT1 (N25021, N25005);
not NOT1 (N25022, N24989);
and AND2 (N25023, N25008, N11186);
or OR3 (N25024, N25018, N14461, N16199);
not NOT1 (N25025, N25011);
nor NOR4 (N25026, N25007, N3847, N6063, N11313);
nor NOR4 (N25027, N25025, N70, N13948, N24048);
xor XOR2 (N25028, N25017, N3905);
nand NAND2 (N25029, N25003, N2906);
nor NOR4 (N25030, N25022, N3237, N5750, N18979);
or OR3 (N25031, N25023, N9575, N16898);
xor XOR2 (N25032, N25026, N3727);
or OR4 (N25033, N25024, N14737, N17092, N22389);
nand NAND4 (N25034, N25032, N22824, N10419, N11036);
nand NAND4 (N25035, N25033, N11059, N7136, N20083);
or OR3 (N25036, N25028, N524, N5213);
not NOT1 (N25037, N25036);
nand NAND4 (N25038, N25020, N18296, N8258, N5950);
nand NAND4 (N25039, N25016, N7228, N9866, N19421);
nand NAND3 (N25040, N25037, N10202, N19732);
and AND4 (N25041, N25034, N4194, N19640, N13993);
nor NOR2 (N25042, N25035, N23350);
buf BUF1 (N25043, N25038);
or OR4 (N25044, N25040, N2859, N18037, N2976);
xor XOR2 (N25045, N25043, N11161);
or OR3 (N25046, N25029, N1651, N9841);
and AND3 (N25047, N25042, N18613, N16882);
and AND2 (N25048, N25039, N1285);
and AND4 (N25049, N25030, N1930, N12843, N17719);
xor XOR2 (N25050, N25046, N23032);
nand NAND3 (N25051, N25048, N20575, N9107);
or OR2 (N25052, N25047, N14795);
and AND2 (N25053, N25052, N24304);
nand NAND3 (N25054, N25044, N5454, N15906);
buf BUF1 (N25055, N25049);
or OR2 (N25056, N25045, N7226);
not NOT1 (N25057, N25051);
and AND4 (N25058, N25050, N10949, N20515, N21473);
and AND3 (N25059, N25058, N21998, N718);
and AND3 (N25060, N25031, N16031, N12196);
xor XOR2 (N25061, N25056, N1031);
or OR2 (N25062, N25060, N18655);
xor XOR2 (N25063, N25054, N17056);
not NOT1 (N25064, N25062);
buf BUF1 (N25065, N25021);
nand NAND4 (N25066, N25059, N12055, N10659, N193);
or OR2 (N25067, N25055, N12312);
xor XOR2 (N25068, N25041, N5873);
xor XOR2 (N25069, N25063, N22064);
not NOT1 (N25070, N25027);
or OR4 (N25071, N25070, N22587, N5443, N7965);
buf BUF1 (N25072, N25061);
not NOT1 (N25073, N25057);
or OR2 (N25074, N25067, N21422);
nand NAND3 (N25075, N25064, N22533, N2502);
and AND4 (N25076, N25053, N7411, N7435, N20030);
nor NOR4 (N25077, N25076, N13908, N13723, N10205);
and AND4 (N25078, N25077, N10339, N3299, N14354);
nand NAND4 (N25079, N25068, N7266, N2618, N13846);
nor NOR3 (N25080, N25079, N10907, N13214);
not NOT1 (N25081, N25065);
not NOT1 (N25082, N25074);
or OR2 (N25083, N25082, N24456);
buf BUF1 (N25084, N25075);
buf BUF1 (N25085, N25081);
not NOT1 (N25086, N25069);
or OR2 (N25087, N25080, N9279);
buf BUF1 (N25088, N25066);
nand NAND3 (N25089, N25083, N19918, N22444);
not NOT1 (N25090, N25086);
xor XOR2 (N25091, N25088, N10039);
or OR2 (N25092, N25089, N4413);
or OR2 (N25093, N25073, N17625);
xor XOR2 (N25094, N25090, N21677);
and AND2 (N25095, N25087, N20637);
buf BUF1 (N25096, N25091);
nand NAND4 (N25097, N25093, N1033, N8471, N23082);
or OR2 (N25098, N25072, N6140);
nand NAND3 (N25099, N25084, N7156, N3745);
xor XOR2 (N25100, N25094, N5862);
not NOT1 (N25101, N25099);
or OR4 (N25102, N25100, N61, N328, N15616);
or OR4 (N25103, N25098, N19673, N8087, N1082);
or OR3 (N25104, N25095, N7444, N24576);
nand NAND3 (N25105, N25104, N5595, N10995);
not NOT1 (N25106, N25078);
not NOT1 (N25107, N25102);
not NOT1 (N25108, N25085);
or OR4 (N25109, N25071, N14845, N5873, N215);
nor NOR3 (N25110, N25108, N14381, N13888);
and AND2 (N25111, N25110, N9139);
nor NOR4 (N25112, N25106, N17286, N15674, N8359);
buf BUF1 (N25113, N25097);
and AND4 (N25114, N25101, N9836, N17426, N19850);
and AND2 (N25115, N25109, N1078);
xor XOR2 (N25116, N25112, N17317);
nand NAND4 (N25117, N25113, N2100, N43, N23330);
or OR2 (N25118, N25114, N870);
xor XOR2 (N25119, N25115, N464);
nand NAND4 (N25120, N25117, N1807, N19377, N19072);
xor XOR2 (N25121, N25116, N11952);
nand NAND2 (N25122, N25119, N18271);
or OR4 (N25123, N25118, N17805, N612, N23694);
not NOT1 (N25124, N25092);
buf BUF1 (N25125, N25124);
nor NOR2 (N25126, N25123, N22870);
nor NOR2 (N25127, N25125, N13373);
xor XOR2 (N25128, N25096, N2023);
nor NOR3 (N25129, N25128, N22263, N12702);
xor XOR2 (N25130, N25122, N4162);
not NOT1 (N25131, N25120);
buf BUF1 (N25132, N25111);
xor XOR2 (N25133, N25107, N24631);
buf BUF1 (N25134, N25131);
nor NOR3 (N25135, N25126, N11291, N12307);
or OR3 (N25136, N25127, N6486, N7334);
nor NOR4 (N25137, N25130, N2917, N9548, N23666);
and AND4 (N25138, N25103, N7716, N12276, N13500);
xor XOR2 (N25139, N25138, N24120);
xor XOR2 (N25140, N25134, N5985);
or OR3 (N25141, N25136, N16414, N6814);
not NOT1 (N25142, N25132);
and AND2 (N25143, N25142, N12790);
buf BUF1 (N25144, N25105);
xor XOR2 (N25145, N25141, N17900);
nand NAND4 (N25146, N25129, N17072, N5078, N25059);
and AND3 (N25147, N25133, N3769, N11502);
buf BUF1 (N25148, N25140);
and AND4 (N25149, N25135, N3714, N21521, N1117);
and AND2 (N25150, N25148, N24507);
or OR4 (N25151, N25146, N7281, N8019, N22032);
not NOT1 (N25152, N25139);
nor NOR3 (N25153, N25150, N19294, N15081);
and AND3 (N25154, N25143, N17970, N20436);
not NOT1 (N25155, N25152);
nand NAND3 (N25156, N25154, N20240, N7856);
nor NOR4 (N25157, N25147, N23282, N13698, N5311);
xor XOR2 (N25158, N25155, N11461);
and AND4 (N25159, N25151, N11873, N19121, N23055);
not NOT1 (N25160, N25145);
xor XOR2 (N25161, N25156, N14665);
nor NOR4 (N25162, N25144, N23499, N19800, N2114);
nand NAND2 (N25163, N25159, N24125);
xor XOR2 (N25164, N25121, N5120);
buf BUF1 (N25165, N25153);
not NOT1 (N25166, N25160);
or OR2 (N25167, N25157, N17772);
xor XOR2 (N25168, N25165, N14711);
or OR4 (N25169, N25137, N17711, N24038, N7585);
nand NAND3 (N25170, N25167, N15979, N13812);
xor XOR2 (N25171, N25162, N18064);
xor XOR2 (N25172, N25164, N19985);
or OR2 (N25173, N25161, N21648);
and AND2 (N25174, N25149, N24709);
not NOT1 (N25175, N25171);
and AND4 (N25176, N25168, N5074, N25150, N16118);
nor NOR2 (N25177, N25172, N6520);
nor NOR3 (N25178, N25174, N3016, N11947);
not NOT1 (N25179, N25176);
not NOT1 (N25180, N25177);
xor XOR2 (N25181, N25179, N19237);
buf BUF1 (N25182, N25170);
xor XOR2 (N25183, N25166, N11442);
or OR2 (N25184, N25182, N22312);
and AND4 (N25185, N25175, N629, N15642, N15532);
buf BUF1 (N25186, N25183);
not NOT1 (N25187, N25163);
nor NOR4 (N25188, N25180, N24748, N10015, N8292);
or OR3 (N25189, N25178, N14305, N2111);
nand NAND3 (N25190, N25188, N9431, N14883);
buf BUF1 (N25191, N25186);
and AND2 (N25192, N25189, N9128);
and AND4 (N25193, N25187, N23523, N2118, N19673);
nand NAND3 (N25194, N25191, N13283, N18975);
or OR3 (N25195, N25190, N8053, N17973);
not NOT1 (N25196, N25195);
not NOT1 (N25197, N25192);
buf BUF1 (N25198, N25158);
and AND2 (N25199, N25197, N7233);
not NOT1 (N25200, N25198);
and AND4 (N25201, N25196, N7039, N5477, N18421);
or OR2 (N25202, N25201, N12288);
nor NOR2 (N25203, N25194, N6578);
not NOT1 (N25204, N25193);
or OR2 (N25205, N25199, N9850);
nand NAND4 (N25206, N25205, N17762, N301, N820);
buf BUF1 (N25207, N25203);
or OR4 (N25208, N25202, N22369, N24365, N23625);
nand NAND4 (N25209, N25206, N15130, N10176, N21926);
or OR2 (N25210, N25207, N17194);
xor XOR2 (N25211, N25204, N21461);
and AND2 (N25212, N25210, N2321);
and AND3 (N25213, N25212, N7187, N8765);
or OR3 (N25214, N25211, N12223, N24804);
xor XOR2 (N25215, N25181, N6959);
nand NAND2 (N25216, N25215, N20260);
xor XOR2 (N25217, N25216, N19400);
xor XOR2 (N25218, N25213, N14356);
not NOT1 (N25219, N25209);
not NOT1 (N25220, N25218);
and AND2 (N25221, N25208, N16942);
buf BUF1 (N25222, N25219);
not NOT1 (N25223, N25185);
or OR4 (N25224, N25221, N15399, N16789, N13792);
nand NAND4 (N25225, N25184, N1475, N6697, N16400);
nand NAND3 (N25226, N25222, N4037, N488);
not NOT1 (N25227, N25223);
nand NAND3 (N25228, N25220, N11335, N5331);
nand NAND2 (N25229, N25228, N1606);
buf BUF1 (N25230, N25214);
xor XOR2 (N25231, N25225, N18863);
nand NAND2 (N25232, N25231, N657);
nor NOR3 (N25233, N25224, N15256, N23406);
not NOT1 (N25234, N25229);
nor NOR4 (N25235, N25230, N9468, N463, N22733);
xor XOR2 (N25236, N25173, N11849);
xor XOR2 (N25237, N25169, N5207);
buf BUF1 (N25238, N25234);
buf BUF1 (N25239, N25227);
nor NOR3 (N25240, N25235, N19302, N4689);
buf BUF1 (N25241, N25240);
or OR2 (N25242, N25239, N21449);
not NOT1 (N25243, N25242);
and AND3 (N25244, N25233, N8630, N23896);
xor XOR2 (N25245, N25244, N4238);
nand NAND4 (N25246, N25232, N1892, N14359, N8711);
buf BUF1 (N25247, N25246);
or OR2 (N25248, N25226, N24497);
or OR3 (N25249, N25248, N23532, N13203);
not NOT1 (N25250, N25238);
not NOT1 (N25251, N25245);
xor XOR2 (N25252, N25243, N15698);
and AND3 (N25253, N25252, N24343, N19216);
or OR2 (N25254, N25250, N24283);
and AND4 (N25255, N25217, N6442, N9059, N15242);
not NOT1 (N25256, N25236);
not NOT1 (N25257, N25255);
xor XOR2 (N25258, N25251, N20405);
nand NAND4 (N25259, N25253, N24921, N21286, N24049);
and AND4 (N25260, N25237, N19014, N6573, N2234);
or OR3 (N25261, N25259, N14918, N15232);
and AND2 (N25262, N25241, N24681);
nand NAND4 (N25263, N25262, N23147, N11059, N14724);
xor XOR2 (N25264, N25200, N4545);
xor XOR2 (N25265, N25260, N11660);
buf BUF1 (N25266, N25265);
or OR4 (N25267, N25264, N8524, N3987, N6550);
and AND4 (N25268, N25267, N23739, N7590, N15505);
or OR2 (N25269, N25261, N10034);
or OR4 (N25270, N25263, N19134, N13477, N18891);
xor XOR2 (N25271, N25257, N11547);
nand NAND3 (N25272, N25254, N23876, N13335);
nor NOR2 (N25273, N25272, N17214);
buf BUF1 (N25274, N25269);
not NOT1 (N25275, N25258);
buf BUF1 (N25276, N25275);
not NOT1 (N25277, N25268);
and AND3 (N25278, N25270, N5253, N11477);
buf BUF1 (N25279, N25247);
xor XOR2 (N25280, N25256, N16480);
not NOT1 (N25281, N25279);
xor XOR2 (N25282, N25278, N13012);
not NOT1 (N25283, N25276);
buf BUF1 (N25284, N25283);
not NOT1 (N25285, N25277);
xor XOR2 (N25286, N25280, N22785);
or OR2 (N25287, N25285, N12300);
and AND3 (N25288, N25286, N23985, N3977);
and AND2 (N25289, N25249, N6510);
buf BUF1 (N25290, N25274);
nor NOR3 (N25291, N25290, N18210, N9494);
nor NOR3 (N25292, N25266, N14416, N14834);
not NOT1 (N25293, N25273);
and AND4 (N25294, N25292, N24558, N7607, N3461);
nand NAND4 (N25295, N25287, N22731, N10203, N2074);
nor NOR3 (N25296, N25282, N24467, N5682);
nand NAND4 (N25297, N25295, N20308, N14673, N18448);
nand NAND3 (N25298, N25271, N8950, N4260);
buf BUF1 (N25299, N25293);
or OR3 (N25300, N25284, N13230, N21218);
and AND4 (N25301, N25299, N1053, N21231, N12694);
nand NAND3 (N25302, N25289, N16329, N18348);
nor NOR2 (N25303, N25302, N11509);
nand NAND2 (N25304, N25300, N21574);
buf BUF1 (N25305, N25303);
and AND4 (N25306, N25297, N6438, N1447, N18536);
and AND4 (N25307, N25304, N5632, N13650, N5449);
and AND2 (N25308, N25296, N16359);
not NOT1 (N25309, N25306);
not NOT1 (N25310, N25305);
nand NAND3 (N25311, N25301, N11366, N20211);
xor XOR2 (N25312, N25309, N6666);
xor XOR2 (N25313, N25298, N15604);
not NOT1 (N25314, N25291);
nor NOR2 (N25315, N25288, N8058);
not NOT1 (N25316, N25312);
and AND3 (N25317, N25313, N24180, N4548);
or OR2 (N25318, N25307, N17440);
or OR3 (N25319, N25294, N6191, N12885);
not NOT1 (N25320, N25310);
nand NAND4 (N25321, N25315, N1386, N10234, N22307);
and AND4 (N25322, N25318, N3129, N12230, N1720);
xor XOR2 (N25323, N25319, N5011);
xor XOR2 (N25324, N25314, N11727);
and AND3 (N25325, N25320, N1616, N10548);
xor XOR2 (N25326, N25321, N16945);
nand NAND3 (N25327, N25326, N14454, N17628);
xor XOR2 (N25328, N25281, N1853);
nor NOR3 (N25329, N25323, N17438, N24050);
or OR3 (N25330, N25316, N1330, N8370);
nor NOR3 (N25331, N25327, N1442, N9024);
or OR2 (N25332, N25322, N22491);
not NOT1 (N25333, N25330);
or OR4 (N25334, N25311, N8472, N13434, N19828);
or OR3 (N25335, N25328, N11387, N19874);
nand NAND4 (N25336, N25317, N22300, N4815, N15781);
nand NAND3 (N25337, N25334, N2497, N16185);
nand NAND4 (N25338, N25336, N9042, N10363, N18346);
or OR2 (N25339, N25331, N7368);
nor NOR3 (N25340, N25332, N11338, N19634);
nor NOR4 (N25341, N25338, N8259, N12921, N12993);
nor NOR2 (N25342, N25333, N12514);
and AND2 (N25343, N25339, N23613);
xor XOR2 (N25344, N25337, N21288);
and AND3 (N25345, N25342, N9065, N11017);
buf BUF1 (N25346, N25340);
nor NOR2 (N25347, N25344, N11302);
or OR3 (N25348, N25346, N3329, N10812);
xor XOR2 (N25349, N25341, N2879);
and AND4 (N25350, N25335, N8240, N13730, N24067);
xor XOR2 (N25351, N25345, N6353);
xor XOR2 (N25352, N25349, N17364);
buf BUF1 (N25353, N25308);
nor NOR4 (N25354, N25352, N14461, N16917, N15292);
xor XOR2 (N25355, N25348, N17295);
not NOT1 (N25356, N25350);
buf BUF1 (N25357, N25356);
or OR2 (N25358, N25354, N2763);
nand NAND3 (N25359, N25347, N9310, N13736);
nand NAND4 (N25360, N25343, N1411, N17708, N2243);
and AND3 (N25361, N25324, N15135, N9009);
buf BUF1 (N25362, N25355);
or OR4 (N25363, N25357, N1344, N2115, N24355);
not NOT1 (N25364, N25325);
not NOT1 (N25365, N25363);
or OR4 (N25366, N25351, N20359, N21847, N443);
and AND3 (N25367, N25329, N1349, N5239);
nand NAND4 (N25368, N25359, N6511, N16816, N24337);
buf BUF1 (N25369, N25368);
xor XOR2 (N25370, N25366, N13318);
buf BUF1 (N25371, N25369);
buf BUF1 (N25372, N25367);
or OR3 (N25373, N25358, N1402, N12356);
and AND4 (N25374, N25353, N3478, N1955, N153);
nor NOR4 (N25375, N25373, N15807, N8458, N25253);
not NOT1 (N25376, N25362);
and AND4 (N25377, N25364, N21076, N7573, N7986);
xor XOR2 (N25378, N25377, N12265);
buf BUF1 (N25379, N25376);
nand NAND2 (N25380, N25361, N9840);
buf BUF1 (N25381, N25375);
and AND2 (N25382, N25381, N24322);
buf BUF1 (N25383, N25360);
nor NOR2 (N25384, N25371, N16218);
buf BUF1 (N25385, N25380);
nand NAND2 (N25386, N25370, N12747);
or OR3 (N25387, N25365, N23839, N5178);
xor XOR2 (N25388, N25387, N3465);
xor XOR2 (N25389, N25386, N355);
or OR2 (N25390, N25382, N4707);
nand NAND3 (N25391, N25372, N19235, N8168);
buf BUF1 (N25392, N25389);
nand NAND2 (N25393, N25379, N2922);
nor NOR3 (N25394, N25393, N19321, N21978);
not NOT1 (N25395, N25392);
nand NAND2 (N25396, N25383, N15811);
and AND2 (N25397, N25394, N18337);
nand NAND3 (N25398, N25395, N22585, N20477);
or OR4 (N25399, N25385, N15885, N21187, N6978);
nand NAND2 (N25400, N25391, N20728);
nor NOR3 (N25401, N25397, N20963, N24555);
nand NAND4 (N25402, N25388, N12301, N16736, N3244);
or OR2 (N25403, N25399, N20952);
or OR4 (N25404, N25378, N1906, N23113, N1262);
nor NOR4 (N25405, N25396, N19243, N23821, N10481);
or OR2 (N25406, N25401, N24421);
nor NOR2 (N25407, N25406, N19528);
and AND3 (N25408, N25384, N21279, N14969);
nor NOR2 (N25409, N25407, N19373);
not NOT1 (N25410, N25404);
not NOT1 (N25411, N25400);
xor XOR2 (N25412, N25374, N5558);
xor XOR2 (N25413, N25398, N9727);
or OR3 (N25414, N25402, N8800, N4803);
nor NOR2 (N25415, N25411, N7453);
nand NAND3 (N25416, N25405, N14247, N5579);
buf BUF1 (N25417, N25414);
nor NOR4 (N25418, N25413, N18179, N8745, N5940);
nor NOR4 (N25419, N25408, N22314, N20495, N8660);
buf BUF1 (N25420, N25416);
xor XOR2 (N25421, N25409, N13078);
nand NAND4 (N25422, N25420, N25169, N21760, N24194);
not NOT1 (N25423, N25421);
or OR4 (N25424, N25390, N24404, N964, N12100);
not NOT1 (N25425, N25418);
and AND4 (N25426, N25419, N15618, N22017, N16506);
nand NAND2 (N25427, N25423, N24742);
or OR2 (N25428, N25415, N12569);
not NOT1 (N25429, N25425);
buf BUF1 (N25430, N25428);
not NOT1 (N25431, N25424);
nor NOR3 (N25432, N25422, N24856, N5112);
buf BUF1 (N25433, N25417);
buf BUF1 (N25434, N25431);
not NOT1 (N25435, N25410);
nor NOR2 (N25436, N25412, N17054);
nand NAND3 (N25437, N25432, N7097, N19938);
nand NAND2 (N25438, N25403, N605);
not NOT1 (N25439, N25435);
not NOT1 (N25440, N25434);
nor NOR3 (N25441, N25429, N7215, N3786);
buf BUF1 (N25442, N25438);
nand NAND4 (N25443, N25430, N15562, N922, N21029);
buf BUF1 (N25444, N25427);
xor XOR2 (N25445, N25437, N16402);
and AND4 (N25446, N25444, N7292, N5289, N9389);
and AND4 (N25447, N25439, N10539, N5463, N5202);
nand NAND2 (N25448, N25447, N25144);
nand NAND4 (N25449, N25440, N20120, N1565, N6139);
buf BUF1 (N25450, N25436);
nand NAND2 (N25451, N25442, N18585);
nor NOR4 (N25452, N25451, N13623, N22776, N23084);
or OR2 (N25453, N25446, N16669);
nand NAND2 (N25454, N25441, N6932);
and AND4 (N25455, N25443, N7024, N18219, N9816);
not NOT1 (N25456, N25453);
nand NAND4 (N25457, N25449, N10983, N14804, N12413);
nand NAND3 (N25458, N25445, N10137, N13360);
not NOT1 (N25459, N25426);
xor XOR2 (N25460, N25457, N15216);
xor XOR2 (N25461, N25460, N5279);
nor NOR4 (N25462, N25454, N19697, N21537, N22580);
xor XOR2 (N25463, N25461, N23654);
nor NOR4 (N25464, N25450, N13084, N5251, N3247);
or OR2 (N25465, N25464, N5599);
not NOT1 (N25466, N25455);
buf BUF1 (N25467, N25456);
xor XOR2 (N25468, N25467, N9923);
buf BUF1 (N25469, N25459);
or OR3 (N25470, N25462, N4978, N7161);
nand NAND2 (N25471, N25468, N12674);
nor NOR2 (N25472, N25452, N11596);
buf BUF1 (N25473, N25463);
xor XOR2 (N25474, N25433, N1338);
nand NAND3 (N25475, N25466, N18619, N17527);
nor NOR4 (N25476, N25475, N21830, N17760, N14065);
not NOT1 (N25477, N25465);
xor XOR2 (N25478, N25470, N16086);
and AND4 (N25479, N25471, N17673, N11037, N374);
nor NOR4 (N25480, N25477, N12657, N17447, N22543);
nand NAND2 (N25481, N25474, N11333);
buf BUF1 (N25482, N25469);
or OR4 (N25483, N25458, N19523, N830, N12238);
buf BUF1 (N25484, N25476);
xor XOR2 (N25485, N25479, N18064);
buf BUF1 (N25486, N25481);
not NOT1 (N25487, N25472);
buf BUF1 (N25488, N25483);
or OR2 (N25489, N25487, N3473);
nor NOR4 (N25490, N25486, N19110, N5781, N23225);
nor NOR3 (N25491, N25480, N6834, N6090);
nand NAND4 (N25492, N25489, N2158, N20639, N20372);
or OR2 (N25493, N25485, N5385);
or OR2 (N25494, N25493, N5148);
not NOT1 (N25495, N25484);
nand NAND4 (N25496, N25482, N13779, N17392, N4597);
nand NAND2 (N25497, N25491, N20442);
or OR3 (N25498, N25497, N4096, N4709);
not NOT1 (N25499, N25492);
or OR3 (N25500, N25498, N12479, N5624);
or OR3 (N25501, N25494, N20297, N19916);
nand NAND4 (N25502, N25496, N20515, N9929, N11003);
and AND3 (N25503, N25495, N1166, N4516);
not NOT1 (N25504, N25503);
not NOT1 (N25505, N25473);
buf BUF1 (N25506, N25499);
or OR4 (N25507, N25502, N5488, N8683, N11274);
and AND3 (N25508, N25501, N20678, N19233);
and AND2 (N25509, N25448, N14442);
or OR2 (N25510, N25478, N22045);
buf BUF1 (N25511, N25505);
xor XOR2 (N25512, N25490, N9626);
and AND3 (N25513, N25507, N24157, N767);
nor NOR3 (N25514, N25488, N5546, N13668);
or OR2 (N25515, N25510, N3761);
and AND2 (N25516, N25509, N18192);
nand NAND2 (N25517, N25508, N1029);
buf BUF1 (N25518, N25513);
nor NOR2 (N25519, N25500, N341);
nor NOR4 (N25520, N25517, N10900, N2268, N19788);
and AND2 (N25521, N25514, N7252);
nand NAND2 (N25522, N25519, N14133);
nor NOR4 (N25523, N25518, N2093, N3796, N19004);
and AND4 (N25524, N25504, N13276, N10387, N6234);
nor NOR2 (N25525, N25511, N17253);
xor XOR2 (N25526, N25512, N14754);
and AND2 (N25527, N25522, N15066);
and AND3 (N25528, N25521, N8017, N21147);
nor NOR3 (N25529, N25527, N3163, N23227);
not NOT1 (N25530, N25523);
or OR4 (N25531, N25506, N5523, N10286, N13172);
buf BUF1 (N25532, N25531);
and AND3 (N25533, N25525, N3934, N7145);
nand NAND3 (N25534, N25515, N2867, N19649);
xor XOR2 (N25535, N25529, N16039);
not NOT1 (N25536, N25534);
xor XOR2 (N25537, N25530, N25438);
nand NAND4 (N25538, N25528, N11004, N18194, N21238);
nor NOR3 (N25539, N25538, N15259, N316);
xor XOR2 (N25540, N25524, N18519);
or OR2 (N25541, N25520, N16923);
nand NAND2 (N25542, N25535, N3588);
nor NOR2 (N25543, N25537, N14549);
not NOT1 (N25544, N25526);
nand NAND3 (N25545, N25544, N8916, N2070);
buf BUF1 (N25546, N25542);
and AND2 (N25547, N25532, N5570);
or OR2 (N25548, N25541, N2207);
or OR3 (N25549, N25540, N21461, N18411);
or OR2 (N25550, N25539, N24972);
buf BUF1 (N25551, N25536);
nand NAND3 (N25552, N25547, N21972, N21206);
not NOT1 (N25553, N25549);
and AND2 (N25554, N25552, N12321);
buf BUF1 (N25555, N25554);
not NOT1 (N25556, N25533);
or OR3 (N25557, N25548, N3730, N2543);
buf BUF1 (N25558, N25543);
and AND4 (N25559, N25555, N4979, N4231, N6990);
or OR4 (N25560, N25559, N1211, N21601, N8062);
and AND4 (N25561, N25560, N6145, N23278, N5911);
nand NAND2 (N25562, N25556, N13857);
nor NOR2 (N25563, N25562, N560);
not NOT1 (N25564, N25545);
and AND2 (N25565, N25557, N17087);
buf BUF1 (N25566, N25550);
xor XOR2 (N25567, N25561, N1073);
not NOT1 (N25568, N25553);
nand NAND4 (N25569, N25566, N3004, N13818, N12183);
or OR3 (N25570, N25569, N22500, N13467);
and AND3 (N25571, N25516, N18574, N1440);
nor NOR4 (N25572, N25564, N17969, N22901, N22538);
nand NAND4 (N25573, N25568, N23973, N14077, N2108);
not NOT1 (N25574, N25551);
or OR3 (N25575, N25565, N11808, N18822);
and AND4 (N25576, N25574, N4727, N15393, N19383);
buf BUF1 (N25577, N25571);
not NOT1 (N25578, N25563);
buf BUF1 (N25579, N25558);
buf BUF1 (N25580, N25577);
nor NOR4 (N25581, N25572, N9188, N15739, N20054);
or OR4 (N25582, N25576, N1621, N6889, N17913);
buf BUF1 (N25583, N25546);
or OR3 (N25584, N25578, N14485, N7870);
not NOT1 (N25585, N25582);
and AND2 (N25586, N25573, N24213);
or OR3 (N25587, N25579, N6644, N8720);
buf BUF1 (N25588, N25584);
not NOT1 (N25589, N25575);
or OR3 (N25590, N25588, N11185, N25086);
xor XOR2 (N25591, N25570, N24797);
not NOT1 (N25592, N25585);
not NOT1 (N25593, N25591);
xor XOR2 (N25594, N25593, N4475);
buf BUF1 (N25595, N25586);
xor XOR2 (N25596, N25583, N22664);
not NOT1 (N25597, N25594);
buf BUF1 (N25598, N25595);
nand NAND4 (N25599, N25598, N2114, N18843, N4776);
not NOT1 (N25600, N25580);
not NOT1 (N25601, N25590);
xor XOR2 (N25602, N25597, N21401);
and AND3 (N25603, N25600, N7948, N12758);
nor NOR2 (N25604, N25602, N5473);
or OR2 (N25605, N25603, N1597);
and AND4 (N25606, N25596, N21587, N15300, N4758);
buf BUF1 (N25607, N25599);
xor XOR2 (N25608, N25604, N18743);
not NOT1 (N25609, N25592);
xor XOR2 (N25610, N25587, N19936);
nor NOR4 (N25611, N25608, N24506, N17284, N15888);
not NOT1 (N25612, N25609);
nand NAND3 (N25613, N25589, N8224, N22253);
nand NAND2 (N25614, N25567, N12044);
and AND3 (N25615, N25613, N18128, N5839);
xor XOR2 (N25616, N25606, N3966);
and AND3 (N25617, N25612, N4994, N2248);
and AND3 (N25618, N25615, N5082, N4428);
buf BUF1 (N25619, N25610);
buf BUF1 (N25620, N25618);
nor NOR4 (N25621, N25607, N17093, N4350, N9263);
nand NAND2 (N25622, N25616, N13507);
and AND2 (N25623, N25614, N15423);
not NOT1 (N25624, N25601);
not NOT1 (N25625, N25622);
nand NAND2 (N25626, N25623, N23440);
xor XOR2 (N25627, N25625, N3765);
nor NOR4 (N25628, N25611, N16846, N15046, N5792);
xor XOR2 (N25629, N25621, N5013);
and AND4 (N25630, N25617, N11913, N3700, N23538);
and AND4 (N25631, N25620, N13098, N23928, N1767);
xor XOR2 (N25632, N25581, N4534);
buf BUF1 (N25633, N25632);
not NOT1 (N25634, N25631);
and AND4 (N25635, N25633, N4364, N9692, N7495);
nor NOR3 (N25636, N25605, N103, N20799);
not NOT1 (N25637, N25635);
and AND2 (N25638, N25624, N14329);
and AND3 (N25639, N25628, N18133, N177);
nand NAND3 (N25640, N25634, N724, N9044);
and AND3 (N25641, N25639, N10113, N538);
buf BUF1 (N25642, N25626);
buf BUF1 (N25643, N25637);
buf BUF1 (N25644, N25630);
buf BUF1 (N25645, N25638);
not NOT1 (N25646, N25644);
xor XOR2 (N25647, N25641, N23999);
or OR3 (N25648, N25636, N24214, N16201);
not NOT1 (N25649, N25642);
or OR4 (N25650, N25648, N2573, N15570, N12717);
and AND4 (N25651, N25627, N12750, N14054, N7722);
and AND3 (N25652, N25619, N7257, N15046);
or OR3 (N25653, N25651, N9891, N23574);
buf BUF1 (N25654, N25640);
and AND2 (N25655, N25645, N18324);
nand NAND2 (N25656, N25647, N7803);
nor NOR2 (N25657, N25652, N24485);
nand NAND3 (N25658, N25646, N19132, N843);
nand NAND2 (N25659, N25643, N14396);
or OR4 (N25660, N25653, N10790, N22979, N2386);
or OR3 (N25661, N25656, N20264, N6841);
buf BUF1 (N25662, N25660);
not NOT1 (N25663, N25650);
nand NAND3 (N25664, N25629, N6810, N2102);
xor XOR2 (N25665, N25663, N20893);
xor XOR2 (N25666, N25654, N8658);
buf BUF1 (N25667, N25657);
or OR3 (N25668, N25659, N5552, N2798);
xor XOR2 (N25669, N25658, N8875);
xor XOR2 (N25670, N25668, N10399);
nor NOR2 (N25671, N25670, N1444);
nand NAND3 (N25672, N25671, N25179, N20869);
xor XOR2 (N25673, N25661, N5322);
nor NOR3 (N25674, N25665, N22093, N1215);
and AND4 (N25675, N25673, N22280, N22955, N584);
nand NAND2 (N25676, N25662, N14028);
xor XOR2 (N25677, N25664, N13701);
or OR4 (N25678, N25666, N15335, N11068, N11192);
and AND2 (N25679, N25672, N23138);
not NOT1 (N25680, N25655);
and AND3 (N25681, N25678, N2752, N7335);
nand NAND2 (N25682, N25680, N22457);
nor NOR2 (N25683, N25674, N7086);
nand NAND4 (N25684, N25667, N23159, N10018, N819);
buf BUF1 (N25685, N25679);
buf BUF1 (N25686, N25676);
not NOT1 (N25687, N25682);
and AND2 (N25688, N25684, N1502);
xor XOR2 (N25689, N25688, N9606);
nand NAND4 (N25690, N25669, N22176, N12133, N20269);
nand NAND2 (N25691, N25683, N19251);
xor XOR2 (N25692, N25677, N14186);
nand NAND4 (N25693, N25692, N1892, N22774, N8997);
nor NOR3 (N25694, N25690, N13511, N9254);
xor XOR2 (N25695, N25686, N25376);
or OR3 (N25696, N25691, N22295, N12384);
nand NAND2 (N25697, N25695, N6605);
nor NOR2 (N25698, N25693, N6452);
not NOT1 (N25699, N25698);
nand NAND2 (N25700, N25694, N9103);
buf BUF1 (N25701, N25687);
buf BUF1 (N25702, N25675);
xor XOR2 (N25703, N25685, N9616);
not NOT1 (N25704, N25681);
not NOT1 (N25705, N25689);
nand NAND3 (N25706, N25703, N24539, N6072);
and AND3 (N25707, N25697, N2937, N4195);
xor XOR2 (N25708, N25649, N338);
and AND3 (N25709, N25700, N13005, N13407);
buf BUF1 (N25710, N25707);
not NOT1 (N25711, N25699);
nor NOR2 (N25712, N25696, N452);
nor NOR3 (N25713, N25704, N25342, N2854);
xor XOR2 (N25714, N25702, N8749);
and AND4 (N25715, N25708, N7561, N12745, N221);
xor XOR2 (N25716, N25701, N14443);
not NOT1 (N25717, N25716);
nor NOR4 (N25718, N25712, N15465, N16029, N24265);
not NOT1 (N25719, N25717);
or OR2 (N25720, N25719, N6766);
xor XOR2 (N25721, N25711, N1150);
or OR4 (N25722, N25706, N16913, N19480, N10018);
buf BUF1 (N25723, N25713);
or OR2 (N25724, N25715, N10041);
not NOT1 (N25725, N25718);
or OR3 (N25726, N25710, N17949, N14183);
nor NOR3 (N25727, N25714, N12530, N991);
nand NAND4 (N25728, N25720, N25201, N15563, N19678);
nand NAND2 (N25729, N25725, N6884);
and AND2 (N25730, N25705, N9876);
or OR2 (N25731, N25727, N11138);
buf BUF1 (N25732, N25729);
or OR3 (N25733, N25723, N10508, N19555);
buf BUF1 (N25734, N25726);
and AND4 (N25735, N25734, N2801, N2707, N2266);
xor XOR2 (N25736, N25733, N4001);
buf BUF1 (N25737, N25732);
buf BUF1 (N25738, N25709);
buf BUF1 (N25739, N25737);
buf BUF1 (N25740, N25730);
not NOT1 (N25741, N25739);
or OR3 (N25742, N25738, N21645, N19883);
buf BUF1 (N25743, N25728);
nand NAND4 (N25744, N25741, N8777, N8996, N18255);
or OR2 (N25745, N25742, N13887);
nand NAND2 (N25746, N25744, N8665);
not NOT1 (N25747, N25735);
not NOT1 (N25748, N25747);
nand NAND2 (N25749, N25731, N16726);
nor NOR2 (N25750, N25746, N24765);
nor NOR3 (N25751, N25740, N22864, N12044);
not NOT1 (N25752, N25751);
or OR3 (N25753, N25745, N14863, N13145);
buf BUF1 (N25754, N25724);
nand NAND2 (N25755, N25749, N15999);
and AND3 (N25756, N25755, N1282, N7285);
nor NOR2 (N25757, N25748, N17044);
or OR4 (N25758, N25750, N3470, N14449, N6894);
or OR4 (N25759, N25754, N13479, N25281, N3237);
and AND4 (N25760, N25736, N12262, N5452, N23384);
nor NOR4 (N25761, N25757, N2765, N3499, N3913);
nand NAND2 (N25762, N25722, N22756);
nand NAND3 (N25763, N25743, N21693, N30);
nor NOR3 (N25764, N25760, N13371, N2962);
and AND3 (N25765, N25721, N15053, N2895);
nand NAND2 (N25766, N25759, N7841);
nand NAND3 (N25767, N25753, N4408, N5921);
and AND4 (N25768, N25752, N761, N14406, N22796);
nor NOR2 (N25769, N25764, N16562);
buf BUF1 (N25770, N25765);
nor NOR4 (N25771, N25761, N9838, N4641, N14142);
nand NAND3 (N25772, N25756, N1546, N16774);
or OR3 (N25773, N25758, N9276, N1656);
not NOT1 (N25774, N25766);
xor XOR2 (N25775, N25767, N7203);
buf BUF1 (N25776, N25769);
and AND4 (N25777, N25770, N20374, N14336, N11932);
xor XOR2 (N25778, N25774, N13059);
and AND3 (N25779, N25777, N10021, N12567);
or OR4 (N25780, N25776, N16850, N14864, N1720);
nand NAND4 (N25781, N25780, N13416, N3522, N22116);
xor XOR2 (N25782, N25771, N5773);
not NOT1 (N25783, N25773);
and AND4 (N25784, N25783, N11512, N19426, N8486);
and AND2 (N25785, N25775, N11814);
xor XOR2 (N25786, N25785, N18241);
nor NOR2 (N25787, N25763, N1985);
or OR3 (N25788, N25768, N11254, N21973);
or OR2 (N25789, N25778, N9210);
buf BUF1 (N25790, N25762);
and AND4 (N25791, N25789, N20919, N6761, N2299);
not NOT1 (N25792, N25772);
xor XOR2 (N25793, N25788, N8116);
nor NOR2 (N25794, N25784, N24546);
not NOT1 (N25795, N25790);
nor NOR2 (N25796, N25793, N20090);
and AND3 (N25797, N25791, N23561, N8143);
xor XOR2 (N25798, N25797, N9473);
not NOT1 (N25799, N25786);
not NOT1 (N25800, N25799);
nor NOR4 (N25801, N25782, N8832, N4911, N5263);
nand NAND4 (N25802, N25795, N15041, N9317, N2084);
or OR3 (N25803, N25800, N6747, N12352);
xor XOR2 (N25804, N25794, N7463);
nand NAND4 (N25805, N25803, N4383, N6688, N11755);
xor XOR2 (N25806, N25779, N24732);
xor XOR2 (N25807, N25787, N25363);
nor NOR2 (N25808, N25806, N5672);
nand NAND2 (N25809, N25798, N24394);
nor NOR2 (N25810, N25805, N10920);
nand NAND4 (N25811, N25807, N9719, N17195, N11894);
buf BUF1 (N25812, N25792);
or OR4 (N25813, N25801, N16508, N9786, N23843);
nor NOR4 (N25814, N25804, N18718, N24819, N13551);
and AND4 (N25815, N25811, N15814, N15972, N18982);
xor XOR2 (N25816, N25802, N7033);
nand NAND4 (N25817, N25813, N25125, N571, N3059);
nand NAND3 (N25818, N25810, N20584, N5615);
nor NOR4 (N25819, N25808, N2168, N21123, N1112);
xor XOR2 (N25820, N25812, N19386);
and AND4 (N25821, N25814, N24316, N14286, N9953);
buf BUF1 (N25822, N25796);
nand NAND2 (N25823, N25822, N18555);
nand NAND2 (N25824, N25815, N23641);
nor NOR2 (N25825, N25818, N11111);
and AND4 (N25826, N25821, N22891, N598, N12142);
not NOT1 (N25827, N25819);
xor XOR2 (N25828, N25820, N9958);
or OR3 (N25829, N25824, N18116, N22901);
or OR4 (N25830, N25816, N13995, N1888, N312);
and AND2 (N25831, N25823, N18650);
not NOT1 (N25832, N25825);
nor NOR3 (N25833, N25831, N10056, N7316);
and AND3 (N25834, N25832, N11746, N2563);
nor NOR3 (N25835, N25781, N10854, N13774);
or OR2 (N25836, N25828, N7408);
and AND3 (N25837, N25836, N9878, N7696);
not NOT1 (N25838, N25826);
xor XOR2 (N25839, N25835, N16412);
xor XOR2 (N25840, N25834, N1132);
and AND2 (N25841, N25839, N21184);
nand NAND2 (N25842, N25837, N17733);
buf BUF1 (N25843, N25809);
nor NOR3 (N25844, N25841, N21766, N4410);
buf BUF1 (N25845, N25817);
xor XOR2 (N25846, N25838, N1145);
nand NAND2 (N25847, N25845, N5368);
xor XOR2 (N25848, N25844, N10481);
nand NAND2 (N25849, N25829, N2140);
or OR3 (N25850, N25833, N18297, N24932);
or OR2 (N25851, N25827, N11752);
xor XOR2 (N25852, N25851, N17321);
and AND3 (N25853, N25849, N6355, N3201);
buf BUF1 (N25854, N25840);
xor XOR2 (N25855, N25846, N16197);
nor NOR3 (N25856, N25852, N16116, N8778);
and AND2 (N25857, N25854, N25505);
xor XOR2 (N25858, N25830, N17626);
nand NAND3 (N25859, N25855, N9201, N10457);
or OR3 (N25860, N25842, N6737, N9515);
buf BUF1 (N25861, N25843);
and AND4 (N25862, N25857, N9897, N19414, N7085);
and AND2 (N25863, N25860, N19088);
nor NOR2 (N25864, N25863, N409);
nor NOR4 (N25865, N25862, N8117, N24676, N22019);
nand NAND2 (N25866, N25847, N17384);
buf BUF1 (N25867, N25858);
or OR4 (N25868, N25848, N11892, N15260, N24806);
not NOT1 (N25869, N25864);
not NOT1 (N25870, N25869);
and AND3 (N25871, N25853, N25562, N15117);
buf BUF1 (N25872, N25865);
not NOT1 (N25873, N25868);
or OR3 (N25874, N25861, N23846, N6632);
or OR2 (N25875, N25850, N3471);
not NOT1 (N25876, N25856);
nor NOR2 (N25877, N25871, N7418);
and AND4 (N25878, N25876, N23613, N21684, N23473);
xor XOR2 (N25879, N25870, N3562);
nor NOR3 (N25880, N25878, N21502, N24946);
not NOT1 (N25881, N25880);
nor NOR3 (N25882, N25877, N7851, N5067);
or OR2 (N25883, N25875, N11181);
nor NOR2 (N25884, N25879, N13905);
nor NOR2 (N25885, N25884, N22280);
or OR4 (N25886, N25859, N4384, N6345, N3984);
or OR4 (N25887, N25882, N18894, N19554, N13342);
buf BUF1 (N25888, N25883);
not NOT1 (N25889, N25866);
and AND3 (N25890, N25889, N15390, N11745);
xor XOR2 (N25891, N25867, N3823);
nor NOR2 (N25892, N25891, N16560);
nor NOR3 (N25893, N25872, N1119, N3435);
nor NOR4 (N25894, N25886, N17676, N17497, N15007);
or OR3 (N25895, N25881, N14356, N18283);
or OR2 (N25896, N25893, N11821);
buf BUF1 (N25897, N25874);
nand NAND3 (N25898, N25896, N1630, N25299);
and AND2 (N25899, N25892, N10117);
and AND2 (N25900, N25899, N15025);
nand NAND4 (N25901, N25897, N22900, N297, N21324);
buf BUF1 (N25902, N25895);
nand NAND3 (N25903, N25888, N20699, N2338);
or OR2 (N25904, N25903, N8568);
or OR3 (N25905, N25901, N13670, N16486);
nand NAND4 (N25906, N25905, N5364, N9569, N15222);
nand NAND4 (N25907, N25873, N9774, N15797, N202);
buf BUF1 (N25908, N25900);
xor XOR2 (N25909, N25908, N17103);
buf BUF1 (N25910, N25887);
and AND3 (N25911, N25909, N17193, N24134);
buf BUF1 (N25912, N25904);
nor NOR4 (N25913, N25910, N20201, N10504, N7127);
and AND3 (N25914, N25890, N15585, N21118);
and AND3 (N25915, N25907, N6990, N13247);
endmodule