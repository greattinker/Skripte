// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21;

output N2514,N2502,N2503,N2520,N2505,N2511,N2513,N2516,N2519,N2521;

not NOT1 (N22, N11);
xor XOR2 (N23, N21, N3);
and AND4 (N24, N7, N20, N3, N17);
buf BUF1 (N25, N24);
buf BUF1 (N26, N17);
buf BUF1 (N27, N25);
xor XOR2 (N28, N2, N27);
or OR4 (N29, N6, N3, N10, N9);
or OR3 (N30, N14, N16, N1);
nor NOR4 (N31, N27, N10, N24, N18);
nand NAND2 (N32, N22, N8);
nand NAND4 (N33, N30, N16, N25, N4);
nand NAND4 (N34, N2, N12, N9, N2);
or OR3 (N35, N21, N14, N5);
xor XOR2 (N36, N15, N33);
nor NOR4 (N37, N30, N6, N5, N1);
nor NOR4 (N38, N23, N35, N23, N30);
nand NAND3 (N39, N27, N17, N2);
not NOT1 (N40, N29);
not NOT1 (N41, N31);
nand NAND4 (N42, N37, N29, N30, N24);
buf BUF1 (N43, N36);
and AND3 (N44, N28, N40, N40);
not NOT1 (N45, N27);
or OR3 (N46, N38, N17, N24);
or OR3 (N47, N45, N14, N43);
nor NOR4 (N48, N35, N1, N46, N27);
not NOT1 (N49, N4);
and AND4 (N50, N34, N46, N29, N1);
or OR4 (N51, N49, N3, N27, N41);
buf BUF1 (N52, N49);
or OR2 (N53, N48, N51);
nor NOR3 (N54, N23, N33, N34);
buf BUF1 (N55, N26);
buf BUF1 (N56, N39);
nor NOR4 (N57, N56, N47, N46, N15);
buf BUF1 (N58, N17);
or OR2 (N59, N32, N12);
or OR2 (N60, N52, N25);
buf BUF1 (N61, N60);
or OR3 (N62, N55, N45, N46);
xor XOR2 (N63, N59, N51);
and AND3 (N64, N54, N4, N57);
not NOT1 (N65, N11);
nand NAND3 (N66, N42, N32, N56);
nand NAND4 (N67, N50, N34, N41, N56);
nor NOR4 (N68, N66, N2, N56, N28);
or OR3 (N69, N67, N67, N62);
nor NOR3 (N70, N5, N18, N7);
buf BUF1 (N71, N65);
or OR3 (N72, N53, N31, N13);
not NOT1 (N73, N64);
not NOT1 (N74, N44);
or OR4 (N75, N70, N12, N20, N66);
not NOT1 (N76, N68);
and AND2 (N77, N63, N62);
or OR4 (N78, N71, N3, N59, N34);
xor XOR2 (N79, N77, N49);
and AND4 (N80, N58, N7, N7, N62);
or OR3 (N81, N78, N48, N29);
buf BUF1 (N82, N79);
nand NAND2 (N83, N61, N68);
nand NAND2 (N84, N81, N7);
and AND2 (N85, N84, N68);
nand NAND2 (N86, N80, N77);
and AND4 (N87, N73, N22, N70, N23);
and AND2 (N88, N85, N59);
or OR4 (N89, N76, N55, N11, N3);
or OR2 (N90, N86, N51);
not NOT1 (N91, N82);
buf BUF1 (N92, N90);
nand NAND4 (N93, N91, N35, N41, N68);
and AND3 (N94, N87, N62, N1);
xor XOR2 (N95, N92, N67);
and AND4 (N96, N95, N65, N46, N26);
and AND3 (N97, N94, N9, N74);
or OR4 (N98, N22, N45, N68, N83);
not NOT1 (N99, N28);
and AND4 (N100, N99, N21, N26, N6);
and AND3 (N101, N89, N99, N1);
and AND4 (N102, N101, N23, N35, N2);
buf BUF1 (N103, N72);
buf BUF1 (N104, N75);
nand NAND4 (N105, N102, N40, N37, N61);
and AND4 (N106, N98, N103, N91, N11);
or OR4 (N107, N53, N101, N79, N42);
nand NAND3 (N108, N88, N78, N71);
nor NOR2 (N109, N96, N3);
buf BUF1 (N110, N104);
or OR2 (N111, N109, N10);
xor XOR2 (N112, N93, N106);
nand NAND2 (N113, N19, N31);
and AND4 (N114, N97, N97, N12, N19);
and AND3 (N115, N105, N97, N103);
nand NAND2 (N116, N111, N27);
buf BUF1 (N117, N108);
and AND3 (N118, N114, N63, N55);
not NOT1 (N119, N107);
or OR2 (N120, N119, N87);
and AND3 (N121, N113, N112, N14);
nand NAND4 (N122, N36, N69, N66, N19);
buf BUF1 (N123, N29);
or OR3 (N124, N116, N4, N46);
or OR3 (N125, N121, N17, N121);
nand NAND3 (N126, N110, N33, N22);
xor XOR2 (N127, N117, N106);
xor XOR2 (N128, N115, N103);
and AND3 (N129, N120, N37, N88);
nand NAND4 (N130, N126, N95, N5, N48);
and AND2 (N131, N100, N55);
or OR4 (N132, N125, N115, N95, N63);
nor NOR4 (N133, N124, N43, N42, N68);
not NOT1 (N134, N127);
and AND2 (N135, N129, N12);
nor NOR3 (N136, N133, N1, N105);
buf BUF1 (N137, N136);
xor XOR2 (N138, N128, N84);
nand NAND2 (N139, N137, N56);
not NOT1 (N140, N118);
nand NAND2 (N141, N123, N32);
nor NOR2 (N142, N122, N65);
nor NOR4 (N143, N132, N133, N126, N28);
not NOT1 (N144, N140);
buf BUF1 (N145, N135);
or OR3 (N146, N143, N85, N56);
buf BUF1 (N147, N141);
and AND3 (N148, N142, N21, N78);
and AND2 (N149, N144, N69);
nor NOR2 (N150, N148, N136);
and AND4 (N151, N147, N61, N120, N80);
nand NAND4 (N152, N138, N120, N16, N44);
and AND3 (N153, N145, N15, N23);
buf BUF1 (N154, N152);
nand NAND3 (N155, N134, N2, N133);
not NOT1 (N156, N155);
buf BUF1 (N157, N130);
buf BUF1 (N158, N151);
and AND2 (N159, N139, N43);
not NOT1 (N160, N156);
and AND4 (N161, N157, N138, N88, N6);
not NOT1 (N162, N154);
nand NAND2 (N163, N131, N63);
and AND2 (N164, N146, N93);
buf BUF1 (N165, N149);
and AND4 (N166, N161, N24, N51, N103);
xor XOR2 (N167, N165, N165);
or OR3 (N168, N163, N142, N75);
not NOT1 (N169, N158);
nand NAND4 (N170, N168, N76, N158, N98);
xor XOR2 (N171, N150, N57);
and AND3 (N172, N164, N136, N97);
nor NOR4 (N173, N160, N16, N74, N141);
buf BUF1 (N174, N171);
xor XOR2 (N175, N174, N157);
xor XOR2 (N176, N173, N143);
nor NOR4 (N177, N169, N105, N140, N112);
nand NAND4 (N178, N153, N107, N16, N74);
xor XOR2 (N179, N178, N159);
nand NAND4 (N180, N102, N64, N25, N10);
not NOT1 (N181, N167);
and AND2 (N182, N180, N39);
and AND3 (N183, N176, N84, N119);
nor NOR3 (N184, N179, N138, N162);
xor XOR2 (N185, N132, N115);
buf BUF1 (N186, N184);
xor XOR2 (N187, N170, N64);
not NOT1 (N188, N175);
nand NAND2 (N189, N185, N129);
or OR2 (N190, N181, N24);
nand NAND2 (N191, N172, N95);
buf BUF1 (N192, N177);
buf BUF1 (N193, N186);
nand NAND4 (N194, N189, N188, N54, N54);
nand NAND3 (N195, N129, N178, N111);
or OR3 (N196, N193, N109, N179);
xor XOR2 (N197, N166, N41);
not NOT1 (N198, N192);
not NOT1 (N199, N196);
and AND4 (N200, N182, N147, N127, N63);
nor NOR3 (N201, N198, N141, N29);
not NOT1 (N202, N200);
nor NOR2 (N203, N183, N100);
nor NOR2 (N204, N197, N135);
xor XOR2 (N205, N191, N191);
nor NOR4 (N206, N204, N173, N61, N103);
buf BUF1 (N207, N187);
nand NAND3 (N208, N203, N88, N174);
not NOT1 (N209, N202);
or OR4 (N210, N195, N107, N142, N144);
buf BUF1 (N211, N205);
xor XOR2 (N212, N194, N58);
or OR2 (N213, N207, N148);
and AND4 (N214, N209, N96, N94, N183);
nand NAND2 (N215, N213, N100);
buf BUF1 (N216, N214);
buf BUF1 (N217, N208);
or OR4 (N218, N215, N136, N112, N78);
or OR4 (N219, N217, N12, N174, N68);
nor NOR2 (N220, N218, N196);
xor XOR2 (N221, N210, N29);
xor XOR2 (N222, N221, N5);
nor NOR3 (N223, N190, N124, N222);
not NOT1 (N224, N115);
or OR2 (N225, N199, N119);
not NOT1 (N226, N224);
or OR3 (N227, N225, N175, N141);
nor NOR2 (N228, N220, N49);
nor NOR2 (N229, N212, N177);
xor XOR2 (N230, N226, N35);
and AND4 (N231, N228, N83, N36, N7);
or OR4 (N232, N223, N46, N25, N28);
or OR4 (N233, N216, N8, N97, N66);
nand NAND4 (N234, N233, N202, N122, N208);
and AND3 (N235, N219, N224, N60);
xor XOR2 (N236, N235, N232);
or OR2 (N237, N61, N229);
xor XOR2 (N238, N214, N43);
xor XOR2 (N239, N211, N131);
nor NOR4 (N240, N230, N43, N109, N57);
or OR2 (N241, N238, N186);
xor XOR2 (N242, N206, N227);
buf BUF1 (N243, N173);
nand NAND3 (N244, N242, N8, N163);
or OR2 (N245, N237, N53);
or OR2 (N246, N231, N90);
xor XOR2 (N247, N236, N138);
nor NOR2 (N248, N234, N215);
buf BUF1 (N249, N247);
xor XOR2 (N250, N240, N108);
or OR3 (N251, N239, N185, N156);
buf BUF1 (N252, N250);
nand NAND2 (N253, N251, N49);
or OR2 (N254, N201, N167);
or OR2 (N255, N245, N242);
nor NOR4 (N256, N244, N232, N3, N67);
not NOT1 (N257, N241);
xor XOR2 (N258, N246, N58);
buf BUF1 (N259, N254);
buf BUF1 (N260, N259);
nor NOR4 (N261, N258, N142, N51, N19);
not NOT1 (N262, N257);
xor XOR2 (N263, N256, N1);
and AND3 (N264, N261, N12, N93);
not NOT1 (N265, N249);
and AND3 (N266, N255, N258, N240);
xor XOR2 (N267, N243, N42);
not NOT1 (N268, N260);
or OR3 (N269, N265, N164, N263);
and AND3 (N270, N122, N191, N44);
nor NOR4 (N271, N248, N252, N127, N158);
or OR4 (N272, N27, N199, N237, N217);
xor XOR2 (N273, N272, N164);
xor XOR2 (N274, N253, N142);
or OR3 (N275, N267, N104, N33);
nor NOR4 (N276, N271, N167, N198, N87);
nor NOR2 (N277, N276, N33);
or OR2 (N278, N266, N19);
and AND3 (N279, N262, N187, N241);
nand NAND2 (N280, N279, N234);
and AND2 (N281, N268, N127);
buf BUF1 (N282, N275);
xor XOR2 (N283, N269, N217);
or OR4 (N284, N280, N237, N273, N93);
not NOT1 (N285, N257);
nand NAND4 (N286, N270, N226, N129, N211);
not NOT1 (N287, N277);
xor XOR2 (N288, N282, N42);
nand NAND2 (N289, N284, N163);
and AND2 (N290, N281, N105);
or OR2 (N291, N287, N120);
and AND4 (N292, N290, N231, N224, N73);
buf BUF1 (N293, N286);
buf BUF1 (N294, N289);
xor XOR2 (N295, N283, N26);
xor XOR2 (N296, N264, N36);
xor XOR2 (N297, N291, N222);
nand NAND2 (N298, N293, N58);
nor NOR3 (N299, N297, N216, N64);
xor XOR2 (N300, N298, N22);
and AND4 (N301, N296, N8, N184, N99);
or OR2 (N302, N300, N205);
nand NAND2 (N303, N292, N88);
not NOT1 (N304, N301);
nor NOR4 (N305, N295, N175, N97, N241);
and AND4 (N306, N278, N41, N38, N257);
nor NOR4 (N307, N274, N253, N1, N66);
nor NOR2 (N308, N304, N7);
xor XOR2 (N309, N294, N307);
nand NAND3 (N310, N239, N129, N291);
not NOT1 (N311, N299);
xor XOR2 (N312, N305, N177);
buf BUF1 (N313, N303);
nor NOR4 (N314, N285, N223, N77, N306);
nand NAND3 (N315, N103, N222, N253);
buf BUF1 (N316, N312);
nand NAND3 (N317, N314, N89, N38);
nand NAND3 (N318, N316, N221, N83);
nor NOR2 (N319, N310, N79);
buf BUF1 (N320, N318);
xor XOR2 (N321, N302, N161);
buf BUF1 (N322, N308);
nand NAND2 (N323, N313, N205);
not NOT1 (N324, N321);
nor NOR4 (N325, N309, N198, N45, N3);
xor XOR2 (N326, N315, N200);
or OR2 (N327, N319, N285);
nor NOR3 (N328, N323, N58, N143);
buf BUF1 (N329, N288);
not NOT1 (N330, N327);
and AND4 (N331, N325, N180, N305, N279);
or OR4 (N332, N317, N207, N117, N49);
buf BUF1 (N333, N320);
nand NAND3 (N334, N328, N3, N22);
or OR4 (N335, N326, N276, N118, N259);
and AND3 (N336, N335, N277, N209);
or OR3 (N337, N330, N77, N253);
xor XOR2 (N338, N332, N95);
nor NOR2 (N339, N311, N191);
and AND3 (N340, N334, N92, N138);
nor NOR3 (N341, N338, N291, N296);
and AND4 (N342, N337, N335, N166, N283);
nor NOR3 (N343, N322, N67, N301);
or OR4 (N344, N342, N333, N298, N242);
and AND3 (N345, N261, N332, N141);
nand NAND4 (N346, N344, N333, N329, N138);
not NOT1 (N347, N289);
buf BUF1 (N348, N336);
xor XOR2 (N349, N346, N190);
xor XOR2 (N350, N348, N175);
buf BUF1 (N351, N341);
and AND2 (N352, N339, N214);
or OR3 (N353, N340, N318, N251);
xor XOR2 (N354, N349, N288);
buf BUF1 (N355, N343);
xor XOR2 (N356, N345, N113);
buf BUF1 (N357, N354);
nor NOR4 (N358, N357, N153, N110, N23);
or OR2 (N359, N352, N339);
and AND3 (N360, N331, N195, N167);
nor NOR4 (N361, N360, N286, N184, N1);
nand NAND2 (N362, N356, N151);
and AND3 (N363, N359, N270, N158);
buf BUF1 (N364, N358);
and AND3 (N365, N324, N176, N72);
nor NOR3 (N366, N350, N30, N168);
and AND4 (N367, N362, N254, N217, N28);
and AND2 (N368, N367, N60);
xor XOR2 (N369, N353, N320);
xor XOR2 (N370, N365, N228);
buf BUF1 (N371, N347);
buf BUF1 (N372, N370);
nand NAND4 (N373, N351, N42, N146, N192);
xor XOR2 (N374, N373, N345);
not NOT1 (N375, N372);
buf BUF1 (N376, N374);
and AND4 (N377, N361, N173, N100, N322);
or OR2 (N378, N355, N68);
not NOT1 (N379, N366);
not NOT1 (N380, N363);
and AND4 (N381, N380, N284, N106, N112);
nor NOR3 (N382, N368, N133, N179);
and AND4 (N383, N381, N313, N157, N69);
and AND3 (N384, N379, N37, N163);
or OR4 (N385, N378, N71, N373, N232);
nand NAND3 (N386, N371, N155, N226);
xor XOR2 (N387, N375, N190);
and AND3 (N388, N377, N216, N333);
or OR3 (N389, N386, N299, N17);
xor XOR2 (N390, N387, N176);
xor XOR2 (N391, N364, N89);
not NOT1 (N392, N391);
or OR2 (N393, N382, N285);
nor NOR4 (N394, N384, N329, N196, N339);
or OR2 (N395, N393, N377);
nor NOR3 (N396, N376, N296, N154);
xor XOR2 (N397, N395, N362);
not NOT1 (N398, N392);
not NOT1 (N399, N394);
and AND2 (N400, N383, N377);
not NOT1 (N401, N389);
or OR4 (N402, N397, N390, N169, N254);
not NOT1 (N403, N276);
nor NOR2 (N404, N403, N147);
nand NAND2 (N405, N400, N140);
xor XOR2 (N406, N369, N310);
nor NOR4 (N407, N385, N209, N21, N14);
and AND3 (N408, N401, N86, N189);
xor XOR2 (N409, N396, N43);
and AND2 (N410, N408, N86);
or OR2 (N411, N405, N163);
nand NAND3 (N412, N409, N233, N141);
not NOT1 (N413, N399);
or OR3 (N414, N412, N382, N19);
buf BUF1 (N415, N404);
and AND2 (N416, N415, N268);
xor XOR2 (N417, N402, N158);
and AND2 (N418, N417, N258);
nor NOR2 (N419, N414, N72);
and AND4 (N420, N413, N149, N224, N44);
buf BUF1 (N421, N411);
or OR3 (N422, N410, N393, N104);
buf BUF1 (N423, N418);
xor XOR2 (N424, N420, N77);
nand NAND2 (N425, N398, N225);
nor NOR2 (N426, N388, N61);
buf BUF1 (N427, N425);
xor XOR2 (N428, N423, N267);
xor XOR2 (N429, N426, N91);
buf BUF1 (N430, N419);
nand NAND4 (N431, N416, N425, N402, N328);
and AND3 (N432, N428, N340, N382);
or OR4 (N433, N406, N223, N390, N63);
and AND3 (N434, N407, N228, N398);
or OR2 (N435, N430, N338);
not NOT1 (N436, N431);
buf BUF1 (N437, N421);
nand NAND3 (N438, N436, N50, N3);
xor XOR2 (N439, N434, N423);
or OR3 (N440, N427, N207, N333);
or OR2 (N441, N433, N274);
not NOT1 (N442, N437);
nand NAND3 (N443, N435, N105, N432);
or OR4 (N444, N300, N153, N202, N35);
xor XOR2 (N445, N440, N27);
and AND2 (N446, N438, N168);
nor NOR4 (N447, N444, N83, N164, N99);
not NOT1 (N448, N439);
nand NAND2 (N449, N448, N305);
xor XOR2 (N450, N429, N330);
nor NOR4 (N451, N443, N400, N36, N315);
not NOT1 (N452, N441);
nand NAND4 (N453, N424, N40, N319, N293);
nor NOR2 (N454, N452, N320);
nor NOR4 (N455, N447, N211, N319, N422);
xor XOR2 (N456, N403, N16);
nor NOR2 (N457, N446, N345);
buf BUF1 (N458, N442);
buf BUF1 (N459, N451);
and AND3 (N460, N445, N330, N36);
nor NOR2 (N461, N457, N94);
nor NOR2 (N462, N458, N70);
and AND2 (N463, N461, N267);
nor NOR3 (N464, N455, N140, N330);
not NOT1 (N465, N462);
buf BUF1 (N466, N456);
or OR3 (N467, N459, N236, N86);
nand NAND4 (N468, N449, N3, N457, N322);
buf BUF1 (N469, N460);
xor XOR2 (N470, N465, N231);
nor NOR4 (N471, N467, N309, N117, N378);
and AND4 (N472, N453, N125, N164, N69);
buf BUF1 (N473, N450);
buf BUF1 (N474, N470);
xor XOR2 (N475, N468, N83);
nand NAND3 (N476, N472, N370, N464);
xor XOR2 (N477, N307, N219);
not NOT1 (N478, N463);
xor XOR2 (N479, N471, N350);
not NOT1 (N480, N477);
or OR4 (N481, N476, N166, N104, N427);
and AND4 (N482, N480, N410, N220, N243);
or OR4 (N483, N482, N305, N149, N243);
nand NAND2 (N484, N481, N366);
and AND3 (N485, N474, N150, N33);
buf BUF1 (N486, N469);
and AND4 (N487, N454, N38, N103, N282);
or OR4 (N488, N487, N412, N422, N313);
and AND4 (N489, N478, N375, N25, N435);
and AND3 (N490, N484, N485, N196);
nor NOR4 (N491, N408, N487, N368, N299);
buf BUF1 (N492, N486);
xor XOR2 (N493, N483, N238);
nor NOR4 (N494, N479, N361, N220, N41);
xor XOR2 (N495, N494, N52);
xor XOR2 (N496, N492, N133);
not NOT1 (N497, N493);
not NOT1 (N498, N490);
not NOT1 (N499, N496);
xor XOR2 (N500, N495, N384);
and AND3 (N501, N499, N156, N301);
or OR4 (N502, N497, N314, N208, N251);
buf BUF1 (N503, N473);
or OR2 (N504, N502, N166);
buf BUF1 (N505, N466);
xor XOR2 (N506, N503, N302);
not NOT1 (N507, N501);
buf BUF1 (N508, N491);
nor NOR4 (N509, N489, N492, N247, N401);
and AND3 (N510, N500, N69, N446);
nor NOR4 (N511, N507, N451, N406, N16);
nand NAND3 (N512, N510, N395, N383);
xor XOR2 (N513, N488, N52);
not NOT1 (N514, N505);
and AND3 (N515, N498, N391, N410);
or OR3 (N516, N508, N375, N181);
xor XOR2 (N517, N516, N453);
buf BUF1 (N518, N515);
nor NOR3 (N519, N511, N26, N135);
xor XOR2 (N520, N513, N212);
buf BUF1 (N521, N504);
nor NOR4 (N522, N512, N54, N191, N427);
nand NAND4 (N523, N518, N403, N517, N1);
xor XOR2 (N524, N237, N28);
buf BUF1 (N525, N520);
xor XOR2 (N526, N523, N104);
or OR2 (N527, N524, N398);
or OR4 (N528, N521, N328, N244, N73);
xor XOR2 (N529, N506, N291);
nand NAND2 (N530, N514, N270);
not NOT1 (N531, N528);
buf BUF1 (N532, N527);
nor NOR3 (N533, N531, N416, N106);
nand NAND2 (N534, N509, N445);
and AND4 (N535, N475, N433, N179, N208);
nor NOR2 (N536, N532, N89);
nand NAND4 (N537, N530, N381, N481, N93);
or OR2 (N538, N526, N529);
or OR4 (N539, N52, N123, N418, N33);
xor XOR2 (N540, N533, N121);
xor XOR2 (N541, N535, N405);
and AND2 (N542, N534, N93);
or OR2 (N543, N519, N172);
not NOT1 (N544, N541);
xor XOR2 (N545, N542, N416);
and AND2 (N546, N537, N516);
buf BUF1 (N547, N536);
not NOT1 (N548, N522);
nor NOR2 (N549, N547, N105);
nand NAND4 (N550, N525, N133, N344, N135);
not NOT1 (N551, N544);
not NOT1 (N552, N551);
nor NOR3 (N553, N548, N264, N305);
not NOT1 (N554, N553);
not NOT1 (N555, N552);
not NOT1 (N556, N540);
and AND2 (N557, N555, N56);
and AND2 (N558, N539, N89);
or OR4 (N559, N546, N530, N494, N444);
xor XOR2 (N560, N557, N348);
or OR4 (N561, N550, N510, N391, N42);
buf BUF1 (N562, N558);
buf BUF1 (N563, N556);
not NOT1 (N564, N538);
nand NAND2 (N565, N559, N563);
or OR3 (N566, N237, N109, N246);
nand NAND4 (N567, N565, N92, N96, N402);
nor NOR3 (N568, N554, N12, N186);
xor XOR2 (N569, N564, N544);
or OR3 (N570, N545, N263, N62);
not NOT1 (N571, N549);
nor NOR2 (N572, N569, N279);
or OR4 (N573, N566, N187, N36, N567);
nand NAND4 (N574, N420, N363, N73, N273);
xor XOR2 (N575, N573, N502);
or OR3 (N576, N560, N355, N450);
or OR4 (N577, N571, N153, N396, N62);
nor NOR3 (N578, N562, N559, N197);
nor NOR4 (N579, N577, N46, N282, N564);
buf BUF1 (N580, N543);
nand NAND2 (N581, N578, N340);
buf BUF1 (N582, N568);
and AND4 (N583, N576, N326, N313, N346);
and AND4 (N584, N575, N20, N235, N21);
and AND2 (N585, N580, N86);
buf BUF1 (N586, N583);
not NOT1 (N587, N579);
and AND4 (N588, N582, N357, N3, N579);
xor XOR2 (N589, N588, N294);
nor NOR4 (N590, N572, N316, N574, N195);
xor XOR2 (N591, N412, N147);
nor NOR4 (N592, N586, N388, N384, N49);
not NOT1 (N593, N591);
not NOT1 (N594, N581);
or OR2 (N595, N585, N138);
and AND4 (N596, N590, N382, N5, N159);
not NOT1 (N597, N596);
nand NAND2 (N598, N587, N161);
nand NAND4 (N599, N561, N265, N383, N103);
buf BUF1 (N600, N595);
nand NAND3 (N601, N599, N337, N309);
nand NAND4 (N602, N601, N231, N360, N463);
nand NAND3 (N603, N584, N14, N18);
buf BUF1 (N604, N592);
xor XOR2 (N605, N602, N275);
xor XOR2 (N606, N594, N79);
and AND2 (N607, N600, N81);
or OR3 (N608, N606, N3, N69);
not NOT1 (N609, N603);
xor XOR2 (N610, N608, N152);
xor XOR2 (N611, N604, N596);
xor XOR2 (N612, N598, N163);
and AND2 (N613, N612, N59);
nor NOR4 (N614, N611, N315, N475, N507);
and AND4 (N615, N570, N546, N389, N463);
nor NOR4 (N616, N613, N492, N425, N530);
nand NAND2 (N617, N615, N309);
nand NAND3 (N618, N614, N577, N586);
not NOT1 (N619, N609);
and AND3 (N620, N618, N73, N475);
and AND2 (N621, N607, N23);
buf BUF1 (N622, N617);
not NOT1 (N623, N621);
buf BUF1 (N624, N619);
and AND3 (N625, N605, N68, N353);
xor XOR2 (N626, N625, N569);
buf BUF1 (N627, N624);
buf BUF1 (N628, N610);
buf BUF1 (N629, N627);
nand NAND4 (N630, N626, N211, N171, N262);
not NOT1 (N631, N620);
not NOT1 (N632, N623);
not NOT1 (N633, N616);
nor NOR3 (N634, N631, N286, N276);
or OR3 (N635, N633, N191, N68);
nand NAND2 (N636, N589, N442);
xor XOR2 (N637, N628, N107);
not NOT1 (N638, N629);
or OR3 (N639, N597, N598, N35);
and AND4 (N640, N622, N349, N424, N259);
nand NAND2 (N641, N634, N224);
buf BUF1 (N642, N641);
and AND4 (N643, N632, N355, N126, N419);
xor XOR2 (N644, N637, N175);
buf BUF1 (N645, N630);
xor XOR2 (N646, N640, N401);
buf BUF1 (N647, N642);
xor XOR2 (N648, N635, N157);
nand NAND3 (N649, N639, N613, N93);
or OR2 (N650, N649, N244);
nor NOR2 (N651, N648, N315);
not NOT1 (N652, N647);
and AND3 (N653, N643, N51, N548);
xor XOR2 (N654, N651, N40);
buf BUF1 (N655, N644);
or OR4 (N656, N645, N34, N638, N320);
buf BUF1 (N657, N160);
nor NOR4 (N658, N652, N613, N193, N461);
and AND3 (N659, N646, N218, N283);
or OR4 (N660, N654, N425, N93, N32);
xor XOR2 (N661, N593, N291);
xor XOR2 (N662, N661, N154);
not NOT1 (N663, N636);
xor XOR2 (N664, N659, N132);
not NOT1 (N665, N656);
buf BUF1 (N666, N660);
not NOT1 (N667, N664);
not NOT1 (N668, N653);
xor XOR2 (N669, N666, N140);
nor NOR4 (N670, N667, N26, N11, N40);
or OR4 (N671, N655, N523, N308, N289);
and AND2 (N672, N658, N292);
buf BUF1 (N673, N671);
and AND2 (N674, N670, N280);
or OR2 (N675, N657, N571);
nand NAND3 (N676, N662, N302, N613);
and AND4 (N677, N650, N313, N8, N473);
xor XOR2 (N678, N669, N271);
and AND4 (N679, N678, N623, N606, N10);
not NOT1 (N680, N672);
or OR2 (N681, N676, N606);
nor NOR2 (N682, N681, N671);
nand NAND4 (N683, N665, N306, N252, N64);
or OR3 (N684, N677, N630, N152);
nor NOR2 (N685, N675, N532);
nor NOR4 (N686, N683, N645, N412, N292);
xor XOR2 (N687, N685, N594);
buf BUF1 (N688, N668);
or OR2 (N689, N663, N72);
not NOT1 (N690, N673);
buf BUF1 (N691, N679);
not NOT1 (N692, N684);
xor XOR2 (N693, N688, N323);
not NOT1 (N694, N690);
buf BUF1 (N695, N686);
nand NAND2 (N696, N680, N452);
nand NAND2 (N697, N689, N236);
nor NOR2 (N698, N682, N402);
buf BUF1 (N699, N696);
or OR2 (N700, N695, N162);
and AND4 (N701, N691, N659, N437, N84);
and AND4 (N702, N687, N502, N296, N375);
buf BUF1 (N703, N698);
or OR2 (N704, N702, N381);
nand NAND2 (N705, N704, N171);
and AND3 (N706, N700, N233, N34);
not NOT1 (N707, N674);
nand NAND2 (N708, N701, N18);
not NOT1 (N709, N706);
buf BUF1 (N710, N697);
or OR4 (N711, N709, N27, N568, N603);
and AND4 (N712, N692, N181, N446, N317);
buf BUF1 (N713, N708);
nor NOR4 (N714, N707, N411, N604, N408);
not NOT1 (N715, N710);
nand NAND4 (N716, N703, N526, N75, N650);
nand NAND3 (N717, N693, N611, N598);
and AND2 (N718, N714, N377);
xor XOR2 (N719, N718, N315);
xor XOR2 (N720, N705, N636);
buf BUF1 (N721, N717);
xor XOR2 (N722, N720, N52);
nor NOR4 (N723, N721, N79, N547, N41);
and AND4 (N724, N722, N71, N156, N228);
buf BUF1 (N725, N716);
nor NOR3 (N726, N724, N469, N499);
xor XOR2 (N727, N713, N519);
or OR2 (N728, N727, N717);
and AND2 (N729, N728, N319);
xor XOR2 (N730, N719, N165);
buf BUF1 (N731, N715);
nand NAND3 (N732, N711, N109, N449);
or OR2 (N733, N732, N21);
xor XOR2 (N734, N726, N141);
and AND4 (N735, N730, N308, N419, N617);
nand NAND4 (N736, N723, N219, N242, N523);
not NOT1 (N737, N734);
nand NAND4 (N738, N725, N686, N685, N670);
nor NOR4 (N739, N733, N296, N523, N400);
and AND3 (N740, N731, N738, N693);
nor NOR4 (N741, N445, N490, N474, N445);
and AND3 (N742, N740, N524, N407);
or OR2 (N743, N694, N659);
buf BUF1 (N744, N699);
or OR3 (N745, N744, N59, N726);
and AND3 (N746, N739, N720, N316);
and AND3 (N747, N742, N218, N25);
xor XOR2 (N748, N735, N492);
nor NOR3 (N749, N736, N477, N59);
and AND2 (N750, N712, N705);
buf BUF1 (N751, N737);
nand NAND4 (N752, N749, N647, N563, N225);
nor NOR2 (N753, N748, N543);
and AND3 (N754, N745, N180, N40);
nor NOR2 (N755, N746, N13);
and AND3 (N756, N743, N565, N354);
xor XOR2 (N757, N747, N630);
or OR3 (N758, N756, N256, N583);
not NOT1 (N759, N751);
not NOT1 (N760, N752);
xor XOR2 (N761, N757, N639);
xor XOR2 (N762, N761, N486);
or OR3 (N763, N762, N366, N433);
nor NOR3 (N764, N754, N564, N197);
xor XOR2 (N765, N741, N580);
and AND3 (N766, N765, N140, N220);
buf BUF1 (N767, N755);
not NOT1 (N768, N767);
and AND2 (N769, N750, N33);
nand NAND2 (N770, N766, N276);
and AND2 (N771, N764, N695);
nand NAND3 (N772, N771, N723, N209);
or OR2 (N773, N772, N514);
buf BUF1 (N774, N769);
not NOT1 (N775, N768);
nor NOR4 (N776, N759, N253, N171, N419);
xor XOR2 (N777, N763, N500);
buf BUF1 (N778, N773);
xor XOR2 (N779, N776, N79);
or OR3 (N780, N774, N33, N21);
not NOT1 (N781, N779);
not NOT1 (N782, N758);
or OR4 (N783, N782, N47, N9, N701);
not NOT1 (N784, N753);
or OR3 (N785, N784, N154, N74);
or OR3 (N786, N780, N729, N74);
not NOT1 (N787, N381);
xor XOR2 (N788, N785, N583);
nand NAND3 (N789, N781, N479, N334);
nor NOR2 (N790, N786, N394);
nand NAND4 (N791, N790, N78, N760, N3);
xor XOR2 (N792, N295, N528);
and AND3 (N793, N788, N760, N418);
and AND2 (N794, N775, N300);
nand NAND4 (N795, N787, N92, N442, N304);
nand NAND2 (N796, N789, N501);
xor XOR2 (N797, N796, N765);
buf BUF1 (N798, N778);
nand NAND2 (N799, N797, N571);
xor XOR2 (N800, N783, N438);
and AND2 (N801, N777, N665);
xor XOR2 (N802, N800, N703);
or OR2 (N803, N770, N74);
not NOT1 (N804, N803);
and AND2 (N805, N801, N294);
nand NAND3 (N806, N792, N469, N280);
xor XOR2 (N807, N806, N151);
or OR3 (N808, N795, N705, N377);
nor NOR3 (N809, N805, N247, N33);
and AND4 (N810, N799, N46, N445, N312);
not NOT1 (N811, N804);
buf BUF1 (N812, N791);
or OR4 (N813, N798, N303, N507, N385);
buf BUF1 (N814, N811);
buf BUF1 (N815, N802);
and AND4 (N816, N813, N41, N536, N372);
xor XOR2 (N817, N810, N648);
nor NOR4 (N818, N809, N333, N631, N146);
buf BUF1 (N819, N816);
xor XOR2 (N820, N812, N628);
buf BUF1 (N821, N820);
and AND2 (N822, N793, N702);
not NOT1 (N823, N819);
nor NOR4 (N824, N817, N660, N604, N573);
nand NAND4 (N825, N814, N563, N21, N35);
nand NAND4 (N826, N821, N708, N85, N453);
xor XOR2 (N827, N825, N6);
nor NOR3 (N828, N815, N503, N513);
and AND4 (N829, N823, N153, N593, N6);
not NOT1 (N830, N794);
and AND4 (N831, N829, N244, N613, N419);
and AND4 (N832, N827, N738, N640, N122);
not NOT1 (N833, N830);
xor XOR2 (N834, N828, N785);
buf BUF1 (N835, N818);
nor NOR2 (N836, N807, N291);
nand NAND2 (N837, N834, N522);
nand NAND2 (N838, N835, N290);
nand NAND3 (N839, N831, N809, N551);
xor XOR2 (N840, N822, N31);
or OR2 (N841, N839, N431);
not NOT1 (N842, N841);
not NOT1 (N843, N832);
nand NAND2 (N844, N840, N211);
nor NOR2 (N845, N833, N702);
not NOT1 (N846, N838);
and AND3 (N847, N837, N110, N118);
nand NAND2 (N848, N843, N473);
xor XOR2 (N849, N808, N724);
buf BUF1 (N850, N826);
and AND4 (N851, N824, N820, N801, N252);
or OR3 (N852, N851, N503, N541);
nand NAND3 (N853, N842, N795, N144);
or OR2 (N854, N848, N359);
xor XOR2 (N855, N852, N588);
buf BUF1 (N856, N836);
xor XOR2 (N857, N856, N206);
or OR2 (N858, N854, N477);
and AND3 (N859, N858, N219, N221);
or OR3 (N860, N846, N272, N362);
nand NAND2 (N861, N855, N129);
and AND3 (N862, N847, N245, N477);
xor XOR2 (N863, N861, N343);
nand NAND4 (N864, N850, N784, N66, N293);
buf BUF1 (N865, N863);
buf BUF1 (N866, N844);
nand NAND4 (N867, N857, N657, N298, N68);
and AND4 (N868, N862, N138, N465, N403);
and AND2 (N869, N867, N165);
or OR2 (N870, N860, N841);
or OR3 (N871, N869, N494, N675);
buf BUF1 (N872, N859);
xor XOR2 (N873, N872, N736);
nor NOR4 (N874, N871, N665, N324, N35);
not NOT1 (N875, N864);
nand NAND4 (N876, N849, N256, N615, N161);
buf BUF1 (N877, N845);
and AND3 (N878, N875, N208, N830);
buf BUF1 (N879, N868);
and AND3 (N880, N873, N192, N131);
nor NOR3 (N881, N877, N337, N702);
buf BUF1 (N882, N880);
or OR3 (N883, N882, N666, N30);
or OR2 (N884, N874, N583);
xor XOR2 (N885, N870, N435);
not NOT1 (N886, N866);
nand NAND4 (N887, N876, N3, N53, N656);
or OR2 (N888, N853, N721);
xor XOR2 (N889, N888, N138);
and AND4 (N890, N883, N594, N720, N857);
nand NAND2 (N891, N885, N475);
or OR4 (N892, N878, N821, N211, N51);
buf BUF1 (N893, N865);
or OR4 (N894, N884, N563, N430, N719);
nor NOR4 (N895, N893, N866, N702, N487);
and AND2 (N896, N891, N153);
xor XOR2 (N897, N889, N523);
and AND4 (N898, N886, N105, N684, N122);
not NOT1 (N899, N892);
not NOT1 (N900, N881);
nand NAND3 (N901, N879, N145, N149);
nand NAND3 (N902, N896, N155, N206);
buf BUF1 (N903, N887);
buf BUF1 (N904, N895);
or OR4 (N905, N900, N95, N836, N568);
and AND3 (N906, N901, N230, N391);
buf BUF1 (N907, N902);
not NOT1 (N908, N894);
not NOT1 (N909, N904);
or OR2 (N910, N908, N514);
xor XOR2 (N911, N899, N887);
xor XOR2 (N912, N909, N392);
xor XOR2 (N913, N907, N551);
buf BUF1 (N914, N911);
and AND3 (N915, N898, N46, N157);
nand NAND2 (N916, N914, N175);
or OR4 (N917, N915, N372, N48, N247);
nor NOR3 (N918, N890, N102, N467);
nand NAND4 (N919, N918, N589, N312, N884);
buf BUF1 (N920, N903);
or OR4 (N921, N906, N579, N456, N795);
and AND3 (N922, N912, N412, N498);
nand NAND2 (N923, N913, N386);
not NOT1 (N924, N905);
nor NOR2 (N925, N919, N659);
not NOT1 (N926, N920);
or OR4 (N927, N916, N598, N895, N431);
and AND3 (N928, N924, N520, N901);
nand NAND3 (N929, N923, N116, N413);
or OR3 (N930, N922, N134, N389);
or OR3 (N931, N910, N23, N407);
xor XOR2 (N932, N897, N567);
nor NOR3 (N933, N921, N466, N354);
buf BUF1 (N934, N929);
buf BUF1 (N935, N925);
nor NOR4 (N936, N932, N687, N123, N471);
not NOT1 (N937, N933);
xor XOR2 (N938, N931, N744);
nor NOR2 (N939, N927, N798);
nor NOR4 (N940, N928, N448, N770, N753);
xor XOR2 (N941, N940, N288);
buf BUF1 (N942, N938);
nor NOR4 (N943, N937, N386, N781, N798);
not NOT1 (N944, N943);
or OR4 (N945, N934, N603, N497, N868);
and AND4 (N946, N936, N47, N619, N66);
not NOT1 (N947, N917);
nor NOR2 (N948, N947, N649);
or OR4 (N949, N942, N586, N7, N702);
xor XOR2 (N950, N944, N594);
nor NOR2 (N951, N926, N257);
xor XOR2 (N952, N945, N898);
not NOT1 (N953, N950);
xor XOR2 (N954, N952, N486);
nor NOR2 (N955, N948, N267);
xor XOR2 (N956, N949, N781);
and AND4 (N957, N951, N576, N896, N178);
buf BUF1 (N958, N946);
or OR2 (N959, N935, N764);
xor XOR2 (N960, N957, N761);
nand NAND4 (N961, N956, N196, N384, N738);
or OR4 (N962, N960, N508, N657, N255);
not NOT1 (N963, N962);
nor NOR3 (N964, N961, N388, N637);
and AND2 (N965, N964, N278);
buf BUF1 (N966, N958);
not NOT1 (N967, N954);
not NOT1 (N968, N966);
nand NAND2 (N969, N930, N547);
not NOT1 (N970, N941);
not NOT1 (N971, N967);
not NOT1 (N972, N968);
buf BUF1 (N973, N969);
nor NOR4 (N974, N955, N499, N653, N175);
and AND3 (N975, N973, N216, N865);
buf BUF1 (N976, N971);
and AND3 (N977, N953, N286, N526);
nand NAND2 (N978, N972, N956);
or OR4 (N979, N978, N819, N876, N303);
and AND4 (N980, N975, N786, N233, N529);
xor XOR2 (N981, N939, N605);
nand NAND4 (N982, N965, N133, N65, N725);
xor XOR2 (N983, N976, N814);
nand NAND3 (N984, N981, N416, N63);
not NOT1 (N985, N959);
not NOT1 (N986, N985);
and AND3 (N987, N983, N259, N205);
not NOT1 (N988, N974);
or OR2 (N989, N984, N124);
not NOT1 (N990, N988);
xor XOR2 (N991, N970, N898);
not NOT1 (N992, N982);
nand NAND2 (N993, N980, N210);
nor NOR4 (N994, N990, N960, N456, N631);
not NOT1 (N995, N963);
nor NOR4 (N996, N979, N225, N832, N551);
xor XOR2 (N997, N992, N25);
xor XOR2 (N998, N995, N654);
and AND3 (N999, N989, N746, N37);
nor NOR4 (N1000, N994, N928, N565, N355);
nor NOR2 (N1001, N998, N517);
nor NOR2 (N1002, N997, N277);
xor XOR2 (N1003, N977, N347);
xor XOR2 (N1004, N996, N316);
or OR3 (N1005, N1004, N362, N933);
or OR2 (N1006, N993, N159);
not NOT1 (N1007, N986);
not NOT1 (N1008, N987);
and AND2 (N1009, N1002, N166);
nor NOR4 (N1010, N991, N850, N964, N424);
and AND4 (N1011, N1008, N581, N841, N864);
not NOT1 (N1012, N1001);
or OR4 (N1013, N1009, N14, N374, N430);
nor NOR3 (N1014, N999, N206, N453);
and AND3 (N1015, N1010, N792, N975);
not NOT1 (N1016, N1006);
nand NAND4 (N1017, N1011, N547, N291, N925);
nand NAND3 (N1018, N1003, N976, N139);
xor XOR2 (N1019, N1012, N418);
nand NAND3 (N1020, N1019, N278, N815);
nor NOR4 (N1021, N1007, N574, N36, N93);
nor NOR2 (N1022, N1016, N263);
xor XOR2 (N1023, N1020, N224);
or OR4 (N1024, N1021, N773, N464, N1003);
not NOT1 (N1025, N1000);
or OR3 (N1026, N1017, N782, N738);
nand NAND2 (N1027, N1023, N533);
and AND2 (N1028, N1015, N669);
nand NAND4 (N1029, N1014, N828, N193, N611);
and AND3 (N1030, N1013, N59, N222);
nor NOR2 (N1031, N1028, N154);
nor NOR2 (N1032, N1022, N716);
or OR4 (N1033, N1032, N18, N370, N793);
not NOT1 (N1034, N1029);
or OR2 (N1035, N1005, N1032);
not NOT1 (N1036, N1033);
buf BUF1 (N1037, N1027);
buf BUF1 (N1038, N1024);
not NOT1 (N1039, N1025);
or OR2 (N1040, N1030, N5);
nor NOR2 (N1041, N1035, N534);
nand NAND3 (N1042, N1031, N744, N822);
or OR2 (N1043, N1026, N778);
nor NOR4 (N1044, N1034, N42, N824, N96);
or OR4 (N1045, N1038, N928, N199, N1010);
xor XOR2 (N1046, N1043, N6);
or OR2 (N1047, N1046, N370);
not NOT1 (N1048, N1037);
xor XOR2 (N1049, N1042, N1034);
not NOT1 (N1050, N1039);
and AND4 (N1051, N1050, N787, N398, N55);
or OR4 (N1052, N1018, N128, N848, N274);
nor NOR2 (N1053, N1045, N1023);
and AND4 (N1054, N1049, N164, N419, N589);
nand NAND2 (N1055, N1047, N702);
and AND4 (N1056, N1053, N434, N102, N935);
buf BUF1 (N1057, N1052);
nor NOR3 (N1058, N1055, N678, N195);
buf BUF1 (N1059, N1036);
nand NAND2 (N1060, N1057, N46);
and AND3 (N1061, N1054, N794, N100);
not NOT1 (N1062, N1041);
buf BUF1 (N1063, N1060);
buf BUF1 (N1064, N1059);
not NOT1 (N1065, N1056);
and AND4 (N1066, N1063, N781, N183, N747);
or OR4 (N1067, N1051, N349, N994, N660);
or OR2 (N1068, N1065, N1047);
xor XOR2 (N1069, N1067, N1060);
nor NOR4 (N1070, N1044, N487, N381, N750);
nand NAND2 (N1071, N1061, N270);
xor XOR2 (N1072, N1070, N910);
buf BUF1 (N1073, N1068);
nand NAND4 (N1074, N1073, N1061, N764, N16);
or OR4 (N1075, N1062, N461, N299, N941);
or OR3 (N1076, N1040, N877, N205);
or OR3 (N1077, N1069, N501, N225);
or OR2 (N1078, N1074, N620);
buf BUF1 (N1079, N1071);
xor XOR2 (N1080, N1075, N936);
and AND3 (N1081, N1076, N108, N822);
not NOT1 (N1082, N1079);
and AND4 (N1083, N1082, N411, N325, N619);
and AND3 (N1084, N1080, N674, N109);
xor XOR2 (N1085, N1066, N1017);
nor NOR2 (N1086, N1084, N1006);
nand NAND4 (N1087, N1085, N876, N977, N640);
or OR3 (N1088, N1081, N646, N718);
and AND2 (N1089, N1077, N450);
nand NAND2 (N1090, N1058, N277);
buf BUF1 (N1091, N1088);
nor NOR3 (N1092, N1083, N772, N936);
not NOT1 (N1093, N1048);
not NOT1 (N1094, N1086);
or OR3 (N1095, N1078, N274, N487);
xor XOR2 (N1096, N1092, N73);
buf BUF1 (N1097, N1095);
and AND4 (N1098, N1093, N331, N342, N237);
nand NAND4 (N1099, N1072, N869, N138, N98);
not NOT1 (N1100, N1091);
nor NOR3 (N1101, N1090, N1044, N854);
nand NAND4 (N1102, N1097, N528, N303, N213);
or OR2 (N1103, N1099, N360);
not NOT1 (N1104, N1089);
or OR4 (N1105, N1101, N911, N396, N283);
xor XOR2 (N1106, N1094, N376);
nand NAND4 (N1107, N1087, N451, N269, N915);
xor XOR2 (N1108, N1103, N157);
nand NAND2 (N1109, N1098, N175);
or OR2 (N1110, N1109, N607);
buf BUF1 (N1111, N1105);
or OR3 (N1112, N1111, N217, N844);
and AND3 (N1113, N1064, N414, N960);
and AND3 (N1114, N1096, N994, N369);
not NOT1 (N1115, N1114);
buf BUF1 (N1116, N1106);
nand NAND4 (N1117, N1102, N675, N789, N1097);
and AND3 (N1118, N1100, N916, N440);
buf BUF1 (N1119, N1116);
not NOT1 (N1120, N1115);
nor NOR3 (N1121, N1108, N235, N559);
or OR3 (N1122, N1104, N795, N457);
xor XOR2 (N1123, N1119, N729);
and AND2 (N1124, N1122, N511);
or OR3 (N1125, N1120, N334, N106);
nand NAND2 (N1126, N1113, N962);
buf BUF1 (N1127, N1118);
not NOT1 (N1128, N1127);
xor XOR2 (N1129, N1112, N422);
or OR2 (N1130, N1107, N916);
buf BUF1 (N1131, N1121);
and AND4 (N1132, N1126, N378, N625, N813);
or OR3 (N1133, N1129, N746, N245);
or OR3 (N1134, N1110, N593, N215);
or OR3 (N1135, N1123, N984, N212);
nor NOR3 (N1136, N1125, N305, N451);
nand NAND4 (N1137, N1132, N922, N114, N392);
xor XOR2 (N1138, N1130, N855);
nand NAND3 (N1139, N1117, N258, N661);
nand NAND4 (N1140, N1134, N796, N1021, N951);
and AND3 (N1141, N1124, N804, N242);
not NOT1 (N1142, N1136);
nand NAND2 (N1143, N1141, N1067);
or OR3 (N1144, N1128, N1025, N419);
nor NOR4 (N1145, N1138, N1076, N739, N1107);
nand NAND3 (N1146, N1139, N68, N90);
or OR2 (N1147, N1146, N790);
buf BUF1 (N1148, N1133);
not NOT1 (N1149, N1148);
not NOT1 (N1150, N1149);
nand NAND4 (N1151, N1150, N964, N416, N809);
nor NOR4 (N1152, N1144, N179, N663, N157);
buf BUF1 (N1153, N1135);
not NOT1 (N1154, N1147);
and AND4 (N1155, N1140, N44, N1023, N172);
nand NAND2 (N1156, N1131, N32);
nor NOR3 (N1157, N1152, N618, N369);
not NOT1 (N1158, N1157);
and AND4 (N1159, N1145, N946, N290, N687);
nand NAND3 (N1160, N1159, N801, N53);
buf BUF1 (N1161, N1151);
and AND2 (N1162, N1160, N487);
and AND3 (N1163, N1156, N266, N990);
xor XOR2 (N1164, N1153, N742);
and AND3 (N1165, N1142, N735, N717);
not NOT1 (N1166, N1158);
nor NOR3 (N1167, N1154, N225, N935);
buf BUF1 (N1168, N1155);
nor NOR3 (N1169, N1161, N371, N300);
buf BUF1 (N1170, N1168);
nor NOR2 (N1171, N1169, N847);
buf BUF1 (N1172, N1170);
nor NOR2 (N1173, N1167, N220);
xor XOR2 (N1174, N1137, N86);
or OR4 (N1175, N1166, N488, N147, N961);
xor XOR2 (N1176, N1174, N559);
nor NOR4 (N1177, N1143, N198, N899, N149);
not NOT1 (N1178, N1164);
nand NAND2 (N1179, N1162, N107);
buf BUF1 (N1180, N1171);
or OR3 (N1181, N1165, N785, N726);
nor NOR4 (N1182, N1181, N57, N513, N723);
or OR2 (N1183, N1180, N319);
not NOT1 (N1184, N1178);
or OR2 (N1185, N1163, N638);
nand NAND2 (N1186, N1182, N488);
nand NAND4 (N1187, N1184, N534, N253, N933);
and AND3 (N1188, N1175, N366, N51);
and AND4 (N1189, N1185, N295, N371, N1158);
nand NAND3 (N1190, N1172, N726, N886);
or OR4 (N1191, N1173, N867, N818, N1130);
nand NAND4 (N1192, N1176, N764, N222, N1104);
nand NAND2 (N1193, N1192, N211);
xor XOR2 (N1194, N1193, N403);
not NOT1 (N1195, N1183);
xor XOR2 (N1196, N1187, N1066);
not NOT1 (N1197, N1186);
nor NOR3 (N1198, N1177, N472, N1045);
xor XOR2 (N1199, N1179, N1034);
buf BUF1 (N1200, N1199);
buf BUF1 (N1201, N1195);
buf BUF1 (N1202, N1197);
not NOT1 (N1203, N1200);
xor XOR2 (N1204, N1190, N722);
not NOT1 (N1205, N1196);
buf BUF1 (N1206, N1194);
nor NOR2 (N1207, N1204, N519);
nor NOR3 (N1208, N1191, N82, N137);
nor NOR3 (N1209, N1205, N693, N838);
xor XOR2 (N1210, N1206, N103);
and AND3 (N1211, N1207, N965, N164);
nand NAND2 (N1212, N1209, N82);
or OR4 (N1213, N1201, N666, N214, N277);
nand NAND4 (N1214, N1203, N181, N726, N1029);
not NOT1 (N1215, N1208);
not NOT1 (N1216, N1188);
nand NAND2 (N1217, N1189, N556);
nor NOR3 (N1218, N1212, N1116, N365);
nand NAND4 (N1219, N1198, N874, N55, N121);
nand NAND2 (N1220, N1202, N1058);
xor XOR2 (N1221, N1220, N420);
nand NAND2 (N1222, N1211, N950);
nor NOR4 (N1223, N1219, N347, N94, N573);
nor NOR2 (N1224, N1213, N1209);
or OR4 (N1225, N1210, N340, N68, N815);
xor XOR2 (N1226, N1216, N119);
nand NAND2 (N1227, N1221, N810);
buf BUF1 (N1228, N1226);
xor XOR2 (N1229, N1222, N402);
and AND2 (N1230, N1217, N1015);
or OR2 (N1231, N1229, N922);
and AND3 (N1232, N1224, N330, N938);
buf BUF1 (N1233, N1232);
nor NOR3 (N1234, N1218, N570, N336);
buf BUF1 (N1235, N1231);
nand NAND2 (N1236, N1215, N845);
nand NAND3 (N1237, N1235, N950, N419);
or OR3 (N1238, N1223, N1092, N1033);
or OR2 (N1239, N1230, N447);
nand NAND2 (N1240, N1228, N1091);
or OR3 (N1241, N1233, N561, N410);
xor XOR2 (N1242, N1237, N646);
not NOT1 (N1243, N1214);
and AND2 (N1244, N1242, N1090);
not NOT1 (N1245, N1241);
buf BUF1 (N1246, N1238);
not NOT1 (N1247, N1240);
or OR3 (N1248, N1239, N314, N1072);
nor NOR3 (N1249, N1236, N125, N873);
or OR4 (N1250, N1243, N1177, N103, N219);
not NOT1 (N1251, N1225);
or OR2 (N1252, N1251, N1238);
xor XOR2 (N1253, N1248, N313);
not NOT1 (N1254, N1253);
buf BUF1 (N1255, N1227);
not NOT1 (N1256, N1245);
and AND3 (N1257, N1244, N914, N432);
buf BUF1 (N1258, N1249);
not NOT1 (N1259, N1256);
or OR4 (N1260, N1234, N1094, N1224, N766);
nand NAND3 (N1261, N1258, N813, N218);
nand NAND2 (N1262, N1261, N436);
not NOT1 (N1263, N1262);
nor NOR4 (N1264, N1255, N622, N1223, N408);
or OR4 (N1265, N1263, N96, N276, N1094);
nor NOR4 (N1266, N1260, N1250, N1154, N803);
buf BUF1 (N1267, N658);
and AND2 (N1268, N1246, N1061);
buf BUF1 (N1269, N1259);
nor NOR3 (N1270, N1268, N1253, N920);
xor XOR2 (N1271, N1264, N179);
nor NOR4 (N1272, N1252, N1018, N792, N924);
and AND2 (N1273, N1270, N1154);
buf BUF1 (N1274, N1254);
nand NAND4 (N1275, N1266, N1137, N250, N1181);
not NOT1 (N1276, N1257);
xor XOR2 (N1277, N1247, N164);
nand NAND2 (N1278, N1269, N510);
and AND4 (N1279, N1277, N1170, N146, N32);
nor NOR3 (N1280, N1267, N794, N510);
nor NOR4 (N1281, N1275, N769, N1038, N960);
nor NOR2 (N1282, N1278, N596);
nor NOR3 (N1283, N1273, N339, N1073);
xor XOR2 (N1284, N1274, N185);
buf BUF1 (N1285, N1271);
buf BUF1 (N1286, N1265);
nand NAND4 (N1287, N1284, N818, N333, N184);
buf BUF1 (N1288, N1286);
not NOT1 (N1289, N1279);
and AND3 (N1290, N1283, N819, N62);
or OR4 (N1291, N1280, N1091, N116, N989);
or OR4 (N1292, N1287, N984, N1248, N1143);
buf BUF1 (N1293, N1291);
not NOT1 (N1294, N1293);
or OR4 (N1295, N1288, N489, N1224, N140);
and AND2 (N1296, N1272, N497);
buf BUF1 (N1297, N1292);
nand NAND2 (N1298, N1295, N949);
not NOT1 (N1299, N1276);
xor XOR2 (N1300, N1294, N859);
buf BUF1 (N1301, N1300);
and AND2 (N1302, N1281, N541);
or OR3 (N1303, N1299, N1107, N598);
not NOT1 (N1304, N1297);
and AND3 (N1305, N1303, N419, N107);
nand NAND4 (N1306, N1304, N879, N709, N1280);
nor NOR4 (N1307, N1296, N160, N514, N412);
nor NOR3 (N1308, N1290, N122, N1127);
xor XOR2 (N1309, N1306, N735);
and AND3 (N1310, N1307, N599, N535);
not NOT1 (N1311, N1282);
and AND3 (N1312, N1302, N1207, N910);
or OR2 (N1313, N1311, N161);
xor XOR2 (N1314, N1301, N504);
or OR4 (N1315, N1310, N489, N1021, N326);
nor NOR3 (N1316, N1313, N163, N655);
nor NOR3 (N1317, N1305, N285, N1025);
nand NAND4 (N1318, N1316, N469, N1084, N503);
nand NAND4 (N1319, N1289, N1122, N358, N331);
nand NAND2 (N1320, N1319, N267);
buf BUF1 (N1321, N1318);
and AND4 (N1322, N1315, N9, N1252, N321);
nand NAND2 (N1323, N1314, N168);
and AND2 (N1324, N1308, N309);
buf BUF1 (N1325, N1320);
and AND2 (N1326, N1317, N989);
nand NAND3 (N1327, N1326, N441, N832);
xor XOR2 (N1328, N1322, N1153);
or OR2 (N1329, N1325, N106);
nand NAND2 (N1330, N1312, N1273);
nor NOR4 (N1331, N1328, N1200, N671, N574);
nand NAND4 (N1332, N1298, N431, N1035, N391);
and AND3 (N1333, N1285, N659, N60);
not NOT1 (N1334, N1321);
xor XOR2 (N1335, N1330, N472);
not NOT1 (N1336, N1335);
nand NAND3 (N1337, N1323, N117, N936);
buf BUF1 (N1338, N1337);
not NOT1 (N1339, N1334);
not NOT1 (N1340, N1324);
and AND2 (N1341, N1340, N424);
not NOT1 (N1342, N1309);
not NOT1 (N1343, N1336);
buf BUF1 (N1344, N1331);
nor NOR4 (N1345, N1339, N1125, N1256, N1125);
not NOT1 (N1346, N1327);
nor NOR3 (N1347, N1345, N441, N472);
not NOT1 (N1348, N1338);
nor NOR4 (N1349, N1342, N602, N668, N1076);
or OR3 (N1350, N1347, N319, N730);
buf BUF1 (N1351, N1329);
or OR2 (N1352, N1349, N617);
nor NOR2 (N1353, N1341, N1027);
or OR3 (N1354, N1332, N995, N1293);
xor XOR2 (N1355, N1352, N770);
xor XOR2 (N1356, N1351, N1167);
nand NAND3 (N1357, N1353, N194, N1282);
not NOT1 (N1358, N1357);
or OR3 (N1359, N1343, N466, N815);
nor NOR2 (N1360, N1356, N132);
or OR4 (N1361, N1355, N1186, N254, N523);
nand NAND4 (N1362, N1361, N1004, N639, N356);
not NOT1 (N1363, N1360);
nor NOR3 (N1364, N1348, N844, N381);
or OR3 (N1365, N1344, N706, N836);
buf BUF1 (N1366, N1350);
and AND3 (N1367, N1354, N965, N1292);
buf BUF1 (N1368, N1365);
xor XOR2 (N1369, N1362, N4);
nor NOR3 (N1370, N1346, N516, N303);
nor NOR3 (N1371, N1363, N447, N913);
nand NAND3 (N1372, N1367, N842, N435);
xor XOR2 (N1373, N1369, N274);
xor XOR2 (N1374, N1359, N310);
nor NOR4 (N1375, N1373, N1323, N30, N218);
not NOT1 (N1376, N1375);
or OR3 (N1377, N1368, N1311, N688);
nand NAND2 (N1378, N1374, N1162);
buf BUF1 (N1379, N1333);
or OR2 (N1380, N1358, N209);
xor XOR2 (N1381, N1377, N893);
not NOT1 (N1382, N1366);
nand NAND3 (N1383, N1370, N913, N792);
nand NAND2 (N1384, N1364, N968);
and AND2 (N1385, N1371, N1159);
and AND4 (N1386, N1381, N580, N404, N1253);
nor NOR2 (N1387, N1379, N341);
and AND3 (N1388, N1378, N221, N1318);
and AND2 (N1389, N1386, N514);
or OR3 (N1390, N1383, N656, N602);
nor NOR2 (N1391, N1380, N1115);
or OR2 (N1392, N1385, N1148);
xor XOR2 (N1393, N1388, N535);
nor NOR3 (N1394, N1392, N1252, N95);
and AND4 (N1395, N1394, N1365, N1339, N601);
not NOT1 (N1396, N1395);
not NOT1 (N1397, N1382);
and AND3 (N1398, N1390, N286, N947);
nor NOR4 (N1399, N1397, N410, N1227, N635);
and AND4 (N1400, N1399, N451, N636, N996);
nor NOR2 (N1401, N1391, N1083);
or OR2 (N1402, N1389, N922);
not NOT1 (N1403, N1400);
xor XOR2 (N1404, N1387, N122);
xor XOR2 (N1405, N1372, N44);
not NOT1 (N1406, N1376);
and AND4 (N1407, N1402, N711, N467, N289);
xor XOR2 (N1408, N1384, N319);
nor NOR2 (N1409, N1403, N272);
xor XOR2 (N1410, N1406, N163);
not NOT1 (N1411, N1401);
nand NAND3 (N1412, N1411, N532, N870);
or OR4 (N1413, N1412, N591, N460, N1121);
buf BUF1 (N1414, N1404);
not NOT1 (N1415, N1408);
or OR2 (N1416, N1407, N14);
xor XOR2 (N1417, N1416, N1334);
or OR2 (N1418, N1415, N1212);
or OR4 (N1419, N1413, N1006, N772, N1246);
or OR3 (N1420, N1405, N344, N91);
xor XOR2 (N1421, N1393, N87);
buf BUF1 (N1422, N1414);
nor NOR2 (N1423, N1421, N1303);
buf BUF1 (N1424, N1417);
nor NOR2 (N1425, N1420, N118);
buf BUF1 (N1426, N1419);
xor XOR2 (N1427, N1410, N127);
xor XOR2 (N1428, N1427, N977);
or OR4 (N1429, N1418, N233, N466, N772);
buf BUF1 (N1430, N1423);
not NOT1 (N1431, N1424);
buf BUF1 (N1432, N1428);
nor NOR2 (N1433, N1396, N392);
or OR2 (N1434, N1426, N23);
buf BUF1 (N1435, N1431);
xor XOR2 (N1436, N1409, N1006);
buf BUF1 (N1437, N1430);
or OR3 (N1438, N1432, N930, N1127);
or OR4 (N1439, N1425, N1025, N314, N615);
buf BUF1 (N1440, N1437);
buf BUF1 (N1441, N1436);
xor XOR2 (N1442, N1429, N1278);
and AND2 (N1443, N1438, N75);
and AND4 (N1444, N1440, N835, N1000, N99);
and AND3 (N1445, N1434, N626, N677);
xor XOR2 (N1446, N1435, N1227);
or OR3 (N1447, N1422, N758, N423);
and AND3 (N1448, N1447, N39, N285);
not NOT1 (N1449, N1446);
buf BUF1 (N1450, N1442);
or OR4 (N1451, N1433, N897, N316, N981);
or OR2 (N1452, N1450, N1309);
nor NOR2 (N1453, N1439, N59);
not NOT1 (N1454, N1448);
nor NOR2 (N1455, N1453, N1228);
xor XOR2 (N1456, N1441, N1432);
buf BUF1 (N1457, N1455);
not NOT1 (N1458, N1451);
buf BUF1 (N1459, N1452);
buf BUF1 (N1460, N1454);
and AND2 (N1461, N1444, N177);
nor NOR4 (N1462, N1461, N782, N822, N98);
nand NAND4 (N1463, N1457, N1262, N1202, N486);
buf BUF1 (N1464, N1458);
nand NAND4 (N1465, N1445, N416, N650, N1205);
nor NOR2 (N1466, N1463, N1396);
and AND4 (N1467, N1398, N1065, N104, N253);
or OR2 (N1468, N1466, N782);
and AND4 (N1469, N1465, N103, N379, N538);
buf BUF1 (N1470, N1464);
buf BUF1 (N1471, N1443);
nand NAND4 (N1472, N1449, N836, N1246, N472);
xor XOR2 (N1473, N1460, N565);
xor XOR2 (N1474, N1456, N241);
or OR2 (N1475, N1468, N1101);
and AND2 (N1476, N1473, N531);
xor XOR2 (N1477, N1472, N315);
or OR2 (N1478, N1474, N768);
buf BUF1 (N1479, N1475);
nor NOR4 (N1480, N1462, N1364, N969, N828);
nor NOR3 (N1481, N1476, N227, N13);
not NOT1 (N1482, N1470);
buf BUF1 (N1483, N1467);
not NOT1 (N1484, N1480);
buf BUF1 (N1485, N1477);
or OR4 (N1486, N1482, N528, N953, N929);
not NOT1 (N1487, N1459);
or OR3 (N1488, N1487, N982, N1430);
not NOT1 (N1489, N1471);
and AND2 (N1490, N1488, N1261);
nand NAND3 (N1491, N1481, N583, N697);
not NOT1 (N1492, N1489);
not NOT1 (N1493, N1484);
not NOT1 (N1494, N1479);
xor XOR2 (N1495, N1483, N577);
buf BUF1 (N1496, N1486);
xor XOR2 (N1497, N1478, N1019);
or OR2 (N1498, N1485, N994);
and AND4 (N1499, N1497, N1470, N374, N408);
or OR4 (N1500, N1498, N726, N1139, N1411);
xor XOR2 (N1501, N1490, N1489);
buf BUF1 (N1502, N1494);
and AND4 (N1503, N1469, N137, N828, N1001);
buf BUF1 (N1504, N1492);
not NOT1 (N1505, N1502);
nor NOR3 (N1506, N1500, N663, N454);
and AND2 (N1507, N1506, N678);
nand NAND3 (N1508, N1496, N405, N1500);
not NOT1 (N1509, N1504);
xor XOR2 (N1510, N1495, N1295);
nand NAND3 (N1511, N1510, N428, N634);
and AND4 (N1512, N1509, N1219, N195, N62);
nand NAND2 (N1513, N1501, N608);
nand NAND4 (N1514, N1507, N794, N806, N1360);
and AND3 (N1515, N1511, N764, N995);
or OR4 (N1516, N1508, N930, N999, N778);
buf BUF1 (N1517, N1503);
nand NAND2 (N1518, N1515, N161);
nor NOR2 (N1519, N1514, N669);
or OR4 (N1520, N1512, N39, N880, N291);
and AND2 (N1521, N1516, N790);
nand NAND2 (N1522, N1519, N1221);
nor NOR4 (N1523, N1493, N1176, N844, N1370);
buf BUF1 (N1524, N1499);
nand NAND2 (N1525, N1513, N740);
and AND3 (N1526, N1523, N390, N1435);
xor XOR2 (N1527, N1518, N470);
not NOT1 (N1528, N1520);
or OR2 (N1529, N1505, N418);
nor NOR2 (N1530, N1527, N79);
not NOT1 (N1531, N1528);
not NOT1 (N1532, N1530);
and AND3 (N1533, N1526, N1185, N1377);
not NOT1 (N1534, N1491);
not NOT1 (N1535, N1525);
and AND4 (N1536, N1529, N167, N61, N745);
buf BUF1 (N1537, N1532);
or OR4 (N1538, N1536, N99, N1510, N687);
buf BUF1 (N1539, N1521);
not NOT1 (N1540, N1533);
nor NOR4 (N1541, N1531, N652, N1381, N908);
nor NOR3 (N1542, N1522, N265, N34);
xor XOR2 (N1543, N1542, N1345);
not NOT1 (N1544, N1539);
not NOT1 (N1545, N1534);
not NOT1 (N1546, N1538);
and AND3 (N1547, N1545, N508, N154);
buf BUF1 (N1548, N1546);
xor XOR2 (N1549, N1541, N718);
nand NAND2 (N1550, N1548, N922);
nand NAND4 (N1551, N1524, N1001, N1055, N345);
nor NOR3 (N1552, N1547, N498, N1350);
buf BUF1 (N1553, N1544);
xor XOR2 (N1554, N1549, N293);
nand NAND2 (N1555, N1552, N375);
not NOT1 (N1556, N1551);
nand NAND4 (N1557, N1535, N1436, N897, N1458);
nand NAND2 (N1558, N1555, N1480);
buf BUF1 (N1559, N1556);
nand NAND2 (N1560, N1517, N879);
nand NAND3 (N1561, N1557, N892, N541);
buf BUF1 (N1562, N1553);
or OR2 (N1563, N1562, N1256);
or OR4 (N1564, N1563, N158, N632, N1052);
nor NOR4 (N1565, N1558, N534, N841, N447);
nor NOR4 (N1566, N1560, N217, N687, N60);
buf BUF1 (N1567, N1566);
nand NAND3 (N1568, N1543, N1141, N1471);
and AND3 (N1569, N1564, N405, N1206);
or OR4 (N1570, N1569, N331, N1099, N775);
xor XOR2 (N1571, N1559, N1171);
or OR3 (N1572, N1561, N799, N1013);
nor NOR4 (N1573, N1554, N1261, N1297, N597);
nor NOR4 (N1574, N1571, N86, N1066, N1309);
and AND4 (N1575, N1537, N1330, N1162, N1276);
xor XOR2 (N1576, N1540, N1241);
nand NAND3 (N1577, N1573, N218, N499);
xor XOR2 (N1578, N1572, N290);
and AND4 (N1579, N1565, N371, N819, N888);
nor NOR2 (N1580, N1577, N1061);
xor XOR2 (N1581, N1580, N509);
xor XOR2 (N1582, N1550, N198);
or OR2 (N1583, N1570, N744);
nand NAND3 (N1584, N1578, N1177, N1072);
or OR3 (N1585, N1583, N314, N1215);
nor NOR2 (N1586, N1582, N1523);
buf BUF1 (N1587, N1568);
and AND4 (N1588, N1567, N688, N488, N1399);
nand NAND2 (N1589, N1576, N1345);
not NOT1 (N1590, N1581);
nand NAND4 (N1591, N1584, N700, N1507, N1018);
buf BUF1 (N1592, N1590);
nor NOR2 (N1593, N1592, N1324);
or OR4 (N1594, N1589, N1501, N1182, N239);
nand NAND2 (N1595, N1587, N743);
nor NOR2 (N1596, N1588, N805);
and AND3 (N1597, N1593, N1273, N1173);
nand NAND3 (N1598, N1595, N359, N645);
xor XOR2 (N1599, N1597, N757);
xor XOR2 (N1600, N1579, N1541);
not NOT1 (N1601, N1598);
and AND2 (N1602, N1594, N1305);
or OR3 (N1603, N1574, N963, N1076);
not NOT1 (N1604, N1575);
not NOT1 (N1605, N1596);
nor NOR3 (N1606, N1602, N252, N1383);
and AND3 (N1607, N1606, N836, N1268);
nor NOR3 (N1608, N1603, N1575, N810);
or OR2 (N1609, N1591, N1529);
xor XOR2 (N1610, N1585, N924);
buf BUF1 (N1611, N1604);
nor NOR4 (N1612, N1599, N396, N93, N453);
and AND3 (N1613, N1608, N985, N14);
and AND2 (N1614, N1605, N451);
or OR4 (N1615, N1613, N397, N407, N1164);
or OR2 (N1616, N1586, N318);
xor XOR2 (N1617, N1611, N87);
xor XOR2 (N1618, N1614, N375);
and AND3 (N1619, N1600, N90, N1325);
not NOT1 (N1620, N1601);
buf BUF1 (N1621, N1609);
nor NOR2 (N1622, N1621, N446);
buf BUF1 (N1623, N1620);
not NOT1 (N1624, N1616);
nand NAND2 (N1625, N1624, N1409);
not NOT1 (N1626, N1610);
buf BUF1 (N1627, N1626);
buf BUF1 (N1628, N1623);
not NOT1 (N1629, N1618);
nand NAND2 (N1630, N1627, N945);
and AND3 (N1631, N1630, N345, N150);
and AND2 (N1632, N1631, N1312);
or OR2 (N1633, N1615, N1099);
nor NOR3 (N1634, N1633, N1414, N4);
not NOT1 (N1635, N1607);
and AND2 (N1636, N1619, N154);
nand NAND3 (N1637, N1617, N1498, N544);
nand NAND2 (N1638, N1628, N1348);
or OR4 (N1639, N1637, N931, N454, N236);
and AND4 (N1640, N1625, N723, N1560, N1273);
buf BUF1 (N1641, N1639);
or OR3 (N1642, N1638, N875, N1061);
not NOT1 (N1643, N1629);
and AND4 (N1644, N1622, N654, N1209, N1441);
nor NOR3 (N1645, N1642, N408, N741);
buf BUF1 (N1646, N1634);
not NOT1 (N1647, N1636);
nor NOR4 (N1648, N1641, N971, N1606, N1117);
nor NOR2 (N1649, N1612, N587);
or OR4 (N1650, N1644, N606, N1359, N982);
xor XOR2 (N1651, N1647, N372);
and AND2 (N1652, N1650, N602);
and AND2 (N1653, N1649, N159);
not NOT1 (N1654, N1652);
and AND3 (N1655, N1640, N1536, N1139);
or OR3 (N1656, N1653, N872, N752);
xor XOR2 (N1657, N1635, N574);
not NOT1 (N1658, N1656);
buf BUF1 (N1659, N1648);
xor XOR2 (N1660, N1643, N802);
or OR2 (N1661, N1659, N864);
buf BUF1 (N1662, N1657);
nand NAND3 (N1663, N1660, N815, N1473);
not NOT1 (N1664, N1632);
buf BUF1 (N1665, N1664);
xor XOR2 (N1666, N1646, N165);
nand NAND2 (N1667, N1658, N886);
not NOT1 (N1668, N1655);
buf BUF1 (N1669, N1661);
buf BUF1 (N1670, N1666);
not NOT1 (N1671, N1662);
nand NAND4 (N1672, N1668, N138, N681, N1493);
and AND3 (N1673, N1667, N981, N1460);
nand NAND2 (N1674, N1645, N502);
not NOT1 (N1675, N1673);
or OR2 (N1676, N1671, N509);
and AND2 (N1677, N1663, N1041);
not NOT1 (N1678, N1670);
xor XOR2 (N1679, N1651, N933);
nor NOR3 (N1680, N1674, N1353, N1244);
xor XOR2 (N1681, N1679, N506);
or OR3 (N1682, N1672, N725, N421);
nand NAND4 (N1683, N1677, N1351, N1374, N783);
buf BUF1 (N1684, N1676);
buf BUF1 (N1685, N1681);
or OR3 (N1686, N1678, N258, N76);
buf BUF1 (N1687, N1685);
or OR4 (N1688, N1665, N1082, N880, N202);
buf BUF1 (N1689, N1683);
buf BUF1 (N1690, N1684);
or OR4 (N1691, N1675, N754, N597, N1275);
and AND4 (N1692, N1686, N1137, N317, N1306);
nor NOR2 (N1693, N1669, N272);
nor NOR2 (N1694, N1687, N1589);
not NOT1 (N1695, N1693);
xor XOR2 (N1696, N1654, N90);
buf BUF1 (N1697, N1692);
not NOT1 (N1698, N1695);
or OR2 (N1699, N1696, N74);
or OR3 (N1700, N1688, N970, N384);
buf BUF1 (N1701, N1680);
buf BUF1 (N1702, N1691);
xor XOR2 (N1703, N1700, N1130);
nand NAND4 (N1704, N1697, N400, N1155, N236);
not NOT1 (N1705, N1682);
not NOT1 (N1706, N1704);
nand NAND2 (N1707, N1694, N1150);
xor XOR2 (N1708, N1707, N1629);
nand NAND2 (N1709, N1706, N133);
not NOT1 (N1710, N1705);
or OR3 (N1711, N1690, N427, N615);
xor XOR2 (N1712, N1703, N253);
or OR3 (N1713, N1709, N453, N448);
and AND2 (N1714, N1710, N180);
xor XOR2 (N1715, N1689, N567);
nand NAND3 (N1716, N1711, N98, N515);
buf BUF1 (N1717, N1714);
xor XOR2 (N1718, N1701, N1377);
nor NOR2 (N1719, N1699, N1034);
or OR2 (N1720, N1712, N572);
nor NOR3 (N1721, N1708, N1622, N127);
not NOT1 (N1722, N1720);
buf BUF1 (N1723, N1715);
buf BUF1 (N1724, N1713);
xor XOR2 (N1725, N1698, N450);
and AND3 (N1726, N1717, N1413, N324);
not NOT1 (N1727, N1726);
xor XOR2 (N1728, N1719, N1526);
and AND3 (N1729, N1725, N1673, N1018);
xor XOR2 (N1730, N1728, N1090);
nor NOR4 (N1731, N1702, N1130, N896, N1034);
xor XOR2 (N1732, N1730, N799);
buf BUF1 (N1733, N1722);
xor XOR2 (N1734, N1727, N540);
nand NAND2 (N1735, N1731, N1689);
and AND4 (N1736, N1724, N354, N695, N1091);
or OR4 (N1737, N1721, N1198, N1678, N383);
buf BUF1 (N1738, N1737);
not NOT1 (N1739, N1732);
not NOT1 (N1740, N1729);
not NOT1 (N1741, N1735);
not NOT1 (N1742, N1734);
not NOT1 (N1743, N1736);
nor NOR2 (N1744, N1742, N459);
or OR3 (N1745, N1740, N86, N586);
and AND3 (N1746, N1741, N237, N1019);
and AND4 (N1747, N1745, N218, N1235, N581);
and AND2 (N1748, N1716, N1372);
or OR4 (N1749, N1743, N952, N388, N1049);
buf BUF1 (N1750, N1744);
buf BUF1 (N1751, N1723);
nand NAND3 (N1752, N1739, N1182, N193);
not NOT1 (N1753, N1748);
nor NOR4 (N1754, N1750, N1697, N572, N116);
nand NAND4 (N1755, N1749, N506, N576, N1009);
or OR2 (N1756, N1752, N1461);
and AND4 (N1757, N1751, N272, N1492, N483);
not NOT1 (N1758, N1747);
and AND3 (N1759, N1758, N1516, N351);
nand NAND4 (N1760, N1753, N1586, N1387, N226);
or OR2 (N1761, N1718, N939);
nor NOR3 (N1762, N1733, N621, N140);
or OR2 (N1763, N1757, N735);
or OR3 (N1764, N1738, N1269, N1592);
and AND2 (N1765, N1759, N697);
xor XOR2 (N1766, N1760, N494);
xor XOR2 (N1767, N1766, N1449);
buf BUF1 (N1768, N1754);
xor XOR2 (N1769, N1768, N660);
buf BUF1 (N1770, N1756);
nor NOR3 (N1771, N1765, N732, N340);
xor XOR2 (N1772, N1770, N559);
nor NOR3 (N1773, N1761, N101, N1277);
or OR3 (N1774, N1773, N582, N764);
and AND4 (N1775, N1771, N986, N1208, N1359);
and AND4 (N1776, N1767, N1045, N856, N1577);
buf BUF1 (N1777, N1746);
xor XOR2 (N1778, N1774, N1285);
not NOT1 (N1779, N1763);
nand NAND3 (N1780, N1772, N1288, N81);
nor NOR2 (N1781, N1776, N1408);
nor NOR2 (N1782, N1775, N158);
and AND4 (N1783, N1779, N1635, N805, N974);
xor XOR2 (N1784, N1778, N1284);
or OR4 (N1785, N1784, N1382, N1547, N961);
not NOT1 (N1786, N1783);
and AND3 (N1787, N1780, N1063, N1518);
buf BUF1 (N1788, N1769);
or OR3 (N1789, N1764, N164, N1776);
xor XOR2 (N1790, N1786, N1499);
nand NAND3 (N1791, N1777, N122, N323);
buf BUF1 (N1792, N1790);
buf BUF1 (N1793, N1782);
nand NAND3 (N1794, N1762, N345, N1738);
nor NOR4 (N1795, N1785, N404, N1278, N568);
not NOT1 (N1796, N1791);
not NOT1 (N1797, N1781);
nor NOR4 (N1798, N1787, N1451, N112, N1254);
buf BUF1 (N1799, N1794);
and AND4 (N1800, N1755, N358, N401, N1170);
xor XOR2 (N1801, N1800, N828);
or OR4 (N1802, N1801, N1713, N1278, N145);
or OR2 (N1803, N1792, N279);
not NOT1 (N1804, N1795);
xor XOR2 (N1805, N1793, N366);
xor XOR2 (N1806, N1798, N1517);
and AND2 (N1807, N1806, N981);
not NOT1 (N1808, N1797);
not NOT1 (N1809, N1803);
buf BUF1 (N1810, N1788);
buf BUF1 (N1811, N1808);
not NOT1 (N1812, N1811);
xor XOR2 (N1813, N1796, N833);
nand NAND4 (N1814, N1813, N706, N111, N346);
or OR3 (N1815, N1812, N537, N972);
or OR4 (N1816, N1809, N427, N395, N685);
nor NOR3 (N1817, N1816, N1791, N1645);
or OR2 (N1818, N1799, N1014);
nand NAND3 (N1819, N1805, N392, N1355);
and AND4 (N1820, N1810, N43, N327, N734);
not NOT1 (N1821, N1818);
nor NOR4 (N1822, N1802, N1176, N252, N436);
not NOT1 (N1823, N1814);
xor XOR2 (N1824, N1823, N1165);
and AND2 (N1825, N1824, N1692);
nor NOR4 (N1826, N1815, N793, N1102, N1330);
or OR2 (N1827, N1822, N1378);
and AND3 (N1828, N1807, N1249, N1756);
or OR2 (N1829, N1827, N593);
nor NOR2 (N1830, N1789, N1136);
or OR3 (N1831, N1825, N1297, N1555);
buf BUF1 (N1832, N1828);
or OR3 (N1833, N1804, N905, N478);
not NOT1 (N1834, N1829);
not NOT1 (N1835, N1830);
xor XOR2 (N1836, N1835, N1387);
not NOT1 (N1837, N1819);
and AND3 (N1838, N1834, N1414, N1459);
not NOT1 (N1839, N1826);
or OR2 (N1840, N1833, N1190);
xor XOR2 (N1841, N1820, N1013);
buf BUF1 (N1842, N1832);
buf BUF1 (N1843, N1839);
and AND2 (N1844, N1838, N71);
or OR2 (N1845, N1842, N773);
nor NOR4 (N1846, N1845, N1597, N332, N1258);
buf BUF1 (N1847, N1837);
nand NAND2 (N1848, N1821, N812);
not NOT1 (N1849, N1817);
or OR4 (N1850, N1841, N397, N233, N1485);
nand NAND2 (N1851, N1848, N140);
nor NOR3 (N1852, N1836, N1774, N1262);
xor XOR2 (N1853, N1840, N1010);
nand NAND2 (N1854, N1853, N1352);
nand NAND2 (N1855, N1846, N1852);
xor XOR2 (N1856, N15, N258);
xor XOR2 (N1857, N1847, N227);
and AND4 (N1858, N1857, N1610, N1518, N1091);
or OR3 (N1859, N1849, N803, N1759);
nand NAND3 (N1860, N1831, N478, N828);
or OR4 (N1861, N1851, N788, N1052, N1332);
and AND2 (N1862, N1843, N1408);
nand NAND2 (N1863, N1844, N1485);
buf BUF1 (N1864, N1859);
not NOT1 (N1865, N1858);
nor NOR4 (N1866, N1850, N646, N1658, N205);
xor XOR2 (N1867, N1864, N306);
nor NOR2 (N1868, N1855, N242);
buf BUF1 (N1869, N1861);
xor XOR2 (N1870, N1868, N1094);
not NOT1 (N1871, N1867);
buf BUF1 (N1872, N1870);
or OR3 (N1873, N1869, N513, N1371);
and AND4 (N1874, N1866, N335, N554, N145);
not NOT1 (N1875, N1872);
nor NOR2 (N1876, N1862, N1228);
nand NAND3 (N1877, N1876, N1351, N157);
buf BUF1 (N1878, N1877);
nor NOR4 (N1879, N1860, N43, N1272, N1018);
or OR4 (N1880, N1854, N1498, N1594, N158);
buf BUF1 (N1881, N1863);
and AND2 (N1882, N1874, N334);
and AND4 (N1883, N1881, N1858, N55, N494);
nor NOR2 (N1884, N1882, N1451);
or OR3 (N1885, N1883, N324, N372);
nand NAND2 (N1886, N1884, N1722);
buf BUF1 (N1887, N1873);
nor NOR4 (N1888, N1880, N533, N316, N1802);
and AND3 (N1889, N1885, N591, N1279);
nor NOR4 (N1890, N1889, N1481, N202, N1584);
and AND2 (N1891, N1890, N1567);
and AND2 (N1892, N1888, N84);
not NOT1 (N1893, N1886);
nor NOR4 (N1894, N1887, N541, N535, N1632);
xor XOR2 (N1895, N1892, N1177);
or OR4 (N1896, N1893, N712, N1435, N504);
nor NOR2 (N1897, N1875, N38);
nor NOR4 (N1898, N1878, N1298, N686, N1524);
not NOT1 (N1899, N1894);
or OR3 (N1900, N1895, N1060, N197);
buf BUF1 (N1901, N1900);
not NOT1 (N1902, N1856);
and AND4 (N1903, N1898, N223, N1196, N505);
or OR3 (N1904, N1891, N1285, N908);
or OR4 (N1905, N1865, N191, N426, N137);
not NOT1 (N1906, N1879);
xor XOR2 (N1907, N1906, N1267);
nand NAND3 (N1908, N1902, N336, N792);
and AND3 (N1909, N1871, N22, N373);
nor NOR2 (N1910, N1897, N28);
not NOT1 (N1911, N1908);
or OR4 (N1912, N1901, N1215, N677, N1346);
buf BUF1 (N1913, N1912);
or OR3 (N1914, N1910, N159, N266);
nand NAND4 (N1915, N1913, N541, N1895, N870);
buf BUF1 (N1916, N1907);
nand NAND3 (N1917, N1904, N1588, N7);
and AND3 (N1918, N1899, N1319, N469);
not NOT1 (N1919, N1914);
and AND4 (N1920, N1896, N1534, N1405, N1144);
xor XOR2 (N1921, N1918, N846);
nor NOR4 (N1922, N1909, N1240, N770, N738);
nand NAND2 (N1923, N1921, N1643);
or OR2 (N1924, N1920, N1324);
not NOT1 (N1925, N1911);
nor NOR4 (N1926, N1923, N637, N858, N1757);
nor NOR3 (N1927, N1926, N173, N312);
buf BUF1 (N1928, N1916);
buf BUF1 (N1929, N1903);
nand NAND3 (N1930, N1928, N965, N185);
and AND3 (N1931, N1925, N1079, N325);
not NOT1 (N1932, N1915);
and AND3 (N1933, N1919, N882, N1341);
buf BUF1 (N1934, N1931);
xor XOR2 (N1935, N1933, N1289);
nor NOR4 (N1936, N1905, N1882, N406, N865);
nor NOR3 (N1937, N1927, N166, N654);
nand NAND2 (N1938, N1924, N677);
and AND2 (N1939, N1929, N1927);
nand NAND4 (N1940, N1922, N171, N849, N121);
buf BUF1 (N1941, N1932);
and AND3 (N1942, N1938, N954, N1170);
nand NAND2 (N1943, N1942, N480);
buf BUF1 (N1944, N1936);
xor XOR2 (N1945, N1917, N1349);
xor XOR2 (N1946, N1941, N326);
xor XOR2 (N1947, N1943, N22);
xor XOR2 (N1948, N1940, N1459);
buf BUF1 (N1949, N1930);
not NOT1 (N1950, N1939);
or OR2 (N1951, N1945, N902);
buf BUF1 (N1952, N1934);
nand NAND2 (N1953, N1948, N71);
nor NOR3 (N1954, N1949, N1303, N102);
buf BUF1 (N1955, N1937);
buf BUF1 (N1956, N1947);
nand NAND4 (N1957, N1954, N1066, N1241, N700);
or OR2 (N1958, N1955, N1457);
xor XOR2 (N1959, N1953, N1214);
or OR2 (N1960, N1957, N1030);
buf BUF1 (N1961, N1950);
xor XOR2 (N1962, N1935, N77);
xor XOR2 (N1963, N1956, N1097);
nor NOR3 (N1964, N1959, N76, N1668);
xor XOR2 (N1965, N1961, N148);
and AND2 (N1966, N1944, N671);
and AND3 (N1967, N1965, N1904, N334);
and AND4 (N1968, N1952, N785, N128, N1309);
nor NOR3 (N1969, N1960, N986, N1169);
buf BUF1 (N1970, N1958);
or OR4 (N1971, N1946, N1947, N1644, N94);
buf BUF1 (N1972, N1966);
and AND4 (N1973, N1962, N1289, N1946, N1291);
nor NOR4 (N1974, N1970, N1453, N524, N160);
xor XOR2 (N1975, N1973, N1054);
buf BUF1 (N1976, N1968);
not NOT1 (N1977, N1964);
buf BUF1 (N1978, N1977);
or OR2 (N1979, N1974, N522);
nor NOR2 (N1980, N1976, N905);
nand NAND3 (N1981, N1969, N625, N926);
or OR3 (N1982, N1979, N750, N1137);
xor XOR2 (N1983, N1967, N883);
buf BUF1 (N1984, N1978);
or OR2 (N1985, N1971, N839);
not NOT1 (N1986, N1982);
buf BUF1 (N1987, N1981);
xor XOR2 (N1988, N1951, N588);
xor XOR2 (N1989, N1972, N1153);
not NOT1 (N1990, N1988);
nand NAND4 (N1991, N1985, N391, N1726, N1400);
or OR2 (N1992, N1980, N166);
nand NAND3 (N1993, N1990, N1256, N334);
buf BUF1 (N1994, N1983);
buf BUF1 (N1995, N1975);
buf BUF1 (N1996, N1963);
nand NAND4 (N1997, N1992, N1293, N1829, N863);
xor XOR2 (N1998, N1993, N840);
buf BUF1 (N1999, N1989);
nand NAND4 (N2000, N1991, N222, N103, N392);
xor XOR2 (N2001, N1987, N1051);
xor XOR2 (N2002, N2001, N714);
nand NAND4 (N2003, N2000, N951, N1972, N1433);
nor NOR3 (N2004, N2002, N1780, N1679);
and AND2 (N2005, N1984, N444);
nor NOR3 (N2006, N1995, N405, N1270);
or OR4 (N2007, N1994, N1017, N1363, N1158);
and AND2 (N2008, N2003, N1565);
not NOT1 (N2009, N2008);
not NOT1 (N2010, N2005);
or OR4 (N2011, N1997, N697, N143, N378);
not NOT1 (N2012, N1999);
nor NOR3 (N2013, N2009, N64, N320);
nand NAND4 (N2014, N1986, N1133, N1253, N64);
nand NAND3 (N2015, N2006, N1278, N1450);
and AND4 (N2016, N2013, N257, N501, N1529);
buf BUF1 (N2017, N2010);
nor NOR3 (N2018, N2004, N1444, N1278);
nor NOR3 (N2019, N2016, N527, N1198);
nand NAND2 (N2020, N2015, N511);
and AND4 (N2021, N2017, N1206, N818, N718);
nand NAND4 (N2022, N2012, N11, N591, N897);
nor NOR2 (N2023, N2020, N143);
xor XOR2 (N2024, N1996, N171);
not NOT1 (N2025, N2019);
nand NAND4 (N2026, N2022, N1201, N132, N1955);
not NOT1 (N2027, N2007);
and AND3 (N2028, N1998, N1483, N1232);
and AND4 (N2029, N2028, N796, N468, N1069);
not NOT1 (N2030, N2025);
nor NOR3 (N2031, N2011, N1031, N798);
and AND2 (N2032, N2021, N879);
xor XOR2 (N2033, N2024, N1381);
or OR3 (N2034, N2026, N329, N12);
or OR4 (N2035, N2033, N1383, N1332, N1217);
or OR3 (N2036, N2034, N1895, N444);
and AND2 (N2037, N2018, N583);
or OR3 (N2038, N2030, N1806, N1134);
not NOT1 (N2039, N2038);
and AND3 (N2040, N2037, N1735, N1569);
xor XOR2 (N2041, N2040, N1326);
xor XOR2 (N2042, N2029, N1024);
nor NOR3 (N2043, N2042, N54, N385);
buf BUF1 (N2044, N2014);
or OR3 (N2045, N2035, N1835, N1032);
nand NAND4 (N2046, N2043, N231, N1257, N1999);
nand NAND4 (N2047, N2023, N647, N1298, N565);
and AND3 (N2048, N2039, N1853, N117);
nor NOR4 (N2049, N2044, N1825, N1995, N1510);
nand NAND2 (N2050, N2036, N1453);
buf BUF1 (N2051, N2027);
and AND3 (N2052, N2051, N1087, N529);
xor XOR2 (N2053, N2047, N1196);
nand NAND4 (N2054, N2050, N223, N1791, N1043);
xor XOR2 (N2055, N2032, N1189);
not NOT1 (N2056, N2031);
or OR4 (N2057, N2045, N1015, N1549, N1095);
or OR4 (N2058, N2053, N1614, N1577, N96);
buf BUF1 (N2059, N2052);
nor NOR2 (N2060, N2056, N1817);
nor NOR4 (N2061, N2049, N2013, N1792, N1092);
buf BUF1 (N2062, N2060);
nand NAND4 (N2063, N2058, N1813, N1267, N888);
or OR4 (N2064, N2062, N817, N1348, N2028);
and AND3 (N2065, N2059, N863, N627);
not NOT1 (N2066, N2061);
nor NOR4 (N2067, N2064, N76, N674, N452);
nor NOR4 (N2068, N2067, N1299, N549, N822);
not NOT1 (N2069, N2068);
or OR4 (N2070, N2065, N445, N1687, N1879);
or OR4 (N2071, N2066, N2041, N829, N120);
or OR4 (N2072, N1520, N1621, N1761, N1654);
not NOT1 (N2073, N2048);
and AND3 (N2074, N2057, N409, N651);
nor NOR3 (N2075, N2070, N198, N566);
and AND4 (N2076, N2071, N1442, N360, N326);
not NOT1 (N2077, N2054);
not NOT1 (N2078, N2074);
xor XOR2 (N2079, N2077, N1263);
and AND3 (N2080, N2073, N1251, N319);
nand NAND4 (N2081, N2080, N45, N395, N285);
nor NOR3 (N2082, N2078, N210, N647);
or OR4 (N2083, N2082, N28, N989, N300);
nor NOR4 (N2084, N2076, N2077, N732, N1985);
and AND3 (N2085, N2063, N1590, N1491);
nand NAND2 (N2086, N2085, N931);
buf BUF1 (N2087, N2084);
or OR2 (N2088, N2075, N356);
buf BUF1 (N2089, N2046);
nand NAND4 (N2090, N2089, N169, N198, N1499);
or OR2 (N2091, N2087, N661);
or OR3 (N2092, N2086, N462, N2075);
nand NAND4 (N2093, N2091, N66, N277, N250);
not NOT1 (N2094, N2079);
or OR4 (N2095, N2081, N1324, N1120, N810);
xor XOR2 (N2096, N2072, N401);
and AND3 (N2097, N2095, N1644, N525);
xor XOR2 (N2098, N2088, N627);
xor XOR2 (N2099, N2096, N704);
nor NOR3 (N2100, N2093, N1819, N1024);
nand NAND2 (N2101, N2055, N279);
or OR3 (N2102, N2092, N353, N1040);
or OR3 (N2103, N2102, N1869, N363);
buf BUF1 (N2104, N2100);
and AND3 (N2105, N2104, N32, N1840);
nand NAND3 (N2106, N2090, N1322, N1729);
xor XOR2 (N2107, N2098, N233);
nand NAND4 (N2108, N2103, N598, N1470, N1792);
and AND2 (N2109, N2069, N1716);
or OR2 (N2110, N2094, N1454);
buf BUF1 (N2111, N2107);
nand NAND3 (N2112, N2110, N760, N74);
buf BUF1 (N2113, N2112);
xor XOR2 (N2114, N2083, N1912);
and AND2 (N2115, N2106, N1400);
and AND2 (N2116, N2097, N1624);
or OR3 (N2117, N2111, N420, N1872);
and AND3 (N2118, N2116, N158, N438);
nand NAND2 (N2119, N2113, N1204);
nor NOR2 (N2120, N2099, N141);
nand NAND3 (N2121, N2105, N695, N261);
not NOT1 (N2122, N2117);
buf BUF1 (N2123, N2101);
and AND2 (N2124, N2122, N1172);
not NOT1 (N2125, N2109);
and AND3 (N2126, N2121, N1155, N384);
or OR4 (N2127, N2119, N1019, N2027, N1544);
or OR3 (N2128, N2124, N907, N1848);
and AND2 (N2129, N2115, N1181);
nand NAND4 (N2130, N2120, N1396, N1839, N327);
nor NOR3 (N2131, N2127, N280, N2027);
xor XOR2 (N2132, N2129, N1765);
or OR2 (N2133, N2132, N1151);
or OR2 (N2134, N2133, N552);
nand NAND3 (N2135, N2134, N1915, N1192);
nor NOR2 (N2136, N2126, N1895);
buf BUF1 (N2137, N2123);
nand NAND4 (N2138, N2131, N23, N785, N1683);
xor XOR2 (N2139, N2137, N1542);
nand NAND4 (N2140, N2118, N1982, N1658, N371);
nor NOR2 (N2141, N2140, N561);
buf BUF1 (N2142, N2125);
not NOT1 (N2143, N2136);
nand NAND3 (N2144, N2143, N1006, N1886);
xor XOR2 (N2145, N2142, N1943);
nand NAND3 (N2146, N2108, N76, N760);
or OR4 (N2147, N2145, N1800, N889, N1171);
buf BUF1 (N2148, N2144);
buf BUF1 (N2149, N2146);
and AND4 (N2150, N2147, N496, N920, N68);
nand NAND3 (N2151, N2149, N20, N242);
nand NAND2 (N2152, N2151, N544);
and AND2 (N2153, N2135, N1335);
nand NAND3 (N2154, N2139, N205, N461);
nor NOR2 (N2155, N2138, N1131);
or OR3 (N2156, N2154, N1560, N2001);
and AND3 (N2157, N2152, N835, N1845);
and AND4 (N2158, N2148, N789, N236, N620);
buf BUF1 (N2159, N2150);
not NOT1 (N2160, N2155);
buf BUF1 (N2161, N2159);
not NOT1 (N2162, N2156);
nand NAND4 (N2163, N2161, N101, N933, N1318);
not NOT1 (N2164, N2157);
or OR4 (N2165, N2114, N1440, N587, N1694);
and AND2 (N2166, N2160, N1727);
not NOT1 (N2167, N2165);
or OR3 (N2168, N2128, N1392, N1636);
or OR4 (N2169, N2168, N1956, N25, N904);
not NOT1 (N2170, N2167);
buf BUF1 (N2171, N2169);
nor NOR3 (N2172, N2158, N1056, N1960);
not NOT1 (N2173, N2164);
not NOT1 (N2174, N2130);
nor NOR3 (N2175, N2170, N473, N1236);
xor XOR2 (N2176, N2172, N1124);
nand NAND3 (N2177, N2173, N767, N296);
or OR4 (N2178, N2141, N911, N531, N145);
nor NOR2 (N2179, N2153, N1216);
or OR2 (N2180, N2166, N731);
buf BUF1 (N2181, N2178);
or OR4 (N2182, N2179, N147, N467, N1513);
nor NOR2 (N2183, N2162, N850);
not NOT1 (N2184, N2181);
not NOT1 (N2185, N2180);
and AND2 (N2186, N2185, N2133);
nand NAND3 (N2187, N2171, N264, N852);
buf BUF1 (N2188, N2187);
buf BUF1 (N2189, N2175);
not NOT1 (N2190, N2163);
buf BUF1 (N2191, N2188);
nor NOR4 (N2192, N2182, N221, N2095, N1737);
xor XOR2 (N2193, N2176, N669);
nand NAND3 (N2194, N2193, N1060, N1527);
xor XOR2 (N2195, N2192, N1768);
and AND3 (N2196, N2177, N1074, N1752);
xor XOR2 (N2197, N2195, N2150);
xor XOR2 (N2198, N2190, N1425);
nor NOR2 (N2199, N2189, N956);
nand NAND4 (N2200, N2197, N1282, N2047, N1000);
and AND3 (N2201, N2174, N461, N1687);
not NOT1 (N2202, N2198);
and AND2 (N2203, N2194, N1595);
or OR2 (N2204, N2203, N983);
not NOT1 (N2205, N2199);
and AND4 (N2206, N2205, N800, N1531, N2126);
buf BUF1 (N2207, N2200);
nand NAND4 (N2208, N2183, N1089, N243, N805);
and AND2 (N2209, N2196, N1646);
nand NAND4 (N2210, N2184, N1085, N2052, N409);
nand NAND2 (N2211, N2191, N1288);
or OR2 (N2212, N2208, N551);
buf BUF1 (N2213, N2201);
buf BUF1 (N2214, N2211);
buf BUF1 (N2215, N2209);
buf BUF1 (N2216, N2207);
or OR3 (N2217, N2212, N1480, N1399);
xor XOR2 (N2218, N2216, N1780);
nand NAND3 (N2219, N2218, N1902, N285);
nor NOR2 (N2220, N2204, N2152);
nor NOR3 (N2221, N2206, N1147, N2066);
buf BUF1 (N2222, N2202);
and AND3 (N2223, N2221, N1471, N1480);
buf BUF1 (N2224, N2220);
xor XOR2 (N2225, N2222, N1767);
or OR4 (N2226, N2219, N208, N922, N1782);
or OR2 (N2227, N2225, N1422);
nor NOR4 (N2228, N2224, N638, N90, N376);
nor NOR2 (N2229, N2227, N811);
not NOT1 (N2230, N2226);
xor XOR2 (N2231, N2217, N93);
xor XOR2 (N2232, N2231, N2045);
or OR2 (N2233, N2186, N1411);
xor XOR2 (N2234, N2232, N1246);
not NOT1 (N2235, N2210);
nor NOR2 (N2236, N2223, N695);
nand NAND3 (N2237, N2230, N1386, N321);
or OR2 (N2238, N2235, N1505);
buf BUF1 (N2239, N2228);
nand NAND2 (N2240, N2213, N1675);
not NOT1 (N2241, N2238);
buf BUF1 (N2242, N2229);
nand NAND4 (N2243, N2239, N891, N106, N700);
xor XOR2 (N2244, N2233, N743);
nor NOR4 (N2245, N2244, N347, N1657, N1893);
xor XOR2 (N2246, N2234, N1167);
and AND3 (N2247, N2240, N2097, N1352);
nand NAND2 (N2248, N2243, N1607);
not NOT1 (N2249, N2241);
xor XOR2 (N2250, N2249, N2032);
not NOT1 (N2251, N2247);
buf BUF1 (N2252, N2250);
buf BUF1 (N2253, N2237);
not NOT1 (N2254, N2214);
not NOT1 (N2255, N2215);
and AND2 (N2256, N2252, N92);
and AND4 (N2257, N2254, N743, N965, N1480);
not NOT1 (N2258, N2248);
or OR3 (N2259, N2257, N2219, N1299);
buf BUF1 (N2260, N2253);
and AND4 (N2261, N2260, N2051, N1722, N1871);
nor NOR2 (N2262, N2242, N1510);
nor NOR3 (N2263, N2258, N528, N1392);
not NOT1 (N2264, N2245);
xor XOR2 (N2265, N2236, N1174);
nor NOR2 (N2266, N2251, N421);
nor NOR2 (N2267, N2246, N261);
and AND2 (N2268, N2261, N1512);
nor NOR4 (N2269, N2266, N1975, N933, N1821);
xor XOR2 (N2270, N2264, N1739);
and AND2 (N2271, N2262, N491);
nor NOR3 (N2272, N2269, N68, N1354);
buf BUF1 (N2273, N2265);
nand NAND2 (N2274, N2263, N1898);
nor NOR3 (N2275, N2268, N1446, N1086);
xor XOR2 (N2276, N2273, N316);
xor XOR2 (N2277, N2275, N1692);
nand NAND2 (N2278, N2272, N1869);
or OR3 (N2279, N2271, N307, N1435);
and AND2 (N2280, N2270, N213);
not NOT1 (N2281, N2274);
xor XOR2 (N2282, N2277, N1993);
buf BUF1 (N2283, N2281);
or OR4 (N2284, N2280, N1831, N1068, N1047);
buf BUF1 (N2285, N2255);
xor XOR2 (N2286, N2282, N2274);
and AND3 (N2287, N2284, N772, N1391);
and AND4 (N2288, N2283, N1832, N31, N1615);
xor XOR2 (N2289, N2259, N628);
nor NOR3 (N2290, N2289, N2062, N530);
or OR3 (N2291, N2285, N1097, N1937);
not NOT1 (N2292, N2286);
nand NAND2 (N2293, N2290, N735);
buf BUF1 (N2294, N2279);
not NOT1 (N2295, N2287);
nand NAND3 (N2296, N2293, N989, N1547);
not NOT1 (N2297, N2267);
and AND4 (N2298, N2288, N1577, N1785, N364);
buf BUF1 (N2299, N2278);
and AND3 (N2300, N2296, N1145, N1414);
or OR2 (N2301, N2297, N1796);
and AND4 (N2302, N2298, N1494, N1378, N1695);
nor NOR2 (N2303, N2299, N64);
and AND2 (N2304, N2301, N2024);
and AND4 (N2305, N2302, N1832, N1400, N527);
nor NOR2 (N2306, N2300, N1886);
xor XOR2 (N2307, N2294, N1342);
buf BUF1 (N2308, N2291);
and AND3 (N2309, N2292, N8, N2252);
xor XOR2 (N2310, N2308, N2238);
buf BUF1 (N2311, N2256);
xor XOR2 (N2312, N2304, N213);
not NOT1 (N2313, N2311);
buf BUF1 (N2314, N2309);
xor XOR2 (N2315, N2313, N1521);
not NOT1 (N2316, N2295);
and AND3 (N2317, N2315, N1749, N503);
nand NAND2 (N2318, N2314, N2267);
and AND2 (N2319, N2317, N278);
buf BUF1 (N2320, N2307);
or OR2 (N2321, N2306, N2069);
or OR2 (N2322, N2276, N1824);
and AND3 (N2323, N2319, N238, N1731);
xor XOR2 (N2324, N2322, N549);
and AND3 (N2325, N2320, N1086, N422);
nand NAND4 (N2326, N2316, N1309, N1866, N1373);
not NOT1 (N2327, N2325);
buf BUF1 (N2328, N2312);
not NOT1 (N2329, N2324);
not NOT1 (N2330, N2321);
and AND3 (N2331, N2323, N1153, N1343);
not NOT1 (N2332, N2330);
nand NAND3 (N2333, N2332, N787, N1345);
nor NOR2 (N2334, N2318, N1267);
buf BUF1 (N2335, N2305);
nand NAND4 (N2336, N2303, N716, N1100, N219);
xor XOR2 (N2337, N2328, N729);
not NOT1 (N2338, N2334);
nand NAND2 (N2339, N2338, N1920);
buf BUF1 (N2340, N2331);
buf BUF1 (N2341, N2336);
not NOT1 (N2342, N2341);
not NOT1 (N2343, N2333);
or OR4 (N2344, N2335, N2013, N1366, N782);
not NOT1 (N2345, N2329);
xor XOR2 (N2346, N2344, N1846);
not NOT1 (N2347, N2310);
not NOT1 (N2348, N2337);
xor XOR2 (N2349, N2326, N2177);
or OR3 (N2350, N2348, N1973, N1785);
and AND2 (N2351, N2340, N2280);
or OR4 (N2352, N2327, N169, N225, N1104);
nor NOR4 (N2353, N2342, N850, N350, N1547);
not NOT1 (N2354, N2352);
and AND3 (N2355, N2351, N416, N1244);
buf BUF1 (N2356, N2339);
xor XOR2 (N2357, N2347, N1417);
xor XOR2 (N2358, N2356, N1516);
nand NAND4 (N2359, N2350, N1084, N843, N1760);
and AND2 (N2360, N2357, N1989);
xor XOR2 (N2361, N2355, N939);
nand NAND4 (N2362, N2353, N91, N2299, N392);
nand NAND3 (N2363, N2349, N1094, N1856);
and AND2 (N2364, N2362, N1881);
and AND2 (N2365, N2363, N1037);
and AND3 (N2366, N2359, N321, N1539);
nand NAND2 (N2367, N2361, N361);
or OR2 (N2368, N2365, N1162);
xor XOR2 (N2369, N2343, N2152);
or OR4 (N2370, N2345, N2224, N970, N1748);
nand NAND3 (N2371, N2368, N2138, N1856);
and AND3 (N2372, N2366, N2088, N78);
nand NAND4 (N2373, N2360, N467, N393, N1295);
and AND2 (N2374, N2358, N1653);
xor XOR2 (N2375, N2369, N368);
buf BUF1 (N2376, N2371);
or OR3 (N2377, N2372, N310, N1535);
buf BUF1 (N2378, N2370);
xor XOR2 (N2379, N2367, N2082);
nand NAND3 (N2380, N2373, N46, N1746);
or OR4 (N2381, N2378, N779, N1972, N1581);
not NOT1 (N2382, N2354);
and AND4 (N2383, N2380, N1103, N78, N1134);
and AND3 (N2384, N2377, N1239, N1865);
buf BUF1 (N2385, N2376);
xor XOR2 (N2386, N2385, N2062);
or OR2 (N2387, N2379, N772);
or OR4 (N2388, N2387, N1388, N897, N1012);
or OR3 (N2389, N2386, N1133, N2187);
buf BUF1 (N2390, N2389);
xor XOR2 (N2391, N2390, N857);
not NOT1 (N2392, N2391);
xor XOR2 (N2393, N2392, N958);
nor NOR4 (N2394, N2384, N234, N1944, N724);
or OR3 (N2395, N2393, N919, N2328);
or OR2 (N2396, N2374, N532);
nand NAND4 (N2397, N2395, N1649, N1079, N1314);
and AND4 (N2398, N2388, N27, N1447, N1715);
xor XOR2 (N2399, N2394, N2185);
xor XOR2 (N2400, N2398, N393);
nor NOR2 (N2401, N2381, N886);
and AND3 (N2402, N2399, N422, N707);
nand NAND4 (N2403, N2375, N85, N2214, N425);
not NOT1 (N2404, N2397);
buf BUF1 (N2405, N2400);
xor XOR2 (N2406, N2396, N1669);
buf BUF1 (N2407, N2404);
xor XOR2 (N2408, N2402, N1943);
not NOT1 (N2409, N2401);
nand NAND2 (N2410, N2383, N123);
nand NAND3 (N2411, N2407, N395, N1798);
nand NAND2 (N2412, N2409, N873);
xor XOR2 (N2413, N2364, N1162);
not NOT1 (N2414, N2408);
nor NOR4 (N2415, N2406, N1511, N2133, N598);
xor XOR2 (N2416, N2411, N1332);
not NOT1 (N2417, N2405);
nor NOR4 (N2418, N2414, N1360, N852, N306);
xor XOR2 (N2419, N2403, N2107);
or OR4 (N2420, N2419, N2373, N2202, N1456);
or OR4 (N2421, N2410, N33, N1123, N1291);
nand NAND3 (N2422, N2418, N410, N305);
not NOT1 (N2423, N2421);
nor NOR4 (N2424, N2412, N290, N459, N2178);
nand NAND3 (N2425, N2424, N1516, N136);
xor XOR2 (N2426, N2422, N1551);
nand NAND2 (N2427, N2413, N1693);
nor NOR3 (N2428, N2346, N1709, N1056);
not NOT1 (N2429, N2427);
and AND3 (N2430, N2420, N238, N853);
or OR3 (N2431, N2430, N1694, N1831);
nand NAND2 (N2432, N2416, N1397);
xor XOR2 (N2433, N2428, N2270);
xor XOR2 (N2434, N2423, N1767);
not NOT1 (N2435, N2415);
not NOT1 (N2436, N2425);
buf BUF1 (N2437, N2426);
or OR3 (N2438, N2437, N486, N1481);
xor XOR2 (N2439, N2433, N2272);
or OR2 (N2440, N2439, N1072);
xor XOR2 (N2441, N2417, N297);
not NOT1 (N2442, N2438);
xor XOR2 (N2443, N2431, N137);
and AND2 (N2444, N2443, N1204);
buf BUF1 (N2445, N2442);
and AND3 (N2446, N2429, N860, N1173);
or OR4 (N2447, N2382, N26, N2223, N1772);
not NOT1 (N2448, N2432);
or OR2 (N2449, N2436, N2202);
xor XOR2 (N2450, N2444, N367);
or OR2 (N2451, N2450, N1121);
or OR4 (N2452, N2445, N1434, N800, N2047);
not NOT1 (N2453, N2447);
not NOT1 (N2454, N2453);
xor XOR2 (N2455, N2452, N736);
and AND4 (N2456, N2448, N1531, N1326, N2302);
not NOT1 (N2457, N2446);
nand NAND4 (N2458, N2435, N1766, N948, N412);
nand NAND3 (N2459, N2449, N497, N1495);
buf BUF1 (N2460, N2457);
and AND4 (N2461, N2451, N1471, N852, N907);
and AND4 (N2462, N2456, N800, N556, N1772);
or OR4 (N2463, N2454, N326, N1917, N1480);
or OR4 (N2464, N2459, N1190, N2107, N2068);
buf BUF1 (N2465, N2434);
xor XOR2 (N2466, N2463, N524);
or OR2 (N2467, N2440, N635);
and AND3 (N2468, N2464, N1505, N2283);
nand NAND2 (N2469, N2461, N979);
buf BUF1 (N2470, N2467);
and AND2 (N2471, N2455, N2325);
or OR2 (N2472, N2468, N1256);
and AND4 (N2473, N2462, N1630, N2377, N1015);
not NOT1 (N2474, N2465);
xor XOR2 (N2475, N2441, N108);
not NOT1 (N2476, N2475);
xor XOR2 (N2477, N2476, N72);
not NOT1 (N2478, N2460);
and AND3 (N2479, N2466, N1153, N1613);
or OR3 (N2480, N2473, N183, N2099);
nand NAND3 (N2481, N2458, N328, N510);
nor NOR2 (N2482, N2471, N211);
buf BUF1 (N2483, N2477);
nand NAND2 (N2484, N2470, N811);
and AND2 (N2485, N2480, N562);
nand NAND4 (N2486, N2474, N750, N985, N632);
xor XOR2 (N2487, N2469, N1513);
nand NAND3 (N2488, N2487, N525, N704);
buf BUF1 (N2489, N2481);
nor NOR2 (N2490, N2472, N1869);
buf BUF1 (N2491, N2490);
or OR4 (N2492, N2483, N1806, N1840, N1989);
nor NOR2 (N2493, N2484, N1529);
nand NAND4 (N2494, N2491, N1777, N1252, N1503);
and AND2 (N2495, N2494, N597);
nor NOR3 (N2496, N2478, N658, N2130);
xor XOR2 (N2497, N2482, N1806);
or OR2 (N2498, N2489, N1191);
buf BUF1 (N2499, N2492);
buf BUF1 (N2500, N2488);
or OR2 (N2501, N2497, N697);
or OR3 (N2502, N2485, N600, N1944);
or OR2 (N2503, N2498, N108);
or OR4 (N2504, N2496, N147, N1564, N1612);
nand NAND3 (N2505, N2501, N332, N1916);
xor XOR2 (N2506, N2493, N845);
nand NAND4 (N2507, N2500, N1562, N1357, N1057);
and AND2 (N2508, N2507, N198);
not NOT1 (N2509, N2495);
not NOT1 (N2510, N2486);
or OR2 (N2511, N2506, N2346);
xor XOR2 (N2512, N2504, N2415);
not NOT1 (N2513, N2509);
or OR3 (N2514, N2510, N511, N958);
not NOT1 (N2515, N2479);
or OR4 (N2516, N2499, N622, N293, N151);
not NOT1 (N2517, N2512);
nand NAND2 (N2518, N2515, N1656);
or OR2 (N2519, N2508, N440);
buf BUF1 (N2520, N2518);
nand NAND4 (N2521, N2517, N722, N2032, N320);
endmodule