// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12;

output N282,N305,N309,N301,N293,N303,N302,N310,N311,N312;

nand NAND2 (N13, N8, N11);
nand NAND4 (N14, N5, N7, N8, N7);
nor NOR4 (N15, N10, N2, N6, N9);
buf BUF1 (N16, N13);
or OR2 (N17, N10, N4);
not NOT1 (N18, N5);
nand NAND3 (N19, N16, N1, N11);
nor NOR3 (N20, N15, N1, N19);
not NOT1 (N21, N10);
and AND4 (N22, N5, N3, N14, N5);
xor XOR2 (N23, N15, N7);
nand NAND3 (N24, N18, N21, N19);
nand NAND3 (N25, N1, N20, N21);
and AND2 (N26, N8, N24);
buf BUF1 (N27, N23);
or OR3 (N28, N11, N14, N22);
buf BUF1 (N29, N23);
or OR4 (N30, N18, N18, N23, N5);
nand NAND2 (N31, N11, N14);
nand NAND4 (N32, N26, N25, N7, N29);
xor XOR2 (N33, N30, N21);
not NOT1 (N34, N25);
not NOT1 (N35, N11);
buf BUF1 (N36, N32);
or OR2 (N37, N2, N2);
and AND4 (N38, N27, N22, N1, N19);
nand NAND4 (N39, N21, N24, N37, N19);
xor XOR2 (N40, N19, N38);
buf BUF1 (N41, N11);
nand NAND3 (N42, N36, N36, N34);
not NOT1 (N43, N34);
xor XOR2 (N44, N31, N22);
xor XOR2 (N45, N41, N40);
not NOT1 (N46, N12);
and AND4 (N47, N28, N16, N10, N14);
or OR4 (N48, N42, N25, N12, N47);
nand NAND2 (N49, N29, N43);
buf BUF1 (N50, N33);
or OR3 (N51, N2, N42, N37);
buf BUF1 (N52, N49);
or OR2 (N53, N46, N28);
buf BUF1 (N54, N51);
buf BUF1 (N55, N45);
nor NOR3 (N56, N55, N49, N51);
nand NAND3 (N57, N35, N2, N22);
nand NAND4 (N58, N53, N38, N45, N6);
or OR2 (N59, N44, N22);
and AND3 (N60, N39, N23, N20);
or OR2 (N61, N56, N35);
nor NOR2 (N62, N58, N10);
nand NAND2 (N63, N48, N47);
not NOT1 (N64, N62);
nor NOR4 (N65, N52, N36, N47, N4);
xor XOR2 (N66, N50, N19);
or OR4 (N67, N64, N63, N19, N18);
nor NOR4 (N68, N6, N59, N16, N61);
and AND2 (N69, N63, N50);
xor XOR2 (N70, N63, N13);
nand NAND3 (N71, N57, N60, N13);
not NOT1 (N72, N48);
and AND3 (N73, N70, N58, N27);
or OR2 (N74, N71, N68);
or OR2 (N75, N70, N41);
xor XOR2 (N76, N74, N61);
nor NOR4 (N77, N72, N61, N63, N73);
xor XOR2 (N78, N44, N13);
not NOT1 (N79, N69);
nor NOR2 (N80, N65, N71);
not NOT1 (N81, N54);
buf BUF1 (N82, N79);
nor NOR4 (N83, N75, N34, N45, N76);
nand NAND3 (N84, N58, N33, N61);
xor XOR2 (N85, N77, N84);
nor NOR2 (N86, N23, N5);
and AND2 (N87, N83, N27);
xor XOR2 (N88, N66, N71);
or OR2 (N89, N85, N8);
not NOT1 (N90, N67);
nand NAND4 (N91, N78, N89, N23, N25);
and AND4 (N92, N28, N70, N69, N1);
nor NOR4 (N93, N88, N5, N59, N67);
nor NOR4 (N94, N81, N26, N37, N27);
xor XOR2 (N95, N92, N8);
and AND4 (N96, N82, N47, N90, N41);
buf BUF1 (N97, N54);
xor XOR2 (N98, N86, N45);
nand NAND2 (N99, N93, N95);
nor NOR4 (N100, N35, N76, N27, N19);
and AND3 (N101, N94, N89, N56);
not NOT1 (N102, N87);
and AND4 (N103, N91, N62, N71, N50);
xor XOR2 (N104, N97, N94);
buf BUF1 (N105, N96);
nor NOR3 (N106, N104, N90, N70);
buf BUF1 (N107, N103);
and AND2 (N108, N100, N47);
and AND3 (N109, N101, N46, N73);
nand NAND3 (N110, N105, N106, N75);
nand NAND4 (N111, N24, N30, N17, N39);
nand NAND3 (N112, N22, N71, N30);
buf BUF1 (N113, N107);
or OR3 (N114, N98, N32, N27);
nand NAND3 (N115, N80, N63, N60);
nor NOR2 (N116, N114, N77);
not NOT1 (N117, N112);
or OR2 (N118, N115, N32);
and AND2 (N119, N111, N68);
buf BUF1 (N120, N118);
buf BUF1 (N121, N99);
nor NOR3 (N122, N109, N66, N45);
and AND3 (N123, N110, N87, N72);
buf BUF1 (N124, N116);
or OR4 (N125, N113, N56, N92, N8);
xor XOR2 (N126, N124, N76);
xor XOR2 (N127, N125, N60);
nor NOR4 (N128, N120, N59, N48, N23);
not NOT1 (N129, N108);
not NOT1 (N130, N121);
xor XOR2 (N131, N127, N70);
or OR4 (N132, N131, N49, N44, N108);
buf BUF1 (N133, N128);
nand NAND3 (N134, N122, N26, N63);
or OR3 (N135, N123, N9, N13);
or OR4 (N136, N129, N28, N57, N14);
xor XOR2 (N137, N132, N103);
nor NOR3 (N138, N130, N108, N110);
or OR4 (N139, N136, N102, N26, N135);
buf BUF1 (N140, N39);
and AND4 (N141, N86, N59, N93, N121);
or OR2 (N142, N137, N12);
not NOT1 (N143, N126);
nor NOR3 (N144, N139, N139, N64);
and AND2 (N145, N143, N102);
nand NAND3 (N146, N117, N64, N138);
nand NAND2 (N147, N87, N41);
and AND4 (N148, N140, N4, N47, N37);
not NOT1 (N149, N144);
xor XOR2 (N150, N146, N87);
nand NAND4 (N151, N150, N18, N15, N99);
nand NAND2 (N152, N141, N49);
or OR3 (N153, N149, N94, N17);
nor NOR4 (N154, N145, N132, N10, N90);
not NOT1 (N155, N133);
xor XOR2 (N156, N153, N49);
nand NAND3 (N157, N147, N45, N8);
not NOT1 (N158, N119);
or OR4 (N159, N152, N125, N1, N19);
buf BUF1 (N160, N159);
and AND3 (N161, N154, N10, N48);
and AND3 (N162, N142, N16, N29);
nor NOR4 (N163, N162, N127, N137, N22);
xor XOR2 (N164, N134, N159);
and AND4 (N165, N158, N119, N23, N18);
not NOT1 (N166, N151);
xor XOR2 (N167, N156, N74);
xor XOR2 (N168, N164, N5);
not NOT1 (N169, N166);
buf BUF1 (N170, N165);
nor NOR2 (N171, N170, N143);
buf BUF1 (N172, N167);
nor NOR4 (N173, N168, N36, N96, N9);
and AND2 (N174, N163, N30);
nor NOR2 (N175, N148, N107);
xor XOR2 (N176, N161, N74);
buf BUF1 (N177, N173);
not NOT1 (N178, N157);
buf BUF1 (N179, N155);
xor XOR2 (N180, N175, N143);
or OR2 (N181, N180, N111);
or OR3 (N182, N160, N82, N26);
nand NAND3 (N183, N172, N15, N121);
or OR2 (N184, N179, N116);
or OR2 (N185, N176, N112);
not NOT1 (N186, N184);
or OR3 (N187, N178, N97, N149);
or OR3 (N188, N185, N158, N96);
nand NAND4 (N189, N174, N89, N6, N113);
not NOT1 (N190, N182);
not NOT1 (N191, N177);
and AND4 (N192, N186, N157, N22, N64);
nor NOR4 (N193, N169, N173, N55, N58);
nor NOR4 (N194, N190, N84, N12, N9);
not NOT1 (N195, N192);
nor NOR4 (N196, N191, N98, N186, N64);
buf BUF1 (N197, N189);
or OR4 (N198, N187, N109, N38, N124);
and AND3 (N199, N193, N127, N26);
buf BUF1 (N200, N181);
nor NOR3 (N201, N198, N121, N12);
nand NAND3 (N202, N195, N65, N39);
and AND4 (N203, N194, N12, N56, N112);
xor XOR2 (N204, N199, N177);
not NOT1 (N205, N188);
not NOT1 (N206, N204);
buf BUF1 (N207, N196);
nand NAND4 (N208, N207, N52, N57, N164);
buf BUF1 (N209, N202);
or OR3 (N210, N208, N182, N28);
xor XOR2 (N211, N206, N76);
or OR3 (N212, N183, N14, N95);
not NOT1 (N213, N200);
not NOT1 (N214, N210);
xor XOR2 (N215, N212, N40);
xor XOR2 (N216, N201, N71);
nand NAND2 (N217, N214, N120);
nand NAND2 (N218, N197, N92);
nor NOR3 (N219, N205, N136, N94);
and AND2 (N220, N211, N24);
nand NAND4 (N221, N209, N217, N71, N181);
xor XOR2 (N222, N81, N82);
xor XOR2 (N223, N222, N208);
nand NAND3 (N224, N213, N1, N83);
nor NOR4 (N225, N223, N121, N168, N104);
nor NOR3 (N226, N203, N118, N127);
nand NAND2 (N227, N171, N185);
and AND3 (N228, N218, N175, N91);
buf BUF1 (N229, N228);
buf BUF1 (N230, N221);
xor XOR2 (N231, N226, N6);
buf BUF1 (N232, N231);
xor XOR2 (N233, N225, N159);
nor NOR3 (N234, N233, N27, N53);
nand NAND2 (N235, N234, N41);
and AND3 (N236, N232, N114, N228);
buf BUF1 (N237, N219);
or OR3 (N238, N230, N198, N5);
buf BUF1 (N239, N224);
not NOT1 (N240, N220);
or OR4 (N241, N235, N147, N85, N151);
nand NAND4 (N242, N238, N78, N42, N57);
nor NOR4 (N243, N239, N57, N125, N122);
nor NOR4 (N244, N236, N156, N182, N243);
nor NOR3 (N245, N221, N126, N147);
and AND2 (N246, N244, N228);
nand NAND4 (N247, N216, N139, N84, N193);
xor XOR2 (N248, N227, N112);
and AND2 (N249, N241, N100);
xor XOR2 (N250, N247, N33);
nand NAND3 (N251, N242, N233, N96);
buf BUF1 (N252, N249);
and AND3 (N253, N251, N31, N224);
not NOT1 (N254, N229);
nor NOR4 (N255, N253, N211, N84, N218);
buf BUF1 (N256, N248);
nor NOR3 (N257, N255, N43, N223);
not NOT1 (N258, N240);
nor NOR3 (N259, N246, N197, N80);
buf BUF1 (N260, N256);
buf BUF1 (N261, N245);
nor NOR2 (N262, N258, N56);
xor XOR2 (N263, N215, N46);
or OR4 (N264, N237, N35, N230, N263);
not NOT1 (N265, N82);
or OR3 (N266, N264, N151, N65);
nor NOR2 (N267, N262, N100);
buf BUF1 (N268, N265);
nand NAND2 (N269, N259, N249);
and AND3 (N270, N269, N213, N159);
buf BUF1 (N271, N250);
or OR2 (N272, N252, N133);
or OR2 (N273, N254, N106);
and AND2 (N274, N257, N240);
xor XOR2 (N275, N261, N19);
and AND2 (N276, N267, N132);
or OR4 (N277, N266, N133, N202, N142);
not NOT1 (N278, N271);
or OR4 (N279, N272, N48, N230, N93);
or OR4 (N280, N279, N188, N117, N273);
nor NOR3 (N281, N7, N260, N220);
buf BUF1 (N282, N245);
and AND4 (N283, N270, N269, N198, N48);
or OR4 (N284, N277, N121, N28, N34);
nand NAND3 (N285, N274, N27, N128);
not NOT1 (N286, N275);
and AND4 (N287, N280, N240, N275, N3);
or OR3 (N288, N286, N29, N179);
buf BUF1 (N289, N285);
and AND3 (N290, N278, N150, N71);
and AND2 (N291, N284, N286);
or OR4 (N292, N287, N48, N153, N196);
or OR3 (N293, N288, N183, N201);
and AND4 (N294, N289, N193, N125, N55);
and AND2 (N295, N294, N286);
and AND3 (N296, N283, N162, N119);
not NOT1 (N297, N290);
not NOT1 (N298, N297);
buf BUF1 (N299, N295);
not NOT1 (N300, N268);
and AND4 (N301, N299, N185, N88, N211);
xor XOR2 (N302, N281, N90);
nand NAND2 (N303, N296, N83);
not NOT1 (N304, N276);
not NOT1 (N305, N304);
xor XOR2 (N306, N291, N288);
or OR3 (N307, N292, N30, N154);
nor NOR4 (N308, N300, N224, N59, N55);
and AND3 (N309, N307, N222, N29);
not NOT1 (N310, N298);
xor XOR2 (N311, N308, N52);
not NOT1 (N312, N306);
endmodule