// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11;

output N3503,N3509,N3495,N3501,N3508,N3493,N3504,N3510,N3492,N3511;

nand NAND4 (N12, N7, N5, N5, N1);
nand NAND4 (N13, N8, N11, N1, N1);
nor NOR2 (N14, N7, N7);
nor NOR3 (N15, N10, N7, N14);
buf BUF1 (N16, N1);
nor NOR2 (N17, N3, N2);
or OR3 (N18, N2, N16, N14);
xor XOR2 (N19, N15, N14);
or OR2 (N20, N9, N19);
xor XOR2 (N21, N16, N20);
nand NAND2 (N22, N9, N16);
not NOT1 (N23, N1);
or OR4 (N24, N7, N10, N3, N18);
xor XOR2 (N25, N19, N4);
or OR2 (N26, N6, N18);
nor NOR3 (N27, N22, N2, N6);
and AND4 (N28, N26, N27, N22, N20);
not NOT1 (N29, N21);
nand NAND4 (N30, N22, N26, N12, N9);
buf BUF1 (N31, N6);
nor NOR2 (N32, N27, N16);
not NOT1 (N33, N13);
xor XOR2 (N34, N25, N23);
or OR4 (N35, N12, N14, N27, N18);
or OR3 (N36, N31, N3, N17);
buf BUF1 (N37, N20);
xor XOR2 (N38, N28, N6);
nor NOR2 (N39, N37, N16);
and AND4 (N40, N39, N3, N11, N30);
buf BUF1 (N41, N10);
and AND4 (N42, N29, N6, N21, N26);
not NOT1 (N43, N41);
or OR4 (N44, N40, N28, N19, N35);
nor NOR4 (N45, N31, N44, N43, N7);
or OR2 (N46, N42, N14);
not NOT1 (N47, N6);
and AND4 (N48, N18, N1, N25, N4);
buf BUF1 (N49, N48);
or OR2 (N50, N38, N21);
buf BUF1 (N51, N33);
xor XOR2 (N52, N50, N51);
xor XOR2 (N53, N8, N10);
buf BUF1 (N54, N46);
nor NOR4 (N55, N34, N19, N47, N10);
xor XOR2 (N56, N31, N2);
nand NAND3 (N57, N36, N4, N46);
not NOT1 (N58, N57);
xor XOR2 (N59, N45, N54);
nor NOR4 (N60, N6, N31, N46, N19);
and AND3 (N61, N59, N52, N8);
xor XOR2 (N62, N52, N31);
and AND2 (N63, N55, N24);
nand NAND4 (N64, N62, N35, N7, N19);
or OR2 (N65, N52, N19);
and AND3 (N66, N61, N4, N40);
and AND4 (N67, N64, N19, N46, N48);
nand NAND3 (N68, N58, N51, N8);
nand NAND2 (N69, N65, N8);
and AND4 (N70, N60, N18, N31, N7);
not NOT1 (N71, N56);
buf BUF1 (N72, N53);
or OR4 (N73, N66, N5, N37, N43);
not NOT1 (N74, N49);
buf BUF1 (N75, N32);
not NOT1 (N76, N75);
buf BUF1 (N77, N73);
or OR2 (N78, N69, N72);
nor NOR4 (N79, N46, N60, N17, N67);
buf BUF1 (N80, N65);
xor XOR2 (N81, N74, N53);
nand NAND3 (N82, N63, N36, N60);
or OR4 (N83, N78, N74, N72, N54);
or OR2 (N84, N77, N35);
or OR4 (N85, N83, N48, N38, N74);
buf BUF1 (N86, N82);
or OR3 (N87, N85, N53, N24);
xor XOR2 (N88, N71, N79);
and AND3 (N89, N23, N85, N55);
not NOT1 (N90, N87);
xor XOR2 (N91, N89, N73);
buf BUF1 (N92, N88);
xor XOR2 (N93, N80, N33);
buf BUF1 (N94, N84);
and AND3 (N95, N68, N31, N6);
or OR2 (N96, N70, N80);
buf BUF1 (N97, N76);
buf BUF1 (N98, N97);
and AND2 (N99, N86, N60);
buf BUF1 (N100, N93);
nor NOR2 (N101, N98, N15);
or OR4 (N102, N94, N12, N61, N69);
not NOT1 (N103, N102);
or OR4 (N104, N81, N11, N54, N36);
and AND2 (N105, N91, N53);
xor XOR2 (N106, N104, N5);
not NOT1 (N107, N90);
nand NAND4 (N108, N103, N107, N63, N10);
nand NAND3 (N109, N14, N90, N8);
not NOT1 (N110, N100);
nand NAND2 (N111, N96, N24);
xor XOR2 (N112, N110, N103);
nand NAND2 (N113, N108, N66);
xor XOR2 (N114, N99, N30);
or OR2 (N115, N112, N110);
xor XOR2 (N116, N114, N50);
or OR2 (N117, N95, N70);
or OR2 (N118, N105, N43);
nand NAND3 (N119, N116, N115, N69);
not NOT1 (N120, N5);
and AND4 (N121, N92, N37, N45, N87);
xor XOR2 (N122, N101, N62);
nand NAND2 (N123, N122, N98);
or OR4 (N124, N121, N25, N34, N2);
nor NOR3 (N125, N124, N27, N66);
not NOT1 (N126, N123);
nand NAND2 (N127, N120, N121);
nor NOR3 (N128, N119, N47, N42);
xor XOR2 (N129, N113, N32);
xor XOR2 (N130, N125, N28);
xor XOR2 (N131, N109, N76);
not NOT1 (N132, N118);
xor XOR2 (N133, N130, N93);
buf BUF1 (N134, N132);
not NOT1 (N135, N134);
nor NOR4 (N136, N111, N10, N68, N102);
or OR3 (N137, N129, N16, N131);
buf BUF1 (N138, N105);
buf BUF1 (N139, N126);
and AND3 (N140, N106, N132, N89);
nor NOR2 (N141, N136, N93);
and AND2 (N142, N127, N81);
and AND3 (N143, N142, N139, N86);
nand NAND2 (N144, N31, N53);
or OR2 (N145, N128, N111);
and AND3 (N146, N143, N73, N133);
buf BUF1 (N147, N127);
nor NOR4 (N148, N146, N56, N114, N122);
buf BUF1 (N149, N117);
not NOT1 (N150, N148);
and AND4 (N151, N145, N145, N68, N150);
nand NAND4 (N152, N50, N8, N146, N59);
nor NOR3 (N153, N152, N81, N48);
nor NOR4 (N154, N153, N121, N78, N61);
nor NOR3 (N155, N147, N105, N28);
nand NAND4 (N156, N149, N130, N75, N138);
xor XOR2 (N157, N48, N99);
xor XOR2 (N158, N156, N8);
nor NOR3 (N159, N137, N102, N145);
buf BUF1 (N160, N157);
buf BUF1 (N161, N159);
xor XOR2 (N162, N144, N57);
buf BUF1 (N163, N140);
nand NAND4 (N164, N158, N79, N159, N108);
nor NOR3 (N165, N154, N46, N39);
nand NAND4 (N166, N160, N31, N29, N18);
nand NAND4 (N167, N141, N85, N166, N31);
nor NOR4 (N168, N16, N60, N62, N75);
buf BUF1 (N169, N155);
and AND2 (N170, N165, N7);
or OR2 (N171, N151, N70);
not NOT1 (N172, N170);
not NOT1 (N173, N171);
or OR2 (N174, N173, N82);
not NOT1 (N175, N174);
not NOT1 (N176, N135);
nand NAND4 (N177, N161, N136, N24, N165);
xor XOR2 (N178, N167, N87);
or OR4 (N179, N168, N13, N130, N97);
nand NAND4 (N180, N163, N7, N83, N58);
not NOT1 (N181, N175);
buf BUF1 (N182, N176);
xor XOR2 (N183, N177, N156);
nand NAND4 (N184, N182, N78, N181, N108);
buf BUF1 (N185, N13);
buf BUF1 (N186, N184);
nand NAND2 (N187, N186, N79);
nand NAND2 (N188, N178, N157);
nor NOR3 (N189, N179, N36, N79);
and AND3 (N190, N188, N37, N173);
or OR2 (N191, N172, N52);
not NOT1 (N192, N189);
xor XOR2 (N193, N190, N91);
or OR2 (N194, N191, N98);
nor NOR2 (N195, N183, N129);
xor XOR2 (N196, N187, N47);
not NOT1 (N197, N195);
not NOT1 (N198, N185);
xor XOR2 (N199, N180, N37);
nand NAND4 (N200, N199, N97, N90, N26);
nand NAND4 (N201, N162, N71, N44, N127);
or OR3 (N202, N197, N40, N150);
and AND4 (N203, N196, N118, N178, N81);
xor XOR2 (N204, N201, N89);
or OR4 (N205, N192, N189, N15, N92);
and AND3 (N206, N204, N140, N81);
and AND4 (N207, N205, N191, N172, N98);
or OR2 (N208, N164, N103);
buf BUF1 (N209, N207);
or OR4 (N210, N200, N190, N82, N113);
or OR4 (N211, N193, N14, N91, N170);
or OR4 (N212, N208, N106, N106, N153);
nand NAND2 (N213, N203, N204);
and AND4 (N214, N202, N110, N209, N184);
and AND3 (N215, N185, N124, N176);
nor NOR2 (N216, N206, N107);
and AND4 (N217, N211, N26, N114, N134);
nand NAND2 (N218, N214, N78);
or OR2 (N219, N218, N193);
nor NOR2 (N220, N198, N2);
nand NAND3 (N221, N219, N197, N176);
not NOT1 (N222, N215);
or OR4 (N223, N213, N221, N169, N92);
buf BUF1 (N224, N169);
or OR4 (N225, N5, N169, N135, N170);
nor NOR3 (N226, N212, N166, N96);
buf BUF1 (N227, N226);
not NOT1 (N228, N194);
xor XOR2 (N229, N227, N21);
nor NOR4 (N230, N216, N169, N57, N60);
nor NOR3 (N231, N217, N207, N63);
not NOT1 (N232, N210);
nor NOR4 (N233, N232, N117, N54, N15);
xor XOR2 (N234, N233, N214);
and AND3 (N235, N225, N81, N66);
and AND2 (N236, N220, N234);
nand NAND2 (N237, N189, N34);
not NOT1 (N238, N228);
buf BUF1 (N239, N236);
buf BUF1 (N240, N238);
not NOT1 (N241, N237);
or OR3 (N242, N229, N161, N113);
buf BUF1 (N243, N242);
nand NAND2 (N244, N241, N204);
buf BUF1 (N245, N224);
nor NOR2 (N246, N230, N81);
nor NOR2 (N247, N243, N227);
or OR4 (N248, N222, N204, N175, N65);
xor XOR2 (N249, N245, N111);
nor NOR2 (N250, N249, N48);
nand NAND3 (N251, N235, N10, N102);
xor XOR2 (N252, N244, N195);
nor NOR2 (N253, N248, N221);
buf BUF1 (N254, N240);
not NOT1 (N255, N250);
xor XOR2 (N256, N223, N5);
buf BUF1 (N257, N254);
nand NAND3 (N258, N253, N208, N43);
xor XOR2 (N259, N252, N177);
not NOT1 (N260, N239);
nor NOR3 (N261, N247, N64, N136);
buf BUF1 (N262, N231);
and AND4 (N263, N258, N13, N136, N218);
or OR4 (N264, N246, N123, N154, N33);
nand NAND3 (N265, N256, N228, N263);
xor XOR2 (N266, N58, N237);
not NOT1 (N267, N260);
or OR2 (N268, N265, N211);
and AND4 (N269, N266, N48, N4, N237);
nor NOR4 (N270, N255, N255, N181, N89);
and AND2 (N271, N259, N179);
not NOT1 (N272, N267);
buf BUF1 (N273, N270);
or OR4 (N274, N264, N177, N37, N249);
not NOT1 (N275, N261);
xor XOR2 (N276, N274, N247);
or OR4 (N277, N275, N185, N243, N4);
buf BUF1 (N278, N272);
xor XOR2 (N279, N277, N39);
and AND2 (N280, N279, N145);
or OR3 (N281, N280, N136, N255);
xor XOR2 (N282, N257, N72);
buf BUF1 (N283, N262);
nor NOR3 (N284, N269, N77, N238);
buf BUF1 (N285, N273);
or OR4 (N286, N281, N194, N170, N129);
nor NOR4 (N287, N285, N149, N163, N69);
buf BUF1 (N288, N282);
and AND2 (N289, N276, N159);
and AND3 (N290, N289, N114, N75);
not NOT1 (N291, N288);
and AND3 (N292, N278, N134, N178);
xor XOR2 (N293, N286, N124);
not NOT1 (N294, N251);
nor NOR4 (N295, N268, N127, N203, N8);
not NOT1 (N296, N291);
not NOT1 (N297, N294);
not NOT1 (N298, N287);
not NOT1 (N299, N295);
nor NOR3 (N300, N297, N90, N210);
nand NAND4 (N301, N284, N188, N142, N294);
nand NAND2 (N302, N298, N217);
buf BUF1 (N303, N299);
or OR2 (N304, N283, N83);
xor XOR2 (N305, N303, N187);
nor NOR2 (N306, N292, N240);
nor NOR2 (N307, N301, N9);
not NOT1 (N308, N293);
and AND2 (N309, N304, N307);
and AND4 (N310, N265, N305, N302, N151);
and AND3 (N311, N7, N204, N75);
nand NAND4 (N312, N14, N181, N261, N31);
nor NOR3 (N313, N271, N301, N173);
or OR3 (N314, N300, N242, N15);
or OR3 (N315, N306, N15, N141);
not NOT1 (N316, N312);
nand NAND2 (N317, N315, N264);
buf BUF1 (N318, N311);
buf BUF1 (N319, N314);
xor XOR2 (N320, N309, N165);
nor NOR3 (N321, N320, N160, N42);
nor NOR3 (N322, N321, N71, N315);
nor NOR4 (N323, N313, N181, N72, N126);
xor XOR2 (N324, N290, N269);
xor XOR2 (N325, N319, N3);
and AND4 (N326, N318, N105, N23, N267);
nor NOR2 (N327, N317, N196);
nand NAND4 (N328, N310, N78, N243, N294);
nand NAND4 (N329, N308, N309, N62, N149);
nand NAND3 (N330, N325, N70, N246);
and AND2 (N331, N328, N323);
nand NAND4 (N332, N314, N231, N287, N154);
or OR2 (N333, N296, N126);
and AND3 (N334, N333, N91, N178);
nor NOR2 (N335, N327, N21);
nand NAND4 (N336, N324, N273, N229, N167);
nor NOR2 (N337, N322, N249);
buf BUF1 (N338, N330);
not NOT1 (N339, N336);
or OR4 (N340, N339, N274, N161, N47);
and AND4 (N341, N329, N72, N87, N305);
and AND3 (N342, N334, N93, N245);
nor NOR3 (N343, N331, N303, N190);
not NOT1 (N344, N341);
not NOT1 (N345, N340);
nor NOR2 (N346, N316, N23);
xor XOR2 (N347, N332, N346);
or OR2 (N348, N332, N160);
nor NOR4 (N349, N347, N1, N280, N196);
and AND4 (N350, N342, N31, N123, N198);
not NOT1 (N351, N350);
or OR4 (N352, N349, N127, N195, N265);
not NOT1 (N353, N326);
nor NOR2 (N354, N338, N123);
xor XOR2 (N355, N343, N26);
xor XOR2 (N356, N353, N184);
nand NAND3 (N357, N354, N243, N292);
buf BUF1 (N358, N352);
nor NOR3 (N359, N348, N180, N269);
nor NOR2 (N360, N356, N195);
buf BUF1 (N361, N359);
and AND3 (N362, N357, N5, N128);
xor XOR2 (N363, N360, N236);
or OR3 (N364, N351, N346, N227);
xor XOR2 (N365, N363, N285);
nor NOR3 (N366, N345, N209, N77);
nor NOR2 (N367, N337, N277);
not NOT1 (N368, N364);
nor NOR3 (N369, N362, N352, N292);
xor XOR2 (N370, N358, N253);
not NOT1 (N371, N367);
buf BUF1 (N372, N365);
not NOT1 (N373, N370);
and AND4 (N374, N366, N69, N72, N151);
or OR2 (N375, N355, N236);
and AND4 (N376, N375, N57, N308, N239);
or OR3 (N377, N376, N172, N12);
not NOT1 (N378, N372);
nand NAND2 (N379, N377, N6);
and AND2 (N380, N379, N235);
not NOT1 (N381, N373);
not NOT1 (N382, N380);
nand NAND4 (N383, N374, N92, N230, N249);
not NOT1 (N384, N344);
nand NAND3 (N385, N378, N167, N198);
and AND4 (N386, N361, N282, N32, N13);
buf BUF1 (N387, N371);
buf BUF1 (N388, N384);
not NOT1 (N389, N387);
buf BUF1 (N390, N388);
not NOT1 (N391, N383);
or OR2 (N392, N381, N216);
buf BUF1 (N393, N385);
buf BUF1 (N394, N369);
nor NOR4 (N395, N389, N265, N329, N304);
and AND4 (N396, N368, N377, N282, N237);
xor XOR2 (N397, N395, N260);
nand NAND2 (N398, N390, N83);
nor NOR2 (N399, N382, N118);
or OR4 (N400, N391, N197, N339, N115);
or OR2 (N401, N397, N375);
nor NOR4 (N402, N386, N351, N241, N89);
xor XOR2 (N403, N392, N78);
xor XOR2 (N404, N394, N217);
not NOT1 (N405, N403);
nor NOR3 (N406, N335, N214, N103);
buf BUF1 (N407, N401);
xor XOR2 (N408, N399, N126);
nor NOR3 (N409, N408, N9, N282);
xor XOR2 (N410, N400, N393);
or OR4 (N411, N128, N84, N23, N116);
nand NAND2 (N412, N406, N198);
nand NAND4 (N413, N409, N316, N307, N372);
not NOT1 (N414, N396);
nand NAND3 (N415, N413, N339, N93);
xor XOR2 (N416, N404, N292);
nand NAND2 (N417, N405, N25);
nor NOR4 (N418, N414, N215, N122, N397);
xor XOR2 (N419, N402, N374);
nand NAND4 (N420, N419, N84, N315, N358);
and AND4 (N421, N417, N238, N133, N280);
and AND2 (N422, N412, N313);
nand NAND2 (N423, N422, N177);
nand NAND2 (N424, N410, N250);
xor XOR2 (N425, N415, N356);
or OR3 (N426, N416, N355, N413);
nand NAND3 (N427, N420, N383, N147);
and AND2 (N428, N424, N37);
nor NOR2 (N429, N426, N53);
xor XOR2 (N430, N411, N173);
xor XOR2 (N431, N398, N304);
nand NAND3 (N432, N428, N160, N300);
buf BUF1 (N433, N418);
nor NOR4 (N434, N423, N33, N294, N354);
nor NOR4 (N435, N431, N395, N242, N155);
xor XOR2 (N436, N433, N108);
nor NOR2 (N437, N435, N106);
or OR2 (N438, N421, N430);
xor XOR2 (N439, N104, N140);
not NOT1 (N440, N427);
not NOT1 (N441, N440);
buf BUF1 (N442, N429);
not NOT1 (N443, N438);
nor NOR3 (N444, N443, N47, N350);
or OR3 (N445, N442, N125, N11);
or OR2 (N446, N432, N287);
and AND2 (N447, N441, N437);
xor XOR2 (N448, N192, N447);
buf BUF1 (N449, N337);
xor XOR2 (N450, N445, N144);
and AND2 (N451, N407, N434);
xor XOR2 (N452, N40, N129);
nor NOR4 (N453, N436, N276, N278, N360);
or OR2 (N454, N446, N207);
xor XOR2 (N455, N425, N251);
or OR4 (N456, N452, N375, N364, N453);
and AND4 (N457, N35, N6, N299, N353);
or OR3 (N458, N454, N211, N197);
xor XOR2 (N459, N456, N53);
xor XOR2 (N460, N449, N353);
and AND3 (N461, N450, N337, N394);
and AND3 (N462, N461, N238, N136);
or OR4 (N463, N460, N12, N92, N396);
or OR2 (N464, N462, N405);
not NOT1 (N465, N455);
nor NOR4 (N466, N465, N387, N257, N385);
buf BUF1 (N467, N464);
not NOT1 (N468, N448);
and AND2 (N469, N467, N221);
nand NAND3 (N470, N468, N193, N117);
and AND4 (N471, N444, N32, N143, N380);
or OR4 (N472, N470, N468, N199, N285);
not NOT1 (N473, N469);
xor XOR2 (N474, N473, N394);
nand NAND2 (N475, N457, N458);
nand NAND3 (N476, N38, N193, N200);
nor NOR2 (N477, N466, N475);
not NOT1 (N478, N11);
or OR2 (N479, N474, N450);
and AND3 (N480, N463, N18, N24);
and AND3 (N481, N471, N188, N141);
or OR2 (N482, N451, N142);
and AND4 (N483, N479, N91, N58, N418);
xor XOR2 (N484, N439, N309);
not NOT1 (N485, N476);
nand NAND4 (N486, N481, N454, N414, N179);
and AND2 (N487, N486, N468);
and AND3 (N488, N485, N275, N300);
not NOT1 (N489, N477);
and AND3 (N490, N488, N324, N367);
buf BUF1 (N491, N472);
and AND3 (N492, N478, N490, N187);
not NOT1 (N493, N163);
nor NOR4 (N494, N482, N170, N229, N386);
nand NAND3 (N495, N492, N116, N177);
not NOT1 (N496, N493);
nand NAND3 (N497, N484, N346, N326);
buf BUF1 (N498, N489);
nand NAND4 (N499, N487, N8, N32, N187);
or OR2 (N500, N494, N67);
nand NAND4 (N501, N496, N160, N15, N408);
xor XOR2 (N502, N500, N140);
or OR3 (N503, N501, N202, N460);
nor NOR2 (N504, N495, N209);
nand NAND3 (N505, N483, N415, N297);
xor XOR2 (N506, N497, N264);
nand NAND3 (N507, N480, N180, N30);
buf BUF1 (N508, N498);
not NOT1 (N509, N459);
and AND2 (N510, N504, N145);
and AND4 (N511, N502, N70, N64, N85);
nand NAND4 (N512, N503, N308, N207, N185);
or OR2 (N513, N511, N167);
xor XOR2 (N514, N505, N113);
or OR3 (N515, N514, N243, N393);
and AND3 (N516, N506, N309, N189);
and AND2 (N517, N499, N159);
buf BUF1 (N518, N513);
nand NAND2 (N519, N518, N51);
nor NOR2 (N520, N510, N155);
buf BUF1 (N521, N515);
xor XOR2 (N522, N512, N378);
buf BUF1 (N523, N508);
nand NAND2 (N524, N522, N63);
nor NOR4 (N525, N520, N280, N174, N268);
or OR3 (N526, N516, N391, N442);
buf BUF1 (N527, N509);
or OR4 (N528, N524, N13, N280, N266);
nor NOR4 (N529, N526, N366, N393, N319);
xor XOR2 (N530, N527, N182);
nand NAND3 (N531, N507, N395, N316);
nor NOR3 (N532, N531, N105, N501);
and AND2 (N533, N529, N255);
buf BUF1 (N534, N525);
nor NOR3 (N535, N523, N123, N146);
nor NOR4 (N536, N533, N293, N330, N328);
or OR3 (N537, N535, N325, N380);
nand NAND3 (N538, N528, N40, N22);
and AND2 (N539, N532, N251);
not NOT1 (N540, N536);
not NOT1 (N541, N517);
not NOT1 (N542, N521);
not NOT1 (N543, N539);
nor NOR3 (N544, N543, N165, N128);
nand NAND3 (N545, N519, N146, N453);
buf BUF1 (N546, N538);
and AND4 (N547, N540, N435, N449, N476);
nand NAND3 (N548, N547, N491, N49);
and AND3 (N549, N113, N291, N401);
xor XOR2 (N550, N548, N517);
and AND2 (N551, N550, N108);
buf BUF1 (N552, N544);
nand NAND2 (N553, N546, N8);
nand NAND2 (N554, N534, N44);
and AND4 (N555, N549, N136, N536, N367);
buf BUF1 (N556, N554);
xor XOR2 (N557, N541, N523);
not NOT1 (N558, N530);
and AND4 (N559, N542, N184, N359, N541);
or OR3 (N560, N556, N392, N98);
buf BUF1 (N561, N555);
xor XOR2 (N562, N557, N21);
or OR3 (N563, N545, N440, N495);
nand NAND4 (N564, N560, N83, N470, N178);
not NOT1 (N565, N551);
buf BUF1 (N566, N553);
and AND4 (N567, N562, N250, N394, N192);
and AND2 (N568, N564, N215);
or OR4 (N569, N568, N250, N317, N427);
nor NOR3 (N570, N537, N122, N386);
nor NOR2 (N571, N552, N131);
nor NOR4 (N572, N570, N501, N496, N165);
not NOT1 (N573, N563);
nor NOR3 (N574, N567, N356, N508);
nand NAND4 (N575, N565, N85, N398, N116);
nor NOR3 (N576, N571, N460, N105);
nand NAND3 (N577, N558, N163, N294);
xor XOR2 (N578, N573, N549);
nor NOR4 (N579, N578, N262, N274, N298);
nand NAND4 (N580, N566, N476, N507, N133);
or OR4 (N581, N575, N426, N536, N226);
nand NAND4 (N582, N581, N246, N514, N32);
not NOT1 (N583, N580);
buf BUF1 (N584, N574);
or OR4 (N585, N579, N417, N271, N174);
buf BUF1 (N586, N559);
not NOT1 (N587, N585);
not NOT1 (N588, N572);
nand NAND2 (N589, N582, N36);
buf BUF1 (N590, N576);
xor XOR2 (N591, N589, N157);
or OR4 (N592, N590, N527, N37, N72);
buf BUF1 (N593, N577);
and AND4 (N594, N569, N155, N181, N16);
nand NAND3 (N595, N593, N106, N231);
or OR4 (N596, N592, N510, N176, N129);
and AND3 (N597, N586, N320, N196);
nand NAND2 (N598, N588, N501);
or OR2 (N599, N596, N400);
buf BUF1 (N600, N583);
not NOT1 (N601, N598);
nand NAND3 (N602, N591, N492, N115);
nor NOR2 (N603, N600, N493);
buf BUF1 (N604, N584);
xor XOR2 (N605, N561, N373);
buf BUF1 (N606, N603);
or OR4 (N607, N606, N556, N133, N302);
and AND2 (N608, N594, N451);
not NOT1 (N609, N605);
nor NOR3 (N610, N597, N54, N554);
and AND3 (N611, N595, N350, N558);
buf BUF1 (N612, N607);
buf BUF1 (N613, N610);
and AND2 (N614, N608, N412);
and AND2 (N615, N604, N53);
nand NAND3 (N616, N587, N11, N479);
or OR3 (N617, N611, N275, N500);
nand NAND2 (N618, N616, N124);
nand NAND2 (N619, N599, N606);
not NOT1 (N620, N609);
nor NOR4 (N621, N613, N86, N612, N211);
not NOT1 (N622, N494);
nand NAND3 (N623, N601, N108, N552);
buf BUF1 (N624, N617);
not NOT1 (N625, N614);
not NOT1 (N626, N620);
buf BUF1 (N627, N623);
buf BUF1 (N628, N619);
nor NOR4 (N629, N626, N343, N266, N152);
buf BUF1 (N630, N624);
buf BUF1 (N631, N621);
not NOT1 (N632, N602);
not NOT1 (N633, N628);
nand NAND2 (N634, N618, N92);
buf BUF1 (N635, N631);
not NOT1 (N636, N629);
buf BUF1 (N637, N632);
or OR2 (N638, N633, N148);
xor XOR2 (N639, N622, N102);
not NOT1 (N640, N639);
or OR2 (N641, N630, N495);
buf BUF1 (N642, N637);
or OR2 (N643, N615, N538);
or OR3 (N644, N634, N194, N611);
or OR2 (N645, N640, N156);
xor XOR2 (N646, N625, N296);
nor NOR3 (N647, N643, N585, N219);
and AND2 (N648, N638, N611);
or OR3 (N649, N635, N252, N405);
and AND2 (N650, N646, N63);
buf BUF1 (N651, N648);
not NOT1 (N652, N650);
not NOT1 (N653, N641);
buf BUF1 (N654, N642);
or OR2 (N655, N627, N160);
not NOT1 (N656, N645);
and AND3 (N657, N636, N185, N45);
and AND2 (N658, N657, N398);
xor XOR2 (N659, N654, N275);
or OR2 (N660, N658, N658);
and AND3 (N661, N649, N652, N642);
nor NOR4 (N662, N307, N300, N555, N583);
or OR2 (N663, N647, N435);
nand NAND2 (N664, N661, N459);
buf BUF1 (N665, N664);
and AND3 (N666, N651, N204, N519);
buf BUF1 (N667, N655);
and AND2 (N668, N665, N125);
nand NAND3 (N669, N653, N152, N643);
or OR2 (N670, N659, N642);
xor XOR2 (N671, N666, N125);
buf BUF1 (N672, N662);
or OR2 (N673, N656, N233);
and AND4 (N674, N667, N351, N99, N523);
buf BUF1 (N675, N670);
nand NAND2 (N676, N644, N661);
nand NAND4 (N677, N672, N638, N548, N445);
buf BUF1 (N678, N660);
nor NOR3 (N679, N677, N219, N421);
nor NOR2 (N680, N673, N436);
or OR4 (N681, N679, N366, N493, N197);
and AND4 (N682, N668, N137, N452, N444);
nor NOR2 (N683, N680, N494);
nor NOR3 (N684, N663, N371, N597);
and AND3 (N685, N678, N136, N492);
nor NOR3 (N686, N685, N44, N507);
buf BUF1 (N687, N675);
not NOT1 (N688, N682);
xor XOR2 (N689, N684, N583);
buf BUF1 (N690, N674);
nor NOR2 (N691, N689, N235);
buf BUF1 (N692, N686);
xor XOR2 (N693, N683, N182);
nor NOR4 (N694, N692, N39, N31, N279);
xor XOR2 (N695, N688, N268);
xor XOR2 (N696, N687, N70);
xor XOR2 (N697, N696, N181);
nand NAND3 (N698, N694, N566, N417);
xor XOR2 (N699, N695, N167);
or OR3 (N700, N676, N657, N503);
nand NAND3 (N701, N698, N242, N246);
or OR3 (N702, N681, N682, N283);
or OR2 (N703, N701, N517);
and AND3 (N704, N700, N618, N364);
and AND3 (N705, N704, N251, N280);
xor XOR2 (N706, N671, N297);
xor XOR2 (N707, N703, N631);
xor XOR2 (N708, N691, N20);
or OR2 (N709, N690, N193);
and AND3 (N710, N702, N314, N434);
buf BUF1 (N711, N693);
and AND4 (N712, N699, N97, N435, N185);
or OR2 (N713, N706, N260);
and AND3 (N714, N713, N567, N328);
buf BUF1 (N715, N697);
or OR2 (N716, N707, N498);
xor XOR2 (N717, N710, N201);
not NOT1 (N718, N669);
or OR3 (N719, N714, N372, N483);
buf BUF1 (N720, N709);
not NOT1 (N721, N719);
nand NAND4 (N722, N721, N232, N631, N135);
nand NAND4 (N723, N720, N219, N677, N561);
not NOT1 (N724, N708);
nor NOR4 (N725, N718, N260, N724, N555);
not NOT1 (N726, N131);
or OR2 (N727, N705, N636);
nand NAND3 (N728, N712, N678, N587);
nor NOR2 (N729, N715, N408);
nor NOR4 (N730, N726, N285, N503, N408);
not NOT1 (N731, N723);
or OR2 (N732, N711, N27);
nand NAND4 (N733, N731, N658, N296, N190);
and AND3 (N734, N733, N325, N160);
nor NOR4 (N735, N727, N525, N512, N208);
nand NAND3 (N736, N728, N69, N171);
nor NOR2 (N737, N717, N114);
nand NAND2 (N738, N737, N202);
nor NOR3 (N739, N716, N557, N327);
not NOT1 (N740, N734);
not NOT1 (N741, N722);
buf BUF1 (N742, N739);
and AND4 (N743, N738, N198, N426, N730);
xor XOR2 (N744, N624, N705);
not NOT1 (N745, N729);
buf BUF1 (N746, N732);
xor XOR2 (N747, N742, N648);
buf BUF1 (N748, N745);
nand NAND2 (N749, N746, N400);
buf BUF1 (N750, N744);
not NOT1 (N751, N740);
xor XOR2 (N752, N725, N731);
or OR4 (N753, N743, N87, N436, N454);
not NOT1 (N754, N741);
xor XOR2 (N755, N753, N378);
nor NOR3 (N756, N752, N563, N593);
nand NAND3 (N757, N756, N509, N134);
nand NAND4 (N758, N736, N209, N331, N572);
or OR3 (N759, N750, N294, N304);
and AND3 (N760, N749, N526, N42);
not NOT1 (N761, N755);
nor NOR3 (N762, N757, N646, N490);
or OR2 (N763, N748, N6);
nand NAND3 (N764, N751, N653, N652);
buf BUF1 (N765, N763);
nand NAND4 (N766, N747, N324, N309, N93);
nand NAND4 (N767, N765, N677, N564, N171);
nand NAND4 (N768, N761, N690, N246, N209);
or OR3 (N769, N766, N467, N215);
or OR4 (N770, N735, N288, N627, N114);
not NOT1 (N771, N760);
not NOT1 (N772, N762);
buf BUF1 (N773, N772);
not NOT1 (N774, N770);
or OR2 (N775, N768, N252);
not NOT1 (N776, N773);
buf BUF1 (N777, N774);
buf BUF1 (N778, N777);
nand NAND2 (N779, N759, N560);
nor NOR3 (N780, N758, N117, N108);
nor NOR2 (N781, N775, N166);
or OR4 (N782, N769, N454, N733, N428);
and AND4 (N783, N776, N594, N682, N412);
not NOT1 (N784, N764);
xor XOR2 (N785, N780, N697);
nor NOR4 (N786, N782, N18, N574, N260);
not NOT1 (N787, N786);
xor XOR2 (N788, N787, N525);
nor NOR4 (N789, N783, N229, N77, N631);
buf BUF1 (N790, N784);
xor XOR2 (N791, N781, N618);
buf BUF1 (N792, N767);
and AND2 (N793, N789, N417);
nand NAND2 (N794, N788, N748);
xor XOR2 (N795, N778, N773);
nor NOR2 (N796, N771, N574);
xor XOR2 (N797, N754, N1);
and AND2 (N798, N791, N345);
not NOT1 (N799, N792);
or OR2 (N800, N798, N798);
nand NAND4 (N801, N779, N519, N734, N311);
and AND2 (N802, N796, N112);
or OR2 (N803, N794, N202);
and AND4 (N804, N801, N335, N536, N320);
xor XOR2 (N805, N797, N440);
or OR2 (N806, N803, N238);
and AND3 (N807, N793, N55, N172);
or OR3 (N808, N807, N358, N661);
or OR3 (N809, N802, N709, N308);
and AND3 (N810, N795, N369, N168);
xor XOR2 (N811, N808, N44);
or OR2 (N812, N805, N431);
buf BUF1 (N813, N785);
and AND2 (N814, N790, N52);
xor XOR2 (N815, N811, N530);
buf BUF1 (N816, N800);
not NOT1 (N817, N814);
not NOT1 (N818, N809);
not NOT1 (N819, N810);
or OR3 (N820, N817, N777, N776);
xor XOR2 (N821, N806, N133);
or OR4 (N822, N815, N437, N228, N225);
and AND2 (N823, N822, N558);
not NOT1 (N824, N821);
nor NOR3 (N825, N812, N375, N324);
and AND4 (N826, N824, N540, N587, N25);
xor XOR2 (N827, N825, N798);
nand NAND3 (N828, N816, N396, N718);
and AND2 (N829, N823, N461);
not NOT1 (N830, N813);
buf BUF1 (N831, N826);
nand NAND2 (N832, N829, N615);
xor XOR2 (N833, N830, N709);
and AND3 (N834, N833, N274, N282);
not NOT1 (N835, N820);
nor NOR4 (N836, N818, N32, N20, N428);
xor XOR2 (N837, N831, N407);
xor XOR2 (N838, N799, N213);
and AND2 (N839, N804, N325);
or OR2 (N840, N839, N600);
buf BUF1 (N841, N832);
xor XOR2 (N842, N827, N157);
nor NOR2 (N843, N840, N442);
nor NOR3 (N844, N828, N613, N663);
and AND3 (N845, N819, N468, N649);
nand NAND2 (N846, N835, N655);
nor NOR2 (N847, N842, N607);
xor XOR2 (N848, N844, N407);
xor XOR2 (N849, N848, N614);
or OR3 (N850, N834, N482, N779);
or OR4 (N851, N838, N823, N36, N681);
nand NAND3 (N852, N837, N691, N520);
and AND2 (N853, N850, N832);
xor XOR2 (N854, N851, N218);
nor NOR4 (N855, N845, N636, N519, N368);
nor NOR3 (N856, N841, N634, N815);
and AND3 (N857, N855, N473, N576);
buf BUF1 (N858, N853);
nor NOR3 (N859, N836, N832, N393);
and AND3 (N860, N857, N13, N24);
and AND2 (N861, N854, N273);
and AND2 (N862, N858, N362);
or OR3 (N863, N847, N301, N598);
or OR4 (N864, N862, N859, N318, N722);
nand NAND3 (N865, N384, N110, N404);
or OR4 (N866, N863, N133, N61, N112);
not NOT1 (N867, N860);
xor XOR2 (N868, N866, N469);
or OR4 (N869, N864, N363, N351, N775);
and AND2 (N870, N867, N848);
nor NOR2 (N871, N868, N768);
nor NOR2 (N872, N869, N280);
nor NOR2 (N873, N861, N538);
xor XOR2 (N874, N852, N48);
nor NOR2 (N875, N871, N46);
nor NOR2 (N876, N843, N562);
not NOT1 (N877, N849);
buf BUF1 (N878, N846);
nor NOR4 (N879, N870, N687, N811, N672);
or OR3 (N880, N856, N649, N45);
xor XOR2 (N881, N880, N839);
or OR4 (N882, N879, N129, N124, N204);
xor XOR2 (N883, N874, N422);
buf BUF1 (N884, N873);
nand NAND4 (N885, N882, N864, N313, N239);
not NOT1 (N886, N877);
nand NAND4 (N887, N883, N236, N778, N874);
xor XOR2 (N888, N881, N170);
nor NOR3 (N889, N884, N162, N8);
or OR2 (N890, N872, N237);
buf BUF1 (N891, N875);
and AND4 (N892, N865, N600, N708, N370);
buf BUF1 (N893, N888);
and AND3 (N894, N892, N347, N131);
buf BUF1 (N895, N893);
not NOT1 (N896, N876);
buf BUF1 (N897, N887);
or OR2 (N898, N895, N442);
buf BUF1 (N899, N897);
not NOT1 (N900, N889);
xor XOR2 (N901, N878, N542);
nor NOR2 (N902, N886, N729);
not NOT1 (N903, N896);
nand NAND4 (N904, N899, N18, N105, N423);
nor NOR2 (N905, N885, N534);
and AND2 (N906, N898, N339);
not NOT1 (N907, N891);
buf BUF1 (N908, N905);
xor XOR2 (N909, N902, N410);
xor XOR2 (N910, N904, N591);
or OR3 (N911, N908, N822, N457);
buf BUF1 (N912, N910);
nor NOR4 (N913, N903, N231, N711, N742);
nor NOR2 (N914, N913, N500);
and AND2 (N915, N901, N444);
and AND2 (N916, N900, N121);
and AND4 (N917, N907, N497, N25, N753);
xor XOR2 (N918, N906, N200);
xor XOR2 (N919, N890, N235);
nand NAND2 (N920, N894, N575);
and AND4 (N921, N911, N668, N220, N887);
not NOT1 (N922, N912);
nand NAND3 (N923, N920, N651, N762);
nand NAND2 (N924, N923, N616);
xor XOR2 (N925, N924, N222);
and AND4 (N926, N916, N838, N301, N729);
xor XOR2 (N927, N914, N174);
and AND3 (N928, N917, N463, N277);
nand NAND4 (N929, N927, N581, N23, N560);
not NOT1 (N930, N922);
xor XOR2 (N931, N915, N437);
and AND2 (N932, N928, N491);
xor XOR2 (N933, N930, N364);
xor XOR2 (N934, N919, N518);
nand NAND2 (N935, N925, N402);
xor XOR2 (N936, N935, N450);
and AND4 (N937, N929, N291, N2, N733);
xor XOR2 (N938, N932, N546);
xor XOR2 (N939, N933, N667);
and AND4 (N940, N938, N904, N396, N54);
and AND3 (N941, N921, N757, N100);
not NOT1 (N942, N939);
or OR2 (N943, N918, N96);
or OR2 (N944, N937, N414);
not NOT1 (N945, N943);
or OR3 (N946, N931, N200, N922);
buf BUF1 (N947, N941);
or OR2 (N948, N909, N527);
nand NAND4 (N949, N947, N448, N218, N11);
or OR2 (N950, N944, N792);
nand NAND2 (N951, N940, N924);
not NOT1 (N952, N948);
and AND4 (N953, N936, N443, N658, N723);
not NOT1 (N954, N953);
nand NAND3 (N955, N945, N583, N873);
xor XOR2 (N956, N942, N847);
nand NAND3 (N957, N956, N946, N723);
and AND4 (N958, N606, N655, N256, N578);
and AND4 (N959, N954, N101, N949, N762);
nor NOR4 (N960, N654, N492, N139, N397);
nor NOR4 (N961, N958, N263, N199, N117);
or OR3 (N962, N961, N506, N112);
and AND3 (N963, N957, N521, N29);
nand NAND3 (N964, N955, N547, N641);
not NOT1 (N965, N962);
nand NAND3 (N966, N964, N606, N591);
xor XOR2 (N967, N952, N361);
nand NAND3 (N968, N965, N910, N228);
or OR2 (N969, N926, N668);
and AND2 (N970, N950, N693);
and AND3 (N971, N967, N819, N18);
or OR2 (N972, N966, N655);
xor XOR2 (N973, N970, N392);
nor NOR2 (N974, N934, N808);
buf BUF1 (N975, N963);
nor NOR3 (N976, N960, N125, N943);
xor XOR2 (N977, N976, N63);
not NOT1 (N978, N959);
or OR2 (N979, N973, N69);
not NOT1 (N980, N979);
not NOT1 (N981, N980);
nand NAND3 (N982, N971, N439, N25);
or OR4 (N983, N969, N779, N377, N669);
xor XOR2 (N984, N981, N485);
or OR4 (N985, N984, N258, N977, N633);
and AND4 (N986, N341, N574, N875, N810);
buf BUF1 (N987, N972);
xor XOR2 (N988, N983, N293);
nand NAND2 (N989, N951, N143);
not NOT1 (N990, N978);
nor NOR2 (N991, N985, N374);
buf BUF1 (N992, N991);
nor NOR2 (N993, N986, N697);
or OR2 (N994, N990, N331);
not NOT1 (N995, N975);
xor XOR2 (N996, N988, N8);
and AND4 (N997, N982, N978, N557, N866);
xor XOR2 (N998, N987, N12);
and AND2 (N999, N998, N480);
and AND2 (N1000, N997, N544);
xor XOR2 (N1001, N989, N561);
buf BUF1 (N1002, N993);
buf BUF1 (N1003, N968);
nand NAND4 (N1004, N1000, N649, N756, N749);
buf BUF1 (N1005, N974);
not NOT1 (N1006, N1004);
nor NOR2 (N1007, N1006, N86);
or OR2 (N1008, N1002, N59);
or OR3 (N1009, N994, N684, N309);
not NOT1 (N1010, N1005);
xor XOR2 (N1011, N1003, N655);
not NOT1 (N1012, N999);
nand NAND4 (N1013, N1011, N853, N608, N412);
or OR3 (N1014, N1001, N314, N329);
nor NOR2 (N1015, N1008, N677);
buf BUF1 (N1016, N995);
xor XOR2 (N1017, N1014, N638);
buf BUF1 (N1018, N1007);
xor XOR2 (N1019, N1015, N414);
or OR4 (N1020, N1017, N67, N739, N257);
and AND4 (N1021, N1010, N648, N253, N632);
not NOT1 (N1022, N1020);
xor XOR2 (N1023, N996, N668);
and AND4 (N1024, N1023, N773, N197, N126);
nor NOR2 (N1025, N1012, N235);
not NOT1 (N1026, N1018);
buf BUF1 (N1027, N992);
or OR2 (N1028, N1021, N346);
buf BUF1 (N1029, N1022);
nor NOR2 (N1030, N1025, N365);
buf BUF1 (N1031, N1024);
not NOT1 (N1032, N1009);
or OR3 (N1033, N1013, N68, N252);
not NOT1 (N1034, N1029);
not NOT1 (N1035, N1026);
or OR3 (N1036, N1028, N499, N383);
xor XOR2 (N1037, N1035, N169);
or OR3 (N1038, N1034, N347, N252);
nor NOR3 (N1039, N1032, N168, N896);
not NOT1 (N1040, N1016);
nor NOR2 (N1041, N1030, N810);
xor XOR2 (N1042, N1037, N698);
buf BUF1 (N1043, N1039);
nand NAND4 (N1044, N1033, N3, N780, N889);
xor XOR2 (N1045, N1042, N559);
nor NOR2 (N1046, N1044, N210);
nor NOR4 (N1047, N1038, N934, N12, N318);
or OR3 (N1048, N1036, N516, N230);
or OR2 (N1049, N1040, N278);
nand NAND3 (N1050, N1046, N1016, N849);
nor NOR4 (N1051, N1048, N683, N689, N35);
or OR2 (N1052, N1043, N1047);
nor NOR3 (N1053, N5, N62, N706);
or OR4 (N1054, N1053, N29, N484, N521);
xor XOR2 (N1055, N1050, N802);
not NOT1 (N1056, N1045);
buf BUF1 (N1057, N1055);
nor NOR4 (N1058, N1056, N112, N297, N736);
not NOT1 (N1059, N1049);
xor XOR2 (N1060, N1058, N999);
buf BUF1 (N1061, N1057);
buf BUF1 (N1062, N1059);
and AND3 (N1063, N1062, N700, N352);
xor XOR2 (N1064, N1052, N711);
xor XOR2 (N1065, N1064, N140);
and AND4 (N1066, N1065, N1023, N1014, N15);
nand NAND4 (N1067, N1066, N460, N336, N1050);
buf BUF1 (N1068, N1019);
and AND2 (N1069, N1041, N387);
not NOT1 (N1070, N1051);
not NOT1 (N1071, N1054);
and AND2 (N1072, N1031, N862);
nand NAND3 (N1073, N1060, N850, N695);
not NOT1 (N1074, N1063);
nor NOR2 (N1075, N1068, N1022);
buf BUF1 (N1076, N1070);
or OR3 (N1077, N1071, N42, N427);
buf BUF1 (N1078, N1076);
or OR3 (N1079, N1077, N664, N1048);
xor XOR2 (N1080, N1027, N682);
and AND4 (N1081, N1079, N825, N326, N101);
nand NAND4 (N1082, N1080, N331, N408, N434);
nand NAND3 (N1083, N1081, N575, N932);
nor NOR2 (N1084, N1073, N967);
not NOT1 (N1085, N1074);
xor XOR2 (N1086, N1069, N634);
and AND3 (N1087, N1078, N352, N30);
xor XOR2 (N1088, N1067, N142);
not NOT1 (N1089, N1082);
xor XOR2 (N1090, N1085, N625);
buf BUF1 (N1091, N1084);
and AND3 (N1092, N1087, N778, N1075);
not NOT1 (N1093, N303);
nand NAND3 (N1094, N1091, N122, N698);
nor NOR2 (N1095, N1086, N1021);
and AND3 (N1096, N1072, N129, N823);
or OR3 (N1097, N1096, N533, N444);
nand NAND4 (N1098, N1093, N819, N1097, N661);
xor XOR2 (N1099, N417, N912);
xor XOR2 (N1100, N1094, N705);
xor XOR2 (N1101, N1095, N860);
nand NAND2 (N1102, N1083, N305);
nand NAND4 (N1103, N1098, N578, N913, N143);
nor NOR3 (N1104, N1061, N753, N963);
buf BUF1 (N1105, N1104);
not NOT1 (N1106, N1092);
nor NOR4 (N1107, N1088, N578, N328, N510);
xor XOR2 (N1108, N1099, N857);
or OR2 (N1109, N1101, N1091);
buf BUF1 (N1110, N1090);
nand NAND3 (N1111, N1109, N947, N900);
and AND2 (N1112, N1106, N376);
not NOT1 (N1113, N1111);
xor XOR2 (N1114, N1113, N927);
xor XOR2 (N1115, N1110, N772);
not NOT1 (N1116, N1105);
or OR3 (N1117, N1108, N228, N465);
nor NOR3 (N1118, N1089, N544, N757);
or OR2 (N1119, N1112, N190);
xor XOR2 (N1120, N1103, N120);
and AND3 (N1121, N1119, N437, N1102);
nor NOR2 (N1122, N39, N392);
xor XOR2 (N1123, N1107, N395);
xor XOR2 (N1124, N1116, N909);
not NOT1 (N1125, N1115);
nor NOR3 (N1126, N1114, N891, N907);
nor NOR3 (N1127, N1121, N630, N20);
not NOT1 (N1128, N1127);
not NOT1 (N1129, N1123);
or OR3 (N1130, N1118, N757, N230);
and AND4 (N1131, N1129, N222, N542, N319);
nor NOR3 (N1132, N1120, N717, N762);
xor XOR2 (N1133, N1122, N45);
or OR2 (N1134, N1126, N352);
nand NAND3 (N1135, N1131, N634, N60);
buf BUF1 (N1136, N1117);
or OR4 (N1137, N1124, N1129, N420, N1095);
not NOT1 (N1138, N1137);
nor NOR2 (N1139, N1125, N851);
xor XOR2 (N1140, N1132, N499);
not NOT1 (N1141, N1140);
nand NAND4 (N1142, N1130, N204, N520, N206);
nand NAND2 (N1143, N1136, N462);
not NOT1 (N1144, N1139);
nor NOR2 (N1145, N1133, N579);
not NOT1 (N1146, N1144);
and AND3 (N1147, N1143, N413, N119);
xor XOR2 (N1148, N1142, N85);
or OR4 (N1149, N1148, N357, N75, N722);
or OR2 (N1150, N1146, N359);
and AND4 (N1151, N1145, N934, N1088, N266);
and AND3 (N1152, N1150, N391, N192);
or OR2 (N1153, N1149, N1036);
nand NAND2 (N1154, N1100, N1075);
nor NOR3 (N1155, N1134, N211, N80);
or OR3 (N1156, N1155, N102, N990);
nor NOR3 (N1157, N1153, N1092, N243);
not NOT1 (N1158, N1147);
not NOT1 (N1159, N1156);
nand NAND3 (N1160, N1154, N501, N719);
nand NAND4 (N1161, N1157, N333, N1071, N498);
buf BUF1 (N1162, N1151);
not NOT1 (N1163, N1158);
or OR3 (N1164, N1160, N408, N285);
buf BUF1 (N1165, N1128);
and AND4 (N1166, N1162, N312, N252, N527);
and AND3 (N1167, N1165, N796, N439);
xor XOR2 (N1168, N1138, N965);
not NOT1 (N1169, N1152);
or OR3 (N1170, N1163, N125, N313);
or OR4 (N1171, N1161, N937, N524, N737);
not NOT1 (N1172, N1171);
nor NOR3 (N1173, N1168, N620, N155);
not NOT1 (N1174, N1159);
nand NAND2 (N1175, N1173, N1072);
or OR3 (N1176, N1166, N967, N1042);
buf BUF1 (N1177, N1169);
xor XOR2 (N1178, N1175, N63);
nand NAND4 (N1179, N1170, N471, N634, N422);
xor XOR2 (N1180, N1174, N1010);
buf BUF1 (N1181, N1172);
nor NOR2 (N1182, N1177, N498);
nor NOR2 (N1183, N1182, N1013);
xor XOR2 (N1184, N1181, N300);
buf BUF1 (N1185, N1179);
and AND2 (N1186, N1176, N221);
and AND2 (N1187, N1178, N410);
nor NOR4 (N1188, N1167, N352, N32, N64);
or OR2 (N1189, N1184, N160);
or OR3 (N1190, N1188, N530, N1018);
xor XOR2 (N1191, N1185, N314);
and AND4 (N1192, N1190, N561, N707, N1106);
and AND4 (N1193, N1141, N341, N593, N759);
nor NOR2 (N1194, N1180, N806);
buf BUF1 (N1195, N1194);
nor NOR2 (N1196, N1195, N272);
not NOT1 (N1197, N1135);
buf BUF1 (N1198, N1191);
nor NOR2 (N1199, N1198, N217);
not NOT1 (N1200, N1187);
xor XOR2 (N1201, N1193, N288);
xor XOR2 (N1202, N1201, N910);
xor XOR2 (N1203, N1189, N20);
nand NAND3 (N1204, N1199, N754, N276);
xor XOR2 (N1205, N1204, N533);
nand NAND4 (N1206, N1200, N680, N1109, N1045);
and AND2 (N1207, N1202, N481);
xor XOR2 (N1208, N1206, N1121);
and AND2 (N1209, N1192, N1097);
not NOT1 (N1210, N1205);
nand NAND2 (N1211, N1197, N1083);
nor NOR3 (N1212, N1211, N1091, N880);
buf BUF1 (N1213, N1209);
not NOT1 (N1214, N1196);
or OR3 (N1215, N1212, N801, N188);
buf BUF1 (N1216, N1214);
not NOT1 (N1217, N1183);
not NOT1 (N1218, N1203);
nand NAND3 (N1219, N1208, N602, N1075);
or OR4 (N1220, N1210, N274, N840, N466);
buf BUF1 (N1221, N1164);
nand NAND2 (N1222, N1216, N377);
nand NAND2 (N1223, N1221, N53);
not NOT1 (N1224, N1219);
buf BUF1 (N1225, N1215);
not NOT1 (N1226, N1207);
xor XOR2 (N1227, N1213, N146);
or OR2 (N1228, N1227, N159);
nor NOR4 (N1229, N1228, N621, N345, N536);
xor XOR2 (N1230, N1229, N1164);
buf BUF1 (N1231, N1222);
and AND3 (N1232, N1224, N12, N1083);
not NOT1 (N1233, N1232);
buf BUF1 (N1234, N1186);
and AND3 (N1235, N1226, N1136, N768);
xor XOR2 (N1236, N1233, N669);
buf BUF1 (N1237, N1235);
or OR4 (N1238, N1231, N891, N1175, N1191);
and AND3 (N1239, N1218, N66, N1237);
nor NOR3 (N1240, N1002, N130, N51);
and AND2 (N1241, N1236, N1226);
buf BUF1 (N1242, N1225);
nand NAND4 (N1243, N1241, N855, N846, N234);
not NOT1 (N1244, N1240);
xor XOR2 (N1245, N1220, N913);
nor NOR3 (N1246, N1234, N39, N411);
or OR3 (N1247, N1244, N620, N991);
xor XOR2 (N1248, N1242, N929);
nand NAND2 (N1249, N1248, N833);
and AND3 (N1250, N1243, N336, N773);
nand NAND4 (N1251, N1245, N771, N108, N702);
xor XOR2 (N1252, N1250, N631);
xor XOR2 (N1253, N1239, N195);
nand NAND2 (N1254, N1249, N1244);
not NOT1 (N1255, N1217);
and AND4 (N1256, N1255, N327, N1079, N844);
or OR2 (N1257, N1230, N839);
buf BUF1 (N1258, N1252);
and AND3 (N1259, N1253, N441, N237);
xor XOR2 (N1260, N1238, N242);
nor NOR3 (N1261, N1223, N643, N641);
and AND4 (N1262, N1257, N905, N220, N1158);
buf BUF1 (N1263, N1260);
not NOT1 (N1264, N1251);
or OR4 (N1265, N1262, N854, N763, N371);
or OR2 (N1266, N1259, N294);
buf BUF1 (N1267, N1258);
not NOT1 (N1268, N1264);
nor NOR2 (N1269, N1254, N336);
buf BUF1 (N1270, N1246);
nand NAND2 (N1271, N1261, N207);
and AND3 (N1272, N1256, N98, N491);
and AND3 (N1273, N1270, N1134, N236);
nand NAND4 (N1274, N1267, N1083, N236, N558);
xor XOR2 (N1275, N1265, N1063);
nor NOR2 (N1276, N1271, N162);
and AND3 (N1277, N1273, N598, N702);
or OR2 (N1278, N1275, N151);
nand NAND2 (N1279, N1269, N188);
or OR2 (N1280, N1268, N1191);
and AND3 (N1281, N1278, N1231, N1148);
not NOT1 (N1282, N1281);
buf BUF1 (N1283, N1263);
buf BUF1 (N1284, N1247);
nor NOR3 (N1285, N1279, N503, N1072);
and AND3 (N1286, N1266, N587, N1111);
nand NAND4 (N1287, N1280, N1177, N730, N467);
xor XOR2 (N1288, N1284, N130);
buf BUF1 (N1289, N1282);
not NOT1 (N1290, N1283);
not NOT1 (N1291, N1287);
nor NOR2 (N1292, N1289, N354);
and AND3 (N1293, N1277, N192, N370);
xor XOR2 (N1294, N1285, N839);
nor NOR4 (N1295, N1294, N978, N1035, N582);
nand NAND2 (N1296, N1288, N39);
or OR2 (N1297, N1292, N929);
not NOT1 (N1298, N1276);
or OR2 (N1299, N1298, N107);
nor NOR3 (N1300, N1272, N774, N787);
xor XOR2 (N1301, N1286, N198);
or OR3 (N1302, N1301, N467, N1110);
xor XOR2 (N1303, N1274, N746);
buf BUF1 (N1304, N1291);
nor NOR3 (N1305, N1300, N349, N899);
or OR4 (N1306, N1302, N452, N441, N43);
xor XOR2 (N1307, N1306, N35);
xor XOR2 (N1308, N1295, N543);
xor XOR2 (N1309, N1305, N639);
and AND3 (N1310, N1296, N386, N512);
nor NOR2 (N1311, N1297, N615);
nor NOR3 (N1312, N1311, N738, N50);
nand NAND2 (N1313, N1299, N332);
nand NAND4 (N1314, N1307, N251, N451, N134);
nand NAND2 (N1315, N1308, N438);
and AND4 (N1316, N1303, N1266, N1201, N1248);
buf BUF1 (N1317, N1310);
nor NOR4 (N1318, N1293, N760, N574, N185);
and AND2 (N1319, N1315, N218);
nor NOR4 (N1320, N1312, N1279, N579, N477);
buf BUF1 (N1321, N1290);
or OR2 (N1322, N1314, N709);
nor NOR3 (N1323, N1317, N5, N1150);
buf BUF1 (N1324, N1313);
xor XOR2 (N1325, N1321, N471);
xor XOR2 (N1326, N1323, N1277);
or OR2 (N1327, N1316, N1015);
buf BUF1 (N1328, N1304);
xor XOR2 (N1329, N1320, N905);
xor XOR2 (N1330, N1309, N700);
nor NOR2 (N1331, N1319, N375);
or OR2 (N1332, N1327, N574);
xor XOR2 (N1333, N1328, N319);
and AND3 (N1334, N1326, N335, N29);
or OR2 (N1335, N1329, N116);
or OR3 (N1336, N1322, N187, N793);
not NOT1 (N1337, N1330);
nor NOR4 (N1338, N1334, N1017, N677, N509);
nor NOR3 (N1339, N1324, N161, N1080);
not NOT1 (N1340, N1333);
xor XOR2 (N1341, N1340, N719);
xor XOR2 (N1342, N1341, N860);
and AND2 (N1343, N1318, N590);
nor NOR4 (N1344, N1332, N9, N509, N924);
and AND3 (N1345, N1339, N1311, N572);
xor XOR2 (N1346, N1343, N474);
or OR2 (N1347, N1325, N422);
not NOT1 (N1348, N1335);
or OR2 (N1349, N1345, N1067);
and AND3 (N1350, N1331, N937, N1080);
xor XOR2 (N1351, N1338, N1326);
nor NOR4 (N1352, N1344, N836, N679, N202);
xor XOR2 (N1353, N1349, N350);
not NOT1 (N1354, N1348);
nor NOR2 (N1355, N1351, N1025);
nand NAND4 (N1356, N1352, N1314, N493, N1128);
or OR4 (N1357, N1353, N428, N299, N1070);
nor NOR3 (N1358, N1337, N557, N742);
not NOT1 (N1359, N1342);
nor NOR3 (N1360, N1347, N757, N640);
or OR4 (N1361, N1357, N379, N183, N40);
nor NOR3 (N1362, N1361, N993, N703);
nor NOR2 (N1363, N1358, N911);
buf BUF1 (N1364, N1356);
or OR4 (N1365, N1336, N453, N1039, N1113);
nor NOR4 (N1366, N1346, N1299, N937, N263);
xor XOR2 (N1367, N1365, N857);
and AND4 (N1368, N1355, N105, N324, N1106);
and AND3 (N1369, N1362, N550, N922);
buf BUF1 (N1370, N1363);
nand NAND4 (N1371, N1354, N1242, N1210, N275);
or OR3 (N1372, N1350, N184, N102);
xor XOR2 (N1373, N1370, N193);
and AND4 (N1374, N1372, N517, N392, N137);
nor NOR3 (N1375, N1359, N810, N811);
xor XOR2 (N1376, N1371, N538);
nand NAND3 (N1377, N1373, N719, N1348);
and AND3 (N1378, N1374, N489, N1251);
and AND4 (N1379, N1377, N892, N168, N796);
xor XOR2 (N1380, N1367, N635);
and AND2 (N1381, N1380, N130);
buf BUF1 (N1382, N1375);
xor XOR2 (N1383, N1366, N845);
xor XOR2 (N1384, N1383, N57);
and AND3 (N1385, N1382, N760, N403);
buf BUF1 (N1386, N1360);
nor NOR4 (N1387, N1376, N41, N544, N451);
nand NAND4 (N1388, N1364, N1341, N858, N1332);
and AND2 (N1389, N1378, N1001);
or OR2 (N1390, N1386, N1233);
not NOT1 (N1391, N1379);
and AND2 (N1392, N1390, N1330);
nand NAND4 (N1393, N1387, N568, N1258, N120);
xor XOR2 (N1394, N1381, N308);
and AND2 (N1395, N1369, N302);
nand NAND4 (N1396, N1389, N1133, N1001, N955);
xor XOR2 (N1397, N1384, N1364);
nor NOR4 (N1398, N1391, N1053, N996, N239);
nand NAND2 (N1399, N1388, N291);
buf BUF1 (N1400, N1385);
nand NAND4 (N1401, N1396, N1391, N506, N530);
and AND4 (N1402, N1397, N509, N1104, N897);
buf BUF1 (N1403, N1400);
and AND4 (N1404, N1368, N459, N568, N502);
nand NAND3 (N1405, N1401, N397, N600);
nor NOR4 (N1406, N1395, N1320, N412, N122);
or OR2 (N1407, N1393, N720);
not NOT1 (N1408, N1407);
nor NOR2 (N1409, N1404, N1308);
buf BUF1 (N1410, N1394);
xor XOR2 (N1411, N1405, N431);
nor NOR3 (N1412, N1392, N526, N640);
nor NOR2 (N1413, N1412, N839);
and AND3 (N1414, N1413, N719, N652);
nand NAND4 (N1415, N1406, N1237, N292, N1321);
nand NAND4 (N1416, N1410, N376, N255, N922);
and AND3 (N1417, N1411, N465, N711);
nand NAND2 (N1418, N1417, N535);
nand NAND2 (N1419, N1402, N699);
buf BUF1 (N1420, N1419);
xor XOR2 (N1421, N1418, N911);
not NOT1 (N1422, N1416);
nor NOR3 (N1423, N1414, N993, N814);
not NOT1 (N1424, N1422);
not NOT1 (N1425, N1415);
buf BUF1 (N1426, N1408);
or OR2 (N1427, N1399, N266);
xor XOR2 (N1428, N1421, N1106);
xor XOR2 (N1429, N1403, N585);
nor NOR4 (N1430, N1420, N699, N1422, N1072);
and AND3 (N1431, N1423, N450, N693);
nor NOR4 (N1432, N1430, N863, N1272, N641);
or OR4 (N1433, N1424, N498, N254, N149);
or OR4 (N1434, N1432, N393, N1234, N1283);
xor XOR2 (N1435, N1428, N466);
nor NOR2 (N1436, N1398, N519);
or OR3 (N1437, N1427, N315, N107);
nand NAND4 (N1438, N1429, N746, N315, N315);
not NOT1 (N1439, N1438);
or OR4 (N1440, N1437, N31, N790, N1230);
or OR3 (N1441, N1440, N759, N531);
nand NAND3 (N1442, N1441, N1141, N1397);
nand NAND3 (N1443, N1431, N1340, N203);
xor XOR2 (N1444, N1442, N890);
xor XOR2 (N1445, N1426, N491);
or OR4 (N1446, N1434, N363, N1171, N594);
xor XOR2 (N1447, N1443, N731);
not NOT1 (N1448, N1446);
or OR3 (N1449, N1433, N151, N666);
nor NOR2 (N1450, N1436, N852);
nand NAND2 (N1451, N1425, N1074);
xor XOR2 (N1452, N1445, N777);
nand NAND3 (N1453, N1452, N905, N936);
not NOT1 (N1454, N1439);
or OR4 (N1455, N1409, N1090, N462, N406);
nand NAND4 (N1456, N1454, N90, N1406, N1134);
nor NOR2 (N1457, N1450, N1134);
buf BUF1 (N1458, N1457);
nand NAND2 (N1459, N1449, N556);
xor XOR2 (N1460, N1444, N1056);
nand NAND2 (N1461, N1448, N285);
xor XOR2 (N1462, N1451, N277);
buf BUF1 (N1463, N1453);
or OR3 (N1464, N1461, N1417, N1012);
xor XOR2 (N1465, N1458, N486);
nor NOR4 (N1466, N1465, N266, N663, N140);
or OR2 (N1467, N1455, N474);
or OR3 (N1468, N1466, N1186, N697);
or OR4 (N1469, N1460, N402, N714, N1097);
not NOT1 (N1470, N1447);
or OR2 (N1471, N1462, N317);
xor XOR2 (N1472, N1471, N952);
and AND4 (N1473, N1468, N759, N285, N1341);
and AND2 (N1474, N1456, N1195);
nor NOR3 (N1475, N1464, N1295, N7);
nand NAND3 (N1476, N1474, N533, N609);
nor NOR2 (N1477, N1467, N1241);
or OR4 (N1478, N1473, N926, N1261, N957);
buf BUF1 (N1479, N1469);
and AND4 (N1480, N1476, N1200, N1338, N580);
or OR3 (N1481, N1479, N69, N882);
and AND4 (N1482, N1480, N1412, N1125, N516);
xor XOR2 (N1483, N1435, N1208);
buf BUF1 (N1484, N1477);
and AND3 (N1485, N1483, N1388, N760);
nor NOR2 (N1486, N1463, N1459);
and AND4 (N1487, N464, N1138, N247, N182);
buf BUF1 (N1488, N1485);
or OR3 (N1489, N1475, N588, N416);
nand NAND3 (N1490, N1486, N1127, N1170);
nor NOR4 (N1491, N1488, N703, N1235, N668);
nand NAND4 (N1492, N1481, N1321, N1154, N210);
and AND2 (N1493, N1478, N1055);
or OR2 (N1494, N1491, N275);
and AND3 (N1495, N1490, N536, N1255);
or OR2 (N1496, N1472, N328);
not NOT1 (N1497, N1482);
nand NAND2 (N1498, N1495, N1223);
nor NOR3 (N1499, N1470, N1117, N851);
and AND4 (N1500, N1492, N121, N574, N21);
xor XOR2 (N1501, N1498, N799);
nor NOR4 (N1502, N1494, N967, N100, N889);
not NOT1 (N1503, N1487);
and AND3 (N1504, N1501, N1442, N944);
nand NAND2 (N1505, N1504, N767);
nor NOR3 (N1506, N1497, N1222, N990);
or OR3 (N1507, N1500, N727, N1045);
xor XOR2 (N1508, N1499, N1319);
buf BUF1 (N1509, N1505);
or OR3 (N1510, N1493, N1073, N164);
xor XOR2 (N1511, N1503, N1200);
or OR2 (N1512, N1484, N265);
buf BUF1 (N1513, N1508);
xor XOR2 (N1514, N1509, N478);
and AND3 (N1515, N1506, N193, N344);
xor XOR2 (N1516, N1511, N647);
or OR3 (N1517, N1515, N1348, N1056);
nor NOR3 (N1518, N1517, N245, N456);
nand NAND3 (N1519, N1496, N783, N1400);
or OR2 (N1520, N1489, N1307);
nor NOR3 (N1521, N1520, N94, N1341);
nor NOR2 (N1522, N1512, N43);
or OR3 (N1523, N1519, N1116, N1300);
and AND2 (N1524, N1518, N292);
nor NOR3 (N1525, N1514, N1130, N901);
or OR4 (N1526, N1516, N10, N442, N779);
nor NOR3 (N1527, N1502, N656, N1456);
buf BUF1 (N1528, N1513);
not NOT1 (N1529, N1526);
nor NOR3 (N1530, N1523, N808, N1487);
or OR4 (N1531, N1510, N1447, N325, N807);
or OR3 (N1532, N1528, N1060, N757);
and AND4 (N1533, N1527, N737, N1441, N675);
buf BUF1 (N1534, N1533);
nor NOR3 (N1535, N1521, N361, N1365);
not NOT1 (N1536, N1525);
xor XOR2 (N1537, N1529, N955);
not NOT1 (N1538, N1534);
xor XOR2 (N1539, N1532, N172);
xor XOR2 (N1540, N1522, N226);
nor NOR4 (N1541, N1531, N1112, N7, N712);
nand NAND4 (N1542, N1535, N374, N23, N8);
buf BUF1 (N1543, N1541);
not NOT1 (N1544, N1543);
buf BUF1 (N1545, N1539);
and AND3 (N1546, N1524, N1412, N1039);
buf BUF1 (N1547, N1542);
not NOT1 (N1548, N1530);
and AND4 (N1549, N1546, N167, N520, N1115);
not NOT1 (N1550, N1547);
xor XOR2 (N1551, N1544, N1191);
nand NAND2 (N1552, N1545, N1219);
nand NAND3 (N1553, N1537, N200, N613);
xor XOR2 (N1554, N1550, N648);
nand NAND4 (N1555, N1540, N1152, N1381, N451);
not NOT1 (N1556, N1554);
nand NAND3 (N1557, N1538, N1005, N453);
not NOT1 (N1558, N1551);
or OR3 (N1559, N1558, N1409, N484);
buf BUF1 (N1560, N1507);
and AND3 (N1561, N1556, N1180, N287);
or OR3 (N1562, N1549, N262, N677);
buf BUF1 (N1563, N1562);
not NOT1 (N1564, N1536);
not NOT1 (N1565, N1553);
nand NAND4 (N1566, N1557, N1381, N371, N563);
not NOT1 (N1567, N1548);
and AND2 (N1568, N1561, N669);
nor NOR3 (N1569, N1566, N27, N489);
nand NAND2 (N1570, N1564, N1196);
and AND3 (N1571, N1568, N375, N503);
not NOT1 (N1572, N1571);
buf BUF1 (N1573, N1565);
buf BUF1 (N1574, N1567);
buf BUF1 (N1575, N1570);
nor NOR3 (N1576, N1574, N560, N1002);
buf BUF1 (N1577, N1555);
and AND3 (N1578, N1560, N196, N341);
nor NOR2 (N1579, N1573, N511);
not NOT1 (N1580, N1572);
nor NOR4 (N1581, N1563, N1118, N1013, N1143);
buf BUF1 (N1582, N1579);
nor NOR2 (N1583, N1552, N1243);
nor NOR2 (N1584, N1559, N89);
or OR4 (N1585, N1583, N74, N844, N222);
nor NOR2 (N1586, N1581, N649);
and AND2 (N1587, N1585, N174);
and AND4 (N1588, N1578, N1163, N1007, N569);
xor XOR2 (N1589, N1577, N310);
buf BUF1 (N1590, N1586);
not NOT1 (N1591, N1589);
nor NOR4 (N1592, N1584, N1078, N748, N1552);
nor NOR3 (N1593, N1576, N162, N573);
nor NOR3 (N1594, N1582, N1498, N148);
and AND2 (N1595, N1591, N715);
xor XOR2 (N1596, N1595, N5);
buf BUF1 (N1597, N1590);
buf BUF1 (N1598, N1596);
xor XOR2 (N1599, N1594, N96);
nor NOR3 (N1600, N1598, N76, N397);
and AND3 (N1601, N1587, N442, N649);
buf BUF1 (N1602, N1597);
or OR4 (N1603, N1588, N1052, N708, N573);
nand NAND4 (N1604, N1593, N1031, N552, N822);
nor NOR4 (N1605, N1601, N1249, N333, N1366);
nor NOR3 (N1606, N1604, N1424, N292);
and AND2 (N1607, N1605, N137);
nand NAND4 (N1608, N1602, N89, N1040, N550);
nor NOR2 (N1609, N1599, N915);
not NOT1 (N1610, N1592);
buf BUF1 (N1611, N1600);
buf BUF1 (N1612, N1569);
or OR3 (N1613, N1609, N875, N326);
nand NAND3 (N1614, N1610, N1043, N802);
nor NOR2 (N1615, N1611, N1601);
not NOT1 (N1616, N1575);
xor XOR2 (N1617, N1615, N654);
not NOT1 (N1618, N1603);
nand NAND2 (N1619, N1607, N1075);
not NOT1 (N1620, N1612);
buf BUF1 (N1621, N1616);
nand NAND4 (N1622, N1620, N915, N1138, N79);
xor XOR2 (N1623, N1618, N888);
xor XOR2 (N1624, N1622, N283);
buf BUF1 (N1625, N1621);
nor NOR2 (N1626, N1580, N309);
or OR2 (N1627, N1608, N1207);
nor NOR2 (N1628, N1613, N1150);
xor XOR2 (N1629, N1614, N844);
not NOT1 (N1630, N1617);
nand NAND3 (N1631, N1627, N1191, N1593);
nand NAND2 (N1632, N1624, N158);
not NOT1 (N1633, N1623);
not NOT1 (N1634, N1631);
nand NAND4 (N1635, N1634, N274, N1578, N1460);
not NOT1 (N1636, N1629);
buf BUF1 (N1637, N1632);
or OR4 (N1638, N1626, N897, N1146, N490);
and AND2 (N1639, N1628, N503);
buf BUF1 (N1640, N1633);
xor XOR2 (N1641, N1640, N1166);
nand NAND2 (N1642, N1619, N928);
nand NAND2 (N1643, N1638, N383);
or OR4 (N1644, N1637, N1569, N861, N258);
or OR3 (N1645, N1625, N1620, N28);
and AND3 (N1646, N1606, N1586, N401);
buf BUF1 (N1647, N1641);
nor NOR4 (N1648, N1636, N1454, N595, N1059);
and AND3 (N1649, N1635, N1502, N1233);
and AND2 (N1650, N1649, N338);
or OR2 (N1651, N1644, N1290);
buf BUF1 (N1652, N1630);
and AND3 (N1653, N1643, N316, N1017);
nand NAND3 (N1654, N1653, N540, N1293);
nand NAND3 (N1655, N1648, N418, N904);
nand NAND3 (N1656, N1646, N810, N333);
not NOT1 (N1657, N1655);
not NOT1 (N1658, N1657);
buf BUF1 (N1659, N1654);
nor NOR3 (N1660, N1656, N222, N1571);
buf BUF1 (N1661, N1660);
and AND3 (N1662, N1642, N227, N1332);
nand NAND2 (N1663, N1659, N669);
and AND2 (N1664, N1650, N1086);
not NOT1 (N1665, N1645);
nor NOR3 (N1666, N1662, N1051, N507);
xor XOR2 (N1667, N1665, N1496);
xor XOR2 (N1668, N1652, N478);
and AND3 (N1669, N1663, N703, N687);
buf BUF1 (N1670, N1669);
not NOT1 (N1671, N1639);
buf BUF1 (N1672, N1661);
and AND2 (N1673, N1647, N1552);
or OR3 (N1674, N1672, N79, N993);
nor NOR2 (N1675, N1673, N201);
not NOT1 (N1676, N1671);
and AND4 (N1677, N1675, N528, N1176, N1142);
or OR2 (N1678, N1664, N1318);
and AND3 (N1679, N1667, N1250, N1545);
nor NOR4 (N1680, N1678, N779, N646, N1630);
buf BUF1 (N1681, N1676);
nand NAND3 (N1682, N1668, N334, N1328);
and AND2 (N1683, N1682, N695);
buf BUF1 (N1684, N1651);
not NOT1 (N1685, N1670);
or OR4 (N1686, N1684, N873, N657, N364);
nor NOR4 (N1687, N1658, N1371, N432, N1624);
not NOT1 (N1688, N1686);
nand NAND4 (N1689, N1680, N1659, N720, N1134);
nor NOR3 (N1690, N1683, N9, N1347);
nor NOR2 (N1691, N1679, N1575);
and AND3 (N1692, N1691, N1333, N830);
or OR3 (N1693, N1690, N1498, N1621);
nor NOR4 (N1694, N1693, N648, N169, N890);
buf BUF1 (N1695, N1681);
xor XOR2 (N1696, N1677, N726);
not NOT1 (N1697, N1695);
xor XOR2 (N1698, N1697, N281);
not NOT1 (N1699, N1689);
xor XOR2 (N1700, N1687, N1567);
and AND4 (N1701, N1674, N971, N1641, N1131);
or OR4 (N1702, N1699, N1259, N1253, N1272);
xor XOR2 (N1703, N1692, N1533);
not NOT1 (N1704, N1696);
not NOT1 (N1705, N1666);
nor NOR2 (N1706, N1685, N1705);
or OR2 (N1707, N277, N1483);
buf BUF1 (N1708, N1694);
nor NOR4 (N1709, N1703, N466, N326, N690);
xor XOR2 (N1710, N1706, N1315);
and AND4 (N1711, N1708, N892, N8, N988);
xor XOR2 (N1712, N1707, N11);
nand NAND3 (N1713, N1698, N386, N1622);
buf BUF1 (N1714, N1701);
and AND4 (N1715, N1702, N1450, N69, N1598);
and AND3 (N1716, N1704, N1664, N1001);
nor NOR4 (N1717, N1709, N1085, N503, N1419);
nor NOR2 (N1718, N1713, N545);
or OR2 (N1719, N1718, N61);
not NOT1 (N1720, N1716);
or OR2 (N1721, N1717, N1002);
nand NAND3 (N1722, N1720, N87, N685);
buf BUF1 (N1723, N1688);
and AND2 (N1724, N1714, N622);
buf BUF1 (N1725, N1712);
not NOT1 (N1726, N1723);
xor XOR2 (N1727, N1711, N75);
not NOT1 (N1728, N1725);
nor NOR2 (N1729, N1710, N115);
not NOT1 (N1730, N1715);
nor NOR4 (N1731, N1727, N1578, N770, N1704);
nand NAND3 (N1732, N1722, N824, N1205);
nand NAND2 (N1733, N1728, N920);
xor XOR2 (N1734, N1733, N1003);
not NOT1 (N1735, N1724);
and AND4 (N1736, N1730, N461, N51, N1619);
nor NOR3 (N1737, N1731, N1657, N1508);
buf BUF1 (N1738, N1726);
or OR4 (N1739, N1734, N1506, N884, N1072);
nand NAND4 (N1740, N1735, N342, N1600, N333);
buf BUF1 (N1741, N1737);
and AND2 (N1742, N1739, N542);
nor NOR4 (N1743, N1719, N234, N736, N845);
or OR4 (N1744, N1738, N441, N825, N1411);
not NOT1 (N1745, N1700);
nor NOR2 (N1746, N1721, N733);
xor XOR2 (N1747, N1741, N488);
xor XOR2 (N1748, N1742, N1131);
or OR2 (N1749, N1729, N514);
xor XOR2 (N1750, N1746, N419);
nor NOR3 (N1751, N1736, N1565, N847);
nor NOR3 (N1752, N1732, N1326, N1411);
and AND3 (N1753, N1743, N1273, N1100);
and AND3 (N1754, N1747, N1660, N646);
buf BUF1 (N1755, N1750);
nor NOR4 (N1756, N1740, N936, N943, N984);
xor XOR2 (N1757, N1744, N34);
not NOT1 (N1758, N1745);
buf BUF1 (N1759, N1748);
nand NAND3 (N1760, N1759, N1059, N738);
nor NOR2 (N1761, N1756, N1368);
or OR2 (N1762, N1749, N1088);
and AND3 (N1763, N1753, N1238, N1187);
not NOT1 (N1764, N1755);
not NOT1 (N1765, N1760);
and AND2 (N1766, N1764, N415);
nor NOR4 (N1767, N1752, N852, N819, N1402);
xor XOR2 (N1768, N1757, N1413);
or OR4 (N1769, N1754, N1058, N1372, N1036);
nor NOR3 (N1770, N1758, N777, N662);
or OR2 (N1771, N1765, N1226);
xor XOR2 (N1772, N1767, N1753);
buf BUF1 (N1773, N1771);
buf BUF1 (N1774, N1770);
buf BUF1 (N1775, N1751);
xor XOR2 (N1776, N1762, N1015);
nand NAND3 (N1777, N1769, N1380, N740);
buf BUF1 (N1778, N1768);
nand NAND2 (N1779, N1776, N1637);
or OR3 (N1780, N1761, N1549, N512);
or OR3 (N1781, N1773, N392, N1732);
or OR2 (N1782, N1778, N237);
nand NAND4 (N1783, N1772, N1199, N959, N1603);
or OR3 (N1784, N1780, N136, N1067);
nand NAND2 (N1785, N1777, N137);
xor XOR2 (N1786, N1784, N858);
not NOT1 (N1787, N1783);
not NOT1 (N1788, N1781);
xor XOR2 (N1789, N1766, N136);
xor XOR2 (N1790, N1763, N1450);
buf BUF1 (N1791, N1787);
or OR4 (N1792, N1790, N377, N161, N1123);
nor NOR2 (N1793, N1792, N555);
nor NOR3 (N1794, N1785, N813, N1731);
nor NOR3 (N1795, N1775, N51, N52);
not NOT1 (N1796, N1782);
nor NOR4 (N1797, N1789, N1104, N1264, N488);
buf BUF1 (N1798, N1779);
xor XOR2 (N1799, N1797, N1391);
buf BUF1 (N1800, N1774);
nand NAND2 (N1801, N1799, N1725);
nand NAND3 (N1802, N1788, N1053, N615);
nand NAND4 (N1803, N1798, N1243, N9, N976);
not NOT1 (N1804, N1793);
nor NOR4 (N1805, N1800, N638, N1084, N294);
buf BUF1 (N1806, N1805);
xor XOR2 (N1807, N1802, N97);
or OR2 (N1808, N1803, N22);
nor NOR2 (N1809, N1804, N971);
xor XOR2 (N1810, N1806, N86);
and AND2 (N1811, N1809, N1240);
and AND3 (N1812, N1786, N1516, N516);
nand NAND3 (N1813, N1794, N864, N189);
nand NAND3 (N1814, N1813, N673, N1464);
nand NAND2 (N1815, N1814, N70);
xor XOR2 (N1816, N1815, N965);
buf BUF1 (N1817, N1801);
not NOT1 (N1818, N1817);
xor XOR2 (N1819, N1816, N984);
nor NOR3 (N1820, N1795, N541, N536);
not NOT1 (N1821, N1818);
nand NAND4 (N1822, N1808, N738, N1092, N1724);
buf BUF1 (N1823, N1812);
or OR3 (N1824, N1822, N111, N1536);
buf BUF1 (N1825, N1824);
or OR3 (N1826, N1791, N255, N1808);
nand NAND4 (N1827, N1810, N228, N1269, N681);
nand NAND3 (N1828, N1796, N513, N127);
or OR3 (N1829, N1828, N1275, N1653);
not NOT1 (N1830, N1826);
or OR2 (N1831, N1829, N302);
and AND4 (N1832, N1820, N1497, N1064, N1044);
nor NOR2 (N1833, N1830, N508);
not NOT1 (N1834, N1821);
not NOT1 (N1835, N1833);
not NOT1 (N1836, N1835);
buf BUF1 (N1837, N1811);
nand NAND3 (N1838, N1837, N952, N1037);
nor NOR4 (N1839, N1823, N1349, N1265, N1028);
buf BUF1 (N1840, N1819);
not NOT1 (N1841, N1840);
or OR3 (N1842, N1825, N1038, N1475);
xor XOR2 (N1843, N1836, N62);
or OR3 (N1844, N1827, N401, N942);
not NOT1 (N1845, N1839);
nor NOR2 (N1846, N1842, N1040);
nor NOR4 (N1847, N1807, N638, N1398, N435);
nand NAND4 (N1848, N1845, N1512, N932, N1403);
or OR4 (N1849, N1838, N396, N822, N255);
not NOT1 (N1850, N1849);
xor XOR2 (N1851, N1850, N934);
buf BUF1 (N1852, N1832);
buf BUF1 (N1853, N1844);
or OR3 (N1854, N1853, N1166, N217);
not NOT1 (N1855, N1848);
not NOT1 (N1856, N1855);
nand NAND3 (N1857, N1831, N940, N539);
or OR4 (N1858, N1854, N559, N1794, N305);
nor NOR4 (N1859, N1857, N323, N1547, N1033);
nor NOR2 (N1860, N1847, N192);
and AND3 (N1861, N1841, N1786, N1212);
or OR2 (N1862, N1852, N353);
nand NAND4 (N1863, N1859, N1826, N821, N80);
nand NAND4 (N1864, N1860, N1594, N1669, N1713);
xor XOR2 (N1865, N1863, N697);
nand NAND4 (N1866, N1856, N1832, N1830, N404);
and AND4 (N1867, N1866, N1508, N1718, N154);
xor XOR2 (N1868, N1862, N738);
xor XOR2 (N1869, N1851, N194);
nand NAND2 (N1870, N1865, N1703);
not NOT1 (N1871, N1867);
xor XOR2 (N1872, N1843, N552);
nor NOR4 (N1873, N1871, N91, N1730, N724);
nor NOR3 (N1874, N1869, N343, N937);
nand NAND3 (N1875, N1868, N1325, N1776);
nor NOR4 (N1876, N1861, N1529, N778, N345);
buf BUF1 (N1877, N1870);
nor NOR3 (N1878, N1858, N533, N63);
or OR3 (N1879, N1834, N551, N1767);
not NOT1 (N1880, N1877);
xor XOR2 (N1881, N1876, N1216);
or OR2 (N1882, N1879, N55);
not NOT1 (N1883, N1882);
nor NOR4 (N1884, N1881, N1829, N769, N35);
buf BUF1 (N1885, N1875);
and AND4 (N1886, N1884, N570, N1033, N663);
nor NOR4 (N1887, N1885, N1587, N171, N74);
and AND3 (N1888, N1880, N937, N502);
and AND4 (N1889, N1888, N972, N1843, N226);
nand NAND4 (N1890, N1864, N1136, N452, N1858);
nand NAND3 (N1891, N1886, N707, N750);
nor NOR3 (N1892, N1846, N317, N1227);
buf BUF1 (N1893, N1872);
nand NAND3 (N1894, N1890, N71, N475);
nor NOR4 (N1895, N1874, N284, N890, N97);
nand NAND4 (N1896, N1891, N609, N1659, N1509);
or OR2 (N1897, N1883, N314);
nand NAND4 (N1898, N1887, N1590, N819, N1818);
or OR3 (N1899, N1878, N1339, N114);
or OR2 (N1900, N1895, N627);
buf BUF1 (N1901, N1900);
not NOT1 (N1902, N1889);
nor NOR3 (N1903, N1893, N1599, N437);
nor NOR2 (N1904, N1896, N669);
not NOT1 (N1905, N1899);
nor NOR2 (N1906, N1903, N1630);
buf BUF1 (N1907, N1902);
xor XOR2 (N1908, N1873, N386);
not NOT1 (N1909, N1907);
or OR2 (N1910, N1906, N1084);
buf BUF1 (N1911, N1892);
buf BUF1 (N1912, N1905);
buf BUF1 (N1913, N1894);
or OR4 (N1914, N1897, N1256, N1130, N532);
or OR2 (N1915, N1909, N339);
and AND2 (N1916, N1914, N605);
nor NOR2 (N1917, N1913, N69);
nand NAND2 (N1918, N1915, N1271);
not NOT1 (N1919, N1904);
xor XOR2 (N1920, N1916, N535);
buf BUF1 (N1921, N1908);
and AND2 (N1922, N1918, N867);
xor XOR2 (N1923, N1921, N352);
not NOT1 (N1924, N1910);
nor NOR4 (N1925, N1912, N137, N1692, N1017);
and AND2 (N1926, N1925, N634);
buf BUF1 (N1927, N1920);
buf BUF1 (N1928, N1911);
nand NAND4 (N1929, N1901, N252, N1206, N1070);
nor NOR2 (N1930, N1898, N863);
or OR4 (N1931, N1929, N1379, N403, N473);
and AND3 (N1932, N1931, N509, N1395);
and AND4 (N1933, N1932, N1022, N1281, N1281);
nand NAND3 (N1934, N1927, N1466, N1001);
or OR2 (N1935, N1919, N658);
xor XOR2 (N1936, N1917, N665);
nand NAND4 (N1937, N1936, N1347, N754, N452);
nand NAND4 (N1938, N1933, N449, N1240, N399);
nand NAND3 (N1939, N1934, N266, N1704);
and AND3 (N1940, N1938, N137, N1427);
and AND3 (N1941, N1926, N1292, N238);
and AND3 (N1942, N1924, N1393, N361);
not NOT1 (N1943, N1937);
not NOT1 (N1944, N1922);
nor NOR3 (N1945, N1943, N670, N1068);
nand NAND2 (N1946, N1935, N236);
nand NAND3 (N1947, N1928, N381, N776);
and AND3 (N1948, N1947, N465, N22);
and AND2 (N1949, N1946, N1856);
nand NAND3 (N1950, N1923, N352, N1337);
or OR4 (N1951, N1941, N910, N1732, N435);
xor XOR2 (N1952, N1940, N564);
xor XOR2 (N1953, N1930, N288);
not NOT1 (N1954, N1942);
or OR2 (N1955, N1944, N1929);
and AND3 (N1956, N1949, N6, N1402);
xor XOR2 (N1957, N1956, N942);
and AND4 (N1958, N1957, N1507, N943, N496);
xor XOR2 (N1959, N1951, N69);
xor XOR2 (N1960, N1954, N469);
and AND4 (N1961, N1959, N705, N822, N786);
nor NOR3 (N1962, N1950, N1574, N602);
buf BUF1 (N1963, N1962);
xor XOR2 (N1964, N1960, N639);
or OR4 (N1965, N1961, N1038, N950, N189);
buf BUF1 (N1966, N1939);
nor NOR2 (N1967, N1965, N908);
nand NAND2 (N1968, N1964, N967);
nor NOR4 (N1969, N1948, N1097, N685, N1655);
not NOT1 (N1970, N1966);
buf BUF1 (N1971, N1958);
or OR3 (N1972, N1970, N752, N1499);
buf BUF1 (N1973, N1967);
xor XOR2 (N1974, N1963, N1043);
and AND3 (N1975, N1953, N1499, N818);
nand NAND4 (N1976, N1969, N1573, N1685, N669);
nand NAND4 (N1977, N1971, N1644, N660, N1966);
and AND3 (N1978, N1976, N1367, N1658);
buf BUF1 (N1979, N1978);
not NOT1 (N1980, N1952);
or OR2 (N1981, N1955, N1839);
xor XOR2 (N1982, N1945, N1724);
and AND4 (N1983, N1977, N1014, N141, N914);
or OR3 (N1984, N1980, N987, N509);
or OR2 (N1985, N1983, N1616);
or OR3 (N1986, N1982, N235, N79);
nor NOR2 (N1987, N1984, N1052);
nand NAND3 (N1988, N1986, N485, N107);
and AND4 (N1989, N1987, N1055, N1201, N1766);
and AND4 (N1990, N1975, N1796, N735, N1329);
and AND4 (N1991, N1981, N326, N1642, N1235);
and AND3 (N1992, N1972, N1331, N1744);
nand NAND4 (N1993, N1974, N971, N1854, N941);
xor XOR2 (N1994, N1993, N422);
or OR3 (N1995, N1989, N1737, N1880);
nor NOR3 (N1996, N1991, N246, N658);
and AND3 (N1997, N1968, N1555, N1270);
not NOT1 (N1998, N1994);
nand NAND3 (N1999, N1992, N1766, N1467);
and AND3 (N2000, N1979, N1106, N1514);
not NOT1 (N2001, N1999);
nor NOR2 (N2002, N1996, N208);
or OR2 (N2003, N2000, N931);
and AND2 (N2004, N1997, N718);
nor NOR4 (N2005, N1985, N1491, N159, N1162);
and AND2 (N2006, N1988, N973);
buf BUF1 (N2007, N2006);
buf BUF1 (N2008, N2002);
buf BUF1 (N2009, N1995);
xor XOR2 (N2010, N1998, N68);
nor NOR4 (N2011, N1973, N1672, N957, N159);
not NOT1 (N2012, N1990);
xor XOR2 (N2013, N2001, N1685);
or OR4 (N2014, N2011, N430, N846, N710);
xor XOR2 (N2015, N2013, N370);
buf BUF1 (N2016, N2009);
nand NAND2 (N2017, N2007, N845);
buf BUF1 (N2018, N2016);
and AND4 (N2019, N2014, N1278, N769, N1267);
and AND2 (N2020, N2003, N636);
nand NAND3 (N2021, N2004, N1482, N1913);
and AND2 (N2022, N2021, N1613);
and AND2 (N2023, N2010, N131);
nor NOR2 (N2024, N2020, N1974);
xor XOR2 (N2025, N2015, N689);
not NOT1 (N2026, N2022);
and AND3 (N2027, N2005, N706, N342);
xor XOR2 (N2028, N2012, N234);
or OR2 (N2029, N2027, N927);
xor XOR2 (N2030, N2019, N272);
nand NAND4 (N2031, N2025, N347, N1950, N376);
buf BUF1 (N2032, N2026);
xor XOR2 (N2033, N2008, N1507);
and AND4 (N2034, N2018, N1742, N1776, N2025);
or OR2 (N2035, N2029, N1507);
or OR3 (N2036, N2033, N620, N1984);
not NOT1 (N2037, N2032);
nor NOR4 (N2038, N2037, N1301, N1251, N1358);
buf BUF1 (N2039, N2030);
or OR2 (N2040, N2023, N941);
nand NAND3 (N2041, N2028, N538, N747);
buf BUF1 (N2042, N2041);
and AND4 (N2043, N2035, N359, N1430, N1139);
and AND2 (N2044, N2036, N1358);
nor NOR2 (N2045, N2024, N688);
and AND4 (N2046, N2044, N984, N1322, N715);
not NOT1 (N2047, N2034);
not NOT1 (N2048, N2031);
nand NAND3 (N2049, N2038, N1019, N1903);
nand NAND3 (N2050, N2046, N1103, N1865);
and AND3 (N2051, N2050, N686, N625);
xor XOR2 (N2052, N2045, N687);
xor XOR2 (N2053, N2042, N1793);
not NOT1 (N2054, N2039);
xor XOR2 (N2055, N2051, N1899);
or OR4 (N2056, N2054, N2007, N2041, N1652);
buf BUF1 (N2057, N2048);
nor NOR4 (N2058, N2047, N693, N1446, N625);
and AND2 (N2059, N2057, N1251);
nor NOR4 (N2060, N2056, N1109, N1067, N1287);
xor XOR2 (N2061, N2059, N1004);
and AND3 (N2062, N2053, N1176, N1224);
xor XOR2 (N2063, N2052, N1586);
not NOT1 (N2064, N2055);
nand NAND4 (N2065, N2049, N826, N940, N977);
xor XOR2 (N2066, N2040, N65);
or OR4 (N2067, N2062, N48, N1050, N269);
nand NAND2 (N2068, N2064, N2045);
and AND4 (N2069, N2017, N413, N1267, N1006);
or OR4 (N2070, N2058, N712, N1970, N178);
nor NOR4 (N2071, N2065, N373, N755, N208);
buf BUF1 (N2072, N2067);
and AND2 (N2073, N2071, N1606);
and AND4 (N2074, N2068, N494, N1254, N789);
nor NOR3 (N2075, N2069, N124, N1246);
nor NOR3 (N2076, N2061, N1763, N1398);
and AND4 (N2077, N2066, N444, N1101, N1398);
xor XOR2 (N2078, N2077, N2020);
nand NAND4 (N2079, N2076, N959, N145, N40);
nand NAND3 (N2080, N2043, N444, N1260);
and AND3 (N2081, N2078, N272, N1172);
buf BUF1 (N2082, N2063);
buf BUF1 (N2083, N2073);
nor NOR3 (N2084, N2074, N1244, N1292);
not NOT1 (N2085, N2082);
not NOT1 (N2086, N2075);
and AND2 (N2087, N2085, N1499);
xor XOR2 (N2088, N2086, N156);
nor NOR3 (N2089, N2084, N1677, N276);
and AND3 (N2090, N2060, N797, N1737);
xor XOR2 (N2091, N2089, N1129);
or OR2 (N2092, N2083, N1508);
not NOT1 (N2093, N2092);
nand NAND3 (N2094, N2072, N467, N688);
or OR4 (N2095, N2094, N742, N1193, N81);
xor XOR2 (N2096, N2095, N1749);
nand NAND4 (N2097, N2081, N595, N1647, N436);
not NOT1 (N2098, N2097);
not NOT1 (N2099, N2093);
nand NAND2 (N2100, N2079, N958);
xor XOR2 (N2101, N2087, N1613);
or OR2 (N2102, N2080, N1955);
and AND3 (N2103, N2100, N406, N1591);
not NOT1 (N2104, N2096);
not NOT1 (N2105, N2101);
or OR3 (N2106, N2098, N1313, N2010);
not NOT1 (N2107, N2105);
xor XOR2 (N2108, N2103, N1649);
nand NAND3 (N2109, N2107, N984, N1784);
xor XOR2 (N2110, N2106, N509);
nor NOR2 (N2111, N2091, N1974);
and AND4 (N2112, N2109, N501, N522, N992);
and AND3 (N2113, N2088, N1069, N1672);
nand NAND2 (N2114, N2090, N982);
and AND4 (N2115, N2099, N399, N700, N1290);
xor XOR2 (N2116, N2110, N1944);
nor NOR2 (N2117, N2112, N426);
not NOT1 (N2118, N2116);
or OR2 (N2119, N2117, N226);
nand NAND3 (N2120, N2104, N143, N127);
nor NOR2 (N2121, N2113, N1350);
nor NOR2 (N2122, N2115, N422);
nor NOR3 (N2123, N2120, N649, N1457);
buf BUF1 (N2124, N2119);
and AND4 (N2125, N2114, N1484, N2062, N849);
nor NOR2 (N2126, N2125, N622);
or OR2 (N2127, N2123, N1410);
nor NOR2 (N2128, N2121, N415);
nor NOR2 (N2129, N2122, N2122);
and AND3 (N2130, N2070, N1517, N45);
buf BUF1 (N2131, N2128);
or OR4 (N2132, N2124, N612, N348, N1454);
xor XOR2 (N2133, N2129, N349);
nor NOR4 (N2134, N2130, N1684, N834, N1324);
nand NAND3 (N2135, N2127, N1428, N851);
xor XOR2 (N2136, N2135, N1226);
buf BUF1 (N2137, N2131);
nor NOR4 (N2138, N2118, N1444, N1629, N1877);
and AND2 (N2139, N2102, N1629);
buf BUF1 (N2140, N2138);
nor NOR2 (N2141, N2111, N2104);
not NOT1 (N2142, N2132);
nor NOR4 (N2143, N2133, N405, N662, N1097);
nor NOR2 (N2144, N2142, N1581);
buf BUF1 (N2145, N2134);
buf BUF1 (N2146, N2136);
nor NOR3 (N2147, N2139, N1609, N1598);
or OR2 (N2148, N2108, N150);
buf BUF1 (N2149, N2140);
and AND3 (N2150, N2126, N408, N1752);
nand NAND2 (N2151, N2143, N525);
and AND2 (N2152, N2149, N1068);
xor XOR2 (N2153, N2145, N1250);
or OR3 (N2154, N2147, N1399, N1809);
buf BUF1 (N2155, N2153);
and AND2 (N2156, N2155, N1751);
or OR2 (N2157, N2150, N1424);
or OR4 (N2158, N2144, N1723, N85, N1429);
not NOT1 (N2159, N2148);
buf BUF1 (N2160, N2154);
not NOT1 (N2161, N2158);
not NOT1 (N2162, N2151);
nand NAND3 (N2163, N2137, N2001, N31);
nand NAND3 (N2164, N2156, N1111, N712);
xor XOR2 (N2165, N2157, N887);
xor XOR2 (N2166, N2162, N547);
and AND3 (N2167, N2146, N1148, N2123);
or OR2 (N2168, N2161, N867);
nand NAND2 (N2169, N2166, N71);
or OR3 (N2170, N2168, N1290, N763);
not NOT1 (N2171, N2160);
xor XOR2 (N2172, N2141, N1463);
or OR3 (N2173, N2165, N1456, N464);
or OR4 (N2174, N2163, N2101, N1235, N1899);
nor NOR2 (N2175, N2170, N1324);
nor NOR4 (N2176, N2159, N1411, N1749, N1019);
buf BUF1 (N2177, N2167);
not NOT1 (N2178, N2177);
buf BUF1 (N2179, N2171);
not NOT1 (N2180, N2174);
buf BUF1 (N2181, N2169);
nor NOR3 (N2182, N2180, N1230, N1201);
xor XOR2 (N2183, N2182, N282);
nand NAND4 (N2184, N2172, N1592, N1983, N1095);
not NOT1 (N2185, N2184);
and AND3 (N2186, N2183, N927, N1784);
nand NAND3 (N2187, N2186, N1430, N2121);
xor XOR2 (N2188, N2179, N1592);
buf BUF1 (N2189, N2176);
and AND4 (N2190, N2188, N1241, N1774, N1871);
xor XOR2 (N2191, N2190, N962);
nor NOR3 (N2192, N2185, N1628, N865);
buf BUF1 (N2193, N2189);
nand NAND4 (N2194, N2192, N38, N1024, N503);
xor XOR2 (N2195, N2178, N1617);
and AND3 (N2196, N2164, N1615, N234);
nand NAND2 (N2197, N2193, N1607);
nor NOR4 (N2198, N2173, N707, N1652, N1549);
xor XOR2 (N2199, N2198, N1620);
and AND3 (N2200, N2194, N1969, N1387);
xor XOR2 (N2201, N2195, N1232);
xor XOR2 (N2202, N2152, N1041);
nand NAND4 (N2203, N2196, N1500, N875, N220);
not NOT1 (N2204, N2199);
nor NOR2 (N2205, N2197, N1854);
nor NOR2 (N2206, N2204, N1305);
and AND2 (N2207, N2202, N1291);
and AND2 (N2208, N2207, N1668);
not NOT1 (N2209, N2206);
or OR4 (N2210, N2203, N1286, N1142, N1973);
nor NOR4 (N2211, N2181, N730, N745, N105);
xor XOR2 (N2212, N2200, N96);
nor NOR3 (N2213, N2175, N1972, N2051);
not NOT1 (N2214, N2212);
not NOT1 (N2215, N2214);
or OR3 (N2216, N2187, N1024, N869);
nand NAND2 (N2217, N2205, N1401);
not NOT1 (N2218, N2201);
xor XOR2 (N2219, N2191, N544);
nor NOR3 (N2220, N2211, N2199, N1758);
or OR2 (N2221, N2209, N673);
or OR4 (N2222, N2221, N95, N312, N1912);
nor NOR2 (N2223, N2208, N983);
xor XOR2 (N2224, N2213, N1240);
buf BUF1 (N2225, N2210);
or OR2 (N2226, N2222, N1653);
or OR4 (N2227, N2226, N1186, N1160, N634);
and AND3 (N2228, N2223, N581, N221);
or OR3 (N2229, N2217, N546, N2180);
or OR2 (N2230, N2219, N717);
buf BUF1 (N2231, N2224);
nand NAND2 (N2232, N2218, N1742);
or OR2 (N2233, N2225, N442);
nand NAND4 (N2234, N2232, N1973, N2105, N1555);
buf BUF1 (N2235, N2230);
buf BUF1 (N2236, N2235);
xor XOR2 (N2237, N2231, N1550);
xor XOR2 (N2238, N2229, N1903);
xor XOR2 (N2239, N2236, N488);
nand NAND2 (N2240, N2234, N1506);
buf BUF1 (N2241, N2228);
and AND3 (N2242, N2241, N235, N30);
not NOT1 (N2243, N2237);
not NOT1 (N2244, N2216);
or OR2 (N2245, N2220, N1766);
or OR2 (N2246, N2215, N2155);
nand NAND3 (N2247, N2238, N342, N2246);
nor NOR4 (N2248, N61, N589, N775, N1624);
or OR4 (N2249, N2233, N1684, N671, N1576);
nand NAND4 (N2250, N2247, N1379, N1214, N2205);
or OR3 (N2251, N2242, N221, N2020);
not NOT1 (N2252, N2244);
not NOT1 (N2253, N2250);
not NOT1 (N2254, N2243);
or OR3 (N2255, N2253, N905, N1926);
and AND4 (N2256, N2227, N1135, N1582, N1158);
nand NAND3 (N2257, N2252, N950, N2148);
xor XOR2 (N2258, N2245, N1876);
buf BUF1 (N2259, N2254);
and AND3 (N2260, N2259, N851, N923);
nand NAND2 (N2261, N2256, N1573);
buf BUF1 (N2262, N2261);
xor XOR2 (N2263, N2255, N403);
xor XOR2 (N2264, N2263, N1633);
and AND3 (N2265, N2239, N861, N152);
buf BUF1 (N2266, N2258);
or OR2 (N2267, N2265, N1763);
not NOT1 (N2268, N2248);
buf BUF1 (N2269, N2262);
nand NAND4 (N2270, N2268, N1535, N1892, N591);
and AND3 (N2271, N2249, N533, N1544);
nor NOR3 (N2272, N2251, N1421, N673);
nand NAND4 (N2273, N2264, N1323, N1187, N1128);
and AND3 (N2274, N2240, N2128, N324);
xor XOR2 (N2275, N2267, N2117);
nand NAND4 (N2276, N2266, N2147, N1073, N1747);
not NOT1 (N2277, N2260);
nor NOR4 (N2278, N2274, N976, N1419, N1608);
nor NOR3 (N2279, N2277, N941, N1198);
xor XOR2 (N2280, N2272, N1923);
xor XOR2 (N2281, N2280, N125);
nor NOR2 (N2282, N2276, N1848);
not NOT1 (N2283, N2271);
buf BUF1 (N2284, N2273);
xor XOR2 (N2285, N2270, N1668);
buf BUF1 (N2286, N2275);
nand NAND3 (N2287, N2257, N1618, N1911);
nand NAND3 (N2288, N2286, N2130, N576);
xor XOR2 (N2289, N2288, N1437);
nor NOR3 (N2290, N2278, N692, N1419);
nor NOR2 (N2291, N2285, N896);
buf BUF1 (N2292, N2290);
not NOT1 (N2293, N2282);
nor NOR4 (N2294, N2287, N645, N547, N2212);
and AND3 (N2295, N2279, N1547, N2257);
not NOT1 (N2296, N2281);
nand NAND2 (N2297, N2295, N1959);
xor XOR2 (N2298, N2292, N1149);
and AND4 (N2299, N2283, N1825, N355, N1329);
xor XOR2 (N2300, N2296, N2223);
nand NAND4 (N2301, N2293, N942, N2072, N1211);
nand NAND4 (N2302, N2294, N1167, N1496, N1594);
nor NOR3 (N2303, N2269, N310, N1794);
or OR3 (N2304, N2297, N2161, N1643);
or OR3 (N2305, N2301, N2292, N1317);
buf BUF1 (N2306, N2305);
and AND2 (N2307, N2284, N837);
nor NOR3 (N2308, N2289, N370, N125);
xor XOR2 (N2309, N2308, N144);
or OR4 (N2310, N2298, N1092, N984, N1208);
not NOT1 (N2311, N2306);
or OR2 (N2312, N2302, N399);
nand NAND4 (N2313, N2304, N42, N1505, N2061);
nor NOR4 (N2314, N2291, N1844, N122, N1728);
buf BUF1 (N2315, N2300);
nor NOR3 (N2316, N2314, N1258, N1682);
nor NOR3 (N2317, N2313, N983, N310);
not NOT1 (N2318, N2299);
and AND2 (N2319, N2315, N1205);
nor NOR3 (N2320, N2317, N62, N577);
or OR2 (N2321, N2303, N1191);
buf BUF1 (N2322, N2320);
or OR4 (N2323, N2319, N1046, N262, N2240);
and AND3 (N2324, N2311, N1855, N1706);
and AND2 (N2325, N2312, N1181);
buf BUF1 (N2326, N2318);
nor NOR2 (N2327, N2325, N1413);
and AND4 (N2328, N2321, N1451, N1488, N2287);
buf BUF1 (N2329, N2316);
xor XOR2 (N2330, N2322, N1923);
and AND2 (N2331, N2307, N1415);
nor NOR3 (N2332, N2329, N2053, N1619);
xor XOR2 (N2333, N2332, N1074);
xor XOR2 (N2334, N2324, N1606);
xor XOR2 (N2335, N2331, N697);
nand NAND3 (N2336, N2330, N197, N2275);
not NOT1 (N2337, N2328);
buf BUF1 (N2338, N2334);
and AND2 (N2339, N2336, N1789);
and AND3 (N2340, N2333, N1077, N928);
buf BUF1 (N2341, N2335);
xor XOR2 (N2342, N2310, N564);
nand NAND4 (N2343, N2338, N551, N199, N1189);
not NOT1 (N2344, N2340);
nor NOR4 (N2345, N2339, N1902, N147, N1665);
buf BUF1 (N2346, N2342);
nor NOR3 (N2347, N2345, N426, N912);
not NOT1 (N2348, N2323);
or OR2 (N2349, N2309, N2325);
nor NOR3 (N2350, N2337, N1948, N2321);
not NOT1 (N2351, N2348);
buf BUF1 (N2352, N2347);
xor XOR2 (N2353, N2349, N2029);
buf BUF1 (N2354, N2351);
nand NAND4 (N2355, N2350, N187, N1853, N68);
nand NAND3 (N2356, N2327, N2002, N1208);
or OR3 (N2357, N2326, N2041, N1709);
xor XOR2 (N2358, N2346, N1377);
buf BUF1 (N2359, N2356);
buf BUF1 (N2360, N2357);
nand NAND3 (N2361, N2359, N1933, N1531);
nand NAND3 (N2362, N2361, N2054, N845);
xor XOR2 (N2363, N2358, N705);
nand NAND4 (N2364, N2343, N533, N1238, N2075);
buf BUF1 (N2365, N2353);
and AND2 (N2366, N2354, N1630);
buf BUF1 (N2367, N2344);
xor XOR2 (N2368, N2366, N1001);
buf BUF1 (N2369, N2341);
nand NAND2 (N2370, N2352, N2238);
buf BUF1 (N2371, N2363);
xor XOR2 (N2372, N2355, N610);
nor NOR2 (N2373, N2364, N1303);
or OR3 (N2374, N2368, N1490, N282);
buf BUF1 (N2375, N2367);
or OR3 (N2376, N2372, N1980, N1134);
nand NAND4 (N2377, N2373, N410, N478, N2030);
or OR3 (N2378, N2374, N171, N1660);
buf BUF1 (N2379, N2369);
xor XOR2 (N2380, N2371, N817);
xor XOR2 (N2381, N2362, N526);
buf BUF1 (N2382, N2360);
buf BUF1 (N2383, N2377);
nand NAND4 (N2384, N2379, N711, N116, N2074);
xor XOR2 (N2385, N2376, N953);
not NOT1 (N2386, N2385);
and AND3 (N2387, N2382, N1504, N1356);
nor NOR4 (N2388, N2380, N330, N1104, N1959);
and AND2 (N2389, N2383, N1133);
nand NAND2 (N2390, N2387, N410);
and AND3 (N2391, N2389, N1853, N965);
buf BUF1 (N2392, N2384);
and AND4 (N2393, N2375, N1200, N1990, N1670);
or OR4 (N2394, N2381, N1243, N789, N402);
and AND2 (N2395, N2386, N88);
and AND3 (N2396, N2370, N1699, N904);
or OR4 (N2397, N2393, N392, N820, N553);
not NOT1 (N2398, N2395);
nand NAND3 (N2399, N2397, N1273, N20);
nor NOR2 (N2400, N2378, N1476);
not NOT1 (N2401, N2365);
nor NOR3 (N2402, N2390, N1755, N740);
nor NOR4 (N2403, N2400, N2181, N1729, N1700);
xor XOR2 (N2404, N2402, N261);
and AND3 (N2405, N2401, N178, N97);
xor XOR2 (N2406, N2396, N489);
buf BUF1 (N2407, N2394);
or OR3 (N2408, N2388, N1527, N1349);
nor NOR2 (N2409, N2392, N2264);
not NOT1 (N2410, N2408);
nand NAND3 (N2411, N2403, N1659, N2243);
buf BUF1 (N2412, N2399);
xor XOR2 (N2413, N2412, N807);
xor XOR2 (N2414, N2398, N1765);
xor XOR2 (N2415, N2409, N935);
xor XOR2 (N2416, N2407, N17);
buf BUF1 (N2417, N2415);
xor XOR2 (N2418, N2417, N1216);
not NOT1 (N2419, N2410);
nand NAND4 (N2420, N2391, N296, N502, N2354);
or OR2 (N2421, N2406, N2092);
not NOT1 (N2422, N2414);
buf BUF1 (N2423, N2419);
buf BUF1 (N2424, N2411);
buf BUF1 (N2425, N2418);
buf BUF1 (N2426, N2421);
xor XOR2 (N2427, N2416, N681);
nor NOR4 (N2428, N2405, N2189, N2044, N232);
and AND4 (N2429, N2404, N594, N779, N214);
not NOT1 (N2430, N2422);
nor NOR4 (N2431, N2420, N1212, N2106, N1364);
and AND4 (N2432, N2424, N1509, N1684, N1478);
xor XOR2 (N2433, N2430, N886);
or OR3 (N2434, N2431, N536, N982);
xor XOR2 (N2435, N2425, N2303);
not NOT1 (N2436, N2433);
nor NOR4 (N2437, N2432, N151, N1106, N643);
xor XOR2 (N2438, N2434, N414);
or OR3 (N2439, N2435, N1028, N603);
and AND2 (N2440, N2437, N328);
xor XOR2 (N2441, N2429, N138);
buf BUF1 (N2442, N2423);
buf BUF1 (N2443, N2441);
and AND3 (N2444, N2438, N1050, N1700);
or OR4 (N2445, N2426, N402, N390, N1767);
not NOT1 (N2446, N2440);
nor NOR2 (N2447, N2428, N625);
or OR3 (N2448, N2444, N1188, N286);
not NOT1 (N2449, N2447);
or OR3 (N2450, N2445, N1647, N2437);
nor NOR2 (N2451, N2436, N741);
and AND2 (N2452, N2427, N106);
or OR3 (N2453, N2448, N2133, N1341);
or OR3 (N2454, N2452, N2056, N895);
nand NAND2 (N2455, N2451, N4);
not NOT1 (N2456, N2413);
not NOT1 (N2457, N2456);
buf BUF1 (N2458, N2453);
or OR3 (N2459, N2454, N1527, N1628);
nor NOR3 (N2460, N2446, N1484, N334);
nor NOR3 (N2461, N2458, N11, N1953);
buf BUF1 (N2462, N2459);
buf BUF1 (N2463, N2450);
xor XOR2 (N2464, N2455, N1289);
nand NAND3 (N2465, N2461, N1123, N1432);
not NOT1 (N2466, N2460);
or OR4 (N2467, N2466, N2301, N2055, N1634);
nor NOR2 (N2468, N2467, N46);
nand NAND2 (N2469, N2442, N1335);
not NOT1 (N2470, N2463);
or OR4 (N2471, N2464, N1378, N647, N2408);
nor NOR2 (N2472, N2470, N2054);
nor NOR3 (N2473, N2449, N57, N1182);
nand NAND2 (N2474, N2469, N1819);
buf BUF1 (N2475, N2471);
buf BUF1 (N2476, N2474);
nor NOR3 (N2477, N2476, N486, N808);
nand NAND2 (N2478, N2472, N534);
nand NAND4 (N2479, N2462, N2312, N2392, N595);
and AND3 (N2480, N2457, N2435, N570);
buf BUF1 (N2481, N2479);
nand NAND2 (N2482, N2473, N623);
not NOT1 (N2483, N2482);
nand NAND3 (N2484, N2475, N2195, N702);
nor NOR3 (N2485, N2484, N609, N1864);
nor NOR3 (N2486, N2485, N608, N2229);
and AND2 (N2487, N2439, N753);
and AND3 (N2488, N2478, N2459, N1247);
nor NOR2 (N2489, N2468, N885);
and AND4 (N2490, N2465, N707, N722, N1034);
not NOT1 (N2491, N2477);
xor XOR2 (N2492, N2488, N1872);
not NOT1 (N2493, N2491);
not NOT1 (N2494, N2483);
nor NOR4 (N2495, N2494, N2019, N399, N2228);
nor NOR2 (N2496, N2490, N1067);
xor XOR2 (N2497, N2443, N1802);
or OR2 (N2498, N2486, N649);
nand NAND4 (N2499, N2489, N32, N2208, N12);
buf BUF1 (N2500, N2481);
nand NAND4 (N2501, N2497, N114, N1087, N1443);
or OR3 (N2502, N2500, N651, N1347);
xor XOR2 (N2503, N2502, N605);
buf BUF1 (N2504, N2480);
nor NOR2 (N2505, N2493, N1101);
or OR3 (N2506, N2498, N325, N2024);
nand NAND4 (N2507, N2496, N1474, N821, N1550);
xor XOR2 (N2508, N2499, N837);
xor XOR2 (N2509, N2492, N988);
or OR4 (N2510, N2501, N984, N117, N1731);
or OR2 (N2511, N2487, N306);
not NOT1 (N2512, N2511);
and AND4 (N2513, N2510, N39, N1171, N514);
nand NAND4 (N2514, N2505, N2165, N1195, N2421);
nor NOR4 (N2515, N2508, N930, N1941, N1977);
buf BUF1 (N2516, N2503);
nand NAND3 (N2517, N2504, N1188, N539);
nor NOR4 (N2518, N2514, N1421, N986, N545);
or OR2 (N2519, N2506, N361);
not NOT1 (N2520, N2518);
buf BUF1 (N2521, N2517);
or OR3 (N2522, N2509, N2026, N1670);
xor XOR2 (N2523, N2495, N827);
nand NAND3 (N2524, N2520, N977, N184);
or OR2 (N2525, N2524, N1133);
nor NOR4 (N2526, N2507, N2083, N1237, N2316);
buf BUF1 (N2527, N2521);
not NOT1 (N2528, N2523);
and AND4 (N2529, N2515, N2393, N699, N1373);
nor NOR4 (N2530, N2513, N2123, N1818, N151);
or OR3 (N2531, N2525, N1532, N1007);
nor NOR2 (N2532, N2526, N1616);
and AND4 (N2533, N2528, N152, N172, N1918);
nor NOR2 (N2534, N2533, N1576);
or OR3 (N2535, N2519, N711, N1547);
nand NAND4 (N2536, N2530, N1483, N1422, N1004);
xor XOR2 (N2537, N2527, N719);
buf BUF1 (N2538, N2537);
not NOT1 (N2539, N2535);
and AND2 (N2540, N2532, N197);
buf BUF1 (N2541, N2531);
nor NOR4 (N2542, N2541, N2413, N985, N429);
buf BUF1 (N2543, N2522);
nand NAND2 (N2544, N2534, N2380);
nor NOR4 (N2545, N2540, N2500, N1998, N2363);
not NOT1 (N2546, N2542);
buf BUF1 (N2547, N2529);
not NOT1 (N2548, N2516);
xor XOR2 (N2549, N2548, N2211);
nor NOR2 (N2550, N2539, N2516);
nand NAND4 (N2551, N2547, N2492, N1193, N172);
buf BUF1 (N2552, N2543);
xor XOR2 (N2553, N2512, N1828);
or OR4 (N2554, N2544, N758, N1767, N1153);
nand NAND2 (N2555, N2554, N628);
and AND2 (N2556, N2536, N71);
nand NAND2 (N2557, N2552, N1205);
not NOT1 (N2558, N2538);
nand NAND4 (N2559, N2545, N986, N1689, N2019);
or OR3 (N2560, N2559, N1399, N1554);
xor XOR2 (N2561, N2550, N1081);
and AND2 (N2562, N2557, N1548);
nor NOR4 (N2563, N2556, N2328, N1652, N2530);
and AND2 (N2564, N2560, N861);
and AND2 (N2565, N2561, N1414);
nand NAND3 (N2566, N2565, N984, N492);
nor NOR3 (N2567, N2558, N444, N400);
buf BUF1 (N2568, N2566);
xor XOR2 (N2569, N2563, N2484);
xor XOR2 (N2570, N2569, N87);
and AND4 (N2571, N2562, N1882, N1391, N2518);
and AND2 (N2572, N2567, N606);
not NOT1 (N2573, N2551);
nand NAND3 (N2574, N2555, N820, N760);
not NOT1 (N2575, N2553);
nor NOR2 (N2576, N2570, N1772);
xor XOR2 (N2577, N2546, N1916);
nor NOR4 (N2578, N2577, N1439, N1596, N2276);
nor NOR4 (N2579, N2578, N1629, N2285, N508);
and AND4 (N2580, N2564, N281, N1703, N2367);
not NOT1 (N2581, N2580);
not NOT1 (N2582, N2576);
not NOT1 (N2583, N2579);
buf BUF1 (N2584, N2568);
not NOT1 (N2585, N2575);
nor NOR3 (N2586, N2584, N1259, N1453);
or OR2 (N2587, N2582, N1091);
buf BUF1 (N2588, N2549);
nand NAND2 (N2589, N2571, N1229);
buf BUF1 (N2590, N2589);
and AND4 (N2591, N2587, N2222, N201, N2322);
not NOT1 (N2592, N2574);
buf BUF1 (N2593, N2581);
or OR4 (N2594, N2585, N986, N790, N605);
not NOT1 (N2595, N2591);
not NOT1 (N2596, N2586);
nor NOR3 (N2597, N2590, N127, N1972);
and AND2 (N2598, N2588, N472);
xor XOR2 (N2599, N2593, N1724);
buf BUF1 (N2600, N2583);
or OR3 (N2601, N2592, N1749, N1259);
or OR3 (N2602, N2573, N1619, N1841);
or OR3 (N2603, N2597, N482, N2197);
nor NOR2 (N2604, N2572, N2370);
or OR3 (N2605, N2594, N752, N86);
nand NAND2 (N2606, N2603, N812);
buf BUF1 (N2607, N2602);
nor NOR2 (N2608, N2600, N174);
not NOT1 (N2609, N2607);
or OR3 (N2610, N2601, N1808, N405);
not NOT1 (N2611, N2609);
nand NAND2 (N2612, N2610, N199);
and AND2 (N2613, N2595, N875);
nand NAND4 (N2614, N2598, N258, N2398, N2271);
xor XOR2 (N2615, N2608, N2210);
not NOT1 (N2616, N2596);
nand NAND3 (N2617, N2614, N2500, N2011);
xor XOR2 (N2618, N2612, N1499);
and AND3 (N2619, N2606, N952, N1);
not NOT1 (N2620, N2616);
xor XOR2 (N2621, N2599, N160);
not NOT1 (N2622, N2613);
nand NAND3 (N2623, N2622, N779, N1029);
not NOT1 (N2624, N2611);
or OR4 (N2625, N2621, N1724, N2535, N2286);
nand NAND2 (N2626, N2624, N1592);
and AND3 (N2627, N2618, N1246, N1495);
nand NAND4 (N2628, N2620, N2308, N417, N340);
and AND3 (N2629, N2623, N135, N2414);
not NOT1 (N2630, N2627);
buf BUF1 (N2631, N2617);
buf BUF1 (N2632, N2604);
buf BUF1 (N2633, N2619);
nor NOR2 (N2634, N2632, N2441);
xor XOR2 (N2635, N2629, N379);
xor XOR2 (N2636, N2605, N1938);
xor XOR2 (N2637, N2615, N1883);
xor XOR2 (N2638, N2633, N1638);
not NOT1 (N2639, N2628);
or OR2 (N2640, N2625, N1030);
and AND2 (N2641, N2636, N225);
xor XOR2 (N2642, N2626, N1962);
nand NAND3 (N2643, N2631, N1715, N1690);
nor NOR2 (N2644, N2634, N2175);
not NOT1 (N2645, N2644);
xor XOR2 (N2646, N2630, N375);
or OR3 (N2647, N2639, N347, N617);
nor NOR4 (N2648, N2641, N906, N105, N2152);
or OR2 (N2649, N2646, N436);
nand NAND4 (N2650, N2643, N2528, N754, N1855);
nor NOR3 (N2651, N2635, N2630, N654);
buf BUF1 (N2652, N2647);
and AND2 (N2653, N2638, N836);
or OR4 (N2654, N2652, N1591, N700, N945);
buf BUF1 (N2655, N2650);
xor XOR2 (N2656, N2642, N450);
and AND4 (N2657, N2648, N2226, N1957, N2522);
not NOT1 (N2658, N2656);
nor NOR4 (N2659, N2657, N1543, N572, N527);
buf BUF1 (N2660, N2649);
and AND3 (N2661, N2658, N2429, N2403);
or OR3 (N2662, N2640, N1531, N836);
buf BUF1 (N2663, N2645);
nor NOR2 (N2664, N2655, N2228);
xor XOR2 (N2665, N2661, N2032);
nor NOR4 (N2666, N2665, N547, N979, N2034);
nand NAND3 (N2667, N2651, N1149, N68);
nor NOR4 (N2668, N2660, N840, N2172, N2113);
nand NAND3 (N2669, N2654, N2287, N388);
nor NOR4 (N2670, N2669, N1545, N1620, N2647);
nand NAND2 (N2671, N2668, N2601);
nor NOR3 (N2672, N2637, N1950, N1375);
nand NAND4 (N2673, N2662, N1553, N1056, N2021);
xor XOR2 (N2674, N2673, N2633);
not NOT1 (N2675, N2659);
nand NAND4 (N2676, N2670, N2452, N86, N1485);
buf BUF1 (N2677, N2663);
xor XOR2 (N2678, N2674, N1607);
not NOT1 (N2679, N2676);
or OR2 (N2680, N2664, N1487);
xor XOR2 (N2681, N2653, N339);
xor XOR2 (N2682, N2679, N1864);
nand NAND2 (N2683, N2675, N1470);
nor NOR3 (N2684, N2682, N579, N1921);
and AND2 (N2685, N2667, N810);
or OR3 (N2686, N2677, N1593, N1493);
and AND4 (N2687, N2671, N849, N65, N2370);
buf BUF1 (N2688, N2684);
xor XOR2 (N2689, N2678, N2549);
nor NOR2 (N2690, N2685, N2616);
nor NOR2 (N2691, N2686, N1968);
or OR2 (N2692, N2672, N1388);
not NOT1 (N2693, N2688);
not NOT1 (N2694, N2666);
buf BUF1 (N2695, N2694);
xor XOR2 (N2696, N2681, N2089);
nand NAND2 (N2697, N2692, N2321);
nor NOR4 (N2698, N2683, N1724, N2141, N1466);
nor NOR2 (N2699, N2696, N2410);
nand NAND4 (N2700, N2690, N812, N1326, N170);
not NOT1 (N2701, N2680);
not NOT1 (N2702, N2700);
nor NOR2 (N2703, N2693, N2365);
nor NOR3 (N2704, N2698, N2311, N147);
not NOT1 (N2705, N2701);
nor NOR3 (N2706, N2697, N2673, N1732);
xor XOR2 (N2707, N2689, N227);
and AND4 (N2708, N2704, N2272, N2015, N267);
nor NOR2 (N2709, N2691, N2245);
and AND4 (N2710, N2702, N2648, N588, N377);
or OR4 (N2711, N2708, N44, N1949, N2122);
nand NAND3 (N2712, N2709, N1601, N186);
or OR4 (N2713, N2706, N25, N1082, N423);
and AND2 (N2714, N2695, N1759);
not NOT1 (N2715, N2712);
not NOT1 (N2716, N2687);
buf BUF1 (N2717, N2710);
and AND2 (N2718, N2699, N812);
or OR4 (N2719, N2713, N1894, N1078, N1197);
nand NAND3 (N2720, N2711, N621, N1433);
buf BUF1 (N2721, N2717);
or OR2 (N2722, N2718, N2368);
and AND2 (N2723, N2720, N975);
nor NOR3 (N2724, N2719, N2382, N343);
nand NAND2 (N2725, N2714, N2333);
nand NAND3 (N2726, N2703, N1428, N2272);
xor XOR2 (N2727, N2724, N1782);
or OR3 (N2728, N2726, N2075, N797);
and AND3 (N2729, N2721, N1322, N71);
buf BUF1 (N2730, N2716);
xor XOR2 (N2731, N2729, N1689);
buf BUF1 (N2732, N2707);
xor XOR2 (N2733, N2731, N1721);
not NOT1 (N2734, N2723);
not NOT1 (N2735, N2722);
nand NAND3 (N2736, N2735, N594, N1669);
and AND3 (N2737, N2734, N985, N721);
xor XOR2 (N2738, N2727, N683);
nor NOR3 (N2739, N2732, N717, N1475);
xor XOR2 (N2740, N2733, N2308);
nand NAND3 (N2741, N2705, N2607, N1431);
nor NOR2 (N2742, N2738, N55);
xor XOR2 (N2743, N2715, N706);
xor XOR2 (N2744, N2730, N1962);
and AND4 (N2745, N2742, N1280, N1484, N2006);
and AND3 (N2746, N2728, N2478, N1934);
nand NAND2 (N2747, N2746, N1121);
not NOT1 (N2748, N2736);
or OR3 (N2749, N2743, N1036, N2148);
or OR2 (N2750, N2737, N1749);
nand NAND4 (N2751, N2744, N291, N549, N1193);
nand NAND4 (N2752, N2725, N938, N260, N485);
buf BUF1 (N2753, N2749);
xor XOR2 (N2754, N2748, N878);
not NOT1 (N2755, N2754);
or OR2 (N2756, N2739, N2406);
not NOT1 (N2757, N2753);
xor XOR2 (N2758, N2741, N1093);
buf BUF1 (N2759, N2755);
nand NAND4 (N2760, N2759, N496, N372, N1379);
buf BUF1 (N2761, N2747);
nor NOR4 (N2762, N2760, N1116, N1706, N1979);
xor XOR2 (N2763, N2752, N2242);
and AND4 (N2764, N2750, N2241, N2542, N463);
nand NAND4 (N2765, N2758, N1787, N1731, N1265);
nand NAND3 (N2766, N2756, N1066, N2073);
buf BUF1 (N2767, N2764);
xor XOR2 (N2768, N2767, N411);
not NOT1 (N2769, N2761);
nand NAND3 (N2770, N2740, N1661, N1985);
nor NOR3 (N2771, N2745, N2095, N451);
or OR3 (N2772, N2763, N1362, N965);
buf BUF1 (N2773, N2751);
or OR4 (N2774, N2766, N2496, N2533, N1661);
xor XOR2 (N2775, N2769, N2600);
nor NOR4 (N2776, N2757, N2733, N2503, N241);
buf BUF1 (N2777, N2768);
or OR3 (N2778, N2776, N1377, N3);
nor NOR4 (N2779, N2777, N587, N2209, N2336);
nand NAND2 (N2780, N2773, N2548);
buf BUF1 (N2781, N2762);
xor XOR2 (N2782, N2774, N389);
and AND3 (N2783, N2772, N677, N62);
nand NAND4 (N2784, N2765, N1354, N1909, N105);
nand NAND4 (N2785, N2770, N1580, N2049, N2207);
and AND4 (N2786, N2775, N673, N2006, N1872);
nand NAND3 (N2787, N2780, N2514, N917);
and AND2 (N2788, N2785, N762);
buf BUF1 (N2789, N2771);
xor XOR2 (N2790, N2784, N2545);
xor XOR2 (N2791, N2781, N1765);
nand NAND2 (N2792, N2786, N2512);
nor NOR4 (N2793, N2789, N2610, N1961, N663);
buf BUF1 (N2794, N2791);
and AND4 (N2795, N2783, N92, N2282, N1642);
xor XOR2 (N2796, N2779, N679);
or OR4 (N2797, N2782, N1743, N592, N393);
not NOT1 (N2798, N2794);
buf BUF1 (N2799, N2787);
or OR4 (N2800, N2797, N1792, N2197, N853);
nor NOR3 (N2801, N2795, N1470, N1578);
and AND3 (N2802, N2778, N2709, N963);
and AND2 (N2803, N2801, N2028);
nand NAND3 (N2804, N2796, N2708, N1570);
nand NAND4 (N2805, N2788, N1529, N573, N2724);
buf BUF1 (N2806, N2793);
not NOT1 (N2807, N2792);
or OR3 (N2808, N2807, N1166, N1768);
and AND3 (N2809, N2804, N2375, N1356);
xor XOR2 (N2810, N2805, N2657);
or OR3 (N2811, N2803, N2728, N2532);
or OR3 (N2812, N2808, N951, N492);
not NOT1 (N2813, N2811);
and AND4 (N2814, N2800, N2249, N546, N1911);
and AND3 (N2815, N2799, N2801, N2479);
and AND2 (N2816, N2809, N482);
not NOT1 (N2817, N2802);
or OR3 (N2818, N2812, N1810, N2225);
not NOT1 (N2819, N2818);
nand NAND3 (N2820, N2819, N2555, N1787);
nor NOR2 (N2821, N2820, N1383);
or OR3 (N2822, N2806, N1827, N1191);
nand NAND3 (N2823, N2821, N686, N1879);
nand NAND3 (N2824, N2823, N898, N331);
and AND4 (N2825, N2790, N2065, N1362, N974);
nand NAND2 (N2826, N2815, N1524);
nor NOR2 (N2827, N2822, N173);
nor NOR4 (N2828, N2798, N23, N2592, N2396);
nand NAND3 (N2829, N2826, N2269, N487);
xor XOR2 (N2830, N2816, N2256);
nand NAND3 (N2831, N2828, N2106, N514);
buf BUF1 (N2832, N2829);
nand NAND3 (N2833, N2827, N2315, N2396);
and AND4 (N2834, N2833, N245, N1310, N1486);
or OR2 (N2835, N2813, N1999);
or OR3 (N2836, N2810, N2171, N213);
xor XOR2 (N2837, N2825, N326);
nor NOR3 (N2838, N2836, N2813, N2425);
nand NAND2 (N2839, N2831, N1162);
not NOT1 (N2840, N2834);
not NOT1 (N2841, N2824);
and AND4 (N2842, N2830, N899, N551, N1928);
and AND3 (N2843, N2839, N1015, N1698);
xor XOR2 (N2844, N2814, N525);
nor NOR3 (N2845, N2835, N987, N46);
or OR2 (N2846, N2841, N2498);
not NOT1 (N2847, N2845);
not NOT1 (N2848, N2840);
nand NAND4 (N2849, N2837, N2335, N2075, N2031);
xor XOR2 (N2850, N2832, N2652);
nor NOR3 (N2851, N2849, N339, N2825);
xor XOR2 (N2852, N2847, N1276);
nand NAND2 (N2853, N2848, N1198);
not NOT1 (N2854, N2846);
and AND4 (N2855, N2851, N503, N923, N52);
nor NOR4 (N2856, N2844, N2348, N1673, N1076);
or OR3 (N2857, N2850, N663, N2804);
buf BUF1 (N2858, N2857);
and AND2 (N2859, N2853, N1705);
nand NAND2 (N2860, N2817, N2597);
or OR3 (N2861, N2852, N2092, N415);
buf BUF1 (N2862, N2860);
and AND2 (N2863, N2842, N959);
nand NAND3 (N2864, N2856, N905, N1472);
nor NOR3 (N2865, N2863, N2047, N2594);
xor XOR2 (N2866, N2854, N346);
nand NAND4 (N2867, N2865, N1657, N677, N1494);
or OR3 (N2868, N2862, N999, N2117);
xor XOR2 (N2869, N2858, N2190);
nor NOR2 (N2870, N2838, N761);
nand NAND4 (N2871, N2868, N540, N1533, N2420);
nor NOR4 (N2872, N2867, N1637, N1841, N2593);
xor XOR2 (N2873, N2864, N1489);
not NOT1 (N2874, N2872);
xor XOR2 (N2875, N2843, N2496);
buf BUF1 (N2876, N2870);
nand NAND3 (N2877, N2874, N2455, N59);
xor XOR2 (N2878, N2859, N1870);
not NOT1 (N2879, N2873);
nor NOR4 (N2880, N2877, N2376, N157, N1405);
and AND3 (N2881, N2878, N1640, N238);
xor XOR2 (N2882, N2875, N2779);
or OR2 (N2883, N2879, N879);
or OR2 (N2884, N2871, N2841);
and AND4 (N2885, N2866, N1952, N1586, N1210);
xor XOR2 (N2886, N2876, N1724);
nor NOR3 (N2887, N2880, N1843, N1209);
or OR4 (N2888, N2884, N350, N1570, N1178);
not NOT1 (N2889, N2887);
and AND4 (N2890, N2885, N748, N1249, N2101);
buf BUF1 (N2891, N2881);
or OR3 (N2892, N2890, N1785, N2238);
not NOT1 (N2893, N2891);
xor XOR2 (N2894, N2883, N384);
nor NOR3 (N2895, N2855, N1129, N332);
xor XOR2 (N2896, N2869, N255);
and AND2 (N2897, N2886, N1634);
xor XOR2 (N2898, N2889, N2333);
xor XOR2 (N2899, N2888, N1722);
and AND2 (N2900, N2894, N2327);
and AND2 (N2901, N2882, N1345);
and AND3 (N2902, N2897, N2225, N2455);
buf BUF1 (N2903, N2893);
and AND4 (N2904, N2902, N2290, N1330, N1997);
buf BUF1 (N2905, N2903);
not NOT1 (N2906, N2895);
xor XOR2 (N2907, N2892, N454);
nand NAND3 (N2908, N2905, N1664, N2283);
or OR2 (N2909, N2906, N962);
nand NAND2 (N2910, N2908, N2113);
xor XOR2 (N2911, N2901, N2192);
buf BUF1 (N2912, N2910);
not NOT1 (N2913, N2861);
nor NOR4 (N2914, N2912, N1045, N2404, N1075);
xor XOR2 (N2915, N2907, N152);
nor NOR2 (N2916, N2896, N256);
nand NAND2 (N2917, N2916, N1725);
xor XOR2 (N2918, N2904, N2482);
nand NAND4 (N2919, N2899, N1337, N663, N2314);
not NOT1 (N2920, N2919);
and AND2 (N2921, N2914, N1622);
not NOT1 (N2922, N2921);
or OR4 (N2923, N2900, N1114, N650, N260);
not NOT1 (N2924, N2918);
xor XOR2 (N2925, N2915, N2288);
or OR2 (N2926, N2925, N1672);
and AND4 (N2927, N2898, N2313, N1116, N1265);
or OR2 (N2928, N2926, N293);
nor NOR4 (N2929, N2913, N358, N2167, N1039);
not NOT1 (N2930, N2920);
xor XOR2 (N2931, N2928, N1459);
nand NAND4 (N2932, N2931, N821, N1015, N1627);
buf BUF1 (N2933, N2927);
buf BUF1 (N2934, N2922);
or OR3 (N2935, N2909, N2342, N1212);
nor NOR3 (N2936, N2932, N529, N2576);
nand NAND3 (N2937, N2929, N1919, N1881);
or OR2 (N2938, N2911, N1381);
or OR2 (N2939, N2923, N1372);
or OR2 (N2940, N2939, N167);
nor NOR3 (N2941, N2933, N2085, N2368);
nor NOR2 (N2942, N2936, N870);
nand NAND2 (N2943, N2917, N837);
or OR4 (N2944, N2934, N1749, N350, N567);
nand NAND4 (N2945, N2938, N1952, N1760, N2159);
nand NAND2 (N2946, N2944, N2494);
buf BUF1 (N2947, N2941);
and AND3 (N2948, N2947, N1249, N1880);
nor NOR4 (N2949, N2945, N2820, N2742, N452);
nor NOR4 (N2950, N2930, N764, N94, N571);
xor XOR2 (N2951, N2948, N1845);
buf BUF1 (N2952, N2940);
not NOT1 (N2953, N2949);
xor XOR2 (N2954, N2950, N1004);
buf BUF1 (N2955, N2946);
nand NAND4 (N2956, N2924, N765, N575, N1394);
xor XOR2 (N2957, N2935, N2137);
not NOT1 (N2958, N2942);
xor XOR2 (N2959, N2952, N894);
nand NAND2 (N2960, N2957, N1335);
not NOT1 (N2961, N2956);
nor NOR3 (N2962, N2961, N1380, N1267);
nor NOR2 (N2963, N2959, N726);
buf BUF1 (N2964, N2963);
or OR4 (N2965, N2958, N479, N2005, N231);
nor NOR4 (N2966, N2955, N2627, N2860, N1110);
or OR2 (N2967, N2965, N607);
nor NOR2 (N2968, N2937, N2083);
buf BUF1 (N2969, N2954);
buf BUF1 (N2970, N2966);
or OR3 (N2971, N2970, N1994, N2313);
and AND3 (N2972, N2971, N2476, N86);
and AND3 (N2973, N2960, N2180, N1144);
nor NOR4 (N2974, N2951, N432, N1557, N980);
xor XOR2 (N2975, N2968, N1567);
xor XOR2 (N2976, N2953, N502);
nand NAND2 (N2977, N2964, N198);
and AND2 (N2978, N2973, N1199);
or OR4 (N2979, N2978, N1243, N676, N1633);
buf BUF1 (N2980, N2967);
xor XOR2 (N2981, N2962, N2512);
buf BUF1 (N2982, N2976);
nand NAND2 (N2983, N2974, N497);
xor XOR2 (N2984, N2943, N1169);
xor XOR2 (N2985, N2969, N714);
or OR2 (N2986, N2984, N439);
buf BUF1 (N2987, N2977);
nor NOR2 (N2988, N2986, N2260);
nor NOR3 (N2989, N2982, N290, N587);
and AND2 (N2990, N2975, N1024);
buf BUF1 (N2991, N2987);
nand NAND2 (N2992, N2980, N2827);
nor NOR3 (N2993, N2979, N1707, N2985);
xor XOR2 (N2994, N1548, N2929);
xor XOR2 (N2995, N2990, N1092);
not NOT1 (N2996, N2991);
xor XOR2 (N2997, N2993, N2316);
buf BUF1 (N2998, N2992);
and AND4 (N2999, N2997, N1228, N1368, N453);
nor NOR4 (N3000, N2988, N1389, N314, N309);
buf BUF1 (N3001, N2999);
xor XOR2 (N3002, N2998, N2972);
xor XOR2 (N3003, N751, N1732);
nand NAND3 (N3004, N2981, N1967, N977);
xor XOR2 (N3005, N2994, N1713);
buf BUF1 (N3006, N2995);
xor XOR2 (N3007, N3000, N2123);
and AND2 (N3008, N3005, N935);
nand NAND4 (N3009, N2983, N9, N1618, N348);
or OR4 (N3010, N3007, N1507, N967, N1606);
buf BUF1 (N3011, N3001);
nand NAND2 (N3012, N3011, N1120);
and AND2 (N3013, N3008, N2075);
buf BUF1 (N3014, N3013);
buf BUF1 (N3015, N3006);
and AND4 (N3016, N3004, N1868, N1496, N632);
buf BUF1 (N3017, N3012);
or OR2 (N3018, N3015, N2520);
nor NOR2 (N3019, N3010, N1558);
and AND2 (N3020, N2996, N700);
or OR2 (N3021, N3018, N1509);
xor XOR2 (N3022, N3021, N1096);
or OR2 (N3023, N3009, N1962);
or OR4 (N3024, N3014, N2983, N2729, N1514);
buf BUF1 (N3025, N3022);
nand NAND3 (N3026, N3017, N2601, N841);
or OR3 (N3027, N2989, N2798, N829);
nand NAND4 (N3028, N3023, N165, N1018, N2314);
buf BUF1 (N3029, N3016);
buf BUF1 (N3030, N3025);
and AND4 (N3031, N3019, N702, N2741, N1843);
buf BUF1 (N3032, N3031);
xor XOR2 (N3033, N3002, N1135);
not NOT1 (N3034, N3030);
buf BUF1 (N3035, N3027);
and AND2 (N3036, N3029, N1936);
xor XOR2 (N3037, N3032, N624);
nor NOR2 (N3038, N3036, N686);
not NOT1 (N3039, N3033);
not NOT1 (N3040, N3003);
buf BUF1 (N3041, N3020);
nor NOR4 (N3042, N3038, N1749, N1559, N603);
nor NOR2 (N3043, N3028, N2193);
buf BUF1 (N3044, N3043);
nor NOR3 (N3045, N3026, N304, N1927);
nor NOR4 (N3046, N3034, N769, N2872, N2966);
nor NOR4 (N3047, N3041, N1677, N1272, N2862);
nand NAND4 (N3048, N3046, N727, N2357, N657);
nand NAND4 (N3049, N3042, N1955, N1394, N2691);
or OR2 (N3050, N3039, N60);
and AND2 (N3051, N3024, N263);
not NOT1 (N3052, N3050);
nor NOR3 (N3053, N3040, N1993, N233);
and AND3 (N3054, N3045, N1221, N2401);
xor XOR2 (N3055, N3044, N2987);
not NOT1 (N3056, N3055);
buf BUF1 (N3057, N3037);
or OR2 (N3058, N3035, N888);
not NOT1 (N3059, N3054);
nand NAND3 (N3060, N3053, N137, N1323);
nand NAND4 (N3061, N3057, N589, N1877, N2105);
not NOT1 (N3062, N3059);
or OR3 (N3063, N3048, N2679, N2655);
buf BUF1 (N3064, N3060);
not NOT1 (N3065, N3061);
nor NOR4 (N3066, N3058, N1181, N2122, N2129);
nand NAND2 (N3067, N3056, N815);
and AND4 (N3068, N3065, N1031, N715, N961);
xor XOR2 (N3069, N3063, N3016);
not NOT1 (N3070, N3052);
not NOT1 (N3071, N3064);
nor NOR3 (N3072, N3051, N3001, N1719);
and AND2 (N3073, N3066, N754);
and AND3 (N3074, N3068, N161, N2541);
buf BUF1 (N3075, N3074);
not NOT1 (N3076, N3072);
buf BUF1 (N3077, N3076);
or OR4 (N3078, N3070, N2026, N1446, N753);
nand NAND3 (N3079, N3077, N2700, N2571);
not NOT1 (N3080, N3067);
xor XOR2 (N3081, N3080, N1221);
not NOT1 (N3082, N3071);
and AND3 (N3083, N3082, N2344, N2742);
not NOT1 (N3084, N3047);
or OR3 (N3085, N3084, N1518, N711);
buf BUF1 (N3086, N3081);
and AND4 (N3087, N3086, N739, N2137, N1231);
nor NOR2 (N3088, N3083, N3070);
buf BUF1 (N3089, N3073);
not NOT1 (N3090, N3062);
nor NOR2 (N3091, N3090, N152);
buf BUF1 (N3092, N3089);
and AND2 (N3093, N3078, N906);
buf BUF1 (N3094, N3088);
nor NOR2 (N3095, N3094, N2709);
nor NOR2 (N3096, N3093, N2741);
or OR3 (N3097, N3075, N606, N123);
xor XOR2 (N3098, N3091, N2941);
nand NAND4 (N3099, N3092, N3072, N2929, N2033);
nor NOR4 (N3100, N3087, N1447, N2143, N1901);
and AND4 (N3101, N3096, N1119, N2577, N2937);
xor XOR2 (N3102, N3099, N2217);
buf BUF1 (N3103, N3097);
xor XOR2 (N3104, N3085, N1330);
xor XOR2 (N3105, N3104, N979);
xor XOR2 (N3106, N3102, N897);
xor XOR2 (N3107, N3069, N774);
xor XOR2 (N3108, N3095, N269);
or OR2 (N3109, N3100, N180);
nand NAND2 (N3110, N3107, N9);
xor XOR2 (N3111, N3106, N3034);
nor NOR4 (N3112, N3101, N935, N972, N979);
nor NOR3 (N3113, N3049, N875, N2699);
nand NAND3 (N3114, N3098, N360, N2753);
and AND2 (N3115, N3108, N620);
xor XOR2 (N3116, N3115, N57);
or OR2 (N3117, N3110, N948);
buf BUF1 (N3118, N3103);
not NOT1 (N3119, N3111);
and AND2 (N3120, N3079, N1983);
xor XOR2 (N3121, N3116, N438);
xor XOR2 (N3122, N3120, N637);
nand NAND2 (N3123, N3114, N3122);
nor NOR3 (N3124, N937, N2209, N507);
not NOT1 (N3125, N3119);
nor NOR3 (N3126, N3109, N1641, N1490);
and AND3 (N3127, N3124, N316, N239);
or OR3 (N3128, N3117, N250, N1369);
not NOT1 (N3129, N3112);
xor XOR2 (N3130, N3113, N2770);
or OR4 (N3131, N3128, N2966, N1417, N2930);
xor XOR2 (N3132, N3105, N2152);
or OR4 (N3133, N3130, N795, N1228, N834);
nor NOR2 (N3134, N3129, N2545);
xor XOR2 (N3135, N3131, N2405);
or OR2 (N3136, N3127, N2244);
nor NOR4 (N3137, N3134, N1984, N2146, N1690);
nand NAND2 (N3138, N3133, N1608);
not NOT1 (N3139, N3125);
nor NOR4 (N3140, N3123, N3111, N2414, N139);
nand NAND2 (N3141, N3121, N1473);
buf BUF1 (N3142, N3136);
buf BUF1 (N3143, N3139);
buf BUF1 (N3144, N3143);
not NOT1 (N3145, N3126);
and AND2 (N3146, N3141, N2416);
buf BUF1 (N3147, N3118);
and AND3 (N3148, N3145, N1288, N59);
not NOT1 (N3149, N3135);
xor XOR2 (N3150, N3142, N2787);
not NOT1 (N3151, N3137);
buf BUF1 (N3152, N3151);
or OR2 (N3153, N3152, N1006);
and AND4 (N3154, N3144, N2223, N586, N2354);
nand NAND4 (N3155, N3140, N1616, N202, N1081);
nand NAND2 (N3156, N3148, N562);
nand NAND2 (N3157, N3138, N2269);
xor XOR2 (N3158, N3153, N2253);
or OR3 (N3159, N3155, N2687, N1471);
nand NAND4 (N3160, N3132, N2113, N2516, N669);
buf BUF1 (N3161, N3150);
nor NOR4 (N3162, N3161, N403, N1497, N1676);
and AND4 (N3163, N3147, N1582, N1633, N1169);
not NOT1 (N3164, N3146);
nand NAND2 (N3165, N3157, N49);
not NOT1 (N3166, N3159);
xor XOR2 (N3167, N3163, N2459);
buf BUF1 (N3168, N3165);
or OR2 (N3169, N3162, N1321);
xor XOR2 (N3170, N3158, N2625);
and AND3 (N3171, N3156, N799, N3105);
nand NAND3 (N3172, N3168, N1174, N871);
xor XOR2 (N3173, N3167, N938);
buf BUF1 (N3174, N3172);
or OR2 (N3175, N3149, N3056);
buf BUF1 (N3176, N3164);
buf BUF1 (N3177, N3154);
not NOT1 (N3178, N3175);
nand NAND4 (N3179, N3171, N225, N915, N1439);
buf BUF1 (N3180, N3173);
nand NAND3 (N3181, N3174, N229, N1081);
or OR3 (N3182, N3169, N2502, N1198);
nor NOR4 (N3183, N3182, N2152, N2193, N1841);
nand NAND3 (N3184, N3181, N1366, N285);
xor XOR2 (N3185, N3180, N2696);
nor NOR3 (N3186, N3184, N2808, N2270);
xor XOR2 (N3187, N3166, N2171);
nand NAND3 (N3188, N3187, N2270, N2199);
xor XOR2 (N3189, N3177, N2531);
not NOT1 (N3190, N3179);
nand NAND3 (N3191, N3189, N1301, N1792);
buf BUF1 (N3192, N3170);
nor NOR3 (N3193, N3186, N1150, N1389);
and AND4 (N3194, N3185, N500, N2612, N1135);
nor NOR4 (N3195, N3188, N3043, N677, N2912);
nor NOR3 (N3196, N3178, N1795, N1549);
buf BUF1 (N3197, N3195);
and AND3 (N3198, N3193, N146, N100);
not NOT1 (N3199, N3183);
and AND3 (N3200, N3191, N2016, N2847);
buf BUF1 (N3201, N3190);
xor XOR2 (N3202, N3200, N1836);
or OR4 (N3203, N3196, N2275, N25, N274);
nand NAND3 (N3204, N3194, N1302, N2335);
buf BUF1 (N3205, N3199);
and AND4 (N3206, N3176, N2678, N688, N2735);
xor XOR2 (N3207, N3204, N919);
xor XOR2 (N3208, N3160, N3096);
xor XOR2 (N3209, N3206, N915);
nor NOR4 (N3210, N3197, N303, N2595, N2496);
nor NOR2 (N3211, N3202, N2833);
xor XOR2 (N3212, N3203, N2879);
or OR4 (N3213, N3192, N2034, N1520, N2307);
and AND3 (N3214, N3210, N2658, N1087);
nand NAND3 (N3215, N3205, N15, N484);
buf BUF1 (N3216, N3198);
xor XOR2 (N3217, N3208, N659);
not NOT1 (N3218, N3201);
or OR4 (N3219, N3211, N367, N2065, N1840);
nor NOR3 (N3220, N3219, N2135, N2121);
xor XOR2 (N3221, N3215, N1928);
or OR2 (N3222, N3209, N1413);
and AND4 (N3223, N3214, N2893, N2565, N1170);
and AND4 (N3224, N3220, N1288, N2597, N976);
nor NOR2 (N3225, N3207, N3218);
or OR2 (N3226, N2945, N1881);
nand NAND4 (N3227, N3226, N324, N2601, N1556);
or OR4 (N3228, N3225, N2210, N2743, N2448);
and AND3 (N3229, N3217, N1144, N913);
xor XOR2 (N3230, N3223, N1751);
buf BUF1 (N3231, N3212);
or OR4 (N3232, N3230, N113, N1801, N2351);
nor NOR3 (N3233, N3222, N1318, N1217);
or OR4 (N3234, N3231, N2850, N2597, N97);
not NOT1 (N3235, N3229);
nand NAND3 (N3236, N3233, N2845, N2798);
nand NAND3 (N3237, N3227, N2734, N843);
or OR3 (N3238, N3237, N1703, N556);
buf BUF1 (N3239, N3216);
or OR4 (N3240, N3221, N828, N1671, N603);
buf BUF1 (N3241, N3228);
or OR2 (N3242, N3234, N374);
or OR4 (N3243, N3242, N2862, N517, N1199);
and AND2 (N3244, N3239, N3116);
nand NAND2 (N3245, N3238, N1665);
buf BUF1 (N3246, N3241);
xor XOR2 (N3247, N3244, N722);
not NOT1 (N3248, N3246);
or OR3 (N3249, N3240, N2314, N1441);
nand NAND2 (N3250, N3224, N1900);
and AND4 (N3251, N3245, N230, N1666, N2621);
xor XOR2 (N3252, N3248, N3127);
or OR2 (N3253, N3232, N697);
nand NAND3 (N3254, N3236, N1407, N2334);
and AND2 (N3255, N3254, N1670);
buf BUF1 (N3256, N3235);
nand NAND4 (N3257, N3213, N496, N2014, N420);
nor NOR4 (N3258, N3247, N712, N1371, N1699);
and AND3 (N3259, N3258, N407, N1344);
and AND3 (N3260, N3256, N595, N2456);
and AND4 (N3261, N3251, N1333, N255, N251);
and AND4 (N3262, N3255, N1436, N2537, N1349);
or OR4 (N3263, N3261, N308, N3215, N2348);
and AND2 (N3264, N3250, N2758);
buf BUF1 (N3265, N3249);
buf BUF1 (N3266, N3243);
nor NOR3 (N3267, N3262, N668, N1256);
xor XOR2 (N3268, N3263, N1970);
or OR2 (N3269, N3253, N2053);
nor NOR3 (N3270, N3259, N1539, N1500);
or OR4 (N3271, N3266, N395, N1839, N701);
not NOT1 (N3272, N3260);
nand NAND3 (N3273, N3252, N193, N1582);
xor XOR2 (N3274, N3272, N1795);
xor XOR2 (N3275, N3271, N1446);
nor NOR3 (N3276, N3275, N199, N2888);
nor NOR3 (N3277, N3267, N2401, N1324);
or OR4 (N3278, N3257, N2233, N533, N368);
or OR2 (N3279, N3276, N2119);
buf BUF1 (N3280, N3273);
not NOT1 (N3281, N3264);
nor NOR2 (N3282, N3280, N1060);
buf BUF1 (N3283, N3269);
nand NAND4 (N3284, N3268, N2144, N1383, N506);
not NOT1 (N3285, N3279);
nor NOR2 (N3286, N3278, N2144);
not NOT1 (N3287, N3286);
and AND4 (N3288, N3281, N2478, N2170, N248);
not NOT1 (N3289, N3277);
nand NAND3 (N3290, N3285, N42, N2522);
xor XOR2 (N3291, N3289, N1721);
and AND2 (N3292, N3274, N3207);
nand NAND4 (N3293, N3288, N1783, N2926, N2679);
nor NOR3 (N3294, N3293, N1466, N25);
xor XOR2 (N3295, N3294, N2280);
nor NOR2 (N3296, N3292, N2928);
xor XOR2 (N3297, N3265, N1155);
nor NOR2 (N3298, N3296, N519);
buf BUF1 (N3299, N3270);
xor XOR2 (N3300, N3284, N1569);
buf BUF1 (N3301, N3282);
nor NOR4 (N3302, N3290, N2114, N2616, N1889);
xor XOR2 (N3303, N3295, N317);
nand NAND2 (N3304, N3299, N2135);
xor XOR2 (N3305, N3291, N1378);
nor NOR2 (N3306, N3297, N527);
buf BUF1 (N3307, N3300);
nor NOR2 (N3308, N3307, N2581);
not NOT1 (N3309, N3302);
not NOT1 (N3310, N3287);
xor XOR2 (N3311, N3305, N2065);
nand NAND4 (N3312, N3309, N1281, N3108, N1030);
and AND4 (N3313, N3301, N2254, N2734, N136);
xor XOR2 (N3314, N3298, N1902);
not NOT1 (N3315, N3303);
not NOT1 (N3316, N3315);
not NOT1 (N3317, N3311);
not NOT1 (N3318, N3308);
nand NAND2 (N3319, N3310, N3006);
xor XOR2 (N3320, N3313, N45);
nor NOR3 (N3321, N3318, N1674, N490);
not NOT1 (N3322, N3306);
xor XOR2 (N3323, N3314, N2737);
nor NOR2 (N3324, N3317, N756);
nand NAND2 (N3325, N3320, N3136);
nor NOR2 (N3326, N3325, N1007);
and AND3 (N3327, N3312, N1125, N688);
xor XOR2 (N3328, N3322, N2088);
nor NOR3 (N3329, N3304, N669, N2305);
or OR2 (N3330, N3326, N2115);
nand NAND2 (N3331, N3329, N2697);
buf BUF1 (N3332, N3328);
xor XOR2 (N3333, N3323, N1926);
buf BUF1 (N3334, N3330);
nor NOR3 (N3335, N3333, N882, N502);
and AND4 (N3336, N3334, N1999, N1970, N1959);
and AND4 (N3337, N3321, N1899, N408, N1556);
nor NOR4 (N3338, N3332, N1030, N20, N2547);
buf BUF1 (N3339, N3336);
and AND4 (N3340, N3331, N2849, N307, N799);
not NOT1 (N3341, N3316);
nor NOR3 (N3342, N3341, N2459, N72);
xor XOR2 (N3343, N3283, N1090);
or OR4 (N3344, N3327, N1650, N2148, N386);
not NOT1 (N3345, N3343);
xor XOR2 (N3346, N3340, N2310);
and AND2 (N3347, N3335, N2275);
buf BUF1 (N3348, N3345);
nor NOR2 (N3349, N3338, N137);
nor NOR3 (N3350, N3342, N1555, N1471);
nor NOR3 (N3351, N3344, N2396, N462);
buf BUF1 (N3352, N3319);
not NOT1 (N3353, N3337);
not NOT1 (N3354, N3350);
xor XOR2 (N3355, N3324, N2944);
xor XOR2 (N3356, N3348, N7);
not NOT1 (N3357, N3339);
nand NAND2 (N3358, N3352, N1577);
xor XOR2 (N3359, N3358, N2953);
and AND2 (N3360, N3347, N437);
and AND4 (N3361, N3346, N785, N2228, N1182);
nand NAND3 (N3362, N3361, N1025, N2707);
buf BUF1 (N3363, N3351);
xor XOR2 (N3364, N3354, N3361);
not NOT1 (N3365, N3363);
nand NAND3 (N3366, N3356, N2579, N1001);
buf BUF1 (N3367, N3362);
not NOT1 (N3368, N3364);
nor NOR2 (N3369, N3368, N2353);
or OR3 (N3370, N3357, N2261, N2839);
buf BUF1 (N3371, N3366);
not NOT1 (N3372, N3349);
or OR4 (N3373, N3371, N3027, N3188, N1288);
not NOT1 (N3374, N3369);
not NOT1 (N3375, N3374);
nor NOR2 (N3376, N3367, N2628);
not NOT1 (N3377, N3372);
nand NAND3 (N3378, N3359, N2033, N2155);
nor NOR4 (N3379, N3378, N1065, N1886, N2348);
nand NAND3 (N3380, N3360, N495, N1340);
buf BUF1 (N3381, N3375);
and AND3 (N3382, N3376, N1153, N3021);
nor NOR2 (N3383, N3373, N1837);
xor XOR2 (N3384, N3379, N792);
nand NAND3 (N3385, N3355, N3172, N1989);
and AND2 (N3386, N3384, N1466);
or OR3 (N3387, N3370, N1972, N2747);
xor XOR2 (N3388, N3382, N322);
buf BUF1 (N3389, N3388);
buf BUF1 (N3390, N3365);
nor NOR4 (N3391, N3385, N1840, N2447, N3189);
buf BUF1 (N3392, N3380);
or OR3 (N3393, N3389, N1274, N1140);
buf BUF1 (N3394, N3392);
and AND2 (N3395, N3377, N1550);
and AND2 (N3396, N3353, N3183);
or OR2 (N3397, N3396, N1703);
and AND2 (N3398, N3395, N2301);
and AND4 (N3399, N3381, N3121, N2727, N2440);
nand NAND4 (N3400, N3399, N685, N3247, N2294);
not NOT1 (N3401, N3397);
nand NAND4 (N3402, N3391, N191, N1326, N858);
nor NOR2 (N3403, N3390, N1872);
nor NOR4 (N3404, N3403, N2683, N1556, N1370);
or OR3 (N3405, N3383, N745, N123);
nor NOR4 (N3406, N3394, N2237, N366, N2855);
xor XOR2 (N3407, N3401, N3086);
or OR3 (N3408, N3386, N3266, N1277);
nor NOR3 (N3409, N3387, N3375, N2534);
nor NOR4 (N3410, N3406, N1006, N2621, N1117);
not NOT1 (N3411, N3405);
nor NOR4 (N3412, N3409, N36, N3252, N1271);
nand NAND3 (N3413, N3398, N2231, N491);
buf BUF1 (N3414, N3411);
nor NOR3 (N3415, N3393, N1752, N1247);
xor XOR2 (N3416, N3412, N512);
not NOT1 (N3417, N3416);
nor NOR3 (N3418, N3417, N2070, N2706);
or OR4 (N3419, N3402, N3028, N2009, N2466);
buf BUF1 (N3420, N3404);
nand NAND4 (N3421, N3414, N2381, N2481, N1416);
not NOT1 (N3422, N3407);
nand NAND2 (N3423, N3419, N695);
nand NAND2 (N3424, N3421, N1749);
buf BUF1 (N3425, N3408);
nor NOR2 (N3426, N3410, N2948);
or OR3 (N3427, N3418, N1238, N1535);
not NOT1 (N3428, N3424);
not NOT1 (N3429, N3422);
buf BUF1 (N3430, N3427);
xor XOR2 (N3431, N3429, N1488);
not NOT1 (N3432, N3400);
not NOT1 (N3433, N3413);
or OR4 (N3434, N3430, N1671, N1532, N2314);
nand NAND2 (N3435, N3426, N792);
xor XOR2 (N3436, N3415, N1712);
buf BUF1 (N3437, N3431);
nand NAND2 (N3438, N3433, N753);
not NOT1 (N3439, N3438);
nor NOR2 (N3440, N3437, N3354);
not NOT1 (N3441, N3440);
buf BUF1 (N3442, N3434);
xor XOR2 (N3443, N3441, N2375);
and AND4 (N3444, N3443, N929, N706, N164);
nor NOR3 (N3445, N3444, N1202, N20);
buf BUF1 (N3446, N3428);
not NOT1 (N3447, N3432);
buf BUF1 (N3448, N3439);
and AND2 (N3449, N3420, N394);
not NOT1 (N3450, N3435);
buf BUF1 (N3451, N3423);
nand NAND4 (N3452, N3447, N3033, N1433, N2989);
buf BUF1 (N3453, N3452);
buf BUF1 (N3454, N3450);
or OR2 (N3455, N3446, N2230);
nor NOR2 (N3456, N3454, N1414);
or OR4 (N3457, N3456, N504, N1760, N317);
nand NAND4 (N3458, N3449, N2397, N2098, N299);
and AND2 (N3459, N3458, N871);
or OR4 (N3460, N3445, N3194, N519, N1318);
xor XOR2 (N3461, N3455, N157);
and AND4 (N3462, N3453, N2156, N1530, N2432);
and AND2 (N3463, N3442, N1192);
nand NAND3 (N3464, N3436, N161, N28);
nand NAND4 (N3465, N3457, N3224, N2410, N3223);
xor XOR2 (N3466, N3464, N1158);
or OR4 (N3467, N3466, N2990, N542, N2536);
nor NOR3 (N3468, N3467, N3117, N292);
not NOT1 (N3469, N3451);
nor NOR2 (N3470, N3465, N2042);
and AND4 (N3471, N3448, N2422, N2010, N3203);
and AND2 (N3472, N3469, N2362);
or OR2 (N3473, N3470, N1701);
and AND4 (N3474, N3425, N1468, N2472, N2567);
nand NAND4 (N3475, N3461, N600, N1611, N846);
nand NAND3 (N3476, N3462, N3083, N2358);
buf BUF1 (N3477, N3459);
nand NAND2 (N3478, N3473, N1399);
xor XOR2 (N3479, N3477, N1534);
not NOT1 (N3480, N3478);
or OR2 (N3481, N3480, N1163);
nor NOR4 (N3482, N3463, N2942, N1018, N717);
nand NAND4 (N3483, N3482, N684, N740, N1978);
xor XOR2 (N3484, N3476, N1186);
not NOT1 (N3485, N3472);
nor NOR3 (N3486, N3479, N3169, N171);
or OR2 (N3487, N3468, N3198);
and AND3 (N3488, N3471, N2626, N2480);
or OR3 (N3489, N3460, N1849, N2068);
and AND3 (N3490, N3486, N2665, N468);
nand NAND2 (N3491, N3474, N496);
or OR3 (N3492, N3481, N841, N638);
buf BUF1 (N3493, N3483);
xor XOR2 (N3494, N3490, N128);
buf BUF1 (N3495, N3494);
nand NAND3 (N3496, N3485, N1172, N1744);
buf BUF1 (N3497, N3487);
xor XOR2 (N3498, N3497, N2049);
nor NOR4 (N3499, N3484, N83, N1346, N965);
xor XOR2 (N3500, N3491, N1051);
nor NOR2 (N3501, N3489, N236);
nor NOR2 (N3502, N3475, N3320);
and AND3 (N3503, N3499, N1597, N728);
nor NOR3 (N3504, N3498, N3245, N2777);
buf BUF1 (N3505, N3500);
or OR2 (N3506, N3502, N2887);
nand NAND4 (N3507, N3488, N2655, N1855, N935);
xor XOR2 (N3508, N3505, N2659);
and AND4 (N3509, N3496, N560, N2020, N47);
not NOT1 (N3510, N3507);
nand NAND2 (N3511, N3506, N3268);
endmodule