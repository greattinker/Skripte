// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11;

output N2497,N2509,N2471,N2510,N2508,N2507,N2500,N2502,N2505,N2511;

and AND4 (N12, N2, N2, N2, N7);
and AND2 (N13, N10, N7);
nand NAND2 (N14, N6, N4);
nor NOR3 (N15, N1, N6, N6);
not NOT1 (N16, N2);
or OR4 (N17, N12, N11, N8, N15);
and AND2 (N18, N8, N16);
xor XOR2 (N19, N16, N10);
or OR2 (N20, N4, N17);
or OR3 (N21, N11, N16, N20);
and AND3 (N22, N7, N17, N1);
or OR2 (N23, N8, N11);
not NOT1 (N24, N3);
nor NOR4 (N25, N5, N14, N22, N19);
and AND2 (N26, N9, N7);
buf BUF1 (N27, N20);
not NOT1 (N28, N9);
or OR3 (N29, N15, N19, N19);
or OR2 (N30, N13, N1);
nor NOR2 (N31, N28, N29);
xor XOR2 (N32, N13, N21);
nand NAND2 (N33, N26, N16);
buf BUF1 (N34, N20);
or OR2 (N35, N25, N30);
not NOT1 (N36, N20);
nor NOR2 (N37, N35, N24);
nor NOR2 (N38, N9, N11);
nand NAND4 (N39, N32, N31, N10, N8);
xor XOR2 (N40, N37, N11);
and AND2 (N41, N28, N6);
or OR2 (N42, N27, N6);
xor XOR2 (N43, N33, N16);
xor XOR2 (N44, N34, N14);
nor NOR4 (N45, N40, N37, N34, N37);
or OR4 (N46, N43, N14, N29, N25);
buf BUF1 (N47, N42);
xor XOR2 (N48, N44, N43);
buf BUF1 (N49, N41);
nor NOR2 (N50, N18, N28);
buf BUF1 (N51, N39);
nand NAND2 (N52, N23, N48);
buf BUF1 (N53, N18);
and AND3 (N54, N49, N35, N22);
not NOT1 (N55, N45);
or OR2 (N56, N47, N54);
buf BUF1 (N57, N1);
and AND4 (N58, N46, N18, N10, N6);
xor XOR2 (N59, N52, N18);
not NOT1 (N60, N59);
nor NOR2 (N61, N58, N7);
xor XOR2 (N62, N53, N55);
nor NOR2 (N63, N48, N35);
and AND4 (N64, N50, N8, N11, N7);
and AND3 (N65, N61, N30, N43);
xor XOR2 (N66, N63, N44);
or OR2 (N67, N60, N50);
not NOT1 (N68, N38);
buf BUF1 (N69, N66);
not NOT1 (N70, N36);
not NOT1 (N71, N62);
xor XOR2 (N72, N56, N37);
not NOT1 (N73, N69);
and AND2 (N74, N71, N54);
buf BUF1 (N75, N70);
xor XOR2 (N76, N64, N14);
nor NOR2 (N77, N73, N4);
xor XOR2 (N78, N65, N16);
buf BUF1 (N79, N75);
nand NAND2 (N80, N74, N26);
nand NAND4 (N81, N67, N77, N22, N60);
xor XOR2 (N82, N5, N16);
and AND3 (N83, N79, N54, N43);
or OR2 (N84, N57, N44);
nor NOR2 (N85, N51, N52);
and AND3 (N86, N83, N16, N81);
not NOT1 (N87, N47);
and AND3 (N88, N68, N21, N44);
not NOT1 (N89, N72);
and AND2 (N90, N84, N32);
xor XOR2 (N91, N76, N7);
or OR4 (N92, N88, N65, N4, N28);
nor NOR3 (N93, N91, N10, N69);
or OR2 (N94, N93, N9);
or OR4 (N95, N80, N23, N33, N45);
or OR3 (N96, N94, N30, N52);
nand NAND4 (N97, N85, N88, N24, N87);
nand NAND2 (N98, N35, N55);
nor NOR4 (N99, N95, N47, N63, N34);
or OR4 (N100, N78, N28, N92, N52);
not NOT1 (N101, N90);
nand NAND2 (N102, N63, N1);
not NOT1 (N103, N89);
and AND3 (N104, N103, N9, N55);
or OR2 (N105, N86, N11);
nand NAND3 (N106, N105, N49, N50);
nand NAND2 (N107, N102, N44);
or OR2 (N108, N99, N58);
or OR4 (N109, N101, N28, N78, N24);
nand NAND3 (N110, N106, N8, N5);
nand NAND2 (N111, N97, N37);
or OR4 (N112, N107, N4, N84, N15);
and AND3 (N113, N96, N27, N75);
not NOT1 (N114, N110);
nand NAND4 (N115, N113, N91, N54, N27);
xor XOR2 (N116, N98, N31);
nand NAND3 (N117, N111, N45, N14);
nor NOR4 (N118, N112, N58, N75, N87);
not NOT1 (N119, N114);
nand NAND4 (N120, N116, N104, N104, N26);
xor XOR2 (N121, N101, N34);
nor NOR4 (N122, N100, N19, N56, N118);
or OR3 (N123, N23, N55, N27);
xor XOR2 (N124, N115, N17);
and AND4 (N125, N119, N64, N18, N23);
not NOT1 (N126, N125);
or OR4 (N127, N108, N78, N122, N65);
not NOT1 (N128, N81);
buf BUF1 (N129, N120);
or OR2 (N130, N129, N6);
not NOT1 (N131, N117);
and AND4 (N132, N123, N44, N26, N43);
nand NAND4 (N133, N127, N113, N107, N84);
not NOT1 (N134, N132);
xor XOR2 (N135, N131, N102);
nand NAND4 (N136, N126, N125, N104, N118);
buf BUF1 (N137, N133);
nand NAND2 (N138, N124, N65);
and AND3 (N139, N82, N119, N34);
nor NOR3 (N140, N109, N30, N29);
xor XOR2 (N141, N135, N105);
or OR4 (N142, N137, N88, N25, N39);
xor XOR2 (N143, N141, N98);
or OR3 (N144, N130, N94, N135);
or OR2 (N145, N143, N3);
or OR2 (N146, N145, N133);
or OR4 (N147, N128, N109, N32, N90);
not NOT1 (N148, N136);
nor NOR2 (N149, N147, N10);
or OR4 (N150, N149, N62, N106, N60);
not NOT1 (N151, N146);
xor XOR2 (N152, N134, N17);
or OR3 (N153, N121, N14, N79);
or OR3 (N154, N153, N104, N117);
or OR3 (N155, N151, N70, N129);
buf BUF1 (N156, N138);
buf BUF1 (N157, N154);
buf BUF1 (N158, N150);
xor XOR2 (N159, N139, N81);
and AND2 (N160, N158, N29);
nand NAND2 (N161, N140, N131);
or OR2 (N162, N155, N136);
not NOT1 (N163, N161);
nand NAND3 (N164, N163, N127, N84);
xor XOR2 (N165, N142, N124);
buf BUF1 (N166, N162);
buf BUF1 (N167, N160);
and AND3 (N168, N165, N21, N71);
buf BUF1 (N169, N152);
or OR2 (N170, N148, N158);
not NOT1 (N171, N170);
not NOT1 (N172, N166);
buf BUF1 (N173, N168);
xor XOR2 (N174, N157, N34);
and AND4 (N175, N172, N173, N13, N108);
xor XOR2 (N176, N4, N103);
xor XOR2 (N177, N169, N25);
nand NAND2 (N178, N144, N167);
buf BUF1 (N179, N91);
or OR2 (N180, N171, N177);
nand NAND4 (N181, N103, N47, N88, N78);
nand NAND4 (N182, N176, N144, N26, N90);
nor NOR2 (N183, N175, N117);
nor NOR4 (N184, N181, N166, N39, N96);
xor XOR2 (N185, N174, N75);
or OR4 (N186, N164, N45, N54, N163);
not NOT1 (N187, N156);
nor NOR3 (N188, N182, N82, N178);
not NOT1 (N189, N65);
xor XOR2 (N190, N179, N71);
not NOT1 (N191, N159);
not NOT1 (N192, N186);
xor XOR2 (N193, N190, N25);
not NOT1 (N194, N187);
and AND2 (N195, N180, N144);
not NOT1 (N196, N184);
nand NAND2 (N197, N196, N146);
buf BUF1 (N198, N191);
or OR4 (N199, N195, N49, N155, N185);
not NOT1 (N200, N198);
and AND3 (N201, N174, N179, N149);
nand NAND2 (N202, N200, N91);
or OR2 (N203, N183, N122);
or OR2 (N204, N192, N46);
and AND3 (N205, N204, N32, N70);
and AND2 (N206, N202, N32);
or OR3 (N207, N197, N193, N117);
xor XOR2 (N208, N185, N73);
buf BUF1 (N209, N207);
nand NAND3 (N210, N203, N58, N33);
xor XOR2 (N211, N194, N23);
nand NAND4 (N212, N206, N196, N92, N51);
nor NOR3 (N213, N201, N147, N16);
nor NOR4 (N214, N211, N98, N86, N110);
or OR3 (N215, N214, N212, N177);
not NOT1 (N216, N114);
nor NOR4 (N217, N205, N166, N4, N69);
buf BUF1 (N218, N199);
or OR2 (N219, N210, N55);
or OR4 (N220, N216, N210, N73, N172);
not NOT1 (N221, N189);
not NOT1 (N222, N217);
xor XOR2 (N223, N188, N124);
not NOT1 (N224, N222);
and AND2 (N225, N208, N119);
buf BUF1 (N226, N220);
nor NOR3 (N227, N223, N16, N19);
and AND2 (N228, N219, N218);
or OR2 (N229, N87, N138);
xor XOR2 (N230, N228, N70);
nor NOR2 (N231, N226, N209);
not NOT1 (N232, N224);
nor NOR2 (N233, N40, N144);
nand NAND2 (N234, N230, N20);
xor XOR2 (N235, N231, N136);
nand NAND4 (N236, N225, N52, N172, N116);
buf BUF1 (N237, N233);
or OR4 (N238, N229, N116, N75, N34);
xor XOR2 (N239, N235, N37);
xor XOR2 (N240, N238, N66);
xor XOR2 (N241, N237, N183);
xor XOR2 (N242, N239, N148);
buf BUF1 (N243, N236);
xor XOR2 (N244, N241, N161);
and AND4 (N245, N215, N142, N39, N174);
nor NOR3 (N246, N227, N13, N226);
not NOT1 (N247, N213);
buf BUF1 (N248, N221);
xor XOR2 (N249, N245, N24);
not NOT1 (N250, N243);
and AND4 (N251, N247, N73, N240, N90);
buf BUF1 (N252, N124);
nand NAND2 (N253, N250, N78);
not NOT1 (N254, N251);
nand NAND3 (N255, N248, N135, N96);
nor NOR3 (N256, N252, N35, N243);
buf BUF1 (N257, N249);
nand NAND2 (N258, N257, N232);
and AND4 (N259, N28, N11, N218, N220);
xor XOR2 (N260, N242, N203);
or OR3 (N261, N244, N59, N209);
xor XOR2 (N262, N259, N128);
and AND3 (N263, N255, N86, N204);
or OR3 (N264, N262, N133, N233);
nand NAND2 (N265, N258, N40);
nand NAND4 (N266, N265, N92, N193, N17);
not NOT1 (N267, N254);
xor XOR2 (N268, N263, N109);
and AND3 (N269, N246, N84, N41);
not NOT1 (N270, N268);
or OR4 (N271, N266, N153, N206, N214);
nor NOR2 (N272, N269, N12);
xor XOR2 (N273, N261, N3);
or OR4 (N274, N256, N30, N83, N225);
nor NOR2 (N275, N272, N66);
nor NOR3 (N276, N275, N24, N255);
nand NAND3 (N277, N271, N26, N57);
buf BUF1 (N278, N267);
xor XOR2 (N279, N234, N197);
or OR4 (N280, N273, N53, N20, N66);
not NOT1 (N281, N270);
xor XOR2 (N282, N279, N49);
nand NAND3 (N283, N260, N86, N191);
nor NOR4 (N284, N264, N49, N67, N69);
or OR2 (N285, N277, N92);
nand NAND3 (N286, N274, N79, N14);
nand NAND3 (N287, N283, N131, N145);
nand NAND4 (N288, N276, N164, N247, N41);
xor XOR2 (N289, N278, N198);
nor NOR3 (N290, N281, N141, N45);
not NOT1 (N291, N287);
nand NAND3 (N292, N253, N227, N272);
and AND3 (N293, N289, N114, N40);
nor NOR3 (N294, N290, N82, N134);
not NOT1 (N295, N282);
nor NOR4 (N296, N294, N182, N239, N61);
nand NAND2 (N297, N280, N66);
and AND3 (N298, N285, N276, N154);
nor NOR3 (N299, N298, N48, N284);
not NOT1 (N300, N98);
nand NAND4 (N301, N292, N81, N56, N129);
nand NAND2 (N302, N293, N158);
nand NAND3 (N303, N286, N42, N264);
nand NAND4 (N304, N297, N94, N8, N58);
not NOT1 (N305, N299);
and AND4 (N306, N303, N10, N82, N280);
not NOT1 (N307, N300);
not NOT1 (N308, N296);
buf BUF1 (N309, N288);
nand NAND4 (N310, N295, N125, N121, N16);
or OR4 (N311, N304, N257, N26, N79);
or OR4 (N312, N302, N66, N270, N152);
xor XOR2 (N313, N312, N12);
buf BUF1 (N314, N301);
or OR4 (N315, N308, N76, N115, N119);
nand NAND3 (N316, N306, N232, N178);
or OR4 (N317, N310, N262, N309, N13);
xor XOR2 (N318, N145, N78);
xor XOR2 (N319, N291, N221);
buf BUF1 (N320, N319);
or OR2 (N321, N314, N139);
and AND3 (N322, N316, N65, N74);
and AND4 (N323, N321, N96, N18, N282);
xor XOR2 (N324, N318, N256);
not NOT1 (N325, N305);
buf BUF1 (N326, N315);
xor XOR2 (N327, N323, N25);
nand NAND4 (N328, N307, N293, N243, N60);
or OR3 (N329, N328, N103, N103);
nand NAND3 (N330, N322, N4, N260);
and AND4 (N331, N325, N142, N44, N89);
nand NAND3 (N332, N326, N287, N327);
buf BUF1 (N333, N150);
xor XOR2 (N334, N332, N301);
or OR3 (N335, N333, N326, N242);
not NOT1 (N336, N331);
xor XOR2 (N337, N334, N229);
not NOT1 (N338, N337);
buf BUF1 (N339, N324);
xor XOR2 (N340, N336, N112);
xor XOR2 (N341, N330, N222);
nand NAND4 (N342, N339, N306, N316, N163);
buf BUF1 (N343, N341);
buf BUF1 (N344, N340);
xor XOR2 (N345, N317, N203);
buf BUF1 (N346, N343);
xor XOR2 (N347, N346, N154);
nand NAND4 (N348, N335, N322, N57, N315);
and AND2 (N349, N342, N289);
or OR2 (N350, N311, N170);
and AND2 (N351, N347, N33);
buf BUF1 (N352, N351);
nand NAND2 (N353, N344, N300);
nand NAND4 (N354, N352, N315, N234, N71);
not NOT1 (N355, N338);
not NOT1 (N356, N353);
buf BUF1 (N357, N349);
nor NOR3 (N358, N350, N245, N178);
nor NOR3 (N359, N357, N82, N204);
nor NOR3 (N360, N359, N323, N346);
nand NAND3 (N361, N345, N279, N100);
and AND3 (N362, N358, N101, N56);
buf BUF1 (N363, N361);
or OR4 (N364, N363, N242, N134, N1);
not NOT1 (N365, N364);
nor NOR4 (N366, N348, N222, N19, N252);
or OR2 (N367, N356, N340);
xor XOR2 (N368, N367, N109);
xor XOR2 (N369, N354, N91);
nor NOR2 (N370, N355, N127);
xor XOR2 (N371, N365, N227);
or OR2 (N372, N320, N63);
and AND4 (N373, N368, N217, N267, N348);
and AND2 (N374, N371, N297);
buf BUF1 (N375, N362);
buf BUF1 (N376, N360);
nor NOR2 (N377, N366, N319);
and AND3 (N378, N370, N301, N212);
not NOT1 (N379, N378);
not NOT1 (N380, N376);
and AND3 (N381, N380, N203, N2);
nor NOR2 (N382, N372, N59);
nor NOR2 (N383, N329, N129);
nand NAND2 (N384, N381, N180);
buf BUF1 (N385, N375);
nor NOR3 (N386, N379, N305, N73);
or OR3 (N387, N313, N334, N264);
buf BUF1 (N388, N373);
nand NAND4 (N389, N382, N33, N123, N111);
xor XOR2 (N390, N384, N275);
nand NAND3 (N391, N385, N236, N342);
xor XOR2 (N392, N387, N192);
xor XOR2 (N393, N391, N7);
nand NAND4 (N394, N392, N93, N98, N371);
not NOT1 (N395, N394);
nand NAND2 (N396, N395, N260);
buf BUF1 (N397, N386);
nand NAND4 (N398, N383, N173, N324, N164);
not NOT1 (N399, N393);
not NOT1 (N400, N389);
not NOT1 (N401, N397);
not NOT1 (N402, N374);
and AND4 (N403, N399, N226, N88, N112);
not NOT1 (N404, N403);
nand NAND4 (N405, N396, N131, N264, N186);
xor XOR2 (N406, N388, N265);
buf BUF1 (N407, N398);
not NOT1 (N408, N404);
nand NAND4 (N409, N390, N90, N406, N152);
and AND4 (N410, N357, N199, N4, N66);
buf BUF1 (N411, N402);
nand NAND2 (N412, N411, N217);
nor NOR3 (N413, N409, N77, N233);
not NOT1 (N414, N413);
not NOT1 (N415, N414);
nor NOR2 (N416, N412, N103);
nor NOR4 (N417, N377, N296, N28, N214);
nor NOR2 (N418, N415, N358);
nor NOR3 (N419, N408, N56, N19);
nor NOR3 (N420, N401, N403, N316);
not NOT1 (N421, N420);
buf BUF1 (N422, N417);
not NOT1 (N423, N410);
not NOT1 (N424, N416);
nand NAND3 (N425, N369, N139, N138);
buf BUF1 (N426, N419);
nand NAND4 (N427, N424, N257, N360, N411);
and AND2 (N428, N423, N176);
or OR4 (N429, N421, N372, N137, N329);
nand NAND4 (N430, N418, N68, N282, N79);
nor NOR4 (N431, N427, N103, N293, N233);
nand NAND3 (N432, N430, N123, N138);
xor XOR2 (N433, N429, N220);
not NOT1 (N434, N422);
xor XOR2 (N435, N407, N77);
xor XOR2 (N436, N428, N196);
nand NAND4 (N437, N405, N238, N406, N104);
and AND2 (N438, N436, N338);
and AND4 (N439, N431, N278, N91, N351);
nor NOR4 (N440, N400, N96, N363, N403);
nand NAND3 (N441, N435, N109, N8);
not NOT1 (N442, N425);
or OR2 (N443, N440, N195);
not NOT1 (N444, N433);
not NOT1 (N445, N443);
xor XOR2 (N446, N438, N119);
nand NAND4 (N447, N444, N1, N219, N28);
buf BUF1 (N448, N446);
nor NOR3 (N449, N445, N357, N59);
buf BUF1 (N450, N447);
nor NOR2 (N451, N450, N152);
nor NOR2 (N452, N437, N447);
buf BUF1 (N453, N432);
nand NAND2 (N454, N451, N451);
buf BUF1 (N455, N448);
nor NOR4 (N456, N454, N35, N36, N103);
xor XOR2 (N457, N426, N108);
xor XOR2 (N458, N455, N255);
nand NAND4 (N459, N452, N206, N455, N393);
or OR4 (N460, N442, N104, N9, N223);
nand NAND3 (N461, N439, N71, N455);
and AND3 (N462, N434, N215, N382);
and AND3 (N463, N449, N273, N101);
buf BUF1 (N464, N459);
nor NOR3 (N465, N462, N73, N339);
nor NOR2 (N466, N465, N161);
and AND4 (N467, N460, N75, N424, N193);
nor NOR4 (N468, N453, N90, N404, N144);
or OR3 (N469, N468, N33, N172);
buf BUF1 (N470, N458);
not NOT1 (N471, N464);
and AND2 (N472, N463, N83);
xor XOR2 (N473, N461, N240);
xor XOR2 (N474, N441, N184);
and AND3 (N475, N467, N86, N394);
nor NOR3 (N476, N457, N212, N441);
nand NAND4 (N477, N473, N202, N83, N179);
or OR3 (N478, N466, N289, N71);
or OR2 (N479, N472, N345);
nand NAND4 (N480, N471, N386, N76, N173);
xor XOR2 (N481, N469, N136);
nand NAND3 (N482, N456, N296, N248);
or OR2 (N483, N481, N238);
nor NOR4 (N484, N483, N6, N206, N469);
not NOT1 (N485, N477);
not NOT1 (N486, N474);
not NOT1 (N487, N486);
buf BUF1 (N488, N475);
xor XOR2 (N489, N487, N435);
or OR2 (N490, N489, N92);
buf BUF1 (N491, N490);
not NOT1 (N492, N488);
or OR2 (N493, N470, N445);
not NOT1 (N494, N491);
and AND4 (N495, N484, N234, N485, N152);
nand NAND4 (N496, N489, N62, N383, N147);
xor XOR2 (N497, N479, N382);
nor NOR2 (N498, N494, N337);
or OR4 (N499, N480, N153, N317, N426);
buf BUF1 (N500, N497);
buf BUF1 (N501, N499);
xor XOR2 (N502, N478, N163);
nor NOR4 (N503, N502, N104, N98, N37);
xor XOR2 (N504, N476, N501);
xor XOR2 (N505, N345, N345);
buf BUF1 (N506, N498);
not NOT1 (N507, N495);
xor XOR2 (N508, N496, N367);
xor XOR2 (N509, N504, N289);
or OR4 (N510, N493, N265, N24, N95);
buf BUF1 (N511, N503);
not NOT1 (N512, N510);
or OR3 (N513, N505, N261, N344);
and AND2 (N514, N509, N182);
nor NOR4 (N515, N506, N214, N491, N326);
or OR4 (N516, N492, N399, N235, N9);
xor XOR2 (N517, N511, N495);
xor XOR2 (N518, N508, N240);
nand NAND3 (N519, N514, N336, N128);
xor XOR2 (N520, N515, N143);
xor XOR2 (N521, N518, N290);
not NOT1 (N522, N513);
not NOT1 (N523, N507);
buf BUF1 (N524, N517);
and AND4 (N525, N522, N2, N331, N62);
not NOT1 (N526, N523);
nand NAND2 (N527, N482, N50);
xor XOR2 (N528, N521, N20);
nor NOR3 (N529, N525, N440, N337);
nor NOR3 (N530, N500, N220, N391);
or OR2 (N531, N529, N460);
nor NOR2 (N532, N512, N426);
nor NOR3 (N533, N532, N433, N252);
not NOT1 (N534, N516);
nor NOR4 (N535, N533, N283, N356, N437);
not NOT1 (N536, N535);
not NOT1 (N537, N520);
xor XOR2 (N538, N537, N358);
nor NOR2 (N539, N519, N374);
buf BUF1 (N540, N539);
nand NAND2 (N541, N527, N321);
and AND3 (N542, N531, N244, N392);
xor XOR2 (N543, N526, N109);
not NOT1 (N544, N540);
nand NAND3 (N545, N541, N54, N505);
or OR4 (N546, N530, N354, N108, N65);
xor XOR2 (N547, N524, N106);
xor XOR2 (N548, N528, N445);
nand NAND3 (N549, N545, N349, N404);
and AND4 (N550, N538, N179, N455, N334);
or OR3 (N551, N543, N319, N337);
nand NAND2 (N552, N546, N247);
nor NOR3 (N553, N536, N525, N276);
buf BUF1 (N554, N547);
nor NOR4 (N555, N542, N189, N66, N277);
nand NAND2 (N556, N544, N410);
not NOT1 (N557, N556);
nor NOR3 (N558, N534, N210, N121);
nor NOR3 (N559, N554, N190, N258);
nand NAND4 (N560, N557, N354, N405, N79);
nand NAND4 (N561, N560, N155, N294, N48);
buf BUF1 (N562, N559);
not NOT1 (N563, N548);
nand NAND4 (N564, N549, N220, N504, N318);
nor NOR3 (N565, N553, N48, N40);
nor NOR2 (N566, N565, N459);
nor NOR2 (N567, N550, N72);
or OR4 (N568, N558, N186, N540, N351);
xor XOR2 (N569, N555, N78);
nand NAND2 (N570, N551, N373);
nand NAND4 (N571, N570, N148, N247, N497);
and AND2 (N572, N568, N521);
or OR2 (N573, N572, N213);
or OR3 (N574, N564, N140, N458);
or OR3 (N575, N561, N522, N262);
and AND3 (N576, N566, N384, N358);
nor NOR3 (N577, N571, N43, N21);
not NOT1 (N578, N562);
nor NOR3 (N579, N574, N549, N208);
or OR4 (N580, N577, N447, N551, N494);
xor XOR2 (N581, N575, N200);
xor XOR2 (N582, N581, N450);
xor XOR2 (N583, N569, N578);
nor NOR4 (N584, N339, N172, N318, N93);
nand NAND4 (N585, N552, N353, N498, N214);
xor XOR2 (N586, N576, N205);
nand NAND4 (N587, N586, N328, N299, N308);
nor NOR3 (N588, N573, N218, N547);
or OR3 (N589, N582, N349, N56);
and AND3 (N590, N580, N535, N130);
buf BUF1 (N591, N579);
or OR3 (N592, N584, N233, N549);
or OR4 (N593, N588, N239, N489, N352);
not NOT1 (N594, N592);
not NOT1 (N595, N591);
or OR2 (N596, N590, N62);
and AND4 (N597, N596, N235, N320, N536);
not NOT1 (N598, N589);
not NOT1 (N599, N583);
xor XOR2 (N600, N585, N202);
and AND3 (N601, N567, N203, N252);
xor XOR2 (N602, N593, N421);
or OR3 (N603, N602, N218, N260);
and AND4 (N604, N587, N166, N16, N287);
buf BUF1 (N605, N599);
nand NAND2 (N606, N600, N137);
xor XOR2 (N607, N595, N601);
nor NOR3 (N608, N120, N607, N231);
and AND3 (N609, N581, N140, N19);
buf BUF1 (N610, N563);
buf BUF1 (N611, N609);
or OR2 (N612, N594, N36);
and AND3 (N613, N597, N365, N416);
not NOT1 (N614, N608);
or OR3 (N615, N606, N614, N594);
buf BUF1 (N616, N501);
not NOT1 (N617, N603);
xor XOR2 (N618, N613, N452);
not NOT1 (N619, N605);
or OR2 (N620, N610, N557);
not NOT1 (N621, N619);
and AND4 (N622, N620, N490, N100, N406);
nor NOR2 (N623, N617, N424);
nand NAND4 (N624, N616, N340, N90, N530);
and AND3 (N625, N624, N284, N518);
not NOT1 (N626, N604);
buf BUF1 (N627, N598);
xor XOR2 (N628, N621, N608);
buf BUF1 (N629, N628);
nand NAND4 (N630, N626, N256, N251, N495);
nor NOR3 (N631, N629, N304, N452);
nand NAND2 (N632, N627, N406);
and AND2 (N633, N632, N419);
buf BUF1 (N634, N615);
and AND3 (N635, N622, N108, N521);
and AND2 (N636, N611, N48);
xor XOR2 (N637, N625, N131);
not NOT1 (N638, N623);
nand NAND3 (N639, N633, N568, N194);
nand NAND3 (N640, N636, N512, N293);
nor NOR4 (N641, N640, N637, N114, N389);
buf BUF1 (N642, N7);
and AND3 (N643, N631, N259, N405);
xor XOR2 (N644, N630, N267);
not NOT1 (N645, N641);
not NOT1 (N646, N618);
and AND2 (N647, N643, N415);
and AND2 (N648, N635, N395);
or OR4 (N649, N634, N574, N32, N160);
nand NAND3 (N650, N645, N37, N138);
xor XOR2 (N651, N647, N526);
and AND3 (N652, N638, N570, N233);
nor NOR4 (N653, N646, N201, N205, N243);
or OR2 (N654, N648, N388);
nand NAND2 (N655, N639, N374);
xor XOR2 (N656, N654, N413);
not NOT1 (N657, N644);
or OR3 (N658, N649, N420, N470);
xor XOR2 (N659, N653, N287);
buf BUF1 (N660, N612);
nand NAND2 (N661, N660, N67);
nand NAND2 (N662, N655, N567);
xor XOR2 (N663, N662, N425);
buf BUF1 (N664, N652);
nand NAND4 (N665, N650, N258, N172, N395);
nor NOR3 (N666, N664, N532, N231);
nor NOR4 (N667, N642, N567, N593, N178);
nand NAND2 (N668, N656, N328);
xor XOR2 (N669, N658, N264);
xor XOR2 (N670, N668, N307);
and AND2 (N671, N667, N629);
xor XOR2 (N672, N670, N535);
nand NAND4 (N673, N659, N582, N594, N432);
xor XOR2 (N674, N657, N19);
nor NOR3 (N675, N674, N543, N339);
nand NAND3 (N676, N663, N134, N100);
xor XOR2 (N677, N669, N580);
nand NAND3 (N678, N675, N559, N77);
or OR2 (N679, N666, N478);
not NOT1 (N680, N671);
nor NOR2 (N681, N672, N164);
or OR3 (N682, N677, N542, N35);
and AND3 (N683, N651, N578, N92);
xor XOR2 (N684, N682, N207);
xor XOR2 (N685, N681, N179);
nand NAND4 (N686, N665, N676, N120, N670);
or OR4 (N687, N357, N622, N407, N533);
not NOT1 (N688, N684);
not NOT1 (N689, N680);
buf BUF1 (N690, N688);
not NOT1 (N691, N679);
and AND4 (N692, N686, N534, N159, N684);
xor XOR2 (N693, N687, N464);
xor XOR2 (N694, N690, N553);
buf BUF1 (N695, N693);
nor NOR3 (N696, N683, N527, N223);
xor XOR2 (N697, N691, N543);
or OR3 (N698, N678, N635, N357);
nand NAND2 (N699, N661, N18);
or OR3 (N700, N685, N336, N578);
not NOT1 (N701, N700);
not NOT1 (N702, N698);
nand NAND3 (N703, N699, N596, N67);
or OR2 (N704, N695, N177);
nor NOR3 (N705, N703, N692, N335);
buf BUF1 (N706, N680);
buf BUF1 (N707, N702);
nor NOR2 (N708, N707, N121);
xor XOR2 (N709, N689, N684);
nand NAND4 (N710, N697, N203, N582, N411);
buf BUF1 (N711, N694);
and AND3 (N712, N701, N542, N525);
or OR4 (N713, N712, N697, N54, N313);
nand NAND4 (N714, N709, N399, N585, N252);
or OR3 (N715, N705, N693, N470);
and AND4 (N716, N696, N598, N122, N565);
nand NAND2 (N717, N706, N573);
or OR3 (N718, N714, N283, N48);
and AND4 (N719, N673, N120, N39, N480);
nand NAND3 (N720, N717, N362, N442);
xor XOR2 (N721, N715, N155);
and AND2 (N722, N710, N362);
not NOT1 (N723, N721);
or OR4 (N724, N711, N5, N666, N523);
or OR4 (N725, N720, N39, N4, N454);
buf BUF1 (N726, N704);
or OR4 (N727, N722, N334, N400, N141);
nand NAND4 (N728, N725, N448, N561, N499);
not NOT1 (N729, N723);
buf BUF1 (N730, N728);
and AND2 (N731, N718, N384);
buf BUF1 (N732, N730);
and AND4 (N733, N729, N487, N432, N564);
xor XOR2 (N734, N716, N605);
nor NOR3 (N735, N734, N427, N584);
xor XOR2 (N736, N719, N50);
not NOT1 (N737, N726);
nand NAND3 (N738, N735, N551, N494);
not NOT1 (N739, N708);
nand NAND3 (N740, N727, N26, N523);
buf BUF1 (N741, N736);
not NOT1 (N742, N713);
nand NAND2 (N743, N740, N213);
not NOT1 (N744, N739);
buf BUF1 (N745, N741);
not NOT1 (N746, N724);
buf BUF1 (N747, N732);
xor XOR2 (N748, N744, N290);
or OR4 (N749, N737, N433, N373, N315);
buf BUF1 (N750, N738);
not NOT1 (N751, N749);
buf BUF1 (N752, N733);
or OR2 (N753, N731, N621);
or OR4 (N754, N751, N25, N686, N538);
nand NAND3 (N755, N743, N83, N67);
xor XOR2 (N756, N753, N7);
and AND3 (N757, N748, N162, N488);
and AND2 (N758, N755, N128);
and AND3 (N759, N747, N566, N318);
and AND3 (N760, N745, N108, N114);
not NOT1 (N761, N758);
not NOT1 (N762, N761);
or OR4 (N763, N752, N446, N313, N505);
xor XOR2 (N764, N754, N381);
xor XOR2 (N765, N760, N168);
or OR2 (N766, N757, N548);
nor NOR4 (N767, N756, N239, N551, N609);
xor XOR2 (N768, N764, N474);
or OR2 (N769, N750, N516);
or OR4 (N770, N759, N511, N209, N720);
and AND3 (N771, N765, N523, N321);
and AND2 (N772, N770, N75);
xor XOR2 (N773, N742, N171);
buf BUF1 (N774, N768);
nand NAND4 (N775, N767, N489, N369, N673);
or OR2 (N776, N774, N437);
nand NAND2 (N777, N771, N117);
not NOT1 (N778, N773);
buf BUF1 (N779, N766);
nor NOR3 (N780, N763, N217, N520);
nand NAND2 (N781, N778, N236);
buf BUF1 (N782, N777);
xor XOR2 (N783, N769, N40);
or OR3 (N784, N782, N442, N506);
xor XOR2 (N785, N779, N218);
xor XOR2 (N786, N784, N191);
buf BUF1 (N787, N775);
nor NOR2 (N788, N785, N566);
nand NAND3 (N789, N776, N302, N555);
xor XOR2 (N790, N788, N154);
buf BUF1 (N791, N772);
not NOT1 (N792, N791);
and AND4 (N793, N789, N12, N437, N68);
nand NAND2 (N794, N781, N308);
nand NAND4 (N795, N793, N191, N311, N140);
or OR2 (N796, N786, N725);
or OR2 (N797, N794, N145);
nand NAND4 (N798, N795, N557, N482, N678);
or OR4 (N799, N798, N495, N153, N57);
not NOT1 (N800, N783);
buf BUF1 (N801, N790);
xor XOR2 (N802, N746, N707);
nor NOR2 (N803, N801, N481);
and AND2 (N804, N799, N538);
buf BUF1 (N805, N796);
nand NAND3 (N806, N780, N134, N399);
xor XOR2 (N807, N805, N793);
buf BUF1 (N808, N804);
and AND3 (N809, N800, N129, N121);
nor NOR4 (N810, N792, N550, N59, N313);
buf BUF1 (N811, N787);
not NOT1 (N812, N803);
not NOT1 (N813, N812);
xor XOR2 (N814, N802, N808);
buf BUF1 (N815, N779);
not NOT1 (N816, N811);
or OR2 (N817, N813, N562);
not NOT1 (N818, N817);
not NOT1 (N819, N762);
or OR3 (N820, N816, N369, N58);
nor NOR3 (N821, N819, N695, N471);
not NOT1 (N822, N809);
nor NOR4 (N823, N815, N705, N439, N747);
or OR2 (N824, N810, N597);
xor XOR2 (N825, N823, N63);
not NOT1 (N826, N822);
nand NAND4 (N827, N807, N739, N307, N780);
nor NOR4 (N828, N806, N534, N281, N503);
not NOT1 (N829, N821);
nand NAND3 (N830, N829, N723, N110);
nand NAND4 (N831, N797, N431, N424, N433);
nand NAND3 (N832, N830, N426, N828);
xor XOR2 (N833, N813, N621);
not NOT1 (N834, N825);
nor NOR3 (N835, N834, N617, N640);
or OR2 (N836, N824, N807);
nand NAND2 (N837, N831, N547);
xor XOR2 (N838, N833, N302);
buf BUF1 (N839, N837);
or OR4 (N840, N832, N8, N485, N699);
not NOT1 (N841, N826);
and AND3 (N842, N818, N790, N704);
xor XOR2 (N843, N840, N433);
nand NAND2 (N844, N814, N775);
not NOT1 (N845, N839);
buf BUF1 (N846, N836);
nand NAND4 (N847, N846, N190, N32, N484);
not NOT1 (N848, N841);
and AND4 (N849, N835, N708, N722, N85);
nand NAND2 (N850, N849, N513);
buf BUF1 (N851, N820);
buf BUF1 (N852, N843);
xor XOR2 (N853, N847, N807);
and AND4 (N854, N842, N20, N532, N370);
or OR3 (N855, N850, N347, N253);
nor NOR2 (N856, N845, N375);
nor NOR3 (N857, N827, N397, N640);
buf BUF1 (N858, N855);
or OR4 (N859, N853, N12, N106, N814);
buf BUF1 (N860, N858);
not NOT1 (N861, N852);
or OR4 (N862, N860, N211, N376, N135);
nand NAND2 (N863, N856, N100);
nand NAND3 (N864, N854, N789, N154);
not NOT1 (N865, N857);
nor NOR4 (N866, N863, N855, N388, N655);
xor XOR2 (N867, N851, N87);
nand NAND2 (N868, N848, N308);
nor NOR2 (N869, N865, N266);
or OR4 (N870, N861, N181, N231, N422);
or OR3 (N871, N862, N433, N448);
buf BUF1 (N872, N866);
xor XOR2 (N873, N869, N371);
nor NOR4 (N874, N873, N730, N6, N792);
nor NOR2 (N875, N874, N373);
and AND2 (N876, N875, N352);
not NOT1 (N877, N864);
xor XOR2 (N878, N871, N829);
nor NOR2 (N879, N859, N823);
and AND2 (N880, N876, N156);
buf BUF1 (N881, N838);
and AND3 (N882, N878, N522, N481);
xor XOR2 (N883, N872, N263);
nand NAND3 (N884, N867, N91, N48);
and AND2 (N885, N868, N269);
buf BUF1 (N886, N844);
buf BUF1 (N887, N883);
buf BUF1 (N888, N886);
nor NOR2 (N889, N885, N89);
nand NAND2 (N890, N888, N485);
nand NAND3 (N891, N887, N688, N647);
and AND2 (N892, N877, N729);
nand NAND4 (N893, N879, N32, N396, N352);
xor XOR2 (N894, N890, N217);
or OR3 (N895, N870, N749, N554);
buf BUF1 (N896, N884);
and AND4 (N897, N889, N513, N331, N680);
xor XOR2 (N898, N880, N820);
and AND4 (N899, N882, N498, N639, N353);
nand NAND3 (N900, N897, N732, N681);
xor XOR2 (N901, N896, N369);
nand NAND4 (N902, N892, N594, N145, N20);
not NOT1 (N903, N900);
buf BUF1 (N904, N903);
or OR4 (N905, N902, N610, N393, N771);
buf BUF1 (N906, N893);
buf BUF1 (N907, N901);
or OR4 (N908, N904, N403, N261, N119);
nor NOR3 (N909, N891, N308, N848);
buf BUF1 (N910, N898);
not NOT1 (N911, N905);
or OR2 (N912, N907, N89);
or OR3 (N913, N909, N674, N574);
nor NOR2 (N914, N910, N738);
nand NAND3 (N915, N881, N320, N867);
xor XOR2 (N916, N915, N389);
buf BUF1 (N917, N899);
nor NOR4 (N918, N911, N464, N209, N837);
not NOT1 (N919, N912);
nor NOR3 (N920, N918, N710, N450);
nor NOR3 (N921, N914, N27, N862);
nor NOR3 (N922, N919, N581, N842);
nand NAND2 (N923, N895, N557);
nand NAND2 (N924, N906, N662);
nand NAND4 (N925, N923, N184, N516, N505);
nand NAND2 (N926, N894, N337);
nand NAND4 (N927, N921, N751, N148, N557);
not NOT1 (N928, N927);
nand NAND2 (N929, N913, N490);
xor XOR2 (N930, N917, N387);
not NOT1 (N931, N922);
nor NOR2 (N932, N924, N252);
xor XOR2 (N933, N930, N712);
or OR3 (N934, N920, N814, N66);
not NOT1 (N935, N934);
buf BUF1 (N936, N931);
or OR2 (N937, N928, N291);
or OR4 (N938, N908, N868, N116, N383);
and AND3 (N939, N936, N521, N489);
buf BUF1 (N940, N939);
nor NOR4 (N941, N933, N312, N419, N216);
buf BUF1 (N942, N937);
xor XOR2 (N943, N929, N318);
nor NOR4 (N944, N942, N85, N160, N59);
or OR4 (N945, N925, N459, N475, N158);
or OR4 (N946, N935, N154, N3, N235);
and AND2 (N947, N932, N162);
or OR2 (N948, N926, N901);
or OR2 (N949, N947, N550);
and AND2 (N950, N916, N134);
nor NOR2 (N951, N946, N843);
and AND2 (N952, N949, N776);
or OR4 (N953, N952, N603, N663, N642);
and AND4 (N954, N953, N294, N466, N306);
or OR2 (N955, N945, N213);
or OR4 (N956, N954, N788, N223, N878);
or OR2 (N957, N951, N686);
or OR4 (N958, N957, N558, N464, N598);
or OR3 (N959, N948, N484, N395);
nor NOR4 (N960, N940, N696, N882, N546);
not NOT1 (N961, N956);
or OR2 (N962, N955, N508);
buf BUF1 (N963, N960);
xor XOR2 (N964, N941, N877);
nor NOR3 (N965, N943, N469, N820);
nand NAND3 (N966, N950, N575, N314);
xor XOR2 (N967, N966, N441);
nor NOR3 (N968, N965, N431, N692);
xor XOR2 (N969, N944, N899);
and AND3 (N970, N964, N218, N489);
or OR4 (N971, N963, N212, N406, N756);
not NOT1 (N972, N938);
nor NOR4 (N973, N958, N775, N879, N730);
nand NAND3 (N974, N961, N477, N265);
buf BUF1 (N975, N959);
and AND4 (N976, N974, N847, N266, N70);
and AND3 (N977, N967, N731, N850);
or OR2 (N978, N977, N873);
or OR4 (N979, N978, N625, N453, N430);
not NOT1 (N980, N962);
buf BUF1 (N981, N971);
xor XOR2 (N982, N969, N585);
buf BUF1 (N983, N976);
and AND2 (N984, N973, N491);
buf BUF1 (N985, N983);
nand NAND3 (N986, N985, N144, N868);
or OR2 (N987, N986, N945);
not NOT1 (N988, N968);
buf BUF1 (N989, N988);
not NOT1 (N990, N972);
not NOT1 (N991, N990);
nand NAND2 (N992, N989, N315);
not NOT1 (N993, N979);
and AND4 (N994, N993, N29, N902, N776);
nor NOR4 (N995, N981, N301, N939, N789);
nor NOR3 (N996, N975, N290, N362);
and AND2 (N997, N996, N844);
nand NAND2 (N998, N992, N977);
nor NOR2 (N999, N982, N875);
nand NAND2 (N1000, N991, N179);
nand NAND3 (N1001, N998, N821, N522);
nor NOR2 (N1002, N999, N931);
buf BUF1 (N1003, N1000);
and AND4 (N1004, N980, N982, N902, N907);
nand NAND2 (N1005, N987, N343);
buf BUF1 (N1006, N994);
nor NOR3 (N1007, N1005, N91, N223);
xor XOR2 (N1008, N995, N808);
or OR3 (N1009, N1004, N242, N721);
xor XOR2 (N1010, N1001, N719);
and AND4 (N1011, N1006, N877, N273, N398);
buf BUF1 (N1012, N1002);
not NOT1 (N1013, N970);
or OR3 (N1014, N1010, N778, N825);
nor NOR3 (N1015, N1013, N832, N908);
xor XOR2 (N1016, N1009, N450);
buf BUF1 (N1017, N1008);
or OR2 (N1018, N1017, N479);
buf BUF1 (N1019, N1016);
not NOT1 (N1020, N1003);
not NOT1 (N1021, N1020);
buf BUF1 (N1022, N1014);
nand NAND4 (N1023, N1015, N711, N605, N542);
buf BUF1 (N1024, N1018);
xor XOR2 (N1025, N1007, N605);
nor NOR4 (N1026, N1023, N638, N837, N907);
or OR3 (N1027, N1025, N199, N783);
not NOT1 (N1028, N1019);
and AND2 (N1029, N984, N264);
not NOT1 (N1030, N1024);
xor XOR2 (N1031, N1022, N267);
buf BUF1 (N1032, N1012);
xor XOR2 (N1033, N1027, N218);
buf BUF1 (N1034, N997);
nand NAND2 (N1035, N1034, N545);
and AND2 (N1036, N1035, N937);
xor XOR2 (N1037, N1021, N905);
buf BUF1 (N1038, N1011);
buf BUF1 (N1039, N1029);
or OR3 (N1040, N1028, N278, N599);
not NOT1 (N1041, N1038);
nor NOR4 (N1042, N1040, N643, N83, N953);
and AND3 (N1043, N1039, N21, N933);
xor XOR2 (N1044, N1026, N339);
or OR3 (N1045, N1033, N459, N1001);
and AND2 (N1046, N1044, N111);
buf BUF1 (N1047, N1036);
buf BUF1 (N1048, N1045);
nand NAND3 (N1049, N1041, N849, N739);
and AND2 (N1050, N1042, N109);
xor XOR2 (N1051, N1043, N974);
nand NAND4 (N1052, N1050, N274, N1002, N292);
not NOT1 (N1053, N1046);
xor XOR2 (N1054, N1049, N103);
xor XOR2 (N1055, N1054, N554);
nand NAND4 (N1056, N1052, N901, N724, N837);
or OR3 (N1057, N1048, N874, N553);
buf BUF1 (N1058, N1047);
buf BUF1 (N1059, N1037);
or OR3 (N1060, N1055, N803, N28);
nand NAND3 (N1061, N1053, N408, N626);
xor XOR2 (N1062, N1030, N1054);
nor NOR4 (N1063, N1062, N672, N284, N685);
nand NAND2 (N1064, N1059, N878);
xor XOR2 (N1065, N1031, N1041);
nand NAND2 (N1066, N1056, N69);
nor NOR2 (N1067, N1058, N746);
or OR4 (N1068, N1066, N278, N356, N1003);
not NOT1 (N1069, N1032);
xor XOR2 (N1070, N1064, N817);
or OR3 (N1071, N1067, N670, N1021);
or OR3 (N1072, N1071, N153, N518);
and AND3 (N1073, N1065, N1015, N119);
or OR4 (N1074, N1072, N523, N1073, N929);
and AND4 (N1075, N1016, N896, N235, N635);
and AND2 (N1076, N1068, N409);
nor NOR2 (N1077, N1075, N55);
and AND2 (N1078, N1060, N327);
buf BUF1 (N1079, N1078);
and AND3 (N1080, N1070, N340, N64);
and AND2 (N1081, N1079, N157);
buf BUF1 (N1082, N1051);
nor NOR2 (N1083, N1069, N83);
or OR2 (N1084, N1074, N1019);
or OR3 (N1085, N1076, N306, N610);
buf BUF1 (N1086, N1063);
xor XOR2 (N1087, N1084, N446);
or OR3 (N1088, N1081, N635, N768);
buf BUF1 (N1089, N1083);
not NOT1 (N1090, N1085);
nor NOR4 (N1091, N1088, N603, N701, N128);
nor NOR3 (N1092, N1086, N1024, N654);
or OR2 (N1093, N1077, N12);
not NOT1 (N1094, N1087);
and AND2 (N1095, N1061, N396);
nand NAND4 (N1096, N1091, N511, N297, N29);
xor XOR2 (N1097, N1093, N601);
or OR2 (N1098, N1097, N374);
or OR2 (N1099, N1090, N1016);
nor NOR3 (N1100, N1082, N264, N884);
nor NOR3 (N1101, N1099, N694, N23);
nand NAND2 (N1102, N1100, N461);
nand NAND3 (N1103, N1096, N268, N903);
nor NOR3 (N1104, N1102, N138, N612);
or OR4 (N1105, N1080, N223, N532, N619);
and AND4 (N1106, N1103, N295, N229, N141);
buf BUF1 (N1107, N1092);
xor XOR2 (N1108, N1098, N491);
xor XOR2 (N1109, N1101, N572);
not NOT1 (N1110, N1095);
xor XOR2 (N1111, N1106, N788);
nor NOR4 (N1112, N1107, N835, N756, N713);
nand NAND4 (N1113, N1104, N540, N667, N612);
and AND3 (N1114, N1109, N52, N772);
and AND3 (N1115, N1094, N1003, N1069);
buf BUF1 (N1116, N1111);
nand NAND4 (N1117, N1112, N984, N851, N251);
buf BUF1 (N1118, N1110);
not NOT1 (N1119, N1089);
or OR3 (N1120, N1108, N507, N803);
nor NOR4 (N1121, N1114, N132, N344, N834);
nand NAND4 (N1122, N1113, N699, N968, N405);
nand NAND4 (N1123, N1057, N950, N988, N711);
xor XOR2 (N1124, N1122, N480);
or OR3 (N1125, N1121, N525, N42);
or OR4 (N1126, N1119, N738, N299, N206);
not NOT1 (N1127, N1105);
not NOT1 (N1128, N1120);
not NOT1 (N1129, N1126);
nand NAND2 (N1130, N1118, N8);
and AND2 (N1131, N1125, N694);
buf BUF1 (N1132, N1116);
xor XOR2 (N1133, N1129, N1031);
buf BUF1 (N1134, N1124);
and AND3 (N1135, N1127, N1118, N5);
not NOT1 (N1136, N1135);
not NOT1 (N1137, N1130);
buf BUF1 (N1138, N1128);
buf BUF1 (N1139, N1134);
not NOT1 (N1140, N1117);
not NOT1 (N1141, N1115);
xor XOR2 (N1142, N1132, N181);
or OR2 (N1143, N1137, N625);
and AND4 (N1144, N1139, N937, N293, N465);
nor NOR3 (N1145, N1123, N107, N108);
buf BUF1 (N1146, N1140);
not NOT1 (N1147, N1141);
or OR3 (N1148, N1145, N857, N380);
or OR3 (N1149, N1138, N841, N470);
nand NAND2 (N1150, N1136, N451);
or OR3 (N1151, N1144, N782, N21);
not NOT1 (N1152, N1146);
xor XOR2 (N1153, N1131, N644);
nor NOR2 (N1154, N1143, N1027);
xor XOR2 (N1155, N1154, N1034);
xor XOR2 (N1156, N1153, N645);
and AND3 (N1157, N1147, N661, N839);
xor XOR2 (N1158, N1151, N344);
not NOT1 (N1159, N1142);
and AND3 (N1160, N1133, N191, N705);
or OR4 (N1161, N1157, N482, N1, N88);
or OR4 (N1162, N1155, N744, N585, N690);
or OR4 (N1163, N1160, N422, N415, N91);
nand NAND3 (N1164, N1156, N889, N761);
xor XOR2 (N1165, N1150, N845);
buf BUF1 (N1166, N1149);
xor XOR2 (N1167, N1165, N363);
nand NAND4 (N1168, N1161, N1019, N255, N524);
or OR4 (N1169, N1168, N168, N504, N282);
buf BUF1 (N1170, N1167);
or OR2 (N1171, N1169, N383);
and AND4 (N1172, N1158, N1140, N321, N652);
and AND4 (N1173, N1163, N671, N483, N996);
and AND4 (N1174, N1159, N621, N1095, N931);
xor XOR2 (N1175, N1170, N359);
and AND4 (N1176, N1148, N126, N155, N420);
not NOT1 (N1177, N1164);
nand NAND2 (N1178, N1172, N836);
and AND3 (N1179, N1177, N305, N300);
not NOT1 (N1180, N1166);
and AND3 (N1181, N1162, N705, N454);
buf BUF1 (N1182, N1152);
nor NOR3 (N1183, N1178, N139, N276);
and AND4 (N1184, N1173, N328, N416, N78);
buf BUF1 (N1185, N1184);
and AND4 (N1186, N1182, N1132, N231, N592);
nor NOR3 (N1187, N1185, N619, N352);
nor NOR4 (N1188, N1175, N949, N459, N133);
not NOT1 (N1189, N1183);
xor XOR2 (N1190, N1171, N869);
not NOT1 (N1191, N1180);
and AND2 (N1192, N1186, N1041);
xor XOR2 (N1193, N1181, N332);
buf BUF1 (N1194, N1188);
nor NOR2 (N1195, N1194, N207);
nand NAND2 (N1196, N1192, N1064);
not NOT1 (N1197, N1195);
or OR2 (N1198, N1176, N564);
buf BUF1 (N1199, N1193);
not NOT1 (N1200, N1199);
and AND4 (N1201, N1189, N634, N106, N841);
buf BUF1 (N1202, N1174);
buf BUF1 (N1203, N1191);
nor NOR3 (N1204, N1179, N1198, N885);
xor XOR2 (N1205, N308, N406);
nand NAND3 (N1206, N1190, N1179, N507);
not NOT1 (N1207, N1206);
xor XOR2 (N1208, N1200, N524);
not NOT1 (N1209, N1208);
not NOT1 (N1210, N1187);
and AND2 (N1211, N1207, N878);
nor NOR4 (N1212, N1201, N746, N730, N1124);
buf BUF1 (N1213, N1211);
or OR3 (N1214, N1197, N810, N474);
not NOT1 (N1215, N1202);
buf BUF1 (N1216, N1196);
or OR2 (N1217, N1205, N24);
buf BUF1 (N1218, N1213);
nand NAND2 (N1219, N1210, N851);
nand NAND2 (N1220, N1219, N348);
xor XOR2 (N1221, N1209, N627);
not NOT1 (N1222, N1204);
nand NAND4 (N1223, N1218, N210, N528, N250);
nand NAND4 (N1224, N1215, N253, N190, N529);
nand NAND3 (N1225, N1217, N556, N632);
xor XOR2 (N1226, N1224, N1131);
xor XOR2 (N1227, N1223, N188);
not NOT1 (N1228, N1214);
buf BUF1 (N1229, N1227);
or OR4 (N1230, N1203, N99, N134, N474);
nand NAND2 (N1231, N1228, N1064);
nor NOR2 (N1232, N1216, N749);
nand NAND3 (N1233, N1220, N812, N385);
nand NAND3 (N1234, N1225, N615, N1202);
nor NOR4 (N1235, N1229, N263, N1094, N1158);
or OR2 (N1236, N1235, N227);
or OR4 (N1237, N1226, N44, N477, N1219);
nand NAND3 (N1238, N1221, N445, N747);
nand NAND3 (N1239, N1232, N932, N966);
xor XOR2 (N1240, N1212, N1193);
or OR4 (N1241, N1238, N408, N124, N217);
and AND3 (N1242, N1231, N854, N225);
and AND3 (N1243, N1240, N391, N641);
nor NOR4 (N1244, N1230, N758, N202, N451);
xor XOR2 (N1245, N1239, N272);
not NOT1 (N1246, N1234);
nand NAND4 (N1247, N1233, N883, N821, N465);
and AND3 (N1248, N1241, N808, N259);
nor NOR2 (N1249, N1245, N734);
nand NAND4 (N1250, N1247, N142, N529, N974);
or OR4 (N1251, N1237, N396, N457, N235);
and AND3 (N1252, N1248, N418, N32);
or OR4 (N1253, N1242, N1138, N1206, N272);
nand NAND3 (N1254, N1249, N809, N83);
not NOT1 (N1255, N1244);
or OR3 (N1256, N1246, N758, N751);
not NOT1 (N1257, N1251);
xor XOR2 (N1258, N1256, N49);
and AND2 (N1259, N1253, N732);
buf BUF1 (N1260, N1257);
nor NOR3 (N1261, N1250, N1092, N580);
xor XOR2 (N1262, N1236, N1186);
not NOT1 (N1263, N1243);
xor XOR2 (N1264, N1254, N312);
buf BUF1 (N1265, N1260);
not NOT1 (N1266, N1265);
xor XOR2 (N1267, N1262, N784);
not NOT1 (N1268, N1267);
not NOT1 (N1269, N1268);
and AND3 (N1270, N1261, N565, N115);
nor NOR2 (N1271, N1259, N1268);
nor NOR3 (N1272, N1270, N679, N1144);
and AND2 (N1273, N1258, N599);
buf BUF1 (N1274, N1269);
buf BUF1 (N1275, N1272);
nor NOR2 (N1276, N1274, N1245);
nor NOR4 (N1277, N1271, N1163, N930, N1121);
xor XOR2 (N1278, N1277, N468);
buf BUF1 (N1279, N1273);
not NOT1 (N1280, N1276);
and AND4 (N1281, N1278, N1031, N249, N692);
buf BUF1 (N1282, N1266);
not NOT1 (N1283, N1264);
nor NOR2 (N1284, N1263, N498);
not NOT1 (N1285, N1255);
xor XOR2 (N1286, N1281, N414);
nor NOR4 (N1287, N1284, N1095, N512, N297);
buf BUF1 (N1288, N1285);
xor XOR2 (N1289, N1282, N1201);
buf BUF1 (N1290, N1222);
xor XOR2 (N1291, N1252, N1252);
nand NAND4 (N1292, N1283, N435, N478, N314);
not NOT1 (N1293, N1291);
buf BUF1 (N1294, N1279);
or OR3 (N1295, N1294, N927, N277);
nand NAND3 (N1296, N1290, N965, N54);
or OR3 (N1297, N1295, N711, N991);
xor XOR2 (N1298, N1275, N42);
and AND4 (N1299, N1293, N88, N988, N408);
nand NAND2 (N1300, N1297, N953);
not NOT1 (N1301, N1288);
and AND4 (N1302, N1296, N874, N1125, N346);
xor XOR2 (N1303, N1302, N223);
nor NOR2 (N1304, N1289, N1221);
not NOT1 (N1305, N1287);
or OR4 (N1306, N1298, N553, N75, N1138);
nand NAND2 (N1307, N1286, N597);
buf BUF1 (N1308, N1306);
nor NOR3 (N1309, N1307, N1078, N1084);
nand NAND4 (N1310, N1308, N267, N494, N529);
nor NOR4 (N1311, N1280, N767, N784, N841);
nor NOR3 (N1312, N1299, N715, N1301);
nor NOR2 (N1313, N1016, N1139);
xor XOR2 (N1314, N1300, N1268);
xor XOR2 (N1315, N1312, N382);
nor NOR2 (N1316, N1310, N1155);
or OR4 (N1317, N1311, N724, N605, N1108);
xor XOR2 (N1318, N1314, N381);
and AND2 (N1319, N1318, N920);
xor XOR2 (N1320, N1313, N1021);
or OR3 (N1321, N1305, N396, N857);
nand NAND4 (N1322, N1292, N1127, N672, N217);
or OR2 (N1323, N1317, N1132);
and AND2 (N1324, N1316, N922);
nand NAND4 (N1325, N1315, N525, N974, N588);
and AND2 (N1326, N1304, N883);
nor NOR2 (N1327, N1325, N397);
nor NOR2 (N1328, N1324, N552);
nor NOR3 (N1329, N1326, N1048, N92);
and AND4 (N1330, N1319, N10, N192, N353);
xor XOR2 (N1331, N1327, N793);
or OR3 (N1332, N1321, N935, N959);
nand NAND3 (N1333, N1330, N562, N1304);
and AND3 (N1334, N1332, N197, N898);
nor NOR3 (N1335, N1329, N415, N473);
not NOT1 (N1336, N1328);
buf BUF1 (N1337, N1320);
buf BUF1 (N1338, N1333);
buf BUF1 (N1339, N1331);
nor NOR2 (N1340, N1303, N1097);
or OR2 (N1341, N1322, N140);
buf BUF1 (N1342, N1338);
xor XOR2 (N1343, N1339, N1031);
nor NOR3 (N1344, N1343, N44, N646);
xor XOR2 (N1345, N1323, N80);
xor XOR2 (N1346, N1345, N1085);
nor NOR4 (N1347, N1341, N1305, N353, N362);
nor NOR2 (N1348, N1342, N1342);
buf BUF1 (N1349, N1309);
and AND3 (N1350, N1344, N1247, N48);
not NOT1 (N1351, N1336);
and AND3 (N1352, N1349, N1047, N633);
nand NAND2 (N1353, N1334, N741);
or OR4 (N1354, N1350, N68, N585, N824);
xor XOR2 (N1355, N1352, N1190);
or OR4 (N1356, N1340, N1134, N1125, N137);
buf BUF1 (N1357, N1355);
nand NAND2 (N1358, N1354, N139);
or OR2 (N1359, N1347, N908);
buf BUF1 (N1360, N1353);
nand NAND3 (N1361, N1358, N745, N527);
not NOT1 (N1362, N1359);
buf BUF1 (N1363, N1337);
and AND3 (N1364, N1351, N434, N1203);
not NOT1 (N1365, N1364);
nor NOR4 (N1366, N1363, N418, N194, N690);
nor NOR4 (N1367, N1346, N1178, N311, N1191);
nand NAND4 (N1368, N1357, N982, N1132, N580);
not NOT1 (N1369, N1368);
nor NOR2 (N1370, N1361, N259);
buf BUF1 (N1371, N1348);
and AND2 (N1372, N1360, N274);
xor XOR2 (N1373, N1369, N185);
nand NAND2 (N1374, N1356, N1065);
xor XOR2 (N1375, N1370, N683);
and AND4 (N1376, N1372, N1245, N1174, N230);
and AND4 (N1377, N1366, N250, N711, N603);
not NOT1 (N1378, N1375);
nor NOR3 (N1379, N1367, N767, N1094);
nor NOR2 (N1380, N1362, N722);
not NOT1 (N1381, N1374);
not NOT1 (N1382, N1365);
nor NOR2 (N1383, N1377, N881);
nand NAND3 (N1384, N1380, N704, N798);
nor NOR4 (N1385, N1378, N1086, N248, N290);
not NOT1 (N1386, N1376);
buf BUF1 (N1387, N1379);
buf BUF1 (N1388, N1381);
or OR2 (N1389, N1383, N628);
buf BUF1 (N1390, N1384);
and AND3 (N1391, N1371, N314, N654);
not NOT1 (N1392, N1391);
and AND4 (N1393, N1373, N1175, N1135, N23);
buf BUF1 (N1394, N1387);
buf BUF1 (N1395, N1392);
not NOT1 (N1396, N1395);
buf BUF1 (N1397, N1385);
and AND2 (N1398, N1394, N519);
or OR4 (N1399, N1388, N630, N755, N354);
nor NOR3 (N1400, N1399, N23, N347);
nor NOR4 (N1401, N1398, N795, N1205, N967);
or OR4 (N1402, N1382, N1332, N1037, N711);
nand NAND4 (N1403, N1390, N227, N440, N1190);
and AND2 (N1404, N1401, N493);
buf BUF1 (N1405, N1404);
not NOT1 (N1406, N1393);
buf BUF1 (N1407, N1402);
not NOT1 (N1408, N1396);
nand NAND4 (N1409, N1335, N799, N375, N287);
not NOT1 (N1410, N1407);
nor NOR3 (N1411, N1397, N884, N795);
or OR3 (N1412, N1389, N1109, N811);
or OR4 (N1413, N1405, N1259, N488, N351);
nand NAND2 (N1414, N1413, N379);
buf BUF1 (N1415, N1409);
nand NAND4 (N1416, N1403, N481, N518, N1075);
not NOT1 (N1417, N1400);
nor NOR3 (N1418, N1386, N427, N445);
nand NAND4 (N1419, N1414, N1258, N908, N945);
xor XOR2 (N1420, N1419, N1027);
not NOT1 (N1421, N1411);
buf BUF1 (N1422, N1408);
and AND4 (N1423, N1422, N419, N10, N1204);
nor NOR2 (N1424, N1406, N84);
nor NOR2 (N1425, N1412, N246);
and AND4 (N1426, N1423, N742, N1256, N111);
xor XOR2 (N1427, N1425, N405);
nor NOR2 (N1428, N1426, N596);
and AND3 (N1429, N1417, N850, N1350);
nor NOR2 (N1430, N1418, N873);
nor NOR3 (N1431, N1416, N686, N109);
xor XOR2 (N1432, N1429, N624);
nand NAND4 (N1433, N1410, N1382, N504, N401);
nand NAND4 (N1434, N1420, N652, N463, N339);
nor NOR4 (N1435, N1431, N522, N282, N152);
buf BUF1 (N1436, N1427);
buf BUF1 (N1437, N1435);
xor XOR2 (N1438, N1424, N870);
and AND2 (N1439, N1437, N199);
not NOT1 (N1440, N1439);
nor NOR2 (N1441, N1428, N441);
nor NOR2 (N1442, N1421, N1159);
or OR3 (N1443, N1441, N268, N1116);
nor NOR4 (N1444, N1415, N1192, N408, N678);
nor NOR3 (N1445, N1433, N621, N1300);
nand NAND3 (N1446, N1440, N400, N457);
nand NAND3 (N1447, N1443, N1072, N48);
and AND4 (N1448, N1432, N1228, N446, N635);
or OR4 (N1449, N1430, N140, N492, N755);
nor NOR2 (N1450, N1444, N902);
not NOT1 (N1451, N1438);
nor NOR2 (N1452, N1451, N1266);
nand NAND2 (N1453, N1450, N576);
and AND2 (N1454, N1453, N609);
not NOT1 (N1455, N1446);
xor XOR2 (N1456, N1454, N1345);
and AND4 (N1457, N1456, N182, N287, N1210);
nor NOR4 (N1458, N1448, N253, N368, N708);
nor NOR2 (N1459, N1458, N213);
buf BUF1 (N1460, N1449);
buf BUF1 (N1461, N1442);
buf BUF1 (N1462, N1445);
xor XOR2 (N1463, N1447, N749);
and AND3 (N1464, N1455, N465, N316);
or OR2 (N1465, N1457, N593);
and AND3 (N1466, N1461, N1460, N454);
nor NOR3 (N1467, N1461, N495, N966);
xor XOR2 (N1468, N1463, N1332);
nand NAND2 (N1469, N1462, N753);
not NOT1 (N1470, N1436);
nand NAND2 (N1471, N1452, N718);
and AND3 (N1472, N1434, N7, N1194);
nor NOR4 (N1473, N1471, N727, N567, N1469);
and AND3 (N1474, N979, N812, N655);
or OR3 (N1475, N1470, N268, N651);
xor XOR2 (N1476, N1464, N101);
not NOT1 (N1477, N1468);
not NOT1 (N1478, N1459);
nor NOR4 (N1479, N1476, N127, N63, N765);
xor XOR2 (N1480, N1466, N876);
and AND3 (N1481, N1474, N802, N4);
buf BUF1 (N1482, N1465);
not NOT1 (N1483, N1479);
and AND3 (N1484, N1477, N304, N316);
or OR2 (N1485, N1472, N1312);
nor NOR2 (N1486, N1467, N1195);
xor XOR2 (N1487, N1473, N106);
nand NAND3 (N1488, N1482, N103, N735);
buf BUF1 (N1489, N1483);
buf BUF1 (N1490, N1487);
nor NOR3 (N1491, N1488, N767, N801);
or OR2 (N1492, N1489, N239);
xor XOR2 (N1493, N1492, N834);
buf BUF1 (N1494, N1475);
and AND2 (N1495, N1484, N53);
not NOT1 (N1496, N1493);
and AND2 (N1497, N1486, N833);
or OR4 (N1498, N1494, N470, N921, N72);
and AND4 (N1499, N1485, N201, N1323, N298);
buf BUF1 (N1500, N1478);
nand NAND2 (N1501, N1481, N340);
buf BUF1 (N1502, N1500);
or OR3 (N1503, N1496, N1377, N95);
xor XOR2 (N1504, N1491, N2);
not NOT1 (N1505, N1502);
nor NOR2 (N1506, N1503, N356);
nor NOR4 (N1507, N1501, N566, N1463, N710);
xor XOR2 (N1508, N1505, N934);
or OR2 (N1509, N1480, N789);
nor NOR3 (N1510, N1495, N1300, N1479);
not NOT1 (N1511, N1498);
nand NAND3 (N1512, N1508, N914, N79);
nand NAND4 (N1513, N1506, N883, N262, N440);
not NOT1 (N1514, N1504);
not NOT1 (N1515, N1514);
buf BUF1 (N1516, N1513);
not NOT1 (N1517, N1507);
and AND4 (N1518, N1509, N1334, N1031, N1395);
not NOT1 (N1519, N1516);
not NOT1 (N1520, N1519);
not NOT1 (N1521, N1511);
or OR4 (N1522, N1490, N1434, N646, N1439);
and AND2 (N1523, N1518, N1497);
buf BUF1 (N1524, N450);
not NOT1 (N1525, N1510);
and AND2 (N1526, N1521, N1167);
and AND3 (N1527, N1522, N1340, N1269);
or OR4 (N1528, N1525, N16, N756, N162);
buf BUF1 (N1529, N1499);
nor NOR3 (N1530, N1524, N1167, N283);
xor XOR2 (N1531, N1515, N1442);
nor NOR4 (N1532, N1528, N1064, N1483, N465);
buf BUF1 (N1533, N1527);
xor XOR2 (N1534, N1512, N554);
or OR3 (N1535, N1529, N1335, N980);
not NOT1 (N1536, N1532);
and AND4 (N1537, N1535, N735, N483, N921);
or OR2 (N1538, N1526, N1014);
or OR4 (N1539, N1530, N743, N1066, N723);
not NOT1 (N1540, N1520);
and AND2 (N1541, N1531, N1121);
nor NOR2 (N1542, N1540, N282);
xor XOR2 (N1543, N1517, N1448);
nand NAND2 (N1544, N1543, N686);
or OR4 (N1545, N1537, N348, N1121, N978);
xor XOR2 (N1546, N1538, N1039);
buf BUF1 (N1547, N1536);
and AND3 (N1548, N1523, N252, N1374);
nand NAND2 (N1549, N1541, N1499);
nor NOR2 (N1550, N1547, N1232);
not NOT1 (N1551, N1544);
xor XOR2 (N1552, N1546, N166);
xor XOR2 (N1553, N1551, N1523);
nor NOR4 (N1554, N1549, N1038, N986, N1524);
or OR2 (N1555, N1554, N1276);
and AND4 (N1556, N1552, N1156, N883, N1255);
xor XOR2 (N1557, N1556, N854);
and AND4 (N1558, N1550, N955, N722, N1234);
buf BUF1 (N1559, N1542);
or OR2 (N1560, N1559, N460);
buf BUF1 (N1561, N1539);
not NOT1 (N1562, N1558);
nor NOR2 (N1563, N1561, N1072);
not NOT1 (N1564, N1548);
nor NOR4 (N1565, N1563, N1514, N630, N531);
nor NOR2 (N1566, N1533, N839);
not NOT1 (N1567, N1564);
buf BUF1 (N1568, N1557);
xor XOR2 (N1569, N1568, N112);
and AND3 (N1570, N1567, N389, N319);
nand NAND3 (N1571, N1545, N320, N303);
or OR2 (N1572, N1534, N430);
xor XOR2 (N1573, N1553, N11);
not NOT1 (N1574, N1555);
nand NAND4 (N1575, N1574, N1388, N722, N504);
nor NOR3 (N1576, N1573, N418, N444);
or OR3 (N1577, N1566, N16, N114);
nor NOR3 (N1578, N1562, N653, N973);
nor NOR4 (N1579, N1560, N900, N717, N177);
or OR4 (N1580, N1572, N1115, N667, N1178);
buf BUF1 (N1581, N1580);
buf BUF1 (N1582, N1579);
nand NAND2 (N1583, N1565, N769);
nand NAND3 (N1584, N1570, N318, N921);
nor NOR2 (N1585, N1569, N1264);
xor XOR2 (N1586, N1584, N489);
and AND4 (N1587, N1577, N1498, N1409, N1332);
xor XOR2 (N1588, N1583, N1505);
nand NAND4 (N1589, N1587, N190, N52, N1276);
xor XOR2 (N1590, N1578, N597);
nor NOR3 (N1591, N1575, N1223, N1087);
not NOT1 (N1592, N1590);
nand NAND4 (N1593, N1591, N1570, N1258, N626);
and AND2 (N1594, N1582, N284);
buf BUF1 (N1595, N1581);
and AND3 (N1596, N1594, N1016, N297);
nor NOR4 (N1597, N1592, N353, N919, N980);
nor NOR4 (N1598, N1588, N217, N921, N653);
not NOT1 (N1599, N1593);
not NOT1 (N1600, N1585);
not NOT1 (N1601, N1596);
or OR2 (N1602, N1601, N715);
nand NAND4 (N1603, N1576, N233, N1269, N454);
or OR3 (N1604, N1595, N1083, N774);
and AND2 (N1605, N1597, N182);
xor XOR2 (N1606, N1599, N1143);
nand NAND3 (N1607, N1600, N652, N576);
buf BUF1 (N1608, N1604);
nor NOR4 (N1609, N1603, N57, N1015, N485);
not NOT1 (N1610, N1608);
nor NOR4 (N1611, N1586, N173, N432, N120);
nor NOR4 (N1612, N1605, N1328, N1422, N422);
and AND4 (N1613, N1610, N836, N324, N583);
nand NAND2 (N1614, N1612, N53);
buf BUF1 (N1615, N1609);
buf BUF1 (N1616, N1615);
nor NOR4 (N1617, N1611, N1430, N1466, N1167);
xor XOR2 (N1618, N1614, N954);
xor XOR2 (N1619, N1607, N1529);
nor NOR3 (N1620, N1571, N1311, N944);
buf BUF1 (N1621, N1602);
xor XOR2 (N1622, N1616, N264);
buf BUF1 (N1623, N1622);
not NOT1 (N1624, N1617);
buf BUF1 (N1625, N1613);
nand NAND2 (N1626, N1598, N1485);
and AND4 (N1627, N1626, N894, N1141, N930);
and AND2 (N1628, N1627, N111);
nor NOR2 (N1629, N1625, N894);
nand NAND3 (N1630, N1620, N741, N890);
xor XOR2 (N1631, N1623, N1011);
not NOT1 (N1632, N1629);
nand NAND4 (N1633, N1632, N1612, N1123, N1139);
or OR3 (N1634, N1633, N1508, N810);
buf BUF1 (N1635, N1618);
xor XOR2 (N1636, N1619, N877);
not NOT1 (N1637, N1630);
xor XOR2 (N1638, N1606, N98);
buf BUF1 (N1639, N1636);
xor XOR2 (N1640, N1638, N1603);
or OR3 (N1641, N1589, N167, N652);
xor XOR2 (N1642, N1628, N1548);
or OR2 (N1643, N1641, N1396);
buf BUF1 (N1644, N1635);
nand NAND4 (N1645, N1640, N1547, N577, N322);
nand NAND2 (N1646, N1639, N583);
nor NOR3 (N1647, N1646, N1290, N279);
nand NAND3 (N1648, N1634, N551, N694);
xor XOR2 (N1649, N1637, N591);
not NOT1 (N1650, N1649);
buf BUF1 (N1651, N1631);
not NOT1 (N1652, N1647);
not NOT1 (N1653, N1624);
nand NAND2 (N1654, N1652, N1598);
and AND4 (N1655, N1643, N575, N250, N696);
nor NOR3 (N1656, N1653, N1055, N1483);
buf BUF1 (N1657, N1642);
and AND4 (N1658, N1621, N1093, N568, N332);
or OR4 (N1659, N1645, N373, N10, N1386);
or OR2 (N1660, N1650, N910);
xor XOR2 (N1661, N1656, N815);
nand NAND2 (N1662, N1654, N1452);
buf BUF1 (N1663, N1648);
and AND3 (N1664, N1651, N1138, N1169);
xor XOR2 (N1665, N1664, N27);
nand NAND3 (N1666, N1655, N662, N6);
xor XOR2 (N1667, N1659, N1437);
nand NAND3 (N1668, N1644, N450, N500);
nand NAND2 (N1669, N1663, N882);
buf BUF1 (N1670, N1660);
and AND3 (N1671, N1657, N107, N227);
xor XOR2 (N1672, N1669, N980);
buf BUF1 (N1673, N1671);
and AND3 (N1674, N1672, N1320, N1124);
nand NAND3 (N1675, N1661, N1107, N1410);
buf BUF1 (N1676, N1658);
not NOT1 (N1677, N1675);
nor NOR4 (N1678, N1667, N1615, N1366, N288);
nand NAND2 (N1679, N1674, N596);
not NOT1 (N1680, N1662);
buf BUF1 (N1681, N1677);
nor NOR2 (N1682, N1680, N447);
not NOT1 (N1683, N1679);
nand NAND3 (N1684, N1676, N1047, N386);
buf BUF1 (N1685, N1683);
and AND3 (N1686, N1682, N1096, N1268);
buf BUF1 (N1687, N1668);
nor NOR2 (N1688, N1687, N8);
not NOT1 (N1689, N1684);
buf BUF1 (N1690, N1666);
not NOT1 (N1691, N1670);
not NOT1 (N1692, N1685);
nor NOR4 (N1693, N1690, N1598, N740, N1273);
xor XOR2 (N1694, N1665, N1045);
nand NAND2 (N1695, N1694, N1637);
and AND2 (N1696, N1692, N1450);
xor XOR2 (N1697, N1673, N941);
nand NAND3 (N1698, N1688, N446, N150);
and AND3 (N1699, N1689, N1211, N466);
or OR4 (N1700, N1698, N1194, N977, N1061);
nor NOR2 (N1701, N1681, N499);
or OR3 (N1702, N1699, N1511, N324);
or OR2 (N1703, N1697, N1089);
xor XOR2 (N1704, N1701, N760);
nor NOR4 (N1705, N1691, N203, N563, N991);
buf BUF1 (N1706, N1702);
and AND3 (N1707, N1678, N992, N930);
not NOT1 (N1708, N1686);
not NOT1 (N1709, N1693);
and AND2 (N1710, N1705, N274);
and AND4 (N1711, N1703, N756, N400, N1458);
buf BUF1 (N1712, N1711);
nor NOR2 (N1713, N1707, N260);
and AND2 (N1714, N1700, N924);
nor NOR2 (N1715, N1695, N744);
nand NAND3 (N1716, N1710, N671, N1216);
and AND3 (N1717, N1708, N647, N93);
buf BUF1 (N1718, N1706);
not NOT1 (N1719, N1718);
nor NOR3 (N1720, N1714, N801, N1421);
buf BUF1 (N1721, N1719);
and AND2 (N1722, N1704, N1590);
nand NAND2 (N1723, N1713, N9);
not NOT1 (N1724, N1720);
or OR3 (N1725, N1709, N1468, N634);
nor NOR3 (N1726, N1721, N1716, N1695);
xor XOR2 (N1727, N954, N1664);
xor XOR2 (N1728, N1725, N226);
xor XOR2 (N1729, N1712, N968);
buf BUF1 (N1730, N1723);
or OR4 (N1731, N1730, N1638, N1559, N1204);
and AND4 (N1732, N1696, N967, N582, N972);
and AND2 (N1733, N1729, N1700);
xor XOR2 (N1734, N1726, N477);
and AND4 (N1735, N1724, N716, N194, N1318);
or OR2 (N1736, N1733, N553);
or OR2 (N1737, N1722, N1178);
and AND2 (N1738, N1717, N495);
nand NAND2 (N1739, N1727, N1643);
nand NAND4 (N1740, N1734, N730, N1401, N1098);
or OR4 (N1741, N1715, N1022, N1546, N1099);
xor XOR2 (N1742, N1741, N680);
or OR2 (N1743, N1735, N467);
or OR2 (N1744, N1738, N1735);
nand NAND2 (N1745, N1732, N321);
nor NOR2 (N1746, N1745, N163);
or OR2 (N1747, N1731, N1237);
not NOT1 (N1748, N1746);
nand NAND3 (N1749, N1740, N786, N1015);
xor XOR2 (N1750, N1736, N321);
nand NAND4 (N1751, N1747, N1309, N920, N1266);
buf BUF1 (N1752, N1751);
buf BUF1 (N1753, N1750);
buf BUF1 (N1754, N1728);
nor NOR2 (N1755, N1748, N39);
not NOT1 (N1756, N1739);
and AND2 (N1757, N1744, N516);
or OR4 (N1758, N1755, N756, N131, N939);
nor NOR2 (N1759, N1754, N1438);
nand NAND3 (N1760, N1758, N624, N1340);
buf BUF1 (N1761, N1752);
or OR2 (N1762, N1737, N1005);
xor XOR2 (N1763, N1756, N1687);
xor XOR2 (N1764, N1757, N593);
not NOT1 (N1765, N1743);
xor XOR2 (N1766, N1749, N1223);
nor NOR4 (N1767, N1762, N474, N1636, N567);
and AND2 (N1768, N1753, N1423);
buf BUF1 (N1769, N1765);
and AND2 (N1770, N1768, N1736);
xor XOR2 (N1771, N1767, N504);
or OR2 (N1772, N1763, N1547);
nor NOR2 (N1773, N1766, N267);
xor XOR2 (N1774, N1769, N709);
xor XOR2 (N1775, N1759, N924);
and AND3 (N1776, N1761, N871, N7);
and AND2 (N1777, N1760, N961);
buf BUF1 (N1778, N1764);
and AND4 (N1779, N1776, N865, N1130, N77);
nor NOR2 (N1780, N1775, N347);
xor XOR2 (N1781, N1777, N948);
and AND3 (N1782, N1770, N55, N1156);
xor XOR2 (N1783, N1778, N781);
and AND4 (N1784, N1742, N504, N1726, N1494);
or OR2 (N1785, N1780, N1664);
xor XOR2 (N1786, N1783, N1202);
nand NAND3 (N1787, N1785, N968, N1059);
nor NOR3 (N1788, N1773, N930, N464);
nor NOR3 (N1789, N1772, N1173, N1407);
and AND2 (N1790, N1781, N960);
buf BUF1 (N1791, N1784);
and AND2 (N1792, N1791, N779);
nor NOR3 (N1793, N1771, N185, N795);
nor NOR4 (N1794, N1774, N219, N1436, N628);
or OR3 (N1795, N1793, N1032, N1273);
nor NOR4 (N1796, N1788, N268, N1358, N500);
xor XOR2 (N1797, N1792, N578);
and AND2 (N1798, N1794, N12);
buf BUF1 (N1799, N1796);
nand NAND4 (N1800, N1799, N1753, N362, N54);
and AND3 (N1801, N1789, N1795, N645);
nand NAND4 (N1802, N114, N1105, N992, N1055);
nor NOR2 (N1803, N1798, N124);
or OR4 (N1804, N1787, N341, N1530, N1314);
nand NAND4 (N1805, N1800, N1537, N1552, N863);
buf BUF1 (N1806, N1803);
nor NOR2 (N1807, N1804, N1393);
and AND4 (N1808, N1779, N313, N1689, N521);
nor NOR4 (N1809, N1808, N239, N1523, N1228);
xor XOR2 (N1810, N1809, N1012);
or OR4 (N1811, N1807, N696, N1721, N233);
and AND2 (N1812, N1811, N1331);
and AND2 (N1813, N1810, N161);
buf BUF1 (N1814, N1790);
not NOT1 (N1815, N1814);
or OR2 (N1816, N1813, N220);
buf BUF1 (N1817, N1805);
or OR3 (N1818, N1797, N542, N798);
and AND4 (N1819, N1782, N795, N436, N646);
nor NOR3 (N1820, N1819, N1495, N682);
not NOT1 (N1821, N1802);
or OR3 (N1822, N1815, N1234, N323);
nand NAND2 (N1823, N1816, N1537);
buf BUF1 (N1824, N1817);
nand NAND3 (N1825, N1824, N1637, N1594);
nor NOR4 (N1826, N1823, N1063, N688, N1369);
nor NOR3 (N1827, N1826, N1560, N145);
nor NOR3 (N1828, N1825, N1342, N1068);
nor NOR3 (N1829, N1827, N1145, N1474);
xor XOR2 (N1830, N1821, N625);
not NOT1 (N1831, N1820);
xor XOR2 (N1832, N1812, N641);
not NOT1 (N1833, N1806);
nor NOR3 (N1834, N1828, N910, N1379);
nor NOR2 (N1835, N1832, N1416);
buf BUF1 (N1836, N1833);
not NOT1 (N1837, N1831);
nor NOR3 (N1838, N1829, N1523, N1473);
buf BUF1 (N1839, N1786);
or OR4 (N1840, N1834, N82, N1428, N1589);
or OR2 (N1841, N1822, N1808);
and AND3 (N1842, N1840, N998, N1355);
and AND3 (N1843, N1841, N47, N579);
nand NAND2 (N1844, N1818, N325);
or OR4 (N1845, N1836, N503, N41, N906);
buf BUF1 (N1846, N1830);
or OR4 (N1847, N1842, N1078, N702, N863);
or OR2 (N1848, N1839, N1067);
buf BUF1 (N1849, N1801);
buf BUF1 (N1850, N1843);
xor XOR2 (N1851, N1850, N1367);
or OR3 (N1852, N1835, N635, N151);
nor NOR4 (N1853, N1845, N361, N1175, N1288);
buf BUF1 (N1854, N1837);
xor XOR2 (N1855, N1847, N1709);
buf BUF1 (N1856, N1852);
nand NAND2 (N1857, N1856, N348);
xor XOR2 (N1858, N1849, N674);
not NOT1 (N1859, N1857);
buf BUF1 (N1860, N1854);
buf BUF1 (N1861, N1859);
nor NOR2 (N1862, N1858, N1066);
not NOT1 (N1863, N1861);
not NOT1 (N1864, N1848);
nor NOR2 (N1865, N1864, N1129);
not NOT1 (N1866, N1863);
xor XOR2 (N1867, N1862, N1548);
not NOT1 (N1868, N1844);
or OR4 (N1869, N1860, N929, N515, N1134);
buf BUF1 (N1870, N1868);
buf BUF1 (N1871, N1853);
xor XOR2 (N1872, N1855, N216);
xor XOR2 (N1873, N1867, N1570);
nand NAND2 (N1874, N1871, N34);
nor NOR3 (N1875, N1866, N1279, N6);
nor NOR3 (N1876, N1865, N405, N580);
nand NAND3 (N1877, N1838, N1073, N1519);
not NOT1 (N1878, N1875);
not NOT1 (N1879, N1874);
buf BUF1 (N1880, N1846);
nand NAND2 (N1881, N1879, N583);
nand NAND2 (N1882, N1880, N1449);
not NOT1 (N1883, N1882);
buf BUF1 (N1884, N1873);
or OR4 (N1885, N1869, N1052, N1780, N286);
not NOT1 (N1886, N1883);
buf BUF1 (N1887, N1881);
not NOT1 (N1888, N1870);
nor NOR2 (N1889, N1877, N521);
nor NOR4 (N1890, N1888, N267, N94, N1319);
nand NAND2 (N1891, N1872, N160);
not NOT1 (N1892, N1887);
buf BUF1 (N1893, N1886);
xor XOR2 (N1894, N1889, N1538);
xor XOR2 (N1895, N1891, N1167);
not NOT1 (N1896, N1894);
xor XOR2 (N1897, N1895, N1067);
buf BUF1 (N1898, N1878);
xor XOR2 (N1899, N1876, N794);
nand NAND4 (N1900, N1892, N688, N565, N1615);
nand NAND3 (N1901, N1851, N1665, N213);
or OR4 (N1902, N1899, N1769, N381, N496);
nand NAND2 (N1903, N1901, N543);
or OR4 (N1904, N1885, N1685, N1465, N1717);
not NOT1 (N1905, N1890);
or OR4 (N1906, N1902, N1676, N1503, N1716);
nand NAND2 (N1907, N1896, N1010);
or OR4 (N1908, N1893, N1296, N240, N1258);
and AND3 (N1909, N1884, N1603, N747);
buf BUF1 (N1910, N1903);
not NOT1 (N1911, N1908);
and AND3 (N1912, N1900, N1159, N1749);
nand NAND2 (N1913, N1905, N280);
xor XOR2 (N1914, N1906, N1651);
not NOT1 (N1915, N1898);
not NOT1 (N1916, N1911);
and AND4 (N1917, N1916, N1173, N453, N891);
and AND4 (N1918, N1897, N1269, N1657, N1052);
buf BUF1 (N1919, N1910);
not NOT1 (N1920, N1914);
not NOT1 (N1921, N1918);
not NOT1 (N1922, N1920);
or OR2 (N1923, N1915, N1618);
or OR3 (N1924, N1912, N636, N861);
xor XOR2 (N1925, N1923, N253);
and AND3 (N1926, N1913, N535, N871);
or OR4 (N1927, N1909, N586, N1458, N420);
buf BUF1 (N1928, N1925);
or OR4 (N1929, N1924, N1858, N1277, N660);
buf BUF1 (N1930, N1917);
and AND2 (N1931, N1921, N1598);
and AND4 (N1932, N1929, N1548, N1199, N1874);
or OR4 (N1933, N1922, N410, N1682, N162);
xor XOR2 (N1934, N1926, N887);
nor NOR2 (N1935, N1904, N1207);
not NOT1 (N1936, N1927);
not NOT1 (N1937, N1936);
xor XOR2 (N1938, N1934, N1806);
xor XOR2 (N1939, N1930, N572);
not NOT1 (N1940, N1928);
xor XOR2 (N1941, N1938, N1607);
nand NAND3 (N1942, N1935, N1090, N504);
nor NOR3 (N1943, N1940, N1322, N464);
xor XOR2 (N1944, N1907, N1674);
not NOT1 (N1945, N1933);
nor NOR3 (N1946, N1944, N1605, N1631);
xor XOR2 (N1947, N1932, N1148);
or OR4 (N1948, N1945, N1138, N1523, N122);
nand NAND4 (N1949, N1948, N397, N245, N82);
or OR2 (N1950, N1931, N280);
buf BUF1 (N1951, N1937);
or OR4 (N1952, N1950, N1747, N1452, N1180);
and AND2 (N1953, N1946, N1394);
nand NAND3 (N1954, N1939, N972, N1659);
and AND3 (N1955, N1943, N861, N1634);
not NOT1 (N1956, N1953);
buf BUF1 (N1957, N1954);
not NOT1 (N1958, N1951);
nand NAND2 (N1959, N1949, N1622);
nor NOR4 (N1960, N1941, N1057, N1883, N1669);
not NOT1 (N1961, N1960);
xor XOR2 (N1962, N1961, N978);
not NOT1 (N1963, N1955);
xor XOR2 (N1964, N1952, N1504);
buf BUF1 (N1965, N1956);
buf BUF1 (N1966, N1958);
nand NAND2 (N1967, N1963, N380);
not NOT1 (N1968, N1957);
xor XOR2 (N1969, N1967, N1605);
nand NAND4 (N1970, N1942, N396, N1863, N972);
or OR3 (N1971, N1968, N262, N1465);
xor XOR2 (N1972, N1966, N678);
buf BUF1 (N1973, N1947);
xor XOR2 (N1974, N1962, N1789);
not NOT1 (N1975, N1959);
xor XOR2 (N1976, N1974, N1821);
and AND3 (N1977, N1971, N214, N503);
not NOT1 (N1978, N1970);
and AND3 (N1979, N1969, N800, N1849);
nor NOR2 (N1980, N1975, N869);
xor XOR2 (N1981, N1964, N1637);
and AND4 (N1982, N1976, N1707, N1159, N501);
not NOT1 (N1983, N1982);
nand NAND4 (N1984, N1965, N905, N1333, N1829);
xor XOR2 (N1985, N1972, N625);
nor NOR4 (N1986, N1978, N1864, N704, N562);
nand NAND2 (N1987, N1984, N198);
buf BUF1 (N1988, N1979);
buf BUF1 (N1989, N1987);
and AND3 (N1990, N1988, N765, N202);
buf BUF1 (N1991, N1990);
nor NOR4 (N1992, N1989, N732, N264, N1786);
buf BUF1 (N1993, N1985);
or OR3 (N1994, N1992, N348, N172);
nand NAND3 (N1995, N1991, N12, N1337);
or OR4 (N1996, N1980, N1312, N1987, N1762);
buf BUF1 (N1997, N1986);
nor NOR4 (N1998, N1973, N1186, N1783, N747);
and AND4 (N1999, N1919, N1901, N586, N531);
xor XOR2 (N2000, N1998, N916);
not NOT1 (N2001, N1993);
not NOT1 (N2002, N2000);
nor NOR2 (N2003, N2002, N20);
xor XOR2 (N2004, N1994, N1898);
nor NOR3 (N2005, N2001, N1856, N163);
buf BUF1 (N2006, N1983);
not NOT1 (N2007, N1981);
and AND2 (N2008, N1999, N205);
xor XOR2 (N2009, N2007, N175);
not NOT1 (N2010, N2008);
nand NAND3 (N2011, N2009, N1463, N154);
and AND4 (N2012, N2010, N752, N1990, N1914);
and AND3 (N2013, N1977, N1139, N733);
xor XOR2 (N2014, N2006, N695);
and AND3 (N2015, N2014, N865, N418);
and AND2 (N2016, N1996, N373);
or OR3 (N2017, N2013, N1623, N72);
xor XOR2 (N2018, N2012, N1614);
buf BUF1 (N2019, N2017);
not NOT1 (N2020, N2011);
xor XOR2 (N2021, N1995, N497);
and AND4 (N2022, N2016, N551, N1961, N864);
xor XOR2 (N2023, N2003, N696);
buf BUF1 (N2024, N2005);
nand NAND4 (N2025, N2024, N1323, N1233, N1875);
or OR2 (N2026, N2023, N1583);
buf BUF1 (N2027, N1997);
not NOT1 (N2028, N2018);
nand NAND3 (N2029, N2028, N1773, N1365);
not NOT1 (N2030, N2021);
nand NAND2 (N2031, N2029, N1879);
not NOT1 (N2032, N2019);
or OR3 (N2033, N2020, N1662, N1975);
xor XOR2 (N2034, N2015, N1168);
nand NAND4 (N2035, N2030, N538, N895, N1751);
and AND2 (N2036, N2034, N902);
nor NOR4 (N2037, N2035, N584, N829, N657);
xor XOR2 (N2038, N2025, N193);
and AND3 (N2039, N2036, N1706, N708);
nor NOR2 (N2040, N2038, N496);
not NOT1 (N2041, N2037);
not NOT1 (N2042, N2041);
nor NOR3 (N2043, N2039, N543, N142);
xor XOR2 (N2044, N2031, N691);
nand NAND3 (N2045, N2032, N119, N1214);
nor NOR3 (N2046, N2044, N1819, N447);
or OR4 (N2047, N2040, N1338, N1619, N1449);
not NOT1 (N2048, N2033);
nand NAND2 (N2049, N2046, N616);
not NOT1 (N2050, N2026);
or OR4 (N2051, N2042, N536, N656, N1318);
nand NAND4 (N2052, N2022, N1960, N1284, N1824);
or OR3 (N2053, N2051, N297, N888);
buf BUF1 (N2054, N2004);
or OR3 (N2055, N2052, N1079, N1359);
or OR4 (N2056, N2047, N1693, N1418, N1772);
xor XOR2 (N2057, N2056, N976);
xor XOR2 (N2058, N2043, N1337);
buf BUF1 (N2059, N2053);
nor NOR2 (N2060, N2058, N918);
nand NAND4 (N2061, N2027, N620, N563, N735);
not NOT1 (N2062, N2057);
nand NAND2 (N2063, N2055, N1921);
and AND4 (N2064, N2062, N811, N670, N1995);
nor NOR4 (N2065, N2049, N128, N1502, N1882);
xor XOR2 (N2066, N2061, N65);
nand NAND2 (N2067, N2064, N781);
nor NOR3 (N2068, N2059, N1367, N21);
xor XOR2 (N2069, N2067, N1235);
not NOT1 (N2070, N2069);
and AND3 (N2071, N2068, N952, N1973);
or OR2 (N2072, N2054, N1325);
or OR3 (N2073, N2048, N200, N1956);
and AND4 (N2074, N2065, N1257, N651, N1919);
not NOT1 (N2075, N2066);
not NOT1 (N2076, N2045);
not NOT1 (N2077, N2050);
buf BUF1 (N2078, N2076);
xor XOR2 (N2079, N2078, N1044);
not NOT1 (N2080, N2074);
buf BUF1 (N2081, N2072);
buf BUF1 (N2082, N2071);
and AND2 (N2083, N2073, N871);
nor NOR4 (N2084, N2082, N1532, N2034, N1184);
buf BUF1 (N2085, N2084);
nand NAND3 (N2086, N2080, N73, N1477);
nand NAND4 (N2087, N2075, N1354, N1861, N43);
not NOT1 (N2088, N2085);
or OR2 (N2089, N2070, N299);
xor XOR2 (N2090, N2060, N636);
nor NOR3 (N2091, N2081, N1064, N1068);
nor NOR4 (N2092, N2083, N1705, N684, N918);
buf BUF1 (N2093, N2089);
nand NAND2 (N2094, N2092, N301);
xor XOR2 (N2095, N2091, N1076);
or OR4 (N2096, N2077, N1559, N1779, N586);
nand NAND2 (N2097, N2087, N787);
not NOT1 (N2098, N2090);
not NOT1 (N2099, N2086);
nand NAND3 (N2100, N2063, N345, N881);
or OR3 (N2101, N2096, N1691, N1996);
not NOT1 (N2102, N2095);
nand NAND4 (N2103, N2088, N132, N1049, N429);
not NOT1 (N2104, N2097);
nor NOR4 (N2105, N2093, N6, N1108, N716);
not NOT1 (N2106, N2105);
nand NAND4 (N2107, N2079, N1086, N276, N800);
buf BUF1 (N2108, N2107);
and AND3 (N2109, N2101, N365, N1396);
buf BUF1 (N2110, N2094);
nor NOR2 (N2111, N2103, N2027);
and AND3 (N2112, N2109, N1994, N1255);
not NOT1 (N2113, N2112);
buf BUF1 (N2114, N2098);
not NOT1 (N2115, N2111);
nand NAND3 (N2116, N2102, N2012, N1820);
nand NAND2 (N2117, N2108, N804);
nor NOR3 (N2118, N2110, N934, N171);
and AND3 (N2119, N2099, N395, N845);
xor XOR2 (N2120, N2100, N1244);
or OR3 (N2121, N2117, N1997, N117);
and AND2 (N2122, N2106, N1475);
xor XOR2 (N2123, N2104, N1311);
xor XOR2 (N2124, N2120, N1425);
buf BUF1 (N2125, N2124);
or OR3 (N2126, N2114, N1860, N1002);
or OR3 (N2127, N2115, N1086, N144);
or OR4 (N2128, N2119, N791, N457, N1930);
buf BUF1 (N2129, N2116);
xor XOR2 (N2130, N2127, N483);
or OR3 (N2131, N2126, N506, N904);
or OR2 (N2132, N2125, N1916);
not NOT1 (N2133, N2122);
not NOT1 (N2134, N2123);
and AND2 (N2135, N2132, N608);
xor XOR2 (N2136, N2129, N1171);
or OR2 (N2137, N2135, N1949);
not NOT1 (N2138, N2134);
nor NOR2 (N2139, N2131, N591);
nor NOR3 (N2140, N2113, N1916, N1667);
or OR4 (N2141, N2118, N942, N1524, N237);
nand NAND3 (N2142, N2130, N389, N1348);
nor NOR2 (N2143, N2136, N1733);
xor XOR2 (N2144, N2137, N1220);
nand NAND2 (N2145, N2133, N2013);
or OR3 (N2146, N2143, N277, N1677);
or OR4 (N2147, N2128, N1384, N1918, N1650);
not NOT1 (N2148, N2141);
nand NAND3 (N2149, N2138, N1010, N1681);
and AND2 (N2150, N2145, N1905);
xor XOR2 (N2151, N2146, N1662);
xor XOR2 (N2152, N2149, N1159);
nand NAND2 (N2153, N2142, N1901);
and AND2 (N2154, N2150, N1612);
and AND2 (N2155, N2139, N1970);
nor NOR4 (N2156, N2153, N1567, N2090, N160);
nand NAND4 (N2157, N2155, N2153, N2073, N1593);
and AND4 (N2158, N2156, N849, N1796, N1458);
nor NOR2 (N2159, N2147, N1662);
nor NOR2 (N2160, N2148, N351);
or OR3 (N2161, N2154, N697, N1581);
nand NAND2 (N2162, N2158, N1506);
nand NAND3 (N2163, N2151, N637, N1845);
not NOT1 (N2164, N2144);
and AND4 (N2165, N2160, N1876, N1661, N185);
not NOT1 (N2166, N2164);
and AND4 (N2167, N2157, N686, N1156, N167);
nand NAND2 (N2168, N2140, N159);
not NOT1 (N2169, N2167);
not NOT1 (N2170, N2161);
not NOT1 (N2171, N2152);
buf BUF1 (N2172, N2165);
and AND3 (N2173, N2159, N1833, N1233);
or OR3 (N2174, N2163, N129, N1644);
nand NAND2 (N2175, N2171, N1239);
or OR2 (N2176, N2166, N608);
not NOT1 (N2177, N2162);
and AND4 (N2178, N2170, N465, N1792, N1877);
and AND4 (N2179, N2177, N1792, N50, N1178);
buf BUF1 (N2180, N2172);
not NOT1 (N2181, N2180);
xor XOR2 (N2182, N2181, N113);
xor XOR2 (N2183, N2178, N1112);
not NOT1 (N2184, N2182);
xor XOR2 (N2185, N2183, N1206);
not NOT1 (N2186, N2168);
nand NAND4 (N2187, N2173, N1136, N1352, N793);
nor NOR2 (N2188, N2179, N1684);
or OR2 (N2189, N2176, N856);
xor XOR2 (N2190, N2184, N1301);
nor NOR2 (N2191, N2175, N1687);
or OR2 (N2192, N2190, N1193);
xor XOR2 (N2193, N2192, N353);
nor NOR3 (N2194, N2174, N2131, N1527);
nand NAND3 (N2195, N2187, N1431, N82);
nand NAND4 (N2196, N2185, N1774, N29, N120);
nand NAND3 (N2197, N2186, N1484, N1201);
not NOT1 (N2198, N2196);
or OR2 (N2199, N2188, N868);
or OR4 (N2200, N2121, N192, N445, N911);
and AND4 (N2201, N2197, N1172, N383, N1042);
xor XOR2 (N2202, N2169, N928);
nand NAND2 (N2203, N2191, N522);
nor NOR4 (N2204, N2201, N664, N494, N1662);
not NOT1 (N2205, N2189);
not NOT1 (N2206, N2198);
not NOT1 (N2207, N2202);
and AND3 (N2208, N2200, N914, N1262);
nor NOR4 (N2209, N2206, N1212, N742, N888);
or OR2 (N2210, N2194, N1561);
xor XOR2 (N2211, N2207, N1454);
and AND3 (N2212, N2211, N129, N1456);
and AND4 (N2213, N2205, N2204, N2010, N1922);
nand NAND3 (N2214, N2024, N1236, N2007);
and AND4 (N2215, N2212, N1362, N486, N1223);
xor XOR2 (N2216, N2210, N1931);
buf BUF1 (N2217, N2215);
and AND2 (N2218, N2195, N901);
buf BUF1 (N2219, N2218);
buf BUF1 (N2220, N2213);
buf BUF1 (N2221, N2199);
xor XOR2 (N2222, N2214, N64);
and AND4 (N2223, N2209, N1378, N541, N1615);
and AND3 (N2224, N2221, N1941, N1138);
or OR4 (N2225, N2208, N338, N619, N1257);
not NOT1 (N2226, N2223);
buf BUF1 (N2227, N2224);
or OR4 (N2228, N2219, N505, N1695, N1414);
not NOT1 (N2229, N2228);
and AND2 (N2230, N2217, N527);
and AND3 (N2231, N2227, N1702, N22);
or OR2 (N2232, N2226, N1122);
nand NAND2 (N2233, N2231, N1930);
xor XOR2 (N2234, N2220, N456);
not NOT1 (N2235, N2229);
nor NOR3 (N2236, N2222, N812, N679);
nand NAND2 (N2237, N2193, N942);
xor XOR2 (N2238, N2234, N398);
nand NAND3 (N2239, N2232, N1309, N902);
and AND4 (N2240, N2230, N446, N96, N1080);
and AND2 (N2241, N2240, N1821);
buf BUF1 (N2242, N2236);
nor NOR2 (N2243, N2241, N1325);
xor XOR2 (N2244, N2235, N1222);
xor XOR2 (N2245, N2225, N1553);
not NOT1 (N2246, N2245);
nor NOR3 (N2247, N2239, N886, N695);
nand NAND2 (N2248, N2237, N1811);
not NOT1 (N2249, N2238);
and AND4 (N2250, N2216, N1083, N1402, N1083);
and AND2 (N2251, N2243, N537);
or OR2 (N2252, N2249, N2054);
nor NOR4 (N2253, N2244, N300, N551, N861);
or OR2 (N2254, N2248, N118);
nand NAND2 (N2255, N2252, N2176);
or OR3 (N2256, N2255, N1519, N1915);
not NOT1 (N2257, N2256);
nand NAND3 (N2258, N2257, N1025, N1972);
nand NAND3 (N2259, N2242, N590, N1065);
not NOT1 (N2260, N2259);
not NOT1 (N2261, N2258);
nand NAND3 (N2262, N2247, N635, N655);
nand NAND4 (N2263, N2254, N2223, N1570, N1547);
not NOT1 (N2264, N2251);
or OR3 (N2265, N2260, N1808, N199);
not NOT1 (N2266, N2253);
not NOT1 (N2267, N2264);
nand NAND3 (N2268, N2265, N1404, N534);
and AND4 (N2269, N2268, N464, N1649, N1464);
xor XOR2 (N2270, N2267, N59);
nand NAND4 (N2271, N2263, N21, N789, N1429);
nand NAND2 (N2272, N2269, N2259);
nand NAND2 (N2273, N2262, N1966);
buf BUF1 (N2274, N2266);
nor NOR4 (N2275, N2233, N854, N1387, N1688);
not NOT1 (N2276, N2273);
nand NAND3 (N2277, N2276, N452, N1515);
buf BUF1 (N2278, N2277);
and AND4 (N2279, N2272, N1372, N1367, N681);
not NOT1 (N2280, N2261);
or OR2 (N2281, N2279, N27);
nor NOR3 (N2282, N2246, N756, N53);
nand NAND2 (N2283, N2281, N378);
buf BUF1 (N2284, N2270);
nand NAND3 (N2285, N2282, N2001, N501);
nand NAND3 (N2286, N2250, N636, N192);
buf BUF1 (N2287, N2278);
buf BUF1 (N2288, N2287);
buf BUF1 (N2289, N2280);
nand NAND2 (N2290, N2275, N196);
xor XOR2 (N2291, N2203, N1856);
not NOT1 (N2292, N2286);
nand NAND3 (N2293, N2290, N973, N458);
and AND2 (N2294, N2288, N456);
or OR3 (N2295, N2285, N330, N376);
nand NAND4 (N2296, N2294, N2092, N913, N2145);
buf BUF1 (N2297, N2291);
not NOT1 (N2298, N2283);
buf BUF1 (N2299, N2295);
and AND4 (N2300, N2292, N879, N71, N711);
and AND4 (N2301, N2284, N389, N690, N408);
xor XOR2 (N2302, N2274, N1294);
or OR2 (N2303, N2299, N1018);
buf BUF1 (N2304, N2302);
or OR3 (N2305, N2297, N1914, N1706);
nor NOR4 (N2306, N2305, N671, N397, N2138);
nor NOR4 (N2307, N2303, N1235, N942, N843);
xor XOR2 (N2308, N2306, N1267);
buf BUF1 (N2309, N2304);
xor XOR2 (N2310, N2301, N1021);
nor NOR4 (N2311, N2293, N163, N1299, N1070);
nor NOR4 (N2312, N2311, N86, N1201, N1166);
not NOT1 (N2313, N2271);
xor XOR2 (N2314, N2289, N353);
nand NAND3 (N2315, N2312, N442, N1559);
or OR2 (N2316, N2314, N1871);
or OR2 (N2317, N2300, N2273);
nor NOR2 (N2318, N2315, N2135);
or OR3 (N2319, N2298, N2174, N1976);
nand NAND4 (N2320, N2310, N996, N1084, N2118);
nor NOR3 (N2321, N2318, N49, N691);
nand NAND3 (N2322, N2307, N1560, N2150);
xor XOR2 (N2323, N2313, N2268);
not NOT1 (N2324, N2323);
or OR3 (N2325, N2309, N1865, N468);
nand NAND2 (N2326, N2316, N1030);
not NOT1 (N2327, N2322);
and AND2 (N2328, N2326, N1025);
and AND3 (N2329, N2328, N1000, N596);
nor NOR2 (N2330, N2321, N969);
buf BUF1 (N2331, N2296);
nand NAND2 (N2332, N2324, N1796);
not NOT1 (N2333, N2331);
xor XOR2 (N2334, N2330, N1467);
nor NOR2 (N2335, N2333, N1014);
buf BUF1 (N2336, N2319);
xor XOR2 (N2337, N2325, N1425);
or OR4 (N2338, N2317, N787, N1805, N630);
nand NAND2 (N2339, N2336, N1435);
nor NOR4 (N2340, N2332, N2139, N897, N1380);
xor XOR2 (N2341, N2327, N1691);
nor NOR4 (N2342, N2340, N2128, N41, N1197);
and AND2 (N2343, N2335, N1042);
xor XOR2 (N2344, N2343, N413);
not NOT1 (N2345, N2329);
buf BUF1 (N2346, N2334);
nand NAND2 (N2347, N2320, N182);
or OR2 (N2348, N2308, N1267);
nand NAND2 (N2349, N2337, N1737);
or OR2 (N2350, N2341, N2311);
nand NAND4 (N2351, N2338, N1183, N798, N254);
nor NOR4 (N2352, N2351, N1045, N2206, N419);
xor XOR2 (N2353, N2344, N990);
xor XOR2 (N2354, N2348, N874);
nand NAND2 (N2355, N2353, N2339);
nand NAND2 (N2356, N921, N2048);
nor NOR3 (N2357, N2345, N417, N217);
or OR2 (N2358, N2349, N723);
nand NAND4 (N2359, N2342, N658, N236, N1371);
buf BUF1 (N2360, N2347);
nand NAND4 (N2361, N2356, N1771, N225, N324);
not NOT1 (N2362, N2354);
not NOT1 (N2363, N2360);
nand NAND4 (N2364, N2361, N1898, N1269, N2059);
nand NAND2 (N2365, N2364, N253);
not NOT1 (N2366, N2362);
not NOT1 (N2367, N2352);
or OR2 (N2368, N2365, N300);
not NOT1 (N2369, N2366);
buf BUF1 (N2370, N2350);
or OR2 (N2371, N2346, N118);
nand NAND2 (N2372, N2359, N1525);
not NOT1 (N2373, N2357);
buf BUF1 (N2374, N2373);
buf BUF1 (N2375, N2371);
nor NOR2 (N2376, N2369, N579);
xor XOR2 (N2377, N2372, N848);
nand NAND2 (N2378, N2374, N1243);
xor XOR2 (N2379, N2378, N1047);
nor NOR3 (N2380, N2379, N1997, N848);
nor NOR4 (N2381, N2375, N46, N1361, N1739);
not NOT1 (N2382, N2380);
nand NAND2 (N2383, N2358, N240);
or OR2 (N2384, N2363, N321);
or OR4 (N2385, N2381, N2290, N1460, N2238);
buf BUF1 (N2386, N2383);
not NOT1 (N2387, N2377);
and AND2 (N2388, N2367, N47);
xor XOR2 (N2389, N2355, N881);
nor NOR2 (N2390, N2388, N961);
or OR2 (N2391, N2386, N1853);
and AND3 (N2392, N2368, N2156, N584);
nor NOR2 (N2393, N2392, N1627);
and AND3 (N2394, N2387, N478, N1504);
or OR3 (N2395, N2382, N850, N100);
and AND3 (N2396, N2390, N2087, N416);
or OR2 (N2397, N2394, N1264);
nand NAND2 (N2398, N2389, N222);
xor XOR2 (N2399, N2391, N1065);
or OR2 (N2400, N2370, N2351);
buf BUF1 (N2401, N2385);
not NOT1 (N2402, N2400);
or OR2 (N2403, N2384, N132);
or OR3 (N2404, N2403, N920, N1741);
or OR3 (N2405, N2397, N2276, N1213);
xor XOR2 (N2406, N2404, N665);
xor XOR2 (N2407, N2406, N122);
buf BUF1 (N2408, N2402);
xor XOR2 (N2409, N2396, N369);
nand NAND2 (N2410, N2405, N285);
nor NOR3 (N2411, N2408, N1893, N482);
nor NOR3 (N2412, N2401, N313, N163);
xor XOR2 (N2413, N2410, N998);
buf BUF1 (N2414, N2409);
not NOT1 (N2415, N2411);
nand NAND4 (N2416, N2412, N16, N1586, N1312);
nand NAND4 (N2417, N2407, N1659, N128, N1081);
and AND4 (N2418, N2417, N85, N1982, N2110);
nor NOR2 (N2419, N2393, N663);
and AND2 (N2420, N2376, N1365);
nor NOR4 (N2421, N2395, N1520, N664, N596);
buf BUF1 (N2422, N2398);
nor NOR4 (N2423, N2419, N1902, N2235, N1577);
nand NAND3 (N2424, N2423, N834, N336);
buf BUF1 (N2425, N2415);
not NOT1 (N2426, N2399);
not NOT1 (N2427, N2421);
nand NAND4 (N2428, N2425, N33, N103, N1702);
nand NAND4 (N2429, N2416, N774, N1623, N1173);
not NOT1 (N2430, N2422);
not NOT1 (N2431, N2429);
or OR4 (N2432, N2427, N1769, N2123, N224);
nor NOR3 (N2433, N2418, N1976, N2104);
nor NOR3 (N2434, N2428, N271, N738);
nor NOR4 (N2435, N2420, N1992, N1543, N2098);
or OR3 (N2436, N2432, N448, N813);
nand NAND4 (N2437, N2430, N1952, N272, N1642);
or OR2 (N2438, N2436, N453);
nor NOR4 (N2439, N2424, N1923, N769, N2115);
or OR3 (N2440, N2439, N918, N139);
or OR3 (N2441, N2434, N608, N124);
buf BUF1 (N2442, N2440);
not NOT1 (N2443, N2435);
not NOT1 (N2444, N2414);
xor XOR2 (N2445, N2433, N1281);
or OR2 (N2446, N2444, N2129);
not NOT1 (N2447, N2438);
buf BUF1 (N2448, N2443);
buf BUF1 (N2449, N2448);
buf BUF1 (N2450, N2449);
not NOT1 (N2451, N2446);
xor XOR2 (N2452, N2437, N2038);
and AND4 (N2453, N2426, N1519, N2209, N2363);
xor XOR2 (N2454, N2450, N1191);
nand NAND2 (N2455, N2451, N137);
not NOT1 (N2456, N2413);
xor XOR2 (N2457, N2441, N646);
nand NAND2 (N2458, N2452, N178);
or OR3 (N2459, N2453, N457, N2287);
nand NAND2 (N2460, N2445, N479);
not NOT1 (N2461, N2442);
not NOT1 (N2462, N2455);
and AND4 (N2463, N2458, N1074, N442, N2174);
not NOT1 (N2464, N2462);
buf BUF1 (N2465, N2464);
nor NOR3 (N2466, N2447, N247, N2128);
xor XOR2 (N2467, N2459, N1392);
and AND4 (N2468, N2465, N2030, N1681, N972);
or OR3 (N2469, N2466, N1867, N1252);
not NOT1 (N2470, N2468);
or OR3 (N2471, N2454, N1484, N2386);
and AND4 (N2472, N2460, N1757, N540, N1979);
xor XOR2 (N2473, N2461, N1042);
not NOT1 (N2474, N2457);
and AND3 (N2475, N2474, N305, N727);
nor NOR3 (N2476, N2475, N1948, N2389);
and AND2 (N2477, N2467, N1813);
or OR3 (N2478, N2473, N2470, N671);
buf BUF1 (N2479, N1146);
or OR3 (N2480, N2479, N1932, N2035);
not NOT1 (N2481, N2469);
or OR4 (N2482, N2472, N797, N2458, N902);
nand NAND3 (N2483, N2431, N226, N1317);
not NOT1 (N2484, N2456);
nor NOR2 (N2485, N2477, N185);
or OR4 (N2486, N2481, N1150, N196, N468);
nor NOR4 (N2487, N2480, N1978, N2472, N1190);
nand NAND2 (N2488, N2486, N1797);
nand NAND3 (N2489, N2488, N333, N2212);
nand NAND4 (N2490, N2487, N257, N1618, N1654);
xor XOR2 (N2491, N2482, N1327);
not NOT1 (N2492, N2489);
xor XOR2 (N2493, N2484, N893);
nor NOR3 (N2494, N2491, N2108, N1731);
or OR4 (N2495, N2476, N358, N2475, N366);
nor NOR3 (N2496, N2483, N2188, N63);
not NOT1 (N2497, N2494);
nand NAND3 (N2498, N2478, N270, N1136);
nor NOR3 (N2499, N2493, N1315, N1187);
or OR3 (N2500, N2496, N965, N546);
nand NAND4 (N2501, N2495, N487, N1427, N1402);
and AND2 (N2502, N2501, N1263);
buf BUF1 (N2503, N2492);
and AND3 (N2504, N2485, N1787, N1205);
not NOT1 (N2505, N2503);
buf BUF1 (N2506, N2490);
nand NAND2 (N2507, N2506, N1700);
and AND2 (N2508, N2463, N1336);
or OR4 (N2509, N2504, N1067, N1586, N277);
buf BUF1 (N2510, N2499);
buf BUF1 (N2511, N2498);
endmodule