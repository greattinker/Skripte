// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17;

output N3506,N3512,N3515,N3516,N3510,N3511,N3513,N3509,N3484,N3517;

buf BUF1 (N18, N10);
and AND3 (N19, N10, N13, N6);
xor XOR2 (N20, N2, N13);
buf BUF1 (N21, N1);
buf BUF1 (N22, N3);
nor NOR4 (N23, N17, N13, N15, N1);
not NOT1 (N24, N14);
nor NOR2 (N25, N9, N9);
or OR4 (N26, N10, N14, N1, N19);
xor XOR2 (N27, N15, N24);
nand NAND2 (N28, N2, N25);
or OR2 (N29, N2, N19);
nand NAND3 (N30, N9, N25, N26);
or OR4 (N31, N5, N12, N13, N11);
not NOT1 (N32, N29);
nor NOR2 (N33, N20, N19);
and AND2 (N34, N33, N12);
buf BUF1 (N35, N32);
nand NAND3 (N36, N31, N28, N18);
not NOT1 (N37, N16);
xor XOR2 (N38, N5, N8);
and AND3 (N39, N37, N30, N32);
and AND3 (N40, N3, N22, N5);
nand NAND2 (N41, N3, N28);
not NOT1 (N42, N34);
nor NOR3 (N43, N41, N28, N30);
nor NOR2 (N44, N27, N39);
buf BUF1 (N45, N19);
nand NAND2 (N46, N21, N25);
nor NOR4 (N47, N45, N31, N8, N17);
buf BUF1 (N48, N44);
nor NOR2 (N49, N43, N47);
not NOT1 (N50, N18);
nor NOR4 (N51, N40, N35, N27, N33);
or OR4 (N52, N34, N21, N13, N19);
and AND2 (N53, N23, N45);
or OR2 (N54, N48, N52);
xor XOR2 (N55, N33, N46);
nand NAND2 (N56, N54, N16);
nor NOR2 (N57, N16, N52);
or OR4 (N58, N49, N53, N48, N46);
xor XOR2 (N59, N12, N22);
or OR4 (N60, N42, N10, N27, N42);
and AND3 (N61, N57, N50, N19);
nand NAND2 (N62, N56, N12);
not NOT1 (N63, N7);
buf BUF1 (N64, N51);
or OR3 (N65, N36, N63, N2);
nor NOR2 (N66, N25, N57);
and AND2 (N67, N61, N23);
or OR2 (N68, N66, N34);
and AND2 (N69, N38, N68);
nor NOR2 (N70, N50, N6);
and AND2 (N71, N62, N11);
nor NOR2 (N72, N69, N33);
or OR3 (N73, N65, N66, N60);
not NOT1 (N74, N68);
or OR4 (N75, N64, N7, N56, N31);
nor NOR2 (N76, N59, N8);
nor NOR3 (N77, N73, N45, N61);
nand NAND2 (N78, N76, N45);
not NOT1 (N79, N77);
not NOT1 (N80, N67);
nand NAND2 (N81, N72, N32);
xor XOR2 (N82, N80, N9);
and AND4 (N83, N82, N14, N41, N55);
nand NAND4 (N84, N65, N4, N3, N74);
or OR3 (N85, N61, N11, N4);
nor NOR2 (N86, N70, N34);
buf BUF1 (N87, N58);
or OR3 (N88, N79, N18, N74);
buf BUF1 (N89, N71);
not NOT1 (N90, N83);
nor NOR2 (N91, N90, N8);
nor NOR4 (N92, N89, N70, N46, N22);
buf BUF1 (N93, N84);
nor NOR4 (N94, N81, N3, N41, N13);
not NOT1 (N95, N75);
nand NAND4 (N96, N78, N47, N32, N62);
buf BUF1 (N97, N85);
not NOT1 (N98, N96);
nor NOR3 (N99, N88, N98, N29);
xor XOR2 (N100, N97, N6);
buf BUF1 (N101, N57);
not NOT1 (N102, N99);
or OR3 (N103, N102, N55, N70);
buf BUF1 (N104, N95);
or OR3 (N105, N104, N34, N5);
or OR2 (N106, N92, N86);
nor NOR4 (N107, N49, N23, N65, N87);
or OR4 (N108, N100, N89, N75, N73);
buf BUF1 (N109, N56);
nand NAND3 (N110, N108, N63, N70);
or OR4 (N111, N109, N110, N54, N41);
xor XOR2 (N112, N11, N99);
and AND4 (N113, N94, N112, N67, N87);
xor XOR2 (N114, N35, N50);
nor NOR4 (N115, N103, N81, N35, N18);
not NOT1 (N116, N93);
buf BUF1 (N117, N115);
nand NAND3 (N118, N114, N67, N39);
not NOT1 (N119, N107);
xor XOR2 (N120, N105, N86);
or OR4 (N121, N91, N119, N78, N62);
or OR2 (N122, N12, N77);
not NOT1 (N123, N121);
nor NOR3 (N124, N123, N111, N84);
or OR3 (N125, N63, N122, N76);
and AND2 (N126, N1, N123);
nand NAND4 (N127, N117, N45, N43, N99);
nor NOR4 (N128, N127, N119, N40, N70);
not NOT1 (N129, N116);
nand NAND4 (N130, N128, N110, N106, N37);
nor NOR4 (N131, N23, N10, N52, N93);
not NOT1 (N132, N130);
and AND4 (N133, N132, N28, N111, N110);
or OR3 (N134, N113, N119, N17);
nand NAND4 (N135, N101, N83, N53, N42);
buf BUF1 (N136, N124);
not NOT1 (N137, N135);
or OR4 (N138, N134, N17, N127, N122);
and AND3 (N139, N129, N66, N92);
buf BUF1 (N140, N133);
nor NOR4 (N141, N137, N9, N78, N6);
xor XOR2 (N142, N138, N92);
or OR3 (N143, N131, N105, N133);
not NOT1 (N144, N120);
nand NAND3 (N145, N141, N86, N90);
nand NAND2 (N146, N126, N102);
not NOT1 (N147, N139);
xor XOR2 (N148, N144, N56);
or OR4 (N149, N148, N78, N49, N34);
and AND2 (N150, N147, N75);
not NOT1 (N151, N125);
xor XOR2 (N152, N146, N46);
and AND2 (N153, N151, N152);
xor XOR2 (N154, N145, N57);
xor XOR2 (N155, N86, N56);
buf BUF1 (N156, N118);
nor NOR2 (N157, N140, N132);
xor XOR2 (N158, N143, N157);
nor NOR3 (N159, N81, N49, N29);
nor NOR2 (N160, N149, N125);
nor NOR4 (N161, N160, N93, N34, N140);
xor XOR2 (N162, N158, N17);
buf BUF1 (N163, N161);
buf BUF1 (N164, N162);
buf BUF1 (N165, N159);
nor NOR2 (N166, N142, N27);
and AND3 (N167, N163, N114, N15);
or OR2 (N168, N167, N126);
and AND3 (N169, N153, N52, N68);
nand NAND2 (N170, N165, N30);
xor XOR2 (N171, N170, N92);
or OR4 (N172, N155, N51, N170, N49);
or OR3 (N173, N164, N69, N87);
nand NAND3 (N174, N173, N63, N82);
not NOT1 (N175, N172);
and AND3 (N176, N174, N162, N40);
buf BUF1 (N177, N136);
and AND2 (N178, N168, N167);
or OR3 (N179, N176, N174, N71);
buf BUF1 (N180, N154);
not NOT1 (N181, N180);
and AND4 (N182, N177, N34, N48, N103);
or OR2 (N183, N178, N118);
xor XOR2 (N184, N182, N173);
nand NAND4 (N185, N171, N15, N17, N30);
and AND3 (N186, N184, N90, N134);
not NOT1 (N187, N166);
not NOT1 (N188, N181);
xor XOR2 (N189, N188, N180);
xor XOR2 (N190, N189, N123);
not NOT1 (N191, N190);
buf BUF1 (N192, N169);
nand NAND4 (N193, N150, N2, N157, N173);
nand NAND3 (N194, N193, N122, N79);
xor XOR2 (N195, N187, N71);
not NOT1 (N196, N195);
nand NAND3 (N197, N186, N102, N76);
xor XOR2 (N198, N196, N141);
and AND3 (N199, N191, N22, N85);
xor XOR2 (N200, N175, N151);
buf BUF1 (N201, N200);
nor NOR4 (N202, N185, N134, N90, N176);
or OR4 (N203, N202, N6, N38, N111);
xor XOR2 (N204, N199, N170);
nand NAND3 (N205, N183, N26, N38);
nand NAND2 (N206, N198, N101);
and AND3 (N207, N179, N37, N183);
nor NOR2 (N208, N203, N36);
nor NOR4 (N209, N208, N179, N181, N3);
or OR2 (N210, N205, N96);
nand NAND2 (N211, N201, N177);
nor NOR2 (N212, N209, N89);
or OR4 (N213, N156, N55, N54, N99);
and AND2 (N214, N211, N64);
not NOT1 (N215, N214);
buf BUF1 (N216, N204);
xor XOR2 (N217, N215, N56);
not NOT1 (N218, N206);
and AND2 (N219, N192, N96);
buf BUF1 (N220, N197);
or OR3 (N221, N217, N96, N125);
nor NOR2 (N222, N220, N212);
and AND3 (N223, N38, N28, N97);
buf BUF1 (N224, N222);
and AND3 (N225, N224, N159, N41);
nand NAND2 (N226, N207, N197);
not NOT1 (N227, N218);
buf BUF1 (N228, N227);
or OR2 (N229, N219, N88);
nand NAND4 (N230, N228, N196, N54, N120);
nand NAND4 (N231, N194, N66, N129, N8);
and AND4 (N232, N210, N35, N222, N177);
nand NAND4 (N233, N221, N199, N13, N126);
nor NOR3 (N234, N232, N69, N44);
buf BUF1 (N235, N230);
xor XOR2 (N236, N234, N134);
nand NAND2 (N237, N235, N38);
nor NOR4 (N238, N226, N161, N161, N160);
not NOT1 (N239, N238);
not NOT1 (N240, N236);
nor NOR4 (N241, N223, N135, N125, N224);
nand NAND2 (N242, N239, N46);
nand NAND3 (N243, N229, N153, N67);
nor NOR4 (N244, N240, N133, N14, N10);
and AND2 (N245, N216, N157);
nand NAND4 (N246, N237, N230, N46, N134);
buf BUF1 (N247, N233);
buf BUF1 (N248, N241);
not NOT1 (N249, N213);
xor XOR2 (N250, N243, N27);
nor NOR2 (N251, N244, N223);
nor NOR2 (N252, N247, N24);
nand NAND3 (N253, N245, N203, N143);
not NOT1 (N254, N252);
and AND3 (N255, N225, N83, N85);
not NOT1 (N256, N242);
not NOT1 (N257, N249);
not NOT1 (N258, N253);
xor XOR2 (N259, N258, N212);
xor XOR2 (N260, N248, N97);
nor NOR2 (N261, N260, N94);
nor NOR4 (N262, N250, N148, N245, N100);
and AND4 (N263, N257, N157, N47, N47);
and AND2 (N264, N255, N75);
nand NAND3 (N265, N262, N247, N246);
nand NAND2 (N266, N84, N230);
or OR3 (N267, N256, N194, N75);
buf BUF1 (N268, N254);
and AND2 (N269, N261, N100);
not NOT1 (N270, N231);
xor XOR2 (N271, N259, N171);
not NOT1 (N272, N268);
not NOT1 (N273, N269);
and AND2 (N274, N266, N108);
not NOT1 (N275, N274);
buf BUF1 (N276, N267);
nor NOR4 (N277, N273, N191, N200, N30);
buf BUF1 (N278, N276);
nor NOR3 (N279, N270, N185, N203);
nand NAND3 (N280, N271, N162, N94);
and AND4 (N281, N280, N84, N137, N224);
buf BUF1 (N282, N251);
or OR3 (N283, N282, N88, N92);
xor XOR2 (N284, N272, N203);
nand NAND2 (N285, N265, N282);
not NOT1 (N286, N279);
and AND3 (N287, N275, N70, N161);
xor XOR2 (N288, N284, N25);
buf BUF1 (N289, N278);
or OR3 (N290, N285, N199, N237);
or OR2 (N291, N288, N239);
buf BUF1 (N292, N290);
nor NOR2 (N293, N264, N233);
nor NOR3 (N294, N287, N165, N240);
not NOT1 (N295, N292);
nand NAND2 (N296, N263, N62);
nor NOR4 (N297, N296, N106, N139, N136);
nand NAND3 (N298, N289, N3, N100);
and AND4 (N299, N283, N211, N170, N42);
or OR2 (N300, N298, N37);
xor XOR2 (N301, N294, N251);
buf BUF1 (N302, N297);
xor XOR2 (N303, N300, N234);
not NOT1 (N304, N299);
and AND3 (N305, N291, N7, N54);
and AND3 (N306, N281, N280, N282);
and AND2 (N307, N302, N271);
and AND3 (N308, N301, N195, N57);
or OR4 (N309, N304, N193, N66, N29);
nand NAND2 (N310, N306, N265);
or OR3 (N311, N277, N176, N77);
buf BUF1 (N312, N309);
not NOT1 (N313, N295);
nor NOR2 (N314, N303, N91);
xor XOR2 (N315, N311, N78);
not NOT1 (N316, N293);
and AND2 (N317, N307, N170);
not NOT1 (N318, N314);
xor XOR2 (N319, N308, N315);
nor NOR4 (N320, N170, N317, N311, N7);
nand NAND2 (N321, N313, N142);
nor NOR2 (N322, N65, N240);
and AND2 (N323, N312, N5);
and AND3 (N324, N319, N197, N71);
nand NAND2 (N325, N318, N140);
nand NAND4 (N326, N325, N117, N152, N24);
nor NOR3 (N327, N324, N55, N201);
or OR4 (N328, N327, N33, N211, N167);
not NOT1 (N329, N328);
not NOT1 (N330, N316);
buf BUF1 (N331, N326);
nand NAND3 (N332, N329, N114, N80);
and AND3 (N333, N305, N171, N75);
not NOT1 (N334, N310);
buf BUF1 (N335, N321);
nand NAND4 (N336, N332, N217, N142, N23);
xor XOR2 (N337, N336, N261);
xor XOR2 (N338, N330, N141);
not NOT1 (N339, N337);
or OR4 (N340, N339, N166, N160, N280);
nor NOR4 (N341, N335, N71, N188, N95);
or OR4 (N342, N340, N118, N148, N282);
buf BUF1 (N343, N320);
buf BUF1 (N344, N333);
or OR3 (N345, N344, N34, N181);
nor NOR3 (N346, N286, N297, N330);
and AND4 (N347, N343, N148, N81, N200);
buf BUF1 (N348, N347);
buf BUF1 (N349, N322);
nor NOR4 (N350, N346, N77, N330, N321);
and AND4 (N351, N323, N187, N187, N334);
not NOT1 (N352, N68);
nand NAND3 (N353, N338, N299, N20);
not NOT1 (N354, N351);
xor XOR2 (N355, N345, N267);
nand NAND4 (N356, N354, N159, N297, N50);
not NOT1 (N357, N341);
nand NAND2 (N358, N356, N255);
and AND4 (N359, N350, N308, N138, N67);
nand NAND4 (N360, N357, N252, N244, N198);
nor NOR4 (N361, N349, N118, N104, N162);
nand NAND4 (N362, N353, N100, N337, N143);
or OR4 (N363, N361, N114, N318, N68);
and AND2 (N364, N359, N278);
and AND3 (N365, N362, N165, N201);
nor NOR2 (N366, N358, N122);
not NOT1 (N367, N364);
or OR3 (N368, N367, N46, N176);
not NOT1 (N369, N331);
not NOT1 (N370, N348);
xor XOR2 (N371, N370, N285);
buf BUF1 (N372, N371);
nor NOR4 (N373, N355, N232, N262, N59);
and AND4 (N374, N369, N181, N104, N24);
buf BUF1 (N375, N360);
xor XOR2 (N376, N352, N172);
buf BUF1 (N377, N366);
and AND4 (N378, N377, N103, N249, N355);
not NOT1 (N379, N374);
xor XOR2 (N380, N379, N347);
not NOT1 (N381, N372);
nor NOR3 (N382, N375, N69, N214);
nand NAND3 (N383, N363, N285, N228);
nand NAND3 (N384, N376, N61, N382);
buf BUF1 (N385, N308);
xor XOR2 (N386, N368, N70);
nor NOR2 (N387, N342, N17);
nor NOR4 (N388, N378, N201, N366, N118);
buf BUF1 (N389, N373);
not NOT1 (N390, N386);
nand NAND3 (N391, N385, N101, N21);
nor NOR3 (N392, N389, N164, N187);
or OR3 (N393, N380, N334, N54);
and AND3 (N394, N384, N70, N105);
nand NAND3 (N395, N392, N358, N351);
and AND4 (N396, N388, N67, N156, N189);
not NOT1 (N397, N381);
and AND2 (N398, N391, N339);
not NOT1 (N399, N393);
and AND4 (N400, N365, N260, N253, N37);
and AND2 (N401, N383, N86);
or OR2 (N402, N390, N179);
or OR3 (N403, N401, N96, N160);
and AND3 (N404, N398, N9, N156);
buf BUF1 (N405, N402);
xor XOR2 (N406, N387, N368);
and AND3 (N407, N399, N34, N35);
xor XOR2 (N408, N407, N265);
or OR4 (N409, N396, N262, N149, N66);
buf BUF1 (N410, N403);
not NOT1 (N411, N404);
nor NOR2 (N412, N411, N34);
nand NAND2 (N413, N412, N257);
nor NOR4 (N414, N405, N322, N137, N369);
buf BUF1 (N415, N409);
nor NOR4 (N416, N408, N200, N197, N101);
nand NAND3 (N417, N394, N278, N260);
or OR4 (N418, N395, N276, N88, N93);
nor NOR2 (N419, N406, N65);
nor NOR2 (N420, N418, N345);
buf BUF1 (N421, N397);
not NOT1 (N422, N416);
nand NAND3 (N423, N415, N109, N335);
not NOT1 (N424, N410);
nor NOR4 (N425, N400, N102, N317, N146);
or OR4 (N426, N417, N238, N260, N323);
xor XOR2 (N427, N420, N113);
xor XOR2 (N428, N414, N19);
not NOT1 (N429, N425);
and AND4 (N430, N424, N13, N400, N251);
xor XOR2 (N431, N421, N29);
and AND2 (N432, N429, N330);
buf BUF1 (N433, N428);
and AND2 (N434, N431, N179);
nor NOR4 (N435, N413, N128, N104, N252);
and AND4 (N436, N433, N334, N32, N78);
nor NOR4 (N437, N422, N29, N130, N176);
nand NAND3 (N438, N423, N224, N48);
nand NAND3 (N439, N435, N182, N380);
and AND2 (N440, N439, N59);
and AND3 (N441, N430, N322, N138);
not NOT1 (N442, N437);
or OR3 (N443, N432, N274, N354);
and AND3 (N444, N426, N44, N168);
nor NOR4 (N445, N443, N383, N171, N102);
buf BUF1 (N446, N438);
nor NOR4 (N447, N441, N367, N286, N13);
xor XOR2 (N448, N445, N261);
or OR2 (N449, N444, N281);
and AND3 (N450, N447, N307, N173);
nor NOR3 (N451, N450, N336, N424);
not NOT1 (N452, N442);
buf BUF1 (N453, N452);
buf BUF1 (N454, N427);
and AND4 (N455, N453, N160, N43, N11);
nor NOR4 (N456, N419, N173, N454, N148);
nand NAND4 (N457, N62, N361, N388, N336);
xor XOR2 (N458, N446, N20);
nand NAND4 (N459, N440, N29, N83, N379);
buf BUF1 (N460, N451);
nand NAND2 (N461, N448, N60);
buf BUF1 (N462, N449);
xor XOR2 (N463, N459, N393);
buf BUF1 (N464, N457);
not NOT1 (N465, N464);
not NOT1 (N466, N465);
and AND3 (N467, N456, N358, N106);
and AND4 (N468, N434, N464, N383, N464);
and AND4 (N469, N458, N84, N247, N397);
and AND4 (N470, N469, N373, N360, N303);
xor XOR2 (N471, N467, N96);
buf BUF1 (N472, N460);
nand NAND3 (N473, N455, N56, N359);
nand NAND2 (N474, N436, N253);
and AND2 (N475, N468, N71);
or OR4 (N476, N470, N78, N321, N75);
or OR3 (N477, N462, N415, N354);
and AND4 (N478, N475, N42, N421, N124);
xor XOR2 (N479, N472, N327);
and AND3 (N480, N461, N408, N200);
buf BUF1 (N481, N471);
nand NAND3 (N482, N473, N95, N29);
nand NAND3 (N483, N480, N185, N395);
nand NAND3 (N484, N477, N45, N84);
xor XOR2 (N485, N466, N40);
nand NAND3 (N486, N474, N22, N85);
not NOT1 (N487, N483);
or OR4 (N488, N476, N140, N153, N134);
nand NAND2 (N489, N478, N349);
not NOT1 (N490, N487);
nor NOR4 (N491, N485, N118, N17, N335);
xor XOR2 (N492, N490, N300);
and AND3 (N493, N488, N272, N417);
and AND2 (N494, N493, N360);
and AND4 (N495, N491, N493, N37, N308);
not NOT1 (N496, N463);
not NOT1 (N497, N482);
xor XOR2 (N498, N479, N64);
or OR4 (N499, N484, N126, N285, N429);
buf BUF1 (N500, N486);
nor NOR3 (N501, N492, N316, N201);
nor NOR4 (N502, N495, N389, N194, N196);
or OR4 (N503, N499, N298, N240, N155);
nor NOR2 (N504, N481, N457);
and AND3 (N505, N496, N330, N137);
not NOT1 (N506, N504);
xor XOR2 (N507, N500, N48);
buf BUF1 (N508, N501);
xor XOR2 (N509, N497, N57);
nor NOR2 (N510, N498, N268);
xor XOR2 (N511, N509, N97);
xor XOR2 (N512, N510, N210);
nand NAND3 (N513, N494, N433, N194);
or OR4 (N514, N507, N184, N174, N341);
nand NAND3 (N515, N511, N17, N90);
nor NOR2 (N516, N513, N311);
xor XOR2 (N517, N515, N186);
buf BUF1 (N518, N514);
nand NAND3 (N519, N505, N133, N316);
or OR3 (N520, N508, N113, N134);
xor XOR2 (N521, N503, N443);
nor NOR2 (N522, N512, N414);
nor NOR3 (N523, N519, N331, N374);
xor XOR2 (N524, N502, N367);
buf BUF1 (N525, N489);
nor NOR3 (N526, N516, N229, N425);
buf BUF1 (N527, N526);
nand NAND4 (N528, N518, N438, N182, N142);
nand NAND4 (N529, N523, N340, N16, N117);
nor NOR4 (N530, N524, N376, N172, N27);
nor NOR4 (N531, N529, N460, N270, N10);
or OR2 (N532, N530, N102);
xor XOR2 (N533, N531, N325);
or OR3 (N534, N520, N126, N111);
and AND4 (N535, N521, N529, N69, N51);
or OR4 (N536, N528, N450, N450, N321);
and AND4 (N537, N506, N310, N60, N262);
not NOT1 (N538, N532);
xor XOR2 (N539, N537, N403);
nor NOR3 (N540, N535, N398, N395);
nand NAND4 (N541, N527, N27, N312, N536);
nand NAND3 (N542, N166, N269, N25);
nor NOR3 (N543, N517, N133, N523);
not NOT1 (N544, N525);
or OR2 (N545, N522, N326);
and AND3 (N546, N538, N88, N349);
buf BUF1 (N547, N542);
or OR4 (N548, N534, N425, N419, N346);
nand NAND2 (N549, N545, N79);
xor XOR2 (N550, N533, N33);
not NOT1 (N551, N541);
nor NOR3 (N552, N544, N480, N130);
or OR3 (N553, N550, N409, N331);
buf BUF1 (N554, N549);
xor XOR2 (N555, N546, N336);
or OR4 (N556, N555, N320, N312, N206);
and AND4 (N557, N552, N256, N324, N5);
nand NAND2 (N558, N547, N402);
and AND3 (N559, N558, N43, N164);
xor XOR2 (N560, N543, N242);
buf BUF1 (N561, N557);
xor XOR2 (N562, N554, N198);
nor NOR4 (N563, N551, N5, N25, N412);
and AND4 (N564, N559, N232, N207, N446);
nand NAND4 (N565, N556, N39, N479, N363);
or OR4 (N566, N540, N266, N182, N426);
nand NAND3 (N567, N548, N446, N165);
and AND4 (N568, N564, N305, N203, N245);
nand NAND3 (N569, N565, N373, N457);
not NOT1 (N570, N566);
xor XOR2 (N571, N563, N445);
buf BUF1 (N572, N570);
not NOT1 (N573, N553);
and AND4 (N574, N568, N73, N7, N362);
nand NAND2 (N575, N572, N120);
and AND3 (N576, N573, N561, N538);
or OR3 (N577, N407, N522, N69);
nand NAND4 (N578, N571, N193, N122, N170);
buf BUF1 (N579, N560);
not NOT1 (N580, N539);
nand NAND4 (N581, N578, N282, N116, N558);
nand NAND3 (N582, N581, N128, N502);
or OR4 (N583, N569, N130, N243, N271);
or OR2 (N584, N582, N255);
buf BUF1 (N585, N575);
or OR2 (N586, N562, N444);
xor XOR2 (N587, N576, N264);
and AND3 (N588, N583, N30, N56);
nor NOR3 (N589, N580, N491, N501);
or OR2 (N590, N588, N8);
not NOT1 (N591, N587);
and AND3 (N592, N567, N500, N350);
and AND4 (N593, N586, N339, N185, N558);
nand NAND3 (N594, N584, N322, N156);
buf BUF1 (N595, N574);
xor XOR2 (N596, N595, N260);
buf BUF1 (N597, N577);
nand NAND4 (N598, N593, N448, N53, N478);
not NOT1 (N599, N579);
xor XOR2 (N600, N590, N354);
not NOT1 (N601, N598);
buf BUF1 (N602, N585);
and AND3 (N603, N596, N446, N210);
nor NOR3 (N604, N594, N399, N358);
xor XOR2 (N605, N600, N184);
buf BUF1 (N606, N597);
not NOT1 (N607, N601);
xor XOR2 (N608, N592, N529);
buf BUF1 (N609, N608);
nor NOR4 (N610, N604, N32, N367, N242);
and AND3 (N611, N602, N71, N388);
or OR2 (N612, N603, N140);
or OR4 (N613, N589, N256, N280, N305);
nor NOR2 (N614, N610, N106);
buf BUF1 (N615, N609);
and AND2 (N616, N614, N316);
nor NOR4 (N617, N613, N144, N436, N413);
nor NOR3 (N618, N605, N62, N416);
nand NAND4 (N619, N618, N228, N31, N44);
nor NOR2 (N620, N617, N128);
xor XOR2 (N621, N606, N504);
buf BUF1 (N622, N621);
and AND2 (N623, N619, N236);
xor XOR2 (N624, N616, N431);
nor NOR3 (N625, N599, N479, N122);
nand NAND2 (N626, N624, N522);
nor NOR3 (N627, N615, N272, N42);
xor XOR2 (N628, N607, N106);
not NOT1 (N629, N620);
nand NAND2 (N630, N612, N363);
nor NOR4 (N631, N630, N606, N584, N37);
nand NAND2 (N632, N622, N292);
nand NAND2 (N633, N627, N472);
or OR3 (N634, N633, N131, N544);
nor NOR4 (N635, N631, N11, N496, N166);
xor XOR2 (N636, N635, N314);
or OR2 (N637, N636, N95);
nor NOR4 (N638, N628, N602, N374, N190);
nand NAND3 (N639, N591, N280, N297);
xor XOR2 (N640, N625, N53);
buf BUF1 (N641, N638);
buf BUF1 (N642, N639);
not NOT1 (N643, N629);
or OR4 (N644, N634, N40, N544, N442);
nor NOR3 (N645, N642, N608, N27);
buf BUF1 (N646, N611);
nor NOR4 (N647, N643, N553, N84, N115);
buf BUF1 (N648, N640);
buf BUF1 (N649, N645);
not NOT1 (N650, N646);
nor NOR3 (N651, N649, N71, N182);
buf BUF1 (N652, N641);
xor XOR2 (N653, N637, N147);
xor XOR2 (N654, N648, N465);
and AND4 (N655, N654, N244, N606, N415);
xor XOR2 (N656, N651, N172);
or OR4 (N657, N647, N72, N154, N98);
nand NAND3 (N658, N655, N99, N310);
or OR4 (N659, N626, N580, N172, N349);
not NOT1 (N660, N656);
not NOT1 (N661, N650);
or OR3 (N662, N652, N33, N377);
buf BUF1 (N663, N659);
or OR4 (N664, N632, N223, N210, N522);
and AND2 (N665, N623, N146);
and AND3 (N666, N657, N59, N321);
nand NAND3 (N667, N665, N648, N308);
and AND4 (N668, N662, N480, N521, N6);
and AND2 (N669, N661, N597);
and AND3 (N670, N667, N17, N597);
nand NAND3 (N671, N669, N337, N654);
not NOT1 (N672, N666);
not NOT1 (N673, N663);
not NOT1 (N674, N664);
xor XOR2 (N675, N658, N570);
or OR3 (N676, N668, N305, N123);
or OR3 (N677, N673, N344, N383);
and AND2 (N678, N670, N572);
buf BUF1 (N679, N677);
xor XOR2 (N680, N679, N633);
nand NAND3 (N681, N678, N129, N264);
not NOT1 (N682, N674);
nor NOR2 (N683, N682, N258);
and AND3 (N684, N680, N491, N611);
and AND3 (N685, N676, N19, N404);
xor XOR2 (N686, N683, N17);
nor NOR4 (N687, N672, N261, N365, N186);
nand NAND2 (N688, N681, N676);
nor NOR4 (N689, N644, N205, N86, N540);
not NOT1 (N690, N653);
nand NAND2 (N691, N675, N509);
buf BUF1 (N692, N688);
xor XOR2 (N693, N689, N190);
nand NAND2 (N694, N685, N268);
nand NAND4 (N695, N660, N501, N545, N145);
nand NAND2 (N696, N692, N183);
and AND4 (N697, N687, N182, N189, N468);
nor NOR3 (N698, N693, N56, N123);
nand NAND4 (N699, N671, N307, N177, N316);
nor NOR3 (N700, N691, N100, N470);
and AND4 (N701, N699, N234, N213, N73);
xor XOR2 (N702, N698, N141);
or OR2 (N703, N695, N231);
and AND3 (N704, N702, N288, N541);
nand NAND4 (N705, N696, N605, N372, N393);
buf BUF1 (N706, N700);
or OR4 (N707, N686, N584, N598, N270);
or OR3 (N708, N706, N146, N223);
not NOT1 (N709, N708);
nor NOR2 (N710, N684, N433);
xor XOR2 (N711, N705, N178);
buf BUF1 (N712, N710);
or OR4 (N713, N690, N7, N624, N701);
nand NAND3 (N714, N419, N218, N374);
nor NOR3 (N715, N714, N11, N373);
nand NAND2 (N716, N709, N147);
nor NOR4 (N717, N707, N22, N191, N306);
nand NAND2 (N718, N712, N549);
nand NAND3 (N719, N717, N5, N496);
buf BUF1 (N720, N694);
buf BUF1 (N721, N720);
xor XOR2 (N722, N711, N113);
buf BUF1 (N723, N718);
and AND3 (N724, N721, N68, N104);
nand NAND4 (N725, N724, N453, N574, N501);
buf BUF1 (N726, N704);
nand NAND3 (N727, N703, N625, N47);
and AND4 (N728, N719, N14, N488, N604);
and AND4 (N729, N722, N636, N246, N523);
xor XOR2 (N730, N727, N142);
and AND2 (N731, N715, N385);
not NOT1 (N732, N723);
not NOT1 (N733, N732);
not NOT1 (N734, N697);
and AND3 (N735, N713, N704, N603);
not NOT1 (N736, N730);
nor NOR3 (N737, N728, N253, N418);
and AND3 (N738, N731, N711, N680);
not NOT1 (N739, N733);
nor NOR4 (N740, N734, N310, N675, N7);
buf BUF1 (N741, N736);
and AND2 (N742, N740, N481);
or OR3 (N743, N726, N152, N189);
buf BUF1 (N744, N739);
nand NAND3 (N745, N729, N346, N718);
buf BUF1 (N746, N744);
nor NOR4 (N747, N745, N292, N4, N535);
xor XOR2 (N748, N725, N514);
not NOT1 (N749, N737);
not NOT1 (N750, N716);
nor NOR4 (N751, N742, N2, N35, N436);
xor XOR2 (N752, N750, N176);
or OR4 (N753, N749, N744, N645, N448);
or OR4 (N754, N753, N445, N609, N132);
or OR3 (N755, N743, N376, N173);
nand NAND2 (N756, N741, N127);
not NOT1 (N757, N735);
nand NAND3 (N758, N757, N721, N598);
buf BUF1 (N759, N747);
xor XOR2 (N760, N752, N744);
nand NAND2 (N761, N738, N476);
nand NAND4 (N762, N746, N11, N106, N349);
buf BUF1 (N763, N760);
and AND3 (N764, N751, N47, N685);
or OR3 (N765, N754, N335, N275);
and AND2 (N766, N764, N326);
xor XOR2 (N767, N761, N306);
and AND4 (N768, N755, N623, N176, N79);
buf BUF1 (N769, N759);
and AND4 (N770, N765, N545, N592, N493);
nor NOR2 (N771, N758, N550);
and AND3 (N772, N763, N758, N342);
nor NOR2 (N773, N770, N624);
nand NAND3 (N774, N771, N96, N75);
nor NOR4 (N775, N769, N189, N715, N650);
nor NOR2 (N776, N774, N96);
nor NOR3 (N777, N756, N278, N701);
nor NOR3 (N778, N748, N124, N745);
nand NAND2 (N779, N775, N91);
nand NAND3 (N780, N772, N93, N294);
nor NOR4 (N781, N779, N229, N738, N568);
buf BUF1 (N782, N778);
xor XOR2 (N783, N768, N188);
or OR3 (N784, N773, N300, N332);
nor NOR3 (N785, N776, N59, N383);
nor NOR3 (N786, N767, N164, N307);
not NOT1 (N787, N783);
or OR4 (N788, N777, N22, N83, N515);
nor NOR2 (N789, N780, N432);
xor XOR2 (N790, N784, N525);
nor NOR2 (N791, N781, N221);
nor NOR2 (N792, N766, N521);
buf BUF1 (N793, N762);
nor NOR4 (N794, N789, N37, N745, N742);
and AND2 (N795, N788, N419);
buf BUF1 (N796, N791);
not NOT1 (N797, N790);
nor NOR4 (N798, N797, N147, N314, N637);
not NOT1 (N799, N794);
and AND3 (N800, N792, N772, N664);
or OR2 (N801, N800, N673);
not NOT1 (N802, N785);
nor NOR2 (N803, N801, N226);
and AND2 (N804, N803, N136);
buf BUF1 (N805, N793);
not NOT1 (N806, N786);
not NOT1 (N807, N806);
buf BUF1 (N808, N796);
nand NAND3 (N809, N805, N112, N315);
not NOT1 (N810, N804);
not NOT1 (N811, N802);
not NOT1 (N812, N810);
buf BUF1 (N813, N795);
and AND2 (N814, N811, N265);
nor NOR4 (N815, N782, N232, N84, N586);
not NOT1 (N816, N814);
xor XOR2 (N817, N809, N529);
or OR4 (N818, N816, N119, N555, N160);
nand NAND2 (N819, N798, N730);
not NOT1 (N820, N799);
nor NOR2 (N821, N812, N376);
and AND4 (N822, N808, N352, N682, N680);
and AND2 (N823, N815, N753);
not NOT1 (N824, N818);
xor XOR2 (N825, N817, N159);
and AND2 (N826, N819, N221);
nor NOR2 (N827, N813, N235);
xor XOR2 (N828, N821, N691);
and AND2 (N829, N824, N368);
nor NOR3 (N830, N828, N329, N619);
not NOT1 (N831, N826);
and AND4 (N832, N830, N542, N28, N707);
nor NOR4 (N833, N787, N303, N696, N756);
xor XOR2 (N834, N832, N832);
buf BUF1 (N835, N834);
or OR3 (N836, N822, N597, N660);
not NOT1 (N837, N823);
buf BUF1 (N838, N831);
not NOT1 (N839, N835);
nor NOR2 (N840, N807, N758);
not NOT1 (N841, N837);
and AND4 (N842, N840, N472, N119, N41);
or OR4 (N843, N833, N587, N721, N370);
nor NOR2 (N844, N843, N303);
and AND3 (N845, N839, N780, N361);
not NOT1 (N846, N844);
nor NOR4 (N847, N842, N493, N572, N359);
or OR2 (N848, N841, N735);
and AND4 (N849, N838, N480, N113, N496);
buf BUF1 (N850, N829);
buf BUF1 (N851, N820);
nor NOR3 (N852, N845, N807, N404);
buf BUF1 (N853, N848);
buf BUF1 (N854, N849);
or OR3 (N855, N846, N839, N557);
or OR2 (N856, N825, N690);
nor NOR2 (N857, N853, N238);
xor XOR2 (N858, N855, N5);
buf BUF1 (N859, N854);
and AND4 (N860, N858, N31, N24, N725);
nor NOR4 (N861, N847, N591, N79, N322);
or OR3 (N862, N836, N828, N305);
xor XOR2 (N863, N859, N594);
nand NAND4 (N864, N857, N283, N629, N386);
buf BUF1 (N865, N851);
buf BUF1 (N866, N852);
xor XOR2 (N867, N864, N834);
and AND2 (N868, N863, N51);
nand NAND2 (N869, N850, N274);
and AND3 (N870, N868, N564, N237);
and AND4 (N871, N860, N129, N116, N617);
buf BUF1 (N872, N867);
xor XOR2 (N873, N869, N186);
nor NOR3 (N874, N861, N323, N230);
buf BUF1 (N875, N873);
not NOT1 (N876, N866);
xor XOR2 (N877, N876, N752);
nand NAND4 (N878, N875, N498, N533, N350);
nor NOR4 (N879, N827, N6, N551, N552);
and AND3 (N880, N865, N695, N485);
nand NAND2 (N881, N870, N542);
or OR2 (N882, N879, N657);
nor NOR2 (N883, N872, N823);
or OR2 (N884, N862, N322);
not NOT1 (N885, N871);
xor XOR2 (N886, N882, N247);
xor XOR2 (N887, N884, N145);
xor XOR2 (N888, N881, N563);
not NOT1 (N889, N885);
not NOT1 (N890, N886);
buf BUF1 (N891, N887);
buf BUF1 (N892, N878);
or OR3 (N893, N888, N285, N286);
or OR2 (N894, N883, N123);
nand NAND4 (N895, N889, N702, N403, N452);
buf BUF1 (N896, N894);
nor NOR2 (N897, N890, N582);
not NOT1 (N898, N874);
buf BUF1 (N899, N897);
not NOT1 (N900, N899);
buf BUF1 (N901, N900);
nor NOR4 (N902, N877, N641, N158, N582);
and AND3 (N903, N896, N641, N218);
buf BUF1 (N904, N892);
or OR4 (N905, N903, N36, N457, N182);
nand NAND4 (N906, N880, N133, N610, N16);
or OR4 (N907, N906, N399, N68, N101);
or OR4 (N908, N891, N319, N786, N432);
and AND4 (N909, N907, N191, N271, N23);
not NOT1 (N910, N909);
not NOT1 (N911, N898);
nand NAND3 (N912, N856, N707, N141);
or OR3 (N913, N901, N553, N897);
or OR2 (N914, N902, N517);
and AND2 (N915, N913, N566);
and AND2 (N916, N914, N597);
nand NAND4 (N917, N908, N125, N392, N416);
and AND4 (N918, N915, N855, N190, N681);
not NOT1 (N919, N911);
xor XOR2 (N920, N910, N611);
buf BUF1 (N921, N912);
xor XOR2 (N922, N893, N781);
xor XOR2 (N923, N920, N825);
nor NOR4 (N924, N916, N915, N626, N440);
or OR3 (N925, N922, N320, N277);
or OR4 (N926, N905, N38, N598, N743);
not NOT1 (N927, N919);
xor XOR2 (N928, N924, N71);
and AND4 (N929, N917, N223, N80, N290);
nor NOR2 (N930, N928, N140);
and AND4 (N931, N926, N55, N323, N645);
buf BUF1 (N932, N918);
and AND3 (N933, N929, N772, N303);
nand NAND3 (N934, N930, N372, N889);
nand NAND3 (N935, N925, N55, N583);
nand NAND2 (N936, N934, N821);
nand NAND4 (N937, N936, N328, N708, N181);
and AND2 (N938, N937, N192);
buf BUF1 (N939, N938);
not NOT1 (N940, N939);
nand NAND2 (N941, N933, N797);
nor NOR4 (N942, N932, N712, N152, N620);
or OR2 (N943, N931, N440);
not NOT1 (N944, N927);
and AND4 (N945, N895, N397, N572, N443);
or OR4 (N946, N944, N609, N617, N35);
nand NAND4 (N947, N942, N868, N487, N744);
xor XOR2 (N948, N941, N148);
not NOT1 (N949, N945);
not NOT1 (N950, N947);
not NOT1 (N951, N935);
buf BUF1 (N952, N948);
and AND3 (N953, N940, N108, N322);
nand NAND3 (N954, N949, N853, N146);
nor NOR2 (N955, N923, N725);
not NOT1 (N956, N955);
nand NAND2 (N957, N951, N420);
nand NAND4 (N958, N952, N848, N397, N230);
not NOT1 (N959, N943);
xor XOR2 (N960, N950, N255);
and AND2 (N961, N956, N542);
not NOT1 (N962, N957);
buf BUF1 (N963, N958);
buf BUF1 (N964, N961);
or OR2 (N965, N921, N63);
buf BUF1 (N966, N959);
xor XOR2 (N967, N960, N257);
xor XOR2 (N968, N953, N813);
and AND3 (N969, N966, N138, N703);
nor NOR2 (N970, N964, N832);
buf BUF1 (N971, N967);
and AND3 (N972, N971, N792, N40);
xor XOR2 (N973, N965, N899);
xor XOR2 (N974, N963, N944);
xor XOR2 (N975, N968, N613);
nand NAND2 (N976, N973, N422);
not NOT1 (N977, N962);
buf BUF1 (N978, N954);
xor XOR2 (N979, N974, N411);
and AND4 (N980, N946, N774, N177, N831);
buf BUF1 (N981, N980);
nand NAND4 (N982, N981, N264, N940, N609);
buf BUF1 (N983, N975);
and AND2 (N984, N983, N415);
not NOT1 (N985, N976);
nand NAND4 (N986, N969, N884, N470, N798);
not NOT1 (N987, N985);
and AND2 (N988, N978, N101);
not NOT1 (N989, N982);
xor XOR2 (N990, N979, N370);
buf BUF1 (N991, N987);
not NOT1 (N992, N988);
buf BUF1 (N993, N970);
xor XOR2 (N994, N984, N760);
buf BUF1 (N995, N992);
and AND3 (N996, N990, N120, N352);
or OR2 (N997, N995, N929);
and AND3 (N998, N994, N32, N140);
nor NOR2 (N999, N977, N397);
nand NAND3 (N1000, N998, N524, N330);
nor NOR4 (N1001, N999, N557, N406, N532);
nand NAND4 (N1002, N1001, N188, N579, N677);
buf BUF1 (N1003, N972);
buf BUF1 (N1004, N904);
and AND2 (N1005, N997, N691);
not NOT1 (N1006, N993);
buf BUF1 (N1007, N1003);
or OR2 (N1008, N989, N133);
not NOT1 (N1009, N1007);
buf BUF1 (N1010, N991);
nor NOR3 (N1011, N986, N451, N522);
not NOT1 (N1012, N1000);
nor NOR3 (N1013, N1006, N583, N856);
xor XOR2 (N1014, N1009, N353);
nor NOR3 (N1015, N1008, N346, N474);
and AND3 (N1016, N1014, N778, N773);
not NOT1 (N1017, N1011);
xor XOR2 (N1018, N1005, N856);
not NOT1 (N1019, N1017);
nor NOR2 (N1020, N1018, N143);
and AND4 (N1021, N1002, N764, N671, N738);
xor XOR2 (N1022, N996, N207);
nand NAND4 (N1023, N1022, N122, N793, N39);
xor XOR2 (N1024, N1010, N1006);
nor NOR4 (N1025, N1024, N371, N605, N286);
nor NOR4 (N1026, N1025, N237, N662, N230);
not NOT1 (N1027, N1020);
nand NAND4 (N1028, N1026, N339, N255, N16);
or OR2 (N1029, N1023, N1020);
nand NAND2 (N1030, N1016, N1024);
nand NAND4 (N1031, N1019, N687, N323, N187);
not NOT1 (N1032, N1015);
xor XOR2 (N1033, N1028, N668);
buf BUF1 (N1034, N1029);
xor XOR2 (N1035, N1013, N179);
nand NAND2 (N1036, N1035, N14);
xor XOR2 (N1037, N1034, N336);
xor XOR2 (N1038, N1012, N469);
not NOT1 (N1039, N1027);
not NOT1 (N1040, N1036);
xor XOR2 (N1041, N1030, N775);
and AND4 (N1042, N1033, N920, N136, N669);
not NOT1 (N1043, N1042);
buf BUF1 (N1044, N1039);
xor XOR2 (N1045, N1038, N836);
or OR3 (N1046, N1037, N601, N113);
buf BUF1 (N1047, N1044);
nor NOR4 (N1048, N1032, N360, N622, N492);
nand NAND3 (N1049, N1041, N568, N186);
or OR3 (N1050, N1021, N282, N83);
and AND4 (N1051, N1031, N714, N36, N859);
nand NAND2 (N1052, N1040, N222);
or OR4 (N1053, N1049, N35, N975, N515);
nor NOR2 (N1054, N1004, N323);
xor XOR2 (N1055, N1051, N685);
not NOT1 (N1056, N1053);
nand NAND2 (N1057, N1043, N192);
and AND3 (N1058, N1048, N983, N744);
buf BUF1 (N1059, N1056);
buf BUF1 (N1060, N1058);
nor NOR4 (N1061, N1059, N931, N412, N467);
nand NAND2 (N1062, N1052, N705);
nand NAND2 (N1063, N1061, N541);
not NOT1 (N1064, N1062);
and AND4 (N1065, N1064, N346, N664, N343);
or OR3 (N1066, N1050, N736, N464);
buf BUF1 (N1067, N1065);
xor XOR2 (N1068, N1066, N922);
or OR2 (N1069, N1063, N238);
nand NAND2 (N1070, N1068, N530);
and AND4 (N1071, N1055, N226, N839, N930);
and AND2 (N1072, N1060, N626);
or OR4 (N1073, N1067, N59, N791, N902);
not NOT1 (N1074, N1046);
nor NOR4 (N1075, N1074, N726, N861, N699);
xor XOR2 (N1076, N1045, N296);
buf BUF1 (N1077, N1075);
nand NAND2 (N1078, N1077, N531);
or OR4 (N1079, N1072, N361, N784, N402);
nand NAND2 (N1080, N1057, N579);
nor NOR2 (N1081, N1047, N903);
buf BUF1 (N1082, N1079);
nand NAND2 (N1083, N1076, N1002);
or OR4 (N1084, N1054, N652, N742, N16);
and AND3 (N1085, N1070, N940, N663);
or OR4 (N1086, N1071, N462, N714, N357);
not NOT1 (N1087, N1085);
or OR2 (N1088, N1073, N696);
not NOT1 (N1089, N1083);
and AND3 (N1090, N1082, N761, N77);
xor XOR2 (N1091, N1084, N490);
buf BUF1 (N1092, N1080);
buf BUF1 (N1093, N1087);
and AND2 (N1094, N1078, N166);
or OR2 (N1095, N1093, N1060);
not NOT1 (N1096, N1089);
xor XOR2 (N1097, N1069, N76);
nand NAND4 (N1098, N1096, N187, N190, N563);
xor XOR2 (N1099, N1088, N458);
nand NAND2 (N1100, N1092, N944);
or OR4 (N1101, N1097, N1025, N159, N66);
buf BUF1 (N1102, N1095);
xor XOR2 (N1103, N1101, N641);
not NOT1 (N1104, N1081);
buf BUF1 (N1105, N1098);
and AND4 (N1106, N1103, N696, N683, N630);
xor XOR2 (N1107, N1099, N303);
or OR3 (N1108, N1107, N221, N741);
not NOT1 (N1109, N1086);
xor XOR2 (N1110, N1105, N821);
not NOT1 (N1111, N1094);
not NOT1 (N1112, N1102);
or OR3 (N1113, N1110, N1033, N406);
not NOT1 (N1114, N1091);
nor NOR3 (N1115, N1114, N9, N990);
not NOT1 (N1116, N1111);
xor XOR2 (N1117, N1109, N530);
nor NOR2 (N1118, N1113, N407);
xor XOR2 (N1119, N1116, N490);
xor XOR2 (N1120, N1108, N157);
xor XOR2 (N1121, N1115, N252);
not NOT1 (N1122, N1106);
buf BUF1 (N1123, N1121);
or OR4 (N1124, N1100, N585, N416, N458);
nand NAND4 (N1125, N1120, N394, N146, N552);
not NOT1 (N1126, N1090);
buf BUF1 (N1127, N1119);
nand NAND3 (N1128, N1126, N939, N579);
nor NOR3 (N1129, N1117, N638, N1049);
or OR4 (N1130, N1125, N170, N140, N105);
nor NOR4 (N1131, N1129, N990, N916, N366);
nand NAND3 (N1132, N1118, N373, N278);
nand NAND4 (N1133, N1122, N758, N216, N1056);
or OR3 (N1134, N1124, N1027, N882);
nor NOR4 (N1135, N1134, N752, N227, N1080);
nor NOR3 (N1136, N1128, N756, N829);
or OR4 (N1137, N1136, N1117, N274, N1081);
not NOT1 (N1138, N1104);
not NOT1 (N1139, N1123);
not NOT1 (N1140, N1135);
and AND4 (N1141, N1140, N1016, N864, N217);
nor NOR2 (N1142, N1139, N512);
not NOT1 (N1143, N1133);
xor XOR2 (N1144, N1112, N1132);
nand NAND4 (N1145, N214, N194, N985, N113);
or OR4 (N1146, N1145, N1023, N189, N701);
nand NAND4 (N1147, N1131, N1080, N590, N687);
xor XOR2 (N1148, N1147, N1142);
buf BUF1 (N1149, N401);
xor XOR2 (N1150, N1138, N869);
and AND3 (N1151, N1127, N52, N407);
and AND3 (N1152, N1130, N475, N269);
buf BUF1 (N1153, N1151);
nor NOR2 (N1154, N1143, N811);
nor NOR4 (N1155, N1144, N301, N574, N742);
buf BUF1 (N1156, N1154);
xor XOR2 (N1157, N1149, N77);
nor NOR4 (N1158, N1150, N31, N301, N465);
and AND3 (N1159, N1156, N445, N1130);
and AND3 (N1160, N1152, N911, N30);
or OR4 (N1161, N1148, N526, N255, N194);
not NOT1 (N1162, N1146);
or OR2 (N1163, N1153, N282);
nor NOR2 (N1164, N1141, N240);
not NOT1 (N1165, N1163);
nor NOR2 (N1166, N1162, N902);
xor XOR2 (N1167, N1155, N438);
buf BUF1 (N1168, N1167);
not NOT1 (N1169, N1164);
not NOT1 (N1170, N1160);
nand NAND2 (N1171, N1159, N181);
buf BUF1 (N1172, N1158);
nor NOR4 (N1173, N1161, N389, N43, N350);
xor XOR2 (N1174, N1173, N936);
nand NAND3 (N1175, N1166, N1116, N138);
buf BUF1 (N1176, N1171);
or OR4 (N1177, N1170, N508, N858, N963);
or OR3 (N1178, N1157, N332, N157);
nand NAND2 (N1179, N1169, N937);
nor NOR4 (N1180, N1177, N978, N276, N1157);
and AND4 (N1181, N1137, N1118, N222, N839);
xor XOR2 (N1182, N1172, N929);
xor XOR2 (N1183, N1168, N489);
xor XOR2 (N1184, N1180, N264);
or OR3 (N1185, N1179, N286, N1013);
not NOT1 (N1186, N1182);
or OR4 (N1187, N1175, N643, N19, N1165);
xor XOR2 (N1188, N341, N1021);
nand NAND2 (N1189, N1186, N1038);
not NOT1 (N1190, N1183);
nand NAND3 (N1191, N1187, N1120, N692);
not NOT1 (N1192, N1191);
not NOT1 (N1193, N1188);
or OR3 (N1194, N1181, N1132, N82);
xor XOR2 (N1195, N1193, N1024);
or OR2 (N1196, N1174, N50);
and AND4 (N1197, N1189, N726, N1116, N1009);
not NOT1 (N1198, N1176);
or OR2 (N1199, N1196, N648);
nand NAND4 (N1200, N1184, N103, N1126, N244);
and AND2 (N1201, N1197, N920);
nand NAND3 (N1202, N1198, N1053, N120);
and AND3 (N1203, N1185, N164, N622);
buf BUF1 (N1204, N1202);
not NOT1 (N1205, N1204);
nor NOR4 (N1206, N1199, N128, N342, N345);
and AND2 (N1207, N1178, N165);
nor NOR2 (N1208, N1195, N372);
nor NOR3 (N1209, N1205, N697, N888);
xor XOR2 (N1210, N1209, N964);
nand NAND2 (N1211, N1192, N739);
not NOT1 (N1212, N1200);
xor XOR2 (N1213, N1190, N537);
nand NAND3 (N1214, N1203, N723, N292);
nand NAND4 (N1215, N1212, N1125, N1052, N375);
nand NAND3 (N1216, N1207, N820, N932);
buf BUF1 (N1217, N1210);
xor XOR2 (N1218, N1206, N1045);
buf BUF1 (N1219, N1214);
nand NAND2 (N1220, N1213, N1102);
buf BUF1 (N1221, N1208);
xor XOR2 (N1222, N1218, N810);
and AND2 (N1223, N1221, N772);
xor XOR2 (N1224, N1216, N486);
not NOT1 (N1225, N1215);
or OR3 (N1226, N1222, N975, N1112);
xor XOR2 (N1227, N1226, N1000);
or OR3 (N1228, N1219, N785, N18);
nand NAND2 (N1229, N1211, N725);
buf BUF1 (N1230, N1227);
nor NOR3 (N1231, N1217, N45, N927);
xor XOR2 (N1232, N1194, N1112);
nor NOR4 (N1233, N1224, N511, N630, N731);
and AND2 (N1234, N1220, N1057);
xor XOR2 (N1235, N1223, N438);
nand NAND2 (N1236, N1230, N195);
or OR3 (N1237, N1225, N42, N309);
or OR2 (N1238, N1201, N1096);
or OR2 (N1239, N1235, N994);
not NOT1 (N1240, N1237);
nand NAND2 (N1241, N1231, N177);
nor NOR2 (N1242, N1241, N1220);
not NOT1 (N1243, N1242);
or OR2 (N1244, N1234, N791);
and AND3 (N1245, N1239, N709, N167);
or OR2 (N1246, N1244, N159);
and AND4 (N1247, N1246, N1228, N1219, N1246);
nand NAND3 (N1248, N853, N696, N1017);
xor XOR2 (N1249, N1233, N1182);
xor XOR2 (N1250, N1248, N765);
buf BUF1 (N1251, N1249);
and AND3 (N1252, N1251, N1176, N100);
nor NOR2 (N1253, N1252, N233);
and AND2 (N1254, N1238, N325);
nor NOR2 (N1255, N1245, N536);
nor NOR3 (N1256, N1254, N633, N388);
not NOT1 (N1257, N1253);
nor NOR2 (N1258, N1257, N425);
buf BUF1 (N1259, N1243);
not NOT1 (N1260, N1232);
not NOT1 (N1261, N1258);
or OR2 (N1262, N1259, N372);
xor XOR2 (N1263, N1236, N461);
or OR3 (N1264, N1263, N1086, N1103);
nand NAND3 (N1265, N1264, N380, N1013);
not NOT1 (N1266, N1229);
or OR2 (N1267, N1265, N1025);
and AND3 (N1268, N1256, N500, N70);
nand NAND3 (N1269, N1240, N707, N138);
xor XOR2 (N1270, N1262, N733);
and AND2 (N1271, N1269, N1209);
xor XOR2 (N1272, N1255, N337);
xor XOR2 (N1273, N1272, N1203);
xor XOR2 (N1274, N1268, N447);
not NOT1 (N1275, N1273);
buf BUF1 (N1276, N1250);
not NOT1 (N1277, N1270);
nand NAND3 (N1278, N1260, N266, N11);
nand NAND3 (N1279, N1267, N184, N658);
nor NOR4 (N1280, N1275, N144, N1103, N175);
nand NAND4 (N1281, N1279, N424, N423, N506);
xor XOR2 (N1282, N1274, N192);
buf BUF1 (N1283, N1276);
nand NAND3 (N1284, N1247, N916, N196);
xor XOR2 (N1285, N1278, N95);
not NOT1 (N1286, N1282);
xor XOR2 (N1287, N1277, N1251);
buf BUF1 (N1288, N1283);
buf BUF1 (N1289, N1280);
not NOT1 (N1290, N1285);
nor NOR2 (N1291, N1286, N786);
nand NAND3 (N1292, N1281, N835, N475);
not NOT1 (N1293, N1271);
or OR4 (N1294, N1292, N39, N678, N147);
nand NAND4 (N1295, N1284, N58, N607, N94);
or OR4 (N1296, N1287, N1254, N1043, N396);
buf BUF1 (N1297, N1289);
or OR4 (N1298, N1295, N962, N803, N1263);
not NOT1 (N1299, N1261);
nand NAND2 (N1300, N1293, N623);
nand NAND2 (N1301, N1296, N880);
nand NAND2 (N1302, N1294, N82);
buf BUF1 (N1303, N1301);
not NOT1 (N1304, N1302);
not NOT1 (N1305, N1304);
or OR2 (N1306, N1303, N1152);
or OR2 (N1307, N1306, N1287);
and AND2 (N1308, N1291, N1230);
xor XOR2 (N1309, N1300, N87);
buf BUF1 (N1310, N1308);
or OR2 (N1311, N1298, N1039);
buf BUF1 (N1312, N1299);
not NOT1 (N1313, N1290);
nor NOR2 (N1314, N1307, N555);
or OR3 (N1315, N1309, N1289, N928);
nor NOR4 (N1316, N1311, N1186, N935, N1282);
and AND4 (N1317, N1305, N634, N1156, N856);
nor NOR3 (N1318, N1316, N202, N739);
and AND4 (N1319, N1313, N590, N1183, N626);
and AND3 (N1320, N1319, N665, N1301);
nor NOR4 (N1321, N1314, N1298, N1223, N1212);
and AND4 (N1322, N1320, N1147, N14, N415);
and AND2 (N1323, N1321, N529);
or OR4 (N1324, N1288, N523, N887, N1110);
and AND3 (N1325, N1322, N83, N1204);
buf BUF1 (N1326, N1312);
nor NOR3 (N1327, N1315, N1139, N416);
nor NOR3 (N1328, N1326, N175, N1308);
and AND3 (N1329, N1317, N733, N839);
not NOT1 (N1330, N1266);
not NOT1 (N1331, N1329);
not NOT1 (N1332, N1330);
nand NAND2 (N1333, N1297, N875);
not NOT1 (N1334, N1325);
buf BUF1 (N1335, N1310);
and AND2 (N1336, N1323, N1116);
or OR4 (N1337, N1324, N842, N616, N475);
or OR2 (N1338, N1331, N1218);
buf BUF1 (N1339, N1318);
nor NOR2 (N1340, N1337, N931);
and AND4 (N1341, N1340, N677, N1147, N924);
or OR2 (N1342, N1328, N268);
xor XOR2 (N1343, N1335, N446);
or OR4 (N1344, N1341, N176, N1188, N1138);
xor XOR2 (N1345, N1342, N318);
nor NOR4 (N1346, N1334, N290, N505, N798);
nand NAND4 (N1347, N1345, N664, N935, N913);
not NOT1 (N1348, N1343);
buf BUF1 (N1349, N1347);
and AND3 (N1350, N1344, N858, N483);
nor NOR4 (N1351, N1350, N976, N628, N265);
or OR4 (N1352, N1346, N1323, N726, N313);
not NOT1 (N1353, N1338);
not NOT1 (N1354, N1336);
nor NOR4 (N1355, N1352, N122, N846, N90);
nor NOR2 (N1356, N1353, N29);
nor NOR2 (N1357, N1354, N5);
xor XOR2 (N1358, N1332, N492);
xor XOR2 (N1359, N1356, N1164);
nor NOR4 (N1360, N1358, N689, N855, N943);
and AND3 (N1361, N1360, N110, N247);
buf BUF1 (N1362, N1327);
and AND2 (N1363, N1351, N1296);
xor XOR2 (N1364, N1362, N281);
buf BUF1 (N1365, N1333);
or OR4 (N1366, N1355, N157, N1209, N1348);
buf BUF1 (N1367, N476);
and AND4 (N1368, N1367, N701, N863, N1333);
buf BUF1 (N1369, N1357);
and AND2 (N1370, N1364, N849);
nand NAND2 (N1371, N1368, N395);
xor XOR2 (N1372, N1361, N1359);
xor XOR2 (N1373, N1192, N758);
nand NAND4 (N1374, N1363, N324, N1046, N96);
not NOT1 (N1375, N1374);
and AND4 (N1376, N1373, N502, N248, N1046);
not NOT1 (N1377, N1339);
and AND3 (N1378, N1370, N726, N236);
or OR4 (N1379, N1378, N1368, N964, N940);
buf BUF1 (N1380, N1372);
and AND2 (N1381, N1371, N219);
or OR3 (N1382, N1366, N21, N1225);
nor NOR2 (N1383, N1349, N392);
nand NAND2 (N1384, N1380, N1265);
xor XOR2 (N1385, N1377, N936);
nand NAND4 (N1386, N1379, N1354, N728, N1165);
or OR2 (N1387, N1383, N174);
or OR4 (N1388, N1384, N605, N755, N989);
buf BUF1 (N1389, N1385);
and AND2 (N1390, N1388, N68);
or OR2 (N1391, N1375, N392);
nor NOR2 (N1392, N1389, N352);
xor XOR2 (N1393, N1387, N846);
xor XOR2 (N1394, N1386, N1066);
nor NOR4 (N1395, N1381, N1220, N286, N646);
nor NOR4 (N1396, N1382, N472, N250, N618);
not NOT1 (N1397, N1392);
not NOT1 (N1398, N1393);
nand NAND2 (N1399, N1397, N483);
xor XOR2 (N1400, N1399, N534);
buf BUF1 (N1401, N1391);
nand NAND4 (N1402, N1400, N617, N809, N1300);
not NOT1 (N1403, N1396);
and AND2 (N1404, N1390, N494);
xor XOR2 (N1405, N1376, N640);
not NOT1 (N1406, N1365);
or OR4 (N1407, N1394, N677, N257, N363);
buf BUF1 (N1408, N1403);
xor XOR2 (N1409, N1395, N299);
nor NOR3 (N1410, N1409, N191, N1151);
nand NAND3 (N1411, N1369, N381, N527);
and AND2 (N1412, N1401, N115);
and AND4 (N1413, N1402, N210, N772, N1254);
xor XOR2 (N1414, N1411, N310);
or OR2 (N1415, N1408, N988);
buf BUF1 (N1416, N1413);
xor XOR2 (N1417, N1410, N967);
or OR2 (N1418, N1414, N993);
nand NAND3 (N1419, N1404, N1255, N357);
and AND2 (N1420, N1419, N581);
nor NOR3 (N1421, N1406, N1311, N65);
or OR4 (N1422, N1421, N42, N547, N745);
nor NOR4 (N1423, N1417, N524, N1064, N854);
or OR4 (N1424, N1420, N574, N1150, N71);
buf BUF1 (N1425, N1423);
nor NOR4 (N1426, N1415, N752, N884, N750);
and AND4 (N1427, N1426, N760, N319, N658);
or OR2 (N1428, N1424, N896);
or OR4 (N1429, N1416, N776, N423, N972);
or OR4 (N1430, N1427, N13, N760, N1350);
xor XOR2 (N1431, N1405, N1028);
and AND2 (N1432, N1431, N1335);
nand NAND2 (N1433, N1412, N535);
xor XOR2 (N1434, N1428, N1423);
or OR3 (N1435, N1434, N253, N485);
not NOT1 (N1436, N1433);
and AND4 (N1437, N1422, N1194, N92, N685);
nand NAND3 (N1438, N1436, N1347, N737);
xor XOR2 (N1439, N1437, N1226);
xor XOR2 (N1440, N1438, N266);
buf BUF1 (N1441, N1432);
buf BUF1 (N1442, N1429);
not NOT1 (N1443, N1430);
nand NAND2 (N1444, N1441, N480);
nor NOR4 (N1445, N1442, N74, N448, N963);
and AND2 (N1446, N1407, N378);
and AND4 (N1447, N1443, N250, N1144, N46);
nand NAND2 (N1448, N1447, N348);
buf BUF1 (N1449, N1448);
not NOT1 (N1450, N1446);
and AND2 (N1451, N1439, N359);
nand NAND4 (N1452, N1451, N324, N1443, N1089);
or OR2 (N1453, N1435, N653);
nand NAND3 (N1454, N1425, N907, N1101);
nor NOR4 (N1455, N1454, N547, N857, N996);
nor NOR3 (N1456, N1445, N1125, N1139);
and AND4 (N1457, N1440, N605, N1172, N304);
buf BUF1 (N1458, N1456);
buf BUF1 (N1459, N1418);
buf BUF1 (N1460, N1458);
and AND3 (N1461, N1459, N967, N697);
xor XOR2 (N1462, N1461, N564);
xor XOR2 (N1463, N1449, N1242);
xor XOR2 (N1464, N1460, N223);
and AND4 (N1465, N1463, N935, N714, N1077);
nor NOR4 (N1466, N1398, N314, N78, N103);
buf BUF1 (N1467, N1466);
or OR4 (N1468, N1464, N962, N1451, N20);
nand NAND3 (N1469, N1465, N752, N322);
and AND4 (N1470, N1455, N438, N14, N75);
xor XOR2 (N1471, N1462, N368);
buf BUF1 (N1472, N1467);
or OR4 (N1473, N1450, N103, N1034, N639);
xor XOR2 (N1474, N1452, N12);
nand NAND4 (N1475, N1468, N631, N1043, N820);
nor NOR2 (N1476, N1457, N1391);
not NOT1 (N1477, N1470);
buf BUF1 (N1478, N1475);
and AND3 (N1479, N1471, N796, N1381);
nand NAND3 (N1480, N1444, N532, N363);
or OR4 (N1481, N1469, N611, N503, N106);
or OR3 (N1482, N1478, N1126, N530);
and AND4 (N1483, N1477, N324, N1473, N126);
not NOT1 (N1484, N99);
or OR2 (N1485, N1481, N1484);
nand NAND2 (N1486, N1021, N111);
or OR4 (N1487, N1486, N1168, N1473, N445);
and AND2 (N1488, N1482, N246);
or OR3 (N1489, N1453, N300, N387);
not NOT1 (N1490, N1476);
and AND4 (N1491, N1490, N1466, N756, N1325);
buf BUF1 (N1492, N1474);
nand NAND2 (N1493, N1485, N1319);
nand NAND4 (N1494, N1493, N1421, N1423, N545);
buf BUF1 (N1495, N1494);
not NOT1 (N1496, N1495);
nand NAND2 (N1497, N1487, N6);
or OR3 (N1498, N1491, N380, N348);
buf BUF1 (N1499, N1489);
nand NAND3 (N1500, N1492, N941, N1341);
or OR2 (N1501, N1499, N88);
nor NOR2 (N1502, N1483, N728);
nand NAND3 (N1503, N1498, N1040, N311);
buf BUF1 (N1504, N1500);
not NOT1 (N1505, N1503);
nand NAND2 (N1506, N1497, N843);
xor XOR2 (N1507, N1506, N918);
not NOT1 (N1508, N1502);
xor XOR2 (N1509, N1504, N1243);
buf BUF1 (N1510, N1508);
buf BUF1 (N1511, N1480);
nor NOR2 (N1512, N1511, N1316);
or OR4 (N1513, N1488, N193, N1215, N1273);
nand NAND2 (N1514, N1507, N167);
not NOT1 (N1515, N1510);
nor NOR3 (N1516, N1509, N1301, N919);
or OR2 (N1517, N1496, N666);
and AND3 (N1518, N1517, N917, N1179);
and AND3 (N1519, N1512, N111, N1041);
buf BUF1 (N1520, N1518);
nor NOR4 (N1521, N1515, N550, N6, N123);
not NOT1 (N1522, N1513);
buf BUF1 (N1523, N1522);
xor XOR2 (N1524, N1520, N1395);
not NOT1 (N1525, N1514);
xor XOR2 (N1526, N1516, N1091);
buf BUF1 (N1527, N1525);
xor XOR2 (N1528, N1527, N970);
xor XOR2 (N1529, N1521, N911);
not NOT1 (N1530, N1479);
or OR3 (N1531, N1501, N542, N559);
xor XOR2 (N1532, N1472, N583);
nor NOR3 (N1533, N1531, N359, N701);
and AND2 (N1534, N1505, N888);
nand NAND4 (N1535, N1534, N368, N353, N869);
not NOT1 (N1536, N1528);
buf BUF1 (N1537, N1524);
and AND4 (N1538, N1526, N981, N98, N413);
buf BUF1 (N1539, N1535);
or OR3 (N1540, N1538, N1461, N8);
and AND3 (N1541, N1530, N1125, N695);
buf BUF1 (N1542, N1519);
xor XOR2 (N1543, N1541, N1024);
buf BUF1 (N1544, N1529);
nand NAND2 (N1545, N1523, N1382);
or OR3 (N1546, N1537, N993, N370);
and AND3 (N1547, N1532, N25, N761);
and AND4 (N1548, N1543, N922, N812, N34);
nor NOR2 (N1549, N1545, N377);
or OR3 (N1550, N1536, N1499, N993);
nor NOR2 (N1551, N1542, N1318);
nor NOR4 (N1552, N1539, N518, N1204, N392);
or OR2 (N1553, N1547, N357);
or OR3 (N1554, N1548, N93, N298);
and AND4 (N1555, N1549, N844, N112, N1513);
nand NAND4 (N1556, N1550, N898, N1404, N940);
nand NAND3 (N1557, N1556, N472, N745);
nand NAND3 (N1558, N1553, N1370, N1492);
not NOT1 (N1559, N1540);
or OR2 (N1560, N1558, N205);
nand NAND3 (N1561, N1533, N1021, N525);
buf BUF1 (N1562, N1559);
xor XOR2 (N1563, N1562, N715);
not NOT1 (N1564, N1555);
buf BUF1 (N1565, N1551);
nor NOR4 (N1566, N1564, N786, N741, N488);
or OR2 (N1567, N1566, N246);
nor NOR3 (N1568, N1546, N257, N1227);
or OR3 (N1569, N1552, N1228, N752);
xor XOR2 (N1570, N1554, N1564);
buf BUF1 (N1571, N1568);
nand NAND4 (N1572, N1565, N1185, N1138, N104);
nand NAND2 (N1573, N1544, N1371);
not NOT1 (N1574, N1573);
xor XOR2 (N1575, N1571, N1162);
and AND4 (N1576, N1561, N663, N1219, N483);
xor XOR2 (N1577, N1560, N348);
nand NAND4 (N1578, N1576, N1464, N30, N1068);
buf BUF1 (N1579, N1570);
xor XOR2 (N1580, N1557, N473);
xor XOR2 (N1581, N1567, N714);
xor XOR2 (N1582, N1577, N555);
xor XOR2 (N1583, N1575, N1094);
buf BUF1 (N1584, N1574);
xor XOR2 (N1585, N1578, N100);
nand NAND4 (N1586, N1569, N1289, N1242, N1039);
xor XOR2 (N1587, N1563, N11);
buf BUF1 (N1588, N1584);
or OR4 (N1589, N1583, N857, N899, N1204);
or OR3 (N1590, N1589, N213, N123);
nor NOR3 (N1591, N1579, N716, N1063);
not NOT1 (N1592, N1591);
or OR3 (N1593, N1581, N1418, N719);
not NOT1 (N1594, N1593);
or OR3 (N1595, N1582, N1101, N1021);
buf BUF1 (N1596, N1586);
nand NAND3 (N1597, N1590, N1324, N1384);
not NOT1 (N1598, N1572);
or OR4 (N1599, N1587, N1113, N1491, N553);
xor XOR2 (N1600, N1594, N1413);
not NOT1 (N1601, N1588);
or OR3 (N1602, N1598, N158, N182);
not NOT1 (N1603, N1601);
nor NOR3 (N1604, N1603, N1407, N933);
and AND2 (N1605, N1599, N907);
nand NAND4 (N1606, N1604, N581, N175, N1437);
and AND3 (N1607, N1600, N201, N1008);
nor NOR3 (N1608, N1585, N149, N1359);
nor NOR4 (N1609, N1592, N755, N1128, N54);
or OR4 (N1610, N1595, N1214, N537, N386);
buf BUF1 (N1611, N1597);
xor XOR2 (N1612, N1611, N1440);
nor NOR2 (N1613, N1608, N1461);
and AND2 (N1614, N1613, N1053);
nand NAND3 (N1615, N1602, N336, N1224);
or OR2 (N1616, N1612, N728);
nand NAND4 (N1617, N1610, N301, N1282, N1017);
nor NOR3 (N1618, N1615, N935, N208);
and AND3 (N1619, N1607, N918, N492);
and AND3 (N1620, N1619, N1056, N757);
buf BUF1 (N1621, N1605);
nand NAND4 (N1622, N1617, N1399, N73, N521);
nor NOR2 (N1623, N1609, N1582);
buf BUF1 (N1624, N1614);
not NOT1 (N1625, N1616);
xor XOR2 (N1626, N1618, N995);
or OR2 (N1627, N1621, N1274);
buf BUF1 (N1628, N1625);
xor XOR2 (N1629, N1624, N59);
xor XOR2 (N1630, N1628, N365);
nand NAND3 (N1631, N1630, N766, N447);
or OR3 (N1632, N1627, N15, N1423);
not NOT1 (N1633, N1596);
or OR3 (N1634, N1622, N1092, N30);
not NOT1 (N1635, N1634);
or OR4 (N1636, N1632, N1005, N838, N435);
xor XOR2 (N1637, N1633, N1580);
not NOT1 (N1638, N648);
not NOT1 (N1639, N1637);
not NOT1 (N1640, N1639);
nor NOR2 (N1641, N1638, N1002);
nand NAND3 (N1642, N1606, N482, N173);
nor NOR3 (N1643, N1635, N108, N179);
not NOT1 (N1644, N1640);
buf BUF1 (N1645, N1636);
nand NAND3 (N1646, N1629, N423, N1615);
or OR3 (N1647, N1646, N338, N573);
buf BUF1 (N1648, N1642);
buf BUF1 (N1649, N1648);
nand NAND2 (N1650, N1631, N1636);
or OR4 (N1651, N1649, N923, N1615, N1094);
not NOT1 (N1652, N1643);
not NOT1 (N1653, N1626);
nand NAND2 (N1654, N1641, N476);
nor NOR2 (N1655, N1620, N603);
nand NAND2 (N1656, N1653, N1622);
xor XOR2 (N1657, N1647, N35);
nor NOR2 (N1658, N1623, N1641);
nor NOR3 (N1659, N1655, N319, N790);
and AND2 (N1660, N1657, N85);
buf BUF1 (N1661, N1660);
nor NOR4 (N1662, N1661, N67, N831, N476);
xor XOR2 (N1663, N1645, N1294);
buf BUF1 (N1664, N1662);
or OR3 (N1665, N1651, N709, N1309);
nor NOR2 (N1666, N1652, N1565);
buf BUF1 (N1667, N1663);
nand NAND4 (N1668, N1656, N683, N1229, N1180);
or OR4 (N1669, N1668, N192, N616, N1568);
xor XOR2 (N1670, N1644, N1413);
not NOT1 (N1671, N1659);
or OR2 (N1672, N1658, N1649);
xor XOR2 (N1673, N1667, N238);
xor XOR2 (N1674, N1672, N805);
and AND2 (N1675, N1664, N1522);
nand NAND2 (N1676, N1654, N75);
nor NOR3 (N1677, N1650, N145, N1235);
not NOT1 (N1678, N1675);
nor NOR4 (N1679, N1678, N532, N1231, N1378);
xor XOR2 (N1680, N1670, N566);
buf BUF1 (N1681, N1676);
xor XOR2 (N1682, N1680, N1285);
nor NOR3 (N1683, N1665, N1194, N679);
xor XOR2 (N1684, N1681, N1366);
not NOT1 (N1685, N1669);
and AND4 (N1686, N1684, N1379, N1609, N1046);
not NOT1 (N1687, N1671);
buf BUF1 (N1688, N1687);
not NOT1 (N1689, N1666);
not NOT1 (N1690, N1679);
buf BUF1 (N1691, N1677);
and AND2 (N1692, N1685, N539);
or OR2 (N1693, N1673, N1376);
not NOT1 (N1694, N1690);
or OR4 (N1695, N1693, N1428, N253, N141);
xor XOR2 (N1696, N1683, N24);
xor XOR2 (N1697, N1674, N324);
buf BUF1 (N1698, N1696);
nand NAND4 (N1699, N1686, N1520, N1672, N840);
not NOT1 (N1700, N1692);
nor NOR2 (N1701, N1689, N484);
or OR3 (N1702, N1691, N1178, N362);
or OR4 (N1703, N1699, N564, N313, N1580);
xor XOR2 (N1704, N1688, N1164);
nand NAND2 (N1705, N1682, N1693);
or OR2 (N1706, N1705, N529);
or OR2 (N1707, N1702, N1226);
buf BUF1 (N1708, N1700);
and AND3 (N1709, N1708, N97, N319);
and AND2 (N1710, N1694, N1669);
not NOT1 (N1711, N1706);
not NOT1 (N1712, N1711);
nor NOR4 (N1713, N1707, N1653, N923, N1694);
nor NOR3 (N1714, N1704, N157, N466);
buf BUF1 (N1715, N1712);
nand NAND2 (N1716, N1709, N900);
nor NOR3 (N1717, N1697, N511, N1505);
nand NAND2 (N1718, N1716, N1020);
buf BUF1 (N1719, N1698);
not NOT1 (N1720, N1703);
buf BUF1 (N1721, N1717);
nor NOR4 (N1722, N1710, N381, N802, N930);
nand NAND3 (N1723, N1720, N1246, N131);
or OR2 (N1724, N1719, N346);
nand NAND3 (N1725, N1718, N1635, N158);
buf BUF1 (N1726, N1715);
nor NOR2 (N1727, N1726, N989);
nor NOR4 (N1728, N1714, N505, N1245, N940);
nand NAND4 (N1729, N1725, N381, N1146, N370);
and AND3 (N1730, N1713, N1519, N11);
and AND3 (N1731, N1730, N264, N922);
nand NAND3 (N1732, N1724, N497, N304);
nand NAND4 (N1733, N1727, N1347, N811, N462);
and AND4 (N1734, N1723, N160, N202, N436);
buf BUF1 (N1735, N1729);
xor XOR2 (N1736, N1701, N920);
and AND3 (N1737, N1728, N197, N703);
not NOT1 (N1738, N1721);
and AND2 (N1739, N1731, N232);
buf BUF1 (N1740, N1695);
xor XOR2 (N1741, N1734, N1446);
buf BUF1 (N1742, N1739);
nand NAND3 (N1743, N1738, N797, N1575);
not NOT1 (N1744, N1741);
or OR4 (N1745, N1733, N1261, N1009, N576);
nor NOR2 (N1746, N1737, N1268);
buf BUF1 (N1747, N1743);
nor NOR3 (N1748, N1722, N896, N90);
and AND4 (N1749, N1746, N1412, N708, N260);
buf BUF1 (N1750, N1740);
xor XOR2 (N1751, N1735, N894);
buf BUF1 (N1752, N1736);
nor NOR4 (N1753, N1744, N579, N1394, N451);
or OR4 (N1754, N1745, N629, N1376, N1471);
nor NOR3 (N1755, N1752, N1420, N1736);
or OR4 (N1756, N1750, N1472, N420, N1050);
and AND2 (N1757, N1732, N1118);
and AND3 (N1758, N1747, N1567, N556);
or OR2 (N1759, N1748, N968);
xor XOR2 (N1760, N1742, N629);
nor NOR2 (N1761, N1756, N91);
and AND4 (N1762, N1749, N1434, N249, N1016);
or OR2 (N1763, N1760, N712);
and AND2 (N1764, N1758, N1486);
or OR2 (N1765, N1761, N1096);
nor NOR4 (N1766, N1763, N88, N313, N1490);
or OR4 (N1767, N1759, N855, N1137, N59);
or OR3 (N1768, N1762, N1493, N1241);
not NOT1 (N1769, N1768);
and AND4 (N1770, N1764, N111, N613, N742);
not NOT1 (N1771, N1766);
xor XOR2 (N1772, N1765, N531);
xor XOR2 (N1773, N1772, N927);
buf BUF1 (N1774, N1757);
buf BUF1 (N1775, N1774);
xor XOR2 (N1776, N1775, N811);
not NOT1 (N1777, N1767);
xor XOR2 (N1778, N1751, N606);
not NOT1 (N1779, N1754);
or OR3 (N1780, N1753, N1169, N1018);
buf BUF1 (N1781, N1780);
nor NOR4 (N1782, N1769, N707, N65, N107);
buf BUF1 (N1783, N1778);
xor XOR2 (N1784, N1755, N997);
buf BUF1 (N1785, N1783);
and AND4 (N1786, N1770, N1515, N121, N439);
nand NAND2 (N1787, N1784, N258);
buf BUF1 (N1788, N1785);
not NOT1 (N1789, N1776);
xor XOR2 (N1790, N1777, N740);
nand NAND4 (N1791, N1788, N1296, N642, N776);
not NOT1 (N1792, N1781);
and AND3 (N1793, N1782, N1183, N636);
not NOT1 (N1794, N1787);
buf BUF1 (N1795, N1773);
not NOT1 (N1796, N1786);
or OR2 (N1797, N1779, N972);
nand NAND3 (N1798, N1789, N1530, N380);
not NOT1 (N1799, N1791);
nand NAND3 (N1800, N1797, N950, N1779);
not NOT1 (N1801, N1796);
and AND4 (N1802, N1801, N1533, N563, N1743);
or OR2 (N1803, N1792, N1078);
nor NOR4 (N1804, N1799, N1791, N1791, N237);
or OR4 (N1805, N1771, N1544, N20, N1306);
xor XOR2 (N1806, N1800, N1130);
not NOT1 (N1807, N1806);
not NOT1 (N1808, N1798);
not NOT1 (N1809, N1807);
buf BUF1 (N1810, N1802);
nor NOR2 (N1811, N1795, N386);
not NOT1 (N1812, N1805);
and AND3 (N1813, N1793, N577, N327);
xor XOR2 (N1814, N1790, N807);
nor NOR2 (N1815, N1810, N1301);
nand NAND4 (N1816, N1813, N1505, N1271, N333);
xor XOR2 (N1817, N1811, N1416);
xor XOR2 (N1818, N1804, N886);
nand NAND3 (N1819, N1808, N130, N878);
xor XOR2 (N1820, N1817, N1263);
and AND4 (N1821, N1816, N1546, N764, N1155);
buf BUF1 (N1822, N1815);
nand NAND4 (N1823, N1819, N140, N818, N651);
and AND4 (N1824, N1803, N1122, N883, N1531);
and AND3 (N1825, N1823, N1089, N1546);
and AND2 (N1826, N1794, N1074);
not NOT1 (N1827, N1825);
and AND4 (N1828, N1822, N689, N1751, N73);
or OR3 (N1829, N1827, N780, N320);
nand NAND4 (N1830, N1814, N1794, N942, N1399);
not NOT1 (N1831, N1829);
nor NOR4 (N1832, N1821, N316, N986, N1229);
and AND4 (N1833, N1824, N1120, N488, N924);
nor NOR4 (N1834, N1831, N1234, N1286, N845);
nand NAND2 (N1835, N1834, N241);
buf BUF1 (N1836, N1833);
buf BUF1 (N1837, N1828);
or OR4 (N1838, N1836, N408, N502, N602);
buf BUF1 (N1839, N1818);
xor XOR2 (N1840, N1809, N403);
nand NAND3 (N1841, N1840, N1741, N991);
not NOT1 (N1842, N1837);
buf BUF1 (N1843, N1841);
not NOT1 (N1844, N1843);
and AND3 (N1845, N1838, N1633, N1192);
xor XOR2 (N1846, N1830, N169);
not NOT1 (N1847, N1835);
and AND3 (N1848, N1845, N790, N1562);
buf BUF1 (N1849, N1820);
not NOT1 (N1850, N1844);
xor XOR2 (N1851, N1847, N1383);
buf BUF1 (N1852, N1839);
nor NOR4 (N1853, N1812, N1636, N12, N841);
or OR4 (N1854, N1853, N339, N1541, N1552);
not NOT1 (N1855, N1846);
nor NOR2 (N1856, N1851, N622);
not NOT1 (N1857, N1852);
buf BUF1 (N1858, N1849);
not NOT1 (N1859, N1826);
nor NOR2 (N1860, N1858, N1176);
not NOT1 (N1861, N1848);
xor XOR2 (N1862, N1842, N29);
buf BUF1 (N1863, N1857);
not NOT1 (N1864, N1855);
xor XOR2 (N1865, N1864, N1135);
nand NAND4 (N1866, N1860, N1808, N1421, N1029);
nand NAND3 (N1867, N1850, N1426, N18);
not NOT1 (N1868, N1866);
and AND4 (N1869, N1863, N1821, N1773, N1823);
buf BUF1 (N1870, N1869);
xor XOR2 (N1871, N1854, N608);
nor NOR2 (N1872, N1868, N496);
and AND3 (N1873, N1862, N420, N1275);
not NOT1 (N1874, N1856);
nand NAND4 (N1875, N1870, N1218, N668, N1115);
and AND3 (N1876, N1865, N817, N724);
and AND2 (N1877, N1861, N1654);
xor XOR2 (N1878, N1859, N1556);
nand NAND3 (N1879, N1867, N1192, N18);
nor NOR4 (N1880, N1879, N572, N74, N1560);
or OR2 (N1881, N1878, N1575);
not NOT1 (N1882, N1880);
nand NAND2 (N1883, N1876, N472);
nor NOR3 (N1884, N1872, N1265, N1541);
nand NAND2 (N1885, N1883, N481);
buf BUF1 (N1886, N1873);
and AND4 (N1887, N1875, N249, N981, N428);
not NOT1 (N1888, N1882);
nand NAND4 (N1889, N1884, N866, N87, N71);
and AND4 (N1890, N1832, N1024, N495, N964);
buf BUF1 (N1891, N1888);
and AND3 (N1892, N1886, N1350, N135);
nor NOR2 (N1893, N1892, N636);
and AND2 (N1894, N1874, N469);
buf BUF1 (N1895, N1885);
nand NAND3 (N1896, N1887, N1868, N786);
not NOT1 (N1897, N1871);
xor XOR2 (N1898, N1894, N501);
not NOT1 (N1899, N1895);
xor XOR2 (N1900, N1896, N1718);
xor XOR2 (N1901, N1881, N1397);
nand NAND3 (N1902, N1898, N1878, N1479);
and AND3 (N1903, N1899, N602, N492);
xor XOR2 (N1904, N1893, N1469);
nor NOR2 (N1905, N1900, N1129);
nand NAND4 (N1906, N1903, N1850, N25, N82);
buf BUF1 (N1907, N1901);
not NOT1 (N1908, N1906);
not NOT1 (N1909, N1891);
xor XOR2 (N1910, N1908, N1634);
buf BUF1 (N1911, N1905);
buf BUF1 (N1912, N1904);
xor XOR2 (N1913, N1909, N238);
nor NOR3 (N1914, N1913, N392, N1659);
xor XOR2 (N1915, N1911, N1611);
xor XOR2 (N1916, N1915, N1898);
and AND2 (N1917, N1912, N1445);
or OR2 (N1918, N1916, N243);
and AND2 (N1919, N1914, N1126);
nor NOR4 (N1920, N1897, N27, N1366, N878);
or OR4 (N1921, N1889, N1517, N427, N1797);
buf BUF1 (N1922, N1877);
and AND2 (N1923, N1917, N1225);
buf BUF1 (N1924, N1910);
nand NAND4 (N1925, N1921, N984, N1055, N469);
not NOT1 (N1926, N1923);
xor XOR2 (N1927, N1924, N883);
xor XOR2 (N1928, N1922, N1802);
nor NOR2 (N1929, N1902, N1559);
and AND2 (N1930, N1907, N1703);
xor XOR2 (N1931, N1919, N1045);
not NOT1 (N1932, N1930);
buf BUF1 (N1933, N1890);
and AND2 (N1934, N1933, N1399);
xor XOR2 (N1935, N1920, N1006);
and AND3 (N1936, N1926, N299, N915);
nor NOR3 (N1937, N1929, N206, N900);
xor XOR2 (N1938, N1936, N1159);
nand NAND3 (N1939, N1931, N1245, N800);
or OR2 (N1940, N1928, N1385);
nand NAND2 (N1941, N1918, N605);
buf BUF1 (N1942, N1925);
nand NAND3 (N1943, N1939, N1315, N1717);
and AND2 (N1944, N1935, N1626);
not NOT1 (N1945, N1944);
or OR3 (N1946, N1945, N1572, N1382);
xor XOR2 (N1947, N1927, N1691);
not NOT1 (N1948, N1937);
or OR2 (N1949, N1932, N244);
not NOT1 (N1950, N1941);
xor XOR2 (N1951, N1949, N62);
nand NAND3 (N1952, N1938, N349, N770);
nand NAND3 (N1953, N1943, N1572, N973);
nor NOR4 (N1954, N1934, N1168, N931, N489);
and AND2 (N1955, N1942, N592);
xor XOR2 (N1956, N1955, N519);
nand NAND2 (N1957, N1952, N1478);
nand NAND3 (N1958, N1957, N781, N46);
not NOT1 (N1959, N1950);
not NOT1 (N1960, N1959);
buf BUF1 (N1961, N1946);
xor XOR2 (N1962, N1948, N1426);
buf BUF1 (N1963, N1947);
xor XOR2 (N1964, N1958, N86);
not NOT1 (N1965, N1956);
nand NAND4 (N1966, N1962, N844, N1624, N872);
not NOT1 (N1967, N1963);
or OR4 (N1968, N1965, N793, N1134, N1029);
xor XOR2 (N1969, N1951, N409);
and AND3 (N1970, N1953, N392, N467);
buf BUF1 (N1971, N1967);
not NOT1 (N1972, N1961);
nor NOR3 (N1973, N1968, N585, N391);
not NOT1 (N1974, N1973);
and AND2 (N1975, N1970, N1931);
nor NOR4 (N1976, N1940, N1622, N574, N731);
nor NOR2 (N1977, N1954, N998);
or OR3 (N1978, N1975, N1243, N876);
not NOT1 (N1979, N1969);
not NOT1 (N1980, N1977);
and AND3 (N1981, N1978, N1888, N1854);
not NOT1 (N1982, N1966);
buf BUF1 (N1983, N1981);
and AND2 (N1984, N1960, N566);
buf BUF1 (N1985, N1972);
xor XOR2 (N1986, N1982, N260);
and AND4 (N1987, N1984, N521, N781, N308);
and AND2 (N1988, N1985, N1838);
or OR4 (N1989, N1983, N1984, N1484, N1103);
xor XOR2 (N1990, N1987, N1950);
xor XOR2 (N1991, N1989, N173);
and AND3 (N1992, N1980, N1990, N252);
xor XOR2 (N1993, N709, N1579);
nand NAND3 (N1994, N1964, N1344, N393);
nor NOR3 (N1995, N1986, N776, N1293);
not NOT1 (N1996, N1994);
and AND3 (N1997, N1995, N735, N663);
not NOT1 (N1998, N1979);
and AND4 (N1999, N1976, N1798, N1472, N1295);
and AND4 (N2000, N1988, N251, N182, N51);
and AND2 (N2001, N1992, N16);
or OR4 (N2002, N1997, N80, N709, N460);
not NOT1 (N2003, N1974);
and AND3 (N2004, N1998, N264, N831);
or OR4 (N2005, N2002, N1404, N1578, N792);
not NOT1 (N2006, N1999);
nand NAND3 (N2007, N2001, N1043, N423);
or OR3 (N2008, N1991, N543, N597);
not NOT1 (N2009, N2003);
or OR2 (N2010, N2007, N1412);
buf BUF1 (N2011, N2010);
xor XOR2 (N2012, N1996, N1756);
xor XOR2 (N2013, N2000, N457);
not NOT1 (N2014, N2004);
xor XOR2 (N2015, N1971, N346);
nand NAND4 (N2016, N2008, N243, N124, N301);
or OR2 (N2017, N2014, N876);
buf BUF1 (N2018, N2012);
buf BUF1 (N2019, N2013);
or OR2 (N2020, N2005, N1221);
nor NOR3 (N2021, N2006, N514, N286);
and AND4 (N2022, N2009, N928, N1152, N1848);
nor NOR3 (N2023, N2020, N1424, N1173);
xor XOR2 (N2024, N2022, N1820);
xor XOR2 (N2025, N2023, N577);
and AND2 (N2026, N2024, N798);
not NOT1 (N2027, N2025);
and AND2 (N2028, N2018, N838);
and AND2 (N2029, N2026, N394);
or OR4 (N2030, N2016, N1775, N1582, N490);
or OR4 (N2031, N2029, N1994, N1667, N588);
or OR3 (N2032, N1993, N1727, N825);
xor XOR2 (N2033, N2032, N1134);
and AND2 (N2034, N2030, N796);
xor XOR2 (N2035, N2031, N1469);
nand NAND4 (N2036, N2019, N601, N423, N1505);
nand NAND4 (N2037, N2027, N1676, N380, N660);
not NOT1 (N2038, N2034);
nand NAND2 (N2039, N2021, N1960);
or OR3 (N2040, N2015, N1430, N1038);
buf BUF1 (N2041, N2038);
or OR4 (N2042, N2041, N693, N75, N1419);
nor NOR2 (N2043, N2017, N1324);
or OR2 (N2044, N2039, N465);
nor NOR2 (N2045, N2035, N142);
and AND4 (N2046, N2011, N332, N595, N434);
or OR4 (N2047, N2042, N397, N780, N1553);
not NOT1 (N2048, N2043);
or OR2 (N2049, N2028, N834);
nand NAND2 (N2050, N2040, N138);
xor XOR2 (N2051, N2047, N263);
nor NOR2 (N2052, N2049, N1665);
and AND3 (N2053, N2033, N1639, N479);
xor XOR2 (N2054, N2036, N860);
not NOT1 (N2055, N2054);
buf BUF1 (N2056, N2046);
nor NOR2 (N2057, N2050, N686);
or OR4 (N2058, N2051, N1696, N1315, N1504);
or OR3 (N2059, N2044, N321, N1453);
not NOT1 (N2060, N2056);
nor NOR4 (N2061, N2058, N1580, N1073, N1737);
buf BUF1 (N2062, N2057);
or OR2 (N2063, N2053, N1766);
buf BUF1 (N2064, N2055);
buf BUF1 (N2065, N2061);
not NOT1 (N2066, N2048);
or OR4 (N2067, N2052, N1746, N652, N41);
not NOT1 (N2068, N2067);
nor NOR2 (N2069, N2037, N2045);
buf BUF1 (N2070, N501);
and AND2 (N2071, N2059, N1509);
xor XOR2 (N2072, N2068, N1789);
buf BUF1 (N2073, N2062);
or OR3 (N2074, N2071, N1423, N286);
xor XOR2 (N2075, N2063, N1103);
nor NOR2 (N2076, N2070, N822);
or OR3 (N2077, N2065, N1754, N1347);
xor XOR2 (N2078, N2069, N203);
not NOT1 (N2079, N2077);
and AND4 (N2080, N2076, N1067, N992, N190);
not NOT1 (N2081, N2080);
and AND2 (N2082, N2078, N938);
xor XOR2 (N2083, N2073, N94);
or OR3 (N2084, N2075, N2009, N678);
nor NOR3 (N2085, N2082, N1420, N1630);
buf BUF1 (N2086, N2060);
nand NAND4 (N2087, N2072, N1591, N1217, N623);
or OR3 (N2088, N2084, N939, N1109);
or OR2 (N2089, N2079, N665);
and AND2 (N2090, N2088, N1231);
buf BUF1 (N2091, N2081);
or OR3 (N2092, N2066, N1297, N298);
nand NAND4 (N2093, N2091, N1231, N1868, N503);
xor XOR2 (N2094, N2083, N1640);
buf BUF1 (N2095, N2092);
buf BUF1 (N2096, N2095);
nor NOR4 (N2097, N2085, N1951, N835, N1361);
and AND4 (N2098, N2087, N1709, N894, N312);
xor XOR2 (N2099, N2074, N233);
and AND2 (N2100, N2098, N1397);
or OR3 (N2101, N2094, N1098, N973);
not NOT1 (N2102, N2064);
and AND3 (N2103, N2086, N1638, N982);
xor XOR2 (N2104, N2096, N57);
buf BUF1 (N2105, N2093);
xor XOR2 (N2106, N2099, N1707);
or OR2 (N2107, N2089, N863);
nor NOR4 (N2108, N2102, N559, N408, N1947);
buf BUF1 (N2109, N2108);
not NOT1 (N2110, N2109);
or OR4 (N2111, N2107, N2032, N910, N1434);
buf BUF1 (N2112, N2105);
xor XOR2 (N2113, N2110, N204);
not NOT1 (N2114, N2106);
nand NAND4 (N2115, N2103, N337, N859, N1500);
nor NOR2 (N2116, N2113, N35);
nand NAND4 (N2117, N2100, N407, N496, N217);
nor NOR4 (N2118, N2090, N931, N664, N2113);
or OR4 (N2119, N2111, N2103, N416, N1430);
not NOT1 (N2120, N2104);
and AND4 (N2121, N2116, N271, N204, N1856);
nand NAND4 (N2122, N2119, N1427, N1448, N1098);
nor NOR3 (N2123, N2118, N635, N902);
buf BUF1 (N2124, N2101);
or OR3 (N2125, N2122, N2100, N152);
and AND2 (N2126, N2120, N2063);
not NOT1 (N2127, N2125);
not NOT1 (N2128, N2097);
nand NAND4 (N2129, N2115, N762, N951, N686);
xor XOR2 (N2130, N2129, N843);
nor NOR3 (N2131, N2127, N596, N1450);
nand NAND4 (N2132, N2114, N1769, N588, N2048);
or OR3 (N2133, N2130, N1539, N1754);
or OR4 (N2134, N2126, N1945, N550, N1399);
or OR4 (N2135, N2124, N1003, N1532, N1772);
xor XOR2 (N2136, N2135, N2124);
nor NOR3 (N2137, N2134, N750, N210);
buf BUF1 (N2138, N2128);
nand NAND4 (N2139, N2112, N2110, N1431, N679);
nor NOR2 (N2140, N2138, N1168);
nand NAND4 (N2141, N2132, N157, N1943, N1493);
nor NOR4 (N2142, N2123, N377, N511, N1117);
nand NAND2 (N2143, N2131, N777);
and AND3 (N2144, N2117, N1246, N639);
and AND4 (N2145, N2137, N2100, N967, N1946);
xor XOR2 (N2146, N2139, N330);
buf BUF1 (N2147, N2146);
nand NAND2 (N2148, N2147, N1592);
or OR4 (N2149, N2144, N439, N2016, N1872);
xor XOR2 (N2150, N2148, N733);
not NOT1 (N2151, N2121);
nor NOR4 (N2152, N2151, N174, N1367, N727);
nand NAND4 (N2153, N2143, N589, N1833, N827);
not NOT1 (N2154, N2141);
nand NAND3 (N2155, N2142, N2132, N1084);
and AND2 (N2156, N2133, N2065);
or OR3 (N2157, N2140, N1257, N1045);
not NOT1 (N2158, N2157);
and AND3 (N2159, N2153, N1509, N206);
xor XOR2 (N2160, N2136, N411);
not NOT1 (N2161, N2145);
nor NOR2 (N2162, N2161, N1169);
nor NOR2 (N2163, N2162, N1366);
or OR3 (N2164, N2152, N1970, N294);
xor XOR2 (N2165, N2159, N431);
not NOT1 (N2166, N2158);
buf BUF1 (N2167, N2160);
or OR3 (N2168, N2150, N2018, N687);
xor XOR2 (N2169, N2149, N1104);
buf BUF1 (N2170, N2155);
nand NAND4 (N2171, N2165, N1386, N370, N1708);
buf BUF1 (N2172, N2164);
nand NAND4 (N2173, N2167, N526, N1211, N1368);
and AND2 (N2174, N2169, N777);
nor NOR2 (N2175, N2156, N1907);
and AND3 (N2176, N2154, N2137, N652);
or OR3 (N2177, N2171, N900, N1973);
buf BUF1 (N2178, N2170);
nand NAND2 (N2179, N2178, N1574);
buf BUF1 (N2180, N2173);
nor NOR2 (N2181, N2163, N866);
not NOT1 (N2182, N2168);
or OR4 (N2183, N2166, N124, N646, N700);
xor XOR2 (N2184, N2181, N1530);
buf BUF1 (N2185, N2183);
or OR2 (N2186, N2184, N1100);
nand NAND4 (N2187, N2176, N725, N383, N451);
buf BUF1 (N2188, N2186);
nor NOR3 (N2189, N2187, N1006, N665);
or OR2 (N2190, N2189, N596);
or OR4 (N2191, N2174, N177, N1988, N34);
buf BUF1 (N2192, N2177);
or OR4 (N2193, N2192, N1408, N520, N1562);
xor XOR2 (N2194, N2190, N394);
buf BUF1 (N2195, N2193);
or OR4 (N2196, N2180, N204, N490, N906);
nand NAND3 (N2197, N2175, N1334, N1474);
buf BUF1 (N2198, N2188);
nor NOR3 (N2199, N2182, N1970, N1235);
buf BUF1 (N2200, N2194);
nand NAND4 (N2201, N2197, N476, N1355, N1358);
not NOT1 (N2202, N2196);
not NOT1 (N2203, N2191);
or OR3 (N2204, N2203, N930, N1372);
and AND2 (N2205, N2204, N790);
nand NAND2 (N2206, N2198, N2032);
nand NAND4 (N2207, N2202, N357, N996, N846);
buf BUF1 (N2208, N2179);
not NOT1 (N2209, N2205);
nand NAND2 (N2210, N2185, N1778);
or OR3 (N2211, N2199, N1923, N553);
and AND3 (N2212, N2200, N1702, N1080);
or OR4 (N2213, N2195, N885, N1911, N1027);
buf BUF1 (N2214, N2213);
not NOT1 (N2215, N2211);
xor XOR2 (N2216, N2215, N832);
nand NAND4 (N2217, N2201, N136, N1005, N284);
or OR2 (N2218, N2210, N1032);
xor XOR2 (N2219, N2207, N425);
not NOT1 (N2220, N2216);
nand NAND4 (N2221, N2220, N130, N1243, N751);
buf BUF1 (N2222, N2221);
nand NAND2 (N2223, N2206, N94);
and AND2 (N2224, N2223, N945);
nand NAND2 (N2225, N2218, N682);
and AND2 (N2226, N2208, N1174);
xor XOR2 (N2227, N2225, N619);
not NOT1 (N2228, N2224);
not NOT1 (N2229, N2212);
or OR3 (N2230, N2229, N686, N1389);
buf BUF1 (N2231, N2222);
or OR3 (N2232, N2226, N1613, N1277);
buf BUF1 (N2233, N2230);
and AND2 (N2234, N2214, N1970);
or OR4 (N2235, N2232, N1883, N804, N642);
nor NOR4 (N2236, N2235, N1069, N943, N416);
not NOT1 (N2237, N2209);
nor NOR4 (N2238, N2219, N1751, N805, N494);
not NOT1 (N2239, N2234);
xor XOR2 (N2240, N2228, N1273);
not NOT1 (N2241, N2238);
nand NAND2 (N2242, N2237, N650);
xor XOR2 (N2243, N2227, N833);
and AND4 (N2244, N2241, N636, N921, N597);
nand NAND4 (N2245, N2242, N1354, N791, N1178);
not NOT1 (N2246, N2217);
buf BUF1 (N2247, N2239);
nor NOR3 (N2248, N2236, N1097, N1784);
and AND2 (N2249, N2233, N1126);
nor NOR4 (N2250, N2240, N1355, N1950, N680);
nor NOR2 (N2251, N2244, N518);
nor NOR4 (N2252, N2250, N1007, N418, N59);
nor NOR2 (N2253, N2252, N363);
or OR4 (N2254, N2251, N2244, N770, N1170);
buf BUF1 (N2255, N2254);
or OR2 (N2256, N2231, N2039);
xor XOR2 (N2257, N2256, N858);
nand NAND3 (N2258, N2246, N1568, N1573);
nor NOR3 (N2259, N2247, N1872, N751);
and AND2 (N2260, N2249, N2097);
nor NOR2 (N2261, N2260, N764);
not NOT1 (N2262, N2253);
and AND4 (N2263, N2248, N903, N1351, N1302);
nand NAND2 (N2264, N2255, N2240);
xor XOR2 (N2265, N2259, N1531);
or OR4 (N2266, N2264, N672, N364, N103);
nand NAND2 (N2267, N2262, N1204);
buf BUF1 (N2268, N2267);
nand NAND2 (N2269, N2266, N1082);
not NOT1 (N2270, N2268);
nor NOR2 (N2271, N2263, N1934);
nand NAND4 (N2272, N2261, N1369, N73, N985);
or OR2 (N2273, N2243, N124);
not NOT1 (N2274, N2265);
buf BUF1 (N2275, N2272);
and AND2 (N2276, N2245, N1511);
nor NOR4 (N2277, N2276, N2070, N350, N1247);
nand NAND4 (N2278, N2273, N1384, N1922, N80);
and AND2 (N2279, N2258, N1008);
nand NAND2 (N2280, N2269, N1628);
buf BUF1 (N2281, N2280);
xor XOR2 (N2282, N2271, N1999);
not NOT1 (N2283, N2274);
or OR4 (N2284, N2257, N147, N1113, N239);
nand NAND3 (N2285, N2284, N1673, N2253);
xor XOR2 (N2286, N2282, N1534);
nand NAND4 (N2287, N2283, N1537, N2148, N114);
nand NAND3 (N2288, N2281, N848, N2267);
buf BUF1 (N2289, N2285);
buf BUF1 (N2290, N2289);
and AND4 (N2291, N2288, N283, N361, N2215);
or OR4 (N2292, N2279, N535, N2089, N158);
and AND4 (N2293, N2286, N2088, N146, N279);
xor XOR2 (N2294, N2293, N2228);
and AND3 (N2295, N2278, N2226, N592);
buf BUF1 (N2296, N2291);
xor XOR2 (N2297, N2277, N1397);
not NOT1 (N2298, N2290);
not NOT1 (N2299, N2297);
xor XOR2 (N2300, N2294, N646);
and AND4 (N2301, N2292, N1745, N736, N1202);
buf BUF1 (N2302, N2301);
xor XOR2 (N2303, N2296, N391);
xor XOR2 (N2304, N2300, N2146);
xor XOR2 (N2305, N2295, N1677);
and AND2 (N2306, N2299, N1456);
and AND4 (N2307, N2302, N964, N361, N797);
nor NOR4 (N2308, N2304, N2111, N734, N3);
not NOT1 (N2309, N2307);
not NOT1 (N2310, N2270);
or OR3 (N2311, N2308, N1014, N151);
nand NAND4 (N2312, N2311, N293, N994, N1625);
nor NOR3 (N2313, N2306, N2280, N1959);
buf BUF1 (N2314, N2305);
and AND2 (N2315, N2313, N2223);
and AND3 (N2316, N2303, N913, N1518);
xor XOR2 (N2317, N2275, N1565);
and AND3 (N2318, N2172, N180, N883);
and AND3 (N2319, N2314, N1177, N2118);
nand NAND3 (N2320, N2298, N213, N1093);
nor NOR4 (N2321, N2320, N2224, N1167, N1419);
xor XOR2 (N2322, N2321, N500);
or OR3 (N2323, N2287, N1161, N1942);
and AND2 (N2324, N2318, N1953);
not NOT1 (N2325, N2323);
and AND2 (N2326, N2322, N1339);
nand NAND2 (N2327, N2326, N95);
nand NAND4 (N2328, N2325, N118, N904, N2087);
not NOT1 (N2329, N2319);
not NOT1 (N2330, N2312);
nand NAND4 (N2331, N2324, N235, N191, N1485);
xor XOR2 (N2332, N2327, N122);
nor NOR3 (N2333, N2310, N1352, N467);
buf BUF1 (N2334, N2316);
nor NOR2 (N2335, N2331, N1948);
xor XOR2 (N2336, N2332, N266);
nand NAND2 (N2337, N2333, N1136);
buf BUF1 (N2338, N2335);
or OR3 (N2339, N2328, N316, N44);
nand NAND2 (N2340, N2334, N1784);
xor XOR2 (N2341, N2336, N1455);
nor NOR3 (N2342, N2330, N567, N1665);
or OR2 (N2343, N2329, N1100);
and AND3 (N2344, N2317, N1718, N1269);
nand NAND3 (N2345, N2339, N1451, N249);
and AND4 (N2346, N2337, N327, N306, N129);
not NOT1 (N2347, N2309);
xor XOR2 (N2348, N2342, N24);
or OR4 (N2349, N2315, N1343, N911, N1239);
nand NAND2 (N2350, N2345, N1583);
buf BUF1 (N2351, N2346);
buf BUF1 (N2352, N2341);
nor NOR4 (N2353, N2350, N1576, N1582, N1782);
nor NOR2 (N2354, N2340, N615);
xor XOR2 (N2355, N2353, N1576);
xor XOR2 (N2356, N2349, N2253);
and AND4 (N2357, N2347, N1786, N925, N854);
nand NAND3 (N2358, N2348, N2141, N1586);
not NOT1 (N2359, N2355);
not NOT1 (N2360, N2351);
nor NOR3 (N2361, N2343, N2178, N186);
nand NAND4 (N2362, N2338, N2243, N1386, N843);
not NOT1 (N2363, N2352);
not NOT1 (N2364, N2357);
or OR4 (N2365, N2360, N571, N533, N1042);
or OR4 (N2366, N2362, N1516, N573, N1214);
xor XOR2 (N2367, N2359, N765);
xor XOR2 (N2368, N2363, N482);
not NOT1 (N2369, N2367);
or OR2 (N2370, N2369, N65);
buf BUF1 (N2371, N2361);
and AND2 (N2372, N2365, N2065);
nand NAND3 (N2373, N2371, N64, N1885);
buf BUF1 (N2374, N2373);
buf BUF1 (N2375, N2366);
buf BUF1 (N2376, N2356);
xor XOR2 (N2377, N2344, N4);
xor XOR2 (N2378, N2364, N372);
buf BUF1 (N2379, N2372);
buf BUF1 (N2380, N2368);
and AND3 (N2381, N2379, N901, N2197);
and AND4 (N2382, N2376, N1818, N2174, N2238);
xor XOR2 (N2383, N2374, N2204);
nor NOR3 (N2384, N2381, N1807, N253);
xor XOR2 (N2385, N2382, N1307);
nor NOR2 (N2386, N2377, N2124);
xor XOR2 (N2387, N2354, N100);
or OR4 (N2388, N2383, N741, N2074, N2286);
not NOT1 (N2389, N2370);
nand NAND2 (N2390, N2387, N382);
and AND3 (N2391, N2389, N329, N972);
not NOT1 (N2392, N2378);
xor XOR2 (N2393, N2358, N1635);
nor NOR3 (N2394, N2385, N1295, N193);
nand NAND2 (N2395, N2375, N1374);
xor XOR2 (N2396, N2380, N1141);
nor NOR4 (N2397, N2390, N2305, N1296, N1027);
xor XOR2 (N2398, N2396, N334);
nand NAND2 (N2399, N2394, N731);
and AND2 (N2400, N2388, N740);
or OR2 (N2401, N2393, N1765);
buf BUF1 (N2402, N2386);
nand NAND2 (N2403, N2391, N1579);
nor NOR3 (N2404, N2403, N2204, N50);
xor XOR2 (N2405, N2400, N737);
nand NAND3 (N2406, N2397, N372, N624);
nand NAND4 (N2407, N2395, N2241, N2252, N1787);
not NOT1 (N2408, N2399);
buf BUF1 (N2409, N2402);
xor XOR2 (N2410, N2405, N734);
or OR2 (N2411, N2409, N1504);
buf BUF1 (N2412, N2401);
buf BUF1 (N2413, N2392);
not NOT1 (N2414, N2384);
or OR3 (N2415, N2398, N739, N920);
nand NAND3 (N2416, N2415, N2234, N2052);
and AND3 (N2417, N2413, N688, N1193);
and AND3 (N2418, N2410, N1339, N1843);
or OR3 (N2419, N2406, N2325, N234);
xor XOR2 (N2420, N2416, N689);
nor NOR2 (N2421, N2417, N1551);
not NOT1 (N2422, N2407);
nor NOR4 (N2423, N2408, N1307, N792, N497);
nand NAND2 (N2424, N2411, N689);
buf BUF1 (N2425, N2424);
nor NOR3 (N2426, N2421, N263, N1170);
buf BUF1 (N2427, N2425);
xor XOR2 (N2428, N2426, N193);
or OR4 (N2429, N2404, N482, N321, N697);
buf BUF1 (N2430, N2422);
nor NOR2 (N2431, N2420, N616);
and AND4 (N2432, N2430, N1407, N1183, N65);
buf BUF1 (N2433, N2423);
not NOT1 (N2434, N2418);
not NOT1 (N2435, N2414);
xor XOR2 (N2436, N2434, N2054);
xor XOR2 (N2437, N2427, N1613);
nand NAND4 (N2438, N2431, N1114, N1301, N278);
buf BUF1 (N2439, N2433);
buf BUF1 (N2440, N2436);
buf BUF1 (N2441, N2437);
not NOT1 (N2442, N2429);
nor NOR3 (N2443, N2432, N2378, N828);
xor XOR2 (N2444, N2440, N1981);
or OR3 (N2445, N2444, N1400, N2136);
or OR3 (N2446, N2438, N2162, N2095);
nor NOR2 (N2447, N2439, N2164);
buf BUF1 (N2448, N2443);
buf BUF1 (N2449, N2435);
or OR3 (N2450, N2428, N2127, N1141);
and AND4 (N2451, N2445, N1486, N1617, N2307);
nand NAND2 (N2452, N2441, N939);
xor XOR2 (N2453, N2412, N1526);
or OR4 (N2454, N2450, N474, N1661, N333);
nor NOR2 (N2455, N2419, N1294);
buf BUF1 (N2456, N2448);
buf BUF1 (N2457, N2447);
and AND4 (N2458, N2452, N477, N1840, N222);
nor NOR3 (N2459, N2456, N2007, N126);
nand NAND3 (N2460, N2457, N1781, N2307);
or OR4 (N2461, N2451, N186, N911, N1159);
xor XOR2 (N2462, N2454, N1297);
nor NOR4 (N2463, N2449, N903, N625, N694);
nor NOR3 (N2464, N2460, N572, N521);
not NOT1 (N2465, N2462);
or OR4 (N2466, N2464, N544, N2310, N80);
and AND4 (N2467, N2458, N617, N1063, N1151);
buf BUF1 (N2468, N2465);
and AND4 (N2469, N2468, N2238, N1029, N1005);
or OR2 (N2470, N2455, N1422);
not NOT1 (N2471, N2466);
xor XOR2 (N2472, N2470, N1514);
xor XOR2 (N2473, N2442, N426);
buf BUF1 (N2474, N2473);
not NOT1 (N2475, N2467);
buf BUF1 (N2476, N2446);
not NOT1 (N2477, N2476);
nand NAND2 (N2478, N2475, N1073);
or OR4 (N2479, N2471, N1356, N546, N252);
not NOT1 (N2480, N2478);
or OR3 (N2481, N2472, N1279, N1718);
or OR2 (N2482, N2479, N2417);
nor NOR4 (N2483, N2482, N697, N678, N69);
nor NOR4 (N2484, N2474, N2471, N1640, N1323);
and AND3 (N2485, N2483, N690, N2245);
nor NOR3 (N2486, N2481, N276, N811);
buf BUF1 (N2487, N2463);
nor NOR2 (N2488, N2484, N605);
and AND4 (N2489, N2477, N1856, N808, N1826);
or OR2 (N2490, N2488, N2383);
buf BUF1 (N2491, N2486);
and AND3 (N2492, N2487, N623, N2042);
nand NAND4 (N2493, N2461, N536, N1866, N962);
xor XOR2 (N2494, N2480, N2111);
buf BUF1 (N2495, N2459);
or OR3 (N2496, N2494, N1510, N2053);
not NOT1 (N2497, N2492);
buf BUF1 (N2498, N2485);
nor NOR3 (N2499, N2493, N891, N1993);
xor XOR2 (N2500, N2496, N1756);
not NOT1 (N2501, N2499);
nor NOR2 (N2502, N2497, N2200);
not NOT1 (N2503, N2491);
nor NOR4 (N2504, N2495, N1390, N457, N300);
nand NAND3 (N2505, N2503, N1541, N41);
xor XOR2 (N2506, N2453, N2206);
or OR4 (N2507, N2490, N416, N859, N2350);
nand NAND4 (N2508, N2507, N560, N2016, N1761);
nor NOR2 (N2509, N2469, N2275);
nor NOR3 (N2510, N2506, N551, N392);
and AND2 (N2511, N2502, N580);
buf BUF1 (N2512, N2509);
buf BUF1 (N2513, N2504);
not NOT1 (N2514, N2489);
nor NOR4 (N2515, N2514, N1910, N562, N138);
buf BUF1 (N2516, N2508);
or OR2 (N2517, N2510, N1048);
and AND3 (N2518, N2516, N76, N1585);
or OR3 (N2519, N2517, N691, N2084);
not NOT1 (N2520, N2515);
buf BUF1 (N2521, N2512);
buf BUF1 (N2522, N2513);
buf BUF1 (N2523, N2498);
and AND4 (N2524, N2523, N629, N1610, N2458);
or OR2 (N2525, N2505, N735);
not NOT1 (N2526, N2511);
and AND3 (N2527, N2519, N1358, N1854);
xor XOR2 (N2528, N2525, N612);
nand NAND3 (N2529, N2527, N1917, N1873);
nand NAND3 (N2530, N2524, N1199, N1474);
xor XOR2 (N2531, N2530, N2288);
and AND2 (N2532, N2531, N2047);
xor XOR2 (N2533, N2501, N539);
xor XOR2 (N2534, N2522, N1997);
nor NOR4 (N2535, N2533, N2408, N1103, N1255);
nor NOR4 (N2536, N2518, N22, N1349, N1687);
nor NOR2 (N2537, N2520, N556);
and AND4 (N2538, N2532, N167, N2372, N552);
not NOT1 (N2539, N2529);
nand NAND3 (N2540, N2528, N943, N2332);
xor XOR2 (N2541, N2521, N2469);
buf BUF1 (N2542, N2537);
and AND3 (N2543, N2526, N1019, N104);
not NOT1 (N2544, N2538);
xor XOR2 (N2545, N2542, N28);
not NOT1 (N2546, N2545);
or OR2 (N2547, N2500, N1396);
not NOT1 (N2548, N2539);
or OR2 (N2549, N2544, N439);
xor XOR2 (N2550, N2541, N561);
or OR4 (N2551, N2536, N2434, N1924, N777);
not NOT1 (N2552, N2534);
nor NOR4 (N2553, N2540, N77, N533, N2232);
or OR3 (N2554, N2547, N216, N713);
xor XOR2 (N2555, N2535, N313);
not NOT1 (N2556, N2548);
not NOT1 (N2557, N2551);
and AND4 (N2558, N2556, N1500, N639, N210);
nor NOR4 (N2559, N2553, N2414, N921, N1208);
buf BUF1 (N2560, N2555);
xor XOR2 (N2561, N2554, N924);
nand NAND3 (N2562, N2549, N1381, N2232);
buf BUF1 (N2563, N2550);
xor XOR2 (N2564, N2562, N1962);
or OR4 (N2565, N2561, N1333, N1934, N670);
or OR4 (N2566, N2552, N59, N2047, N57);
and AND2 (N2567, N2543, N2472);
not NOT1 (N2568, N2558);
not NOT1 (N2569, N2560);
buf BUF1 (N2570, N2567);
nand NAND4 (N2571, N2568, N1760, N1827, N1205);
and AND2 (N2572, N2559, N877);
and AND3 (N2573, N2565, N1636, N1334);
and AND3 (N2574, N2571, N2235, N467);
or OR2 (N2575, N2546, N1952);
nand NAND4 (N2576, N2574, N2115, N1617, N1106);
buf BUF1 (N2577, N2576);
buf BUF1 (N2578, N2573);
nor NOR3 (N2579, N2563, N2202, N1682);
not NOT1 (N2580, N2564);
and AND4 (N2581, N2579, N1194, N863, N2419);
buf BUF1 (N2582, N2557);
or OR4 (N2583, N2575, N2120, N220, N1935);
not NOT1 (N2584, N2580);
and AND3 (N2585, N2572, N1241, N275);
xor XOR2 (N2586, N2566, N294);
and AND3 (N2587, N2585, N878, N1169);
not NOT1 (N2588, N2581);
nand NAND2 (N2589, N2584, N598);
xor XOR2 (N2590, N2569, N665);
buf BUF1 (N2591, N2586);
not NOT1 (N2592, N2578);
xor XOR2 (N2593, N2588, N2037);
buf BUF1 (N2594, N2590);
nor NOR4 (N2595, N2570, N1005, N955, N823);
not NOT1 (N2596, N2582);
not NOT1 (N2597, N2577);
xor XOR2 (N2598, N2591, N2233);
or OR3 (N2599, N2583, N530, N904);
and AND2 (N2600, N2589, N1085);
and AND3 (N2601, N2595, N719, N835);
nand NAND2 (N2602, N2596, N1564);
and AND2 (N2603, N2599, N2345);
buf BUF1 (N2604, N2602);
xor XOR2 (N2605, N2604, N918);
nand NAND2 (N2606, N2605, N1195);
not NOT1 (N2607, N2594);
nand NAND3 (N2608, N2603, N2358, N1248);
or OR3 (N2609, N2608, N495, N1684);
or OR3 (N2610, N2592, N2426, N1096);
nor NOR3 (N2611, N2587, N1215, N190);
nor NOR4 (N2612, N2607, N1371, N1179, N206);
not NOT1 (N2613, N2598);
nand NAND3 (N2614, N2600, N1314, N305);
buf BUF1 (N2615, N2613);
buf BUF1 (N2616, N2609);
xor XOR2 (N2617, N2593, N190);
not NOT1 (N2618, N2597);
nor NOR4 (N2619, N2618, N2248, N1152, N1433);
xor XOR2 (N2620, N2612, N285);
or OR4 (N2621, N2606, N1656, N1389, N368);
or OR2 (N2622, N2617, N733);
nor NOR4 (N2623, N2622, N1682, N1890, N2215);
not NOT1 (N2624, N2614);
buf BUF1 (N2625, N2624);
nor NOR2 (N2626, N2610, N814);
buf BUF1 (N2627, N2616);
not NOT1 (N2628, N2620);
and AND3 (N2629, N2619, N1546, N869);
xor XOR2 (N2630, N2626, N1674);
xor XOR2 (N2631, N2623, N339);
xor XOR2 (N2632, N2615, N1355);
xor XOR2 (N2633, N2629, N1285);
buf BUF1 (N2634, N2627);
and AND4 (N2635, N2621, N2287, N893, N1118);
nand NAND4 (N2636, N2601, N1703, N93, N1990);
or OR2 (N2637, N2632, N20);
nand NAND2 (N2638, N2611, N1094);
xor XOR2 (N2639, N2633, N152);
and AND4 (N2640, N2639, N2274, N1576, N1841);
or OR2 (N2641, N2637, N1778);
xor XOR2 (N2642, N2630, N1599);
not NOT1 (N2643, N2638);
nor NOR3 (N2644, N2631, N1687, N348);
nor NOR3 (N2645, N2625, N1942, N1405);
or OR4 (N2646, N2628, N368, N1942, N337);
not NOT1 (N2647, N2640);
not NOT1 (N2648, N2634);
nor NOR2 (N2649, N2648, N1183);
buf BUF1 (N2650, N2647);
not NOT1 (N2651, N2644);
buf BUF1 (N2652, N2635);
buf BUF1 (N2653, N2649);
and AND3 (N2654, N2636, N2494, N311);
not NOT1 (N2655, N2641);
and AND3 (N2656, N2643, N1498, N1940);
or OR3 (N2657, N2651, N602, N611);
not NOT1 (N2658, N2656);
or OR4 (N2659, N2654, N2425, N2518, N1947);
or OR3 (N2660, N2653, N1381, N1687);
xor XOR2 (N2661, N2645, N478);
xor XOR2 (N2662, N2658, N2648);
buf BUF1 (N2663, N2646);
and AND2 (N2664, N2650, N1252);
not NOT1 (N2665, N2642);
not NOT1 (N2666, N2657);
nor NOR3 (N2667, N2659, N2111, N1902);
not NOT1 (N2668, N2666);
not NOT1 (N2669, N2665);
buf BUF1 (N2670, N2668);
not NOT1 (N2671, N2663);
xor XOR2 (N2672, N2655, N1919);
xor XOR2 (N2673, N2671, N1617);
xor XOR2 (N2674, N2667, N15);
nand NAND3 (N2675, N2662, N470, N1887);
xor XOR2 (N2676, N2674, N2164);
nor NOR3 (N2677, N2670, N310, N670);
buf BUF1 (N2678, N2660);
buf BUF1 (N2679, N2661);
nand NAND4 (N2680, N2672, N227, N996, N1582);
nor NOR3 (N2681, N2669, N545, N1341);
buf BUF1 (N2682, N2676);
or OR3 (N2683, N2673, N1634, N1135);
nand NAND4 (N2684, N2652, N1404, N376, N556);
buf BUF1 (N2685, N2664);
or OR2 (N2686, N2675, N2469);
nand NAND4 (N2687, N2678, N2479, N1391, N2221);
buf BUF1 (N2688, N2687);
nor NOR3 (N2689, N2688, N24, N483);
or OR3 (N2690, N2677, N235, N78);
not NOT1 (N2691, N2683);
xor XOR2 (N2692, N2690, N2655);
buf BUF1 (N2693, N2682);
nand NAND2 (N2694, N2679, N2128);
buf BUF1 (N2695, N2680);
nand NAND3 (N2696, N2691, N307, N1840);
nor NOR2 (N2697, N2686, N61);
or OR4 (N2698, N2685, N2412, N1564, N369);
nand NAND2 (N2699, N2684, N1576);
xor XOR2 (N2700, N2692, N1998);
or OR4 (N2701, N2681, N1516, N2672, N424);
nor NOR3 (N2702, N2694, N2102, N1790);
buf BUF1 (N2703, N2701);
or OR3 (N2704, N2699, N63, N2122);
not NOT1 (N2705, N2700);
xor XOR2 (N2706, N2698, N2475);
and AND2 (N2707, N2705, N1725);
not NOT1 (N2708, N2697);
buf BUF1 (N2709, N2695);
nor NOR3 (N2710, N2709, N93, N590);
and AND2 (N2711, N2704, N2342);
nor NOR4 (N2712, N2707, N2185, N2097, N2154);
nor NOR4 (N2713, N2696, N1494, N272, N1097);
nor NOR4 (N2714, N2702, N1244, N2545, N827);
buf BUF1 (N2715, N2713);
not NOT1 (N2716, N2710);
not NOT1 (N2717, N2706);
buf BUF1 (N2718, N2717);
not NOT1 (N2719, N2711);
nor NOR4 (N2720, N2715, N2297, N1659, N113);
nand NAND2 (N2721, N2708, N258);
or OR2 (N2722, N2703, N2543);
nand NAND2 (N2723, N2720, N678);
not NOT1 (N2724, N2712);
nand NAND2 (N2725, N2718, N1941);
or OR4 (N2726, N2721, N897, N118, N2467);
not NOT1 (N2727, N2724);
buf BUF1 (N2728, N2722);
nor NOR4 (N2729, N2723, N2668, N769, N490);
buf BUF1 (N2730, N2727);
not NOT1 (N2731, N2725);
xor XOR2 (N2732, N2689, N1543);
nor NOR2 (N2733, N2693, N1320);
or OR3 (N2734, N2716, N1626, N1262);
nand NAND3 (N2735, N2733, N2309, N392);
and AND3 (N2736, N2731, N746, N2124);
xor XOR2 (N2737, N2732, N2181);
not NOT1 (N2738, N2719);
nand NAND2 (N2739, N2734, N256);
nor NOR4 (N2740, N2735, N2085, N2122, N1124);
not NOT1 (N2741, N2730);
not NOT1 (N2742, N2736);
and AND4 (N2743, N2714, N46, N1209, N134);
and AND4 (N2744, N2740, N1067, N371, N1714);
buf BUF1 (N2745, N2741);
xor XOR2 (N2746, N2742, N1799);
or OR2 (N2747, N2744, N2465);
buf BUF1 (N2748, N2726);
nor NOR4 (N2749, N2737, N828, N1000, N2507);
nand NAND3 (N2750, N2745, N40, N472);
xor XOR2 (N2751, N2729, N1951);
buf BUF1 (N2752, N2748);
buf BUF1 (N2753, N2739);
not NOT1 (N2754, N2746);
nor NOR2 (N2755, N2743, N1157);
not NOT1 (N2756, N2755);
nor NOR3 (N2757, N2747, N1803, N1473);
xor XOR2 (N2758, N2738, N627);
buf BUF1 (N2759, N2753);
and AND3 (N2760, N2752, N2665, N421);
nor NOR2 (N2761, N2756, N905);
or OR4 (N2762, N2759, N2729, N2109, N1578);
nand NAND4 (N2763, N2758, N1217, N2480, N472);
and AND2 (N2764, N2751, N1941);
nor NOR3 (N2765, N2749, N1557, N1103);
and AND2 (N2766, N2763, N1397);
nand NAND3 (N2767, N2762, N991, N569);
nor NOR4 (N2768, N2728, N498, N2767, N309);
buf BUF1 (N2769, N438);
nand NAND3 (N2770, N2757, N2546, N1710);
xor XOR2 (N2771, N2766, N2325);
or OR4 (N2772, N2770, N1959, N2252, N2689);
not NOT1 (N2773, N2768);
not NOT1 (N2774, N2754);
buf BUF1 (N2775, N2771);
buf BUF1 (N2776, N2773);
not NOT1 (N2777, N2769);
buf BUF1 (N2778, N2775);
or OR4 (N2779, N2765, N203, N350, N1620);
or OR4 (N2780, N2772, N451, N1392, N279);
nand NAND4 (N2781, N2776, N1365, N1613, N1061);
buf BUF1 (N2782, N2780);
not NOT1 (N2783, N2781);
or OR4 (N2784, N2761, N2079, N1988, N2290);
not NOT1 (N2785, N2779);
nor NOR3 (N2786, N2782, N329, N937);
buf BUF1 (N2787, N2760);
xor XOR2 (N2788, N2787, N1805);
nor NOR3 (N2789, N2778, N1389, N1923);
nand NAND4 (N2790, N2783, N407, N1263, N629);
or OR2 (N2791, N2750, N2062);
or OR2 (N2792, N2791, N907);
buf BUF1 (N2793, N2785);
or OR2 (N2794, N2789, N1507);
not NOT1 (N2795, N2794);
buf BUF1 (N2796, N2764);
and AND2 (N2797, N2777, N779);
or OR2 (N2798, N2795, N2268);
or OR4 (N2799, N2786, N224, N755, N177);
or OR2 (N2800, N2788, N690);
not NOT1 (N2801, N2800);
and AND2 (N2802, N2793, N493);
and AND4 (N2803, N2802, N2742, N2318, N2255);
not NOT1 (N2804, N2784);
not NOT1 (N2805, N2799);
nand NAND4 (N2806, N2774, N2575, N990, N2079);
nand NAND3 (N2807, N2803, N1147, N1806);
xor XOR2 (N2808, N2807, N857);
or OR3 (N2809, N2796, N2756, N1688);
nor NOR3 (N2810, N2809, N2760, N1581);
buf BUF1 (N2811, N2808);
and AND4 (N2812, N2801, N240, N2552, N1215);
nor NOR2 (N2813, N2797, N77);
xor XOR2 (N2814, N2805, N2064);
buf BUF1 (N2815, N2810);
and AND2 (N2816, N2814, N1301);
buf BUF1 (N2817, N2811);
and AND3 (N2818, N2817, N975, N246);
not NOT1 (N2819, N2804);
buf BUF1 (N2820, N2812);
nor NOR2 (N2821, N2818, N841);
and AND3 (N2822, N2815, N979, N1001);
or OR4 (N2823, N2813, N398, N350, N481);
xor XOR2 (N2824, N2806, N169);
nor NOR4 (N2825, N2822, N2678, N2193, N2441);
or OR4 (N2826, N2820, N389, N1480, N2612);
nor NOR4 (N2827, N2825, N537, N1045, N2176);
and AND2 (N2828, N2823, N595);
or OR3 (N2829, N2792, N1501, N124);
xor XOR2 (N2830, N2826, N1033);
nor NOR3 (N2831, N2829, N1357, N2612);
nor NOR4 (N2832, N2828, N1906, N722, N1818);
not NOT1 (N2833, N2798);
or OR2 (N2834, N2830, N2792);
or OR2 (N2835, N2790, N529);
nor NOR2 (N2836, N2827, N1866);
and AND2 (N2837, N2819, N2038);
and AND3 (N2838, N2836, N1375, N228);
buf BUF1 (N2839, N2821);
or OR2 (N2840, N2834, N678);
buf BUF1 (N2841, N2835);
not NOT1 (N2842, N2831);
buf BUF1 (N2843, N2838);
nand NAND4 (N2844, N2833, N903, N870, N2161);
xor XOR2 (N2845, N2844, N2684);
nand NAND2 (N2846, N2839, N1004);
or OR2 (N2847, N2837, N1748);
and AND4 (N2848, N2846, N2734, N553, N1992);
nand NAND4 (N2849, N2847, N2824, N1686, N277);
xor XOR2 (N2850, N1742, N2731);
xor XOR2 (N2851, N2849, N436);
nor NOR3 (N2852, N2816, N2575, N2229);
nor NOR3 (N2853, N2832, N297, N799);
nor NOR4 (N2854, N2850, N2234, N1622, N1338);
buf BUF1 (N2855, N2843);
and AND3 (N2856, N2842, N2336, N989);
nor NOR3 (N2857, N2856, N334, N538);
nor NOR2 (N2858, N2848, N2492);
not NOT1 (N2859, N2854);
nor NOR4 (N2860, N2841, N633, N1891, N1948);
nand NAND2 (N2861, N2855, N2525);
or OR4 (N2862, N2857, N1216, N1200, N1562);
xor XOR2 (N2863, N2845, N2179);
and AND3 (N2864, N2859, N1691, N1303);
not NOT1 (N2865, N2862);
xor XOR2 (N2866, N2852, N1753);
xor XOR2 (N2867, N2858, N2240);
nand NAND4 (N2868, N2860, N467, N1230, N1839);
nor NOR4 (N2869, N2863, N828, N212, N581);
not NOT1 (N2870, N2840);
xor XOR2 (N2871, N2869, N2421);
not NOT1 (N2872, N2851);
nor NOR4 (N2873, N2870, N65, N1694, N623);
nand NAND3 (N2874, N2867, N326, N1841);
nand NAND4 (N2875, N2853, N15, N1490, N1280);
or OR3 (N2876, N2861, N2475, N2276);
nand NAND2 (N2877, N2866, N87);
not NOT1 (N2878, N2877);
nand NAND2 (N2879, N2878, N1432);
buf BUF1 (N2880, N2868);
and AND3 (N2881, N2871, N1902, N2769);
and AND2 (N2882, N2872, N2039);
nor NOR2 (N2883, N2882, N1479);
buf BUF1 (N2884, N2875);
not NOT1 (N2885, N2879);
or OR3 (N2886, N2873, N1575, N794);
buf BUF1 (N2887, N2864);
and AND4 (N2888, N2884, N1875, N1837, N928);
nand NAND2 (N2889, N2881, N1051);
and AND2 (N2890, N2883, N600);
nor NOR3 (N2891, N2886, N148, N1949);
and AND4 (N2892, N2880, N2461, N1750, N2626);
buf BUF1 (N2893, N2865);
and AND3 (N2894, N2885, N1165, N1128);
xor XOR2 (N2895, N2894, N1586);
xor XOR2 (N2896, N2890, N1429);
nand NAND3 (N2897, N2896, N206, N2605);
not NOT1 (N2898, N2888);
buf BUF1 (N2899, N2892);
buf BUF1 (N2900, N2876);
or OR2 (N2901, N2900, N464);
nand NAND4 (N2902, N2897, N2522, N2361, N2520);
nand NAND2 (N2903, N2874, N588);
nand NAND2 (N2904, N2898, N817);
and AND2 (N2905, N2895, N494);
and AND2 (N2906, N2891, N309);
nand NAND3 (N2907, N2887, N1254, N453);
nor NOR3 (N2908, N2893, N2068, N488);
xor XOR2 (N2909, N2908, N1688);
xor XOR2 (N2910, N2905, N1199);
nor NOR2 (N2911, N2904, N266);
and AND2 (N2912, N2911, N2755);
and AND2 (N2913, N2910, N828);
nand NAND2 (N2914, N2903, N2384);
nor NOR2 (N2915, N2912, N262);
nor NOR2 (N2916, N2906, N2818);
nand NAND3 (N2917, N2909, N478, N1394);
xor XOR2 (N2918, N2914, N1363);
or OR2 (N2919, N2915, N1381);
or OR3 (N2920, N2919, N276, N2673);
xor XOR2 (N2921, N2920, N1117);
or OR3 (N2922, N2916, N839, N1752);
not NOT1 (N2923, N2899);
nand NAND2 (N2924, N2889, N2440);
and AND4 (N2925, N2901, N2718, N455, N2776);
nand NAND3 (N2926, N2922, N785, N448);
buf BUF1 (N2927, N2917);
not NOT1 (N2928, N2924);
nand NAND2 (N2929, N2907, N368);
xor XOR2 (N2930, N2929, N1174);
nand NAND4 (N2931, N2913, N1817, N29, N627);
and AND3 (N2932, N2931, N1163, N803);
and AND2 (N2933, N2930, N2169);
and AND4 (N2934, N2932, N1687, N1999, N1023);
and AND3 (N2935, N2934, N170, N1133);
nor NOR4 (N2936, N2935, N1139, N1412, N2189);
nand NAND3 (N2937, N2926, N1093, N19);
buf BUF1 (N2938, N2902);
and AND4 (N2939, N2933, N2729, N2230, N618);
buf BUF1 (N2940, N2918);
nand NAND4 (N2941, N2940, N2764, N238, N2454);
nor NOR2 (N2942, N2923, N719);
nor NOR2 (N2943, N2939, N2428);
xor XOR2 (N2944, N2936, N1002);
nor NOR3 (N2945, N2943, N797, N527);
nand NAND2 (N2946, N2925, N988);
nand NAND3 (N2947, N2944, N2912, N1802);
and AND2 (N2948, N2928, N572);
buf BUF1 (N2949, N2945);
nor NOR2 (N2950, N2938, N2280);
nand NAND2 (N2951, N2948, N292);
nor NOR2 (N2952, N2947, N2718);
nand NAND3 (N2953, N2952, N461, N1586);
nand NAND4 (N2954, N2953, N49, N2671, N481);
nor NOR2 (N2955, N2942, N2055);
buf BUF1 (N2956, N2950);
buf BUF1 (N2957, N2956);
or OR3 (N2958, N2941, N1706, N1435);
not NOT1 (N2959, N2957);
and AND3 (N2960, N2954, N2221, N1827);
nor NOR2 (N2961, N2927, N957);
nor NOR2 (N2962, N2951, N2310);
buf BUF1 (N2963, N2949);
not NOT1 (N2964, N2961);
and AND3 (N2965, N2964, N1918, N1523);
or OR4 (N2966, N2958, N1433, N950, N240);
or OR4 (N2967, N2962, N467, N537, N212);
xor XOR2 (N2968, N2967, N593);
nor NOR2 (N2969, N2946, N2861);
or OR4 (N2970, N2937, N1659, N2196, N107);
nand NAND3 (N2971, N2955, N2906, N2658);
not NOT1 (N2972, N2966);
not NOT1 (N2973, N2970);
not NOT1 (N2974, N2972);
nor NOR3 (N2975, N2959, N864, N2549);
buf BUF1 (N2976, N2973);
xor XOR2 (N2977, N2971, N2292);
or OR2 (N2978, N2968, N2758);
nand NAND2 (N2979, N2960, N2659);
or OR3 (N2980, N2979, N2537, N734);
and AND2 (N2981, N2976, N2092);
nand NAND2 (N2982, N2969, N85);
and AND4 (N2983, N2978, N285, N1835, N233);
xor XOR2 (N2984, N2980, N412);
xor XOR2 (N2985, N2977, N1938);
and AND2 (N2986, N2984, N1649);
not NOT1 (N2987, N2965);
nor NOR2 (N2988, N2983, N1691);
or OR2 (N2989, N2987, N27);
or OR2 (N2990, N2921, N426);
nor NOR3 (N2991, N2990, N770, N1744);
nand NAND2 (N2992, N2986, N1544);
buf BUF1 (N2993, N2989);
nor NOR4 (N2994, N2992, N1355, N556, N2679);
and AND4 (N2995, N2963, N2537, N1968, N2332);
buf BUF1 (N2996, N2982);
or OR4 (N2997, N2985, N2121, N520, N758);
nor NOR3 (N2998, N2974, N1358, N886);
nor NOR2 (N2999, N2995, N2404);
nor NOR4 (N3000, N2991, N2984, N2126, N2628);
buf BUF1 (N3001, N3000);
buf BUF1 (N3002, N2994);
buf BUF1 (N3003, N3002);
xor XOR2 (N3004, N2997, N2807);
nor NOR2 (N3005, N2998, N2600);
and AND3 (N3006, N3001, N2447, N965);
not NOT1 (N3007, N3004);
nor NOR2 (N3008, N2999, N2906);
buf BUF1 (N3009, N3003);
not NOT1 (N3010, N3007);
and AND4 (N3011, N3009, N1328, N2613, N2958);
xor XOR2 (N3012, N3005, N695);
buf BUF1 (N3013, N3006);
nand NAND4 (N3014, N2996, N1766, N73, N1681);
buf BUF1 (N3015, N3012);
and AND2 (N3016, N3008, N1712);
and AND4 (N3017, N2988, N2454, N2746, N96);
nor NOR2 (N3018, N3014, N1404);
nor NOR4 (N3019, N3016, N1003, N1244, N1313);
buf BUF1 (N3020, N2975);
or OR4 (N3021, N2993, N2158, N1448, N1723);
or OR2 (N3022, N3021, N1438);
nand NAND3 (N3023, N3018, N2778, N965);
nand NAND2 (N3024, N3023, N1952);
xor XOR2 (N3025, N3011, N486);
xor XOR2 (N3026, N3015, N1631);
xor XOR2 (N3027, N3017, N349);
not NOT1 (N3028, N3019);
or OR3 (N3029, N2981, N1795, N2490);
buf BUF1 (N3030, N3013);
not NOT1 (N3031, N3010);
nor NOR3 (N3032, N3024, N2679, N2751);
nand NAND4 (N3033, N3031, N156, N2660, N182);
nand NAND4 (N3034, N3032, N1707, N1999, N2293);
not NOT1 (N3035, N3028);
not NOT1 (N3036, N3025);
nor NOR4 (N3037, N3033, N887, N2644, N432);
or OR3 (N3038, N3030, N1074, N1373);
xor XOR2 (N3039, N3020, N680);
nor NOR4 (N3040, N3026, N2241, N1220, N1964);
or OR4 (N3041, N3039, N1073, N2676, N591);
nand NAND4 (N3042, N3027, N392, N2160, N1842);
buf BUF1 (N3043, N3040);
or OR2 (N3044, N3041, N2434);
nor NOR2 (N3045, N3044, N2876);
nor NOR3 (N3046, N3022, N1715, N1923);
and AND3 (N3047, N3043, N67, N456);
buf BUF1 (N3048, N3035);
xor XOR2 (N3049, N3048, N253);
buf BUF1 (N3050, N3042);
and AND4 (N3051, N3034, N352, N2522, N2756);
or OR4 (N3052, N3037, N2248, N1287, N156);
buf BUF1 (N3053, N3046);
not NOT1 (N3054, N3045);
buf BUF1 (N3055, N3047);
nand NAND2 (N3056, N3053, N2702);
not NOT1 (N3057, N3050);
not NOT1 (N3058, N3056);
nand NAND3 (N3059, N3054, N824, N1925);
buf BUF1 (N3060, N3059);
not NOT1 (N3061, N3055);
xor XOR2 (N3062, N3036, N1952);
not NOT1 (N3063, N3060);
xor XOR2 (N3064, N3061, N848);
and AND2 (N3065, N3029, N1966);
nand NAND2 (N3066, N3065, N2841);
nand NAND3 (N3067, N3063, N1073, N1391);
nand NAND4 (N3068, N3038, N717, N330, N695);
and AND3 (N3069, N3068, N1285, N2746);
buf BUF1 (N3070, N3066);
xor XOR2 (N3071, N3069, N95);
not NOT1 (N3072, N3052);
or OR4 (N3073, N3067, N796, N1983, N636);
nand NAND3 (N3074, N3064, N1287, N471);
xor XOR2 (N3075, N3074, N2519);
buf BUF1 (N3076, N3049);
or OR4 (N3077, N3073, N726, N458, N2034);
xor XOR2 (N3078, N3058, N2225);
buf BUF1 (N3079, N3071);
not NOT1 (N3080, N3070);
nor NOR2 (N3081, N3079, N2366);
nand NAND2 (N3082, N3078, N2101);
not NOT1 (N3083, N3076);
and AND4 (N3084, N3062, N2348, N2184, N2412);
or OR3 (N3085, N3075, N1477, N544);
xor XOR2 (N3086, N3082, N174);
buf BUF1 (N3087, N3084);
nand NAND2 (N3088, N3072, N1994);
nor NOR4 (N3089, N3088, N2867, N1592, N684);
and AND4 (N3090, N3087, N2945, N1399, N2022);
and AND3 (N3091, N3080, N1255, N2504);
and AND4 (N3092, N3090, N2114, N712, N1170);
and AND3 (N3093, N3081, N799, N2949);
buf BUF1 (N3094, N3086);
nand NAND4 (N3095, N3057, N1805, N934, N7);
not NOT1 (N3096, N3092);
nand NAND2 (N3097, N3094, N2564);
and AND3 (N3098, N3095, N283, N180);
nor NOR4 (N3099, N3096, N2949, N2367, N1350);
nor NOR3 (N3100, N3091, N2602, N354);
or OR2 (N3101, N3093, N1742);
nor NOR4 (N3102, N3089, N2610, N1986, N1785);
or OR2 (N3103, N3100, N570);
and AND3 (N3104, N3101, N2946, N2092);
nor NOR2 (N3105, N3077, N706);
and AND2 (N3106, N3085, N312);
or OR2 (N3107, N3105, N1518);
xor XOR2 (N3108, N3103, N680);
or OR3 (N3109, N3104, N900, N2585);
xor XOR2 (N3110, N3102, N1820);
nor NOR2 (N3111, N3110, N1814);
nand NAND2 (N3112, N3107, N2979);
xor XOR2 (N3113, N3098, N927);
buf BUF1 (N3114, N3111);
buf BUF1 (N3115, N3099);
nand NAND4 (N3116, N3083, N1411, N213, N784);
xor XOR2 (N3117, N3116, N1928);
nand NAND4 (N3118, N3117, N858, N1487, N1048);
xor XOR2 (N3119, N3108, N2001);
buf BUF1 (N3120, N3051);
xor XOR2 (N3121, N3114, N3064);
buf BUF1 (N3122, N3118);
not NOT1 (N3123, N3109);
and AND3 (N3124, N3121, N2035, N3042);
buf BUF1 (N3125, N3120);
xor XOR2 (N3126, N3119, N2767);
nand NAND3 (N3127, N3115, N2458, N1444);
nor NOR3 (N3128, N3127, N2322, N2087);
nor NOR2 (N3129, N3124, N546);
nand NAND3 (N3130, N3106, N3129, N1658);
or OR2 (N3131, N834, N1743);
buf BUF1 (N3132, N3122);
xor XOR2 (N3133, N3097, N1845);
nor NOR3 (N3134, N3131, N701, N2456);
buf BUF1 (N3135, N3133);
buf BUF1 (N3136, N3125);
and AND2 (N3137, N3128, N1304);
not NOT1 (N3138, N3112);
and AND3 (N3139, N3134, N2830, N2469);
buf BUF1 (N3140, N3137);
buf BUF1 (N3141, N3135);
nand NAND2 (N3142, N3132, N2828);
buf BUF1 (N3143, N3113);
buf BUF1 (N3144, N3126);
not NOT1 (N3145, N3143);
nor NOR4 (N3146, N3130, N1109, N1360, N2785);
nand NAND2 (N3147, N3140, N1483);
nand NAND3 (N3148, N3141, N97, N2504);
nand NAND2 (N3149, N3146, N685);
nand NAND2 (N3150, N3147, N1665);
buf BUF1 (N3151, N3139);
nand NAND2 (N3152, N3150, N921);
buf BUF1 (N3153, N3149);
and AND2 (N3154, N3136, N218);
or OR4 (N3155, N3151, N245, N774, N142);
xor XOR2 (N3156, N3138, N2441);
nand NAND2 (N3157, N3123, N3106);
nand NAND4 (N3158, N3154, N2487, N2003, N3070);
not NOT1 (N3159, N3156);
or OR4 (N3160, N3142, N896, N1476, N1325);
or OR4 (N3161, N3158, N131, N3096, N2125);
nand NAND4 (N3162, N3145, N2751, N1385, N2194);
xor XOR2 (N3163, N3161, N2538);
and AND4 (N3164, N3155, N727, N2445, N1281);
not NOT1 (N3165, N3160);
and AND2 (N3166, N3159, N352);
or OR4 (N3167, N3166, N1554, N2098, N1406);
buf BUF1 (N3168, N3157);
nor NOR4 (N3169, N3152, N613, N937, N407);
and AND3 (N3170, N3165, N1690, N3052);
nand NAND3 (N3171, N3162, N529, N3170);
xor XOR2 (N3172, N1678, N1579);
and AND4 (N3173, N3153, N485, N521, N2235);
xor XOR2 (N3174, N3171, N2180);
or OR3 (N3175, N3163, N1115, N2856);
xor XOR2 (N3176, N3164, N1662);
nand NAND2 (N3177, N3148, N2651);
or OR2 (N3178, N3172, N641);
xor XOR2 (N3179, N3177, N2932);
and AND4 (N3180, N3174, N1574, N442, N798);
and AND2 (N3181, N3173, N1973);
nor NOR2 (N3182, N3175, N2023);
xor XOR2 (N3183, N3181, N3002);
not NOT1 (N3184, N3176);
xor XOR2 (N3185, N3183, N1501);
and AND2 (N3186, N3167, N183);
nand NAND3 (N3187, N3144, N2503, N1874);
xor XOR2 (N3188, N3182, N499);
and AND4 (N3189, N3185, N650, N407, N211);
not NOT1 (N3190, N3187);
xor XOR2 (N3191, N3178, N2846);
not NOT1 (N3192, N3186);
nor NOR4 (N3193, N3189, N2714, N2675, N2716);
nand NAND3 (N3194, N3191, N33, N2206);
xor XOR2 (N3195, N3169, N923);
buf BUF1 (N3196, N3194);
nor NOR4 (N3197, N3168, N2558, N1117, N978);
nand NAND2 (N3198, N3179, N1940);
xor XOR2 (N3199, N3188, N2890);
not NOT1 (N3200, N3192);
or OR3 (N3201, N3195, N1309, N1023);
nand NAND4 (N3202, N3199, N884, N2922, N2906);
not NOT1 (N3203, N3193);
nor NOR3 (N3204, N3202, N1938, N149);
nor NOR3 (N3205, N3184, N1684, N319);
buf BUF1 (N3206, N3204);
buf BUF1 (N3207, N3206);
or OR2 (N3208, N3200, N564);
xor XOR2 (N3209, N3197, N2178);
not NOT1 (N3210, N3208);
nor NOR2 (N3211, N3198, N2136);
not NOT1 (N3212, N3203);
nand NAND3 (N3213, N3205, N297, N3157);
not NOT1 (N3214, N3213);
and AND3 (N3215, N3209, N2910, N2276);
nand NAND3 (N3216, N3196, N10, N2416);
nand NAND2 (N3217, N3214, N2084);
not NOT1 (N3218, N3212);
or OR3 (N3219, N3190, N2663, N2488);
nor NOR2 (N3220, N3210, N2044);
or OR4 (N3221, N3219, N767, N2808, N1616);
and AND4 (N3222, N3221, N2330, N1345, N2908);
xor XOR2 (N3223, N3217, N2788);
or OR2 (N3224, N3223, N79);
nand NAND3 (N3225, N3180, N2985, N2182);
not NOT1 (N3226, N3211);
nor NOR2 (N3227, N3220, N1928);
nand NAND2 (N3228, N3222, N1048);
buf BUF1 (N3229, N3218);
nand NAND2 (N3230, N3201, N819);
nor NOR2 (N3231, N3224, N1435);
nor NOR2 (N3232, N3216, N594);
and AND2 (N3233, N3232, N1168);
not NOT1 (N3234, N3228);
xor XOR2 (N3235, N3227, N2145);
nand NAND3 (N3236, N3215, N1930, N2158);
buf BUF1 (N3237, N3231);
buf BUF1 (N3238, N3234);
or OR2 (N3239, N3238, N859);
nor NOR3 (N3240, N3207, N1376, N2457);
buf BUF1 (N3241, N3230);
and AND4 (N3242, N3225, N1445, N2430, N228);
and AND4 (N3243, N3229, N1009, N2198, N525);
nor NOR3 (N3244, N3235, N3232, N1052);
buf BUF1 (N3245, N3236);
nor NOR4 (N3246, N3241, N876, N2820, N1638);
nor NOR2 (N3247, N3240, N2755);
and AND3 (N3248, N3244, N873, N2184);
nand NAND4 (N3249, N3248, N581, N1220, N240);
or OR3 (N3250, N3239, N2573, N1419);
nor NOR3 (N3251, N3246, N546, N175);
buf BUF1 (N3252, N3247);
xor XOR2 (N3253, N3226, N1913);
nor NOR2 (N3254, N3243, N203);
not NOT1 (N3255, N3251);
not NOT1 (N3256, N3255);
buf BUF1 (N3257, N3242);
or OR4 (N3258, N3245, N1199, N1865, N2136);
nor NOR3 (N3259, N3233, N2338, N2911);
xor XOR2 (N3260, N3253, N2283);
nor NOR2 (N3261, N3259, N2496);
and AND3 (N3262, N3257, N865, N3088);
not NOT1 (N3263, N3237);
nor NOR3 (N3264, N3254, N2109, N344);
nor NOR2 (N3265, N3262, N1255);
or OR3 (N3266, N3263, N2876, N1501);
and AND4 (N3267, N3264, N1769, N1131, N1906);
xor XOR2 (N3268, N3252, N3017);
xor XOR2 (N3269, N3261, N1921);
nand NAND4 (N3270, N3256, N864, N1885, N2467);
and AND3 (N3271, N3268, N3137, N634);
and AND4 (N3272, N3271, N3240, N2429, N1010);
and AND2 (N3273, N3265, N958);
or OR2 (N3274, N3272, N2919);
nand NAND4 (N3275, N3269, N2815, N996, N1402);
and AND3 (N3276, N3270, N1152, N1855);
nand NAND4 (N3277, N3266, N1312, N355, N1644);
nor NOR3 (N3278, N3275, N2987, N245);
and AND2 (N3279, N3260, N2728);
and AND4 (N3280, N3250, N2389, N659, N2908);
nand NAND3 (N3281, N3267, N2150, N758);
and AND2 (N3282, N3258, N643);
buf BUF1 (N3283, N3277);
buf BUF1 (N3284, N3276);
xor XOR2 (N3285, N3249, N2294);
not NOT1 (N3286, N3284);
not NOT1 (N3287, N3273);
or OR3 (N3288, N3281, N1715, N1731);
not NOT1 (N3289, N3280);
nor NOR3 (N3290, N3289, N2415, N1309);
not NOT1 (N3291, N3287);
xor XOR2 (N3292, N3290, N633);
xor XOR2 (N3293, N3279, N1630);
buf BUF1 (N3294, N3283);
not NOT1 (N3295, N3293);
nor NOR3 (N3296, N3274, N2584, N302);
nand NAND2 (N3297, N3292, N490);
buf BUF1 (N3298, N3296);
or OR4 (N3299, N3298, N1170, N2957, N2734);
and AND4 (N3300, N3291, N693, N683, N1602);
not NOT1 (N3301, N3286);
buf BUF1 (N3302, N3285);
nand NAND4 (N3303, N3297, N920, N2775, N3);
and AND2 (N3304, N3299, N3291);
or OR4 (N3305, N3300, N317, N709, N2231);
xor XOR2 (N3306, N3282, N2994);
xor XOR2 (N3307, N3305, N2042);
not NOT1 (N3308, N3303);
nor NOR2 (N3309, N3308, N3246);
nor NOR2 (N3310, N3309, N454);
buf BUF1 (N3311, N3307);
xor XOR2 (N3312, N3288, N1160);
xor XOR2 (N3313, N3294, N3301);
and AND3 (N3314, N3170, N2843, N3175);
xor XOR2 (N3315, N3314, N796);
buf BUF1 (N3316, N3313);
nand NAND3 (N3317, N3304, N2586, N2245);
or OR4 (N3318, N3317, N1071, N720, N527);
nand NAND3 (N3319, N3278, N950, N458);
nor NOR3 (N3320, N3316, N2594, N567);
xor XOR2 (N3321, N3319, N1834);
xor XOR2 (N3322, N3312, N1559);
xor XOR2 (N3323, N3322, N1669);
buf BUF1 (N3324, N3302);
xor XOR2 (N3325, N3306, N2678);
nor NOR3 (N3326, N3323, N1894, N1937);
not NOT1 (N3327, N3310);
xor XOR2 (N3328, N3320, N1219);
not NOT1 (N3329, N3324);
nor NOR4 (N3330, N3295, N2709, N1806, N2424);
or OR4 (N3331, N3330, N407, N394, N2839);
not NOT1 (N3332, N3318);
xor XOR2 (N3333, N3325, N1875);
nor NOR3 (N3334, N3326, N1164, N2410);
or OR3 (N3335, N3334, N456, N2618);
and AND3 (N3336, N3321, N508, N1622);
xor XOR2 (N3337, N3327, N2624);
nor NOR3 (N3338, N3315, N695, N1878);
nor NOR3 (N3339, N3332, N2161, N478);
xor XOR2 (N3340, N3333, N2087);
buf BUF1 (N3341, N3337);
and AND3 (N3342, N3311, N1957, N1535);
not NOT1 (N3343, N3336);
or OR3 (N3344, N3331, N1031, N2533);
not NOT1 (N3345, N3341);
nand NAND2 (N3346, N3338, N1502);
buf BUF1 (N3347, N3339);
xor XOR2 (N3348, N3328, N662);
buf BUF1 (N3349, N3346);
nand NAND4 (N3350, N3348, N1197, N2559, N2700);
or OR2 (N3351, N3343, N2028);
not NOT1 (N3352, N3347);
buf BUF1 (N3353, N3342);
nor NOR3 (N3354, N3344, N2031, N3281);
buf BUF1 (N3355, N3349);
xor XOR2 (N3356, N3329, N693);
buf BUF1 (N3357, N3335);
not NOT1 (N3358, N3352);
buf BUF1 (N3359, N3358);
not NOT1 (N3360, N3345);
not NOT1 (N3361, N3357);
not NOT1 (N3362, N3360);
buf BUF1 (N3363, N3361);
and AND2 (N3364, N3340, N1038);
xor XOR2 (N3365, N3354, N1879);
not NOT1 (N3366, N3362);
xor XOR2 (N3367, N3356, N2580);
not NOT1 (N3368, N3350);
or OR4 (N3369, N3351, N394, N2990, N90);
or OR2 (N3370, N3367, N326);
and AND4 (N3371, N3366, N2764, N452, N2288);
and AND4 (N3372, N3359, N2011, N3267, N1790);
nand NAND4 (N3373, N3368, N483, N1277, N781);
or OR3 (N3374, N3365, N138, N816);
and AND2 (N3375, N3363, N3101);
nor NOR3 (N3376, N3372, N363, N2367);
and AND3 (N3377, N3376, N604, N2846);
nand NAND2 (N3378, N3370, N2754);
xor XOR2 (N3379, N3374, N1698);
nand NAND3 (N3380, N3355, N189, N380);
nor NOR3 (N3381, N3379, N2760, N2586);
nand NAND4 (N3382, N3373, N2214, N1345, N1924);
nor NOR2 (N3383, N3378, N2113);
xor XOR2 (N3384, N3380, N3077);
buf BUF1 (N3385, N3377);
not NOT1 (N3386, N3385);
and AND4 (N3387, N3386, N11, N3007, N1819);
and AND4 (N3388, N3382, N14, N2058, N2170);
or OR3 (N3389, N3369, N176, N2558);
or OR3 (N3390, N3384, N63, N1981);
nor NOR2 (N3391, N3387, N953);
nand NAND2 (N3392, N3364, N3120);
nand NAND4 (N3393, N3371, N944, N704, N3185);
and AND2 (N3394, N3383, N3019);
nand NAND4 (N3395, N3381, N849, N2242, N964);
nand NAND2 (N3396, N3353, N2700);
not NOT1 (N3397, N3395);
or OR3 (N3398, N3392, N514, N147);
buf BUF1 (N3399, N3394);
xor XOR2 (N3400, N3389, N2150);
nor NOR4 (N3401, N3388, N172, N3272, N918);
not NOT1 (N3402, N3398);
or OR3 (N3403, N3390, N2023, N1076);
not NOT1 (N3404, N3393);
and AND2 (N3405, N3375, N1890);
xor XOR2 (N3406, N3403, N2585);
nand NAND3 (N3407, N3396, N2909, N3067);
xor XOR2 (N3408, N3397, N3058);
not NOT1 (N3409, N3406);
nor NOR2 (N3410, N3402, N2257);
and AND3 (N3411, N3410, N1931, N895);
buf BUF1 (N3412, N3409);
nand NAND4 (N3413, N3404, N2278, N179, N2288);
or OR4 (N3414, N3408, N1800, N847, N2694);
nand NAND2 (N3415, N3412, N521);
buf BUF1 (N3416, N3405);
nor NOR3 (N3417, N3411, N1554, N2063);
nand NAND3 (N3418, N3413, N1615, N1773);
and AND4 (N3419, N3391, N2345, N3241, N3237);
buf BUF1 (N3420, N3415);
buf BUF1 (N3421, N3417);
not NOT1 (N3422, N3401);
not NOT1 (N3423, N3400);
not NOT1 (N3424, N3399);
buf BUF1 (N3425, N3422);
buf BUF1 (N3426, N3421);
not NOT1 (N3427, N3414);
nor NOR2 (N3428, N3423, N813);
not NOT1 (N3429, N3425);
not NOT1 (N3430, N3416);
or OR4 (N3431, N3420, N3365, N355, N2070);
nor NOR3 (N3432, N3427, N148, N3079);
nand NAND2 (N3433, N3407, N2981);
buf BUF1 (N3434, N3418);
nand NAND3 (N3435, N3434, N3419, N1077);
buf BUF1 (N3436, N1659);
nor NOR3 (N3437, N3433, N3181, N1852);
buf BUF1 (N3438, N3436);
nand NAND2 (N3439, N3424, N2557);
nand NAND2 (N3440, N3428, N2073);
not NOT1 (N3441, N3431);
and AND4 (N3442, N3435, N1038, N723, N1621);
buf BUF1 (N3443, N3430);
nor NOR3 (N3444, N3438, N306, N672);
nand NAND2 (N3445, N3437, N3083);
and AND2 (N3446, N3441, N582);
and AND4 (N3447, N3429, N486, N2340, N1239);
or OR2 (N3448, N3446, N1822);
xor XOR2 (N3449, N3440, N2574);
nand NAND4 (N3450, N3432, N289, N3070, N767);
or OR2 (N3451, N3444, N962);
buf BUF1 (N3452, N3445);
buf BUF1 (N3453, N3442);
or OR2 (N3454, N3448, N3266);
nand NAND4 (N3455, N3453, N509, N2030, N2918);
nor NOR3 (N3456, N3451, N3324, N182);
nand NAND3 (N3457, N3456, N1184, N1131);
nand NAND2 (N3458, N3450, N266);
buf BUF1 (N3459, N3452);
buf BUF1 (N3460, N3439);
buf BUF1 (N3461, N3443);
not NOT1 (N3462, N3455);
and AND4 (N3463, N3457, N2207, N1278, N833);
or OR3 (N3464, N3454, N1427, N1092);
buf BUF1 (N3465, N3462);
not NOT1 (N3466, N3465);
buf BUF1 (N3467, N3466);
xor XOR2 (N3468, N3460, N1327);
buf BUF1 (N3469, N3447);
buf BUF1 (N3470, N3469);
not NOT1 (N3471, N3470);
and AND2 (N3472, N3459, N216);
nor NOR2 (N3473, N3472, N3439);
or OR4 (N3474, N3461, N1981, N1521, N1509);
or OR4 (N3475, N3467, N547, N1262, N2135);
and AND3 (N3476, N3463, N3462, N2490);
and AND3 (N3477, N3476, N2718, N2876);
and AND3 (N3478, N3477, N2594, N2614);
and AND4 (N3479, N3473, N2238, N3178, N2236);
and AND3 (N3480, N3468, N2750, N146);
buf BUF1 (N3481, N3474);
not NOT1 (N3482, N3471);
nor NOR4 (N3483, N3449, N572, N1237, N1379);
or OR4 (N3484, N3475, N2288, N971, N3130);
and AND4 (N3485, N3458, N2221, N2219, N961);
nand NAND3 (N3486, N3480, N3179, N1400);
and AND3 (N3487, N3486, N3449, N2045);
xor XOR2 (N3488, N3464, N3065);
nand NAND3 (N3489, N3483, N1669, N664);
or OR2 (N3490, N3482, N1565);
or OR4 (N3491, N3490, N139, N1918, N2748);
nand NAND3 (N3492, N3481, N2405, N444);
and AND4 (N3493, N3478, N3165, N2254, N1150);
buf BUF1 (N3494, N3488);
or OR2 (N3495, N3487, N1295);
and AND4 (N3496, N3479, N188, N1824, N981);
or OR3 (N3497, N3494, N909, N296);
nor NOR4 (N3498, N3426, N56, N2541, N949);
and AND3 (N3499, N3496, N3236, N2809);
xor XOR2 (N3500, N3495, N2715);
xor XOR2 (N3501, N3499, N1642);
and AND3 (N3502, N3489, N2736, N493);
nor NOR2 (N3503, N3500, N1374);
buf BUF1 (N3504, N3497);
nand NAND3 (N3505, N3502, N1864, N2289);
and AND2 (N3506, N3501, N1009);
xor XOR2 (N3507, N3505, N1181);
not NOT1 (N3508, N3498);
xor XOR2 (N3509, N3508, N2454);
and AND4 (N3510, N3485, N552, N1626, N773);
nor NOR2 (N3511, N3491, N881);
and AND2 (N3512, N3493, N98);
buf BUF1 (N3513, N3503);
or OR3 (N3514, N3507, N334, N835);
nor NOR4 (N3515, N3492, N9, N1439, N1036);
buf BUF1 (N3516, N3514);
xor XOR2 (N3517, N3504, N3467);
endmodule