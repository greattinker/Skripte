// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;

output N921,N913,N916,N911,N919,N887,N918,N923,N922,N924;

and AND3 (N25, N18, N17, N11);
nor NOR4 (N26, N21, N20, N25, N6);
or OR3 (N27, N1, N26, N7);
nor NOR4 (N28, N26, N11, N4, N16);
and AND2 (N29, N28, N5);
or OR2 (N30, N26, N19);
or OR2 (N31, N11, N15);
xor XOR2 (N32, N6, N25);
not NOT1 (N33, N5);
or OR2 (N34, N25, N10);
not NOT1 (N35, N25);
and AND2 (N36, N15, N24);
not NOT1 (N37, N23);
or OR2 (N38, N34, N5);
nor NOR2 (N39, N29, N35);
buf BUF1 (N40, N10);
or OR2 (N41, N36, N3);
nand NAND3 (N42, N38, N5, N9);
xor XOR2 (N43, N39, N15);
and AND2 (N44, N41, N5);
xor XOR2 (N45, N27, N36);
not NOT1 (N46, N42);
nand NAND2 (N47, N40, N22);
buf BUF1 (N48, N32);
xor XOR2 (N49, N31, N18);
or OR3 (N50, N48, N46, N48);
buf BUF1 (N51, N10);
and AND4 (N52, N51, N44, N8, N29);
nor NOR3 (N53, N25, N46, N51);
and AND3 (N54, N45, N28, N11);
buf BUF1 (N55, N53);
or OR3 (N56, N33, N39, N21);
or OR4 (N57, N49, N55, N55, N40);
or OR2 (N58, N41, N38);
or OR2 (N59, N54, N3);
and AND3 (N60, N37, N57, N6);
nand NAND4 (N61, N23, N30, N35, N57);
nand NAND2 (N62, N28, N26);
nor NOR3 (N63, N50, N1, N4);
buf BUF1 (N64, N62);
nor NOR4 (N65, N58, N35, N44, N20);
xor XOR2 (N66, N56, N49);
xor XOR2 (N67, N60, N11);
xor XOR2 (N68, N63, N39);
xor XOR2 (N69, N47, N42);
xor XOR2 (N70, N68, N50);
buf BUF1 (N71, N69);
nand NAND2 (N72, N61, N60);
xor XOR2 (N73, N59, N72);
not NOT1 (N74, N6);
xor XOR2 (N75, N73, N8);
nor NOR3 (N76, N71, N3, N2);
and AND2 (N77, N70, N25);
nor NOR4 (N78, N64, N16, N61, N73);
or OR2 (N79, N52, N4);
nor NOR3 (N80, N75, N27, N71);
xor XOR2 (N81, N67, N48);
and AND4 (N82, N81, N52, N22, N13);
nor NOR3 (N83, N82, N15, N39);
not NOT1 (N84, N43);
buf BUF1 (N85, N76);
xor XOR2 (N86, N85, N10);
nand NAND3 (N87, N84, N32, N43);
or OR3 (N88, N79, N18, N69);
or OR4 (N89, N87, N42, N50, N60);
or OR3 (N90, N83, N85, N19);
and AND3 (N91, N80, N38, N70);
buf BUF1 (N92, N74);
nand NAND4 (N93, N77, N9, N2, N44);
nand NAND4 (N94, N93, N82, N73, N37);
and AND3 (N95, N92, N80, N39);
nor NOR3 (N96, N86, N32, N29);
nand NAND2 (N97, N88, N10);
buf BUF1 (N98, N96);
buf BUF1 (N99, N89);
and AND4 (N100, N99, N93, N47, N6);
and AND2 (N101, N100, N20);
buf BUF1 (N102, N90);
buf BUF1 (N103, N78);
buf BUF1 (N104, N95);
nor NOR3 (N105, N66, N92, N39);
nand NAND2 (N106, N105, N102);
nand NAND3 (N107, N103, N79, N50);
xor XOR2 (N108, N67, N65);
not NOT1 (N109, N7);
and AND4 (N110, N107, N41, N39, N35);
buf BUF1 (N111, N104);
xor XOR2 (N112, N101, N49);
not NOT1 (N113, N94);
and AND2 (N114, N106, N18);
or OR2 (N115, N98, N67);
xor XOR2 (N116, N112, N79);
or OR3 (N117, N110, N23, N78);
xor XOR2 (N118, N111, N24);
or OR4 (N119, N113, N49, N25, N29);
buf BUF1 (N120, N109);
nand NAND3 (N121, N120, N109, N69);
and AND4 (N122, N116, N76, N28, N22);
not NOT1 (N123, N114);
or OR3 (N124, N123, N62, N122);
and AND4 (N125, N14, N67, N96, N91);
nor NOR2 (N126, N43, N111);
nand NAND4 (N127, N115, N20, N24, N121);
xor XOR2 (N128, N45, N122);
nor NOR4 (N129, N108, N22, N85, N105);
and AND2 (N130, N125, N58);
nand NAND2 (N131, N117, N63);
and AND4 (N132, N129, N38, N71, N101);
or OR3 (N133, N127, N70, N20);
xor XOR2 (N134, N128, N84);
buf BUF1 (N135, N118);
or OR4 (N136, N134, N6, N17, N131);
and AND3 (N137, N1, N106, N74);
not NOT1 (N138, N136);
buf BUF1 (N139, N132);
buf BUF1 (N140, N138);
not NOT1 (N141, N126);
and AND2 (N142, N141, N21);
nor NOR4 (N143, N124, N19, N48, N122);
or OR3 (N144, N140, N23, N122);
xor XOR2 (N145, N97, N118);
and AND3 (N146, N142, N99, N114);
nand NAND3 (N147, N130, N8, N141);
nor NOR3 (N148, N146, N143, N14);
not NOT1 (N149, N70);
buf BUF1 (N150, N139);
and AND4 (N151, N147, N95, N81, N83);
not NOT1 (N152, N135);
or OR3 (N153, N150, N6, N81);
nand NAND3 (N154, N153, N17, N64);
xor XOR2 (N155, N151, N141);
not NOT1 (N156, N137);
nor NOR2 (N157, N149, N145);
and AND4 (N158, N76, N105, N124, N76);
nand NAND2 (N159, N156, N133);
nor NOR3 (N160, N93, N26, N97);
not NOT1 (N161, N160);
not NOT1 (N162, N157);
xor XOR2 (N163, N162, N157);
buf BUF1 (N164, N159);
or OR4 (N165, N144, N149, N20, N90);
and AND2 (N166, N163, N39);
nor NOR3 (N167, N155, N45, N112);
buf BUF1 (N168, N152);
and AND3 (N169, N168, N153, N19);
nor NOR4 (N170, N154, N148, N162, N86);
nand NAND2 (N171, N71, N65);
nand NAND4 (N172, N164, N78, N98, N46);
xor XOR2 (N173, N158, N151);
not NOT1 (N174, N171);
nor NOR4 (N175, N167, N16, N134, N13);
not NOT1 (N176, N169);
xor XOR2 (N177, N166, N106);
and AND4 (N178, N177, N97, N144, N80);
or OR4 (N179, N161, N87, N117, N114);
xor XOR2 (N180, N175, N131);
or OR3 (N181, N165, N105, N162);
or OR4 (N182, N170, N117, N47, N103);
xor XOR2 (N183, N181, N178);
nor NOR2 (N184, N105, N138);
buf BUF1 (N185, N184);
nand NAND2 (N186, N172, N98);
xor XOR2 (N187, N185, N60);
and AND4 (N188, N187, N104, N127, N50);
and AND2 (N189, N180, N155);
not NOT1 (N190, N173);
or OR4 (N191, N119, N189, N38, N86);
nand NAND3 (N192, N184, N130, N115);
not NOT1 (N193, N191);
xor XOR2 (N194, N188, N186);
nor NOR2 (N195, N137, N32);
nor NOR4 (N196, N183, N146, N152, N57);
not NOT1 (N197, N195);
nor NOR3 (N198, N196, N157, N144);
buf BUF1 (N199, N198);
xor XOR2 (N200, N176, N142);
or OR2 (N201, N190, N167);
buf BUF1 (N202, N174);
or OR3 (N203, N201, N156, N18);
nor NOR3 (N204, N193, N60, N10);
buf BUF1 (N205, N200);
and AND2 (N206, N192, N112);
nand NAND2 (N207, N205, N195);
and AND3 (N208, N179, N142, N70);
buf BUF1 (N209, N206);
and AND4 (N210, N197, N181, N124, N40);
nand NAND2 (N211, N202, N49);
or OR3 (N212, N199, N87, N34);
and AND3 (N213, N182, N29, N47);
nand NAND2 (N214, N194, N210);
or OR3 (N215, N89, N167, N211);
and AND4 (N216, N176, N80, N37, N74);
nand NAND3 (N217, N213, N35, N198);
nor NOR3 (N218, N209, N51, N217);
not NOT1 (N219, N59);
or OR3 (N220, N212, N203, N197);
and AND4 (N221, N35, N118, N103, N169);
nand NAND3 (N222, N207, N109, N20);
nor NOR2 (N223, N220, N201);
buf BUF1 (N224, N222);
xor XOR2 (N225, N224, N107);
nand NAND3 (N226, N214, N82, N26);
nand NAND2 (N227, N225, N166);
not NOT1 (N228, N219);
xor XOR2 (N229, N227, N118);
nand NAND4 (N230, N218, N5, N3, N114);
or OR2 (N231, N228, N213);
nor NOR4 (N232, N223, N23, N49, N34);
nor NOR3 (N233, N231, N207, N209);
nand NAND4 (N234, N216, N153, N104, N3);
or OR4 (N235, N230, N47, N9, N196);
buf BUF1 (N236, N232);
not NOT1 (N237, N235);
or OR4 (N238, N234, N184, N143, N64);
nand NAND4 (N239, N237, N178, N153, N119);
nor NOR4 (N240, N208, N75, N70, N230);
buf BUF1 (N241, N236);
xor XOR2 (N242, N240, N14);
xor XOR2 (N243, N241, N225);
and AND3 (N244, N238, N176, N80);
and AND3 (N245, N243, N244, N233);
buf BUF1 (N246, N149);
buf BUF1 (N247, N107);
or OR3 (N248, N215, N230, N160);
buf BUF1 (N249, N246);
xor XOR2 (N250, N226, N125);
not NOT1 (N251, N204);
or OR3 (N252, N249, N185, N250);
nor NOR3 (N253, N195, N180, N64);
and AND4 (N254, N239, N166, N130, N221);
buf BUF1 (N255, N130);
nor NOR3 (N256, N245, N4, N125);
nor NOR4 (N257, N253, N176, N35, N245);
buf BUF1 (N258, N257);
nor NOR3 (N259, N254, N126, N11);
nand NAND4 (N260, N247, N134, N226, N192);
nand NAND4 (N261, N260, N47, N90, N168);
and AND2 (N262, N252, N51);
not NOT1 (N263, N255);
xor XOR2 (N264, N242, N73);
and AND4 (N265, N229, N22, N129, N106);
nor NOR3 (N266, N248, N259, N49);
xor XOR2 (N267, N6, N165);
nand NAND2 (N268, N267, N208);
and AND4 (N269, N251, N156, N46, N259);
and AND2 (N270, N268, N203);
xor XOR2 (N271, N261, N200);
nor NOR3 (N272, N270, N130, N66);
xor XOR2 (N273, N262, N76);
nand NAND3 (N274, N265, N113, N36);
and AND2 (N275, N272, N9);
not NOT1 (N276, N275);
xor XOR2 (N277, N276, N266);
not NOT1 (N278, N243);
or OR3 (N279, N277, N154, N46);
not NOT1 (N280, N263);
xor XOR2 (N281, N280, N254);
or OR4 (N282, N279, N220, N55, N258);
nand NAND4 (N283, N73, N202, N22, N90);
buf BUF1 (N284, N282);
nor NOR4 (N285, N281, N154, N8, N246);
xor XOR2 (N286, N285, N206);
or OR2 (N287, N284, N39);
xor XOR2 (N288, N278, N203);
nor NOR2 (N289, N264, N136);
nor NOR3 (N290, N256, N132, N10);
not NOT1 (N291, N289);
buf BUF1 (N292, N287);
nor NOR4 (N293, N291, N238, N69, N7);
or OR3 (N294, N286, N100, N226);
nand NAND4 (N295, N273, N42, N22, N208);
not NOT1 (N296, N292);
not NOT1 (N297, N283);
xor XOR2 (N298, N274, N136);
nand NAND2 (N299, N296, N93);
nor NOR3 (N300, N271, N72, N243);
not NOT1 (N301, N295);
nor NOR4 (N302, N301, N38, N3, N144);
nand NAND2 (N303, N298, N119);
buf BUF1 (N304, N299);
buf BUF1 (N305, N304);
nor NOR4 (N306, N302, N64, N154, N42);
buf BUF1 (N307, N303);
buf BUF1 (N308, N300);
and AND4 (N309, N306, N268, N183, N189);
nor NOR4 (N310, N269, N223, N247, N171);
and AND2 (N311, N310, N79);
not NOT1 (N312, N290);
and AND4 (N313, N294, N86, N267, N133);
nand NAND4 (N314, N297, N311, N133, N111);
xor XOR2 (N315, N129, N305);
xor XOR2 (N316, N295, N295);
nand NAND4 (N317, N314, N69, N267, N136);
nor NOR2 (N318, N293, N256);
and AND3 (N319, N309, N190, N304);
not NOT1 (N320, N307);
nand NAND3 (N321, N313, N181, N97);
and AND4 (N322, N315, N140, N14, N296);
xor XOR2 (N323, N288, N42);
and AND2 (N324, N319, N166);
and AND2 (N325, N321, N293);
and AND3 (N326, N323, N281, N305);
and AND4 (N327, N320, N227, N208, N287);
not NOT1 (N328, N327);
not NOT1 (N329, N322);
and AND2 (N330, N325, N48);
nand NAND2 (N331, N316, N244);
xor XOR2 (N332, N324, N116);
buf BUF1 (N333, N329);
nand NAND3 (N334, N330, N171, N275);
nor NOR3 (N335, N328, N119, N214);
nor NOR3 (N336, N308, N240, N151);
xor XOR2 (N337, N331, N309);
nor NOR4 (N338, N335, N16, N213, N16);
or OR3 (N339, N334, N153, N248);
xor XOR2 (N340, N339, N239);
and AND4 (N341, N338, N303, N102, N77);
xor XOR2 (N342, N312, N177);
nor NOR2 (N343, N337, N114);
buf BUF1 (N344, N343);
buf BUF1 (N345, N340);
nor NOR2 (N346, N342, N71);
xor XOR2 (N347, N344, N114);
xor XOR2 (N348, N336, N23);
and AND2 (N349, N346, N21);
not NOT1 (N350, N318);
xor XOR2 (N351, N349, N183);
xor XOR2 (N352, N351, N133);
buf BUF1 (N353, N350);
nor NOR2 (N354, N345, N293);
nor NOR4 (N355, N326, N310, N31, N118);
nor NOR3 (N356, N333, N184, N252);
or OR3 (N357, N332, N146, N42);
and AND4 (N358, N353, N158, N41, N343);
or OR3 (N359, N352, N72, N58);
and AND3 (N360, N356, N87, N72);
nor NOR3 (N361, N347, N73, N236);
or OR2 (N362, N360, N350);
nand NAND3 (N363, N354, N262, N302);
buf BUF1 (N364, N341);
nor NOR4 (N365, N363, N313, N213, N272);
or OR3 (N366, N355, N342, N337);
nand NAND4 (N367, N362, N360, N264, N118);
buf BUF1 (N368, N364);
not NOT1 (N369, N361);
and AND3 (N370, N368, N351, N322);
buf BUF1 (N371, N359);
nor NOR2 (N372, N365, N19);
nand NAND2 (N373, N367, N33);
or OR4 (N374, N369, N191, N205, N146);
xor XOR2 (N375, N366, N55);
nand NAND4 (N376, N373, N337, N177, N112);
nor NOR3 (N377, N370, N254, N295);
and AND3 (N378, N358, N139, N53);
nand NAND4 (N379, N357, N60, N60, N69);
not NOT1 (N380, N379);
nand NAND4 (N381, N378, N176, N27, N242);
not NOT1 (N382, N380);
and AND2 (N383, N376, N153);
xor XOR2 (N384, N372, N249);
or OR2 (N385, N381, N95);
not NOT1 (N386, N385);
buf BUF1 (N387, N382);
buf BUF1 (N388, N386);
buf BUF1 (N389, N374);
nor NOR4 (N390, N389, N362, N147, N156);
and AND3 (N391, N375, N88, N62);
or OR2 (N392, N384, N123);
nand NAND3 (N393, N377, N284, N4);
nor NOR2 (N394, N317, N211);
buf BUF1 (N395, N387);
not NOT1 (N396, N394);
xor XOR2 (N397, N383, N272);
and AND2 (N398, N391, N82);
or OR2 (N399, N395, N232);
not NOT1 (N400, N397);
nor NOR4 (N401, N390, N273, N76, N272);
or OR2 (N402, N392, N61);
or OR2 (N403, N400, N207);
buf BUF1 (N404, N399);
or OR2 (N405, N396, N144);
and AND4 (N406, N371, N374, N104, N1);
or OR2 (N407, N402, N208);
or OR3 (N408, N393, N368, N119);
or OR2 (N409, N406, N322);
not NOT1 (N410, N403);
not NOT1 (N411, N407);
nor NOR4 (N412, N404, N17, N126, N326);
buf BUF1 (N413, N411);
buf BUF1 (N414, N413);
nor NOR3 (N415, N405, N360, N210);
nor NOR4 (N416, N401, N284, N85, N109);
or OR2 (N417, N409, N233);
and AND3 (N418, N408, N322, N250);
or OR3 (N419, N398, N162, N108);
buf BUF1 (N420, N348);
and AND2 (N421, N420, N394);
not NOT1 (N422, N414);
nand NAND3 (N423, N421, N325, N121);
or OR4 (N424, N418, N185, N130, N362);
or OR2 (N425, N417, N317);
nor NOR2 (N426, N424, N131);
nand NAND2 (N427, N415, N1);
buf BUF1 (N428, N419);
and AND3 (N429, N427, N178, N146);
not NOT1 (N430, N422);
or OR4 (N431, N428, N295, N345, N180);
xor XOR2 (N432, N388, N279);
buf BUF1 (N433, N416);
nand NAND3 (N434, N429, N4, N304);
or OR4 (N435, N410, N265, N76, N402);
or OR4 (N436, N412, N280, N412, N93);
not NOT1 (N437, N433);
buf BUF1 (N438, N426);
not NOT1 (N439, N432);
not NOT1 (N440, N425);
xor XOR2 (N441, N440, N106);
xor XOR2 (N442, N436, N235);
nand NAND3 (N443, N441, N89, N211);
or OR3 (N444, N437, N106, N381);
buf BUF1 (N445, N423);
nor NOR3 (N446, N442, N363, N158);
xor XOR2 (N447, N430, N309);
or OR2 (N448, N447, N139);
or OR3 (N449, N438, N343, N272);
and AND3 (N450, N443, N336, N201);
not NOT1 (N451, N431);
not NOT1 (N452, N445);
nor NOR2 (N453, N449, N115);
nor NOR4 (N454, N452, N421, N29, N379);
buf BUF1 (N455, N446);
nor NOR3 (N456, N439, N215, N163);
nor NOR3 (N457, N448, N430, N129);
or OR3 (N458, N434, N207, N437);
buf BUF1 (N459, N435);
or OR3 (N460, N458, N237, N305);
buf BUF1 (N461, N456);
and AND2 (N462, N459, N263);
nor NOR3 (N463, N451, N142, N310);
nor NOR2 (N464, N455, N60);
nor NOR3 (N465, N463, N463, N69);
not NOT1 (N466, N460);
xor XOR2 (N467, N464, N269);
nor NOR3 (N468, N465, N310, N419);
nor NOR2 (N469, N468, N57);
and AND4 (N470, N462, N301, N364, N361);
nand NAND4 (N471, N467, N399, N348, N427);
nand NAND4 (N472, N450, N192, N260, N277);
nand NAND4 (N473, N469, N277, N50, N401);
nor NOR2 (N474, N453, N278);
buf BUF1 (N475, N444);
xor XOR2 (N476, N454, N91);
and AND2 (N477, N466, N343);
not NOT1 (N478, N475);
nand NAND4 (N479, N473, N460, N231, N247);
buf BUF1 (N480, N471);
or OR3 (N481, N470, N205, N316);
buf BUF1 (N482, N476);
buf BUF1 (N483, N461);
nand NAND2 (N484, N472, N53);
nor NOR3 (N485, N483, N125, N482);
xor XOR2 (N486, N322, N81);
nor NOR4 (N487, N457, N302, N384, N318);
nor NOR3 (N488, N487, N340, N10);
buf BUF1 (N489, N485);
not NOT1 (N490, N489);
nand NAND4 (N491, N477, N66, N443, N48);
and AND3 (N492, N490, N59, N133);
nor NOR2 (N493, N484, N12);
and AND3 (N494, N492, N464, N466);
or OR4 (N495, N488, N121, N224, N55);
xor XOR2 (N496, N478, N72);
not NOT1 (N497, N493);
or OR4 (N498, N486, N407, N414, N241);
nand NAND2 (N499, N481, N24);
nand NAND4 (N500, N498, N427, N239, N336);
nand NAND3 (N501, N480, N127, N486);
nand NAND3 (N502, N501, N165, N227);
nand NAND4 (N503, N474, N213, N258, N459);
xor XOR2 (N504, N500, N46);
nor NOR4 (N505, N496, N292, N19, N426);
or OR3 (N506, N491, N213, N432);
not NOT1 (N507, N497);
and AND4 (N508, N502, N57, N457, N64);
and AND3 (N509, N504, N496, N119);
and AND2 (N510, N507, N39);
xor XOR2 (N511, N508, N412);
xor XOR2 (N512, N499, N43);
nand NAND2 (N513, N494, N158);
nor NOR2 (N514, N506, N127);
not NOT1 (N515, N514);
nand NAND4 (N516, N479, N152, N337, N515);
nand NAND2 (N517, N480, N203);
not NOT1 (N518, N513);
xor XOR2 (N519, N512, N57);
nand NAND4 (N520, N503, N510, N114, N186);
or OR2 (N521, N65, N395);
nor NOR4 (N522, N519, N112, N451, N179);
or OR4 (N523, N522, N390, N267, N436);
buf BUF1 (N524, N518);
not NOT1 (N525, N521);
buf BUF1 (N526, N520);
nor NOR4 (N527, N505, N106, N305, N334);
xor XOR2 (N528, N524, N223);
not NOT1 (N529, N527);
nand NAND4 (N530, N526, N312, N472, N521);
or OR2 (N531, N528, N253);
nand NAND4 (N532, N509, N169, N413, N232);
not NOT1 (N533, N531);
not NOT1 (N534, N523);
not NOT1 (N535, N511);
or OR4 (N536, N530, N398, N160, N222);
nand NAND2 (N537, N536, N383);
xor XOR2 (N538, N534, N10);
xor XOR2 (N539, N532, N191);
nor NOR4 (N540, N516, N455, N475, N34);
xor XOR2 (N541, N517, N300);
and AND2 (N542, N535, N87);
xor XOR2 (N543, N533, N522);
buf BUF1 (N544, N543);
not NOT1 (N545, N537);
xor XOR2 (N546, N525, N325);
and AND4 (N547, N542, N323, N460, N510);
buf BUF1 (N548, N546);
or OR2 (N549, N547, N432);
nor NOR4 (N550, N529, N25, N105, N74);
xor XOR2 (N551, N545, N423);
not NOT1 (N552, N495);
and AND2 (N553, N544, N350);
xor XOR2 (N554, N540, N257);
xor XOR2 (N555, N538, N279);
or OR3 (N556, N548, N423, N188);
nand NAND2 (N557, N555, N178);
buf BUF1 (N558, N553);
and AND3 (N559, N554, N113, N25);
or OR4 (N560, N559, N515, N169, N448);
nand NAND3 (N561, N552, N45, N332);
xor XOR2 (N562, N557, N205);
not NOT1 (N563, N556);
nand NAND3 (N564, N558, N390, N499);
nand NAND2 (N565, N539, N82);
buf BUF1 (N566, N564);
and AND4 (N567, N563, N464, N22, N542);
and AND3 (N568, N562, N185, N495);
xor XOR2 (N569, N568, N472);
xor XOR2 (N570, N561, N415);
and AND2 (N571, N549, N179);
buf BUF1 (N572, N569);
not NOT1 (N573, N570);
and AND2 (N574, N541, N323);
nor NOR3 (N575, N565, N225, N61);
nor NOR2 (N576, N574, N358);
nor NOR2 (N577, N572, N334);
xor XOR2 (N578, N560, N12);
or OR4 (N579, N550, N446, N361, N76);
nor NOR2 (N580, N573, N550);
nor NOR3 (N581, N578, N338, N563);
nand NAND3 (N582, N575, N471, N451);
and AND3 (N583, N571, N449, N73);
nor NOR2 (N584, N581, N23);
and AND4 (N585, N551, N252, N341, N162);
buf BUF1 (N586, N582);
not NOT1 (N587, N585);
and AND2 (N588, N583, N75);
not NOT1 (N589, N579);
not NOT1 (N590, N589);
xor XOR2 (N591, N580, N3);
not NOT1 (N592, N588);
nand NAND3 (N593, N577, N72, N43);
not NOT1 (N594, N566);
and AND2 (N595, N567, N225);
and AND3 (N596, N593, N467, N75);
not NOT1 (N597, N592);
not NOT1 (N598, N591);
or OR3 (N599, N598, N422, N483);
nor NOR2 (N600, N597, N571);
buf BUF1 (N601, N587);
and AND2 (N602, N600, N150);
nor NOR4 (N603, N601, N164, N66, N131);
not NOT1 (N604, N596);
nand NAND4 (N605, N603, N248, N272, N555);
or OR2 (N606, N595, N272);
or OR4 (N607, N584, N172, N598, N378);
and AND2 (N608, N599, N285);
or OR3 (N609, N608, N558, N537);
xor XOR2 (N610, N602, N471);
or OR3 (N611, N590, N348, N549);
buf BUF1 (N612, N606);
or OR2 (N613, N607, N383);
not NOT1 (N614, N612);
nor NOR3 (N615, N604, N281, N614);
xor XOR2 (N616, N479, N341);
nand NAND2 (N617, N611, N289);
nand NAND4 (N618, N576, N612, N472, N334);
and AND4 (N619, N605, N374, N599, N459);
not NOT1 (N620, N618);
xor XOR2 (N621, N610, N374);
xor XOR2 (N622, N617, N316);
nand NAND4 (N623, N621, N113, N489, N455);
xor XOR2 (N624, N609, N74);
buf BUF1 (N625, N619);
nand NAND3 (N626, N613, N185, N304);
xor XOR2 (N627, N594, N312);
not NOT1 (N628, N624);
buf BUF1 (N629, N616);
buf BUF1 (N630, N620);
and AND3 (N631, N630, N499, N402);
not NOT1 (N632, N615);
nand NAND4 (N633, N631, N107, N99, N631);
buf BUF1 (N634, N623);
and AND3 (N635, N626, N124, N384);
or OR3 (N636, N625, N96, N144);
nand NAND4 (N637, N628, N26, N560, N118);
and AND2 (N638, N627, N442);
nand NAND2 (N639, N622, N389);
or OR2 (N640, N635, N458);
nand NAND4 (N641, N586, N163, N349, N155);
nand NAND4 (N642, N636, N25, N571, N346);
nand NAND2 (N643, N638, N362);
nor NOR3 (N644, N632, N521, N496);
xor XOR2 (N645, N639, N588);
not NOT1 (N646, N629);
nand NAND4 (N647, N642, N340, N236, N152);
and AND4 (N648, N641, N572, N210, N202);
xor XOR2 (N649, N646, N380);
not NOT1 (N650, N647);
nor NOR2 (N651, N643, N398);
nand NAND4 (N652, N649, N25, N102, N18);
nand NAND4 (N653, N637, N123, N623, N51);
xor XOR2 (N654, N648, N425);
and AND2 (N655, N651, N529);
buf BUF1 (N656, N633);
xor XOR2 (N657, N650, N95);
nand NAND2 (N658, N644, N161);
or OR4 (N659, N645, N616, N99, N385);
and AND4 (N660, N659, N27, N381, N184);
xor XOR2 (N661, N652, N301);
not NOT1 (N662, N634);
nor NOR2 (N663, N662, N163);
nor NOR4 (N664, N640, N36, N47, N31);
nand NAND3 (N665, N653, N173, N322);
nand NAND2 (N666, N656, N255);
and AND4 (N667, N661, N245, N330, N355);
xor XOR2 (N668, N657, N39);
not NOT1 (N669, N655);
xor XOR2 (N670, N654, N527);
and AND2 (N671, N665, N170);
and AND3 (N672, N669, N508, N348);
not NOT1 (N673, N658);
not NOT1 (N674, N673);
nor NOR2 (N675, N666, N345);
not NOT1 (N676, N667);
nand NAND3 (N677, N660, N441, N377);
or OR2 (N678, N664, N239);
or OR2 (N679, N674, N59);
nand NAND3 (N680, N668, N593, N62);
not NOT1 (N681, N677);
xor XOR2 (N682, N681, N240);
buf BUF1 (N683, N671);
xor XOR2 (N684, N676, N615);
xor XOR2 (N685, N678, N464);
buf BUF1 (N686, N675);
nand NAND2 (N687, N670, N320);
nor NOR2 (N688, N685, N679);
nor NOR2 (N689, N362, N635);
nor NOR3 (N690, N688, N86, N353);
or OR4 (N691, N686, N364, N265, N484);
nor NOR2 (N692, N682, N586);
or OR2 (N693, N687, N387);
not NOT1 (N694, N693);
and AND4 (N695, N684, N562, N622, N587);
xor XOR2 (N696, N690, N410);
nor NOR3 (N697, N689, N393, N541);
buf BUF1 (N698, N691);
buf BUF1 (N699, N692);
or OR2 (N700, N699, N422);
nand NAND4 (N701, N695, N489, N130, N14);
nand NAND4 (N702, N683, N190, N76, N612);
nor NOR4 (N703, N698, N208, N255, N319);
not NOT1 (N704, N680);
xor XOR2 (N705, N700, N288);
buf BUF1 (N706, N696);
nand NAND2 (N707, N705, N496);
nand NAND4 (N708, N697, N38, N351, N326);
buf BUF1 (N709, N707);
or OR2 (N710, N708, N437);
nor NOR4 (N711, N702, N248, N67, N438);
xor XOR2 (N712, N709, N287);
or OR2 (N713, N694, N322);
buf BUF1 (N714, N706);
nor NOR4 (N715, N714, N534, N3, N54);
and AND4 (N716, N663, N500, N192, N664);
nor NOR2 (N717, N712, N58);
not NOT1 (N718, N716);
nor NOR3 (N719, N711, N702, N243);
nand NAND3 (N720, N710, N316, N491);
nor NOR4 (N721, N672, N687, N306, N275);
nand NAND2 (N722, N720, N53);
buf BUF1 (N723, N704);
nor NOR4 (N724, N723, N179, N440, N203);
and AND4 (N725, N703, N407, N451, N412);
buf BUF1 (N726, N721);
xor XOR2 (N727, N719, N501);
xor XOR2 (N728, N701, N691);
nand NAND3 (N729, N728, N641, N326);
xor XOR2 (N730, N715, N435);
or OR3 (N731, N727, N401, N232);
xor XOR2 (N732, N713, N188);
nor NOR3 (N733, N724, N171, N223);
nand NAND2 (N734, N732, N415);
or OR4 (N735, N725, N240, N602, N727);
nor NOR4 (N736, N735, N76, N405, N433);
not NOT1 (N737, N733);
nand NAND2 (N738, N736, N618);
xor XOR2 (N739, N717, N3);
xor XOR2 (N740, N730, N455);
nor NOR4 (N741, N726, N609, N276, N468);
xor XOR2 (N742, N740, N484);
not NOT1 (N743, N734);
and AND2 (N744, N743, N234);
nor NOR2 (N745, N718, N652);
nand NAND3 (N746, N741, N426, N56);
not NOT1 (N747, N729);
or OR2 (N748, N746, N418);
nand NAND4 (N749, N739, N587, N353, N667);
or OR4 (N750, N731, N722, N300, N200);
nor NOR4 (N751, N253, N300, N10, N380);
not NOT1 (N752, N737);
nor NOR3 (N753, N752, N317, N507);
not NOT1 (N754, N742);
not NOT1 (N755, N747);
not NOT1 (N756, N745);
nor NOR4 (N757, N748, N657, N73, N548);
xor XOR2 (N758, N749, N721);
buf BUF1 (N759, N754);
nand NAND2 (N760, N757, N87);
or OR3 (N761, N760, N573, N484);
nand NAND4 (N762, N753, N240, N32, N571);
and AND2 (N763, N755, N122);
nand NAND3 (N764, N751, N606, N275);
xor XOR2 (N765, N763, N431);
not NOT1 (N766, N759);
xor XOR2 (N767, N762, N653);
xor XOR2 (N768, N756, N719);
buf BUF1 (N769, N764);
xor XOR2 (N770, N769, N580);
buf BUF1 (N771, N770);
nor NOR2 (N772, N750, N686);
nand NAND4 (N773, N766, N126, N197, N108);
xor XOR2 (N774, N771, N240);
not NOT1 (N775, N773);
nand NAND2 (N776, N767, N206);
nor NOR3 (N777, N768, N579, N37);
nand NAND4 (N778, N761, N639, N613, N92);
and AND3 (N779, N738, N59, N264);
and AND4 (N780, N744, N91, N460, N734);
buf BUF1 (N781, N776);
and AND2 (N782, N778, N157);
or OR3 (N783, N781, N488, N421);
nor NOR2 (N784, N780, N732);
xor XOR2 (N785, N758, N214);
or OR3 (N786, N779, N724, N509);
and AND3 (N787, N774, N86, N8);
nor NOR2 (N788, N765, N424);
nor NOR3 (N789, N783, N496, N438);
and AND3 (N790, N775, N92, N29);
xor XOR2 (N791, N782, N284);
or OR3 (N792, N772, N309, N110);
and AND2 (N793, N789, N235);
and AND4 (N794, N786, N179, N84, N522);
nand NAND3 (N795, N792, N260, N56);
buf BUF1 (N796, N791);
and AND4 (N797, N795, N429, N597, N771);
xor XOR2 (N798, N793, N4);
not NOT1 (N799, N797);
xor XOR2 (N800, N798, N761);
and AND3 (N801, N794, N263, N520);
xor XOR2 (N802, N788, N83);
or OR2 (N803, N796, N157);
buf BUF1 (N804, N784);
buf BUF1 (N805, N785);
not NOT1 (N806, N777);
nor NOR4 (N807, N805, N380, N355, N725);
nand NAND2 (N808, N799, N402);
nand NAND2 (N809, N803, N639);
or OR3 (N810, N807, N415, N18);
or OR3 (N811, N810, N108, N127);
buf BUF1 (N812, N802);
not NOT1 (N813, N811);
nand NAND2 (N814, N812, N89);
or OR4 (N815, N806, N104, N160, N65);
and AND4 (N816, N808, N66, N247, N681);
or OR4 (N817, N809, N275, N221, N160);
nor NOR4 (N818, N800, N168, N353, N263);
buf BUF1 (N819, N815);
xor XOR2 (N820, N804, N39);
buf BUF1 (N821, N813);
or OR3 (N822, N820, N323, N618);
buf BUF1 (N823, N816);
nor NOR4 (N824, N814, N276, N574, N496);
xor XOR2 (N825, N823, N430);
nand NAND3 (N826, N790, N632, N764);
buf BUF1 (N827, N819);
buf BUF1 (N828, N822);
xor XOR2 (N829, N827, N80);
nand NAND4 (N830, N829, N738, N744, N803);
not NOT1 (N831, N824);
or OR3 (N832, N787, N197, N133);
not NOT1 (N833, N826);
nor NOR4 (N834, N831, N306, N321, N710);
xor XOR2 (N835, N825, N509);
xor XOR2 (N836, N828, N184);
or OR4 (N837, N834, N603, N295, N809);
xor XOR2 (N838, N830, N363);
nor NOR2 (N839, N835, N518);
xor XOR2 (N840, N836, N361);
not NOT1 (N841, N833);
not NOT1 (N842, N841);
xor XOR2 (N843, N832, N321);
not NOT1 (N844, N801);
and AND2 (N845, N838, N643);
nand NAND2 (N846, N839, N521);
and AND3 (N847, N842, N793, N720);
and AND3 (N848, N847, N116, N214);
and AND3 (N849, N817, N4, N232);
and AND4 (N850, N818, N793, N618, N794);
xor XOR2 (N851, N845, N730);
nand NAND4 (N852, N850, N472, N354, N650);
and AND3 (N853, N843, N44, N25);
or OR3 (N854, N851, N531, N18);
and AND2 (N855, N854, N478);
or OR3 (N856, N844, N849, N110);
xor XOR2 (N857, N323, N421);
not NOT1 (N858, N821);
nor NOR3 (N859, N840, N450, N404);
buf BUF1 (N860, N853);
and AND2 (N861, N856, N833);
not NOT1 (N862, N860);
and AND3 (N863, N862, N209, N386);
buf BUF1 (N864, N846);
or OR3 (N865, N863, N718, N727);
xor XOR2 (N866, N852, N390);
or OR4 (N867, N864, N89, N136, N348);
nor NOR2 (N868, N861, N413);
or OR2 (N869, N867, N613);
nor NOR3 (N870, N837, N241, N735);
nand NAND3 (N871, N855, N147, N598);
nand NAND3 (N872, N870, N457, N30);
buf BUF1 (N873, N868);
xor XOR2 (N874, N848, N662);
and AND4 (N875, N858, N863, N592, N133);
and AND3 (N876, N871, N4, N92);
or OR3 (N877, N874, N227, N305);
or OR3 (N878, N877, N846, N641);
not NOT1 (N879, N876);
or OR3 (N880, N859, N373, N243);
nand NAND3 (N881, N878, N182, N738);
nand NAND3 (N882, N866, N267, N656);
nor NOR2 (N883, N881, N351);
or OR4 (N884, N879, N610, N762, N351);
and AND4 (N885, N882, N390, N847, N716);
nor NOR3 (N886, N865, N315, N359);
buf BUF1 (N887, N875);
nand NAND3 (N888, N885, N548, N74);
nor NOR2 (N889, N869, N284);
xor XOR2 (N890, N884, N472);
nor NOR4 (N891, N886, N152, N512, N679);
nand NAND2 (N892, N872, N610);
nand NAND4 (N893, N889, N687, N875, N803);
buf BUF1 (N894, N891);
nand NAND3 (N895, N880, N600, N209);
and AND4 (N896, N894, N370, N461, N299);
and AND3 (N897, N896, N440, N736);
nor NOR2 (N898, N888, N653);
or OR2 (N899, N897, N416);
not NOT1 (N900, N898);
and AND4 (N901, N873, N197, N592, N719);
nor NOR3 (N902, N893, N130, N71);
nor NOR4 (N903, N883, N687, N519, N545);
nor NOR2 (N904, N902, N170);
xor XOR2 (N905, N895, N563);
nand NAND2 (N906, N900, N376);
xor XOR2 (N907, N892, N1);
nand NAND3 (N908, N907, N207, N774);
buf BUF1 (N909, N906);
or OR3 (N910, N903, N144, N263);
buf BUF1 (N911, N857);
nand NAND2 (N912, N905, N690);
not NOT1 (N913, N901);
or OR4 (N914, N909, N788, N733, N466);
not NOT1 (N915, N912);
not NOT1 (N916, N910);
not NOT1 (N917, N914);
not NOT1 (N918, N899);
not NOT1 (N919, N890);
xor XOR2 (N920, N917, N224);
not NOT1 (N921, N904);
or OR2 (N922, N920, N739);
nand NAND2 (N923, N908, N232);
not NOT1 (N924, N915);
endmodule