// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15;

output N902,N897,N910,N914,N912,N896,N907,N884,N911,N915;

nand NAND3 (N16, N15, N9, N6);
not NOT1 (N17, N8);
or OR4 (N18, N15, N10, N8, N3);
or OR4 (N19, N11, N17, N7, N3);
not NOT1 (N20, N12);
not NOT1 (N21, N11);
nand NAND2 (N22, N17, N13);
xor XOR2 (N23, N10, N1);
not NOT1 (N24, N8);
xor XOR2 (N25, N14, N6);
nor NOR4 (N26, N6, N10, N10, N7);
not NOT1 (N27, N19);
xor XOR2 (N28, N21, N3);
or OR2 (N29, N20, N11);
nor NOR4 (N30, N25, N16, N14, N12);
and AND3 (N31, N13, N26, N27);
xor XOR2 (N32, N28, N8);
buf BUF1 (N33, N32);
nand NAND4 (N34, N27, N7, N23, N2);
buf BUF1 (N35, N23);
nand NAND2 (N36, N4, N21);
or OR2 (N37, N35, N24);
or OR3 (N38, N32, N10, N25);
nand NAND3 (N39, N36, N22, N2);
buf BUF1 (N40, N24);
or OR3 (N41, N38, N4, N30);
and AND2 (N42, N13, N28);
nor NOR3 (N43, N31, N26, N12);
nand NAND2 (N44, N18, N39);
not NOT1 (N45, N31);
nand NAND2 (N46, N34, N17);
not NOT1 (N47, N33);
and AND2 (N48, N47, N1);
nand NAND4 (N49, N46, N25, N20, N41);
and AND2 (N50, N49, N4);
buf BUF1 (N51, N26);
buf BUF1 (N52, N40);
xor XOR2 (N53, N43, N18);
or OR3 (N54, N45, N37, N43);
not NOT1 (N55, N42);
not NOT1 (N56, N34);
nand NAND3 (N57, N56, N8, N13);
and AND2 (N58, N53, N9);
nand NAND4 (N59, N54, N4, N58, N16);
xor XOR2 (N60, N40, N39);
not NOT1 (N61, N50);
buf BUF1 (N62, N60);
xor XOR2 (N63, N44, N34);
buf BUF1 (N64, N29);
not NOT1 (N65, N61);
not NOT1 (N66, N65);
or OR3 (N67, N66, N57, N50);
xor XOR2 (N68, N44, N67);
nor NOR3 (N69, N22, N44, N25);
buf BUF1 (N70, N68);
or OR3 (N71, N59, N21, N9);
and AND2 (N72, N70, N60);
buf BUF1 (N73, N55);
buf BUF1 (N74, N62);
nand NAND2 (N75, N51, N72);
not NOT1 (N76, N9);
or OR3 (N77, N69, N59, N11);
nor NOR2 (N78, N74, N24);
and AND3 (N79, N75, N43, N36);
nand NAND2 (N80, N71, N19);
xor XOR2 (N81, N79, N77);
nor NOR4 (N82, N31, N21, N55, N22);
xor XOR2 (N83, N78, N37);
not NOT1 (N84, N82);
xor XOR2 (N85, N64, N16);
nor NOR4 (N86, N80, N48, N16, N71);
not NOT1 (N87, N24);
nand NAND3 (N88, N83, N4, N33);
nand NAND4 (N89, N81, N5, N58, N83);
or OR2 (N90, N87, N70);
buf BUF1 (N91, N90);
xor XOR2 (N92, N52, N12);
nand NAND3 (N93, N73, N74, N70);
xor XOR2 (N94, N93, N63);
nor NOR3 (N95, N16, N75, N16);
or OR3 (N96, N95, N76, N79);
and AND3 (N97, N61, N43, N91);
nor NOR4 (N98, N30, N14, N6, N12);
and AND3 (N99, N85, N15, N54);
not NOT1 (N100, N96);
buf BUF1 (N101, N97);
xor XOR2 (N102, N100, N67);
xor XOR2 (N103, N92, N64);
not NOT1 (N104, N86);
or OR2 (N105, N101, N7);
buf BUF1 (N106, N104);
nand NAND4 (N107, N105, N44, N51, N69);
buf BUF1 (N108, N107);
or OR2 (N109, N102, N54);
not NOT1 (N110, N84);
xor XOR2 (N111, N106, N41);
nand NAND3 (N112, N89, N29, N15);
nor NOR2 (N113, N88, N12);
not NOT1 (N114, N94);
nand NAND4 (N115, N99, N107, N107, N13);
buf BUF1 (N116, N113);
nand NAND3 (N117, N108, N69, N18);
and AND3 (N118, N115, N13, N79);
buf BUF1 (N119, N109);
xor XOR2 (N120, N116, N31);
buf BUF1 (N121, N112);
or OR2 (N122, N114, N3);
buf BUF1 (N123, N122);
nor NOR4 (N124, N121, N33, N108, N111);
nor NOR4 (N125, N121, N99, N78, N11);
xor XOR2 (N126, N125, N121);
and AND3 (N127, N123, N126, N64);
and AND3 (N128, N70, N15, N54);
or OR3 (N129, N128, N73, N114);
buf BUF1 (N130, N120);
buf BUF1 (N131, N117);
and AND2 (N132, N119, N57);
and AND4 (N133, N103, N117, N14, N82);
buf BUF1 (N134, N130);
xor XOR2 (N135, N133, N58);
xor XOR2 (N136, N118, N97);
xor XOR2 (N137, N129, N76);
buf BUF1 (N138, N131);
not NOT1 (N139, N135);
buf BUF1 (N140, N110);
nor NOR4 (N141, N134, N89, N41, N21);
and AND2 (N142, N140, N31);
or OR3 (N143, N136, N19, N135);
buf BUF1 (N144, N143);
or OR2 (N145, N127, N62);
and AND3 (N146, N144, N80, N10);
or OR2 (N147, N142, N77);
nor NOR2 (N148, N137, N39);
or OR4 (N149, N138, N118, N10, N49);
or OR3 (N150, N147, N25, N107);
xor XOR2 (N151, N145, N132);
or OR2 (N152, N1, N20);
nor NOR2 (N153, N152, N116);
not NOT1 (N154, N150);
and AND2 (N155, N154, N112);
not NOT1 (N156, N155);
nand NAND2 (N157, N98, N39);
buf BUF1 (N158, N151);
or OR4 (N159, N124, N44, N88, N135);
and AND2 (N160, N159, N58);
or OR2 (N161, N139, N68);
buf BUF1 (N162, N146);
not NOT1 (N163, N153);
buf BUF1 (N164, N158);
nand NAND2 (N165, N161, N17);
not NOT1 (N166, N148);
or OR2 (N167, N157, N35);
nor NOR3 (N168, N165, N69, N86);
not NOT1 (N169, N141);
xor XOR2 (N170, N168, N96);
not NOT1 (N171, N149);
and AND3 (N172, N162, N10, N14);
nor NOR4 (N173, N166, N6, N17, N133);
and AND4 (N174, N160, N2, N42, N119);
xor XOR2 (N175, N163, N46);
and AND3 (N176, N167, N157, N42);
or OR3 (N177, N164, N109, N16);
nor NOR4 (N178, N172, N144, N36, N27);
or OR2 (N179, N178, N142);
nand NAND4 (N180, N176, N91, N83, N6);
or OR4 (N181, N177, N49, N166, N61);
xor XOR2 (N182, N169, N11);
or OR3 (N183, N180, N137, N69);
buf BUF1 (N184, N181);
xor XOR2 (N185, N171, N124);
or OR3 (N186, N179, N63, N103);
not NOT1 (N187, N182);
nand NAND4 (N188, N173, N46, N78, N169);
buf BUF1 (N189, N188);
not NOT1 (N190, N183);
and AND3 (N191, N189, N115, N142);
buf BUF1 (N192, N185);
or OR2 (N193, N175, N189);
not NOT1 (N194, N191);
not NOT1 (N195, N187);
not NOT1 (N196, N156);
nor NOR2 (N197, N196, N143);
not NOT1 (N198, N192);
not NOT1 (N199, N184);
xor XOR2 (N200, N194, N77);
not NOT1 (N201, N198);
or OR3 (N202, N190, N108, N14);
or OR3 (N203, N174, N2, N194);
buf BUF1 (N204, N193);
buf BUF1 (N205, N195);
xor XOR2 (N206, N203, N23);
not NOT1 (N207, N197);
or OR2 (N208, N201, N129);
buf BUF1 (N209, N202);
or OR3 (N210, N199, N180, N102);
or OR4 (N211, N186, N65, N38, N65);
xor XOR2 (N212, N211, N51);
nand NAND3 (N213, N209, N173, N33);
and AND2 (N214, N170, N43);
not NOT1 (N215, N212);
xor XOR2 (N216, N207, N82);
or OR3 (N217, N216, N102, N99);
or OR2 (N218, N217, N153);
not NOT1 (N219, N214);
and AND3 (N220, N213, N56, N72);
buf BUF1 (N221, N215);
xor XOR2 (N222, N210, N185);
not NOT1 (N223, N221);
xor XOR2 (N224, N205, N140);
xor XOR2 (N225, N224, N104);
or OR4 (N226, N222, N218, N136, N112);
xor XOR2 (N227, N143, N33);
and AND3 (N228, N226, N154, N98);
not NOT1 (N229, N204);
buf BUF1 (N230, N225);
nor NOR4 (N231, N208, N181, N118, N149);
or OR3 (N232, N219, N112, N177);
nand NAND3 (N233, N231, N41, N187);
nor NOR3 (N234, N200, N100, N127);
not NOT1 (N235, N206);
xor XOR2 (N236, N232, N4);
not NOT1 (N237, N220);
nand NAND2 (N238, N234, N138);
and AND4 (N239, N223, N152, N197, N138);
nand NAND3 (N240, N238, N7, N86);
buf BUF1 (N241, N228);
xor XOR2 (N242, N241, N204);
not NOT1 (N243, N235);
buf BUF1 (N244, N230);
and AND2 (N245, N229, N56);
buf BUF1 (N246, N245);
or OR2 (N247, N243, N52);
or OR2 (N248, N244, N144);
not NOT1 (N249, N239);
nor NOR2 (N250, N237, N14);
nand NAND3 (N251, N242, N85, N33);
nand NAND2 (N252, N251, N110);
nor NOR3 (N253, N247, N156, N131);
xor XOR2 (N254, N252, N60);
xor XOR2 (N255, N233, N195);
or OR3 (N256, N246, N72, N18);
not NOT1 (N257, N248);
xor XOR2 (N258, N240, N230);
nor NOR2 (N259, N257, N143);
buf BUF1 (N260, N253);
buf BUF1 (N261, N255);
nor NOR3 (N262, N256, N76, N258);
nand NAND2 (N263, N131, N261);
xor XOR2 (N264, N63, N168);
and AND3 (N265, N249, N61, N55);
or OR3 (N266, N254, N134, N57);
or OR2 (N267, N227, N188);
or OR4 (N268, N266, N57, N139, N70);
not NOT1 (N269, N262);
nor NOR3 (N270, N268, N267, N173);
buf BUF1 (N271, N10);
or OR4 (N272, N265, N77, N153, N12);
or OR4 (N273, N269, N52, N149, N25);
or OR4 (N274, N260, N224, N124, N219);
or OR4 (N275, N250, N183, N35, N74);
nand NAND3 (N276, N273, N71, N160);
nand NAND2 (N277, N272, N20);
not NOT1 (N278, N259);
not NOT1 (N279, N274);
xor XOR2 (N280, N279, N20);
and AND4 (N281, N275, N182, N81, N134);
nor NOR4 (N282, N281, N159, N170, N270);
and AND3 (N283, N116, N11, N183);
or OR3 (N284, N283, N248, N20);
and AND2 (N285, N276, N33);
not NOT1 (N286, N282);
not NOT1 (N287, N236);
nand NAND3 (N288, N286, N38, N20);
not NOT1 (N289, N264);
nand NAND4 (N290, N289, N27, N131, N238);
and AND2 (N291, N278, N104);
not NOT1 (N292, N263);
nand NAND2 (N293, N285, N74);
not NOT1 (N294, N292);
and AND2 (N295, N294, N58);
xor XOR2 (N296, N290, N223);
buf BUF1 (N297, N288);
xor XOR2 (N298, N280, N16);
nand NAND4 (N299, N291, N282, N297, N17);
nor NOR2 (N300, N61, N252);
and AND3 (N301, N277, N110, N238);
or OR2 (N302, N287, N88);
nor NOR2 (N303, N284, N191);
nor NOR4 (N304, N302, N104, N118, N19);
xor XOR2 (N305, N301, N160);
xor XOR2 (N306, N300, N294);
nor NOR3 (N307, N303, N56, N111);
and AND3 (N308, N307, N277, N145);
nand NAND3 (N309, N304, N69, N176);
and AND4 (N310, N306, N69, N159, N36);
nand NAND2 (N311, N299, N61);
xor XOR2 (N312, N311, N270);
not NOT1 (N313, N308);
buf BUF1 (N314, N271);
xor XOR2 (N315, N313, N266);
nor NOR4 (N316, N295, N82, N203, N15);
and AND4 (N317, N314, N100, N241, N250);
xor XOR2 (N318, N305, N301);
or OR2 (N319, N316, N109);
not NOT1 (N320, N310);
xor XOR2 (N321, N309, N148);
buf BUF1 (N322, N317);
or OR2 (N323, N312, N178);
nor NOR2 (N324, N323, N67);
not NOT1 (N325, N324);
buf BUF1 (N326, N320);
nor NOR4 (N327, N318, N229, N306, N224);
buf BUF1 (N328, N326);
buf BUF1 (N329, N319);
buf BUF1 (N330, N315);
or OR4 (N331, N322, N61, N40, N154);
nand NAND2 (N332, N330, N169);
and AND2 (N333, N321, N69);
not NOT1 (N334, N298);
nor NOR3 (N335, N327, N307, N226);
or OR2 (N336, N329, N34);
xor XOR2 (N337, N335, N155);
and AND2 (N338, N293, N148);
nor NOR2 (N339, N338, N82);
xor XOR2 (N340, N331, N160);
and AND3 (N341, N325, N173, N146);
and AND2 (N342, N296, N335);
not NOT1 (N343, N339);
nand NAND3 (N344, N341, N50, N228);
or OR4 (N345, N334, N299, N126, N323);
not NOT1 (N346, N342);
not NOT1 (N347, N336);
xor XOR2 (N348, N340, N164);
or OR4 (N349, N333, N44, N113, N39);
nand NAND4 (N350, N344, N299, N278, N87);
buf BUF1 (N351, N328);
nor NOR2 (N352, N343, N143);
and AND3 (N353, N337, N171, N287);
or OR2 (N354, N349, N48);
or OR3 (N355, N346, N109, N351);
or OR4 (N356, N128, N87, N28, N31);
nand NAND2 (N357, N348, N169);
buf BUF1 (N358, N332);
and AND2 (N359, N358, N69);
and AND2 (N360, N345, N296);
not NOT1 (N361, N356);
xor XOR2 (N362, N361, N39);
and AND2 (N363, N359, N244);
buf BUF1 (N364, N362);
buf BUF1 (N365, N353);
or OR2 (N366, N363, N196);
buf BUF1 (N367, N357);
not NOT1 (N368, N364);
or OR4 (N369, N355, N33, N1, N182);
xor XOR2 (N370, N369, N57);
not NOT1 (N371, N350);
not NOT1 (N372, N365);
buf BUF1 (N373, N366);
or OR2 (N374, N373, N18);
or OR2 (N375, N368, N14);
buf BUF1 (N376, N354);
and AND4 (N377, N352, N89, N17, N237);
buf BUF1 (N378, N360);
buf BUF1 (N379, N375);
or OR3 (N380, N372, N342, N139);
not NOT1 (N381, N380);
nand NAND4 (N382, N378, N279, N339, N226);
or OR2 (N383, N371, N111);
nor NOR2 (N384, N382, N164);
nor NOR4 (N385, N384, N336, N139, N274);
xor XOR2 (N386, N376, N236);
nand NAND4 (N387, N370, N22, N211, N229);
not NOT1 (N388, N383);
nor NOR3 (N389, N387, N16, N316);
buf BUF1 (N390, N367);
not NOT1 (N391, N347);
not NOT1 (N392, N390);
not NOT1 (N393, N385);
and AND4 (N394, N386, N178, N105, N336);
nand NAND3 (N395, N374, N392, N40);
buf BUF1 (N396, N367);
buf BUF1 (N397, N381);
xor XOR2 (N398, N396, N163);
not NOT1 (N399, N379);
buf BUF1 (N400, N388);
or OR3 (N401, N394, N231, N166);
nor NOR2 (N402, N400, N345);
nand NAND2 (N403, N401, N323);
buf BUF1 (N404, N403);
nor NOR2 (N405, N395, N388);
xor XOR2 (N406, N399, N251);
nor NOR3 (N407, N404, N17, N257);
xor XOR2 (N408, N398, N4);
nand NAND2 (N409, N397, N255);
not NOT1 (N410, N405);
and AND3 (N411, N389, N30, N369);
nor NOR3 (N412, N409, N201, N351);
not NOT1 (N413, N393);
xor XOR2 (N414, N406, N65);
or OR3 (N415, N410, N30, N262);
nor NOR4 (N416, N414, N307, N297, N131);
or OR3 (N417, N413, N145, N270);
or OR2 (N418, N407, N396);
or OR3 (N419, N417, N33, N294);
or OR3 (N420, N415, N116, N63);
and AND4 (N421, N420, N11, N134, N147);
not NOT1 (N422, N418);
nand NAND3 (N423, N411, N170, N367);
xor XOR2 (N424, N402, N31);
nand NAND3 (N425, N424, N132, N136);
not NOT1 (N426, N421);
nand NAND4 (N427, N412, N39, N283, N129);
nor NOR3 (N428, N423, N58, N251);
nand NAND4 (N429, N419, N327, N297, N105);
nor NOR3 (N430, N408, N423, N26);
or OR2 (N431, N429, N111);
and AND4 (N432, N377, N171, N94, N384);
and AND2 (N433, N425, N368);
xor XOR2 (N434, N428, N292);
nand NAND4 (N435, N391, N354, N220, N133);
xor XOR2 (N436, N426, N89);
and AND4 (N437, N422, N355, N335, N203);
buf BUF1 (N438, N432);
or OR4 (N439, N435, N7, N290, N211);
nor NOR2 (N440, N439, N410);
nand NAND4 (N441, N434, N195, N294, N104);
nand NAND2 (N442, N441, N290);
or OR2 (N443, N436, N86);
buf BUF1 (N444, N438);
buf BUF1 (N445, N444);
or OR3 (N446, N433, N95, N259);
xor XOR2 (N447, N446, N78);
and AND3 (N448, N430, N60, N266);
buf BUF1 (N449, N440);
xor XOR2 (N450, N443, N446);
not NOT1 (N451, N450);
buf BUF1 (N452, N442);
xor XOR2 (N453, N452, N388);
nor NOR3 (N454, N447, N179, N213);
not NOT1 (N455, N416);
buf BUF1 (N456, N449);
xor XOR2 (N457, N451, N203);
nor NOR4 (N458, N453, N285, N10, N433);
nor NOR3 (N459, N427, N77, N330);
xor XOR2 (N460, N454, N192);
nor NOR3 (N461, N455, N149, N430);
xor XOR2 (N462, N457, N183);
buf BUF1 (N463, N458);
buf BUF1 (N464, N456);
not NOT1 (N465, N448);
xor XOR2 (N466, N462, N392);
nor NOR4 (N467, N431, N410, N92, N277);
not NOT1 (N468, N467);
or OR4 (N469, N468, N199, N335, N83);
nand NAND2 (N470, N464, N259);
and AND3 (N471, N470, N389, N433);
and AND4 (N472, N466, N187, N404, N213);
nand NAND3 (N473, N471, N111, N119);
nand NAND2 (N474, N461, N175);
xor XOR2 (N475, N472, N127);
nand NAND3 (N476, N465, N8, N307);
xor XOR2 (N477, N459, N188);
nand NAND4 (N478, N473, N211, N129, N431);
nor NOR4 (N479, N437, N398, N283, N370);
and AND3 (N480, N445, N467, N253);
nor NOR2 (N481, N479, N411);
nand NAND4 (N482, N474, N343, N407, N225);
nand NAND4 (N483, N460, N145, N11, N198);
xor XOR2 (N484, N480, N452);
nand NAND4 (N485, N469, N82, N107, N327);
xor XOR2 (N486, N463, N56);
nor NOR4 (N487, N475, N156, N4, N346);
buf BUF1 (N488, N484);
and AND2 (N489, N485, N442);
nand NAND3 (N490, N476, N221, N27);
buf BUF1 (N491, N486);
or OR3 (N492, N478, N260, N428);
buf BUF1 (N493, N492);
or OR3 (N494, N488, N266, N114);
or OR2 (N495, N477, N121);
xor XOR2 (N496, N483, N176);
xor XOR2 (N497, N496, N30);
buf BUF1 (N498, N481);
or OR3 (N499, N494, N33, N137);
and AND3 (N500, N497, N211, N409);
nand NAND2 (N501, N491, N351);
not NOT1 (N502, N487);
nor NOR3 (N503, N500, N343, N103);
and AND2 (N504, N489, N497);
or OR2 (N505, N501, N298);
nor NOR3 (N506, N498, N312, N225);
and AND2 (N507, N505, N391);
or OR3 (N508, N506, N98, N267);
or OR4 (N509, N507, N239, N315, N322);
or OR3 (N510, N502, N451, N395);
not NOT1 (N511, N509);
nor NOR3 (N512, N511, N508, N350);
or OR2 (N513, N310, N370);
not NOT1 (N514, N482);
nand NAND2 (N515, N503, N187);
nand NAND3 (N516, N514, N402, N306);
not NOT1 (N517, N499);
not NOT1 (N518, N512);
and AND3 (N519, N504, N302, N217);
xor XOR2 (N520, N513, N139);
not NOT1 (N521, N495);
xor XOR2 (N522, N493, N27);
not NOT1 (N523, N522);
not NOT1 (N524, N523);
buf BUF1 (N525, N516);
or OR3 (N526, N515, N360, N33);
or OR2 (N527, N519, N149);
and AND2 (N528, N527, N222);
nand NAND4 (N529, N524, N170, N244, N342);
nand NAND4 (N530, N518, N194, N285, N451);
xor XOR2 (N531, N521, N229);
and AND4 (N532, N531, N228, N282, N281);
not NOT1 (N533, N530);
nand NAND3 (N534, N517, N142, N196);
not NOT1 (N535, N526);
and AND4 (N536, N534, N347, N200, N259);
nand NAND3 (N537, N520, N418, N21);
not NOT1 (N538, N535);
and AND2 (N539, N538, N103);
buf BUF1 (N540, N533);
nand NAND2 (N541, N490, N148);
nand NAND2 (N542, N541, N183);
and AND3 (N543, N539, N341, N442);
not NOT1 (N544, N543);
or OR4 (N545, N537, N264, N179, N196);
buf BUF1 (N546, N529);
nand NAND4 (N547, N546, N546, N92, N428);
nand NAND3 (N548, N536, N366, N291);
buf BUF1 (N549, N545);
buf BUF1 (N550, N540);
and AND3 (N551, N542, N11, N71);
or OR4 (N552, N528, N164, N366, N289);
and AND2 (N553, N549, N306);
nor NOR2 (N554, N552, N211);
and AND3 (N555, N548, N329, N471);
nor NOR3 (N556, N544, N55, N531);
nor NOR3 (N557, N532, N1, N234);
nor NOR3 (N558, N554, N94, N224);
nor NOR4 (N559, N558, N366, N329, N316);
or OR4 (N560, N557, N461, N6, N163);
and AND2 (N561, N560, N213);
buf BUF1 (N562, N550);
nand NAND3 (N563, N559, N549, N214);
and AND4 (N564, N547, N116, N251, N381);
buf BUF1 (N565, N510);
and AND4 (N566, N561, N254, N145, N108);
nand NAND3 (N567, N564, N505, N390);
xor XOR2 (N568, N556, N33);
nand NAND4 (N569, N553, N346, N320, N444);
buf BUF1 (N570, N569);
nand NAND3 (N571, N562, N490, N404);
nand NAND4 (N572, N525, N220, N512, N270);
nor NOR4 (N573, N571, N511, N359, N65);
or OR4 (N574, N551, N115, N374, N100);
nor NOR3 (N575, N572, N92, N512);
nand NAND2 (N576, N574, N313);
buf BUF1 (N577, N567);
nor NOR2 (N578, N565, N235);
and AND3 (N579, N570, N530, N456);
xor XOR2 (N580, N563, N499);
xor XOR2 (N581, N580, N126);
not NOT1 (N582, N579);
xor XOR2 (N583, N568, N167);
not NOT1 (N584, N577);
and AND4 (N585, N573, N383, N302, N13);
xor XOR2 (N586, N581, N569);
nor NOR4 (N587, N585, N331, N150, N419);
xor XOR2 (N588, N583, N532);
buf BUF1 (N589, N586);
xor XOR2 (N590, N576, N302);
nor NOR2 (N591, N588, N120);
nand NAND4 (N592, N575, N440, N427, N137);
nor NOR2 (N593, N589, N321);
buf BUF1 (N594, N566);
xor XOR2 (N595, N591, N152);
not NOT1 (N596, N590);
and AND2 (N597, N595, N313);
and AND3 (N598, N587, N27, N293);
not NOT1 (N599, N596);
not NOT1 (N600, N593);
not NOT1 (N601, N600);
and AND2 (N602, N601, N128);
or OR3 (N603, N597, N298, N17);
buf BUF1 (N604, N602);
and AND4 (N605, N598, N285, N337, N126);
and AND2 (N606, N594, N226);
and AND3 (N607, N599, N99, N185);
nor NOR4 (N608, N578, N274, N352, N595);
or OR2 (N609, N584, N155);
buf BUF1 (N610, N604);
or OR4 (N611, N592, N187, N26, N450);
nor NOR3 (N612, N606, N288, N498);
or OR4 (N613, N607, N523, N98, N600);
nor NOR4 (N614, N582, N392, N597, N62);
or OR4 (N615, N611, N176, N63, N229);
buf BUF1 (N616, N609);
or OR3 (N617, N614, N227, N544);
not NOT1 (N618, N603);
and AND2 (N619, N608, N518);
nand NAND2 (N620, N613, N7);
not NOT1 (N621, N620);
or OR3 (N622, N610, N503, N449);
not NOT1 (N623, N615);
or OR4 (N624, N621, N176, N140, N581);
or OR2 (N625, N617, N227);
not NOT1 (N626, N619);
and AND2 (N627, N623, N296);
buf BUF1 (N628, N626);
not NOT1 (N629, N612);
buf BUF1 (N630, N616);
or OR4 (N631, N630, N15, N497, N391);
nand NAND2 (N632, N629, N310);
or OR4 (N633, N555, N374, N147, N532);
xor XOR2 (N634, N633, N620);
buf BUF1 (N635, N625);
and AND3 (N636, N628, N341, N510);
nand NAND4 (N637, N605, N394, N381, N348);
buf BUF1 (N638, N622);
not NOT1 (N639, N636);
not NOT1 (N640, N634);
buf BUF1 (N641, N632);
xor XOR2 (N642, N635, N586);
nand NAND4 (N643, N641, N445, N131, N136);
not NOT1 (N644, N618);
xor XOR2 (N645, N640, N245);
or OR2 (N646, N637, N449);
nand NAND3 (N647, N644, N41, N215);
nor NOR4 (N648, N624, N450, N645, N550);
xor XOR2 (N649, N45, N57);
not NOT1 (N650, N649);
not NOT1 (N651, N627);
buf BUF1 (N652, N631);
nor NOR4 (N653, N648, N490, N137, N371);
xor XOR2 (N654, N647, N487);
not NOT1 (N655, N639);
nand NAND2 (N656, N646, N173);
buf BUF1 (N657, N653);
xor XOR2 (N658, N638, N613);
xor XOR2 (N659, N656, N160);
nand NAND3 (N660, N642, N245, N445);
nand NAND2 (N661, N657, N5);
or OR2 (N662, N650, N644);
nor NOR4 (N663, N658, N51, N397, N382);
xor XOR2 (N664, N651, N563);
xor XOR2 (N665, N652, N54);
nand NAND2 (N666, N661, N620);
or OR3 (N667, N643, N101, N374);
nand NAND4 (N668, N654, N145, N508, N305);
nand NAND4 (N669, N664, N583, N108, N67);
buf BUF1 (N670, N663);
not NOT1 (N671, N659);
and AND4 (N672, N662, N624, N65, N113);
or OR4 (N673, N669, N652, N381, N294);
and AND4 (N674, N655, N322, N278, N68);
and AND3 (N675, N668, N616, N608);
nand NAND3 (N676, N673, N71, N5);
nand NAND4 (N677, N666, N12, N530, N133);
nor NOR4 (N678, N672, N662, N57, N608);
buf BUF1 (N679, N674);
buf BUF1 (N680, N665);
nor NOR3 (N681, N676, N15, N208);
xor XOR2 (N682, N667, N249);
not NOT1 (N683, N679);
nand NAND3 (N684, N680, N74, N528);
not NOT1 (N685, N670);
nor NOR4 (N686, N685, N570, N163, N486);
xor XOR2 (N687, N677, N20);
xor XOR2 (N688, N660, N138);
and AND2 (N689, N681, N101);
nor NOR3 (N690, N688, N591, N103);
nand NAND3 (N691, N687, N488, N261);
nand NAND3 (N692, N690, N45, N103);
or OR3 (N693, N678, N504, N668);
and AND4 (N694, N692, N464, N409, N262);
xor XOR2 (N695, N683, N677);
xor XOR2 (N696, N691, N363);
or OR4 (N697, N675, N421, N374, N44);
nand NAND3 (N698, N671, N127, N555);
nor NOR3 (N699, N696, N122, N672);
or OR4 (N700, N694, N484, N194, N15);
xor XOR2 (N701, N684, N275);
nand NAND4 (N702, N701, N348, N473, N531);
buf BUF1 (N703, N693);
and AND2 (N704, N703, N30);
xor XOR2 (N705, N695, N51);
nand NAND4 (N706, N705, N501, N130, N10);
not NOT1 (N707, N698);
not NOT1 (N708, N707);
xor XOR2 (N709, N686, N436);
not NOT1 (N710, N689);
xor XOR2 (N711, N682, N704);
nand NAND4 (N712, N12, N560, N527, N574);
not NOT1 (N713, N702);
buf BUF1 (N714, N710);
or OR3 (N715, N711, N243, N33);
nand NAND2 (N716, N706, N152);
and AND4 (N717, N709, N490, N174, N362);
and AND3 (N718, N712, N36, N172);
and AND3 (N719, N713, N53, N365);
nor NOR2 (N720, N718, N167);
and AND4 (N721, N719, N568, N403, N689);
nand NAND4 (N722, N714, N36, N660, N277);
and AND3 (N723, N697, N571, N119);
nand NAND3 (N724, N715, N634, N141);
nor NOR4 (N725, N716, N1, N20, N657);
not NOT1 (N726, N720);
or OR3 (N727, N717, N130, N196);
or OR2 (N728, N700, N3);
buf BUF1 (N729, N726);
nand NAND4 (N730, N722, N714, N691, N57);
and AND2 (N731, N725, N424);
and AND3 (N732, N723, N82, N183);
and AND2 (N733, N731, N232);
nor NOR2 (N734, N729, N169);
not NOT1 (N735, N708);
and AND2 (N736, N734, N621);
nor NOR4 (N737, N699, N81, N660, N565);
not NOT1 (N738, N732);
nand NAND3 (N739, N738, N128, N436);
nand NAND3 (N740, N728, N224, N219);
nor NOR4 (N741, N735, N606, N201, N309);
buf BUF1 (N742, N736);
nor NOR4 (N743, N737, N240, N145, N497);
xor XOR2 (N744, N741, N2);
buf BUF1 (N745, N727);
nor NOR2 (N746, N744, N236);
not NOT1 (N747, N724);
not NOT1 (N748, N740);
or OR3 (N749, N743, N441, N79);
buf BUF1 (N750, N742);
buf BUF1 (N751, N730);
xor XOR2 (N752, N751, N138);
and AND3 (N753, N749, N199, N517);
buf BUF1 (N754, N752);
nand NAND3 (N755, N733, N75, N73);
xor XOR2 (N756, N753, N215);
nand NAND2 (N757, N754, N335);
not NOT1 (N758, N750);
buf BUF1 (N759, N721);
and AND2 (N760, N739, N391);
not NOT1 (N761, N758);
not NOT1 (N762, N748);
or OR3 (N763, N756, N488, N512);
xor XOR2 (N764, N760, N253);
nand NAND2 (N765, N763, N67);
nor NOR3 (N766, N755, N476, N454);
not NOT1 (N767, N762);
xor XOR2 (N768, N757, N445);
and AND4 (N769, N745, N575, N641, N2);
nand NAND3 (N770, N759, N146, N657);
or OR2 (N771, N746, N90);
and AND2 (N772, N771, N120);
or OR4 (N773, N766, N382, N535, N195);
or OR2 (N774, N772, N765);
buf BUF1 (N775, N523);
nor NOR4 (N776, N774, N771, N132, N207);
nand NAND3 (N777, N773, N604, N306);
not NOT1 (N778, N770);
and AND4 (N779, N764, N656, N157, N619);
and AND4 (N780, N747, N43, N165, N137);
nor NOR4 (N781, N778, N573, N275, N238);
nor NOR2 (N782, N776, N390);
buf BUF1 (N783, N781);
not NOT1 (N784, N761);
not NOT1 (N785, N768);
xor XOR2 (N786, N775, N549);
nand NAND3 (N787, N767, N575, N120);
or OR2 (N788, N779, N600);
and AND3 (N789, N786, N466, N257);
and AND2 (N790, N784, N58);
and AND3 (N791, N787, N760, N667);
not NOT1 (N792, N791);
buf BUF1 (N793, N788);
or OR4 (N794, N792, N20, N491, N362);
buf BUF1 (N795, N782);
or OR2 (N796, N795, N479);
and AND4 (N797, N769, N366, N437, N681);
not NOT1 (N798, N780);
nand NAND2 (N799, N796, N139);
not NOT1 (N800, N790);
buf BUF1 (N801, N797);
or OR3 (N802, N798, N207, N53);
nor NOR3 (N803, N789, N666, N336);
nand NAND4 (N804, N794, N84, N787, N216);
nor NOR3 (N805, N801, N160, N355);
not NOT1 (N806, N805);
xor XOR2 (N807, N793, N263);
xor XOR2 (N808, N802, N384);
buf BUF1 (N809, N785);
or OR3 (N810, N803, N181, N586);
nor NOR2 (N811, N804, N379);
nor NOR3 (N812, N783, N175, N378);
nor NOR3 (N813, N811, N113, N244);
and AND3 (N814, N808, N325, N256);
nand NAND4 (N815, N813, N703, N206, N594);
nand NAND2 (N816, N806, N65);
or OR2 (N817, N777, N645);
buf BUF1 (N818, N810);
nor NOR4 (N819, N815, N631, N633, N322);
or OR2 (N820, N819, N126);
or OR2 (N821, N820, N681);
xor XOR2 (N822, N821, N35);
xor XOR2 (N823, N817, N53);
buf BUF1 (N824, N814);
buf BUF1 (N825, N822);
or OR2 (N826, N807, N55);
nor NOR4 (N827, N799, N382, N269, N102);
and AND3 (N828, N818, N58, N48);
buf BUF1 (N829, N825);
and AND2 (N830, N812, N676);
not NOT1 (N831, N800);
nand NAND4 (N832, N831, N733, N35, N713);
or OR2 (N833, N827, N408);
not NOT1 (N834, N809);
nand NAND3 (N835, N834, N1, N249);
not NOT1 (N836, N833);
buf BUF1 (N837, N826);
or OR3 (N838, N837, N706, N573);
or OR3 (N839, N823, N327, N187);
nor NOR3 (N840, N835, N335, N420);
xor XOR2 (N841, N829, N490);
xor XOR2 (N842, N828, N180);
buf BUF1 (N843, N839);
buf BUF1 (N844, N840);
buf BUF1 (N845, N842);
nor NOR4 (N846, N843, N555, N97, N158);
xor XOR2 (N847, N845, N765);
xor XOR2 (N848, N838, N427);
nor NOR2 (N849, N841, N96);
nor NOR4 (N850, N846, N111, N584, N726);
not NOT1 (N851, N836);
nand NAND3 (N852, N849, N212, N739);
or OR3 (N853, N830, N716, N199);
nor NOR3 (N854, N816, N759, N261);
buf BUF1 (N855, N848);
xor XOR2 (N856, N824, N318);
not NOT1 (N857, N852);
nand NAND2 (N858, N844, N127);
not NOT1 (N859, N853);
buf BUF1 (N860, N850);
nand NAND4 (N861, N860, N789, N222, N250);
xor XOR2 (N862, N851, N106);
nand NAND3 (N863, N861, N784, N580);
and AND4 (N864, N857, N403, N633, N8);
nand NAND2 (N865, N862, N347);
xor XOR2 (N866, N859, N484);
and AND3 (N867, N847, N349, N123);
buf BUF1 (N868, N866);
nand NAND2 (N869, N865, N453);
and AND2 (N870, N856, N405);
not NOT1 (N871, N858);
nor NOR2 (N872, N871, N280);
nand NAND2 (N873, N872, N322);
nor NOR4 (N874, N873, N45, N675, N32);
buf BUF1 (N875, N864);
nand NAND2 (N876, N868, N646);
nand NAND3 (N877, N875, N171, N42);
nand NAND4 (N878, N854, N668, N552, N217);
nand NAND4 (N879, N877, N482, N839, N681);
not NOT1 (N880, N867);
nor NOR2 (N881, N855, N824);
xor XOR2 (N882, N880, N705);
nand NAND3 (N883, N876, N182, N255);
and AND3 (N884, N874, N671, N432);
or OR2 (N885, N869, N80);
nor NOR2 (N886, N870, N618);
nor NOR4 (N887, N883, N309, N716, N538);
buf BUF1 (N888, N863);
or OR3 (N889, N882, N685, N233);
nor NOR4 (N890, N887, N391, N48, N544);
nor NOR2 (N891, N881, N772);
buf BUF1 (N892, N890);
nor NOR2 (N893, N889, N862);
buf BUF1 (N894, N893);
xor XOR2 (N895, N894, N653);
nor NOR4 (N896, N878, N108, N269, N251);
nand NAND3 (N897, N879, N855, N582);
nor NOR4 (N898, N895, N552, N154, N262);
and AND2 (N899, N888, N84);
nand NAND3 (N900, N886, N340, N49);
xor XOR2 (N901, N885, N738);
buf BUF1 (N902, N892);
or OR2 (N903, N900, N109);
xor XOR2 (N904, N891, N861);
nand NAND3 (N905, N898, N830, N551);
xor XOR2 (N906, N901, N192);
and AND3 (N907, N905, N598, N597);
not NOT1 (N908, N904);
xor XOR2 (N909, N899, N144);
and AND2 (N910, N903, N854);
or OR4 (N911, N909, N599, N383, N527);
xor XOR2 (N912, N832, N50);
buf BUF1 (N913, N906);
buf BUF1 (N914, N908);
or OR3 (N915, N913, N715, N735);
endmodule