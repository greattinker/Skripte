// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16;

output N711,N707,N713,N710,N712,N709,N714,N715,N704,N716;

or OR2 (N17, N13, N1);
nand NAND2 (N18, N8, N6);
and AND3 (N19, N1, N7, N14);
not NOT1 (N20, N14);
not NOT1 (N21, N16);
xor XOR2 (N22, N16, N13);
buf BUF1 (N23, N8);
nor NOR4 (N24, N4, N9, N22, N13);
nor NOR2 (N25, N5, N8);
or OR3 (N26, N5, N2, N19);
not NOT1 (N27, N5);
not NOT1 (N28, N9);
not NOT1 (N29, N24);
not NOT1 (N30, N17);
nor NOR3 (N31, N28, N20, N28);
nand NAND3 (N32, N31, N9, N28);
not NOT1 (N33, N12);
nor NOR3 (N34, N18, N13, N28);
xor XOR2 (N35, N34, N27);
and AND4 (N36, N34, N31, N12, N13);
and AND4 (N37, N30, N8, N2, N24);
nand NAND4 (N38, N32, N7, N4, N13);
buf BUF1 (N39, N36);
nand NAND4 (N40, N39, N30, N21, N36);
nor NOR3 (N41, N26, N33, N32);
not NOT1 (N42, N26);
nand NAND4 (N43, N30, N32, N20, N22);
nand NAND4 (N44, N43, N37, N8, N8);
xor XOR2 (N45, N42, N6);
xor XOR2 (N46, N32, N33);
not NOT1 (N47, N25);
and AND2 (N48, N23, N47);
xor XOR2 (N49, N21, N41);
xor XOR2 (N50, N7, N14);
xor XOR2 (N51, N35, N20);
and AND2 (N52, N45, N25);
not NOT1 (N53, N40);
nand NAND2 (N54, N48, N12);
buf BUF1 (N55, N46);
xor XOR2 (N56, N44, N8);
xor XOR2 (N57, N38, N22);
xor XOR2 (N58, N52, N14);
not NOT1 (N59, N51);
nor NOR3 (N60, N54, N42, N5);
buf BUF1 (N61, N58);
not NOT1 (N62, N60);
nand NAND2 (N63, N29, N9);
xor XOR2 (N64, N59, N25);
not NOT1 (N65, N63);
xor XOR2 (N66, N49, N44);
and AND3 (N67, N53, N40, N21);
buf BUF1 (N68, N66);
not NOT1 (N69, N64);
not NOT1 (N70, N55);
not NOT1 (N71, N61);
xor XOR2 (N72, N67, N17);
and AND3 (N73, N50, N58, N39);
nor NOR2 (N74, N72, N31);
not NOT1 (N75, N68);
not NOT1 (N76, N70);
nor NOR3 (N77, N69, N45, N15);
not NOT1 (N78, N56);
buf BUF1 (N79, N76);
not NOT1 (N80, N75);
not NOT1 (N81, N77);
xor XOR2 (N82, N57, N53);
xor XOR2 (N83, N81, N1);
or OR4 (N84, N65, N44, N27, N56);
not NOT1 (N85, N62);
or OR4 (N86, N84, N78, N61, N73);
buf BUF1 (N87, N86);
or OR4 (N88, N70, N55, N79, N2);
nor NOR2 (N89, N24, N11);
nand NAND2 (N90, N68, N61);
and AND3 (N91, N90, N61, N36);
buf BUF1 (N92, N88);
not NOT1 (N93, N71);
not NOT1 (N94, N83);
nor NOR3 (N95, N92, N77, N1);
and AND4 (N96, N80, N81, N50, N30);
buf BUF1 (N97, N91);
xor XOR2 (N98, N96, N28);
buf BUF1 (N99, N94);
nand NAND2 (N100, N95, N93);
nand NAND3 (N101, N63, N61, N1);
not NOT1 (N102, N100);
xor XOR2 (N103, N101, N74);
and AND2 (N104, N30, N65);
buf BUF1 (N105, N103);
nand NAND3 (N106, N87, N104, N27);
xor XOR2 (N107, N27, N24);
or OR2 (N108, N98, N56);
nor NOR3 (N109, N97, N76, N59);
nor NOR3 (N110, N106, N91, N57);
not NOT1 (N111, N89);
nor NOR2 (N112, N107, N12);
nand NAND3 (N113, N105, N50, N5);
and AND3 (N114, N112, N59, N67);
or OR3 (N115, N82, N7, N41);
buf BUF1 (N116, N109);
not NOT1 (N117, N108);
or OR2 (N118, N115, N76);
not NOT1 (N119, N99);
or OR4 (N120, N110, N111, N10, N82);
nor NOR4 (N121, N115, N110, N100, N50);
and AND3 (N122, N118, N47, N109);
xor XOR2 (N123, N116, N9);
buf BUF1 (N124, N113);
and AND3 (N125, N117, N66, N76);
not NOT1 (N126, N114);
or OR3 (N127, N122, N61, N123);
and AND2 (N128, N98, N25);
nor NOR3 (N129, N102, N80, N23);
not NOT1 (N130, N125);
nand NAND4 (N131, N127, N110, N47, N88);
buf BUF1 (N132, N124);
not NOT1 (N133, N121);
or OR2 (N134, N128, N7);
xor XOR2 (N135, N129, N26);
nor NOR2 (N136, N85, N56);
or OR3 (N137, N126, N45, N40);
xor XOR2 (N138, N136, N49);
nand NAND4 (N139, N135, N3, N123, N4);
xor XOR2 (N140, N119, N104);
xor XOR2 (N141, N131, N55);
and AND2 (N142, N134, N37);
or OR3 (N143, N132, N76, N123);
xor XOR2 (N144, N133, N85);
not NOT1 (N145, N120);
buf BUF1 (N146, N140);
nor NOR2 (N147, N146, N113);
nand NAND2 (N148, N142, N18);
buf BUF1 (N149, N147);
buf BUF1 (N150, N139);
xor XOR2 (N151, N137, N51);
nand NAND2 (N152, N149, N121);
xor XOR2 (N153, N152, N139);
or OR3 (N154, N143, N132, N30);
buf BUF1 (N155, N138);
or OR2 (N156, N144, N70);
nand NAND2 (N157, N145, N118);
nor NOR4 (N158, N154, N98, N143, N134);
or OR4 (N159, N158, N119, N20, N34);
not NOT1 (N160, N148);
or OR3 (N161, N155, N47, N106);
xor XOR2 (N162, N153, N150);
nor NOR4 (N163, N19, N159, N130, N153);
not NOT1 (N164, N71);
buf BUF1 (N165, N65);
not NOT1 (N166, N141);
and AND3 (N167, N163, N88, N134);
buf BUF1 (N168, N161);
nand NAND2 (N169, N167, N44);
buf BUF1 (N170, N164);
or OR4 (N171, N165, N106, N18, N45);
not NOT1 (N172, N168);
not NOT1 (N173, N170);
not NOT1 (N174, N169);
xor XOR2 (N175, N174, N15);
not NOT1 (N176, N173);
nor NOR3 (N177, N160, N122, N125);
buf BUF1 (N178, N162);
and AND2 (N179, N175, N143);
nand NAND4 (N180, N178, N62, N59, N10);
and AND4 (N181, N179, N110, N73, N110);
nor NOR3 (N182, N176, N142, N94);
xor XOR2 (N183, N180, N18);
nor NOR3 (N184, N177, N8, N25);
buf BUF1 (N185, N156);
nor NOR3 (N186, N181, N108, N182);
buf BUF1 (N187, N138);
xor XOR2 (N188, N185, N174);
or OR4 (N189, N157, N91, N60, N66);
xor XOR2 (N190, N189, N83);
buf BUF1 (N191, N151);
and AND4 (N192, N191, N60, N67, N118);
nor NOR3 (N193, N187, N61, N69);
nand NAND4 (N194, N183, N103, N184, N123);
nor NOR3 (N195, N182, N42, N72);
nand NAND2 (N196, N171, N40);
xor XOR2 (N197, N192, N102);
nand NAND4 (N198, N197, N21, N45, N69);
not NOT1 (N199, N190);
or OR4 (N200, N196, N155, N89, N180);
and AND3 (N201, N200, N49, N27);
nor NOR3 (N202, N186, N66, N59);
xor XOR2 (N203, N198, N156);
not NOT1 (N204, N188);
or OR3 (N205, N202, N101, N30);
and AND4 (N206, N172, N138, N13, N148);
and AND3 (N207, N201, N126, N193);
nand NAND2 (N208, N16, N153);
buf BUF1 (N209, N205);
buf BUF1 (N210, N206);
nor NOR2 (N211, N204, N47);
not NOT1 (N212, N166);
not NOT1 (N213, N208);
buf BUF1 (N214, N211);
nor NOR3 (N215, N209, N177, N88);
nor NOR4 (N216, N207, N86, N58, N210);
buf BUF1 (N217, N176);
xor XOR2 (N218, N217, N129);
nor NOR3 (N219, N215, N69, N186);
xor XOR2 (N220, N194, N160);
xor XOR2 (N221, N203, N91);
buf BUF1 (N222, N216);
nand NAND4 (N223, N219, N11, N141, N26);
and AND3 (N224, N223, N21, N148);
nor NOR2 (N225, N199, N193);
or OR2 (N226, N222, N88);
xor XOR2 (N227, N218, N88);
not NOT1 (N228, N220);
or OR2 (N229, N212, N62);
nand NAND2 (N230, N225, N61);
xor XOR2 (N231, N229, N1);
or OR3 (N232, N224, N122, N119);
not NOT1 (N233, N221);
xor XOR2 (N234, N233, N226);
xor XOR2 (N235, N69, N7);
nand NAND2 (N236, N228, N25);
buf BUF1 (N237, N227);
buf BUF1 (N238, N234);
or OR4 (N239, N237, N174, N17, N167);
nand NAND2 (N240, N195, N62);
nor NOR2 (N241, N213, N140);
or OR4 (N242, N214, N85, N18, N165);
xor XOR2 (N243, N242, N219);
nor NOR4 (N244, N232, N213, N128, N38);
nor NOR2 (N245, N240, N186);
xor XOR2 (N246, N239, N241);
buf BUF1 (N247, N72);
nor NOR4 (N248, N231, N187, N100, N176);
buf BUF1 (N249, N247);
and AND4 (N250, N246, N131, N54, N143);
and AND4 (N251, N243, N161, N207, N180);
nor NOR3 (N252, N251, N90, N57);
and AND4 (N253, N252, N192, N55, N247);
nor NOR2 (N254, N230, N130);
and AND4 (N255, N248, N156, N201, N36);
or OR2 (N256, N250, N97);
not NOT1 (N257, N245);
buf BUF1 (N258, N244);
not NOT1 (N259, N249);
nand NAND2 (N260, N254, N205);
not NOT1 (N261, N258);
buf BUF1 (N262, N259);
buf BUF1 (N263, N257);
not NOT1 (N264, N238);
and AND3 (N265, N253, N61, N34);
xor XOR2 (N266, N260, N54);
xor XOR2 (N267, N265, N61);
nor NOR3 (N268, N256, N92, N214);
buf BUF1 (N269, N264);
nor NOR4 (N270, N236, N58, N165, N169);
or OR4 (N271, N266, N119, N49, N209);
or OR4 (N272, N268, N79, N135, N265);
buf BUF1 (N273, N269);
xor XOR2 (N274, N255, N43);
buf BUF1 (N275, N271);
and AND3 (N276, N274, N120, N141);
or OR2 (N277, N261, N256);
buf BUF1 (N278, N275);
and AND2 (N279, N235, N202);
not NOT1 (N280, N278);
not NOT1 (N281, N267);
buf BUF1 (N282, N270);
buf BUF1 (N283, N262);
nor NOR4 (N284, N282, N275, N81, N6);
and AND3 (N285, N273, N211, N124);
not NOT1 (N286, N263);
and AND3 (N287, N272, N252, N79);
or OR4 (N288, N285, N264, N7, N44);
or OR4 (N289, N280, N11, N230, N202);
and AND4 (N290, N289, N62, N122, N48);
xor XOR2 (N291, N279, N60);
buf BUF1 (N292, N291);
not NOT1 (N293, N277);
buf BUF1 (N294, N293);
xor XOR2 (N295, N288, N51);
not NOT1 (N296, N283);
nor NOR3 (N297, N292, N261, N114);
or OR4 (N298, N296, N261, N290, N58);
buf BUF1 (N299, N22);
or OR4 (N300, N276, N256, N114, N222);
xor XOR2 (N301, N298, N58);
not NOT1 (N302, N294);
xor XOR2 (N303, N295, N91);
and AND4 (N304, N286, N159, N100, N201);
buf BUF1 (N305, N287);
nand NAND4 (N306, N284, N229, N192, N248);
nor NOR2 (N307, N304, N236);
and AND4 (N308, N307, N271, N98, N221);
nor NOR4 (N309, N306, N208, N281, N219);
nor NOR2 (N310, N208, N269);
and AND4 (N311, N305, N294, N294, N172);
not NOT1 (N312, N302);
nor NOR2 (N313, N310, N46);
not NOT1 (N314, N308);
nand NAND2 (N315, N312, N302);
or OR2 (N316, N303, N82);
and AND4 (N317, N301, N183, N92, N65);
not NOT1 (N318, N309);
or OR3 (N319, N311, N16, N186);
buf BUF1 (N320, N317);
nand NAND2 (N321, N319, N13);
and AND4 (N322, N320, N92, N59, N304);
nand NAND2 (N323, N318, N179);
or OR3 (N324, N316, N173, N177);
not NOT1 (N325, N300);
nand NAND3 (N326, N299, N52, N218);
xor XOR2 (N327, N324, N87);
nor NOR3 (N328, N322, N267, N47);
nor NOR4 (N329, N327, N14, N312, N61);
nand NAND2 (N330, N315, N317);
nor NOR3 (N331, N323, N269, N216);
nand NAND4 (N332, N321, N130, N319, N130);
nand NAND3 (N333, N314, N119, N294);
nor NOR4 (N334, N325, N270, N253, N60);
buf BUF1 (N335, N334);
xor XOR2 (N336, N313, N188);
not NOT1 (N337, N331);
not NOT1 (N338, N335);
buf BUF1 (N339, N338);
and AND4 (N340, N337, N76, N244, N226);
nand NAND2 (N341, N340, N250);
xor XOR2 (N342, N328, N55);
not NOT1 (N343, N341);
nor NOR2 (N344, N333, N140);
xor XOR2 (N345, N326, N261);
nand NAND2 (N346, N345, N121);
or OR2 (N347, N332, N266);
nand NAND2 (N348, N344, N312);
buf BUF1 (N349, N343);
buf BUF1 (N350, N348);
buf BUF1 (N351, N350);
nand NAND3 (N352, N349, N187, N280);
buf BUF1 (N353, N330);
xor XOR2 (N354, N336, N132);
and AND4 (N355, N297, N161, N327, N58);
nand NAND4 (N356, N347, N243, N339, N183);
or OR3 (N357, N96, N331, N206);
or OR2 (N358, N351, N128);
buf BUF1 (N359, N342);
nand NAND2 (N360, N357, N83);
not NOT1 (N361, N356);
not NOT1 (N362, N359);
not NOT1 (N363, N353);
nand NAND4 (N364, N329, N43, N140, N59);
xor XOR2 (N365, N358, N108);
not NOT1 (N366, N365);
nor NOR2 (N367, N366, N321);
and AND4 (N368, N352, N227, N8, N250);
and AND2 (N369, N346, N235);
nor NOR4 (N370, N361, N56, N353, N65);
not NOT1 (N371, N370);
xor XOR2 (N372, N360, N319);
buf BUF1 (N373, N371);
nor NOR2 (N374, N363, N112);
buf BUF1 (N375, N355);
nor NOR4 (N376, N373, N252, N332, N67);
and AND4 (N377, N372, N299, N369, N10);
or OR2 (N378, N265, N301);
or OR2 (N379, N367, N287);
nand NAND3 (N380, N377, N379, N268);
xor XOR2 (N381, N78, N361);
nor NOR2 (N382, N380, N363);
xor XOR2 (N383, N374, N230);
nand NAND4 (N384, N375, N382, N341, N50);
nand NAND4 (N385, N346, N324, N352, N322);
and AND3 (N386, N362, N150, N206);
not NOT1 (N387, N364);
xor XOR2 (N388, N381, N172);
and AND3 (N389, N378, N120, N197);
and AND2 (N390, N387, N79);
or OR4 (N391, N354, N115, N158, N329);
xor XOR2 (N392, N383, N211);
and AND2 (N393, N390, N97);
and AND2 (N394, N376, N101);
buf BUF1 (N395, N368);
buf BUF1 (N396, N391);
xor XOR2 (N397, N384, N37);
buf BUF1 (N398, N385);
xor XOR2 (N399, N395, N47);
not NOT1 (N400, N397);
or OR2 (N401, N399, N93);
or OR4 (N402, N396, N240, N82, N249);
nand NAND4 (N403, N398, N360, N13, N177);
not NOT1 (N404, N400);
not NOT1 (N405, N388);
or OR3 (N406, N392, N302, N337);
nand NAND3 (N407, N402, N116, N22);
buf BUF1 (N408, N386);
or OR4 (N409, N403, N271, N393, N332);
nand NAND3 (N410, N219, N242, N327);
nand NAND4 (N411, N405, N246, N352, N48);
nand NAND4 (N412, N410, N349, N371, N162);
and AND3 (N413, N411, N357, N235);
not NOT1 (N414, N412);
buf BUF1 (N415, N406);
nor NOR4 (N416, N389, N406, N213, N284);
nand NAND4 (N417, N404, N36, N397, N256);
and AND2 (N418, N414, N336);
nand NAND2 (N419, N415, N262);
and AND2 (N420, N408, N344);
or OR2 (N421, N407, N124);
nand NAND2 (N422, N417, N333);
nor NOR4 (N423, N420, N107, N293, N88);
nor NOR4 (N424, N418, N26, N3, N156);
nor NOR4 (N425, N423, N228, N145, N205);
nand NAND4 (N426, N421, N210, N94, N184);
not NOT1 (N427, N409);
and AND4 (N428, N401, N22, N118, N237);
buf BUF1 (N429, N428);
nand NAND2 (N430, N429, N300);
buf BUF1 (N431, N425);
not NOT1 (N432, N419);
buf BUF1 (N433, N426);
not NOT1 (N434, N394);
buf BUF1 (N435, N424);
nand NAND2 (N436, N422, N123);
not NOT1 (N437, N431);
buf BUF1 (N438, N427);
xor XOR2 (N439, N430, N300);
buf BUF1 (N440, N435);
and AND3 (N441, N436, N216, N395);
xor XOR2 (N442, N439, N69);
not NOT1 (N443, N434);
and AND4 (N444, N442, N105, N261, N64);
xor XOR2 (N445, N440, N295);
and AND4 (N446, N432, N374, N201, N202);
xor XOR2 (N447, N437, N261);
nand NAND3 (N448, N433, N87, N366);
not NOT1 (N449, N444);
or OR4 (N450, N449, N412, N63, N42);
or OR2 (N451, N447, N387);
buf BUF1 (N452, N443);
or OR3 (N453, N416, N6, N293);
and AND3 (N454, N445, N358, N34);
xor XOR2 (N455, N451, N196);
nor NOR4 (N456, N441, N126, N412, N397);
nand NAND4 (N457, N454, N371, N429, N299);
not NOT1 (N458, N452);
nand NAND2 (N459, N413, N391);
nand NAND2 (N460, N456, N454);
nor NOR2 (N461, N455, N47);
xor XOR2 (N462, N457, N326);
nor NOR4 (N463, N446, N332, N179, N193);
or OR3 (N464, N459, N253, N175);
or OR4 (N465, N460, N115, N78, N136);
xor XOR2 (N466, N462, N375);
or OR3 (N467, N461, N438, N390);
not NOT1 (N468, N254);
nor NOR4 (N469, N463, N75, N458, N400);
and AND3 (N470, N82, N413, N426);
xor XOR2 (N471, N469, N380);
nand NAND4 (N472, N465, N449, N352, N377);
buf BUF1 (N473, N450);
buf BUF1 (N474, N453);
xor XOR2 (N475, N448, N344);
xor XOR2 (N476, N475, N466);
buf BUF1 (N477, N86);
nor NOR2 (N478, N474, N64);
not NOT1 (N479, N472);
buf BUF1 (N480, N467);
or OR4 (N481, N480, N66, N220, N383);
or OR3 (N482, N481, N280, N68);
and AND3 (N483, N468, N279, N424);
or OR3 (N484, N483, N14, N202);
nand NAND3 (N485, N473, N381, N317);
and AND2 (N486, N471, N7);
xor XOR2 (N487, N478, N379);
xor XOR2 (N488, N484, N149);
or OR4 (N489, N486, N120, N271, N166);
buf BUF1 (N490, N489);
nor NOR4 (N491, N476, N287, N214, N218);
not NOT1 (N492, N487);
buf BUF1 (N493, N485);
or OR4 (N494, N477, N219, N22, N312);
not NOT1 (N495, N490);
buf BUF1 (N496, N488);
or OR4 (N497, N493, N431, N257, N85);
or OR4 (N498, N495, N9, N213, N15);
or OR3 (N499, N496, N180, N15);
nand NAND2 (N500, N499, N115);
and AND3 (N501, N470, N284, N234);
buf BUF1 (N502, N500);
or OR4 (N503, N464, N450, N155, N321);
not NOT1 (N504, N503);
nor NOR3 (N505, N491, N420, N260);
not NOT1 (N506, N497);
not NOT1 (N507, N506);
xor XOR2 (N508, N507, N289);
xor XOR2 (N509, N494, N208);
and AND2 (N510, N498, N296);
or OR2 (N511, N509, N84);
buf BUF1 (N512, N508);
and AND2 (N513, N502, N134);
or OR4 (N514, N492, N177, N295, N155);
nand NAND4 (N515, N504, N212, N443, N63);
or OR2 (N516, N512, N85);
buf BUF1 (N517, N514);
and AND4 (N518, N505, N80, N358, N272);
and AND2 (N519, N510, N122);
nor NOR2 (N520, N511, N486);
and AND4 (N521, N482, N163, N452, N483);
and AND4 (N522, N479, N379, N211, N193);
buf BUF1 (N523, N521);
buf BUF1 (N524, N501);
or OR3 (N525, N513, N138, N9);
nand NAND4 (N526, N525, N349, N299, N418);
buf BUF1 (N527, N515);
not NOT1 (N528, N526);
buf BUF1 (N529, N524);
buf BUF1 (N530, N529);
and AND4 (N531, N530, N371, N58, N256);
nor NOR3 (N532, N519, N488, N318);
and AND4 (N533, N532, N169, N13, N191);
and AND4 (N534, N518, N512, N1, N113);
and AND4 (N535, N523, N57, N474, N277);
nand NAND3 (N536, N516, N478, N324);
not NOT1 (N537, N528);
not NOT1 (N538, N527);
or OR2 (N539, N536, N279);
xor XOR2 (N540, N522, N4);
and AND3 (N541, N539, N490, N39);
xor XOR2 (N542, N535, N482);
and AND3 (N543, N534, N71, N389);
buf BUF1 (N544, N542);
buf BUF1 (N545, N520);
and AND2 (N546, N540, N14);
or OR3 (N547, N544, N171, N404);
buf BUF1 (N548, N541);
xor XOR2 (N549, N537, N540);
not NOT1 (N550, N531);
and AND4 (N551, N543, N434, N377, N549);
and AND3 (N552, N318, N316, N168);
xor XOR2 (N553, N538, N550);
and AND2 (N554, N178, N150);
nor NOR3 (N555, N554, N259, N120);
xor XOR2 (N556, N533, N323);
and AND2 (N557, N545, N524);
nor NOR4 (N558, N552, N116, N447, N434);
buf BUF1 (N559, N551);
nor NOR4 (N560, N558, N327, N212, N215);
and AND3 (N561, N555, N131, N321);
nor NOR2 (N562, N556, N545);
buf BUF1 (N563, N517);
nand NAND2 (N564, N548, N415);
not NOT1 (N565, N564);
nor NOR2 (N566, N559, N509);
xor XOR2 (N567, N547, N108);
nand NAND3 (N568, N563, N40, N14);
nor NOR4 (N569, N562, N60, N390, N491);
not NOT1 (N570, N568);
nand NAND3 (N571, N561, N376, N387);
not NOT1 (N572, N553);
or OR2 (N573, N566, N67);
nor NOR4 (N574, N573, N4, N119, N105);
xor XOR2 (N575, N570, N19);
not NOT1 (N576, N572);
and AND2 (N577, N560, N519);
and AND3 (N578, N567, N131, N554);
nor NOR4 (N579, N574, N343, N155, N267);
buf BUF1 (N580, N569);
xor XOR2 (N581, N565, N87);
buf BUF1 (N582, N576);
and AND3 (N583, N581, N354, N275);
xor XOR2 (N584, N579, N329);
nor NOR4 (N585, N571, N104, N445, N345);
nand NAND2 (N586, N583, N465);
xor XOR2 (N587, N584, N101);
xor XOR2 (N588, N580, N315);
xor XOR2 (N589, N582, N235);
or OR3 (N590, N546, N410, N120);
not NOT1 (N591, N578);
or OR2 (N592, N591, N374);
nor NOR3 (N593, N586, N434, N408);
nor NOR2 (N594, N577, N47);
nand NAND2 (N595, N592, N429);
and AND3 (N596, N588, N262, N226);
xor XOR2 (N597, N585, N219);
buf BUF1 (N598, N593);
buf BUF1 (N599, N587);
nand NAND2 (N600, N598, N169);
buf BUF1 (N601, N599);
or OR4 (N602, N590, N560, N86, N296);
buf BUF1 (N603, N596);
and AND3 (N604, N557, N537, N566);
not NOT1 (N605, N603);
xor XOR2 (N606, N601, N587);
buf BUF1 (N607, N606);
or OR3 (N608, N595, N230, N90);
nor NOR3 (N609, N589, N209, N57);
buf BUF1 (N610, N605);
nor NOR3 (N611, N594, N261, N221);
nor NOR4 (N612, N575, N197, N602, N230);
buf BUF1 (N613, N330);
buf BUF1 (N614, N600);
or OR2 (N615, N614, N583);
xor XOR2 (N616, N611, N102);
and AND3 (N617, N597, N523, N28);
nand NAND3 (N618, N609, N217, N579);
not NOT1 (N619, N612);
xor XOR2 (N620, N610, N479);
xor XOR2 (N621, N618, N408);
and AND3 (N622, N616, N388, N251);
xor XOR2 (N623, N604, N83);
or OR3 (N624, N623, N416, N369);
and AND4 (N625, N617, N18, N193, N42);
buf BUF1 (N626, N613);
or OR2 (N627, N615, N592);
and AND3 (N628, N607, N142, N116);
xor XOR2 (N629, N620, N300);
nor NOR4 (N630, N622, N433, N83, N559);
xor XOR2 (N631, N621, N266);
nor NOR4 (N632, N628, N588, N494, N373);
buf BUF1 (N633, N631);
buf BUF1 (N634, N608);
buf BUF1 (N635, N634);
buf BUF1 (N636, N619);
and AND2 (N637, N629, N500);
xor XOR2 (N638, N637, N523);
nand NAND3 (N639, N630, N33, N410);
xor XOR2 (N640, N633, N541);
nor NOR2 (N641, N632, N533);
and AND2 (N642, N635, N271);
and AND4 (N643, N626, N164, N137, N159);
and AND2 (N644, N625, N153);
not NOT1 (N645, N639);
xor XOR2 (N646, N627, N442);
not NOT1 (N647, N646);
or OR3 (N648, N645, N276, N278);
not NOT1 (N649, N641);
xor XOR2 (N650, N636, N4);
or OR4 (N651, N647, N8, N451, N165);
and AND2 (N652, N649, N127);
or OR4 (N653, N642, N75, N45, N309);
not NOT1 (N654, N652);
not NOT1 (N655, N643);
and AND2 (N656, N644, N359);
not NOT1 (N657, N651);
buf BUF1 (N658, N653);
and AND4 (N659, N656, N259, N104, N163);
or OR2 (N660, N648, N253);
not NOT1 (N661, N654);
and AND3 (N662, N660, N382, N654);
or OR2 (N663, N624, N554);
and AND2 (N664, N650, N143);
nor NOR2 (N665, N664, N658);
or OR3 (N666, N413, N605, N397);
xor XOR2 (N667, N657, N55);
buf BUF1 (N668, N655);
nor NOR2 (N669, N667, N174);
not NOT1 (N670, N669);
xor XOR2 (N671, N663, N511);
buf BUF1 (N672, N666);
nand NAND2 (N673, N672, N360);
nor NOR3 (N674, N671, N180, N93);
buf BUF1 (N675, N665);
or OR2 (N676, N670, N314);
nor NOR2 (N677, N674, N313);
buf BUF1 (N678, N638);
xor XOR2 (N679, N659, N342);
not NOT1 (N680, N662);
not NOT1 (N681, N673);
buf BUF1 (N682, N679);
nor NOR3 (N683, N678, N130, N49);
xor XOR2 (N684, N680, N174);
and AND4 (N685, N640, N481, N647, N285);
buf BUF1 (N686, N675);
not NOT1 (N687, N683);
or OR2 (N688, N677, N262);
or OR4 (N689, N682, N327, N215, N462);
buf BUF1 (N690, N661);
nand NAND2 (N691, N687, N154);
buf BUF1 (N692, N689);
nor NOR3 (N693, N688, N299, N308);
and AND4 (N694, N668, N425, N54, N120);
nor NOR4 (N695, N692, N571, N667, N100);
and AND4 (N696, N694, N99, N220, N327);
nor NOR2 (N697, N686, N624);
and AND4 (N698, N695, N203, N241, N93);
not NOT1 (N699, N691);
buf BUF1 (N700, N684);
and AND2 (N701, N697, N185);
or OR2 (N702, N685, N65);
buf BUF1 (N703, N698);
nand NAND2 (N704, N700, N126);
nor NOR2 (N705, N702, N9);
nor NOR4 (N706, N681, N137, N129, N521);
or OR2 (N707, N699, N11);
nor NOR3 (N708, N703, N27, N505);
buf BUF1 (N709, N701);
xor XOR2 (N710, N676, N683);
and AND2 (N711, N708, N573);
nor NOR3 (N712, N705, N193, N339);
not NOT1 (N713, N693);
buf BUF1 (N714, N706);
xor XOR2 (N715, N696, N449);
or OR3 (N716, N690, N581, N322);
endmodule