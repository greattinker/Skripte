// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16;

output N2507,N2515,N2483,N2511,N2498,N2510,N2514,N2474,N2493,N2516;

nor NOR2 (N17, N3, N8);
not NOT1 (N18, N9);
or OR3 (N19, N8, N17, N14);
buf BUF1 (N20, N9);
nand NAND2 (N21, N4, N10);
xor XOR2 (N22, N8, N9);
or OR3 (N23, N9, N16, N16);
nand NAND4 (N24, N17, N11, N13, N19);
nor NOR2 (N25, N14, N12);
buf BUF1 (N26, N4);
and AND2 (N27, N7, N9);
or OR4 (N28, N3, N12, N21, N9);
or OR4 (N29, N4, N10, N18, N25);
xor XOR2 (N30, N27, N11);
or OR4 (N31, N7, N22, N21, N1);
nand NAND4 (N32, N30, N27, N8, N23);
and AND4 (N33, N32, N25, N23, N22);
buf BUF1 (N34, N20);
xor XOR2 (N35, N30, N28);
xor XOR2 (N36, N9, N12);
xor XOR2 (N37, N21, N17);
nor NOR3 (N38, N15, N30, N15);
not NOT1 (N39, N24);
buf BUF1 (N40, N39);
not NOT1 (N41, N34);
xor XOR2 (N42, N33, N10);
buf BUF1 (N43, N36);
xor XOR2 (N44, N26, N17);
buf BUF1 (N45, N31);
or OR2 (N46, N37, N35);
not NOT1 (N47, N24);
nor NOR3 (N48, N38, N31, N21);
not NOT1 (N49, N48);
nand NAND2 (N50, N44, N24);
not NOT1 (N51, N40);
nor NOR2 (N52, N29, N16);
or OR4 (N53, N51, N15, N26, N48);
nor NOR2 (N54, N43, N33);
not NOT1 (N55, N46);
not NOT1 (N56, N41);
not NOT1 (N57, N53);
nor NOR3 (N58, N49, N40, N22);
and AND3 (N59, N54, N26, N39);
xor XOR2 (N60, N57, N45);
nand NAND2 (N61, N7, N53);
or OR2 (N62, N52, N31);
nand NAND2 (N63, N58, N56);
buf BUF1 (N64, N34);
not NOT1 (N65, N63);
and AND4 (N66, N61, N40, N15, N46);
nand NAND3 (N67, N55, N57, N2);
not NOT1 (N68, N66);
not NOT1 (N69, N68);
xor XOR2 (N70, N50, N58);
buf BUF1 (N71, N59);
nand NAND2 (N72, N64, N39);
xor XOR2 (N73, N72, N13);
and AND3 (N74, N67, N15, N6);
or OR4 (N75, N73, N49, N11, N67);
buf BUF1 (N76, N75);
and AND2 (N77, N71, N24);
or OR2 (N78, N74, N31);
not NOT1 (N79, N78);
not NOT1 (N80, N42);
or OR3 (N81, N69, N17, N32);
nand NAND3 (N82, N79, N29, N80);
nand NAND2 (N83, N77, N5);
buf BUF1 (N84, N53);
and AND2 (N85, N76, N44);
xor XOR2 (N86, N62, N43);
and AND3 (N87, N83, N12, N82);
or OR2 (N88, N83, N52);
nor NOR4 (N89, N85, N69, N2, N81);
or OR2 (N90, N30, N70);
nand NAND3 (N91, N54, N49, N42);
nor NOR2 (N92, N87, N42);
and AND2 (N93, N89, N43);
or OR4 (N94, N84, N26, N64, N10);
nor NOR4 (N95, N94, N30, N29, N78);
or OR3 (N96, N90, N29, N72);
buf BUF1 (N97, N92);
not NOT1 (N98, N60);
xor XOR2 (N99, N95, N93);
nor NOR3 (N100, N14, N59, N57);
and AND2 (N101, N91, N12);
nor NOR2 (N102, N47, N38);
not NOT1 (N103, N96);
buf BUF1 (N104, N86);
buf BUF1 (N105, N97);
nor NOR3 (N106, N99, N46, N4);
buf BUF1 (N107, N100);
xor XOR2 (N108, N104, N22);
nor NOR3 (N109, N88, N25, N53);
nand NAND3 (N110, N109, N94, N11);
or OR4 (N111, N65, N45, N56, N82);
buf BUF1 (N112, N101);
nand NAND3 (N113, N106, N90, N104);
nor NOR3 (N114, N111, N75, N58);
buf BUF1 (N115, N110);
not NOT1 (N116, N112);
nor NOR3 (N117, N116, N70, N89);
or OR3 (N118, N108, N54, N5);
not NOT1 (N119, N102);
not NOT1 (N120, N114);
not NOT1 (N121, N118);
or OR4 (N122, N117, N12, N96, N103);
and AND4 (N123, N21, N1, N55, N122);
or OR2 (N124, N110, N31);
nand NAND4 (N125, N107, N43, N56, N119);
buf BUF1 (N126, N83);
not NOT1 (N127, N123);
not NOT1 (N128, N121);
nor NOR2 (N129, N127, N38);
nand NAND3 (N130, N126, N29, N20);
or OR3 (N131, N125, N120, N114);
nor NOR4 (N132, N5, N118, N64, N40);
xor XOR2 (N133, N113, N29);
buf BUF1 (N134, N124);
not NOT1 (N135, N98);
nand NAND2 (N136, N135, N4);
nor NOR3 (N137, N129, N96, N33);
or OR4 (N138, N136, N121, N45, N116);
and AND2 (N139, N134, N13);
nand NAND4 (N140, N137, N81, N32, N70);
and AND4 (N141, N133, N61, N17, N109);
or OR2 (N142, N105, N56);
or OR2 (N143, N128, N141);
buf BUF1 (N144, N1);
nand NAND4 (N145, N142, N9, N128, N109);
not NOT1 (N146, N131);
nand NAND2 (N147, N138, N82);
nor NOR4 (N148, N115, N95, N81, N79);
nand NAND2 (N149, N132, N89);
not NOT1 (N150, N149);
or OR2 (N151, N143, N80);
or OR2 (N152, N150, N40);
xor XOR2 (N153, N139, N124);
nand NAND4 (N154, N145, N29, N120, N34);
buf BUF1 (N155, N130);
or OR2 (N156, N155, N105);
nor NOR3 (N157, N144, N111, N85);
or OR4 (N158, N148, N75, N111, N111);
nor NOR4 (N159, N151, N79, N118, N150);
and AND4 (N160, N157, N151, N121, N106);
buf BUF1 (N161, N147);
xor XOR2 (N162, N159, N2);
and AND4 (N163, N161, N126, N20, N159);
and AND2 (N164, N153, N17);
nand NAND4 (N165, N154, N102, N99, N3);
xor XOR2 (N166, N158, N164);
xor XOR2 (N167, N144, N47);
and AND2 (N168, N167, N115);
and AND4 (N169, N140, N40, N114, N41);
xor XOR2 (N170, N168, N168);
and AND4 (N171, N146, N154, N79, N68);
xor XOR2 (N172, N170, N164);
nor NOR2 (N173, N160, N48);
or OR2 (N174, N169, N49);
buf BUF1 (N175, N165);
buf BUF1 (N176, N152);
xor XOR2 (N177, N162, N62);
nand NAND2 (N178, N172, N132);
and AND4 (N179, N178, N66, N31, N149);
buf BUF1 (N180, N174);
buf BUF1 (N181, N156);
nor NOR2 (N182, N180, N173);
or OR3 (N183, N65, N149, N182);
and AND2 (N184, N52, N7);
nor NOR2 (N185, N171, N107);
xor XOR2 (N186, N176, N160);
xor XOR2 (N187, N185, N79);
nor NOR4 (N188, N181, N122, N63, N164);
buf BUF1 (N189, N179);
and AND3 (N190, N183, N40, N29);
not NOT1 (N191, N187);
and AND3 (N192, N189, N2, N130);
xor XOR2 (N193, N184, N140);
nor NOR2 (N194, N186, N60);
buf BUF1 (N195, N188);
xor XOR2 (N196, N194, N159);
nor NOR2 (N197, N195, N155);
not NOT1 (N198, N190);
and AND4 (N199, N192, N147, N42, N191);
nor NOR2 (N200, N44, N85);
or OR4 (N201, N200, N149, N33, N134);
or OR3 (N202, N196, N54, N196);
buf BUF1 (N203, N166);
and AND4 (N204, N201, N41, N166, N149);
nor NOR2 (N205, N202, N94);
not NOT1 (N206, N204);
buf BUF1 (N207, N197);
nor NOR4 (N208, N175, N3, N117, N57);
not NOT1 (N209, N203);
and AND3 (N210, N206, N90, N162);
xor XOR2 (N211, N193, N201);
not NOT1 (N212, N177);
nor NOR3 (N213, N198, N171, N22);
nand NAND2 (N214, N205, N6);
not NOT1 (N215, N210);
and AND2 (N216, N213, N208);
nand NAND2 (N217, N144, N97);
buf BUF1 (N218, N214);
nor NOR3 (N219, N211, N27, N47);
nor NOR3 (N220, N217, N211, N97);
nand NAND4 (N221, N215, N173, N59, N22);
nor NOR2 (N222, N212, N195);
buf BUF1 (N223, N199);
buf BUF1 (N224, N218);
buf BUF1 (N225, N163);
or OR2 (N226, N220, N82);
and AND2 (N227, N225, N137);
and AND3 (N228, N224, N16, N7);
and AND3 (N229, N216, N143, N174);
not NOT1 (N230, N207);
and AND3 (N231, N226, N204, N184);
xor XOR2 (N232, N229, N13);
buf BUF1 (N233, N219);
buf BUF1 (N234, N209);
or OR4 (N235, N232, N154, N101, N81);
not NOT1 (N236, N235);
buf BUF1 (N237, N236);
and AND4 (N238, N231, N75, N26, N190);
nand NAND2 (N239, N228, N24);
and AND2 (N240, N234, N106);
not NOT1 (N241, N222);
nor NOR3 (N242, N237, N121, N64);
and AND4 (N243, N221, N95, N222, N72);
xor XOR2 (N244, N238, N105);
nor NOR3 (N245, N242, N177, N208);
or OR4 (N246, N240, N5, N23, N174);
and AND2 (N247, N233, N229);
not NOT1 (N248, N244);
nor NOR2 (N249, N223, N36);
xor XOR2 (N250, N239, N11);
nor NOR2 (N251, N243, N153);
xor XOR2 (N252, N247, N150);
buf BUF1 (N253, N249);
and AND2 (N254, N227, N84);
nand NAND4 (N255, N250, N233, N152, N231);
xor XOR2 (N256, N230, N146);
nor NOR4 (N257, N256, N156, N113, N34);
and AND4 (N258, N257, N66, N144, N115);
or OR2 (N259, N246, N188);
nor NOR2 (N260, N241, N5);
nand NAND2 (N261, N255, N46);
buf BUF1 (N262, N252);
nor NOR4 (N263, N253, N167, N146, N228);
xor XOR2 (N264, N254, N230);
nor NOR3 (N265, N262, N207, N160);
xor XOR2 (N266, N258, N191);
nand NAND3 (N267, N251, N206, N231);
buf BUF1 (N268, N266);
not NOT1 (N269, N248);
or OR2 (N270, N265, N206);
not NOT1 (N271, N269);
nand NAND3 (N272, N263, N207, N31);
or OR4 (N273, N261, N187, N42, N177);
or OR3 (N274, N245, N136, N251);
nand NAND3 (N275, N270, N15, N142);
nand NAND4 (N276, N275, N258, N222, N154);
and AND2 (N277, N274, N95);
buf BUF1 (N278, N264);
nand NAND2 (N279, N273, N229);
nor NOR3 (N280, N259, N163, N261);
nand NAND3 (N281, N278, N14, N127);
xor XOR2 (N282, N276, N245);
not NOT1 (N283, N267);
and AND2 (N284, N272, N65);
buf BUF1 (N285, N284);
and AND4 (N286, N260, N157, N190, N280);
xor XOR2 (N287, N238, N59);
or OR4 (N288, N285, N107, N141, N35);
buf BUF1 (N289, N282);
xor XOR2 (N290, N286, N183);
nor NOR3 (N291, N268, N221, N18);
nand NAND3 (N292, N291, N45, N67);
nor NOR2 (N293, N279, N291);
xor XOR2 (N294, N277, N188);
nand NAND4 (N295, N294, N118, N198, N18);
and AND4 (N296, N281, N5, N249, N31);
and AND4 (N297, N293, N151, N253, N286);
xor XOR2 (N298, N271, N9);
nor NOR3 (N299, N295, N198, N20);
xor XOR2 (N300, N289, N212);
buf BUF1 (N301, N290);
xor XOR2 (N302, N292, N14);
xor XOR2 (N303, N298, N206);
and AND2 (N304, N299, N275);
not NOT1 (N305, N302);
buf BUF1 (N306, N283);
or OR2 (N307, N287, N151);
nand NAND2 (N308, N306, N247);
and AND4 (N309, N308, N48, N100, N191);
nor NOR2 (N310, N296, N204);
nor NOR3 (N311, N305, N298, N119);
or OR4 (N312, N297, N124, N266, N103);
buf BUF1 (N313, N309);
nand NAND3 (N314, N313, N6, N166);
xor XOR2 (N315, N310, N27);
nor NOR4 (N316, N315, N152, N70, N315);
and AND3 (N317, N301, N45, N140);
not NOT1 (N318, N300);
buf BUF1 (N319, N314);
xor XOR2 (N320, N303, N121);
buf BUF1 (N321, N311);
nor NOR3 (N322, N318, N117, N85);
and AND3 (N323, N322, N279, N52);
xor XOR2 (N324, N304, N267);
buf BUF1 (N325, N324);
xor XOR2 (N326, N316, N120);
buf BUF1 (N327, N319);
nand NAND2 (N328, N321, N160);
and AND4 (N329, N288, N266, N270, N99);
xor XOR2 (N330, N323, N84);
xor XOR2 (N331, N320, N72);
not NOT1 (N332, N317);
nor NOR2 (N333, N330, N271);
or OR4 (N334, N307, N150, N84, N11);
not NOT1 (N335, N333);
or OR3 (N336, N328, N221, N195);
nand NAND3 (N337, N312, N230, N24);
nor NOR3 (N338, N334, N237, N48);
nor NOR4 (N339, N332, N286, N143, N327);
xor XOR2 (N340, N218, N255);
xor XOR2 (N341, N329, N91);
nand NAND2 (N342, N340, N339);
or OR2 (N343, N45, N265);
or OR4 (N344, N337, N97, N95, N311);
nand NAND3 (N345, N325, N183, N149);
xor XOR2 (N346, N326, N207);
nand NAND3 (N347, N338, N310, N288);
buf BUF1 (N348, N343);
and AND4 (N349, N347, N170, N59, N101);
nand NAND4 (N350, N331, N218, N269, N126);
and AND3 (N351, N349, N17, N196);
xor XOR2 (N352, N344, N136);
buf BUF1 (N353, N351);
nand NAND3 (N354, N352, N19, N352);
or OR4 (N355, N354, N139, N151, N271);
buf BUF1 (N356, N335);
buf BUF1 (N357, N356);
nand NAND4 (N358, N350, N297, N116, N70);
nand NAND2 (N359, N342, N179);
nor NOR3 (N360, N346, N105, N120);
nor NOR4 (N361, N336, N31, N225, N253);
or OR2 (N362, N355, N298);
not NOT1 (N363, N360);
or OR4 (N364, N353, N7, N8, N23);
or OR3 (N365, N361, N71, N166);
or OR2 (N366, N359, N277);
not NOT1 (N367, N366);
or OR2 (N368, N348, N343);
buf BUF1 (N369, N364);
or OR2 (N370, N368, N307);
not NOT1 (N371, N370);
and AND4 (N372, N341, N312, N358, N163);
nand NAND4 (N373, N9, N112, N163, N282);
buf BUF1 (N374, N362);
buf BUF1 (N375, N357);
not NOT1 (N376, N374);
nor NOR4 (N377, N365, N69, N30, N351);
buf BUF1 (N378, N373);
not NOT1 (N379, N345);
or OR3 (N380, N377, N306, N291);
xor XOR2 (N381, N371, N284);
or OR2 (N382, N375, N43);
nor NOR2 (N383, N378, N16);
not NOT1 (N384, N383);
xor XOR2 (N385, N367, N298);
nand NAND4 (N386, N379, N85, N140, N345);
nor NOR3 (N387, N372, N222, N48);
not NOT1 (N388, N387);
xor XOR2 (N389, N382, N192);
not NOT1 (N390, N381);
xor XOR2 (N391, N388, N81);
xor XOR2 (N392, N376, N293);
xor XOR2 (N393, N369, N366);
xor XOR2 (N394, N363, N243);
buf BUF1 (N395, N391);
buf BUF1 (N396, N380);
not NOT1 (N397, N392);
nand NAND4 (N398, N397, N208, N298, N86);
not NOT1 (N399, N384);
and AND3 (N400, N389, N68, N353);
xor XOR2 (N401, N398, N340);
nand NAND2 (N402, N395, N77);
nor NOR2 (N403, N401, N17);
or OR4 (N404, N390, N350, N359, N299);
or OR3 (N405, N394, N328, N254);
not NOT1 (N406, N403);
and AND2 (N407, N385, N258);
buf BUF1 (N408, N406);
not NOT1 (N409, N402);
not NOT1 (N410, N409);
and AND2 (N411, N396, N233);
xor XOR2 (N412, N405, N314);
not NOT1 (N413, N411);
not NOT1 (N414, N386);
buf BUF1 (N415, N393);
not NOT1 (N416, N412);
nor NOR3 (N417, N415, N135, N169);
nor NOR2 (N418, N414, N346);
xor XOR2 (N419, N413, N315);
not NOT1 (N420, N400);
nand NAND4 (N421, N419, N365, N329, N134);
nand NAND4 (N422, N418, N34, N210, N373);
xor XOR2 (N423, N408, N269);
nand NAND3 (N424, N410, N192, N285);
nand NAND4 (N425, N422, N5, N10, N334);
nand NAND3 (N426, N424, N312, N333);
xor XOR2 (N427, N404, N118);
and AND2 (N428, N420, N386);
not NOT1 (N429, N407);
nor NOR2 (N430, N421, N275);
xor XOR2 (N431, N430, N58);
not NOT1 (N432, N429);
nor NOR4 (N433, N425, N80, N402, N277);
nor NOR3 (N434, N399, N231, N418);
not NOT1 (N435, N431);
or OR3 (N436, N433, N50, N272);
buf BUF1 (N437, N426);
buf BUF1 (N438, N437);
nand NAND3 (N439, N423, N82, N179);
or OR3 (N440, N439, N436, N216);
xor XOR2 (N441, N411, N46);
not NOT1 (N442, N441);
nor NOR4 (N443, N435, N90, N12, N249);
nand NAND4 (N444, N434, N291, N418, N303);
buf BUF1 (N445, N438);
and AND2 (N446, N445, N231);
not NOT1 (N447, N442);
nand NAND2 (N448, N432, N167);
or OR2 (N449, N447, N92);
xor XOR2 (N450, N446, N391);
buf BUF1 (N451, N443);
buf BUF1 (N452, N450);
or OR2 (N453, N448, N135);
nor NOR2 (N454, N451, N185);
xor XOR2 (N455, N452, N193);
nor NOR2 (N456, N455, N1);
and AND3 (N457, N454, N222, N210);
buf BUF1 (N458, N453);
nor NOR4 (N459, N417, N221, N359, N200);
or OR3 (N460, N456, N146, N437);
not NOT1 (N461, N416);
not NOT1 (N462, N449);
not NOT1 (N463, N459);
buf BUF1 (N464, N457);
not NOT1 (N465, N463);
xor XOR2 (N466, N427, N258);
nand NAND4 (N467, N444, N368, N327, N406);
nor NOR2 (N468, N464, N398);
and AND3 (N469, N461, N170, N140);
not NOT1 (N470, N465);
xor XOR2 (N471, N462, N44);
nor NOR3 (N472, N469, N60, N261);
or OR2 (N473, N428, N292);
nand NAND3 (N474, N466, N104, N26);
nand NAND3 (N475, N467, N61, N229);
and AND2 (N476, N474, N455);
and AND3 (N477, N458, N210, N253);
nor NOR3 (N478, N477, N109, N128);
nor NOR4 (N479, N460, N397, N66, N132);
nor NOR3 (N480, N468, N316, N366);
buf BUF1 (N481, N480);
xor XOR2 (N482, N440, N68);
not NOT1 (N483, N482);
nand NAND3 (N484, N478, N427, N30);
buf BUF1 (N485, N481);
nor NOR2 (N486, N476, N221);
or OR2 (N487, N471, N4);
and AND3 (N488, N483, N486, N178);
xor XOR2 (N489, N4, N111);
and AND2 (N490, N472, N111);
or OR4 (N491, N473, N172, N296, N273);
nand NAND4 (N492, N484, N397, N196, N332);
and AND3 (N493, N479, N45, N59);
xor XOR2 (N494, N485, N42);
nand NAND2 (N495, N490, N321);
and AND4 (N496, N470, N352, N70, N197);
or OR4 (N497, N493, N149, N163, N375);
xor XOR2 (N498, N495, N478);
xor XOR2 (N499, N489, N19);
buf BUF1 (N500, N492);
nor NOR2 (N501, N491, N121);
not NOT1 (N502, N496);
buf BUF1 (N503, N487);
nor NOR4 (N504, N488, N179, N372, N32);
or OR4 (N505, N497, N470, N419, N133);
and AND3 (N506, N494, N130, N131);
xor XOR2 (N507, N498, N326);
and AND4 (N508, N507, N496, N238, N363);
nand NAND2 (N509, N499, N375);
nor NOR2 (N510, N509, N72);
nor NOR2 (N511, N503, N66);
buf BUF1 (N512, N500);
nor NOR3 (N513, N510, N155, N412);
or OR3 (N514, N512, N7, N105);
buf BUF1 (N515, N475);
and AND2 (N516, N505, N107);
nand NAND2 (N517, N513, N71);
xor XOR2 (N518, N508, N409);
and AND4 (N519, N515, N132, N101, N79);
not NOT1 (N520, N517);
nand NAND4 (N521, N504, N423, N407, N391);
not NOT1 (N522, N511);
and AND3 (N523, N518, N339, N184);
buf BUF1 (N524, N520);
or OR4 (N525, N519, N109, N5, N300);
and AND2 (N526, N525, N7);
and AND2 (N527, N501, N359);
or OR3 (N528, N527, N52, N271);
or OR2 (N529, N516, N227);
xor XOR2 (N530, N522, N20);
and AND2 (N531, N530, N154);
buf BUF1 (N532, N524);
and AND2 (N533, N502, N50);
buf BUF1 (N534, N533);
buf BUF1 (N535, N532);
or OR3 (N536, N521, N202, N133);
buf BUF1 (N537, N536);
nor NOR4 (N538, N537, N36, N257, N188);
or OR3 (N539, N531, N38, N288);
xor XOR2 (N540, N534, N452);
or OR2 (N541, N529, N346);
or OR3 (N542, N538, N306, N63);
and AND2 (N543, N506, N254);
and AND2 (N544, N539, N539);
or OR3 (N545, N544, N161, N158);
nand NAND4 (N546, N543, N364, N545, N121);
nor NOR4 (N547, N312, N86, N439, N292);
nor NOR2 (N548, N523, N371);
and AND2 (N549, N541, N413);
nor NOR3 (N550, N535, N219, N107);
nor NOR4 (N551, N549, N131, N299, N308);
nor NOR2 (N552, N550, N257);
xor XOR2 (N553, N546, N532);
not NOT1 (N554, N547);
not NOT1 (N555, N526);
not NOT1 (N556, N551);
buf BUF1 (N557, N552);
nand NAND2 (N558, N556, N423);
xor XOR2 (N559, N548, N551);
nor NOR3 (N560, N558, N359, N2);
buf BUF1 (N561, N514);
or OR4 (N562, N553, N545, N43, N377);
nor NOR4 (N563, N528, N386, N556, N236);
and AND3 (N564, N554, N339, N254);
not NOT1 (N565, N540);
buf BUF1 (N566, N563);
and AND2 (N567, N557, N329);
buf BUF1 (N568, N564);
nor NOR3 (N569, N565, N390, N417);
nor NOR3 (N570, N568, N288, N432);
and AND3 (N571, N562, N217, N304);
nor NOR4 (N572, N559, N199, N453, N75);
or OR4 (N573, N555, N135, N277, N101);
buf BUF1 (N574, N573);
nand NAND3 (N575, N570, N491, N410);
buf BUF1 (N576, N566);
or OR2 (N577, N574, N412);
not NOT1 (N578, N576);
nand NAND2 (N579, N571, N465);
buf BUF1 (N580, N578);
xor XOR2 (N581, N542, N187);
nor NOR2 (N582, N560, N287);
nand NAND2 (N583, N579, N335);
nand NAND3 (N584, N582, N45, N207);
or OR2 (N585, N569, N100);
xor XOR2 (N586, N583, N146);
not NOT1 (N587, N577);
not NOT1 (N588, N584);
xor XOR2 (N589, N586, N403);
not NOT1 (N590, N589);
not NOT1 (N591, N587);
not NOT1 (N592, N580);
xor XOR2 (N593, N591, N308);
nor NOR3 (N594, N575, N94, N130);
and AND2 (N595, N594, N216);
buf BUF1 (N596, N592);
xor XOR2 (N597, N595, N259);
and AND4 (N598, N590, N37, N303, N153);
and AND4 (N599, N572, N45, N589, N277);
or OR4 (N600, N597, N458, N340, N467);
nand NAND2 (N601, N600, N449);
nor NOR2 (N602, N588, N273);
xor XOR2 (N603, N581, N579);
or OR2 (N604, N585, N390);
xor XOR2 (N605, N602, N431);
xor XOR2 (N606, N596, N491);
buf BUF1 (N607, N567);
buf BUF1 (N608, N604);
nor NOR2 (N609, N606, N449);
xor XOR2 (N610, N603, N327);
or OR2 (N611, N609, N250);
not NOT1 (N612, N607);
nand NAND4 (N613, N605, N409, N534, N134);
and AND3 (N614, N593, N267, N536);
and AND3 (N615, N561, N328, N140);
or OR4 (N616, N611, N357, N34, N585);
buf BUF1 (N617, N598);
nand NAND4 (N618, N617, N212, N273, N8);
nor NOR4 (N619, N599, N430, N296, N150);
nand NAND4 (N620, N613, N354, N105, N26);
xor XOR2 (N621, N608, N605);
buf BUF1 (N622, N601);
and AND4 (N623, N610, N544, N336, N270);
nand NAND3 (N624, N622, N80, N276);
not NOT1 (N625, N624);
not NOT1 (N626, N625);
nand NAND2 (N627, N615, N42);
not NOT1 (N628, N612);
buf BUF1 (N629, N620);
and AND3 (N630, N623, N396, N279);
xor XOR2 (N631, N626, N337);
not NOT1 (N632, N630);
buf BUF1 (N633, N619);
xor XOR2 (N634, N632, N541);
buf BUF1 (N635, N621);
nand NAND3 (N636, N633, N71, N462);
xor XOR2 (N637, N628, N241);
buf BUF1 (N638, N627);
or OR2 (N639, N636, N225);
nand NAND4 (N640, N616, N604, N95, N311);
nand NAND3 (N641, N618, N365, N134);
buf BUF1 (N642, N637);
nor NOR4 (N643, N614, N605, N223, N50);
buf BUF1 (N644, N638);
or OR4 (N645, N640, N145, N138, N549);
nor NOR3 (N646, N642, N577, N413);
or OR4 (N647, N634, N225, N499, N487);
xor XOR2 (N648, N639, N481);
and AND2 (N649, N635, N12);
nand NAND2 (N650, N646, N497);
xor XOR2 (N651, N631, N68);
and AND3 (N652, N648, N221, N577);
nor NOR3 (N653, N649, N25, N57);
xor XOR2 (N654, N651, N112);
nand NAND2 (N655, N650, N7);
nand NAND2 (N656, N652, N323);
not NOT1 (N657, N656);
and AND4 (N658, N647, N533, N331, N226);
and AND2 (N659, N629, N303);
and AND3 (N660, N654, N614, N431);
and AND3 (N661, N660, N494, N308);
nor NOR4 (N662, N643, N599, N339, N545);
buf BUF1 (N663, N645);
or OR3 (N664, N653, N376, N510);
nand NAND2 (N665, N663, N183);
or OR2 (N666, N661, N249);
nor NOR2 (N667, N657, N352);
nand NAND3 (N668, N664, N491, N325);
buf BUF1 (N669, N641);
nand NAND4 (N670, N655, N363, N372, N156);
nor NOR2 (N671, N668, N552);
nand NAND4 (N672, N669, N90, N135, N59);
or OR4 (N673, N666, N572, N531, N36);
or OR4 (N674, N662, N35, N636, N360);
nor NOR4 (N675, N670, N247, N28, N653);
nand NAND2 (N676, N665, N544);
xor XOR2 (N677, N644, N178);
or OR3 (N678, N677, N220, N469);
not NOT1 (N679, N674);
not NOT1 (N680, N672);
xor XOR2 (N681, N676, N436);
xor XOR2 (N682, N667, N491);
and AND4 (N683, N658, N256, N315, N216);
buf BUF1 (N684, N678);
and AND2 (N685, N681, N237);
not NOT1 (N686, N685);
or OR3 (N687, N659, N38, N273);
xor XOR2 (N688, N680, N395);
not NOT1 (N689, N673);
and AND2 (N690, N689, N535);
not NOT1 (N691, N675);
or OR2 (N692, N682, N335);
and AND2 (N693, N671, N58);
buf BUF1 (N694, N679);
and AND2 (N695, N683, N554);
nand NAND2 (N696, N694, N147);
not NOT1 (N697, N691);
and AND4 (N698, N690, N578, N168, N138);
and AND2 (N699, N684, N381);
nand NAND3 (N700, N698, N323, N477);
xor XOR2 (N701, N693, N168);
and AND3 (N702, N686, N146, N35);
nand NAND2 (N703, N699, N101);
not NOT1 (N704, N702);
and AND4 (N705, N701, N144, N265, N561);
nand NAND2 (N706, N687, N271);
or OR3 (N707, N696, N216, N556);
buf BUF1 (N708, N706);
not NOT1 (N709, N695);
not NOT1 (N710, N705);
or OR3 (N711, N704, N1, N516);
nand NAND2 (N712, N692, N128);
nand NAND3 (N713, N708, N563, N594);
nor NOR2 (N714, N709, N316);
nand NAND2 (N715, N697, N376);
nand NAND3 (N716, N710, N486, N253);
and AND2 (N717, N700, N148);
and AND4 (N718, N711, N709, N431, N449);
nand NAND3 (N719, N715, N395, N177);
buf BUF1 (N720, N703);
or OR3 (N721, N714, N299, N719);
nor NOR3 (N722, N628, N237, N335);
and AND2 (N723, N688, N517);
nand NAND3 (N724, N713, N176, N571);
nor NOR3 (N725, N716, N672, N130);
or OR2 (N726, N721, N367);
nor NOR2 (N727, N712, N35);
xor XOR2 (N728, N724, N480);
and AND2 (N729, N722, N27);
buf BUF1 (N730, N723);
not NOT1 (N731, N729);
xor XOR2 (N732, N730, N177);
nor NOR3 (N733, N728, N148, N715);
buf BUF1 (N734, N726);
or OR3 (N735, N734, N522, N534);
buf BUF1 (N736, N735);
xor XOR2 (N737, N720, N505);
or OR3 (N738, N725, N316, N355);
nand NAND3 (N739, N717, N173, N195);
buf BUF1 (N740, N739);
or OR2 (N741, N736, N255);
xor XOR2 (N742, N727, N162);
not NOT1 (N743, N733);
xor XOR2 (N744, N741, N238);
not NOT1 (N745, N742);
not NOT1 (N746, N718);
buf BUF1 (N747, N707);
nand NAND4 (N748, N732, N210, N227, N356);
nor NOR2 (N749, N737, N647);
nand NAND4 (N750, N746, N547, N426, N156);
not NOT1 (N751, N731);
nand NAND2 (N752, N740, N523);
and AND4 (N753, N743, N68, N106, N447);
xor XOR2 (N754, N752, N378);
nand NAND3 (N755, N749, N654, N432);
buf BUF1 (N756, N755);
nor NOR4 (N757, N750, N45, N718, N402);
buf BUF1 (N758, N745);
nor NOR4 (N759, N744, N572, N55, N362);
not NOT1 (N760, N754);
or OR3 (N761, N759, N396, N609);
buf BUF1 (N762, N758);
and AND4 (N763, N748, N571, N496, N455);
xor XOR2 (N764, N753, N359);
nand NAND3 (N765, N760, N100, N230);
nand NAND4 (N766, N762, N420, N338, N529);
nand NAND2 (N767, N756, N678);
or OR3 (N768, N751, N91, N690);
and AND3 (N769, N765, N415, N292);
xor XOR2 (N770, N761, N11);
nor NOR2 (N771, N738, N581);
or OR4 (N772, N769, N249, N582, N396);
xor XOR2 (N773, N771, N334);
not NOT1 (N774, N757);
buf BUF1 (N775, N773);
xor XOR2 (N776, N767, N398);
xor XOR2 (N777, N774, N368);
and AND4 (N778, N747, N694, N194, N726);
or OR2 (N779, N775, N435);
nand NAND4 (N780, N776, N690, N267, N180);
nor NOR4 (N781, N768, N557, N342, N420);
buf BUF1 (N782, N770);
buf BUF1 (N783, N764);
and AND3 (N784, N777, N184, N49);
and AND2 (N785, N782, N715);
buf BUF1 (N786, N766);
not NOT1 (N787, N781);
nand NAND4 (N788, N783, N587, N348, N414);
buf BUF1 (N789, N778);
not NOT1 (N790, N785);
nand NAND2 (N791, N786, N736);
and AND4 (N792, N772, N78, N322, N321);
nand NAND2 (N793, N784, N412);
or OR2 (N794, N787, N652);
nor NOR4 (N795, N789, N515, N60, N394);
xor XOR2 (N796, N794, N62);
not NOT1 (N797, N790);
or OR3 (N798, N797, N214, N377);
nand NAND4 (N799, N763, N527, N272, N122);
or OR3 (N800, N779, N366, N762);
nor NOR4 (N801, N798, N589, N44, N239);
or OR4 (N802, N795, N420, N284, N151);
xor XOR2 (N803, N788, N319);
xor XOR2 (N804, N801, N246);
not NOT1 (N805, N800);
and AND2 (N806, N780, N375);
nor NOR2 (N807, N806, N728);
and AND2 (N808, N802, N751);
or OR2 (N809, N805, N423);
and AND2 (N810, N796, N157);
nand NAND2 (N811, N792, N289);
or OR3 (N812, N791, N216, N564);
nand NAND2 (N813, N810, N812);
xor XOR2 (N814, N169, N221);
nand NAND2 (N815, N814, N314);
buf BUF1 (N816, N811);
buf BUF1 (N817, N807);
or OR4 (N818, N809, N768, N563, N127);
or OR4 (N819, N804, N527, N534, N386);
or OR3 (N820, N818, N409, N651);
buf BUF1 (N821, N813);
xor XOR2 (N822, N817, N408);
not NOT1 (N823, N799);
xor XOR2 (N824, N815, N307);
and AND3 (N825, N803, N738, N511);
or OR2 (N826, N816, N683);
nor NOR3 (N827, N826, N239, N461);
or OR2 (N828, N823, N816);
or OR2 (N829, N793, N733);
buf BUF1 (N830, N828);
and AND4 (N831, N829, N157, N748, N530);
nor NOR2 (N832, N830, N627);
not NOT1 (N833, N832);
nand NAND2 (N834, N822, N706);
buf BUF1 (N835, N808);
nand NAND4 (N836, N825, N662, N412, N87);
nor NOR2 (N837, N833, N49);
xor XOR2 (N838, N836, N130);
not NOT1 (N839, N819);
not NOT1 (N840, N824);
buf BUF1 (N841, N834);
nand NAND4 (N842, N821, N150, N186, N47);
xor XOR2 (N843, N842, N779);
buf BUF1 (N844, N843);
and AND2 (N845, N831, N747);
nand NAND3 (N846, N839, N631, N126);
nor NOR2 (N847, N838, N6);
nor NOR3 (N848, N845, N683, N367);
and AND2 (N849, N844, N415);
xor XOR2 (N850, N841, N324);
not NOT1 (N851, N837);
or OR4 (N852, N847, N96, N394, N481);
or OR3 (N853, N848, N831, N834);
buf BUF1 (N854, N853);
buf BUF1 (N855, N852);
nor NOR2 (N856, N827, N300);
xor XOR2 (N857, N850, N45);
and AND3 (N858, N849, N572, N695);
not NOT1 (N859, N851);
nand NAND4 (N860, N859, N574, N460, N437);
nor NOR3 (N861, N857, N748, N777);
and AND2 (N862, N840, N217);
xor XOR2 (N863, N820, N81);
buf BUF1 (N864, N854);
nor NOR3 (N865, N860, N280, N306);
not NOT1 (N866, N864);
and AND3 (N867, N855, N60, N756);
and AND3 (N868, N835, N202, N228);
or OR2 (N869, N856, N71);
nand NAND4 (N870, N863, N86, N215, N123);
buf BUF1 (N871, N866);
nand NAND2 (N872, N868, N600);
xor XOR2 (N873, N869, N455);
and AND3 (N874, N846, N433, N665);
and AND3 (N875, N861, N401, N628);
buf BUF1 (N876, N870);
or OR4 (N877, N858, N146, N195, N158);
nor NOR2 (N878, N874, N615);
not NOT1 (N879, N876);
nor NOR4 (N880, N865, N309, N706, N571);
xor XOR2 (N881, N867, N578);
and AND4 (N882, N875, N467, N451, N459);
or OR2 (N883, N872, N649);
nor NOR2 (N884, N879, N150);
and AND4 (N885, N871, N315, N512, N740);
and AND4 (N886, N873, N847, N776, N607);
buf BUF1 (N887, N880);
and AND2 (N888, N877, N160);
or OR4 (N889, N884, N301, N723, N421);
nor NOR2 (N890, N889, N285);
or OR2 (N891, N878, N707);
nor NOR4 (N892, N885, N555, N624, N446);
buf BUF1 (N893, N890);
buf BUF1 (N894, N893);
nor NOR4 (N895, N883, N119, N182, N626);
and AND3 (N896, N888, N501, N130);
nand NAND3 (N897, N891, N28, N275);
nor NOR3 (N898, N882, N415, N812);
nand NAND3 (N899, N895, N830, N164);
nor NOR4 (N900, N898, N738, N699, N166);
or OR2 (N901, N896, N594);
or OR2 (N902, N900, N808);
not NOT1 (N903, N892);
buf BUF1 (N904, N881);
and AND3 (N905, N887, N836, N424);
nor NOR4 (N906, N862, N348, N184, N64);
nand NAND3 (N907, N886, N803, N508);
and AND4 (N908, N905, N529, N416, N214);
or OR2 (N909, N907, N276);
and AND2 (N910, N901, N738);
nor NOR2 (N911, N910, N187);
nand NAND4 (N912, N903, N361, N770, N487);
nor NOR2 (N913, N912, N902);
or OR3 (N914, N522, N189, N127);
buf BUF1 (N915, N914);
nor NOR4 (N916, N894, N346, N657, N908);
buf BUF1 (N917, N136);
xor XOR2 (N918, N906, N237);
buf BUF1 (N919, N916);
and AND2 (N920, N899, N444);
nor NOR2 (N921, N909, N99);
and AND4 (N922, N897, N342, N474, N547);
nand NAND4 (N923, N913, N673, N22, N883);
or OR3 (N924, N904, N326, N525);
or OR3 (N925, N911, N677, N658);
not NOT1 (N926, N917);
or OR2 (N927, N918, N419);
and AND2 (N928, N925, N857);
buf BUF1 (N929, N920);
and AND4 (N930, N915, N288, N333, N230);
or OR2 (N931, N926, N278);
or OR2 (N932, N921, N249);
or OR2 (N933, N930, N163);
and AND3 (N934, N928, N912, N538);
or OR3 (N935, N927, N189, N849);
nand NAND4 (N936, N924, N409, N592, N463);
nand NAND4 (N937, N929, N102, N775, N517);
nor NOR2 (N938, N935, N49);
not NOT1 (N939, N934);
xor XOR2 (N940, N932, N35);
nor NOR3 (N941, N931, N570, N790);
not NOT1 (N942, N938);
or OR4 (N943, N940, N678, N784, N237);
buf BUF1 (N944, N919);
buf BUF1 (N945, N941);
nor NOR2 (N946, N945, N70);
xor XOR2 (N947, N936, N946);
nand NAND2 (N948, N665, N843);
buf BUF1 (N949, N943);
not NOT1 (N950, N933);
not NOT1 (N951, N937);
or OR4 (N952, N948, N655, N98, N907);
nand NAND2 (N953, N949, N424);
nor NOR3 (N954, N942, N286, N41);
buf BUF1 (N955, N939);
and AND3 (N956, N923, N163, N190);
xor XOR2 (N957, N950, N920);
or OR2 (N958, N947, N333);
or OR2 (N959, N922, N924);
buf BUF1 (N960, N957);
buf BUF1 (N961, N954);
not NOT1 (N962, N961);
nand NAND2 (N963, N959, N160);
nand NAND2 (N964, N958, N575);
buf BUF1 (N965, N963);
not NOT1 (N966, N964);
buf BUF1 (N967, N951);
buf BUF1 (N968, N956);
not NOT1 (N969, N965);
and AND3 (N970, N968, N518, N519);
nand NAND2 (N971, N960, N205);
or OR3 (N972, N962, N921, N706);
nand NAND4 (N973, N972, N513, N722, N831);
nand NAND4 (N974, N967, N702, N747, N776);
nand NAND4 (N975, N953, N263, N757, N447);
nand NAND4 (N976, N975, N269, N955, N298);
xor XOR2 (N977, N622, N848);
nor NOR4 (N978, N973, N150, N697, N471);
nand NAND4 (N979, N944, N654, N475, N673);
nor NOR4 (N980, N979, N897, N911, N586);
buf BUF1 (N981, N952);
and AND2 (N982, N977, N397);
xor XOR2 (N983, N974, N207);
nor NOR2 (N984, N980, N551);
and AND4 (N985, N984, N2, N455, N267);
not NOT1 (N986, N969);
and AND2 (N987, N981, N501);
nor NOR2 (N988, N976, N212);
nand NAND4 (N989, N966, N487, N266, N846);
buf BUF1 (N990, N985);
xor XOR2 (N991, N970, N130);
nor NOR4 (N992, N989, N148, N212, N65);
not NOT1 (N993, N971);
and AND3 (N994, N978, N264, N387);
and AND4 (N995, N987, N805, N992, N494);
not NOT1 (N996, N55);
nor NOR3 (N997, N990, N324, N595);
or OR3 (N998, N994, N117, N320);
nor NOR3 (N999, N998, N67, N991);
nand NAND4 (N1000, N408, N735, N41, N101);
buf BUF1 (N1001, N993);
and AND3 (N1002, N1001, N296, N336);
nor NOR4 (N1003, N1002, N60, N198, N312);
xor XOR2 (N1004, N1000, N199);
not NOT1 (N1005, N1003);
not NOT1 (N1006, N988);
nor NOR3 (N1007, N982, N361, N498);
nand NAND3 (N1008, N999, N361, N864);
or OR2 (N1009, N995, N196);
xor XOR2 (N1010, N1007, N603);
not NOT1 (N1011, N1008);
nor NOR2 (N1012, N1010, N817);
or OR4 (N1013, N986, N55, N849, N744);
or OR2 (N1014, N1005, N694);
nor NOR3 (N1015, N1012, N811, N551);
or OR4 (N1016, N997, N283, N741, N141);
nand NAND4 (N1017, N1009, N858, N512, N385);
not NOT1 (N1018, N1015);
nor NOR2 (N1019, N1006, N392);
not NOT1 (N1020, N1014);
xor XOR2 (N1021, N1011, N389);
xor XOR2 (N1022, N983, N735);
xor XOR2 (N1023, N1017, N267);
nor NOR3 (N1024, N1023, N595, N594);
nand NAND2 (N1025, N1018, N832);
buf BUF1 (N1026, N1025);
nor NOR4 (N1027, N1026, N643, N301, N328);
nand NAND3 (N1028, N1021, N812, N132);
xor XOR2 (N1029, N1020, N863);
nor NOR4 (N1030, N1022, N520, N771, N777);
and AND2 (N1031, N1030, N532);
and AND2 (N1032, N996, N696);
and AND2 (N1033, N1019, N158);
not NOT1 (N1034, N1028);
or OR4 (N1035, N1029, N3, N80, N585);
or OR3 (N1036, N1033, N432, N85);
xor XOR2 (N1037, N1024, N59);
or OR3 (N1038, N1031, N595, N610);
not NOT1 (N1039, N1038);
not NOT1 (N1040, N1013);
xor XOR2 (N1041, N1040, N970);
not NOT1 (N1042, N1034);
and AND2 (N1043, N1042, N334);
nor NOR2 (N1044, N1004, N120);
and AND3 (N1045, N1016, N891, N574);
xor XOR2 (N1046, N1039, N469);
xor XOR2 (N1047, N1044, N718);
nor NOR2 (N1048, N1027, N907);
buf BUF1 (N1049, N1047);
not NOT1 (N1050, N1045);
buf BUF1 (N1051, N1048);
or OR3 (N1052, N1050, N714, N909);
nand NAND4 (N1053, N1032, N248, N635, N170);
nor NOR2 (N1054, N1043, N644);
or OR3 (N1055, N1046, N465, N856);
nor NOR4 (N1056, N1054, N574, N547, N452);
nor NOR4 (N1057, N1055, N556, N721, N270);
xor XOR2 (N1058, N1035, N754);
not NOT1 (N1059, N1051);
nor NOR4 (N1060, N1057, N506, N220, N878);
not NOT1 (N1061, N1053);
or OR2 (N1062, N1036, N875);
xor XOR2 (N1063, N1056, N21);
xor XOR2 (N1064, N1060, N683);
xor XOR2 (N1065, N1058, N267);
buf BUF1 (N1066, N1037);
nand NAND3 (N1067, N1065, N690, N393);
and AND4 (N1068, N1067, N245, N73, N485);
or OR4 (N1069, N1052, N631, N1062, N743);
not NOT1 (N1070, N630);
nor NOR2 (N1071, N1070, N398);
and AND4 (N1072, N1049, N876, N44, N389);
buf BUF1 (N1073, N1064);
not NOT1 (N1074, N1041);
or OR3 (N1075, N1073, N628, N1057);
nor NOR3 (N1076, N1075, N287, N281);
xor XOR2 (N1077, N1071, N1021);
xor XOR2 (N1078, N1068, N348);
or OR4 (N1079, N1072, N818, N421, N145);
and AND2 (N1080, N1074, N45);
xor XOR2 (N1081, N1069, N185);
xor XOR2 (N1082, N1078, N583);
nand NAND2 (N1083, N1082, N15);
or OR3 (N1084, N1063, N29, N646);
xor XOR2 (N1085, N1077, N364);
and AND2 (N1086, N1066, N604);
nor NOR2 (N1087, N1059, N411);
nor NOR2 (N1088, N1079, N954);
nor NOR4 (N1089, N1083, N867, N927, N1022);
or OR3 (N1090, N1084, N829, N764);
and AND3 (N1091, N1061, N672, N473);
and AND4 (N1092, N1090, N209, N567, N148);
or OR4 (N1093, N1081, N925, N142, N310);
or OR2 (N1094, N1088, N85);
nor NOR3 (N1095, N1080, N911, N336);
not NOT1 (N1096, N1086);
not NOT1 (N1097, N1087);
xor XOR2 (N1098, N1076, N125);
nor NOR3 (N1099, N1085, N294, N403);
nor NOR3 (N1100, N1098, N116, N178);
nor NOR3 (N1101, N1089, N316, N1060);
nand NAND2 (N1102, N1097, N105);
and AND4 (N1103, N1099, N250, N917, N605);
nor NOR3 (N1104, N1092, N1021, N43);
nand NAND4 (N1105, N1096, N874, N147, N447);
xor XOR2 (N1106, N1091, N155);
nand NAND2 (N1107, N1104, N905);
xor XOR2 (N1108, N1100, N12);
nor NOR2 (N1109, N1095, N631);
nor NOR4 (N1110, N1101, N550, N847, N277);
buf BUF1 (N1111, N1109);
xor XOR2 (N1112, N1102, N1018);
buf BUF1 (N1113, N1094);
not NOT1 (N1114, N1111);
nor NOR2 (N1115, N1112, N224);
not NOT1 (N1116, N1108);
or OR2 (N1117, N1113, N1053);
not NOT1 (N1118, N1116);
or OR4 (N1119, N1103, N1118, N742, N219);
nor NOR2 (N1120, N51, N194);
nor NOR4 (N1121, N1120, N501, N310, N378);
nand NAND3 (N1122, N1117, N607, N974);
nor NOR3 (N1123, N1106, N324, N302);
or OR2 (N1124, N1093, N863);
and AND2 (N1125, N1123, N276);
or OR3 (N1126, N1105, N561, N1039);
nor NOR2 (N1127, N1121, N954);
xor XOR2 (N1128, N1122, N92);
or OR4 (N1129, N1107, N1045, N281, N481);
buf BUF1 (N1130, N1129);
and AND3 (N1131, N1115, N538, N466);
xor XOR2 (N1132, N1114, N479);
buf BUF1 (N1133, N1130);
or OR4 (N1134, N1132, N939, N701, N1092);
nand NAND3 (N1135, N1127, N199, N381);
and AND3 (N1136, N1133, N46, N275);
or OR3 (N1137, N1124, N916, N976);
nor NOR2 (N1138, N1110, N708);
buf BUF1 (N1139, N1136);
buf BUF1 (N1140, N1128);
nand NAND4 (N1141, N1137, N1120, N202, N720);
not NOT1 (N1142, N1138);
buf BUF1 (N1143, N1135);
and AND4 (N1144, N1134, N880, N155, N513);
and AND2 (N1145, N1125, N35);
buf BUF1 (N1146, N1145);
or OR4 (N1147, N1144, N1125, N1109, N833);
not NOT1 (N1148, N1142);
and AND2 (N1149, N1147, N627);
nand NAND3 (N1150, N1143, N208, N1032);
nand NAND4 (N1151, N1131, N571, N996, N89);
xor XOR2 (N1152, N1149, N320);
xor XOR2 (N1153, N1139, N940);
and AND2 (N1154, N1151, N282);
or OR2 (N1155, N1154, N273);
and AND3 (N1156, N1148, N324, N392);
xor XOR2 (N1157, N1141, N782);
nor NOR4 (N1158, N1153, N163, N1144, N863);
not NOT1 (N1159, N1155);
xor XOR2 (N1160, N1126, N457);
buf BUF1 (N1161, N1152);
or OR3 (N1162, N1150, N430, N465);
or OR4 (N1163, N1159, N1117, N116, N380);
nor NOR3 (N1164, N1119, N382, N276);
nand NAND3 (N1165, N1161, N536, N276);
and AND2 (N1166, N1164, N445);
nand NAND3 (N1167, N1157, N1027, N1127);
buf BUF1 (N1168, N1163);
or OR4 (N1169, N1156, N1148, N1143, N812);
not NOT1 (N1170, N1158);
not NOT1 (N1171, N1169);
nand NAND2 (N1172, N1171, N439);
or OR3 (N1173, N1167, N604, N876);
not NOT1 (N1174, N1170);
nor NOR2 (N1175, N1174, N1159);
nor NOR2 (N1176, N1173, N722);
buf BUF1 (N1177, N1140);
nand NAND2 (N1178, N1160, N697);
and AND3 (N1179, N1146, N958, N44);
or OR4 (N1180, N1178, N4, N356, N1081);
or OR4 (N1181, N1172, N8, N14, N333);
or OR2 (N1182, N1180, N331);
and AND3 (N1183, N1165, N834, N946);
xor XOR2 (N1184, N1168, N1132);
xor XOR2 (N1185, N1184, N2);
or OR2 (N1186, N1166, N495);
not NOT1 (N1187, N1186);
nor NOR3 (N1188, N1183, N278, N406);
nor NOR4 (N1189, N1179, N798, N405, N35);
not NOT1 (N1190, N1187);
and AND3 (N1191, N1189, N95, N299);
nand NAND2 (N1192, N1188, N522);
xor XOR2 (N1193, N1192, N860);
nor NOR3 (N1194, N1182, N211, N996);
xor XOR2 (N1195, N1162, N712);
buf BUF1 (N1196, N1193);
xor XOR2 (N1197, N1177, N662);
not NOT1 (N1198, N1181);
xor XOR2 (N1199, N1198, N612);
not NOT1 (N1200, N1197);
not NOT1 (N1201, N1199);
nand NAND3 (N1202, N1176, N215, N182);
not NOT1 (N1203, N1175);
and AND2 (N1204, N1201, N357);
nor NOR4 (N1205, N1204, N368, N409, N303);
or OR2 (N1206, N1191, N1162);
nor NOR4 (N1207, N1190, N551, N653, N844);
and AND2 (N1208, N1207, N679);
or OR2 (N1209, N1205, N311);
not NOT1 (N1210, N1206);
not NOT1 (N1211, N1210);
nor NOR3 (N1212, N1202, N246, N466);
nor NOR4 (N1213, N1196, N1210, N25, N1034);
not NOT1 (N1214, N1212);
buf BUF1 (N1215, N1185);
nor NOR4 (N1216, N1194, N994, N1214, N1159);
not NOT1 (N1217, N574);
nand NAND4 (N1218, N1209, N793, N1072, N652);
or OR4 (N1219, N1195, N297, N309, N634);
and AND3 (N1220, N1211, N117, N1063);
xor XOR2 (N1221, N1218, N925);
or OR3 (N1222, N1217, N1100, N732);
not NOT1 (N1223, N1208);
and AND4 (N1224, N1215, N761, N1012, N663);
nand NAND3 (N1225, N1200, N100, N806);
buf BUF1 (N1226, N1222);
and AND2 (N1227, N1226, N1156);
xor XOR2 (N1228, N1225, N922);
xor XOR2 (N1229, N1203, N364);
nand NAND3 (N1230, N1213, N863, N1148);
not NOT1 (N1231, N1223);
buf BUF1 (N1232, N1219);
or OR2 (N1233, N1221, N653);
and AND3 (N1234, N1227, N1146, N259);
nand NAND4 (N1235, N1234, N615, N30, N408);
xor XOR2 (N1236, N1231, N352);
and AND4 (N1237, N1220, N308, N648, N827);
and AND3 (N1238, N1237, N177, N568);
nor NOR2 (N1239, N1232, N350);
nor NOR3 (N1240, N1228, N656, N157);
and AND2 (N1241, N1233, N125);
xor XOR2 (N1242, N1230, N1044);
buf BUF1 (N1243, N1238);
not NOT1 (N1244, N1243);
nand NAND4 (N1245, N1240, N922, N817, N918);
not NOT1 (N1246, N1245);
xor XOR2 (N1247, N1242, N101);
and AND3 (N1248, N1216, N1161, N744);
not NOT1 (N1249, N1229);
nor NOR4 (N1250, N1247, N999, N695, N519);
xor XOR2 (N1251, N1246, N479);
or OR3 (N1252, N1235, N1063, N1247);
and AND4 (N1253, N1249, N89, N105, N840);
xor XOR2 (N1254, N1248, N87);
buf BUF1 (N1255, N1252);
not NOT1 (N1256, N1251);
buf BUF1 (N1257, N1256);
nand NAND3 (N1258, N1244, N527, N701);
not NOT1 (N1259, N1257);
nand NAND2 (N1260, N1254, N175);
and AND3 (N1261, N1250, N460, N967);
nand NAND3 (N1262, N1253, N588, N111);
nand NAND3 (N1263, N1236, N1132, N142);
xor XOR2 (N1264, N1263, N461);
not NOT1 (N1265, N1264);
or OR3 (N1266, N1241, N427, N769);
xor XOR2 (N1267, N1266, N843);
xor XOR2 (N1268, N1239, N233);
or OR4 (N1269, N1267, N929, N1165, N315);
not NOT1 (N1270, N1262);
and AND4 (N1271, N1265, N1042, N928, N1093);
nand NAND3 (N1272, N1260, N142, N206);
and AND3 (N1273, N1261, N518, N1113);
nor NOR4 (N1274, N1273, N28, N1208, N1230);
nor NOR2 (N1275, N1269, N236);
and AND2 (N1276, N1270, N1005);
buf BUF1 (N1277, N1272);
nand NAND2 (N1278, N1277, N345);
nor NOR3 (N1279, N1224, N408, N675);
buf BUF1 (N1280, N1274);
buf BUF1 (N1281, N1278);
buf BUF1 (N1282, N1281);
buf BUF1 (N1283, N1258);
nor NOR4 (N1284, N1276, N339, N920, N536);
buf BUF1 (N1285, N1279);
not NOT1 (N1286, N1271);
nand NAND3 (N1287, N1255, N727, N737);
or OR4 (N1288, N1283, N115, N27, N1047);
and AND4 (N1289, N1259, N1231, N289, N1237);
xor XOR2 (N1290, N1275, N616);
or OR4 (N1291, N1289, N852, N209, N666);
and AND2 (N1292, N1290, N148);
or OR3 (N1293, N1285, N1025, N936);
buf BUF1 (N1294, N1268);
and AND3 (N1295, N1282, N440, N546);
or OR3 (N1296, N1291, N1133, N41);
or OR3 (N1297, N1292, N1287, N549);
nor NOR2 (N1298, N471, N208);
buf BUF1 (N1299, N1298);
nor NOR2 (N1300, N1296, N615);
and AND2 (N1301, N1299, N341);
and AND4 (N1302, N1294, N963, N395, N1048);
not NOT1 (N1303, N1301);
and AND4 (N1304, N1302, N97, N943, N1224);
not NOT1 (N1305, N1295);
not NOT1 (N1306, N1293);
buf BUF1 (N1307, N1304);
xor XOR2 (N1308, N1306, N336);
and AND4 (N1309, N1288, N1130, N842, N477);
not NOT1 (N1310, N1280);
xor XOR2 (N1311, N1303, N71);
xor XOR2 (N1312, N1308, N215);
and AND4 (N1313, N1305, N468, N977, N743);
buf BUF1 (N1314, N1311);
not NOT1 (N1315, N1284);
nor NOR3 (N1316, N1310, N924, N736);
xor XOR2 (N1317, N1286, N814);
xor XOR2 (N1318, N1317, N1172);
xor XOR2 (N1319, N1300, N88);
not NOT1 (N1320, N1313);
xor XOR2 (N1321, N1309, N371);
xor XOR2 (N1322, N1315, N933);
or OR3 (N1323, N1322, N218, N674);
and AND2 (N1324, N1321, N1069);
nor NOR3 (N1325, N1324, N1238, N960);
or OR3 (N1326, N1312, N1068, N1002);
buf BUF1 (N1327, N1297);
xor XOR2 (N1328, N1325, N738);
nor NOR2 (N1329, N1314, N697);
nor NOR4 (N1330, N1328, N714, N52, N290);
nor NOR3 (N1331, N1330, N917, N650);
or OR3 (N1332, N1329, N1152, N756);
not NOT1 (N1333, N1323);
buf BUF1 (N1334, N1326);
nand NAND2 (N1335, N1316, N83);
xor XOR2 (N1336, N1327, N952);
nand NAND3 (N1337, N1332, N483, N93);
buf BUF1 (N1338, N1335);
buf BUF1 (N1339, N1336);
nand NAND4 (N1340, N1318, N960, N854, N104);
nand NAND2 (N1341, N1307, N566);
nor NOR4 (N1342, N1337, N305, N1027, N890);
or OR3 (N1343, N1338, N883, N64);
not NOT1 (N1344, N1320);
buf BUF1 (N1345, N1341);
xor XOR2 (N1346, N1319, N255);
not NOT1 (N1347, N1340);
nor NOR3 (N1348, N1345, N82, N1249);
xor XOR2 (N1349, N1339, N604);
not NOT1 (N1350, N1349);
or OR2 (N1351, N1334, N536);
xor XOR2 (N1352, N1346, N390);
xor XOR2 (N1353, N1342, N65);
not NOT1 (N1354, N1343);
nor NOR4 (N1355, N1333, N588, N1124, N1015);
xor XOR2 (N1356, N1331, N576);
and AND2 (N1357, N1353, N670);
nand NAND4 (N1358, N1348, N766, N295, N768);
nor NOR3 (N1359, N1352, N1127, N1345);
nand NAND3 (N1360, N1356, N1050, N50);
not NOT1 (N1361, N1360);
not NOT1 (N1362, N1357);
or OR2 (N1363, N1361, N1351);
or OR3 (N1364, N1030, N425, N1018);
or OR3 (N1365, N1358, N688, N499);
nor NOR2 (N1366, N1365, N677);
xor XOR2 (N1367, N1347, N767);
buf BUF1 (N1368, N1359);
and AND3 (N1369, N1368, N944, N821);
or OR4 (N1370, N1363, N866, N51, N1073);
nand NAND2 (N1371, N1369, N446);
buf BUF1 (N1372, N1350);
and AND4 (N1373, N1371, N1234, N1049, N794);
and AND3 (N1374, N1355, N936, N552);
nor NOR2 (N1375, N1374, N53);
and AND2 (N1376, N1362, N813);
buf BUF1 (N1377, N1370);
not NOT1 (N1378, N1377);
nor NOR3 (N1379, N1375, N349, N284);
and AND4 (N1380, N1367, N867, N760, N606);
not NOT1 (N1381, N1366);
buf BUF1 (N1382, N1344);
and AND4 (N1383, N1376, N1302, N870, N185);
and AND3 (N1384, N1372, N1161, N538);
nor NOR3 (N1385, N1379, N108, N700);
or OR3 (N1386, N1384, N1210, N1036);
xor XOR2 (N1387, N1373, N648);
and AND4 (N1388, N1381, N1350, N884, N203);
not NOT1 (N1389, N1388);
and AND2 (N1390, N1383, N821);
xor XOR2 (N1391, N1382, N17);
and AND2 (N1392, N1354, N79);
or OR3 (N1393, N1380, N428, N481);
buf BUF1 (N1394, N1378);
or OR3 (N1395, N1385, N523, N89);
nor NOR3 (N1396, N1394, N1185, N738);
or OR4 (N1397, N1391, N1079, N421, N104);
nand NAND3 (N1398, N1397, N1208, N802);
nor NOR3 (N1399, N1393, N101, N1241);
not NOT1 (N1400, N1387);
or OR2 (N1401, N1400, N1259);
nand NAND4 (N1402, N1389, N278, N213, N75);
not NOT1 (N1403, N1395);
and AND4 (N1404, N1402, N107, N641, N478);
xor XOR2 (N1405, N1403, N860);
xor XOR2 (N1406, N1364, N878);
not NOT1 (N1407, N1386);
buf BUF1 (N1408, N1405);
xor XOR2 (N1409, N1406, N121);
buf BUF1 (N1410, N1401);
buf BUF1 (N1411, N1396);
and AND2 (N1412, N1399, N1362);
buf BUF1 (N1413, N1412);
nand NAND4 (N1414, N1411, N640, N299, N697);
and AND3 (N1415, N1398, N244, N573);
or OR2 (N1416, N1415, N1362);
nand NAND4 (N1417, N1408, N1145, N1283, N202);
nand NAND2 (N1418, N1390, N1070);
or OR3 (N1419, N1410, N1201, N1057);
xor XOR2 (N1420, N1392, N1132);
nand NAND4 (N1421, N1407, N229, N1049, N111);
and AND3 (N1422, N1409, N450, N321);
nand NAND3 (N1423, N1419, N523, N1161);
nor NOR2 (N1424, N1413, N1240);
nand NAND2 (N1425, N1423, N839);
buf BUF1 (N1426, N1421);
and AND3 (N1427, N1420, N358, N1214);
or OR3 (N1428, N1416, N747, N560);
xor XOR2 (N1429, N1414, N405);
nor NOR4 (N1430, N1428, N795, N908, N1093);
nand NAND2 (N1431, N1418, N33);
and AND4 (N1432, N1427, N868, N128, N805);
nor NOR4 (N1433, N1425, N965, N575, N107);
buf BUF1 (N1434, N1430);
buf BUF1 (N1435, N1404);
nor NOR3 (N1436, N1429, N12, N273);
xor XOR2 (N1437, N1434, N146);
nor NOR3 (N1438, N1422, N227, N234);
and AND4 (N1439, N1417, N202, N1157, N1373);
nor NOR3 (N1440, N1426, N198, N313);
xor XOR2 (N1441, N1437, N1417);
or OR3 (N1442, N1424, N193, N1215);
nand NAND3 (N1443, N1440, N1394, N875);
not NOT1 (N1444, N1439);
and AND4 (N1445, N1444, N1225, N1121, N1078);
nor NOR2 (N1446, N1441, N1205);
xor XOR2 (N1447, N1436, N332);
or OR2 (N1448, N1443, N547);
or OR4 (N1449, N1432, N211, N927, N1330);
or OR3 (N1450, N1438, N785, N1189);
not NOT1 (N1451, N1447);
and AND2 (N1452, N1446, N1380);
buf BUF1 (N1453, N1448);
nor NOR2 (N1454, N1449, N766);
and AND2 (N1455, N1451, N1005);
not NOT1 (N1456, N1450);
buf BUF1 (N1457, N1453);
buf BUF1 (N1458, N1457);
buf BUF1 (N1459, N1452);
nor NOR3 (N1460, N1445, N557, N402);
not NOT1 (N1461, N1459);
nand NAND4 (N1462, N1435, N623, N719, N855);
not NOT1 (N1463, N1433);
xor XOR2 (N1464, N1463, N805);
and AND2 (N1465, N1442, N1239);
or OR2 (N1466, N1455, N915);
and AND2 (N1467, N1462, N1153);
or OR4 (N1468, N1461, N879, N1386, N764);
and AND3 (N1469, N1465, N118, N605);
buf BUF1 (N1470, N1454);
nand NAND2 (N1471, N1456, N467);
xor XOR2 (N1472, N1467, N85);
buf BUF1 (N1473, N1464);
nor NOR4 (N1474, N1431, N885, N16, N927);
nor NOR2 (N1475, N1473, N1065);
and AND3 (N1476, N1468, N142, N820);
nand NAND4 (N1477, N1460, N858, N465, N132);
nor NOR3 (N1478, N1477, N1457, N75);
and AND4 (N1479, N1469, N420, N198, N62);
nand NAND4 (N1480, N1458, N1466, N262, N505);
not NOT1 (N1481, N441);
nand NAND2 (N1482, N1471, N115);
xor XOR2 (N1483, N1482, N670);
buf BUF1 (N1484, N1475);
nand NAND4 (N1485, N1479, N628, N945, N1413);
or OR4 (N1486, N1474, N1096, N287, N1328);
nor NOR3 (N1487, N1480, N1368, N168);
not NOT1 (N1488, N1485);
nor NOR2 (N1489, N1483, N1202);
and AND2 (N1490, N1478, N693);
xor XOR2 (N1491, N1488, N624);
nor NOR4 (N1492, N1472, N412, N96, N559);
xor XOR2 (N1493, N1484, N111);
not NOT1 (N1494, N1490);
xor XOR2 (N1495, N1487, N1063);
or OR3 (N1496, N1486, N192, N1048);
buf BUF1 (N1497, N1493);
xor XOR2 (N1498, N1496, N721);
xor XOR2 (N1499, N1492, N30);
or OR4 (N1500, N1476, N945, N88, N1302);
and AND3 (N1501, N1498, N941, N1096);
not NOT1 (N1502, N1494);
or OR4 (N1503, N1497, N125, N1302, N1452);
xor XOR2 (N1504, N1491, N451);
xor XOR2 (N1505, N1470, N1358);
nand NAND4 (N1506, N1495, N107, N1364, N684);
buf BUF1 (N1507, N1506);
nor NOR4 (N1508, N1481, N1451, N1193, N1207);
xor XOR2 (N1509, N1501, N99);
nand NAND3 (N1510, N1509, N177, N898);
nand NAND3 (N1511, N1507, N98, N259);
xor XOR2 (N1512, N1510, N1129);
and AND2 (N1513, N1500, N1163);
nor NOR3 (N1514, N1503, N557, N404);
buf BUF1 (N1515, N1512);
or OR4 (N1516, N1504, N32, N1347, N1435);
xor XOR2 (N1517, N1511, N327);
nand NAND4 (N1518, N1508, N912, N164, N671);
not NOT1 (N1519, N1513);
buf BUF1 (N1520, N1499);
nand NAND3 (N1521, N1517, N132, N1046);
and AND3 (N1522, N1489, N1262, N602);
and AND3 (N1523, N1518, N1377, N655);
nand NAND2 (N1524, N1521, N315);
xor XOR2 (N1525, N1520, N444);
not NOT1 (N1526, N1525);
and AND2 (N1527, N1505, N791);
buf BUF1 (N1528, N1502);
buf BUF1 (N1529, N1519);
not NOT1 (N1530, N1516);
buf BUF1 (N1531, N1529);
buf BUF1 (N1532, N1522);
xor XOR2 (N1533, N1523, N567);
buf BUF1 (N1534, N1514);
and AND4 (N1535, N1531, N188, N1148, N392);
xor XOR2 (N1536, N1515, N59);
nand NAND2 (N1537, N1536, N1392);
nand NAND4 (N1538, N1534, N112, N377, N1064);
buf BUF1 (N1539, N1538);
or OR4 (N1540, N1526, N1033, N772, N628);
or OR4 (N1541, N1540, N1193, N278, N1395);
not NOT1 (N1542, N1537);
nor NOR2 (N1543, N1539, N459);
not NOT1 (N1544, N1528);
nor NOR2 (N1545, N1542, N171);
buf BUF1 (N1546, N1530);
nor NOR3 (N1547, N1533, N1250, N838);
buf BUF1 (N1548, N1546);
nor NOR2 (N1549, N1543, N803);
buf BUF1 (N1550, N1547);
nor NOR3 (N1551, N1550, N1228, N831);
nand NAND3 (N1552, N1549, N733, N673);
or OR4 (N1553, N1552, N433, N1140, N567);
nand NAND4 (N1554, N1524, N19, N82, N249);
and AND4 (N1555, N1548, N498, N378, N1150);
xor XOR2 (N1556, N1553, N28);
xor XOR2 (N1557, N1544, N464);
nor NOR4 (N1558, N1541, N901, N858, N1277);
nand NAND2 (N1559, N1551, N546);
and AND3 (N1560, N1555, N1371, N906);
nand NAND2 (N1561, N1532, N1442);
xor XOR2 (N1562, N1560, N1198);
and AND3 (N1563, N1527, N751, N1174);
and AND4 (N1564, N1535, N645, N1308, N1087);
buf BUF1 (N1565, N1545);
or OR3 (N1566, N1563, N502, N1183);
nor NOR2 (N1567, N1556, N74);
xor XOR2 (N1568, N1558, N1340);
buf BUF1 (N1569, N1559);
nor NOR3 (N1570, N1569, N867, N348);
and AND2 (N1571, N1568, N798);
nor NOR4 (N1572, N1554, N924, N1539, N358);
or OR3 (N1573, N1572, N567, N1510);
nor NOR2 (N1574, N1562, N1113);
not NOT1 (N1575, N1565);
or OR3 (N1576, N1557, N838, N1452);
nand NAND4 (N1577, N1575, N212, N106, N800);
xor XOR2 (N1578, N1576, N1043);
nor NOR3 (N1579, N1561, N625, N1347);
nor NOR2 (N1580, N1567, N814);
or OR4 (N1581, N1571, N1196, N448, N108);
and AND2 (N1582, N1564, N1489);
xor XOR2 (N1583, N1580, N812);
not NOT1 (N1584, N1579);
buf BUF1 (N1585, N1570);
nor NOR4 (N1586, N1578, N1192, N1163, N363);
and AND2 (N1587, N1585, N1340);
not NOT1 (N1588, N1577);
nand NAND2 (N1589, N1582, N1145);
and AND3 (N1590, N1574, N983, N700);
buf BUF1 (N1591, N1590);
not NOT1 (N1592, N1587);
nor NOR3 (N1593, N1592, N478, N55);
buf BUF1 (N1594, N1581);
xor XOR2 (N1595, N1589, N1323);
nand NAND4 (N1596, N1586, N452, N212, N146);
buf BUF1 (N1597, N1588);
and AND2 (N1598, N1573, N640);
buf BUF1 (N1599, N1591);
or OR4 (N1600, N1566, N367, N807, N1113);
or OR2 (N1601, N1598, N1475);
nor NOR3 (N1602, N1595, N1423, N911);
nand NAND4 (N1603, N1597, N1397, N932, N906);
not NOT1 (N1604, N1603);
or OR4 (N1605, N1596, N1256, N1325, N1255);
or OR4 (N1606, N1583, N1343, N1222, N590);
nand NAND4 (N1607, N1606, N2, N495, N819);
and AND4 (N1608, N1605, N1355, N524, N1436);
nor NOR2 (N1609, N1604, N1399);
or OR4 (N1610, N1584, N1106, N608, N1561);
buf BUF1 (N1611, N1602);
nand NAND3 (N1612, N1609, N1155, N258);
not NOT1 (N1613, N1607);
or OR3 (N1614, N1610, N675, N198);
or OR2 (N1615, N1599, N873);
not NOT1 (N1616, N1614);
nor NOR4 (N1617, N1594, N729, N388, N904);
or OR2 (N1618, N1600, N1478);
and AND4 (N1619, N1616, N338, N1031, N1269);
or OR3 (N1620, N1618, N415, N347);
xor XOR2 (N1621, N1619, N1609);
nor NOR3 (N1622, N1620, N311, N1486);
and AND2 (N1623, N1593, N526);
xor XOR2 (N1624, N1612, N1376);
xor XOR2 (N1625, N1615, N365);
not NOT1 (N1626, N1625);
xor XOR2 (N1627, N1601, N271);
nand NAND2 (N1628, N1627, N242);
and AND2 (N1629, N1628, N1540);
nand NAND4 (N1630, N1617, N91, N1052, N57);
nand NAND3 (N1631, N1608, N751, N534);
nand NAND2 (N1632, N1611, N445);
buf BUF1 (N1633, N1621);
and AND2 (N1634, N1624, N1114);
nand NAND4 (N1635, N1634, N812, N1228, N1491);
nor NOR3 (N1636, N1631, N1547, N1114);
nor NOR2 (N1637, N1630, N1092);
or OR4 (N1638, N1636, N995, N1086, N347);
nand NAND3 (N1639, N1633, N1593, N656);
xor XOR2 (N1640, N1632, N257);
or OR2 (N1641, N1623, N1449);
or OR2 (N1642, N1641, N1461);
not NOT1 (N1643, N1638);
nand NAND4 (N1644, N1613, N1156, N1631, N659);
xor XOR2 (N1645, N1629, N888);
nand NAND2 (N1646, N1640, N622);
not NOT1 (N1647, N1645);
nand NAND4 (N1648, N1642, N1146, N616, N26);
nor NOR3 (N1649, N1646, N736, N1265);
not NOT1 (N1650, N1637);
buf BUF1 (N1651, N1622);
and AND4 (N1652, N1626, N1614, N849, N30);
xor XOR2 (N1653, N1649, N1602);
and AND2 (N1654, N1647, N1253);
nand NAND3 (N1655, N1639, N1374, N1538);
not NOT1 (N1656, N1655);
not NOT1 (N1657, N1653);
not NOT1 (N1658, N1654);
nand NAND2 (N1659, N1635, N552);
nor NOR4 (N1660, N1658, N1096, N37, N1252);
or OR2 (N1661, N1657, N1404);
or OR4 (N1662, N1648, N380, N830, N1163);
xor XOR2 (N1663, N1651, N1235);
xor XOR2 (N1664, N1643, N545);
or OR4 (N1665, N1661, N1058, N1194, N274);
xor XOR2 (N1666, N1652, N1323);
buf BUF1 (N1667, N1660);
nand NAND2 (N1668, N1644, N1511);
nor NOR4 (N1669, N1663, N1577, N1071, N1303);
buf BUF1 (N1670, N1650);
nor NOR3 (N1671, N1668, N609, N615);
and AND2 (N1672, N1669, N874);
nor NOR3 (N1673, N1666, N1080, N1356);
nor NOR2 (N1674, N1656, N409);
nor NOR3 (N1675, N1662, N341, N1174);
buf BUF1 (N1676, N1672);
buf BUF1 (N1677, N1673);
nand NAND2 (N1678, N1665, N100);
not NOT1 (N1679, N1659);
nor NOR2 (N1680, N1671, N124);
xor XOR2 (N1681, N1678, N1333);
nand NAND4 (N1682, N1680, N589, N1389, N927);
xor XOR2 (N1683, N1667, N43);
not NOT1 (N1684, N1681);
or OR2 (N1685, N1684, N131);
xor XOR2 (N1686, N1685, N602);
buf BUF1 (N1687, N1677);
nand NAND2 (N1688, N1686, N997);
and AND3 (N1689, N1675, N595, N214);
nor NOR2 (N1690, N1664, N1317);
buf BUF1 (N1691, N1690);
nand NAND4 (N1692, N1676, N271, N1427, N577);
xor XOR2 (N1693, N1691, N910);
not NOT1 (N1694, N1689);
xor XOR2 (N1695, N1693, N754);
nand NAND4 (N1696, N1687, N456, N41, N70);
buf BUF1 (N1697, N1670);
and AND4 (N1698, N1692, N1575, N357, N1006);
nor NOR4 (N1699, N1698, N453, N1520, N1125);
nand NAND2 (N1700, N1682, N61);
nand NAND4 (N1701, N1700, N501, N1050, N1160);
buf BUF1 (N1702, N1696);
nor NOR3 (N1703, N1701, N986, N1492);
not NOT1 (N1704, N1697);
nor NOR3 (N1705, N1688, N552, N194);
not NOT1 (N1706, N1702);
nor NOR4 (N1707, N1699, N1644, N1052, N1692);
or OR3 (N1708, N1674, N183, N967);
and AND3 (N1709, N1705, N1481, N812);
xor XOR2 (N1710, N1703, N1210);
and AND2 (N1711, N1683, N1205);
nor NOR3 (N1712, N1710, N604, N1267);
buf BUF1 (N1713, N1708);
and AND4 (N1714, N1694, N1544, N1140, N1327);
buf BUF1 (N1715, N1707);
and AND2 (N1716, N1679, N1016);
buf BUF1 (N1717, N1715);
or OR3 (N1718, N1716, N968, N803);
nor NOR3 (N1719, N1709, N1519, N1366);
nand NAND3 (N1720, N1706, N1152, N1437);
xor XOR2 (N1721, N1718, N548);
and AND4 (N1722, N1720, N451, N63, N332);
buf BUF1 (N1723, N1712);
and AND2 (N1724, N1719, N1477);
and AND4 (N1725, N1723, N1666, N934, N302);
and AND4 (N1726, N1721, N1332, N334, N1243);
xor XOR2 (N1727, N1714, N383);
buf BUF1 (N1728, N1713);
buf BUF1 (N1729, N1724);
or OR3 (N1730, N1725, N257, N146);
buf BUF1 (N1731, N1729);
buf BUF1 (N1732, N1722);
buf BUF1 (N1733, N1704);
xor XOR2 (N1734, N1733, N171);
buf BUF1 (N1735, N1727);
nand NAND2 (N1736, N1731, N1200);
nor NOR3 (N1737, N1730, N1721, N1161);
xor XOR2 (N1738, N1736, N23);
or OR4 (N1739, N1735, N421, N1231, N1082);
nor NOR2 (N1740, N1695, N1332);
or OR4 (N1741, N1738, N1090, N546, N1531);
and AND4 (N1742, N1726, N373, N419, N1315);
xor XOR2 (N1743, N1741, N1166);
and AND4 (N1744, N1732, N1177, N1137, N965);
not NOT1 (N1745, N1737);
not NOT1 (N1746, N1743);
and AND4 (N1747, N1744, N1645, N488, N943);
and AND4 (N1748, N1745, N1419, N1059, N1450);
and AND2 (N1749, N1728, N1444);
xor XOR2 (N1750, N1717, N1714);
buf BUF1 (N1751, N1734);
nor NOR2 (N1752, N1747, N285);
xor XOR2 (N1753, N1746, N1094);
nor NOR4 (N1754, N1750, N1032, N1239, N664);
nor NOR4 (N1755, N1749, N435, N1000, N540);
or OR4 (N1756, N1740, N470, N793, N1210);
and AND3 (N1757, N1739, N574, N219);
or OR4 (N1758, N1756, N1033, N1585, N1078);
nor NOR2 (N1759, N1758, N1464);
nand NAND2 (N1760, N1752, N1217);
xor XOR2 (N1761, N1760, N1128);
nor NOR2 (N1762, N1754, N1533);
and AND2 (N1763, N1753, N1204);
or OR3 (N1764, N1711, N405, N1672);
nor NOR3 (N1765, N1762, N1102, N1103);
nor NOR2 (N1766, N1763, N287);
nand NAND4 (N1767, N1748, N574, N1656, N1633);
buf BUF1 (N1768, N1765);
buf BUF1 (N1769, N1767);
nand NAND2 (N1770, N1751, N719);
xor XOR2 (N1771, N1755, N92);
buf BUF1 (N1772, N1761);
xor XOR2 (N1773, N1759, N128);
not NOT1 (N1774, N1766);
nand NAND4 (N1775, N1768, N1181, N1571, N958);
or OR3 (N1776, N1770, N1255, N745);
and AND3 (N1777, N1772, N932, N451);
xor XOR2 (N1778, N1771, N798);
nor NOR4 (N1779, N1742, N514, N1438, N380);
xor XOR2 (N1780, N1776, N669);
nand NAND3 (N1781, N1780, N1490, N1152);
xor XOR2 (N1782, N1778, N675);
buf BUF1 (N1783, N1764);
or OR4 (N1784, N1783, N201, N332, N1651);
nor NOR4 (N1785, N1777, N261, N392, N1321);
and AND3 (N1786, N1757, N1036, N1347);
nor NOR4 (N1787, N1784, N570, N1443, N1501);
nor NOR2 (N1788, N1782, N1312);
buf BUF1 (N1789, N1786);
buf BUF1 (N1790, N1779);
not NOT1 (N1791, N1769);
nor NOR4 (N1792, N1789, N238, N1233, N1584);
or OR2 (N1793, N1792, N545);
not NOT1 (N1794, N1791);
xor XOR2 (N1795, N1774, N922);
nand NAND3 (N1796, N1794, N104, N981);
nand NAND2 (N1797, N1785, N1580);
nor NOR2 (N1798, N1787, N1477);
or OR2 (N1799, N1775, N1649);
buf BUF1 (N1800, N1799);
and AND2 (N1801, N1781, N1085);
not NOT1 (N1802, N1793);
buf BUF1 (N1803, N1798);
not NOT1 (N1804, N1795);
and AND3 (N1805, N1801, N497, N1370);
xor XOR2 (N1806, N1788, N1039);
nor NOR2 (N1807, N1802, N273);
or OR3 (N1808, N1803, N1171, N585);
or OR3 (N1809, N1797, N997, N643);
nor NOR4 (N1810, N1804, N433, N119, N1076);
not NOT1 (N1811, N1806);
buf BUF1 (N1812, N1810);
and AND3 (N1813, N1808, N1520, N1286);
or OR2 (N1814, N1796, N999);
or OR4 (N1815, N1800, N1754, N446, N1128);
or OR2 (N1816, N1812, N1441);
buf BUF1 (N1817, N1813);
and AND3 (N1818, N1816, N596, N1369);
or OR4 (N1819, N1815, N1799, N1436, N335);
nor NOR2 (N1820, N1773, N1729);
nand NAND3 (N1821, N1819, N1609, N1407);
and AND4 (N1822, N1817, N811, N1552, N1236);
and AND4 (N1823, N1809, N125, N1715, N813);
nand NAND4 (N1824, N1822, N1308, N170, N708);
buf BUF1 (N1825, N1818);
nor NOR4 (N1826, N1805, N145, N1622, N1172);
buf BUF1 (N1827, N1807);
not NOT1 (N1828, N1814);
nor NOR4 (N1829, N1823, N754, N116, N985);
not NOT1 (N1830, N1821);
buf BUF1 (N1831, N1827);
nand NAND4 (N1832, N1820, N846, N957, N1492);
not NOT1 (N1833, N1825);
or OR2 (N1834, N1833, N511);
or OR4 (N1835, N1829, N401, N1641, N796);
xor XOR2 (N1836, N1835, N942);
buf BUF1 (N1837, N1831);
buf BUF1 (N1838, N1811);
xor XOR2 (N1839, N1828, N802);
nand NAND2 (N1840, N1834, N1157);
nand NAND2 (N1841, N1840, N1060);
xor XOR2 (N1842, N1832, N167);
nand NAND3 (N1843, N1824, N1746, N1266);
nor NOR2 (N1844, N1790, N639);
nand NAND2 (N1845, N1844, N614);
or OR2 (N1846, N1842, N544);
xor XOR2 (N1847, N1837, N47);
nor NOR4 (N1848, N1830, N1736, N1138, N1144);
nand NAND4 (N1849, N1845, N566, N1627, N1773);
not NOT1 (N1850, N1849);
nand NAND3 (N1851, N1826, N406, N744);
nand NAND2 (N1852, N1836, N345);
and AND3 (N1853, N1843, N1340, N557);
nor NOR4 (N1854, N1848, N1346, N1129, N1748);
or OR4 (N1855, N1838, N518, N1366, N364);
nor NOR3 (N1856, N1841, N1556, N1828);
and AND2 (N1857, N1852, N258);
nand NAND4 (N1858, N1853, N871, N1568, N1151);
xor XOR2 (N1859, N1846, N536);
nor NOR2 (N1860, N1855, N1638);
xor XOR2 (N1861, N1850, N77);
nand NAND2 (N1862, N1861, N1329);
not NOT1 (N1863, N1851);
nand NAND2 (N1864, N1857, N1396);
or OR2 (N1865, N1858, N1467);
buf BUF1 (N1866, N1847);
and AND2 (N1867, N1854, N137);
buf BUF1 (N1868, N1859);
and AND3 (N1869, N1867, N397, N638);
nor NOR2 (N1870, N1866, N1226);
not NOT1 (N1871, N1868);
and AND3 (N1872, N1863, N986, N381);
nand NAND3 (N1873, N1860, N46, N1838);
nor NOR4 (N1874, N1873, N1289, N554, N1314);
nor NOR3 (N1875, N1874, N1491, N982);
nor NOR3 (N1876, N1864, N664, N1725);
not NOT1 (N1877, N1872);
buf BUF1 (N1878, N1869);
buf BUF1 (N1879, N1856);
nand NAND4 (N1880, N1865, N1299, N379, N1823);
and AND2 (N1881, N1862, N587);
and AND3 (N1882, N1879, N17, N1779);
nor NOR4 (N1883, N1875, N274, N235, N1738);
xor XOR2 (N1884, N1883, N238);
and AND4 (N1885, N1870, N853, N31, N1566);
not NOT1 (N1886, N1839);
and AND3 (N1887, N1885, N1456, N1237);
not NOT1 (N1888, N1886);
nor NOR3 (N1889, N1881, N1691, N1182);
xor XOR2 (N1890, N1878, N709);
and AND4 (N1891, N1877, N1499, N761, N1423);
xor XOR2 (N1892, N1880, N397);
xor XOR2 (N1893, N1871, N193);
and AND3 (N1894, N1882, N34, N1013);
or OR4 (N1895, N1884, N1614, N1186, N328);
and AND2 (N1896, N1895, N189);
buf BUF1 (N1897, N1889);
buf BUF1 (N1898, N1891);
buf BUF1 (N1899, N1892);
nand NAND4 (N1900, N1888, N1076, N1354, N907);
nor NOR4 (N1901, N1898, N558, N1121, N1383);
nand NAND3 (N1902, N1876, N940, N764);
or OR2 (N1903, N1894, N1799);
nor NOR2 (N1904, N1890, N1772);
not NOT1 (N1905, N1897);
and AND3 (N1906, N1903, N57, N1641);
nor NOR3 (N1907, N1900, N1765, N1808);
and AND3 (N1908, N1896, N1773, N547);
and AND4 (N1909, N1887, N1626, N781, N286);
or OR4 (N1910, N1909, N412, N367, N103);
nor NOR2 (N1911, N1910, N946);
nor NOR2 (N1912, N1902, N1348);
xor XOR2 (N1913, N1908, N1857);
nand NAND4 (N1914, N1905, N110, N1572, N789);
nand NAND4 (N1915, N1912, N652, N1291, N1656);
buf BUF1 (N1916, N1914);
xor XOR2 (N1917, N1899, N601);
xor XOR2 (N1918, N1907, N181);
and AND4 (N1919, N1911, N1488, N1649, N1620);
or OR2 (N1920, N1917, N488);
not NOT1 (N1921, N1919);
buf BUF1 (N1922, N1918);
or OR3 (N1923, N1901, N1326, N778);
nor NOR3 (N1924, N1904, N470, N702);
nand NAND3 (N1925, N1906, N1738, N241);
and AND2 (N1926, N1920, N1094);
xor XOR2 (N1927, N1923, N937);
xor XOR2 (N1928, N1927, N247);
nor NOR3 (N1929, N1916, N1420, N979);
and AND3 (N1930, N1926, N1302, N545);
buf BUF1 (N1931, N1913);
not NOT1 (N1932, N1925);
xor XOR2 (N1933, N1932, N194);
not NOT1 (N1934, N1893);
or OR2 (N1935, N1929, N865);
not NOT1 (N1936, N1915);
buf BUF1 (N1937, N1924);
nand NAND3 (N1938, N1935, N1350, N187);
or OR4 (N1939, N1922, N1372, N1281, N265);
not NOT1 (N1940, N1936);
and AND2 (N1941, N1933, N1251);
or OR4 (N1942, N1930, N438, N1797, N872);
nand NAND4 (N1943, N1931, N618, N1054, N730);
not NOT1 (N1944, N1940);
nor NOR4 (N1945, N1934, N1546, N1049, N204);
xor XOR2 (N1946, N1945, N1687);
nand NAND4 (N1947, N1938, N1796, N1526, N474);
or OR2 (N1948, N1942, N714);
not NOT1 (N1949, N1941);
and AND2 (N1950, N1939, N1743);
nand NAND2 (N1951, N1949, N547);
xor XOR2 (N1952, N1950, N1324);
nor NOR4 (N1953, N1946, N22, N1486, N1444);
nor NOR4 (N1954, N1944, N1451, N819, N1773);
not NOT1 (N1955, N1948);
nor NOR4 (N1956, N1921, N1252, N816, N606);
nand NAND4 (N1957, N1943, N1385, N404, N650);
xor XOR2 (N1958, N1952, N160);
nand NAND2 (N1959, N1953, N1028);
and AND2 (N1960, N1947, N267);
not NOT1 (N1961, N1954);
and AND3 (N1962, N1951, N1155, N630);
xor XOR2 (N1963, N1958, N1638);
xor XOR2 (N1964, N1961, N429);
or OR2 (N1965, N1956, N1186);
or OR4 (N1966, N1963, N461, N1916, N202);
buf BUF1 (N1967, N1965);
or OR3 (N1968, N1937, N687, N400);
nor NOR4 (N1969, N1967, N1308, N847, N1761);
xor XOR2 (N1970, N1962, N363);
and AND2 (N1971, N1959, N127);
not NOT1 (N1972, N1971);
buf BUF1 (N1973, N1960);
buf BUF1 (N1974, N1928);
and AND2 (N1975, N1969, N130);
or OR2 (N1976, N1968, N297);
buf BUF1 (N1977, N1974);
xor XOR2 (N1978, N1973, N9);
nand NAND2 (N1979, N1978, N838);
buf BUF1 (N1980, N1977);
and AND3 (N1981, N1975, N1524, N851);
buf BUF1 (N1982, N1976);
nand NAND4 (N1983, N1982, N1603, N1410, N1472);
not NOT1 (N1984, N1980);
buf BUF1 (N1985, N1955);
buf BUF1 (N1986, N1964);
buf BUF1 (N1987, N1972);
and AND3 (N1988, N1957, N1032, N739);
and AND3 (N1989, N1985, N381, N115);
and AND3 (N1990, N1966, N94, N71);
nand NAND2 (N1991, N1987, N1752);
nor NOR2 (N1992, N1970, N329);
and AND3 (N1993, N1990, N1156, N537);
or OR3 (N1994, N1979, N731, N215);
nor NOR4 (N1995, N1993, N1372, N644, N1922);
nand NAND3 (N1996, N1981, N1226, N423);
nand NAND2 (N1997, N1984, N1084);
and AND2 (N1998, N1995, N658);
xor XOR2 (N1999, N1989, N181);
and AND4 (N2000, N1994, N17, N314, N979);
and AND4 (N2001, N1988, N1874, N555, N1861);
nand NAND3 (N2002, N2000, N924, N563);
not NOT1 (N2003, N1998);
and AND3 (N2004, N2003, N707, N723);
not NOT1 (N2005, N2004);
or OR3 (N2006, N1983, N1728, N387);
buf BUF1 (N2007, N1999);
and AND2 (N2008, N1986, N1850);
or OR3 (N2009, N2001, N884, N961);
not NOT1 (N2010, N2009);
not NOT1 (N2011, N1991);
xor XOR2 (N2012, N2007, N1373);
nor NOR3 (N2013, N2012, N564, N1869);
xor XOR2 (N2014, N1997, N400);
nor NOR2 (N2015, N2014, N1902);
nand NAND2 (N2016, N2002, N1229);
buf BUF1 (N2017, N2005);
and AND4 (N2018, N1996, N198, N1498, N1602);
nand NAND2 (N2019, N2016, N496);
not NOT1 (N2020, N2008);
and AND2 (N2021, N2013, N181);
buf BUF1 (N2022, N2006);
not NOT1 (N2023, N2011);
buf BUF1 (N2024, N2021);
and AND2 (N2025, N2017, N1069);
nand NAND3 (N2026, N1992, N660, N317);
or OR3 (N2027, N2026, N327, N1176);
xor XOR2 (N2028, N2027, N532);
or OR2 (N2029, N2022, N638);
and AND4 (N2030, N2028, N674, N260, N1377);
xor XOR2 (N2031, N2019, N480);
buf BUF1 (N2032, N2020);
and AND3 (N2033, N2010, N169, N1095);
xor XOR2 (N2034, N2031, N1847);
or OR4 (N2035, N2015, N1783, N1341, N1538);
buf BUF1 (N2036, N2025);
nand NAND2 (N2037, N2036, N712);
xor XOR2 (N2038, N2029, N1390);
buf BUF1 (N2039, N2023);
xor XOR2 (N2040, N2030, N1685);
buf BUF1 (N2041, N2039);
buf BUF1 (N2042, N2037);
and AND2 (N2043, N2041, N429);
buf BUF1 (N2044, N2040);
xor XOR2 (N2045, N2032, N212);
and AND3 (N2046, N2038, N516, N2014);
xor XOR2 (N2047, N2042, N1707);
and AND2 (N2048, N2045, N265);
xor XOR2 (N2049, N2018, N1264);
nand NAND4 (N2050, N2048, N1478, N1866, N1026);
and AND2 (N2051, N2043, N208);
not NOT1 (N2052, N2035);
not NOT1 (N2053, N2033);
and AND4 (N2054, N2046, N139, N965, N77);
nor NOR3 (N2055, N2047, N202, N1508);
xor XOR2 (N2056, N2051, N424);
or OR3 (N2057, N2055, N486, N517);
buf BUF1 (N2058, N2057);
not NOT1 (N2059, N2044);
or OR4 (N2060, N2059, N1713, N1384, N627);
nor NOR3 (N2061, N2056, N1723, N1600);
or OR3 (N2062, N2060, N1920, N1393);
and AND3 (N2063, N2062, N119, N333);
or OR2 (N2064, N2024, N757);
and AND3 (N2065, N2058, N112, N25);
or OR4 (N2066, N2050, N145, N1850, N1917);
and AND2 (N2067, N2061, N576);
nand NAND3 (N2068, N2064, N210, N876);
nor NOR4 (N2069, N2054, N1274, N674, N1824);
and AND2 (N2070, N2034, N1339);
xor XOR2 (N2071, N2053, N1402);
nor NOR4 (N2072, N2049, N1054, N639, N1630);
buf BUF1 (N2073, N2072);
nand NAND2 (N2074, N2067, N240);
and AND2 (N2075, N2071, N2072);
nand NAND3 (N2076, N2066, N4, N806);
not NOT1 (N2077, N2075);
xor XOR2 (N2078, N2065, N1287);
xor XOR2 (N2079, N2076, N872);
or OR3 (N2080, N2070, N1061, N1029);
and AND2 (N2081, N2074, N304);
nor NOR4 (N2082, N2063, N1923, N1681, N867);
or OR4 (N2083, N2080, N1421, N291, N244);
and AND4 (N2084, N2052, N1487, N1063, N764);
not NOT1 (N2085, N2082);
xor XOR2 (N2086, N2085, N793);
not NOT1 (N2087, N2086);
not NOT1 (N2088, N2078);
nor NOR2 (N2089, N2084, N757);
nor NOR3 (N2090, N2068, N1242, N1385);
xor XOR2 (N2091, N2077, N886);
not NOT1 (N2092, N2073);
nand NAND3 (N2093, N2069, N1851, N359);
or OR4 (N2094, N2089, N1028, N1921, N1598);
not NOT1 (N2095, N2091);
and AND4 (N2096, N2087, N419, N1796, N1128);
and AND3 (N2097, N2088, N1480, N645);
xor XOR2 (N2098, N2092, N2042);
or OR4 (N2099, N2090, N1107, N2017, N1996);
nor NOR3 (N2100, N2095, N1976, N479);
xor XOR2 (N2101, N2099, N1548);
or OR4 (N2102, N2101, N533, N1842, N1422);
buf BUF1 (N2103, N2100);
nand NAND3 (N2104, N2079, N1218, N284);
not NOT1 (N2105, N2083);
nor NOR2 (N2106, N2104, N1620);
buf BUF1 (N2107, N2093);
nor NOR4 (N2108, N2096, N1819, N18, N575);
or OR3 (N2109, N2094, N388, N1289);
or OR3 (N2110, N2097, N1478, N775);
not NOT1 (N2111, N2108);
and AND2 (N2112, N2105, N1614);
and AND3 (N2113, N2109, N442, N1830);
not NOT1 (N2114, N2113);
and AND2 (N2115, N2112, N1479);
buf BUF1 (N2116, N2081);
not NOT1 (N2117, N2115);
or OR4 (N2118, N2106, N1982, N712, N684);
nand NAND2 (N2119, N2118, N239);
and AND2 (N2120, N2116, N1988);
xor XOR2 (N2121, N2119, N217);
buf BUF1 (N2122, N2117);
buf BUF1 (N2123, N2111);
buf BUF1 (N2124, N2103);
xor XOR2 (N2125, N2098, N844);
nand NAND4 (N2126, N2120, N348, N864, N165);
buf BUF1 (N2127, N2126);
or OR3 (N2128, N2122, N589, N1005);
nor NOR4 (N2129, N2107, N1256, N423, N1579);
or OR4 (N2130, N2129, N1898, N435, N885);
nor NOR4 (N2131, N2128, N90, N224, N2054);
nor NOR2 (N2132, N2121, N880);
buf BUF1 (N2133, N2114);
nand NAND2 (N2134, N2123, N1110);
nand NAND3 (N2135, N2132, N1104, N1349);
and AND3 (N2136, N2102, N767, N1455);
nor NOR2 (N2137, N2127, N1466);
not NOT1 (N2138, N2136);
nor NOR2 (N2139, N2133, N1201);
buf BUF1 (N2140, N2130);
nor NOR2 (N2141, N2125, N1139);
xor XOR2 (N2142, N2141, N2039);
nand NAND2 (N2143, N2142, N1328);
nor NOR2 (N2144, N2131, N637);
nor NOR4 (N2145, N2140, N785, N1338, N421);
xor XOR2 (N2146, N2134, N2104);
not NOT1 (N2147, N2137);
and AND3 (N2148, N2135, N823, N1754);
buf BUF1 (N2149, N2148);
and AND3 (N2150, N2144, N851, N1623);
nand NAND4 (N2151, N2147, N756, N1365, N1861);
nand NAND3 (N2152, N2150, N525, N1119);
xor XOR2 (N2153, N2124, N1423);
buf BUF1 (N2154, N2146);
buf BUF1 (N2155, N2153);
nand NAND2 (N2156, N2155, N1284);
buf BUF1 (N2157, N2151);
xor XOR2 (N2158, N2110, N552);
buf BUF1 (N2159, N2158);
xor XOR2 (N2160, N2143, N757);
xor XOR2 (N2161, N2156, N1747);
nand NAND4 (N2162, N2145, N2123, N527, N1961);
nand NAND3 (N2163, N2162, N443, N612);
and AND4 (N2164, N2157, N1636, N350, N185);
nand NAND3 (N2165, N2154, N1688, N1346);
xor XOR2 (N2166, N2163, N1123);
and AND2 (N2167, N2159, N734);
buf BUF1 (N2168, N2165);
nor NOR4 (N2169, N2168, N1109, N664, N100);
buf BUF1 (N2170, N2169);
not NOT1 (N2171, N2149);
nand NAND2 (N2172, N2160, N1043);
nor NOR2 (N2173, N2171, N577);
not NOT1 (N2174, N2172);
buf BUF1 (N2175, N2166);
nor NOR3 (N2176, N2174, N819, N1792);
not NOT1 (N2177, N2138);
not NOT1 (N2178, N2175);
or OR2 (N2179, N2164, N122);
nand NAND3 (N2180, N2173, N1841, N1739);
or OR4 (N2181, N2170, N1, N34, N1220);
and AND3 (N2182, N2167, N1832, N819);
xor XOR2 (N2183, N2179, N1065);
buf BUF1 (N2184, N2182);
or OR3 (N2185, N2177, N880, N384);
or OR2 (N2186, N2183, N1127);
nand NAND4 (N2187, N2152, N1491, N1, N1813);
xor XOR2 (N2188, N2181, N1736);
and AND4 (N2189, N2180, N518, N177, N2178);
xor XOR2 (N2190, N1686, N856);
nor NOR2 (N2191, N2176, N139);
or OR4 (N2192, N2139, N1389, N1632, N739);
and AND2 (N2193, N2186, N692);
or OR2 (N2194, N2193, N1358);
xor XOR2 (N2195, N2191, N1329);
not NOT1 (N2196, N2185);
or OR3 (N2197, N2188, N886, N503);
not NOT1 (N2198, N2161);
and AND3 (N2199, N2196, N589, N757);
or OR4 (N2200, N2194, N132, N1031, N883);
or OR2 (N2201, N2189, N1782);
not NOT1 (N2202, N2195);
not NOT1 (N2203, N2184);
nor NOR4 (N2204, N2199, N1500, N1120, N1492);
not NOT1 (N2205, N2200);
or OR3 (N2206, N2201, N1925, N1143);
buf BUF1 (N2207, N2198);
buf BUF1 (N2208, N2204);
or OR3 (N2209, N2187, N465, N32);
or OR4 (N2210, N2207, N40, N2016, N1836);
not NOT1 (N2211, N2206);
and AND3 (N2212, N2192, N1863, N1864);
not NOT1 (N2213, N2205);
buf BUF1 (N2214, N2202);
nand NAND2 (N2215, N2197, N545);
nor NOR4 (N2216, N2203, N1740, N398, N703);
nand NAND4 (N2217, N2215, N1863, N435, N1561);
not NOT1 (N2218, N2211);
nor NOR4 (N2219, N2218, N489, N917, N696);
or OR2 (N2220, N2209, N2043);
and AND4 (N2221, N2220, N1404, N1485, N2057);
not NOT1 (N2222, N2221);
nand NAND2 (N2223, N2219, N1550);
buf BUF1 (N2224, N2216);
nor NOR2 (N2225, N2222, N1829);
and AND3 (N2226, N2208, N496, N421);
or OR2 (N2227, N2212, N1581);
xor XOR2 (N2228, N2210, N1311);
buf BUF1 (N2229, N2227);
nand NAND3 (N2230, N2223, N142, N1845);
xor XOR2 (N2231, N2190, N230);
or OR4 (N2232, N2231, N612, N145, N1513);
and AND4 (N2233, N2213, N1525, N1075, N2056);
buf BUF1 (N2234, N2230);
xor XOR2 (N2235, N2217, N192);
nand NAND4 (N2236, N2233, N811, N1480, N1611);
or OR3 (N2237, N2224, N122, N180);
not NOT1 (N2238, N2237);
buf BUF1 (N2239, N2226);
buf BUF1 (N2240, N2234);
nor NOR4 (N2241, N2214, N2010, N2155, N2042);
buf BUF1 (N2242, N2240);
buf BUF1 (N2243, N2229);
xor XOR2 (N2244, N2232, N518);
and AND2 (N2245, N2239, N31);
nand NAND2 (N2246, N2228, N1456);
buf BUF1 (N2247, N2244);
or OR2 (N2248, N2241, N545);
nand NAND2 (N2249, N2246, N1809);
nand NAND3 (N2250, N2248, N1145, N15);
and AND2 (N2251, N2242, N1227);
not NOT1 (N2252, N2235);
and AND4 (N2253, N2225, N1351, N2178, N2231);
or OR2 (N2254, N2252, N423);
and AND2 (N2255, N2253, N24);
or OR2 (N2256, N2250, N96);
not NOT1 (N2257, N2255);
xor XOR2 (N2258, N2245, N1941);
nand NAND3 (N2259, N2249, N2024, N434);
buf BUF1 (N2260, N2257);
or OR2 (N2261, N2247, N125);
and AND2 (N2262, N2256, N919);
and AND2 (N2263, N2243, N1381);
buf BUF1 (N2264, N2262);
not NOT1 (N2265, N2254);
xor XOR2 (N2266, N2263, N1160);
nor NOR2 (N2267, N2259, N1340);
buf BUF1 (N2268, N2236);
nor NOR3 (N2269, N2258, N366, N137);
not NOT1 (N2270, N2260);
and AND2 (N2271, N2267, N773);
buf BUF1 (N2272, N2265);
not NOT1 (N2273, N2251);
nand NAND2 (N2274, N2272, N100);
not NOT1 (N2275, N2274);
or OR2 (N2276, N2270, N1393);
or OR4 (N2277, N2268, N801, N102, N1064);
nand NAND4 (N2278, N2273, N1037, N894, N1076);
nor NOR3 (N2279, N2238, N341, N1981);
xor XOR2 (N2280, N2275, N550);
nor NOR3 (N2281, N2278, N1488, N1307);
or OR3 (N2282, N2279, N692, N712);
nand NAND2 (N2283, N2280, N1068);
or OR4 (N2284, N2271, N281, N103, N1498);
and AND4 (N2285, N2261, N524, N657, N384);
and AND3 (N2286, N2284, N1600, N900);
or OR4 (N2287, N2277, N1821, N1677, N1666);
not NOT1 (N2288, N2269);
and AND2 (N2289, N2264, N667);
xor XOR2 (N2290, N2286, N1183);
nor NOR2 (N2291, N2285, N1806);
and AND2 (N2292, N2288, N64);
nand NAND3 (N2293, N2266, N2038, N934);
xor XOR2 (N2294, N2282, N992);
buf BUF1 (N2295, N2292);
xor XOR2 (N2296, N2289, N1501);
xor XOR2 (N2297, N2293, N1824);
not NOT1 (N2298, N2281);
xor XOR2 (N2299, N2297, N1625);
or OR2 (N2300, N2287, N1351);
nor NOR3 (N2301, N2290, N2050, N42);
and AND2 (N2302, N2301, N2199);
and AND4 (N2303, N2294, N1092, N738, N1962);
not NOT1 (N2304, N2298);
not NOT1 (N2305, N2296);
nand NAND3 (N2306, N2305, N1579, N914);
nand NAND4 (N2307, N2291, N493, N799, N145);
xor XOR2 (N2308, N2304, N1755);
nor NOR4 (N2309, N2307, N1067, N2279, N1609);
and AND3 (N2310, N2302, N704, N791);
xor XOR2 (N2311, N2306, N1809);
not NOT1 (N2312, N2283);
buf BUF1 (N2313, N2312);
not NOT1 (N2314, N2303);
not NOT1 (N2315, N2300);
not NOT1 (N2316, N2276);
nand NAND4 (N2317, N2315, N1219, N1774, N1416);
nor NOR4 (N2318, N2314, N1298, N1275, N1255);
xor XOR2 (N2319, N2299, N74);
xor XOR2 (N2320, N2319, N819);
and AND2 (N2321, N2311, N844);
xor XOR2 (N2322, N2313, N2144);
nor NOR3 (N2323, N2318, N1742, N779);
nor NOR3 (N2324, N2316, N124, N2112);
or OR2 (N2325, N2310, N976);
buf BUF1 (N2326, N2317);
or OR3 (N2327, N2324, N2308, N1643);
buf BUF1 (N2328, N585);
and AND4 (N2329, N2323, N1080, N963, N2236);
or OR4 (N2330, N2325, N1219, N1468, N504);
buf BUF1 (N2331, N2295);
buf BUF1 (N2332, N2321);
nor NOR3 (N2333, N2329, N1018, N543);
nand NAND2 (N2334, N2333, N1542);
nand NAND2 (N2335, N2334, N252);
and AND4 (N2336, N2327, N788, N712, N2055);
and AND4 (N2337, N2330, N1059, N30, N933);
nand NAND3 (N2338, N2331, N2110, N570);
not NOT1 (N2339, N2332);
buf BUF1 (N2340, N2337);
buf BUF1 (N2341, N2328);
nor NOR3 (N2342, N2338, N1796, N2289);
not NOT1 (N2343, N2340);
buf BUF1 (N2344, N2309);
nor NOR2 (N2345, N2336, N2178);
or OR2 (N2346, N2344, N1163);
buf BUF1 (N2347, N2326);
buf BUF1 (N2348, N2341);
and AND2 (N2349, N2339, N1687);
nor NOR2 (N2350, N2320, N1283);
buf BUF1 (N2351, N2346);
or OR2 (N2352, N2343, N1197);
nand NAND2 (N2353, N2342, N687);
buf BUF1 (N2354, N2353);
xor XOR2 (N2355, N2349, N625);
xor XOR2 (N2356, N2322, N2328);
not NOT1 (N2357, N2356);
nand NAND3 (N2358, N2355, N2210, N456);
or OR2 (N2359, N2350, N2141);
xor XOR2 (N2360, N2347, N201);
xor XOR2 (N2361, N2354, N991);
and AND2 (N2362, N2358, N23);
and AND3 (N2363, N2359, N2290, N2208);
nand NAND2 (N2364, N2361, N1100);
and AND4 (N2365, N2351, N1274, N187, N233);
not NOT1 (N2366, N2352);
buf BUF1 (N2367, N2357);
not NOT1 (N2368, N2363);
or OR2 (N2369, N2348, N1213);
or OR4 (N2370, N2362, N63, N2140, N1972);
nor NOR3 (N2371, N2368, N1492, N297);
not NOT1 (N2372, N2360);
nand NAND4 (N2373, N2367, N40, N838, N1487);
xor XOR2 (N2374, N2373, N565);
xor XOR2 (N2375, N2335, N1643);
not NOT1 (N2376, N2364);
not NOT1 (N2377, N2376);
buf BUF1 (N2378, N2345);
not NOT1 (N2379, N2371);
not NOT1 (N2380, N2379);
xor XOR2 (N2381, N2369, N694);
nor NOR4 (N2382, N2377, N2079, N299, N1733);
buf BUF1 (N2383, N2378);
nor NOR3 (N2384, N2366, N1047, N2326);
buf BUF1 (N2385, N2381);
or OR3 (N2386, N2374, N1136, N1155);
nand NAND2 (N2387, N2370, N1312);
nor NOR3 (N2388, N2382, N1189, N423);
nor NOR3 (N2389, N2388, N1086, N672);
or OR4 (N2390, N2380, N722, N78, N1453);
nand NAND3 (N2391, N2375, N1101, N278);
or OR3 (N2392, N2372, N621, N969);
and AND3 (N2393, N2365, N1754, N1656);
xor XOR2 (N2394, N2387, N1470);
buf BUF1 (N2395, N2392);
buf BUF1 (N2396, N2395);
nand NAND4 (N2397, N2389, N769, N1312, N2025);
nor NOR3 (N2398, N2384, N2327, N441);
and AND3 (N2399, N2385, N1596, N1275);
and AND3 (N2400, N2397, N1758, N834);
or OR2 (N2401, N2390, N2215);
or OR3 (N2402, N2398, N653, N432);
or OR3 (N2403, N2399, N1292, N398);
xor XOR2 (N2404, N2393, N897);
and AND3 (N2405, N2402, N84, N283);
and AND3 (N2406, N2396, N251, N1140);
not NOT1 (N2407, N2401);
or OR2 (N2408, N2405, N880);
buf BUF1 (N2409, N2403);
buf BUF1 (N2410, N2394);
or OR3 (N2411, N2404, N1074, N1339);
nor NOR3 (N2412, N2406, N903, N1580);
or OR3 (N2413, N2400, N2166, N2024);
or OR2 (N2414, N2409, N2325);
not NOT1 (N2415, N2408);
nor NOR2 (N2416, N2413, N5);
buf BUF1 (N2417, N2412);
nor NOR2 (N2418, N2414, N692);
or OR3 (N2419, N2391, N325, N713);
buf BUF1 (N2420, N2407);
not NOT1 (N2421, N2411);
xor XOR2 (N2422, N2410, N2033);
not NOT1 (N2423, N2421);
nor NOR3 (N2424, N2420, N2335, N1518);
buf BUF1 (N2425, N2383);
buf BUF1 (N2426, N2423);
nand NAND2 (N2427, N2386, N735);
nand NAND3 (N2428, N2417, N1177, N764);
buf BUF1 (N2429, N2419);
or OR4 (N2430, N2422, N1408, N1880, N731);
and AND2 (N2431, N2418, N1625);
not NOT1 (N2432, N2427);
buf BUF1 (N2433, N2415);
or OR3 (N2434, N2429, N2115, N2237);
buf BUF1 (N2435, N2431);
buf BUF1 (N2436, N2416);
nand NAND3 (N2437, N2434, N1215, N1385);
buf BUF1 (N2438, N2428);
not NOT1 (N2439, N2424);
and AND2 (N2440, N2436, N470);
nand NAND4 (N2441, N2440, N1352, N1829, N1932);
not NOT1 (N2442, N2432);
not NOT1 (N2443, N2433);
and AND3 (N2444, N2430, N535, N1408);
and AND2 (N2445, N2442, N1057);
xor XOR2 (N2446, N2438, N1224);
and AND3 (N2447, N2435, N812, N677);
nor NOR3 (N2448, N2425, N1095, N1231);
and AND3 (N2449, N2445, N2403, N2068);
nand NAND2 (N2450, N2447, N1306);
buf BUF1 (N2451, N2448);
buf BUF1 (N2452, N2441);
nor NOR4 (N2453, N2452, N2328, N2332, N420);
buf BUF1 (N2454, N2439);
and AND3 (N2455, N2443, N1400, N1383);
xor XOR2 (N2456, N2437, N1391);
not NOT1 (N2457, N2449);
and AND2 (N2458, N2426, N253);
buf BUF1 (N2459, N2451);
and AND3 (N2460, N2450, N127, N690);
not NOT1 (N2461, N2444);
buf BUF1 (N2462, N2461);
not NOT1 (N2463, N2455);
or OR3 (N2464, N2459, N184, N2437);
not NOT1 (N2465, N2457);
or OR2 (N2466, N2465, N1903);
nand NAND4 (N2467, N2454, N2315, N2384, N1210);
nand NAND3 (N2468, N2456, N2188, N2338);
and AND4 (N2469, N2463, N1118, N1758, N2074);
nand NAND2 (N2470, N2462, N105);
not NOT1 (N2471, N2460);
not NOT1 (N2472, N2466);
buf BUF1 (N2473, N2469);
buf BUF1 (N2474, N2446);
xor XOR2 (N2475, N2464, N1614);
nor NOR4 (N2476, N2473, N2253, N2141, N1878);
or OR2 (N2477, N2472, N2358);
nor NOR3 (N2478, N2468, N1054, N885);
xor XOR2 (N2479, N2475, N1040);
not NOT1 (N2480, N2479);
not NOT1 (N2481, N2476);
or OR2 (N2482, N2467, N371);
nor NOR4 (N2483, N2458, N1423, N239, N666);
nand NAND2 (N2484, N2482, N2365);
and AND2 (N2485, N2453, N2115);
or OR3 (N2486, N2480, N1003, N2440);
nand NAND3 (N2487, N2471, N2041, N2339);
xor XOR2 (N2488, N2481, N213);
and AND2 (N2489, N2478, N1021);
nand NAND3 (N2490, N2470, N801, N372);
or OR3 (N2491, N2490, N604, N1622);
not NOT1 (N2492, N2484);
or OR4 (N2493, N2477, N869, N2068, N1854);
buf BUF1 (N2494, N2489);
not NOT1 (N2495, N2485);
xor XOR2 (N2496, N2491, N532);
not NOT1 (N2497, N2492);
and AND4 (N2498, N2494, N1176, N159, N2344);
not NOT1 (N2499, N2487);
and AND4 (N2500, N2496, N2063, N119, N1014);
nand NAND2 (N2501, N2497, N1029);
nor NOR4 (N2502, N2486, N226, N429, N800);
nor NOR4 (N2503, N2495, N1850, N820, N1758);
or OR3 (N2504, N2499, N272, N567);
buf BUF1 (N2505, N2488);
and AND3 (N2506, N2503, N1846, N2191);
nor NOR3 (N2507, N2506, N1296, N602);
nor NOR3 (N2508, N2504, N426, N1770);
and AND4 (N2509, N2500, N463, N2096, N1021);
nand NAND3 (N2510, N2502, N1843, N241);
buf BUF1 (N2511, N2501);
nand NAND3 (N2512, N2509, N778, N2400);
not NOT1 (N2513, N2508);
xor XOR2 (N2514, N2505, N433);
xor XOR2 (N2515, N2513, N57);
nand NAND4 (N2516, N2512, N1832, N2440, N782);
endmodule