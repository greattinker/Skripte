// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15;

output N4012,N4001,N4010,N4009,N4014,N4013,N4011,N3981,N4007,N4015;

nand NAND3 (N16, N12, N7, N7);
and AND2 (N17, N13, N9);
and AND4 (N18, N7, N10, N4, N9);
nor NOR4 (N19, N18, N18, N18, N4);
xor XOR2 (N20, N4, N8);
and AND4 (N21, N4, N2, N18, N18);
nand NAND2 (N22, N2, N17);
nor NOR4 (N23, N21, N5, N8, N1);
nor NOR4 (N24, N18, N2, N5, N2);
nor NOR3 (N25, N7, N23, N7);
nand NAND2 (N26, N14, N13);
nor NOR2 (N27, N9, N19);
or OR3 (N28, N10, N1, N18);
not NOT1 (N29, N4);
buf BUF1 (N30, N8);
not NOT1 (N31, N29);
nor NOR4 (N32, N31, N22, N25, N4);
not NOT1 (N33, N25);
not NOT1 (N34, N8);
not NOT1 (N35, N34);
xor XOR2 (N36, N20, N6);
or OR4 (N37, N32, N28, N5, N32);
and AND3 (N38, N9, N36, N19);
nor NOR3 (N39, N37, N15, N12);
and AND2 (N40, N11, N16);
and AND4 (N41, N38, N17, N1, N37);
nor NOR4 (N42, N2, N5, N12, N40);
and AND3 (N43, N36, N1, N18);
or OR3 (N44, N41, N28, N39);
xor XOR2 (N45, N25, N43);
nand NAND2 (N46, N2, N5);
and AND4 (N47, N26, N43, N45, N4);
nor NOR2 (N48, N18, N17);
or OR4 (N49, N33, N21, N35, N31);
not NOT1 (N50, N45);
xor XOR2 (N51, N46, N35);
and AND2 (N52, N42, N19);
nand NAND3 (N53, N50, N7, N45);
not NOT1 (N54, N49);
not NOT1 (N55, N27);
buf BUF1 (N56, N55);
not NOT1 (N57, N48);
buf BUF1 (N58, N24);
buf BUF1 (N59, N51);
nor NOR4 (N60, N56, N42, N30, N14);
or OR3 (N61, N36, N27, N59);
nand NAND2 (N62, N27, N54);
or OR4 (N63, N2, N6, N24, N4);
xor XOR2 (N64, N58, N49);
not NOT1 (N65, N57);
not NOT1 (N66, N44);
and AND3 (N67, N53, N45, N9);
nor NOR4 (N68, N66, N40, N2, N66);
or OR2 (N69, N61, N68);
or OR4 (N70, N1, N27, N62, N40);
xor XOR2 (N71, N14, N9);
buf BUF1 (N72, N69);
or OR2 (N73, N60, N1);
or OR2 (N74, N73, N8);
nand NAND2 (N75, N70, N20);
or OR2 (N76, N67, N39);
xor XOR2 (N77, N52, N60);
and AND2 (N78, N64, N46);
nor NOR4 (N79, N71, N9, N37, N75);
or OR4 (N80, N10, N23, N52, N42);
not NOT1 (N81, N79);
buf BUF1 (N82, N78);
not NOT1 (N83, N63);
nand NAND2 (N84, N83, N36);
nand NAND4 (N85, N77, N83, N10, N15);
or OR2 (N86, N82, N32);
nand NAND2 (N87, N84, N74);
and AND3 (N88, N69, N69, N10);
not NOT1 (N89, N86);
nor NOR4 (N90, N47, N63, N32, N10);
xor XOR2 (N91, N87, N75);
and AND2 (N92, N90, N57);
or OR3 (N93, N65, N30, N92);
xor XOR2 (N94, N31, N90);
nand NAND4 (N95, N91, N16, N90, N71);
xor XOR2 (N96, N81, N10);
buf BUF1 (N97, N80);
or OR2 (N98, N94, N43);
and AND2 (N99, N95, N52);
xor XOR2 (N100, N99, N24);
nor NOR4 (N101, N97, N72, N99, N21);
and AND3 (N102, N3, N26, N43);
and AND3 (N103, N76, N94, N92);
nand NAND3 (N104, N93, N24, N57);
xor XOR2 (N105, N98, N5);
nand NAND4 (N106, N101, N74, N83, N5);
nand NAND2 (N107, N105, N35);
nor NOR3 (N108, N103, N9, N23);
xor XOR2 (N109, N107, N50);
nand NAND3 (N110, N108, N16, N17);
not NOT1 (N111, N110);
xor XOR2 (N112, N106, N91);
nor NOR3 (N113, N96, N77, N27);
nand NAND2 (N114, N102, N97);
and AND3 (N115, N113, N35, N90);
not NOT1 (N116, N104);
nor NOR4 (N117, N114, N82, N90, N22);
and AND2 (N118, N109, N69);
nand NAND4 (N119, N117, N3, N27, N9);
not NOT1 (N120, N112);
nor NOR4 (N121, N118, N32, N38, N85);
and AND4 (N122, N23, N39, N71, N93);
buf BUF1 (N123, N88);
or OR3 (N124, N119, N3, N60);
nand NAND4 (N125, N122, N70, N25, N55);
and AND3 (N126, N125, N121, N84);
xor XOR2 (N127, N59, N18);
xor XOR2 (N128, N120, N4);
and AND4 (N129, N111, N6, N75, N17);
or OR2 (N130, N127, N16);
nand NAND4 (N131, N130, N8, N106, N55);
buf BUF1 (N132, N123);
not NOT1 (N133, N128);
nor NOR4 (N134, N129, N34, N44, N83);
not NOT1 (N135, N132);
and AND2 (N136, N133, N22);
or OR3 (N137, N124, N20, N11);
and AND4 (N138, N136, N58, N137, N59);
xor XOR2 (N139, N83, N79);
and AND2 (N140, N89, N24);
or OR4 (N141, N116, N104, N137, N56);
nand NAND4 (N142, N115, N14, N47, N20);
nand NAND2 (N143, N139, N31);
nor NOR4 (N144, N134, N82, N133, N69);
nand NAND2 (N145, N131, N44);
and AND4 (N146, N126, N27, N141, N36);
or OR4 (N147, N109, N27, N63, N26);
and AND3 (N148, N143, N107, N33);
and AND2 (N149, N138, N2);
buf BUF1 (N150, N100);
or OR2 (N151, N149, N99);
or OR3 (N152, N146, N129, N13);
and AND3 (N153, N142, N9, N132);
nand NAND4 (N154, N152, N66, N57, N14);
buf BUF1 (N155, N150);
or OR2 (N156, N153, N90);
xor XOR2 (N157, N156, N1);
nor NOR3 (N158, N151, N123, N11);
or OR4 (N159, N155, N87, N98, N93);
nand NAND3 (N160, N148, N54, N40);
buf BUF1 (N161, N159);
buf BUF1 (N162, N144);
nor NOR3 (N163, N145, N99, N101);
or OR3 (N164, N158, N149, N10);
buf BUF1 (N165, N162);
nand NAND2 (N166, N163, N34);
and AND4 (N167, N166, N135, N127, N14);
nand NAND4 (N168, N149, N132, N91, N78);
buf BUF1 (N169, N154);
and AND2 (N170, N161, N52);
or OR3 (N171, N168, N40, N31);
or OR2 (N172, N167, N99);
xor XOR2 (N173, N147, N54);
not NOT1 (N174, N164);
nand NAND4 (N175, N174, N134, N30, N99);
and AND3 (N176, N165, N18, N36);
nor NOR4 (N177, N173, N8, N11, N34);
or OR4 (N178, N169, N46, N122, N19);
xor XOR2 (N179, N171, N152);
not NOT1 (N180, N140);
not NOT1 (N181, N172);
not NOT1 (N182, N180);
buf BUF1 (N183, N176);
or OR3 (N184, N183, N143, N123);
and AND4 (N185, N170, N168, N71, N96);
nor NOR4 (N186, N157, N75, N69, N81);
or OR3 (N187, N177, N171, N39);
nand NAND3 (N188, N179, N145, N152);
buf BUF1 (N189, N184);
not NOT1 (N190, N187);
xor XOR2 (N191, N160, N111);
and AND4 (N192, N190, N164, N184, N151);
not NOT1 (N193, N188);
nand NAND3 (N194, N189, N154, N114);
xor XOR2 (N195, N193, N3);
and AND4 (N196, N181, N82, N71, N91);
nor NOR4 (N197, N186, N179, N159, N156);
or OR3 (N198, N185, N130, N83);
nor NOR4 (N199, N197, N87, N122, N46);
and AND2 (N200, N194, N96);
or OR4 (N201, N192, N33, N176, N200);
and AND2 (N202, N182, N120);
nor NOR2 (N203, N89, N202);
nor NOR2 (N204, N15, N30);
not NOT1 (N205, N191);
or OR4 (N206, N201, N9, N5, N116);
nor NOR4 (N207, N203, N177, N58, N52);
not NOT1 (N208, N207);
xor XOR2 (N209, N204, N55);
nor NOR3 (N210, N199, N7, N111);
buf BUF1 (N211, N206);
buf BUF1 (N212, N205);
nand NAND4 (N213, N175, N149, N127, N101);
not NOT1 (N214, N209);
nand NAND2 (N215, N210, N153);
buf BUF1 (N216, N211);
not NOT1 (N217, N196);
not NOT1 (N218, N208);
and AND4 (N219, N212, N125, N208, N187);
xor XOR2 (N220, N195, N66);
buf BUF1 (N221, N198);
buf BUF1 (N222, N221);
nor NOR2 (N223, N219, N54);
nor NOR3 (N224, N213, N165, N204);
and AND2 (N225, N217, N137);
xor XOR2 (N226, N178, N51);
not NOT1 (N227, N215);
nor NOR2 (N228, N214, N70);
nor NOR2 (N229, N224, N137);
nand NAND2 (N230, N228, N57);
and AND2 (N231, N218, N47);
xor XOR2 (N232, N231, N76);
not NOT1 (N233, N216);
xor XOR2 (N234, N225, N173);
and AND4 (N235, N226, N17, N64, N112);
and AND2 (N236, N220, N68);
or OR3 (N237, N230, N29, N41);
nand NAND4 (N238, N237, N71, N75, N228);
not NOT1 (N239, N227);
and AND4 (N240, N232, N41, N140, N68);
nand NAND3 (N241, N229, N204, N162);
and AND2 (N242, N222, N228);
buf BUF1 (N243, N242);
buf BUF1 (N244, N235);
nor NOR3 (N245, N233, N39, N5);
xor XOR2 (N246, N241, N74);
not NOT1 (N247, N234);
xor XOR2 (N248, N223, N111);
xor XOR2 (N249, N244, N109);
and AND2 (N250, N243, N90);
or OR4 (N251, N236, N195, N52, N213);
buf BUF1 (N252, N239);
nor NOR2 (N253, N251, N94);
or OR4 (N254, N238, N145, N81, N158);
xor XOR2 (N255, N253, N171);
nand NAND4 (N256, N250, N148, N203, N35);
nand NAND4 (N257, N252, N142, N170, N129);
nor NOR4 (N258, N257, N31, N194, N206);
not NOT1 (N259, N245);
not NOT1 (N260, N258);
or OR3 (N261, N248, N203, N2);
not NOT1 (N262, N240);
or OR2 (N263, N255, N131);
and AND2 (N264, N256, N22);
and AND2 (N265, N264, N135);
not NOT1 (N266, N261);
not NOT1 (N267, N263);
and AND3 (N268, N259, N258, N132);
nor NOR3 (N269, N247, N214, N232);
buf BUF1 (N270, N249);
not NOT1 (N271, N254);
and AND4 (N272, N246, N224, N250, N72);
buf BUF1 (N273, N268);
buf BUF1 (N274, N260);
buf BUF1 (N275, N266);
nor NOR2 (N276, N270, N117);
or OR2 (N277, N273, N38);
nand NAND4 (N278, N276, N158, N81, N192);
not NOT1 (N279, N274);
nor NOR2 (N280, N262, N248);
and AND4 (N281, N279, N153, N101, N18);
nand NAND4 (N282, N269, N139, N128, N262);
or OR2 (N283, N271, N280);
buf BUF1 (N284, N87);
nor NOR4 (N285, N281, N54, N224, N80);
not NOT1 (N286, N277);
nand NAND4 (N287, N284, N244, N60, N90);
and AND2 (N288, N285, N223);
and AND3 (N289, N275, N36, N199);
nor NOR3 (N290, N289, N203, N54);
and AND2 (N291, N282, N52);
nor NOR3 (N292, N291, N266, N282);
and AND2 (N293, N288, N55);
nor NOR3 (N294, N267, N176, N137);
xor XOR2 (N295, N290, N287);
and AND3 (N296, N150, N83, N168);
nor NOR3 (N297, N293, N14, N180);
xor XOR2 (N298, N278, N200);
nand NAND4 (N299, N294, N289, N188, N186);
not NOT1 (N300, N295);
nor NOR3 (N301, N300, N298, N288);
nand NAND3 (N302, N119, N80, N234);
xor XOR2 (N303, N297, N49);
and AND4 (N304, N283, N213, N102, N127);
nor NOR2 (N305, N302, N160);
nand NAND4 (N306, N292, N67, N12, N183);
not NOT1 (N307, N306);
nor NOR2 (N308, N286, N119);
xor XOR2 (N309, N272, N169);
nand NAND3 (N310, N301, N223, N93);
xor XOR2 (N311, N307, N309);
not NOT1 (N312, N248);
buf BUF1 (N313, N312);
not NOT1 (N314, N265);
nand NAND2 (N315, N305, N99);
xor XOR2 (N316, N304, N225);
buf BUF1 (N317, N316);
nand NAND3 (N318, N296, N166, N153);
or OR2 (N319, N310, N14);
not NOT1 (N320, N317);
xor XOR2 (N321, N320, N312);
or OR3 (N322, N303, N168, N144);
or OR3 (N323, N314, N231, N139);
nor NOR3 (N324, N308, N306, N160);
nor NOR2 (N325, N299, N43);
nor NOR3 (N326, N321, N122, N10);
buf BUF1 (N327, N313);
nand NAND4 (N328, N322, N271, N81, N301);
not NOT1 (N329, N311);
or OR3 (N330, N329, N47, N16);
nand NAND2 (N331, N315, N313);
not NOT1 (N332, N326);
and AND2 (N333, N323, N99);
or OR4 (N334, N331, N125, N212, N110);
not NOT1 (N335, N327);
nor NOR4 (N336, N319, N324, N196, N327);
nor NOR4 (N337, N127, N318, N257, N159);
or OR2 (N338, N61, N255);
nor NOR3 (N339, N337, N171, N204);
or OR2 (N340, N333, N281);
nand NAND4 (N341, N328, N150, N285, N205);
nand NAND2 (N342, N341, N247);
nand NAND3 (N343, N342, N71, N129);
xor XOR2 (N344, N343, N305);
xor XOR2 (N345, N344, N140);
nand NAND3 (N346, N325, N343, N305);
nand NAND2 (N347, N336, N212);
or OR2 (N348, N340, N129);
nor NOR3 (N349, N335, N322, N30);
xor XOR2 (N350, N334, N347);
or OR4 (N351, N28, N125, N156, N308);
nand NAND4 (N352, N338, N211, N173, N37);
nand NAND3 (N353, N330, N283, N279);
not NOT1 (N354, N349);
and AND2 (N355, N348, N278);
nand NAND3 (N356, N353, N232, N234);
nand NAND2 (N357, N355, N75);
buf BUF1 (N358, N332);
nand NAND3 (N359, N356, N229, N76);
buf BUF1 (N360, N345);
nand NAND3 (N361, N339, N13, N245);
buf BUF1 (N362, N357);
and AND4 (N363, N351, N26, N186, N360);
or OR2 (N364, N263, N342);
nand NAND4 (N365, N352, N307, N51, N46);
xor XOR2 (N366, N362, N20);
nand NAND3 (N367, N364, N261, N236);
xor XOR2 (N368, N359, N10);
xor XOR2 (N369, N368, N247);
buf BUF1 (N370, N363);
not NOT1 (N371, N350);
buf BUF1 (N372, N370);
and AND4 (N373, N371, N182, N332, N311);
and AND4 (N374, N369, N236, N301, N205);
xor XOR2 (N375, N346, N116);
xor XOR2 (N376, N361, N352);
nor NOR2 (N377, N367, N20);
nand NAND2 (N378, N354, N311);
nand NAND2 (N379, N378, N120);
xor XOR2 (N380, N365, N66);
nor NOR2 (N381, N376, N27);
xor XOR2 (N382, N379, N75);
nand NAND3 (N383, N375, N367, N8);
xor XOR2 (N384, N383, N44);
not NOT1 (N385, N381);
buf BUF1 (N386, N374);
not NOT1 (N387, N377);
xor XOR2 (N388, N382, N328);
nand NAND3 (N389, N380, N88, N54);
xor XOR2 (N390, N387, N328);
nor NOR2 (N391, N384, N317);
nor NOR2 (N392, N390, N91);
and AND4 (N393, N366, N253, N148, N36);
not NOT1 (N394, N358);
xor XOR2 (N395, N388, N255);
nand NAND4 (N396, N373, N145, N337, N291);
xor XOR2 (N397, N393, N279);
xor XOR2 (N398, N392, N255);
buf BUF1 (N399, N386);
and AND2 (N400, N385, N378);
nor NOR4 (N401, N399, N388, N340, N110);
nor NOR2 (N402, N400, N313);
nor NOR2 (N403, N398, N310);
buf BUF1 (N404, N402);
or OR4 (N405, N395, N57, N262, N202);
buf BUF1 (N406, N397);
nor NOR3 (N407, N394, N124, N33);
nor NOR2 (N408, N389, N83);
not NOT1 (N409, N391);
nand NAND3 (N410, N407, N309, N170);
nor NOR4 (N411, N403, N255, N139, N2);
nor NOR3 (N412, N409, N107, N357);
not NOT1 (N413, N412);
and AND4 (N414, N404, N202, N383, N318);
nor NOR4 (N415, N408, N99, N377, N413);
nand NAND4 (N416, N331, N157, N267, N392);
nor NOR2 (N417, N415, N65);
or OR3 (N418, N406, N186, N85);
not NOT1 (N419, N418);
xor XOR2 (N420, N396, N305);
and AND2 (N421, N416, N80);
buf BUF1 (N422, N421);
or OR2 (N423, N419, N9);
nand NAND3 (N424, N401, N345, N326);
xor XOR2 (N425, N423, N150);
or OR2 (N426, N410, N376);
xor XOR2 (N427, N417, N240);
or OR3 (N428, N424, N183, N45);
nor NOR2 (N429, N427, N259);
not NOT1 (N430, N425);
or OR3 (N431, N372, N220, N252);
nand NAND3 (N432, N430, N145, N53);
not NOT1 (N433, N422);
xor XOR2 (N434, N414, N408);
buf BUF1 (N435, N411);
and AND3 (N436, N434, N137, N386);
buf BUF1 (N437, N426);
and AND4 (N438, N432, N321, N437, N59);
nand NAND4 (N439, N363, N2, N35, N345);
nand NAND4 (N440, N435, N344, N152, N150);
and AND4 (N441, N438, N319, N219, N37);
nor NOR4 (N442, N440, N184, N74, N403);
buf BUF1 (N443, N428);
buf BUF1 (N444, N443);
nand NAND4 (N445, N441, N343, N379, N348);
nand NAND4 (N446, N420, N42, N374, N259);
nand NAND2 (N447, N445, N25);
and AND3 (N448, N429, N273, N297);
buf BUF1 (N449, N448);
xor XOR2 (N450, N442, N163);
nor NOR2 (N451, N450, N163);
nor NOR3 (N452, N431, N254, N117);
xor XOR2 (N453, N449, N180);
nand NAND2 (N454, N405, N130);
nand NAND3 (N455, N436, N328, N150);
nor NOR3 (N456, N446, N206, N343);
xor XOR2 (N457, N447, N416);
nand NAND4 (N458, N452, N108, N139, N117);
and AND2 (N459, N457, N108);
nor NOR2 (N460, N455, N331);
xor XOR2 (N461, N453, N101);
or OR4 (N462, N444, N169, N21, N3);
buf BUF1 (N463, N459);
not NOT1 (N464, N454);
buf BUF1 (N465, N458);
nand NAND4 (N466, N451, N332, N261, N209);
buf BUF1 (N467, N439);
or OR4 (N468, N463, N442, N459, N317);
nor NOR4 (N469, N456, N196, N463, N422);
nor NOR4 (N470, N433, N108, N320, N404);
or OR3 (N471, N465, N330, N29);
xor XOR2 (N472, N469, N456);
buf BUF1 (N473, N460);
not NOT1 (N474, N471);
xor XOR2 (N475, N470, N165);
or OR3 (N476, N475, N124, N38);
nor NOR3 (N477, N476, N11, N414);
and AND4 (N478, N466, N398, N410, N157);
buf BUF1 (N479, N478);
xor XOR2 (N480, N472, N179);
and AND2 (N481, N474, N171);
nand NAND4 (N482, N462, N399, N266, N250);
nand NAND2 (N483, N461, N187);
and AND4 (N484, N473, N312, N221, N250);
and AND2 (N485, N467, N44);
nor NOR3 (N486, N481, N213, N213);
or OR3 (N487, N485, N481, N233);
nand NAND2 (N488, N483, N17);
buf BUF1 (N489, N479);
nand NAND2 (N490, N484, N43);
not NOT1 (N491, N488);
and AND2 (N492, N477, N323);
xor XOR2 (N493, N492, N459);
nand NAND2 (N494, N491, N236);
nand NAND4 (N495, N480, N325, N122, N479);
or OR4 (N496, N493, N25, N469, N102);
and AND4 (N497, N490, N321, N402, N217);
nor NOR3 (N498, N468, N468, N73);
or OR4 (N499, N464, N232, N343, N141);
buf BUF1 (N500, N496);
xor XOR2 (N501, N486, N285);
nor NOR4 (N502, N497, N5, N217, N125);
or OR3 (N503, N500, N309, N160);
or OR4 (N504, N495, N360, N389, N391);
nand NAND2 (N505, N489, N434);
nand NAND4 (N506, N487, N389, N342, N371);
and AND3 (N507, N505, N252, N231);
buf BUF1 (N508, N502);
nor NOR2 (N509, N507, N288);
or OR2 (N510, N501, N115);
and AND2 (N511, N498, N233);
nor NOR4 (N512, N506, N467, N47, N297);
nor NOR3 (N513, N508, N469, N277);
or OR3 (N514, N511, N429, N484);
and AND3 (N515, N509, N1, N88);
not NOT1 (N516, N512);
or OR3 (N517, N513, N313, N142);
nand NAND3 (N518, N514, N284, N462);
nor NOR2 (N519, N499, N365);
nor NOR2 (N520, N519, N433);
nand NAND4 (N521, N504, N272, N463, N5);
nand NAND4 (N522, N518, N62, N24, N236);
nand NAND3 (N523, N522, N468, N486);
buf BUF1 (N524, N523);
nand NAND2 (N525, N515, N58);
nand NAND3 (N526, N520, N319, N92);
xor XOR2 (N527, N510, N192);
or OR4 (N528, N482, N28, N129, N263);
buf BUF1 (N529, N525);
nand NAND2 (N530, N516, N422);
or OR2 (N531, N521, N490);
or OR2 (N532, N528, N476);
xor XOR2 (N533, N527, N404);
not NOT1 (N534, N517);
xor XOR2 (N535, N526, N11);
or OR4 (N536, N532, N289, N96, N391);
nand NAND3 (N537, N533, N66, N54);
nand NAND4 (N538, N530, N132, N202, N382);
nand NAND3 (N539, N536, N184, N354);
not NOT1 (N540, N538);
nor NOR3 (N541, N534, N169, N435);
buf BUF1 (N542, N541);
buf BUF1 (N543, N503);
and AND4 (N544, N531, N12, N181, N491);
or OR4 (N545, N542, N389, N336, N278);
nor NOR2 (N546, N524, N447);
or OR2 (N547, N535, N454);
and AND2 (N548, N540, N379);
buf BUF1 (N549, N529);
or OR2 (N550, N545, N374);
buf BUF1 (N551, N548);
or OR4 (N552, N547, N239, N428, N334);
or OR3 (N553, N551, N545, N36);
nor NOR3 (N554, N546, N85, N397);
nand NAND3 (N555, N552, N461, N482);
or OR4 (N556, N550, N531, N456, N23);
buf BUF1 (N557, N539);
or OR4 (N558, N549, N358, N380, N216);
or OR2 (N559, N537, N303);
or OR2 (N560, N553, N471);
xor XOR2 (N561, N543, N187);
nor NOR3 (N562, N559, N117, N159);
xor XOR2 (N563, N562, N188);
and AND2 (N564, N555, N176);
and AND4 (N565, N554, N136, N39, N262);
and AND3 (N566, N561, N7, N22);
not NOT1 (N567, N544);
nand NAND4 (N568, N556, N538, N63, N65);
not NOT1 (N569, N564);
and AND2 (N570, N568, N195);
nand NAND4 (N571, N567, N71, N534, N388);
xor XOR2 (N572, N558, N519);
nand NAND3 (N573, N571, N353, N423);
buf BUF1 (N574, N566);
nor NOR4 (N575, N570, N550, N31, N376);
not NOT1 (N576, N569);
buf BUF1 (N577, N563);
not NOT1 (N578, N576);
nor NOR4 (N579, N574, N3, N430, N218);
nand NAND2 (N580, N560, N496);
nand NAND3 (N581, N557, N304, N563);
nand NAND2 (N582, N581, N252);
and AND3 (N583, N577, N475, N113);
buf BUF1 (N584, N578);
not NOT1 (N585, N582);
nor NOR3 (N586, N580, N584, N242);
nand NAND4 (N587, N43, N61, N539, N534);
nand NAND3 (N588, N583, N364, N323);
buf BUF1 (N589, N575);
nor NOR4 (N590, N586, N407, N131, N307);
nor NOR4 (N591, N573, N45, N548, N148);
or OR4 (N592, N590, N183, N317, N76);
not NOT1 (N593, N572);
buf BUF1 (N594, N585);
or OR2 (N595, N592, N593);
not NOT1 (N596, N78);
xor XOR2 (N597, N594, N518);
nor NOR2 (N598, N588, N458);
or OR2 (N599, N589, N583);
nand NAND3 (N600, N565, N95, N497);
or OR3 (N601, N595, N354, N38);
buf BUF1 (N602, N591);
xor XOR2 (N603, N494, N365);
or OR4 (N604, N598, N343, N83, N452);
or OR2 (N605, N602, N153);
and AND3 (N606, N604, N460, N140);
buf BUF1 (N607, N603);
xor XOR2 (N608, N600, N144);
nor NOR2 (N609, N599, N234);
or OR2 (N610, N606, N38);
nor NOR4 (N611, N608, N428, N494, N192);
nand NAND3 (N612, N611, N534, N1);
not NOT1 (N613, N601);
nand NAND3 (N614, N612, N570, N495);
not NOT1 (N615, N596);
buf BUF1 (N616, N614);
nand NAND3 (N617, N587, N524, N407);
nand NAND3 (N618, N597, N162, N449);
not NOT1 (N619, N615);
xor XOR2 (N620, N609, N60);
nor NOR3 (N621, N605, N13, N569);
buf BUF1 (N622, N579);
and AND3 (N623, N622, N114, N294);
xor XOR2 (N624, N610, N155);
and AND3 (N625, N616, N432, N401);
buf BUF1 (N626, N624);
nor NOR2 (N627, N626, N519);
nand NAND3 (N628, N627, N340, N442);
and AND4 (N629, N619, N584, N323, N553);
buf BUF1 (N630, N625);
nand NAND3 (N631, N623, N336, N43);
buf BUF1 (N632, N628);
and AND3 (N633, N620, N504, N138);
nor NOR4 (N634, N618, N630, N299, N465);
nor NOR2 (N635, N277, N40);
buf BUF1 (N636, N631);
or OR4 (N637, N632, N421, N333, N157);
nand NAND3 (N638, N617, N1, N520);
not NOT1 (N639, N613);
not NOT1 (N640, N635);
buf BUF1 (N641, N629);
nand NAND2 (N642, N639, N134);
xor XOR2 (N643, N641, N637);
buf BUF1 (N644, N563);
nor NOR2 (N645, N644, N450);
buf BUF1 (N646, N621);
nand NAND2 (N647, N633, N6);
xor XOR2 (N648, N642, N76);
or OR3 (N649, N638, N615, N342);
and AND3 (N650, N640, N381, N59);
nor NOR3 (N651, N646, N134, N295);
xor XOR2 (N652, N650, N326);
buf BUF1 (N653, N651);
nand NAND3 (N654, N649, N560, N319);
nand NAND4 (N655, N654, N167, N149, N48);
not NOT1 (N656, N647);
or OR4 (N657, N656, N577, N165, N208);
nor NOR2 (N658, N643, N355);
buf BUF1 (N659, N652);
nand NAND2 (N660, N655, N353);
not NOT1 (N661, N657);
not NOT1 (N662, N634);
xor XOR2 (N663, N661, N600);
nand NAND2 (N664, N645, N253);
buf BUF1 (N665, N662);
buf BUF1 (N666, N664);
and AND4 (N667, N663, N252, N542, N109);
and AND4 (N668, N658, N387, N413, N477);
nand NAND2 (N669, N668, N435);
nand NAND2 (N670, N667, N3);
nand NAND4 (N671, N666, N108, N309, N630);
and AND4 (N672, N648, N393, N83, N96);
xor XOR2 (N673, N671, N324);
buf BUF1 (N674, N636);
xor XOR2 (N675, N659, N24);
nor NOR3 (N676, N672, N559, N466);
or OR4 (N677, N670, N435, N178, N117);
nand NAND4 (N678, N660, N78, N459, N186);
and AND3 (N679, N674, N353, N478);
and AND4 (N680, N653, N578, N376, N146);
or OR2 (N681, N677, N355);
not NOT1 (N682, N681);
and AND2 (N683, N680, N672);
nor NOR2 (N684, N673, N148);
nand NAND3 (N685, N683, N417, N359);
nor NOR4 (N686, N665, N128, N48, N574);
xor XOR2 (N687, N684, N408);
nor NOR4 (N688, N675, N460, N467, N128);
or OR3 (N689, N685, N592, N573);
or OR3 (N690, N689, N592, N204);
xor XOR2 (N691, N690, N116);
not NOT1 (N692, N676);
not NOT1 (N693, N669);
buf BUF1 (N694, N686);
nor NOR2 (N695, N679, N326);
xor XOR2 (N696, N682, N119);
nor NOR3 (N697, N688, N200, N160);
and AND3 (N698, N678, N685, N161);
not NOT1 (N699, N687);
not NOT1 (N700, N691);
xor XOR2 (N701, N607, N521);
nand NAND3 (N702, N694, N442, N388);
buf BUF1 (N703, N702);
not NOT1 (N704, N695);
buf BUF1 (N705, N696);
nand NAND2 (N706, N705, N366);
nor NOR3 (N707, N693, N598, N393);
or OR2 (N708, N692, N680);
nand NAND4 (N709, N698, N633, N381, N597);
and AND3 (N710, N700, N423, N97);
or OR4 (N711, N706, N615, N570, N66);
xor XOR2 (N712, N703, N276);
buf BUF1 (N713, N711);
xor XOR2 (N714, N709, N168);
and AND4 (N715, N697, N200, N228, N117);
xor XOR2 (N716, N714, N16);
nand NAND3 (N717, N708, N4, N604);
nand NAND4 (N718, N716, N401, N388, N676);
not NOT1 (N719, N713);
xor XOR2 (N720, N699, N414);
not NOT1 (N721, N720);
buf BUF1 (N722, N717);
or OR2 (N723, N710, N142);
nor NOR3 (N724, N704, N433, N637);
and AND4 (N725, N701, N650, N249, N328);
xor XOR2 (N726, N718, N182);
not NOT1 (N727, N707);
and AND2 (N728, N724, N544);
nor NOR2 (N729, N722, N517);
and AND4 (N730, N726, N292, N447, N326);
xor XOR2 (N731, N727, N624);
nor NOR2 (N732, N730, N117);
xor XOR2 (N733, N728, N579);
buf BUF1 (N734, N732);
buf BUF1 (N735, N719);
buf BUF1 (N736, N715);
and AND2 (N737, N731, N675);
nand NAND3 (N738, N734, N211, N245);
nand NAND3 (N739, N729, N347, N117);
or OR3 (N740, N712, N171, N408);
not NOT1 (N741, N721);
nand NAND4 (N742, N737, N550, N321, N257);
nand NAND2 (N743, N735, N480);
and AND3 (N744, N743, N574, N529);
nand NAND3 (N745, N740, N659, N439);
or OR2 (N746, N739, N258);
or OR2 (N747, N744, N152);
and AND4 (N748, N741, N280, N302, N289);
and AND4 (N749, N742, N509, N614, N265);
or OR3 (N750, N738, N320, N119);
and AND2 (N751, N749, N587);
nor NOR4 (N752, N750, N161, N579, N522);
and AND4 (N753, N747, N158, N82, N543);
and AND4 (N754, N751, N590, N130, N731);
and AND2 (N755, N748, N137);
xor XOR2 (N756, N723, N702);
nand NAND2 (N757, N746, N570);
xor XOR2 (N758, N757, N608);
buf BUF1 (N759, N725);
buf BUF1 (N760, N754);
nor NOR3 (N761, N736, N309, N647);
nor NOR2 (N762, N756, N269);
xor XOR2 (N763, N759, N541);
not NOT1 (N764, N758);
and AND3 (N765, N752, N484, N456);
buf BUF1 (N766, N764);
and AND3 (N767, N745, N614, N706);
or OR4 (N768, N753, N736, N680, N72);
and AND4 (N769, N767, N374, N740, N763);
and AND3 (N770, N356, N195, N435);
nor NOR3 (N771, N755, N709, N699);
or OR2 (N772, N762, N685);
not NOT1 (N773, N766);
nor NOR2 (N774, N773, N561);
or OR3 (N775, N733, N244, N110);
and AND4 (N776, N768, N529, N394, N224);
nand NAND3 (N777, N776, N237, N470);
buf BUF1 (N778, N765);
nand NAND3 (N779, N769, N95, N264);
and AND3 (N780, N760, N552, N424);
nor NOR4 (N781, N761, N349, N292, N229);
and AND3 (N782, N778, N218, N51);
buf BUF1 (N783, N775);
nor NOR2 (N784, N777, N477);
nand NAND4 (N785, N774, N83, N452, N781);
not NOT1 (N786, N374);
and AND3 (N787, N782, N730, N187);
not NOT1 (N788, N772);
buf BUF1 (N789, N770);
buf BUF1 (N790, N785);
nor NOR4 (N791, N789, N569, N39, N136);
xor XOR2 (N792, N784, N62);
and AND3 (N793, N788, N570, N611);
not NOT1 (N794, N793);
not NOT1 (N795, N794);
nor NOR2 (N796, N779, N498);
buf BUF1 (N797, N790);
or OR3 (N798, N771, N660, N413);
xor XOR2 (N799, N795, N35);
nand NAND4 (N800, N780, N263, N244, N612);
buf BUF1 (N801, N798);
buf BUF1 (N802, N791);
nor NOR3 (N803, N796, N204, N28);
and AND4 (N804, N783, N449, N503, N62);
xor XOR2 (N805, N803, N431);
nor NOR4 (N806, N802, N193, N529, N556);
or OR3 (N807, N805, N345, N13);
buf BUF1 (N808, N801);
not NOT1 (N809, N804);
buf BUF1 (N810, N786);
and AND4 (N811, N797, N403, N329, N213);
or OR2 (N812, N810, N34);
not NOT1 (N813, N809);
and AND3 (N814, N806, N633, N190);
buf BUF1 (N815, N814);
not NOT1 (N816, N787);
buf BUF1 (N817, N813);
nand NAND2 (N818, N816, N788);
nand NAND2 (N819, N792, N374);
or OR3 (N820, N800, N671, N331);
nor NOR3 (N821, N808, N621, N670);
nor NOR2 (N822, N807, N799);
and AND4 (N823, N461, N194, N586, N394);
nor NOR3 (N824, N822, N511, N247);
or OR2 (N825, N812, N424);
nor NOR3 (N826, N819, N529, N351);
not NOT1 (N827, N811);
nor NOR2 (N828, N826, N657);
not NOT1 (N829, N823);
nand NAND2 (N830, N827, N764);
nand NAND4 (N831, N820, N380, N714, N458);
or OR2 (N832, N815, N581);
xor XOR2 (N833, N825, N734);
xor XOR2 (N834, N830, N136);
nand NAND2 (N835, N828, N22);
and AND3 (N836, N834, N430, N524);
nor NOR4 (N837, N818, N202, N623, N653);
not NOT1 (N838, N829);
nor NOR2 (N839, N824, N141);
and AND4 (N840, N835, N509, N456, N463);
buf BUF1 (N841, N837);
nand NAND4 (N842, N841, N687, N838, N605);
xor XOR2 (N843, N808, N584);
nand NAND3 (N844, N831, N583, N218);
and AND3 (N845, N821, N68, N618);
or OR4 (N846, N844, N799, N558, N318);
nor NOR3 (N847, N843, N143, N597);
nand NAND2 (N848, N845, N485);
buf BUF1 (N849, N836);
not NOT1 (N850, N817);
nor NOR3 (N851, N846, N173, N389);
nand NAND4 (N852, N840, N810, N248, N579);
not NOT1 (N853, N849);
not NOT1 (N854, N842);
xor XOR2 (N855, N852, N264);
nand NAND2 (N856, N847, N177);
nand NAND4 (N857, N833, N195, N356, N100);
nand NAND4 (N858, N856, N48, N101, N675);
buf BUF1 (N859, N857);
and AND4 (N860, N854, N354, N497, N856);
or OR3 (N861, N853, N264, N186);
buf BUF1 (N862, N851);
not NOT1 (N863, N858);
and AND4 (N864, N859, N581, N111, N546);
not NOT1 (N865, N864);
or OR2 (N866, N865, N584);
xor XOR2 (N867, N855, N17);
nor NOR2 (N868, N860, N654);
nor NOR4 (N869, N862, N321, N76, N639);
xor XOR2 (N870, N868, N9);
and AND3 (N871, N869, N831, N213);
buf BUF1 (N872, N839);
not NOT1 (N873, N870);
nand NAND2 (N874, N871, N775);
or OR2 (N875, N867, N766);
xor XOR2 (N876, N861, N156);
not NOT1 (N877, N875);
or OR3 (N878, N850, N253, N156);
and AND3 (N879, N873, N699, N226);
buf BUF1 (N880, N872);
or OR2 (N881, N879, N47);
or OR3 (N882, N832, N613, N364);
nor NOR2 (N883, N848, N572);
nor NOR4 (N884, N881, N882, N339, N252);
or OR3 (N885, N162, N263, N428);
nand NAND4 (N886, N866, N640, N219, N20);
not NOT1 (N887, N878);
buf BUF1 (N888, N874);
nor NOR2 (N889, N877, N41);
xor XOR2 (N890, N889, N51);
or OR3 (N891, N885, N853, N23);
and AND2 (N892, N886, N206);
nor NOR3 (N893, N884, N467, N245);
xor XOR2 (N894, N890, N351);
buf BUF1 (N895, N891);
nor NOR3 (N896, N863, N585, N530);
and AND2 (N897, N893, N321);
or OR3 (N898, N888, N633, N39);
nor NOR3 (N899, N876, N827, N318);
or OR4 (N900, N897, N504, N714, N862);
nand NAND3 (N901, N887, N697, N86);
nor NOR2 (N902, N896, N309);
and AND4 (N903, N883, N825, N810, N673);
or OR3 (N904, N903, N231, N414);
not NOT1 (N905, N894);
nand NAND4 (N906, N901, N668, N500, N31);
and AND2 (N907, N902, N453);
nand NAND3 (N908, N906, N333, N121);
buf BUF1 (N909, N904);
xor XOR2 (N910, N908, N111);
nor NOR4 (N911, N899, N6, N780, N399);
nand NAND2 (N912, N909, N890);
nor NOR3 (N913, N892, N388, N107);
xor XOR2 (N914, N900, N268);
nor NOR3 (N915, N913, N4, N375);
nor NOR4 (N916, N914, N134, N799, N37);
nand NAND4 (N917, N910, N795, N759, N744);
buf BUF1 (N918, N905);
or OR2 (N919, N916, N188);
or OR2 (N920, N912, N872);
nor NOR4 (N921, N895, N835, N82, N220);
and AND4 (N922, N918, N79, N234, N526);
not NOT1 (N923, N911);
nor NOR3 (N924, N919, N776, N48);
or OR2 (N925, N880, N294);
and AND3 (N926, N923, N758, N385);
not NOT1 (N927, N922);
nand NAND3 (N928, N921, N421, N877);
nand NAND3 (N929, N920, N407, N326);
nand NAND2 (N930, N926, N220);
xor XOR2 (N931, N928, N292);
buf BUF1 (N932, N930);
or OR3 (N933, N929, N258, N530);
nand NAND4 (N934, N898, N444, N470, N870);
and AND4 (N935, N907, N53, N703, N42);
buf BUF1 (N936, N924);
xor XOR2 (N937, N925, N254);
nand NAND4 (N938, N933, N676, N207, N351);
nor NOR4 (N939, N936, N511, N119, N895);
and AND3 (N940, N937, N147, N612);
xor XOR2 (N941, N934, N584);
and AND3 (N942, N927, N637, N430);
nand NAND3 (N943, N941, N414, N287);
xor XOR2 (N944, N939, N79);
buf BUF1 (N945, N931);
xor XOR2 (N946, N940, N395);
xor XOR2 (N947, N915, N469);
nand NAND3 (N948, N946, N532, N615);
xor XOR2 (N949, N938, N228);
and AND3 (N950, N945, N574, N780);
not NOT1 (N951, N950);
not NOT1 (N952, N943);
not NOT1 (N953, N942);
nor NOR3 (N954, N917, N252, N54);
not NOT1 (N955, N932);
not NOT1 (N956, N955);
nor NOR3 (N957, N956, N842, N184);
or OR3 (N958, N944, N872, N683);
and AND3 (N959, N951, N428, N27);
and AND2 (N960, N959, N645);
or OR4 (N961, N948, N96, N37, N807);
and AND3 (N962, N957, N93, N437);
nand NAND3 (N963, N960, N424, N62);
nand NAND3 (N964, N963, N295, N153);
nand NAND4 (N965, N947, N884, N765, N654);
xor XOR2 (N966, N935, N857);
nor NOR3 (N967, N949, N395, N136);
nor NOR4 (N968, N966, N831, N500, N552);
and AND4 (N969, N964, N871, N963, N876);
nand NAND4 (N970, N962, N199, N808, N135);
nand NAND4 (N971, N968, N485, N168, N408);
nor NOR4 (N972, N970, N308, N675, N578);
xor XOR2 (N973, N965, N112);
and AND4 (N974, N953, N646, N763, N403);
buf BUF1 (N975, N967);
or OR2 (N976, N969, N19);
nor NOR4 (N977, N974, N887, N714, N387);
nor NOR3 (N978, N975, N936, N430);
not NOT1 (N979, N978);
or OR2 (N980, N961, N362);
not NOT1 (N981, N972);
nand NAND2 (N982, N971, N52);
xor XOR2 (N983, N976, N910);
and AND4 (N984, N973, N624, N759, N874);
nand NAND2 (N985, N983, N342);
or OR4 (N986, N977, N832, N746, N839);
buf BUF1 (N987, N984);
xor XOR2 (N988, N958, N495);
nor NOR2 (N989, N954, N185);
and AND4 (N990, N987, N7, N290, N673);
nor NOR3 (N991, N986, N628, N781);
or OR2 (N992, N990, N382);
or OR2 (N993, N982, N664);
not NOT1 (N994, N980);
nor NOR3 (N995, N952, N632, N280);
not NOT1 (N996, N995);
not NOT1 (N997, N994);
nand NAND2 (N998, N992, N27);
xor XOR2 (N999, N988, N84);
xor XOR2 (N1000, N989, N58);
and AND3 (N1001, N996, N745, N529);
not NOT1 (N1002, N993);
nor NOR2 (N1003, N985, N332);
buf BUF1 (N1004, N997);
not NOT1 (N1005, N998);
buf BUF1 (N1006, N1000);
buf BUF1 (N1007, N1005);
nand NAND3 (N1008, N981, N231, N136);
or OR4 (N1009, N1006, N288, N152, N13);
nor NOR4 (N1010, N999, N733, N695, N209);
or OR3 (N1011, N1003, N765, N468);
or OR3 (N1012, N1001, N823, N543);
or OR2 (N1013, N1012, N331);
and AND4 (N1014, N1002, N258, N946, N642);
or OR2 (N1015, N1010, N535);
or OR3 (N1016, N1009, N762, N784);
nand NAND4 (N1017, N991, N715, N348, N111);
buf BUF1 (N1018, N1013);
not NOT1 (N1019, N1008);
or OR2 (N1020, N1015, N548);
nor NOR4 (N1021, N1004, N630, N797, N391);
nor NOR4 (N1022, N1020, N201, N200, N260);
xor XOR2 (N1023, N979, N126);
nand NAND2 (N1024, N1007, N532);
nor NOR2 (N1025, N1017, N798);
and AND2 (N1026, N1021, N925);
xor XOR2 (N1027, N1019, N714);
xor XOR2 (N1028, N1011, N911);
xor XOR2 (N1029, N1026, N71);
xor XOR2 (N1030, N1029, N186);
or OR4 (N1031, N1023, N878, N885, N893);
not NOT1 (N1032, N1024);
and AND3 (N1033, N1016, N380, N121);
or OR4 (N1034, N1030, N314, N936, N207);
nor NOR3 (N1035, N1018, N628, N512);
xor XOR2 (N1036, N1028, N214);
not NOT1 (N1037, N1022);
or OR4 (N1038, N1035, N1017, N12, N1034);
xor XOR2 (N1039, N536, N442);
or OR3 (N1040, N1027, N868, N818);
nand NAND4 (N1041, N1036, N509, N997, N633);
nand NAND2 (N1042, N1025, N380);
nor NOR2 (N1043, N1039, N238);
not NOT1 (N1044, N1032);
not NOT1 (N1045, N1014);
buf BUF1 (N1046, N1031);
and AND4 (N1047, N1045, N757, N761, N93);
nor NOR4 (N1048, N1043, N959, N494, N2);
buf BUF1 (N1049, N1040);
or OR2 (N1050, N1044, N697);
nor NOR4 (N1051, N1046, N298, N544, N327);
xor XOR2 (N1052, N1038, N700);
nand NAND2 (N1053, N1052, N523);
not NOT1 (N1054, N1037);
nor NOR2 (N1055, N1041, N384);
nor NOR2 (N1056, N1049, N623);
or OR2 (N1057, N1055, N156);
buf BUF1 (N1058, N1051);
not NOT1 (N1059, N1042);
and AND4 (N1060, N1058, N1046, N160, N1031);
or OR4 (N1061, N1033, N638, N392, N712);
nor NOR2 (N1062, N1057, N83);
buf BUF1 (N1063, N1059);
xor XOR2 (N1064, N1062, N435);
nor NOR3 (N1065, N1048, N440, N570);
and AND2 (N1066, N1056, N480);
not NOT1 (N1067, N1054);
or OR3 (N1068, N1065, N336, N1006);
xor XOR2 (N1069, N1066, N259);
nor NOR2 (N1070, N1069, N412);
xor XOR2 (N1071, N1063, N358);
and AND4 (N1072, N1067, N207, N241, N3);
buf BUF1 (N1073, N1047);
xor XOR2 (N1074, N1050, N800);
nor NOR3 (N1075, N1068, N655, N914);
or OR2 (N1076, N1071, N686);
and AND2 (N1077, N1061, N187);
nand NAND2 (N1078, N1064, N62);
or OR2 (N1079, N1078, N969);
nand NAND4 (N1080, N1074, N633, N928, N225);
buf BUF1 (N1081, N1053);
xor XOR2 (N1082, N1072, N287);
not NOT1 (N1083, N1075);
or OR3 (N1084, N1076, N472, N897);
nand NAND4 (N1085, N1060, N709, N189, N723);
and AND3 (N1086, N1083, N163, N236);
buf BUF1 (N1087, N1080);
buf BUF1 (N1088, N1070);
or OR2 (N1089, N1081, N430);
not NOT1 (N1090, N1073);
nor NOR2 (N1091, N1084, N271);
nor NOR4 (N1092, N1088, N70, N125, N88);
buf BUF1 (N1093, N1089);
nor NOR2 (N1094, N1077, N433);
or OR3 (N1095, N1086, N1071, N626);
nor NOR4 (N1096, N1094, N987, N367, N747);
buf BUF1 (N1097, N1087);
buf BUF1 (N1098, N1092);
nand NAND2 (N1099, N1079, N848);
not NOT1 (N1100, N1099);
buf BUF1 (N1101, N1095);
nor NOR2 (N1102, N1090, N200);
or OR4 (N1103, N1100, N1070, N241, N354);
nor NOR2 (N1104, N1093, N88);
or OR2 (N1105, N1096, N956);
and AND4 (N1106, N1102, N486, N957, N97);
not NOT1 (N1107, N1105);
or OR2 (N1108, N1097, N297);
not NOT1 (N1109, N1107);
buf BUF1 (N1110, N1108);
buf BUF1 (N1111, N1104);
and AND2 (N1112, N1098, N417);
not NOT1 (N1113, N1111);
buf BUF1 (N1114, N1082);
xor XOR2 (N1115, N1091, N336);
xor XOR2 (N1116, N1106, N855);
buf BUF1 (N1117, N1116);
nor NOR2 (N1118, N1112, N136);
xor XOR2 (N1119, N1114, N55);
or OR3 (N1120, N1113, N1067, N992);
buf BUF1 (N1121, N1109);
not NOT1 (N1122, N1120);
nand NAND4 (N1123, N1117, N576, N613, N999);
xor XOR2 (N1124, N1101, N49);
and AND4 (N1125, N1118, N736, N130, N205);
nor NOR4 (N1126, N1115, N202, N960, N719);
or OR2 (N1127, N1119, N317);
buf BUF1 (N1128, N1123);
not NOT1 (N1129, N1124);
nor NOR3 (N1130, N1127, N479, N107);
buf BUF1 (N1131, N1125);
buf BUF1 (N1132, N1122);
buf BUF1 (N1133, N1121);
and AND2 (N1134, N1133, N979);
or OR4 (N1135, N1131, N1082, N778, N1128);
nand NAND2 (N1136, N133, N477);
nor NOR3 (N1137, N1132, N969, N588);
xor XOR2 (N1138, N1136, N384);
or OR2 (N1139, N1085, N510);
nor NOR2 (N1140, N1137, N311);
or OR2 (N1141, N1135, N432);
or OR2 (N1142, N1129, N377);
buf BUF1 (N1143, N1142);
and AND2 (N1144, N1134, N213);
buf BUF1 (N1145, N1141);
nand NAND3 (N1146, N1138, N947, N245);
buf BUF1 (N1147, N1146);
nand NAND3 (N1148, N1130, N275, N533);
and AND2 (N1149, N1126, N839);
or OR2 (N1150, N1145, N310);
nor NOR4 (N1151, N1140, N615, N694, N293);
buf BUF1 (N1152, N1143);
xor XOR2 (N1153, N1110, N506);
or OR2 (N1154, N1152, N117);
and AND3 (N1155, N1150, N384, N803);
not NOT1 (N1156, N1103);
nor NOR4 (N1157, N1139, N509, N1118, N723);
xor XOR2 (N1158, N1157, N1004);
not NOT1 (N1159, N1158);
not NOT1 (N1160, N1148);
xor XOR2 (N1161, N1151, N555);
and AND4 (N1162, N1147, N920, N898, N502);
or OR2 (N1163, N1160, N719);
xor XOR2 (N1164, N1156, N290);
nand NAND3 (N1165, N1159, N22, N813);
not NOT1 (N1166, N1162);
not NOT1 (N1167, N1153);
not NOT1 (N1168, N1154);
buf BUF1 (N1169, N1149);
xor XOR2 (N1170, N1155, N524);
xor XOR2 (N1171, N1169, N921);
nor NOR4 (N1172, N1166, N464, N573, N521);
nor NOR4 (N1173, N1172, N597, N8, N205);
nand NAND4 (N1174, N1170, N957, N788, N699);
buf BUF1 (N1175, N1163);
nor NOR4 (N1176, N1174, N104, N185, N768);
xor XOR2 (N1177, N1165, N865);
not NOT1 (N1178, N1167);
nor NOR3 (N1179, N1178, N985, N519);
not NOT1 (N1180, N1168);
buf BUF1 (N1181, N1161);
nand NAND4 (N1182, N1144, N741, N327, N731);
xor XOR2 (N1183, N1181, N609);
not NOT1 (N1184, N1176);
xor XOR2 (N1185, N1180, N1144);
or OR3 (N1186, N1179, N275, N956);
xor XOR2 (N1187, N1183, N313);
not NOT1 (N1188, N1173);
or OR4 (N1189, N1171, N274, N849, N409);
not NOT1 (N1190, N1189);
nand NAND2 (N1191, N1188, N464);
xor XOR2 (N1192, N1164, N347);
and AND4 (N1193, N1192, N57, N744, N232);
or OR2 (N1194, N1177, N65);
or OR2 (N1195, N1175, N704);
not NOT1 (N1196, N1193);
buf BUF1 (N1197, N1186);
buf BUF1 (N1198, N1184);
xor XOR2 (N1199, N1191, N85);
or OR3 (N1200, N1199, N490, N903);
or OR2 (N1201, N1197, N1057);
xor XOR2 (N1202, N1195, N958);
xor XOR2 (N1203, N1202, N1155);
and AND4 (N1204, N1190, N102, N482, N165);
not NOT1 (N1205, N1203);
xor XOR2 (N1206, N1185, N613);
or OR4 (N1207, N1206, N933, N157, N492);
nor NOR2 (N1208, N1200, N1001);
nand NAND3 (N1209, N1201, N330, N1068);
and AND4 (N1210, N1204, N1113, N802, N1172);
and AND3 (N1211, N1182, N715, N378);
not NOT1 (N1212, N1210);
nand NAND4 (N1213, N1207, N681, N1046, N1084);
not NOT1 (N1214, N1198);
not NOT1 (N1215, N1187);
and AND4 (N1216, N1211, N241, N646, N542);
xor XOR2 (N1217, N1196, N548);
nor NOR3 (N1218, N1215, N897, N319);
nor NOR3 (N1219, N1212, N369, N1216);
nor NOR4 (N1220, N1079, N45, N253, N294);
nand NAND4 (N1221, N1213, N380, N575, N820);
not NOT1 (N1222, N1194);
xor XOR2 (N1223, N1218, N472);
nor NOR3 (N1224, N1205, N1049, N409);
nand NAND4 (N1225, N1208, N1000, N507, N122);
buf BUF1 (N1226, N1225);
buf BUF1 (N1227, N1223);
and AND2 (N1228, N1221, N653);
or OR2 (N1229, N1220, N692);
nand NAND2 (N1230, N1228, N1106);
nor NOR2 (N1231, N1229, N1227);
or OR2 (N1232, N419, N1012);
and AND4 (N1233, N1222, N1130, N518, N494);
or OR3 (N1234, N1230, N633, N2);
and AND3 (N1235, N1224, N87, N962);
buf BUF1 (N1236, N1235);
nor NOR3 (N1237, N1233, N426, N608);
nor NOR4 (N1238, N1231, N1027, N460, N29);
nor NOR2 (N1239, N1219, N983);
and AND4 (N1240, N1236, N1189, N64, N353);
or OR4 (N1241, N1239, N1007, N207, N1135);
nor NOR4 (N1242, N1234, N242, N290, N1078);
or OR2 (N1243, N1226, N931);
nand NAND3 (N1244, N1232, N998, N829);
nand NAND2 (N1245, N1214, N796);
xor XOR2 (N1246, N1242, N543);
buf BUF1 (N1247, N1240);
nor NOR3 (N1248, N1238, N1056, N842);
or OR3 (N1249, N1217, N887, N751);
nand NAND2 (N1250, N1246, N58);
not NOT1 (N1251, N1245);
and AND4 (N1252, N1249, N496, N691, N1172);
or OR3 (N1253, N1209, N989, N1252);
nor NOR3 (N1254, N434, N30, N1251);
nor NOR4 (N1255, N1068, N1221, N987, N1082);
and AND3 (N1256, N1248, N240, N857);
buf BUF1 (N1257, N1255);
nor NOR4 (N1258, N1247, N582, N504, N242);
not NOT1 (N1259, N1244);
not NOT1 (N1260, N1257);
or OR4 (N1261, N1241, N911, N281, N563);
xor XOR2 (N1262, N1250, N1062);
nand NAND2 (N1263, N1254, N940);
or OR4 (N1264, N1261, N150, N254, N970);
or OR4 (N1265, N1262, N975, N1255, N96);
nand NAND3 (N1266, N1264, N311, N913);
and AND4 (N1267, N1259, N335, N373, N542);
buf BUF1 (N1268, N1263);
xor XOR2 (N1269, N1265, N622);
and AND4 (N1270, N1253, N831, N140, N249);
xor XOR2 (N1271, N1269, N350);
or OR2 (N1272, N1258, N1021);
not NOT1 (N1273, N1266);
buf BUF1 (N1274, N1256);
and AND4 (N1275, N1274, N916, N564, N794);
buf BUF1 (N1276, N1271);
nor NOR2 (N1277, N1273, N1012);
and AND3 (N1278, N1276, N455, N314);
not NOT1 (N1279, N1272);
and AND3 (N1280, N1237, N482, N39);
nor NOR3 (N1281, N1275, N228, N602);
and AND2 (N1282, N1267, N821);
and AND4 (N1283, N1260, N979, N545, N89);
or OR4 (N1284, N1243, N190, N713, N533);
xor XOR2 (N1285, N1279, N344);
nor NOR2 (N1286, N1270, N1227);
nor NOR2 (N1287, N1280, N1107);
xor XOR2 (N1288, N1281, N690);
nor NOR3 (N1289, N1278, N1154, N1246);
buf BUF1 (N1290, N1268);
nor NOR4 (N1291, N1290, N346, N212, N257);
nor NOR2 (N1292, N1277, N47);
nor NOR3 (N1293, N1288, N1056, N426);
buf BUF1 (N1294, N1283);
or OR3 (N1295, N1284, N1019, N1270);
and AND3 (N1296, N1289, N920, N747);
or OR3 (N1297, N1295, N1144, N325);
nand NAND2 (N1298, N1287, N254);
buf BUF1 (N1299, N1294);
not NOT1 (N1300, N1297);
and AND4 (N1301, N1285, N996, N1150, N2);
or OR3 (N1302, N1293, N230, N835);
xor XOR2 (N1303, N1296, N959);
buf BUF1 (N1304, N1299);
nor NOR3 (N1305, N1282, N545, N1045);
xor XOR2 (N1306, N1301, N1060);
and AND2 (N1307, N1298, N33);
nor NOR2 (N1308, N1292, N1009);
nand NAND2 (N1309, N1286, N584);
nor NOR4 (N1310, N1306, N763, N1141, N617);
or OR3 (N1311, N1291, N489, N1104);
or OR4 (N1312, N1311, N265, N1232, N770);
nand NAND4 (N1313, N1302, N1277, N394, N131);
xor XOR2 (N1314, N1305, N858);
nor NOR2 (N1315, N1312, N434);
or OR3 (N1316, N1307, N520, N146);
xor XOR2 (N1317, N1308, N930);
xor XOR2 (N1318, N1303, N115);
or OR4 (N1319, N1300, N1072, N672, N38);
or OR3 (N1320, N1318, N561, N758);
nor NOR2 (N1321, N1313, N865);
buf BUF1 (N1322, N1314);
or OR3 (N1323, N1319, N1093, N46);
xor XOR2 (N1324, N1315, N977);
or OR3 (N1325, N1309, N454, N148);
nand NAND3 (N1326, N1322, N53, N659);
or OR2 (N1327, N1320, N240);
and AND2 (N1328, N1316, N909);
nor NOR3 (N1329, N1326, N582, N1262);
buf BUF1 (N1330, N1325);
nand NAND2 (N1331, N1324, N127);
not NOT1 (N1332, N1329);
or OR3 (N1333, N1323, N472, N550);
buf BUF1 (N1334, N1304);
xor XOR2 (N1335, N1327, N1202);
nor NOR4 (N1336, N1335, N314, N670, N87);
nand NAND3 (N1337, N1332, N1065, N1186);
xor XOR2 (N1338, N1330, N45);
nor NOR2 (N1339, N1321, N206);
buf BUF1 (N1340, N1339);
nand NAND2 (N1341, N1338, N576);
and AND2 (N1342, N1337, N889);
not NOT1 (N1343, N1328);
and AND4 (N1344, N1340, N1094, N1044, N218);
buf BUF1 (N1345, N1310);
nand NAND3 (N1346, N1317, N781, N828);
xor XOR2 (N1347, N1334, N514);
not NOT1 (N1348, N1336);
not NOT1 (N1349, N1341);
xor XOR2 (N1350, N1331, N179);
nand NAND3 (N1351, N1342, N999, N830);
buf BUF1 (N1352, N1346);
nor NOR3 (N1353, N1333, N990, N478);
buf BUF1 (N1354, N1349);
not NOT1 (N1355, N1350);
nand NAND3 (N1356, N1351, N301, N343);
and AND4 (N1357, N1352, N465, N825, N436);
not NOT1 (N1358, N1355);
not NOT1 (N1359, N1347);
and AND2 (N1360, N1348, N915);
not NOT1 (N1361, N1359);
or OR3 (N1362, N1344, N668, N1301);
buf BUF1 (N1363, N1343);
nor NOR2 (N1364, N1357, N301);
nor NOR2 (N1365, N1353, N757);
or OR2 (N1366, N1365, N729);
not NOT1 (N1367, N1358);
buf BUF1 (N1368, N1367);
not NOT1 (N1369, N1366);
or OR4 (N1370, N1369, N1081, N642, N633);
or OR3 (N1371, N1356, N734, N791);
not NOT1 (N1372, N1364);
and AND2 (N1373, N1370, N177);
nand NAND2 (N1374, N1354, N287);
nor NOR2 (N1375, N1371, N709);
and AND2 (N1376, N1363, N482);
not NOT1 (N1377, N1345);
buf BUF1 (N1378, N1373);
nor NOR2 (N1379, N1372, N721);
buf BUF1 (N1380, N1378);
buf BUF1 (N1381, N1375);
nor NOR4 (N1382, N1362, N895, N700, N305);
nor NOR3 (N1383, N1374, N905, N221);
nand NAND4 (N1384, N1361, N77, N634, N1278);
not NOT1 (N1385, N1384);
or OR2 (N1386, N1381, N48);
xor XOR2 (N1387, N1379, N1311);
and AND3 (N1388, N1386, N1051, N404);
nor NOR3 (N1389, N1360, N475, N1077);
xor XOR2 (N1390, N1382, N1182);
nand NAND4 (N1391, N1368, N1156, N1179, N74);
xor XOR2 (N1392, N1380, N587);
not NOT1 (N1393, N1385);
buf BUF1 (N1394, N1393);
not NOT1 (N1395, N1390);
or OR4 (N1396, N1388, N1055, N960, N373);
or OR2 (N1397, N1392, N189);
xor XOR2 (N1398, N1389, N446);
buf BUF1 (N1399, N1377);
xor XOR2 (N1400, N1399, N335);
nand NAND4 (N1401, N1376, N571, N627, N988);
buf BUF1 (N1402, N1387);
xor XOR2 (N1403, N1401, N513);
xor XOR2 (N1404, N1403, N358);
nand NAND2 (N1405, N1383, N16);
xor XOR2 (N1406, N1391, N871);
nor NOR4 (N1407, N1396, N675, N458, N1048);
nand NAND3 (N1408, N1407, N1231, N160);
and AND4 (N1409, N1408, N930, N1240, N528);
xor XOR2 (N1410, N1395, N1312);
xor XOR2 (N1411, N1394, N810);
xor XOR2 (N1412, N1397, N575);
buf BUF1 (N1413, N1405);
not NOT1 (N1414, N1398);
and AND4 (N1415, N1402, N153, N1361, N338);
buf BUF1 (N1416, N1400);
not NOT1 (N1417, N1404);
and AND2 (N1418, N1413, N284);
or OR2 (N1419, N1410, N153);
and AND3 (N1420, N1414, N197, N121);
buf BUF1 (N1421, N1415);
xor XOR2 (N1422, N1406, N1122);
buf BUF1 (N1423, N1417);
or OR2 (N1424, N1419, N304);
or OR3 (N1425, N1418, N182, N293);
and AND3 (N1426, N1409, N768, N366);
buf BUF1 (N1427, N1425);
not NOT1 (N1428, N1422);
buf BUF1 (N1429, N1427);
buf BUF1 (N1430, N1429);
nand NAND3 (N1431, N1416, N734, N189);
xor XOR2 (N1432, N1421, N307);
and AND4 (N1433, N1426, N597, N834, N513);
nor NOR3 (N1434, N1433, N412, N18);
and AND2 (N1435, N1428, N959);
not NOT1 (N1436, N1432);
and AND4 (N1437, N1431, N1026, N596, N989);
nor NOR2 (N1438, N1412, N345);
and AND4 (N1439, N1430, N1036, N616, N1132);
buf BUF1 (N1440, N1435);
xor XOR2 (N1441, N1423, N1361);
nor NOR4 (N1442, N1440, N227, N1329, N574);
nand NAND3 (N1443, N1441, N1245, N1239);
nor NOR3 (N1444, N1443, N550, N743);
nor NOR3 (N1445, N1420, N401, N807);
not NOT1 (N1446, N1411);
or OR4 (N1447, N1445, N238, N744, N1309);
and AND2 (N1448, N1438, N256);
nor NOR2 (N1449, N1437, N628);
nand NAND3 (N1450, N1448, N476, N195);
nand NAND2 (N1451, N1446, N1287);
xor XOR2 (N1452, N1442, N251);
buf BUF1 (N1453, N1447);
not NOT1 (N1454, N1439);
nor NOR2 (N1455, N1424, N488);
buf BUF1 (N1456, N1454);
nand NAND3 (N1457, N1451, N317, N611);
or OR4 (N1458, N1456, N1062, N1292, N362);
nand NAND4 (N1459, N1453, N1001, N1098, N401);
or OR4 (N1460, N1444, N1326, N479, N184);
not NOT1 (N1461, N1459);
and AND2 (N1462, N1452, N554);
and AND2 (N1463, N1460, N1329);
buf BUF1 (N1464, N1434);
and AND4 (N1465, N1464, N30, N320, N1047);
nor NOR3 (N1466, N1463, N1427, N37);
xor XOR2 (N1467, N1458, N1277);
not NOT1 (N1468, N1466);
or OR3 (N1469, N1436, N1314, N1277);
buf BUF1 (N1470, N1467);
nand NAND2 (N1471, N1450, N572);
not NOT1 (N1472, N1455);
not NOT1 (N1473, N1471);
xor XOR2 (N1474, N1470, N865);
nand NAND4 (N1475, N1462, N467, N531, N571);
buf BUF1 (N1476, N1461);
xor XOR2 (N1477, N1449, N605);
and AND3 (N1478, N1457, N696, N91);
nand NAND2 (N1479, N1473, N672);
nand NAND3 (N1480, N1477, N252, N611);
xor XOR2 (N1481, N1474, N382);
nor NOR4 (N1482, N1465, N985, N3, N856);
not NOT1 (N1483, N1479);
not NOT1 (N1484, N1480);
nor NOR2 (N1485, N1472, N489);
buf BUF1 (N1486, N1476);
nand NAND2 (N1487, N1468, N1111);
and AND4 (N1488, N1478, N1260, N172, N1393);
nand NAND3 (N1489, N1469, N396, N245);
xor XOR2 (N1490, N1484, N404);
and AND2 (N1491, N1487, N1047);
not NOT1 (N1492, N1488);
nand NAND4 (N1493, N1492, N1047, N703, N915);
nor NOR4 (N1494, N1485, N1087, N949, N993);
buf BUF1 (N1495, N1490);
nand NAND3 (N1496, N1481, N1208, N23);
buf BUF1 (N1497, N1475);
buf BUF1 (N1498, N1482);
nand NAND4 (N1499, N1483, N1378, N349, N85);
and AND2 (N1500, N1497, N1262);
and AND2 (N1501, N1493, N782);
and AND2 (N1502, N1498, N527);
not NOT1 (N1503, N1495);
and AND4 (N1504, N1499, N635, N1366, N496);
nor NOR4 (N1505, N1503, N494, N1436, N1435);
xor XOR2 (N1506, N1486, N1271);
nor NOR4 (N1507, N1506, N1497, N1379, N658);
or OR3 (N1508, N1505, N1063, N743);
nand NAND3 (N1509, N1501, N258, N143);
nor NOR3 (N1510, N1509, N865, N752);
nand NAND2 (N1511, N1508, N1136);
xor XOR2 (N1512, N1489, N1008);
or OR2 (N1513, N1512, N119);
buf BUF1 (N1514, N1502);
or OR4 (N1515, N1504, N555, N1015, N570);
xor XOR2 (N1516, N1514, N77);
buf BUF1 (N1517, N1491);
nand NAND3 (N1518, N1507, N1469, N1097);
nor NOR2 (N1519, N1510, N984);
xor XOR2 (N1520, N1511, N1457);
xor XOR2 (N1521, N1516, N947);
not NOT1 (N1522, N1520);
and AND3 (N1523, N1522, N1384, N680);
not NOT1 (N1524, N1494);
buf BUF1 (N1525, N1500);
or OR2 (N1526, N1515, N1119);
xor XOR2 (N1527, N1521, N285);
xor XOR2 (N1528, N1517, N612);
and AND3 (N1529, N1527, N1521, N1121);
xor XOR2 (N1530, N1525, N1267);
not NOT1 (N1531, N1529);
nand NAND4 (N1532, N1530, N315, N1229, N112);
not NOT1 (N1533, N1496);
nand NAND3 (N1534, N1513, N1064, N453);
nand NAND2 (N1535, N1519, N638);
and AND2 (N1536, N1526, N464);
and AND3 (N1537, N1536, N1060, N222);
and AND4 (N1538, N1534, N1320, N1240, N934);
nor NOR3 (N1539, N1537, N1168, N112);
buf BUF1 (N1540, N1524);
nand NAND2 (N1541, N1533, N190);
not NOT1 (N1542, N1531);
nand NAND2 (N1543, N1518, N504);
not NOT1 (N1544, N1523);
nor NOR4 (N1545, N1538, N436, N1328, N620);
nand NAND3 (N1546, N1540, N1483, N1414);
or OR4 (N1547, N1535, N104, N954, N1338);
xor XOR2 (N1548, N1547, N638);
nor NOR2 (N1549, N1544, N1470);
nand NAND2 (N1550, N1532, N485);
or OR4 (N1551, N1545, N131, N453, N86);
xor XOR2 (N1552, N1551, N420);
buf BUF1 (N1553, N1542);
nand NAND2 (N1554, N1553, N516);
xor XOR2 (N1555, N1554, N352);
and AND4 (N1556, N1549, N1055, N34, N1294);
or OR4 (N1557, N1543, N554, N1404, N1374);
nand NAND3 (N1558, N1552, N1389, N350);
nor NOR4 (N1559, N1558, N1475, N902, N698);
buf BUF1 (N1560, N1528);
xor XOR2 (N1561, N1560, N875);
nand NAND4 (N1562, N1557, N1462, N826, N1364);
nor NOR2 (N1563, N1550, N1027);
nor NOR2 (N1564, N1548, N991);
nor NOR2 (N1565, N1563, N1274);
buf BUF1 (N1566, N1541);
not NOT1 (N1567, N1539);
or OR2 (N1568, N1556, N242);
buf BUF1 (N1569, N1555);
and AND4 (N1570, N1564, N1330, N1427, N93);
or OR2 (N1571, N1562, N1350);
xor XOR2 (N1572, N1561, N1429);
buf BUF1 (N1573, N1572);
buf BUF1 (N1574, N1568);
and AND2 (N1575, N1565, N1224);
xor XOR2 (N1576, N1546, N1141);
xor XOR2 (N1577, N1567, N678);
buf BUF1 (N1578, N1577);
buf BUF1 (N1579, N1573);
nand NAND2 (N1580, N1559, N37);
nand NAND3 (N1581, N1575, N1311, N1179);
nor NOR2 (N1582, N1570, N89);
buf BUF1 (N1583, N1569);
not NOT1 (N1584, N1582);
buf BUF1 (N1585, N1584);
or OR3 (N1586, N1566, N1558, N1401);
xor XOR2 (N1587, N1583, N1496);
and AND4 (N1588, N1578, N687, N849, N399);
and AND3 (N1589, N1579, N406, N579);
and AND3 (N1590, N1587, N1280, N1379);
xor XOR2 (N1591, N1576, N836);
or OR4 (N1592, N1581, N622, N1225, N979);
buf BUF1 (N1593, N1592);
or OR2 (N1594, N1588, N475);
or OR4 (N1595, N1580, N166, N511, N277);
not NOT1 (N1596, N1593);
or OR2 (N1597, N1571, N876);
not NOT1 (N1598, N1594);
not NOT1 (N1599, N1586);
or OR2 (N1600, N1596, N211);
xor XOR2 (N1601, N1574, N861);
nand NAND4 (N1602, N1591, N956, N717, N622);
buf BUF1 (N1603, N1589);
nand NAND4 (N1604, N1585, N512, N1220, N1560);
xor XOR2 (N1605, N1598, N1199);
and AND4 (N1606, N1604, N1202, N1542, N955);
buf BUF1 (N1607, N1590);
nor NOR2 (N1608, N1599, N930);
not NOT1 (N1609, N1595);
nor NOR4 (N1610, N1608, N1172, N213, N1170);
and AND2 (N1611, N1597, N1130);
xor XOR2 (N1612, N1602, N1068);
nand NAND2 (N1613, N1612, N866);
not NOT1 (N1614, N1605);
and AND2 (N1615, N1614, N8);
and AND3 (N1616, N1615, N1272, N1564);
not NOT1 (N1617, N1606);
or OR4 (N1618, N1616, N1529, N1155, N1291);
not NOT1 (N1619, N1613);
buf BUF1 (N1620, N1617);
nor NOR3 (N1621, N1620, N1037, N1264);
nand NAND4 (N1622, N1600, N1327, N1163, N818);
xor XOR2 (N1623, N1618, N1584);
buf BUF1 (N1624, N1609);
nand NAND4 (N1625, N1622, N1457, N1575, N1015);
not NOT1 (N1626, N1624);
or OR3 (N1627, N1603, N612, N115);
not NOT1 (N1628, N1607);
xor XOR2 (N1629, N1628, N581);
not NOT1 (N1630, N1610);
not NOT1 (N1631, N1625);
nor NOR3 (N1632, N1611, N731, N1564);
not NOT1 (N1633, N1627);
nor NOR4 (N1634, N1630, N145, N698, N85);
nand NAND4 (N1635, N1634, N1117, N1405, N843);
buf BUF1 (N1636, N1632);
or OR2 (N1637, N1623, N614);
buf BUF1 (N1638, N1631);
nand NAND2 (N1639, N1629, N933);
and AND4 (N1640, N1638, N542, N1283, N284);
nand NAND2 (N1641, N1619, N219);
xor XOR2 (N1642, N1637, N1114);
not NOT1 (N1643, N1635);
xor XOR2 (N1644, N1639, N637);
nand NAND3 (N1645, N1640, N479, N587);
and AND4 (N1646, N1643, N1194, N741, N886);
and AND4 (N1647, N1644, N780, N231, N1513);
and AND3 (N1648, N1633, N27, N1645);
buf BUF1 (N1649, N537);
not NOT1 (N1650, N1636);
or OR4 (N1651, N1601, N572, N1267, N1131);
or OR3 (N1652, N1621, N1109, N1081);
buf BUF1 (N1653, N1648);
and AND3 (N1654, N1626, N423, N593);
and AND3 (N1655, N1647, N521, N798);
buf BUF1 (N1656, N1652);
or OR3 (N1657, N1656, N325, N622);
not NOT1 (N1658, N1657);
not NOT1 (N1659, N1642);
and AND3 (N1660, N1649, N172, N529);
buf BUF1 (N1661, N1653);
nand NAND3 (N1662, N1650, N985, N218);
nand NAND3 (N1663, N1641, N1345, N452);
buf BUF1 (N1664, N1662);
buf BUF1 (N1665, N1655);
buf BUF1 (N1666, N1646);
nor NOR3 (N1667, N1665, N1553, N248);
nor NOR4 (N1668, N1654, N479, N199, N1193);
and AND3 (N1669, N1659, N1099, N1301);
not NOT1 (N1670, N1658);
nand NAND4 (N1671, N1660, N665, N784, N1565);
xor XOR2 (N1672, N1669, N1365);
buf BUF1 (N1673, N1672);
xor XOR2 (N1674, N1663, N789);
nand NAND3 (N1675, N1674, N908, N886);
nor NOR4 (N1676, N1661, N831, N1385, N90);
buf BUF1 (N1677, N1668);
and AND4 (N1678, N1664, N1098, N995, N1036);
nand NAND3 (N1679, N1677, N1319, N1372);
nand NAND2 (N1680, N1679, N1254);
nand NAND2 (N1681, N1673, N1083);
or OR4 (N1682, N1680, N1047, N1028, N1143);
buf BUF1 (N1683, N1676);
or OR4 (N1684, N1670, N195, N1165, N618);
nand NAND3 (N1685, N1684, N954, N565);
and AND4 (N1686, N1683, N1137, N758, N1357);
not NOT1 (N1687, N1685);
not NOT1 (N1688, N1678);
nor NOR4 (N1689, N1671, N258, N1023, N200);
not NOT1 (N1690, N1681);
and AND2 (N1691, N1682, N1416);
xor XOR2 (N1692, N1666, N615);
xor XOR2 (N1693, N1686, N1493);
not NOT1 (N1694, N1687);
or OR2 (N1695, N1694, N244);
not NOT1 (N1696, N1691);
nand NAND4 (N1697, N1692, N968, N1149, N1599);
nand NAND2 (N1698, N1696, N1125);
nor NOR4 (N1699, N1667, N1284, N25, N436);
nand NAND3 (N1700, N1698, N204, N651);
or OR2 (N1701, N1699, N163);
xor XOR2 (N1702, N1689, N516);
nor NOR3 (N1703, N1688, N1503, N1044);
xor XOR2 (N1704, N1701, N435);
or OR2 (N1705, N1651, N343);
and AND4 (N1706, N1703, N580, N1080, N482);
nor NOR3 (N1707, N1705, N1202, N909);
nor NOR4 (N1708, N1675, N669, N1681, N960);
xor XOR2 (N1709, N1697, N946);
xor XOR2 (N1710, N1706, N852);
nor NOR3 (N1711, N1690, N147, N1640);
buf BUF1 (N1712, N1695);
xor XOR2 (N1713, N1712, N751);
buf BUF1 (N1714, N1709);
nand NAND4 (N1715, N1702, N447, N399, N1163);
nor NOR2 (N1716, N1710, N640);
buf BUF1 (N1717, N1716);
xor XOR2 (N1718, N1704, N1684);
nor NOR2 (N1719, N1707, N923);
nor NOR4 (N1720, N1719, N1302, N365, N582);
buf BUF1 (N1721, N1711);
and AND3 (N1722, N1717, N1419, N1018);
buf BUF1 (N1723, N1713);
or OR4 (N1724, N1718, N1123, N413, N15);
not NOT1 (N1725, N1722);
not NOT1 (N1726, N1715);
xor XOR2 (N1727, N1720, N1613);
buf BUF1 (N1728, N1725);
nand NAND3 (N1729, N1714, N819, N1427);
and AND2 (N1730, N1724, N945);
nor NOR4 (N1731, N1708, N282, N563, N1260);
xor XOR2 (N1732, N1730, N1522);
buf BUF1 (N1733, N1723);
not NOT1 (N1734, N1721);
and AND4 (N1735, N1729, N76, N1061, N388);
or OR4 (N1736, N1700, N331, N1324, N1652);
not NOT1 (N1737, N1693);
nand NAND3 (N1738, N1733, N1260, N1307);
buf BUF1 (N1739, N1738);
and AND2 (N1740, N1737, N387);
or OR4 (N1741, N1735, N1173, N764, N1608);
not NOT1 (N1742, N1728);
or OR4 (N1743, N1731, N1411, N1632, N382);
or OR4 (N1744, N1727, N384, N1452, N567);
nand NAND4 (N1745, N1739, N889, N1318, N1427);
nor NOR4 (N1746, N1726, N882, N924, N465);
nand NAND2 (N1747, N1734, N301);
or OR4 (N1748, N1746, N708, N426, N623);
xor XOR2 (N1749, N1748, N1131);
or OR2 (N1750, N1740, N488);
and AND4 (N1751, N1747, N1655, N1655, N765);
not NOT1 (N1752, N1749);
xor XOR2 (N1753, N1742, N1203);
nand NAND4 (N1754, N1732, N210, N146, N402);
and AND2 (N1755, N1743, N1680);
buf BUF1 (N1756, N1755);
nand NAND2 (N1757, N1754, N529);
nand NAND2 (N1758, N1751, N652);
not NOT1 (N1759, N1752);
and AND4 (N1760, N1756, N1064, N1002, N1039);
not NOT1 (N1761, N1757);
buf BUF1 (N1762, N1744);
nand NAND3 (N1763, N1758, N984, N535);
nor NOR2 (N1764, N1763, N896);
nor NOR3 (N1765, N1762, N972, N856);
nor NOR2 (N1766, N1741, N1070);
or OR4 (N1767, N1761, N1358, N1212, N830);
and AND4 (N1768, N1753, N365, N114, N1568);
or OR4 (N1769, N1736, N966, N35, N1026);
and AND2 (N1770, N1767, N1586);
not NOT1 (N1771, N1769);
or OR4 (N1772, N1759, N947, N1320, N1685);
xor XOR2 (N1773, N1770, N1363);
nor NOR2 (N1774, N1768, N1470);
or OR3 (N1775, N1766, N819, N93);
not NOT1 (N1776, N1771);
or OR4 (N1777, N1750, N167, N568, N1360);
nor NOR3 (N1778, N1774, N1671, N1309);
nand NAND2 (N1779, N1775, N1280);
not NOT1 (N1780, N1777);
or OR4 (N1781, N1772, N563, N53, N1266);
buf BUF1 (N1782, N1776);
nand NAND4 (N1783, N1764, N1289, N1033, N984);
or OR2 (N1784, N1760, N529);
nand NAND4 (N1785, N1783, N341, N1573, N117);
xor XOR2 (N1786, N1781, N924);
buf BUF1 (N1787, N1780);
nand NAND2 (N1788, N1745, N1531);
nor NOR3 (N1789, N1788, N1288, N264);
xor XOR2 (N1790, N1789, N44);
and AND2 (N1791, N1785, N1758);
not NOT1 (N1792, N1787);
xor XOR2 (N1793, N1765, N1018);
nand NAND3 (N1794, N1786, N1323, N300);
xor XOR2 (N1795, N1778, N508);
buf BUF1 (N1796, N1790);
nand NAND4 (N1797, N1795, N45, N1023, N1324);
nand NAND2 (N1798, N1782, N1649);
and AND2 (N1799, N1797, N1520);
nor NOR4 (N1800, N1798, N40, N920, N1290);
or OR4 (N1801, N1773, N392, N613, N841);
xor XOR2 (N1802, N1779, N1678);
or OR4 (N1803, N1792, N968, N1089, N1555);
nand NAND4 (N1804, N1796, N551, N767, N737);
xor XOR2 (N1805, N1804, N1173);
and AND4 (N1806, N1794, N1647, N868, N74);
nand NAND2 (N1807, N1806, N735);
nand NAND3 (N1808, N1793, N1453, N1647);
or OR3 (N1809, N1799, N899, N349);
buf BUF1 (N1810, N1801);
not NOT1 (N1811, N1810);
or OR2 (N1812, N1809, N963);
and AND4 (N1813, N1805, N1016, N1625, N273);
buf BUF1 (N1814, N1803);
or OR3 (N1815, N1814, N518, N357);
xor XOR2 (N1816, N1791, N522);
and AND4 (N1817, N1784, N678, N424, N1000);
nor NOR3 (N1818, N1811, N158, N378);
nor NOR2 (N1819, N1802, N1026);
nor NOR2 (N1820, N1818, N382);
nand NAND2 (N1821, N1816, N1320);
nor NOR3 (N1822, N1820, N236, N246);
not NOT1 (N1823, N1815);
nand NAND2 (N1824, N1819, N1615);
and AND2 (N1825, N1822, N259);
and AND4 (N1826, N1817, N1141, N381, N718);
not NOT1 (N1827, N1813);
nand NAND2 (N1828, N1826, N407);
or OR2 (N1829, N1808, N159);
or OR4 (N1830, N1800, N1001, N318, N211);
nand NAND2 (N1831, N1821, N140);
buf BUF1 (N1832, N1827);
xor XOR2 (N1833, N1828, N404);
or OR3 (N1834, N1807, N478, N1366);
nand NAND3 (N1835, N1834, N1185, N1673);
not NOT1 (N1836, N1831);
xor XOR2 (N1837, N1829, N1250);
xor XOR2 (N1838, N1833, N15);
nand NAND4 (N1839, N1823, N1633, N177, N522);
buf BUF1 (N1840, N1837);
xor XOR2 (N1841, N1825, N1806);
xor XOR2 (N1842, N1832, N1447);
not NOT1 (N1843, N1824);
not NOT1 (N1844, N1839);
or OR3 (N1845, N1836, N1519, N1333);
nand NAND3 (N1846, N1812, N1315, N1004);
xor XOR2 (N1847, N1838, N847);
not NOT1 (N1848, N1847);
buf BUF1 (N1849, N1846);
nand NAND2 (N1850, N1848, N790);
or OR3 (N1851, N1830, N298, N53);
buf BUF1 (N1852, N1842);
and AND4 (N1853, N1845, N1692, N1668, N1254);
or OR2 (N1854, N1843, N1646);
buf BUF1 (N1855, N1840);
buf BUF1 (N1856, N1835);
nand NAND2 (N1857, N1844, N1103);
xor XOR2 (N1858, N1851, N757);
nand NAND3 (N1859, N1856, N1820, N1454);
not NOT1 (N1860, N1849);
nand NAND2 (N1861, N1860, N660);
buf BUF1 (N1862, N1841);
not NOT1 (N1863, N1852);
nor NOR4 (N1864, N1854, N1664, N306, N715);
not NOT1 (N1865, N1857);
or OR2 (N1866, N1861, N417);
xor XOR2 (N1867, N1863, N1330);
or OR3 (N1868, N1859, N320, N1698);
and AND3 (N1869, N1850, N609, N420);
buf BUF1 (N1870, N1864);
buf BUF1 (N1871, N1858);
not NOT1 (N1872, N1870);
nand NAND2 (N1873, N1865, N643);
nand NAND3 (N1874, N1855, N1238, N1046);
xor XOR2 (N1875, N1872, N1615);
or OR3 (N1876, N1869, N615, N253);
xor XOR2 (N1877, N1867, N316);
buf BUF1 (N1878, N1868);
buf BUF1 (N1879, N1876);
xor XOR2 (N1880, N1878, N785);
not NOT1 (N1881, N1879);
buf BUF1 (N1882, N1873);
xor XOR2 (N1883, N1880, N1823);
and AND2 (N1884, N1881, N1673);
not NOT1 (N1885, N1884);
xor XOR2 (N1886, N1875, N419);
nand NAND2 (N1887, N1883, N1533);
nor NOR4 (N1888, N1862, N1009, N1164, N1491);
xor XOR2 (N1889, N1882, N236);
buf BUF1 (N1890, N1887);
nand NAND4 (N1891, N1874, N648, N1198, N1468);
nor NOR3 (N1892, N1886, N370, N622);
nand NAND2 (N1893, N1866, N1749);
xor XOR2 (N1894, N1891, N502);
nand NAND3 (N1895, N1892, N174, N1267);
buf BUF1 (N1896, N1885);
nand NAND3 (N1897, N1896, N152, N1151);
xor XOR2 (N1898, N1871, N728);
nor NOR4 (N1899, N1877, N83, N1370, N742);
not NOT1 (N1900, N1895);
not NOT1 (N1901, N1853);
nand NAND3 (N1902, N1898, N1124, N1703);
nand NAND3 (N1903, N1890, N1393, N2);
xor XOR2 (N1904, N1888, N14);
not NOT1 (N1905, N1902);
nor NOR2 (N1906, N1903, N1211);
buf BUF1 (N1907, N1905);
buf BUF1 (N1908, N1899);
nand NAND3 (N1909, N1897, N1715, N1133);
buf BUF1 (N1910, N1904);
nand NAND2 (N1911, N1889, N670);
or OR4 (N1912, N1908, N1197, N1020, N1498);
or OR2 (N1913, N1912, N1523);
buf BUF1 (N1914, N1909);
not NOT1 (N1915, N1911);
or OR4 (N1916, N1894, N1288, N1031, N155);
buf BUF1 (N1917, N1915);
and AND3 (N1918, N1914, N251, N85);
nand NAND2 (N1919, N1907, N1866);
xor XOR2 (N1920, N1893, N1502);
or OR3 (N1921, N1916, N26, N880);
nand NAND2 (N1922, N1919, N200);
xor XOR2 (N1923, N1910, N587);
or OR2 (N1924, N1906, N1332);
nand NAND4 (N1925, N1920, N1360, N649, N1315);
nand NAND4 (N1926, N1900, N834, N489, N100);
nor NOR3 (N1927, N1924, N315, N1531);
nor NOR2 (N1928, N1925, N1223);
buf BUF1 (N1929, N1926);
buf BUF1 (N1930, N1922);
nand NAND4 (N1931, N1929, N44, N124, N116);
buf BUF1 (N1932, N1918);
and AND2 (N1933, N1913, N249);
and AND2 (N1934, N1930, N1834);
buf BUF1 (N1935, N1932);
nand NAND3 (N1936, N1927, N631, N935);
xor XOR2 (N1937, N1935, N1509);
or OR3 (N1938, N1931, N1592, N650);
nand NAND2 (N1939, N1917, N421);
or OR4 (N1940, N1934, N1140, N1644, N1727);
nor NOR4 (N1941, N1939, N987, N1097, N308);
xor XOR2 (N1942, N1933, N1801);
xor XOR2 (N1943, N1921, N204);
or OR4 (N1944, N1901, N352, N914, N408);
or OR3 (N1945, N1938, N186, N278);
nand NAND2 (N1946, N1940, N1234);
xor XOR2 (N1947, N1923, N1553);
and AND4 (N1948, N1945, N21, N378, N1531);
not NOT1 (N1949, N1936);
nand NAND2 (N1950, N1942, N1866);
buf BUF1 (N1951, N1946);
not NOT1 (N1952, N1943);
not NOT1 (N1953, N1947);
not NOT1 (N1954, N1952);
nor NOR3 (N1955, N1949, N266, N102);
buf BUF1 (N1956, N1944);
nand NAND3 (N1957, N1928, N105, N1168);
buf BUF1 (N1958, N1950);
buf BUF1 (N1959, N1953);
nand NAND4 (N1960, N1954, N956, N895, N46);
nand NAND3 (N1961, N1955, N1663, N884);
nand NAND2 (N1962, N1961, N959);
or OR2 (N1963, N1951, N1650);
buf BUF1 (N1964, N1963);
not NOT1 (N1965, N1937);
or OR3 (N1966, N1958, N521, N1787);
and AND2 (N1967, N1962, N263);
nor NOR3 (N1968, N1956, N1842, N249);
or OR3 (N1969, N1967, N1013, N1020);
not NOT1 (N1970, N1948);
xor XOR2 (N1971, N1966, N1021);
not NOT1 (N1972, N1957);
and AND4 (N1973, N1941, N1711, N1167, N799);
nor NOR2 (N1974, N1973, N143);
not NOT1 (N1975, N1970);
nor NOR3 (N1976, N1969, N638, N1449);
and AND3 (N1977, N1972, N1450, N1882);
and AND3 (N1978, N1964, N1015, N1544);
or OR3 (N1979, N1965, N1603, N291);
nor NOR3 (N1980, N1978, N628, N1697);
and AND3 (N1981, N1968, N1440, N979);
or OR3 (N1982, N1979, N694, N1161);
buf BUF1 (N1983, N1980);
or OR4 (N1984, N1983, N1278, N900, N1484);
buf BUF1 (N1985, N1982);
not NOT1 (N1986, N1971);
nand NAND4 (N1987, N1960, N474, N700, N34);
and AND2 (N1988, N1984, N800);
nor NOR4 (N1989, N1987, N126, N1142, N1897);
nand NAND2 (N1990, N1977, N141);
nand NAND2 (N1991, N1989, N1685);
nand NAND4 (N1992, N1959, N1464, N1769, N485);
xor XOR2 (N1993, N1991, N169);
buf BUF1 (N1994, N1981);
and AND4 (N1995, N1993, N1092, N84, N106);
buf BUF1 (N1996, N1992);
nor NOR2 (N1997, N1975, N1339);
xor XOR2 (N1998, N1990, N1133);
nor NOR2 (N1999, N1998, N954);
xor XOR2 (N2000, N1999, N274);
nand NAND2 (N2001, N2000, N1776);
or OR3 (N2002, N1986, N1705, N562);
nor NOR3 (N2003, N1997, N141, N12);
and AND4 (N2004, N1976, N1322, N504, N988);
nand NAND2 (N2005, N2003, N1710);
and AND3 (N2006, N1996, N1649, N328);
not NOT1 (N2007, N2004);
or OR3 (N2008, N2001, N1700, N159);
buf BUF1 (N2009, N2007);
and AND4 (N2010, N2008, N715, N1944, N339);
buf BUF1 (N2011, N1988);
and AND2 (N2012, N1974, N1522);
nand NAND2 (N2013, N2011, N1972);
nand NAND3 (N2014, N2012, N1420, N46);
and AND2 (N2015, N1995, N732);
xor XOR2 (N2016, N2005, N1047);
and AND2 (N2017, N2016, N419);
not NOT1 (N2018, N2009);
xor XOR2 (N2019, N2010, N534);
or OR3 (N2020, N1985, N608, N704);
not NOT1 (N2021, N2006);
xor XOR2 (N2022, N2018, N415);
nor NOR2 (N2023, N2017, N802);
xor XOR2 (N2024, N2002, N184);
buf BUF1 (N2025, N2022);
nand NAND2 (N2026, N2015, N1633);
or OR2 (N2027, N2020, N1256);
nor NOR3 (N2028, N2026, N1007, N844);
or OR3 (N2029, N2025, N908, N1270);
xor XOR2 (N2030, N2013, N38);
nor NOR3 (N2031, N2030, N1434, N565);
nor NOR2 (N2032, N2028, N1452);
xor XOR2 (N2033, N2014, N913);
not NOT1 (N2034, N2023);
nor NOR3 (N2035, N2019, N932, N1976);
or OR4 (N2036, N2029, N1813, N506, N1439);
and AND3 (N2037, N2021, N286, N1626);
not NOT1 (N2038, N2035);
buf BUF1 (N2039, N2038);
buf BUF1 (N2040, N2027);
not NOT1 (N2041, N1994);
buf BUF1 (N2042, N2031);
nand NAND4 (N2043, N2039, N1403, N1895, N1352);
nor NOR3 (N2044, N2024, N1892, N1172);
and AND3 (N2045, N2042, N1069, N1903);
not NOT1 (N2046, N2043);
not NOT1 (N2047, N2036);
xor XOR2 (N2048, N2040, N489);
nand NAND3 (N2049, N2032, N1149, N635);
xor XOR2 (N2050, N2048, N518);
xor XOR2 (N2051, N2044, N1698);
buf BUF1 (N2052, N2033);
not NOT1 (N2053, N2046);
buf BUF1 (N2054, N2053);
nand NAND2 (N2055, N2052, N1079);
xor XOR2 (N2056, N2047, N1557);
not NOT1 (N2057, N2049);
or OR3 (N2058, N2050, N498, N2021);
or OR3 (N2059, N2056, N1564, N887);
buf BUF1 (N2060, N2045);
nand NAND3 (N2061, N2055, N66, N1093);
nor NOR4 (N2062, N2034, N1354, N281, N1744);
nor NOR4 (N2063, N2061, N823, N1741, N493);
not NOT1 (N2064, N2063);
and AND3 (N2065, N2058, N804, N619);
not NOT1 (N2066, N2041);
nor NOR3 (N2067, N2054, N659, N1172);
xor XOR2 (N2068, N2051, N360);
xor XOR2 (N2069, N2060, N755);
not NOT1 (N2070, N2065);
xor XOR2 (N2071, N2062, N899);
buf BUF1 (N2072, N2037);
nor NOR4 (N2073, N2069, N368, N236, N1695);
and AND4 (N2074, N2072, N937, N1994, N879);
or OR3 (N2075, N2071, N177, N347);
not NOT1 (N2076, N2068);
buf BUF1 (N2077, N2076);
not NOT1 (N2078, N2074);
nor NOR4 (N2079, N2077, N600, N728, N1724);
buf BUF1 (N2080, N2064);
nand NAND3 (N2081, N2079, N1936, N371);
not NOT1 (N2082, N2067);
buf BUF1 (N2083, N2080);
nand NAND2 (N2084, N2059, N1025);
buf BUF1 (N2085, N2073);
not NOT1 (N2086, N2070);
xor XOR2 (N2087, N2085, N1681);
and AND3 (N2088, N2086, N1166, N571);
or OR2 (N2089, N2057, N665);
or OR2 (N2090, N2081, N142);
and AND4 (N2091, N2066, N1140, N1705, N926);
buf BUF1 (N2092, N2078);
xor XOR2 (N2093, N2092, N143);
or OR4 (N2094, N2083, N426, N450, N1085);
or OR3 (N2095, N2089, N185, N1418);
buf BUF1 (N2096, N2090);
nand NAND4 (N2097, N2096, N816, N1244, N1478);
nand NAND2 (N2098, N2091, N312);
nand NAND3 (N2099, N2098, N472, N1058);
nand NAND4 (N2100, N2099, N2002, N2054, N725);
and AND2 (N2101, N2095, N741);
xor XOR2 (N2102, N2094, N653);
and AND3 (N2103, N2087, N67, N773);
not NOT1 (N2104, N2082);
nand NAND3 (N2105, N2084, N1854, N746);
nand NAND3 (N2106, N2103, N1719, N2023);
or OR3 (N2107, N2075, N1502, N42);
and AND3 (N2108, N2101, N943, N725);
not NOT1 (N2109, N2100);
buf BUF1 (N2110, N2088);
and AND4 (N2111, N2106, N1574, N857, N1542);
not NOT1 (N2112, N2108);
or OR2 (N2113, N2105, N1955);
buf BUF1 (N2114, N2097);
nand NAND4 (N2115, N2112, N498, N1778, N1795);
nor NOR2 (N2116, N2107, N806);
and AND2 (N2117, N2111, N1602);
not NOT1 (N2118, N2114);
xor XOR2 (N2119, N2118, N125);
or OR2 (N2120, N2102, N1432);
buf BUF1 (N2121, N2119);
buf BUF1 (N2122, N2109);
and AND2 (N2123, N2122, N665);
nand NAND4 (N2124, N2113, N1482, N126, N189);
not NOT1 (N2125, N2120);
not NOT1 (N2126, N2123);
buf BUF1 (N2127, N2121);
nor NOR3 (N2128, N2115, N1411, N1293);
nand NAND4 (N2129, N2126, N869, N766, N963);
and AND4 (N2130, N2104, N1719, N1512, N163);
xor XOR2 (N2131, N2110, N415);
and AND2 (N2132, N2124, N1350);
and AND3 (N2133, N2125, N1261, N984);
nor NOR4 (N2134, N2130, N1155, N1077, N1249);
nor NOR3 (N2135, N2132, N1880, N1578);
not NOT1 (N2136, N2116);
buf BUF1 (N2137, N2134);
xor XOR2 (N2138, N2137, N328);
nor NOR2 (N2139, N2128, N2008);
and AND3 (N2140, N2138, N1378, N1615);
and AND2 (N2141, N2136, N1975);
and AND4 (N2142, N2141, N24, N1820, N1826);
or OR2 (N2143, N2140, N1524);
or OR4 (N2144, N2127, N1281, N1882, N1784);
nor NOR4 (N2145, N2139, N1101, N2037, N1497);
not NOT1 (N2146, N2143);
nor NOR2 (N2147, N2135, N1158);
buf BUF1 (N2148, N2133);
nand NAND4 (N2149, N2117, N195, N1684, N571);
and AND4 (N2150, N2144, N1602, N1591, N612);
nor NOR3 (N2151, N2131, N2134, N147);
or OR4 (N2152, N2142, N637, N1968, N286);
and AND2 (N2153, N2148, N1161);
nand NAND2 (N2154, N2146, N2045);
buf BUF1 (N2155, N2129);
nand NAND4 (N2156, N2152, N2058, N412, N1926);
nor NOR3 (N2157, N2156, N236, N134);
or OR2 (N2158, N2145, N1798);
nor NOR4 (N2159, N2153, N775, N303, N1032);
nand NAND2 (N2160, N2154, N1769);
not NOT1 (N2161, N2147);
nand NAND4 (N2162, N2151, N1991, N1924, N1023);
and AND4 (N2163, N2150, N1263, N1110, N496);
buf BUF1 (N2164, N2163);
buf BUF1 (N2165, N2162);
xor XOR2 (N2166, N2157, N477);
and AND4 (N2167, N2161, N681, N680, N71);
and AND4 (N2168, N2167, N996, N740, N1286);
or OR2 (N2169, N2166, N352);
not NOT1 (N2170, N2164);
and AND2 (N2171, N2160, N295);
and AND3 (N2172, N2170, N142, N991);
xor XOR2 (N2173, N2165, N1345);
xor XOR2 (N2174, N2173, N733);
nor NOR4 (N2175, N2172, N1487, N861, N769);
or OR3 (N2176, N2174, N1279, N222);
nor NOR2 (N2177, N2158, N1998);
buf BUF1 (N2178, N2169);
or OR4 (N2179, N2155, N1346, N1965, N777);
not NOT1 (N2180, N2177);
nor NOR3 (N2181, N2175, N260, N231);
nand NAND2 (N2182, N2181, N1488);
buf BUF1 (N2183, N2149);
buf BUF1 (N2184, N2180);
not NOT1 (N2185, N2168);
not NOT1 (N2186, N2182);
or OR3 (N2187, N2183, N2172, N591);
not NOT1 (N2188, N2186);
nor NOR2 (N2189, N2179, N30);
xor XOR2 (N2190, N2176, N1016);
xor XOR2 (N2191, N2159, N1385);
or OR3 (N2192, N2093, N1883, N2013);
xor XOR2 (N2193, N2188, N1935);
buf BUF1 (N2194, N2190);
nand NAND3 (N2195, N2171, N693, N1822);
xor XOR2 (N2196, N2194, N2161);
nand NAND4 (N2197, N2184, N2073, N990, N1047);
or OR4 (N2198, N2195, N404, N507, N1188);
nand NAND3 (N2199, N2185, N1200, N559);
nand NAND3 (N2200, N2197, N1598, N100);
nor NOR3 (N2201, N2178, N2179, N1132);
xor XOR2 (N2202, N2199, N1717);
xor XOR2 (N2203, N2196, N1726);
buf BUF1 (N2204, N2191);
nand NAND4 (N2205, N2193, N801, N37, N900);
buf BUF1 (N2206, N2205);
or OR4 (N2207, N2203, N1649, N1532, N1973);
nor NOR2 (N2208, N2189, N742);
nand NAND2 (N2209, N2206, N1262);
nand NAND2 (N2210, N2198, N596);
nand NAND4 (N2211, N2209, N1104, N657, N144);
xor XOR2 (N2212, N2201, N1385);
not NOT1 (N2213, N2187);
buf BUF1 (N2214, N2202);
and AND3 (N2215, N2200, N2096, N1038);
not NOT1 (N2216, N2214);
not NOT1 (N2217, N2210);
nand NAND4 (N2218, N2217, N1279, N1307, N878);
nand NAND3 (N2219, N2213, N31, N972);
nor NOR4 (N2220, N2215, N1180, N1003, N1619);
xor XOR2 (N2221, N2207, N336);
nor NOR3 (N2222, N2218, N871, N851);
or OR4 (N2223, N2219, N588, N391, N849);
xor XOR2 (N2224, N2211, N1280);
and AND3 (N2225, N2221, N1246, N545);
and AND3 (N2226, N2220, N288, N1950);
nand NAND3 (N2227, N2225, N1652, N147);
not NOT1 (N2228, N2224);
buf BUF1 (N2229, N2222);
not NOT1 (N2230, N2228);
nand NAND2 (N2231, N2223, N143);
and AND2 (N2232, N2192, N1906);
nand NAND4 (N2233, N2232, N632, N824, N1641);
xor XOR2 (N2234, N2226, N917);
or OR2 (N2235, N2229, N2087);
not NOT1 (N2236, N2216);
or OR3 (N2237, N2204, N203, N738);
and AND4 (N2238, N2237, N864, N1568, N881);
xor XOR2 (N2239, N2238, N1814);
nand NAND4 (N2240, N2208, N2085, N1635, N937);
and AND2 (N2241, N2231, N74);
or OR3 (N2242, N2240, N2173, N78);
nand NAND2 (N2243, N2242, N442);
and AND2 (N2244, N2233, N434);
not NOT1 (N2245, N2243);
xor XOR2 (N2246, N2236, N854);
and AND3 (N2247, N2227, N1686, N443);
xor XOR2 (N2248, N2239, N306);
or OR3 (N2249, N2234, N1547, N1285);
not NOT1 (N2250, N2212);
or OR4 (N2251, N2245, N1303, N1480, N1522);
nand NAND3 (N2252, N2247, N419, N297);
nor NOR2 (N2253, N2241, N701);
or OR4 (N2254, N2230, N310, N1564, N811);
xor XOR2 (N2255, N2250, N1527);
buf BUF1 (N2256, N2244);
buf BUF1 (N2257, N2235);
or OR2 (N2258, N2254, N798);
and AND4 (N2259, N2257, N195, N1764, N2028);
nor NOR3 (N2260, N2255, N1767, N1312);
and AND4 (N2261, N2259, N340, N605, N1503);
buf BUF1 (N2262, N2253);
or OR2 (N2263, N2256, N1876);
nor NOR4 (N2264, N2249, N2127, N1800, N1123);
xor XOR2 (N2265, N2263, N795);
nand NAND3 (N2266, N2261, N736, N371);
and AND3 (N2267, N2258, N1826, N1767);
and AND3 (N2268, N2246, N1820, N2194);
and AND4 (N2269, N2268, N2160, N132, N1401);
nand NAND3 (N2270, N2252, N2174, N1328);
nor NOR4 (N2271, N2269, N31, N2193, N280);
and AND2 (N2272, N2264, N524);
nor NOR2 (N2273, N2270, N1080);
or OR4 (N2274, N2262, N1973, N1484, N731);
or OR3 (N2275, N2274, N1103, N1999);
or OR4 (N2276, N2265, N1686, N1075, N1752);
or OR3 (N2277, N2273, N231, N394);
and AND2 (N2278, N2272, N1938);
xor XOR2 (N2279, N2276, N767);
or OR4 (N2280, N2275, N882, N1012, N1961);
nor NOR3 (N2281, N2279, N992, N1597);
or OR3 (N2282, N2280, N881, N1392);
or OR3 (N2283, N2248, N1063, N223);
or OR3 (N2284, N2260, N540, N2161);
or OR2 (N2285, N2271, N1322);
xor XOR2 (N2286, N2267, N1861);
nor NOR4 (N2287, N2283, N1971, N1233, N415);
buf BUF1 (N2288, N2282);
and AND3 (N2289, N2284, N1906, N1195);
nand NAND4 (N2290, N2285, N1145, N1768, N1152);
nand NAND4 (N2291, N2266, N665, N725, N1167);
xor XOR2 (N2292, N2281, N130);
buf BUF1 (N2293, N2292);
nor NOR3 (N2294, N2288, N1052, N891);
nor NOR4 (N2295, N2291, N1130, N389, N262);
not NOT1 (N2296, N2295);
nand NAND3 (N2297, N2294, N1937, N1468);
nor NOR2 (N2298, N2297, N1743);
not NOT1 (N2299, N2296);
xor XOR2 (N2300, N2251, N2267);
nand NAND3 (N2301, N2298, N467, N1055);
xor XOR2 (N2302, N2278, N1857);
and AND2 (N2303, N2277, N33);
or OR4 (N2304, N2300, N1716, N1058, N1082);
nand NAND4 (N2305, N2289, N248, N2244, N2088);
nor NOR2 (N2306, N2303, N5);
nand NAND2 (N2307, N2301, N1537);
nand NAND4 (N2308, N2304, N2208, N173, N1120);
not NOT1 (N2309, N2305);
nor NOR2 (N2310, N2286, N437);
nor NOR2 (N2311, N2287, N1789);
not NOT1 (N2312, N2302);
or OR3 (N2313, N2308, N164, N1206);
nor NOR4 (N2314, N2306, N1236, N1729, N1073);
nor NOR3 (N2315, N2312, N1296, N166);
nor NOR4 (N2316, N2314, N657, N929, N312);
xor XOR2 (N2317, N2293, N1600);
or OR2 (N2318, N2290, N1768);
nor NOR2 (N2319, N2316, N1576);
and AND4 (N2320, N2310, N2128, N228, N1773);
nand NAND3 (N2321, N2319, N12, N1772);
buf BUF1 (N2322, N2320);
not NOT1 (N2323, N2299);
and AND2 (N2324, N2315, N668);
nor NOR4 (N2325, N2318, N1209, N1236, N1940);
nor NOR2 (N2326, N2311, N2271);
buf BUF1 (N2327, N2324);
xor XOR2 (N2328, N2313, N587);
nand NAND4 (N2329, N2317, N904, N97, N2146);
nand NAND4 (N2330, N2323, N42, N861, N1904);
not NOT1 (N2331, N2330);
nor NOR4 (N2332, N2325, N1726, N517, N1082);
nor NOR4 (N2333, N2332, N1519, N1768, N1881);
buf BUF1 (N2334, N2329);
buf BUF1 (N2335, N2328);
not NOT1 (N2336, N2326);
buf BUF1 (N2337, N2309);
and AND3 (N2338, N2322, N254, N2081);
nand NAND2 (N2339, N2327, N161);
buf BUF1 (N2340, N2337);
not NOT1 (N2341, N2336);
nand NAND4 (N2342, N2334, N882, N2110, N13);
xor XOR2 (N2343, N2321, N1511);
not NOT1 (N2344, N2342);
not NOT1 (N2345, N2343);
or OR4 (N2346, N2331, N1102, N22, N2034);
or OR4 (N2347, N2338, N2322, N1602, N375);
or OR2 (N2348, N2340, N2167);
buf BUF1 (N2349, N2339);
buf BUF1 (N2350, N2347);
xor XOR2 (N2351, N2345, N341);
xor XOR2 (N2352, N2344, N604);
nand NAND4 (N2353, N2346, N1285, N763, N1727);
not NOT1 (N2354, N2353);
nand NAND3 (N2355, N2348, N1828, N2184);
xor XOR2 (N2356, N2355, N1415);
or OR3 (N2357, N2356, N142, N2282);
xor XOR2 (N2358, N2351, N1062);
nand NAND4 (N2359, N2341, N1045, N808, N623);
xor XOR2 (N2360, N2352, N1908);
buf BUF1 (N2361, N2349);
buf BUF1 (N2362, N2357);
xor XOR2 (N2363, N2333, N1402);
buf BUF1 (N2364, N2362);
or OR3 (N2365, N2335, N1835, N574);
nor NOR3 (N2366, N2358, N176, N1121);
xor XOR2 (N2367, N2359, N1476);
xor XOR2 (N2368, N2361, N1943);
buf BUF1 (N2369, N2367);
xor XOR2 (N2370, N2350, N2156);
xor XOR2 (N2371, N2370, N1657);
not NOT1 (N2372, N2366);
nand NAND4 (N2373, N2363, N683, N722, N726);
not NOT1 (N2374, N2369);
and AND2 (N2375, N2372, N60);
buf BUF1 (N2376, N2364);
buf BUF1 (N2377, N2365);
buf BUF1 (N2378, N2368);
nand NAND4 (N2379, N2374, N1142, N1065, N1424);
not NOT1 (N2380, N2373);
and AND3 (N2381, N2376, N596, N781);
or OR3 (N2382, N2354, N600, N1045);
not NOT1 (N2383, N2379);
buf BUF1 (N2384, N2380);
buf BUF1 (N2385, N2378);
nand NAND3 (N2386, N2377, N94, N1090);
not NOT1 (N2387, N2375);
xor XOR2 (N2388, N2371, N261);
or OR2 (N2389, N2384, N2059);
or OR4 (N2390, N2307, N272, N496, N1229);
buf BUF1 (N2391, N2385);
xor XOR2 (N2392, N2387, N450);
and AND2 (N2393, N2383, N1891);
nor NOR3 (N2394, N2360, N196, N1622);
or OR2 (N2395, N2393, N841);
nor NOR4 (N2396, N2392, N490, N911, N1494);
nand NAND3 (N2397, N2381, N2165, N538);
nand NAND2 (N2398, N2388, N1674);
or OR3 (N2399, N2390, N1396, N2165);
nand NAND2 (N2400, N2389, N2156);
not NOT1 (N2401, N2396);
xor XOR2 (N2402, N2386, N1071);
buf BUF1 (N2403, N2391);
xor XOR2 (N2404, N2401, N124);
xor XOR2 (N2405, N2398, N2224);
nor NOR3 (N2406, N2405, N503, N876);
nand NAND4 (N2407, N2404, N1158, N2345, N524);
nor NOR3 (N2408, N2395, N1469, N1712);
nand NAND2 (N2409, N2394, N2324);
nand NAND3 (N2410, N2382, N65, N1546);
or OR2 (N2411, N2410, N668);
and AND3 (N2412, N2407, N113, N2279);
nor NOR2 (N2413, N2397, N1163);
not NOT1 (N2414, N2400);
nor NOR4 (N2415, N2403, N1441, N1761, N1833);
buf BUF1 (N2416, N2414);
or OR2 (N2417, N2412, N86);
or OR3 (N2418, N2415, N1251, N1570);
and AND3 (N2419, N2408, N769, N832);
not NOT1 (N2420, N2399);
buf BUF1 (N2421, N2409);
nand NAND3 (N2422, N2421, N2245, N33);
not NOT1 (N2423, N2418);
or OR4 (N2424, N2420, N632, N2283, N112);
or OR3 (N2425, N2422, N565, N2197);
nand NAND4 (N2426, N2419, N1592, N1806, N1679);
not NOT1 (N2427, N2425);
nor NOR2 (N2428, N2427, N1501);
nor NOR2 (N2429, N2406, N62);
nor NOR4 (N2430, N2416, N2058, N2339, N1773);
buf BUF1 (N2431, N2423);
or OR4 (N2432, N2429, N973, N96, N1793);
or OR3 (N2433, N2411, N2152, N1591);
or OR4 (N2434, N2417, N1231, N2201, N1112);
not NOT1 (N2435, N2402);
nor NOR2 (N2436, N2413, N51);
xor XOR2 (N2437, N2426, N213);
xor XOR2 (N2438, N2436, N936);
buf BUF1 (N2439, N2431);
xor XOR2 (N2440, N2433, N1701);
nand NAND4 (N2441, N2438, N1369, N952, N1313);
buf BUF1 (N2442, N2437);
not NOT1 (N2443, N2442);
and AND4 (N2444, N2424, N526, N868, N2013);
nor NOR4 (N2445, N2443, N1935, N1280, N1795);
nor NOR3 (N2446, N2428, N1515, N711);
nor NOR2 (N2447, N2435, N2085);
and AND4 (N2448, N2434, N1819, N1039, N2305);
or OR3 (N2449, N2445, N1736, N2331);
not NOT1 (N2450, N2446);
xor XOR2 (N2451, N2430, N152);
buf BUF1 (N2452, N2440);
buf BUF1 (N2453, N2444);
nand NAND4 (N2454, N2451, N187, N2208, N813);
not NOT1 (N2455, N2432);
nand NAND4 (N2456, N2450, N791, N1800, N762);
or OR2 (N2457, N2454, N2322);
and AND3 (N2458, N2456, N962, N1374);
or OR2 (N2459, N2452, N464);
buf BUF1 (N2460, N2448);
and AND2 (N2461, N2458, N2407);
and AND2 (N2462, N2441, N698);
nor NOR2 (N2463, N2461, N2016);
not NOT1 (N2464, N2463);
not NOT1 (N2465, N2459);
buf BUF1 (N2466, N2449);
nor NOR2 (N2467, N2464, N1358);
xor XOR2 (N2468, N2453, N1015);
nand NAND3 (N2469, N2457, N1871, N20);
nand NAND2 (N2470, N2465, N416);
and AND2 (N2471, N2466, N85);
and AND4 (N2472, N2447, N683, N1993, N220);
or OR2 (N2473, N2472, N568);
or OR4 (N2474, N2471, N332, N2035, N1548);
and AND4 (N2475, N2467, N2053, N220, N1958);
nor NOR2 (N2476, N2474, N1558);
xor XOR2 (N2477, N2455, N1477);
and AND3 (N2478, N2439, N1221, N893);
nor NOR4 (N2479, N2469, N1142, N2131, N1323);
and AND4 (N2480, N2468, N2033, N1351, N29);
xor XOR2 (N2481, N2462, N2284);
or OR4 (N2482, N2479, N1232, N230, N2476);
not NOT1 (N2483, N508);
and AND2 (N2484, N2470, N151);
xor XOR2 (N2485, N2473, N526);
or OR2 (N2486, N2475, N2456);
not NOT1 (N2487, N2477);
nand NAND2 (N2488, N2487, N1581);
xor XOR2 (N2489, N2480, N755);
or OR3 (N2490, N2483, N1994, N1345);
buf BUF1 (N2491, N2478);
nor NOR4 (N2492, N2460, N1148, N2209, N1346);
nand NAND2 (N2493, N2491, N1789);
and AND4 (N2494, N2485, N1289, N726, N1624);
and AND2 (N2495, N2494, N2090);
or OR4 (N2496, N2493, N2440, N396, N1688);
nor NOR4 (N2497, N2482, N251, N1998, N2437);
buf BUF1 (N2498, N2490);
not NOT1 (N2499, N2492);
buf BUF1 (N2500, N2486);
nor NOR2 (N2501, N2481, N427);
and AND3 (N2502, N2500, N386, N444);
xor XOR2 (N2503, N2484, N224);
or OR4 (N2504, N2497, N1618, N1839, N2343);
not NOT1 (N2505, N2501);
nand NAND2 (N2506, N2498, N455);
not NOT1 (N2507, N2506);
and AND3 (N2508, N2504, N2342, N507);
nand NAND4 (N2509, N2499, N1170, N1362, N529);
and AND3 (N2510, N2507, N797, N2420);
and AND3 (N2511, N2502, N1693, N1085);
nor NOR4 (N2512, N2495, N2434, N375, N2429);
xor XOR2 (N2513, N2511, N2380);
xor XOR2 (N2514, N2509, N379);
not NOT1 (N2515, N2508);
buf BUF1 (N2516, N2496);
nand NAND3 (N2517, N2489, N1769, N2158);
nand NAND2 (N2518, N2488, N1006);
not NOT1 (N2519, N2512);
and AND4 (N2520, N2503, N1789, N859, N590);
xor XOR2 (N2521, N2510, N2168);
nor NOR4 (N2522, N2520, N1815, N599, N1263);
not NOT1 (N2523, N2513);
buf BUF1 (N2524, N2522);
and AND4 (N2525, N2505, N1363, N2317, N2430);
nor NOR4 (N2526, N2514, N1386, N1349, N1042);
nor NOR3 (N2527, N2523, N1687, N994);
xor XOR2 (N2528, N2521, N455);
xor XOR2 (N2529, N2526, N220);
buf BUF1 (N2530, N2516);
not NOT1 (N2531, N2527);
xor XOR2 (N2532, N2518, N941);
nand NAND3 (N2533, N2525, N2273, N66);
xor XOR2 (N2534, N2519, N1212);
not NOT1 (N2535, N2531);
and AND2 (N2536, N2515, N1351);
or OR2 (N2537, N2534, N502);
not NOT1 (N2538, N2532);
not NOT1 (N2539, N2517);
nand NAND4 (N2540, N2530, N1613, N627, N1493);
buf BUF1 (N2541, N2540);
buf BUF1 (N2542, N2536);
not NOT1 (N2543, N2541);
buf BUF1 (N2544, N2528);
or OR4 (N2545, N2533, N2399, N35, N2143);
or OR3 (N2546, N2524, N952, N1728);
nand NAND3 (N2547, N2538, N631, N1961);
and AND2 (N2548, N2546, N1755);
and AND3 (N2549, N2542, N2335, N2211);
xor XOR2 (N2550, N2545, N693);
not NOT1 (N2551, N2529);
and AND4 (N2552, N2539, N2103, N1199, N1985);
nand NAND3 (N2553, N2552, N899, N915);
buf BUF1 (N2554, N2551);
xor XOR2 (N2555, N2549, N722);
buf BUF1 (N2556, N2554);
not NOT1 (N2557, N2550);
and AND2 (N2558, N2543, N2134);
xor XOR2 (N2559, N2558, N1055);
or OR3 (N2560, N2535, N1224, N100);
nor NOR4 (N2561, N2553, N700, N138, N1725);
nand NAND4 (N2562, N2544, N22, N1153, N1898);
nand NAND3 (N2563, N2547, N1606, N1416);
xor XOR2 (N2564, N2562, N1898);
not NOT1 (N2565, N2563);
or OR3 (N2566, N2565, N476, N1319);
nor NOR2 (N2567, N2560, N1605);
or OR3 (N2568, N2556, N677, N250);
buf BUF1 (N2569, N2564);
nand NAND2 (N2570, N2568, N1921);
xor XOR2 (N2571, N2548, N585);
not NOT1 (N2572, N2566);
not NOT1 (N2573, N2571);
or OR2 (N2574, N2572, N1279);
not NOT1 (N2575, N2557);
and AND2 (N2576, N2574, N1558);
nand NAND3 (N2577, N2555, N12, N33);
buf BUF1 (N2578, N2561);
and AND4 (N2579, N2577, N2029, N1504, N1839);
and AND3 (N2580, N2567, N2561, N1963);
or OR2 (N2581, N2575, N964);
not NOT1 (N2582, N2580);
and AND2 (N2583, N2569, N973);
not NOT1 (N2584, N2570);
buf BUF1 (N2585, N2573);
and AND3 (N2586, N2583, N651, N2453);
xor XOR2 (N2587, N2559, N1113);
nand NAND3 (N2588, N2581, N577, N1659);
nor NOR3 (N2589, N2579, N1303, N862);
buf BUF1 (N2590, N2578);
buf BUF1 (N2591, N2582);
not NOT1 (N2592, N2585);
nand NAND2 (N2593, N2590, N1489);
xor XOR2 (N2594, N2537, N1282);
nor NOR2 (N2595, N2589, N1858);
nand NAND4 (N2596, N2594, N1684, N65, N2042);
not NOT1 (N2597, N2587);
or OR3 (N2598, N2595, N1253, N2092);
nor NOR3 (N2599, N2586, N1711, N1803);
nor NOR4 (N2600, N2596, N848, N1038, N208);
xor XOR2 (N2601, N2599, N1977);
nor NOR3 (N2602, N2600, N754, N441);
nor NOR2 (N2603, N2597, N772);
not NOT1 (N2604, N2602);
nand NAND4 (N2605, N2593, N1476, N1265, N2505);
not NOT1 (N2606, N2584);
or OR4 (N2607, N2598, N1442, N1710, N1565);
not NOT1 (N2608, N2603);
nor NOR2 (N2609, N2605, N1212);
not NOT1 (N2610, N2592);
and AND4 (N2611, N2609, N1235, N347, N1286);
buf BUF1 (N2612, N2610);
not NOT1 (N2613, N2611);
and AND4 (N2614, N2612, N2014, N592, N2351);
and AND4 (N2615, N2607, N1953, N746, N2335);
xor XOR2 (N2616, N2588, N1848);
and AND2 (N2617, N2613, N907);
and AND4 (N2618, N2606, N12, N1325, N1735);
xor XOR2 (N2619, N2616, N2423);
not NOT1 (N2620, N2614);
and AND4 (N2621, N2618, N2141, N1340, N2187);
not NOT1 (N2622, N2591);
nand NAND2 (N2623, N2617, N2065);
xor XOR2 (N2624, N2620, N18);
or OR4 (N2625, N2623, N1391, N785, N553);
nor NOR3 (N2626, N2619, N1205, N2138);
xor XOR2 (N2627, N2625, N1566);
nand NAND2 (N2628, N2627, N1436);
nand NAND4 (N2629, N2622, N678, N1188, N2002);
not NOT1 (N2630, N2628);
and AND3 (N2631, N2601, N752, N1038);
buf BUF1 (N2632, N2624);
not NOT1 (N2633, N2631);
xor XOR2 (N2634, N2604, N845);
xor XOR2 (N2635, N2608, N1859);
not NOT1 (N2636, N2629);
nand NAND4 (N2637, N2630, N1324, N1859, N1831);
buf BUF1 (N2638, N2633);
xor XOR2 (N2639, N2637, N1397);
nor NOR4 (N2640, N2638, N2315, N1931, N1620);
or OR3 (N2641, N2632, N1597, N732);
buf BUF1 (N2642, N2640);
and AND3 (N2643, N2635, N1264, N1181);
buf BUF1 (N2644, N2621);
and AND2 (N2645, N2636, N1802);
buf BUF1 (N2646, N2634);
and AND4 (N2647, N2644, N1819, N1485, N695);
nand NAND3 (N2648, N2615, N2317, N1736);
or OR3 (N2649, N2645, N380, N922);
nor NOR2 (N2650, N2643, N2526);
nand NAND2 (N2651, N2641, N1885);
not NOT1 (N2652, N2639);
xor XOR2 (N2653, N2576, N831);
or OR3 (N2654, N2652, N804, N1351);
or OR3 (N2655, N2642, N771, N2650);
or OR2 (N2656, N2394, N933);
or OR2 (N2657, N2649, N2083);
or OR3 (N2658, N2655, N1843, N1242);
not NOT1 (N2659, N2647);
or OR2 (N2660, N2659, N208);
buf BUF1 (N2661, N2651);
nand NAND4 (N2662, N2654, N2642, N1004, N1601);
nor NOR3 (N2663, N2657, N410, N2387);
nand NAND3 (N2664, N2662, N1643, N212);
or OR2 (N2665, N2646, N2414);
xor XOR2 (N2666, N2663, N1616);
not NOT1 (N2667, N2665);
buf BUF1 (N2668, N2667);
buf BUF1 (N2669, N2656);
buf BUF1 (N2670, N2653);
xor XOR2 (N2671, N2660, N1361);
xor XOR2 (N2672, N2670, N1323);
and AND3 (N2673, N2666, N2531, N729);
buf BUF1 (N2674, N2673);
nand NAND2 (N2675, N2626, N1208);
xor XOR2 (N2676, N2664, N834);
nor NOR4 (N2677, N2675, N200, N1250, N434);
and AND2 (N2678, N2658, N53);
not NOT1 (N2679, N2648);
nand NAND4 (N2680, N2669, N2621, N99, N1456);
or OR3 (N2681, N2668, N1493, N87);
buf BUF1 (N2682, N2680);
nand NAND4 (N2683, N2672, N1353, N1482, N2561);
buf BUF1 (N2684, N2674);
or OR4 (N2685, N2683, N325, N1631, N949);
nor NOR2 (N2686, N2679, N439);
and AND2 (N2687, N2681, N683);
nor NOR2 (N2688, N2671, N773);
not NOT1 (N2689, N2685);
nor NOR3 (N2690, N2661, N2538, N845);
not NOT1 (N2691, N2684);
buf BUF1 (N2692, N2676);
xor XOR2 (N2693, N2687, N676);
xor XOR2 (N2694, N2688, N2293);
nor NOR2 (N2695, N2693, N1727);
and AND4 (N2696, N2692, N1613, N1102, N1629);
or OR4 (N2697, N2690, N1226, N2225, N1059);
not NOT1 (N2698, N2694);
and AND4 (N2699, N2677, N2687, N1336, N1405);
buf BUF1 (N2700, N2696);
buf BUF1 (N2701, N2686);
nor NOR2 (N2702, N2682, N162);
not NOT1 (N2703, N2697);
not NOT1 (N2704, N2698);
not NOT1 (N2705, N2689);
and AND2 (N2706, N2704, N344);
nor NOR4 (N2707, N2703, N1374, N1355, N661);
not NOT1 (N2708, N2700);
xor XOR2 (N2709, N2708, N753);
or OR3 (N2710, N2705, N837, N2662);
not NOT1 (N2711, N2699);
not NOT1 (N2712, N2702);
or OR3 (N2713, N2709, N2007, N360);
nand NAND3 (N2714, N2701, N1750, N62);
or OR2 (N2715, N2710, N579);
nand NAND3 (N2716, N2691, N1990, N664);
nor NOR3 (N2717, N2695, N476, N419);
buf BUF1 (N2718, N2716);
nor NOR4 (N2719, N2707, N1191, N1414, N1369);
nand NAND4 (N2720, N2714, N317, N2381, N2323);
nor NOR2 (N2721, N2718, N1801);
and AND2 (N2722, N2715, N73);
xor XOR2 (N2723, N2722, N955);
or OR3 (N2724, N2723, N1408, N2322);
xor XOR2 (N2725, N2719, N414);
nand NAND2 (N2726, N2725, N233);
or OR4 (N2727, N2712, N1264, N896, N1586);
not NOT1 (N2728, N2713);
xor XOR2 (N2729, N2720, N1020);
nor NOR3 (N2730, N2729, N1121, N799);
and AND3 (N2731, N2678, N2327, N758);
and AND3 (N2732, N2730, N2614, N644);
and AND4 (N2733, N2728, N836, N551, N2238);
or OR4 (N2734, N2717, N1735, N1699, N435);
xor XOR2 (N2735, N2733, N962);
buf BUF1 (N2736, N2727);
buf BUF1 (N2737, N2732);
buf BUF1 (N2738, N2734);
or OR3 (N2739, N2721, N2584, N2260);
and AND3 (N2740, N2739, N504, N1843);
xor XOR2 (N2741, N2731, N42);
buf BUF1 (N2742, N2741);
or OR4 (N2743, N2735, N220, N974, N2351);
or OR3 (N2744, N2740, N2717, N2352);
nor NOR3 (N2745, N2726, N56, N1070);
and AND3 (N2746, N2738, N1047, N2528);
nor NOR3 (N2747, N2711, N24, N2611);
not NOT1 (N2748, N2742);
nor NOR3 (N2749, N2744, N1633, N212);
nor NOR3 (N2750, N2706, N1936, N693);
xor XOR2 (N2751, N2736, N1557);
and AND3 (N2752, N2745, N2397, N2583);
buf BUF1 (N2753, N2737);
xor XOR2 (N2754, N2743, N375);
and AND3 (N2755, N2754, N1208, N2364);
nand NAND2 (N2756, N2752, N1273);
nor NOR2 (N2757, N2750, N2180);
or OR3 (N2758, N2747, N637, N1600);
buf BUF1 (N2759, N2753);
nor NOR4 (N2760, N2751, N536, N1629, N975);
and AND3 (N2761, N2758, N1100, N762);
and AND4 (N2762, N2755, N362, N928, N2727);
nand NAND4 (N2763, N2748, N1959, N1738, N540);
not NOT1 (N2764, N2757);
nand NAND4 (N2765, N2764, N1485, N2718, N1864);
nand NAND3 (N2766, N2765, N2460, N370);
not NOT1 (N2767, N2724);
not NOT1 (N2768, N2756);
nor NOR2 (N2769, N2749, N303);
nand NAND4 (N2770, N2768, N1891, N2648, N1804);
buf BUF1 (N2771, N2761);
not NOT1 (N2772, N2771);
and AND3 (N2773, N2762, N761, N2409);
buf BUF1 (N2774, N2772);
nand NAND2 (N2775, N2767, N899);
or OR4 (N2776, N2774, N1714, N1817, N2438);
and AND2 (N2777, N2746, N857);
xor XOR2 (N2778, N2766, N119);
buf BUF1 (N2779, N2759);
xor XOR2 (N2780, N2769, N2332);
buf BUF1 (N2781, N2773);
xor XOR2 (N2782, N2770, N1604);
and AND3 (N2783, N2777, N811, N377);
not NOT1 (N2784, N2775);
xor XOR2 (N2785, N2760, N1958);
nand NAND2 (N2786, N2783, N2492);
not NOT1 (N2787, N2785);
xor XOR2 (N2788, N2781, N2104);
nor NOR4 (N2789, N2763, N1285, N2290, N2717);
and AND4 (N2790, N2779, N992, N2671, N1771);
buf BUF1 (N2791, N2776);
not NOT1 (N2792, N2791);
and AND2 (N2793, N2792, N2015);
not NOT1 (N2794, N2784);
not NOT1 (N2795, N2793);
nor NOR4 (N2796, N2782, N1983, N2448, N2328);
nor NOR4 (N2797, N2796, N1538, N1747, N2173);
and AND2 (N2798, N2789, N2723);
nand NAND4 (N2799, N2795, N1720, N2506, N685);
not NOT1 (N2800, N2797);
not NOT1 (N2801, N2787);
buf BUF1 (N2802, N2788);
nand NAND4 (N2803, N2780, N1228, N1411, N2583);
and AND4 (N2804, N2800, N1035, N2385, N340);
buf BUF1 (N2805, N2798);
or OR4 (N2806, N2786, N2597, N668, N551);
or OR3 (N2807, N2794, N534, N1012);
nand NAND2 (N2808, N2803, N1826);
nand NAND2 (N2809, N2799, N697);
not NOT1 (N2810, N2806);
not NOT1 (N2811, N2778);
nor NOR4 (N2812, N2804, N156, N729, N662);
buf BUF1 (N2813, N2812);
nand NAND4 (N2814, N2808, N236, N1601, N1543);
nor NOR3 (N2815, N2807, N1088, N1203);
and AND3 (N2816, N2810, N2445, N1585);
or OR2 (N2817, N2816, N1901);
nand NAND3 (N2818, N2817, N1700, N1906);
xor XOR2 (N2819, N2815, N493);
xor XOR2 (N2820, N2805, N940);
xor XOR2 (N2821, N2820, N622);
or OR2 (N2822, N2821, N739);
xor XOR2 (N2823, N2802, N1722);
nor NOR3 (N2824, N2790, N801, N1735);
buf BUF1 (N2825, N2822);
nor NOR2 (N2826, N2814, N676);
or OR4 (N2827, N2818, N855, N773, N1448);
and AND2 (N2828, N2827, N226);
xor XOR2 (N2829, N2825, N840);
xor XOR2 (N2830, N2813, N2236);
or OR2 (N2831, N2830, N828);
xor XOR2 (N2832, N2826, N2797);
and AND2 (N2833, N2832, N613);
and AND3 (N2834, N2831, N30, N1724);
or OR3 (N2835, N2828, N762, N1293);
and AND3 (N2836, N2819, N2273, N2604);
nor NOR3 (N2837, N2809, N704, N2232);
not NOT1 (N2838, N2834);
nand NAND4 (N2839, N2833, N616, N684, N1926);
not NOT1 (N2840, N2835);
not NOT1 (N2841, N2824);
not NOT1 (N2842, N2829);
nor NOR3 (N2843, N2801, N1520, N892);
and AND4 (N2844, N2823, N2667, N1914, N2691);
nor NOR3 (N2845, N2811, N2471, N482);
not NOT1 (N2846, N2845);
and AND2 (N2847, N2841, N165);
or OR4 (N2848, N2837, N2220, N1596, N680);
xor XOR2 (N2849, N2846, N2);
xor XOR2 (N2850, N2843, N1579);
not NOT1 (N2851, N2842);
buf BUF1 (N2852, N2839);
nand NAND3 (N2853, N2844, N825, N466);
buf BUF1 (N2854, N2836);
or OR2 (N2855, N2847, N2564);
or OR3 (N2856, N2853, N392, N819);
nor NOR2 (N2857, N2849, N516);
xor XOR2 (N2858, N2838, N2710);
not NOT1 (N2859, N2852);
not NOT1 (N2860, N2859);
and AND3 (N2861, N2857, N2240, N1557);
not NOT1 (N2862, N2858);
xor XOR2 (N2863, N2840, N151);
xor XOR2 (N2864, N2854, N691);
not NOT1 (N2865, N2862);
buf BUF1 (N2866, N2861);
buf BUF1 (N2867, N2855);
nand NAND4 (N2868, N2866, N1611, N2373, N557);
or OR3 (N2869, N2850, N1037, N335);
nand NAND3 (N2870, N2865, N870, N521);
and AND4 (N2871, N2860, N57, N2309, N138);
and AND3 (N2872, N2868, N248, N1670);
xor XOR2 (N2873, N2848, N691);
nand NAND4 (N2874, N2864, N451, N977, N760);
and AND2 (N2875, N2872, N444);
xor XOR2 (N2876, N2867, N2087);
nor NOR4 (N2877, N2876, N1674, N215, N580);
not NOT1 (N2878, N2874);
nand NAND3 (N2879, N2878, N1353, N1667);
nor NOR3 (N2880, N2870, N2879, N2871);
and AND3 (N2881, N610, N1428, N540);
not NOT1 (N2882, N2455);
buf BUF1 (N2883, N2875);
xor XOR2 (N2884, N2856, N2604);
not NOT1 (N2885, N2881);
and AND2 (N2886, N2882, N62);
not NOT1 (N2887, N2884);
not NOT1 (N2888, N2863);
not NOT1 (N2889, N2873);
xor XOR2 (N2890, N2851, N2791);
nor NOR2 (N2891, N2869, N2268);
nand NAND4 (N2892, N2883, N598, N633, N1706);
buf BUF1 (N2893, N2892);
or OR4 (N2894, N2889, N1761, N2398, N2167);
or OR2 (N2895, N2885, N684);
xor XOR2 (N2896, N2886, N790);
xor XOR2 (N2897, N2894, N2315);
nor NOR4 (N2898, N2896, N918, N1780, N2271);
nand NAND3 (N2899, N2890, N543, N1608);
nor NOR3 (N2900, N2877, N1998, N318);
xor XOR2 (N2901, N2893, N1100);
buf BUF1 (N2902, N2900);
xor XOR2 (N2903, N2901, N1746);
nand NAND3 (N2904, N2903, N2001, N1998);
xor XOR2 (N2905, N2898, N1087);
xor XOR2 (N2906, N2895, N165);
and AND4 (N2907, N2902, N989, N2462, N314);
not NOT1 (N2908, N2907);
or OR4 (N2909, N2904, N1818, N2749, N2475);
not NOT1 (N2910, N2908);
not NOT1 (N2911, N2880);
buf BUF1 (N2912, N2905);
xor XOR2 (N2913, N2887, N2397);
and AND4 (N2914, N2899, N56, N2169, N1281);
or OR4 (N2915, N2911, N1594, N2171, N694);
xor XOR2 (N2916, N2897, N2305);
buf BUF1 (N2917, N2891);
not NOT1 (N2918, N2910);
nand NAND2 (N2919, N2909, N2508);
nand NAND2 (N2920, N2912, N1349);
and AND2 (N2921, N2919, N2732);
nand NAND3 (N2922, N2918, N182, N2655);
nor NOR3 (N2923, N2913, N1361, N2119);
and AND2 (N2924, N2920, N479);
buf BUF1 (N2925, N2923);
buf BUF1 (N2926, N2925);
nor NOR4 (N2927, N2914, N927, N205, N2326);
and AND3 (N2928, N2921, N517, N2921);
nor NOR3 (N2929, N2917, N2747, N1825);
xor XOR2 (N2930, N2924, N1252);
xor XOR2 (N2931, N2926, N849);
xor XOR2 (N2932, N2906, N727);
or OR4 (N2933, N2927, N1402, N1128, N2740);
and AND4 (N2934, N2931, N1689, N2547, N2776);
nor NOR2 (N2935, N2930, N1838);
or OR4 (N2936, N2932, N2598, N2040, N2748);
nor NOR3 (N2937, N2915, N988, N178);
nand NAND4 (N2938, N2922, N2063, N2342, N1518);
nor NOR3 (N2939, N2916, N379, N1793);
or OR2 (N2940, N2934, N2522);
or OR2 (N2941, N2928, N1866);
and AND2 (N2942, N2936, N1362);
buf BUF1 (N2943, N2937);
and AND3 (N2944, N2940, N760, N592);
nand NAND3 (N2945, N2938, N1844, N46);
nand NAND3 (N2946, N2929, N143, N549);
nand NAND2 (N2947, N2941, N1396);
xor XOR2 (N2948, N2942, N1676);
and AND2 (N2949, N2943, N1333);
nand NAND2 (N2950, N2945, N543);
nor NOR3 (N2951, N2939, N552, N294);
nand NAND2 (N2952, N2951, N1932);
not NOT1 (N2953, N2948);
xor XOR2 (N2954, N2946, N188);
nor NOR3 (N2955, N2933, N2926, N1283);
buf BUF1 (N2956, N2944);
nand NAND3 (N2957, N2953, N2117, N838);
and AND3 (N2958, N2888, N2511, N1917);
nand NAND2 (N2959, N2956, N338);
or OR3 (N2960, N2935, N2653, N1080);
and AND2 (N2961, N2950, N252);
or OR4 (N2962, N2947, N532, N2487, N1588);
nor NOR2 (N2963, N2955, N1619);
buf BUF1 (N2964, N2959);
xor XOR2 (N2965, N2964, N2006);
nand NAND4 (N2966, N2952, N2079, N533, N842);
xor XOR2 (N2967, N2954, N2373);
buf BUF1 (N2968, N2949);
and AND2 (N2969, N2963, N775);
not NOT1 (N2970, N2969);
and AND4 (N2971, N2967, N653, N1102, N2196);
nor NOR4 (N2972, N2971, N2576, N1709, N910);
buf BUF1 (N2973, N2966);
nand NAND3 (N2974, N2965, N2269, N209);
or OR3 (N2975, N2961, N700, N2188);
xor XOR2 (N2976, N2968, N2368);
buf BUF1 (N2977, N2960);
nand NAND4 (N2978, N2976, N1965, N1514, N1204);
or OR4 (N2979, N2962, N1963, N2198, N364);
and AND2 (N2980, N2977, N514);
nand NAND4 (N2981, N2972, N2405, N2892, N1254);
or OR4 (N2982, N2979, N622, N496, N920);
or OR3 (N2983, N2981, N2504, N922);
xor XOR2 (N2984, N2957, N123);
and AND2 (N2985, N2980, N625);
nor NOR3 (N2986, N2958, N2617, N2912);
and AND3 (N2987, N2973, N1360, N2621);
buf BUF1 (N2988, N2978);
nor NOR3 (N2989, N2982, N2036, N1499);
nand NAND3 (N2990, N2983, N2955, N2761);
and AND3 (N2991, N2988, N2544, N2773);
nand NAND4 (N2992, N2984, N2705, N809, N2232);
nand NAND2 (N2993, N2975, N1394);
nor NOR2 (N2994, N2993, N1973);
xor XOR2 (N2995, N2989, N1989);
and AND2 (N2996, N2991, N613);
or OR2 (N2997, N2996, N2396);
and AND2 (N2998, N2997, N1145);
xor XOR2 (N2999, N2990, N1276);
and AND3 (N3000, N2999, N1451, N393);
nor NOR4 (N3001, N2998, N2485, N2446, N2738);
not NOT1 (N3002, N2970);
or OR4 (N3003, N2994, N2225, N294, N449);
buf BUF1 (N3004, N2987);
or OR2 (N3005, N2992, N2827);
not NOT1 (N3006, N2995);
or OR3 (N3007, N3005, N1218, N1147);
xor XOR2 (N3008, N3000, N2092);
buf BUF1 (N3009, N3002);
and AND3 (N3010, N3003, N2935, N448);
buf BUF1 (N3011, N2986);
nand NAND2 (N3012, N3006, N195);
xor XOR2 (N3013, N3001, N245);
nand NAND2 (N3014, N2985, N1035);
not NOT1 (N3015, N3009);
buf BUF1 (N3016, N2974);
buf BUF1 (N3017, N3010);
or OR3 (N3018, N3013, N358, N428);
nand NAND3 (N3019, N3008, N2405, N2438);
or OR4 (N3020, N3018, N1283, N222, N169);
or OR2 (N3021, N3020, N499);
nand NAND3 (N3022, N3014, N1673, N277);
nand NAND3 (N3023, N3017, N1044, N932);
or OR3 (N3024, N3004, N1867, N2261);
nor NOR4 (N3025, N3015, N698, N2723, N489);
and AND2 (N3026, N3021, N148);
or OR2 (N3027, N3016, N2850);
buf BUF1 (N3028, N3022);
buf BUF1 (N3029, N3011);
or OR3 (N3030, N3028, N163, N332);
xor XOR2 (N3031, N3007, N2035);
xor XOR2 (N3032, N3030, N2400);
buf BUF1 (N3033, N3023);
nor NOR4 (N3034, N3031, N1441, N1423, N934);
nor NOR3 (N3035, N3026, N1839, N2444);
nand NAND2 (N3036, N3029, N2387);
nand NAND4 (N3037, N3024, N228, N238, N1832);
xor XOR2 (N3038, N3036, N1500);
nor NOR4 (N3039, N3019, N2760, N450, N1656);
nor NOR3 (N3040, N3032, N465, N1091);
xor XOR2 (N3041, N3038, N81);
nand NAND3 (N3042, N3037, N875, N890);
not NOT1 (N3043, N3040);
not NOT1 (N3044, N3025);
or OR3 (N3045, N3012, N1802, N2398);
or OR3 (N3046, N3041, N197, N698);
not NOT1 (N3047, N3042);
not NOT1 (N3048, N3047);
nand NAND3 (N3049, N3044, N259, N2870);
xor XOR2 (N3050, N3039, N2702);
nand NAND2 (N3051, N3045, N1247);
and AND3 (N3052, N3027, N1298, N2906);
nor NOR2 (N3053, N3034, N528);
xor XOR2 (N3054, N3051, N2615);
nand NAND3 (N3055, N3052, N617, N1006);
nand NAND2 (N3056, N3048, N207);
or OR2 (N3057, N3049, N1285);
xor XOR2 (N3058, N3033, N78);
not NOT1 (N3059, N3053);
not NOT1 (N3060, N3054);
and AND4 (N3061, N3035, N359, N155, N1300);
buf BUF1 (N3062, N3046);
not NOT1 (N3063, N3043);
not NOT1 (N3064, N3060);
nand NAND2 (N3065, N3059, N133);
nand NAND3 (N3066, N3063, N2801, N998);
not NOT1 (N3067, N3057);
or OR2 (N3068, N3055, N1116);
nand NAND2 (N3069, N3050, N1830);
not NOT1 (N3070, N3062);
nand NAND2 (N3071, N3064, N353);
not NOT1 (N3072, N3056);
or OR4 (N3073, N3067, N1941, N1071, N2900);
buf BUF1 (N3074, N3068);
nor NOR2 (N3075, N3074, N704);
not NOT1 (N3076, N3075);
or OR2 (N3077, N3070, N338);
buf BUF1 (N3078, N3066);
buf BUF1 (N3079, N3061);
and AND4 (N3080, N3069, N2701, N2135, N1453);
and AND4 (N3081, N3058, N2730, N1630, N475);
and AND3 (N3082, N3073, N2528, N348);
buf BUF1 (N3083, N3065);
buf BUF1 (N3084, N3080);
buf BUF1 (N3085, N3084);
not NOT1 (N3086, N3082);
or OR2 (N3087, N3086, N541);
buf BUF1 (N3088, N3077);
nor NOR3 (N3089, N3085, N1762, N1955);
buf BUF1 (N3090, N3076);
nor NOR3 (N3091, N3089, N1821, N586);
buf BUF1 (N3092, N3091);
not NOT1 (N3093, N3088);
nor NOR2 (N3094, N3087, N2448);
buf BUF1 (N3095, N3093);
nand NAND4 (N3096, N3083, N1236, N1552, N3002);
not NOT1 (N3097, N3071);
and AND2 (N3098, N3094, N2316);
or OR3 (N3099, N3096, N206, N2964);
nand NAND3 (N3100, N3078, N611, N632);
buf BUF1 (N3101, N3090);
not NOT1 (N3102, N3098);
nor NOR3 (N3103, N3081, N2845, N1850);
or OR4 (N3104, N3101, N220, N791, N406);
not NOT1 (N3105, N3099);
nor NOR4 (N3106, N3103, N1482, N155, N1456);
nand NAND2 (N3107, N3104, N2391);
buf BUF1 (N3108, N3072);
xor XOR2 (N3109, N3097, N2879);
buf BUF1 (N3110, N3106);
nor NOR3 (N3111, N3108, N2262, N809);
buf BUF1 (N3112, N3105);
nor NOR4 (N3113, N3107, N3019, N217, N1652);
or OR2 (N3114, N3092, N2406);
buf BUF1 (N3115, N3113);
or OR4 (N3116, N3095, N2854, N838, N1794);
xor XOR2 (N3117, N3079, N2283);
nand NAND2 (N3118, N3110, N1687);
and AND4 (N3119, N3111, N692, N2054, N477);
nand NAND2 (N3120, N3109, N2621);
nor NOR3 (N3121, N3114, N2488, N78);
nand NAND4 (N3122, N3112, N2033, N2805, N1055);
nand NAND3 (N3123, N3120, N189, N1708);
nor NOR3 (N3124, N3116, N330, N87);
and AND3 (N3125, N3119, N1412, N1316);
or OR2 (N3126, N3122, N2294);
xor XOR2 (N3127, N3117, N2125);
or OR2 (N3128, N3125, N1457);
not NOT1 (N3129, N3115);
nor NOR4 (N3130, N3126, N138, N2157, N710);
buf BUF1 (N3131, N3123);
or OR3 (N3132, N3130, N2216, N3031);
or OR4 (N3133, N3131, N1836, N2969, N545);
xor XOR2 (N3134, N3118, N1711);
or OR3 (N3135, N3129, N1612, N3097);
xor XOR2 (N3136, N3133, N2520);
nand NAND3 (N3137, N3134, N656, N2881);
xor XOR2 (N3138, N3102, N151);
or OR4 (N3139, N3135, N1633, N135, N1344);
nand NAND2 (N3140, N3121, N453);
buf BUF1 (N3141, N3132);
not NOT1 (N3142, N3100);
and AND2 (N3143, N3138, N1970);
nand NAND4 (N3144, N3141, N13, N1999, N2095);
nor NOR3 (N3145, N3143, N1599, N738);
and AND4 (N3146, N3142, N2271, N2697, N416);
not NOT1 (N3147, N3128);
or OR3 (N3148, N3124, N782, N698);
or OR3 (N3149, N3145, N45, N1983);
buf BUF1 (N3150, N3139);
or OR4 (N3151, N3150, N2545, N1488, N430);
or OR4 (N3152, N3148, N2211, N1525, N1323);
nor NOR3 (N3153, N3137, N102, N1609);
buf BUF1 (N3154, N3147);
not NOT1 (N3155, N3127);
or OR2 (N3156, N3154, N1142);
and AND4 (N3157, N3153, N1510, N659, N3030);
not NOT1 (N3158, N3155);
and AND4 (N3159, N3149, N453, N2079, N1621);
or OR3 (N3160, N3151, N1308, N1552);
and AND4 (N3161, N3152, N71, N2284, N2464);
nand NAND4 (N3162, N3146, N1811, N2762, N2306);
nor NOR3 (N3163, N3162, N2876, N173);
xor XOR2 (N3164, N3156, N378);
buf BUF1 (N3165, N3140);
nor NOR3 (N3166, N3165, N1220, N437);
xor XOR2 (N3167, N3160, N1762);
or OR2 (N3168, N3166, N1347);
nor NOR3 (N3169, N3168, N1573, N2127);
nand NAND4 (N3170, N3161, N742, N2284, N2439);
or OR4 (N3171, N3157, N2254, N612, N274);
nand NAND4 (N3172, N3144, N1675, N1602, N1944);
and AND2 (N3173, N3163, N2087);
xor XOR2 (N3174, N3169, N835);
nor NOR2 (N3175, N3136, N551);
and AND3 (N3176, N3158, N1109, N1382);
buf BUF1 (N3177, N3167);
nand NAND2 (N3178, N3159, N2115);
buf BUF1 (N3179, N3176);
nor NOR4 (N3180, N3173, N1715, N2003, N826);
xor XOR2 (N3181, N3177, N1662);
nand NAND4 (N3182, N3178, N118, N1383, N396);
buf BUF1 (N3183, N3181);
buf BUF1 (N3184, N3180);
nor NOR3 (N3185, N3179, N2552, N1163);
xor XOR2 (N3186, N3171, N2940);
and AND2 (N3187, N3164, N723);
or OR3 (N3188, N3185, N3044, N2303);
nor NOR4 (N3189, N3172, N1903, N97, N2228);
xor XOR2 (N3190, N3189, N3046);
nor NOR4 (N3191, N3187, N688, N2870, N1170);
nor NOR3 (N3192, N3186, N291, N1880);
nand NAND3 (N3193, N3174, N1636, N2421);
not NOT1 (N3194, N3182);
nand NAND3 (N3195, N3170, N461, N2767);
and AND4 (N3196, N3191, N837, N577, N775);
nand NAND2 (N3197, N3195, N192);
not NOT1 (N3198, N3196);
nand NAND2 (N3199, N3184, N873);
buf BUF1 (N3200, N3192);
nor NOR3 (N3201, N3193, N2162, N3095);
buf BUF1 (N3202, N3201);
and AND2 (N3203, N3202, N232);
and AND2 (N3204, N3194, N3055);
buf BUF1 (N3205, N3183);
xor XOR2 (N3206, N3175, N2116);
or OR2 (N3207, N3190, N160);
buf BUF1 (N3208, N3198);
or OR4 (N3209, N3204, N1951, N2378, N427);
not NOT1 (N3210, N3199);
nand NAND2 (N3211, N3206, N1658);
and AND3 (N3212, N3207, N1515, N51);
or OR4 (N3213, N3211, N2834, N2435, N1874);
xor XOR2 (N3214, N3203, N342);
xor XOR2 (N3215, N3197, N1309);
and AND4 (N3216, N3209, N2871, N192, N2887);
not NOT1 (N3217, N3212);
nand NAND4 (N3218, N3188, N3108, N601, N135);
not NOT1 (N3219, N3217);
nand NAND4 (N3220, N3200, N2696, N1201, N2844);
xor XOR2 (N3221, N3205, N1631);
not NOT1 (N3222, N3221);
not NOT1 (N3223, N3220);
not NOT1 (N3224, N3208);
xor XOR2 (N3225, N3223, N2168);
nor NOR3 (N3226, N3210, N2594, N2409);
nand NAND4 (N3227, N3226, N2630, N2786, N633);
nor NOR2 (N3228, N3222, N469);
nor NOR4 (N3229, N3219, N450, N926, N3087);
buf BUF1 (N3230, N3229);
xor XOR2 (N3231, N3218, N718);
nor NOR4 (N3232, N3224, N20, N3036, N3194);
and AND3 (N3233, N3216, N1211, N2855);
nand NAND3 (N3234, N3225, N2929, N3151);
nand NAND2 (N3235, N3231, N419);
not NOT1 (N3236, N3235);
nand NAND3 (N3237, N3228, N28, N2076);
and AND3 (N3238, N3232, N619, N2705);
xor XOR2 (N3239, N3236, N1736);
or OR2 (N3240, N3237, N2193);
xor XOR2 (N3241, N3238, N2257);
nor NOR4 (N3242, N3230, N381, N2777, N325);
not NOT1 (N3243, N3215);
or OR2 (N3244, N3241, N555);
or OR3 (N3245, N3244, N33, N935);
and AND4 (N3246, N3234, N721, N2, N1476);
xor XOR2 (N3247, N3227, N2639);
xor XOR2 (N3248, N3247, N2319);
nor NOR4 (N3249, N3245, N1807, N104, N1031);
nand NAND2 (N3250, N3248, N516);
nand NAND2 (N3251, N3213, N1546);
nand NAND3 (N3252, N3249, N2288, N687);
and AND3 (N3253, N3239, N2027, N1884);
and AND3 (N3254, N3250, N1550, N2621);
nor NOR3 (N3255, N3240, N2448, N2043);
not NOT1 (N3256, N3233);
xor XOR2 (N3257, N3252, N2067);
not NOT1 (N3258, N3214);
xor XOR2 (N3259, N3251, N3047);
or OR3 (N3260, N3258, N773, N2986);
nor NOR3 (N3261, N3243, N1582, N2633);
nor NOR3 (N3262, N3253, N3092, N677);
buf BUF1 (N3263, N3254);
and AND4 (N3264, N3261, N279, N674, N2481);
buf BUF1 (N3265, N3255);
nor NOR3 (N3266, N3259, N76, N2758);
not NOT1 (N3267, N3242);
nor NOR3 (N3268, N3265, N3215, N1673);
and AND4 (N3269, N3264, N799, N3232, N2154);
not NOT1 (N3270, N3246);
and AND4 (N3271, N3257, N1584, N2477, N1912);
nor NOR4 (N3272, N3263, N3009, N3151, N938);
or OR4 (N3273, N3266, N880, N1230, N2179);
buf BUF1 (N3274, N3273);
nand NAND4 (N3275, N3272, N2360, N2077, N589);
or OR3 (N3276, N3274, N1023, N2644);
or OR4 (N3277, N3268, N2705, N151, N1143);
nor NOR2 (N3278, N3271, N504);
and AND4 (N3279, N3267, N1157, N828, N2007);
or OR3 (N3280, N3276, N2494, N823);
xor XOR2 (N3281, N3280, N743);
xor XOR2 (N3282, N3260, N2220);
not NOT1 (N3283, N3269);
or OR2 (N3284, N3282, N893);
not NOT1 (N3285, N3284);
or OR4 (N3286, N3275, N958, N2905, N1003);
not NOT1 (N3287, N3281);
buf BUF1 (N3288, N3262);
buf BUF1 (N3289, N3277);
xor XOR2 (N3290, N3256, N227);
not NOT1 (N3291, N3270);
and AND3 (N3292, N3291, N955, N837);
xor XOR2 (N3293, N3285, N1543);
nor NOR2 (N3294, N3278, N1205);
not NOT1 (N3295, N3279);
and AND2 (N3296, N3292, N2080);
nand NAND3 (N3297, N3293, N1968, N1409);
nand NAND2 (N3298, N3286, N2974);
nand NAND2 (N3299, N3298, N1129);
not NOT1 (N3300, N3295);
nand NAND4 (N3301, N3300, N2217, N1131, N1356);
or OR3 (N3302, N3290, N27, N2456);
nor NOR2 (N3303, N3283, N2842);
xor XOR2 (N3304, N3287, N99);
buf BUF1 (N3305, N3299);
xor XOR2 (N3306, N3301, N2432);
xor XOR2 (N3307, N3303, N2802);
nor NOR4 (N3308, N3304, N2123, N753, N1808);
and AND3 (N3309, N3294, N480, N899);
nand NAND3 (N3310, N3302, N3262, N43);
xor XOR2 (N3311, N3297, N384);
or OR3 (N3312, N3308, N1027, N98);
nand NAND2 (N3313, N3289, N2360);
xor XOR2 (N3314, N3305, N1255);
not NOT1 (N3315, N3309);
buf BUF1 (N3316, N3311);
nand NAND3 (N3317, N3313, N3286, N2960);
and AND3 (N3318, N3296, N2536, N1900);
or OR3 (N3319, N3314, N2141, N1839);
xor XOR2 (N3320, N3315, N467);
nand NAND3 (N3321, N3312, N2195, N2265);
or OR2 (N3322, N3316, N820);
not NOT1 (N3323, N3307);
nand NAND4 (N3324, N3317, N3073, N2025, N3078);
xor XOR2 (N3325, N3323, N1949);
buf BUF1 (N3326, N3306);
buf BUF1 (N3327, N3310);
not NOT1 (N3328, N3318);
nand NAND2 (N3329, N3328, N2254);
not NOT1 (N3330, N3325);
not NOT1 (N3331, N3329);
buf BUF1 (N3332, N3324);
not NOT1 (N3333, N3320);
xor XOR2 (N3334, N3330, N1543);
and AND4 (N3335, N3288, N511, N2568, N2655);
not NOT1 (N3336, N3334);
nand NAND2 (N3337, N3333, N806);
nand NAND3 (N3338, N3336, N3014, N3128);
xor XOR2 (N3339, N3335, N126);
or OR4 (N3340, N3319, N1033, N1713, N3261);
not NOT1 (N3341, N3337);
xor XOR2 (N3342, N3327, N2243);
buf BUF1 (N3343, N3331);
not NOT1 (N3344, N3332);
nor NOR4 (N3345, N3344, N2919, N379, N2384);
not NOT1 (N3346, N3342);
or OR4 (N3347, N3341, N339, N146, N2626);
xor XOR2 (N3348, N3347, N3142);
not NOT1 (N3349, N3343);
nand NAND2 (N3350, N3348, N2804);
or OR2 (N3351, N3345, N2165);
not NOT1 (N3352, N3321);
nand NAND4 (N3353, N3338, N2583, N1632, N2663);
nand NAND4 (N3354, N3350, N3290, N1016, N194);
not NOT1 (N3355, N3351);
or OR2 (N3356, N3349, N813);
and AND4 (N3357, N3339, N1821, N642, N1227);
buf BUF1 (N3358, N3352);
nor NOR3 (N3359, N3326, N2444, N3296);
and AND4 (N3360, N3359, N253, N2031, N2189);
and AND4 (N3361, N3354, N1553, N3038, N2885);
and AND4 (N3362, N3360, N589, N1441, N1225);
nor NOR2 (N3363, N3362, N2316);
or OR3 (N3364, N3358, N464, N799);
nor NOR2 (N3365, N3363, N2150);
xor XOR2 (N3366, N3356, N2804);
xor XOR2 (N3367, N3361, N77);
nand NAND3 (N3368, N3346, N3154, N2028);
or OR4 (N3369, N3365, N2082, N2439, N1492);
nor NOR3 (N3370, N3368, N1864, N1222);
nand NAND3 (N3371, N3322, N407, N3162);
nand NAND4 (N3372, N3366, N2155, N2757, N1169);
xor XOR2 (N3373, N3340, N589);
nand NAND3 (N3374, N3370, N1499, N1396);
or OR2 (N3375, N3357, N435);
not NOT1 (N3376, N3364);
not NOT1 (N3377, N3373);
buf BUF1 (N3378, N3355);
buf BUF1 (N3379, N3367);
xor XOR2 (N3380, N3369, N1443);
or OR4 (N3381, N3371, N1554, N1931, N1161);
nor NOR2 (N3382, N3375, N2912);
xor XOR2 (N3383, N3378, N621);
not NOT1 (N3384, N3382);
xor XOR2 (N3385, N3383, N2715);
and AND4 (N3386, N3353, N349, N3361, N702);
not NOT1 (N3387, N3385);
buf BUF1 (N3388, N3381);
xor XOR2 (N3389, N3377, N2149);
nor NOR3 (N3390, N3386, N1474, N856);
buf BUF1 (N3391, N3372);
nand NAND2 (N3392, N3380, N282);
or OR3 (N3393, N3391, N1170, N2256);
and AND3 (N3394, N3387, N1830, N2123);
or OR4 (N3395, N3379, N2296, N663, N859);
buf BUF1 (N3396, N3384);
nor NOR3 (N3397, N3396, N9, N2424);
or OR2 (N3398, N3395, N2530);
not NOT1 (N3399, N3393);
nor NOR2 (N3400, N3374, N3327);
not NOT1 (N3401, N3389);
not NOT1 (N3402, N3388);
xor XOR2 (N3403, N3398, N55);
not NOT1 (N3404, N3390);
nor NOR3 (N3405, N3397, N683, N3111);
xor XOR2 (N3406, N3405, N1231);
xor XOR2 (N3407, N3406, N1841);
buf BUF1 (N3408, N3407);
or OR3 (N3409, N3403, N386, N2367);
nand NAND3 (N3410, N3409, N1388, N3133);
buf BUF1 (N3411, N3394);
nor NOR2 (N3412, N3411, N2289);
xor XOR2 (N3413, N3399, N1066);
xor XOR2 (N3414, N3401, N1041);
nand NAND3 (N3415, N3404, N1434, N3299);
nor NOR2 (N3416, N3413, N3167);
nor NOR2 (N3417, N3392, N546);
not NOT1 (N3418, N3415);
buf BUF1 (N3419, N3418);
and AND4 (N3420, N3408, N2573, N225, N407);
not NOT1 (N3421, N3402);
not NOT1 (N3422, N3400);
nor NOR3 (N3423, N3419, N384, N1406);
or OR2 (N3424, N3421, N697);
xor XOR2 (N3425, N3417, N535);
or OR4 (N3426, N3414, N2574, N3200, N1074);
or OR3 (N3427, N3422, N1907, N2171);
xor XOR2 (N3428, N3425, N3360);
or OR3 (N3429, N3410, N3099, N1114);
or OR2 (N3430, N3424, N2390);
nand NAND3 (N3431, N3429, N825, N1868);
nand NAND3 (N3432, N3430, N3403, N1333);
or OR3 (N3433, N3423, N347, N1759);
not NOT1 (N3434, N3416);
nand NAND4 (N3435, N3426, N2957, N433, N3131);
nand NAND3 (N3436, N3376, N441, N2950);
xor XOR2 (N3437, N3428, N471);
or OR2 (N3438, N3432, N2889);
and AND4 (N3439, N3438, N3363, N1199, N1545);
and AND3 (N3440, N3420, N244, N1819);
nor NOR4 (N3441, N3439, N2316, N2934, N3353);
and AND4 (N3442, N3436, N2120, N3023, N2018);
nand NAND3 (N3443, N3440, N2504, N3055);
buf BUF1 (N3444, N3435);
nor NOR3 (N3445, N3443, N3440, N768);
and AND2 (N3446, N3437, N1562);
and AND4 (N3447, N3427, N1810, N1383, N95);
nor NOR4 (N3448, N3445, N3196, N254, N2052);
nand NAND4 (N3449, N3447, N3385, N3237, N2761);
not NOT1 (N3450, N3434);
nor NOR4 (N3451, N3433, N13, N2066, N2985);
or OR3 (N3452, N3444, N1028, N1469);
buf BUF1 (N3453, N3451);
xor XOR2 (N3454, N3442, N2118);
buf BUF1 (N3455, N3446);
and AND2 (N3456, N3453, N3163);
and AND2 (N3457, N3412, N3063);
nor NOR2 (N3458, N3441, N3118);
xor XOR2 (N3459, N3448, N1699);
and AND3 (N3460, N3455, N749, N2260);
nand NAND3 (N3461, N3450, N951, N148);
buf BUF1 (N3462, N3456);
nor NOR2 (N3463, N3449, N897);
not NOT1 (N3464, N3460);
buf BUF1 (N3465, N3461);
xor XOR2 (N3466, N3458, N2611);
nand NAND2 (N3467, N3466, N184);
not NOT1 (N3468, N3467);
xor XOR2 (N3469, N3463, N2654);
nor NOR2 (N3470, N3457, N1116);
and AND2 (N3471, N3452, N1230);
or OR4 (N3472, N3465, N2881, N1685, N1635);
buf BUF1 (N3473, N3454);
or OR4 (N3474, N3470, N1427, N2173, N1141);
nand NAND4 (N3475, N3468, N579, N2728, N2795);
and AND3 (N3476, N3462, N756, N2565);
xor XOR2 (N3477, N3431, N705);
nor NOR3 (N3478, N3464, N1509, N1763);
nor NOR4 (N3479, N3477, N2903, N3161, N1196);
xor XOR2 (N3480, N3471, N1589);
not NOT1 (N3481, N3469);
buf BUF1 (N3482, N3479);
xor XOR2 (N3483, N3475, N1250);
and AND3 (N3484, N3478, N170, N1694);
xor XOR2 (N3485, N3480, N2718);
nor NOR2 (N3486, N3459, N2404);
nand NAND3 (N3487, N3485, N3450, N3179);
not NOT1 (N3488, N3487);
or OR4 (N3489, N3472, N2535, N2416, N794);
nor NOR4 (N3490, N3476, N1764, N605, N315);
nor NOR4 (N3491, N3484, N2869, N3423, N3267);
and AND3 (N3492, N3482, N2349, N492);
nor NOR2 (N3493, N3489, N377);
and AND4 (N3494, N3473, N2827, N264, N1777);
xor XOR2 (N3495, N3493, N856);
nand NAND3 (N3496, N3491, N2721, N2157);
not NOT1 (N3497, N3495);
or OR2 (N3498, N3488, N686);
nor NOR3 (N3499, N3497, N3158, N1707);
nand NAND4 (N3500, N3498, N3467, N3318, N438);
nand NAND4 (N3501, N3486, N2522, N1027, N3385);
or OR3 (N3502, N3490, N3132, N885);
nor NOR2 (N3503, N3481, N2468);
xor XOR2 (N3504, N3499, N1939);
not NOT1 (N3505, N3501);
not NOT1 (N3506, N3474);
buf BUF1 (N3507, N3494);
and AND3 (N3508, N3483, N82, N2561);
or OR2 (N3509, N3507, N1774);
or OR3 (N3510, N3503, N64, N2573);
and AND3 (N3511, N3492, N2820, N2673);
and AND2 (N3512, N3500, N1959);
xor XOR2 (N3513, N3502, N823);
nand NAND2 (N3514, N3496, N1201);
and AND4 (N3515, N3509, N400, N1778, N1715);
xor XOR2 (N3516, N3512, N1546);
nor NOR4 (N3517, N3511, N2375, N2119, N1085);
and AND4 (N3518, N3517, N49, N1275, N2508);
or OR4 (N3519, N3518, N1803, N442, N2567);
and AND2 (N3520, N3510, N616);
nor NOR4 (N3521, N3515, N1356, N1863, N3332);
nor NOR4 (N3522, N3506, N1890, N960, N2036);
buf BUF1 (N3523, N3520);
xor XOR2 (N3524, N3504, N909);
buf BUF1 (N3525, N3523);
nand NAND4 (N3526, N3514, N2078, N963, N3278);
buf BUF1 (N3527, N3525);
nand NAND3 (N3528, N3505, N3204, N1462);
nor NOR4 (N3529, N3521, N935, N9, N341);
and AND4 (N3530, N3508, N1874, N1148, N2323);
and AND4 (N3531, N3519, N466, N3337, N416);
and AND2 (N3532, N3526, N2684);
xor XOR2 (N3533, N3528, N1438);
buf BUF1 (N3534, N3524);
xor XOR2 (N3535, N3534, N1671);
nand NAND4 (N3536, N3522, N1790, N2963, N2811);
not NOT1 (N3537, N3529);
or OR4 (N3538, N3531, N3272, N2373, N1262);
nand NAND3 (N3539, N3533, N1474, N730);
or OR4 (N3540, N3539, N2385, N2994, N3093);
or OR4 (N3541, N3540, N1920, N2360, N2031);
buf BUF1 (N3542, N3532);
nor NOR4 (N3543, N3541, N3147, N862, N1245);
xor XOR2 (N3544, N3538, N2708);
xor XOR2 (N3545, N3516, N1305);
buf BUF1 (N3546, N3513);
or OR2 (N3547, N3535, N2301);
xor XOR2 (N3548, N3527, N1922);
nor NOR2 (N3549, N3530, N1331);
buf BUF1 (N3550, N3536);
not NOT1 (N3551, N3550);
or OR3 (N3552, N3542, N1436, N2870);
nand NAND3 (N3553, N3537, N2072, N3212);
nor NOR3 (N3554, N3552, N2193, N449);
xor XOR2 (N3555, N3554, N2971);
nor NOR2 (N3556, N3548, N321);
buf BUF1 (N3557, N3553);
or OR4 (N3558, N3555, N3064, N264, N3343);
and AND3 (N3559, N3556, N1619, N482);
xor XOR2 (N3560, N3545, N1452);
xor XOR2 (N3561, N3560, N1387);
and AND3 (N3562, N3559, N2213, N558);
nand NAND4 (N3563, N3543, N480, N2817, N232);
buf BUF1 (N3564, N3546);
nand NAND3 (N3565, N3561, N2883, N2942);
or OR3 (N3566, N3558, N2584, N3239);
or OR4 (N3567, N3551, N3091, N587, N1361);
buf BUF1 (N3568, N3547);
and AND2 (N3569, N3564, N1540);
or OR3 (N3570, N3563, N2875, N2463);
or OR3 (N3571, N3566, N731, N341);
and AND4 (N3572, N3569, N3372, N2360, N2153);
or OR4 (N3573, N3557, N2582, N1123, N693);
or OR2 (N3574, N3567, N1363);
nor NOR3 (N3575, N3568, N1904, N2341);
buf BUF1 (N3576, N3574);
nand NAND4 (N3577, N3575, N1502, N3126, N3175);
nand NAND4 (N3578, N3544, N2431, N1663, N2859);
xor XOR2 (N3579, N3576, N1396);
xor XOR2 (N3580, N3570, N1862);
not NOT1 (N3581, N3572);
xor XOR2 (N3582, N3577, N2242);
and AND3 (N3583, N3565, N1839, N2401);
nand NAND2 (N3584, N3581, N1762);
buf BUF1 (N3585, N3583);
and AND3 (N3586, N3578, N1802, N772);
not NOT1 (N3587, N3580);
buf BUF1 (N3588, N3573);
or OR3 (N3589, N3571, N2402, N672);
xor XOR2 (N3590, N3586, N2037);
buf BUF1 (N3591, N3589);
and AND4 (N3592, N3562, N1576, N1280, N2111);
not NOT1 (N3593, N3549);
buf BUF1 (N3594, N3585);
xor XOR2 (N3595, N3587, N2202);
nor NOR3 (N3596, N3592, N1509, N2950);
and AND4 (N3597, N3582, N1671, N3312, N2670);
nor NOR2 (N3598, N3596, N2946);
and AND2 (N3599, N3591, N789);
or OR4 (N3600, N3598, N2679, N3463, N636);
nor NOR3 (N3601, N3600, N920, N1586);
or OR2 (N3602, N3594, N1005);
nor NOR2 (N3603, N3595, N3229);
nor NOR2 (N3604, N3579, N1783);
and AND4 (N3605, N3599, N3069, N280, N2796);
xor XOR2 (N3606, N3605, N1823);
xor XOR2 (N3607, N3606, N3260);
not NOT1 (N3608, N3588);
or OR2 (N3609, N3604, N1279);
nor NOR2 (N3610, N3603, N681);
or OR3 (N3611, N3610, N207, N2177);
nor NOR3 (N3612, N3611, N1360, N2748);
and AND4 (N3613, N3590, N2561, N1483, N3366);
or OR3 (N3614, N3609, N2188, N2704);
xor XOR2 (N3615, N3602, N311);
xor XOR2 (N3616, N3608, N3239);
buf BUF1 (N3617, N3615);
buf BUF1 (N3618, N3616);
buf BUF1 (N3619, N3614);
buf BUF1 (N3620, N3584);
not NOT1 (N3621, N3619);
or OR4 (N3622, N3621, N2976, N809, N1149);
and AND2 (N3623, N3622, N417);
xor XOR2 (N3624, N3607, N1945);
not NOT1 (N3625, N3623);
xor XOR2 (N3626, N3612, N3363);
xor XOR2 (N3627, N3613, N3196);
not NOT1 (N3628, N3618);
or OR4 (N3629, N3624, N2848, N638, N1976);
nand NAND4 (N3630, N3629, N117, N3602, N2460);
nor NOR3 (N3631, N3593, N335, N2507);
nor NOR4 (N3632, N3630, N636, N2710, N2285);
nand NAND3 (N3633, N3626, N3568, N1352);
and AND3 (N3634, N3617, N773, N3133);
or OR2 (N3635, N3627, N338);
nand NAND2 (N3636, N3632, N2409);
xor XOR2 (N3637, N3628, N1447);
nor NOR4 (N3638, N3635, N3010, N2152, N3391);
nand NAND3 (N3639, N3636, N2874, N2564);
or OR3 (N3640, N3601, N1266, N1195);
xor XOR2 (N3641, N3631, N1293);
and AND2 (N3642, N3625, N1678);
not NOT1 (N3643, N3597);
xor XOR2 (N3644, N3643, N691);
or OR4 (N3645, N3641, N1448, N1600, N796);
buf BUF1 (N3646, N3645);
xor XOR2 (N3647, N3642, N2517);
nand NAND2 (N3648, N3639, N1348);
nand NAND4 (N3649, N3637, N3202, N865, N370);
buf BUF1 (N3650, N3648);
not NOT1 (N3651, N3646);
or OR2 (N3652, N3633, N884);
and AND2 (N3653, N3651, N2674);
nand NAND2 (N3654, N3650, N2555);
or OR3 (N3655, N3638, N1290, N428);
nand NAND2 (N3656, N3644, N9);
nor NOR4 (N3657, N3652, N3535, N2447, N348);
nand NAND3 (N3658, N3640, N2146, N871);
and AND2 (N3659, N3620, N1570);
nor NOR4 (N3660, N3654, N1999, N2566, N1941);
nand NAND2 (N3661, N3634, N3023);
not NOT1 (N3662, N3658);
or OR2 (N3663, N3647, N2837);
not NOT1 (N3664, N3649);
xor XOR2 (N3665, N3664, N2388);
nor NOR2 (N3666, N3653, N3178);
nor NOR2 (N3667, N3663, N760);
buf BUF1 (N3668, N3659);
nand NAND3 (N3669, N3665, N2182, N38);
not NOT1 (N3670, N3656);
xor XOR2 (N3671, N3668, N3521);
nand NAND2 (N3672, N3666, N1188);
and AND3 (N3673, N3661, N320, N3502);
not NOT1 (N3674, N3670);
nor NOR3 (N3675, N3669, N376, N517);
buf BUF1 (N3676, N3662);
buf BUF1 (N3677, N3676);
buf BUF1 (N3678, N3657);
buf BUF1 (N3679, N3674);
buf BUF1 (N3680, N3675);
or OR2 (N3681, N3671, N614);
xor XOR2 (N3682, N3680, N2051);
not NOT1 (N3683, N3672);
not NOT1 (N3684, N3667);
not NOT1 (N3685, N3660);
nor NOR4 (N3686, N3678, N3362, N44, N86);
and AND2 (N3687, N3684, N1593);
nor NOR2 (N3688, N3679, N1402);
xor XOR2 (N3689, N3686, N3500);
nand NAND3 (N3690, N3682, N2784, N3591);
not NOT1 (N3691, N3673);
nand NAND3 (N3692, N3689, N2951, N2778);
nand NAND2 (N3693, N3692, N1256);
and AND4 (N3694, N3688, N3402, N2998, N2001);
and AND2 (N3695, N3693, N1630);
or OR2 (N3696, N3655, N2542);
nor NOR3 (N3697, N3683, N506, N398);
nor NOR2 (N3698, N3681, N3091);
not NOT1 (N3699, N3687);
not NOT1 (N3700, N3694);
xor XOR2 (N3701, N3685, N219);
buf BUF1 (N3702, N3695);
nand NAND2 (N3703, N3697, N1470);
and AND3 (N3704, N3699, N2762, N3079);
xor XOR2 (N3705, N3704, N3136);
and AND4 (N3706, N3690, N208, N2436, N1328);
nand NAND3 (N3707, N3696, N649, N1348);
and AND4 (N3708, N3700, N272, N3392, N2470);
buf BUF1 (N3709, N3701);
nor NOR4 (N3710, N3705, N2824, N1788, N1942);
nand NAND4 (N3711, N3703, N905, N2643, N45);
and AND4 (N3712, N3677, N1608, N35, N3061);
nand NAND4 (N3713, N3707, N1334, N3529, N892);
nor NOR2 (N3714, N3712, N3025);
not NOT1 (N3715, N3709);
nor NOR4 (N3716, N3713, N3356, N2651, N176);
or OR3 (N3717, N3691, N1447, N665);
or OR2 (N3718, N3717, N1637);
and AND2 (N3719, N3702, N2981);
not NOT1 (N3720, N3698);
xor XOR2 (N3721, N3720, N663);
nor NOR4 (N3722, N3718, N2095, N472, N3336);
not NOT1 (N3723, N3722);
nand NAND3 (N3724, N3706, N2274, N1073);
buf BUF1 (N3725, N3715);
xor XOR2 (N3726, N3719, N2365);
and AND3 (N3727, N3721, N2880, N1861);
nand NAND2 (N3728, N3710, N1169);
nor NOR3 (N3729, N3727, N2172, N1069);
and AND4 (N3730, N3729, N579, N2004, N2638);
nand NAND3 (N3731, N3711, N400, N3708);
buf BUF1 (N3732, N2494);
nand NAND2 (N3733, N3726, N1991);
not NOT1 (N3734, N3723);
nand NAND2 (N3735, N3730, N2833);
xor XOR2 (N3736, N3716, N1703);
nand NAND2 (N3737, N3724, N70);
buf BUF1 (N3738, N3728);
buf BUF1 (N3739, N3714);
buf BUF1 (N3740, N3738);
xor XOR2 (N3741, N3733, N1231);
buf BUF1 (N3742, N3739);
not NOT1 (N3743, N3740);
and AND2 (N3744, N3741, N1138);
nand NAND2 (N3745, N3744, N1580);
nand NAND4 (N3746, N3736, N3577, N1774, N3541);
nand NAND3 (N3747, N3745, N604, N3581);
nor NOR2 (N3748, N3743, N1258);
not NOT1 (N3749, N3742);
nor NOR2 (N3750, N3732, N3508);
nand NAND3 (N3751, N3748, N2991, N3746);
buf BUF1 (N3752, N2904);
buf BUF1 (N3753, N3751);
nand NAND3 (N3754, N3737, N649, N3659);
buf BUF1 (N3755, N3735);
nand NAND3 (N3756, N3754, N286, N1085);
buf BUF1 (N3757, N3756);
buf BUF1 (N3758, N3752);
not NOT1 (N3759, N3758);
nand NAND2 (N3760, N3759, N902);
nor NOR4 (N3761, N3750, N2928, N56, N2963);
or OR4 (N3762, N3734, N2673, N1469, N980);
and AND4 (N3763, N3755, N508, N619, N1490);
xor XOR2 (N3764, N3762, N541);
and AND4 (N3765, N3725, N123, N3015, N3520);
xor XOR2 (N3766, N3731, N2382);
and AND3 (N3767, N3765, N2729, N1455);
nor NOR2 (N3768, N3764, N3039);
or OR3 (N3769, N3757, N2934, N1450);
nor NOR2 (N3770, N3766, N1103);
or OR4 (N3771, N3761, N2401, N3285, N1802);
buf BUF1 (N3772, N3767);
nor NOR2 (N3773, N3771, N2381);
not NOT1 (N3774, N3763);
nand NAND4 (N3775, N3774, N1887, N1647, N2317);
nand NAND2 (N3776, N3772, N503);
and AND2 (N3777, N3747, N1);
nand NAND4 (N3778, N3777, N3192, N328, N1235);
or OR3 (N3779, N3776, N2283, N498);
and AND4 (N3780, N3768, N1965, N3532, N2621);
or OR2 (N3781, N3780, N3589);
or OR2 (N3782, N3769, N3606);
or OR4 (N3783, N3782, N322, N1403, N3555);
and AND3 (N3784, N3781, N3651, N3105);
nor NOR2 (N3785, N3779, N2140);
and AND2 (N3786, N3778, N2447);
and AND3 (N3787, N3753, N3318, N2313);
or OR2 (N3788, N3770, N3311);
xor XOR2 (N3789, N3787, N411);
nor NOR3 (N3790, N3789, N439, N2999);
not NOT1 (N3791, N3788);
and AND4 (N3792, N3749, N1057, N254, N3083);
and AND3 (N3793, N3792, N1491, N1581);
and AND3 (N3794, N3783, N3102, N3473);
or OR4 (N3795, N3790, N1380, N1765, N3725);
buf BUF1 (N3796, N3793);
nor NOR4 (N3797, N3786, N1206, N750, N2326);
nand NAND4 (N3798, N3784, N1023, N2838, N2185);
xor XOR2 (N3799, N3796, N1133);
nor NOR4 (N3800, N3785, N1910, N171, N599);
not NOT1 (N3801, N3773);
nand NAND3 (N3802, N3791, N840, N737);
or OR2 (N3803, N3802, N2027);
buf BUF1 (N3804, N3798);
buf BUF1 (N3805, N3760);
and AND3 (N3806, N3795, N3171, N551);
xor XOR2 (N3807, N3803, N1615);
or OR2 (N3808, N3805, N2681);
buf BUF1 (N3809, N3806);
nor NOR3 (N3810, N3801, N1254, N3656);
not NOT1 (N3811, N3799);
or OR4 (N3812, N3797, N3484, N1522, N1578);
nor NOR3 (N3813, N3811, N664, N1753);
nor NOR4 (N3814, N3812, N2194, N3430, N3254);
buf BUF1 (N3815, N3775);
not NOT1 (N3816, N3794);
buf BUF1 (N3817, N3813);
or OR2 (N3818, N3808, N1411);
xor XOR2 (N3819, N3800, N862);
not NOT1 (N3820, N3816);
nor NOR4 (N3821, N3809, N1947, N2283, N3819);
nor NOR2 (N3822, N3467, N1980);
nor NOR3 (N3823, N3818, N2100, N42);
nand NAND3 (N3824, N3820, N987, N2425);
or OR4 (N3825, N3810, N3434, N3040, N2514);
or OR3 (N3826, N3807, N3539, N532);
xor XOR2 (N3827, N3814, N848);
or OR4 (N3828, N3825, N3656, N3750, N3094);
and AND4 (N3829, N3826, N2546, N3282, N357);
buf BUF1 (N3830, N3821);
xor XOR2 (N3831, N3815, N52);
buf BUF1 (N3832, N3830);
and AND2 (N3833, N3822, N2259);
nor NOR3 (N3834, N3823, N3757, N1678);
nor NOR3 (N3835, N3829, N64, N1314);
nor NOR3 (N3836, N3834, N520, N3773);
or OR4 (N3837, N3832, N1153, N3835, N1355);
nor NOR2 (N3838, N3792, N1182);
xor XOR2 (N3839, N3831, N1108);
and AND2 (N3840, N3817, N1463);
nor NOR2 (N3841, N3827, N1343);
buf BUF1 (N3842, N3840);
nand NAND4 (N3843, N3841, N2271, N891, N3117);
nand NAND2 (N3844, N3824, N2018);
nand NAND3 (N3845, N3836, N150, N700);
and AND3 (N3846, N3839, N3004, N3181);
xor XOR2 (N3847, N3842, N583);
buf BUF1 (N3848, N3833);
buf BUF1 (N3849, N3837);
nand NAND3 (N3850, N3848, N2691, N2129);
nor NOR2 (N3851, N3843, N1525);
not NOT1 (N3852, N3804);
not NOT1 (N3853, N3849);
xor XOR2 (N3854, N3838, N2470);
not NOT1 (N3855, N3851);
nand NAND3 (N3856, N3852, N1211, N1392);
nand NAND2 (N3857, N3846, N989);
not NOT1 (N3858, N3844);
or OR3 (N3859, N3850, N3802, N3114);
or OR2 (N3860, N3854, N199);
nand NAND2 (N3861, N3847, N571);
buf BUF1 (N3862, N3845);
and AND3 (N3863, N3858, N200, N3459);
buf BUF1 (N3864, N3857);
or OR3 (N3865, N3859, N447, N2021);
or OR4 (N3866, N3865, N2081, N2580, N104);
nand NAND2 (N3867, N3860, N3081);
not NOT1 (N3868, N3863);
and AND4 (N3869, N3853, N473, N3281, N1717);
not NOT1 (N3870, N3867);
nor NOR3 (N3871, N3856, N2850, N338);
buf BUF1 (N3872, N3866);
xor XOR2 (N3873, N3862, N3859);
or OR2 (N3874, N3864, N1929);
xor XOR2 (N3875, N3855, N3199);
nor NOR2 (N3876, N3875, N2567);
nor NOR3 (N3877, N3869, N3415, N2626);
buf BUF1 (N3878, N3874);
xor XOR2 (N3879, N3876, N9);
nand NAND2 (N3880, N3868, N1507);
and AND4 (N3881, N3873, N1446, N944, N1725);
nor NOR4 (N3882, N3871, N920, N757, N1482);
and AND2 (N3883, N3879, N1066);
not NOT1 (N3884, N3878);
xor XOR2 (N3885, N3872, N1945);
nor NOR2 (N3886, N3884, N2890);
or OR4 (N3887, N3870, N537, N1358, N161);
or OR3 (N3888, N3881, N2167, N1147);
buf BUF1 (N3889, N3882);
and AND2 (N3890, N3877, N3141);
nor NOR3 (N3891, N3890, N3849, N959);
buf BUF1 (N3892, N3828);
buf BUF1 (N3893, N3883);
buf BUF1 (N3894, N3888);
and AND4 (N3895, N3891, N1894, N1439, N2219);
or OR2 (N3896, N3893, N3722);
not NOT1 (N3897, N3892);
or OR3 (N3898, N3889, N322, N3585);
nand NAND3 (N3899, N3896, N1729, N1101);
xor XOR2 (N3900, N3885, N3263);
nor NOR3 (N3901, N3861, N928, N1506);
nor NOR2 (N3902, N3895, N2360);
buf BUF1 (N3903, N3898);
or OR4 (N3904, N3901, N3133, N3594, N1207);
and AND3 (N3905, N3897, N1753, N2224);
xor XOR2 (N3906, N3904, N3719);
and AND4 (N3907, N3887, N3096, N1887, N2894);
and AND2 (N3908, N3899, N1935);
not NOT1 (N3909, N3905);
nor NOR2 (N3910, N3880, N2501);
not NOT1 (N3911, N3886);
buf BUF1 (N3912, N3894);
and AND4 (N3913, N3903, N2260, N2985, N2407);
or OR3 (N3914, N3910, N877, N1072);
or OR3 (N3915, N3909, N2868, N2230);
or OR4 (N3916, N3902, N953, N1915, N1053);
not NOT1 (N3917, N3912);
nand NAND3 (N3918, N3907, N2595, N1824);
or OR3 (N3919, N3918, N33, N2326);
buf BUF1 (N3920, N3916);
nor NOR2 (N3921, N3914, N1576);
not NOT1 (N3922, N3908);
and AND3 (N3923, N3915, N2963, N3298);
nor NOR4 (N3924, N3913, N3262, N328, N3283);
and AND4 (N3925, N3900, N307, N2217, N205);
nand NAND4 (N3926, N3925, N1140, N2138, N2555);
or OR4 (N3927, N3923, N302, N2644, N2497);
not NOT1 (N3928, N3921);
xor XOR2 (N3929, N3926, N721);
or OR2 (N3930, N3920, N3682);
buf BUF1 (N3931, N3929);
buf BUF1 (N3932, N3927);
not NOT1 (N3933, N3931);
and AND3 (N3934, N3924, N632, N1446);
xor XOR2 (N3935, N3906, N2148);
not NOT1 (N3936, N3922);
not NOT1 (N3937, N3934);
nor NOR4 (N3938, N3936, N2358, N3286, N3008);
and AND3 (N3939, N3928, N2439, N2938);
nor NOR2 (N3940, N3917, N1778);
nor NOR3 (N3941, N3940, N3685, N1207);
buf BUF1 (N3942, N3911);
xor XOR2 (N3943, N3938, N2190);
or OR3 (N3944, N3919, N2953, N730);
nand NAND2 (N3945, N3935, N3185);
and AND3 (N3946, N3939, N2881, N1708);
and AND3 (N3947, N3942, N1935, N1713);
buf BUF1 (N3948, N3930);
nand NAND3 (N3949, N3945, N1883, N3340);
not NOT1 (N3950, N3946);
nor NOR2 (N3951, N3949, N1602);
and AND2 (N3952, N3937, N3621);
or OR2 (N3953, N3941, N3401);
nand NAND3 (N3954, N3932, N1196, N388);
not NOT1 (N3955, N3953);
not NOT1 (N3956, N3950);
or OR3 (N3957, N3947, N898, N3513);
nand NAND3 (N3958, N3956, N227, N219);
or OR3 (N3959, N3933, N3855, N826);
nand NAND4 (N3960, N3954, N1723, N1575, N3205);
or OR3 (N3961, N3959, N795, N3488);
xor XOR2 (N3962, N3958, N163);
not NOT1 (N3963, N3960);
xor XOR2 (N3964, N3951, N3381);
not NOT1 (N3965, N3962);
or OR3 (N3966, N3948, N1301, N108);
and AND3 (N3967, N3966, N1763, N1940);
xor XOR2 (N3968, N3964, N3847);
nor NOR4 (N3969, N3955, N2190, N3735, N1621);
not NOT1 (N3970, N3968);
and AND3 (N3971, N3952, N188, N403);
not NOT1 (N3972, N3965);
nor NOR4 (N3973, N3969, N2793, N3330, N3090);
xor XOR2 (N3974, N3961, N1661);
not NOT1 (N3975, N3967);
and AND2 (N3976, N3972, N1273);
or OR3 (N3977, N3944, N570, N3231);
nor NOR4 (N3978, N3976, N2783, N3809, N406);
nand NAND4 (N3979, N3978, N2131, N1714, N1198);
nor NOR3 (N3980, N3977, N3764, N2128);
xor XOR2 (N3981, N3975, N876);
and AND4 (N3982, N3970, N3400, N2413, N2585);
not NOT1 (N3983, N3982);
nand NAND2 (N3984, N3980, N1788);
not NOT1 (N3985, N3973);
xor XOR2 (N3986, N3984, N3694);
nor NOR2 (N3987, N3957, N2472);
and AND2 (N3988, N3983, N3699);
xor XOR2 (N3989, N3974, N1120);
not NOT1 (N3990, N3985);
not NOT1 (N3991, N3979);
nor NOR2 (N3992, N3986, N23);
nand NAND3 (N3993, N3963, N3273, N3616);
buf BUF1 (N3994, N3989);
nand NAND2 (N3995, N3992, N3697);
buf BUF1 (N3996, N3943);
and AND2 (N3997, N3987, N864);
xor XOR2 (N3998, N3997, N3022);
and AND3 (N3999, N3995, N2657, N2842);
not NOT1 (N4000, N3994);
xor XOR2 (N4001, N3971, N39);
or OR2 (N4002, N4000, N1179);
nor NOR4 (N4003, N3993, N2558, N3288, N3072);
not NOT1 (N4004, N3990);
buf BUF1 (N4005, N4002);
and AND4 (N4006, N4005, N1929, N575, N315);
not NOT1 (N4007, N3988);
buf BUF1 (N4008, N3991);
and AND4 (N4009, N4003, N1861, N3475, N3554);
buf BUF1 (N4010, N3996);
not NOT1 (N4011, N4004);
not NOT1 (N4012, N4006);
not NOT1 (N4013, N4008);
nor NOR4 (N4014, N3999, N1692, N1128, N3608);
not NOT1 (N4015, N3998);
endmodule