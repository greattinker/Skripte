// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;

output N909,N913,N908,N917,N915,N910,N911,N916,N914,N918;

nor NOR3 (N19, N7, N11, N9);
not NOT1 (N20, N12);
and AND2 (N21, N19, N17);
nand NAND2 (N22, N9, N11);
xor XOR2 (N23, N2, N18);
buf BUF1 (N24, N5);
buf BUF1 (N25, N10);
xor XOR2 (N26, N20, N10);
buf BUF1 (N27, N14);
xor XOR2 (N28, N4, N4);
nor NOR3 (N29, N1, N6, N2);
buf BUF1 (N30, N19);
xor XOR2 (N31, N29, N16);
not NOT1 (N32, N26);
buf BUF1 (N33, N27);
and AND4 (N34, N22, N6, N27, N3);
and AND4 (N35, N28, N30, N4, N18);
xor XOR2 (N36, N14, N20);
and AND3 (N37, N33, N22, N35);
buf BUF1 (N38, N31);
buf BUF1 (N39, N34);
nand NAND2 (N40, N21, N37);
nand NAND4 (N41, N13, N30, N4, N38);
and AND4 (N42, N10, N39, N39, N5);
buf BUF1 (N43, N38);
not NOT1 (N44, N1);
buf BUF1 (N45, N24);
not NOT1 (N46, N32);
not NOT1 (N47, N43);
buf BUF1 (N48, N47);
xor XOR2 (N49, N40, N1);
or OR3 (N50, N46, N40, N42);
nor NOR2 (N51, N47, N26);
not NOT1 (N52, N23);
nand NAND3 (N53, N41, N32, N48);
or OR2 (N54, N47, N38);
nand NAND4 (N55, N53, N7, N34, N28);
buf BUF1 (N56, N54);
or OR2 (N57, N56, N13);
not NOT1 (N58, N50);
xor XOR2 (N59, N51, N52);
nand NAND4 (N60, N22, N29, N10, N55);
nand NAND4 (N61, N56, N26, N15, N27);
not NOT1 (N62, N59);
buf BUF1 (N63, N25);
xor XOR2 (N64, N36, N10);
nand NAND2 (N65, N60, N13);
buf BUF1 (N66, N63);
buf BUF1 (N67, N62);
nor NOR2 (N68, N61, N10);
nor NOR2 (N69, N45, N3);
and AND4 (N70, N67, N16, N22, N60);
xor XOR2 (N71, N57, N10);
and AND4 (N72, N44, N10, N17, N8);
or OR3 (N73, N66, N10, N38);
and AND2 (N74, N71, N55);
nor NOR2 (N75, N49, N58);
and AND2 (N76, N69, N25);
not NOT1 (N77, N13);
or OR2 (N78, N73, N50);
buf BUF1 (N79, N72);
xor XOR2 (N80, N77, N58);
or OR2 (N81, N74, N9);
nor NOR2 (N82, N75, N37);
and AND4 (N83, N64, N21, N19, N69);
buf BUF1 (N84, N68);
not NOT1 (N85, N79);
and AND4 (N86, N65, N56, N17, N85);
nor NOR2 (N87, N37, N86);
nor NOR2 (N88, N80, N43);
nor NOR2 (N89, N9, N2);
nor NOR3 (N90, N76, N84, N40);
not NOT1 (N91, N70);
nand NAND4 (N92, N4, N20, N85, N10);
not NOT1 (N93, N83);
not NOT1 (N94, N87);
xor XOR2 (N95, N92, N83);
or OR4 (N96, N94, N29, N40, N14);
nor NOR3 (N97, N81, N30, N46);
nor NOR4 (N98, N96, N64, N47, N62);
buf BUF1 (N99, N98);
and AND4 (N100, N82, N38, N57, N2);
buf BUF1 (N101, N99);
nand NAND2 (N102, N101, N57);
nand NAND4 (N103, N95, N98, N62, N76);
not NOT1 (N104, N91);
nand NAND3 (N105, N97, N9, N90);
buf BUF1 (N106, N17);
and AND3 (N107, N103, N58, N50);
nand NAND4 (N108, N89, N87, N2, N99);
nand NAND3 (N109, N100, N5, N97);
or OR3 (N110, N102, N65, N32);
nand NAND3 (N111, N106, N86, N29);
not NOT1 (N112, N110);
nand NAND2 (N113, N105, N12);
and AND2 (N114, N78, N82);
not NOT1 (N115, N108);
or OR2 (N116, N107, N80);
nand NAND4 (N117, N115, N77, N71, N76);
nand NAND2 (N118, N114, N73);
xor XOR2 (N119, N111, N3);
nand NAND3 (N120, N116, N38, N71);
xor XOR2 (N121, N113, N43);
and AND4 (N122, N93, N34, N110, N94);
not NOT1 (N123, N118);
buf BUF1 (N124, N120);
and AND3 (N125, N117, N13, N16);
buf BUF1 (N126, N121);
not NOT1 (N127, N112);
nand NAND2 (N128, N126, N43);
buf BUF1 (N129, N88);
buf BUF1 (N130, N127);
nand NAND2 (N131, N122, N2);
buf BUF1 (N132, N104);
nand NAND4 (N133, N123, N11, N97, N20);
buf BUF1 (N134, N129);
not NOT1 (N135, N130);
nor NOR4 (N136, N119, N59, N62, N99);
xor XOR2 (N137, N132, N96);
and AND3 (N138, N133, N86, N6);
nand NAND3 (N139, N138, N111, N110);
xor XOR2 (N140, N109, N27);
not NOT1 (N141, N134);
not NOT1 (N142, N137);
buf BUF1 (N143, N125);
nor NOR4 (N144, N136, N39, N95, N49);
nand NAND2 (N145, N124, N30);
xor XOR2 (N146, N135, N114);
xor XOR2 (N147, N146, N15);
and AND2 (N148, N144, N37);
nand NAND4 (N149, N140, N135, N110, N35);
buf BUF1 (N150, N143);
nand NAND4 (N151, N145, N76, N119, N37);
or OR3 (N152, N142, N30, N142);
and AND2 (N153, N151, N141);
nor NOR4 (N154, N11, N90, N67, N29);
xor XOR2 (N155, N153, N38);
buf BUF1 (N156, N147);
or OR4 (N157, N150, N15, N12, N36);
nand NAND3 (N158, N154, N144, N25);
not NOT1 (N159, N128);
nand NAND4 (N160, N159, N107, N121, N153);
xor XOR2 (N161, N131, N135);
and AND3 (N162, N149, N11, N68);
nor NOR3 (N163, N139, N27, N118);
or OR3 (N164, N163, N68, N73);
buf BUF1 (N165, N161);
xor XOR2 (N166, N152, N15);
or OR2 (N167, N162, N69);
nor NOR4 (N168, N165, N160, N79, N128);
buf BUF1 (N169, N69);
buf BUF1 (N170, N156);
xor XOR2 (N171, N166, N79);
nand NAND2 (N172, N169, N49);
xor XOR2 (N173, N148, N78);
nand NAND4 (N174, N164, N164, N157, N28);
not NOT1 (N175, N171);
xor XOR2 (N176, N23, N66);
xor XOR2 (N177, N176, N103);
not NOT1 (N178, N155);
xor XOR2 (N179, N167, N178);
nor NOR2 (N180, N135, N4);
and AND2 (N181, N179, N62);
nand NAND4 (N182, N175, N105, N152, N4);
buf BUF1 (N183, N174);
nor NOR3 (N184, N182, N19, N106);
nand NAND2 (N185, N183, N123);
nor NOR3 (N186, N173, N1, N12);
not NOT1 (N187, N172);
nor NOR2 (N188, N170, N54);
or OR4 (N189, N187, N178, N60, N182);
nor NOR3 (N190, N158, N95, N88);
buf BUF1 (N191, N185);
not NOT1 (N192, N189);
nor NOR4 (N193, N181, N159, N132, N65);
nand NAND3 (N194, N184, N165, N44);
nor NOR4 (N195, N168, N2, N130, N63);
buf BUF1 (N196, N186);
buf BUF1 (N197, N190);
and AND4 (N198, N195, N92, N114, N41);
or OR2 (N199, N197, N79);
buf BUF1 (N200, N196);
or OR4 (N201, N198, N121, N69, N27);
nor NOR3 (N202, N193, N29, N66);
nand NAND3 (N203, N188, N108, N43);
xor XOR2 (N204, N201, N71);
and AND4 (N205, N192, N144, N108, N61);
not NOT1 (N206, N204);
or OR2 (N207, N191, N130);
xor XOR2 (N208, N202, N70);
not NOT1 (N209, N206);
buf BUF1 (N210, N200);
or OR4 (N211, N199, N116, N130, N76);
xor XOR2 (N212, N194, N149);
and AND2 (N213, N208, N145);
and AND2 (N214, N210, N201);
nand NAND3 (N215, N177, N149, N92);
or OR3 (N216, N203, N26, N176);
or OR2 (N217, N214, N76);
not NOT1 (N218, N205);
nor NOR4 (N219, N218, N82, N164, N206);
not NOT1 (N220, N207);
or OR2 (N221, N215, N127);
nand NAND4 (N222, N221, N15, N33, N153);
nand NAND2 (N223, N217, N118);
buf BUF1 (N224, N216);
and AND2 (N225, N180, N85);
not NOT1 (N226, N212);
and AND2 (N227, N219, N212);
nand NAND3 (N228, N226, N137, N128);
xor XOR2 (N229, N222, N199);
xor XOR2 (N230, N228, N204);
not NOT1 (N231, N220);
or OR4 (N232, N230, N141, N38, N56);
or OR3 (N233, N229, N108, N142);
nand NAND2 (N234, N223, N43);
nand NAND2 (N235, N213, N53);
xor XOR2 (N236, N233, N101);
xor XOR2 (N237, N234, N118);
or OR3 (N238, N232, N229, N205);
nor NOR3 (N239, N231, N116, N151);
and AND4 (N240, N237, N152, N186, N2);
buf BUF1 (N241, N235);
xor XOR2 (N242, N227, N25);
or OR3 (N243, N238, N153, N125);
buf BUF1 (N244, N239);
xor XOR2 (N245, N209, N211);
and AND2 (N246, N146, N74);
buf BUF1 (N247, N242);
nor NOR3 (N248, N244, N214, N107);
nand NAND2 (N249, N241, N29);
nand NAND3 (N250, N245, N179, N2);
or OR4 (N251, N240, N145, N160, N216);
and AND3 (N252, N224, N84, N18);
and AND4 (N253, N246, N224, N79, N16);
or OR2 (N254, N249, N63);
nand NAND3 (N255, N251, N84, N38);
xor XOR2 (N256, N248, N198);
nand NAND3 (N257, N254, N233, N145);
and AND2 (N258, N253, N161);
not NOT1 (N259, N258);
not NOT1 (N260, N257);
nand NAND3 (N261, N259, N189, N27);
nand NAND2 (N262, N261, N182);
not NOT1 (N263, N252);
and AND3 (N264, N263, N221, N145);
buf BUF1 (N265, N236);
buf BUF1 (N266, N260);
or OR2 (N267, N262, N247);
and AND4 (N268, N227, N20, N53, N59);
not NOT1 (N269, N267);
nor NOR2 (N270, N269, N105);
and AND4 (N271, N264, N91, N140, N36);
not NOT1 (N272, N256);
and AND4 (N273, N243, N149, N66, N72);
nand NAND4 (N274, N270, N21, N127, N66);
buf BUF1 (N275, N273);
nor NOR3 (N276, N250, N3, N20);
nor NOR3 (N277, N255, N66, N2);
and AND4 (N278, N275, N208, N263, N29);
or OR2 (N279, N225, N180);
or OR2 (N280, N276, N196);
and AND4 (N281, N277, N76, N83, N116);
or OR3 (N282, N280, N106, N142);
or OR4 (N283, N272, N234, N149, N93);
not NOT1 (N284, N282);
nand NAND3 (N285, N268, N232, N141);
nor NOR2 (N286, N284, N4);
not NOT1 (N287, N266);
nor NOR2 (N288, N287, N80);
nor NOR4 (N289, N274, N239, N84, N202);
not NOT1 (N290, N279);
and AND4 (N291, N265, N234, N174, N255);
nand NAND2 (N292, N283, N6);
not NOT1 (N293, N271);
and AND2 (N294, N288, N79);
nor NOR3 (N295, N286, N155, N35);
buf BUF1 (N296, N281);
nand NAND3 (N297, N293, N166, N51);
xor XOR2 (N298, N295, N289);
xor XOR2 (N299, N84, N156);
xor XOR2 (N300, N299, N80);
nor NOR2 (N301, N278, N169);
xor XOR2 (N302, N291, N217);
nand NAND4 (N303, N296, N70, N197, N219);
or OR2 (N304, N292, N293);
and AND4 (N305, N304, N152, N170, N291);
not NOT1 (N306, N302);
nand NAND3 (N307, N290, N220, N301);
not NOT1 (N308, N245);
xor XOR2 (N309, N298, N300);
buf BUF1 (N310, N246);
xor XOR2 (N311, N285, N243);
buf BUF1 (N312, N309);
buf BUF1 (N313, N306);
buf BUF1 (N314, N312);
or OR3 (N315, N310, N29, N26);
or OR3 (N316, N294, N213, N303);
nand NAND2 (N317, N172, N293);
buf BUF1 (N318, N316);
nor NOR4 (N319, N318, N93, N166, N204);
buf BUF1 (N320, N308);
and AND2 (N321, N307, N129);
xor XOR2 (N322, N320, N148);
nand NAND4 (N323, N317, N240, N287, N77);
not NOT1 (N324, N311);
and AND2 (N325, N305, N139);
and AND2 (N326, N313, N53);
or OR3 (N327, N319, N49, N1);
or OR2 (N328, N323, N286);
not NOT1 (N329, N328);
buf BUF1 (N330, N326);
nand NAND2 (N331, N329, N193);
nor NOR2 (N332, N314, N170);
or OR4 (N333, N325, N303, N141, N104);
buf BUF1 (N334, N315);
and AND2 (N335, N330, N293);
not NOT1 (N336, N297);
or OR4 (N337, N335, N12, N73, N331);
and AND2 (N338, N321, N195);
nor NOR3 (N339, N181, N147, N22);
nand NAND3 (N340, N334, N213, N164);
nand NAND4 (N341, N327, N118, N220, N261);
and AND3 (N342, N333, N33, N240);
xor XOR2 (N343, N339, N160);
not NOT1 (N344, N336);
not NOT1 (N345, N322);
or OR3 (N346, N342, N190, N100);
or OR4 (N347, N324, N55, N134, N185);
nor NOR4 (N348, N343, N150, N282, N209);
or OR2 (N349, N347, N45);
not NOT1 (N350, N338);
nor NOR2 (N351, N348, N292);
and AND3 (N352, N340, N340, N126);
nand NAND3 (N353, N344, N253, N202);
nand NAND2 (N354, N346, N110);
nand NAND3 (N355, N341, N15, N258);
xor XOR2 (N356, N354, N350);
or OR3 (N357, N226, N165, N193);
buf BUF1 (N358, N353);
nor NOR2 (N359, N351, N156);
or OR4 (N360, N337, N227, N59, N2);
and AND2 (N361, N358, N65);
buf BUF1 (N362, N361);
nand NAND3 (N363, N332, N196, N175);
xor XOR2 (N364, N360, N180);
and AND4 (N365, N362, N353, N49, N187);
or OR3 (N366, N345, N247, N124);
and AND4 (N367, N364, N37, N65, N352);
xor XOR2 (N368, N211, N232);
nor NOR4 (N369, N366, N101, N199, N145);
not NOT1 (N370, N365);
buf BUF1 (N371, N363);
nand NAND2 (N372, N371, N229);
not NOT1 (N373, N367);
nand NAND2 (N374, N370, N338);
buf BUF1 (N375, N357);
xor XOR2 (N376, N368, N47);
not NOT1 (N377, N374);
xor XOR2 (N378, N373, N43);
xor XOR2 (N379, N377, N365);
not NOT1 (N380, N372);
and AND2 (N381, N359, N42);
not NOT1 (N382, N380);
not NOT1 (N383, N375);
not NOT1 (N384, N383);
nor NOR3 (N385, N376, N290, N247);
xor XOR2 (N386, N349, N136);
xor XOR2 (N387, N385, N45);
nand NAND3 (N388, N384, N89, N63);
xor XOR2 (N389, N378, N95);
or OR4 (N390, N369, N219, N255, N52);
and AND4 (N391, N388, N332, N73, N232);
not NOT1 (N392, N381);
and AND3 (N393, N356, N134, N108);
nor NOR4 (N394, N382, N39, N231, N103);
xor XOR2 (N395, N355, N16);
not NOT1 (N396, N379);
xor XOR2 (N397, N391, N138);
nor NOR4 (N398, N390, N105, N270, N301);
or OR2 (N399, N396, N201);
not NOT1 (N400, N397);
or OR2 (N401, N394, N356);
nand NAND4 (N402, N393, N107, N378, N388);
or OR2 (N403, N400, N299);
buf BUF1 (N404, N398);
xor XOR2 (N405, N402, N8);
and AND2 (N406, N386, N365);
nor NOR2 (N407, N395, N177);
nand NAND3 (N408, N401, N247, N192);
nand NAND4 (N409, N407, N76, N154, N364);
and AND4 (N410, N403, N186, N310, N205);
nand NAND3 (N411, N410, N312, N187);
buf BUF1 (N412, N406);
nor NOR4 (N413, N412, N195, N5, N311);
and AND3 (N414, N409, N94, N59);
not NOT1 (N415, N405);
xor XOR2 (N416, N404, N16);
nand NAND4 (N417, N392, N379, N122, N242);
and AND2 (N418, N416, N119);
buf BUF1 (N419, N417);
or OR3 (N420, N413, N46, N408);
not NOT1 (N421, N347);
buf BUF1 (N422, N387);
xor XOR2 (N423, N422, N205);
or OR3 (N424, N418, N274, N321);
nor NOR2 (N425, N420, N234);
or OR4 (N426, N414, N12, N421, N103);
nand NAND3 (N427, N244, N354, N200);
nor NOR4 (N428, N389, N379, N75, N386);
or OR2 (N429, N425, N59);
xor XOR2 (N430, N424, N380);
and AND3 (N431, N427, N39, N422);
and AND2 (N432, N426, N106);
nand NAND3 (N433, N431, N315, N158);
not NOT1 (N434, N433);
xor XOR2 (N435, N411, N31);
not NOT1 (N436, N430);
nor NOR3 (N437, N428, N341, N98);
nand NAND3 (N438, N429, N344, N331);
nor NOR3 (N439, N432, N281, N169);
xor XOR2 (N440, N438, N337);
nor NOR4 (N441, N439, N273, N80, N410);
xor XOR2 (N442, N440, N124);
xor XOR2 (N443, N437, N432);
xor XOR2 (N444, N399, N115);
and AND2 (N445, N434, N147);
nor NOR4 (N446, N441, N412, N144, N441);
nor NOR2 (N447, N443, N6);
nand NAND3 (N448, N423, N406, N235);
or OR2 (N449, N446, N312);
xor XOR2 (N450, N435, N443);
nor NOR4 (N451, N442, N38, N264, N315);
not NOT1 (N452, N447);
and AND3 (N453, N436, N230, N369);
xor XOR2 (N454, N453, N3);
or OR4 (N455, N419, N179, N244, N204);
and AND4 (N456, N452, N197, N60, N160);
xor XOR2 (N457, N415, N403);
not NOT1 (N458, N448);
xor XOR2 (N459, N444, N183);
and AND4 (N460, N451, N169, N280, N384);
not NOT1 (N461, N456);
and AND3 (N462, N457, N6, N397);
nor NOR2 (N463, N450, N47);
not NOT1 (N464, N449);
nand NAND2 (N465, N454, N459);
and AND3 (N466, N28, N122, N415);
nand NAND3 (N467, N458, N374, N27);
not NOT1 (N468, N455);
or OR2 (N469, N460, N456);
and AND2 (N470, N465, N419);
xor XOR2 (N471, N461, N21);
nor NOR4 (N472, N470, N378, N150, N170);
and AND4 (N473, N464, N358, N276, N48);
not NOT1 (N474, N473);
or OR3 (N475, N466, N28, N207);
or OR3 (N476, N445, N31, N308);
and AND3 (N477, N469, N356, N34);
xor XOR2 (N478, N462, N41);
xor XOR2 (N479, N463, N380);
and AND2 (N480, N478, N389);
not NOT1 (N481, N472);
nor NOR3 (N482, N468, N131, N414);
not NOT1 (N483, N482);
not NOT1 (N484, N476);
buf BUF1 (N485, N477);
buf BUF1 (N486, N474);
or OR4 (N487, N467, N256, N22, N312);
nor NOR2 (N488, N475, N151);
xor XOR2 (N489, N484, N128);
and AND2 (N490, N471, N30);
nor NOR3 (N491, N485, N140, N26);
not NOT1 (N492, N488);
or OR2 (N493, N486, N139);
not NOT1 (N494, N487);
and AND4 (N495, N492, N31, N423, N47);
not NOT1 (N496, N494);
or OR2 (N497, N483, N298);
not NOT1 (N498, N495);
not NOT1 (N499, N479);
and AND2 (N500, N481, N409);
xor XOR2 (N501, N490, N324);
nand NAND3 (N502, N498, N221, N441);
nand NAND4 (N503, N496, N401, N92, N38);
buf BUF1 (N504, N497);
not NOT1 (N505, N501);
or OR3 (N506, N503, N198, N293);
nor NOR4 (N507, N480, N390, N482, N271);
not NOT1 (N508, N505);
buf BUF1 (N509, N504);
nand NAND2 (N510, N499, N470);
nand NAND4 (N511, N500, N276, N105, N105);
nand NAND2 (N512, N510, N426);
and AND3 (N513, N493, N396, N24);
not NOT1 (N514, N508);
not NOT1 (N515, N511);
and AND2 (N516, N515, N159);
not NOT1 (N517, N509);
not NOT1 (N518, N516);
nor NOR2 (N519, N514, N8);
xor XOR2 (N520, N519, N63);
buf BUF1 (N521, N491);
and AND2 (N522, N507, N201);
or OR4 (N523, N512, N226, N341, N254);
nor NOR3 (N524, N523, N340, N445);
nor NOR3 (N525, N506, N13, N120);
or OR4 (N526, N517, N282, N211, N112);
nand NAND2 (N527, N525, N161);
nor NOR2 (N528, N489, N399);
xor XOR2 (N529, N518, N488);
and AND2 (N530, N522, N443);
nor NOR3 (N531, N502, N152, N340);
and AND3 (N532, N513, N425, N253);
xor XOR2 (N533, N524, N258);
or OR2 (N534, N521, N98);
buf BUF1 (N535, N531);
nor NOR3 (N536, N533, N134, N451);
or OR2 (N537, N520, N524);
nand NAND2 (N538, N529, N203);
and AND2 (N539, N527, N372);
nand NAND3 (N540, N537, N65, N148);
or OR4 (N541, N538, N243, N462, N458);
buf BUF1 (N542, N526);
or OR4 (N543, N535, N341, N51, N469);
or OR3 (N544, N536, N34, N540);
xor XOR2 (N545, N519, N340);
not NOT1 (N546, N530);
nand NAND4 (N547, N539, N465, N344, N507);
not NOT1 (N548, N547);
not NOT1 (N549, N546);
buf BUF1 (N550, N544);
nor NOR4 (N551, N541, N354, N181, N184);
buf BUF1 (N552, N542);
or OR3 (N553, N543, N46, N331);
xor XOR2 (N554, N551, N196);
nor NOR4 (N555, N545, N258, N24, N493);
not NOT1 (N556, N555);
nand NAND2 (N557, N534, N379);
buf BUF1 (N558, N553);
xor XOR2 (N559, N558, N428);
not NOT1 (N560, N532);
nand NAND3 (N561, N557, N538, N215);
buf BUF1 (N562, N550);
nor NOR3 (N563, N560, N177, N26);
nand NAND2 (N564, N549, N177);
or OR4 (N565, N564, N354, N248, N518);
not NOT1 (N566, N528);
not NOT1 (N567, N562);
buf BUF1 (N568, N565);
xor XOR2 (N569, N552, N496);
nand NAND3 (N570, N559, N287, N406);
nor NOR3 (N571, N563, N11, N470);
not NOT1 (N572, N561);
xor XOR2 (N573, N571, N3);
not NOT1 (N574, N569);
and AND3 (N575, N568, N574, N225);
not NOT1 (N576, N457);
nand NAND4 (N577, N554, N130, N117, N18);
not NOT1 (N578, N556);
xor XOR2 (N579, N576, N38);
nand NAND4 (N580, N577, N145, N132, N424);
nand NAND2 (N581, N578, N119);
nor NOR3 (N582, N572, N522, N291);
nor NOR3 (N583, N581, N226, N124);
xor XOR2 (N584, N582, N294);
nand NAND4 (N585, N573, N491, N154, N292);
or OR3 (N586, N579, N312, N422);
nand NAND2 (N587, N583, N112);
or OR4 (N588, N570, N37, N344, N574);
xor XOR2 (N589, N548, N470);
nand NAND2 (N590, N567, N520);
buf BUF1 (N591, N588);
xor XOR2 (N592, N590, N169);
not NOT1 (N593, N584);
xor XOR2 (N594, N593, N171);
xor XOR2 (N595, N594, N36);
or OR4 (N596, N592, N77, N36, N289);
not NOT1 (N597, N575);
and AND2 (N598, N585, N412);
or OR3 (N599, N591, N431, N180);
not NOT1 (N600, N580);
buf BUF1 (N601, N586);
xor XOR2 (N602, N596, N88);
nor NOR2 (N603, N597, N27);
buf BUF1 (N604, N599);
nand NAND3 (N605, N595, N306, N567);
nand NAND2 (N606, N604, N79);
nor NOR4 (N607, N605, N242, N417, N85);
nand NAND4 (N608, N603, N58, N568, N26);
not NOT1 (N609, N601);
nor NOR2 (N610, N602, N559);
and AND3 (N611, N600, N236, N12);
or OR3 (N612, N606, N260, N228);
nand NAND2 (N613, N611, N100);
or OR2 (N614, N598, N16);
nand NAND4 (N615, N613, N494, N509, N81);
buf BUF1 (N616, N607);
nand NAND2 (N617, N610, N409);
not NOT1 (N618, N616);
buf BUF1 (N619, N617);
buf BUF1 (N620, N608);
buf BUF1 (N621, N615);
and AND3 (N622, N609, N203, N246);
nor NOR4 (N623, N612, N530, N483, N10);
or OR3 (N624, N620, N490, N300);
and AND4 (N625, N621, N67, N265, N143);
or OR3 (N626, N589, N499, N542);
not NOT1 (N627, N566);
not NOT1 (N628, N618);
nand NAND4 (N629, N614, N85, N425, N228);
nor NOR3 (N630, N622, N451, N82);
or OR3 (N631, N628, N122, N363);
and AND3 (N632, N630, N232, N264);
and AND4 (N633, N631, N563, N469, N149);
not NOT1 (N634, N624);
or OR2 (N635, N587, N349);
xor XOR2 (N636, N635, N452);
nand NAND3 (N637, N632, N535, N594);
xor XOR2 (N638, N625, N56);
not NOT1 (N639, N637);
nand NAND4 (N640, N633, N63, N398, N238);
nand NAND3 (N641, N623, N638, N528);
xor XOR2 (N642, N381, N311);
xor XOR2 (N643, N640, N394);
not NOT1 (N644, N627);
xor XOR2 (N645, N639, N603);
nor NOR3 (N646, N634, N544, N179);
buf BUF1 (N647, N626);
nor NOR4 (N648, N642, N410, N513, N594);
nor NOR2 (N649, N645, N294);
nand NAND3 (N650, N641, N49, N263);
not NOT1 (N651, N650);
buf BUF1 (N652, N629);
and AND2 (N653, N644, N196);
buf BUF1 (N654, N647);
and AND3 (N655, N648, N195, N152);
not NOT1 (N656, N652);
xor XOR2 (N657, N656, N115);
nand NAND2 (N658, N655, N467);
buf BUF1 (N659, N643);
or OR2 (N660, N654, N174);
not NOT1 (N661, N659);
buf BUF1 (N662, N646);
not NOT1 (N663, N653);
nand NAND2 (N664, N660, N201);
nand NAND3 (N665, N661, N93, N501);
xor XOR2 (N666, N636, N374);
nand NAND4 (N667, N657, N623, N370, N321);
nor NOR2 (N668, N662, N549);
xor XOR2 (N669, N666, N106);
xor XOR2 (N670, N667, N385);
not NOT1 (N671, N619);
not NOT1 (N672, N665);
or OR3 (N673, N668, N275, N53);
xor XOR2 (N674, N669, N239);
nand NAND4 (N675, N663, N342, N246, N353);
and AND2 (N676, N673, N138);
not NOT1 (N677, N674);
nand NAND4 (N678, N671, N386, N444, N486);
and AND4 (N679, N675, N245, N302, N175);
not NOT1 (N680, N658);
buf BUF1 (N681, N649);
xor XOR2 (N682, N681, N110);
and AND4 (N683, N672, N247, N45, N193);
not NOT1 (N684, N677);
buf BUF1 (N685, N678);
buf BUF1 (N686, N684);
not NOT1 (N687, N686);
buf BUF1 (N688, N651);
nand NAND2 (N689, N687, N612);
or OR2 (N690, N679, N90);
nand NAND3 (N691, N689, N476, N315);
nand NAND3 (N692, N680, N28, N636);
nor NOR2 (N693, N692, N283);
xor XOR2 (N694, N670, N168);
or OR2 (N695, N682, N541);
buf BUF1 (N696, N688);
not NOT1 (N697, N664);
or OR3 (N698, N690, N598, N586);
not NOT1 (N699, N683);
and AND4 (N700, N696, N333, N588, N302);
or OR3 (N701, N695, N297, N464);
or OR4 (N702, N685, N10, N140, N321);
not NOT1 (N703, N691);
not NOT1 (N704, N697);
xor XOR2 (N705, N699, N682);
nor NOR2 (N706, N703, N201);
not NOT1 (N707, N693);
xor XOR2 (N708, N705, N117);
or OR4 (N709, N698, N22, N379, N477);
buf BUF1 (N710, N701);
xor XOR2 (N711, N708, N285);
buf BUF1 (N712, N711);
and AND3 (N713, N710, N506, N481);
and AND3 (N714, N704, N111, N660);
xor XOR2 (N715, N712, N637);
buf BUF1 (N716, N706);
buf BUF1 (N717, N694);
not NOT1 (N718, N713);
nor NOR3 (N719, N715, N165, N358);
nand NAND3 (N720, N709, N546, N28);
xor XOR2 (N721, N716, N325);
or OR4 (N722, N676, N500, N364, N707);
xor XOR2 (N723, N533, N366);
not NOT1 (N724, N722);
xor XOR2 (N725, N700, N416);
nor NOR3 (N726, N718, N68, N585);
and AND3 (N727, N702, N687, N127);
buf BUF1 (N728, N720);
xor XOR2 (N729, N727, N381);
nor NOR3 (N730, N726, N659, N193);
not NOT1 (N731, N728);
buf BUF1 (N732, N725);
or OR2 (N733, N732, N560);
not NOT1 (N734, N731);
nand NAND2 (N735, N729, N572);
or OR4 (N736, N734, N190, N650, N46);
not NOT1 (N737, N714);
or OR3 (N738, N721, N536, N342);
xor XOR2 (N739, N737, N268);
and AND4 (N740, N738, N69, N664, N728);
or OR3 (N741, N736, N403, N595);
and AND4 (N742, N735, N358, N55, N85);
not NOT1 (N743, N723);
and AND4 (N744, N724, N84, N244, N415);
not NOT1 (N745, N740);
nor NOR4 (N746, N739, N519, N356, N326);
nor NOR4 (N747, N717, N31, N712, N369);
nor NOR2 (N748, N741, N595);
and AND2 (N749, N747, N178);
nor NOR3 (N750, N743, N342, N566);
or OR4 (N751, N733, N310, N297, N172);
nand NAND2 (N752, N745, N534);
nor NOR4 (N753, N730, N455, N182, N74);
buf BUF1 (N754, N748);
xor XOR2 (N755, N752, N480);
xor XOR2 (N756, N754, N208);
xor XOR2 (N757, N744, N310);
buf BUF1 (N758, N750);
nor NOR3 (N759, N756, N312, N203);
buf BUF1 (N760, N719);
or OR2 (N761, N746, N333);
not NOT1 (N762, N755);
nand NAND4 (N763, N751, N501, N414, N46);
buf BUF1 (N764, N762);
not NOT1 (N765, N764);
xor XOR2 (N766, N742, N421);
xor XOR2 (N767, N763, N218);
xor XOR2 (N768, N760, N753);
and AND3 (N769, N32, N479, N640);
not NOT1 (N770, N765);
and AND2 (N771, N759, N75);
buf BUF1 (N772, N766);
and AND3 (N773, N772, N639, N197);
nand NAND3 (N774, N768, N764, N718);
and AND4 (N775, N761, N763, N409, N554);
nand NAND2 (N776, N775, N514);
not NOT1 (N777, N749);
not NOT1 (N778, N770);
not NOT1 (N779, N757);
or OR3 (N780, N779, N629, N147);
or OR2 (N781, N780, N501);
and AND4 (N782, N767, N748, N582, N668);
buf BUF1 (N783, N771);
nor NOR4 (N784, N773, N193, N544, N396);
not NOT1 (N785, N781);
or OR2 (N786, N782, N189);
buf BUF1 (N787, N778);
and AND3 (N788, N784, N242, N416);
not NOT1 (N789, N785);
not NOT1 (N790, N777);
not NOT1 (N791, N790);
nor NOR4 (N792, N787, N698, N259, N120);
not NOT1 (N793, N791);
nor NOR3 (N794, N776, N244, N14);
or OR4 (N795, N783, N27, N455, N580);
buf BUF1 (N796, N774);
buf BUF1 (N797, N758);
buf BUF1 (N798, N795);
nor NOR2 (N799, N788, N398);
nand NAND4 (N800, N798, N694, N383, N415);
xor XOR2 (N801, N799, N598);
not NOT1 (N802, N769);
xor XOR2 (N803, N802, N792);
and AND2 (N804, N307, N607);
buf BUF1 (N805, N789);
xor XOR2 (N806, N801, N682);
xor XOR2 (N807, N794, N701);
nand NAND4 (N808, N804, N714, N787, N101);
buf BUF1 (N809, N800);
or OR4 (N810, N807, N262, N57, N407);
xor XOR2 (N811, N786, N399);
nand NAND3 (N812, N810, N55, N171);
xor XOR2 (N813, N797, N658);
not NOT1 (N814, N813);
xor XOR2 (N815, N793, N88);
not NOT1 (N816, N814);
and AND3 (N817, N809, N554, N13);
nand NAND2 (N818, N803, N694);
nand NAND3 (N819, N815, N510, N719);
not NOT1 (N820, N806);
or OR3 (N821, N819, N204, N284);
not NOT1 (N822, N821);
not NOT1 (N823, N805);
nor NOR4 (N824, N823, N763, N263, N527);
nor NOR4 (N825, N816, N441, N757, N760);
nor NOR3 (N826, N820, N289, N249);
and AND2 (N827, N812, N246);
and AND4 (N828, N811, N156, N91, N735);
xor XOR2 (N829, N826, N349);
not NOT1 (N830, N818);
and AND3 (N831, N824, N663, N668);
nand NAND3 (N832, N830, N309, N237);
buf BUF1 (N833, N808);
or OR3 (N834, N822, N728, N549);
nand NAND3 (N835, N796, N570, N617);
nand NAND3 (N836, N817, N362, N566);
not NOT1 (N837, N835);
nor NOR4 (N838, N831, N518, N465, N739);
xor XOR2 (N839, N837, N302);
and AND2 (N840, N827, N358);
xor XOR2 (N841, N833, N798);
and AND2 (N842, N840, N257);
xor XOR2 (N843, N825, N41);
buf BUF1 (N844, N838);
nand NAND4 (N845, N832, N283, N64, N700);
buf BUF1 (N846, N828);
or OR4 (N847, N836, N457, N743, N425);
buf BUF1 (N848, N839);
buf BUF1 (N849, N846);
nor NOR4 (N850, N842, N762, N106, N360);
buf BUF1 (N851, N848);
nor NOR3 (N852, N829, N117, N711);
and AND3 (N853, N845, N404, N160);
nand NAND3 (N854, N850, N439, N676);
or OR3 (N855, N853, N490, N618);
and AND4 (N856, N849, N435, N820, N357);
or OR4 (N857, N841, N626, N557, N117);
nand NAND3 (N858, N856, N731, N585);
and AND2 (N859, N855, N329);
xor XOR2 (N860, N854, N695);
not NOT1 (N861, N852);
not NOT1 (N862, N834);
buf BUF1 (N863, N859);
nand NAND3 (N864, N843, N224, N446);
nor NOR2 (N865, N847, N313);
or OR4 (N866, N844, N71, N835, N569);
not NOT1 (N867, N864);
or OR4 (N868, N865, N258, N103, N796);
not NOT1 (N869, N861);
buf BUF1 (N870, N858);
xor XOR2 (N871, N862, N557);
xor XOR2 (N872, N870, N94);
not NOT1 (N873, N860);
nand NAND2 (N874, N857, N223);
nor NOR4 (N875, N869, N376, N44, N734);
buf BUF1 (N876, N871);
xor XOR2 (N877, N868, N455);
nor NOR3 (N878, N872, N691, N515);
nor NOR4 (N879, N873, N260, N106, N461);
nand NAND2 (N880, N879, N211);
buf BUF1 (N881, N863);
and AND3 (N882, N874, N92, N225);
or OR2 (N883, N866, N597);
and AND4 (N884, N875, N594, N244, N542);
and AND3 (N885, N877, N749, N654);
nor NOR3 (N886, N876, N747, N325);
or OR3 (N887, N878, N7, N705);
not NOT1 (N888, N882);
not NOT1 (N889, N886);
or OR2 (N890, N889, N762);
and AND3 (N891, N881, N852, N647);
and AND2 (N892, N851, N378);
nand NAND2 (N893, N891, N446);
buf BUF1 (N894, N885);
buf BUF1 (N895, N887);
and AND4 (N896, N892, N194, N737, N7);
xor XOR2 (N897, N883, N666);
nand NAND2 (N898, N880, N517);
nor NOR4 (N899, N898, N759, N547, N419);
xor XOR2 (N900, N867, N72);
and AND2 (N901, N896, N806);
or OR2 (N902, N894, N682);
nand NAND2 (N903, N902, N470);
nand NAND2 (N904, N893, N173);
nor NOR2 (N905, N890, N455);
nand NAND2 (N906, N903, N799);
nand NAND2 (N907, N906, N811);
not NOT1 (N908, N897);
xor XOR2 (N909, N901, N80);
and AND2 (N910, N895, N354);
nand NAND2 (N911, N884, N825);
and AND4 (N912, N899, N213, N804, N650);
xor XOR2 (N913, N907, N345);
not NOT1 (N914, N900);
xor XOR2 (N915, N905, N737);
nor NOR2 (N916, N912, N876);
not NOT1 (N917, N904);
or OR4 (N918, N888, N102, N567, N809);
endmodule