// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19;

output N25612,N25614,N25615,N25569,N25613,N25601,N25618,N25617,N25611,N25619;

or OR4 (N20, N9, N3, N16, N3);
xor XOR2 (N21, N20, N1);
buf BUF1 (N22, N20);
and AND4 (N23, N2, N22, N14, N12);
xor XOR2 (N24, N15, N15);
buf BUF1 (N25, N18);
xor XOR2 (N26, N18, N1);
not NOT1 (N27, N18);
or OR4 (N28, N3, N23, N15, N14);
nand NAND2 (N29, N15, N26);
not NOT1 (N30, N2);
nor NOR2 (N31, N29, N16);
nor NOR2 (N32, N29, N4);
xor XOR2 (N33, N21, N30);
or OR2 (N34, N17, N14);
nand NAND3 (N35, N8, N27, N32);
buf BUF1 (N36, N12);
xor XOR2 (N37, N31, N11);
xor XOR2 (N38, N33, N20);
and AND3 (N39, N30, N25, N34);
buf BUF1 (N40, N25);
or OR2 (N41, N21, N39);
not NOT1 (N42, N1);
xor XOR2 (N43, N32, N10);
not NOT1 (N44, N40);
buf BUF1 (N45, N28);
and AND2 (N46, N45, N7);
nor NOR3 (N47, N44, N12, N42);
nor NOR3 (N48, N34, N32, N15);
nor NOR3 (N49, N48, N28, N9);
xor XOR2 (N50, N46, N11);
nor NOR4 (N51, N47, N43, N22, N46);
nand NAND4 (N52, N17, N18, N9, N42);
or OR4 (N53, N50, N28, N30, N14);
and AND3 (N54, N38, N8, N47);
nor NOR3 (N55, N53, N8, N29);
buf BUF1 (N56, N41);
not NOT1 (N57, N49);
and AND3 (N58, N56, N56, N6);
nor NOR3 (N59, N24, N11, N21);
not NOT1 (N60, N57);
xor XOR2 (N61, N35, N14);
nor NOR3 (N62, N61, N9, N37);
buf BUF1 (N63, N56);
buf BUF1 (N64, N51);
nor NOR4 (N65, N63, N5, N58, N20);
not NOT1 (N66, N24);
nor NOR4 (N67, N62, N32, N12, N25);
xor XOR2 (N68, N65, N61);
not NOT1 (N69, N54);
and AND2 (N70, N67, N65);
buf BUF1 (N71, N36);
nand NAND2 (N72, N68, N20);
nor NOR4 (N73, N52, N4, N32, N40);
nand NAND3 (N74, N73, N34, N30);
buf BUF1 (N75, N69);
and AND3 (N76, N59, N20, N16);
nor NOR2 (N77, N74, N64);
and AND2 (N78, N58, N11);
or OR3 (N79, N78, N11, N62);
or OR3 (N80, N77, N13, N20);
and AND2 (N81, N80, N68);
buf BUF1 (N82, N79);
and AND4 (N83, N72, N6, N82, N55);
nand NAND3 (N84, N68, N68, N66);
not NOT1 (N85, N16);
nor NOR3 (N86, N13, N2, N67);
and AND4 (N87, N86, N31, N69, N83);
nand NAND4 (N88, N28, N3, N35, N5);
nor NOR3 (N89, N75, N72, N66);
not NOT1 (N90, N60);
not NOT1 (N91, N84);
xor XOR2 (N92, N87, N26);
or OR4 (N93, N70, N76, N49, N66);
nor NOR3 (N94, N79, N48, N80);
buf BUF1 (N95, N91);
and AND4 (N96, N92, N80, N92, N48);
nand NAND3 (N97, N89, N19, N16);
and AND3 (N98, N85, N38, N34);
xor XOR2 (N99, N95, N51);
nand NAND2 (N100, N99, N64);
xor XOR2 (N101, N88, N15);
nand NAND2 (N102, N101, N10);
and AND2 (N103, N98, N70);
buf BUF1 (N104, N103);
or OR4 (N105, N96, N15, N84, N7);
buf BUF1 (N106, N93);
buf BUF1 (N107, N71);
not NOT1 (N108, N97);
nand NAND4 (N109, N105, N95, N89, N74);
or OR4 (N110, N100, N65, N55, N37);
buf BUF1 (N111, N106);
and AND3 (N112, N102, N25, N2);
not NOT1 (N113, N108);
nor NOR3 (N114, N104, N16, N92);
nor NOR2 (N115, N94, N14);
xor XOR2 (N116, N112, N27);
and AND3 (N117, N115, N51, N29);
xor XOR2 (N118, N111, N95);
nor NOR2 (N119, N90, N76);
xor XOR2 (N120, N119, N9);
buf BUF1 (N121, N109);
buf BUF1 (N122, N116);
buf BUF1 (N123, N107);
nor NOR2 (N124, N123, N77);
nand NAND3 (N125, N118, N117, N100);
nand NAND2 (N126, N91, N70);
nand NAND3 (N127, N121, N53, N126);
or OR2 (N128, N74, N18);
xor XOR2 (N129, N120, N111);
nor NOR3 (N130, N127, N123, N4);
nand NAND4 (N131, N114, N120, N98, N56);
nand NAND4 (N132, N110, N84, N2, N122);
and AND4 (N133, N47, N90, N20, N94);
not NOT1 (N134, N124);
nand NAND3 (N135, N129, N42, N72);
or OR3 (N136, N128, N120, N62);
or OR3 (N137, N133, N83, N113);
or OR3 (N138, N129, N131, N29);
or OR2 (N139, N133, N26);
and AND3 (N140, N135, N137, N102);
xor XOR2 (N141, N42, N70);
and AND2 (N142, N136, N49);
and AND4 (N143, N141, N137, N120, N134);
nor NOR2 (N144, N87, N66);
buf BUF1 (N145, N140);
nand NAND3 (N146, N142, N40, N93);
buf BUF1 (N147, N125);
nand NAND2 (N148, N144, N67);
or OR4 (N149, N143, N92, N148, N38);
buf BUF1 (N150, N13);
buf BUF1 (N151, N138);
and AND3 (N152, N132, N69, N134);
nand NAND3 (N153, N139, N46, N44);
or OR4 (N154, N150, N1, N33, N79);
not NOT1 (N155, N147);
or OR3 (N156, N155, N96, N15);
xor XOR2 (N157, N81, N58);
not NOT1 (N158, N149);
xor XOR2 (N159, N151, N28);
nand NAND4 (N160, N153, N66, N64, N123);
and AND2 (N161, N156, N53);
xor XOR2 (N162, N154, N58);
buf BUF1 (N163, N162);
nand NAND3 (N164, N145, N131, N39);
nand NAND3 (N165, N158, N74, N8);
nand NAND2 (N166, N159, N65);
not NOT1 (N167, N166);
buf BUF1 (N168, N152);
and AND2 (N169, N168, N77);
or OR4 (N170, N164, N86, N26, N77);
nor NOR4 (N171, N161, N150, N106, N82);
buf BUF1 (N172, N167);
and AND4 (N173, N171, N94, N54, N77);
not NOT1 (N174, N157);
nor NOR4 (N175, N146, N169, N7, N161);
buf BUF1 (N176, N7);
and AND3 (N177, N175, N33, N81);
buf BUF1 (N178, N170);
or OR2 (N179, N178, N35);
buf BUF1 (N180, N172);
not NOT1 (N181, N176);
or OR3 (N182, N163, N98, N77);
not NOT1 (N183, N179);
xor XOR2 (N184, N181, N11);
buf BUF1 (N185, N180);
and AND4 (N186, N184, N79, N139, N149);
and AND4 (N187, N182, N96, N74, N62);
xor XOR2 (N188, N183, N82);
nand NAND3 (N189, N177, N180, N86);
xor XOR2 (N190, N173, N78);
and AND2 (N191, N187, N92);
buf BUF1 (N192, N191);
nand NAND3 (N193, N165, N73, N19);
buf BUF1 (N194, N189);
nor NOR3 (N195, N194, N31, N139);
not NOT1 (N196, N185);
or OR2 (N197, N160, N94);
and AND3 (N198, N190, N113, N75);
buf BUF1 (N199, N193);
nand NAND2 (N200, N130, N97);
nand NAND2 (N201, N186, N200);
nand NAND2 (N202, N28, N36);
or OR4 (N203, N174, N74, N116, N52);
nor NOR3 (N204, N203, N115, N19);
buf BUF1 (N205, N202);
xor XOR2 (N206, N196, N21);
nor NOR4 (N207, N188, N177, N82, N118);
nor NOR3 (N208, N206, N102, N188);
or OR4 (N209, N208, N37, N136, N37);
not NOT1 (N210, N198);
nand NAND2 (N211, N199, N125);
not NOT1 (N212, N209);
or OR4 (N213, N211, N80, N84, N33);
xor XOR2 (N214, N207, N81);
not NOT1 (N215, N214);
and AND3 (N216, N213, N38, N93);
buf BUF1 (N217, N210);
xor XOR2 (N218, N197, N90);
and AND4 (N219, N216, N179, N210, N195);
xor XOR2 (N220, N206, N211);
not NOT1 (N221, N220);
and AND4 (N222, N192, N99, N76, N156);
xor XOR2 (N223, N218, N105);
nor NOR2 (N224, N204, N149);
buf BUF1 (N225, N222);
not NOT1 (N226, N219);
xor XOR2 (N227, N224, N203);
nand NAND3 (N228, N221, N174, N48);
nor NOR2 (N229, N228, N136);
nand NAND2 (N230, N223, N181);
nand NAND2 (N231, N225, N228);
and AND2 (N232, N212, N175);
not NOT1 (N233, N232);
not NOT1 (N234, N205);
nand NAND4 (N235, N226, N57, N188, N201);
nor NOR3 (N236, N95, N92, N214);
not NOT1 (N237, N215);
xor XOR2 (N238, N227, N179);
or OR2 (N239, N233, N144);
xor XOR2 (N240, N235, N219);
buf BUF1 (N241, N229);
nor NOR4 (N242, N231, N64, N119, N236);
nor NOR4 (N243, N2, N132, N82, N41);
or OR2 (N244, N234, N112);
not NOT1 (N245, N240);
xor XOR2 (N246, N242, N105);
not NOT1 (N247, N238);
and AND4 (N248, N230, N93, N211, N243);
nor NOR2 (N249, N244, N62);
not NOT1 (N250, N44);
buf BUF1 (N251, N217);
buf BUF1 (N252, N249);
or OR4 (N253, N237, N33, N203, N32);
not NOT1 (N254, N250);
nand NAND4 (N255, N245, N24, N202, N213);
not NOT1 (N256, N253);
not NOT1 (N257, N252);
xor XOR2 (N258, N239, N23);
and AND4 (N259, N248, N154, N74, N178);
nor NOR3 (N260, N247, N161, N94);
buf BUF1 (N261, N258);
and AND3 (N262, N257, N190, N131);
or OR3 (N263, N256, N64, N250);
or OR4 (N264, N259, N121, N175, N250);
nor NOR4 (N265, N261, N264, N140, N19);
nand NAND4 (N266, N153, N230, N110, N130);
xor XOR2 (N267, N254, N41);
buf BUF1 (N268, N241);
nand NAND2 (N269, N263, N163);
nand NAND4 (N270, N255, N31, N20, N114);
buf BUF1 (N271, N246);
nand NAND2 (N272, N266, N140);
not NOT1 (N273, N269);
and AND4 (N274, N270, N69, N243, N80);
nor NOR4 (N275, N267, N251, N194, N70);
and AND2 (N276, N54, N209);
and AND2 (N277, N273, N256);
or OR4 (N278, N265, N132, N37, N57);
nor NOR2 (N279, N262, N181);
xor XOR2 (N280, N272, N217);
buf BUF1 (N281, N278);
xor XOR2 (N282, N277, N208);
nor NOR4 (N283, N268, N210, N213, N42);
or OR4 (N284, N279, N125, N32, N114);
nand NAND4 (N285, N271, N162, N48, N107);
nor NOR2 (N286, N276, N226);
or OR3 (N287, N274, N256, N218);
nor NOR3 (N288, N260, N116, N251);
or OR2 (N289, N287, N111);
buf BUF1 (N290, N282);
nand NAND4 (N291, N283, N98, N134, N263);
and AND3 (N292, N288, N98, N142);
or OR3 (N293, N291, N94, N249);
or OR3 (N294, N292, N137, N176);
not NOT1 (N295, N289);
nor NOR3 (N296, N286, N158, N223);
or OR2 (N297, N294, N239);
or OR3 (N298, N295, N230, N130);
xor XOR2 (N299, N296, N79);
buf BUF1 (N300, N293);
or OR2 (N301, N290, N4);
buf BUF1 (N302, N281);
nand NAND4 (N303, N275, N173, N296, N38);
not NOT1 (N304, N285);
xor XOR2 (N305, N299, N168);
not NOT1 (N306, N300);
not NOT1 (N307, N297);
buf BUF1 (N308, N303);
or OR3 (N309, N305, N123, N137);
nand NAND4 (N310, N308, N93, N74, N263);
xor XOR2 (N311, N309, N36);
not NOT1 (N312, N310);
nand NAND2 (N313, N301, N83);
not NOT1 (N314, N313);
buf BUF1 (N315, N298);
not NOT1 (N316, N302);
nand NAND3 (N317, N311, N144, N73);
or OR2 (N318, N317, N214);
xor XOR2 (N319, N315, N276);
or OR4 (N320, N316, N195, N15, N137);
nand NAND2 (N321, N314, N283);
nand NAND3 (N322, N307, N194, N167);
nor NOR3 (N323, N320, N237, N83);
or OR4 (N324, N318, N73, N211, N224);
and AND4 (N325, N324, N211, N4, N286);
nor NOR3 (N326, N321, N147, N71);
nand NAND4 (N327, N284, N136, N60, N125);
nor NOR2 (N328, N312, N103);
and AND2 (N329, N323, N98);
and AND2 (N330, N304, N213);
not NOT1 (N331, N322);
xor XOR2 (N332, N325, N114);
buf BUF1 (N333, N326);
nand NAND2 (N334, N333, N9);
not NOT1 (N335, N330);
buf BUF1 (N336, N280);
xor XOR2 (N337, N327, N131);
not NOT1 (N338, N329);
nand NAND3 (N339, N328, N196, N201);
nand NAND4 (N340, N332, N154, N330, N166);
not NOT1 (N341, N338);
xor XOR2 (N342, N331, N184);
and AND4 (N343, N334, N102, N279, N39);
and AND2 (N344, N341, N139);
buf BUF1 (N345, N342);
or OR4 (N346, N319, N37, N122, N344);
and AND3 (N347, N320, N34, N336);
buf BUF1 (N348, N212);
buf BUF1 (N349, N343);
and AND4 (N350, N347, N104, N197, N331);
nor NOR4 (N351, N340, N347, N35, N275);
xor XOR2 (N352, N351, N326);
or OR4 (N353, N352, N150, N333, N26);
and AND4 (N354, N353, N191, N37, N299);
and AND4 (N355, N346, N123, N160, N269);
nand NAND2 (N356, N339, N54);
nand NAND4 (N357, N306, N188, N179, N262);
buf BUF1 (N358, N335);
or OR3 (N359, N358, N211, N206);
buf BUF1 (N360, N354);
xor XOR2 (N361, N356, N267);
xor XOR2 (N362, N359, N135);
nor NOR4 (N363, N350, N84, N108, N88);
and AND3 (N364, N345, N272, N304);
xor XOR2 (N365, N348, N148);
nor NOR2 (N366, N349, N319);
nand NAND2 (N367, N364, N217);
buf BUF1 (N368, N361);
buf BUF1 (N369, N367);
and AND4 (N370, N363, N364, N268, N75);
nand NAND4 (N371, N370, N307, N74, N17);
nand NAND3 (N372, N371, N73, N105);
xor XOR2 (N373, N337, N271);
or OR2 (N374, N372, N215);
or OR3 (N375, N374, N84, N29);
buf BUF1 (N376, N355);
xor XOR2 (N377, N373, N44);
not NOT1 (N378, N366);
buf BUF1 (N379, N378);
not NOT1 (N380, N379);
and AND3 (N381, N377, N271, N173);
nand NAND2 (N382, N381, N96);
nor NOR3 (N383, N369, N30, N303);
nor NOR4 (N384, N368, N309, N338, N201);
nor NOR4 (N385, N357, N70, N52, N367);
buf BUF1 (N386, N362);
nor NOR3 (N387, N365, N247, N352);
not NOT1 (N388, N380);
buf BUF1 (N389, N360);
buf BUF1 (N390, N387);
or OR4 (N391, N386, N49, N231, N201);
not NOT1 (N392, N391);
not NOT1 (N393, N385);
buf BUF1 (N394, N384);
not NOT1 (N395, N390);
and AND2 (N396, N389, N221);
nand NAND3 (N397, N395, N344, N209);
and AND2 (N398, N382, N329);
xor XOR2 (N399, N394, N365);
and AND2 (N400, N396, N113);
xor XOR2 (N401, N398, N82);
and AND2 (N402, N388, N130);
and AND2 (N403, N399, N156);
buf BUF1 (N404, N401);
and AND4 (N405, N400, N90, N35, N12);
and AND4 (N406, N405, N41, N185, N280);
buf BUF1 (N407, N376);
nand NAND2 (N408, N383, N291);
and AND3 (N409, N375, N323, N332);
buf BUF1 (N410, N397);
buf BUF1 (N411, N403);
and AND4 (N412, N406, N68, N60, N388);
xor XOR2 (N413, N407, N43);
nor NOR4 (N414, N402, N167, N4, N155);
xor XOR2 (N415, N413, N144);
buf BUF1 (N416, N409);
nand NAND2 (N417, N393, N402);
and AND3 (N418, N416, N252, N328);
buf BUF1 (N419, N417);
nand NAND4 (N420, N412, N268, N387, N260);
buf BUF1 (N421, N392);
nand NAND3 (N422, N408, N270, N52);
nand NAND2 (N423, N414, N110);
buf BUF1 (N424, N421);
nor NOR2 (N425, N410, N83);
nor NOR2 (N426, N419, N339);
nor NOR3 (N427, N422, N166, N99);
not NOT1 (N428, N411);
buf BUF1 (N429, N424);
buf BUF1 (N430, N415);
nand NAND4 (N431, N427, N269, N85, N71);
nor NOR2 (N432, N431, N385);
or OR3 (N433, N420, N339, N173);
and AND3 (N434, N428, N128, N150);
or OR4 (N435, N404, N76, N255, N217);
nand NAND2 (N436, N435, N106);
buf BUF1 (N437, N433);
nor NOR4 (N438, N430, N348, N410, N243);
not NOT1 (N439, N436);
nand NAND2 (N440, N438, N387);
nand NAND4 (N441, N425, N144, N197, N227);
not NOT1 (N442, N429);
buf BUF1 (N443, N434);
nor NOR2 (N444, N442, N231);
and AND3 (N445, N423, N80, N15);
not NOT1 (N446, N441);
nand NAND2 (N447, N440, N371);
and AND2 (N448, N444, N418);
xor XOR2 (N449, N179, N204);
xor XOR2 (N450, N447, N135);
not NOT1 (N451, N445);
nor NOR3 (N452, N450, N103, N312);
not NOT1 (N453, N439);
not NOT1 (N454, N448);
and AND2 (N455, N426, N113);
xor XOR2 (N456, N455, N382);
not NOT1 (N457, N453);
and AND4 (N458, N452, N168, N443, N287);
and AND2 (N459, N82, N325);
and AND2 (N460, N449, N270);
xor XOR2 (N461, N458, N21);
nand NAND2 (N462, N457, N130);
not NOT1 (N463, N432);
buf BUF1 (N464, N437);
and AND3 (N465, N456, N191, N358);
xor XOR2 (N466, N461, N12);
nand NAND2 (N467, N464, N125);
xor XOR2 (N468, N446, N106);
or OR3 (N469, N454, N86, N372);
or OR3 (N470, N463, N282, N340);
xor XOR2 (N471, N469, N267);
xor XOR2 (N472, N460, N297);
xor XOR2 (N473, N472, N42);
and AND4 (N474, N467, N399, N2, N215);
xor XOR2 (N475, N462, N263);
and AND2 (N476, N471, N319);
xor XOR2 (N477, N470, N149);
xor XOR2 (N478, N465, N121);
xor XOR2 (N479, N476, N204);
not NOT1 (N480, N477);
nor NOR2 (N481, N468, N124);
nor NOR4 (N482, N473, N27, N185, N316);
nor NOR2 (N483, N475, N215);
xor XOR2 (N484, N481, N460);
nor NOR4 (N485, N451, N366, N39, N417);
and AND4 (N486, N482, N233, N263, N366);
xor XOR2 (N487, N478, N72);
and AND4 (N488, N485, N454, N347, N478);
not NOT1 (N489, N466);
nor NOR3 (N490, N489, N239, N456);
buf BUF1 (N491, N479);
xor XOR2 (N492, N488, N350);
not NOT1 (N493, N484);
buf BUF1 (N494, N492);
or OR3 (N495, N490, N231, N458);
buf BUF1 (N496, N474);
not NOT1 (N497, N493);
nor NOR2 (N498, N486, N320);
and AND4 (N499, N483, N229, N30, N101);
buf BUF1 (N500, N480);
and AND4 (N501, N499, N54, N55, N469);
or OR3 (N502, N496, N487, N221);
nor NOR3 (N503, N276, N267, N310);
nor NOR3 (N504, N497, N275, N218);
not NOT1 (N505, N502);
or OR3 (N506, N495, N171, N350);
nand NAND3 (N507, N506, N378, N504);
xor XOR2 (N508, N489, N21);
nor NOR3 (N509, N505, N452, N190);
nand NAND2 (N510, N507, N342);
buf BUF1 (N511, N500);
and AND2 (N512, N498, N244);
buf BUF1 (N513, N512);
and AND2 (N514, N508, N436);
nor NOR2 (N515, N510, N231);
not NOT1 (N516, N515);
or OR4 (N517, N511, N6, N171, N216);
and AND2 (N518, N513, N390);
not NOT1 (N519, N501);
nand NAND4 (N520, N517, N21, N264, N201);
nor NOR3 (N521, N491, N198, N154);
or OR4 (N522, N503, N281, N485, N26);
buf BUF1 (N523, N518);
buf BUF1 (N524, N520);
nand NAND2 (N525, N514, N26);
or OR2 (N526, N524, N220);
xor XOR2 (N527, N509, N110);
or OR2 (N528, N516, N248);
or OR3 (N529, N527, N333, N273);
xor XOR2 (N530, N459, N472);
nor NOR2 (N531, N519, N303);
and AND4 (N532, N525, N365, N121, N81);
nand NAND4 (N533, N532, N506, N489, N188);
nand NAND4 (N534, N530, N174, N489, N467);
nand NAND4 (N535, N529, N228, N309, N416);
nor NOR4 (N536, N523, N473, N523, N228);
not NOT1 (N537, N536);
nand NAND3 (N538, N537, N89, N190);
buf BUF1 (N539, N528);
and AND2 (N540, N539, N491);
or OR4 (N541, N526, N444, N12, N438);
and AND4 (N542, N494, N4, N383, N489);
and AND2 (N543, N522, N202);
buf BUF1 (N544, N534);
or OR2 (N545, N533, N137);
buf BUF1 (N546, N544);
not NOT1 (N547, N543);
buf BUF1 (N548, N541);
buf BUF1 (N549, N547);
or OR4 (N550, N542, N236, N386, N189);
nor NOR4 (N551, N540, N137, N306, N376);
or OR4 (N552, N546, N1, N262, N551);
and AND4 (N553, N63, N534, N296, N269);
not NOT1 (N554, N538);
buf BUF1 (N555, N535);
and AND4 (N556, N554, N548, N462, N251);
not NOT1 (N557, N265);
not NOT1 (N558, N553);
not NOT1 (N559, N557);
xor XOR2 (N560, N521, N254);
or OR3 (N561, N559, N56, N119);
nand NAND4 (N562, N556, N381, N202, N502);
buf BUF1 (N563, N550);
or OR2 (N564, N555, N511);
not NOT1 (N565, N558);
or OR2 (N566, N564, N169);
nor NOR2 (N567, N531, N105);
nor NOR3 (N568, N561, N110, N357);
buf BUF1 (N569, N560);
nand NAND3 (N570, N565, N385, N390);
not NOT1 (N571, N570);
nor NOR4 (N572, N545, N344, N139, N146);
buf BUF1 (N573, N572);
and AND3 (N574, N563, N101, N108);
nor NOR2 (N575, N571, N253);
xor XOR2 (N576, N549, N231);
and AND4 (N577, N568, N147, N257, N177);
not NOT1 (N578, N562);
nand NAND3 (N579, N575, N344, N435);
and AND2 (N580, N579, N548);
nor NOR2 (N581, N577, N355);
nor NOR3 (N582, N581, N21, N570);
nor NOR4 (N583, N582, N557, N418, N481);
xor XOR2 (N584, N574, N269);
buf BUF1 (N585, N567);
or OR2 (N586, N576, N374);
not NOT1 (N587, N573);
buf BUF1 (N588, N569);
or OR3 (N589, N586, N278, N554);
buf BUF1 (N590, N583);
buf BUF1 (N591, N552);
and AND2 (N592, N585, N90);
and AND4 (N593, N578, N288, N225, N120);
nor NOR4 (N594, N566, N426, N359, N16);
or OR4 (N595, N592, N211, N313, N208);
not NOT1 (N596, N589);
or OR2 (N597, N594, N343);
and AND3 (N598, N597, N1, N404);
not NOT1 (N599, N587);
buf BUF1 (N600, N599);
nand NAND4 (N601, N596, N552, N525, N41);
xor XOR2 (N602, N595, N389);
not NOT1 (N603, N588);
not NOT1 (N604, N580);
and AND4 (N605, N603, N461, N485, N378);
buf BUF1 (N606, N602);
buf BUF1 (N607, N601);
and AND3 (N608, N590, N147, N422);
or OR3 (N609, N608, N557, N401);
and AND4 (N610, N584, N47, N186, N590);
xor XOR2 (N611, N593, N551);
not NOT1 (N612, N600);
nand NAND2 (N613, N598, N493);
or OR2 (N614, N613, N380);
nor NOR3 (N615, N607, N450, N492);
not NOT1 (N616, N604);
xor XOR2 (N617, N611, N100);
or OR3 (N618, N605, N128, N237);
not NOT1 (N619, N612);
not NOT1 (N620, N591);
or OR4 (N621, N620, N108, N560, N326);
buf BUF1 (N622, N615);
or OR4 (N623, N610, N466, N251, N556);
buf BUF1 (N624, N621);
nand NAND2 (N625, N617, N130);
and AND2 (N626, N616, N578);
nand NAND4 (N627, N609, N557, N375, N420);
nor NOR3 (N628, N619, N328, N572);
xor XOR2 (N629, N626, N298);
not NOT1 (N630, N625);
and AND4 (N631, N606, N64, N362, N402);
or OR4 (N632, N622, N185, N225, N347);
not NOT1 (N633, N614);
xor XOR2 (N634, N623, N292);
or OR2 (N635, N633, N369);
buf BUF1 (N636, N635);
nor NOR3 (N637, N627, N428, N454);
nor NOR4 (N638, N631, N198, N226, N143);
xor XOR2 (N639, N636, N291);
nand NAND4 (N640, N639, N234, N171, N398);
and AND4 (N641, N640, N463, N234, N471);
nor NOR2 (N642, N637, N475);
nand NAND3 (N643, N642, N500, N594);
buf BUF1 (N644, N624);
buf BUF1 (N645, N634);
nor NOR4 (N646, N628, N89, N53, N308);
nand NAND3 (N647, N641, N561, N254);
buf BUF1 (N648, N630);
nand NAND2 (N649, N629, N118);
nor NOR2 (N650, N644, N226);
not NOT1 (N651, N638);
nor NOR4 (N652, N643, N488, N529, N415);
and AND2 (N653, N649, N381);
buf BUF1 (N654, N648);
nand NAND3 (N655, N654, N433, N57);
and AND2 (N656, N632, N540);
nor NOR3 (N657, N645, N13, N592);
and AND3 (N658, N618, N29, N58);
xor XOR2 (N659, N647, N570);
nor NOR3 (N660, N655, N506, N421);
nand NAND3 (N661, N660, N141, N110);
nor NOR4 (N662, N651, N328, N192, N111);
and AND4 (N663, N652, N628, N378, N477);
buf BUF1 (N664, N661);
nor NOR4 (N665, N663, N343, N628, N259);
and AND3 (N666, N658, N273, N67);
nand NAND2 (N667, N646, N195);
and AND4 (N668, N659, N137, N342, N481);
nor NOR3 (N669, N665, N506, N337);
buf BUF1 (N670, N650);
or OR4 (N671, N669, N23, N151, N175);
or OR4 (N672, N671, N406, N82, N231);
or OR2 (N673, N672, N109);
buf BUF1 (N674, N662);
and AND4 (N675, N668, N612, N542, N483);
nor NOR2 (N676, N657, N491);
buf BUF1 (N677, N674);
buf BUF1 (N678, N673);
not NOT1 (N679, N678);
or OR4 (N680, N670, N290, N393, N59);
xor XOR2 (N681, N653, N497);
nand NAND4 (N682, N656, N258, N427, N120);
buf BUF1 (N683, N680);
not NOT1 (N684, N666);
xor XOR2 (N685, N675, N481);
xor XOR2 (N686, N676, N369);
or OR3 (N687, N683, N158, N380);
not NOT1 (N688, N679);
nand NAND4 (N689, N677, N608, N598, N387);
xor XOR2 (N690, N682, N222);
or OR3 (N691, N688, N476, N319);
nor NOR4 (N692, N689, N497, N340, N38);
nand NAND3 (N693, N691, N254, N338);
buf BUF1 (N694, N690);
nor NOR2 (N695, N693, N109);
buf BUF1 (N696, N694);
nand NAND4 (N697, N681, N288, N602, N160);
and AND2 (N698, N685, N491);
or OR4 (N699, N687, N545, N448, N635);
buf BUF1 (N700, N664);
buf BUF1 (N701, N697);
and AND4 (N702, N699, N207, N394, N333);
xor XOR2 (N703, N696, N164);
buf BUF1 (N704, N703);
not NOT1 (N705, N692);
xor XOR2 (N706, N702, N550);
not NOT1 (N707, N667);
xor XOR2 (N708, N707, N631);
buf BUF1 (N709, N686);
nor NOR4 (N710, N704, N308, N199, N429);
or OR3 (N711, N709, N180, N220);
and AND4 (N712, N705, N480, N277, N123);
and AND4 (N713, N684, N85, N423, N404);
buf BUF1 (N714, N712);
and AND3 (N715, N706, N63, N713);
buf BUF1 (N716, N506);
not NOT1 (N717, N714);
or OR4 (N718, N711, N245, N287, N50);
or OR4 (N719, N701, N429, N570, N396);
nand NAND3 (N720, N715, N520, N273);
nor NOR3 (N721, N695, N77, N604);
or OR2 (N722, N698, N616);
or OR2 (N723, N710, N9);
or OR4 (N724, N720, N323, N126, N6);
not NOT1 (N725, N721);
xor XOR2 (N726, N722, N387);
and AND3 (N727, N708, N709, N615);
and AND3 (N728, N718, N579, N180);
nand NAND2 (N729, N726, N162);
buf BUF1 (N730, N727);
nand NAND3 (N731, N700, N11, N402);
xor XOR2 (N732, N725, N500);
nand NAND3 (N733, N732, N360, N536);
xor XOR2 (N734, N733, N593);
xor XOR2 (N735, N716, N444);
not NOT1 (N736, N735);
xor XOR2 (N737, N724, N409);
not NOT1 (N738, N729);
nand NAND3 (N739, N737, N682, N711);
nor NOR2 (N740, N736, N108);
not NOT1 (N741, N731);
nor NOR4 (N742, N719, N463, N652, N694);
nand NAND4 (N743, N717, N228, N312, N670);
nand NAND2 (N744, N741, N413);
xor XOR2 (N745, N742, N76);
buf BUF1 (N746, N739);
not NOT1 (N747, N728);
or OR3 (N748, N740, N514, N3);
buf BUF1 (N749, N730);
or OR4 (N750, N743, N143, N273, N268);
xor XOR2 (N751, N750, N53);
xor XOR2 (N752, N747, N323);
not NOT1 (N753, N734);
nand NAND4 (N754, N746, N118, N600, N690);
not NOT1 (N755, N738);
buf BUF1 (N756, N723);
or OR2 (N757, N754, N736);
nand NAND4 (N758, N756, N514, N10, N616);
xor XOR2 (N759, N751, N23);
buf BUF1 (N760, N759);
nor NOR3 (N761, N755, N278, N613);
nand NAND2 (N762, N752, N674);
buf BUF1 (N763, N760);
nor NOR3 (N764, N748, N83, N95);
not NOT1 (N765, N749);
not NOT1 (N766, N753);
buf BUF1 (N767, N761);
or OR2 (N768, N767, N291);
and AND3 (N769, N762, N361, N500);
xor XOR2 (N770, N744, N699);
nand NAND2 (N771, N768, N158);
buf BUF1 (N772, N766);
nand NAND2 (N773, N770, N83);
and AND4 (N774, N773, N523, N349, N20);
or OR2 (N775, N771, N8);
not NOT1 (N776, N769);
and AND2 (N777, N745, N42);
or OR4 (N778, N757, N193, N314, N220);
nand NAND3 (N779, N764, N590, N605);
nand NAND4 (N780, N763, N523, N90, N236);
xor XOR2 (N781, N777, N553);
xor XOR2 (N782, N765, N562);
buf BUF1 (N783, N782);
not NOT1 (N784, N775);
and AND2 (N785, N758, N313);
and AND4 (N786, N779, N163, N234, N646);
nor NOR2 (N787, N778, N685);
not NOT1 (N788, N780);
and AND2 (N789, N787, N192);
buf BUF1 (N790, N781);
not NOT1 (N791, N790);
and AND3 (N792, N774, N210, N133);
or OR2 (N793, N785, N42);
nand NAND4 (N794, N772, N41, N641, N34);
xor XOR2 (N795, N792, N455);
nand NAND3 (N796, N788, N510, N589);
nor NOR2 (N797, N784, N545);
not NOT1 (N798, N786);
nor NOR2 (N799, N798, N386);
nand NAND4 (N800, N794, N647, N242, N508);
not NOT1 (N801, N797);
nor NOR3 (N802, N789, N428, N643);
or OR3 (N803, N791, N588, N757);
or OR2 (N804, N793, N105);
or OR3 (N805, N802, N290, N255);
buf BUF1 (N806, N805);
nand NAND2 (N807, N795, N623);
buf BUF1 (N808, N807);
not NOT1 (N809, N803);
xor XOR2 (N810, N796, N127);
nand NAND4 (N811, N810, N11, N196, N40);
or OR3 (N812, N811, N324, N350);
buf BUF1 (N813, N799);
not NOT1 (N814, N800);
or OR2 (N815, N813, N173);
or OR2 (N816, N815, N236);
xor XOR2 (N817, N809, N785);
buf BUF1 (N818, N801);
nand NAND2 (N819, N776, N174);
nand NAND4 (N820, N818, N663, N307, N610);
xor XOR2 (N821, N812, N625);
not NOT1 (N822, N821);
xor XOR2 (N823, N816, N600);
buf BUF1 (N824, N783);
not NOT1 (N825, N823);
nor NOR3 (N826, N824, N70, N347);
buf BUF1 (N827, N820);
nand NAND2 (N828, N808, N793);
xor XOR2 (N829, N806, N568);
and AND4 (N830, N817, N57, N574, N551);
not NOT1 (N831, N827);
nand NAND3 (N832, N830, N462, N379);
buf BUF1 (N833, N822);
and AND3 (N834, N826, N263, N604);
and AND4 (N835, N804, N28, N314, N35);
nand NAND4 (N836, N831, N479, N352, N62);
nor NOR2 (N837, N834, N553);
nor NOR3 (N838, N832, N63, N311);
buf BUF1 (N839, N825);
xor XOR2 (N840, N838, N309);
buf BUF1 (N841, N814);
and AND3 (N842, N819, N319, N114);
nand NAND2 (N843, N841, N463);
buf BUF1 (N844, N828);
nor NOR3 (N845, N839, N799, N569);
buf BUF1 (N846, N844);
or OR3 (N847, N846, N641, N748);
and AND4 (N848, N833, N467, N692, N476);
nor NOR2 (N849, N837, N489);
nor NOR2 (N850, N848, N125);
nand NAND4 (N851, N840, N213, N570, N410);
and AND3 (N852, N835, N803, N586);
and AND4 (N853, N836, N563, N97, N67);
nor NOR3 (N854, N849, N678, N180);
and AND2 (N855, N842, N213);
nor NOR4 (N856, N852, N673, N403, N218);
or OR3 (N857, N854, N177, N287);
xor XOR2 (N858, N851, N187);
and AND3 (N859, N850, N249, N824);
buf BUF1 (N860, N829);
or OR4 (N861, N843, N476, N82, N172);
and AND3 (N862, N860, N796, N167);
or OR4 (N863, N856, N808, N61, N571);
xor XOR2 (N864, N847, N248);
nor NOR3 (N865, N864, N290, N471);
not NOT1 (N866, N853);
nand NAND3 (N867, N861, N179, N441);
nand NAND3 (N868, N858, N154, N550);
nor NOR2 (N869, N862, N550);
not NOT1 (N870, N865);
nand NAND4 (N871, N859, N276, N697, N270);
nand NAND3 (N872, N845, N763, N310);
buf BUF1 (N873, N868);
nor NOR4 (N874, N871, N665, N431, N685);
not NOT1 (N875, N874);
nor NOR3 (N876, N869, N27, N54);
nand NAND4 (N877, N866, N83, N424, N3);
not NOT1 (N878, N870);
not NOT1 (N879, N877);
or OR2 (N880, N857, N211);
not NOT1 (N881, N878);
xor XOR2 (N882, N880, N441);
nor NOR2 (N883, N879, N708);
nand NAND3 (N884, N855, N775, N557);
or OR4 (N885, N881, N759, N829, N817);
buf BUF1 (N886, N873);
buf BUF1 (N887, N886);
buf BUF1 (N888, N876);
and AND3 (N889, N875, N427, N715);
nand NAND2 (N890, N882, N349);
not NOT1 (N891, N884);
not NOT1 (N892, N872);
buf BUF1 (N893, N890);
xor XOR2 (N894, N867, N66);
nor NOR3 (N895, N863, N136, N685);
or OR2 (N896, N888, N827);
or OR3 (N897, N892, N510, N766);
xor XOR2 (N898, N883, N9);
nand NAND2 (N899, N898, N389);
nor NOR2 (N900, N889, N389);
nand NAND2 (N901, N894, N701);
not NOT1 (N902, N893);
or OR3 (N903, N895, N858, N289);
nor NOR4 (N904, N900, N516, N284, N550);
not NOT1 (N905, N891);
and AND2 (N906, N887, N703);
nand NAND4 (N907, N897, N30, N650, N799);
not NOT1 (N908, N901);
and AND3 (N909, N908, N503, N402);
or OR2 (N910, N905, N481);
nor NOR4 (N911, N896, N670, N514, N103);
xor XOR2 (N912, N910, N589);
nor NOR2 (N913, N906, N456);
and AND2 (N914, N907, N386);
not NOT1 (N915, N903);
not NOT1 (N916, N912);
nand NAND4 (N917, N916, N23, N903, N170);
nand NAND4 (N918, N885, N51, N778, N670);
and AND4 (N919, N911, N847, N134, N830);
and AND3 (N920, N919, N667, N838);
nor NOR4 (N921, N913, N382, N817, N740);
buf BUF1 (N922, N904);
buf BUF1 (N923, N914);
and AND4 (N924, N899, N453, N867, N390);
nor NOR2 (N925, N923, N505);
xor XOR2 (N926, N917, N207);
not NOT1 (N927, N925);
buf BUF1 (N928, N920);
buf BUF1 (N929, N922);
buf BUF1 (N930, N924);
or OR3 (N931, N927, N710, N582);
not NOT1 (N932, N931);
buf BUF1 (N933, N902);
nand NAND4 (N934, N930, N55, N643, N346);
not NOT1 (N935, N926);
buf BUF1 (N936, N928);
nor NOR4 (N937, N918, N346, N624, N631);
not NOT1 (N938, N929);
nand NAND3 (N939, N921, N340, N608);
or OR3 (N940, N909, N568, N715);
not NOT1 (N941, N932);
nor NOR2 (N942, N939, N32);
and AND4 (N943, N938, N508, N206, N84);
buf BUF1 (N944, N943);
buf BUF1 (N945, N942);
and AND3 (N946, N936, N220, N180);
nand NAND2 (N947, N941, N242);
nor NOR3 (N948, N946, N116, N355);
buf BUF1 (N949, N944);
or OR4 (N950, N945, N706, N224, N130);
nand NAND4 (N951, N950, N252, N556, N839);
buf BUF1 (N952, N949);
nand NAND2 (N953, N947, N621);
or OR2 (N954, N915, N251);
buf BUF1 (N955, N934);
not NOT1 (N956, N951);
or OR4 (N957, N937, N373, N71, N277);
and AND3 (N958, N955, N210, N12);
and AND2 (N959, N957, N222);
and AND3 (N960, N933, N554, N502);
buf BUF1 (N961, N952);
buf BUF1 (N962, N940);
nand NAND4 (N963, N961, N568, N476, N184);
or OR4 (N964, N954, N921, N936, N61);
or OR4 (N965, N960, N116, N517, N352);
nor NOR3 (N966, N962, N865, N487);
not NOT1 (N967, N963);
nand NAND4 (N968, N965, N560, N465, N422);
nand NAND2 (N969, N966, N24);
xor XOR2 (N970, N953, N672);
nor NOR2 (N971, N958, N799);
and AND4 (N972, N959, N915, N308, N606);
nor NOR2 (N973, N969, N788);
xor XOR2 (N974, N948, N912);
xor XOR2 (N975, N972, N369);
nor NOR2 (N976, N971, N17);
not NOT1 (N977, N970);
not NOT1 (N978, N935);
nand NAND4 (N979, N977, N333, N944, N932);
buf BUF1 (N980, N956);
nand NAND4 (N981, N979, N697, N481, N576);
xor XOR2 (N982, N964, N511);
buf BUF1 (N983, N982);
buf BUF1 (N984, N967);
nand NAND4 (N985, N981, N755, N43, N704);
xor XOR2 (N986, N985, N605);
and AND4 (N987, N974, N751, N763, N292);
nand NAND3 (N988, N980, N248, N873);
nand NAND3 (N989, N984, N728, N607);
buf BUF1 (N990, N986);
or OR2 (N991, N989, N832);
not NOT1 (N992, N987);
nor NOR2 (N993, N976, N248);
nor NOR4 (N994, N973, N633, N189, N144);
buf BUF1 (N995, N993);
or OR2 (N996, N995, N95);
buf BUF1 (N997, N988);
and AND4 (N998, N968, N583, N896, N747);
and AND3 (N999, N978, N444, N453);
buf BUF1 (N1000, N992);
and AND2 (N1001, N990, N958);
xor XOR2 (N1002, N1001, N973);
nand NAND4 (N1003, N998, N733, N400, N123);
nand NAND3 (N1004, N1000, N983, N121);
buf BUF1 (N1005, N999);
nor NOR4 (N1006, N941, N967, N740, N536);
xor XOR2 (N1007, N1005, N303);
xor XOR2 (N1008, N1002, N933);
not NOT1 (N1009, N994);
and AND2 (N1010, N1004, N790);
nor NOR3 (N1011, N996, N778, N883);
or OR3 (N1012, N1006, N21, N333);
or OR2 (N1013, N1007, N531);
nor NOR4 (N1014, N1010, N807, N566, N639);
nand NAND4 (N1015, N1013, N722, N64, N155);
not NOT1 (N1016, N1008);
or OR3 (N1017, N1003, N488, N115);
or OR2 (N1018, N1015, N846);
nand NAND3 (N1019, N1016, N192, N21);
buf BUF1 (N1020, N1011);
buf BUF1 (N1021, N1020);
buf BUF1 (N1022, N1017);
xor XOR2 (N1023, N1022, N792);
nor NOR4 (N1024, N975, N166, N466, N785);
not NOT1 (N1025, N1014);
nor NOR3 (N1026, N1019, N666, N263);
xor XOR2 (N1027, N1018, N143);
xor XOR2 (N1028, N997, N793);
buf BUF1 (N1029, N1027);
and AND2 (N1030, N1012, N1005);
buf BUF1 (N1031, N991);
buf BUF1 (N1032, N1031);
nor NOR3 (N1033, N1024, N271, N971);
nor NOR3 (N1034, N1026, N912, N845);
nor NOR3 (N1035, N1025, N915, N459);
buf BUF1 (N1036, N1029);
or OR3 (N1037, N1032, N239, N375);
nor NOR4 (N1038, N1009, N814, N667, N785);
not NOT1 (N1039, N1033);
and AND3 (N1040, N1035, N804, N243);
nor NOR4 (N1041, N1034, N924, N449, N1020);
xor XOR2 (N1042, N1023, N534);
not NOT1 (N1043, N1030);
nand NAND2 (N1044, N1021, N570);
buf BUF1 (N1045, N1039);
and AND2 (N1046, N1028, N377);
xor XOR2 (N1047, N1037, N952);
and AND2 (N1048, N1041, N862);
buf BUF1 (N1049, N1036);
xor XOR2 (N1050, N1046, N511);
or OR3 (N1051, N1043, N512, N683);
nand NAND2 (N1052, N1049, N696);
xor XOR2 (N1053, N1047, N1020);
nand NAND4 (N1054, N1044, N106, N181, N654);
xor XOR2 (N1055, N1051, N827);
or OR3 (N1056, N1040, N466, N425);
and AND2 (N1057, N1050, N808);
buf BUF1 (N1058, N1042);
or OR4 (N1059, N1055, N913, N897, N50);
nand NAND2 (N1060, N1056, N849);
and AND3 (N1061, N1059, N448, N592);
xor XOR2 (N1062, N1057, N722);
not NOT1 (N1063, N1062);
xor XOR2 (N1064, N1045, N1040);
not NOT1 (N1065, N1061);
not NOT1 (N1066, N1058);
and AND4 (N1067, N1063, N96, N284, N255);
or OR3 (N1068, N1053, N992, N106);
buf BUF1 (N1069, N1068);
not NOT1 (N1070, N1069);
nand NAND2 (N1071, N1064, N158);
nor NOR3 (N1072, N1052, N230, N710);
buf BUF1 (N1073, N1070);
xor XOR2 (N1074, N1067, N608);
nand NAND2 (N1075, N1066, N10);
nor NOR2 (N1076, N1065, N224);
nand NAND4 (N1077, N1073, N741, N696, N987);
xor XOR2 (N1078, N1048, N96);
xor XOR2 (N1079, N1074, N482);
nor NOR3 (N1080, N1076, N1051, N305);
or OR2 (N1081, N1079, N373);
or OR4 (N1082, N1054, N756, N443, N130);
nand NAND3 (N1083, N1038, N961, N735);
xor XOR2 (N1084, N1077, N331);
not NOT1 (N1085, N1060);
buf BUF1 (N1086, N1072);
nor NOR4 (N1087, N1081, N576, N248, N127);
and AND3 (N1088, N1083, N1019, N56);
and AND2 (N1089, N1085, N745);
buf BUF1 (N1090, N1089);
nand NAND3 (N1091, N1082, N874, N209);
nand NAND2 (N1092, N1078, N289);
xor XOR2 (N1093, N1084, N348);
not NOT1 (N1094, N1080);
nor NOR3 (N1095, N1075, N740, N817);
xor XOR2 (N1096, N1095, N944);
nand NAND4 (N1097, N1088, N472, N1081, N918);
or OR2 (N1098, N1087, N1014);
not NOT1 (N1099, N1098);
and AND2 (N1100, N1086, N23);
or OR3 (N1101, N1096, N167, N303);
and AND3 (N1102, N1071, N310, N503);
and AND4 (N1103, N1097, N36, N370, N93);
or OR3 (N1104, N1102, N739, N329);
nand NAND2 (N1105, N1100, N311);
buf BUF1 (N1106, N1104);
xor XOR2 (N1107, N1099, N1059);
xor XOR2 (N1108, N1094, N157);
and AND4 (N1109, N1093, N611, N876, N248);
nor NOR4 (N1110, N1103, N288, N183, N343);
buf BUF1 (N1111, N1109);
nand NAND2 (N1112, N1091, N246);
nand NAND2 (N1113, N1105, N318);
or OR4 (N1114, N1108, N708, N574, N879);
buf BUF1 (N1115, N1090);
nor NOR3 (N1116, N1110, N150, N442);
and AND2 (N1117, N1106, N514);
xor XOR2 (N1118, N1092, N548);
or OR2 (N1119, N1113, N877);
not NOT1 (N1120, N1107);
buf BUF1 (N1121, N1114);
not NOT1 (N1122, N1115);
nand NAND4 (N1123, N1119, N316, N1068, N428);
nor NOR2 (N1124, N1120, N223);
nand NAND2 (N1125, N1117, N1050);
and AND4 (N1126, N1122, N292, N798, N40);
nand NAND2 (N1127, N1126, N202);
nor NOR4 (N1128, N1116, N385, N612, N793);
buf BUF1 (N1129, N1118);
not NOT1 (N1130, N1128);
xor XOR2 (N1131, N1127, N556);
nor NOR2 (N1132, N1129, N1083);
and AND3 (N1133, N1123, N719, N336);
or OR2 (N1134, N1125, N406);
nor NOR4 (N1135, N1124, N834, N339, N350);
and AND4 (N1136, N1101, N858, N96, N119);
nor NOR4 (N1137, N1130, N1000, N780, N447);
nand NAND2 (N1138, N1112, N620);
or OR2 (N1139, N1121, N424);
nand NAND3 (N1140, N1138, N960, N897);
nand NAND2 (N1141, N1137, N529);
nand NAND4 (N1142, N1111, N690, N861, N238);
not NOT1 (N1143, N1134);
or OR2 (N1144, N1143, N788);
nand NAND2 (N1145, N1135, N121);
buf BUF1 (N1146, N1144);
and AND2 (N1147, N1132, N290);
nand NAND2 (N1148, N1136, N654);
buf BUF1 (N1149, N1139);
or OR4 (N1150, N1141, N1088, N239, N861);
xor XOR2 (N1151, N1133, N329);
xor XOR2 (N1152, N1140, N918);
and AND2 (N1153, N1131, N498);
or OR2 (N1154, N1153, N86);
xor XOR2 (N1155, N1147, N531);
xor XOR2 (N1156, N1146, N852);
buf BUF1 (N1157, N1156);
not NOT1 (N1158, N1157);
nand NAND2 (N1159, N1142, N1131);
not NOT1 (N1160, N1145);
buf BUF1 (N1161, N1150);
buf BUF1 (N1162, N1152);
nand NAND2 (N1163, N1149, N256);
or OR4 (N1164, N1158, N739, N828, N237);
xor XOR2 (N1165, N1162, N347);
buf BUF1 (N1166, N1154);
not NOT1 (N1167, N1166);
buf BUF1 (N1168, N1159);
or OR3 (N1169, N1163, N159, N970);
and AND4 (N1170, N1169, N588, N970, N953);
xor XOR2 (N1171, N1148, N988);
and AND2 (N1172, N1167, N87);
buf BUF1 (N1173, N1161);
not NOT1 (N1174, N1155);
or OR3 (N1175, N1171, N529, N83);
and AND3 (N1176, N1164, N872, N879);
xor XOR2 (N1177, N1165, N1025);
xor XOR2 (N1178, N1151, N997);
not NOT1 (N1179, N1172);
xor XOR2 (N1180, N1179, N144);
and AND2 (N1181, N1176, N660);
xor XOR2 (N1182, N1173, N1157);
nand NAND3 (N1183, N1182, N1158, N23);
buf BUF1 (N1184, N1183);
buf BUF1 (N1185, N1184);
buf BUF1 (N1186, N1160);
or OR4 (N1187, N1186, N202, N866, N450);
nor NOR3 (N1188, N1170, N1039, N911);
or OR4 (N1189, N1187, N29, N928, N580);
buf BUF1 (N1190, N1175);
xor XOR2 (N1191, N1168, N731);
not NOT1 (N1192, N1185);
buf BUF1 (N1193, N1192);
and AND4 (N1194, N1177, N195, N739, N935);
or OR4 (N1195, N1181, N630, N617, N1148);
xor XOR2 (N1196, N1174, N160);
xor XOR2 (N1197, N1180, N917);
xor XOR2 (N1198, N1190, N69);
not NOT1 (N1199, N1188);
not NOT1 (N1200, N1194);
or OR4 (N1201, N1197, N711, N972, N1192);
buf BUF1 (N1202, N1178);
xor XOR2 (N1203, N1200, N707);
and AND4 (N1204, N1196, N516, N566, N392);
not NOT1 (N1205, N1193);
xor XOR2 (N1206, N1202, N604);
buf BUF1 (N1207, N1198);
not NOT1 (N1208, N1195);
or OR4 (N1209, N1208, N654, N92, N83);
and AND2 (N1210, N1203, N763);
and AND4 (N1211, N1205, N1136, N1108, N724);
buf BUF1 (N1212, N1211);
and AND2 (N1213, N1199, N284);
not NOT1 (N1214, N1209);
nand NAND3 (N1215, N1210, N313, N850);
xor XOR2 (N1216, N1207, N51);
nand NAND3 (N1217, N1191, N734, N1131);
nand NAND3 (N1218, N1204, N693, N263);
nor NOR2 (N1219, N1214, N890);
buf BUF1 (N1220, N1213);
not NOT1 (N1221, N1216);
xor XOR2 (N1222, N1219, N601);
nand NAND4 (N1223, N1215, N490, N704, N889);
xor XOR2 (N1224, N1217, N1186);
nor NOR4 (N1225, N1206, N126, N1208, N1011);
buf BUF1 (N1226, N1221);
nand NAND2 (N1227, N1226, N446);
xor XOR2 (N1228, N1227, N1028);
buf BUF1 (N1229, N1212);
xor XOR2 (N1230, N1222, N785);
and AND2 (N1231, N1224, N397);
buf BUF1 (N1232, N1218);
nand NAND2 (N1233, N1231, N1198);
not NOT1 (N1234, N1189);
xor XOR2 (N1235, N1233, N1035);
xor XOR2 (N1236, N1220, N1138);
nand NAND3 (N1237, N1236, N770, N928);
nand NAND4 (N1238, N1225, N865, N1017, N531);
not NOT1 (N1239, N1234);
nor NOR3 (N1240, N1230, N93, N357);
not NOT1 (N1241, N1239);
or OR2 (N1242, N1238, N517);
nor NOR4 (N1243, N1229, N33, N415, N542);
and AND3 (N1244, N1228, N596, N441);
xor XOR2 (N1245, N1232, N266);
nand NAND2 (N1246, N1240, N411);
or OR2 (N1247, N1243, N688);
nand NAND2 (N1248, N1247, N306);
nand NAND3 (N1249, N1242, N816, N70);
and AND2 (N1250, N1241, N967);
buf BUF1 (N1251, N1250);
xor XOR2 (N1252, N1244, N231);
and AND2 (N1253, N1245, N662);
nor NOR2 (N1254, N1253, N114);
and AND3 (N1255, N1248, N443, N688);
and AND3 (N1256, N1201, N1024, N543);
or OR2 (N1257, N1249, N1148);
xor XOR2 (N1258, N1237, N465);
buf BUF1 (N1259, N1258);
xor XOR2 (N1260, N1257, N108);
nand NAND3 (N1261, N1235, N521, N412);
nand NAND3 (N1262, N1261, N969, N73);
not NOT1 (N1263, N1251);
nor NOR2 (N1264, N1223, N983);
buf BUF1 (N1265, N1262);
and AND4 (N1266, N1246, N452, N686, N743);
not NOT1 (N1267, N1263);
or OR3 (N1268, N1254, N912, N807);
nand NAND2 (N1269, N1256, N379);
and AND3 (N1270, N1265, N554, N627);
or OR3 (N1271, N1255, N301, N42);
and AND4 (N1272, N1252, N557, N670, N242);
nand NAND4 (N1273, N1264, N784, N854, N262);
nor NOR2 (N1274, N1273, N795);
buf BUF1 (N1275, N1267);
nor NOR4 (N1276, N1268, N1180, N1006, N1016);
not NOT1 (N1277, N1266);
buf BUF1 (N1278, N1274);
and AND3 (N1279, N1260, N1031, N11);
not NOT1 (N1280, N1277);
xor XOR2 (N1281, N1270, N1003);
and AND3 (N1282, N1280, N672, N1260);
or OR2 (N1283, N1272, N1244);
buf BUF1 (N1284, N1275);
xor XOR2 (N1285, N1281, N705);
buf BUF1 (N1286, N1285);
buf BUF1 (N1287, N1282);
and AND2 (N1288, N1283, N710);
or OR3 (N1289, N1286, N1211, N524);
nand NAND3 (N1290, N1269, N610, N266);
and AND3 (N1291, N1259, N84, N693);
nor NOR4 (N1292, N1276, N373, N529, N335);
buf BUF1 (N1293, N1279);
xor XOR2 (N1294, N1288, N1015);
nand NAND3 (N1295, N1294, N86, N366);
nor NOR4 (N1296, N1292, N319, N1250, N673);
nand NAND3 (N1297, N1291, N4, N218);
xor XOR2 (N1298, N1271, N1207);
and AND3 (N1299, N1297, N723, N326);
xor XOR2 (N1300, N1299, N1290);
nor NOR4 (N1301, N215, N1211, N690, N818);
or OR4 (N1302, N1289, N262, N407, N1012);
and AND2 (N1303, N1302, N1216);
and AND4 (N1304, N1284, N1275, N1134, N784);
nand NAND3 (N1305, N1301, N762, N720);
xor XOR2 (N1306, N1287, N9);
not NOT1 (N1307, N1306);
not NOT1 (N1308, N1296);
xor XOR2 (N1309, N1305, N1102);
nor NOR3 (N1310, N1293, N920, N1000);
xor XOR2 (N1311, N1310, N417);
not NOT1 (N1312, N1303);
not NOT1 (N1313, N1304);
nand NAND2 (N1314, N1298, N874);
not NOT1 (N1315, N1300);
xor XOR2 (N1316, N1307, N836);
not NOT1 (N1317, N1278);
nor NOR3 (N1318, N1308, N124, N771);
nor NOR3 (N1319, N1313, N467, N583);
xor XOR2 (N1320, N1319, N367);
buf BUF1 (N1321, N1320);
not NOT1 (N1322, N1318);
nand NAND3 (N1323, N1311, N479, N456);
nand NAND3 (N1324, N1312, N690, N415);
and AND2 (N1325, N1309, N1015);
or OR4 (N1326, N1324, N687, N46, N769);
and AND4 (N1327, N1321, N155, N438, N493);
and AND3 (N1328, N1315, N661, N471);
xor XOR2 (N1329, N1328, N973);
xor XOR2 (N1330, N1295, N303);
nor NOR2 (N1331, N1323, N25);
not NOT1 (N1332, N1329);
and AND3 (N1333, N1325, N970, N729);
nor NOR4 (N1334, N1326, N958, N302, N1009);
or OR3 (N1335, N1334, N907, N629);
xor XOR2 (N1336, N1330, N468);
or OR4 (N1337, N1336, N1033, N414, N221);
and AND3 (N1338, N1335, N144, N491);
xor XOR2 (N1339, N1338, N1312);
nor NOR3 (N1340, N1317, N163, N864);
and AND4 (N1341, N1316, N223, N1273, N1291);
not NOT1 (N1342, N1331);
nand NAND4 (N1343, N1327, N1025, N576, N655);
xor XOR2 (N1344, N1341, N1324);
not NOT1 (N1345, N1339);
or OR2 (N1346, N1314, N782);
and AND3 (N1347, N1346, N97, N366);
nand NAND4 (N1348, N1337, N952, N1032, N542);
not NOT1 (N1349, N1343);
not NOT1 (N1350, N1322);
nor NOR3 (N1351, N1347, N1049, N1267);
and AND4 (N1352, N1333, N980, N773, N1092);
and AND3 (N1353, N1351, N84, N1161);
xor XOR2 (N1354, N1352, N833);
nand NAND3 (N1355, N1342, N1109, N872);
xor XOR2 (N1356, N1355, N136);
xor XOR2 (N1357, N1353, N396);
xor XOR2 (N1358, N1356, N687);
and AND3 (N1359, N1348, N793, N788);
nor NOR2 (N1360, N1354, N556);
not NOT1 (N1361, N1360);
xor XOR2 (N1362, N1358, N547);
not NOT1 (N1363, N1349);
or OR3 (N1364, N1357, N561, N436);
not NOT1 (N1365, N1364);
buf BUF1 (N1366, N1340);
nor NOR3 (N1367, N1362, N291, N750);
buf BUF1 (N1368, N1345);
and AND3 (N1369, N1361, N216, N54);
nor NOR4 (N1370, N1365, N720, N778, N1357);
and AND2 (N1371, N1363, N1356);
and AND2 (N1372, N1369, N971);
nand NAND3 (N1373, N1344, N447, N226);
xor XOR2 (N1374, N1373, N645);
not NOT1 (N1375, N1359);
or OR3 (N1376, N1368, N478, N993);
nand NAND3 (N1377, N1366, N108, N887);
not NOT1 (N1378, N1375);
not NOT1 (N1379, N1376);
nor NOR3 (N1380, N1350, N531, N762);
nand NAND3 (N1381, N1379, N898, N1338);
not NOT1 (N1382, N1370);
or OR2 (N1383, N1371, N921);
nand NAND2 (N1384, N1383, N589);
nor NOR3 (N1385, N1377, N1213, N82);
nand NAND4 (N1386, N1378, N1261, N67, N801);
nand NAND4 (N1387, N1382, N395, N1317, N604);
nor NOR3 (N1388, N1380, N793, N766);
buf BUF1 (N1389, N1367);
nand NAND3 (N1390, N1389, N1240, N985);
and AND3 (N1391, N1388, N1200, N44);
nand NAND3 (N1392, N1372, N1132, N203);
nand NAND4 (N1393, N1385, N1390, N615, N896);
or OR3 (N1394, N454, N352, N975);
or OR4 (N1395, N1387, N961, N36, N1272);
nand NAND3 (N1396, N1384, N611, N1020);
buf BUF1 (N1397, N1386);
xor XOR2 (N1398, N1374, N1293);
nand NAND4 (N1399, N1393, N300, N833, N1250);
not NOT1 (N1400, N1332);
not NOT1 (N1401, N1381);
xor XOR2 (N1402, N1395, N796);
buf BUF1 (N1403, N1401);
buf BUF1 (N1404, N1396);
buf BUF1 (N1405, N1394);
and AND4 (N1406, N1391, N1025, N542, N129);
xor XOR2 (N1407, N1400, N932);
not NOT1 (N1408, N1399);
nand NAND2 (N1409, N1404, N199);
nand NAND4 (N1410, N1398, N165, N1282, N832);
nor NOR2 (N1411, N1402, N16);
nor NOR2 (N1412, N1405, N1264);
and AND2 (N1413, N1408, N1176);
buf BUF1 (N1414, N1403);
or OR3 (N1415, N1407, N1022, N1079);
xor XOR2 (N1416, N1413, N561);
buf BUF1 (N1417, N1415);
or OR2 (N1418, N1392, N873);
nor NOR4 (N1419, N1406, N540, N595, N716);
nand NAND3 (N1420, N1410, N660, N1002);
and AND2 (N1421, N1411, N787);
not NOT1 (N1422, N1416);
not NOT1 (N1423, N1412);
or OR3 (N1424, N1419, N1132, N278);
and AND2 (N1425, N1417, N1034);
or OR3 (N1426, N1420, N159, N455);
or OR3 (N1427, N1423, N209, N682);
and AND3 (N1428, N1414, N281, N532);
or OR3 (N1429, N1421, N227, N131);
nand NAND2 (N1430, N1427, N955);
nand NAND2 (N1431, N1424, N860);
or OR2 (N1432, N1397, N832);
buf BUF1 (N1433, N1430);
buf BUF1 (N1434, N1425);
nand NAND3 (N1435, N1418, N165, N1295);
nand NAND2 (N1436, N1435, N401);
xor XOR2 (N1437, N1426, N476);
or OR2 (N1438, N1429, N1266);
buf BUF1 (N1439, N1431);
nor NOR3 (N1440, N1439, N90, N307);
xor XOR2 (N1441, N1434, N1051);
buf BUF1 (N1442, N1433);
xor XOR2 (N1443, N1436, N45);
nor NOR2 (N1444, N1409, N1024);
nand NAND2 (N1445, N1441, N146);
buf BUF1 (N1446, N1444);
nand NAND3 (N1447, N1428, N500, N712);
nand NAND4 (N1448, N1437, N211, N334, N801);
not NOT1 (N1449, N1438);
not NOT1 (N1450, N1422);
nand NAND2 (N1451, N1447, N875);
buf BUF1 (N1452, N1451);
not NOT1 (N1453, N1432);
xor XOR2 (N1454, N1445, N135);
buf BUF1 (N1455, N1450);
not NOT1 (N1456, N1442);
buf BUF1 (N1457, N1443);
xor XOR2 (N1458, N1454, N1072);
and AND4 (N1459, N1457, N995, N581, N838);
nand NAND2 (N1460, N1440, N399);
nand NAND2 (N1461, N1452, N1249);
and AND3 (N1462, N1446, N1355, N5);
nor NOR3 (N1463, N1460, N863, N984);
buf BUF1 (N1464, N1461);
or OR4 (N1465, N1448, N109, N923, N51);
nor NOR3 (N1466, N1456, N577, N525);
buf BUF1 (N1467, N1464);
nand NAND3 (N1468, N1459, N195, N838);
buf BUF1 (N1469, N1455);
or OR3 (N1470, N1453, N327, N1227);
xor XOR2 (N1471, N1465, N1152);
not NOT1 (N1472, N1466);
nand NAND3 (N1473, N1471, N1066, N467);
xor XOR2 (N1474, N1468, N808);
not NOT1 (N1475, N1472);
or OR2 (N1476, N1469, N251);
and AND4 (N1477, N1470, N967, N532, N350);
nor NOR4 (N1478, N1463, N711, N38, N120);
xor XOR2 (N1479, N1449, N957);
buf BUF1 (N1480, N1458);
not NOT1 (N1481, N1467);
nor NOR3 (N1482, N1475, N17, N678);
not NOT1 (N1483, N1480);
xor XOR2 (N1484, N1483, N979);
nand NAND4 (N1485, N1462, N1291, N404, N102);
nand NAND2 (N1486, N1481, N664);
buf BUF1 (N1487, N1476);
buf BUF1 (N1488, N1473);
nor NOR3 (N1489, N1477, N103, N16);
nor NOR4 (N1490, N1482, N528, N708, N879);
or OR2 (N1491, N1489, N513);
nand NAND2 (N1492, N1485, N901);
xor XOR2 (N1493, N1479, N791);
or OR4 (N1494, N1491, N1328, N1212, N1023);
nand NAND2 (N1495, N1492, N1024);
xor XOR2 (N1496, N1494, N1466);
xor XOR2 (N1497, N1493, N726);
or OR4 (N1498, N1488, N887, N285, N1303);
buf BUF1 (N1499, N1495);
xor XOR2 (N1500, N1498, N114);
nor NOR2 (N1501, N1474, N286);
or OR3 (N1502, N1486, N987, N1110);
buf BUF1 (N1503, N1499);
or OR4 (N1504, N1503, N112, N950, N1046);
xor XOR2 (N1505, N1504, N983);
buf BUF1 (N1506, N1496);
nor NOR3 (N1507, N1506, N233, N920);
xor XOR2 (N1508, N1490, N1396);
not NOT1 (N1509, N1487);
not NOT1 (N1510, N1509);
xor XOR2 (N1511, N1510, N1173);
xor XOR2 (N1512, N1497, N798);
nor NOR4 (N1513, N1501, N1035, N488, N1406);
or OR4 (N1514, N1478, N570, N705, N333);
not NOT1 (N1515, N1514);
not NOT1 (N1516, N1511);
buf BUF1 (N1517, N1500);
xor XOR2 (N1518, N1512, N116);
nor NOR3 (N1519, N1507, N1291, N1070);
nand NAND2 (N1520, N1502, N1008);
and AND4 (N1521, N1508, N1128, N181, N430);
nor NOR4 (N1522, N1516, N262, N12, N594);
and AND3 (N1523, N1519, N1368, N110);
nor NOR4 (N1524, N1520, N1121, N642, N367);
xor XOR2 (N1525, N1515, N460);
nor NOR3 (N1526, N1518, N1128, N402);
and AND2 (N1527, N1524, N1518);
buf BUF1 (N1528, N1484);
and AND2 (N1529, N1513, N583);
buf BUF1 (N1530, N1522);
buf BUF1 (N1531, N1527);
and AND2 (N1532, N1517, N1294);
buf BUF1 (N1533, N1505);
and AND3 (N1534, N1526, N1375, N482);
nand NAND3 (N1535, N1533, N191, N33);
nand NAND4 (N1536, N1529, N401, N398, N478);
and AND2 (N1537, N1531, N238);
and AND3 (N1538, N1537, N1159, N1362);
not NOT1 (N1539, N1535);
and AND2 (N1540, N1532, N1393);
nand NAND4 (N1541, N1539, N1229, N885, N779);
buf BUF1 (N1542, N1534);
not NOT1 (N1543, N1530);
nor NOR3 (N1544, N1528, N1091, N557);
or OR3 (N1545, N1541, N438, N1512);
xor XOR2 (N1546, N1525, N1368);
buf BUF1 (N1547, N1545);
or OR3 (N1548, N1536, N13, N1258);
or OR2 (N1549, N1542, N1453);
buf BUF1 (N1550, N1548);
xor XOR2 (N1551, N1540, N1024);
nand NAND4 (N1552, N1547, N153, N37, N782);
or OR3 (N1553, N1538, N1079, N576);
not NOT1 (N1554, N1552);
and AND4 (N1555, N1543, N572, N90, N556);
or OR4 (N1556, N1551, N199, N598, N1421);
xor XOR2 (N1557, N1555, N1304);
nand NAND2 (N1558, N1544, N703);
not NOT1 (N1559, N1558);
nor NOR3 (N1560, N1559, N1520, N486);
not NOT1 (N1561, N1560);
nor NOR4 (N1562, N1546, N386, N1234, N616);
not NOT1 (N1563, N1549);
buf BUF1 (N1564, N1553);
buf BUF1 (N1565, N1556);
not NOT1 (N1566, N1557);
xor XOR2 (N1567, N1563, N1246);
xor XOR2 (N1568, N1523, N827);
xor XOR2 (N1569, N1562, N1532);
nor NOR2 (N1570, N1567, N667);
not NOT1 (N1571, N1554);
or OR4 (N1572, N1566, N986, N1570, N760);
and AND4 (N1573, N1259, N270, N158, N329);
nor NOR4 (N1574, N1521, N960, N576, N543);
and AND3 (N1575, N1571, N957, N112);
nand NAND2 (N1576, N1565, N320);
buf BUF1 (N1577, N1572);
nor NOR2 (N1578, N1569, N119);
nand NAND4 (N1579, N1576, N1087, N443, N1423);
and AND3 (N1580, N1577, N1141, N1093);
nor NOR4 (N1581, N1550, N1463, N658, N1509);
not NOT1 (N1582, N1581);
buf BUF1 (N1583, N1582);
not NOT1 (N1584, N1579);
nand NAND3 (N1585, N1583, N1171, N1232);
nor NOR3 (N1586, N1568, N682, N644);
buf BUF1 (N1587, N1585);
nand NAND4 (N1588, N1575, N208, N816, N166);
buf BUF1 (N1589, N1586);
nor NOR2 (N1590, N1564, N57);
buf BUF1 (N1591, N1587);
nor NOR3 (N1592, N1561, N590, N873);
xor XOR2 (N1593, N1578, N53);
not NOT1 (N1594, N1590);
and AND4 (N1595, N1588, N1453, N888, N1373);
nor NOR4 (N1596, N1595, N1552, N1562, N327);
or OR4 (N1597, N1593, N394, N1106, N974);
nor NOR4 (N1598, N1597, N711, N737, N458);
nand NAND2 (N1599, N1591, N562);
nor NOR4 (N1600, N1592, N1281, N551, N1349);
and AND3 (N1601, N1598, N1485, N35);
not NOT1 (N1602, N1599);
not NOT1 (N1603, N1594);
nor NOR2 (N1604, N1596, N612);
not NOT1 (N1605, N1601);
buf BUF1 (N1606, N1603);
and AND4 (N1607, N1584, N326, N735, N263);
buf BUF1 (N1608, N1574);
nor NOR3 (N1609, N1602, N1450, N1012);
xor XOR2 (N1610, N1608, N1400);
not NOT1 (N1611, N1573);
nor NOR2 (N1612, N1609, N484);
nand NAND2 (N1613, N1605, N1540);
xor XOR2 (N1614, N1580, N239);
nand NAND2 (N1615, N1607, N1082);
or OR2 (N1616, N1589, N751);
or OR4 (N1617, N1615, N18, N766, N535);
and AND3 (N1618, N1613, N1427, N178);
buf BUF1 (N1619, N1610);
and AND3 (N1620, N1617, N453, N1550);
nand NAND3 (N1621, N1618, N1234, N854);
nand NAND3 (N1622, N1606, N443, N463);
or OR4 (N1623, N1620, N298, N1565, N15);
or OR3 (N1624, N1616, N155, N58);
and AND4 (N1625, N1621, N874, N84, N1106);
and AND3 (N1626, N1614, N989, N484);
xor XOR2 (N1627, N1612, N1571);
xor XOR2 (N1628, N1626, N1270);
xor XOR2 (N1629, N1611, N527);
not NOT1 (N1630, N1623);
nor NOR4 (N1631, N1604, N702, N224, N781);
nor NOR3 (N1632, N1631, N64, N99);
nor NOR4 (N1633, N1632, N167, N797, N426);
xor XOR2 (N1634, N1630, N1);
or OR2 (N1635, N1627, N1025);
or OR2 (N1636, N1628, N72);
xor XOR2 (N1637, N1636, N338);
xor XOR2 (N1638, N1634, N1157);
and AND4 (N1639, N1624, N355, N783, N538);
or OR4 (N1640, N1600, N769, N829, N1222);
or OR2 (N1641, N1622, N757);
or OR4 (N1642, N1633, N939, N1322, N960);
xor XOR2 (N1643, N1637, N1631);
or OR3 (N1644, N1643, N334, N807);
and AND3 (N1645, N1640, N1031, N1221);
buf BUF1 (N1646, N1625);
nand NAND2 (N1647, N1644, N227);
nand NAND2 (N1648, N1619, N303);
buf BUF1 (N1649, N1645);
buf BUF1 (N1650, N1639);
xor XOR2 (N1651, N1649, N668);
nor NOR4 (N1652, N1651, N1567, N1640, N986);
or OR3 (N1653, N1652, N505, N1414);
and AND4 (N1654, N1638, N51, N1073, N408);
nand NAND4 (N1655, N1648, N380, N956, N615);
buf BUF1 (N1656, N1653);
not NOT1 (N1657, N1655);
not NOT1 (N1658, N1629);
buf BUF1 (N1659, N1656);
not NOT1 (N1660, N1650);
buf BUF1 (N1661, N1642);
and AND4 (N1662, N1654, N508, N1413, N1);
nand NAND2 (N1663, N1647, N1167);
nand NAND4 (N1664, N1659, N1284, N1098, N558);
nor NOR4 (N1665, N1664, N1080, N91, N164);
nor NOR4 (N1666, N1641, N1640, N392, N638);
xor XOR2 (N1667, N1661, N1315);
xor XOR2 (N1668, N1646, N927);
not NOT1 (N1669, N1663);
not NOT1 (N1670, N1669);
and AND3 (N1671, N1657, N303, N1429);
xor XOR2 (N1672, N1660, N730);
buf BUF1 (N1673, N1665);
and AND3 (N1674, N1667, N126, N1526);
and AND2 (N1675, N1662, N1052);
and AND3 (N1676, N1672, N1002, N800);
and AND4 (N1677, N1674, N387, N27, N175);
buf BUF1 (N1678, N1635);
nand NAND2 (N1679, N1677, N1057);
nor NOR3 (N1680, N1671, N1145, N346);
xor XOR2 (N1681, N1666, N711);
and AND3 (N1682, N1676, N14, N232);
or OR3 (N1683, N1678, N773, N1299);
not NOT1 (N1684, N1673);
not NOT1 (N1685, N1683);
and AND4 (N1686, N1670, N835, N392, N1005);
not NOT1 (N1687, N1658);
and AND2 (N1688, N1679, N1393);
not NOT1 (N1689, N1682);
xor XOR2 (N1690, N1675, N743);
and AND4 (N1691, N1690, N1476, N1641, N430);
or OR4 (N1692, N1688, N390, N595, N938);
not NOT1 (N1693, N1689);
nand NAND2 (N1694, N1680, N808);
nor NOR2 (N1695, N1684, N537);
nor NOR4 (N1696, N1687, N1391, N1370, N381);
and AND2 (N1697, N1695, N1192);
xor XOR2 (N1698, N1681, N684);
xor XOR2 (N1699, N1696, N1330);
nor NOR2 (N1700, N1698, N1543);
or OR3 (N1701, N1691, N973, N1677);
xor XOR2 (N1702, N1694, N1619);
buf BUF1 (N1703, N1697);
nand NAND4 (N1704, N1692, N599, N114, N193);
buf BUF1 (N1705, N1702);
buf BUF1 (N1706, N1686);
xor XOR2 (N1707, N1668, N1669);
buf BUF1 (N1708, N1705);
nor NOR3 (N1709, N1700, N1087, N190);
buf BUF1 (N1710, N1703);
buf BUF1 (N1711, N1701);
nand NAND3 (N1712, N1685, N1401, N399);
xor XOR2 (N1713, N1710, N128);
buf BUF1 (N1714, N1712);
nor NOR3 (N1715, N1708, N598, N1692);
nand NAND4 (N1716, N1713, N972, N340, N1236);
buf BUF1 (N1717, N1699);
nor NOR4 (N1718, N1716, N638, N869, N450);
xor XOR2 (N1719, N1704, N449);
not NOT1 (N1720, N1706);
not NOT1 (N1721, N1714);
not NOT1 (N1722, N1721);
buf BUF1 (N1723, N1722);
buf BUF1 (N1724, N1715);
not NOT1 (N1725, N1707);
and AND3 (N1726, N1723, N1697, N354);
nand NAND2 (N1727, N1718, N964);
and AND4 (N1728, N1725, N1629, N884, N1344);
not NOT1 (N1729, N1717);
and AND4 (N1730, N1729, N760, N401, N23);
buf BUF1 (N1731, N1730);
and AND2 (N1732, N1719, N1679);
nand NAND4 (N1733, N1726, N1524, N1661, N680);
and AND3 (N1734, N1709, N1215, N1414);
buf BUF1 (N1735, N1727);
not NOT1 (N1736, N1732);
and AND2 (N1737, N1733, N1675);
buf BUF1 (N1738, N1711);
xor XOR2 (N1739, N1728, N711);
nor NOR3 (N1740, N1731, N1279, N1683);
and AND2 (N1741, N1740, N194);
or OR2 (N1742, N1736, N1040);
nor NOR2 (N1743, N1741, N1063);
nor NOR4 (N1744, N1724, N504, N1259, N837);
buf BUF1 (N1745, N1738);
nand NAND2 (N1746, N1739, N895);
and AND3 (N1747, N1745, N1291, N416);
xor XOR2 (N1748, N1747, N1731);
nor NOR2 (N1749, N1743, N6);
buf BUF1 (N1750, N1735);
not NOT1 (N1751, N1744);
nor NOR2 (N1752, N1750, N1665);
xor XOR2 (N1753, N1748, N734);
nand NAND2 (N1754, N1751, N512);
and AND3 (N1755, N1693, N379, N82);
or OR4 (N1756, N1755, N1671, N1621, N280);
and AND4 (N1757, N1746, N1020, N1667, N1609);
xor XOR2 (N1758, N1756, N1710);
xor XOR2 (N1759, N1742, N1170);
nor NOR4 (N1760, N1720, N1174, N1088, N1714);
nor NOR4 (N1761, N1759, N566, N529, N1123);
nor NOR3 (N1762, N1749, N184, N504);
nand NAND4 (N1763, N1752, N1720, N1142, N1036);
nor NOR4 (N1764, N1763, N266, N935, N572);
nor NOR2 (N1765, N1762, N1225);
not NOT1 (N1766, N1753);
not NOT1 (N1767, N1760);
xor XOR2 (N1768, N1754, N350);
xor XOR2 (N1769, N1768, N69);
and AND4 (N1770, N1757, N801, N1561, N954);
nand NAND3 (N1771, N1767, N637, N1251);
not NOT1 (N1772, N1770);
and AND3 (N1773, N1772, N1346, N970);
and AND4 (N1774, N1769, N1623, N375, N363);
nand NAND3 (N1775, N1771, N1550, N561);
not NOT1 (N1776, N1774);
nand NAND4 (N1777, N1764, N515, N4, N224);
or OR4 (N1778, N1773, N1712, N270, N1438);
and AND2 (N1779, N1775, N1191);
or OR4 (N1780, N1761, N937, N587, N335);
buf BUF1 (N1781, N1777);
nor NOR3 (N1782, N1737, N352, N1561);
and AND2 (N1783, N1782, N802);
not NOT1 (N1784, N1766);
nor NOR4 (N1785, N1734, N966, N745, N582);
xor XOR2 (N1786, N1781, N1491);
nand NAND2 (N1787, N1784, N727);
nor NOR3 (N1788, N1786, N1475, N569);
or OR3 (N1789, N1758, N1169, N1086);
buf BUF1 (N1790, N1783);
and AND4 (N1791, N1778, N949, N810, N1013);
nor NOR4 (N1792, N1787, N1229, N1340, N86);
buf BUF1 (N1793, N1765);
buf BUF1 (N1794, N1791);
nor NOR4 (N1795, N1794, N215, N348, N168);
buf BUF1 (N1796, N1780);
buf BUF1 (N1797, N1790);
nor NOR3 (N1798, N1797, N696, N1671);
and AND3 (N1799, N1796, N380, N1494);
nor NOR3 (N1800, N1798, N1228, N1746);
xor XOR2 (N1801, N1792, N783);
or OR3 (N1802, N1793, N588, N1017);
or OR4 (N1803, N1779, N1792, N1553, N587);
or OR4 (N1804, N1803, N486, N215, N597);
nand NAND4 (N1805, N1788, N723, N695, N27);
xor XOR2 (N1806, N1776, N1754);
xor XOR2 (N1807, N1789, N114);
and AND3 (N1808, N1800, N2, N71);
buf BUF1 (N1809, N1802);
xor XOR2 (N1810, N1807, N493);
or OR3 (N1811, N1795, N1623, N356);
and AND2 (N1812, N1785, N199);
or OR2 (N1813, N1809, N922);
buf BUF1 (N1814, N1811);
nand NAND2 (N1815, N1808, N304);
buf BUF1 (N1816, N1806);
and AND3 (N1817, N1804, N1588, N207);
xor XOR2 (N1818, N1812, N1544);
xor XOR2 (N1819, N1801, N515);
nor NOR3 (N1820, N1814, N1781, N1396);
xor XOR2 (N1821, N1817, N388);
nor NOR2 (N1822, N1816, N1188);
xor XOR2 (N1823, N1819, N977);
or OR2 (N1824, N1820, N43);
nor NOR4 (N1825, N1823, N34, N840, N964);
nand NAND4 (N1826, N1813, N44, N1337, N415);
buf BUF1 (N1827, N1805);
buf BUF1 (N1828, N1825);
or OR4 (N1829, N1826, N349, N1071, N622);
xor XOR2 (N1830, N1815, N773);
nor NOR3 (N1831, N1821, N550, N1531);
not NOT1 (N1832, N1810);
buf BUF1 (N1833, N1832);
not NOT1 (N1834, N1833);
nor NOR2 (N1835, N1822, N1017);
not NOT1 (N1836, N1831);
nand NAND4 (N1837, N1830, N225, N613, N1380);
nor NOR3 (N1838, N1835, N1389, N28);
or OR2 (N1839, N1829, N999);
or OR2 (N1840, N1827, N697);
or OR3 (N1841, N1838, N858, N922);
xor XOR2 (N1842, N1818, N406);
xor XOR2 (N1843, N1841, N1318);
or OR4 (N1844, N1839, N361, N682, N282);
or OR3 (N1845, N1836, N182, N1429);
or OR2 (N1846, N1845, N595);
not NOT1 (N1847, N1844);
nand NAND4 (N1848, N1840, N1614, N320, N324);
nand NAND4 (N1849, N1846, N391, N1197, N1213);
or OR2 (N1850, N1848, N1327);
and AND4 (N1851, N1837, N985, N1693, N869);
nand NAND4 (N1852, N1828, N114, N228, N1729);
xor XOR2 (N1853, N1850, N454);
nand NAND3 (N1854, N1852, N662, N1327);
buf BUF1 (N1855, N1851);
not NOT1 (N1856, N1854);
or OR4 (N1857, N1799, N59, N18, N134);
xor XOR2 (N1858, N1842, N1210);
buf BUF1 (N1859, N1857);
xor XOR2 (N1860, N1859, N1199);
nand NAND2 (N1861, N1858, N503);
xor XOR2 (N1862, N1861, N1076);
nand NAND4 (N1863, N1847, N594, N37, N101);
not NOT1 (N1864, N1853);
buf BUF1 (N1865, N1824);
buf BUF1 (N1866, N1860);
buf BUF1 (N1867, N1863);
not NOT1 (N1868, N1867);
not NOT1 (N1869, N1849);
not NOT1 (N1870, N1866);
buf BUF1 (N1871, N1834);
nor NOR4 (N1872, N1864, N1349, N1009, N992);
nor NOR4 (N1873, N1843, N841, N636, N1865);
xor XOR2 (N1874, N1609, N1482);
nand NAND3 (N1875, N1872, N1065, N1213);
nor NOR4 (N1876, N1874, N1033, N36, N1828);
not NOT1 (N1877, N1862);
buf BUF1 (N1878, N1869);
not NOT1 (N1879, N1871);
or OR2 (N1880, N1877, N741);
nor NOR2 (N1881, N1878, N1162);
or OR2 (N1882, N1868, N261);
or OR4 (N1883, N1876, N1139, N1682, N1583);
nor NOR3 (N1884, N1880, N1191, N1004);
and AND2 (N1885, N1856, N113);
or OR4 (N1886, N1883, N597, N256, N974);
buf BUF1 (N1887, N1879);
nor NOR4 (N1888, N1855, N125, N348, N32);
nand NAND4 (N1889, N1885, N421, N1258, N832);
nand NAND3 (N1890, N1881, N1428, N23);
or OR3 (N1891, N1870, N1468, N801);
buf BUF1 (N1892, N1882);
xor XOR2 (N1893, N1891, N620);
nor NOR2 (N1894, N1873, N1145);
nand NAND4 (N1895, N1890, N1355, N1480, N1364);
nand NAND4 (N1896, N1888, N676, N401, N1209);
nand NAND2 (N1897, N1893, N471);
and AND2 (N1898, N1895, N1746);
nor NOR2 (N1899, N1889, N1267);
not NOT1 (N1900, N1899);
xor XOR2 (N1901, N1896, N336);
nand NAND2 (N1902, N1884, N173);
not NOT1 (N1903, N1887);
nor NOR3 (N1904, N1875, N873, N537);
not NOT1 (N1905, N1900);
not NOT1 (N1906, N1892);
nand NAND4 (N1907, N1904, N872, N972, N193);
not NOT1 (N1908, N1898);
not NOT1 (N1909, N1908);
nand NAND4 (N1910, N1906, N1380, N104, N1587);
and AND4 (N1911, N1886, N685, N1721, N759);
not NOT1 (N1912, N1902);
nand NAND3 (N1913, N1901, N1676, N1351);
not NOT1 (N1914, N1910);
and AND2 (N1915, N1914, N871);
buf BUF1 (N1916, N1915);
buf BUF1 (N1917, N1903);
buf BUF1 (N1918, N1911);
nand NAND3 (N1919, N1894, N1328, N1890);
buf BUF1 (N1920, N1916);
nor NOR3 (N1921, N1897, N1171, N342);
nand NAND2 (N1922, N1907, N526);
nor NOR3 (N1923, N1922, N606, N698);
not NOT1 (N1924, N1918);
and AND4 (N1925, N1909, N895, N40, N780);
nand NAND2 (N1926, N1905, N385);
xor XOR2 (N1927, N1921, N1558);
or OR4 (N1928, N1912, N930, N962, N195);
and AND4 (N1929, N1923, N850, N331, N717);
nor NOR3 (N1930, N1919, N491, N393);
and AND4 (N1931, N1913, N1864, N1727, N1361);
nor NOR4 (N1932, N1917, N504, N1562, N1918);
nor NOR3 (N1933, N1924, N521, N786);
buf BUF1 (N1934, N1920);
nand NAND2 (N1935, N1932, N524);
or OR3 (N1936, N1933, N1102, N1419);
not NOT1 (N1937, N1935);
xor XOR2 (N1938, N1931, N915);
or OR2 (N1939, N1937, N1787);
nor NOR4 (N1940, N1929, N1885, N952, N545);
and AND4 (N1941, N1925, N888, N197, N694);
buf BUF1 (N1942, N1938);
xor XOR2 (N1943, N1936, N1);
and AND2 (N1944, N1927, N462);
not NOT1 (N1945, N1934);
xor XOR2 (N1946, N1928, N1557);
and AND4 (N1947, N1944, N1353, N1328, N816);
xor XOR2 (N1948, N1930, N1693);
xor XOR2 (N1949, N1926, N1295);
xor XOR2 (N1950, N1948, N1546);
nor NOR3 (N1951, N1950, N370, N57);
buf BUF1 (N1952, N1941);
and AND2 (N1953, N1945, N1853);
nand NAND3 (N1954, N1952, N833, N334);
buf BUF1 (N1955, N1939);
or OR4 (N1956, N1949, N1328, N1820, N92);
buf BUF1 (N1957, N1955);
and AND4 (N1958, N1951, N1576, N1180, N1601);
nand NAND3 (N1959, N1953, N159, N571);
and AND4 (N1960, N1959, N149, N745, N753);
or OR4 (N1961, N1940, N400, N1384, N962);
xor XOR2 (N1962, N1954, N1763);
xor XOR2 (N1963, N1957, N772);
and AND4 (N1964, N1946, N1113, N1259, N323);
nor NOR4 (N1965, N1961, N638, N1244, N1358);
xor XOR2 (N1966, N1956, N1640);
nor NOR3 (N1967, N1942, N863, N302);
nand NAND3 (N1968, N1966, N1005, N1927);
buf BUF1 (N1969, N1963);
and AND3 (N1970, N1964, N1186, N1174);
not NOT1 (N1971, N1958);
nor NOR2 (N1972, N1947, N282);
not NOT1 (N1973, N1968);
buf BUF1 (N1974, N1969);
nand NAND4 (N1975, N1971, N1445, N1510, N770);
nor NOR2 (N1976, N1960, N108);
nor NOR4 (N1977, N1976, N983, N1415, N94);
buf BUF1 (N1978, N1962);
not NOT1 (N1979, N1974);
nor NOR4 (N1980, N1965, N817, N1700, N1179);
not NOT1 (N1981, N1943);
not NOT1 (N1982, N1977);
nand NAND2 (N1983, N1970, N58);
or OR4 (N1984, N1981, N1276, N1320, N470);
and AND4 (N1985, N1984, N707, N548, N709);
nor NOR2 (N1986, N1978, N1549);
xor XOR2 (N1987, N1983, N327);
or OR3 (N1988, N1975, N471, N294);
xor XOR2 (N1989, N1982, N619);
not NOT1 (N1990, N1980);
nor NOR3 (N1991, N1989, N1843, N1742);
nand NAND2 (N1992, N1972, N408);
or OR3 (N1993, N1973, N1971, N685);
or OR4 (N1994, N1985, N1508, N1052, N698);
buf BUF1 (N1995, N1994);
and AND2 (N1996, N1993, N1972);
xor XOR2 (N1997, N1995, N1145);
or OR4 (N1998, N1991, N1401, N1036, N1363);
nor NOR4 (N1999, N1990, N1902, N1631, N1010);
and AND4 (N2000, N1987, N883, N1677, N1150);
xor XOR2 (N2001, N1997, N1743);
buf BUF1 (N2002, N1996);
nor NOR4 (N2003, N1992, N1960, N1390, N491);
and AND4 (N2004, N2002, N1200, N1660, N1457);
not NOT1 (N2005, N2003);
buf BUF1 (N2006, N1988);
not NOT1 (N2007, N1967);
nor NOR3 (N2008, N1999, N1211, N525);
nor NOR3 (N2009, N2007, N1036, N306);
or OR3 (N2010, N2001, N689, N1756);
nand NAND4 (N2011, N2004, N196, N18, N340);
buf BUF1 (N2012, N1979);
xor XOR2 (N2013, N2005, N1203);
nor NOR2 (N2014, N2013, N1790);
buf BUF1 (N2015, N2014);
not NOT1 (N2016, N2015);
buf BUF1 (N2017, N2016);
buf BUF1 (N2018, N1986);
xor XOR2 (N2019, N2012, N1759);
buf BUF1 (N2020, N2017);
and AND3 (N2021, N2020, N1387, N1833);
nor NOR2 (N2022, N2019, N221);
and AND2 (N2023, N2009, N1456);
xor XOR2 (N2024, N2008, N1067);
nand NAND2 (N2025, N2022, N1874);
and AND2 (N2026, N2025, N1617);
or OR4 (N2027, N2006, N715, N86, N1209);
nand NAND3 (N2028, N2026, N757, N1970);
not NOT1 (N2029, N2010);
buf BUF1 (N2030, N2023);
or OR3 (N2031, N2000, N167, N673);
nor NOR2 (N2032, N1998, N932);
xor XOR2 (N2033, N2028, N534);
not NOT1 (N2034, N2011);
buf BUF1 (N2035, N2024);
not NOT1 (N2036, N2032);
not NOT1 (N2037, N2027);
xor XOR2 (N2038, N2029, N1437);
and AND2 (N2039, N2038, N1418);
not NOT1 (N2040, N2033);
xor XOR2 (N2041, N2037, N1518);
nor NOR4 (N2042, N2035, N1596, N358, N950);
not NOT1 (N2043, N2018);
buf BUF1 (N2044, N2043);
nor NOR4 (N2045, N2034, N1985, N1980, N1050);
nor NOR4 (N2046, N2041, N1386, N223, N1991);
buf BUF1 (N2047, N2021);
not NOT1 (N2048, N2046);
or OR4 (N2049, N2039, N1334, N1645, N1382);
xor XOR2 (N2050, N2031, N1190);
nor NOR4 (N2051, N2050, N147, N656, N741);
nor NOR2 (N2052, N2036, N471);
or OR2 (N2053, N2049, N780);
buf BUF1 (N2054, N2042);
not NOT1 (N2055, N2054);
nor NOR3 (N2056, N2047, N1952, N1617);
buf BUF1 (N2057, N2053);
buf BUF1 (N2058, N2040);
not NOT1 (N2059, N2048);
or OR3 (N2060, N2055, N347, N1045);
nor NOR4 (N2061, N2045, N1233, N1806, N281);
buf BUF1 (N2062, N2060);
or OR2 (N2063, N2062, N411);
and AND3 (N2064, N2056, N713, N1843);
nand NAND4 (N2065, N2061, N429, N342, N1732);
xor XOR2 (N2066, N2065, N1056);
or OR3 (N2067, N2058, N1212, N1029);
nand NAND3 (N2068, N2052, N1068, N1256);
nand NAND4 (N2069, N2030, N1339, N1875, N1472);
or OR4 (N2070, N2067, N308, N2043, N1097);
or OR2 (N2071, N2059, N748);
not NOT1 (N2072, N2064);
nand NAND3 (N2073, N2044, N1540, N1954);
or OR4 (N2074, N2073, N1732, N1386, N39);
nor NOR2 (N2075, N2057, N658);
nand NAND4 (N2076, N2070, N2019, N212, N735);
nand NAND3 (N2077, N2063, N274, N1704);
xor XOR2 (N2078, N2069, N850);
or OR3 (N2079, N2074, N429, N1834);
or OR3 (N2080, N2068, N1925, N1218);
or OR4 (N2081, N2071, N371, N1172, N412);
xor XOR2 (N2082, N2051, N594);
buf BUF1 (N2083, N2080);
nand NAND4 (N2084, N2078, N1287, N1872, N1656);
xor XOR2 (N2085, N2084, N702);
nand NAND4 (N2086, N2072, N477, N653, N981);
nor NOR3 (N2087, N2075, N782, N840);
not NOT1 (N2088, N2086);
buf BUF1 (N2089, N2088);
not NOT1 (N2090, N2082);
not NOT1 (N2091, N2087);
and AND2 (N2092, N2085, N1627);
xor XOR2 (N2093, N2092, N1191);
nor NOR3 (N2094, N2077, N367, N1777);
or OR3 (N2095, N2090, N1342, N882);
xor XOR2 (N2096, N2089, N466);
or OR4 (N2097, N2076, N1185, N840, N1728);
buf BUF1 (N2098, N2083);
and AND2 (N2099, N2081, N1738);
and AND3 (N2100, N2094, N1232, N1355);
nand NAND3 (N2101, N2091, N702, N629);
or OR3 (N2102, N2093, N763, N318);
nand NAND2 (N2103, N2096, N681);
buf BUF1 (N2104, N2079);
nand NAND4 (N2105, N2104, N1673, N1419, N459);
not NOT1 (N2106, N2100);
and AND4 (N2107, N2106, N2102, N1916, N724);
or OR2 (N2108, N1736, N1503);
not NOT1 (N2109, N2097);
nor NOR4 (N2110, N2105, N1624, N459, N1857);
nand NAND3 (N2111, N2107, N413, N815);
not NOT1 (N2112, N2109);
not NOT1 (N2113, N2111);
buf BUF1 (N2114, N2113);
buf BUF1 (N2115, N2112);
and AND4 (N2116, N2114, N1314, N762, N1097);
nand NAND2 (N2117, N2095, N378);
nor NOR3 (N2118, N2101, N1882, N2074);
or OR3 (N2119, N2103, N647, N1833);
nand NAND2 (N2120, N2117, N458);
or OR4 (N2121, N2118, N1282, N939, N982);
or OR4 (N2122, N2116, N455, N1866, N1146);
or OR4 (N2123, N2066, N565, N793, N1332);
or OR3 (N2124, N2119, N1520, N788);
buf BUF1 (N2125, N2098);
or OR3 (N2126, N2123, N149, N1508);
nand NAND2 (N2127, N2122, N1312);
xor XOR2 (N2128, N2120, N896);
and AND3 (N2129, N2110, N1161, N1553);
xor XOR2 (N2130, N2121, N510);
nand NAND2 (N2131, N2126, N1424);
or OR2 (N2132, N2124, N1886);
buf BUF1 (N2133, N2128);
nand NAND2 (N2134, N2130, N1902);
buf BUF1 (N2135, N2115);
nor NOR3 (N2136, N2131, N257, N894);
or OR4 (N2137, N2136, N1681, N1022, N977);
nor NOR3 (N2138, N2127, N1039, N1977);
or OR3 (N2139, N2129, N885, N244);
buf BUF1 (N2140, N2132);
not NOT1 (N2141, N2140);
not NOT1 (N2142, N2139);
nor NOR2 (N2143, N2142, N143);
xor XOR2 (N2144, N2108, N1992);
and AND4 (N2145, N2135, N1071, N1977, N608);
nor NOR4 (N2146, N2141, N1120, N90, N1528);
not NOT1 (N2147, N2134);
buf BUF1 (N2148, N2146);
nor NOR4 (N2149, N2143, N318, N1752, N111);
xor XOR2 (N2150, N2125, N496);
nor NOR4 (N2151, N2149, N1730, N1513, N965);
not NOT1 (N2152, N2133);
buf BUF1 (N2153, N2144);
nand NAND4 (N2154, N2145, N882, N1781, N1822);
nand NAND2 (N2155, N2152, N105);
or OR2 (N2156, N2155, N412);
xor XOR2 (N2157, N2148, N149);
xor XOR2 (N2158, N2099, N1389);
not NOT1 (N2159, N2158);
xor XOR2 (N2160, N2151, N1020);
buf BUF1 (N2161, N2153);
buf BUF1 (N2162, N2150);
xor XOR2 (N2163, N2138, N1060);
buf BUF1 (N2164, N2161);
xor XOR2 (N2165, N2164, N1846);
xor XOR2 (N2166, N2162, N1405);
buf BUF1 (N2167, N2166);
buf BUF1 (N2168, N2167);
or OR3 (N2169, N2154, N1303, N634);
and AND3 (N2170, N2137, N1143, N2014);
or OR4 (N2171, N2165, N1401, N1176, N1230);
or OR3 (N2172, N2170, N1921, N1427);
not NOT1 (N2173, N2168);
not NOT1 (N2174, N2172);
not NOT1 (N2175, N2159);
buf BUF1 (N2176, N2171);
nor NOR4 (N2177, N2175, N2155, N1023, N984);
nor NOR3 (N2178, N2147, N1874, N168);
buf BUF1 (N2179, N2173);
nor NOR2 (N2180, N2179, N1783);
buf BUF1 (N2181, N2169);
or OR2 (N2182, N2160, N592);
and AND2 (N2183, N2157, N1681);
buf BUF1 (N2184, N2181);
buf BUF1 (N2185, N2178);
not NOT1 (N2186, N2184);
not NOT1 (N2187, N2182);
or OR3 (N2188, N2183, N2123, N45);
xor XOR2 (N2189, N2188, N1947);
nand NAND2 (N2190, N2174, N361);
buf BUF1 (N2191, N2185);
nor NOR3 (N2192, N2187, N1899, N1385);
nor NOR4 (N2193, N2176, N1516, N1397, N39);
nand NAND2 (N2194, N2193, N172);
nand NAND3 (N2195, N2190, N138, N912);
and AND3 (N2196, N2192, N1932, N1743);
buf BUF1 (N2197, N2194);
or OR4 (N2198, N2195, N569, N339, N2150);
buf BUF1 (N2199, N2191);
not NOT1 (N2200, N2186);
xor XOR2 (N2201, N2196, N1962);
xor XOR2 (N2202, N2199, N979);
xor XOR2 (N2203, N2198, N2180);
nand NAND2 (N2204, N501, N1875);
xor XOR2 (N2205, N2156, N1621);
xor XOR2 (N2206, N2204, N109);
and AND4 (N2207, N2189, N44, N1212, N907);
nor NOR3 (N2208, N2207, N1173, N1044);
not NOT1 (N2209, N2206);
nor NOR4 (N2210, N2197, N1724, N1101, N329);
xor XOR2 (N2211, N2208, N1823);
nand NAND4 (N2212, N2163, N1943, N391, N70);
or OR2 (N2213, N2177, N1872);
buf BUF1 (N2214, N2211);
buf BUF1 (N2215, N2203);
buf BUF1 (N2216, N2210);
buf BUF1 (N2217, N2209);
and AND3 (N2218, N2215, N1956, N1570);
not NOT1 (N2219, N2213);
buf BUF1 (N2220, N2218);
and AND4 (N2221, N2201, N2155, N700, N1443);
and AND4 (N2222, N2216, N67, N1014, N220);
or OR2 (N2223, N2202, N1524);
buf BUF1 (N2224, N2205);
xor XOR2 (N2225, N2214, N912);
or OR4 (N2226, N2221, N332, N374, N158);
and AND4 (N2227, N2224, N2081, N1315, N1371);
xor XOR2 (N2228, N2226, N608);
and AND3 (N2229, N2222, N1073, N731);
buf BUF1 (N2230, N2223);
not NOT1 (N2231, N2217);
nor NOR4 (N2232, N2219, N1815, N315, N1910);
nand NAND2 (N2233, N2230, N1587);
and AND4 (N2234, N2228, N1947, N884, N1854);
buf BUF1 (N2235, N2200);
nand NAND4 (N2236, N2231, N866, N299, N1357);
buf BUF1 (N2237, N2235);
or OR2 (N2238, N2227, N636);
and AND4 (N2239, N2236, N928, N957, N1732);
or OR4 (N2240, N2237, N777, N386, N1130);
nand NAND2 (N2241, N2229, N1537);
and AND3 (N2242, N2212, N371, N940);
nor NOR4 (N2243, N2242, N1670, N338, N1615);
buf BUF1 (N2244, N2241);
nand NAND2 (N2245, N2243, N784);
buf BUF1 (N2246, N2232);
buf BUF1 (N2247, N2220);
buf BUF1 (N2248, N2234);
xor XOR2 (N2249, N2245, N1005);
nand NAND4 (N2250, N2249, N1326, N1907, N2227);
nor NOR4 (N2251, N2248, N2157, N686, N341);
or OR4 (N2252, N2244, N1647, N102, N10);
buf BUF1 (N2253, N2225);
not NOT1 (N2254, N2253);
nand NAND2 (N2255, N2254, N739);
not NOT1 (N2256, N2240);
nor NOR4 (N2257, N2238, N1524, N859, N1473);
or OR4 (N2258, N2257, N1473, N1864, N990);
buf BUF1 (N2259, N2256);
nand NAND2 (N2260, N2259, N217);
nor NOR2 (N2261, N2247, N528);
not NOT1 (N2262, N2261);
or OR2 (N2263, N2252, N2247);
nand NAND2 (N2264, N2233, N1885);
not NOT1 (N2265, N2260);
or OR2 (N2266, N2265, N652);
or OR2 (N2267, N2263, N1118);
nand NAND3 (N2268, N2246, N1677, N615);
nor NOR4 (N2269, N2262, N184, N1131, N1505);
nor NOR4 (N2270, N2269, N669, N1429, N2233);
buf BUF1 (N2271, N2264);
nor NOR4 (N2272, N2251, N575, N399, N424);
or OR3 (N2273, N2268, N624, N1350);
buf BUF1 (N2274, N2270);
xor XOR2 (N2275, N2271, N1954);
nor NOR3 (N2276, N2239, N1960, N383);
xor XOR2 (N2277, N2255, N1051);
xor XOR2 (N2278, N2277, N266);
xor XOR2 (N2279, N2274, N369);
and AND3 (N2280, N2258, N1507, N169);
xor XOR2 (N2281, N2276, N1204);
buf BUF1 (N2282, N2273);
nor NOR2 (N2283, N2275, N1906);
buf BUF1 (N2284, N2279);
and AND2 (N2285, N2283, N2096);
nand NAND3 (N2286, N2280, N926, N1900);
and AND3 (N2287, N2267, N533, N1726);
nand NAND2 (N2288, N2287, N2081);
and AND4 (N2289, N2250, N1747, N129, N1281);
or OR2 (N2290, N2289, N2223);
buf BUF1 (N2291, N2282);
nand NAND3 (N2292, N2281, N784, N2183);
nor NOR4 (N2293, N2286, N1288, N894, N1113);
xor XOR2 (N2294, N2285, N759);
or OR3 (N2295, N2266, N1144, N783);
and AND2 (N2296, N2284, N14);
or OR3 (N2297, N2290, N1169, N971);
and AND3 (N2298, N2294, N839, N1931);
or OR2 (N2299, N2288, N1570);
xor XOR2 (N2300, N2295, N1135);
buf BUF1 (N2301, N2272);
xor XOR2 (N2302, N2298, N292);
and AND3 (N2303, N2299, N1861, N644);
buf BUF1 (N2304, N2296);
or OR2 (N2305, N2303, N490);
nor NOR2 (N2306, N2291, N686);
or OR2 (N2307, N2306, N500);
or OR3 (N2308, N2300, N1108, N877);
or OR2 (N2309, N2278, N858);
buf BUF1 (N2310, N2293);
or OR2 (N2311, N2305, N920);
nand NAND2 (N2312, N2292, N993);
nand NAND3 (N2313, N2302, N1188, N1151);
xor XOR2 (N2314, N2311, N1462);
buf BUF1 (N2315, N2308);
not NOT1 (N2316, N2307);
not NOT1 (N2317, N2297);
not NOT1 (N2318, N2304);
buf BUF1 (N2319, N2316);
buf BUF1 (N2320, N2315);
or OR4 (N2321, N2301, N2193, N1781, N2146);
xor XOR2 (N2322, N2312, N1831);
buf BUF1 (N2323, N2313);
buf BUF1 (N2324, N2319);
not NOT1 (N2325, N2322);
and AND3 (N2326, N2314, N2270, N101);
not NOT1 (N2327, N2320);
xor XOR2 (N2328, N2323, N297);
xor XOR2 (N2329, N2328, N1228);
not NOT1 (N2330, N2317);
and AND2 (N2331, N2324, N159);
and AND2 (N2332, N2325, N1147);
and AND2 (N2333, N2327, N2045);
nor NOR2 (N2334, N2333, N2153);
nand NAND2 (N2335, N2330, N336);
or OR4 (N2336, N2329, N1307, N1299, N1616);
nor NOR4 (N2337, N2309, N140, N2239, N244);
nor NOR3 (N2338, N2337, N1343, N1584);
buf BUF1 (N2339, N2326);
or OR2 (N2340, N2336, N1838);
buf BUF1 (N2341, N2310);
nor NOR2 (N2342, N2318, N2014);
buf BUF1 (N2343, N2342);
xor XOR2 (N2344, N2334, N654);
not NOT1 (N2345, N2341);
xor XOR2 (N2346, N2344, N186);
and AND2 (N2347, N2340, N2318);
buf BUF1 (N2348, N2321);
buf BUF1 (N2349, N2332);
buf BUF1 (N2350, N2346);
and AND4 (N2351, N2347, N574, N1868, N190);
nor NOR4 (N2352, N2348, N474, N886, N1608);
or OR2 (N2353, N2352, N1581);
xor XOR2 (N2354, N2338, N1176);
buf BUF1 (N2355, N2335);
and AND3 (N2356, N2351, N1018, N119);
nand NAND4 (N2357, N2345, N1839, N2230, N675);
buf BUF1 (N2358, N2349);
nor NOR2 (N2359, N2358, N1112);
xor XOR2 (N2360, N2350, N469);
buf BUF1 (N2361, N2354);
or OR3 (N2362, N2331, N366, N386);
nand NAND2 (N2363, N2339, N1875);
and AND3 (N2364, N2353, N33, N521);
nand NAND2 (N2365, N2343, N641);
nand NAND2 (N2366, N2364, N1546);
xor XOR2 (N2367, N2363, N287);
not NOT1 (N2368, N2366);
xor XOR2 (N2369, N2360, N1183);
not NOT1 (N2370, N2356);
and AND2 (N2371, N2367, N1179);
or OR2 (N2372, N2357, N1354);
nand NAND2 (N2373, N2368, N1944);
xor XOR2 (N2374, N2361, N1643);
xor XOR2 (N2375, N2371, N1173);
not NOT1 (N2376, N2375);
nor NOR2 (N2377, N2359, N2197);
buf BUF1 (N2378, N2373);
not NOT1 (N2379, N2370);
buf BUF1 (N2380, N2379);
or OR3 (N2381, N2378, N2067, N969);
or OR2 (N2382, N2381, N2012);
buf BUF1 (N2383, N2355);
or OR4 (N2384, N2365, N2035, N561, N1932);
not NOT1 (N2385, N2382);
and AND3 (N2386, N2362, N541, N995);
not NOT1 (N2387, N2380);
not NOT1 (N2388, N2386);
not NOT1 (N2389, N2377);
or OR4 (N2390, N2384, N634, N707, N1199);
not NOT1 (N2391, N2385);
xor XOR2 (N2392, N2387, N1486);
not NOT1 (N2393, N2374);
nor NOR3 (N2394, N2376, N1167, N932);
buf BUF1 (N2395, N2390);
nand NAND2 (N2396, N2383, N414);
xor XOR2 (N2397, N2396, N333);
not NOT1 (N2398, N2394);
buf BUF1 (N2399, N2393);
or OR3 (N2400, N2392, N1244, N435);
not NOT1 (N2401, N2388);
not NOT1 (N2402, N2400);
not NOT1 (N2403, N2369);
or OR4 (N2404, N2403, N689, N248, N698);
nand NAND2 (N2405, N2372, N1669);
nor NOR3 (N2406, N2401, N1236, N1521);
nor NOR3 (N2407, N2389, N978, N2277);
and AND4 (N2408, N2395, N1673, N1113, N101);
or OR2 (N2409, N2397, N338);
and AND3 (N2410, N2406, N702, N2092);
and AND4 (N2411, N2409, N582, N306, N1480);
not NOT1 (N2412, N2404);
buf BUF1 (N2413, N2391);
nand NAND2 (N2414, N2412, N379);
and AND2 (N2415, N2408, N1849);
and AND4 (N2416, N2410, N2057, N1615, N2408);
xor XOR2 (N2417, N2414, N1124);
not NOT1 (N2418, N2416);
xor XOR2 (N2419, N2411, N2393);
not NOT1 (N2420, N2413);
buf BUF1 (N2421, N2405);
xor XOR2 (N2422, N2407, N318);
nand NAND2 (N2423, N2420, N450);
buf BUF1 (N2424, N2418);
or OR4 (N2425, N2421, N1130, N406, N1624);
or OR4 (N2426, N2425, N1711, N1765, N960);
xor XOR2 (N2427, N2417, N147);
not NOT1 (N2428, N2426);
nand NAND4 (N2429, N2402, N359, N1034, N1236);
and AND3 (N2430, N2415, N289, N749);
not NOT1 (N2431, N2419);
nand NAND4 (N2432, N2398, N677, N426, N266);
xor XOR2 (N2433, N2429, N322);
not NOT1 (N2434, N2431);
nand NAND3 (N2435, N2428, N711, N643);
buf BUF1 (N2436, N2433);
or OR2 (N2437, N2424, N2402);
not NOT1 (N2438, N2430);
and AND2 (N2439, N2437, N104);
and AND2 (N2440, N2439, N1327);
or OR4 (N2441, N2422, N1391, N2418, N401);
xor XOR2 (N2442, N2423, N863);
and AND2 (N2443, N2438, N369);
buf BUF1 (N2444, N2442);
or OR3 (N2445, N2399, N1060, N1689);
nor NOR4 (N2446, N2445, N517, N2293, N339);
not NOT1 (N2447, N2443);
or OR2 (N2448, N2435, N372);
and AND2 (N2449, N2444, N2232);
or OR2 (N2450, N2447, N105);
or OR2 (N2451, N2441, N2305);
and AND4 (N2452, N2449, N2187, N2208, N2343);
or OR4 (N2453, N2432, N762, N77, N1839);
buf BUF1 (N2454, N2427);
not NOT1 (N2455, N2440);
not NOT1 (N2456, N2454);
buf BUF1 (N2457, N2451);
nor NOR3 (N2458, N2452, N1511, N414);
not NOT1 (N2459, N2436);
or OR3 (N2460, N2448, N1555, N2150);
buf BUF1 (N2461, N2460);
nor NOR3 (N2462, N2456, N78, N1079);
xor XOR2 (N2463, N2457, N594);
not NOT1 (N2464, N2455);
xor XOR2 (N2465, N2446, N1459);
xor XOR2 (N2466, N2459, N2052);
nor NOR3 (N2467, N2458, N198, N1596);
and AND2 (N2468, N2450, N1600);
nor NOR2 (N2469, N2468, N1527);
and AND2 (N2470, N2463, N1563);
nand NAND2 (N2471, N2467, N1219);
not NOT1 (N2472, N2453);
nand NAND4 (N2473, N2469, N1411, N869, N408);
nand NAND2 (N2474, N2464, N2275);
not NOT1 (N2475, N2465);
and AND2 (N2476, N2462, N144);
not NOT1 (N2477, N2473);
nor NOR2 (N2478, N2474, N351);
xor XOR2 (N2479, N2434, N1461);
nor NOR3 (N2480, N2461, N1893, N1653);
xor XOR2 (N2481, N2472, N515);
or OR3 (N2482, N2478, N1252, N1727);
and AND2 (N2483, N2470, N499);
buf BUF1 (N2484, N2480);
nand NAND3 (N2485, N2476, N2158, N1247);
buf BUF1 (N2486, N2477);
nor NOR4 (N2487, N2482, N601, N839, N1749);
nand NAND4 (N2488, N2466, N1689, N1774, N1764);
xor XOR2 (N2489, N2475, N1384);
buf BUF1 (N2490, N2484);
or OR2 (N2491, N2485, N2466);
not NOT1 (N2492, N2471);
not NOT1 (N2493, N2483);
nand NAND2 (N2494, N2490, N1134);
xor XOR2 (N2495, N2486, N2320);
nor NOR3 (N2496, N2481, N948, N1774);
nand NAND2 (N2497, N2496, N1625);
buf BUF1 (N2498, N2487);
xor XOR2 (N2499, N2493, N1949);
buf BUF1 (N2500, N2488);
xor XOR2 (N2501, N2495, N2409);
nand NAND3 (N2502, N2498, N579, N2199);
nand NAND2 (N2503, N2494, N499);
xor XOR2 (N2504, N2489, N1956);
not NOT1 (N2505, N2497);
or OR3 (N2506, N2499, N1973, N1889);
and AND4 (N2507, N2506, N1786, N112, N1822);
not NOT1 (N2508, N2501);
nand NAND2 (N2509, N2491, N280);
nand NAND4 (N2510, N2503, N882, N2295, N2394);
nor NOR4 (N2511, N2505, N2490, N1189, N2419);
xor XOR2 (N2512, N2500, N2451);
nor NOR4 (N2513, N2507, N1835, N2263, N1860);
not NOT1 (N2514, N2511);
nor NOR4 (N2515, N2479, N139, N1803, N2027);
buf BUF1 (N2516, N2508);
and AND2 (N2517, N2512, N1368);
buf BUF1 (N2518, N2516);
or OR2 (N2519, N2514, N2138);
xor XOR2 (N2520, N2517, N569);
xor XOR2 (N2521, N2504, N1276);
nand NAND3 (N2522, N2509, N495, N1535);
xor XOR2 (N2523, N2510, N221);
xor XOR2 (N2524, N2520, N1967);
buf BUF1 (N2525, N2523);
buf BUF1 (N2526, N2518);
buf BUF1 (N2527, N2519);
or OR3 (N2528, N2502, N1957, N1171);
and AND2 (N2529, N2527, N1155);
xor XOR2 (N2530, N2513, N2398);
nand NAND3 (N2531, N2515, N2324, N1149);
buf BUF1 (N2532, N2526);
and AND3 (N2533, N2525, N575, N1466);
nor NOR2 (N2534, N2492, N2064);
nor NOR2 (N2535, N2533, N2072);
or OR2 (N2536, N2522, N581);
nand NAND3 (N2537, N2536, N1052, N2138);
nand NAND4 (N2538, N2531, N73, N9, N1340);
not NOT1 (N2539, N2528);
or OR4 (N2540, N2524, N1392, N1420, N2017);
not NOT1 (N2541, N2534);
not NOT1 (N2542, N2537);
or OR2 (N2543, N2532, N8);
buf BUF1 (N2544, N2542);
buf BUF1 (N2545, N2529);
buf BUF1 (N2546, N2538);
or OR4 (N2547, N2541, N1898, N1104, N171);
not NOT1 (N2548, N2535);
not NOT1 (N2549, N2544);
xor XOR2 (N2550, N2549, N1117);
and AND3 (N2551, N2540, N780, N1444);
xor XOR2 (N2552, N2551, N783);
buf BUF1 (N2553, N2546);
buf BUF1 (N2554, N2548);
or OR3 (N2555, N2543, N2375, N2126);
xor XOR2 (N2556, N2553, N150);
nor NOR2 (N2557, N2547, N1404);
or OR4 (N2558, N2545, N2120, N504, N610);
not NOT1 (N2559, N2554);
buf BUF1 (N2560, N2558);
nor NOR4 (N2561, N2556, N1789, N1490, N456);
nand NAND4 (N2562, N2521, N788, N1316, N2465);
not NOT1 (N2563, N2561);
and AND4 (N2564, N2560, N1537, N1719, N2242);
nand NAND4 (N2565, N2539, N2422, N884, N963);
nand NAND2 (N2566, N2565, N2269);
not NOT1 (N2567, N2552);
buf BUF1 (N2568, N2557);
xor XOR2 (N2569, N2564, N1801);
buf BUF1 (N2570, N2568);
nor NOR2 (N2571, N2550, N208);
xor XOR2 (N2572, N2530, N2198);
not NOT1 (N2573, N2559);
or OR2 (N2574, N2570, N1354);
nor NOR3 (N2575, N2569, N546, N1429);
nor NOR2 (N2576, N2571, N1541);
buf BUF1 (N2577, N2566);
nor NOR4 (N2578, N2576, N1260, N10, N828);
nand NAND2 (N2579, N2567, N693);
and AND3 (N2580, N2577, N2219, N276);
nand NAND4 (N2581, N2555, N214, N500, N37);
not NOT1 (N2582, N2580);
not NOT1 (N2583, N2574);
buf BUF1 (N2584, N2572);
xor XOR2 (N2585, N2584, N887);
not NOT1 (N2586, N2585);
nor NOR3 (N2587, N2562, N1438, N733);
or OR3 (N2588, N2563, N114, N93);
nor NOR4 (N2589, N2582, N1697, N1754, N2366);
xor XOR2 (N2590, N2581, N2098);
xor XOR2 (N2591, N2589, N2569);
nand NAND3 (N2592, N2586, N207, N1483);
not NOT1 (N2593, N2592);
or OR4 (N2594, N2573, N1774, N967, N1827);
and AND3 (N2595, N2594, N2153, N778);
not NOT1 (N2596, N2593);
and AND2 (N2597, N2590, N1315);
buf BUF1 (N2598, N2583);
not NOT1 (N2599, N2579);
nand NAND4 (N2600, N2598, N455, N98, N356);
not NOT1 (N2601, N2591);
or OR3 (N2602, N2601, N2031, N1944);
nand NAND2 (N2603, N2600, N1829);
nor NOR4 (N2604, N2602, N1720, N1914, N601);
and AND2 (N2605, N2587, N2478);
not NOT1 (N2606, N2578);
buf BUF1 (N2607, N2597);
not NOT1 (N2608, N2606);
xor XOR2 (N2609, N2603, N2313);
not NOT1 (N2610, N2596);
xor XOR2 (N2611, N2608, N2068);
nand NAND3 (N2612, N2607, N768, N860);
not NOT1 (N2613, N2575);
or OR2 (N2614, N2611, N1975);
buf BUF1 (N2615, N2605);
buf BUF1 (N2616, N2610);
nand NAND4 (N2617, N2588, N2079, N894, N981);
buf BUF1 (N2618, N2604);
buf BUF1 (N2619, N2609);
not NOT1 (N2620, N2595);
nand NAND4 (N2621, N2613, N1620, N933, N989);
xor XOR2 (N2622, N2614, N1344);
or OR3 (N2623, N2620, N962, N299);
xor XOR2 (N2624, N2599, N386);
or OR2 (N2625, N2623, N2518);
buf BUF1 (N2626, N2622);
xor XOR2 (N2627, N2624, N203);
nand NAND4 (N2628, N2616, N1429, N2531, N168);
xor XOR2 (N2629, N2628, N2031);
xor XOR2 (N2630, N2618, N928);
nor NOR4 (N2631, N2629, N2298, N2401, N945);
not NOT1 (N2632, N2612);
or OR4 (N2633, N2626, N2150, N2598, N1910);
xor XOR2 (N2634, N2631, N1773);
and AND4 (N2635, N2617, N517, N2238, N2214);
or OR2 (N2636, N2632, N1200);
nor NOR3 (N2637, N2619, N2559, N2049);
nor NOR2 (N2638, N2636, N2475);
nand NAND4 (N2639, N2627, N1760, N2079, N2373);
nand NAND3 (N2640, N2637, N530, N7);
nand NAND3 (N2641, N2630, N1883, N2036);
and AND3 (N2642, N2639, N1048, N1286);
nor NOR2 (N2643, N2634, N342);
xor XOR2 (N2644, N2625, N1703);
nor NOR4 (N2645, N2638, N746, N567, N310);
not NOT1 (N2646, N2645);
not NOT1 (N2647, N2635);
nor NOR2 (N2648, N2644, N1221);
buf BUF1 (N2649, N2646);
nand NAND4 (N2650, N2640, N38, N592, N525);
xor XOR2 (N2651, N2650, N1111);
or OR4 (N2652, N2648, N2376, N108, N1416);
nand NAND2 (N2653, N2633, N1284);
buf BUF1 (N2654, N2642);
xor XOR2 (N2655, N2641, N915);
nor NOR4 (N2656, N2652, N464, N1158, N1372);
not NOT1 (N2657, N2647);
xor XOR2 (N2658, N2656, N1444);
nand NAND3 (N2659, N2658, N2547, N788);
and AND3 (N2660, N2653, N91, N1754);
buf BUF1 (N2661, N2615);
not NOT1 (N2662, N2654);
not NOT1 (N2663, N2643);
xor XOR2 (N2664, N2657, N1339);
and AND3 (N2665, N2660, N2553, N2534);
nand NAND2 (N2666, N2665, N1374);
or OR3 (N2667, N2621, N894, N670);
nand NAND3 (N2668, N2649, N497, N2463);
nand NAND3 (N2669, N2661, N1758, N814);
not NOT1 (N2670, N2666);
and AND2 (N2671, N2667, N1926);
buf BUF1 (N2672, N2651);
not NOT1 (N2673, N2669);
xor XOR2 (N2674, N2655, N848);
nor NOR3 (N2675, N2662, N2340, N594);
nor NOR3 (N2676, N2668, N1476, N589);
nand NAND2 (N2677, N2673, N1101);
and AND2 (N2678, N2677, N402);
buf BUF1 (N2679, N2659);
xor XOR2 (N2680, N2675, N2458);
not NOT1 (N2681, N2663);
buf BUF1 (N2682, N2670);
nor NOR2 (N2683, N2678, N381);
and AND3 (N2684, N2682, N1692, N2393);
or OR2 (N2685, N2679, N977);
not NOT1 (N2686, N2684);
buf BUF1 (N2687, N2680);
nand NAND3 (N2688, N2672, N869, N2632);
or OR3 (N2689, N2687, N2402, N401);
xor XOR2 (N2690, N2671, N640);
buf BUF1 (N2691, N2688);
or OR4 (N2692, N2674, N843, N2125, N1741);
xor XOR2 (N2693, N2690, N165);
not NOT1 (N2694, N2686);
nand NAND4 (N2695, N2685, N1320, N666, N2635);
nand NAND4 (N2696, N2681, N382, N1022, N576);
nand NAND4 (N2697, N2683, N426, N1003, N1362);
nand NAND2 (N2698, N2692, N1460);
or OR4 (N2699, N2696, N1717, N1591, N1147);
xor XOR2 (N2700, N2697, N135);
xor XOR2 (N2701, N2700, N665);
and AND2 (N2702, N2691, N1217);
not NOT1 (N2703, N2699);
nand NAND2 (N2704, N2695, N255);
xor XOR2 (N2705, N2664, N213);
or OR3 (N2706, N2705, N6, N1043);
or OR2 (N2707, N2698, N1978);
not NOT1 (N2708, N2706);
not NOT1 (N2709, N2708);
not NOT1 (N2710, N2694);
nor NOR3 (N2711, N2702, N576, N702);
xor XOR2 (N2712, N2709, N418);
or OR2 (N2713, N2703, N1079);
and AND3 (N2714, N2707, N1296, N2482);
xor XOR2 (N2715, N2676, N937);
xor XOR2 (N2716, N2689, N2074);
or OR4 (N2717, N2693, N832, N2167, N1894);
buf BUF1 (N2718, N2713);
not NOT1 (N2719, N2716);
nor NOR4 (N2720, N2710, N310, N2680, N652);
nor NOR4 (N2721, N2704, N2011, N1501, N72);
buf BUF1 (N2722, N2717);
not NOT1 (N2723, N2720);
nor NOR2 (N2724, N2715, N1198);
or OR2 (N2725, N2719, N1759);
nand NAND2 (N2726, N2721, N2544);
or OR3 (N2727, N2711, N2079, N2225);
and AND4 (N2728, N2725, N2336, N86, N2250);
not NOT1 (N2729, N2724);
buf BUF1 (N2730, N2714);
nand NAND2 (N2731, N2701, N1857);
or OR3 (N2732, N2730, N2143, N667);
buf BUF1 (N2733, N2729);
not NOT1 (N2734, N2722);
nor NOR2 (N2735, N2726, N1179);
and AND4 (N2736, N2718, N1283, N500, N2442);
nor NOR2 (N2737, N2732, N242);
nand NAND3 (N2738, N2736, N1197, N2727);
and AND4 (N2739, N2572, N1942, N33, N895);
xor XOR2 (N2740, N2731, N2186);
or OR3 (N2741, N2739, N995, N800);
or OR3 (N2742, N2723, N2148, N848);
or OR2 (N2743, N2712, N594);
nand NAND4 (N2744, N2733, N1240, N2596, N2405);
and AND3 (N2745, N2737, N487, N520);
or OR2 (N2746, N2735, N2477);
not NOT1 (N2747, N2742);
buf BUF1 (N2748, N2728);
xor XOR2 (N2749, N2747, N2096);
or OR3 (N2750, N2749, N89, N1278);
not NOT1 (N2751, N2745);
not NOT1 (N2752, N2751);
and AND3 (N2753, N2738, N926, N152);
and AND4 (N2754, N2753, N1882, N2672, N1516);
or OR4 (N2755, N2734, N2134, N675, N1727);
nor NOR2 (N2756, N2750, N1221);
not NOT1 (N2757, N2748);
and AND4 (N2758, N2757, N1014, N1917, N1061);
not NOT1 (N2759, N2756);
not NOT1 (N2760, N2740);
xor XOR2 (N2761, N2741, N537);
buf BUF1 (N2762, N2755);
and AND2 (N2763, N2758, N2536);
and AND4 (N2764, N2761, N1984, N2009, N2532);
nand NAND2 (N2765, N2752, N715);
and AND3 (N2766, N2759, N1639, N453);
xor XOR2 (N2767, N2764, N38);
or OR3 (N2768, N2766, N1426, N1464);
not NOT1 (N2769, N2765);
nand NAND2 (N2770, N2768, N2115);
and AND2 (N2771, N2767, N1190);
not NOT1 (N2772, N2744);
nor NOR2 (N2773, N2754, N1240);
not NOT1 (N2774, N2772);
or OR3 (N2775, N2746, N2516, N524);
nand NAND2 (N2776, N2775, N1666);
nand NAND3 (N2777, N2770, N78, N225);
nor NOR4 (N2778, N2771, N335, N2746, N58);
nand NAND4 (N2779, N2760, N2017, N2292, N1189);
nand NAND2 (N2780, N2776, N1560);
buf BUF1 (N2781, N2762);
not NOT1 (N2782, N2780);
and AND3 (N2783, N2743, N2235, N1903);
and AND3 (N2784, N2769, N1206, N487);
buf BUF1 (N2785, N2777);
nor NOR2 (N2786, N2773, N564);
not NOT1 (N2787, N2763);
nand NAND3 (N2788, N2786, N1368, N2391);
buf BUF1 (N2789, N2787);
nor NOR2 (N2790, N2789, N1398);
nand NAND4 (N2791, N2784, N756, N1155, N2360);
nand NAND3 (N2792, N2783, N1118, N2667);
xor XOR2 (N2793, N2792, N1011);
buf BUF1 (N2794, N2793);
xor XOR2 (N2795, N2782, N1947);
nand NAND2 (N2796, N2778, N2030);
and AND3 (N2797, N2790, N888, N609);
nand NAND2 (N2798, N2779, N2585);
or OR3 (N2799, N2796, N664, N1625);
buf BUF1 (N2800, N2797);
nand NAND4 (N2801, N2800, N657, N3, N2451);
nand NAND4 (N2802, N2791, N2396, N533, N1924);
xor XOR2 (N2803, N2785, N934);
nand NAND2 (N2804, N2803, N1737);
and AND3 (N2805, N2799, N788, N290);
and AND2 (N2806, N2805, N1899);
buf BUF1 (N2807, N2806);
buf BUF1 (N2808, N2807);
not NOT1 (N2809, N2802);
xor XOR2 (N2810, N2808, N2024);
not NOT1 (N2811, N2801);
nor NOR3 (N2812, N2811, N1612, N2492);
nand NAND2 (N2813, N2804, N1702);
nand NAND3 (N2814, N2781, N119, N328);
not NOT1 (N2815, N2812);
buf BUF1 (N2816, N2794);
xor XOR2 (N2817, N2816, N70);
nor NOR2 (N2818, N2810, N2170);
buf BUF1 (N2819, N2788);
nor NOR2 (N2820, N2774, N1847);
xor XOR2 (N2821, N2819, N2238);
and AND2 (N2822, N2813, N1614);
buf BUF1 (N2823, N2820);
or OR2 (N2824, N2798, N1505);
nand NAND3 (N2825, N2818, N1188, N1509);
nor NOR2 (N2826, N2821, N844);
nand NAND3 (N2827, N2822, N612, N1088);
nor NOR4 (N2828, N2814, N686, N475, N2501);
nand NAND2 (N2829, N2825, N230);
nand NAND2 (N2830, N2823, N1460);
nand NAND4 (N2831, N2826, N1066, N1625, N113);
nor NOR2 (N2832, N2827, N2036);
or OR4 (N2833, N2829, N270, N2587, N1685);
or OR3 (N2834, N2795, N1958, N1460);
and AND4 (N2835, N2834, N909, N2823, N1892);
not NOT1 (N2836, N2824);
xor XOR2 (N2837, N2832, N2674);
not NOT1 (N2838, N2833);
or OR2 (N2839, N2815, N2084);
or OR4 (N2840, N2828, N1136, N2366, N516);
nand NAND2 (N2841, N2839, N1167);
not NOT1 (N2842, N2831);
nor NOR4 (N2843, N2817, N1283, N2236, N2732);
nor NOR3 (N2844, N2835, N1011, N1553);
buf BUF1 (N2845, N2840);
nand NAND2 (N2846, N2842, N2735);
or OR2 (N2847, N2846, N1213);
buf BUF1 (N2848, N2845);
nand NAND2 (N2849, N2837, N1199);
not NOT1 (N2850, N2838);
nor NOR2 (N2851, N2841, N637);
xor XOR2 (N2852, N2847, N1183);
and AND2 (N2853, N2844, N1120);
buf BUF1 (N2854, N2830);
and AND2 (N2855, N2848, N2473);
nand NAND4 (N2856, N2851, N45, N1631, N327);
and AND4 (N2857, N2809, N2672, N2206, N1009);
nand NAND3 (N2858, N2836, N1043, N902);
nand NAND4 (N2859, N2843, N524, N2330, N1967);
buf BUF1 (N2860, N2854);
or OR4 (N2861, N2849, N354, N688, N660);
nand NAND4 (N2862, N2853, N59, N2508, N2198);
not NOT1 (N2863, N2862);
xor XOR2 (N2864, N2863, N2612);
nand NAND2 (N2865, N2858, N1809);
xor XOR2 (N2866, N2855, N207);
and AND2 (N2867, N2850, N841);
nand NAND4 (N2868, N2857, N468, N1069, N1713);
and AND2 (N2869, N2861, N2671);
nor NOR2 (N2870, N2866, N30);
xor XOR2 (N2871, N2864, N1460);
nor NOR2 (N2872, N2860, N1927);
nand NAND4 (N2873, N2867, N2644, N1248, N310);
nor NOR4 (N2874, N2869, N993, N1806, N2725);
nor NOR2 (N2875, N2874, N1130);
not NOT1 (N2876, N2873);
and AND4 (N2877, N2871, N965, N2131, N2317);
nor NOR2 (N2878, N2868, N468);
not NOT1 (N2879, N2875);
buf BUF1 (N2880, N2872);
buf BUF1 (N2881, N2856);
xor XOR2 (N2882, N2879, N1554);
not NOT1 (N2883, N2870);
and AND3 (N2884, N2878, N1165, N2320);
not NOT1 (N2885, N2852);
nand NAND3 (N2886, N2880, N451, N2506);
nor NOR2 (N2887, N2876, N258);
nand NAND3 (N2888, N2877, N865, N320);
xor XOR2 (N2889, N2859, N339);
not NOT1 (N2890, N2889);
nor NOR3 (N2891, N2888, N825, N1514);
nor NOR4 (N2892, N2883, N39, N1533, N1180);
and AND4 (N2893, N2890, N2703, N296, N2458);
nor NOR4 (N2894, N2887, N2661, N2680, N1247);
or OR2 (N2895, N2894, N1394);
not NOT1 (N2896, N2895);
nor NOR2 (N2897, N2896, N1593);
xor XOR2 (N2898, N2882, N346);
or OR2 (N2899, N2885, N1538);
not NOT1 (N2900, N2886);
or OR4 (N2901, N2900, N2820, N1446, N1827);
nor NOR3 (N2902, N2865, N2032, N2623);
nor NOR2 (N2903, N2902, N937);
nand NAND3 (N2904, N2899, N2580, N2902);
and AND3 (N2905, N2898, N1859, N1562);
or OR2 (N2906, N2897, N144);
nor NOR3 (N2907, N2881, N2330, N2792);
or OR4 (N2908, N2891, N2196, N467, N1783);
or OR4 (N2909, N2892, N2337, N1871, N362);
or OR2 (N2910, N2901, N239);
nor NOR3 (N2911, N2904, N2109, N330);
nor NOR2 (N2912, N2907, N2024);
not NOT1 (N2913, N2905);
and AND4 (N2914, N2906, N656, N222, N1286);
nand NAND4 (N2915, N2913, N2868, N2412, N868);
nand NAND2 (N2916, N2915, N116);
buf BUF1 (N2917, N2884);
buf BUF1 (N2918, N2912);
nand NAND4 (N2919, N2908, N2621, N1531, N2910);
not NOT1 (N2920, N2814);
buf BUF1 (N2921, N2914);
nand NAND4 (N2922, N2920, N2298, N2152, N2292);
buf BUF1 (N2923, N2918);
and AND2 (N2924, N2922, N2644);
not NOT1 (N2925, N2903);
or OR3 (N2926, N2909, N2874, N372);
nand NAND3 (N2927, N2919, N104, N1063);
xor XOR2 (N2928, N2916, N78);
xor XOR2 (N2929, N2928, N1097);
nand NAND4 (N2930, N2921, N1222, N2603, N1032);
xor XOR2 (N2931, N2923, N464);
and AND2 (N2932, N2911, N821);
xor XOR2 (N2933, N2930, N1341);
and AND2 (N2934, N2927, N781);
or OR3 (N2935, N2924, N1728, N808);
xor XOR2 (N2936, N2925, N1462);
nor NOR4 (N2937, N2934, N133, N1024, N390);
nand NAND2 (N2938, N2929, N436);
or OR4 (N2939, N2935, N2219, N2906, N1271);
nand NAND2 (N2940, N2936, N2359);
not NOT1 (N2941, N2940);
nand NAND2 (N2942, N2917, N2866);
nand NAND2 (N2943, N2932, N2596);
and AND3 (N2944, N2926, N1805, N2738);
or OR2 (N2945, N2939, N142);
xor XOR2 (N2946, N2933, N80);
nand NAND3 (N2947, N2893, N2604, N685);
nand NAND2 (N2948, N2946, N1470);
xor XOR2 (N2949, N2944, N707);
not NOT1 (N2950, N2947);
nor NOR2 (N2951, N2937, N2251);
or OR2 (N2952, N2938, N1572);
buf BUF1 (N2953, N2950);
xor XOR2 (N2954, N2951, N1214);
nand NAND3 (N2955, N2952, N1171, N2435);
not NOT1 (N2956, N2954);
and AND4 (N2957, N2955, N1806, N225, N1353);
buf BUF1 (N2958, N2942);
and AND3 (N2959, N2943, N1123, N274);
not NOT1 (N2960, N2941);
buf BUF1 (N2961, N2949);
not NOT1 (N2962, N2945);
nor NOR3 (N2963, N2962, N506, N2084);
nor NOR3 (N2964, N2953, N1126, N2156);
xor XOR2 (N2965, N2963, N1349);
or OR3 (N2966, N2959, N2120, N2153);
xor XOR2 (N2967, N2948, N1601);
nand NAND4 (N2968, N2965, N1442, N1767, N366);
or OR2 (N2969, N2964, N421);
xor XOR2 (N2970, N2931, N764);
or OR3 (N2971, N2966, N1869, N2591);
and AND4 (N2972, N2961, N1252, N1083, N553);
xor XOR2 (N2973, N2960, N745);
nand NAND4 (N2974, N2957, N235, N378, N1837);
not NOT1 (N2975, N2956);
xor XOR2 (N2976, N2969, N1911);
buf BUF1 (N2977, N2968);
buf BUF1 (N2978, N2973);
nor NOR3 (N2979, N2971, N932, N1496);
and AND2 (N2980, N2976, N2224);
and AND3 (N2981, N2972, N990, N2082);
and AND2 (N2982, N2958, N522);
or OR4 (N2983, N2982, N1494, N9, N2524);
buf BUF1 (N2984, N2979);
or OR3 (N2985, N2983, N519, N641);
and AND2 (N2986, N2984, N2766);
nand NAND3 (N2987, N2967, N1922, N2404);
nor NOR3 (N2988, N2980, N1025, N725);
and AND4 (N2989, N2987, N1436, N390, N783);
buf BUF1 (N2990, N2974);
or OR2 (N2991, N2977, N2634);
not NOT1 (N2992, N2978);
nand NAND2 (N2993, N2991, N2719);
xor XOR2 (N2994, N2990, N1632);
and AND4 (N2995, N2985, N1455, N1369, N2231);
nor NOR2 (N2996, N2988, N1090);
and AND3 (N2997, N2996, N2447, N1085);
and AND2 (N2998, N2992, N1098);
nand NAND3 (N2999, N2995, N129, N712);
buf BUF1 (N3000, N2994);
nor NOR4 (N3001, N2970, N1831, N1433, N149);
buf BUF1 (N3002, N2999);
xor XOR2 (N3003, N2975, N1086);
xor XOR2 (N3004, N2981, N70);
or OR4 (N3005, N3003, N1968, N1859, N2468);
and AND2 (N3006, N2998, N1512);
or OR3 (N3007, N2989, N2650, N1142);
nor NOR4 (N3008, N3001, N2548, N1329, N1021);
and AND2 (N3009, N3002, N1918);
buf BUF1 (N3010, N2993);
buf BUF1 (N3011, N3000);
not NOT1 (N3012, N3011);
xor XOR2 (N3013, N2986, N523);
nor NOR2 (N3014, N2997, N175);
and AND4 (N3015, N3006, N2989, N2911, N760);
nand NAND4 (N3016, N3014, N1706, N2198, N1571);
or OR2 (N3017, N3005, N2767);
and AND2 (N3018, N3009, N211);
nor NOR3 (N3019, N3007, N268, N1574);
xor XOR2 (N3020, N3013, N1547);
nand NAND2 (N3021, N3008, N750);
nand NAND2 (N3022, N3010, N489);
buf BUF1 (N3023, N3021);
or OR3 (N3024, N3016, N2258, N2316);
not NOT1 (N3025, N3020);
buf BUF1 (N3026, N3019);
nand NAND2 (N3027, N3004, N129);
nor NOR3 (N3028, N3024, N2180, N2222);
xor XOR2 (N3029, N3018, N2171);
not NOT1 (N3030, N3015);
nor NOR2 (N3031, N3017, N402);
buf BUF1 (N3032, N3027);
xor XOR2 (N3033, N3026, N1155);
and AND3 (N3034, N3033, N827, N2705);
or OR4 (N3035, N3029, N2102, N491, N747);
nor NOR2 (N3036, N3028, N683);
or OR3 (N3037, N3032, N1313, N84);
not NOT1 (N3038, N3031);
or OR3 (N3039, N3023, N1332, N1563);
nand NAND4 (N3040, N3034, N431, N1819, N2100);
not NOT1 (N3041, N3022);
or OR2 (N3042, N3036, N1579);
or OR2 (N3043, N3030, N1363);
and AND3 (N3044, N3025, N2946, N2395);
not NOT1 (N3045, N3044);
and AND3 (N3046, N3037, N1863, N893);
not NOT1 (N3047, N3035);
nand NAND4 (N3048, N3038, N1532, N1146, N2163);
and AND2 (N3049, N3046, N2846);
or OR2 (N3050, N3047, N2800);
nand NAND2 (N3051, N3050, N2534);
not NOT1 (N3052, N3041);
not NOT1 (N3053, N3039);
or OR3 (N3054, N3042, N248, N1635);
and AND2 (N3055, N3040, N472);
not NOT1 (N3056, N3052);
and AND4 (N3057, N3055, N560, N102, N1779);
and AND2 (N3058, N3043, N2477);
nand NAND4 (N3059, N3045, N1426, N897, N2960);
and AND3 (N3060, N3053, N2386, N1144);
buf BUF1 (N3061, N3056);
xor XOR2 (N3062, N3058, N1785);
buf BUF1 (N3063, N3054);
or OR4 (N3064, N3063, N2136, N1214, N2505);
buf BUF1 (N3065, N3064);
nand NAND4 (N3066, N3059, N2405, N26, N249);
not NOT1 (N3067, N3062);
or OR3 (N3068, N3051, N1283, N1581);
or OR4 (N3069, N3049, N524, N735, N3066);
nand NAND4 (N3070, N1203, N1125, N472, N1053);
nor NOR4 (N3071, N3067, N101, N1357, N1496);
not NOT1 (N3072, N3069);
and AND4 (N3073, N3068, N1918, N1909, N2308);
and AND3 (N3074, N3065, N2957, N3065);
buf BUF1 (N3075, N3071);
and AND4 (N3076, N3060, N36, N667, N1037);
nand NAND3 (N3077, N3072, N942, N2021);
buf BUF1 (N3078, N3070);
or OR4 (N3079, N3048, N1606, N1654, N2549);
nand NAND4 (N3080, N3075, N751, N2713, N986);
buf BUF1 (N3081, N3057);
not NOT1 (N3082, N3074);
xor XOR2 (N3083, N3077, N555);
not NOT1 (N3084, N3081);
xor XOR2 (N3085, N3076, N223);
and AND3 (N3086, N3078, N1914, N1348);
and AND2 (N3087, N3073, N289);
xor XOR2 (N3088, N3084, N1735);
xor XOR2 (N3089, N3088, N2977);
nand NAND4 (N3090, N3082, N341, N2079, N1995);
and AND4 (N3091, N3089, N2735, N2086, N1198);
nor NOR2 (N3092, N3080, N327);
or OR4 (N3093, N3092, N2477, N1649, N563);
and AND4 (N3094, N3093, N902, N2497, N760);
not NOT1 (N3095, N3079);
buf BUF1 (N3096, N3087);
xor XOR2 (N3097, N3091, N1773);
not NOT1 (N3098, N3083);
nand NAND4 (N3099, N3095, N2547, N1926, N1469);
buf BUF1 (N3100, N3086);
buf BUF1 (N3101, N3094);
buf BUF1 (N3102, N3012);
nor NOR3 (N3103, N3099, N4, N51);
nand NAND3 (N3104, N3097, N1072, N425);
nand NAND3 (N3105, N3101, N2886, N3069);
nand NAND3 (N3106, N3102, N2667, N1029);
nor NOR3 (N3107, N3100, N3095, N2801);
not NOT1 (N3108, N3103);
nor NOR3 (N3109, N3061, N3029, N2588);
not NOT1 (N3110, N3090);
buf BUF1 (N3111, N3096);
or OR3 (N3112, N3110, N1469, N266);
not NOT1 (N3113, N3109);
or OR4 (N3114, N3112, N906, N2267, N1275);
and AND4 (N3115, N3098, N2015, N403, N2037);
nor NOR4 (N3116, N3105, N1543, N433, N2661);
or OR3 (N3117, N3106, N614, N61);
nand NAND3 (N3118, N3117, N950, N2281);
nand NAND4 (N3119, N3118, N2018, N2352, N2183);
not NOT1 (N3120, N3104);
buf BUF1 (N3121, N3107);
nor NOR3 (N3122, N3116, N2544, N2114);
nor NOR2 (N3123, N3120, N788);
nor NOR3 (N3124, N3085, N2334, N609);
xor XOR2 (N3125, N3108, N2684);
nor NOR3 (N3126, N3115, N498, N1364);
nor NOR2 (N3127, N3113, N2783);
buf BUF1 (N3128, N3127);
and AND3 (N3129, N3121, N2401, N1771);
not NOT1 (N3130, N3111);
nor NOR3 (N3131, N3124, N1318, N1321);
nand NAND4 (N3132, N3119, N2441, N1216, N2133);
not NOT1 (N3133, N3129);
not NOT1 (N3134, N3133);
and AND2 (N3135, N3122, N85);
nand NAND3 (N3136, N3135, N1647, N2123);
buf BUF1 (N3137, N3136);
and AND4 (N3138, N3134, N1636, N1239, N1946);
nand NAND4 (N3139, N3130, N1176, N1637, N1568);
xor XOR2 (N3140, N3137, N1947);
or OR2 (N3141, N3131, N1112);
nor NOR3 (N3142, N3128, N469, N1565);
nor NOR4 (N3143, N3139, N1288, N510, N947);
nand NAND3 (N3144, N3141, N2365, N187);
nor NOR4 (N3145, N3132, N2808, N2097, N823);
buf BUF1 (N3146, N3145);
and AND4 (N3147, N3142, N824, N365, N2219);
nor NOR2 (N3148, N3126, N2869);
and AND2 (N3149, N3114, N2021);
buf BUF1 (N3150, N3147);
nand NAND2 (N3151, N3138, N2435);
not NOT1 (N3152, N3149);
xor XOR2 (N3153, N3151, N1753);
xor XOR2 (N3154, N3152, N261);
nand NAND4 (N3155, N3154, N2757, N1347, N679);
not NOT1 (N3156, N3143);
or OR3 (N3157, N3123, N2472, N2880);
xor XOR2 (N3158, N3148, N1830);
or OR4 (N3159, N3153, N2989, N3075, N1369);
xor XOR2 (N3160, N3140, N749);
nand NAND2 (N3161, N3146, N3129);
nor NOR4 (N3162, N3157, N1509, N757, N642);
or OR3 (N3163, N3161, N443, N632);
or OR2 (N3164, N3155, N2819);
buf BUF1 (N3165, N3150);
or OR2 (N3166, N3163, N527);
not NOT1 (N3167, N3159);
not NOT1 (N3168, N3166);
and AND2 (N3169, N3160, N1344);
and AND3 (N3170, N3125, N2620, N2679);
and AND3 (N3171, N3169, N1164, N2924);
xor XOR2 (N3172, N3167, N2193);
nor NOR2 (N3173, N3172, N1113);
nand NAND3 (N3174, N3158, N688, N2849);
not NOT1 (N3175, N3174);
not NOT1 (N3176, N3171);
or OR4 (N3177, N3173, N771, N1344, N147);
and AND3 (N3178, N3176, N1415, N3009);
or OR2 (N3179, N3177, N194);
xor XOR2 (N3180, N3178, N784);
nor NOR3 (N3181, N3175, N1588, N281);
and AND3 (N3182, N3181, N2124, N1129);
xor XOR2 (N3183, N3162, N1708);
not NOT1 (N3184, N3179);
nand NAND2 (N3185, N3182, N2686);
xor XOR2 (N3186, N3165, N2513);
nand NAND2 (N3187, N3183, N310);
xor XOR2 (N3188, N3156, N207);
buf BUF1 (N3189, N3184);
xor XOR2 (N3190, N3189, N266);
xor XOR2 (N3191, N3190, N2878);
xor XOR2 (N3192, N3191, N1325);
and AND3 (N3193, N3185, N208, N2514);
xor XOR2 (N3194, N3170, N2629);
nor NOR2 (N3195, N3194, N966);
xor XOR2 (N3196, N3187, N1088);
nor NOR3 (N3197, N3180, N2345, N1939);
nand NAND3 (N3198, N3188, N2470, N2767);
not NOT1 (N3199, N3195);
not NOT1 (N3200, N3144);
buf BUF1 (N3201, N3168);
not NOT1 (N3202, N3201);
nor NOR3 (N3203, N3199, N459, N371);
xor XOR2 (N3204, N3196, N1920);
nor NOR4 (N3205, N3198, N1843, N2554, N2893);
nand NAND4 (N3206, N3202, N2690, N2284, N2302);
or OR2 (N3207, N3206, N891);
or OR3 (N3208, N3186, N1422, N1839);
not NOT1 (N3209, N3164);
or OR2 (N3210, N3204, N2953);
buf BUF1 (N3211, N3200);
or OR2 (N3212, N3192, N2048);
not NOT1 (N3213, N3203);
xor XOR2 (N3214, N3197, N3078);
and AND4 (N3215, N3205, N3200, N652, N2897);
not NOT1 (N3216, N3215);
buf BUF1 (N3217, N3213);
and AND4 (N3218, N3217, N1353, N1664, N949);
or OR4 (N3219, N3209, N1000, N2901, N134);
nand NAND2 (N3220, N3214, N2085);
or OR4 (N3221, N3207, N2559, N2532, N261);
nand NAND3 (N3222, N3210, N1879, N2791);
or OR2 (N3223, N3216, N1198);
buf BUF1 (N3224, N3212);
buf BUF1 (N3225, N3220);
nand NAND4 (N3226, N3222, N2605, N2579, N1581);
not NOT1 (N3227, N3193);
nor NOR2 (N3228, N3221, N2587);
or OR2 (N3229, N3227, N1526);
and AND2 (N3230, N3218, N1530);
and AND3 (N3231, N3226, N1285, N3025);
and AND4 (N3232, N3229, N1034, N786, N915);
nand NAND2 (N3233, N3228, N51);
buf BUF1 (N3234, N3232);
and AND2 (N3235, N3219, N1824);
or OR3 (N3236, N3211, N2439, N2194);
buf BUF1 (N3237, N3236);
nand NAND2 (N3238, N3224, N3035);
not NOT1 (N3239, N3231);
not NOT1 (N3240, N3235);
or OR2 (N3241, N3237, N1677);
or OR3 (N3242, N3223, N690, N928);
or OR3 (N3243, N3241, N1037, N293);
buf BUF1 (N3244, N3240);
or OR4 (N3245, N3234, N1945, N371, N1560);
xor XOR2 (N3246, N3233, N55);
buf BUF1 (N3247, N3242);
buf BUF1 (N3248, N3246);
buf BUF1 (N3249, N3238);
xor XOR2 (N3250, N3208, N1036);
not NOT1 (N3251, N3245);
and AND4 (N3252, N3248, N975, N1001, N1621);
buf BUF1 (N3253, N3244);
and AND2 (N3254, N3239, N2638);
xor XOR2 (N3255, N3251, N1465);
or OR4 (N3256, N3252, N182, N1498, N1558);
nand NAND2 (N3257, N3243, N306);
nand NAND2 (N3258, N3247, N2038);
buf BUF1 (N3259, N3256);
or OR3 (N3260, N3250, N1671, N14);
buf BUF1 (N3261, N3257);
xor XOR2 (N3262, N3254, N2535);
nand NAND2 (N3263, N3253, N3089);
nor NOR4 (N3264, N3258, N2177, N439, N1690);
nand NAND2 (N3265, N3261, N14);
nor NOR3 (N3266, N3259, N3092, N1598);
xor XOR2 (N3267, N3260, N660);
xor XOR2 (N3268, N3262, N3023);
nor NOR3 (N3269, N3263, N1387, N1602);
nand NAND2 (N3270, N3265, N485);
and AND3 (N3271, N3230, N269, N1594);
xor XOR2 (N3272, N3266, N1787);
nor NOR3 (N3273, N3268, N513, N785);
xor XOR2 (N3274, N3269, N1885);
or OR4 (N3275, N3267, N3143, N2688, N1556);
nor NOR2 (N3276, N3249, N2503);
xor XOR2 (N3277, N3275, N3104);
nor NOR4 (N3278, N3272, N2219, N564, N121);
and AND4 (N3279, N3225, N1007, N1454, N3247);
nor NOR2 (N3280, N3274, N2021);
buf BUF1 (N3281, N3279);
xor XOR2 (N3282, N3264, N1487);
xor XOR2 (N3283, N3278, N1599);
buf BUF1 (N3284, N3277);
nand NAND3 (N3285, N3271, N1964, N2839);
xor XOR2 (N3286, N3255, N1692);
and AND2 (N3287, N3276, N2203);
nand NAND2 (N3288, N3273, N1273);
nand NAND3 (N3289, N3282, N1812, N737);
or OR2 (N3290, N3288, N1796);
nor NOR2 (N3291, N3289, N1669);
or OR4 (N3292, N3290, N2612, N36, N753);
not NOT1 (N3293, N3287);
not NOT1 (N3294, N3286);
not NOT1 (N3295, N3270);
and AND3 (N3296, N3294, N1576, N1904);
nor NOR4 (N3297, N3295, N367, N488, N736);
nor NOR4 (N3298, N3284, N67, N2466, N2646);
not NOT1 (N3299, N3293);
or OR3 (N3300, N3299, N2934, N3255);
and AND4 (N3301, N3280, N1435, N3, N1699);
buf BUF1 (N3302, N3281);
xor XOR2 (N3303, N3291, N1392);
buf BUF1 (N3304, N3297);
xor XOR2 (N3305, N3285, N1695);
nor NOR4 (N3306, N3296, N1919, N917, N1291);
nand NAND4 (N3307, N3304, N851, N2730, N230);
and AND3 (N3308, N3306, N423, N1651);
not NOT1 (N3309, N3298);
buf BUF1 (N3310, N3308);
not NOT1 (N3311, N3300);
and AND4 (N3312, N3292, N1083, N3130, N1172);
nand NAND4 (N3313, N3311, N276, N1029, N1182);
not NOT1 (N3314, N3312);
nor NOR3 (N3315, N3313, N1275, N1364);
or OR2 (N3316, N3301, N815);
not NOT1 (N3317, N3309);
nor NOR4 (N3318, N3307, N3021, N1167, N3147);
nand NAND3 (N3319, N3305, N2368, N2031);
not NOT1 (N3320, N3310);
xor XOR2 (N3321, N3314, N2598);
and AND3 (N3322, N3319, N2234, N1899);
nor NOR3 (N3323, N3283, N940, N3193);
nand NAND3 (N3324, N3302, N324, N2985);
xor XOR2 (N3325, N3317, N64);
buf BUF1 (N3326, N3322);
not NOT1 (N3327, N3315);
nand NAND3 (N3328, N3327, N915, N1);
and AND3 (N3329, N3320, N1788, N1439);
xor XOR2 (N3330, N3318, N80);
nor NOR4 (N3331, N3328, N368, N10, N2913);
nand NAND3 (N3332, N3324, N3134, N756);
nand NAND3 (N3333, N3330, N2155, N619);
buf BUF1 (N3334, N3303);
or OR4 (N3335, N3325, N1921, N3027, N196);
not NOT1 (N3336, N3332);
buf BUF1 (N3337, N3335);
not NOT1 (N3338, N3329);
not NOT1 (N3339, N3323);
nand NAND2 (N3340, N3316, N2777);
nand NAND3 (N3341, N3331, N1198, N3339);
or OR2 (N3342, N985, N2537);
not NOT1 (N3343, N3337);
or OR2 (N3344, N3342, N2578);
and AND2 (N3345, N3334, N1581);
nand NAND2 (N3346, N3338, N148);
nand NAND3 (N3347, N3340, N865, N1119);
or OR4 (N3348, N3336, N666, N3137, N46);
nand NAND2 (N3349, N3347, N1029);
buf BUF1 (N3350, N3321);
xor XOR2 (N3351, N3344, N3255);
not NOT1 (N3352, N3346);
or OR2 (N3353, N3345, N2734);
and AND2 (N3354, N3341, N1241);
nor NOR3 (N3355, N3353, N1723, N2895);
buf BUF1 (N3356, N3348);
xor XOR2 (N3357, N3356, N1549);
not NOT1 (N3358, N3351);
nor NOR4 (N3359, N3352, N123, N838, N1403);
nor NOR3 (N3360, N3350, N137, N1591);
not NOT1 (N3361, N3357);
not NOT1 (N3362, N3333);
or OR3 (N3363, N3358, N2699, N2583);
nor NOR2 (N3364, N3360, N1548);
nand NAND3 (N3365, N3362, N1753, N2367);
nand NAND2 (N3366, N3365, N334);
not NOT1 (N3367, N3364);
or OR2 (N3368, N3354, N2294);
nor NOR4 (N3369, N3368, N3013, N922, N2911);
or OR3 (N3370, N3363, N1043, N1632);
not NOT1 (N3371, N3361);
and AND4 (N3372, N3349, N1270, N2001, N3194);
nand NAND2 (N3373, N3371, N482);
and AND3 (N3374, N3326, N1970, N1617);
or OR4 (N3375, N3374, N976, N3339, N2047);
buf BUF1 (N3376, N3366);
not NOT1 (N3377, N3355);
and AND2 (N3378, N3376, N1241);
xor XOR2 (N3379, N3373, N3220);
or OR2 (N3380, N3379, N1057);
buf BUF1 (N3381, N3377);
nand NAND2 (N3382, N3380, N793);
not NOT1 (N3383, N3375);
nor NOR3 (N3384, N3381, N2472, N61);
and AND4 (N3385, N3369, N1962, N1140, N43);
buf BUF1 (N3386, N3384);
not NOT1 (N3387, N3382);
buf BUF1 (N3388, N3359);
or OR2 (N3389, N3370, N2973);
or OR2 (N3390, N3378, N1082);
xor XOR2 (N3391, N3343, N1411);
not NOT1 (N3392, N3386);
buf BUF1 (N3393, N3388);
nand NAND4 (N3394, N3387, N42, N724, N673);
nor NOR2 (N3395, N3367, N1257);
nand NAND3 (N3396, N3385, N2158, N1659);
nor NOR2 (N3397, N3394, N1242);
nor NOR2 (N3398, N3393, N1333);
nand NAND3 (N3399, N3398, N3180, N518);
xor XOR2 (N3400, N3391, N1491);
nand NAND2 (N3401, N3389, N695);
and AND2 (N3402, N3395, N1858);
nor NOR4 (N3403, N3392, N1700, N211, N2939);
nand NAND2 (N3404, N3400, N662);
buf BUF1 (N3405, N3401);
and AND3 (N3406, N3405, N1819, N2963);
xor XOR2 (N3407, N3397, N1074);
and AND4 (N3408, N3399, N2821, N551, N2989);
or OR4 (N3409, N3403, N2492, N542, N1413);
and AND4 (N3410, N3372, N2086, N1874, N1887);
and AND4 (N3411, N3396, N1616, N425, N1074);
nor NOR3 (N3412, N3402, N1041, N2290);
nand NAND3 (N3413, N3412, N1196, N2160);
nor NOR3 (N3414, N3407, N2812, N53);
xor XOR2 (N3415, N3413, N2259);
nor NOR3 (N3416, N3408, N235, N1206);
or OR2 (N3417, N3409, N2281);
not NOT1 (N3418, N3415);
nor NOR2 (N3419, N3390, N2389);
xor XOR2 (N3420, N3404, N1221);
not NOT1 (N3421, N3417);
or OR3 (N3422, N3383, N9, N2103);
buf BUF1 (N3423, N3416);
or OR3 (N3424, N3421, N2398, N2752);
buf BUF1 (N3425, N3420);
buf BUF1 (N3426, N3406);
nor NOR3 (N3427, N3418, N2282, N389);
xor XOR2 (N3428, N3414, N2603);
xor XOR2 (N3429, N3422, N1311);
or OR3 (N3430, N3410, N626, N2533);
and AND3 (N3431, N3428, N1617, N442);
and AND3 (N3432, N3429, N1754, N1873);
buf BUF1 (N3433, N3427);
nor NOR4 (N3434, N3432, N1279, N1006, N1547);
and AND2 (N3435, N3434, N1468);
nand NAND2 (N3436, N3425, N3334);
nor NOR2 (N3437, N3430, N880);
buf BUF1 (N3438, N3436);
buf BUF1 (N3439, N3419);
and AND2 (N3440, N3438, N951);
nand NAND4 (N3441, N3423, N979, N1030, N3393);
nor NOR3 (N3442, N3439, N1834, N1093);
not NOT1 (N3443, N3411);
nor NOR3 (N3444, N3443, N966, N2768);
not NOT1 (N3445, N3424);
buf BUF1 (N3446, N3444);
xor XOR2 (N3447, N3442, N1388);
nor NOR2 (N3448, N3440, N1718);
xor XOR2 (N3449, N3437, N2190);
nand NAND4 (N3450, N3435, N1491, N41, N1133);
and AND4 (N3451, N3431, N1631, N2917, N1615);
not NOT1 (N3452, N3445);
nor NOR2 (N3453, N3446, N1423);
or OR2 (N3454, N3426, N45);
xor XOR2 (N3455, N3454, N1957);
xor XOR2 (N3456, N3451, N2970);
or OR2 (N3457, N3453, N3311);
xor XOR2 (N3458, N3433, N3149);
and AND3 (N3459, N3458, N2733, N1927);
and AND4 (N3460, N3447, N1001, N3033, N1066);
or OR4 (N3461, N3452, N960, N2794, N2135);
nand NAND4 (N3462, N3455, N1775, N2769, N3276);
buf BUF1 (N3463, N3457);
not NOT1 (N3464, N3461);
nor NOR3 (N3465, N3441, N2305, N1623);
nand NAND4 (N3466, N3456, N229, N2656, N2071);
nor NOR3 (N3467, N3449, N3445, N288);
and AND3 (N3468, N3464, N1019, N1815);
and AND2 (N3469, N3467, N635);
or OR3 (N3470, N3450, N3046, N1290);
buf BUF1 (N3471, N3469);
buf BUF1 (N3472, N3460);
and AND4 (N3473, N3462, N2415, N3002, N218);
buf BUF1 (N3474, N3463);
nand NAND3 (N3475, N3474, N1873, N524);
nor NOR2 (N3476, N3468, N1818);
buf BUF1 (N3477, N3448);
nand NAND2 (N3478, N3470, N1185);
buf BUF1 (N3479, N3459);
buf BUF1 (N3480, N3479);
or OR4 (N3481, N3475, N2033, N1436, N314);
nor NOR3 (N3482, N3466, N1827, N118);
xor XOR2 (N3483, N3480, N312);
or OR2 (N3484, N3478, N247);
xor XOR2 (N3485, N3484, N2190);
or OR2 (N3486, N3485, N1743);
or OR4 (N3487, N3476, N881, N1340, N3006);
and AND2 (N3488, N3473, N2185);
and AND3 (N3489, N3465, N1836, N1899);
nand NAND4 (N3490, N3486, N1858, N2125, N3310);
xor XOR2 (N3491, N3477, N3098);
xor XOR2 (N3492, N3489, N2197);
nor NOR4 (N3493, N3490, N3279, N2515, N3058);
xor XOR2 (N3494, N3482, N416);
not NOT1 (N3495, N3471);
or OR4 (N3496, N3481, N1500, N2294, N1236);
or OR4 (N3497, N3472, N789, N443, N2389);
not NOT1 (N3498, N3487);
nor NOR3 (N3499, N3483, N1482, N3496);
xor XOR2 (N3500, N2817, N3286);
not NOT1 (N3501, N3499);
nor NOR2 (N3502, N3500, N64);
and AND4 (N3503, N3501, N506, N3318, N541);
nor NOR3 (N3504, N3494, N443, N1997);
not NOT1 (N3505, N3498);
xor XOR2 (N3506, N3497, N1515);
and AND4 (N3507, N3495, N140, N1964, N1727);
buf BUF1 (N3508, N3493);
not NOT1 (N3509, N3488);
buf BUF1 (N3510, N3507);
or OR4 (N3511, N3506, N575, N619, N281);
nor NOR2 (N3512, N3491, N348);
or OR4 (N3513, N3505, N122, N391, N3271);
or OR2 (N3514, N3513, N2550);
or OR4 (N3515, N3511, N1626, N2470, N3398);
not NOT1 (N3516, N3509);
nor NOR4 (N3517, N3502, N2054, N1308, N3007);
nand NAND4 (N3518, N3492, N3027, N66, N2584);
nor NOR3 (N3519, N3512, N1231, N1305);
and AND4 (N3520, N3515, N570, N1494, N2355);
buf BUF1 (N3521, N3519);
buf BUF1 (N3522, N3517);
or OR3 (N3523, N3522, N2919, N3009);
xor XOR2 (N3524, N3520, N275);
buf BUF1 (N3525, N3516);
or OR4 (N3526, N3504, N622, N2244, N586);
and AND4 (N3527, N3523, N1129, N1435, N1301);
or OR2 (N3528, N3524, N703);
nand NAND3 (N3529, N3525, N2677, N2513);
nor NOR2 (N3530, N3529, N2752);
xor XOR2 (N3531, N3527, N735);
or OR3 (N3532, N3518, N651, N2967);
nand NAND2 (N3533, N3528, N1811);
and AND3 (N3534, N3532, N318, N2003);
not NOT1 (N3535, N3534);
not NOT1 (N3536, N3526);
nor NOR2 (N3537, N3531, N821);
buf BUF1 (N3538, N3530);
nor NOR4 (N3539, N3536, N3475, N3522, N3310);
buf BUF1 (N3540, N3521);
not NOT1 (N3541, N3538);
buf BUF1 (N3542, N3535);
buf BUF1 (N3543, N3514);
nor NOR3 (N3544, N3539, N1660, N123);
xor XOR2 (N3545, N3503, N920);
or OR2 (N3546, N3542, N2531);
not NOT1 (N3547, N3546);
nor NOR3 (N3548, N3547, N101, N2782);
nor NOR2 (N3549, N3544, N1285);
buf BUF1 (N3550, N3541);
and AND3 (N3551, N3508, N2013, N1503);
or OR3 (N3552, N3533, N3029, N36);
buf BUF1 (N3553, N3551);
buf BUF1 (N3554, N3510);
and AND3 (N3555, N3543, N40, N947);
nor NOR2 (N3556, N3550, N469);
not NOT1 (N3557, N3537);
buf BUF1 (N3558, N3553);
or OR2 (N3559, N3549, N315);
not NOT1 (N3560, N3555);
not NOT1 (N3561, N3558);
xor XOR2 (N3562, N3548, N3006);
nor NOR2 (N3563, N3561, N1312);
or OR4 (N3564, N3559, N664, N455, N723);
and AND4 (N3565, N3556, N3443, N2222, N768);
or OR4 (N3566, N3560, N529, N316, N435);
nor NOR4 (N3567, N3545, N887, N1238, N3173);
buf BUF1 (N3568, N3566);
and AND2 (N3569, N3564, N3016);
nor NOR4 (N3570, N3557, N1161, N1894, N2412);
or OR3 (N3571, N3568, N2504, N2831);
not NOT1 (N3572, N3554);
nor NOR3 (N3573, N3567, N1209, N1341);
nand NAND2 (N3574, N3572, N3004);
not NOT1 (N3575, N3563);
xor XOR2 (N3576, N3552, N724);
nand NAND3 (N3577, N3571, N71, N1297);
or OR3 (N3578, N3577, N1003, N1995);
nor NOR4 (N3579, N3574, N150, N356, N1441);
not NOT1 (N3580, N3562);
and AND2 (N3581, N3575, N1593);
and AND3 (N3582, N3578, N2006, N2216);
not NOT1 (N3583, N3565);
buf BUF1 (N3584, N3583);
and AND4 (N3585, N3573, N1722, N1567, N415);
buf BUF1 (N3586, N3579);
not NOT1 (N3587, N3581);
and AND3 (N3588, N3586, N902, N1093);
or OR4 (N3589, N3576, N802, N1652, N332);
nor NOR2 (N3590, N3584, N2168);
xor XOR2 (N3591, N3569, N1740);
not NOT1 (N3592, N3589);
not NOT1 (N3593, N3588);
or OR4 (N3594, N3582, N61, N1048, N113);
not NOT1 (N3595, N3580);
buf BUF1 (N3596, N3585);
or OR3 (N3597, N3570, N810, N442);
xor XOR2 (N3598, N3594, N633);
nor NOR4 (N3599, N3596, N743, N327, N1565);
not NOT1 (N3600, N3593);
not NOT1 (N3601, N3600);
buf BUF1 (N3602, N3595);
xor XOR2 (N3603, N3601, N1651);
or OR2 (N3604, N3590, N263);
buf BUF1 (N3605, N3599);
not NOT1 (N3606, N3587);
or OR2 (N3607, N3591, N3475);
and AND4 (N3608, N3540, N791, N2829, N102);
buf BUF1 (N3609, N3604);
nor NOR4 (N3610, N3609, N2519, N3316, N2453);
or OR4 (N3611, N3605, N3406, N2543, N1155);
nand NAND2 (N3612, N3597, N470);
not NOT1 (N3613, N3611);
xor XOR2 (N3614, N3606, N2881);
nor NOR4 (N3615, N3612, N232, N2088, N3220);
nand NAND3 (N3616, N3603, N1619, N1461);
or OR2 (N3617, N3608, N2107);
not NOT1 (N3618, N3617);
buf BUF1 (N3619, N3592);
and AND2 (N3620, N3607, N1948);
or OR4 (N3621, N3613, N3426, N2318, N1492);
and AND4 (N3622, N3615, N3484, N3284, N227);
buf BUF1 (N3623, N3622);
and AND3 (N3624, N3623, N3376, N1193);
buf BUF1 (N3625, N3618);
nand NAND2 (N3626, N3616, N1984);
nand NAND2 (N3627, N3625, N1809);
and AND2 (N3628, N3598, N2963);
nand NAND4 (N3629, N3624, N968, N822, N584);
xor XOR2 (N3630, N3614, N1346);
and AND3 (N3631, N3626, N373, N2850);
xor XOR2 (N3632, N3619, N1994);
nor NOR4 (N3633, N3630, N3217, N26, N2299);
buf BUF1 (N3634, N3602);
not NOT1 (N3635, N3620);
and AND3 (N3636, N3627, N1225, N871);
nand NAND4 (N3637, N3636, N2313, N180, N3209);
and AND4 (N3638, N3629, N925, N3033, N602);
and AND4 (N3639, N3634, N821, N971, N1632);
nor NOR3 (N3640, N3628, N1935, N3415);
nor NOR4 (N3641, N3610, N788, N3128, N2680);
buf BUF1 (N3642, N3640);
nor NOR2 (N3643, N3621, N3122);
nand NAND3 (N3644, N3642, N2347, N323);
or OR4 (N3645, N3631, N3148, N1411, N289);
xor XOR2 (N3646, N3633, N2855);
or OR2 (N3647, N3637, N3449);
or OR2 (N3648, N3639, N3338);
and AND3 (N3649, N3638, N839, N1096);
and AND4 (N3650, N3646, N3160, N2869, N2100);
nor NOR3 (N3651, N3635, N758, N1298);
xor XOR2 (N3652, N3644, N2465);
buf BUF1 (N3653, N3652);
nor NOR2 (N3654, N3632, N2887);
not NOT1 (N3655, N3645);
and AND2 (N3656, N3649, N2697);
or OR4 (N3657, N3656, N3107, N139, N2329);
or OR2 (N3658, N3641, N2915);
nand NAND2 (N3659, N3643, N2447);
buf BUF1 (N3660, N3654);
buf BUF1 (N3661, N3657);
nand NAND3 (N3662, N3648, N2437, N1506);
xor XOR2 (N3663, N3660, N3133);
and AND3 (N3664, N3655, N3020, N2494);
xor XOR2 (N3665, N3650, N1418);
xor XOR2 (N3666, N3659, N816);
not NOT1 (N3667, N3663);
buf BUF1 (N3668, N3647);
or OR3 (N3669, N3665, N3425, N2827);
and AND2 (N3670, N3669, N2956);
xor XOR2 (N3671, N3670, N3150);
or OR2 (N3672, N3667, N862);
nor NOR2 (N3673, N3653, N2008);
and AND3 (N3674, N3664, N3537, N2622);
nand NAND3 (N3675, N3668, N825, N198);
not NOT1 (N3676, N3672);
xor XOR2 (N3677, N3661, N624);
and AND3 (N3678, N3671, N1149, N622);
not NOT1 (N3679, N3658);
and AND3 (N3680, N3666, N1537, N220);
or OR3 (N3681, N3675, N3159, N195);
not NOT1 (N3682, N3680);
nor NOR2 (N3683, N3678, N15);
nand NAND2 (N3684, N3682, N1789);
not NOT1 (N3685, N3681);
not NOT1 (N3686, N3683);
or OR2 (N3687, N3684, N902);
nor NOR4 (N3688, N3685, N1105, N1046, N1769);
nand NAND3 (N3689, N3662, N2396, N2610);
nand NAND3 (N3690, N3679, N952, N530);
not NOT1 (N3691, N3674);
nand NAND4 (N3692, N3676, N846, N2105, N1564);
and AND4 (N3693, N3687, N2529, N2186, N147);
not NOT1 (N3694, N3692);
xor XOR2 (N3695, N3673, N2628);
xor XOR2 (N3696, N3694, N2803);
and AND2 (N3697, N3696, N3640);
buf BUF1 (N3698, N3695);
buf BUF1 (N3699, N3686);
xor XOR2 (N3700, N3697, N1761);
nand NAND4 (N3701, N3651, N3413, N774, N2541);
not NOT1 (N3702, N3698);
and AND2 (N3703, N3690, N1861);
buf BUF1 (N3704, N3699);
nor NOR2 (N3705, N3703, N1507);
xor XOR2 (N3706, N3705, N3420);
nor NOR3 (N3707, N3704, N1510, N2001);
xor XOR2 (N3708, N3700, N1);
and AND3 (N3709, N3706, N65, N435);
not NOT1 (N3710, N3702);
nand NAND4 (N3711, N3707, N1949, N3352, N2951);
xor XOR2 (N3712, N3701, N2805);
nor NOR4 (N3713, N3677, N2076, N2544, N3022);
not NOT1 (N3714, N3711);
and AND2 (N3715, N3712, N1007);
nor NOR3 (N3716, N3713, N958, N1218);
nor NOR4 (N3717, N3714, N3199, N3153, N2228);
or OR4 (N3718, N3689, N1312, N963, N352);
buf BUF1 (N3719, N3693);
not NOT1 (N3720, N3715);
xor XOR2 (N3721, N3710, N1075);
nor NOR3 (N3722, N3719, N1417, N2544);
not NOT1 (N3723, N3709);
or OR2 (N3724, N3691, N3297);
xor XOR2 (N3725, N3716, N2061);
nor NOR4 (N3726, N3688, N1545, N1795, N613);
not NOT1 (N3727, N3726);
or OR4 (N3728, N3720, N1808, N1697, N271);
buf BUF1 (N3729, N3721);
buf BUF1 (N3730, N3722);
and AND2 (N3731, N3729, N2107);
not NOT1 (N3732, N3723);
not NOT1 (N3733, N3724);
xor XOR2 (N3734, N3732, N2788);
nand NAND4 (N3735, N3718, N2610, N2339, N2006);
not NOT1 (N3736, N3717);
buf BUF1 (N3737, N3731);
and AND4 (N3738, N3725, N2164, N2865, N137);
buf BUF1 (N3739, N3736);
and AND2 (N3740, N3708, N1699);
buf BUF1 (N3741, N3727);
xor XOR2 (N3742, N3733, N2368);
nor NOR2 (N3743, N3742, N2328);
nor NOR3 (N3744, N3730, N3560, N3431);
nor NOR4 (N3745, N3737, N2890, N1675, N1347);
xor XOR2 (N3746, N3728, N1235);
nand NAND3 (N3747, N3735, N491, N753);
xor XOR2 (N3748, N3744, N141);
or OR3 (N3749, N3740, N1321, N749);
nand NAND4 (N3750, N3747, N1578, N2044, N1173);
xor XOR2 (N3751, N3748, N1965);
buf BUF1 (N3752, N3743);
not NOT1 (N3753, N3745);
and AND4 (N3754, N3751, N1237, N282, N1560);
or OR4 (N3755, N3749, N1285, N3171, N987);
buf BUF1 (N3756, N3750);
or OR4 (N3757, N3738, N419, N3520, N3388);
not NOT1 (N3758, N3757);
or OR4 (N3759, N3739, N1413, N2434, N2861);
or OR3 (N3760, N3754, N650, N1576);
or OR2 (N3761, N3755, N2191);
not NOT1 (N3762, N3760);
nor NOR3 (N3763, N3761, N2031, N3426);
xor XOR2 (N3764, N3759, N1129);
and AND4 (N3765, N3753, N222, N3591, N1255);
and AND3 (N3766, N3752, N754, N663);
or OR4 (N3767, N3756, N410, N781, N1203);
and AND4 (N3768, N3765, N2400, N2996, N749);
nor NOR4 (N3769, N3767, N2662, N3226, N3206);
buf BUF1 (N3770, N3764);
nor NOR3 (N3771, N3746, N3453, N1231);
or OR4 (N3772, N3763, N1567, N502, N1379);
or OR2 (N3773, N3766, N2787);
and AND4 (N3774, N3734, N590, N2120, N2914);
nor NOR3 (N3775, N3762, N707, N3075);
not NOT1 (N3776, N3770);
and AND4 (N3777, N3769, N2864, N1945, N3034);
xor XOR2 (N3778, N3741, N3731);
and AND3 (N3779, N3777, N1077, N1094);
xor XOR2 (N3780, N3773, N3108);
or OR3 (N3781, N3772, N993, N651);
buf BUF1 (N3782, N3774);
nor NOR3 (N3783, N3782, N2642, N2254);
not NOT1 (N3784, N3780);
xor XOR2 (N3785, N3779, N3779);
and AND4 (N3786, N3785, N3519, N2004, N3554);
or OR3 (N3787, N3758, N2509, N1597);
or OR4 (N3788, N3778, N2144, N1883, N2458);
nor NOR4 (N3789, N3783, N2603, N1092, N415);
or OR3 (N3790, N3784, N2395, N397);
nand NAND4 (N3791, N3789, N2755, N1975, N2715);
or OR2 (N3792, N3775, N1495);
and AND3 (N3793, N3776, N1198, N1496);
nand NAND2 (N3794, N3771, N1400);
nor NOR3 (N3795, N3786, N1108, N2725);
not NOT1 (N3796, N3791);
nand NAND2 (N3797, N3792, N2408);
xor XOR2 (N3798, N3797, N1261);
or OR2 (N3799, N3787, N1965);
nor NOR3 (N3800, N3794, N1818, N1317);
and AND2 (N3801, N3799, N2202);
nand NAND2 (N3802, N3796, N1944);
not NOT1 (N3803, N3802);
nor NOR3 (N3804, N3801, N1006, N931);
nand NAND3 (N3805, N3798, N440, N1449);
buf BUF1 (N3806, N3805);
buf BUF1 (N3807, N3804);
or OR3 (N3808, N3790, N320, N594);
nand NAND3 (N3809, N3793, N2598, N3384);
buf BUF1 (N3810, N3781);
buf BUF1 (N3811, N3808);
not NOT1 (N3812, N3803);
and AND2 (N3813, N3800, N3630);
and AND2 (N3814, N3810, N300);
and AND3 (N3815, N3768, N1594, N3361);
and AND4 (N3816, N3814, N1710, N2555, N167);
or OR4 (N3817, N3788, N1063, N1145, N1095);
nand NAND4 (N3818, N3812, N1889, N1611, N3343);
buf BUF1 (N3819, N3806);
not NOT1 (N3820, N3811);
and AND3 (N3821, N3815, N981, N2644);
xor XOR2 (N3822, N3820, N744);
and AND2 (N3823, N3818, N1739);
xor XOR2 (N3824, N3795, N3036);
or OR3 (N3825, N3821, N789, N2681);
nand NAND2 (N3826, N3817, N486);
not NOT1 (N3827, N3819);
and AND2 (N3828, N3813, N2955);
nand NAND4 (N3829, N3824, N189, N486, N3629);
xor XOR2 (N3830, N3807, N1940);
and AND4 (N3831, N3809, N2192, N2774, N2444);
nor NOR4 (N3832, N3823, N1961, N142, N3352);
xor XOR2 (N3833, N3816, N2007);
or OR2 (N3834, N3828, N1468);
or OR2 (N3835, N3832, N2991);
buf BUF1 (N3836, N3831);
nor NOR4 (N3837, N3826, N2160, N485, N1545);
and AND4 (N3838, N3829, N245, N1654, N2737);
buf BUF1 (N3839, N3827);
buf BUF1 (N3840, N3838);
or OR2 (N3841, N3834, N607);
buf BUF1 (N3842, N3836);
or OR3 (N3843, N3822, N3174, N803);
and AND2 (N3844, N3843, N2533);
or OR3 (N3845, N3835, N1755, N2608);
xor XOR2 (N3846, N3825, N2669);
xor XOR2 (N3847, N3830, N2157);
and AND2 (N3848, N3837, N2368);
xor XOR2 (N3849, N3844, N2015);
and AND3 (N3850, N3847, N2424, N1415);
and AND2 (N3851, N3833, N2132);
nor NOR2 (N3852, N3842, N3190);
or OR3 (N3853, N3850, N659, N2929);
not NOT1 (N3854, N3846);
nor NOR4 (N3855, N3845, N1737, N243, N634);
xor XOR2 (N3856, N3852, N2357);
and AND3 (N3857, N3856, N2408, N2202);
buf BUF1 (N3858, N3849);
and AND4 (N3859, N3839, N178, N419, N1121);
buf BUF1 (N3860, N3853);
xor XOR2 (N3861, N3848, N269);
not NOT1 (N3862, N3859);
nand NAND3 (N3863, N3854, N3798, N347);
buf BUF1 (N3864, N3863);
or OR2 (N3865, N3864, N1515);
or OR2 (N3866, N3840, N509);
not NOT1 (N3867, N3861);
or OR2 (N3868, N3862, N1798);
or OR3 (N3869, N3851, N1042, N982);
or OR2 (N3870, N3868, N809);
buf BUF1 (N3871, N3865);
xor XOR2 (N3872, N3866, N1134);
and AND2 (N3873, N3869, N2303);
nand NAND4 (N3874, N3855, N1050, N139, N1275);
not NOT1 (N3875, N3858);
not NOT1 (N3876, N3867);
nor NOR2 (N3877, N3841, N2584);
nand NAND2 (N3878, N3877, N1865);
not NOT1 (N3879, N3876);
xor XOR2 (N3880, N3870, N3877);
xor XOR2 (N3881, N3874, N3130);
not NOT1 (N3882, N3875);
or OR4 (N3883, N3881, N762, N3607, N2795);
nand NAND2 (N3884, N3882, N1631);
buf BUF1 (N3885, N3883);
nor NOR2 (N3886, N3860, N1515);
and AND2 (N3887, N3879, N3854);
or OR4 (N3888, N3857, N3038, N1037, N2945);
or OR3 (N3889, N3880, N1106, N1449);
and AND2 (N3890, N3888, N1821);
or OR4 (N3891, N3889, N2620, N101, N592);
nor NOR2 (N3892, N3890, N1679);
nor NOR3 (N3893, N3871, N3020, N681);
or OR4 (N3894, N3873, N1175, N2599, N897);
xor XOR2 (N3895, N3872, N3254);
xor XOR2 (N3896, N3891, N778);
and AND2 (N3897, N3878, N2085);
nand NAND2 (N3898, N3885, N1428);
nor NOR3 (N3899, N3886, N2181, N3490);
and AND4 (N3900, N3893, N1622, N1428, N136);
not NOT1 (N3901, N3896);
xor XOR2 (N3902, N3900, N1235);
nand NAND4 (N3903, N3901, N3431, N1466, N3538);
buf BUF1 (N3904, N3892);
nand NAND2 (N3905, N3904, N3191);
xor XOR2 (N3906, N3903, N3417);
and AND2 (N3907, N3887, N3240);
nand NAND4 (N3908, N3906, N3451, N2872, N1703);
nor NOR2 (N3909, N3884, N487);
or OR3 (N3910, N3898, N3130, N3587);
nor NOR2 (N3911, N3895, N2807);
xor XOR2 (N3912, N3910, N562);
buf BUF1 (N3913, N3908);
not NOT1 (N3914, N3913);
nand NAND3 (N3915, N3905, N485, N537);
buf BUF1 (N3916, N3902);
buf BUF1 (N3917, N3894);
not NOT1 (N3918, N3911);
or OR2 (N3919, N3899, N3722);
nor NOR4 (N3920, N3909, N1209, N2388, N519);
or OR4 (N3921, N3916, N195, N2638, N3265);
xor XOR2 (N3922, N3907, N2398);
xor XOR2 (N3923, N3912, N3726);
not NOT1 (N3924, N3922);
buf BUF1 (N3925, N3921);
nand NAND2 (N3926, N3917, N1331);
not NOT1 (N3927, N3925);
xor XOR2 (N3928, N3918, N3071);
and AND3 (N3929, N3923, N3449, N416);
nor NOR4 (N3930, N3927, N2161, N1840, N2049);
nor NOR3 (N3931, N3928, N3478, N60);
not NOT1 (N3932, N3926);
and AND3 (N3933, N3931, N1693, N529);
not NOT1 (N3934, N3915);
and AND3 (N3935, N3930, N1111, N1934);
nand NAND2 (N3936, N3933, N1514);
xor XOR2 (N3937, N3914, N97);
nor NOR3 (N3938, N3897, N1549, N772);
nor NOR2 (N3939, N3932, N1112);
xor XOR2 (N3940, N3939, N2026);
and AND3 (N3941, N3935, N394, N3234);
and AND3 (N3942, N3934, N2677, N865);
nand NAND2 (N3943, N3919, N313);
nand NAND4 (N3944, N3940, N3774, N1761, N2721);
not NOT1 (N3945, N3943);
and AND2 (N3946, N3929, N1340);
nand NAND2 (N3947, N3924, N3171);
nand NAND4 (N3948, N3920, N3577, N3471, N315);
xor XOR2 (N3949, N3941, N3852);
nand NAND4 (N3950, N3949, N575, N1897, N1505);
and AND2 (N3951, N3945, N2609);
buf BUF1 (N3952, N3946);
nand NAND4 (N3953, N3951, N1004, N1659, N2891);
or OR2 (N3954, N3948, N1123);
and AND2 (N3955, N3954, N132);
nand NAND4 (N3956, N3942, N902, N1183, N1792);
or OR3 (N3957, N3950, N3422, N908);
xor XOR2 (N3958, N3957, N2626);
xor XOR2 (N3959, N3938, N3634);
not NOT1 (N3960, N3959);
not NOT1 (N3961, N3952);
nand NAND2 (N3962, N3944, N298);
nor NOR2 (N3963, N3937, N2342);
buf BUF1 (N3964, N3958);
nand NAND3 (N3965, N3955, N1856, N1476);
nor NOR3 (N3966, N3953, N3104, N2708);
nor NOR3 (N3967, N3966, N3853, N2610);
buf BUF1 (N3968, N3963);
or OR2 (N3969, N3962, N2711);
or OR2 (N3970, N3968, N1558);
xor XOR2 (N3971, N3969, N2258);
nand NAND4 (N3972, N3961, N1204, N1030, N3553);
nor NOR4 (N3973, N3956, N134, N402, N369);
xor XOR2 (N3974, N3936, N441);
xor XOR2 (N3975, N3964, N1738);
or OR4 (N3976, N3975, N21, N326, N928);
xor XOR2 (N3977, N3973, N1658);
buf BUF1 (N3978, N3972);
not NOT1 (N3979, N3976);
xor XOR2 (N3980, N3971, N1092);
not NOT1 (N3981, N3979);
and AND3 (N3982, N3974, N2493, N2861);
not NOT1 (N3983, N3965);
xor XOR2 (N3984, N3967, N3129);
xor XOR2 (N3985, N3977, N2057);
or OR4 (N3986, N3982, N1511, N2870, N595);
or OR4 (N3987, N3947, N1589, N1706, N2593);
nor NOR2 (N3988, N3986, N2655);
nand NAND2 (N3989, N3984, N1519);
nand NAND2 (N3990, N3978, N752);
nand NAND2 (N3991, N3981, N400);
and AND2 (N3992, N3985, N1704);
nand NAND3 (N3993, N3987, N2303, N674);
or OR3 (N3994, N3988, N2160, N2009);
not NOT1 (N3995, N3989);
nand NAND3 (N3996, N3960, N3234, N945);
buf BUF1 (N3997, N3995);
buf BUF1 (N3998, N3992);
nor NOR4 (N3999, N3996, N2855, N3073, N3353);
or OR3 (N4000, N3970, N2957, N3933);
buf BUF1 (N4001, N3991);
nor NOR2 (N4002, N3994, N2638);
xor XOR2 (N4003, N3990, N3953);
nor NOR3 (N4004, N4000, N532, N2207);
or OR2 (N4005, N4002, N121);
not NOT1 (N4006, N3998);
buf BUF1 (N4007, N4003);
nand NAND2 (N4008, N3993, N2598);
buf BUF1 (N4009, N4005);
nand NAND3 (N4010, N3999, N3048, N2007);
nand NAND2 (N4011, N3983, N2163);
or OR4 (N4012, N4010, N1884, N263, N1257);
or OR3 (N4013, N3980, N1234, N3840);
nand NAND2 (N4014, N4011, N3437);
buf BUF1 (N4015, N4001);
buf BUF1 (N4016, N4012);
and AND2 (N4017, N4004, N2689);
nand NAND2 (N4018, N4013, N1759);
buf BUF1 (N4019, N4014);
xor XOR2 (N4020, N4017, N2105);
buf BUF1 (N4021, N4018);
and AND4 (N4022, N3997, N3568, N980, N679);
or OR2 (N4023, N4016, N3805);
buf BUF1 (N4024, N4008);
or OR3 (N4025, N4007, N4002, N1966);
and AND4 (N4026, N4020, N1103, N1310, N1859);
nand NAND3 (N4027, N4022, N439, N660);
and AND4 (N4028, N4009, N1582, N1062, N217);
nor NOR4 (N4029, N4023, N213, N2737, N1240);
not NOT1 (N4030, N4028);
or OR3 (N4031, N4029, N864, N2146);
nand NAND4 (N4032, N4031, N2944, N3330, N1719);
buf BUF1 (N4033, N4032);
or OR3 (N4034, N4015, N2407, N1051);
nor NOR2 (N4035, N4027, N304);
buf BUF1 (N4036, N4024);
or OR4 (N4037, N4035, N2343, N3071, N1220);
and AND3 (N4038, N4030, N1478, N1611);
xor XOR2 (N4039, N4037, N2034);
not NOT1 (N4040, N4026);
not NOT1 (N4041, N4036);
not NOT1 (N4042, N4040);
xor XOR2 (N4043, N4021, N1039);
buf BUF1 (N4044, N4006);
nand NAND2 (N4045, N4043, N397);
xor XOR2 (N4046, N4034, N3076);
or OR2 (N4047, N4033, N230);
xor XOR2 (N4048, N4042, N4009);
or OR3 (N4049, N4025, N3846, N3484);
nor NOR3 (N4050, N4041, N3511, N2158);
nor NOR3 (N4051, N4044, N4032, N2130);
nor NOR3 (N4052, N4019, N680, N2199);
xor XOR2 (N4053, N4046, N3417);
xor XOR2 (N4054, N4045, N2787);
nor NOR2 (N4055, N4051, N107);
not NOT1 (N4056, N4050);
not NOT1 (N4057, N4038);
or OR4 (N4058, N4056, N713, N3399, N38);
nand NAND3 (N4059, N4054, N696, N1671);
buf BUF1 (N4060, N4058);
nor NOR2 (N4061, N4057, N2367);
nand NAND4 (N4062, N4061, N532, N1810, N1175);
xor XOR2 (N4063, N4052, N4012);
buf BUF1 (N4064, N4060);
nand NAND4 (N4065, N4049, N413, N3097, N1902);
or OR3 (N4066, N4064, N3881, N1948);
nor NOR4 (N4067, N4055, N1631, N805, N2385);
nand NAND2 (N4068, N4053, N3583);
and AND4 (N4069, N4039, N2457, N2077, N3839);
nand NAND4 (N4070, N4068, N523, N3441, N2246);
and AND2 (N4071, N4063, N3180);
nand NAND3 (N4072, N4062, N397, N1748);
not NOT1 (N4073, N4072);
nor NOR4 (N4074, N4059, N3679, N1845, N509);
xor XOR2 (N4075, N4047, N795);
xor XOR2 (N4076, N4070, N706);
nand NAND4 (N4077, N4069, N3772, N2230, N2286);
nor NOR4 (N4078, N4076, N1409, N2214, N354);
and AND2 (N4079, N4075, N1931);
not NOT1 (N4080, N4074);
nand NAND4 (N4081, N4071, N2376, N797, N2221);
xor XOR2 (N4082, N4048, N1344);
nand NAND3 (N4083, N4080, N778, N3535);
xor XOR2 (N4084, N4083, N2560);
buf BUF1 (N4085, N4073);
or OR2 (N4086, N4077, N1378);
nor NOR3 (N4087, N4079, N950, N2338);
xor XOR2 (N4088, N4065, N3068);
not NOT1 (N4089, N4066);
nor NOR3 (N4090, N4088, N1261, N1819);
not NOT1 (N4091, N4090);
buf BUF1 (N4092, N4087);
or OR4 (N4093, N4085, N1075, N1720, N3622);
not NOT1 (N4094, N4093);
xor XOR2 (N4095, N4067, N2501);
buf BUF1 (N4096, N4091);
buf BUF1 (N4097, N4092);
nand NAND2 (N4098, N4095, N3935);
and AND2 (N4099, N4081, N2191);
and AND4 (N4100, N4098, N3649, N1050, N731);
buf BUF1 (N4101, N4097);
or OR2 (N4102, N4101, N3809);
xor XOR2 (N4103, N4094, N1449);
buf BUF1 (N4104, N4096);
and AND4 (N4105, N4084, N1778, N1816, N2905);
xor XOR2 (N4106, N4099, N1634);
xor XOR2 (N4107, N4103, N3214);
or OR2 (N4108, N4082, N1950);
nor NOR3 (N4109, N4086, N3172, N4101);
and AND4 (N4110, N4108, N1908, N2545, N1980);
nand NAND4 (N4111, N4104, N1016, N2662, N2436);
nor NOR3 (N4112, N4102, N1704, N1217);
buf BUF1 (N4113, N4109);
and AND2 (N4114, N4106, N3168);
and AND2 (N4115, N4114, N2096);
buf BUF1 (N4116, N4105);
nor NOR3 (N4117, N4112, N2423, N800);
or OR4 (N4118, N4110, N557, N723, N740);
and AND4 (N4119, N4118, N612, N318, N1550);
not NOT1 (N4120, N4116);
buf BUF1 (N4121, N4117);
and AND2 (N4122, N4089, N2031);
nand NAND2 (N4123, N4115, N1805);
or OR3 (N4124, N4100, N3834, N3462);
or OR2 (N4125, N4078, N1258);
not NOT1 (N4126, N4124);
xor XOR2 (N4127, N4125, N2272);
or OR2 (N4128, N4122, N2148);
nand NAND4 (N4129, N4123, N2142, N3222, N147);
xor XOR2 (N4130, N4129, N580);
nand NAND4 (N4131, N4113, N2277, N2493, N3617);
nor NOR3 (N4132, N4119, N758, N3893);
buf BUF1 (N4133, N4107);
nor NOR2 (N4134, N4127, N3289);
buf BUF1 (N4135, N4126);
not NOT1 (N4136, N4121);
not NOT1 (N4137, N4133);
buf BUF1 (N4138, N4120);
buf BUF1 (N4139, N4131);
xor XOR2 (N4140, N4138, N3059);
buf BUF1 (N4141, N4140);
and AND4 (N4142, N4111, N2348, N3317, N2518);
and AND3 (N4143, N4132, N2468, N3525);
or OR4 (N4144, N4135, N2965, N1530, N1157);
buf BUF1 (N4145, N4134);
buf BUF1 (N4146, N4142);
or OR3 (N4147, N4141, N739, N682);
xor XOR2 (N4148, N4146, N526);
or OR4 (N4149, N4147, N550, N2038, N2530);
xor XOR2 (N4150, N4139, N1640);
and AND2 (N4151, N4144, N1795);
nor NOR2 (N4152, N4151, N1920);
nor NOR2 (N4153, N4130, N3071);
or OR3 (N4154, N4150, N3840, N2001);
and AND4 (N4155, N4136, N3455, N1138, N1763);
not NOT1 (N4156, N4154);
nand NAND3 (N4157, N4152, N303, N2566);
or OR4 (N4158, N4128, N2088, N682, N923);
nor NOR3 (N4159, N4153, N1159, N885);
not NOT1 (N4160, N4157);
xor XOR2 (N4161, N4145, N3993);
nand NAND4 (N4162, N4155, N3165, N4014, N1690);
or OR2 (N4163, N4156, N1130);
xor XOR2 (N4164, N4149, N3604);
not NOT1 (N4165, N4161);
xor XOR2 (N4166, N4164, N350);
not NOT1 (N4167, N4159);
not NOT1 (N4168, N4158);
xor XOR2 (N4169, N4162, N459);
xor XOR2 (N4170, N4166, N400);
xor XOR2 (N4171, N4143, N2014);
nand NAND3 (N4172, N4170, N2809, N2523);
not NOT1 (N4173, N4168);
nor NOR2 (N4174, N4160, N128);
xor XOR2 (N4175, N4171, N16);
or OR4 (N4176, N4175, N739, N4104, N1588);
nand NAND2 (N4177, N4173, N617);
buf BUF1 (N4178, N4165);
nor NOR4 (N4179, N4148, N2492, N1748, N2428);
and AND4 (N4180, N4174, N2873, N849, N2791);
or OR4 (N4181, N4179, N1483, N809, N3274);
buf BUF1 (N4182, N4167);
buf BUF1 (N4183, N4182);
nand NAND4 (N4184, N4172, N946, N1882, N3581);
not NOT1 (N4185, N4180);
buf BUF1 (N4186, N4177);
nor NOR3 (N4187, N4184, N459, N3555);
buf BUF1 (N4188, N4187);
nand NAND2 (N4189, N4185, N3367);
buf BUF1 (N4190, N4137);
xor XOR2 (N4191, N4176, N2212);
not NOT1 (N4192, N4178);
buf BUF1 (N4193, N4191);
or OR4 (N4194, N4193, N657, N1807, N927);
not NOT1 (N4195, N4163);
nor NOR2 (N4196, N4192, N1018);
nand NAND4 (N4197, N4190, N790, N773, N3505);
buf BUF1 (N4198, N4197);
buf BUF1 (N4199, N4186);
or OR3 (N4200, N4199, N3931, N800);
buf BUF1 (N4201, N4195);
xor XOR2 (N4202, N4196, N3712);
and AND2 (N4203, N4183, N2609);
and AND3 (N4204, N4201, N4167, N456);
buf BUF1 (N4205, N4188);
buf BUF1 (N4206, N4200);
not NOT1 (N4207, N4206);
not NOT1 (N4208, N4207);
and AND2 (N4209, N4198, N1898);
or OR2 (N4210, N4194, N2256);
not NOT1 (N4211, N4189);
not NOT1 (N4212, N4210);
nand NAND4 (N4213, N4181, N1518, N1381, N3795);
not NOT1 (N4214, N4212);
not NOT1 (N4215, N4203);
and AND2 (N4216, N4204, N908);
or OR4 (N4217, N4216, N3853, N1002, N1132);
not NOT1 (N4218, N4211);
or OR2 (N4219, N4169, N492);
buf BUF1 (N4220, N4214);
buf BUF1 (N4221, N4202);
buf BUF1 (N4222, N4215);
or OR2 (N4223, N4222, N312);
nor NOR4 (N4224, N4219, N3196, N2081, N4039);
nor NOR3 (N4225, N4221, N3464, N520);
not NOT1 (N4226, N4217);
xor XOR2 (N4227, N4220, N2684);
nor NOR2 (N4228, N4226, N2628);
nand NAND2 (N4229, N4208, N1092);
not NOT1 (N4230, N4213);
not NOT1 (N4231, N4205);
xor XOR2 (N4232, N4225, N2601);
or OR3 (N4233, N4229, N518, N2694);
nand NAND4 (N4234, N4230, N1790, N2935, N3771);
buf BUF1 (N4235, N4223);
nor NOR3 (N4236, N4209, N305, N3606);
not NOT1 (N4237, N4234);
nand NAND2 (N4238, N4231, N2738);
buf BUF1 (N4239, N4236);
or OR3 (N4240, N4232, N3634, N1649);
nor NOR4 (N4241, N4224, N2180, N3885, N901);
and AND3 (N4242, N4227, N2758, N3380);
nand NAND2 (N4243, N4240, N3368);
buf BUF1 (N4244, N4235);
and AND2 (N4245, N4237, N1454);
nand NAND4 (N4246, N4218, N2071, N488, N3926);
not NOT1 (N4247, N4228);
or OR3 (N4248, N4243, N4064, N3012);
nand NAND3 (N4249, N4239, N2295, N3569);
or OR2 (N4250, N4244, N4047);
or OR3 (N4251, N4233, N1133, N3766);
not NOT1 (N4252, N4242);
and AND2 (N4253, N4251, N501);
not NOT1 (N4254, N4238);
buf BUF1 (N4255, N4245);
or OR2 (N4256, N4254, N167);
and AND3 (N4257, N4247, N562, N87);
nand NAND4 (N4258, N4248, N2307, N2912, N3688);
not NOT1 (N4259, N4256);
and AND4 (N4260, N4259, N244, N842, N893);
nand NAND3 (N4261, N4250, N1350, N3426);
nand NAND2 (N4262, N4249, N2189);
nor NOR3 (N4263, N4241, N961, N3113);
not NOT1 (N4264, N4255);
xor XOR2 (N4265, N4263, N2091);
or OR4 (N4266, N4258, N2119, N1171, N2821);
nand NAND3 (N4267, N4252, N2785, N601);
nor NOR2 (N4268, N4265, N1820);
buf BUF1 (N4269, N4257);
and AND4 (N4270, N4261, N3956, N1702, N1594);
nand NAND4 (N4271, N4270, N966, N3534, N1742);
and AND2 (N4272, N4246, N96);
or OR2 (N4273, N4253, N2027);
nor NOR4 (N4274, N4271, N1394, N3751, N689);
not NOT1 (N4275, N4266);
and AND3 (N4276, N4275, N801, N790);
nor NOR4 (N4277, N4268, N3107, N3526, N1946);
nor NOR3 (N4278, N4260, N140, N2069);
not NOT1 (N4279, N4277);
nand NAND2 (N4280, N4267, N3715);
buf BUF1 (N4281, N4280);
nand NAND3 (N4282, N4279, N3512, N2266);
or OR4 (N4283, N4281, N2325, N16, N200);
not NOT1 (N4284, N4264);
nand NAND3 (N4285, N4262, N3119, N5);
buf BUF1 (N4286, N4278);
buf BUF1 (N4287, N4282);
nor NOR3 (N4288, N4284, N3320, N3437);
not NOT1 (N4289, N4285);
buf BUF1 (N4290, N4269);
and AND2 (N4291, N4276, N2713);
nand NAND3 (N4292, N4288, N2997, N4101);
buf BUF1 (N4293, N4273);
nand NAND4 (N4294, N4291, N1382, N1555, N4086);
nor NOR2 (N4295, N4286, N2568);
nor NOR2 (N4296, N4272, N2148);
buf BUF1 (N4297, N4289);
nor NOR2 (N4298, N4295, N2260);
buf BUF1 (N4299, N4297);
buf BUF1 (N4300, N4294);
buf BUF1 (N4301, N4300);
and AND3 (N4302, N4287, N1752, N402);
nand NAND2 (N4303, N4283, N2479);
and AND2 (N4304, N4302, N847);
buf BUF1 (N4305, N4290);
not NOT1 (N4306, N4305);
buf BUF1 (N4307, N4274);
nor NOR3 (N4308, N4307, N327, N4015);
and AND2 (N4309, N4304, N1621);
and AND3 (N4310, N4299, N2686, N1669);
not NOT1 (N4311, N4308);
and AND2 (N4312, N4301, N2289);
or OR2 (N4313, N4292, N960);
xor XOR2 (N4314, N4298, N3767);
and AND3 (N4315, N4314, N838, N73);
buf BUF1 (N4316, N4296);
nor NOR3 (N4317, N4306, N3537, N2631);
buf BUF1 (N4318, N4303);
and AND2 (N4319, N4318, N2446);
not NOT1 (N4320, N4293);
buf BUF1 (N4321, N4311);
xor XOR2 (N4322, N4309, N1774);
not NOT1 (N4323, N4319);
nor NOR3 (N4324, N4315, N4276, N2232);
nor NOR2 (N4325, N4310, N1565);
buf BUF1 (N4326, N4323);
not NOT1 (N4327, N4324);
or OR4 (N4328, N4312, N531, N480, N493);
nor NOR4 (N4329, N4322, N3410, N602, N2186);
and AND3 (N4330, N4329, N2045, N151);
nand NAND2 (N4331, N4328, N1517);
or OR4 (N4332, N4330, N2956, N1850, N2804);
nand NAND3 (N4333, N4317, N1787, N1904);
not NOT1 (N4334, N4326);
or OR3 (N4335, N4333, N921, N2173);
buf BUF1 (N4336, N4313);
buf BUF1 (N4337, N4321);
xor XOR2 (N4338, N4327, N692);
not NOT1 (N4339, N4331);
not NOT1 (N4340, N4325);
and AND4 (N4341, N4335, N3106, N1197, N454);
or OR3 (N4342, N4341, N62, N3430);
buf BUF1 (N4343, N4334);
nor NOR4 (N4344, N4332, N2609, N3768, N2614);
buf BUF1 (N4345, N4340);
xor XOR2 (N4346, N4337, N3780);
nor NOR4 (N4347, N4344, N342, N1893, N3977);
nor NOR2 (N4348, N4346, N1183);
nand NAND3 (N4349, N4345, N627, N1111);
and AND2 (N4350, N4338, N1704);
not NOT1 (N4351, N4347);
xor XOR2 (N4352, N4348, N230);
nor NOR2 (N4353, N4342, N289);
or OR4 (N4354, N4351, N1195, N3553, N246);
buf BUF1 (N4355, N4354);
not NOT1 (N4356, N4350);
buf BUF1 (N4357, N4352);
xor XOR2 (N4358, N4339, N400);
xor XOR2 (N4359, N4316, N2606);
buf BUF1 (N4360, N4355);
or OR3 (N4361, N4349, N3679, N2105);
nor NOR3 (N4362, N4361, N1241, N3540);
or OR3 (N4363, N4343, N563, N802);
xor XOR2 (N4364, N4353, N3449);
and AND2 (N4365, N4362, N1137);
nor NOR2 (N4366, N4356, N1051);
or OR3 (N4367, N4360, N1325, N1263);
xor XOR2 (N4368, N4363, N2662);
or OR4 (N4369, N4358, N2817, N2388, N2675);
nor NOR3 (N4370, N4366, N2633, N3386);
buf BUF1 (N4371, N4336);
or OR3 (N4372, N4365, N3171, N1167);
nand NAND4 (N4373, N4320, N3780, N3237, N1420);
nand NAND3 (N4374, N4372, N2414, N3785);
and AND4 (N4375, N4367, N3605, N1280, N2211);
buf BUF1 (N4376, N4371);
or OR2 (N4377, N4375, N2487);
nor NOR2 (N4378, N4377, N3292);
buf BUF1 (N4379, N4373);
nand NAND2 (N4380, N4364, N3671);
nor NOR3 (N4381, N4357, N4002, N1268);
not NOT1 (N4382, N4359);
or OR2 (N4383, N4369, N967);
xor XOR2 (N4384, N4380, N4228);
nor NOR3 (N4385, N4378, N1613, N1440);
and AND3 (N4386, N4382, N2889, N98);
or OR4 (N4387, N4384, N921, N4032, N283);
and AND3 (N4388, N4368, N2618, N2770);
or OR3 (N4389, N4386, N2831, N3678);
xor XOR2 (N4390, N4374, N613);
and AND3 (N4391, N4389, N3231, N1998);
xor XOR2 (N4392, N4391, N3715);
nor NOR3 (N4393, N4383, N3633, N745);
or OR4 (N4394, N4370, N4287, N2852, N1086);
not NOT1 (N4395, N4376);
nor NOR2 (N4396, N4381, N2230);
nand NAND4 (N4397, N4393, N1056, N3008, N3351);
and AND4 (N4398, N4379, N2137, N2911, N2835);
and AND3 (N4399, N4397, N3793, N4183);
and AND4 (N4400, N4385, N2165, N1626, N369);
nand NAND3 (N4401, N4400, N3085, N2934);
buf BUF1 (N4402, N4388);
and AND3 (N4403, N4390, N198, N2066);
nand NAND3 (N4404, N4394, N4187, N70);
xor XOR2 (N4405, N4387, N2396);
or OR4 (N4406, N4398, N619, N1417, N2111);
xor XOR2 (N4407, N4392, N3926);
and AND3 (N4408, N4406, N3953, N2647);
xor XOR2 (N4409, N4405, N857);
xor XOR2 (N4410, N4407, N986);
xor XOR2 (N4411, N4399, N816);
not NOT1 (N4412, N4395);
xor XOR2 (N4413, N4409, N4401);
buf BUF1 (N4414, N1691);
nand NAND3 (N4415, N4412, N1237, N4146);
and AND2 (N4416, N4410, N4082);
not NOT1 (N4417, N4414);
and AND2 (N4418, N4396, N4324);
or OR4 (N4419, N4417, N2149, N2127, N2409);
buf BUF1 (N4420, N4404);
or OR4 (N4421, N4413, N2242, N4352, N3446);
xor XOR2 (N4422, N4416, N1949);
and AND3 (N4423, N4418, N1769, N4089);
or OR3 (N4424, N4422, N1866, N1374);
xor XOR2 (N4425, N4402, N816);
xor XOR2 (N4426, N4421, N296);
not NOT1 (N4427, N4415);
not NOT1 (N4428, N4427);
not NOT1 (N4429, N4419);
xor XOR2 (N4430, N4403, N4315);
or OR3 (N4431, N4430, N2732, N575);
nand NAND2 (N4432, N4428, N3653);
or OR2 (N4433, N4424, N3352);
or OR2 (N4434, N4408, N2145);
not NOT1 (N4435, N4425);
and AND2 (N4436, N4429, N287);
xor XOR2 (N4437, N4431, N714);
buf BUF1 (N4438, N4435);
xor XOR2 (N4439, N4426, N752);
nand NAND4 (N4440, N4439, N2514, N2871, N3005);
not NOT1 (N4441, N4411);
nor NOR4 (N4442, N4423, N347, N210, N4285);
nor NOR4 (N4443, N4434, N4198, N2962, N3500);
and AND4 (N4444, N4420, N2450, N1915, N1165);
nand NAND2 (N4445, N4441, N392);
buf BUF1 (N4446, N4437);
and AND2 (N4447, N4440, N1053);
and AND2 (N4448, N4444, N2809);
or OR2 (N4449, N4446, N1595);
buf BUF1 (N4450, N4438);
or OR2 (N4451, N4445, N637);
or OR3 (N4452, N4436, N1007, N615);
nor NOR4 (N4453, N4447, N497, N2823, N3303);
or OR3 (N4454, N4432, N989, N367);
nor NOR3 (N4455, N4448, N909, N2713);
xor XOR2 (N4456, N4443, N1529);
or OR2 (N4457, N4453, N1180);
nor NOR4 (N4458, N4433, N3022, N175, N4171);
xor XOR2 (N4459, N4451, N563);
xor XOR2 (N4460, N4452, N2614);
or OR2 (N4461, N4456, N1479);
not NOT1 (N4462, N4449);
nor NOR3 (N4463, N4442, N644, N326);
not NOT1 (N4464, N4454);
buf BUF1 (N4465, N4450);
and AND3 (N4466, N4458, N1371, N2831);
xor XOR2 (N4467, N4461, N1564);
or OR4 (N4468, N4460, N3705, N1639, N4433);
xor XOR2 (N4469, N4459, N215);
buf BUF1 (N4470, N4463);
or OR2 (N4471, N4465, N3547);
or OR2 (N4472, N4470, N1047);
not NOT1 (N4473, N4467);
or OR4 (N4474, N4455, N2547, N4150, N1745);
xor XOR2 (N4475, N4457, N21);
xor XOR2 (N4476, N4474, N3833);
buf BUF1 (N4477, N4473);
not NOT1 (N4478, N4468);
and AND2 (N4479, N4478, N3666);
or OR3 (N4480, N4464, N3994, N2224);
nor NOR3 (N4481, N4476, N873, N1065);
buf BUF1 (N4482, N4481);
buf BUF1 (N4483, N4466);
buf BUF1 (N4484, N4479);
xor XOR2 (N4485, N4483, N932);
buf BUF1 (N4486, N4475);
xor XOR2 (N4487, N4484, N2229);
or OR2 (N4488, N4485, N3331);
or OR2 (N4489, N4471, N2427);
not NOT1 (N4490, N4489);
xor XOR2 (N4491, N4469, N1739);
or OR3 (N4492, N4462, N2651, N1342);
buf BUF1 (N4493, N4482);
nand NAND4 (N4494, N4472, N1421, N553, N1648);
not NOT1 (N4495, N4477);
and AND3 (N4496, N4493, N4092, N3932);
not NOT1 (N4497, N4491);
nand NAND3 (N4498, N4494, N1069, N4032);
xor XOR2 (N4499, N4487, N1461);
and AND2 (N4500, N4490, N1626);
or OR4 (N4501, N4499, N1801, N58, N3465);
nand NAND4 (N4502, N4500, N787, N1284, N2139);
nand NAND2 (N4503, N4492, N4005);
xor XOR2 (N4504, N4497, N4249);
not NOT1 (N4505, N4496);
nand NAND3 (N4506, N4486, N4486, N2748);
nand NAND2 (N4507, N4505, N2752);
and AND4 (N4508, N4501, N1085, N1195, N1402);
nor NOR4 (N4509, N4508, N984, N3265, N1202);
and AND4 (N4510, N4488, N3623, N1627, N2476);
or OR4 (N4511, N4503, N4129, N499, N750);
and AND2 (N4512, N4506, N1026);
or OR2 (N4513, N4512, N3678);
xor XOR2 (N4514, N4480, N2995);
buf BUF1 (N4515, N4495);
xor XOR2 (N4516, N4513, N3534);
buf BUF1 (N4517, N4509);
nor NOR3 (N4518, N4516, N3873, N3861);
xor XOR2 (N4519, N4498, N3138);
or OR4 (N4520, N4518, N4480, N4267, N301);
and AND2 (N4521, N4502, N2336);
and AND3 (N4522, N4515, N1936, N3168);
or OR2 (N4523, N4514, N1286);
nand NAND2 (N4524, N4523, N3573);
nand NAND2 (N4525, N4519, N2766);
buf BUF1 (N4526, N4521);
buf BUF1 (N4527, N4517);
nor NOR3 (N4528, N4527, N167, N1619);
xor XOR2 (N4529, N4507, N2527);
nand NAND2 (N4530, N4504, N2675);
or OR3 (N4531, N4520, N734, N2884);
or OR3 (N4532, N4531, N4150, N1331);
not NOT1 (N4533, N4522);
or OR3 (N4534, N4524, N1525, N3814);
or OR3 (N4535, N4533, N3273, N971);
or OR3 (N4536, N4528, N2150, N162);
nand NAND2 (N4537, N4510, N3139);
not NOT1 (N4538, N4526);
and AND3 (N4539, N4532, N868, N176);
not NOT1 (N4540, N4511);
nand NAND3 (N4541, N4530, N1454, N3031);
buf BUF1 (N4542, N4529);
xor XOR2 (N4543, N4537, N4201);
xor XOR2 (N4544, N4535, N1908);
or OR4 (N4545, N4544, N4073, N229, N3006);
nand NAND3 (N4546, N4538, N2784, N1022);
nor NOR2 (N4547, N4536, N2171);
not NOT1 (N4548, N4541);
nor NOR3 (N4549, N4546, N3276, N31);
not NOT1 (N4550, N4543);
buf BUF1 (N4551, N4550);
buf BUF1 (N4552, N4542);
and AND4 (N4553, N4548, N1025, N2925, N2553);
xor XOR2 (N4554, N4553, N3806);
and AND3 (N4555, N4540, N4202, N3013);
not NOT1 (N4556, N4534);
not NOT1 (N4557, N4549);
buf BUF1 (N4558, N4525);
and AND4 (N4559, N4556, N38, N1248, N1045);
or OR3 (N4560, N4559, N4386, N4115);
nor NOR2 (N4561, N4560, N718);
not NOT1 (N4562, N4554);
xor XOR2 (N4563, N4552, N558);
nand NAND4 (N4564, N4562, N3209, N3174, N2536);
buf BUF1 (N4565, N4551);
buf BUF1 (N4566, N4565);
nor NOR4 (N4567, N4561, N502, N606, N3199);
buf BUF1 (N4568, N4545);
nor NOR3 (N4569, N4539, N573, N898);
nand NAND2 (N4570, N4569, N1122);
or OR2 (N4571, N4568, N904);
nand NAND4 (N4572, N4563, N3879, N48, N3748);
and AND3 (N4573, N4564, N60, N333);
xor XOR2 (N4574, N4567, N596);
or OR3 (N4575, N4555, N3348, N3330);
not NOT1 (N4576, N4574);
buf BUF1 (N4577, N4573);
nand NAND2 (N4578, N4557, N813);
nand NAND2 (N4579, N4578, N998);
xor XOR2 (N4580, N4571, N3227);
xor XOR2 (N4581, N4547, N1743);
buf BUF1 (N4582, N4575);
xor XOR2 (N4583, N4577, N946);
buf BUF1 (N4584, N4572);
and AND2 (N4585, N4566, N3822);
nand NAND4 (N4586, N4581, N598, N3392, N2901);
nand NAND2 (N4587, N4584, N3188);
nand NAND2 (N4588, N4583, N415);
nand NAND4 (N4589, N4586, N3102, N4093, N456);
not NOT1 (N4590, N4580);
buf BUF1 (N4591, N4570);
nor NOR2 (N4592, N4591, N1046);
and AND4 (N4593, N4590, N844, N1456, N3113);
buf BUF1 (N4594, N4587);
buf BUF1 (N4595, N4592);
nand NAND4 (N4596, N4595, N1408, N10, N2600);
xor XOR2 (N4597, N4585, N1869);
buf BUF1 (N4598, N4582);
not NOT1 (N4599, N4579);
and AND3 (N4600, N4598, N3847, N1472);
nor NOR3 (N4601, N4597, N979, N2889);
xor XOR2 (N4602, N4594, N3694);
not NOT1 (N4603, N4593);
or OR3 (N4604, N4576, N1502, N1030);
xor XOR2 (N4605, N4558, N3900);
xor XOR2 (N4606, N4605, N1353);
not NOT1 (N4607, N4599);
nor NOR2 (N4608, N4601, N1967);
and AND3 (N4609, N4596, N1173, N1388);
nand NAND4 (N4610, N4603, N1548, N441, N1866);
buf BUF1 (N4611, N4608);
or OR3 (N4612, N4600, N752, N177);
nand NAND4 (N4613, N4589, N1464, N2000, N3155);
nor NOR2 (N4614, N4602, N1399);
and AND3 (N4615, N4606, N1950, N229);
not NOT1 (N4616, N4609);
nor NOR3 (N4617, N4612, N2932, N1187);
or OR4 (N4618, N4615, N1967, N1657, N1181);
nand NAND4 (N4619, N4618, N1025, N4200, N2056);
or OR3 (N4620, N4607, N671, N1782);
and AND4 (N4621, N4611, N4547, N4228, N3097);
xor XOR2 (N4622, N4610, N3987);
buf BUF1 (N4623, N4616);
nor NOR4 (N4624, N4620, N175, N1111, N2841);
not NOT1 (N4625, N4621);
or OR4 (N4626, N4614, N3317, N1701, N4204);
or OR3 (N4627, N4623, N3470, N82);
and AND3 (N4628, N4622, N1690, N4241);
nor NOR4 (N4629, N4617, N290, N2476, N1113);
or OR4 (N4630, N4613, N1120, N3162, N2290);
buf BUF1 (N4631, N4588);
xor XOR2 (N4632, N4630, N189);
and AND3 (N4633, N4624, N4312, N4039);
xor XOR2 (N4634, N4629, N2678);
xor XOR2 (N4635, N4619, N1694);
xor XOR2 (N4636, N4625, N2794);
and AND2 (N4637, N4636, N3514);
xor XOR2 (N4638, N4627, N1907);
not NOT1 (N4639, N4632);
and AND3 (N4640, N4604, N4101, N2082);
nand NAND3 (N4641, N4633, N976, N1654);
xor XOR2 (N4642, N4634, N4248);
buf BUF1 (N4643, N4637);
nand NAND3 (N4644, N4631, N1794, N364);
xor XOR2 (N4645, N4639, N1330);
nor NOR2 (N4646, N4642, N2508);
not NOT1 (N4647, N4641);
or OR2 (N4648, N4628, N2587);
nand NAND2 (N4649, N4646, N462);
and AND3 (N4650, N4645, N3622, N913);
nand NAND2 (N4651, N4638, N1804);
and AND3 (N4652, N4640, N4486, N3393);
or OR4 (N4653, N4643, N2426, N2124, N3991);
and AND3 (N4654, N4626, N4158, N3208);
buf BUF1 (N4655, N4647);
and AND2 (N4656, N4648, N2460);
xor XOR2 (N4657, N4650, N1832);
and AND3 (N4658, N4635, N2446, N4088);
xor XOR2 (N4659, N4652, N3649);
nor NOR3 (N4660, N4657, N4507, N1321);
nand NAND4 (N4661, N4658, N1922, N4654, N1425);
xor XOR2 (N4662, N1507, N3294);
or OR2 (N4663, N4656, N64);
buf BUF1 (N4664, N4659);
xor XOR2 (N4665, N4662, N4032);
nor NOR2 (N4666, N4649, N2303);
and AND2 (N4667, N4665, N1913);
xor XOR2 (N4668, N4667, N4120);
not NOT1 (N4669, N4668);
xor XOR2 (N4670, N4653, N3941);
nor NOR3 (N4671, N4669, N2714, N1641);
nand NAND3 (N4672, N4651, N1561, N1599);
nand NAND4 (N4673, N4661, N1679, N1010, N985);
not NOT1 (N4674, N4666);
xor XOR2 (N4675, N4671, N1732);
nor NOR4 (N4676, N4674, N1734, N3748, N2751);
or OR3 (N4677, N4673, N4137, N4291);
xor XOR2 (N4678, N4664, N843);
nor NOR4 (N4679, N4678, N3449, N3426, N3673);
nor NOR3 (N4680, N4655, N3029, N3530);
not NOT1 (N4681, N4670);
or OR2 (N4682, N4676, N3954);
xor XOR2 (N4683, N4679, N1762);
xor XOR2 (N4684, N4644, N1062);
and AND3 (N4685, N4677, N4425, N4461);
nor NOR2 (N4686, N4672, N470);
nor NOR2 (N4687, N4683, N2429);
or OR3 (N4688, N4687, N1999, N3079);
not NOT1 (N4689, N4682);
not NOT1 (N4690, N4685);
buf BUF1 (N4691, N4663);
nor NOR3 (N4692, N4690, N3, N4365);
nand NAND3 (N4693, N4680, N4255, N3141);
nor NOR2 (N4694, N4675, N4367);
nand NAND3 (N4695, N4692, N2793, N4036);
buf BUF1 (N4696, N4681);
buf BUF1 (N4697, N4686);
buf BUF1 (N4698, N4695);
or OR3 (N4699, N4697, N715, N4158);
buf BUF1 (N4700, N4694);
xor XOR2 (N4701, N4700, N4400);
nand NAND4 (N4702, N4689, N4247, N289, N2276);
or OR3 (N4703, N4698, N120, N676);
nor NOR3 (N4704, N4660, N1747, N1550);
or OR2 (N4705, N4699, N4034);
xor XOR2 (N4706, N4688, N96);
and AND2 (N4707, N4705, N1284);
nand NAND2 (N4708, N4703, N1133);
nand NAND2 (N4709, N4701, N2371);
nor NOR4 (N4710, N4684, N3729, N2109, N1522);
and AND2 (N4711, N4691, N2770);
nor NOR2 (N4712, N4711, N634);
and AND3 (N4713, N4708, N1688, N4402);
xor XOR2 (N4714, N4704, N1329);
xor XOR2 (N4715, N4707, N3624);
nor NOR2 (N4716, N4715, N4683);
nor NOR4 (N4717, N4710, N265, N187, N802);
or OR4 (N4718, N4712, N1798, N4398, N3428);
buf BUF1 (N4719, N4716);
not NOT1 (N4720, N4717);
not NOT1 (N4721, N4713);
or OR2 (N4722, N4702, N2540);
or OR2 (N4723, N4693, N2741);
or OR2 (N4724, N4719, N2182);
nand NAND2 (N4725, N4718, N1854);
nand NAND2 (N4726, N4709, N2078);
nor NOR4 (N4727, N4723, N1150, N4319, N3977);
not NOT1 (N4728, N4696);
xor XOR2 (N4729, N4721, N4145);
xor XOR2 (N4730, N4729, N2546);
and AND3 (N4731, N4730, N1123, N131);
and AND4 (N4732, N4714, N3332, N707, N871);
nor NOR2 (N4733, N4720, N3646);
and AND3 (N4734, N4733, N3063, N1617);
nor NOR3 (N4735, N4722, N283, N155);
nand NAND2 (N4736, N4731, N4405);
nand NAND3 (N4737, N4727, N1087, N1946);
nand NAND3 (N4738, N4706, N894, N4212);
nor NOR2 (N4739, N4737, N2517);
buf BUF1 (N4740, N4736);
xor XOR2 (N4741, N4726, N1552);
not NOT1 (N4742, N4725);
or OR2 (N4743, N4735, N2165);
nand NAND3 (N4744, N4741, N875, N894);
not NOT1 (N4745, N4739);
xor XOR2 (N4746, N4744, N2798);
nor NOR4 (N4747, N4724, N3955, N3113, N3819);
xor XOR2 (N4748, N4745, N1740);
nand NAND3 (N4749, N4743, N1855, N4663);
buf BUF1 (N4750, N4746);
nand NAND3 (N4751, N4728, N4651, N2552);
nor NOR2 (N4752, N4750, N985);
not NOT1 (N4753, N4751);
nor NOR4 (N4754, N4742, N1651, N3015, N3093);
xor XOR2 (N4755, N4749, N4092);
or OR2 (N4756, N4753, N3442);
not NOT1 (N4757, N4738);
or OR2 (N4758, N4748, N768);
nor NOR2 (N4759, N4734, N1691);
nand NAND2 (N4760, N4740, N1041);
not NOT1 (N4761, N4754);
and AND2 (N4762, N4760, N4460);
not NOT1 (N4763, N4757);
and AND3 (N4764, N4759, N4543, N983);
buf BUF1 (N4765, N4755);
not NOT1 (N4766, N4764);
xor XOR2 (N4767, N4762, N507);
buf BUF1 (N4768, N4763);
buf BUF1 (N4769, N4765);
and AND3 (N4770, N4769, N163, N525);
not NOT1 (N4771, N4767);
nand NAND2 (N4772, N4761, N3107);
and AND4 (N4773, N4772, N4770, N737, N1458);
and AND4 (N4774, N144, N950, N2414, N968);
nor NOR3 (N4775, N4747, N2135, N2925);
not NOT1 (N4776, N4766);
xor XOR2 (N4777, N4776, N1144);
and AND4 (N4778, N4775, N3704, N2976, N1091);
buf BUF1 (N4779, N4756);
buf BUF1 (N4780, N4732);
nor NOR2 (N4781, N4780, N261);
buf BUF1 (N4782, N4768);
not NOT1 (N4783, N4781);
not NOT1 (N4784, N4782);
nand NAND3 (N4785, N4774, N4541, N3524);
xor XOR2 (N4786, N4771, N4670);
xor XOR2 (N4787, N4777, N2359);
nand NAND4 (N4788, N4752, N572, N2155, N1139);
and AND2 (N4789, N4787, N3579);
not NOT1 (N4790, N4778);
buf BUF1 (N4791, N4783);
or OR3 (N4792, N4779, N2243, N2);
nand NAND4 (N4793, N4786, N711, N121, N4582);
nor NOR2 (N4794, N4789, N3262);
or OR4 (N4795, N4758, N582, N1556, N2799);
or OR4 (N4796, N4785, N1096, N3476, N327);
nor NOR4 (N4797, N4794, N460, N4289, N2993);
and AND2 (N4798, N4784, N2453);
xor XOR2 (N4799, N4788, N3434);
nor NOR3 (N4800, N4798, N3000, N3229);
nand NAND4 (N4801, N4773, N3895, N3273, N3422);
nand NAND3 (N4802, N4800, N2561, N2823);
xor XOR2 (N4803, N4793, N4294);
xor XOR2 (N4804, N4803, N1996);
nor NOR2 (N4805, N4795, N4038);
buf BUF1 (N4806, N4797);
xor XOR2 (N4807, N4792, N3593);
buf BUF1 (N4808, N4791);
xor XOR2 (N4809, N4799, N4165);
not NOT1 (N4810, N4808);
and AND3 (N4811, N4806, N2500, N4557);
nand NAND3 (N4812, N4809, N2033, N4773);
or OR2 (N4813, N4804, N600);
and AND4 (N4814, N4807, N4067, N1982, N1513);
buf BUF1 (N4815, N4796);
xor XOR2 (N4816, N4810, N1491);
xor XOR2 (N4817, N4816, N1005);
nand NAND2 (N4818, N4813, N4817);
not NOT1 (N4819, N1327);
buf BUF1 (N4820, N4790);
not NOT1 (N4821, N4801);
not NOT1 (N4822, N4818);
or OR4 (N4823, N4821, N2667, N4563, N2970);
or OR4 (N4824, N4823, N43, N1440, N88);
nand NAND3 (N4825, N4812, N4566, N321);
buf BUF1 (N4826, N4815);
nor NOR4 (N4827, N4824, N3427, N3578, N3043);
nor NOR4 (N4828, N4814, N1278, N1971, N1290);
nor NOR2 (N4829, N4827, N148);
or OR3 (N4830, N4826, N3017, N237);
nor NOR3 (N4831, N4820, N2801, N892);
or OR3 (N4832, N4829, N2634, N4212);
xor XOR2 (N4833, N4802, N4790);
nand NAND4 (N4834, N4825, N3313, N1147, N2288);
buf BUF1 (N4835, N4828);
buf BUF1 (N4836, N4832);
buf BUF1 (N4837, N4822);
not NOT1 (N4838, N4831);
or OR3 (N4839, N4837, N4202, N3269);
and AND2 (N4840, N4833, N2905);
buf BUF1 (N4841, N4805);
nand NAND3 (N4842, N4839, N3624, N3330);
not NOT1 (N4843, N4811);
or OR4 (N4844, N4840, N228, N812, N2082);
xor XOR2 (N4845, N4834, N2253);
or OR2 (N4846, N4836, N4777);
xor XOR2 (N4847, N4844, N2123);
buf BUF1 (N4848, N4835);
nor NOR3 (N4849, N4843, N4721, N1975);
or OR4 (N4850, N4842, N302, N1265, N3571);
xor XOR2 (N4851, N4838, N3349);
and AND2 (N4852, N4851, N2514);
nor NOR4 (N4853, N4849, N1469, N2164, N582);
nor NOR2 (N4854, N4846, N661);
or OR4 (N4855, N4830, N4434, N919, N3621);
nor NOR2 (N4856, N4850, N4723);
nand NAND4 (N4857, N4854, N19, N759, N2740);
or OR3 (N4858, N4841, N4405, N3401);
buf BUF1 (N4859, N4853);
or OR2 (N4860, N4859, N3545);
and AND4 (N4861, N4857, N4654, N4275, N461);
nor NOR4 (N4862, N4847, N2712, N2693, N4447);
buf BUF1 (N4863, N4852);
not NOT1 (N4864, N4856);
not NOT1 (N4865, N4862);
nand NAND4 (N4866, N4864, N773, N3208, N1370);
nand NAND4 (N4867, N4863, N4666, N4774, N2884);
nand NAND4 (N4868, N4845, N3862, N4382, N2346);
xor XOR2 (N4869, N4861, N3117);
or OR2 (N4870, N4865, N4541);
not NOT1 (N4871, N4848);
xor XOR2 (N4872, N4869, N3892);
nand NAND3 (N4873, N4867, N22, N2993);
buf BUF1 (N4874, N4866);
nor NOR2 (N4875, N4873, N585);
nor NOR4 (N4876, N4860, N1211, N2742, N4376);
nand NAND4 (N4877, N4871, N1022, N482, N3930);
nand NAND4 (N4878, N4876, N454, N4234, N3301);
not NOT1 (N4879, N4872);
buf BUF1 (N4880, N4878);
nor NOR3 (N4881, N4819, N1686, N4828);
nand NAND3 (N4882, N4868, N647, N1266);
nand NAND4 (N4883, N4870, N263, N4430, N3758);
or OR3 (N4884, N4858, N1903, N145);
nor NOR2 (N4885, N4884, N1550);
nor NOR4 (N4886, N4880, N2853, N221, N2098);
not NOT1 (N4887, N4855);
nor NOR3 (N4888, N4875, N2185, N4020);
and AND3 (N4889, N4877, N882, N2070);
not NOT1 (N4890, N4889);
and AND2 (N4891, N4883, N3394);
and AND2 (N4892, N4885, N236);
not NOT1 (N4893, N4890);
buf BUF1 (N4894, N4882);
xor XOR2 (N4895, N4894, N4143);
buf BUF1 (N4896, N4891);
nor NOR2 (N4897, N4886, N1323);
nor NOR2 (N4898, N4887, N1502);
xor XOR2 (N4899, N4874, N1871);
not NOT1 (N4900, N4895);
not NOT1 (N4901, N4888);
buf BUF1 (N4902, N4899);
nor NOR4 (N4903, N4896, N989, N1601, N467);
xor XOR2 (N4904, N4898, N4121);
xor XOR2 (N4905, N4881, N2666);
nor NOR3 (N4906, N4902, N4276, N4159);
nand NAND4 (N4907, N4906, N4411, N4337, N2950);
not NOT1 (N4908, N4900);
nand NAND4 (N4909, N4903, N3387, N2254, N2666);
xor XOR2 (N4910, N4901, N3487);
xor XOR2 (N4911, N4904, N3456);
nor NOR4 (N4912, N4905, N1619, N75, N4777);
nand NAND2 (N4913, N4910, N2904);
nand NAND3 (N4914, N4912, N2556, N4145);
nor NOR2 (N4915, N4879, N2043);
not NOT1 (N4916, N4911);
nand NAND3 (N4917, N4897, N1278, N4860);
nand NAND4 (N4918, N4909, N4455, N3144, N3857);
xor XOR2 (N4919, N4907, N262);
and AND3 (N4920, N4913, N3392, N130);
buf BUF1 (N4921, N4892);
and AND3 (N4922, N4918, N2133, N3366);
buf BUF1 (N4923, N4920);
not NOT1 (N4924, N4917);
or OR3 (N4925, N4924, N3758, N2744);
or OR4 (N4926, N4914, N128, N3763, N140);
xor XOR2 (N4927, N4921, N2764);
xor XOR2 (N4928, N4922, N321);
or OR2 (N4929, N4927, N1443);
and AND2 (N4930, N4923, N915);
buf BUF1 (N4931, N4928);
nand NAND2 (N4932, N4930, N3970);
xor XOR2 (N4933, N4893, N115);
and AND3 (N4934, N4926, N2581, N4910);
buf BUF1 (N4935, N4919);
or OR3 (N4936, N4935, N1883, N3579);
not NOT1 (N4937, N4936);
buf BUF1 (N4938, N4925);
not NOT1 (N4939, N4933);
nand NAND3 (N4940, N4934, N141, N3588);
buf BUF1 (N4941, N4932);
or OR4 (N4942, N4929, N4367, N3724, N3110);
not NOT1 (N4943, N4938);
nand NAND3 (N4944, N4941, N1397, N339);
nand NAND3 (N4945, N4937, N278, N712);
and AND2 (N4946, N4931, N709);
xor XOR2 (N4947, N4943, N1979);
or OR4 (N4948, N4939, N2490, N1984, N1152);
nand NAND3 (N4949, N4948, N1227, N1329);
nand NAND2 (N4950, N4944, N309);
or OR2 (N4951, N4946, N4620);
not NOT1 (N4952, N4951);
not NOT1 (N4953, N4950);
nor NOR4 (N4954, N4952, N4476, N1512, N720);
or OR2 (N4955, N4947, N4779);
not NOT1 (N4956, N4945);
not NOT1 (N4957, N4954);
not NOT1 (N4958, N4956);
buf BUF1 (N4959, N4942);
buf BUF1 (N4960, N4908);
xor XOR2 (N4961, N4957, N3802);
buf BUF1 (N4962, N4915);
or OR4 (N4963, N4959, N4139, N4730, N3185);
nand NAND4 (N4964, N4955, N1730, N2369, N3357);
and AND3 (N4965, N4963, N2402, N4890);
nor NOR4 (N4966, N4916, N1809, N4906, N443);
xor XOR2 (N4967, N4960, N1524);
xor XOR2 (N4968, N4940, N1344);
buf BUF1 (N4969, N4962);
xor XOR2 (N4970, N4965, N4460);
not NOT1 (N4971, N4964);
or OR4 (N4972, N4953, N3414, N1248, N4454);
or OR3 (N4973, N4958, N1408, N943);
nand NAND3 (N4974, N4967, N3142, N2966);
or OR3 (N4975, N4974, N4307, N4013);
not NOT1 (N4976, N4970);
xor XOR2 (N4977, N4949, N3614);
nor NOR3 (N4978, N4961, N975, N611);
xor XOR2 (N4979, N4971, N4445);
xor XOR2 (N4980, N4979, N3296);
and AND3 (N4981, N4978, N1949, N3962);
buf BUF1 (N4982, N4966);
buf BUF1 (N4983, N4972);
nor NOR4 (N4984, N4982, N3555, N563, N1393);
buf BUF1 (N4985, N4975);
not NOT1 (N4986, N4980);
and AND2 (N4987, N4968, N2164);
or OR4 (N4988, N4981, N803, N3991, N3812);
xor XOR2 (N4989, N4987, N135);
not NOT1 (N4990, N4989);
nor NOR2 (N4991, N4977, N2460);
xor XOR2 (N4992, N4983, N3359);
nor NOR2 (N4993, N4988, N3619);
nand NAND3 (N4994, N4993, N540, N4743);
not NOT1 (N4995, N4969);
nor NOR4 (N4996, N4984, N2238, N2353, N4961);
buf BUF1 (N4997, N4996);
or OR4 (N4998, N4976, N3057, N4986, N1004);
or OR2 (N4999, N2957, N1287);
xor XOR2 (N5000, N4997, N116);
nand NAND2 (N5001, N4994, N2313);
nand NAND4 (N5002, N4992, N2209, N4413, N398);
and AND4 (N5003, N4999, N2885, N2898, N3027);
not NOT1 (N5004, N5000);
or OR3 (N5005, N4985, N4461, N2605);
not NOT1 (N5006, N5002);
nand NAND2 (N5007, N5004, N906);
xor XOR2 (N5008, N5001, N4502);
nor NOR4 (N5009, N4991, N1016, N3134, N3321);
not NOT1 (N5010, N5003);
nand NAND2 (N5011, N5005, N1459);
buf BUF1 (N5012, N5010);
nor NOR3 (N5013, N4998, N246, N1577);
and AND2 (N5014, N5007, N423);
and AND3 (N5015, N5013, N1629, N4152);
nand NAND3 (N5016, N5008, N1078, N2575);
nand NAND4 (N5017, N5011, N2536, N1776, N3065);
xor XOR2 (N5018, N5017, N4619);
xor XOR2 (N5019, N5018, N604);
not NOT1 (N5020, N5015);
not NOT1 (N5021, N5020);
not NOT1 (N5022, N5006);
nor NOR3 (N5023, N4995, N2235, N3685);
buf BUF1 (N5024, N4990);
and AND4 (N5025, N4973, N1665, N3342, N2571);
and AND4 (N5026, N5024, N4575, N4812, N855);
or OR3 (N5027, N5025, N934, N4087);
not NOT1 (N5028, N5021);
buf BUF1 (N5029, N5023);
not NOT1 (N5030, N5026);
and AND3 (N5031, N5016, N1366, N267);
or OR3 (N5032, N5012, N2336, N148);
nor NOR2 (N5033, N5019, N189);
buf BUF1 (N5034, N5009);
nand NAND2 (N5035, N5034, N1191);
or OR3 (N5036, N5029, N4907, N5011);
or OR4 (N5037, N5036, N1896, N2404, N3689);
or OR2 (N5038, N5014, N4188);
nor NOR2 (N5039, N5032, N820);
or OR4 (N5040, N5038, N4493, N701, N2167);
or OR4 (N5041, N5040, N2867, N2370, N452);
nand NAND3 (N5042, N5031, N3394, N315);
xor XOR2 (N5043, N5030, N1022);
nor NOR2 (N5044, N5035, N2318);
buf BUF1 (N5045, N5022);
nand NAND2 (N5046, N5044, N206);
nor NOR3 (N5047, N5041, N3258, N3325);
buf BUF1 (N5048, N5039);
xor XOR2 (N5049, N5046, N4563);
nor NOR2 (N5050, N5027, N3795);
xor XOR2 (N5051, N5047, N4359);
or OR4 (N5052, N5037, N1562, N3826, N3004);
xor XOR2 (N5053, N5048, N343);
or OR2 (N5054, N5042, N2935);
not NOT1 (N5055, N5053);
buf BUF1 (N5056, N5033);
and AND2 (N5057, N5045, N1311);
or OR3 (N5058, N5052, N1918, N1768);
or OR3 (N5059, N5050, N341, N2706);
not NOT1 (N5060, N5043);
nand NAND2 (N5061, N5058, N4211);
nand NAND2 (N5062, N5051, N2108);
or OR2 (N5063, N5057, N2012);
and AND2 (N5064, N5049, N2756);
or OR3 (N5065, N5055, N2392, N2400);
nor NOR2 (N5066, N5054, N3351);
or OR2 (N5067, N5028, N2007);
or OR4 (N5068, N5065, N1063, N1237, N2270);
xor XOR2 (N5069, N5064, N994);
and AND4 (N5070, N5068, N4917, N4303, N571);
or OR2 (N5071, N5067, N1371);
buf BUF1 (N5072, N5063);
or OR4 (N5073, N5066, N3488, N3756, N4703);
buf BUF1 (N5074, N5056);
xor XOR2 (N5075, N5073, N4519);
not NOT1 (N5076, N5070);
buf BUF1 (N5077, N5071);
and AND4 (N5078, N5074, N3652, N1462, N603);
nor NOR3 (N5079, N5062, N854, N4244);
xor XOR2 (N5080, N5077, N3263);
buf BUF1 (N5081, N5075);
or OR3 (N5082, N5076, N1563, N4391);
nand NAND3 (N5083, N5078, N4008, N4165);
nor NOR3 (N5084, N5060, N4015, N4744);
xor XOR2 (N5085, N5069, N4017);
and AND3 (N5086, N5082, N1942, N1718);
nand NAND3 (N5087, N5081, N440, N939);
buf BUF1 (N5088, N5086);
buf BUF1 (N5089, N5084);
or OR2 (N5090, N5085, N1754);
buf BUF1 (N5091, N5083);
buf BUF1 (N5092, N5090);
nor NOR4 (N5093, N5089, N1711, N1217, N1591);
or OR4 (N5094, N5080, N4676, N176, N3322);
or OR2 (N5095, N5059, N3670);
nand NAND4 (N5096, N5079, N1398, N4073, N3437);
xor XOR2 (N5097, N5095, N5023);
nand NAND4 (N5098, N5096, N3587, N544, N2041);
nand NAND2 (N5099, N5091, N1791);
buf BUF1 (N5100, N5088);
not NOT1 (N5101, N5099);
and AND3 (N5102, N5087, N3109, N151);
buf BUF1 (N5103, N5100);
xor XOR2 (N5104, N5061, N1387);
xor XOR2 (N5105, N5103, N634);
and AND4 (N5106, N5102, N391, N3880, N599);
nand NAND4 (N5107, N5105, N1862, N3979, N3779);
nand NAND2 (N5108, N5106, N3617);
buf BUF1 (N5109, N5108);
or OR4 (N5110, N5093, N2045, N3646, N3375);
xor XOR2 (N5111, N5110, N126);
nor NOR4 (N5112, N5107, N2212, N538, N4649);
buf BUF1 (N5113, N5072);
or OR3 (N5114, N5094, N1416, N1892);
not NOT1 (N5115, N5111);
buf BUF1 (N5116, N5113);
not NOT1 (N5117, N5104);
not NOT1 (N5118, N5109);
or OR4 (N5119, N5101, N4018, N3021, N3515);
xor XOR2 (N5120, N5115, N3116);
nand NAND2 (N5121, N5119, N4252);
not NOT1 (N5122, N5116);
and AND2 (N5123, N5121, N3972);
nor NOR3 (N5124, N5117, N1173, N215);
nand NAND4 (N5125, N5098, N3990, N5123, N2480);
nor NOR2 (N5126, N985, N2965);
xor XOR2 (N5127, N5122, N5103);
and AND2 (N5128, N5118, N529);
xor XOR2 (N5129, N5128, N2879);
and AND4 (N5130, N5126, N2775, N554, N2701);
buf BUF1 (N5131, N5112);
nor NOR4 (N5132, N5114, N3679, N3179, N4604);
nor NOR4 (N5133, N5092, N2308, N3140, N3779);
not NOT1 (N5134, N5130);
nand NAND4 (N5135, N5125, N4584, N107, N4512);
buf BUF1 (N5136, N5134);
xor XOR2 (N5137, N5131, N5);
xor XOR2 (N5138, N5133, N1918);
buf BUF1 (N5139, N5137);
nor NOR2 (N5140, N5135, N2172);
and AND2 (N5141, N5097, N4324);
nand NAND3 (N5142, N5127, N1353, N4657);
or OR3 (N5143, N5120, N537, N2690);
not NOT1 (N5144, N5138);
buf BUF1 (N5145, N5124);
and AND3 (N5146, N5140, N1812, N4667);
or OR2 (N5147, N5146, N2345);
or OR3 (N5148, N5144, N1553, N1649);
and AND4 (N5149, N5136, N3806, N3716, N1244);
or OR4 (N5150, N5148, N3407, N3715, N373);
not NOT1 (N5151, N5150);
and AND2 (N5152, N5142, N2831);
or OR2 (N5153, N5152, N4014);
nor NOR3 (N5154, N5147, N2537, N1786);
not NOT1 (N5155, N5139);
and AND2 (N5156, N5151, N3348);
buf BUF1 (N5157, N5145);
and AND4 (N5158, N5153, N3099, N3438, N4470);
not NOT1 (N5159, N5141);
nand NAND3 (N5160, N5157, N2392, N4461);
or OR3 (N5161, N5132, N1471, N5156);
or OR2 (N5162, N1994, N2146);
nand NAND2 (N5163, N5160, N3407);
buf BUF1 (N5164, N5159);
and AND2 (N5165, N5149, N3949);
not NOT1 (N5166, N5154);
buf BUF1 (N5167, N5143);
buf BUF1 (N5168, N5165);
nand NAND4 (N5169, N5167, N36, N1021, N430);
and AND2 (N5170, N5169, N677);
not NOT1 (N5171, N5170);
xor XOR2 (N5172, N5158, N974);
and AND4 (N5173, N5172, N2975, N3374, N2304);
or OR2 (N5174, N5171, N5068);
nor NOR4 (N5175, N5162, N2059, N2124, N3152);
nand NAND3 (N5176, N5161, N4318, N4004);
nand NAND2 (N5177, N5174, N1272);
not NOT1 (N5178, N5164);
xor XOR2 (N5179, N5155, N3269);
not NOT1 (N5180, N5178);
not NOT1 (N5181, N5129);
or OR2 (N5182, N5180, N720);
or OR4 (N5183, N5176, N4512, N914, N117);
nand NAND4 (N5184, N5166, N1659, N3606, N3879);
xor XOR2 (N5185, N5181, N469);
or OR4 (N5186, N5179, N3328, N4222, N3165);
and AND3 (N5187, N5173, N566, N3370);
not NOT1 (N5188, N5183);
not NOT1 (N5189, N5163);
nor NOR3 (N5190, N5177, N2728, N4566);
buf BUF1 (N5191, N5185);
nand NAND2 (N5192, N5175, N1579);
nor NOR4 (N5193, N5188, N3729, N2335, N4721);
and AND4 (N5194, N5191, N4392, N1559, N4161);
and AND4 (N5195, N5190, N1292, N2067, N1102);
nand NAND4 (N5196, N5194, N4077, N555, N4050);
xor XOR2 (N5197, N5186, N324);
and AND4 (N5198, N5193, N5149, N3374, N291);
xor XOR2 (N5199, N5189, N1648);
or OR3 (N5200, N5182, N2458, N4465);
and AND2 (N5201, N5187, N2915);
or OR2 (N5202, N5168, N80);
or OR3 (N5203, N5201, N872, N718);
xor XOR2 (N5204, N5192, N929);
and AND2 (N5205, N5195, N3804);
nor NOR2 (N5206, N5202, N2615);
buf BUF1 (N5207, N5206);
and AND4 (N5208, N5200, N893, N881, N1932);
not NOT1 (N5209, N5207);
and AND3 (N5210, N5209, N2707, N26);
xor XOR2 (N5211, N5197, N4574);
or OR4 (N5212, N5205, N4306, N826, N2551);
nand NAND4 (N5213, N5196, N3298, N3817, N1548);
nor NOR3 (N5214, N5213, N1446, N5139);
not NOT1 (N5215, N5214);
nor NOR4 (N5216, N5204, N3354, N2454, N458);
buf BUF1 (N5217, N5215);
nand NAND4 (N5218, N5198, N922, N1348, N1930);
nand NAND2 (N5219, N5212, N3763);
and AND4 (N5220, N5184, N4891, N4320, N1098);
xor XOR2 (N5221, N5216, N2400);
or OR3 (N5222, N5208, N809, N3189);
nor NOR3 (N5223, N5210, N336, N3402);
not NOT1 (N5224, N5219);
nand NAND3 (N5225, N5222, N3252, N87);
nor NOR4 (N5226, N5223, N7, N249, N1973);
and AND3 (N5227, N5218, N738, N4963);
and AND3 (N5228, N5225, N3718, N1321);
xor XOR2 (N5229, N5228, N1111);
not NOT1 (N5230, N5211);
buf BUF1 (N5231, N5221);
not NOT1 (N5232, N5203);
or OR2 (N5233, N5231, N513);
and AND4 (N5234, N5220, N2301, N1377, N918);
nand NAND3 (N5235, N5232, N2507, N2074);
xor XOR2 (N5236, N5227, N646);
nor NOR3 (N5237, N5233, N4358, N3856);
nor NOR2 (N5238, N5235, N3744);
not NOT1 (N5239, N5217);
buf BUF1 (N5240, N5226);
buf BUF1 (N5241, N5229);
or OR4 (N5242, N5240, N146, N873, N4280);
nand NAND3 (N5243, N5239, N296, N5175);
xor XOR2 (N5244, N5238, N1079);
buf BUF1 (N5245, N5236);
nand NAND2 (N5246, N5241, N2522);
not NOT1 (N5247, N5230);
buf BUF1 (N5248, N5244);
not NOT1 (N5249, N5247);
buf BUF1 (N5250, N5248);
not NOT1 (N5251, N5234);
and AND4 (N5252, N5243, N288, N3673, N5234);
nand NAND2 (N5253, N5252, N2080);
and AND4 (N5254, N5249, N4737, N2016, N784);
nor NOR2 (N5255, N5253, N502);
nand NAND4 (N5256, N5255, N3301, N1738, N3216);
nand NAND4 (N5257, N5254, N2296, N2968, N263);
xor XOR2 (N5258, N5199, N3617);
or OR4 (N5259, N5237, N5009, N65, N911);
nand NAND4 (N5260, N5256, N5031, N3200, N1636);
not NOT1 (N5261, N5224);
buf BUF1 (N5262, N5258);
nor NOR3 (N5263, N5242, N1190, N5045);
or OR2 (N5264, N5250, N4610);
and AND4 (N5265, N5257, N3182, N1517, N4509);
buf BUF1 (N5266, N5265);
nor NOR3 (N5267, N5260, N2044, N4535);
not NOT1 (N5268, N5262);
buf BUF1 (N5269, N5261);
or OR2 (N5270, N5266, N436);
nor NOR2 (N5271, N5245, N3103);
not NOT1 (N5272, N5264);
nand NAND3 (N5273, N5268, N3636, N4276);
buf BUF1 (N5274, N5271);
and AND4 (N5275, N5267, N4254, N955, N2403);
not NOT1 (N5276, N5246);
buf BUF1 (N5277, N5272);
nor NOR4 (N5278, N5275, N517, N852, N3113);
or OR2 (N5279, N5269, N3481);
xor XOR2 (N5280, N5259, N1820);
nor NOR4 (N5281, N5276, N1895, N3082, N1552);
xor XOR2 (N5282, N5280, N3943);
xor XOR2 (N5283, N5279, N1583);
not NOT1 (N5284, N5282);
and AND2 (N5285, N5284, N2280);
not NOT1 (N5286, N5251);
nand NAND4 (N5287, N5273, N5012, N4770, N2943);
buf BUF1 (N5288, N5286);
buf BUF1 (N5289, N5285);
and AND4 (N5290, N5263, N3038, N3367, N5096);
buf BUF1 (N5291, N5289);
xor XOR2 (N5292, N5281, N1406);
not NOT1 (N5293, N5290);
not NOT1 (N5294, N5277);
xor XOR2 (N5295, N5283, N4340);
nand NAND4 (N5296, N5293, N1727, N3089, N2215);
nor NOR4 (N5297, N5296, N2289, N1919, N487);
buf BUF1 (N5298, N5287);
nor NOR2 (N5299, N5291, N4472);
nor NOR4 (N5300, N5298, N1854, N1026, N407);
buf BUF1 (N5301, N5299);
nor NOR2 (N5302, N5278, N2159);
nand NAND2 (N5303, N5301, N1156);
nand NAND4 (N5304, N5288, N990, N2267, N4045);
not NOT1 (N5305, N5300);
not NOT1 (N5306, N5295);
and AND2 (N5307, N5305, N3774);
nor NOR2 (N5308, N5297, N322);
xor XOR2 (N5309, N5303, N3113);
or OR3 (N5310, N5274, N2230, N2129);
buf BUF1 (N5311, N5308);
buf BUF1 (N5312, N5304);
and AND2 (N5313, N5294, N694);
or OR3 (N5314, N5307, N1304, N4714);
not NOT1 (N5315, N5313);
or OR2 (N5316, N5302, N2574);
and AND4 (N5317, N5314, N405, N658, N4870);
buf BUF1 (N5318, N5311);
and AND4 (N5319, N5312, N4100, N323, N2402);
buf BUF1 (N5320, N5310);
nand NAND3 (N5321, N5320, N5265, N3879);
nor NOR2 (N5322, N5306, N3253);
nand NAND4 (N5323, N5270, N2, N4039, N4942);
nor NOR3 (N5324, N5321, N562, N5054);
xor XOR2 (N5325, N5316, N4396);
nor NOR4 (N5326, N5292, N258, N2113, N2836);
or OR2 (N5327, N5315, N3926);
or OR4 (N5328, N5319, N924, N1274, N5079);
nand NAND2 (N5329, N5327, N3907);
nand NAND3 (N5330, N5329, N207, N2307);
buf BUF1 (N5331, N5325);
and AND3 (N5332, N5328, N5165, N173);
nor NOR2 (N5333, N5309, N2065);
or OR3 (N5334, N5318, N292, N127);
nor NOR2 (N5335, N5330, N3874);
not NOT1 (N5336, N5333);
buf BUF1 (N5337, N5326);
not NOT1 (N5338, N5334);
nor NOR4 (N5339, N5336, N1656, N3927, N1119);
nand NAND2 (N5340, N5339, N4914);
xor XOR2 (N5341, N5324, N2369);
and AND2 (N5342, N5338, N3767);
or OR2 (N5343, N5340, N813);
buf BUF1 (N5344, N5323);
not NOT1 (N5345, N5344);
buf BUF1 (N5346, N5331);
not NOT1 (N5347, N5341);
nor NOR2 (N5348, N5343, N2432);
nor NOR3 (N5349, N5322, N4252, N1657);
not NOT1 (N5350, N5345);
xor XOR2 (N5351, N5332, N411);
nand NAND3 (N5352, N5347, N3484, N3317);
not NOT1 (N5353, N5349);
and AND2 (N5354, N5351, N3532);
xor XOR2 (N5355, N5346, N4471);
not NOT1 (N5356, N5348);
xor XOR2 (N5357, N5337, N1536);
nand NAND3 (N5358, N5357, N4843, N990);
or OR4 (N5359, N5355, N634, N4636, N2902);
or OR3 (N5360, N5359, N552, N2702);
not NOT1 (N5361, N5335);
and AND2 (N5362, N5350, N583);
and AND2 (N5363, N5358, N1348);
and AND2 (N5364, N5353, N2284);
and AND4 (N5365, N5360, N236, N5046, N4164);
not NOT1 (N5366, N5365);
and AND3 (N5367, N5363, N3285, N1991);
not NOT1 (N5368, N5362);
xor XOR2 (N5369, N5352, N3139);
buf BUF1 (N5370, N5368);
buf BUF1 (N5371, N5366);
nand NAND4 (N5372, N5361, N1818, N4841, N3595);
nand NAND2 (N5373, N5354, N2676);
xor XOR2 (N5374, N5370, N5154);
nand NAND4 (N5375, N5356, N3452, N3073, N119);
or OR2 (N5376, N5317, N3132);
not NOT1 (N5377, N5375);
or OR3 (N5378, N5364, N1256, N1867);
or OR2 (N5379, N5369, N470);
nor NOR2 (N5380, N5342, N5034);
nand NAND3 (N5381, N5377, N5149, N1603);
not NOT1 (N5382, N5374);
buf BUF1 (N5383, N5376);
xor XOR2 (N5384, N5383, N1308);
xor XOR2 (N5385, N5371, N2416);
or OR3 (N5386, N5385, N3567, N4445);
nor NOR2 (N5387, N5367, N4293);
not NOT1 (N5388, N5387);
buf BUF1 (N5389, N5372);
xor XOR2 (N5390, N5378, N3083);
not NOT1 (N5391, N5384);
nor NOR3 (N5392, N5390, N5244, N3188);
or OR2 (N5393, N5379, N1783);
and AND3 (N5394, N5381, N987, N3862);
xor XOR2 (N5395, N5391, N920);
and AND4 (N5396, N5380, N4296, N1035, N5244);
and AND3 (N5397, N5386, N2897, N5137);
nand NAND3 (N5398, N5373, N2119, N3056);
not NOT1 (N5399, N5392);
nor NOR2 (N5400, N5389, N3550);
not NOT1 (N5401, N5399);
not NOT1 (N5402, N5396);
nand NAND2 (N5403, N5382, N1920);
buf BUF1 (N5404, N5400);
xor XOR2 (N5405, N5393, N4192);
nor NOR2 (N5406, N5403, N3002);
not NOT1 (N5407, N5406);
nor NOR3 (N5408, N5398, N498, N570);
buf BUF1 (N5409, N5402);
buf BUF1 (N5410, N5405);
or OR2 (N5411, N5410, N4169);
xor XOR2 (N5412, N5407, N4273);
or OR2 (N5413, N5404, N2390);
and AND2 (N5414, N5388, N3033);
not NOT1 (N5415, N5412);
nor NOR3 (N5416, N5409, N4321, N3984);
and AND3 (N5417, N5397, N4565, N424);
nor NOR4 (N5418, N5394, N122, N4329, N3295);
not NOT1 (N5419, N5413);
nor NOR3 (N5420, N5419, N4769, N3630);
or OR2 (N5421, N5415, N481);
not NOT1 (N5422, N5416);
nor NOR2 (N5423, N5420, N2240);
buf BUF1 (N5424, N5418);
xor XOR2 (N5425, N5424, N646);
not NOT1 (N5426, N5401);
nand NAND4 (N5427, N5417, N3314, N3281, N889);
not NOT1 (N5428, N5422);
buf BUF1 (N5429, N5414);
buf BUF1 (N5430, N5427);
xor XOR2 (N5431, N5411, N4896);
and AND4 (N5432, N5423, N4146, N2067, N2028);
not NOT1 (N5433, N5430);
and AND2 (N5434, N5395, N4827);
nand NAND4 (N5435, N5425, N2209, N565, N3717);
and AND4 (N5436, N5431, N1220, N1931, N1545);
buf BUF1 (N5437, N5432);
not NOT1 (N5438, N5421);
xor XOR2 (N5439, N5426, N2747);
nand NAND4 (N5440, N5435, N3178, N4463, N1304);
nor NOR2 (N5441, N5437, N5050);
nand NAND3 (N5442, N5441, N4333, N1219);
not NOT1 (N5443, N5408);
not NOT1 (N5444, N5429);
nor NOR3 (N5445, N5440, N409, N809);
not NOT1 (N5446, N5444);
nand NAND3 (N5447, N5443, N3656, N1439);
and AND2 (N5448, N5436, N2868);
xor XOR2 (N5449, N5445, N3592);
xor XOR2 (N5450, N5442, N1757);
buf BUF1 (N5451, N5447);
xor XOR2 (N5452, N5433, N449);
and AND2 (N5453, N5446, N3129);
nand NAND4 (N5454, N5439, N1004, N4557, N5356);
or OR4 (N5455, N5452, N4484, N3978, N3450);
nor NOR2 (N5456, N5438, N4042);
buf BUF1 (N5457, N5455);
or OR2 (N5458, N5451, N3546);
xor XOR2 (N5459, N5456, N4063);
buf BUF1 (N5460, N5454);
buf BUF1 (N5461, N5428);
xor XOR2 (N5462, N5449, N2475);
nor NOR4 (N5463, N5448, N351, N649, N4766);
or OR2 (N5464, N5453, N2443);
and AND3 (N5465, N5457, N296, N3942);
and AND3 (N5466, N5458, N5410, N4572);
and AND4 (N5467, N5459, N207, N517, N2938);
buf BUF1 (N5468, N5463);
nand NAND4 (N5469, N5434, N2819, N51, N3486);
xor XOR2 (N5470, N5460, N1924);
xor XOR2 (N5471, N5464, N2243);
or OR4 (N5472, N5462, N641, N985, N2035);
nor NOR3 (N5473, N5466, N585, N3863);
nand NAND2 (N5474, N5471, N1036);
or OR4 (N5475, N5465, N4119, N4380, N5266);
buf BUF1 (N5476, N5469);
not NOT1 (N5477, N5475);
and AND2 (N5478, N5450, N4386);
not NOT1 (N5479, N5477);
nand NAND2 (N5480, N5472, N2785);
nor NOR4 (N5481, N5468, N2120, N4484, N1725);
buf BUF1 (N5482, N5474);
xor XOR2 (N5483, N5482, N2651);
not NOT1 (N5484, N5479);
or OR4 (N5485, N5476, N2676, N5353, N2167);
not NOT1 (N5486, N5485);
nand NAND2 (N5487, N5483, N107);
xor XOR2 (N5488, N5487, N86);
and AND3 (N5489, N5480, N3372, N1834);
not NOT1 (N5490, N5489);
or OR2 (N5491, N5490, N234);
nor NOR3 (N5492, N5484, N5447, N3991);
xor XOR2 (N5493, N5478, N1742);
buf BUF1 (N5494, N5493);
not NOT1 (N5495, N5488);
nand NAND2 (N5496, N5481, N2525);
and AND3 (N5497, N5486, N5439, N3944);
nand NAND4 (N5498, N5491, N4944, N4047, N4445);
buf BUF1 (N5499, N5470);
nor NOR2 (N5500, N5497, N5462);
not NOT1 (N5501, N5461);
nor NOR2 (N5502, N5495, N4238);
xor XOR2 (N5503, N5494, N4259);
nor NOR4 (N5504, N5499, N5446, N4714, N4266);
nand NAND3 (N5505, N5500, N4587, N705);
nand NAND3 (N5506, N5502, N4171, N1840);
buf BUF1 (N5507, N5506);
xor XOR2 (N5508, N5473, N1728);
buf BUF1 (N5509, N5492);
or OR2 (N5510, N5496, N1267);
not NOT1 (N5511, N5504);
nand NAND4 (N5512, N5505, N4282, N74, N951);
and AND3 (N5513, N5508, N380, N1335);
and AND2 (N5514, N5509, N170);
not NOT1 (N5515, N5467);
not NOT1 (N5516, N5514);
nor NOR2 (N5517, N5498, N3684);
nand NAND2 (N5518, N5503, N1222);
buf BUF1 (N5519, N5518);
xor XOR2 (N5520, N5513, N792);
or OR2 (N5521, N5516, N3920);
xor XOR2 (N5522, N5519, N4625);
buf BUF1 (N5523, N5511);
or OR4 (N5524, N5501, N314, N1342, N1000);
nor NOR2 (N5525, N5523, N3840);
and AND2 (N5526, N5525, N3931);
xor XOR2 (N5527, N5520, N3737);
and AND4 (N5528, N5515, N3961, N2922, N1686);
nor NOR2 (N5529, N5528, N3717);
nor NOR4 (N5530, N5524, N4052, N1714, N4880);
xor XOR2 (N5531, N5530, N746);
nand NAND4 (N5532, N5527, N3729, N3060, N155);
xor XOR2 (N5533, N5517, N3402);
nand NAND4 (N5534, N5526, N1216, N4017, N4210);
buf BUF1 (N5535, N5529);
or OR2 (N5536, N5522, N5121);
not NOT1 (N5537, N5521);
nand NAND2 (N5538, N5532, N3217);
buf BUF1 (N5539, N5531);
nor NOR4 (N5540, N5512, N5158, N2905, N8);
not NOT1 (N5541, N5534);
and AND4 (N5542, N5537, N4146, N4864, N3633);
and AND3 (N5543, N5541, N2961, N4384);
not NOT1 (N5544, N5533);
and AND3 (N5545, N5544, N601, N2467);
nand NAND4 (N5546, N5536, N3131, N4106, N4977);
nor NOR4 (N5547, N5535, N4766, N3983, N5029);
nand NAND2 (N5548, N5538, N2581);
buf BUF1 (N5549, N5510);
and AND2 (N5550, N5545, N3677);
or OR4 (N5551, N5540, N719, N2296, N5351);
nand NAND4 (N5552, N5546, N5022, N3880, N3575);
nor NOR4 (N5553, N5548, N3175, N2838, N2082);
not NOT1 (N5554, N5539);
or OR2 (N5555, N5547, N1605);
and AND3 (N5556, N5549, N3088, N3245);
xor XOR2 (N5557, N5542, N1892);
not NOT1 (N5558, N5556);
or OR4 (N5559, N5551, N339, N771, N471);
xor XOR2 (N5560, N5553, N1157);
or OR2 (N5561, N5559, N3847);
nand NAND2 (N5562, N5507, N5161);
buf BUF1 (N5563, N5561);
and AND2 (N5564, N5560, N1058);
nand NAND2 (N5565, N5558, N66);
and AND2 (N5566, N5552, N97);
buf BUF1 (N5567, N5554);
or OR4 (N5568, N5565, N2912, N5406, N968);
nor NOR2 (N5569, N5557, N1986);
nand NAND2 (N5570, N5564, N2223);
nand NAND3 (N5571, N5555, N1250, N5252);
buf BUF1 (N5572, N5562);
and AND4 (N5573, N5572, N1437, N602, N4904);
nand NAND2 (N5574, N5571, N2054);
nand NAND3 (N5575, N5550, N1602, N3705);
not NOT1 (N5576, N5574);
nand NAND4 (N5577, N5568, N1864, N4012, N3525);
buf BUF1 (N5578, N5543);
nand NAND2 (N5579, N5576, N3153);
buf BUF1 (N5580, N5566);
buf BUF1 (N5581, N5579);
and AND2 (N5582, N5567, N2527);
buf BUF1 (N5583, N5569);
not NOT1 (N5584, N5581);
or OR4 (N5585, N5575, N5356, N4324, N3282);
nand NAND2 (N5586, N5585, N2968);
nand NAND2 (N5587, N5584, N4998);
or OR3 (N5588, N5586, N2974, N2659);
buf BUF1 (N5589, N5580);
and AND2 (N5590, N5563, N4994);
buf BUF1 (N5591, N5577);
and AND4 (N5592, N5582, N2640, N4940, N1620);
buf BUF1 (N5593, N5570);
xor XOR2 (N5594, N5591, N1914);
and AND2 (N5595, N5593, N1579);
not NOT1 (N5596, N5595);
and AND2 (N5597, N5590, N1989);
xor XOR2 (N5598, N5588, N3420);
and AND3 (N5599, N5596, N2686, N4837);
and AND4 (N5600, N5599, N3049, N1119, N4883);
and AND2 (N5601, N5573, N5548);
or OR2 (N5602, N5578, N1840);
xor XOR2 (N5603, N5600, N3282);
not NOT1 (N5604, N5589);
xor XOR2 (N5605, N5603, N2791);
nor NOR4 (N5606, N5597, N4133, N1858, N4556);
or OR4 (N5607, N5606, N5159, N5122, N3830);
nand NAND4 (N5608, N5604, N1597, N5386, N2499);
xor XOR2 (N5609, N5587, N5454);
nand NAND3 (N5610, N5601, N401, N3241);
and AND2 (N5611, N5609, N4321);
not NOT1 (N5612, N5608);
nor NOR2 (N5613, N5583, N5337);
nand NAND4 (N5614, N5592, N4653, N1397, N4204);
nand NAND3 (N5615, N5605, N5611, N2605);
buf BUF1 (N5616, N318);
or OR4 (N5617, N5614, N2788, N1521, N1139);
nor NOR3 (N5618, N5613, N1579, N3491);
not NOT1 (N5619, N5607);
buf BUF1 (N5620, N5598);
and AND4 (N5621, N5619, N2195, N4512, N3741);
xor XOR2 (N5622, N5620, N1382);
or OR2 (N5623, N5615, N4159);
nor NOR3 (N5624, N5594, N4560, N4301);
or OR3 (N5625, N5622, N2270, N25);
xor XOR2 (N5626, N5624, N1285);
not NOT1 (N5627, N5610);
not NOT1 (N5628, N5612);
or OR3 (N5629, N5616, N2920, N2391);
and AND4 (N5630, N5602, N267, N1387, N469);
buf BUF1 (N5631, N5626);
xor XOR2 (N5632, N5623, N2438);
nand NAND3 (N5633, N5630, N1205, N802);
nor NOR4 (N5634, N5631, N5267, N3220, N1205);
nor NOR3 (N5635, N5632, N3309, N5071);
nor NOR2 (N5636, N5629, N810);
buf BUF1 (N5637, N5618);
buf BUF1 (N5638, N5636);
xor XOR2 (N5639, N5634, N1157);
xor XOR2 (N5640, N5625, N3225);
xor XOR2 (N5641, N5633, N3487);
not NOT1 (N5642, N5617);
buf BUF1 (N5643, N5637);
and AND2 (N5644, N5643, N4743);
buf BUF1 (N5645, N5635);
and AND3 (N5646, N5621, N2161, N4046);
or OR2 (N5647, N5627, N3075);
nand NAND4 (N5648, N5647, N2398, N5045, N2177);
nor NOR3 (N5649, N5641, N3650, N5390);
and AND3 (N5650, N5648, N4110, N285);
xor XOR2 (N5651, N5638, N5602);
nor NOR3 (N5652, N5640, N1065, N2753);
nor NOR2 (N5653, N5650, N5430);
nor NOR2 (N5654, N5639, N5293);
nand NAND4 (N5655, N5652, N3593, N5068, N2729);
not NOT1 (N5656, N5628);
not NOT1 (N5657, N5645);
xor XOR2 (N5658, N5649, N970);
not NOT1 (N5659, N5653);
or OR3 (N5660, N5644, N1037, N5190);
not NOT1 (N5661, N5655);
nand NAND4 (N5662, N5661, N4223, N3732, N736);
nand NAND2 (N5663, N5646, N4636);
nand NAND2 (N5664, N5642, N3639);
or OR2 (N5665, N5654, N3316);
or OR3 (N5666, N5665, N4122, N2059);
nand NAND3 (N5667, N5651, N822, N5326);
or OR3 (N5668, N5667, N2963, N3794);
and AND4 (N5669, N5657, N2420, N4873, N1522);
or OR2 (N5670, N5660, N2306);
nand NAND2 (N5671, N5658, N4996);
buf BUF1 (N5672, N5662);
buf BUF1 (N5673, N5670);
buf BUF1 (N5674, N5664);
nor NOR3 (N5675, N5656, N3113, N909);
xor XOR2 (N5676, N5663, N793);
not NOT1 (N5677, N5668);
xor XOR2 (N5678, N5666, N4824);
not NOT1 (N5679, N5659);
nor NOR3 (N5680, N5678, N1278, N4283);
nor NOR2 (N5681, N5676, N5005);
xor XOR2 (N5682, N5672, N3224);
buf BUF1 (N5683, N5673);
xor XOR2 (N5684, N5669, N1025);
nand NAND2 (N5685, N5683, N2979);
xor XOR2 (N5686, N5685, N3671);
and AND2 (N5687, N5674, N2785);
nand NAND3 (N5688, N5681, N4236, N2749);
or OR4 (N5689, N5677, N4165, N3198, N572);
and AND3 (N5690, N5675, N3464, N30);
buf BUF1 (N5691, N5671);
nor NOR3 (N5692, N5684, N459, N2474);
buf BUF1 (N5693, N5686);
and AND4 (N5694, N5679, N3662, N2764, N1275);
nand NAND4 (N5695, N5682, N5196, N765, N876);
buf BUF1 (N5696, N5688);
or OR3 (N5697, N5689, N3289, N4888);
or OR2 (N5698, N5696, N4392);
buf BUF1 (N5699, N5690);
buf BUF1 (N5700, N5687);
xor XOR2 (N5701, N5693, N4789);
nor NOR2 (N5702, N5680, N521);
xor XOR2 (N5703, N5695, N3036);
not NOT1 (N5704, N5698);
buf BUF1 (N5705, N5701);
nor NOR3 (N5706, N5702, N3213, N2317);
nor NOR3 (N5707, N5692, N1946, N43);
and AND2 (N5708, N5706, N2443);
not NOT1 (N5709, N5707);
buf BUF1 (N5710, N5708);
not NOT1 (N5711, N5700);
and AND3 (N5712, N5711, N5423, N4422);
not NOT1 (N5713, N5709);
and AND2 (N5714, N5705, N4233);
nor NOR2 (N5715, N5691, N2666);
and AND2 (N5716, N5699, N2899);
nand NAND4 (N5717, N5713, N289, N4957, N3172);
and AND3 (N5718, N5694, N4158, N4532);
buf BUF1 (N5719, N5703);
not NOT1 (N5720, N5714);
and AND2 (N5721, N5720, N1339);
nand NAND3 (N5722, N5697, N1792, N2391);
not NOT1 (N5723, N5718);
not NOT1 (N5724, N5712);
xor XOR2 (N5725, N5721, N221);
and AND2 (N5726, N5704, N528);
and AND2 (N5727, N5724, N5335);
not NOT1 (N5728, N5722);
and AND4 (N5729, N5717, N1528, N3049, N2965);
or OR4 (N5730, N5715, N1080, N1641, N3686);
and AND3 (N5731, N5725, N4382, N2155);
not NOT1 (N5732, N5719);
buf BUF1 (N5733, N5710);
buf BUF1 (N5734, N5729);
buf BUF1 (N5735, N5734);
nand NAND2 (N5736, N5716, N4977);
buf BUF1 (N5737, N5726);
nor NOR2 (N5738, N5730, N5061);
buf BUF1 (N5739, N5735);
not NOT1 (N5740, N5739);
nor NOR3 (N5741, N5736, N1082, N4648);
buf BUF1 (N5742, N5733);
or OR2 (N5743, N5732, N4405);
nand NAND2 (N5744, N5742, N1520);
nand NAND2 (N5745, N5740, N5699);
buf BUF1 (N5746, N5737);
nor NOR4 (N5747, N5743, N1799, N4485, N3843);
xor XOR2 (N5748, N5746, N2460);
or OR2 (N5749, N5728, N2755);
nand NAND3 (N5750, N5749, N784, N2399);
nand NAND2 (N5751, N5723, N2965);
or OR3 (N5752, N5748, N5621, N3765);
or OR3 (N5753, N5731, N1001, N4674);
not NOT1 (N5754, N5727);
or OR4 (N5755, N5753, N4218, N4049, N3424);
not NOT1 (N5756, N5744);
nor NOR2 (N5757, N5754, N5249);
nor NOR4 (N5758, N5755, N3274, N5348, N1827);
xor XOR2 (N5759, N5747, N3830);
and AND4 (N5760, N5759, N1234, N5169, N1209);
or OR4 (N5761, N5750, N3433, N2838, N924);
nor NOR2 (N5762, N5756, N342);
xor XOR2 (N5763, N5758, N2395);
buf BUF1 (N5764, N5752);
buf BUF1 (N5765, N5757);
and AND2 (N5766, N5751, N2904);
buf BUF1 (N5767, N5745);
xor XOR2 (N5768, N5741, N4052);
buf BUF1 (N5769, N5766);
or OR3 (N5770, N5764, N3962, N947);
not NOT1 (N5771, N5763);
and AND3 (N5772, N5771, N2254, N934);
nor NOR3 (N5773, N5767, N3301, N1654);
xor XOR2 (N5774, N5762, N2665);
not NOT1 (N5775, N5774);
or OR3 (N5776, N5765, N2295, N2056);
xor XOR2 (N5777, N5770, N3282);
buf BUF1 (N5778, N5777);
or OR2 (N5779, N5768, N4608);
not NOT1 (N5780, N5761);
nor NOR4 (N5781, N5769, N5177, N295, N4404);
not NOT1 (N5782, N5781);
or OR3 (N5783, N5779, N594, N3860);
not NOT1 (N5784, N5775);
xor XOR2 (N5785, N5780, N3779);
nor NOR2 (N5786, N5778, N3190);
not NOT1 (N5787, N5784);
not NOT1 (N5788, N5738);
not NOT1 (N5789, N5782);
not NOT1 (N5790, N5760);
not NOT1 (N5791, N5788);
not NOT1 (N5792, N5772);
nand NAND2 (N5793, N5789, N4914);
and AND4 (N5794, N5785, N5737, N2622, N820);
xor XOR2 (N5795, N5793, N2089);
nand NAND3 (N5796, N5790, N4823, N2380);
not NOT1 (N5797, N5795);
nand NAND3 (N5798, N5792, N2331, N4866);
and AND4 (N5799, N5796, N2224, N4042, N1252);
not NOT1 (N5800, N5798);
and AND4 (N5801, N5787, N131, N1690, N220);
or OR3 (N5802, N5776, N3567, N5472);
nand NAND4 (N5803, N5801, N2360, N3340, N3796);
xor XOR2 (N5804, N5791, N1548);
and AND3 (N5805, N5794, N3005, N4293);
nand NAND3 (N5806, N5797, N5791, N3000);
xor XOR2 (N5807, N5800, N4492);
buf BUF1 (N5808, N5805);
and AND4 (N5809, N5773, N3245, N4588, N4189);
not NOT1 (N5810, N5786);
and AND2 (N5811, N5799, N499);
not NOT1 (N5812, N5808);
nand NAND2 (N5813, N5812, N528);
or OR2 (N5814, N5804, N5129);
or OR4 (N5815, N5814, N3227, N4798, N5568);
nor NOR3 (N5816, N5807, N4398, N544);
or OR3 (N5817, N5783, N3975, N2949);
buf BUF1 (N5818, N5802);
or OR4 (N5819, N5811, N3030, N750, N5000);
xor XOR2 (N5820, N5816, N5435);
nor NOR3 (N5821, N5803, N1038, N5690);
nand NAND3 (N5822, N5820, N108, N615);
buf BUF1 (N5823, N5821);
or OR4 (N5824, N5822, N240, N4195, N3004);
xor XOR2 (N5825, N5815, N2604);
not NOT1 (N5826, N5806);
nand NAND3 (N5827, N5809, N1980, N4386);
xor XOR2 (N5828, N5827, N1781);
not NOT1 (N5829, N5818);
or OR2 (N5830, N5823, N4337);
nand NAND4 (N5831, N5813, N2520, N745, N298);
nor NOR3 (N5832, N5829, N507, N504);
xor XOR2 (N5833, N5817, N2020);
nor NOR4 (N5834, N5828, N991, N609, N3921);
nand NAND3 (N5835, N5832, N1021, N3071);
buf BUF1 (N5836, N5833);
nand NAND4 (N5837, N5826, N2772, N3314, N1024);
and AND4 (N5838, N5825, N1735, N5293, N4647);
nor NOR2 (N5839, N5819, N2262);
or OR3 (N5840, N5836, N283, N3290);
and AND3 (N5841, N5837, N1656, N3997);
xor XOR2 (N5842, N5835, N4295);
nand NAND2 (N5843, N5838, N215);
or OR3 (N5844, N5830, N3042, N3272);
buf BUF1 (N5845, N5834);
and AND2 (N5846, N5840, N2873);
nor NOR4 (N5847, N5844, N3894, N897, N1416);
nand NAND2 (N5848, N5810, N5148);
nand NAND3 (N5849, N5824, N857, N2720);
or OR4 (N5850, N5842, N4349, N167, N821);
buf BUF1 (N5851, N5849);
not NOT1 (N5852, N5850);
and AND2 (N5853, N5843, N4188);
xor XOR2 (N5854, N5839, N4656);
xor XOR2 (N5855, N5847, N1592);
and AND3 (N5856, N5854, N5730, N4528);
or OR3 (N5857, N5845, N512, N3985);
nor NOR2 (N5858, N5848, N472);
not NOT1 (N5859, N5856);
nor NOR4 (N5860, N5855, N4992, N4172, N1773);
nor NOR2 (N5861, N5860, N1667);
buf BUF1 (N5862, N5859);
nor NOR4 (N5863, N5846, N5746, N4238, N1368);
nor NOR4 (N5864, N5861, N5669, N4581, N1218);
buf BUF1 (N5865, N5853);
nand NAND2 (N5866, N5862, N2427);
buf BUF1 (N5867, N5866);
and AND3 (N5868, N5865, N1321, N5853);
and AND2 (N5869, N5867, N5773);
xor XOR2 (N5870, N5868, N1544);
and AND2 (N5871, N5870, N1803);
or OR3 (N5872, N5857, N2405, N953);
nor NOR3 (N5873, N5864, N969, N1869);
nor NOR3 (N5874, N5873, N5849, N2832);
xor XOR2 (N5875, N5851, N4695);
xor XOR2 (N5876, N5831, N2091);
xor XOR2 (N5877, N5874, N2573);
nor NOR4 (N5878, N5872, N5203, N26, N817);
not NOT1 (N5879, N5863);
not NOT1 (N5880, N5841);
not NOT1 (N5881, N5878);
buf BUF1 (N5882, N5871);
nor NOR4 (N5883, N5880, N5213, N292, N3994);
nor NOR3 (N5884, N5882, N2311, N2786);
and AND3 (N5885, N5877, N3658, N77);
nand NAND4 (N5886, N5881, N3671, N833, N4567);
and AND4 (N5887, N5885, N3367, N4936, N5670);
buf BUF1 (N5888, N5869);
nor NOR4 (N5889, N5876, N220, N3260, N705);
and AND4 (N5890, N5852, N3023, N4002, N977);
nor NOR2 (N5891, N5879, N2615);
buf BUF1 (N5892, N5889);
nor NOR2 (N5893, N5884, N1945);
or OR3 (N5894, N5893, N1655, N3178);
and AND3 (N5895, N5883, N4146, N5448);
xor XOR2 (N5896, N5888, N4466);
or OR2 (N5897, N5892, N2054);
nand NAND3 (N5898, N5896, N2344, N4189);
or OR3 (N5899, N5891, N751, N2555);
not NOT1 (N5900, N5895);
xor XOR2 (N5901, N5898, N2809);
and AND4 (N5902, N5886, N3541, N2681, N3305);
xor XOR2 (N5903, N5901, N1949);
or OR3 (N5904, N5903, N5842, N3746);
nand NAND3 (N5905, N5875, N5016, N3154);
buf BUF1 (N5906, N5904);
nand NAND4 (N5907, N5900, N694, N4918, N4292);
nand NAND3 (N5908, N5906, N2460, N443);
and AND2 (N5909, N5899, N1793);
nor NOR2 (N5910, N5905, N387);
not NOT1 (N5911, N5894);
nand NAND3 (N5912, N5902, N2913, N3854);
nand NAND3 (N5913, N5897, N3194, N3090);
nor NOR2 (N5914, N5887, N3172);
buf BUF1 (N5915, N5912);
nor NOR2 (N5916, N5914, N1773);
and AND4 (N5917, N5858, N5465, N2917, N1055);
nor NOR3 (N5918, N5917, N1874, N5188);
not NOT1 (N5919, N5908);
nor NOR4 (N5920, N5918, N759, N5427, N5404);
xor XOR2 (N5921, N5911, N192);
xor XOR2 (N5922, N5890, N883);
not NOT1 (N5923, N5916);
nor NOR2 (N5924, N5913, N2729);
and AND4 (N5925, N5907, N1337, N4078, N4284);
or OR2 (N5926, N5923, N4748);
or OR4 (N5927, N5922, N4683, N2402, N2907);
buf BUF1 (N5928, N5924);
and AND3 (N5929, N5926, N3753, N4174);
and AND3 (N5930, N5929, N5612, N4639);
or OR2 (N5931, N5909, N2758);
not NOT1 (N5932, N5915);
not NOT1 (N5933, N5932);
or OR3 (N5934, N5920, N2034, N862);
xor XOR2 (N5935, N5930, N1271);
and AND4 (N5936, N5919, N2162, N5768, N2996);
nor NOR4 (N5937, N5910, N2860, N3250, N5802);
nor NOR4 (N5938, N5934, N5567, N824, N91);
nor NOR3 (N5939, N5925, N4128, N1388);
and AND4 (N5940, N5931, N4117, N548, N996);
buf BUF1 (N5941, N5927);
nor NOR4 (N5942, N5921, N1562, N5229, N3767);
not NOT1 (N5943, N5940);
and AND2 (N5944, N5939, N662);
nor NOR3 (N5945, N5937, N2623, N3860);
and AND3 (N5946, N5941, N4931, N5477);
or OR2 (N5947, N5938, N262);
buf BUF1 (N5948, N5935);
nor NOR4 (N5949, N5947, N1771, N4602, N4384);
and AND2 (N5950, N5948, N4258);
or OR2 (N5951, N5933, N4643);
xor XOR2 (N5952, N5949, N4954);
or OR3 (N5953, N5950, N5336, N1492);
nor NOR3 (N5954, N5928, N2395, N4269);
buf BUF1 (N5955, N5946);
and AND4 (N5956, N5951, N5563, N5434, N3345);
xor XOR2 (N5957, N5945, N2534);
and AND4 (N5958, N5953, N5586, N820, N1479);
and AND4 (N5959, N5943, N973, N2867, N4903);
and AND3 (N5960, N5955, N3322, N1656);
not NOT1 (N5961, N5959);
nand NAND3 (N5962, N5960, N2655, N5594);
not NOT1 (N5963, N5956);
nor NOR4 (N5964, N5954, N793, N5598, N906);
nand NAND4 (N5965, N5942, N759, N244, N5927);
and AND4 (N5966, N5957, N5746, N2206, N1821);
buf BUF1 (N5967, N5952);
nand NAND2 (N5968, N5944, N1407);
xor XOR2 (N5969, N5968, N3361);
or OR4 (N5970, N5967, N3250, N4970, N2024);
buf BUF1 (N5971, N5963);
not NOT1 (N5972, N5961);
and AND3 (N5973, N5972, N1272, N477);
or OR2 (N5974, N5966, N5493);
nand NAND2 (N5975, N5936, N384);
not NOT1 (N5976, N5974);
nor NOR4 (N5977, N5958, N528, N3780, N5971);
and AND2 (N5978, N1892, N4166);
not NOT1 (N5979, N5975);
or OR2 (N5980, N5970, N2800);
buf BUF1 (N5981, N5962);
nand NAND2 (N5982, N5981, N2044);
buf BUF1 (N5983, N5964);
nor NOR4 (N5984, N5983, N1129, N4354, N3605);
xor XOR2 (N5985, N5976, N976);
xor XOR2 (N5986, N5969, N3502);
nor NOR3 (N5987, N5982, N4248, N3374);
and AND3 (N5988, N5984, N1495, N3362);
not NOT1 (N5989, N5973);
buf BUF1 (N5990, N5989);
not NOT1 (N5991, N5987);
nor NOR3 (N5992, N5978, N2962, N5405);
not NOT1 (N5993, N5965);
and AND4 (N5994, N5992, N1375, N2032, N3400);
buf BUF1 (N5995, N5991);
and AND2 (N5996, N5988, N3013);
buf BUF1 (N5997, N5985);
xor XOR2 (N5998, N5996, N4623);
or OR2 (N5999, N5977, N3309);
nand NAND4 (N6000, N5990, N4055, N178, N5924);
xor XOR2 (N6001, N5998, N4576);
xor XOR2 (N6002, N5979, N2113);
or OR2 (N6003, N6001, N1866);
and AND3 (N6004, N5995, N4507, N2382);
buf BUF1 (N6005, N5994);
or OR3 (N6006, N5986, N359, N4028);
and AND2 (N6007, N5997, N5156);
or OR4 (N6008, N6002, N5013, N47, N424);
not NOT1 (N6009, N6005);
buf BUF1 (N6010, N6003);
nand NAND3 (N6011, N6009, N4193, N3068);
buf BUF1 (N6012, N6011);
nor NOR2 (N6013, N6007, N4879);
nor NOR3 (N6014, N6006, N4605, N668);
xor XOR2 (N6015, N5999, N5237);
and AND2 (N6016, N6008, N2458);
and AND2 (N6017, N6016, N4211);
and AND4 (N6018, N6010, N5028, N3728, N2798);
nor NOR2 (N6019, N6018, N3266);
not NOT1 (N6020, N6012);
and AND3 (N6021, N6000, N1745, N2056);
and AND3 (N6022, N6020, N3101, N5627);
nand NAND3 (N6023, N6015, N945, N749);
and AND3 (N6024, N6021, N580, N3469);
not NOT1 (N6025, N6013);
or OR2 (N6026, N6019, N4322);
nand NAND2 (N6027, N5980, N1758);
buf BUF1 (N6028, N5993);
nor NOR3 (N6029, N6004, N4397, N853);
nand NAND4 (N6030, N6028, N6008, N2997, N5169);
or OR3 (N6031, N6025, N3369, N3867);
xor XOR2 (N6032, N6017, N2835);
and AND2 (N6033, N6031, N351);
nor NOR2 (N6034, N6029, N2627);
or OR3 (N6035, N6027, N1722, N4199);
buf BUF1 (N6036, N6014);
nand NAND4 (N6037, N6033, N709, N1933, N2233);
xor XOR2 (N6038, N6032, N4732);
or OR3 (N6039, N6034, N2268, N1778);
buf BUF1 (N6040, N6039);
and AND3 (N6041, N6036, N1447, N2634);
and AND2 (N6042, N6022, N270);
nor NOR4 (N6043, N6037, N190, N3427, N1164);
and AND4 (N6044, N6030, N4254, N5177, N762);
nand NAND2 (N6045, N6023, N1094);
and AND2 (N6046, N6038, N3880);
and AND3 (N6047, N6026, N4834, N3209);
buf BUF1 (N6048, N6041);
xor XOR2 (N6049, N6046, N5799);
buf BUF1 (N6050, N6047);
nand NAND2 (N6051, N6024, N5676);
nor NOR3 (N6052, N6045, N1169, N5668);
and AND3 (N6053, N6042, N4241, N900);
and AND2 (N6054, N6050, N3841);
and AND3 (N6055, N6052, N3428, N1909);
or OR4 (N6056, N6040, N2723, N2253, N4646);
xor XOR2 (N6057, N6055, N3529);
not NOT1 (N6058, N6043);
or OR2 (N6059, N6056, N3918);
not NOT1 (N6060, N6044);
nand NAND3 (N6061, N6051, N5496, N2486);
xor XOR2 (N6062, N6061, N193);
and AND4 (N6063, N6057, N2837, N2876, N5169);
buf BUF1 (N6064, N6059);
buf BUF1 (N6065, N6062);
not NOT1 (N6066, N6048);
buf BUF1 (N6067, N6054);
or OR3 (N6068, N6060, N1470, N5195);
and AND3 (N6069, N6064, N5791, N1647);
not NOT1 (N6070, N6058);
xor XOR2 (N6071, N6065, N3826);
nor NOR2 (N6072, N6063, N125);
nor NOR2 (N6073, N6070, N3269);
buf BUF1 (N6074, N6073);
nor NOR2 (N6075, N6068, N6040);
nand NAND4 (N6076, N6066, N140, N2746, N3541);
not NOT1 (N6077, N6067);
or OR3 (N6078, N6069, N2624, N4446);
nor NOR4 (N6079, N6035, N2432, N4359, N1312);
buf BUF1 (N6080, N6078);
xor XOR2 (N6081, N6077, N618);
and AND4 (N6082, N6080, N2232, N4087, N4054);
nor NOR4 (N6083, N6079, N2002, N4350, N5888);
xor XOR2 (N6084, N6049, N2600);
not NOT1 (N6085, N6081);
xor XOR2 (N6086, N6084, N1924);
buf BUF1 (N6087, N6085);
xor XOR2 (N6088, N6087, N4284);
or OR2 (N6089, N6086, N4742);
xor XOR2 (N6090, N6083, N4734);
nand NAND3 (N6091, N6089, N2311, N2573);
not NOT1 (N6092, N6082);
xor XOR2 (N6093, N6053, N3230);
not NOT1 (N6094, N6092);
buf BUF1 (N6095, N6076);
buf BUF1 (N6096, N6071);
xor XOR2 (N6097, N6091, N4719);
buf BUF1 (N6098, N6094);
not NOT1 (N6099, N6095);
nand NAND2 (N6100, N6090, N478);
xor XOR2 (N6101, N6100, N2316);
or OR4 (N6102, N6088, N5407, N2746, N4698);
or OR3 (N6103, N6101, N6057, N2806);
or OR2 (N6104, N6103, N2723);
or OR3 (N6105, N6072, N2975, N3535);
and AND2 (N6106, N6097, N1416);
nand NAND2 (N6107, N6075, N5945);
xor XOR2 (N6108, N6106, N4518);
nor NOR4 (N6109, N6093, N362, N4904, N2338);
xor XOR2 (N6110, N6099, N5095);
nor NOR2 (N6111, N6110, N3337);
nand NAND2 (N6112, N6074, N1854);
or OR3 (N6113, N6111, N2836, N4014);
nand NAND2 (N6114, N6098, N388);
or OR4 (N6115, N6113, N1224, N92, N5785);
nor NOR2 (N6116, N6104, N1813);
not NOT1 (N6117, N6096);
xor XOR2 (N6118, N6114, N1206);
or OR4 (N6119, N6109, N5926, N1424, N2487);
buf BUF1 (N6120, N6107);
buf BUF1 (N6121, N6117);
nor NOR3 (N6122, N6120, N5913, N2088);
and AND3 (N6123, N6119, N4298, N161);
or OR4 (N6124, N6115, N3428, N1745, N2114);
nor NOR4 (N6125, N6118, N5902, N4355, N3082);
not NOT1 (N6126, N6122);
buf BUF1 (N6127, N6123);
xor XOR2 (N6128, N6125, N673);
and AND2 (N6129, N6102, N5960);
nand NAND2 (N6130, N6126, N5768);
or OR4 (N6131, N6116, N1545, N978, N661);
buf BUF1 (N6132, N6129);
nand NAND4 (N6133, N6130, N968, N802, N293);
nand NAND2 (N6134, N6133, N6108);
buf BUF1 (N6135, N4699);
or OR4 (N6136, N6132, N5660, N3708, N3078);
or OR4 (N6137, N6124, N2239, N2438, N4378);
and AND4 (N6138, N6127, N5154, N4973, N3025);
buf BUF1 (N6139, N6135);
buf BUF1 (N6140, N6139);
and AND2 (N6141, N6137, N4526);
nor NOR2 (N6142, N6141, N3618);
and AND2 (N6143, N6138, N3659);
not NOT1 (N6144, N6105);
not NOT1 (N6145, N6136);
nand NAND4 (N6146, N6143, N2179, N4847, N5559);
nor NOR3 (N6147, N6134, N5776, N183);
nor NOR4 (N6148, N6121, N4047, N4475, N2451);
and AND2 (N6149, N6147, N4134);
nand NAND4 (N6150, N6145, N4717, N2673, N2794);
nor NOR2 (N6151, N6149, N5625);
or OR2 (N6152, N6150, N3266);
and AND3 (N6153, N6151, N4228, N5496);
not NOT1 (N6154, N6153);
or OR2 (N6155, N6140, N3899);
xor XOR2 (N6156, N6142, N6102);
nor NOR3 (N6157, N6152, N5132, N4595);
xor XOR2 (N6158, N6146, N2382);
and AND3 (N6159, N6131, N5264, N894);
nor NOR3 (N6160, N6158, N4310, N751);
or OR2 (N6161, N6148, N3977);
and AND2 (N6162, N6144, N3369);
and AND2 (N6163, N6159, N3314);
buf BUF1 (N6164, N6156);
buf BUF1 (N6165, N6112);
nor NOR3 (N6166, N6155, N4227, N1138);
xor XOR2 (N6167, N6164, N619);
nor NOR3 (N6168, N6154, N2866, N1382);
xor XOR2 (N6169, N6166, N3209);
nand NAND3 (N6170, N6168, N2738, N3621);
nand NAND4 (N6171, N6163, N2730, N5464, N2204);
and AND2 (N6172, N6167, N4718);
nor NOR2 (N6173, N6172, N3246);
nand NAND4 (N6174, N6165, N2910, N2512, N807);
or OR4 (N6175, N6173, N3184, N708, N4840);
and AND4 (N6176, N6170, N4308, N661, N6104);
and AND4 (N6177, N6171, N1914, N5886, N538);
nand NAND2 (N6178, N6157, N1711);
nand NAND2 (N6179, N6161, N881);
nand NAND4 (N6180, N6175, N5223, N1997, N3062);
or OR4 (N6181, N6180, N3654, N2165, N3515);
xor XOR2 (N6182, N6162, N274);
buf BUF1 (N6183, N6181);
nor NOR4 (N6184, N6128, N5952, N2109, N1310);
not NOT1 (N6185, N6169);
or OR4 (N6186, N6176, N5644, N2669, N581);
xor XOR2 (N6187, N6160, N3925);
nand NAND2 (N6188, N6178, N3299);
xor XOR2 (N6189, N6187, N385);
xor XOR2 (N6190, N6174, N2956);
xor XOR2 (N6191, N6182, N1503);
buf BUF1 (N6192, N6189);
not NOT1 (N6193, N6177);
nand NAND4 (N6194, N6188, N3510, N5673, N436);
or OR4 (N6195, N6194, N5590, N4978, N5527);
xor XOR2 (N6196, N6192, N1145);
nand NAND3 (N6197, N6193, N1317, N6070);
not NOT1 (N6198, N6179);
xor XOR2 (N6199, N6183, N2247);
or OR4 (N6200, N6186, N2896, N6132, N2166);
or OR2 (N6201, N6200, N244);
not NOT1 (N6202, N6198);
and AND2 (N6203, N6197, N2309);
nor NOR2 (N6204, N6202, N3668);
not NOT1 (N6205, N6195);
and AND4 (N6206, N6201, N1794, N867, N3130);
and AND2 (N6207, N6199, N1584);
buf BUF1 (N6208, N6185);
or OR4 (N6209, N6207, N723, N341, N5902);
not NOT1 (N6210, N6184);
xor XOR2 (N6211, N6206, N1453);
or OR2 (N6212, N6203, N2818);
nand NAND2 (N6213, N6209, N5349);
not NOT1 (N6214, N6205);
xor XOR2 (N6215, N6212, N1354);
and AND2 (N6216, N6215, N2320);
xor XOR2 (N6217, N6216, N3374);
nand NAND4 (N6218, N6213, N5834, N1617, N4876);
nor NOR2 (N6219, N6191, N2369);
buf BUF1 (N6220, N6214);
or OR4 (N6221, N6211, N4002, N5160, N3395);
xor XOR2 (N6222, N6219, N5673);
nor NOR4 (N6223, N6190, N2280, N212, N3865);
buf BUF1 (N6224, N6220);
xor XOR2 (N6225, N6221, N3521);
xor XOR2 (N6226, N6204, N807);
and AND4 (N6227, N6196, N633, N873, N1835);
xor XOR2 (N6228, N6218, N2);
buf BUF1 (N6229, N6217);
buf BUF1 (N6230, N6229);
nor NOR2 (N6231, N6228, N2969);
or OR4 (N6232, N6224, N2, N1967, N6023);
not NOT1 (N6233, N6232);
not NOT1 (N6234, N6210);
nor NOR3 (N6235, N6231, N1727, N3335);
buf BUF1 (N6236, N6230);
xor XOR2 (N6237, N6223, N4628);
and AND3 (N6238, N6208, N3859, N353);
xor XOR2 (N6239, N6222, N1656);
not NOT1 (N6240, N6238);
and AND3 (N6241, N6239, N88, N4916);
or OR3 (N6242, N6234, N3584, N4161);
or OR2 (N6243, N6227, N759);
buf BUF1 (N6244, N6233);
nand NAND3 (N6245, N6244, N2, N620);
buf BUF1 (N6246, N6225);
nor NOR2 (N6247, N6246, N4220);
nand NAND3 (N6248, N6226, N3081, N3112);
nor NOR3 (N6249, N6243, N6222, N2672);
xor XOR2 (N6250, N6242, N1237);
nor NOR4 (N6251, N6235, N430, N3371, N2363);
and AND4 (N6252, N6240, N4501, N394, N3036);
buf BUF1 (N6253, N6250);
nor NOR4 (N6254, N6237, N5011, N2312, N233);
and AND3 (N6255, N6251, N5343, N519);
not NOT1 (N6256, N6253);
xor XOR2 (N6257, N6256, N113);
nand NAND3 (N6258, N6252, N6176, N3130);
and AND3 (N6259, N6245, N5405, N6084);
nor NOR4 (N6260, N6249, N5057, N3575, N1125);
nand NAND2 (N6261, N6260, N3329);
or OR2 (N6262, N6241, N5410);
buf BUF1 (N6263, N6248);
xor XOR2 (N6264, N6259, N1871);
not NOT1 (N6265, N6264);
or OR3 (N6266, N6254, N2738, N4313);
or OR2 (N6267, N6262, N5125);
nor NOR2 (N6268, N6263, N3526);
buf BUF1 (N6269, N6236);
nand NAND4 (N6270, N6261, N3353, N1588, N5414);
and AND4 (N6271, N6266, N5228, N5069, N2152);
or OR3 (N6272, N6255, N5362, N1323);
nand NAND4 (N6273, N6268, N4553, N3586, N5625);
buf BUF1 (N6274, N6258);
xor XOR2 (N6275, N6273, N5965);
xor XOR2 (N6276, N6247, N2541);
nand NAND2 (N6277, N6276, N5);
buf BUF1 (N6278, N6267);
nand NAND3 (N6279, N6272, N3828, N4540);
not NOT1 (N6280, N6269);
or OR3 (N6281, N6274, N790, N5005);
nand NAND2 (N6282, N6280, N4658);
nor NOR4 (N6283, N6281, N2467, N1932, N887);
or OR4 (N6284, N6275, N2894, N2253, N6161);
or OR3 (N6285, N6282, N5812, N2449);
xor XOR2 (N6286, N6285, N1083);
not NOT1 (N6287, N6284);
and AND4 (N6288, N6270, N3902, N1569, N2327);
or OR4 (N6289, N6279, N3388, N504, N4879);
nand NAND3 (N6290, N6278, N4362, N4344);
not NOT1 (N6291, N6257);
or OR4 (N6292, N6291, N1471, N3994, N2360);
not NOT1 (N6293, N6290);
nand NAND3 (N6294, N6293, N5069, N5778);
xor XOR2 (N6295, N6288, N5783);
not NOT1 (N6296, N6295);
or OR3 (N6297, N6292, N5278, N1668);
and AND2 (N6298, N6286, N1623);
or OR3 (N6299, N6271, N2105, N5184);
not NOT1 (N6300, N6265);
and AND4 (N6301, N6297, N5194, N4684, N3446);
or OR2 (N6302, N6287, N3272);
and AND4 (N6303, N6289, N3265, N2676, N3002);
nor NOR4 (N6304, N6300, N2381, N4537, N1291);
not NOT1 (N6305, N6304);
or OR3 (N6306, N6296, N5460, N1482);
xor XOR2 (N6307, N6299, N1912);
and AND3 (N6308, N6298, N3232, N5705);
buf BUF1 (N6309, N6307);
or OR4 (N6310, N6283, N2363, N2549, N3904);
nor NOR2 (N6311, N6277, N266);
not NOT1 (N6312, N6310);
nor NOR3 (N6313, N6308, N5469, N1208);
not NOT1 (N6314, N6302);
buf BUF1 (N6315, N6311);
nor NOR3 (N6316, N6294, N130, N1288);
and AND3 (N6317, N6301, N5276, N6219);
xor XOR2 (N6318, N6315, N1250);
and AND2 (N6319, N6313, N2645);
and AND4 (N6320, N6314, N1287, N3504, N239);
xor XOR2 (N6321, N6319, N1837);
not NOT1 (N6322, N6317);
or OR2 (N6323, N6306, N1677);
buf BUF1 (N6324, N6312);
nand NAND4 (N6325, N6309, N4118, N5407, N3965);
and AND4 (N6326, N6325, N3648, N5076, N5542);
buf BUF1 (N6327, N6320);
buf BUF1 (N6328, N6322);
not NOT1 (N6329, N6323);
or OR2 (N6330, N6327, N2139);
not NOT1 (N6331, N6303);
xor XOR2 (N6332, N6326, N1149);
nor NOR3 (N6333, N6328, N5135, N1471);
or OR3 (N6334, N6305, N4559, N6281);
not NOT1 (N6335, N6330);
nor NOR4 (N6336, N6324, N3814, N4044, N6090);
or OR4 (N6337, N6332, N4899, N4772, N1942);
nand NAND3 (N6338, N6337, N1586, N2979);
or OR2 (N6339, N6318, N2494);
or OR2 (N6340, N6336, N6286);
or OR4 (N6341, N6339, N3114, N1105, N926);
not NOT1 (N6342, N6341);
nand NAND3 (N6343, N6338, N2457, N6340);
buf BUF1 (N6344, N1766);
not NOT1 (N6345, N6316);
xor XOR2 (N6346, N6342, N5397);
nand NAND2 (N6347, N6329, N4608);
or OR3 (N6348, N6331, N2933, N4073);
nor NOR3 (N6349, N6347, N4011, N1069);
or OR3 (N6350, N6335, N478, N87);
nand NAND2 (N6351, N6344, N6281);
not NOT1 (N6352, N6350);
or OR2 (N6353, N6348, N1912);
nor NOR2 (N6354, N6352, N4840);
not NOT1 (N6355, N6351);
buf BUF1 (N6356, N6349);
or OR4 (N6357, N6321, N6338, N5762, N755);
nand NAND2 (N6358, N6356, N6295);
nor NOR2 (N6359, N6333, N2978);
xor XOR2 (N6360, N6346, N2899);
nand NAND3 (N6361, N6358, N227, N1824);
or OR4 (N6362, N6359, N458, N2081, N5965);
buf BUF1 (N6363, N6345);
and AND3 (N6364, N6354, N4769, N1963);
nand NAND2 (N6365, N6355, N5956);
not NOT1 (N6366, N6365);
xor XOR2 (N6367, N6364, N6074);
or OR3 (N6368, N6362, N1351, N5633);
or OR2 (N6369, N6357, N3439);
not NOT1 (N6370, N6363);
or OR3 (N6371, N6370, N122, N5476);
not NOT1 (N6372, N6367);
or OR3 (N6373, N6371, N762, N5907);
and AND4 (N6374, N6334, N1537, N4660, N1280);
or OR3 (N6375, N6360, N5117, N315);
nor NOR4 (N6376, N6372, N1397, N4971, N4799);
nand NAND3 (N6377, N6374, N5354, N4553);
xor XOR2 (N6378, N6373, N3808);
nand NAND3 (N6379, N6366, N190, N4568);
or OR2 (N6380, N6353, N711);
nor NOR3 (N6381, N6375, N5433, N1363);
xor XOR2 (N6382, N6378, N4069);
nand NAND2 (N6383, N6377, N876);
nand NAND3 (N6384, N6368, N6149, N5004);
xor XOR2 (N6385, N6343, N2133);
or OR3 (N6386, N6369, N4175, N2396);
buf BUF1 (N6387, N6381);
or OR2 (N6388, N6380, N6168);
and AND4 (N6389, N6382, N3400, N5256, N4387);
and AND3 (N6390, N6383, N815, N3562);
nand NAND2 (N6391, N6384, N2745);
and AND2 (N6392, N6387, N1768);
and AND2 (N6393, N6386, N6106);
or OR2 (N6394, N6389, N4313);
buf BUF1 (N6395, N6394);
not NOT1 (N6396, N6395);
xor XOR2 (N6397, N6396, N1219);
buf BUF1 (N6398, N6391);
buf BUF1 (N6399, N6392);
nand NAND2 (N6400, N6388, N2247);
nor NOR3 (N6401, N6400, N3212, N4115);
nor NOR4 (N6402, N6401, N1762, N5248, N2243);
nor NOR2 (N6403, N6399, N396);
and AND2 (N6404, N6403, N6375);
buf BUF1 (N6405, N6404);
not NOT1 (N6406, N6397);
nand NAND4 (N6407, N6376, N3488, N4297, N6027);
nor NOR3 (N6408, N6361, N4662, N920);
xor XOR2 (N6409, N6407, N1375);
buf BUF1 (N6410, N6402);
not NOT1 (N6411, N6379);
and AND3 (N6412, N6409, N5124, N4519);
and AND3 (N6413, N6406, N2123, N181);
buf BUF1 (N6414, N6405);
nand NAND4 (N6415, N6410, N3678, N2383, N3018);
or OR4 (N6416, N6393, N1638, N3538, N1924);
and AND4 (N6417, N6416, N5886, N3334, N2698);
or OR3 (N6418, N6390, N5211, N4465);
xor XOR2 (N6419, N6413, N2559);
or OR3 (N6420, N6411, N5788, N4583);
nand NAND2 (N6421, N6419, N5543);
nor NOR3 (N6422, N6421, N5809, N1695);
or OR3 (N6423, N6408, N2760, N212);
nand NAND3 (N6424, N6417, N5976, N2552);
nand NAND3 (N6425, N6398, N5856, N1034);
nor NOR2 (N6426, N6412, N4529);
nand NAND3 (N6427, N6426, N35, N1236);
or OR3 (N6428, N6414, N5130, N4043);
nand NAND4 (N6429, N6425, N1326, N1603, N4417);
or OR3 (N6430, N6424, N1204, N4354);
xor XOR2 (N6431, N6428, N1353);
not NOT1 (N6432, N6427);
or OR3 (N6433, N6423, N610, N318);
or OR2 (N6434, N6385, N3033);
xor XOR2 (N6435, N6434, N395);
and AND2 (N6436, N6430, N2193);
nor NOR4 (N6437, N6415, N4160, N5883, N5875);
buf BUF1 (N6438, N6437);
nor NOR2 (N6439, N6436, N856);
nand NAND4 (N6440, N6435, N5308, N4934, N5265);
buf BUF1 (N6441, N6429);
buf BUF1 (N6442, N6433);
buf BUF1 (N6443, N6432);
xor XOR2 (N6444, N6431, N3230);
xor XOR2 (N6445, N6442, N5932);
nor NOR3 (N6446, N6440, N1903, N1496);
not NOT1 (N6447, N6441);
nor NOR3 (N6448, N6447, N5367, N2114);
and AND2 (N6449, N6439, N3006);
and AND2 (N6450, N6438, N3068);
not NOT1 (N6451, N6449);
nand NAND3 (N6452, N6420, N689, N4003);
nand NAND4 (N6453, N6418, N2159, N6113, N1794);
xor XOR2 (N6454, N6452, N5784);
xor XOR2 (N6455, N6446, N220);
nor NOR4 (N6456, N6422, N6435, N4437, N1819);
not NOT1 (N6457, N6453);
buf BUF1 (N6458, N6454);
buf BUF1 (N6459, N6448);
and AND3 (N6460, N6455, N134, N4469);
xor XOR2 (N6461, N6458, N449);
or OR2 (N6462, N6460, N3428);
and AND3 (N6463, N6456, N4337, N1366);
or OR3 (N6464, N6462, N6141, N1170);
buf BUF1 (N6465, N6457);
or OR2 (N6466, N6464, N4877);
and AND2 (N6467, N6465, N1046);
nor NOR3 (N6468, N6443, N2311, N4400);
nor NOR2 (N6469, N6467, N5426);
or OR2 (N6470, N6461, N2239);
xor XOR2 (N6471, N6445, N4496);
nand NAND3 (N6472, N6451, N5130, N3695);
nand NAND2 (N6473, N6444, N4411);
buf BUF1 (N6474, N6469);
or OR2 (N6475, N6474, N1255);
not NOT1 (N6476, N6475);
and AND2 (N6477, N6450, N5591);
nand NAND4 (N6478, N6473, N2410, N704, N4866);
buf BUF1 (N6479, N6476);
not NOT1 (N6480, N6479);
xor XOR2 (N6481, N6471, N5483);
buf BUF1 (N6482, N6468);
nand NAND3 (N6483, N6466, N1803, N4570);
and AND4 (N6484, N6478, N2636, N2337, N4770);
buf BUF1 (N6485, N6483);
and AND3 (N6486, N6459, N1630, N6379);
nand NAND2 (N6487, N6485, N4473);
nand NAND3 (N6488, N6463, N6231, N240);
buf BUF1 (N6489, N6481);
and AND4 (N6490, N6487, N3876, N2834, N684);
xor XOR2 (N6491, N6472, N2922);
nor NOR2 (N6492, N6477, N5175);
nor NOR4 (N6493, N6488, N3796, N3883, N274);
xor XOR2 (N6494, N6480, N3045);
xor XOR2 (N6495, N6486, N4058);
nand NAND4 (N6496, N6484, N2977, N2256, N6265);
nor NOR2 (N6497, N6482, N5167);
buf BUF1 (N6498, N6489);
and AND3 (N6499, N6491, N586, N1156);
xor XOR2 (N6500, N6499, N3329);
nor NOR2 (N6501, N6494, N1733);
not NOT1 (N6502, N6498);
and AND3 (N6503, N6501, N2781, N1219);
xor XOR2 (N6504, N6492, N1183);
not NOT1 (N6505, N6504);
and AND2 (N6506, N6496, N194);
nor NOR2 (N6507, N6503, N4771);
or OR3 (N6508, N6506, N5042, N6472);
and AND2 (N6509, N6495, N3694);
or OR2 (N6510, N6505, N5210);
xor XOR2 (N6511, N6507, N4189);
or OR4 (N6512, N6497, N2525, N6188, N6235);
or OR4 (N6513, N6470, N1753, N3690, N6169);
not NOT1 (N6514, N6512);
nor NOR4 (N6515, N6502, N1681, N4868, N1825);
and AND4 (N6516, N6509, N6091, N4685, N5747);
and AND3 (N6517, N6516, N3664, N3910);
and AND3 (N6518, N6493, N5023, N6361);
nor NOR4 (N6519, N6518, N2933, N4771, N4151);
not NOT1 (N6520, N6513);
xor XOR2 (N6521, N6520, N482);
and AND3 (N6522, N6508, N6050, N1818);
and AND4 (N6523, N6514, N2587, N3821, N3529);
nor NOR2 (N6524, N6490, N4196);
not NOT1 (N6525, N6500);
or OR3 (N6526, N6522, N4283, N576);
nor NOR2 (N6527, N6519, N5245);
and AND4 (N6528, N6517, N3706, N1084, N4713);
nor NOR2 (N6529, N6524, N4903);
buf BUF1 (N6530, N6527);
nand NAND3 (N6531, N6515, N5330, N1046);
not NOT1 (N6532, N6523);
and AND2 (N6533, N6531, N4399);
nand NAND4 (N6534, N6532, N35, N1748, N29);
not NOT1 (N6535, N6521);
buf BUF1 (N6536, N6529);
nor NOR3 (N6537, N6510, N5630, N3555);
or OR3 (N6538, N6525, N2774, N226);
nand NAND4 (N6539, N6511, N4428, N1798, N1654);
xor XOR2 (N6540, N6533, N2700);
nor NOR2 (N6541, N6538, N2980);
or OR3 (N6542, N6540, N4043, N2971);
not NOT1 (N6543, N6530);
not NOT1 (N6544, N6539);
nand NAND2 (N6545, N6528, N2569);
xor XOR2 (N6546, N6537, N2312);
xor XOR2 (N6547, N6542, N4608);
buf BUF1 (N6548, N6543);
xor XOR2 (N6549, N6541, N4826);
nand NAND2 (N6550, N6545, N6423);
and AND3 (N6551, N6550, N5973, N6280);
xor XOR2 (N6552, N6544, N5232);
not NOT1 (N6553, N6551);
nand NAND2 (N6554, N6546, N2042);
not NOT1 (N6555, N6554);
and AND3 (N6556, N6549, N3967, N3048);
nand NAND4 (N6557, N6535, N3282, N3612, N3272);
xor XOR2 (N6558, N6547, N2863);
and AND2 (N6559, N6552, N5348);
nand NAND4 (N6560, N6558, N1081, N3595, N1121);
nand NAND2 (N6561, N6559, N686);
nand NAND2 (N6562, N6561, N1754);
xor XOR2 (N6563, N6556, N469);
not NOT1 (N6564, N6563);
or OR3 (N6565, N6553, N5884, N1868);
xor XOR2 (N6566, N6557, N3931);
and AND2 (N6567, N6564, N3205);
and AND4 (N6568, N6566, N6355, N6107, N3780);
nand NAND4 (N6569, N6568, N3773, N610, N5735);
nor NOR4 (N6570, N6536, N90, N995, N3617);
nand NAND2 (N6571, N6567, N6303);
not NOT1 (N6572, N6526);
buf BUF1 (N6573, N6548);
and AND4 (N6574, N6565, N5022, N5170, N3518);
buf BUF1 (N6575, N6555);
not NOT1 (N6576, N6574);
nor NOR2 (N6577, N6575, N4189);
nand NAND3 (N6578, N6562, N6074, N6429);
nand NAND2 (N6579, N6573, N457);
and AND4 (N6580, N6577, N1523, N1978, N5107);
and AND2 (N6581, N6572, N2979);
not NOT1 (N6582, N6576);
and AND2 (N6583, N6534, N1735);
nor NOR2 (N6584, N6570, N3472);
buf BUF1 (N6585, N6582);
and AND2 (N6586, N6578, N3400);
nor NOR4 (N6587, N6586, N2153, N2057, N5436);
nor NOR3 (N6588, N6583, N419, N1246);
xor XOR2 (N6589, N6587, N1091);
nor NOR2 (N6590, N6581, N6383);
nand NAND2 (N6591, N6580, N3300);
and AND2 (N6592, N6584, N6517);
or OR4 (N6593, N6569, N2865, N4977, N2518);
xor XOR2 (N6594, N6579, N5007);
xor XOR2 (N6595, N6590, N2146);
and AND2 (N6596, N6592, N4099);
buf BUF1 (N6597, N6595);
and AND2 (N6598, N6571, N4029);
or OR4 (N6599, N6585, N2721, N5051, N1547);
and AND2 (N6600, N6588, N2354);
buf BUF1 (N6601, N6600);
or OR3 (N6602, N6597, N3003, N2323);
and AND3 (N6603, N6593, N2308, N2925);
not NOT1 (N6604, N6601);
not NOT1 (N6605, N6599);
buf BUF1 (N6606, N6560);
nand NAND3 (N6607, N6603, N160, N3709);
xor XOR2 (N6608, N6598, N5583);
not NOT1 (N6609, N6608);
xor XOR2 (N6610, N6606, N2552);
and AND4 (N6611, N6589, N1775, N218, N2899);
and AND4 (N6612, N6591, N4574, N6042, N2785);
not NOT1 (N6613, N6609);
or OR4 (N6614, N6604, N4904, N3964, N582);
xor XOR2 (N6615, N6613, N3981);
buf BUF1 (N6616, N6605);
buf BUF1 (N6617, N6616);
or OR4 (N6618, N6612, N187, N5132, N4469);
or OR4 (N6619, N6602, N53, N4247, N3017);
xor XOR2 (N6620, N6615, N4903);
nand NAND4 (N6621, N6594, N2991, N4402, N4158);
and AND3 (N6622, N6610, N401, N5182);
buf BUF1 (N6623, N6620);
or OR2 (N6624, N6622, N3145);
not NOT1 (N6625, N6624);
not NOT1 (N6626, N6611);
nand NAND2 (N6627, N6614, N57);
xor XOR2 (N6628, N6618, N1782);
not NOT1 (N6629, N6628);
buf BUF1 (N6630, N6623);
and AND3 (N6631, N6607, N2398, N2091);
buf BUF1 (N6632, N6629);
nand NAND2 (N6633, N6627, N2427);
nand NAND3 (N6634, N6625, N5871, N2534);
not NOT1 (N6635, N6630);
and AND4 (N6636, N6632, N410, N2899, N324);
or OR4 (N6637, N6636, N4594, N1555, N550);
nor NOR3 (N6638, N6596, N4023, N3170);
nand NAND3 (N6639, N6638, N3306, N4801);
xor XOR2 (N6640, N6619, N1864);
nor NOR3 (N6641, N6637, N967, N6427);
nor NOR3 (N6642, N6639, N801, N5905);
nand NAND2 (N6643, N6635, N2019);
or OR2 (N6644, N6640, N4874);
not NOT1 (N6645, N6626);
nor NOR4 (N6646, N6641, N6330, N5772, N2579);
xor XOR2 (N6647, N6633, N5390);
nor NOR2 (N6648, N6631, N3853);
nor NOR4 (N6649, N6648, N6134, N6557, N2055);
and AND3 (N6650, N6647, N5918, N2067);
buf BUF1 (N6651, N6644);
xor XOR2 (N6652, N6650, N3735);
xor XOR2 (N6653, N6617, N2378);
or OR4 (N6654, N6649, N4369, N3900, N1268);
and AND4 (N6655, N6654, N265, N2389, N5130);
buf BUF1 (N6656, N6653);
or OR4 (N6657, N6655, N6457, N4163, N692);
buf BUF1 (N6658, N6643);
buf BUF1 (N6659, N6656);
nor NOR2 (N6660, N6657, N5654);
xor XOR2 (N6661, N6634, N2906);
nand NAND4 (N6662, N6651, N4588, N4602, N5140);
buf BUF1 (N6663, N6645);
or OR4 (N6664, N6662, N1135, N613, N1630);
not NOT1 (N6665, N6652);
not NOT1 (N6666, N6646);
or OR2 (N6667, N6663, N4519);
nand NAND4 (N6668, N6660, N5146, N4673, N763);
nor NOR2 (N6669, N6665, N4070);
buf BUF1 (N6670, N6666);
not NOT1 (N6671, N6661);
not NOT1 (N6672, N6642);
and AND3 (N6673, N6667, N1414, N1431);
not NOT1 (N6674, N6664);
and AND4 (N6675, N6669, N6440, N6589, N2666);
buf BUF1 (N6676, N6658);
not NOT1 (N6677, N6621);
or OR3 (N6678, N6672, N507, N3514);
nand NAND3 (N6679, N6671, N5053, N2650);
nand NAND2 (N6680, N6678, N5271);
and AND3 (N6681, N6670, N1960, N1117);
nand NAND4 (N6682, N6659, N4547, N4790, N3629);
nand NAND3 (N6683, N6681, N1706, N3765);
nand NAND2 (N6684, N6677, N1300);
nor NOR2 (N6685, N6673, N5201);
not NOT1 (N6686, N6684);
nor NOR3 (N6687, N6680, N6534, N2958);
or OR2 (N6688, N6676, N783);
xor XOR2 (N6689, N6668, N4266);
or OR3 (N6690, N6689, N4433, N1920);
not NOT1 (N6691, N6690);
xor XOR2 (N6692, N6682, N1205);
buf BUF1 (N6693, N6685);
xor XOR2 (N6694, N6687, N5720);
nand NAND3 (N6695, N6693, N5283, N3178);
nor NOR2 (N6696, N6692, N889);
nor NOR4 (N6697, N6694, N6050, N226, N6559);
and AND4 (N6698, N6695, N1628, N650, N6103);
not NOT1 (N6699, N6697);
nor NOR4 (N6700, N6679, N1739, N478, N4676);
buf BUF1 (N6701, N6688);
not NOT1 (N6702, N6675);
or OR2 (N6703, N6691, N4514);
or OR4 (N6704, N6686, N5987, N4210, N39);
not NOT1 (N6705, N6699);
nand NAND3 (N6706, N6683, N6629, N2332);
or OR2 (N6707, N6698, N1799);
not NOT1 (N6708, N6701);
or OR3 (N6709, N6707, N790, N3656);
or OR2 (N6710, N6696, N6021);
not NOT1 (N6711, N6674);
buf BUF1 (N6712, N6703);
not NOT1 (N6713, N6712);
buf BUF1 (N6714, N6709);
not NOT1 (N6715, N6700);
xor XOR2 (N6716, N6713, N3021);
and AND2 (N6717, N6705, N6355);
or OR2 (N6718, N6717, N5459);
nor NOR4 (N6719, N6710, N5821, N6449, N3841);
xor XOR2 (N6720, N6719, N1772);
nand NAND3 (N6721, N6720, N344, N4981);
not NOT1 (N6722, N6708);
not NOT1 (N6723, N6718);
not NOT1 (N6724, N6706);
buf BUF1 (N6725, N6702);
buf BUF1 (N6726, N6725);
and AND2 (N6727, N6704, N5867);
nand NAND2 (N6728, N6724, N5238);
not NOT1 (N6729, N6723);
or OR3 (N6730, N6722, N2212, N6173);
or OR3 (N6731, N6728, N217, N3559);
nor NOR4 (N6732, N6711, N5221, N5236, N1183);
buf BUF1 (N6733, N6715);
not NOT1 (N6734, N6731);
xor XOR2 (N6735, N6732, N1178);
xor XOR2 (N6736, N6733, N4515);
buf BUF1 (N6737, N6730);
nand NAND2 (N6738, N6721, N5250);
not NOT1 (N6739, N6714);
not NOT1 (N6740, N6734);
or OR4 (N6741, N6736, N680, N6669, N3845);
xor XOR2 (N6742, N6739, N1611);
buf BUF1 (N6743, N6729);
and AND2 (N6744, N6716, N4520);
buf BUF1 (N6745, N6738);
nand NAND2 (N6746, N6737, N4233);
nand NAND4 (N6747, N6727, N191, N3631, N4040);
and AND3 (N6748, N6740, N3471, N242);
or OR3 (N6749, N6747, N3402, N4476);
nor NOR2 (N6750, N6749, N1964);
buf BUF1 (N6751, N6750);
nand NAND3 (N6752, N6741, N3019, N6201);
xor XOR2 (N6753, N6746, N5039);
nor NOR3 (N6754, N6752, N3233, N4943);
buf BUF1 (N6755, N6748);
nor NOR4 (N6756, N6754, N4348, N6640, N3987);
and AND3 (N6757, N6755, N2153, N4685);
xor XOR2 (N6758, N6745, N4134);
not NOT1 (N6759, N6726);
nand NAND2 (N6760, N6759, N3859);
xor XOR2 (N6761, N6743, N1459);
nor NOR4 (N6762, N6751, N4872, N3298, N4847);
and AND2 (N6763, N6735, N343);
nand NAND2 (N6764, N6756, N5682);
not NOT1 (N6765, N6757);
not NOT1 (N6766, N6762);
nand NAND4 (N6767, N6765, N2782, N2958, N4626);
and AND2 (N6768, N6763, N1156);
xor XOR2 (N6769, N6742, N5897);
nand NAND3 (N6770, N6769, N4291, N2690);
nand NAND2 (N6771, N6767, N6170);
not NOT1 (N6772, N6768);
or OR4 (N6773, N6771, N2117, N6379, N4141);
not NOT1 (N6774, N6744);
not NOT1 (N6775, N6758);
nand NAND3 (N6776, N6764, N3668, N5725);
not NOT1 (N6777, N6772);
not NOT1 (N6778, N6774);
nand NAND3 (N6779, N6777, N4846, N1527);
nand NAND4 (N6780, N6776, N500, N4851, N6744);
or OR3 (N6781, N6761, N692, N1669);
buf BUF1 (N6782, N6780);
buf BUF1 (N6783, N6775);
xor XOR2 (N6784, N6781, N5946);
nand NAND4 (N6785, N6760, N6214, N5118, N3205);
buf BUF1 (N6786, N6783);
nand NAND4 (N6787, N6784, N6703, N4476, N5381);
and AND3 (N6788, N6766, N4453, N125);
xor XOR2 (N6789, N6785, N4532);
buf BUF1 (N6790, N6782);
or OR4 (N6791, N6790, N1781, N3854, N3376);
nand NAND2 (N6792, N6786, N2471);
buf BUF1 (N6793, N6789);
xor XOR2 (N6794, N6792, N4656);
not NOT1 (N6795, N6787);
xor XOR2 (N6796, N6793, N1671);
nand NAND4 (N6797, N6778, N5492, N1858, N2002);
xor XOR2 (N6798, N6779, N2106);
xor XOR2 (N6799, N6797, N3762);
not NOT1 (N6800, N6798);
and AND2 (N6801, N6770, N1272);
and AND3 (N6802, N6773, N853, N1386);
nand NAND2 (N6803, N6753, N365);
buf BUF1 (N6804, N6799);
buf BUF1 (N6805, N6801);
nor NOR4 (N6806, N6803, N3343, N1289, N5233);
and AND2 (N6807, N6806, N2042);
xor XOR2 (N6808, N6800, N5879);
nor NOR3 (N6809, N6808, N747, N3712);
not NOT1 (N6810, N6802);
nor NOR4 (N6811, N6807, N3715, N4687, N4843);
nand NAND3 (N6812, N6788, N4336, N6287);
or OR2 (N6813, N6795, N4312);
xor XOR2 (N6814, N6791, N1895);
buf BUF1 (N6815, N6812);
xor XOR2 (N6816, N6815, N3928);
or OR4 (N6817, N6809, N3301, N3946, N3606);
or OR4 (N6818, N6816, N203, N4442, N6216);
and AND3 (N6819, N6796, N5726, N5324);
nand NAND2 (N6820, N6817, N2507);
buf BUF1 (N6821, N6804);
xor XOR2 (N6822, N6794, N5539);
or OR2 (N6823, N6819, N314);
not NOT1 (N6824, N6813);
xor XOR2 (N6825, N6818, N1157);
nand NAND4 (N6826, N6810, N508, N4661, N5011);
buf BUF1 (N6827, N6822);
not NOT1 (N6828, N6820);
and AND3 (N6829, N6825, N4676, N2239);
buf BUF1 (N6830, N6811);
nor NOR3 (N6831, N6805, N338, N2354);
or OR4 (N6832, N6829, N664, N5864, N5462);
nor NOR4 (N6833, N6824, N4840, N3871, N3486);
nand NAND4 (N6834, N6823, N4259, N894, N3322);
buf BUF1 (N6835, N6832);
not NOT1 (N6836, N6828);
xor XOR2 (N6837, N6827, N214);
and AND2 (N6838, N6831, N5320);
nand NAND4 (N6839, N6834, N5079, N62, N3366);
or OR2 (N6840, N6838, N4919);
nor NOR2 (N6841, N6840, N2610);
nor NOR2 (N6842, N6839, N6277);
xor XOR2 (N6843, N6821, N3146);
nand NAND3 (N6844, N6833, N1620, N4770);
xor XOR2 (N6845, N6837, N5551);
not NOT1 (N6846, N6830);
buf BUF1 (N6847, N6844);
xor XOR2 (N6848, N6841, N6280);
or OR2 (N6849, N6826, N1057);
nand NAND2 (N6850, N6848, N1376);
buf BUF1 (N6851, N6850);
and AND2 (N6852, N6843, N2632);
and AND3 (N6853, N6835, N6112, N4042);
not NOT1 (N6854, N6836);
buf BUF1 (N6855, N6854);
or OR3 (N6856, N6845, N5960, N920);
nand NAND2 (N6857, N6846, N313);
nand NAND2 (N6858, N6847, N1908);
buf BUF1 (N6859, N6852);
xor XOR2 (N6860, N6858, N5180);
and AND3 (N6861, N6856, N5773, N2587);
buf BUF1 (N6862, N6861);
nand NAND2 (N6863, N6814, N116);
not NOT1 (N6864, N6857);
nor NOR3 (N6865, N6851, N6302, N4402);
or OR4 (N6866, N6863, N3907, N4886, N2865);
buf BUF1 (N6867, N6853);
nand NAND2 (N6868, N6866, N4610);
or OR3 (N6869, N6855, N1280, N5967);
xor XOR2 (N6870, N6860, N4442);
nor NOR4 (N6871, N6867, N5113, N4566, N6782);
and AND2 (N6872, N6849, N3453);
nand NAND3 (N6873, N6872, N4145, N1940);
not NOT1 (N6874, N6865);
nand NAND2 (N6875, N6859, N49);
xor XOR2 (N6876, N6864, N5615);
not NOT1 (N6877, N6862);
and AND3 (N6878, N6875, N2374, N2933);
nand NAND4 (N6879, N6842, N5029, N2017, N6014);
nor NOR2 (N6880, N6873, N1291);
not NOT1 (N6881, N6879);
not NOT1 (N6882, N6869);
xor XOR2 (N6883, N6870, N2391);
not NOT1 (N6884, N6871);
not NOT1 (N6885, N6880);
not NOT1 (N6886, N6877);
nand NAND2 (N6887, N6868, N3807);
not NOT1 (N6888, N6887);
nand NAND3 (N6889, N6874, N2028, N4689);
nand NAND2 (N6890, N6883, N3914);
or OR4 (N6891, N6885, N2145, N3939, N5357);
or OR3 (N6892, N6876, N2502, N3594);
not NOT1 (N6893, N6886);
and AND3 (N6894, N6878, N2291, N6595);
or OR2 (N6895, N6888, N5075);
xor XOR2 (N6896, N6891, N2218);
nand NAND2 (N6897, N6881, N2336);
buf BUF1 (N6898, N6893);
and AND2 (N6899, N6895, N1428);
and AND2 (N6900, N6898, N5239);
or OR2 (N6901, N6884, N6615);
and AND3 (N6902, N6894, N3607, N505);
and AND2 (N6903, N6892, N1775);
nor NOR2 (N6904, N6890, N1433);
and AND3 (N6905, N6904, N1023, N170);
nor NOR3 (N6906, N6889, N2370, N6724);
buf BUF1 (N6907, N6903);
nor NOR3 (N6908, N6901, N5444, N5241);
or OR2 (N6909, N6908, N2581);
or OR3 (N6910, N6899, N2427, N343);
nand NAND2 (N6911, N6902, N4466);
not NOT1 (N6912, N6911);
nor NOR3 (N6913, N6909, N1216, N6648);
buf BUF1 (N6914, N6882);
and AND3 (N6915, N6897, N4790, N1180);
nand NAND4 (N6916, N6896, N3237, N1954, N5663);
nor NOR2 (N6917, N6914, N1267);
nor NOR4 (N6918, N6916, N3723, N4107, N6);
nor NOR4 (N6919, N6912, N3095, N6188, N4317);
not NOT1 (N6920, N6918);
nand NAND2 (N6921, N6905, N2780);
xor XOR2 (N6922, N6921, N6893);
and AND4 (N6923, N6906, N5251, N3339, N6541);
and AND2 (N6924, N6910, N1854);
nand NAND3 (N6925, N6922, N4820, N6863);
nand NAND4 (N6926, N6917, N3945, N909, N568);
not NOT1 (N6927, N6925);
not NOT1 (N6928, N6923);
and AND4 (N6929, N6913, N6151, N325, N3384);
or OR3 (N6930, N6929, N6925, N1487);
or OR3 (N6931, N6924, N4204, N4185);
or OR4 (N6932, N6915, N4482, N4320, N1537);
buf BUF1 (N6933, N6907);
and AND2 (N6934, N6919, N3325);
or OR2 (N6935, N6930, N6390);
nor NOR2 (N6936, N6926, N1828);
and AND2 (N6937, N6933, N6721);
xor XOR2 (N6938, N6932, N1219);
not NOT1 (N6939, N6927);
buf BUF1 (N6940, N6900);
buf BUF1 (N6941, N6935);
or OR2 (N6942, N6920, N661);
nand NAND3 (N6943, N6940, N1362, N1160);
nand NAND2 (N6944, N6937, N6081);
buf BUF1 (N6945, N6943);
or OR4 (N6946, N6942, N5784, N2261, N1696);
nand NAND2 (N6947, N6939, N2638);
buf BUF1 (N6948, N6931);
xor XOR2 (N6949, N6946, N111);
nand NAND2 (N6950, N6944, N1106);
buf BUF1 (N6951, N6928);
nand NAND4 (N6952, N6936, N4467, N3152, N2252);
nand NAND3 (N6953, N6950, N6049, N1848);
or OR3 (N6954, N6951, N5529, N706);
nand NAND3 (N6955, N6938, N3114, N3623);
or OR3 (N6956, N6953, N6290, N202);
nand NAND2 (N6957, N6955, N1395);
nand NAND4 (N6958, N6956, N5399, N3320, N216);
nor NOR3 (N6959, N6947, N3053, N2765);
nor NOR2 (N6960, N6945, N5631);
and AND3 (N6961, N6954, N839, N1285);
and AND4 (N6962, N6941, N6214, N3090, N1069);
or OR4 (N6963, N6948, N4618, N5598, N2826);
buf BUF1 (N6964, N6934);
not NOT1 (N6965, N6957);
nand NAND3 (N6966, N6965, N2853, N4188);
xor XOR2 (N6967, N6952, N5957);
and AND2 (N6968, N6949, N2453);
nand NAND4 (N6969, N6963, N2592, N6508, N5368);
buf BUF1 (N6970, N6962);
not NOT1 (N6971, N6958);
nand NAND2 (N6972, N6966, N608);
nand NAND2 (N6973, N6969, N1805);
or OR3 (N6974, N6964, N952, N1730);
or OR4 (N6975, N6967, N6286, N462, N3838);
nand NAND4 (N6976, N6959, N6591, N2809, N4387);
nor NOR2 (N6977, N6961, N4852);
nand NAND4 (N6978, N6960, N689, N3437, N4252);
nor NOR2 (N6979, N6976, N6025);
nand NAND4 (N6980, N6973, N2034, N4385, N3994);
buf BUF1 (N6981, N6970);
buf BUF1 (N6982, N6974);
xor XOR2 (N6983, N6981, N3766);
or OR3 (N6984, N6968, N3885, N4717);
and AND4 (N6985, N6982, N5341, N1302, N1855);
xor XOR2 (N6986, N6975, N2303);
not NOT1 (N6987, N6986);
not NOT1 (N6988, N6984);
and AND3 (N6989, N6971, N3937, N2272);
and AND3 (N6990, N6979, N5693, N710);
xor XOR2 (N6991, N6987, N956);
or OR3 (N6992, N6978, N5517, N4688);
nor NOR2 (N6993, N6988, N3761);
and AND3 (N6994, N6993, N1785, N5227);
nand NAND2 (N6995, N6985, N2552);
nand NAND2 (N6996, N6994, N5797);
nor NOR4 (N6997, N6995, N6480, N5752, N1671);
buf BUF1 (N6998, N6992);
buf BUF1 (N6999, N6972);
buf BUF1 (N7000, N6980);
buf BUF1 (N7001, N6997);
and AND2 (N7002, N7001, N6020);
xor XOR2 (N7003, N6998, N5887);
not NOT1 (N7004, N6996);
xor XOR2 (N7005, N6977, N4589);
nor NOR3 (N7006, N7002, N3150, N1114);
not NOT1 (N7007, N6983);
nor NOR4 (N7008, N6999, N2869, N6415, N1809);
nor NOR3 (N7009, N7007, N3612, N652);
and AND2 (N7010, N7008, N2288);
xor XOR2 (N7011, N7009, N6373);
not NOT1 (N7012, N7000);
and AND3 (N7013, N6989, N1070, N690);
xor XOR2 (N7014, N6991, N3363);
or OR3 (N7015, N7005, N634, N34);
nor NOR4 (N7016, N7012, N3324, N3034, N406);
xor XOR2 (N7017, N7014, N5928);
and AND2 (N7018, N7006, N6378);
xor XOR2 (N7019, N7003, N5354);
xor XOR2 (N7020, N7010, N4387);
and AND4 (N7021, N7015, N1298, N1579, N2376);
or OR4 (N7022, N6990, N5921, N849, N3921);
or OR3 (N7023, N7013, N5456, N2887);
nor NOR3 (N7024, N7023, N689, N3279);
nor NOR4 (N7025, N7004, N5540, N1932, N2257);
nand NAND2 (N7026, N7018, N220);
xor XOR2 (N7027, N7017, N4916);
not NOT1 (N7028, N7020);
buf BUF1 (N7029, N7016);
nand NAND3 (N7030, N7019, N579, N2751);
or OR4 (N7031, N7028, N2535, N2009, N6424);
buf BUF1 (N7032, N7030);
and AND3 (N7033, N7025, N6675, N5301);
nand NAND4 (N7034, N7011, N2521, N5883, N2018);
nand NAND4 (N7035, N7034, N2978, N3899, N4567);
not NOT1 (N7036, N7021);
not NOT1 (N7037, N7036);
nor NOR2 (N7038, N7024, N1531);
nand NAND3 (N7039, N7037, N2485, N4752);
and AND4 (N7040, N7035, N3150, N5069, N4582);
xor XOR2 (N7041, N7038, N6640);
buf BUF1 (N7042, N7031);
buf BUF1 (N7043, N7040);
xor XOR2 (N7044, N7032, N4836);
buf BUF1 (N7045, N7027);
xor XOR2 (N7046, N7026, N5889);
buf BUF1 (N7047, N7022);
nand NAND2 (N7048, N7042, N1632);
xor XOR2 (N7049, N7048, N1066);
xor XOR2 (N7050, N7049, N4581);
xor XOR2 (N7051, N7045, N6707);
nand NAND3 (N7052, N7050, N3712, N905);
and AND3 (N7053, N7041, N1184, N6548);
or OR3 (N7054, N7052, N136, N2022);
buf BUF1 (N7055, N7046);
xor XOR2 (N7056, N7033, N592);
xor XOR2 (N7057, N7044, N2454);
not NOT1 (N7058, N7054);
nand NAND4 (N7059, N7047, N1374, N122, N2295);
nor NOR2 (N7060, N7051, N1241);
xor XOR2 (N7061, N7029, N4608);
buf BUF1 (N7062, N7039);
nand NAND2 (N7063, N7055, N3846);
not NOT1 (N7064, N7056);
nand NAND3 (N7065, N7060, N326, N63);
not NOT1 (N7066, N7059);
nor NOR3 (N7067, N7063, N3509, N4126);
nor NOR2 (N7068, N7061, N1663);
not NOT1 (N7069, N7058);
not NOT1 (N7070, N7066);
and AND2 (N7071, N7069, N1789);
not NOT1 (N7072, N7053);
nand NAND3 (N7073, N7071, N1341, N6471);
not NOT1 (N7074, N7064);
and AND3 (N7075, N7068, N3606, N1699);
not NOT1 (N7076, N7065);
or OR2 (N7077, N7074, N2967);
nor NOR2 (N7078, N7077, N4775);
nor NOR2 (N7079, N7043, N6317);
buf BUF1 (N7080, N7075);
or OR2 (N7081, N7078, N1822);
buf BUF1 (N7082, N7070);
not NOT1 (N7083, N7062);
and AND2 (N7084, N7082, N4722);
or OR2 (N7085, N7073, N1021);
buf BUF1 (N7086, N7083);
xor XOR2 (N7087, N7081, N2342);
xor XOR2 (N7088, N7072, N4495);
nor NOR3 (N7089, N7086, N1830, N5642);
nor NOR3 (N7090, N7076, N1974, N1165);
nand NAND2 (N7091, N7089, N6681);
nor NOR2 (N7092, N7090, N5178);
nor NOR3 (N7093, N7088, N2962, N5414);
nand NAND3 (N7094, N7085, N4659, N4314);
nor NOR4 (N7095, N7092, N614, N6721, N4685);
nand NAND3 (N7096, N7067, N6460, N5246);
nor NOR2 (N7097, N7057, N6734);
xor XOR2 (N7098, N7080, N6899);
nand NAND4 (N7099, N7098, N2065, N2647, N2053);
buf BUF1 (N7100, N7079);
buf BUF1 (N7101, N7099);
or OR4 (N7102, N7093, N3264, N2475, N2154);
and AND4 (N7103, N7101, N1093, N1687, N1575);
and AND3 (N7104, N7084, N4441, N2826);
or OR2 (N7105, N7102, N2648);
xor XOR2 (N7106, N7100, N4233);
or OR3 (N7107, N7095, N5745, N4783);
or OR2 (N7108, N7097, N7);
not NOT1 (N7109, N7087);
buf BUF1 (N7110, N7109);
buf BUF1 (N7111, N7107);
buf BUF1 (N7112, N7091);
buf BUF1 (N7113, N7104);
buf BUF1 (N7114, N7105);
or OR4 (N7115, N7110, N3492, N2619, N2660);
not NOT1 (N7116, N7106);
xor XOR2 (N7117, N7116, N6145);
xor XOR2 (N7118, N7113, N6603);
not NOT1 (N7119, N7117);
or OR3 (N7120, N7115, N2645, N6965);
and AND4 (N7121, N7120, N7116, N6737, N5536);
xor XOR2 (N7122, N7118, N2508);
buf BUF1 (N7123, N7119);
not NOT1 (N7124, N7103);
buf BUF1 (N7125, N7108);
and AND4 (N7126, N7094, N245, N2347, N1940);
or OR4 (N7127, N7111, N6974, N5665, N1254);
not NOT1 (N7128, N7125);
xor XOR2 (N7129, N7121, N4261);
xor XOR2 (N7130, N7126, N605);
xor XOR2 (N7131, N7122, N1162);
xor XOR2 (N7132, N7124, N466);
xor XOR2 (N7133, N7131, N5642);
not NOT1 (N7134, N7114);
nor NOR4 (N7135, N7132, N5977, N6387, N1558);
nor NOR3 (N7136, N7128, N4524, N2661);
not NOT1 (N7137, N7112);
nor NOR3 (N7138, N7129, N388, N2952);
nor NOR2 (N7139, N7096, N6861);
nand NAND4 (N7140, N7135, N52, N2124, N830);
xor XOR2 (N7141, N7123, N1408);
buf BUF1 (N7142, N7137);
nor NOR3 (N7143, N7138, N681, N6154);
or OR4 (N7144, N7136, N732, N2223, N4807);
nor NOR2 (N7145, N7139, N6966);
and AND4 (N7146, N7142, N5663, N7007, N5528);
nor NOR2 (N7147, N7144, N1186);
and AND4 (N7148, N7145, N4482, N6458, N4338);
or OR4 (N7149, N7133, N3808, N3150, N6474);
nor NOR3 (N7150, N7147, N2523, N3905);
nand NAND4 (N7151, N7140, N2528, N4760, N3812);
xor XOR2 (N7152, N7141, N1018);
nand NAND3 (N7153, N7150, N3119, N1976);
buf BUF1 (N7154, N7151);
nand NAND2 (N7155, N7127, N3836);
not NOT1 (N7156, N7155);
xor XOR2 (N7157, N7149, N4827);
xor XOR2 (N7158, N7143, N3632);
not NOT1 (N7159, N7157);
and AND2 (N7160, N7134, N6369);
buf BUF1 (N7161, N7158);
buf BUF1 (N7162, N7153);
and AND4 (N7163, N7162, N723, N356, N3524);
buf BUF1 (N7164, N7160);
nand NAND4 (N7165, N7159, N478, N6199, N977);
nor NOR3 (N7166, N7130, N2079, N1721);
xor XOR2 (N7167, N7156, N6510);
or OR3 (N7168, N7152, N6497, N1469);
nand NAND4 (N7169, N7163, N2750, N4695, N6273);
or OR4 (N7170, N7165, N6719, N3505, N1002);
or OR3 (N7171, N7148, N2219, N6485);
xor XOR2 (N7172, N7171, N5364);
nand NAND2 (N7173, N7164, N3164);
buf BUF1 (N7174, N7166);
nor NOR3 (N7175, N7161, N5217, N5726);
nand NAND2 (N7176, N7146, N3159);
and AND3 (N7177, N7175, N3084, N2452);
and AND4 (N7178, N7172, N3248, N2511, N3526);
and AND4 (N7179, N7176, N1444, N5490, N972);
buf BUF1 (N7180, N7178);
nand NAND4 (N7181, N7173, N5869, N4997, N2964);
not NOT1 (N7182, N7168);
nor NOR3 (N7183, N7174, N6651, N4748);
nand NAND4 (N7184, N7167, N5573, N3036, N6013);
nand NAND3 (N7185, N7179, N4016, N3117);
buf BUF1 (N7186, N7170);
xor XOR2 (N7187, N7154, N1589);
nor NOR2 (N7188, N7181, N1680);
not NOT1 (N7189, N7180);
not NOT1 (N7190, N7183);
and AND4 (N7191, N7187, N4436, N4293, N5723);
buf BUF1 (N7192, N7185);
xor XOR2 (N7193, N7188, N4191);
and AND4 (N7194, N7177, N745, N4383, N2924);
nand NAND4 (N7195, N7182, N4549, N6472, N4944);
buf BUF1 (N7196, N7186);
or OR4 (N7197, N7189, N6236, N5132, N3602);
nor NOR2 (N7198, N7169, N6643);
not NOT1 (N7199, N7192);
nand NAND3 (N7200, N7197, N6486, N5923);
and AND4 (N7201, N7184, N529, N2300, N6462);
buf BUF1 (N7202, N7198);
nor NOR2 (N7203, N7202, N4342);
nand NAND4 (N7204, N7203, N4189, N2132, N6876);
nor NOR4 (N7205, N7195, N5743, N43, N3439);
or OR4 (N7206, N7196, N3992, N1795, N3460);
and AND4 (N7207, N7205, N3706, N6460, N5262);
or OR2 (N7208, N7207, N130);
buf BUF1 (N7209, N7204);
and AND3 (N7210, N7208, N2110, N2051);
or OR3 (N7211, N7200, N5393, N1742);
and AND3 (N7212, N7194, N2226, N4473);
or OR2 (N7213, N7193, N4123);
not NOT1 (N7214, N7199);
or OR2 (N7215, N7191, N1932);
or OR3 (N7216, N7209, N6209, N2291);
buf BUF1 (N7217, N7212);
nand NAND2 (N7218, N7217, N7152);
nand NAND3 (N7219, N7211, N2825, N5382);
nor NOR4 (N7220, N7206, N2926, N5988, N3111);
nor NOR2 (N7221, N7201, N885);
nor NOR4 (N7222, N7210, N807, N309, N5759);
and AND4 (N7223, N7220, N2703, N2810, N6896);
nand NAND4 (N7224, N7215, N129, N646, N5604);
and AND4 (N7225, N7223, N3373, N2787, N4212);
buf BUF1 (N7226, N7224);
and AND4 (N7227, N7225, N5166, N221, N1675);
buf BUF1 (N7228, N7221);
nor NOR2 (N7229, N7214, N958);
nor NOR4 (N7230, N7229, N756, N5050, N6541);
buf BUF1 (N7231, N7222);
xor XOR2 (N7232, N7190, N2877);
xor XOR2 (N7233, N7228, N897);
or OR2 (N7234, N7230, N964);
or OR2 (N7235, N7233, N4071);
xor XOR2 (N7236, N7231, N3334);
not NOT1 (N7237, N7219);
nor NOR4 (N7238, N7232, N5388, N5752, N6420);
buf BUF1 (N7239, N7235);
buf BUF1 (N7240, N7236);
nand NAND3 (N7241, N7227, N1970, N3869);
xor XOR2 (N7242, N7226, N3038);
and AND2 (N7243, N7237, N5828);
nand NAND4 (N7244, N7240, N2364, N5953, N5132);
and AND2 (N7245, N7242, N6115);
buf BUF1 (N7246, N7243);
xor XOR2 (N7247, N7239, N3665);
xor XOR2 (N7248, N7216, N3962);
buf BUF1 (N7249, N7248);
nor NOR4 (N7250, N7234, N7118, N6193, N2122);
buf BUF1 (N7251, N7247);
and AND3 (N7252, N7241, N4731, N5182);
nand NAND2 (N7253, N7250, N1756);
nand NAND3 (N7254, N7251, N1626, N1755);
xor XOR2 (N7255, N7249, N3042);
xor XOR2 (N7256, N7246, N2876);
xor XOR2 (N7257, N7254, N4423);
or OR2 (N7258, N7252, N5445);
not NOT1 (N7259, N7245);
and AND2 (N7260, N7238, N3436);
not NOT1 (N7261, N7256);
nor NOR2 (N7262, N7259, N4764);
nand NAND3 (N7263, N7218, N1534, N4588);
nand NAND2 (N7264, N7244, N5038);
and AND4 (N7265, N7213, N597, N5159, N2690);
or OR3 (N7266, N7261, N934, N4083);
or OR4 (N7267, N7263, N5969, N793, N1272);
xor XOR2 (N7268, N7267, N3138);
nand NAND2 (N7269, N7262, N855);
not NOT1 (N7270, N7253);
not NOT1 (N7271, N7269);
nand NAND4 (N7272, N7264, N1747, N6937, N4244);
and AND2 (N7273, N7265, N2485);
and AND3 (N7274, N7268, N3758, N4081);
and AND2 (N7275, N7255, N4890);
nand NAND4 (N7276, N7266, N5998, N4309, N5255);
and AND3 (N7277, N7276, N2229, N5532);
nand NAND2 (N7278, N7275, N1725);
nor NOR4 (N7279, N7278, N3314, N2130, N4851);
nand NAND2 (N7280, N7258, N5846);
nand NAND2 (N7281, N7257, N891);
nand NAND3 (N7282, N7273, N2531, N6609);
nor NOR2 (N7283, N7280, N3059);
xor XOR2 (N7284, N7274, N2949);
xor XOR2 (N7285, N7272, N3235);
not NOT1 (N7286, N7271);
xor XOR2 (N7287, N7279, N5332);
not NOT1 (N7288, N7285);
not NOT1 (N7289, N7286);
or OR2 (N7290, N7277, N3173);
xor XOR2 (N7291, N7260, N4560);
buf BUF1 (N7292, N7281);
or OR2 (N7293, N7282, N6634);
and AND2 (N7294, N7270, N2935);
buf BUF1 (N7295, N7287);
not NOT1 (N7296, N7293);
not NOT1 (N7297, N7292);
nor NOR4 (N7298, N7289, N6655, N4479, N1278);
buf BUF1 (N7299, N7291);
nor NOR2 (N7300, N7294, N5591);
nor NOR2 (N7301, N7299, N4713);
or OR3 (N7302, N7283, N1210, N2604);
and AND2 (N7303, N7300, N1614);
and AND4 (N7304, N7284, N6467, N413, N1718);
buf BUF1 (N7305, N7290);
not NOT1 (N7306, N7304);
and AND4 (N7307, N7303, N260, N591, N505);
buf BUF1 (N7308, N7295);
buf BUF1 (N7309, N7301);
xor XOR2 (N7310, N7307, N55);
xor XOR2 (N7311, N7298, N4817);
not NOT1 (N7312, N7296);
buf BUF1 (N7313, N7306);
not NOT1 (N7314, N7297);
buf BUF1 (N7315, N7305);
nand NAND2 (N7316, N7311, N494);
xor XOR2 (N7317, N7314, N3039);
xor XOR2 (N7318, N7309, N411);
or OR3 (N7319, N7310, N2494, N906);
not NOT1 (N7320, N7318);
or OR3 (N7321, N7315, N2151, N2821);
nand NAND2 (N7322, N7316, N109);
and AND4 (N7323, N7302, N5777, N4719, N3945);
buf BUF1 (N7324, N7288);
nor NOR3 (N7325, N7320, N4392, N3176);
buf BUF1 (N7326, N7308);
xor XOR2 (N7327, N7325, N1991);
nand NAND3 (N7328, N7326, N6957, N4351);
or OR3 (N7329, N7327, N1199, N5723);
nor NOR3 (N7330, N7322, N2178, N7210);
and AND3 (N7331, N7323, N6391, N5478);
buf BUF1 (N7332, N7313);
nor NOR2 (N7333, N7324, N3278);
nand NAND3 (N7334, N7330, N3490, N2405);
nand NAND3 (N7335, N7329, N1529, N670);
xor XOR2 (N7336, N7319, N2114);
nor NOR4 (N7337, N7317, N3289, N3971, N7);
nor NOR4 (N7338, N7334, N1127, N4318, N390);
nor NOR3 (N7339, N7321, N5019, N6153);
or OR3 (N7340, N7339, N6745, N2014);
and AND4 (N7341, N7331, N2559, N4922, N4802);
not NOT1 (N7342, N7333);
xor XOR2 (N7343, N7341, N5206);
and AND4 (N7344, N7332, N29, N3665, N2984);
and AND2 (N7345, N7344, N2406);
or OR2 (N7346, N7342, N5528);
nand NAND4 (N7347, N7345, N6053, N5373, N578);
nand NAND4 (N7348, N7347, N6704, N1124, N6819);
and AND4 (N7349, N7340, N3286, N105, N974);
or OR3 (N7350, N7335, N283, N270);
and AND3 (N7351, N7337, N852, N2348);
buf BUF1 (N7352, N7346);
nand NAND4 (N7353, N7312, N5585, N1076, N5552);
nand NAND2 (N7354, N7343, N2554);
xor XOR2 (N7355, N7338, N834);
xor XOR2 (N7356, N7351, N2221);
and AND3 (N7357, N7353, N3562, N5767);
buf BUF1 (N7358, N7350);
not NOT1 (N7359, N7357);
nand NAND4 (N7360, N7358, N6547, N7316, N7261);
xor XOR2 (N7361, N7336, N3408);
buf BUF1 (N7362, N7360);
buf BUF1 (N7363, N7349);
and AND2 (N7364, N7348, N3757);
buf BUF1 (N7365, N7356);
nor NOR3 (N7366, N7362, N56, N3859);
nor NOR2 (N7367, N7364, N6087);
buf BUF1 (N7368, N7365);
or OR4 (N7369, N7361, N2755, N780, N4818);
buf BUF1 (N7370, N7367);
not NOT1 (N7371, N7368);
not NOT1 (N7372, N7354);
and AND2 (N7373, N7366, N2777);
buf BUF1 (N7374, N7369);
not NOT1 (N7375, N7352);
nand NAND2 (N7376, N7373, N1600);
nor NOR2 (N7377, N7374, N6581);
nand NAND2 (N7378, N7355, N4657);
nand NAND2 (N7379, N7375, N3491);
or OR3 (N7380, N7359, N6084, N407);
xor XOR2 (N7381, N7370, N4729);
or OR3 (N7382, N7376, N5033, N6539);
and AND2 (N7383, N7378, N3692);
not NOT1 (N7384, N7383);
and AND2 (N7385, N7377, N2698);
and AND3 (N7386, N7384, N269, N6990);
and AND3 (N7387, N7381, N3088, N1841);
nor NOR2 (N7388, N7385, N1072);
nand NAND4 (N7389, N7371, N6369, N3456, N2481);
buf BUF1 (N7390, N7379);
not NOT1 (N7391, N7386);
or OR4 (N7392, N7387, N1327, N6919, N3092);
not NOT1 (N7393, N7380);
nor NOR4 (N7394, N7389, N723, N3624, N81);
buf BUF1 (N7395, N7363);
and AND4 (N7396, N7391, N91, N4991, N3116);
buf BUF1 (N7397, N7396);
nand NAND3 (N7398, N7388, N5223, N4072);
not NOT1 (N7399, N7394);
nor NOR2 (N7400, N7328, N2431);
buf BUF1 (N7401, N7395);
xor XOR2 (N7402, N7397, N1513);
or OR2 (N7403, N7390, N784);
buf BUF1 (N7404, N7403);
xor XOR2 (N7405, N7404, N5245);
and AND2 (N7406, N7392, N970);
not NOT1 (N7407, N7372);
buf BUF1 (N7408, N7382);
buf BUF1 (N7409, N7405);
nand NAND3 (N7410, N7408, N6595, N348);
buf BUF1 (N7411, N7407);
not NOT1 (N7412, N7398);
not NOT1 (N7413, N7402);
xor XOR2 (N7414, N7393, N7037);
buf BUF1 (N7415, N7401);
nor NOR2 (N7416, N7410, N3416);
or OR4 (N7417, N7406, N6062, N6485, N6893);
xor XOR2 (N7418, N7400, N4934);
not NOT1 (N7419, N7412);
nor NOR2 (N7420, N7411, N6932);
nand NAND3 (N7421, N7420, N6189, N1262);
and AND3 (N7422, N7409, N1883, N5903);
xor XOR2 (N7423, N7413, N1989);
and AND3 (N7424, N7418, N895, N7375);
or OR4 (N7425, N7415, N2036, N1870, N658);
and AND3 (N7426, N7399, N7242, N3252);
buf BUF1 (N7427, N7422);
xor XOR2 (N7428, N7414, N3095);
not NOT1 (N7429, N7424);
and AND2 (N7430, N7416, N2333);
or OR3 (N7431, N7423, N2210, N2017);
buf BUF1 (N7432, N7430);
or OR4 (N7433, N7426, N4189, N4661, N4289);
nand NAND3 (N7434, N7431, N3886, N24);
and AND3 (N7435, N7433, N1276, N3612);
or OR4 (N7436, N7434, N74, N6937, N1969);
xor XOR2 (N7437, N7436, N118);
and AND2 (N7438, N7428, N5065);
nor NOR2 (N7439, N7435, N3738);
xor XOR2 (N7440, N7432, N1391);
buf BUF1 (N7441, N7429);
or OR2 (N7442, N7438, N2085);
xor XOR2 (N7443, N7441, N1795);
xor XOR2 (N7444, N7425, N6189);
and AND2 (N7445, N7439, N4048);
or OR4 (N7446, N7421, N7348, N6793, N1171);
nor NOR4 (N7447, N7443, N3104, N4069, N4608);
not NOT1 (N7448, N7446);
and AND4 (N7449, N7448, N3683, N3793, N2927);
and AND4 (N7450, N7449, N2640, N2642, N3171);
and AND4 (N7451, N7417, N3130, N5496, N1078);
xor XOR2 (N7452, N7440, N4502);
not NOT1 (N7453, N7442);
xor XOR2 (N7454, N7452, N6594);
not NOT1 (N7455, N7419);
xor XOR2 (N7456, N7444, N6251);
buf BUF1 (N7457, N7455);
or OR2 (N7458, N7454, N6687);
or OR4 (N7459, N7457, N4141, N5318, N6160);
or OR4 (N7460, N7458, N7203, N6525, N3949);
xor XOR2 (N7461, N7427, N6450);
nand NAND2 (N7462, N7447, N513);
and AND3 (N7463, N7462, N5392, N2067);
and AND4 (N7464, N7456, N7397, N2575, N385);
and AND4 (N7465, N7445, N3687, N3418, N327);
nor NOR4 (N7466, N7465, N6590, N532, N1871);
or OR4 (N7467, N7437, N6374, N789, N1344);
buf BUF1 (N7468, N7463);
not NOT1 (N7469, N7453);
not NOT1 (N7470, N7464);
buf BUF1 (N7471, N7467);
nand NAND3 (N7472, N7469, N3785, N4297);
nor NOR4 (N7473, N7468, N538, N6013, N1242);
nand NAND3 (N7474, N7470, N5223, N3947);
buf BUF1 (N7475, N7471);
not NOT1 (N7476, N7461);
or OR4 (N7477, N7475, N6887, N3100, N4241);
and AND4 (N7478, N7451, N3561, N6943, N1159);
buf BUF1 (N7479, N7460);
buf BUF1 (N7480, N7473);
xor XOR2 (N7481, N7472, N2342);
buf BUF1 (N7482, N7476);
or OR4 (N7483, N7466, N5873, N4876, N437);
and AND2 (N7484, N7478, N1226);
buf BUF1 (N7485, N7482);
and AND2 (N7486, N7484, N7218);
nand NAND4 (N7487, N7481, N348, N1946, N5253);
not NOT1 (N7488, N7474);
or OR3 (N7489, N7459, N5363, N5020);
or OR3 (N7490, N7485, N1213, N2600);
or OR4 (N7491, N7479, N848, N2547, N4955);
or OR2 (N7492, N7486, N3405);
xor XOR2 (N7493, N7480, N1120);
not NOT1 (N7494, N7490);
nor NOR3 (N7495, N7493, N7178, N5560);
and AND4 (N7496, N7488, N452, N6935, N3089);
nor NOR3 (N7497, N7477, N3542, N3184);
or OR3 (N7498, N7492, N3273, N3624);
or OR3 (N7499, N7489, N6753, N3212);
nand NAND3 (N7500, N7491, N3591, N2249);
nand NAND3 (N7501, N7499, N6557, N4277);
nor NOR3 (N7502, N7495, N7132, N4055);
and AND2 (N7503, N7494, N6119);
xor XOR2 (N7504, N7483, N1120);
nor NOR2 (N7505, N7450, N7308);
and AND3 (N7506, N7487, N67, N6245);
xor XOR2 (N7507, N7501, N6803);
xor XOR2 (N7508, N7504, N4358);
nor NOR2 (N7509, N7505, N1494);
buf BUF1 (N7510, N7497);
and AND4 (N7511, N7507, N5920, N1462, N1213);
xor XOR2 (N7512, N7496, N2003);
not NOT1 (N7513, N7502);
nand NAND2 (N7514, N7509, N4656);
and AND2 (N7515, N7503, N1366);
nand NAND4 (N7516, N7500, N2074, N1303, N5225);
xor XOR2 (N7517, N7514, N2630);
not NOT1 (N7518, N7506);
or OR2 (N7519, N7513, N7015);
buf BUF1 (N7520, N7508);
not NOT1 (N7521, N7520);
and AND2 (N7522, N7516, N3260);
or OR2 (N7523, N7522, N7201);
nand NAND2 (N7524, N7521, N6676);
not NOT1 (N7525, N7517);
buf BUF1 (N7526, N7498);
not NOT1 (N7527, N7510);
buf BUF1 (N7528, N7525);
buf BUF1 (N7529, N7518);
nand NAND4 (N7530, N7529, N2307, N7457, N6060);
buf BUF1 (N7531, N7527);
and AND3 (N7532, N7515, N2076, N7322);
xor XOR2 (N7533, N7528, N133);
nor NOR3 (N7534, N7532, N6450, N2922);
xor XOR2 (N7535, N7531, N3447);
nand NAND4 (N7536, N7534, N1075, N176, N5133);
nand NAND2 (N7537, N7519, N4100);
and AND2 (N7538, N7512, N6677);
and AND3 (N7539, N7511, N2691, N1097);
and AND2 (N7540, N7537, N558);
or OR2 (N7541, N7540, N4701);
and AND4 (N7542, N7523, N4715, N7034, N3601);
nand NAND3 (N7543, N7526, N3386, N4853);
nor NOR4 (N7544, N7538, N4644, N2411, N4590);
and AND4 (N7545, N7530, N2588, N6552, N7264);
buf BUF1 (N7546, N7539);
buf BUF1 (N7547, N7541);
and AND2 (N7548, N7542, N6237);
or OR2 (N7549, N7524, N4167);
nor NOR2 (N7550, N7544, N6308);
or OR4 (N7551, N7550, N4576, N2823, N4453);
not NOT1 (N7552, N7548);
and AND4 (N7553, N7543, N4337, N5072, N6751);
nor NOR2 (N7554, N7533, N5274);
buf BUF1 (N7555, N7547);
or OR2 (N7556, N7553, N2947);
nor NOR3 (N7557, N7536, N1016, N2287);
and AND2 (N7558, N7557, N7440);
and AND3 (N7559, N7555, N1976, N4162);
buf BUF1 (N7560, N7545);
and AND3 (N7561, N7535, N5768, N1756);
nand NAND3 (N7562, N7551, N6141, N7092);
not NOT1 (N7563, N7558);
and AND2 (N7564, N7549, N1520);
and AND3 (N7565, N7556, N2590, N2783);
and AND4 (N7566, N7554, N1901, N7551, N629);
nor NOR4 (N7567, N7563, N819, N4393, N1756);
nand NAND4 (N7568, N7566, N2516, N1479, N1104);
or OR4 (N7569, N7568, N7532, N5674, N7083);
nor NOR2 (N7570, N7560, N309);
nor NOR2 (N7571, N7546, N2205);
buf BUF1 (N7572, N7567);
not NOT1 (N7573, N7570);
and AND2 (N7574, N7569, N2878);
nor NOR4 (N7575, N7572, N6339, N757, N4096);
nand NAND4 (N7576, N7571, N1624, N4574, N3127);
not NOT1 (N7577, N7559);
and AND2 (N7578, N7564, N5650);
not NOT1 (N7579, N7561);
or OR3 (N7580, N7576, N3779, N395);
not NOT1 (N7581, N7579);
and AND3 (N7582, N7575, N2862, N1868);
or OR3 (N7583, N7577, N6439, N5973);
not NOT1 (N7584, N7562);
nand NAND4 (N7585, N7578, N6521, N484, N6843);
buf BUF1 (N7586, N7573);
nor NOR3 (N7587, N7582, N5998, N2214);
nor NOR4 (N7588, N7552, N3437, N3145, N5445);
nand NAND2 (N7589, N7588, N336);
not NOT1 (N7590, N7574);
not NOT1 (N7591, N7585);
and AND2 (N7592, N7584, N7347);
and AND4 (N7593, N7565, N1536, N7008, N5473);
buf BUF1 (N7594, N7592);
or OR4 (N7595, N7593, N4565, N4633, N1599);
and AND3 (N7596, N7580, N2253, N214);
nand NAND4 (N7597, N7594, N4224, N5471, N4815);
nor NOR3 (N7598, N7596, N4157, N1182);
nor NOR3 (N7599, N7587, N3071, N4682);
not NOT1 (N7600, N7591);
xor XOR2 (N7601, N7583, N1450);
xor XOR2 (N7602, N7586, N3937);
buf BUF1 (N7603, N7601);
and AND3 (N7604, N7598, N139, N1516);
or OR4 (N7605, N7603, N3849, N6608, N5440);
nor NOR3 (N7606, N7599, N2988, N3410);
buf BUF1 (N7607, N7604);
and AND2 (N7608, N7600, N2237);
nand NAND3 (N7609, N7589, N7225, N3318);
and AND2 (N7610, N7609, N6844);
or OR2 (N7611, N7590, N2415);
not NOT1 (N7612, N7602);
and AND3 (N7613, N7605, N6448, N3140);
nor NOR3 (N7614, N7612, N6916, N3027);
xor XOR2 (N7615, N7610, N5114);
xor XOR2 (N7616, N7615, N7378);
xor XOR2 (N7617, N7595, N143);
or OR4 (N7618, N7614, N4997, N3388, N837);
or OR4 (N7619, N7608, N5327, N259, N3433);
and AND2 (N7620, N7597, N6614);
nand NAND4 (N7621, N7617, N838, N3536, N6395);
not NOT1 (N7622, N7618);
nor NOR2 (N7623, N7616, N438);
nor NOR4 (N7624, N7620, N2640, N6596, N1957);
not NOT1 (N7625, N7613);
xor XOR2 (N7626, N7607, N3772);
nand NAND4 (N7627, N7622, N7287, N1129, N5397);
and AND3 (N7628, N7611, N3709, N1694);
nand NAND2 (N7629, N7628, N1495);
nand NAND2 (N7630, N7581, N803);
nand NAND4 (N7631, N7606, N2259, N4953, N5816);
and AND2 (N7632, N7626, N2093);
or OR4 (N7633, N7631, N6817, N4047, N1752);
and AND2 (N7634, N7624, N645);
buf BUF1 (N7635, N7633);
xor XOR2 (N7636, N7635, N5879);
or OR3 (N7637, N7630, N2431, N7317);
xor XOR2 (N7638, N7634, N7194);
nor NOR2 (N7639, N7637, N6029);
nand NAND3 (N7640, N7636, N2847, N7076);
or OR3 (N7641, N7632, N3458, N370);
and AND4 (N7642, N7640, N1416, N3229, N1369);
nand NAND4 (N7643, N7642, N1607, N4953, N6279);
xor XOR2 (N7644, N7638, N2531);
nand NAND3 (N7645, N7623, N1214, N2670);
not NOT1 (N7646, N7639);
nand NAND3 (N7647, N7625, N4102, N1204);
buf BUF1 (N7648, N7641);
xor XOR2 (N7649, N7646, N5877);
nand NAND3 (N7650, N7629, N4189, N6457);
or OR3 (N7651, N7619, N5866, N1278);
or OR2 (N7652, N7645, N775);
nand NAND2 (N7653, N7648, N1149);
buf BUF1 (N7654, N7652);
buf BUF1 (N7655, N7649);
and AND3 (N7656, N7644, N7266, N6542);
nand NAND2 (N7657, N7643, N7199);
and AND2 (N7658, N7653, N4414);
not NOT1 (N7659, N7651);
xor XOR2 (N7660, N7656, N6654);
and AND4 (N7661, N7654, N2500, N977, N6938);
or OR3 (N7662, N7627, N2012, N1784);
xor XOR2 (N7663, N7661, N1452);
buf BUF1 (N7664, N7621);
and AND4 (N7665, N7663, N1778, N7274, N1858);
xor XOR2 (N7666, N7650, N4055);
buf BUF1 (N7667, N7660);
nand NAND2 (N7668, N7659, N2309);
xor XOR2 (N7669, N7662, N2728);
and AND3 (N7670, N7667, N6667, N4796);
xor XOR2 (N7671, N7664, N2400);
and AND3 (N7672, N7658, N2535, N6823);
nor NOR3 (N7673, N7671, N2748, N1218);
not NOT1 (N7674, N7666);
nor NOR2 (N7675, N7665, N1925);
and AND4 (N7676, N7672, N54, N3175, N3900);
or OR2 (N7677, N7675, N5337);
buf BUF1 (N7678, N7669);
nor NOR4 (N7679, N7657, N7518, N2852, N5912);
or OR4 (N7680, N7678, N4952, N5267, N6766);
xor XOR2 (N7681, N7647, N3042);
and AND4 (N7682, N7681, N4074, N3227, N2446);
and AND3 (N7683, N7682, N6066, N786);
nand NAND2 (N7684, N7655, N3498);
buf BUF1 (N7685, N7683);
and AND2 (N7686, N7674, N4003);
not NOT1 (N7687, N7679);
and AND4 (N7688, N7686, N4747, N5671, N292);
nand NAND2 (N7689, N7673, N1870);
not NOT1 (N7690, N7689);
nor NOR3 (N7691, N7668, N5020, N4098);
buf BUF1 (N7692, N7670);
nor NOR3 (N7693, N7688, N5055, N2584);
xor XOR2 (N7694, N7693, N6562);
nand NAND2 (N7695, N7691, N2822);
or OR4 (N7696, N7690, N2929, N4202, N3502);
nor NOR4 (N7697, N7680, N7215, N5903, N4507);
nor NOR3 (N7698, N7687, N4367, N823);
nor NOR2 (N7699, N7695, N750);
and AND2 (N7700, N7685, N3973);
or OR2 (N7701, N7694, N4372);
buf BUF1 (N7702, N7676);
and AND4 (N7703, N7700, N5417, N4605, N1444);
nor NOR4 (N7704, N7692, N2591, N556, N3965);
xor XOR2 (N7705, N7697, N3186);
xor XOR2 (N7706, N7704, N923);
nor NOR3 (N7707, N7703, N5317, N6745);
nor NOR4 (N7708, N7702, N2224, N7371, N1544);
xor XOR2 (N7709, N7701, N1127);
xor XOR2 (N7710, N7708, N2053);
nor NOR3 (N7711, N7698, N195, N7107);
and AND2 (N7712, N7711, N1001);
not NOT1 (N7713, N7699);
not NOT1 (N7714, N7696);
not NOT1 (N7715, N7684);
nand NAND3 (N7716, N7715, N3709, N6292);
buf BUF1 (N7717, N7709);
or OR2 (N7718, N7705, N6748);
nand NAND4 (N7719, N7712, N3411, N163, N305);
nand NAND3 (N7720, N7717, N4055, N3740);
not NOT1 (N7721, N7716);
xor XOR2 (N7722, N7707, N2767);
and AND4 (N7723, N7718, N7479, N1910, N1922);
and AND2 (N7724, N7721, N6772);
nor NOR3 (N7725, N7723, N6872, N5473);
or OR4 (N7726, N7713, N2, N5069, N4472);
nand NAND4 (N7727, N7722, N590, N1652, N6691);
nand NAND2 (N7728, N7724, N4172);
or OR2 (N7729, N7727, N462);
xor XOR2 (N7730, N7728, N5651);
nand NAND3 (N7731, N7706, N1929, N531);
buf BUF1 (N7732, N7731);
and AND3 (N7733, N7720, N3706, N615);
xor XOR2 (N7734, N7726, N1215);
buf BUF1 (N7735, N7714);
not NOT1 (N7736, N7733);
nor NOR3 (N7737, N7732, N3539, N1117);
or OR2 (N7738, N7735, N7202);
not NOT1 (N7739, N7677);
and AND2 (N7740, N7725, N4085);
nor NOR4 (N7741, N7738, N7441, N287, N4317);
nand NAND2 (N7742, N7734, N3386);
and AND2 (N7743, N7741, N876);
xor XOR2 (N7744, N7736, N1237);
or OR2 (N7745, N7740, N3376);
not NOT1 (N7746, N7729);
buf BUF1 (N7747, N7737);
buf BUF1 (N7748, N7744);
buf BUF1 (N7749, N7719);
buf BUF1 (N7750, N7749);
not NOT1 (N7751, N7710);
not NOT1 (N7752, N7745);
not NOT1 (N7753, N7742);
buf BUF1 (N7754, N7753);
buf BUF1 (N7755, N7754);
not NOT1 (N7756, N7751);
xor XOR2 (N7757, N7750, N364);
or OR2 (N7758, N7752, N2434);
nand NAND4 (N7759, N7756, N3376, N1278, N7086);
buf BUF1 (N7760, N7755);
xor XOR2 (N7761, N7748, N3734);
xor XOR2 (N7762, N7739, N1902);
xor XOR2 (N7763, N7759, N2815);
not NOT1 (N7764, N7760);
not NOT1 (N7765, N7757);
buf BUF1 (N7766, N7743);
buf BUF1 (N7767, N7762);
nand NAND3 (N7768, N7747, N6895, N1642);
xor XOR2 (N7769, N7768, N3369);
nand NAND2 (N7770, N7746, N644);
nor NOR3 (N7771, N7761, N2659, N6651);
xor XOR2 (N7772, N7771, N6322);
not NOT1 (N7773, N7767);
nand NAND3 (N7774, N7770, N1810, N5058);
not NOT1 (N7775, N7772);
not NOT1 (N7776, N7769);
nor NOR4 (N7777, N7730, N797, N4482, N7487);
xor XOR2 (N7778, N7763, N2043);
and AND4 (N7779, N7765, N3801, N3989, N7655);
nand NAND4 (N7780, N7776, N7338, N3381, N800);
xor XOR2 (N7781, N7778, N7126);
buf BUF1 (N7782, N7781);
nand NAND3 (N7783, N7773, N5446, N4024);
not NOT1 (N7784, N7774);
and AND2 (N7785, N7780, N4770);
buf BUF1 (N7786, N7764);
or OR3 (N7787, N7782, N3925, N168);
buf BUF1 (N7788, N7785);
nand NAND4 (N7789, N7784, N3004, N3012, N1559);
nand NAND3 (N7790, N7758, N5653, N4417);
nor NOR3 (N7791, N7786, N4884, N2638);
and AND3 (N7792, N7789, N5932, N4202);
buf BUF1 (N7793, N7779);
xor XOR2 (N7794, N7790, N5055);
xor XOR2 (N7795, N7794, N529);
xor XOR2 (N7796, N7777, N7757);
nor NOR2 (N7797, N7788, N6535);
or OR3 (N7798, N7791, N2032, N2805);
or OR3 (N7799, N7793, N2043, N6024);
or OR3 (N7800, N7799, N5979, N1454);
or OR4 (N7801, N7783, N6610, N5775, N3593);
xor XOR2 (N7802, N7797, N5089);
xor XOR2 (N7803, N7792, N5021);
not NOT1 (N7804, N7775);
not NOT1 (N7805, N7800);
xor XOR2 (N7806, N7805, N5216);
xor XOR2 (N7807, N7806, N5310);
xor XOR2 (N7808, N7807, N1869);
and AND3 (N7809, N7808, N5041, N2126);
not NOT1 (N7810, N7787);
buf BUF1 (N7811, N7801);
or OR2 (N7812, N7766, N2274);
nand NAND4 (N7813, N7809, N7624, N938, N6246);
nor NOR4 (N7814, N7796, N2247, N4941, N3358);
not NOT1 (N7815, N7795);
nand NAND2 (N7816, N7815, N2867);
or OR3 (N7817, N7813, N2308, N3310);
nand NAND4 (N7818, N7810, N5806, N6210, N3229);
xor XOR2 (N7819, N7817, N7290);
or OR2 (N7820, N7802, N2787);
buf BUF1 (N7821, N7804);
nor NOR3 (N7822, N7798, N5598, N3739);
and AND2 (N7823, N7822, N2350);
or OR2 (N7824, N7821, N5512);
nand NAND2 (N7825, N7816, N7533);
nor NOR2 (N7826, N7820, N4417);
nor NOR3 (N7827, N7818, N1498, N5390);
xor XOR2 (N7828, N7819, N6898);
nor NOR4 (N7829, N7812, N7756, N5876, N7017);
not NOT1 (N7830, N7829);
xor XOR2 (N7831, N7824, N2114);
xor XOR2 (N7832, N7830, N7078);
or OR4 (N7833, N7831, N6037, N2059, N750);
not NOT1 (N7834, N7832);
and AND4 (N7835, N7834, N1258, N4606, N5608);
nor NOR4 (N7836, N7803, N3492, N53, N4918);
xor XOR2 (N7837, N7825, N2210);
xor XOR2 (N7838, N7836, N141);
nand NAND2 (N7839, N7811, N1612);
nor NOR4 (N7840, N7838, N5769, N6218, N1236);
buf BUF1 (N7841, N7835);
nand NAND3 (N7842, N7827, N2158, N6699);
or OR4 (N7843, N7842, N7787, N2307, N370);
nor NOR2 (N7844, N7826, N1751);
not NOT1 (N7845, N7839);
xor XOR2 (N7846, N7837, N7361);
nor NOR2 (N7847, N7833, N6410);
and AND2 (N7848, N7814, N4731);
or OR3 (N7849, N7847, N4691, N284);
nor NOR3 (N7850, N7848, N7086, N5566);
buf BUF1 (N7851, N7828);
not NOT1 (N7852, N7841);
not NOT1 (N7853, N7844);
and AND3 (N7854, N7851, N1772, N5740);
nand NAND4 (N7855, N7852, N997, N7468, N7161);
xor XOR2 (N7856, N7853, N458);
nor NOR4 (N7857, N7854, N4149, N3030, N4996);
not NOT1 (N7858, N7856);
nand NAND4 (N7859, N7850, N3721, N3728, N7318);
not NOT1 (N7860, N7823);
and AND3 (N7861, N7859, N5526, N1622);
buf BUF1 (N7862, N7843);
or OR4 (N7863, N7849, N879, N6118, N4075);
xor XOR2 (N7864, N7861, N1728);
buf BUF1 (N7865, N7864);
nor NOR3 (N7866, N7862, N859, N3591);
buf BUF1 (N7867, N7858);
or OR2 (N7868, N7866, N1642);
and AND3 (N7869, N7863, N2514, N7096);
not NOT1 (N7870, N7865);
nor NOR4 (N7871, N7845, N4715, N5025, N6314);
buf BUF1 (N7872, N7860);
not NOT1 (N7873, N7869);
nand NAND2 (N7874, N7846, N2273);
xor XOR2 (N7875, N7840, N1133);
buf BUF1 (N7876, N7874);
not NOT1 (N7877, N7868);
xor XOR2 (N7878, N7867, N3056);
not NOT1 (N7879, N7877);
not NOT1 (N7880, N7879);
xor XOR2 (N7881, N7873, N3219);
xor XOR2 (N7882, N7881, N4240);
or OR3 (N7883, N7871, N456, N6569);
nor NOR3 (N7884, N7878, N3339, N1051);
buf BUF1 (N7885, N7880);
or OR3 (N7886, N7857, N4359, N6555);
or OR4 (N7887, N7875, N5196, N4768, N7430);
xor XOR2 (N7888, N7886, N3841);
nand NAND2 (N7889, N7885, N3444);
nand NAND3 (N7890, N7888, N6754, N4786);
or OR2 (N7891, N7889, N2360);
nor NOR3 (N7892, N7883, N3504, N1701);
or OR2 (N7893, N7876, N2433);
nor NOR3 (N7894, N7890, N3393, N5135);
and AND3 (N7895, N7882, N2407, N4595);
buf BUF1 (N7896, N7895);
and AND2 (N7897, N7870, N3634);
buf BUF1 (N7898, N7872);
and AND3 (N7899, N7891, N6226, N3159);
not NOT1 (N7900, N7894);
nand NAND2 (N7901, N7855, N631);
not NOT1 (N7902, N7884);
not NOT1 (N7903, N7897);
and AND2 (N7904, N7896, N2835);
nor NOR4 (N7905, N7893, N44, N4496, N790);
or OR4 (N7906, N7903, N989, N7364, N2531);
and AND2 (N7907, N7892, N2619);
or OR3 (N7908, N7902, N2227, N1082);
nor NOR3 (N7909, N7906, N1046, N383);
xor XOR2 (N7910, N7887, N4730);
or OR4 (N7911, N7900, N6149, N666, N7165);
nor NOR3 (N7912, N7901, N6671, N1063);
not NOT1 (N7913, N7908);
nor NOR4 (N7914, N7905, N5255, N7329, N6383);
nand NAND4 (N7915, N7904, N6088, N6748, N2524);
and AND2 (N7916, N7913, N2465);
nor NOR4 (N7917, N7910, N4117, N3219, N1033);
xor XOR2 (N7918, N7898, N515);
and AND3 (N7919, N7899, N5082, N2404);
buf BUF1 (N7920, N7907);
or OR3 (N7921, N7918, N3994, N4574);
or OR3 (N7922, N7919, N5565, N7108);
nand NAND2 (N7923, N7915, N6924);
not NOT1 (N7924, N7909);
not NOT1 (N7925, N7921);
nor NOR4 (N7926, N7920, N3090, N4178, N563);
nand NAND3 (N7927, N7926, N3520, N4819);
nand NAND2 (N7928, N7917, N5974);
buf BUF1 (N7929, N7928);
buf BUF1 (N7930, N7911);
not NOT1 (N7931, N7930);
nand NAND4 (N7932, N7922, N4203, N3340, N3171);
and AND2 (N7933, N7931, N12);
and AND4 (N7934, N7924, N6829, N1560, N2146);
nand NAND3 (N7935, N7929, N4006, N6296);
not NOT1 (N7936, N7914);
buf BUF1 (N7937, N7935);
nor NOR2 (N7938, N7923, N1143);
not NOT1 (N7939, N7925);
nand NAND2 (N7940, N7937, N7052);
and AND2 (N7941, N7912, N317);
nand NAND4 (N7942, N7933, N3798, N2022, N5985);
nand NAND4 (N7943, N7934, N4575, N1673, N6843);
and AND4 (N7944, N7938, N6737, N7711, N7663);
and AND3 (N7945, N7943, N5410, N5725);
xor XOR2 (N7946, N7936, N3600);
not NOT1 (N7947, N7944);
not NOT1 (N7948, N7939);
and AND3 (N7949, N7940, N5364, N707);
nor NOR4 (N7950, N7927, N4209, N7773, N1279);
and AND4 (N7951, N7942, N6133, N7023, N341);
and AND3 (N7952, N7949, N432, N3863);
not NOT1 (N7953, N7916);
buf BUF1 (N7954, N7945);
xor XOR2 (N7955, N7953, N6643);
and AND4 (N7956, N7947, N4951, N7174, N7367);
nand NAND3 (N7957, N7946, N7313, N1251);
nor NOR4 (N7958, N7955, N4845, N5778, N3439);
nand NAND3 (N7959, N7956, N3322, N7502);
nor NOR4 (N7960, N7958, N6407, N7017, N572);
nor NOR3 (N7961, N7950, N6982, N6799);
nand NAND3 (N7962, N7954, N5214, N3067);
and AND2 (N7963, N7960, N113);
or OR3 (N7964, N7952, N1065, N6797);
buf BUF1 (N7965, N7941);
not NOT1 (N7966, N7965);
and AND2 (N7967, N7957, N1468);
nor NOR3 (N7968, N7961, N5167, N6316);
xor XOR2 (N7969, N7948, N6420);
or OR2 (N7970, N7959, N244);
buf BUF1 (N7971, N7970);
xor XOR2 (N7972, N7966, N7519);
not NOT1 (N7973, N7964);
buf BUF1 (N7974, N7951);
nor NOR4 (N7975, N7968, N53, N5818, N2989);
or OR2 (N7976, N7974, N3418);
buf BUF1 (N7977, N7971);
or OR4 (N7978, N7932, N4782, N5427, N5147);
xor XOR2 (N7979, N7976, N6307);
not NOT1 (N7980, N7973);
nand NAND3 (N7981, N7963, N3256, N6598);
xor XOR2 (N7982, N7981, N5671);
and AND2 (N7983, N7979, N812);
or OR2 (N7984, N7983, N659);
nor NOR2 (N7985, N7978, N1119);
buf BUF1 (N7986, N7984);
or OR3 (N7987, N7969, N3056, N6051);
not NOT1 (N7988, N7985);
buf BUF1 (N7989, N7980);
nand NAND4 (N7990, N7982, N7630, N3101, N5795);
nand NAND2 (N7991, N7975, N6699);
xor XOR2 (N7992, N7989, N6988);
or OR2 (N7993, N7962, N667);
nor NOR2 (N7994, N7992, N3403);
or OR2 (N7995, N7991, N6081);
nand NAND3 (N7996, N7993, N5440, N7041);
nand NAND4 (N7997, N7967, N755, N6494, N1245);
not NOT1 (N7998, N7986);
buf BUF1 (N7999, N7995);
nand NAND3 (N8000, N7972, N1209, N3404);
nor NOR4 (N8001, N7988, N6168, N7268, N1045);
nand NAND3 (N8002, N7977, N5905, N2629);
not NOT1 (N8003, N7987);
not NOT1 (N8004, N8001);
buf BUF1 (N8005, N7999);
or OR2 (N8006, N7994, N1825);
xor XOR2 (N8007, N7997, N745);
not NOT1 (N8008, N8006);
or OR2 (N8009, N8002, N379);
xor XOR2 (N8010, N8003, N3009);
or OR2 (N8011, N8005, N4871);
buf BUF1 (N8012, N7998);
nand NAND3 (N8013, N7996, N3335, N4025);
buf BUF1 (N8014, N8008);
nand NAND3 (N8015, N8011, N5393, N318);
nand NAND2 (N8016, N8007, N2199);
not NOT1 (N8017, N8009);
or OR2 (N8018, N8010, N669);
and AND3 (N8019, N8015, N363, N7699);
and AND3 (N8020, N7990, N336, N797);
nand NAND3 (N8021, N8000, N6736, N3664);
xor XOR2 (N8022, N8012, N3942);
xor XOR2 (N8023, N8022, N7421);
or OR4 (N8024, N8004, N3723, N6893, N5296);
not NOT1 (N8025, N8013);
nor NOR2 (N8026, N8019, N3954);
xor XOR2 (N8027, N8018, N4358);
not NOT1 (N8028, N8024);
not NOT1 (N8029, N8028);
and AND2 (N8030, N8020, N7651);
nand NAND3 (N8031, N8027, N6844, N3075);
buf BUF1 (N8032, N8030);
buf BUF1 (N8033, N8017);
nand NAND3 (N8034, N8025, N3716, N4251);
buf BUF1 (N8035, N8023);
xor XOR2 (N8036, N8026, N2903);
nand NAND3 (N8037, N8032, N3443, N932);
not NOT1 (N8038, N8014);
not NOT1 (N8039, N8033);
and AND3 (N8040, N8016, N3823, N6709);
xor XOR2 (N8041, N8039, N6352);
nor NOR3 (N8042, N8021, N2424, N5118);
and AND4 (N8043, N8040, N4915, N5686, N2091);
not NOT1 (N8044, N8035);
buf BUF1 (N8045, N8036);
xor XOR2 (N8046, N8029, N7262);
buf BUF1 (N8047, N8044);
buf BUF1 (N8048, N8031);
and AND2 (N8049, N8038, N280);
xor XOR2 (N8050, N8043, N3103);
and AND2 (N8051, N8048, N1451);
not NOT1 (N8052, N8045);
nand NAND4 (N8053, N8034, N7401, N7240, N385);
and AND4 (N8054, N8046, N5089, N1135, N894);
nand NAND2 (N8055, N8053, N3850);
buf BUF1 (N8056, N8042);
xor XOR2 (N8057, N8055, N5017);
buf BUF1 (N8058, N8051);
xor XOR2 (N8059, N8047, N2187);
not NOT1 (N8060, N8054);
nand NAND3 (N8061, N8059, N7622, N6627);
buf BUF1 (N8062, N8037);
xor XOR2 (N8063, N8057, N1528);
buf BUF1 (N8064, N8056);
nand NAND3 (N8065, N8049, N5313, N3909);
nor NOR4 (N8066, N8062, N1648, N5726, N5955);
and AND2 (N8067, N8061, N6085);
buf BUF1 (N8068, N8064);
xor XOR2 (N8069, N8041, N6102);
nand NAND3 (N8070, N8066, N1059, N2240);
nor NOR2 (N8071, N8052, N1543);
not NOT1 (N8072, N8050);
and AND3 (N8073, N8069, N1499, N4899);
buf BUF1 (N8074, N8068);
xor XOR2 (N8075, N8065, N7361);
nand NAND4 (N8076, N8072, N383, N6785, N5278);
and AND3 (N8077, N8075, N2457, N5372);
buf BUF1 (N8078, N8074);
nor NOR2 (N8079, N8076, N3974);
nand NAND4 (N8080, N8073, N7149, N1547, N4640);
nand NAND4 (N8081, N8067, N8052, N2898, N33);
nand NAND2 (N8082, N8077, N7783);
or OR4 (N8083, N8079, N6173, N3248, N1305);
or OR2 (N8084, N8060, N5980);
nor NOR2 (N8085, N8084, N229);
or OR2 (N8086, N8063, N6624);
nand NAND2 (N8087, N8080, N482);
not NOT1 (N8088, N8083);
or OR2 (N8089, N8070, N6348);
or OR3 (N8090, N8082, N1436, N596);
nor NOR2 (N8091, N8085, N6882);
xor XOR2 (N8092, N8081, N4761);
or OR4 (N8093, N8087, N6451, N5625, N1038);
nor NOR4 (N8094, N8090, N4088, N4954, N734);
not NOT1 (N8095, N8088);
nand NAND4 (N8096, N8095, N1584, N4684, N3993);
xor XOR2 (N8097, N8089, N7905);
and AND2 (N8098, N8096, N4620);
buf BUF1 (N8099, N8097);
not NOT1 (N8100, N8092);
xor XOR2 (N8101, N8091, N3313);
not NOT1 (N8102, N8100);
and AND3 (N8103, N8098, N5621, N5741);
not NOT1 (N8104, N8102);
or OR4 (N8105, N8078, N1025, N2990, N6879);
xor XOR2 (N8106, N8058, N7961);
nand NAND2 (N8107, N8099, N1913);
buf BUF1 (N8108, N8101);
and AND2 (N8109, N8107, N1849);
not NOT1 (N8110, N8109);
and AND2 (N8111, N8104, N3635);
not NOT1 (N8112, N8111);
or OR3 (N8113, N8086, N3898, N2619);
nand NAND2 (N8114, N8103, N3713);
nor NOR2 (N8115, N8106, N738);
not NOT1 (N8116, N8114);
nor NOR3 (N8117, N8116, N545, N31);
nor NOR4 (N8118, N8105, N1482, N156, N4029);
or OR2 (N8119, N8108, N4745);
xor XOR2 (N8120, N8094, N3779);
and AND2 (N8121, N8120, N7964);
and AND2 (N8122, N8113, N179);
or OR3 (N8123, N8112, N6410, N1042);
and AND2 (N8124, N8117, N4111);
nor NOR2 (N8125, N8121, N3191);
nor NOR3 (N8126, N8123, N8007, N134);
nand NAND3 (N8127, N8125, N7218, N6334);
nor NOR3 (N8128, N8127, N1150, N4952);
or OR2 (N8129, N8115, N648);
and AND2 (N8130, N8119, N3177);
xor XOR2 (N8131, N8124, N6730);
xor XOR2 (N8132, N8126, N4421);
or OR4 (N8133, N8118, N3858, N6700, N4671);
xor XOR2 (N8134, N8132, N4507);
buf BUF1 (N8135, N8110);
xor XOR2 (N8136, N8129, N5826);
nand NAND3 (N8137, N8136, N2793, N7686);
or OR3 (N8138, N8130, N3300, N869);
not NOT1 (N8139, N8071);
xor XOR2 (N8140, N8131, N7706);
xor XOR2 (N8141, N8122, N1273);
xor XOR2 (N8142, N8138, N4569);
nor NOR4 (N8143, N8139, N465, N4186, N7507);
or OR2 (N8144, N8128, N2850);
nor NOR2 (N8145, N8144, N4284);
nor NOR2 (N8146, N8135, N2790);
not NOT1 (N8147, N8141);
and AND3 (N8148, N8145, N4920, N3304);
buf BUF1 (N8149, N8147);
and AND2 (N8150, N8148, N3147);
or OR4 (N8151, N8140, N1123, N5132, N5281);
not NOT1 (N8152, N8137);
or OR3 (N8153, N8134, N1368, N1383);
buf BUF1 (N8154, N8153);
or OR2 (N8155, N8154, N2799);
and AND3 (N8156, N8155, N6091, N1109);
or OR4 (N8157, N8146, N528, N3066, N2065);
buf BUF1 (N8158, N8157);
nor NOR3 (N8159, N8152, N7384, N7816);
and AND3 (N8160, N8158, N6039, N751);
xor XOR2 (N8161, N8142, N2455);
nor NOR3 (N8162, N8093, N3043, N6453);
xor XOR2 (N8163, N8162, N4109);
nand NAND2 (N8164, N8150, N2734);
nand NAND4 (N8165, N8163, N6290, N3514, N264);
nand NAND4 (N8166, N8143, N2789, N7518, N1139);
nand NAND2 (N8167, N8151, N7576);
nor NOR2 (N8168, N8159, N1627);
and AND2 (N8169, N8161, N7135);
or OR2 (N8170, N8149, N7677);
not NOT1 (N8171, N8160);
not NOT1 (N8172, N8165);
nor NOR2 (N8173, N8170, N2512);
xor XOR2 (N8174, N8164, N1944);
xor XOR2 (N8175, N8156, N8047);
and AND4 (N8176, N8173, N2829, N3833, N5865);
buf BUF1 (N8177, N8172);
xor XOR2 (N8178, N8133, N1199);
xor XOR2 (N8179, N8169, N5428);
and AND3 (N8180, N8177, N185, N5298);
nand NAND2 (N8181, N8167, N2085);
nand NAND2 (N8182, N8168, N4059);
not NOT1 (N8183, N8181);
not NOT1 (N8184, N8175);
nand NAND4 (N8185, N8166, N4635, N61, N6084);
not NOT1 (N8186, N8179);
nand NAND3 (N8187, N8180, N2620, N7929);
nor NOR2 (N8188, N8176, N3233);
not NOT1 (N8189, N8185);
not NOT1 (N8190, N8186);
nor NOR2 (N8191, N8183, N4712);
not NOT1 (N8192, N8174);
nand NAND4 (N8193, N8178, N7720, N432, N1727);
buf BUF1 (N8194, N8189);
and AND4 (N8195, N8171, N1960, N303, N112);
nand NAND3 (N8196, N8184, N6155, N43);
nand NAND4 (N8197, N8191, N182, N3092, N2838);
not NOT1 (N8198, N8192);
buf BUF1 (N8199, N8195);
and AND3 (N8200, N8187, N1119, N2971);
or OR3 (N8201, N8194, N8084, N2914);
buf BUF1 (N8202, N8182);
or OR3 (N8203, N8199, N6342, N3216);
xor XOR2 (N8204, N8203, N1829);
nor NOR2 (N8205, N8190, N7027);
and AND2 (N8206, N8202, N4567);
buf BUF1 (N8207, N8201);
buf BUF1 (N8208, N8198);
nand NAND4 (N8209, N8208, N3509, N6014, N7121);
and AND3 (N8210, N8209, N527, N3541);
buf BUF1 (N8211, N8193);
buf BUF1 (N8212, N8188);
nor NOR2 (N8213, N8200, N2347);
nor NOR2 (N8214, N8210, N4951);
xor XOR2 (N8215, N8211, N55);
not NOT1 (N8216, N8215);
and AND3 (N8217, N8206, N2038, N2933);
buf BUF1 (N8218, N8212);
nand NAND4 (N8219, N8204, N1922, N8094, N5047);
nor NOR4 (N8220, N8218, N5472, N1213, N7281);
nor NOR4 (N8221, N8197, N5803, N7153, N7551);
not NOT1 (N8222, N8216);
nor NOR2 (N8223, N8196, N3108);
or OR2 (N8224, N8217, N1416);
or OR4 (N8225, N8213, N7998, N6842, N63);
and AND2 (N8226, N8220, N3454);
nor NOR4 (N8227, N8224, N2590, N1396, N3215);
or OR4 (N8228, N8207, N7708, N5191, N255);
not NOT1 (N8229, N8205);
xor XOR2 (N8230, N8222, N4514);
buf BUF1 (N8231, N8230);
buf BUF1 (N8232, N8225);
nor NOR4 (N8233, N8226, N7183, N5444, N3248);
xor XOR2 (N8234, N8232, N5223);
nand NAND2 (N8235, N8228, N252);
xor XOR2 (N8236, N8221, N1624);
nand NAND3 (N8237, N8235, N2937, N7346);
nor NOR3 (N8238, N8214, N5538, N3443);
or OR2 (N8239, N8231, N2242);
nand NAND3 (N8240, N8236, N2819, N7269);
nand NAND3 (N8241, N8219, N2928, N2649);
and AND2 (N8242, N8241, N393);
nor NOR2 (N8243, N8223, N3053);
and AND2 (N8244, N8242, N5509);
nor NOR2 (N8245, N8234, N5715);
nor NOR4 (N8246, N8237, N1427, N2773, N2652);
xor XOR2 (N8247, N8233, N5085);
nand NAND2 (N8248, N8247, N6601);
nor NOR2 (N8249, N8243, N5674);
or OR3 (N8250, N8246, N5968, N8007);
xor XOR2 (N8251, N8245, N3547);
not NOT1 (N8252, N8249);
nor NOR2 (N8253, N8244, N5396);
xor XOR2 (N8254, N8239, N3374);
nand NAND3 (N8255, N8253, N6759, N1544);
not NOT1 (N8256, N8252);
nand NAND3 (N8257, N8251, N5685, N3697);
nand NAND3 (N8258, N8250, N3873, N1919);
or OR3 (N8259, N8227, N7501, N2294);
and AND2 (N8260, N8258, N7313);
nor NOR2 (N8261, N8254, N2503);
nor NOR2 (N8262, N8261, N2038);
or OR4 (N8263, N8257, N3445, N6933, N4976);
nand NAND3 (N8264, N8240, N1542, N2492);
nor NOR3 (N8265, N8262, N5168, N3310);
nand NAND2 (N8266, N8248, N5941);
not NOT1 (N8267, N8255);
and AND3 (N8268, N8264, N2665, N5470);
nor NOR2 (N8269, N8267, N6712);
nor NOR4 (N8270, N8238, N1700, N6424, N594);
or OR4 (N8271, N8260, N3086, N6391, N6979);
not NOT1 (N8272, N8229);
nand NAND3 (N8273, N8268, N6688, N3661);
xor XOR2 (N8274, N8265, N1960);
and AND3 (N8275, N8270, N4949, N5650);
or OR3 (N8276, N8275, N758, N7517);
and AND4 (N8277, N8274, N474, N3712, N1496);
or OR2 (N8278, N8263, N7265);
and AND4 (N8279, N8277, N87, N433, N2407);
xor XOR2 (N8280, N8272, N6384);
xor XOR2 (N8281, N8278, N7048);
nor NOR3 (N8282, N8256, N3811, N2861);
not NOT1 (N8283, N8282);
xor XOR2 (N8284, N8281, N5252);
not NOT1 (N8285, N8269);
nor NOR4 (N8286, N8266, N7481, N7116, N8032);
nor NOR2 (N8287, N8280, N6701);
nor NOR2 (N8288, N8283, N3289);
nor NOR3 (N8289, N8288, N7646, N3953);
or OR4 (N8290, N8279, N3911, N6534, N2674);
or OR4 (N8291, N8284, N3869, N6052, N4182);
xor XOR2 (N8292, N8259, N6055);
and AND3 (N8293, N8271, N2136, N498);
nor NOR3 (N8294, N8276, N6241, N3367);
nand NAND2 (N8295, N8285, N3168);
not NOT1 (N8296, N8286);
buf BUF1 (N8297, N8287);
and AND3 (N8298, N8297, N2101, N1395);
not NOT1 (N8299, N8294);
and AND2 (N8300, N8299, N7520);
buf BUF1 (N8301, N8289);
xor XOR2 (N8302, N8290, N6585);
not NOT1 (N8303, N8301);
and AND2 (N8304, N8303, N7494);
xor XOR2 (N8305, N8296, N8000);
nor NOR2 (N8306, N8302, N4422);
buf BUF1 (N8307, N8305);
nand NAND4 (N8308, N8273, N2551, N4262, N5958);
nand NAND2 (N8309, N8306, N6806);
and AND3 (N8310, N8298, N6315, N7389);
not NOT1 (N8311, N8292);
xor XOR2 (N8312, N8291, N6827);
or OR2 (N8313, N8309, N6995);
or OR4 (N8314, N8312, N1840, N5698, N2585);
not NOT1 (N8315, N8300);
not NOT1 (N8316, N8293);
nand NAND4 (N8317, N8311, N1585, N5533, N1817);
not NOT1 (N8318, N8316);
buf BUF1 (N8319, N8318);
nor NOR2 (N8320, N8307, N1884);
and AND4 (N8321, N8313, N6618, N538, N5028);
not NOT1 (N8322, N8310);
buf BUF1 (N8323, N8304);
and AND4 (N8324, N8315, N1468, N1187, N6543);
buf BUF1 (N8325, N8295);
xor XOR2 (N8326, N8322, N1866);
nor NOR2 (N8327, N8314, N4491);
and AND4 (N8328, N8323, N3556, N1716, N3289);
nor NOR4 (N8329, N8317, N5451, N5978, N5143);
xor XOR2 (N8330, N8308, N3207);
nand NAND2 (N8331, N8326, N5679);
nand NAND4 (N8332, N8330, N793, N5224, N7764);
nand NAND3 (N8333, N8324, N6021, N6625);
not NOT1 (N8334, N8332);
or OR3 (N8335, N8329, N2792, N7072);
not NOT1 (N8336, N8335);
not NOT1 (N8337, N8325);
nand NAND2 (N8338, N8320, N7540);
or OR2 (N8339, N8333, N5879);
not NOT1 (N8340, N8327);
buf BUF1 (N8341, N8339);
or OR3 (N8342, N8334, N1748, N2547);
nor NOR2 (N8343, N8342, N2045);
xor XOR2 (N8344, N8343, N6507);
not NOT1 (N8345, N8328);
nor NOR4 (N8346, N8341, N5392, N2197, N5844);
xor XOR2 (N8347, N8336, N7116);
nor NOR3 (N8348, N8344, N4148, N2461);
or OR4 (N8349, N8348, N4478, N183, N5282);
nand NAND2 (N8350, N8319, N4526);
nor NOR2 (N8351, N8338, N8058);
not NOT1 (N8352, N8349);
and AND2 (N8353, N8345, N4562);
xor XOR2 (N8354, N8351, N4638);
not NOT1 (N8355, N8354);
nand NAND4 (N8356, N8340, N7278, N7280, N6429);
and AND4 (N8357, N8350, N6134, N537, N919);
and AND3 (N8358, N8346, N8259, N6925);
and AND3 (N8359, N8355, N5450, N5043);
and AND4 (N8360, N8321, N1288, N6033, N4818);
buf BUF1 (N8361, N8359);
and AND3 (N8362, N8331, N4209, N2003);
nand NAND3 (N8363, N8357, N4169, N7218);
nand NAND4 (N8364, N8358, N3036, N433, N3569);
and AND2 (N8365, N8352, N7129);
and AND3 (N8366, N8361, N3370, N4214);
xor XOR2 (N8367, N8360, N410);
nand NAND2 (N8368, N8362, N6132);
nand NAND4 (N8369, N8365, N8297, N4489, N1995);
and AND3 (N8370, N8363, N6859, N1852);
xor XOR2 (N8371, N8369, N6495);
not NOT1 (N8372, N8368);
nor NOR3 (N8373, N8356, N7059, N6296);
or OR3 (N8374, N8370, N4763, N1778);
nand NAND2 (N8375, N8347, N4779);
buf BUF1 (N8376, N8337);
nand NAND3 (N8377, N8376, N657, N3138);
and AND4 (N8378, N8353, N2401, N1681, N1813);
xor XOR2 (N8379, N8366, N1377);
xor XOR2 (N8380, N8371, N4811);
or OR4 (N8381, N8380, N1832, N4056, N2230);
and AND3 (N8382, N8381, N5129, N7877);
buf BUF1 (N8383, N8378);
or OR4 (N8384, N8377, N389, N2863, N4502);
and AND3 (N8385, N8373, N4920, N7875);
buf BUF1 (N8386, N8367);
xor XOR2 (N8387, N8375, N4614);
xor XOR2 (N8388, N8383, N1909);
nor NOR3 (N8389, N8387, N6855, N252);
not NOT1 (N8390, N8382);
and AND2 (N8391, N8364, N5921);
buf BUF1 (N8392, N8374);
xor XOR2 (N8393, N8385, N2337);
and AND2 (N8394, N8384, N4475);
nand NAND3 (N8395, N8394, N6382, N1826);
xor XOR2 (N8396, N8390, N2786);
nand NAND4 (N8397, N8396, N8084, N1180, N8092);
buf BUF1 (N8398, N8379);
and AND4 (N8399, N8395, N3920, N4176, N5501);
not NOT1 (N8400, N8389);
xor XOR2 (N8401, N8399, N2426);
and AND4 (N8402, N8388, N6243, N5414, N6361);
xor XOR2 (N8403, N8386, N87);
nand NAND2 (N8404, N8393, N413);
nor NOR4 (N8405, N8402, N8170, N1239, N2538);
buf BUF1 (N8406, N8397);
buf BUF1 (N8407, N8401);
xor XOR2 (N8408, N8403, N1093);
buf BUF1 (N8409, N8405);
nand NAND3 (N8410, N8409, N6659, N2959);
nor NOR4 (N8411, N8391, N4785, N4726, N2717);
or OR2 (N8412, N8411, N2737);
and AND3 (N8413, N8372, N7055, N6489);
not NOT1 (N8414, N8392);
and AND4 (N8415, N8404, N4190, N736, N7720);
or OR3 (N8416, N8414, N7674, N4169);
buf BUF1 (N8417, N8410);
buf BUF1 (N8418, N8408);
nand NAND4 (N8419, N8407, N1824, N1627, N5885);
not NOT1 (N8420, N8412);
xor XOR2 (N8421, N8400, N2251);
and AND2 (N8422, N8406, N8369);
and AND3 (N8423, N8421, N2359, N5381);
and AND4 (N8424, N8423, N8010, N23, N3048);
nand NAND3 (N8425, N8419, N8244, N4997);
buf BUF1 (N8426, N8425);
buf BUF1 (N8427, N8426);
nor NOR4 (N8428, N8417, N6058, N2983, N7796);
buf BUF1 (N8429, N8420);
nand NAND2 (N8430, N8413, N2854);
and AND2 (N8431, N8416, N4917);
not NOT1 (N8432, N8431);
not NOT1 (N8433, N8422);
nor NOR3 (N8434, N8429, N2215, N5519);
not NOT1 (N8435, N8398);
buf BUF1 (N8436, N8427);
and AND4 (N8437, N8435, N3029, N2819, N5654);
and AND4 (N8438, N8437, N8060, N7991, N7057);
or OR3 (N8439, N8424, N3363, N5693);
nand NAND3 (N8440, N8415, N364, N1334);
not NOT1 (N8441, N8440);
and AND2 (N8442, N8439, N7977);
not NOT1 (N8443, N8430);
nor NOR4 (N8444, N8432, N3461, N8233, N3207);
not NOT1 (N8445, N8428);
buf BUF1 (N8446, N8441);
nand NAND2 (N8447, N8434, N3934);
and AND3 (N8448, N8433, N4298, N3072);
nor NOR2 (N8449, N8446, N3935);
nand NAND2 (N8450, N8436, N3569);
not NOT1 (N8451, N8442);
buf BUF1 (N8452, N8447);
and AND4 (N8453, N8445, N2919, N2803, N3206);
xor XOR2 (N8454, N8451, N3546);
buf BUF1 (N8455, N8454);
and AND3 (N8456, N8453, N794, N5768);
not NOT1 (N8457, N8418);
nand NAND4 (N8458, N8443, N4536, N4623, N1980);
and AND3 (N8459, N8458, N1046, N5550);
nand NAND4 (N8460, N8455, N2395, N8406, N2280);
nor NOR3 (N8461, N8459, N916, N2502);
nand NAND4 (N8462, N8449, N5380, N2677, N3650);
and AND4 (N8463, N8438, N1621, N2138, N4645);
and AND4 (N8464, N8460, N5678, N868, N7003);
buf BUF1 (N8465, N8463);
and AND2 (N8466, N8465, N89);
xor XOR2 (N8467, N8456, N5);
nand NAND4 (N8468, N8467, N6660, N1002, N5984);
nand NAND2 (N8469, N8462, N379);
not NOT1 (N8470, N8450);
nand NAND3 (N8471, N8470, N7131, N3678);
and AND4 (N8472, N8457, N6484, N801, N8302);
and AND4 (N8473, N8466, N7703, N4144, N877);
xor XOR2 (N8474, N8472, N6854);
or OR3 (N8475, N8474, N4991, N6116);
not NOT1 (N8476, N8464);
nor NOR4 (N8477, N8444, N174, N4554, N290);
buf BUF1 (N8478, N8448);
nand NAND2 (N8479, N8471, N3179);
nand NAND2 (N8480, N8461, N1946);
nor NOR2 (N8481, N8478, N6568);
xor XOR2 (N8482, N8476, N6544);
and AND4 (N8483, N8477, N8434, N6510, N113);
not NOT1 (N8484, N8469);
nor NOR2 (N8485, N8468, N3840);
or OR2 (N8486, N8484, N5179);
buf BUF1 (N8487, N8475);
nor NOR3 (N8488, N8480, N4913, N3747);
not NOT1 (N8489, N8487);
xor XOR2 (N8490, N8481, N7565);
xor XOR2 (N8491, N8452, N2784);
xor XOR2 (N8492, N8485, N3358);
and AND4 (N8493, N8473, N2558, N6834, N2915);
or OR2 (N8494, N8483, N3125);
nor NOR3 (N8495, N8488, N2278, N2269);
xor XOR2 (N8496, N8493, N5430);
nor NOR3 (N8497, N8496, N7042, N5394);
not NOT1 (N8498, N8491);
xor XOR2 (N8499, N8486, N2716);
nor NOR3 (N8500, N8489, N6121, N5024);
nand NAND4 (N8501, N8482, N6566, N7092, N5727);
xor XOR2 (N8502, N8494, N1477);
nand NAND4 (N8503, N8501, N3697, N2924, N5316);
nor NOR2 (N8504, N8492, N3397);
not NOT1 (N8505, N8479);
nand NAND2 (N8506, N8505, N7758);
not NOT1 (N8507, N8498);
or OR4 (N8508, N8502, N5896, N2438, N1673);
nand NAND3 (N8509, N8504, N7856, N4922);
nor NOR4 (N8510, N8497, N7889, N1593, N3002);
buf BUF1 (N8511, N8507);
and AND3 (N8512, N8495, N1008, N8114);
not NOT1 (N8513, N8499);
not NOT1 (N8514, N8512);
nor NOR4 (N8515, N8508, N1721, N7748, N7300);
or OR2 (N8516, N8500, N1464);
nand NAND3 (N8517, N8503, N7888, N5568);
and AND4 (N8518, N8490, N6866, N3514, N1852);
nor NOR2 (N8519, N8510, N2159);
not NOT1 (N8520, N8516);
nor NOR2 (N8521, N8514, N4670);
and AND3 (N8522, N8509, N3205, N5518);
and AND2 (N8523, N8517, N5804);
xor XOR2 (N8524, N8521, N7238);
xor XOR2 (N8525, N8506, N3862);
or OR2 (N8526, N8513, N1566);
nand NAND4 (N8527, N8524, N841, N7604, N3827);
buf BUF1 (N8528, N8511);
not NOT1 (N8529, N8526);
not NOT1 (N8530, N8527);
buf BUF1 (N8531, N8519);
nand NAND3 (N8532, N8520, N5305, N2909);
nand NAND2 (N8533, N8515, N823);
nand NAND3 (N8534, N8525, N1195, N1284);
and AND2 (N8535, N8523, N7488);
nor NOR3 (N8536, N8532, N961, N3093);
not NOT1 (N8537, N8536);
nor NOR3 (N8538, N8529, N3974, N5933);
and AND3 (N8539, N8533, N7737, N5825);
nor NOR2 (N8540, N8530, N7541);
xor XOR2 (N8541, N8534, N7105);
and AND2 (N8542, N8522, N7569);
or OR2 (N8543, N8542, N6465);
xor XOR2 (N8544, N8528, N7139);
nand NAND4 (N8545, N8518, N461, N3886, N338);
xor XOR2 (N8546, N8538, N1603);
xor XOR2 (N8547, N8545, N4085);
xor XOR2 (N8548, N8535, N5442);
nand NAND4 (N8549, N8548, N4123, N2935, N7795);
xor XOR2 (N8550, N8547, N3114);
xor XOR2 (N8551, N8531, N6136);
or OR2 (N8552, N8550, N7143);
buf BUF1 (N8553, N8546);
nand NAND3 (N8554, N8541, N2634, N1379);
xor XOR2 (N8555, N8537, N139);
nand NAND3 (N8556, N8543, N5288, N6973);
nand NAND4 (N8557, N8549, N3090, N5698, N5);
or OR2 (N8558, N8557, N311);
xor XOR2 (N8559, N8558, N7027);
nor NOR4 (N8560, N8540, N6133, N3223, N8079);
not NOT1 (N8561, N8544);
buf BUF1 (N8562, N8554);
buf BUF1 (N8563, N8556);
xor XOR2 (N8564, N8563, N5154);
or OR2 (N8565, N8562, N651);
nand NAND3 (N8566, N8555, N1119, N1749);
or OR4 (N8567, N8539, N706, N3551, N5094);
and AND4 (N8568, N8560, N6226, N6880, N132);
nand NAND2 (N8569, N8559, N4079);
not NOT1 (N8570, N8564);
or OR4 (N8571, N8561, N7059, N6751, N7704);
and AND3 (N8572, N8568, N2553, N6274);
buf BUF1 (N8573, N8567);
and AND4 (N8574, N8572, N2468, N7726, N2584);
nand NAND2 (N8575, N8565, N3317);
buf BUF1 (N8576, N8573);
buf BUF1 (N8577, N8551);
not NOT1 (N8578, N8552);
nand NAND3 (N8579, N8571, N4958, N7313);
buf BUF1 (N8580, N8574);
not NOT1 (N8581, N8579);
nor NOR4 (N8582, N8576, N1536, N5034, N1519);
nor NOR2 (N8583, N8580, N4075);
and AND4 (N8584, N8578, N1505, N7252, N4866);
not NOT1 (N8585, N8575);
nor NOR3 (N8586, N8582, N4272, N1948);
buf BUF1 (N8587, N8553);
or OR4 (N8588, N8577, N3304, N384, N54);
and AND3 (N8589, N8583, N1111, N5418);
nand NAND4 (N8590, N8566, N5147, N5479, N7994);
and AND2 (N8591, N8569, N6670);
buf BUF1 (N8592, N8590);
not NOT1 (N8593, N8570);
or OR4 (N8594, N8581, N3498, N2449, N6240);
xor XOR2 (N8595, N8584, N1744);
and AND3 (N8596, N8594, N1916, N5596);
nand NAND3 (N8597, N8588, N1927, N6286);
buf BUF1 (N8598, N8596);
nor NOR4 (N8599, N8598, N2983, N6792, N6757);
buf BUF1 (N8600, N8599);
and AND4 (N8601, N8585, N1684, N2185, N5822);
and AND3 (N8602, N8587, N7380, N4440);
nor NOR2 (N8603, N8602, N5378);
buf BUF1 (N8604, N8593);
xor XOR2 (N8605, N8597, N2692);
not NOT1 (N8606, N8605);
or OR2 (N8607, N8606, N5917);
or OR3 (N8608, N8591, N507, N1427);
or OR4 (N8609, N8604, N1352, N3304, N1243);
buf BUF1 (N8610, N8607);
or OR4 (N8611, N8595, N1459, N5673, N3821);
not NOT1 (N8612, N8600);
xor XOR2 (N8613, N8608, N5440);
not NOT1 (N8614, N8610);
xor XOR2 (N8615, N8601, N461);
or OR3 (N8616, N8603, N5595, N2924);
and AND4 (N8617, N8614, N235, N8505, N701);
and AND2 (N8618, N8611, N2312);
xor XOR2 (N8619, N8613, N7274);
xor XOR2 (N8620, N8616, N4033);
or OR2 (N8621, N8592, N8372);
nand NAND2 (N8622, N8609, N4767);
not NOT1 (N8623, N8615);
buf BUF1 (N8624, N8586);
nor NOR3 (N8625, N8617, N6074, N3409);
nand NAND3 (N8626, N8618, N6632, N4639);
and AND3 (N8627, N8625, N2946, N755);
xor XOR2 (N8628, N8620, N7942);
xor XOR2 (N8629, N8619, N6010);
xor XOR2 (N8630, N8612, N4327);
and AND4 (N8631, N8626, N2392, N1417, N1934);
nor NOR4 (N8632, N8630, N263, N2803, N3421);
nor NOR4 (N8633, N8629, N4001, N8355, N830);
buf BUF1 (N8634, N8632);
not NOT1 (N8635, N8589);
xor XOR2 (N8636, N8634, N1952);
buf BUF1 (N8637, N8623);
nand NAND2 (N8638, N8622, N2354);
nor NOR3 (N8639, N8635, N8455, N6862);
not NOT1 (N8640, N8621);
xor XOR2 (N8641, N8637, N5941);
nand NAND2 (N8642, N8640, N3632);
nor NOR4 (N8643, N8641, N2547, N822, N3124);
nand NAND4 (N8644, N8624, N6260, N2015, N8316);
not NOT1 (N8645, N8631);
nor NOR4 (N8646, N8643, N2220, N3022, N3401);
nor NOR2 (N8647, N8644, N1326);
or OR4 (N8648, N8639, N4908, N6393, N8463);
not NOT1 (N8649, N8638);
nand NAND3 (N8650, N8648, N7866, N4475);
or OR3 (N8651, N8636, N4381, N6282);
nand NAND3 (N8652, N8647, N6670, N2539);
nand NAND2 (N8653, N8651, N8204);
xor XOR2 (N8654, N8645, N2061);
nor NOR3 (N8655, N8633, N8011, N5211);
nand NAND3 (N8656, N8653, N814, N5987);
nor NOR4 (N8657, N8649, N2626, N4, N1120);
nor NOR3 (N8658, N8654, N4971, N6501);
or OR3 (N8659, N8627, N4360, N3509);
and AND3 (N8660, N8646, N7830, N8050);
buf BUF1 (N8661, N8628);
nand NAND2 (N8662, N8661, N2957);
nand NAND4 (N8663, N8658, N1242, N3688, N1885);
not NOT1 (N8664, N8662);
nand NAND4 (N8665, N8657, N1547, N3105, N6311);
nand NAND3 (N8666, N8656, N5285, N3136);
buf BUF1 (N8667, N8665);
or OR3 (N8668, N8660, N7732, N2725);
or OR3 (N8669, N8650, N3556, N6037);
and AND4 (N8670, N8667, N7412, N4390, N2538);
or OR4 (N8671, N8652, N368, N8641, N639);
nor NOR4 (N8672, N8663, N2636, N1001, N2889);
xor XOR2 (N8673, N8642, N3344);
xor XOR2 (N8674, N8672, N8582);
and AND3 (N8675, N8664, N6410, N4296);
nand NAND4 (N8676, N8674, N3518, N3598, N7934);
nor NOR2 (N8677, N8670, N6168);
not NOT1 (N8678, N8659);
and AND2 (N8679, N8655, N4665);
xor XOR2 (N8680, N8675, N1819);
not NOT1 (N8681, N8676);
nor NOR2 (N8682, N8680, N8466);
and AND2 (N8683, N8666, N5524);
buf BUF1 (N8684, N8682);
buf BUF1 (N8685, N8677);
not NOT1 (N8686, N8668);
xor XOR2 (N8687, N8685, N7155);
buf BUF1 (N8688, N8678);
xor XOR2 (N8689, N8671, N8629);
nand NAND2 (N8690, N8683, N7615);
xor XOR2 (N8691, N8673, N567);
xor XOR2 (N8692, N8688, N8586);
or OR2 (N8693, N8669, N7040);
nor NOR2 (N8694, N8681, N5867);
nand NAND2 (N8695, N8689, N8529);
buf BUF1 (N8696, N8684);
buf BUF1 (N8697, N8695);
and AND2 (N8698, N8693, N4624);
nand NAND4 (N8699, N8687, N4687, N6638, N4839);
and AND3 (N8700, N8679, N2764, N2549);
nor NOR2 (N8701, N8699, N5534);
buf BUF1 (N8702, N8692);
not NOT1 (N8703, N8698);
buf BUF1 (N8704, N8700);
and AND4 (N8705, N8703, N4381, N715, N8610);
not NOT1 (N8706, N8690);
nand NAND2 (N8707, N8691, N8307);
and AND4 (N8708, N8706, N6241, N7402, N6360);
nand NAND4 (N8709, N8708, N6234, N6372, N6788);
xor XOR2 (N8710, N8694, N5313);
not NOT1 (N8711, N8709);
nand NAND2 (N8712, N8710, N7076);
nand NAND3 (N8713, N8707, N6881, N2990);
buf BUF1 (N8714, N8697);
nor NOR3 (N8715, N8711, N5567, N8266);
and AND3 (N8716, N8714, N3750, N1418);
nor NOR3 (N8717, N8686, N2595, N8261);
or OR3 (N8718, N8704, N4320, N7265);
not NOT1 (N8719, N8713);
not NOT1 (N8720, N8702);
buf BUF1 (N8721, N8716);
buf BUF1 (N8722, N8705);
and AND3 (N8723, N8715, N8228, N6177);
and AND4 (N8724, N8696, N1264, N3302, N1980);
not NOT1 (N8725, N8724);
and AND3 (N8726, N8717, N621, N434);
and AND3 (N8727, N8719, N7936, N5338);
buf BUF1 (N8728, N8722);
nor NOR3 (N8729, N8701, N3648, N7980);
not NOT1 (N8730, N8718);
buf BUF1 (N8731, N8727);
nor NOR4 (N8732, N8730, N4988, N5321, N2663);
buf BUF1 (N8733, N8723);
or OR4 (N8734, N8726, N8315, N7318, N5328);
nand NAND3 (N8735, N8725, N7040, N8216);
xor XOR2 (N8736, N8712, N2096);
buf BUF1 (N8737, N8731);
or OR2 (N8738, N8732, N97);
nor NOR3 (N8739, N8733, N4126, N6058);
buf BUF1 (N8740, N8737);
buf BUF1 (N8741, N8739);
xor XOR2 (N8742, N8735, N4211);
xor XOR2 (N8743, N8738, N2703);
nor NOR2 (N8744, N8729, N3313);
and AND4 (N8745, N8741, N7168, N1706, N6141);
or OR4 (N8746, N8720, N8739, N7276, N3003);
xor XOR2 (N8747, N8745, N4060);
nand NAND2 (N8748, N8734, N69);
or OR3 (N8749, N8748, N7888, N2843);
or OR4 (N8750, N8736, N2720, N50, N8403);
or OR4 (N8751, N8742, N5800, N6917, N3319);
and AND2 (N8752, N8740, N147);
xor XOR2 (N8753, N8721, N2801);
nor NOR2 (N8754, N8743, N5164);
and AND3 (N8755, N8754, N5858, N6619);
nor NOR3 (N8756, N8744, N1348, N7953);
xor XOR2 (N8757, N8728, N2715);
nor NOR2 (N8758, N8753, N669);
xor XOR2 (N8759, N8751, N5539);
or OR2 (N8760, N8746, N5654);
xor XOR2 (N8761, N8747, N8306);
and AND3 (N8762, N8752, N7700, N6722);
buf BUF1 (N8763, N8755);
xor XOR2 (N8764, N8759, N349);
nor NOR4 (N8765, N8763, N4096, N3338, N19);
not NOT1 (N8766, N8761);
xor XOR2 (N8767, N8764, N3795);
or OR4 (N8768, N8758, N6125, N5304, N3696);
nand NAND4 (N8769, N8750, N2878, N2843, N1276);
nor NOR4 (N8770, N8766, N6406, N4731, N5604);
xor XOR2 (N8771, N8749, N7633);
xor XOR2 (N8772, N8767, N6242);
buf BUF1 (N8773, N8765);
not NOT1 (N8774, N8757);
nand NAND2 (N8775, N8772, N7290);
buf BUF1 (N8776, N8774);
or OR2 (N8777, N8773, N4739);
or OR2 (N8778, N8776, N7900);
nor NOR3 (N8779, N8769, N293, N7134);
xor XOR2 (N8780, N8775, N4105);
and AND4 (N8781, N8779, N2999, N3299, N6479);
nand NAND2 (N8782, N8760, N4658);
or OR4 (N8783, N8782, N2138, N1635, N8732);
nor NOR4 (N8784, N8756, N8622, N3496, N992);
not NOT1 (N8785, N8771);
and AND3 (N8786, N8768, N7215, N5629);
xor XOR2 (N8787, N8780, N6587);
or OR2 (N8788, N8783, N7337);
not NOT1 (N8789, N8781);
or OR3 (N8790, N8762, N3492, N2218);
nor NOR4 (N8791, N8787, N6861, N5418, N4761);
nand NAND4 (N8792, N8784, N6013, N2451, N6414);
nand NAND4 (N8793, N8791, N831, N7225, N6223);
nor NOR3 (N8794, N8786, N7801, N3138);
buf BUF1 (N8795, N8770);
xor XOR2 (N8796, N8788, N8710);
not NOT1 (N8797, N8795);
and AND2 (N8798, N8789, N7207);
nor NOR2 (N8799, N8778, N4984);
not NOT1 (N8800, N8799);
nor NOR2 (N8801, N8794, N3014);
nand NAND2 (N8802, N8777, N4424);
not NOT1 (N8803, N8802);
not NOT1 (N8804, N8785);
nand NAND2 (N8805, N8793, N5245);
xor XOR2 (N8806, N8798, N1414);
not NOT1 (N8807, N8800);
not NOT1 (N8808, N8792);
nor NOR3 (N8809, N8805, N5995, N6335);
nand NAND3 (N8810, N8801, N6615, N6488);
or OR3 (N8811, N8803, N7000, N7995);
and AND4 (N8812, N8807, N7588, N1116, N8809);
nor NOR2 (N8813, N4957, N2851);
or OR3 (N8814, N8811, N7455, N1963);
nor NOR2 (N8815, N8806, N3156);
nor NOR3 (N8816, N8796, N8465, N1290);
buf BUF1 (N8817, N8790);
or OR4 (N8818, N8817, N8462, N6909, N179);
or OR2 (N8819, N8818, N2236);
nand NAND2 (N8820, N8813, N1744);
nand NAND3 (N8821, N8804, N5611, N2922);
not NOT1 (N8822, N8808);
or OR2 (N8823, N8812, N3333);
nand NAND3 (N8824, N8822, N3729, N6019);
nor NOR2 (N8825, N8797, N5804);
nand NAND3 (N8826, N8816, N3070, N7296);
xor XOR2 (N8827, N8810, N7663);
nand NAND2 (N8828, N8825, N2074);
not NOT1 (N8829, N8820);
or OR2 (N8830, N8815, N4424);
buf BUF1 (N8831, N8828);
nor NOR2 (N8832, N8819, N1057);
nand NAND4 (N8833, N8826, N6088, N2249, N5429);
buf BUF1 (N8834, N8833);
not NOT1 (N8835, N8831);
xor XOR2 (N8836, N8821, N1581);
and AND3 (N8837, N8823, N2599, N8549);
not NOT1 (N8838, N8834);
xor XOR2 (N8839, N8814, N8591);
or OR3 (N8840, N8824, N7306, N7495);
nor NOR4 (N8841, N8836, N6478, N1097, N4412);
nor NOR4 (N8842, N8830, N2331, N6493, N7997);
not NOT1 (N8843, N8827);
or OR3 (N8844, N8838, N8270, N3067);
nand NAND4 (N8845, N8837, N129, N3440, N1876);
xor XOR2 (N8846, N8839, N2071);
not NOT1 (N8847, N8841);
nor NOR2 (N8848, N8845, N6499);
or OR2 (N8849, N8835, N2236);
nand NAND4 (N8850, N8844, N52, N6365, N2248);
nand NAND4 (N8851, N8848, N2143, N1001, N8135);
nand NAND2 (N8852, N8843, N5286);
or OR2 (N8853, N8840, N425);
nor NOR4 (N8854, N8847, N4944, N1555, N5843);
not NOT1 (N8855, N8852);
or OR3 (N8856, N8849, N7496, N667);
and AND2 (N8857, N8846, N1693);
xor XOR2 (N8858, N8857, N5098);
nand NAND3 (N8859, N8853, N5688, N3596);
nor NOR2 (N8860, N8858, N7814);
xor XOR2 (N8861, N8842, N4309);
not NOT1 (N8862, N8854);
buf BUF1 (N8863, N8861);
buf BUF1 (N8864, N8859);
xor XOR2 (N8865, N8863, N8053);
nor NOR4 (N8866, N8860, N2947, N3375, N4844);
and AND2 (N8867, N8855, N5055);
not NOT1 (N8868, N8829);
nor NOR2 (N8869, N8832, N2443);
or OR2 (N8870, N8865, N3344);
xor XOR2 (N8871, N8851, N1039);
buf BUF1 (N8872, N8867);
xor XOR2 (N8873, N8870, N5509);
nand NAND2 (N8874, N8869, N3825);
and AND3 (N8875, N8864, N2043, N3750);
nand NAND2 (N8876, N8868, N1489);
buf BUF1 (N8877, N8850);
and AND3 (N8878, N8877, N7510, N690);
and AND2 (N8879, N8872, N7914);
not NOT1 (N8880, N8879);
not NOT1 (N8881, N8873);
xor XOR2 (N8882, N8878, N4662);
or OR2 (N8883, N8881, N6031);
buf BUF1 (N8884, N8874);
or OR3 (N8885, N8884, N4014, N7608);
nor NOR4 (N8886, N8880, N2256, N7871, N8688);
xor XOR2 (N8887, N8886, N8042);
nand NAND4 (N8888, N8871, N2108, N2016, N5620);
buf BUF1 (N8889, N8866);
and AND2 (N8890, N8889, N3472);
and AND3 (N8891, N8887, N7006, N7069);
or OR3 (N8892, N8883, N2697, N1691);
xor XOR2 (N8893, N8862, N6996);
buf BUF1 (N8894, N8892);
nand NAND3 (N8895, N8856, N2677, N2798);
nor NOR3 (N8896, N8885, N5106, N6676);
and AND2 (N8897, N8894, N3725);
nand NAND2 (N8898, N8896, N7582);
nand NAND2 (N8899, N8891, N7781);
and AND2 (N8900, N8899, N2879);
and AND2 (N8901, N8895, N3786);
or OR3 (N8902, N8900, N6012, N6900);
and AND4 (N8903, N8898, N480, N2090, N4909);
xor XOR2 (N8904, N8897, N3000);
nor NOR4 (N8905, N8893, N139, N1195, N1932);
nand NAND2 (N8906, N8888, N4771);
and AND2 (N8907, N8905, N7504);
nor NOR4 (N8908, N8901, N6238, N5625, N3531);
not NOT1 (N8909, N8875);
buf BUF1 (N8910, N8909);
xor XOR2 (N8911, N8907, N4277);
or OR3 (N8912, N8904, N6298, N3016);
nor NOR2 (N8913, N8912, N5750);
xor XOR2 (N8914, N8890, N1615);
buf BUF1 (N8915, N8882);
not NOT1 (N8916, N8915);
nor NOR4 (N8917, N8908, N6869, N1559, N4472);
or OR3 (N8918, N8917, N4001, N3910);
and AND2 (N8919, N8918, N4572);
or OR4 (N8920, N8903, N6377, N441, N188);
and AND2 (N8921, N8910, N4475);
xor XOR2 (N8922, N8919, N7072);
nand NAND4 (N8923, N8902, N5499, N2465, N8562);
not NOT1 (N8924, N8920);
not NOT1 (N8925, N8876);
nand NAND3 (N8926, N8921, N3445, N8253);
nand NAND4 (N8927, N8924, N4075, N3204, N4946);
not NOT1 (N8928, N8911);
or OR2 (N8929, N8923, N8132);
nand NAND4 (N8930, N8929, N3881, N979, N3358);
nor NOR2 (N8931, N8925, N6410);
and AND3 (N8932, N8922, N3313, N7465);
nor NOR3 (N8933, N8930, N5471, N6530);
nand NAND2 (N8934, N8932, N5909);
and AND4 (N8935, N8933, N4353, N345, N1473);
nor NOR4 (N8936, N8934, N6416, N4254, N8182);
or OR4 (N8937, N8914, N2635, N6974, N6971);
nor NOR3 (N8938, N8913, N8796, N3738);
or OR3 (N8939, N8935, N153, N7505);
not NOT1 (N8940, N8931);
not NOT1 (N8941, N8906);
not NOT1 (N8942, N8927);
buf BUF1 (N8943, N8941);
or OR3 (N8944, N8943, N4467, N5159);
buf BUF1 (N8945, N8944);
and AND3 (N8946, N8942, N3729, N491);
nand NAND2 (N8947, N8937, N132);
xor XOR2 (N8948, N8936, N5912);
nor NOR4 (N8949, N8945, N5092, N3937, N8162);
and AND4 (N8950, N8938, N6737, N3963, N134);
buf BUF1 (N8951, N8949);
buf BUF1 (N8952, N8948);
nor NOR3 (N8953, N8939, N2266, N6435);
buf BUF1 (N8954, N8916);
xor XOR2 (N8955, N8953, N5324);
nand NAND4 (N8956, N8952, N4177, N3786, N873);
not NOT1 (N8957, N8940);
nor NOR3 (N8958, N8957, N8770, N7759);
xor XOR2 (N8959, N8954, N6846);
or OR3 (N8960, N8956, N6620, N1084);
buf BUF1 (N8961, N8959);
or OR3 (N8962, N8946, N7607, N6099);
nor NOR4 (N8963, N8961, N6911, N5335, N816);
nor NOR4 (N8964, N8947, N5167, N1722, N1316);
buf BUF1 (N8965, N8960);
nor NOR4 (N8966, N8964, N7702, N2909, N1548);
and AND4 (N8967, N8965, N1247, N5305, N731);
buf BUF1 (N8968, N8962);
and AND4 (N8969, N8928, N2536, N3586, N3516);
or OR2 (N8970, N8969, N8160);
and AND3 (N8971, N8966, N7360, N8298);
or OR3 (N8972, N8950, N5098, N5707);
and AND3 (N8973, N8958, N2382, N8567);
xor XOR2 (N8974, N8951, N5934);
and AND2 (N8975, N8968, N2842);
buf BUF1 (N8976, N8973);
xor XOR2 (N8977, N8972, N4047);
and AND2 (N8978, N8974, N4287);
nor NOR3 (N8979, N8978, N857, N7673);
and AND4 (N8980, N8955, N3344, N332, N8664);
nand NAND3 (N8981, N8970, N8042, N7932);
or OR3 (N8982, N8926, N543, N6030);
not NOT1 (N8983, N8977);
not NOT1 (N8984, N8983);
not NOT1 (N8985, N8980);
not NOT1 (N8986, N8975);
not NOT1 (N8987, N8976);
and AND2 (N8988, N8979, N6592);
buf BUF1 (N8989, N8982);
or OR4 (N8990, N8981, N5474, N4953, N7837);
xor XOR2 (N8991, N8987, N3072);
buf BUF1 (N8992, N8990);
nor NOR2 (N8993, N8985, N7003);
or OR3 (N8994, N8989, N6461, N2552);
nor NOR3 (N8995, N8963, N5012, N2926);
and AND2 (N8996, N8984, N814);
not NOT1 (N8997, N8971);
xor XOR2 (N8998, N8967, N4978);
not NOT1 (N8999, N8996);
and AND2 (N9000, N8994, N1268);
and AND4 (N9001, N8999, N2505, N8786, N8179);
or OR2 (N9002, N8993, N3161);
buf BUF1 (N9003, N9000);
and AND4 (N9004, N8986, N6898, N4341, N3289);
nor NOR3 (N9005, N9001, N3225, N829);
not NOT1 (N9006, N9002);
nor NOR4 (N9007, N8995, N2368, N472, N1375);
xor XOR2 (N9008, N9004, N8409);
xor XOR2 (N9009, N9008, N6078);
nor NOR2 (N9010, N9006, N3251);
nand NAND2 (N9011, N8988, N7677);
or OR3 (N9012, N9009, N242, N6018);
xor XOR2 (N9013, N8998, N2182);
and AND4 (N9014, N9012, N1859, N3375, N5592);
nor NOR2 (N9015, N9010, N4572);
or OR2 (N9016, N9003, N3251);
or OR4 (N9017, N9016, N2522, N6404, N1910);
nand NAND3 (N9018, N8991, N8388, N7990);
and AND2 (N9019, N9005, N709);
not NOT1 (N9020, N9017);
and AND3 (N9021, N9013, N5479, N3566);
buf BUF1 (N9022, N9020);
nor NOR3 (N9023, N9018, N6198, N3462);
or OR2 (N9024, N9014, N3714);
nor NOR2 (N9025, N9019, N3126);
buf BUF1 (N9026, N9015);
buf BUF1 (N9027, N9007);
buf BUF1 (N9028, N9022);
or OR2 (N9029, N9027, N4080);
nand NAND4 (N9030, N9024, N3711, N7548, N4969);
xor XOR2 (N9031, N9029, N8348);
and AND2 (N9032, N9031, N7151);
or OR3 (N9033, N9030, N7927, N8689);
buf BUF1 (N9034, N9033);
or OR3 (N9035, N9034, N2604, N1902);
and AND2 (N9036, N9026, N7993);
and AND4 (N9037, N8997, N8341, N6568, N1818);
xor XOR2 (N9038, N9032, N1624);
or OR2 (N9039, N9025, N8147);
or OR4 (N9040, N9038, N7903, N8236, N3406);
nor NOR3 (N9041, N9011, N5039, N4553);
nor NOR2 (N9042, N9021, N522);
not NOT1 (N9043, N8992);
and AND3 (N9044, N9041, N28, N1837);
not NOT1 (N9045, N9043);
buf BUF1 (N9046, N9036);
not NOT1 (N9047, N9035);
not NOT1 (N9048, N9042);
xor XOR2 (N9049, N9040, N5180);
or OR2 (N9050, N9037, N1173);
xor XOR2 (N9051, N9039, N6729);
or OR2 (N9052, N9050, N7160);
xor XOR2 (N9053, N9028, N1469);
buf BUF1 (N9054, N9045);
nand NAND2 (N9055, N9046, N3672);
and AND4 (N9056, N9049, N285, N5323, N3688);
not NOT1 (N9057, N9056);
and AND4 (N9058, N9052, N2994, N2375, N2365);
xor XOR2 (N9059, N9051, N1785);
xor XOR2 (N9060, N9057, N2299);
and AND3 (N9061, N9053, N1860, N8044);
or OR3 (N9062, N9061, N8797, N5544);
not NOT1 (N9063, N9048);
nand NAND2 (N9064, N9063, N8730);
not NOT1 (N9065, N9054);
nand NAND4 (N9066, N9060, N4504, N1841, N4133);
nand NAND4 (N9067, N9044, N5644, N1076, N7057);
nand NAND4 (N9068, N9067, N2745, N3314, N4643);
nand NAND2 (N9069, N9065, N5052);
or OR3 (N9070, N9064, N2584, N7981);
or OR2 (N9071, N9059, N7383);
or OR2 (N9072, N9062, N3427);
nor NOR2 (N9073, N9072, N1529);
buf BUF1 (N9074, N9058);
buf BUF1 (N9075, N9068);
nor NOR3 (N9076, N9069, N7543, N3934);
buf BUF1 (N9077, N9071);
xor XOR2 (N9078, N9066, N7893);
nand NAND4 (N9079, N9070, N3652, N1716, N1892);
not NOT1 (N9080, N9077);
not NOT1 (N9081, N9075);
xor XOR2 (N9082, N9074, N7274);
buf BUF1 (N9083, N9079);
buf BUF1 (N9084, N9023);
nand NAND2 (N9085, N9080, N988);
xor XOR2 (N9086, N9073, N7025);
and AND2 (N9087, N9076, N3495);
and AND3 (N9088, N9055, N8856, N3158);
buf BUF1 (N9089, N9082);
or OR4 (N9090, N9087, N3365, N6733, N1026);
xor XOR2 (N9091, N9090, N9);
nand NAND3 (N9092, N9091, N8431, N5571);
nor NOR2 (N9093, N9088, N1230);
xor XOR2 (N9094, N9078, N7562);
xor XOR2 (N9095, N9086, N7870);
nand NAND4 (N9096, N9093, N7360, N5937, N3962);
nor NOR3 (N9097, N9094, N1288, N1844);
not NOT1 (N9098, N9081);
not NOT1 (N9099, N9092);
not NOT1 (N9100, N9095);
nor NOR4 (N9101, N9098, N1264, N2628, N3969);
and AND3 (N9102, N9096, N6908, N3110);
xor XOR2 (N9103, N9099, N6558);
nand NAND4 (N9104, N9102, N2825, N4613, N6663);
buf BUF1 (N9105, N9083);
nor NOR2 (N9106, N9085, N2631);
nor NOR4 (N9107, N9100, N3212, N1352, N8424);
not NOT1 (N9108, N9047);
xor XOR2 (N9109, N9104, N3558);
xor XOR2 (N9110, N9106, N1663);
xor XOR2 (N9111, N9097, N2293);
not NOT1 (N9112, N9089);
buf BUF1 (N9113, N9105);
nor NOR4 (N9114, N9108, N6049, N6353, N970);
and AND4 (N9115, N9101, N3071, N6609, N4267);
or OR2 (N9116, N9114, N7129);
not NOT1 (N9117, N9112);
or OR2 (N9118, N9116, N1905);
or OR4 (N9119, N9103, N8685, N5723, N185);
buf BUF1 (N9120, N9084);
nor NOR2 (N9121, N9113, N4814);
nand NAND2 (N9122, N9117, N6058);
not NOT1 (N9123, N9110);
xor XOR2 (N9124, N9123, N135);
buf BUF1 (N9125, N9121);
nor NOR4 (N9126, N9119, N5261, N2875, N604);
xor XOR2 (N9127, N9122, N6806);
buf BUF1 (N9128, N9124);
buf BUF1 (N9129, N9118);
or OR4 (N9130, N9127, N7215, N8107, N5061);
not NOT1 (N9131, N9109);
nand NAND4 (N9132, N9129, N5161, N444, N2266);
or OR4 (N9133, N9131, N7257, N6129, N4974);
nor NOR2 (N9134, N9128, N1825);
nor NOR4 (N9135, N9133, N7091, N3115, N5670);
buf BUF1 (N9136, N9120);
not NOT1 (N9137, N9107);
nor NOR4 (N9138, N9111, N6158, N8542, N3645);
not NOT1 (N9139, N9132);
nor NOR3 (N9140, N9125, N1741, N2742);
nor NOR3 (N9141, N9135, N4711, N1408);
nand NAND2 (N9142, N9130, N216);
nor NOR4 (N9143, N9139, N3313, N1523, N7632);
not NOT1 (N9144, N9136);
nor NOR4 (N9145, N9126, N3126, N6276, N2628);
xor XOR2 (N9146, N9140, N7204);
not NOT1 (N9147, N9138);
or OR2 (N9148, N9146, N8461);
nand NAND3 (N9149, N9115, N5347, N1816);
not NOT1 (N9150, N9148);
not NOT1 (N9151, N9149);
nand NAND2 (N9152, N9150, N6420);
buf BUF1 (N9153, N9152);
nand NAND3 (N9154, N9147, N164, N6311);
and AND4 (N9155, N9153, N5372, N2831, N7455);
nand NAND4 (N9156, N9137, N15, N6151, N3243);
xor XOR2 (N9157, N9154, N4191);
xor XOR2 (N9158, N9134, N108);
not NOT1 (N9159, N9142);
not NOT1 (N9160, N9141);
nand NAND4 (N9161, N9144, N8474, N5505, N2883);
xor XOR2 (N9162, N9155, N4306);
nor NOR3 (N9163, N9143, N6990, N2634);
and AND4 (N9164, N9158, N2358, N5421, N5144);
or OR2 (N9165, N9163, N7496);
or OR4 (N9166, N9156, N5337, N3423, N4864);
not NOT1 (N9167, N9145);
or OR2 (N9168, N9167, N1858);
not NOT1 (N9169, N9157);
xor XOR2 (N9170, N9160, N7240);
nor NOR3 (N9171, N9170, N2894, N8316);
and AND4 (N9172, N9171, N1683, N2867, N912);
not NOT1 (N9173, N9164);
not NOT1 (N9174, N9168);
buf BUF1 (N9175, N9169);
or OR2 (N9176, N9162, N4585);
and AND4 (N9177, N9172, N5445, N4833, N389);
or OR4 (N9178, N9165, N8660, N2758, N8061);
nand NAND2 (N9179, N9176, N7217);
or OR3 (N9180, N9151, N628, N6566);
nor NOR4 (N9181, N9179, N675, N544, N3821);
and AND3 (N9182, N9173, N3466, N28);
nor NOR4 (N9183, N9175, N5940, N8865, N8612);
xor XOR2 (N9184, N9174, N8557);
nor NOR3 (N9185, N9178, N2402, N5551);
and AND2 (N9186, N9181, N7371);
buf BUF1 (N9187, N9180);
buf BUF1 (N9188, N9183);
nand NAND3 (N9189, N9185, N5680, N3714);
and AND3 (N9190, N9184, N1650, N6831);
and AND2 (N9191, N9177, N8363);
nor NOR3 (N9192, N9182, N1684, N6165);
and AND4 (N9193, N9192, N6506, N3059, N8658);
or OR2 (N9194, N9191, N953);
and AND3 (N9195, N9189, N1625, N4226);
not NOT1 (N9196, N9195);
buf BUF1 (N9197, N9188);
or OR4 (N9198, N9186, N4653, N2241, N5367);
nand NAND3 (N9199, N9159, N1100, N3736);
nand NAND4 (N9200, N9190, N8102, N4566, N3974);
or OR3 (N9201, N9200, N7939, N175);
xor XOR2 (N9202, N9198, N6071);
and AND4 (N9203, N9187, N616, N7306, N2922);
xor XOR2 (N9204, N9203, N2163);
nor NOR2 (N9205, N9161, N2334);
and AND2 (N9206, N9197, N3400);
buf BUF1 (N9207, N9202);
xor XOR2 (N9208, N9205, N2612);
nand NAND3 (N9209, N9194, N5040, N7396);
nand NAND4 (N9210, N9208, N3595, N1961, N3612);
nand NAND3 (N9211, N9206, N7534, N7773);
not NOT1 (N9212, N9166);
not NOT1 (N9213, N9211);
xor XOR2 (N9214, N9207, N4731);
xor XOR2 (N9215, N9199, N6480);
or OR4 (N9216, N9196, N2351, N5994, N4129);
or OR2 (N9217, N9209, N8076);
not NOT1 (N9218, N9204);
xor XOR2 (N9219, N9218, N6358);
buf BUF1 (N9220, N9201);
xor XOR2 (N9221, N9220, N4911);
or OR4 (N9222, N9193, N2301, N7582, N2528);
nor NOR2 (N9223, N9210, N5305);
nor NOR2 (N9224, N9219, N8141);
or OR2 (N9225, N9224, N6576);
xor XOR2 (N9226, N9223, N3718);
or OR2 (N9227, N9216, N2557);
not NOT1 (N9228, N9212);
xor XOR2 (N9229, N9214, N8237);
and AND3 (N9230, N9225, N3706, N2060);
nand NAND2 (N9231, N9217, N4895);
buf BUF1 (N9232, N9221);
nor NOR4 (N9233, N9228, N8673, N4407, N8718);
and AND2 (N9234, N9222, N6722);
and AND2 (N9235, N9233, N8449);
not NOT1 (N9236, N9231);
nor NOR3 (N9237, N9236, N9042, N8421);
buf BUF1 (N9238, N9229);
not NOT1 (N9239, N9234);
or OR2 (N9240, N9238, N6479);
xor XOR2 (N9241, N9227, N2569);
or OR4 (N9242, N9230, N7479, N8848, N3470);
not NOT1 (N9243, N9235);
or OR2 (N9244, N9215, N8414);
buf BUF1 (N9245, N9240);
nor NOR2 (N9246, N9239, N7940);
or OR4 (N9247, N9241, N4159, N2297, N5734);
buf BUF1 (N9248, N9242);
nor NOR2 (N9249, N9248, N838);
buf BUF1 (N9250, N9213);
buf BUF1 (N9251, N9250);
nand NAND4 (N9252, N9247, N2420, N1896, N5127);
nand NAND3 (N9253, N9249, N6497, N8449);
and AND3 (N9254, N9252, N7591, N4313);
xor XOR2 (N9255, N9246, N5900);
buf BUF1 (N9256, N9254);
buf BUF1 (N9257, N9256);
nor NOR2 (N9258, N9232, N5287);
or OR2 (N9259, N9226, N3139);
not NOT1 (N9260, N9258);
or OR3 (N9261, N9251, N5251, N7153);
and AND2 (N9262, N9245, N3342);
nand NAND4 (N9263, N9244, N2977, N1437, N6979);
not NOT1 (N9264, N9237);
nand NAND2 (N9265, N9263, N949);
nor NOR2 (N9266, N9255, N6031);
not NOT1 (N9267, N9266);
not NOT1 (N9268, N9259);
not NOT1 (N9269, N9268);
nor NOR3 (N9270, N9253, N8423, N1433);
or OR2 (N9271, N9264, N5759);
xor XOR2 (N9272, N9262, N4069);
xor XOR2 (N9273, N9269, N1105);
buf BUF1 (N9274, N9267);
buf BUF1 (N9275, N9261);
and AND4 (N9276, N9274, N9013, N568, N6420);
buf BUF1 (N9277, N9273);
not NOT1 (N9278, N9260);
nor NOR2 (N9279, N9278, N200);
nand NAND2 (N9280, N9277, N7106);
buf BUF1 (N9281, N9275);
or OR3 (N9282, N9257, N5957, N6947);
or OR4 (N9283, N9276, N6962, N3944, N5304);
buf BUF1 (N9284, N9271);
not NOT1 (N9285, N9283);
not NOT1 (N9286, N9270);
xor XOR2 (N9287, N9285, N712);
or OR3 (N9288, N9265, N571, N3833);
nand NAND2 (N9289, N9287, N6536);
buf BUF1 (N9290, N9272);
nand NAND4 (N9291, N9288, N4560, N4233, N4698);
or OR2 (N9292, N9280, N7801);
nand NAND2 (N9293, N9279, N954);
nand NAND4 (N9294, N9291, N5481, N5018, N8035);
nor NOR2 (N9295, N9289, N9111);
or OR4 (N9296, N9293, N7903, N7112, N5185);
not NOT1 (N9297, N9286);
xor XOR2 (N9298, N9297, N988);
nor NOR2 (N9299, N9243, N4624);
buf BUF1 (N9300, N9292);
buf BUF1 (N9301, N9281);
nor NOR4 (N9302, N9282, N5439, N3931, N5386);
or OR4 (N9303, N9295, N3505, N4742, N5191);
nand NAND2 (N9304, N9290, N3695);
buf BUF1 (N9305, N9303);
or OR2 (N9306, N9296, N5330);
or OR4 (N9307, N9298, N6059, N6946, N6499);
buf BUF1 (N9308, N9305);
xor XOR2 (N9309, N9300, N8654);
nor NOR2 (N9310, N9304, N8553);
or OR3 (N9311, N9284, N668, N2067);
buf BUF1 (N9312, N9310);
nor NOR2 (N9313, N9302, N1131);
nor NOR3 (N9314, N9301, N2399, N6064);
buf BUF1 (N9315, N9294);
not NOT1 (N9316, N9313);
nor NOR3 (N9317, N9315, N9046, N2953);
nand NAND4 (N9318, N9306, N6213, N6420, N1341);
xor XOR2 (N9319, N9299, N8306);
and AND2 (N9320, N9309, N1773);
or OR3 (N9321, N9307, N5203, N3635);
nor NOR3 (N9322, N9321, N2741, N5000);
and AND2 (N9323, N9318, N3640);
buf BUF1 (N9324, N9317);
or OR3 (N9325, N9312, N7780, N865);
or OR2 (N9326, N9311, N6448);
nor NOR3 (N9327, N9324, N2867, N5977);
buf BUF1 (N9328, N9308);
nand NAND2 (N9329, N9316, N2109);
xor XOR2 (N9330, N9323, N6312);
or OR4 (N9331, N9326, N825, N8360, N3964);
not NOT1 (N9332, N9327);
xor XOR2 (N9333, N9320, N2422);
or OR3 (N9334, N9330, N7136, N4795);
and AND2 (N9335, N9331, N4492);
and AND2 (N9336, N9319, N5657);
and AND4 (N9337, N9328, N6395, N3969, N2079);
xor XOR2 (N9338, N9322, N3960);
not NOT1 (N9339, N9335);
xor XOR2 (N9340, N9332, N7339);
nor NOR3 (N9341, N9340, N9318, N4031);
nor NOR4 (N9342, N9329, N4984, N4313, N6117);
or OR4 (N9343, N9342, N1450, N7953, N471);
buf BUF1 (N9344, N9333);
nand NAND3 (N9345, N9343, N4648, N8018);
buf BUF1 (N9346, N9338);
or OR4 (N9347, N9345, N7322, N5638, N7667);
nor NOR3 (N9348, N9337, N188, N8774);
buf BUF1 (N9349, N9339);
or OR3 (N9350, N9334, N2996, N1864);
buf BUF1 (N9351, N9336);
not NOT1 (N9352, N9348);
nor NOR3 (N9353, N9314, N1622, N7822);
not NOT1 (N9354, N9349);
or OR3 (N9355, N9347, N3236, N4243);
nand NAND3 (N9356, N9352, N3772, N6472);
and AND3 (N9357, N9325, N4568, N8414);
or OR4 (N9358, N9355, N6826, N9237, N4348);
nand NAND3 (N9359, N9346, N5414, N4568);
or OR4 (N9360, N9354, N7997, N4014, N7680);
not NOT1 (N9361, N9353);
buf BUF1 (N9362, N9359);
nor NOR4 (N9363, N9360, N9071, N6836, N5886);
xor XOR2 (N9364, N9341, N6962);
or OR2 (N9365, N9350, N6839);
nand NAND3 (N9366, N9358, N2370, N5978);
nand NAND4 (N9367, N9361, N183, N5275, N8761);
nor NOR3 (N9368, N9356, N1338, N6076);
nand NAND3 (N9369, N9351, N212, N8312);
nor NOR3 (N9370, N9366, N5140, N4968);
xor XOR2 (N9371, N9368, N4873);
buf BUF1 (N9372, N9371);
xor XOR2 (N9373, N9370, N1512);
nand NAND4 (N9374, N9362, N5966, N6883, N8800);
and AND2 (N9375, N9357, N7198);
buf BUF1 (N9376, N9372);
buf BUF1 (N9377, N9374);
nand NAND2 (N9378, N9373, N4115);
buf BUF1 (N9379, N9365);
and AND4 (N9380, N9377, N8447, N4199, N1827);
or OR4 (N9381, N9380, N4096, N7406, N3415);
buf BUF1 (N9382, N9379);
or OR3 (N9383, N9367, N243, N985);
or OR4 (N9384, N9381, N5195, N1801, N8855);
buf BUF1 (N9385, N9344);
nand NAND4 (N9386, N9378, N4805, N8386, N801);
xor XOR2 (N9387, N9384, N4098);
or OR4 (N9388, N9369, N2647, N7202, N5945);
and AND2 (N9389, N9383, N5813);
nor NOR3 (N9390, N9389, N8669, N4700);
nor NOR3 (N9391, N9387, N798, N3830);
and AND4 (N9392, N9391, N5028, N5227, N5121);
not NOT1 (N9393, N9364);
xor XOR2 (N9394, N9388, N8580);
and AND4 (N9395, N9392, N8879, N6031, N7237);
buf BUF1 (N9396, N9393);
nand NAND3 (N9397, N9390, N8503, N2241);
not NOT1 (N9398, N9394);
and AND3 (N9399, N9386, N8006, N1085);
or OR3 (N9400, N9399, N4039, N2463);
or OR2 (N9401, N9376, N8198);
xor XOR2 (N9402, N9395, N4246);
or OR4 (N9403, N9396, N3618, N5995, N3529);
and AND2 (N9404, N9397, N8846);
buf BUF1 (N9405, N9363);
or OR4 (N9406, N9382, N5626, N778, N2035);
and AND4 (N9407, N9385, N8119, N5251, N37);
and AND2 (N9408, N9407, N4117);
or OR3 (N9409, N9403, N7799, N8371);
xor XOR2 (N9410, N9400, N6226);
xor XOR2 (N9411, N9406, N1498);
not NOT1 (N9412, N9405);
or OR3 (N9413, N9411, N5444, N5951);
xor XOR2 (N9414, N9412, N8836);
and AND3 (N9415, N9404, N3286, N86);
nor NOR3 (N9416, N9375, N4325, N7327);
and AND4 (N9417, N9413, N8137, N2954, N6255);
and AND4 (N9418, N9398, N3557, N9298, N8199);
and AND2 (N9419, N9414, N1852);
xor XOR2 (N9420, N9401, N6908);
xor XOR2 (N9421, N9409, N8468);
nand NAND2 (N9422, N9421, N3500);
not NOT1 (N9423, N9402);
buf BUF1 (N9424, N9408);
nor NOR4 (N9425, N9423, N1694, N2029, N6295);
or OR4 (N9426, N9420, N4122, N3972, N798);
buf BUF1 (N9427, N9415);
nor NOR4 (N9428, N9422, N2799, N6231, N3507);
nor NOR2 (N9429, N9425, N7459);
and AND2 (N9430, N9419, N351);
nor NOR2 (N9431, N9429, N3543);
xor XOR2 (N9432, N9431, N4348);
xor XOR2 (N9433, N9417, N498);
nor NOR2 (N9434, N9424, N8615);
nand NAND4 (N9435, N9418, N2645, N2921, N4613);
buf BUF1 (N9436, N9433);
buf BUF1 (N9437, N9432);
and AND4 (N9438, N9434, N7922, N1462, N2585);
and AND4 (N9439, N9410, N4851, N5002, N5533);
or OR3 (N9440, N9427, N1739, N4487);
and AND3 (N9441, N9435, N7151, N5234);
xor XOR2 (N9442, N9416, N2904);
nand NAND3 (N9443, N9437, N7876, N1901);
nor NOR2 (N9444, N9426, N5671);
nor NOR4 (N9445, N9441, N9059, N1996, N4841);
buf BUF1 (N9446, N9439);
nand NAND4 (N9447, N9430, N3155, N7549, N8607);
xor XOR2 (N9448, N9436, N5148);
or OR3 (N9449, N9445, N8096, N5865);
xor XOR2 (N9450, N9447, N3378);
not NOT1 (N9451, N9438);
xor XOR2 (N9452, N9444, N7157);
and AND3 (N9453, N9428, N4426, N1537);
nand NAND2 (N9454, N9448, N3482);
buf BUF1 (N9455, N9451);
and AND2 (N9456, N9453, N7658);
or OR3 (N9457, N9454, N1424, N645);
nand NAND3 (N9458, N9449, N4565, N7522);
xor XOR2 (N9459, N9455, N5416);
buf BUF1 (N9460, N9459);
buf BUF1 (N9461, N9446);
nand NAND3 (N9462, N9443, N7937, N4819);
nand NAND3 (N9463, N9442, N8216, N6730);
buf BUF1 (N9464, N9440);
buf BUF1 (N9465, N9463);
nor NOR3 (N9466, N9450, N1297, N5641);
and AND3 (N9467, N9456, N5210, N2404);
or OR3 (N9468, N9465, N6094, N7752);
buf BUF1 (N9469, N9461);
or OR3 (N9470, N9460, N7003, N4116);
and AND2 (N9471, N9458, N4299);
nand NAND2 (N9472, N9470, N8747);
nor NOR4 (N9473, N9471, N1828, N7532, N95);
or OR2 (N9474, N9467, N3539);
buf BUF1 (N9475, N9469);
nand NAND4 (N9476, N9457, N1745, N42, N6507);
xor XOR2 (N9477, N9462, N2166);
xor XOR2 (N9478, N9477, N3481);
and AND4 (N9479, N9478, N4071, N7395, N403);
and AND2 (N9480, N9468, N4086);
buf BUF1 (N9481, N9473);
nand NAND4 (N9482, N9474, N1118, N6840, N823);
nor NOR4 (N9483, N9480, N8117, N3753, N5864);
nand NAND4 (N9484, N9483, N7407, N8643, N8410);
buf BUF1 (N9485, N9466);
and AND4 (N9486, N9484, N7819, N1462, N7687);
not NOT1 (N9487, N9452);
not NOT1 (N9488, N9464);
nand NAND2 (N9489, N9482, N13);
and AND2 (N9490, N9479, N7279);
xor XOR2 (N9491, N9488, N3467);
buf BUF1 (N9492, N9487);
xor XOR2 (N9493, N9492, N2753);
buf BUF1 (N9494, N9472);
and AND4 (N9495, N9485, N466, N7308, N4287);
nand NAND3 (N9496, N9495, N4297, N2486);
and AND2 (N9497, N9486, N4967);
xor XOR2 (N9498, N9491, N1483);
nand NAND4 (N9499, N9481, N2352, N730, N2336);
and AND3 (N9500, N9493, N7292, N4004);
xor XOR2 (N9501, N9489, N8386);
and AND4 (N9502, N9497, N9105, N6021, N7155);
buf BUF1 (N9503, N9499);
not NOT1 (N9504, N9500);
buf BUF1 (N9505, N9504);
buf BUF1 (N9506, N9498);
xor XOR2 (N9507, N9503, N8961);
nor NOR3 (N9508, N9496, N2069, N5668);
nand NAND3 (N9509, N9507, N9192, N8944);
xor XOR2 (N9510, N9501, N5980);
nor NOR3 (N9511, N9490, N6603, N4351);
and AND4 (N9512, N9510, N243, N9394, N8342);
and AND3 (N9513, N9494, N4961, N1068);
buf BUF1 (N9514, N9509);
xor XOR2 (N9515, N9514, N7393);
or OR4 (N9516, N9511, N3962, N3726, N279);
xor XOR2 (N9517, N9508, N1866);
nor NOR2 (N9518, N9506, N4415);
xor XOR2 (N9519, N9513, N5837);
nand NAND2 (N9520, N9476, N4430);
nor NOR3 (N9521, N9475, N2728, N1450);
nand NAND3 (N9522, N9505, N8823, N2222);
xor XOR2 (N9523, N9512, N5770);
buf BUF1 (N9524, N9516);
nand NAND2 (N9525, N9520, N6807);
and AND2 (N9526, N9518, N8592);
and AND4 (N9527, N9519, N7739, N2879, N6480);
xor XOR2 (N9528, N9521, N4964);
nand NAND2 (N9529, N9527, N1585);
nor NOR3 (N9530, N9524, N1608, N5996);
not NOT1 (N9531, N9515);
xor XOR2 (N9532, N9526, N1882);
nor NOR4 (N9533, N9532, N8394, N6928, N4193);
nand NAND3 (N9534, N9533, N2726, N7209);
and AND4 (N9535, N9529, N7053, N745, N3512);
nor NOR2 (N9536, N9522, N4737);
or OR4 (N9537, N9525, N9460, N3600, N4324);
nor NOR2 (N9538, N9536, N1060);
or OR3 (N9539, N9534, N423, N9112);
buf BUF1 (N9540, N9531);
buf BUF1 (N9541, N9528);
and AND2 (N9542, N9538, N2861);
and AND3 (N9543, N9535, N4439, N8770);
and AND4 (N9544, N9523, N6995, N5637, N4688);
buf BUF1 (N9545, N9544);
and AND4 (N9546, N9540, N1757, N7459, N5152);
not NOT1 (N9547, N9541);
xor XOR2 (N9548, N9545, N4569);
or OR4 (N9549, N9548, N1547, N1380, N3039);
and AND3 (N9550, N9549, N3832, N2797);
nor NOR4 (N9551, N9502, N1921, N2861, N5318);
or OR2 (N9552, N9546, N7406);
nor NOR4 (N9553, N9539, N8014, N7342, N109);
buf BUF1 (N9554, N9553);
xor XOR2 (N9555, N9517, N3293);
not NOT1 (N9556, N9537);
not NOT1 (N9557, N9552);
nand NAND2 (N9558, N9542, N6561);
not NOT1 (N9559, N9554);
nor NOR3 (N9560, N9551, N5854, N2436);
or OR4 (N9561, N9556, N4816, N3771, N8479);
buf BUF1 (N9562, N9543);
xor XOR2 (N9563, N9558, N3868);
nor NOR4 (N9564, N9560, N5955, N2726, N3727);
nor NOR4 (N9565, N9563, N5835, N5206, N3655);
buf BUF1 (N9566, N9565);
not NOT1 (N9567, N9547);
xor XOR2 (N9568, N9559, N9038);
xor XOR2 (N9569, N9567, N2892);
nand NAND4 (N9570, N9566, N6049, N1562, N4942);
nand NAND2 (N9571, N9569, N36);
and AND3 (N9572, N9562, N2351, N3780);
buf BUF1 (N9573, N9564);
nand NAND3 (N9574, N9571, N9085, N5978);
or OR2 (N9575, N9561, N8332);
not NOT1 (N9576, N9568);
not NOT1 (N9577, N9572);
and AND2 (N9578, N9550, N5385);
and AND4 (N9579, N9576, N609, N4151, N752);
nand NAND2 (N9580, N9557, N3227);
nand NAND4 (N9581, N9578, N9184, N1355, N3721);
not NOT1 (N9582, N9575);
or OR2 (N9583, N9570, N8700);
and AND3 (N9584, N9583, N2958, N552);
xor XOR2 (N9585, N9574, N1915);
buf BUF1 (N9586, N9555);
and AND3 (N9587, N9586, N4938, N6026);
or OR4 (N9588, N9581, N3924, N2331, N6101);
nand NAND2 (N9589, N9579, N8976);
buf BUF1 (N9590, N9530);
xor XOR2 (N9591, N9573, N1562);
or OR3 (N9592, N9585, N8057, N495);
or OR2 (N9593, N9589, N7429);
and AND4 (N9594, N9580, N8378, N5213, N5698);
nor NOR2 (N9595, N9590, N8482);
buf BUF1 (N9596, N9594);
xor XOR2 (N9597, N9587, N6096);
and AND3 (N9598, N9595, N5099, N9072);
nor NOR4 (N9599, N9588, N8331, N3498, N313);
and AND4 (N9600, N9599, N6612, N6656, N6276);
nor NOR3 (N9601, N9600, N2956, N7920);
buf BUF1 (N9602, N9596);
or OR4 (N9603, N9597, N6020, N7606, N3382);
nor NOR2 (N9604, N9577, N5036);
not NOT1 (N9605, N9584);
or OR3 (N9606, N9598, N3185, N2929);
not NOT1 (N9607, N9593);
nor NOR3 (N9608, N9603, N947, N3624);
or OR4 (N9609, N9591, N1399, N7815, N8686);
nor NOR4 (N9610, N9604, N444, N904, N2362);
and AND4 (N9611, N9608, N9153, N1835, N2557);
xor XOR2 (N9612, N9601, N5186);
not NOT1 (N9613, N9582);
or OR2 (N9614, N9606, N6242);
not NOT1 (N9615, N9614);
not NOT1 (N9616, N9611);
nor NOR2 (N9617, N9609, N5622);
nor NOR4 (N9618, N9605, N1958, N5161, N1109);
not NOT1 (N9619, N9607);
and AND4 (N9620, N9612, N5748, N3294, N3488);
xor XOR2 (N9621, N9602, N1654);
buf BUF1 (N9622, N9616);
nand NAND3 (N9623, N9622, N4881, N210);
not NOT1 (N9624, N9621);
buf BUF1 (N9625, N9624);
not NOT1 (N9626, N9625);
nor NOR4 (N9627, N9618, N7896, N4768, N3920);
buf BUF1 (N9628, N9617);
not NOT1 (N9629, N9619);
or OR3 (N9630, N9628, N8319, N186);
nor NOR2 (N9631, N9630, N9478);
nand NAND3 (N9632, N9592, N395, N839);
not NOT1 (N9633, N9620);
not NOT1 (N9634, N9623);
xor XOR2 (N9635, N9629, N6657);
nor NOR2 (N9636, N9613, N9304);
xor XOR2 (N9637, N9632, N5281);
not NOT1 (N9638, N9634);
nor NOR2 (N9639, N9633, N5546);
buf BUF1 (N9640, N9627);
nor NOR4 (N9641, N9638, N5263, N8677, N9095);
or OR4 (N9642, N9640, N3356, N3112, N8930);
not NOT1 (N9643, N9642);
and AND3 (N9644, N9639, N2423, N7376);
and AND2 (N9645, N9643, N4866);
not NOT1 (N9646, N9645);
buf BUF1 (N9647, N9615);
and AND4 (N9648, N9646, N3871, N6736, N7465);
or OR2 (N9649, N9647, N845);
or OR4 (N9650, N9649, N1285, N3838, N7539);
nor NOR4 (N9651, N9635, N3685, N6850, N910);
not NOT1 (N9652, N9610);
nand NAND3 (N9653, N9652, N4130, N6366);
xor XOR2 (N9654, N9648, N8021);
nand NAND2 (N9655, N9650, N4108);
not NOT1 (N9656, N9644);
not NOT1 (N9657, N9655);
buf BUF1 (N9658, N9631);
nor NOR4 (N9659, N9653, N1902, N2593, N3484);
buf BUF1 (N9660, N9654);
and AND3 (N9661, N9658, N5388, N6507);
and AND3 (N9662, N9660, N8516, N952);
or OR4 (N9663, N9637, N2115, N8739, N1177);
and AND3 (N9664, N9661, N4713, N1035);
and AND4 (N9665, N9662, N8710, N2391, N5899);
buf BUF1 (N9666, N9665);
not NOT1 (N9667, N9659);
nor NOR3 (N9668, N9667, N8578, N2134);
and AND3 (N9669, N9663, N9371, N7459);
buf BUF1 (N9670, N9657);
or OR3 (N9671, N9641, N9073, N2055);
xor XOR2 (N9672, N9656, N9491);
xor XOR2 (N9673, N9668, N6827);
buf BUF1 (N9674, N9636);
nand NAND4 (N9675, N9666, N3957, N3656, N9564);
or OR2 (N9676, N9664, N4572);
nor NOR2 (N9677, N9671, N4918);
nand NAND3 (N9678, N9669, N5905, N2286);
buf BUF1 (N9679, N9626);
nor NOR3 (N9680, N9672, N5149, N7892);
not NOT1 (N9681, N9677);
buf BUF1 (N9682, N9680);
and AND2 (N9683, N9678, N3392);
or OR4 (N9684, N9682, N8202, N20, N1964);
not NOT1 (N9685, N9684);
and AND4 (N9686, N9676, N5458, N5947, N5358);
xor XOR2 (N9687, N9679, N9173);
nor NOR3 (N9688, N9675, N9249, N546);
xor XOR2 (N9689, N9688, N4915);
not NOT1 (N9690, N9670);
and AND4 (N9691, N9651, N4045, N3627, N8787);
not NOT1 (N9692, N9686);
nand NAND2 (N9693, N9674, N4984);
buf BUF1 (N9694, N9681);
not NOT1 (N9695, N9693);
or OR2 (N9696, N9687, N47);
or OR2 (N9697, N9690, N399);
and AND4 (N9698, N9685, N1626, N5574, N4605);
nor NOR3 (N9699, N9694, N7027, N836);
and AND4 (N9700, N9691, N4376, N5545, N5092);
xor XOR2 (N9701, N9692, N3785);
buf BUF1 (N9702, N9673);
nand NAND4 (N9703, N9683, N5071, N9059, N9048);
buf BUF1 (N9704, N9696);
and AND2 (N9705, N9698, N8180);
nor NOR4 (N9706, N9704, N7819, N6377, N3430);
or OR3 (N9707, N9700, N6499, N5306);
or OR2 (N9708, N9689, N7259);
buf BUF1 (N9709, N9699);
buf BUF1 (N9710, N9701);
nor NOR4 (N9711, N9709, N2290, N3511, N1148);
buf BUF1 (N9712, N9703);
not NOT1 (N9713, N9705);
or OR3 (N9714, N9708, N5725, N6471);
not NOT1 (N9715, N9706);
nor NOR4 (N9716, N9715, N1120, N7437, N5599);
buf BUF1 (N9717, N9716);
nor NOR3 (N9718, N9714, N5978, N3333);
xor XOR2 (N9719, N9710, N8203);
buf BUF1 (N9720, N9718);
or OR3 (N9721, N9711, N2515, N4003);
buf BUF1 (N9722, N9713);
nand NAND4 (N9723, N9719, N3429, N6220, N1784);
and AND4 (N9724, N9707, N4029, N734, N3243);
not NOT1 (N9725, N9702);
xor XOR2 (N9726, N9695, N2931);
or OR3 (N9727, N9725, N5832, N4215);
or OR2 (N9728, N9720, N4117);
xor XOR2 (N9729, N9712, N9448);
and AND3 (N9730, N9717, N4151, N6038);
xor XOR2 (N9731, N9728, N125);
xor XOR2 (N9732, N9722, N8570);
or OR2 (N9733, N9723, N3583);
nor NOR2 (N9734, N9732, N2155);
nor NOR2 (N9735, N9724, N8810);
nand NAND3 (N9736, N9721, N56, N1348);
nor NOR4 (N9737, N9729, N1658, N8017, N933);
or OR4 (N9738, N9736, N5424, N7050, N3202);
and AND2 (N9739, N9697, N9663);
and AND4 (N9740, N9733, N6184, N4961, N9212);
nor NOR2 (N9741, N9727, N1473);
or OR3 (N9742, N9740, N8869, N388);
nor NOR3 (N9743, N9735, N7798, N8124);
nor NOR2 (N9744, N9731, N756);
or OR3 (N9745, N9743, N418, N9480);
buf BUF1 (N9746, N9739);
and AND3 (N9747, N9744, N7991, N5447);
or OR2 (N9748, N9742, N481);
or OR2 (N9749, N9726, N9363);
xor XOR2 (N9750, N9730, N8825);
or OR4 (N9751, N9738, N7796, N3493, N1382);
xor XOR2 (N9752, N9749, N2974);
xor XOR2 (N9753, N9748, N1600);
nor NOR2 (N9754, N9746, N77);
nand NAND2 (N9755, N9741, N7269);
not NOT1 (N9756, N9745);
buf BUF1 (N9757, N9737);
or OR4 (N9758, N9750, N4117, N4441, N8803);
buf BUF1 (N9759, N9756);
or OR4 (N9760, N9747, N726, N9638, N6515);
not NOT1 (N9761, N9754);
not NOT1 (N9762, N9760);
xor XOR2 (N9763, N9752, N4882);
nand NAND2 (N9764, N9762, N1130);
nand NAND3 (N9765, N9755, N8707, N5266);
and AND4 (N9766, N9751, N8300, N4638, N4817);
nand NAND4 (N9767, N9761, N7078, N6023, N353);
nor NOR2 (N9768, N9764, N2572);
buf BUF1 (N9769, N9763);
buf BUF1 (N9770, N9768);
nand NAND4 (N9771, N9769, N7629, N4546, N2232);
nand NAND4 (N9772, N9767, N9695, N163, N423);
buf BUF1 (N9773, N9753);
or OR3 (N9774, N9765, N7917, N981);
buf BUF1 (N9775, N9772);
nand NAND4 (N9776, N9774, N4354, N8156, N6562);
xor XOR2 (N9777, N9776, N4352);
nor NOR2 (N9778, N9777, N2014);
and AND2 (N9779, N9734, N1656);
or OR2 (N9780, N9771, N5089);
buf BUF1 (N9781, N9780);
buf BUF1 (N9782, N9773);
nand NAND4 (N9783, N9766, N3960, N6996, N1686);
nor NOR2 (N9784, N9781, N5533);
xor XOR2 (N9785, N9778, N6324);
buf BUF1 (N9786, N9784);
not NOT1 (N9787, N9786);
not NOT1 (N9788, N9782);
or OR3 (N9789, N9787, N8808, N8003);
and AND2 (N9790, N9775, N160);
not NOT1 (N9791, N9790);
not NOT1 (N9792, N9783);
and AND3 (N9793, N9788, N1015, N608);
buf BUF1 (N9794, N9757);
nor NOR2 (N9795, N9785, N5514);
nor NOR2 (N9796, N9789, N8693);
buf BUF1 (N9797, N9759);
or OR3 (N9798, N9797, N646, N4739);
not NOT1 (N9799, N9793);
or OR2 (N9800, N9798, N2938);
nand NAND2 (N9801, N9792, N3201);
or OR2 (N9802, N9801, N8315);
and AND3 (N9803, N9799, N6957, N8807);
buf BUF1 (N9804, N9779);
nand NAND3 (N9805, N9802, N9197, N9532);
not NOT1 (N9806, N9804);
not NOT1 (N9807, N9796);
xor XOR2 (N9808, N9803, N3461);
xor XOR2 (N9809, N9807, N3002);
not NOT1 (N9810, N9770);
nand NAND4 (N9811, N9806, N890, N3831, N1792);
and AND3 (N9812, N9811, N9298, N7047);
or OR2 (N9813, N9800, N2577);
nand NAND3 (N9814, N9813, N4604, N4146);
nor NOR2 (N9815, N9810, N3906);
nor NOR2 (N9816, N9758, N4236);
xor XOR2 (N9817, N9794, N1113);
and AND2 (N9818, N9795, N4451);
and AND2 (N9819, N9814, N7078);
nand NAND2 (N9820, N9817, N4779);
buf BUF1 (N9821, N9820);
buf BUF1 (N9822, N9818);
and AND4 (N9823, N9821, N6919, N7779, N7519);
buf BUF1 (N9824, N9822);
xor XOR2 (N9825, N9816, N9358);
or OR3 (N9826, N9823, N7338, N5798);
nand NAND2 (N9827, N9819, N6226);
or OR4 (N9828, N9805, N2009, N4822, N4740);
buf BUF1 (N9829, N9809);
nand NAND4 (N9830, N9825, N9797, N3950, N6607);
and AND2 (N9831, N9812, N9783);
buf BUF1 (N9832, N9829);
xor XOR2 (N9833, N9831, N7666);
or OR2 (N9834, N9832, N3787);
nand NAND3 (N9835, N9830, N6949, N7640);
nor NOR3 (N9836, N9808, N3691, N9155);
nor NOR2 (N9837, N9827, N8177);
and AND2 (N9838, N9835, N4573);
and AND2 (N9839, N9833, N8350);
or OR2 (N9840, N9834, N4217);
nand NAND2 (N9841, N9840, N7911);
xor XOR2 (N9842, N9836, N3099);
xor XOR2 (N9843, N9841, N6173);
not NOT1 (N9844, N9838);
buf BUF1 (N9845, N9837);
buf BUF1 (N9846, N9842);
buf BUF1 (N9847, N9839);
nand NAND4 (N9848, N9791, N1076, N2486, N6088);
or OR4 (N9849, N9815, N9051, N9396, N2539);
or OR3 (N9850, N9844, N5659, N5345);
nand NAND4 (N9851, N9843, N9060, N1947, N7104);
nor NOR3 (N9852, N9848, N5708, N8);
not NOT1 (N9853, N9846);
nor NOR4 (N9854, N9849, N1471, N2478, N239);
buf BUF1 (N9855, N9828);
or OR3 (N9856, N9854, N7643, N9381);
not NOT1 (N9857, N9847);
buf BUF1 (N9858, N9856);
and AND4 (N9859, N9845, N3629, N3970, N1405);
nor NOR4 (N9860, N9853, N1894, N3623, N4154);
not NOT1 (N9861, N9852);
or OR2 (N9862, N9860, N1470);
nor NOR2 (N9863, N9858, N1941);
nor NOR4 (N9864, N9824, N2217, N6711, N8626);
not NOT1 (N9865, N9863);
not NOT1 (N9866, N9864);
or OR4 (N9867, N9859, N3828, N1232, N2189);
nor NOR4 (N9868, N9866, N9564, N5115, N4707);
buf BUF1 (N9869, N9865);
or OR4 (N9870, N9868, N3703, N4990, N3449);
not NOT1 (N9871, N9851);
xor XOR2 (N9872, N9855, N8900);
or OR4 (N9873, N9862, N7196, N5091, N9739);
or OR3 (N9874, N9871, N5085, N1076);
buf BUF1 (N9875, N9870);
and AND2 (N9876, N9850, N7088);
and AND4 (N9877, N9875, N3966, N7388, N5907);
buf BUF1 (N9878, N9872);
xor XOR2 (N9879, N9857, N564);
xor XOR2 (N9880, N9876, N6018);
buf BUF1 (N9881, N9873);
nor NOR2 (N9882, N9881, N2797);
or OR3 (N9883, N9878, N6582, N9106);
or OR2 (N9884, N9879, N1765);
nand NAND4 (N9885, N9874, N5046, N4837, N5909);
xor XOR2 (N9886, N9882, N9577);
and AND2 (N9887, N9867, N8355);
xor XOR2 (N9888, N9883, N4590);
nand NAND3 (N9889, N9888, N7452, N7867);
buf BUF1 (N9890, N9880);
nand NAND2 (N9891, N9884, N3833);
xor XOR2 (N9892, N9886, N5989);
or OR3 (N9893, N9889, N2839, N5708);
not NOT1 (N9894, N9887);
nand NAND2 (N9895, N9892, N9845);
nor NOR2 (N9896, N9895, N5699);
buf BUF1 (N9897, N9869);
or OR3 (N9898, N9877, N2742, N6889);
xor XOR2 (N9899, N9898, N8133);
and AND4 (N9900, N9890, N2690, N356, N3812);
and AND2 (N9901, N9896, N4613);
not NOT1 (N9902, N9885);
buf BUF1 (N9903, N9826);
xor XOR2 (N9904, N9861, N468);
xor XOR2 (N9905, N9899, N354);
buf BUF1 (N9906, N9894);
and AND4 (N9907, N9897, N7801, N9733, N3177);
and AND2 (N9908, N9904, N9742);
nor NOR3 (N9909, N9903, N4201, N5803);
nor NOR3 (N9910, N9909, N4320, N124);
nor NOR3 (N9911, N9910, N5569, N6175);
buf BUF1 (N9912, N9891);
nand NAND3 (N9913, N9900, N362, N8909);
and AND3 (N9914, N9907, N1808, N5080);
nor NOR3 (N9915, N9906, N5140, N4354);
buf BUF1 (N9916, N9913);
xor XOR2 (N9917, N9905, N3570);
xor XOR2 (N9918, N9911, N6880);
nor NOR4 (N9919, N9916, N2272, N5219, N4852);
not NOT1 (N9920, N9912);
not NOT1 (N9921, N9901);
xor XOR2 (N9922, N9917, N8487);
nand NAND3 (N9923, N9918, N8353, N7023);
xor XOR2 (N9924, N9919, N513);
and AND4 (N9925, N9915, N1162, N8606, N6979);
not NOT1 (N9926, N9921);
and AND4 (N9927, N9908, N5834, N1514, N9732);
buf BUF1 (N9928, N9922);
nor NOR3 (N9929, N9920, N7976, N3079);
and AND2 (N9930, N9927, N1665);
not NOT1 (N9931, N9930);
nor NOR4 (N9932, N9914, N1051, N8077, N5479);
not NOT1 (N9933, N9929);
nor NOR3 (N9934, N9931, N4618, N3592);
xor XOR2 (N9935, N9932, N1933);
nor NOR2 (N9936, N9902, N6727);
xor XOR2 (N9937, N9936, N4136);
nor NOR4 (N9938, N9926, N1820, N7087, N3859);
not NOT1 (N9939, N9924);
buf BUF1 (N9940, N9938);
nand NAND3 (N9941, N9925, N7307, N7330);
nand NAND3 (N9942, N9934, N8407, N5187);
not NOT1 (N9943, N9937);
or OR4 (N9944, N9933, N4816, N6565, N8820);
or OR3 (N9945, N9940, N8138, N2792);
and AND4 (N9946, N9941, N7333, N5721, N4216);
xor XOR2 (N9947, N9935, N944);
nor NOR3 (N9948, N9945, N5619, N8854);
nor NOR2 (N9949, N9923, N46);
or OR4 (N9950, N9893, N3720, N4952, N3258);
buf BUF1 (N9951, N9946);
buf BUF1 (N9952, N9928);
not NOT1 (N9953, N9944);
xor XOR2 (N9954, N9950, N671);
buf BUF1 (N9955, N9943);
or OR2 (N9956, N9947, N2489);
not NOT1 (N9957, N9953);
not NOT1 (N9958, N9951);
buf BUF1 (N9959, N9952);
nor NOR2 (N9960, N9942, N7571);
and AND2 (N9961, N9939, N202);
and AND4 (N9962, N9954, N2685, N21, N29);
xor XOR2 (N9963, N9948, N8538);
and AND3 (N9964, N9955, N689, N5580);
not NOT1 (N9965, N9964);
or OR4 (N9966, N9956, N6314, N4080, N8343);
or OR3 (N9967, N9965, N6001, N4695);
nand NAND2 (N9968, N9958, N6675);
nor NOR4 (N9969, N9968, N2178, N8807, N2771);
not NOT1 (N9970, N9957);
xor XOR2 (N9971, N9960, N5774);
or OR4 (N9972, N9970, N5752, N8773, N134);
nand NAND4 (N9973, N9949, N8757, N3322, N3295);
and AND3 (N9974, N9959, N2560, N9656);
and AND2 (N9975, N9971, N6254);
not NOT1 (N9976, N9963);
buf BUF1 (N9977, N9969);
buf BUF1 (N9978, N9977);
nor NOR2 (N9979, N9973, N2456);
and AND2 (N9980, N9972, N6151);
or OR3 (N9981, N9974, N6353, N6740);
or OR4 (N9982, N9981, N8173, N5179, N3672);
or OR4 (N9983, N9976, N5921, N8409, N316);
nor NOR4 (N9984, N9979, N4228, N3294, N8997);
buf BUF1 (N9985, N9966);
nand NAND3 (N9986, N9961, N1819, N4375);
nand NAND4 (N9987, N9983, N3936, N531, N6893);
xor XOR2 (N9988, N9967, N1902);
nor NOR2 (N9989, N9975, N1414);
xor XOR2 (N9990, N9984, N4528);
xor XOR2 (N9991, N9978, N6638);
not NOT1 (N9992, N9990);
not NOT1 (N9993, N9989);
nand NAND3 (N9994, N9991, N794, N9590);
xor XOR2 (N9995, N9962, N7544);
nor NOR2 (N9996, N9994, N7950);
nor NOR2 (N9997, N9980, N8376);
nor NOR2 (N9998, N9992, N7988);
or OR4 (N9999, N9988, N630, N4995, N7565);
nand NAND4 (N10000, N9996, N5259, N3927, N3760);
or OR3 (N10001, N9999, N6499, N6678);
xor XOR2 (N10002, N9995, N4257);
or OR4 (N10003, N9998, N4570, N7717, N101);
nor NOR2 (N10004, N9993, N4155);
not NOT1 (N10005, N10000);
buf BUF1 (N10006, N10002);
xor XOR2 (N10007, N9986, N5018);
or OR4 (N10008, N9987, N1927, N3340, N8256);
nor NOR2 (N10009, N9982, N2623);
nor NOR3 (N10010, N10007, N6808, N9351);
nand NAND3 (N10011, N9997, N9669, N4297);
not NOT1 (N10012, N10009);
not NOT1 (N10013, N10004);
xor XOR2 (N10014, N10005, N2241);
buf BUF1 (N10015, N10013);
and AND3 (N10016, N10014, N9763, N64);
not NOT1 (N10017, N10003);
and AND3 (N10018, N10011, N2408, N7069);
and AND3 (N10019, N10016, N1023, N9905);
nand NAND2 (N10020, N10006, N1835);
nand NAND3 (N10021, N10001, N7707, N1232);
not NOT1 (N10022, N10021);
or OR4 (N10023, N10010, N2585, N818, N3640);
not NOT1 (N10024, N10018);
nand NAND2 (N10025, N10020, N398);
or OR2 (N10026, N10023, N5731);
xor XOR2 (N10027, N10015, N4467);
not NOT1 (N10028, N10008);
not NOT1 (N10029, N10019);
buf BUF1 (N10030, N10029);
nor NOR2 (N10031, N10026, N1245);
and AND4 (N10032, N9985, N9860, N164, N3731);
or OR3 (N10033, N10028, N2912, N213);
buf BUF1 (N10034, N10012);
nor NOR2 (N10035, N10025, N7842);
not NOT1 (N10036, N10033);
or OR3 (N10037, N10017, N9653, N6413);
buf BUF1 (N10038, N10037);
buf BUF1 (N10039, N10035);
not NOT1 (N10040, N10034);
nor NOR3 (N10041, N10032, N9384, N6003);
xor XOR2 (N10042, N10024, N901);
not NOT1 (N10043, N10027);
nor NOR3 (N10044, N10031, N588, N2965);
buf BUF1 (N10045, N10022);
nor NOR4 (N10046, N10042, N4456, N8952, N4016);
xor XOR2 (N10047, N10030, N346);
and AND3 (N10048, N10039, N4265, N1936);
and AND4 (N10049, N10044, N1771, N6698, N4187);
or OR3 (N10050, N10043, N1426, N8686);
and AND4 (N10051, N10040, N701, N9709, N1360);
and AND3 (N10052, N10036, N4624, N5244);
xor XOR2 (N10053, N10038, N6055);
nor NOR2 (N10054, N10046, N5581);
and AND2 (N10055, N10047, N3768);
xor XOR2 (N10056, N10053, N269);
or OR4 (N10057, N10055, N9975, N5889, N10029);
nand NAND2 (N10058, N10052, N7373);
not NOT1 (N10059, N10049);
not NOT1 (N10060, N10045);
xor XOR2 (N10061, N10048, N2174);
and AND2 (N10062, N10051, N7603);
and AND2 (N10063, N10059, N9144);
or OR4 (N10064, N10058, N7617, N2276, N2431);
not NOT1 (N10065, N10054);
nor NOR3 (N10066, N10060, N9428, N287);
nand NAND2 (N10067, N10062, N121);
and AND3 (N10068, N10066, N142, N2286);
and AND3 (N10069, N10057, N5180, N5313);
not NOT1 (N10070, N10056);
xor XOR2 (N10071, N10067, N7665);
nor NOR2 (N10072, N10070, N8069);
not NOT1 (N10073, N10061);
buf BUF1 (N10074, N10073);
nor NOR3 (N10075, N10074, N7890, N7889);
or OR3 (N10076, N10071, N221, N6017);
buf BUF1 (N10077, N10072);
xor XOR2 (N10078, N10041, N1129);
or OR2 (N10079, N10063, N7900);
and AND3 (N10080, N10069, N6900, N4259);
and AND2 (N10081, N10077, N6289);
nor NOR2 (N10082, N10080, N3566);
nand NAND4 (N10083, N10050, N9664, N4030, N7088);
and AND4 (N10084, N10083, N7009, N645, N1669);
or OR4 (N10085, N10084, N2095, N3095, N6631);
nand NAND2 (N10086, N10078, N7864);
buf BUF1 (N10087, N10065);
or OR3 (N10088, N10079, N8045, N6044);
not NOT1 (N10089, N10064);
or OR4 (N10090, N10082, N5719, N5844, N7146);
or OR2 (N10091, N10076, N3551);
and AND3 (N10092, N10087, N3602, N9051);
not NOT1 (N10093, N10092);
nor NOR3 (N10094, N10075, N9414, N9923);
or OR3 (N10095, N10086, N4442, N4492);
nor NOR3 (N10096, N10094, N1405, N9218);
nor NOR4 (N10097, N10089, N10087, N8196, N6115);
and AND4 (N10098, N10091, N5368, N6806, N9675);
buf BUF1 (N10099, N10096);
not NOT1 (N10100, N10068);
nor NOR2 (N10101, N10093, N8721);
nand NAND4 (N10102, N10098, N7057, N8298, N3448);
nand NAND3 (N10103, N10088, N7631, N7138);
not NOT1 (N10104, N10095);
nor NOR2 (N10105, N10099, N8047);
xor XOR2 (N10106, N10103, N4558);
nor NOR3 (N10107, N10081, N3578, N178);
and AND2 (N10108, N10085, N3234);
xor XOR2 (N10109, N10105, N212);
nand NAND2 (N10110, N10101, N3038);
nor NOR3 (N10111, N10100, N3707, N5774);
and AND3 (N10112, N10106, N7530, N4807);
nor NOR2 (N10113, N10110, N4982);
nand NAND3 (N10114, N10109, N7091, N4085);
nand NAND3 (N10115, N10113, N2408, N3779);
nand NAND2 (N10116, N10112, N696);
and AND4 (N10117, N10107, N8513, N5915, N1480);
and AND4 (N10118, N10116, N2110, N8507, N4909);
nor NOR4 (N10119, N10115, N2821, N3430, N812);
xor XOR2 (N10120, N10111, N5562);
xor XOR2 (N10121, N10097, N3790);
not NOT1 (N10122, N10090);
buf BUF1 (N10123, N10122);
xor XOR2 (N10124, N10108, N7366);
buf BUF1 (N10125, N10119);
and AND3 (N10126, N10120, N2982, N337);
xor XOR2 (N10127, N10114, N2425);
not NOT1 (N10128, N10104);
and AND2 (N10129, N10123, N475);
xor XOR2 (N10130, N10117, N1917);
xor XOR2 (N10131, N10124, N9972);
not NOT1 (N10132, N10126);
nor NOR4 (N10133, N10128, N3448, N5058, N3390);
or OR4 (N10134, N10125, N5691, N5229, N9096);
xor XOR2 (N10135, N10131, N9264);
nor NOR4 (N10136, N10118, N5699, N1721, N1611);
nor NOR4 (N10137, N10134, N9489, N9451, N7173);
and AND4 (N10138, N10130, N9028, N3572, N7858);
buf BUF1 (N10139, N10136);
buf BUF1 (N10140, N10135);
nor NOR3 (N10141, N10139, N1491, N1542);
nand NAND4 (N10142, N10137, N6422, N2490, N3921);
xor XOR2 (N10143, N10138, N8935);
xor XOR2 (N10144, N10132, N590);
or OR2 (N10145, N10144, N4152);
and AND3 (N10146, N10102, N6124, N1139);
not NOT1 (N10147, N10127);
xor XOR2 (N10148, N10143, N2590);
nor NOR2 (N10149, N10148, N5671);
nor NOR4 (N10150, N10133, N7563, N7373, N5571);
and AND4 (N10151, N10142, N9026, N6532, N8210);
not NOT1 (N10152, N10129);
xor XOR2 (N10153, N10152, N3736);
buf BUF1 (N10154, N10146);
xor XOR2 (N10155, N10150, N8625);
or OR3 (N10156, N10153, N8196, N5964);
nand NAND3 (N10157, N10156, N8190, N6185);
xor XOR2 (N10158, N10145, N8900);
nor NOR2 (N10159, N10140, N1945);
nor NOR3 (N10160, N10158, N3737, N2431);
nor NOR3 (N10161, N10141, N1107, N8950);
buf BUF1 (N10162, N10157);
nor NOR4 (N10163, N10160, N5484, N6884, N5716);
nand NAND4 (N10164, N10155, N3950, N4309, N7990);
nand NAND3 (N10165, N10163, N6573, N1626);
or OR3 (N10166, N10159, N9250, N2851);
or OR3 (N10167, N10154, N517, N53);
xor XOR2 (N10168, N10165, N5055);
and AND4 (N10169, N10161, N4590, N767, N5271);
nor NOR3 (N10170, N10121, N2189, N6982);
buf BUF1 (N10171, N10149);
or OR4 (N10172, N10169, N847, N460, N3641);
buf BUF1 (N10173, N10172);
not NOT1 (N10174, N10166);
nor NOR4 (N10175, N10174, N8969, N6852, N8760);
or OR2 (N10176, N10171, N5943);
buf BUF1 (N10177, N10162);
buf BUF1 (N10178, N10173);
buf BUF1 (N10179, N10175);
not NOT1 (N10180, N10179);
nor NOR3 (N10181, N10147, N5097, N8493);
or OR4 (N10182, N10170, N262, N4609, N8005);
nor NOR2 (N10183, N10177, N6121);
buf BUF1 (N10184, N10176);
or OR4 (N10185, N10178, N5284, N1355, N2821);
xor XOR2 (N10186, N10180, N3196);
not NOT1 (N10187, N10182);
or OR2 (N10188, N10184, N9678);
or OR2 (N10189, N10168, N9994);
nand NAND4 (N10190, N10185, N2850, N3869, N5446);
not NOT1 (N10191, N10164);
xor XOR2 (N10192, N10187, N2058);
not NOT1 (N10193, N10181);
buf BUF1 (N10194, N10151);
buf BUF1 (N10195, N10194);
or OR3 (N10196, N10167, N9140, N7787);
not NOT1 (N10197, N10183);
not NOT1 (N10198, N10196);
buf BUF1 (N10199, N10191);
xor XOR2 (N10200, N10197, N9134);
nand NAND4 (N10201, N10195, N6685, N4465, N3756);
xor XOR2 (N10202, N10192, N9321);
nor NOR4 (N10203, N10188, N9462, N2518, N3732);
not NOT1 (N10204, N10193);
xor XOR2 (N10205, N10204, N1773);
and AND4 (N10206, N10200, N3315, N244, N4574);
nor NOR2 (N10207, N10190, N2923);
and AND4 (N10208, N10202, N1659, N9955, N6601);
and AND2 (N10209, N10201, N1020);
buf BUF1 (N10210, N10208);
and AND4 (N10211, N10210, N2260, N5029, N4255);
and AND2 (N10212, N10189, N5248);
buf BUF1 (N10213, N10211);
xor XOR2 (N10214, N10206, N8411);
xor XOR2 (N10215, N10199, N5842);
and AND2 (N10216, N10205, N1956);
nor NOR4 (N10217, N10207, N8212, N1369, N2691);
nor NOR2 (N10218, N10216, N2593);
nand NAND2 (N10219, N10212, N724);
or OR3 (N10220, N10215, N5390, N6771);
nand NAND3 (N10221, N10217, N6045, N3286);
nand NAND4 (N10222, N10186, N6334, N7449, N646);
and AND2 (N10223, N10198, N1736);
nor NOR4 (N10224, N10223, N7985, N2287, N4744);
nor NOR2 (N10225, N10203, N4587);
nand NAND3 (N10226, N10209, N3099, N7101);
nor NOR2 (N10227, N10219, N9370);
nor NOR2 (N10228, N10226, N9492);
nand NAND3 (N10229, N10214, N8185, N6081);
not NOT1 (N10230, N10213);
or OR2 (N10231, N10218, N2258);
buf BUF1 (N10232, N10221);
nand NAND3 (N10233, N10230, N4817, N5363);
nand NAND4 (N10234, N10220, N925, N622, N3867);
or OR3 (N10235, N10232, N8724, N9098);
and AND2 (N10236, N10234, N6558);
nand NAND2 (N10237, N10224, N4482);
xor XOR2 (N10238, N10231, N5008);
nand NAND4 (N10239, N10233, N153, N196, N1592);
not NOT1 (N10240, N10222);
not NOT1 (N10241, N10236);
buf BUF1 (N10242, N10235);
and AND3 (N10243, N10229, N8402, N7656);
nand NAND3 (N10244, N10227, N7374, N4635);
nand NAND3 (N10245, N10240, N1769, N1455);
buf BUF1 (N10246, N10228);
nand NAND2 (N10247, N10237, N7397);
nand NAND3 (N10248, N10247, N5591, N5170);
nand NAND2 (N10249, N10244, N6091);
and AND4 (N10250, N10248, N4844, N5865, N7051);
buf BUF1 (N10251, N10246);
or OR4 (N10252, N10243, N3969, N5385, N842);
or OR4 (N10253, N10249, N232, N2354, N9744);
and AND4 (N10254, N10245, N9604, N8144, N1955);
nor NOR3 (N10255, N10241, N1051, N5123);
xor XOR2 (N10256, N10253, N9704);
or OR3 (N10257, N10242, N3083, N8997);
and AND3 (N10258, N10255, N8430, N2601);
xor XOR2 (N10259, N10251, N3178);
xor XOR2 (N10260, N10254, N3421);
xor XOR2 (N10261, N10238, N5587);
nor NOR3 (N10262, N10257, N9176, N6276);
nor NOR3 (N10263, N10252, N3462, N3232);
buf BUF1 (N10264, N10263);
and AND2 (N10265, N10259, N5294);
nor NOR3 (N10266, N10258, N6029, N2864);
or OR2 (N10267, N10262, N6695);
nand NAND2 (N10268, N10256, N9644);
nor NOR2 (N10269, N10260, N398);
nor NOR3 (N10270, N10261, N1209, N5647);
nor NOR4 (N10271, N10266, N3845, N3731, N2377);
buf BUF1 (N10272, N10270);
nand NAND4 (N10273, N10272, N7089, N7173, N695);
and AND3 (N10274, N10239, N5857, N7083);
not NOT1 (N10275, N10273);
buf BUF1 (N10276, N10264);
and AND2 (N10277, N10268, N5060);
nand NAND4 (N10278, N10225, N9478, N8267, N4381);
or OR3 (N10279, N10250, N3315, N249);
buf BUF1 (N10280, N10269);
and AND3 (N10281, N10274, N375, N1751);
buf BUF1 (N10282, N10280);
and AND2 (N10283, N10265, N7671);
xor XOR2 (N10284, N10279, N3266);
or OR3 (N10285, N10284, N2657, N2856);
xor XOR2 (N10286, N10267, N8716);
nand NAND2 (N10287, N10282, N5336);
or OR2 (N10288, N10285, N9535);
buf BUF1 (N10289, N10286);
or OR4 (N10290, N10283, N4241, N1815, N5187);
xor XOR2 (N10291, N10271, N527);
nand NAND4 (N10292, N10288, N3157, N6068, N2964);
and AND2 (N10293, N10281, N1056);
xor XOR2 (N10294, N10277, N7959);
or OR3 (N10295, N10287, N1709, N8812);
nor NOR4 (N10296, N10278, N2859, N7592, N4482);
xor XOR2 (N10297, N10291, N3075);
nor NOR3 (N10298, N10297, N8192, N2382);
and AND4 (N10299, N10292, N9664, N6377, N2145);
xor XOR2 (N10300, N10290, N9389);
nand NAND3 (N10301, N10299, N9250, N3904);
xor XOR2 (N10302, N10296, N7607);
buf BUF1 (N10303, N10275);
and AND2 (N10304, N10301, N4782);
nor NOR3 (N10305, N10302, N8367, N2604);
buf BUF1 (N10306, N10293);
not NOT1 (N10307, N10295);
nand NAND2 (N10308, N10303, N7349);
xor XOR2 (N10309, N10308, N6649);
or OR4 (N10310, N10276, N7339, N5893, N2611);
buf BUF1 (N10311, N10289);
or OR4 (N10312, N10294, N5170, N35, N10261);
nor NOR3 (N10313, N10307, N2456, N2634);
nand NAND4 (N10314, N10309, N7878, N7731, N9856);
nand NAND3 (N10315, N10314, N10283, N1019);
or OR2 (N10316, N10306, N3206);
nor NOR4 (N10317, N10304, N5516, N7417, N5622);
buf BUF1 (N10318, N10315);
or OR4 (N10319, N10310, N1180, N6207, N8422);
and AND3 (N10320, N10317, N2131, N6059);
nand NAND2 (N10321, N10300, N9141);
and AND2 (N10322, N10319, N3351);
buf BUF1 (N10323, N10298);
or OR2 (N10324, N10320, N7138);
buf BUF1 (N10325, N10322);
or OR4 (N10326, N10313, N7511, N4768, N4630);
or OR4 (N10327, N10324, N6983, N5544, N6970);
xor XOR2 (N10328, N10327, N5259);
nand NAND3 (N10329, N10321, N9929, N7617);
nor NOR4 (N10330, N10329, N9570, N1732, N3878);
nor NOR2 (N10331, N10311, N2182);
buf BUF1 (N10332, N10323);
and AND4 (N10333, N10332, N6975, N4372, N9546);
nor NOR3 (N10334, N10305, N7945, N8429);
and AND4 (N10335, N10328, N5878, N2500, N9660);
nor NOR3 (N10336, N10330, N10184, N5295);
or OR3 (N10337, N10336, N7668, N9282);
or OR4 (N10338, N10326, N3568, N4463, N5984);
nand NAND3 (N10339, N10331, N7435, N9889);
and AND4 (N10340, N10337, N5547, N5487, N7453);
xor XOR2 (N10341, N10333, N8131);
buf BUF1 (N10342, N10316);
buf BUF1 (N10343, N10342);
or OR3 (N10344, N10325, N9730, N3358);
or OR4 (N10345, N10338, N4410, N3281, N4604);
buf BUF1 (N10346, N10340);
nand NAND4 (N10347, N10318, N7712, N34, N2550);
xor XOR2 (N10348, N10339, N9483);
and AND3 (N10349, N10345, N131, N4670);
or OR4 (N10350, N10343, N8711, N3558, N2365);
nand NAND4 (N10351, N10347, N162, N3515, N5361);
not NOT1 (N10352, N10348);
or OR3 (N10353, N10341, N9128, N9669);
nor NOR2 (N10354, N10335, N2108);
not NOT1 (N10355, N10312);
and AND3 (N10356, N10334, N3920, N6614);
nor NOR4 (N10357, N10353, N7567, N8719, N1030);
xor XOR2 (N10358, N10354, N8061);
and AND3 (N10359, N10349, N7400, N6410);
nor NOR3 (N10360, N10358, N5977, N4578);
not NOT1 (N10361, N10350);
nand NAND2 (N10362, N10357, N222);
not NOT1 (N10363, N10362);
nor NOR3 (N10364, N10361, N4288, N1126);
not NOT1 (N10365, N10355);
buf BUF1 (N10366, N10351);
not NOT1 (N10367, N10356);
and AND2 (N10368, N10364, N1725);
buf BUF1 (N10369, N10365);
buf BUF1 (N10370, N10363);
or OR2 (N10371, N10369, N412);
or OR2 (N10372, N10371, N8625);
and AND3 (N10373, N10344, N3659, N6479);
xor XOR2 (N10374, N10366, N6397);
buf BUF1 (N10375, N10374);
and AND2 (N10376, N10368, N6358);
nand NAND3 (N10377, N10373, N5510, N7006);
xor XOR2 (N10378, N10359, N4463);
xor XOR2 (N10379, N10376, N9965);
not NOT1 (N10380, N10372);
nor NOR3 (N10381, N10375, N8672, N9684);
or OR2 (N10382, N10346, N5040);
and AND3 (N10383, N10370, N6756, N1454);
nor NOR3 (N10384, N10367, N1861, N1876);
xor XOR2 (N10385, N10381, N4533);
buf BUF1 (N10386, N10377);
xor XOR2 (N10387, N10378, N9225);
or OR4 (N10388, N10382, N3381, N3638, N7989);
nand NAND4 (N10389, N10385, N6683, N1821, N7391);
nor NOR2 (N10390, N10360, N10054);
buf BUF1 (N10391, N10386);
xor XOR2 (N10392, N10379, N2717);
buf BUF1 (N10393, N10392);
or OR2 (N10394, N10384, N1285);
nor NOR2 (N10395, N10352, N5879);
nor NOR2 (N10396, N10389, N399);
buf BUF1 (N10397, N10393);
nand NAND2 (N10398, N10395, N382);
nor NOR3 (N10399, N10398, N2680, N5315);
or OR3 (N10400, N10383, N3471, N8363);
nand NAND4 (N10401, N10380, N253, N157, N1685);
nand NAND4 (N10402, N10397, N8466, N8466, N7030);
buf BUF1 (N10403, N10399);
buf BUF1 (N10404, N10400);
xor XOR2 (N10405, N10391, N6054);
nand NAND3 (N10406, N10388, N1077, N8756);
or OR4 (N10407, N10403, N772, N1618, N5533);
or OR2 (N10408, N10387, N9993);
xor XOR2 (N10409, N10404, N6785);
xor XOR2 (N10410, N10401, N8678);
buf BUF1 (N10411, N10396);
buf BUF1 (N10412, N10405);
nor NOR4 (N10413, N10408, N8869, N6479, N5849);
nand NAND3 (N10414, N10409, N30, N781);
or OR4 (N10415, N10390, N6268, N7869, N9682);
or OR4 (N10416, N10411, N1590, N9280, N23);
nor NOR3 (N10417, N10414, N2626, N8203);
not NOT1 (N10418, N10407);
or OR4 (N10419, N10415, N8141, N3978, N4857);
and AND3 (N10420, N10417, N7788, N4359);
not NOT1 (N10421, N10418);
buf BUF1 (N10422, N10402);
or OR3 (N10423, N10419, N7074, N2757);
xor XOR2 (N10424, N10412, N2692);
not NOT1 (N10425, N10413);
nor NOR3 (N10426, N10416, N7832, N7185);
xor XOR2 (N10427, N10423, N1645);
not NOT1 (N10428, N10421);
xor XOR2 (N10429, N10394, N710);
nor NOR3 (N10430, N10422, N2898, N6148);
nand NAND2 (N10431, N10424, N9884);
nor NOR4 (N10432, N10427, N8990, N3445, N2735);
buf BUF1 (N10433, N10410);
not NOT1 (N10434, N10433);
nand NAND3 (N10435, N10430, N3886, N6009);
xor XOR2 (N10436, N10431, N10058);
buf BUF1 (N10437, N10425);
or OR2 (N10438, N10428, N377);
xor XOR2 (N10439, N10438, N3320);
not NOT1 (N10440, N10406);
or OR3 (N10441, N10435, N852, N3859);
not NOT1 (N10442, N10420);
not NOT1 (N10443, N10436);
xor XOR2 (N10444, N10434, N5294);
xor XOR2 (N10445, N10432, N10400);
buf BUF1 (N10446, N10426);
or OR3 (N10447, N10441, N4985, N5241);
nor NOR2 (N10448, N10439, N6228);
xor XOR2 (N10449, N10446, N7539);
not NOT1 (N10450, N10445);
and AND4 (N10451, N10450, N3735, N5080, N4660);
or OR4 (N10452, N10447, N1186, N4993, N4799);
nand NAND4 (N10453, N10437, N10132, N8264, N4202);
or OR4 (N10454, N10440, N8646, N8919, N9856);
nor NOR2 (N10455, N10454, N2714);
xor XOR2 (N10456, N10444, N6979);
nor NOR4 (N10457, N10452, N9470, N5586, N6598);
buf BUF1 (N10458, N10455);
and AND2 (N10459, N10453, N1649);
not NOT1 (N10460, N10458);
or OR3 (N10461, N10443, N427, N1032);
and AND2 (N10462, N10442, N6765);
nand NAND3 (N10463, N10429, N4344, N9570);
not NOT1 (N10464, N10460);
not NOT1 (N10465, N10457);
or OR2 (N10466, N10448, N558);
buf BUF1 (N10467, N10456);
buf BUF1 (N10468, N10451);
not NOT1 (N10469, N10466);
xor XOR2 (N10470, N10461, N3465);
nor NOR4 (N10471, N10462, N1427, N3159, N1460);
xor XOR2 (N10472, N10468, N9551);
nor NOR3 (N10473, N10469, N6074, N6455);
or OR3 (N10474, N10465, N10174, N9030);
and AND3 (N10475, N10470, N5695, N8717);
or OR4 (N10476, N10467, N828, N1308, N5381);
or OR2 (N10477, N10473, N1008);
buf BUF1 (N10478, N10471);
not NOT1 (N10479, N10459);
not NOT1 (N10480, N10476);
xor XOR2 (N10481, N10478, N7127);
nor NOR4 (N10482, N10475, N3375, N4666, N1904);
and AND3 (N10483, N10479, N10317, N2136);
nand NAND4 (N10484, N10481, N938, N4670, N3656);
or OR4 (N10485, N10474, N661, N5386, N4601);
or OR4 (N10486, N10482, N9844, N7926, N1144);
or OR3 (N10487, N10464, N8634, N2333);
or OR4 (N10488, N10472, N4840, N10246, N5288);
nor NOR2 (N10489, N10488, N6990);
nor NOR4 (N10490, N10484, N4501, N9688, N4267);
not NOT1 (N10491, N10449);
nor NOR3 (N10492, N10463, N9069, N9226);
buf BUF1 (N10493, N10487);
xor XOR2 (N10494, N10493, N1785);
xor XOR2 (N10495, N10494, N5635);
xor XOR2 (N10496, N10477, N3920);
buf BUF1 (N10497, N10496);
or OR2 (N10498, N10491, N4350);
not NOT1 (N10499, N10492);
nor NOR2 (N10500, N10497, N3773);
nand NAND3 (N10501, N10489, N3745, N1828);
xor XOR2 (N10502, N10483, N2199);
xor XOR2 (N10503, N10495, N3350);
not NOT1 (N10504, N10499);
xor XOR2 (N10505, N10486, N9918);
and AND2 (N10506, N10485, N6020);
or OR4 (N10507, N10506, N3397, N205, N2348);
or OR4 (N10508, N10501, N4790, N2383, N1422);
nor NOR3 (N10509, N10480, N4925, N7523);
and AND4 (N10510, N10505, N1577, N6671, N3890);
not NOT1 (N10511, N10490);
not NOT1 (N10512, N10508);
xor XOR2 (N10513, N10511, N6253);
not NOT1 (N10514, N10500);
or OR4 (N10515, N10514, N8592, N2904, N1688);
xor XOR2 (N10516, N10502, N2514);
and AND4 (N10517, N10510, N2626, N219, N9562);
buf BUF1 (N10518, N10515);
or OR4 (N10519, N10518, N539, N6273, N7198);
xor XOR2 (N10520, N10519, N7527);
and AND4 (N10521, N10516, N4923, N6121, N7585);
and AND2 (N10522, N10498, N9871);
and AND4 (N10523, N10512, N6051, N4312, N6363);
or OR4 (N10524, N10503, N7010, N4388, N5902);
nor NOR3 (N10525, N10504, N5666, N6036);
buf BUF1 (N10526, N10517);
or OR2 (N10527, N10526, N10247);
nand NAND2 (N10528, N10521, N6967);
xor XOR2 (N10529, N10523, N2438);
not NOT1 (N10530, N10527);
nand NAND3 (N10531, N10528, N6177, N1786);
buf BUF1 (N10532, N10520);
buf BUF1 (N10533, N10532);
xor XOR2 (N10534, N10529, N4107);
or OR4 (N10535, N10525, N3301, N803, N2366);
nand NAND4 (N10536, N10513, N5896, N9947, N9247);
buf BUF1 (N10537, N10531);
xor XOR2 (N10538, N10507, N6493);
nand NAND2 (N10539, N10538, N2046);
and AND4 (N10540, N10536, N246, N1141, N4881);
nor NOR3 (N10541, N10540, N6969, N5940);
and AND2 (N10542, N10533, N3337);
xor XOR2 (N10543, N10539, N7465);
buf BUF1 (N10544, N10541);
nand NAND4 (N10545, N10543, N8020, N9465, N8699);
nand NAND4 (N10546, N10535, N6938, N1018, N4764);
xor XOR2 (N10547, N10524, N9348);
xor XOR2 (N10548, N10509, N6301);
buf BUF1 (N10549, N10542);
buf BUF1 (N10550, N10537);
not NOT1 (N10551, N10534);
not NOT1 (N10552, N10545);
xor XOR2 (N10553, N10550, N2506);
nand NAND3 (N10554, N10549, N8056, N5566);
not NOT1 (N10555, N10530);
buf BUF1 (N10556, N10553);
xor XOR2 (N10557, N10552, N2919);
not NOT1 (N10558, N10548);
buf BUF1 (N10559, N10558);
not NOT1 (N10560, N10551);
not NOT1 (N10561, N10556);
nor NOR4 (N10562, N10554, N6199, N3785, N8183);
or OR3 (N10563, N10544, N3118, N9233);
not NOT1 (N10564, N10562);
xor XOR2 (N10565, N10522, N4837);
not NOT1 (N10566, N10546);
nand NAND3 (N10567, N10547, N8578, N6746);
not NOT1 (N10568, N10567);
buf BUF1 (N10569, N10564);
nor NOR4 (N10570, N10557, N10481, N1593, N1002);
nand NAND4 (N10571, N10570, N6950, N3011, N3102);
and AND3 (N10572, N10565, N10537, N9352);
not NOT1 (N10573, N10561);
xor XOR2 (N10574, N10568, N9470);
or OR2 (N10575, N10571, N6485);
not NOT1 (N10576, N10569);
nor NOR2 (N10577, N10563, N5675);
buf BUF1 (N10578, N10577);
xor XOR2 (N10579, N10559, N1326);
not NOT1 (N10580, N10560);
not NOT1 (N10581, N10580);
xor XOR2 (N10582, N10573, N7566);
nor NOR2 (N10583, N10581, N8790);
or OR4 (N10584, N10582, N8564, N10073, N9819);
xor XOR2 (N10585, N10578, N6826);
xor XOR2 (N10586, N10574, N10567);
or OR2 (N10587, N10586, N6483);
nor NOR4 (N10588, N10566, N6971, N8745, N4560);
or OR4 (N10589, N10585, N9057, N5588, N3086);
nand NAND3 (N10590, N10575, N9241, N8712);
xor XOR2 (N10591, N10589, N2290);
buf BUF1 (N10592, N10591);
or OR3 (N10593, N10572, N6174, N9329);
nand NAND4 (N10594, N10590, N10389, N3332, N9013);
nand NAND4 (N10595, N10579, N4325, N4594, N3445);
or OR4 (N10596, N10576, N1399, N4678, N6613);
and AND3 (N10597, N10592, N3301, N5173);
buf BUF1 (N10598, N10583);
buf BUF1 (N10599, N10593);
not NOT1 (N10600, N10596);
not NOT1 (N10601, N10588);
buf BUF1 (N10602, N10584);
xor XOR2 (N10603, N10594, N5139);
nand NAND2 (N10604, N10595, N4399);
and AND2 (N10605, N10604, N8568);
not NOT1 (N10606, N10605);
nand NAND3 (N10607, N10597, N6411, N9475);
nor NOR4 (N10608, N10607, N8199, N5715, N9136);
nor NOR4 (N10609, N10599, N4293, N9493, N421);
buf BUF1 (N10610, N10601);
xor XOR2 (N10611, N10610, N6551);
or OR3 (N10612, N10603, N3997, N5222);
not NOT1 (N10613, N10612);
or OR3 (N10614, N10611, N5539, N2993);
not NOT1 (N10615, N10614);
nand NAND4 (N10616, N10555, N4355, N9981, N2820);
buf BUF1 (N10617, N10613);
not NOT1 (N10618, N10587);
not NOT1 (N10619, N10609);
nor NOR3 (N10620, N10606, N266, N8411);
or OR4 (N10621, N10615, N3691, N4255, N4378);
nand NAND2 (N10622, N10621, N4946);
or OR3 (N10623, N10598, N3393, N3773);
buf BUF1 (N10624, N10600);
or OR3 (N10625, N10616, N8603, N8555);
or OR3 (N10626, N10623, N10024, N6504);
not NOT1 (N10627, N10624);
and AND3 (N10628, N10619, N983, N9418);
nor NOR3 (N10629, N10628, N6534, N8638);
xor XOR2 (N10630, N10620, N7410);
xor XOR2 (N10631, N10617, N2857);
nor NOR3 (N10632, N10622, N3658, N10041);
xor XOR2 (N10633, N10629, N2922);
nor NOR3 (N10634, N10626, N8399, N10129);
buf BUF1 (N10635, N10618);
not NOT1 (N10636, N10634);
or OR2 (N10637, N10632, N7668);
nand NAND4 (N10638, N10608, N4248, N3614, N5869);
nor NOR2 (N10639, N10602, N8527);
xor XOR2 (N10640, N10636, N3510);
not NOT1 (N10641, N10630);
nor NOR2 (N10642, N10639, N10023);
and AND3 (N10643, N10633, N6184, N5632);
xor XOR2 (N10644, N10627, N4741);
and AND4 (N10645, N10644, N5545, N6598, N6197);
buf BUF1 (N10646, N10637);
or OR4 (N10647, N10641, N7008, N2759, N6237);
not NOT1 (N10648, N10635);
and AND3 (N10649, N10648, N8283, N4812);
nor NOR3 (N10650, N10649, N5643, N10273);
or OR2 (N10651, N10645, N8444);
xor XOR2 (N10652, N10638, N1058);
xor XOR2 (N10653, N10651, N7328);
xor XOR2 (N10654, N10647, N7176);
nand NAND2 (N10655, N10652, N749);
or OR3 (N10656, N10625, N3685, N3110);
xor XOR2 (N10657, N10643, N6548);
nand NAND3 (N10658, N10631, N1922, N3279);
and AND2 (N10659, N10655, N3242);
nand NAND4 (N10660, N10659, N6295, N9527, N9141);
nor NOR2 (N10661, N10654, N6833);
and AND3 (N10662, N10657, N3046, N7168);
not NOT1 (N10663, N10662);
nor NOR4 (N10664, N10656, N5094, N2588, N8692);
buf BUF1 (N10665, N10650);
nand NAND2 (N10666, N10664, N468);
or OR3 (N10667, N10642, N3690, N5744);
or OR4 (N10668, N10646, N3238, N4049, N9059);
and AND3 (N10669, N10666, N3655, N6448);
nor NOR3 (N10670, N10668, N7861, N6056);
buf BUF1 (N10671, N10669);
or OR3 (N10672, N10640, N10293, N4792);
or OR4 (N10673, N10658, N527, N8065, N3348);
nor NOR2 (N10674, N10667, N3527);
not NOT1 (N10675, N10665);
or OR4 (N10676, N10671, N68, N7498, N5864);
not NOT1 (N10677, N10675);
xor XOR2 (N10678, N10663, N6204);
buf BUF1 (N10679, N10670);
xor XOR2 (N10680, N10679, N1680);
xor XOR2 (N10681, N10674, N7017);
not NOT1 (N10682, N10677);
or OR2 (N10683, N10676, N7998);
nor NOR3 (N10684, N10661, N6292, N8867);
buf BUF1 (N10685, N10660);
not NOT1 (N10686, N10673);
nand NAND2 (N10687, N10681, N9074);
xor XOR2 (N10688, N10683, N6566);
and AND4 (N10689, N10688, N8931, N5212, N5759);
or OR3 (N10690, N10685, N2150, N6957);
not NOT1 (N10691, N10684);
xor XOR2 (N10692, N10686, N5236);
or OR2 (N10693, N10680, N3391);
and AND2 (N10694, N10690, N1000);
and AND2 (N10695, N10693, N7538);
not NOT1 (N10696, N10692);
nand NAND2 (N10697, N10689, N8914);
nand NAND2 (N10698, N10695, N1262);
buf BUF1 (N10699, N10691);
or OR2 (N10700, N10678, N5018);
nand NAND2 (N10701, N10687, N1850);
buf BUF1 (N10702, N10694);
and AND3 (N10703, N10698, N10656, N7479);
or OR4 (N10704, N10653, N4644, N5774, N8718);
xor XOR2 (N10705, N10704, N1172);
buf BUF1 (N10706, N10682);
xor XOR2 (N10707, N10705, N717);
nor NOR2 (N10708, N10697, N7930);
or OR2 (N10709, N10703, N492);
buf BUF1 (N10710, N10700);
nor NOR3 (N10711, N10708, N7397, N2639);
nor NOR2 (N10712, N10672, N6072);
or OR4 (N10713, N10699, N9943, N2976, N2636);
and AND3 (N10714, N10707, N559, N4110);
and AND2 (N10715, N10702, N2661);
or OR4 (N10716, N10715, N2354, N440, N5889);
buf BUF1 (N10717, N10714);
and AND3 (N10718, N10713, N1351, N8235);
or OR2 (N10719, N10709, N8504);
xor XOR2 (N10720, N10718, N1559);
xor XOR2 (N10721, N10719, N6370);
nand NAND2 (N10722, N10721, N3525);
not NOT1 (N10723, N10712);
nand NAND4 (N10724, N10716, N1269, N954, N4168);
xor XOR2 (N10725, N10701, N8968);
buf BUF1 (N10726, N10706);
xor XOR2 (N10727, N10723, N8587);
nand NAND4 (N10728, N10726, N5529, N9206, N1759);
not NOT1 (N10729, N10696);
and AND4 (N10730, N10725, N6792, N467, N2394);
not NOT1 (N10731, N10727);
and AND2 (N10732, N10710, N9293);
or OR3 (N10733, N10717, N1425, N2975);
xor XOR2 (N10734, N10720, N1784);
nand NAND4 (N10735, N10730, N1498, N8919, N1030);
xor XOR2 (N10736, N10731, N4918);
nand NAND3 (N10737, N10711, N649, N9104);
nand NAND4 (N10738, N10736, N9390, N4801, N6449);
not NOT1 (N10739, N10722);
xor XOR2 (N10740, N10729, N9850);
not NOT1 (N10741, N10738);
nand NAND2 (N10742, N10734, N4619);
buf BUF1 (N10743, N10728);
or OR2 (N10744, N10743, N5579);
not NOT1 (N10745, N10732);
or OR3 (N10746, N10724, N5724, N6339);
xor XOR2 (N10747, N10746, N3622);
nor NOR4 (N10748, N10744, N4214, N668, N341);
or OR4 (N10749, N10739, N6852, N4062, N3513);
or OR3 (N10750, N10747, N3065, N597);
nand NAND3 (N10751, N10749, N3647, N2293);
nand NAND2 (N10752, N10741, N9978);
and AND2 (N10753, N10733, N4075);
or OR3 (N10754, N10748, N10206, N5354);
and AND3 (N10755, N10740, N34, N3508);
nand NAND2 (N10756, N10754, N8751);
nor NOR3 (N10757, N10751, N5279, N3781);
buf BUF1 (N10758, N10742);
not NOT1 (N10759, N10737);
not NOT1 (N10760, N10758);
nor NOR2 (N10761, N10753, N3414);
buf BUF1 (N10762, N10760);
buf BUF1 (N10763, N10745);
not NOT1 (N10764, N10759);
nand NAND3 (N10765, N10752, N2959, N10208);
xor XOR2 (N10766, N10750, N9178);
not NOT1 (N10767, N10757);
or OR4 (N10768, N10735, N5096, N4897, N6819);
and AND3 (N10769, N10755, N9541, N2539);
or OR4 (N10770, N10766, N10195, N4854, N4656);
or OR4 (N10771, N10763, N8112, N10643, N4951);
nor NOR4 (N10772, N10756, N10201, N3176, N2064);
nand NAND3 (N10773, N10767, N3686, N5924);
xor XOR2 (N10774, N10761, N7658);
and AND2 (N10775, N10770, N6216);
and AND3 (N10776, N10775, N203, N8790);
and AND4 (N10777, N10769, N8933, N8369, N7260);
buf BUF1 (N10778, N10768);
nor NOR4 (N10779, N10777, N8872, N4126, N4309);
nand NAND4 (N10780, N10774, N4572, N8971, N2534);
or OR2 (N10781, N10778, N8555);
xor XOR2 (N10782, N10779, N8311);
or OR3 (N10783, N10780, N9913, N5652);
xor XOR2 (N10784, N10771, N5164);
or OR2 (N10785, N10782, N8708);
not NOT1 (N10786, N10784);
and AND4 (N10787, N10776, N5618, N9315, N6585);
buf BUF1 (N10788, N10785);
xor XOR2 (N10789, N10786, N2875);
or OR4 (N10790, N10764, N8239, N889, N411);
buf BUF1 (N10791, N10765);
not NOT1 (N10792, N10787);
and AND2 (N10793, N10791, N3588);
or OR4 (N10794, N10772, N8548, N5697, N1455);
or OR4 (N10795, N10773, N10289, N8217, N1569);
nor NOR3 (N10796, N10783, N3772, N637);
or OR4 (N10797, N10790, N6140, N9781, N2810);
xor XOR2 (N10798, N10789, N3088);
xor XOR2 (N10799, N10793, N4003);
or OR3 (N10800, N10792, N9934, N2054);
or OR3 (N10801, N10799, N8277, N9681);
or OR3 (N10802, N10798, N4224, N2533);
buf BUF1 (N10803, N10797);
buf BUF1 (N10804, N10762);
buf BUF1 (N10805, N10801);
nand NAND4 (N10806, N10796, N8887, N10290, N7844);
not NOT1 (N10807, N10802);
or OR2 (N10808, N10807, N1722);
not NOT1 (N10809, N10806);
not NOT1 (N10810, N10809);
xor XOR2 (N10811, N10810, N9175);
buf BUF1 (N10812, N10804);
or OR2 (N10813, N10795, N9145);
not NOT1 (N10814, N10788);
not NOT1 (N10815, N10781);
buf BUF1 (N10816, N10800);
and AND4 (N10817, N10814, N7794, N4781, N5655);
and AND3 (N10818, N10817, N9765, N6753);
buf BUF1 (N10819, N10794);
buf BUF1 (N10820, N10819);
not NOT1 (N10821, N10813);
not NOT1 (N10822, N10805);
not NOT1 (N10823, N10803);
nand NAND3 (N10824, N10818, N8277, N6362);
buf BUF1 (N10825, N10820);
xor XOR2 (N10826, N10815, N8677);
and AND3 (N10827, N10823, N4345, N9765);
and AND2 (N10828, N10826, N4402);
or OR2 (N10829, N10808, N3910);
and AND3 (N10830, N10828, N9116, N899);
buf BUF1 (N10831, N10822);
or OR2 (N10832, N10829, N2459);
nand NAND4 (N10833, N10811, N4349, N3678, N3898);
and AND3 (N10834, N10832, N3592, N8716);
not NOT1 (N10835, N10812);
buf BUF1 (N10836, N10824);
xor XOR2 (N10837, N10821, N2047);
or OR4 (N10838, N10825, N6615, N2932, N7861);
buf BUF1 (N10839, N10834);
or OR2 (N10840, N10835, N4782);
nand NAND2 (N10841, N10840, N8864);
or OR2 (N10842, N10837, N3325);
not NOT1 (N10843, N10838);
or OR2 (N10844, N10842, N8973);
not NOT1 (N10845, N10839);
not NOT1 (N10846, N10827);
nor NOR3 (N10847, N10833, N4327, N10366);
xor XOR2 (N10848, N10831, N9019);
nand NAND4 (N10849, N10843, N8600, N2500, N5708);
xor XOR2 (N10850, N10836, N7417);
xor XOR2 (N10851, N10849, N5074);
and AND2 (N10852, N10841, N1817);
buf BUF1 (N10853, N10830);
nand NAND3 (N10854, N10846, N10056, N5010);
xor XOR2 (N10855, N10850, N1166);
not NOT1 (N10856, N10816);
xor XOR2 (N10857, N10844, N206);
buf BUF1 (N10858, N10845);
nor NOR4 (N10859, N10851, N4620, N4780, N5443);
buf BUF1 (N10860, N10856);
xor XOR2 (N10861, N10860, N504);
nor NOR4 (N10862, N10852, N181, N167, N1864);
nand NAND3 (N10863, N10848, N3595, N2620);
not NOT1 (N10864, N10854);
and AND3 (N10865, N10857, N9073, N4236);
or OR3 (N10866, N10864, N1504, N4835);
or OR3 (N10867, N10861, N3447, N8828);
xor XOR2 (N10868, N10867, N9940);
not NOT1 (N10869, N10868);
nand NAND4 (N10870, N10865, N2755, N7168, N5789);
buf BUF1 (N10871, N10847);
or OR2 (N10872, N10858, N2354);
nand NAND4 (N10873, N10862, N2649, N2670, N2048);
nor NOR2 (N10874, N10863, N2203);
buf BUF1 (N10875, N10872);
nand NAND2 (N10876, N10869, N5022);
not NOT1 (N10877, N10874);
nor NOR4 (N10878, N10853, N8517, N3999, N8860);
xor XOR2 (N10879, N10873, N5023);
buf BUF1 (N10880, N10871);
and AND4 (N10881, N10876, N4546, N9474, N8050);
nor NOR4 (N10882, N10877, N5789, N315, N4825);
not NOT1 (N10883, N10866);
and AND3 (N10884, N10880, N1667, N1605);
xor XOR2 (N10885, N10878, N10479);
nor NOR2 (N10886, N10882, N1092);
or OR2 (N10887, N10859, N82);
nor NOR2 (N10888, N10875, N939);
nor NOR4 (N10889, N10879, N3441, N4815, N10272);
and AND4 (N10890, N10887, N10656, N4018, N8449);
xor XOR2 (N10891, N10855, N3951);
xor XOR2 (N10892, N10888, N887);
nor NOR4 (N10893, N10885, N9996, N2524, N4408);
nor NOR2 (N10894, N10881, N1053);
nor NOR2 (N10895, N10891, N3062);
buf BUF1 (N10896, N10894);
nor NOR2 (N10897, N10895, N9828);
not NOT1 (N10898, N10883);
nor NOR3 (N10899, N10892, N8464, N8701);
buf BUF1 (N10900, N10886);
and AND2 (N10901, N10889, N3539);
not NOT1 (N10902, N10884);
xor XOR2 (N10903, N10902, N2784);
or OR4 (N10904, N10897, N1265, N4692, N9734);
nand NAND3 (N10905, N10903, N5410, N10224);
nor NOR2 (N10906, N10870, N9456);
buf BUF1 (N10907, N10896);
xor XOR2 (N10908, N10905, N3359);
buf BUF1 (N10909, N10901);
and AND4 (N10910, N10900, N1333, N6218, N8382);
nor NOR2 (N10911, N10906, N10051);
nand NAND2 (N10912, N10908, N6247);
not NOT1 (N10913, N10890);
nand NAND2 (N10914, N10893, N3619);
nand NAND3 (N10915, N10907, N1703, N9897);
not NOT1 (N10916, N10910);
nand NAND3 (N10917, N10912, N1535, N2519);
and AND3 (N10918, N10916, N1374, N4805);
xor XOR2 (N10919, N10909, N7845);
not NOT1 (N10920, N10915);
buf BUF1 (N10921, N10914);
nor NOR4 (N10922, N10913, N625, N375, N9415);
and AND3 (N10923, N10918, N894, N9867);
xor XOR2 (N10924, N10917, N10455);
xor XOR2 (N10925, N10899, N7686);
nor NOR3 (N10926, N10925, N2502, N2832);
not NOT1 (N10927, N10926);
and AND2 (N10928, N10898, N5779);
or OR4 (N10929, N10919, N7404, N10218, N10804);
not NOT1 (N10930, N10928);
nand NAND2 (N10931, N10911, N1425);
nand NAND3 (N10932, N10927, N8887, N1009);
buf BUF1 (N10933, N10930);
not NOT1 (N10934, N10920);
not NOT1 (N10935, N10933);
xor XOR2 (N10936, N10904, N6967);
buf BUF1 (N10937, N10936);
or OR4 (N10938, N10932, N5071, N10229, N4812);
not NOT1 (N10939, N10938);
not NOT1 (N10940, N10934);
not NOT1 (N10941, N10939);
not NOT1 (N10942, N10935);
nor NOR2 (N10943, N10929, N6357);
and AND2 (N10944, N10922, N8460);
nand NAND4 (N10945, N10924, N1507, N8099, N6831);
not NOT1 (N10946, N10940);
xor XOR2 (N10947, N10931, N4836);
not NOT1 (N10948, N10923);
xor XOR2 (N10949, N10947, N4551);
xor XOR2 (N10950, N10948, N1430);
and AND4 (N10951, N10942, N10084, N10405, N817);
nand NAND4 (N10952, N10945, N6533, N5653, N1235);
nor NOR2 (N10953, N10946, N10400);
nor NOR4 (N10954, N10943, N10589, N9092, N6463);
not NOT1 (N10955, N10944);
nor NOR2 (N10956, N10953, N5164);
and AND4 (N10957, N10956, N2827, N3757, N5259);
buf BUF1 (N10958, N10955);
and AND2 (N10959, N10937, N5967);
or OR3 (N10960, N10921, N5014, N1243);
nand NAND4 (N10961, N10957, N5494, N2249, N2839);
buf BUF1 (N10962, N10949);
nor NOR4 (N10963, N10958, N2607, N8381, N1754);
and AND4 (N10964, N10950, N5935, N8799, N9331);
nand NAND3 (N10965, N10962, N1648, N1022);
nor NOR3 (N10966, N10959, N1903, N9298);
xor XOR2 (N10967, N10961, N7664);
buf BUF1 (N10968, N10965);
or OR4 (N10969, N10951, N8941, N6529, N1162);
xor XOR2 (N10970, N10968, N130);
nand NAND4 (N10971, N10954, N10167, N81, N2266);
and AND3 (N10972, N10969, N4618, N9429);
nand NAND4 (N10973, N10941, N3905, N1484, N49);
xor XOR2 (N10974, N10952, N818);
not NOT1 (N10975, N10972);
nand NAND3 (N10976, N10967, N6909, N8318);
buf BUF1 (N10977, N10964);
nand NAND2 (N10978, N10975, N7715);
and AND4 (N10979, N10960, N2335, N9291, N3501);
xor XOR2 (N10980, N10970, N1247);
and AND4 (N10981, N10974, N5892, N3265, N7014);
not NOT1 (N10982, N10973);
nand NAND3 (N10983, N10981, N2610, N10841);
and AND4 (N10984, N10983, N4738, N8147, N5009);
nand NAND4 (N10985, N10963, N5333, N5625, N4880);
nand NAND4 (N10986, N10966, N6781, N8347, N10855);
nor NOR3 (N10987, N10971, N678, N3733);
nor NOR2 (N10988, N10987, N3715);
or OR2 (N10989, N10980, N5147);
or OR3 (N10990, N10978, N7382, N3933);
buf BUF1 (N10991, N10985);
and AND3 (N10992, N10988, N7696, N4301);
xor XOR2 (N10993, N10989, N8806);
and AND3 (N10994, N10982, N9611, N8913);
and AND4 (N10995, N10984, N5117, N368, N4650);
nand NAND4 (N10996, N10977, N10784, N7442, N1854);
and AND3 (N10997, N10995, N4943, N3923);
not NOT1 (N10998, N10979);
and AND3 (N10999, N10986, N8998, N3389);
not NOT1 (N11000, N10976);
and AND2 (N11001, N10992, N1087);
and AND2 (N11002, N10998, N9312);
nor NOR3 (N11003, N10991, N7448, N2257);
nor NOR3 (N11004, N10999, N2770, N3218);
and AND2 (N11005, N11003, N5620);
and AND2 (N11006, N11002, N10220);
xor XOR2 (N11007, N10994, N5829);
and AND3 (N11008, N11007, N6209, N10039);
buf BUF1 (N11009, N11001);
nor NOR2 (N11010, N10990, N3193);
and AND4 (N11011, N10996, N9583, N3895, N3890);
and AND3 (N11012, N11005, N10119, N8866);
or OR3 (N11013, N11009, N5098, N2021);
and AND2 (N11014, N11013, N645);
nor NOR2 (N11015, N11012, N5673);
nand NAND2 (N11016, N10993, N7179);
nand NAND2 (N11017, N11016, N6432);
nand NAND4 (N11018, N11000, N3898, N3244, N7964);
and AND4 (N11019, N10997, N8214, N6451, N5537);
buf BUF1 (N11020, N11014);
not NOT1 (N11021, N11019);
not NOT1 (N11022, N11011);
xor XOR2 (N11023, N11006, N5231);
xor XOR2 (N11024, N11008, N6353);
and AND3 (N11025, N11022, N6677, N1290);
nor NOR2 (N11026, N11018, N1671);
or OR3 (N11027, N11010, N2565, N18);
or OR3 (N11028, N11027, N2235, N3380);
or OR3 (N11029, N11020, N10010, N1060);
buf BUF1 (N11030, N11023);
xor XOR2 (N11031, N11030, N8543);
buf BUF1 (N11032, N11004);
nor NOR3 (N11033, N11028, N10997, N1919);
not NOT1 (N11034, N11026);
and AND4 (N11035, N11015, N2815, N2660, N2934);
buf BUF1 (N11036, N11033);
buf BUF1 (N11037, N11029);
xor XOR2 (N11038, N11017, N1824);
xor XOR2 (N11039, N11025, N1881);
xor XOR2 (N11040, N11039, N9508);
nand NAND4 (N11041, N11034, N365, N10014, N1393);
not NOT1 (N11042, N11040);
nand NAND3 (N11043, N11036, N5135, N6598);
xor XOR2 (N11044, N11035, N7237);
and AND4 (N11045, N11032, N8810, N7188, N7636);
buf BUF1 (N11046, N11044);
and AND3 (N11047, N11024, N219, N9246);
xor XOR2 (N11048, N11042, N1406);
not NOT1 (N11049, N11047);
not NOT1 (N11050, N11048);
or OR4 (N11051, N11043, N10821, N6705, N3187);
or OR2 (N11052, N11031, N3210);
or OR4 (N11053, N11021, N1299, N1814, N8365);
buf BUF1 (N11054, N11051);
nand NAND2 (N11055, N11046, N10958);
not NOT1 (N11056, N11055);
buf BUF1 (N11057, N11056);
buf BUF1 (N11058, N11052);
and AND3 (N11059, N11041, N4205, N1635);
xor XOR2 (N11060, N11054, N53);
and AND2 (N11061, N11057, N4470);
buf BUF1 (N11062, N11049);
nand NAND3 (N11063, N11062, N2831, N2695);
nor NOR4 (N11064, N11050, N3195, N4426, N7085);
nor NOR2 (N11065, N11037, N9267);
not NOT1 (N11066, N11063);
and AND2 (N11067, N11058, N783);
not NOT1 (N11068, N11060);
or OR2 (N11069, N11053, N8249);
and AND4 (N11070, N11045, N5528, N5897, N7594);
or OR2 (N11071, N11066, N10981);
and AND2 (N11072, N11061, N3938);
or OR3 (N11073, N11038, N1230, N6765);
and AND4 (N11074, N11070, N9278, N3116, N10233);
nand NAND4 (N11075, N11059, N1164, N5073, N4219);
buf BUF1 (N11076, N11067);
xor XOR2 (N11077, N11069, N2690);
or OR4 (N11078, N11068, N6272, N11033, N105);
buf BUF1 (N11079, N11074);
xor XOR2 (N11080, N11077, N8157);
not NOT1 (N11081, N11064);
not NOT1 (N11082, N11080);
buf BUF1 (N11083, N11065);
xor XOR2 (N11084, N11073, N11054);
and AND2 (N11085, N11084, N9285);
or OR4 (N11086, N11085, N5151, N6259, N713);
nand NAND2 (N11087, N11076, N9649);
nand NAND2 (N11088, N11072, N185);
not NOT1 (N11089, N11075);
not NOT1 (N11090, N11086);
or OR3 (N11091, N11088, N2805, N2253);
xor XOR2 (N11092, N11087, N3379);
not NOT1 (N11093, N11071);
nand NAND3 (N11094, N11082, N10623, N370);
buf BUF1 (N11095, N11083);
and AND3 (N11096, N11093, N1676, N6227);
nand NAND2 (N11097, N11078, N10907);
or OR4 (N11098, N11095, N163, N8736, N1945);
nand NAND4 (N11099, N11089, N3691, N937, N10017);
not NOT1 (N11100, N11099);
not NOT1 (N11101, N11098);
nand NAND3 (N11102, N11091, N6027, N833);
nor NOR3 (N11103, N11081, N4609, N3535);
or OR3 (N11104, N11096, N9240, N684);
buf BUF1 (N11105, N11102);
not NOT1 (N11106, N11103);
not NOT1 (N11107, N11106);
or OR3 (N11108, N11090, N6807, N5694);
xor XOR2 (N11109, N11101, N2284);
and AND3 (N11110, N11105, N1344, N9846);
nand NAND2 (N11111, N11109, N4874);
or OR2 (N11112, N11079, N1945);
nor NOR3 (N11113, N11111, N1623, N10886);
nor NOR3 (N11114, N11107, N5480, N1347);
not NOT1 (N11115, N11114);
nor NOR4 (N11116, N11115, N4579, N10980, N2401);
xor XOR2 (N11117, N11097, N5570);
or OR3 (N11118, N11112, N6590, N8304);
nor NOR3 (N11119, N11113, N2378, N8433);
nor NOR3 (N11120, N11108, N4214, N6949);
nor NOR4 (N11121, N11104, N8683, N7341, N8543);
not NOT1 (N11122, N11094);
nand NAND2 (N11123, N11120, N5731);
buf BUF1 (N11124, N11092);
and AND4 (N11125, N11121, N8791, N4083, N4429);
nor NOR3 (N11126, N11123, N10596, N9059);
not NOT1 (N11127, N11125);
xor XOR2 (N11128, N11126, N2651);
nor NOR3 (N11129, N11128, N481, N5259);
nand NAND3 (N11130, N11129, N6436, N1930);
and AND2 (N11131, N11124, N3954);
xor XOR2 (N11132, N11122, N3429);
nor NOR3 (N11133, N11117, N10498, N6197);
buf BUF1 (N11134, N11116);
buf BUF1 (N11135, N11130);
or OR4 (N11136, N11119, N2956, N5351, N3796);
not NOT1 (N11137, N11100);
or OR3 (N11138, N11127, N10135, N7505);
xor XOR2 (N11139, N11132, N4808);
xor XOR2 (N11140, N11135, N2636);
not NOT1 (N11141, N11110);
nand NAND2 (N11142, N11136, N10219);
buf BUF1 (N11143, N11142);
not NOT1 (N11144, N11137);
xor XOR2 (N11145, N11118, N4370);
nand NAND3 (N11146, N11133, N3803, N6106);
and AND4 (N11147, N11138, N6121, N3397, N1260);
nor NOR4 (N11148, N11134, N319, N282, N9611);
buf BUF1 (N11149, N11140);
xor XOR2 (N11150, N11147, N1384);
nand NAND4 (N11151, N11131, N7434, N10262, N4546);
not NOT1 (N11152, N11141);
not NOT1 (N11153, N11139);
xor XOR2 (N11154, N11148, N6763);
not NOT1 (N11155, N11146);
nand NAND3 (N11156, N11153, N5207, N10921);
nor NOR2 (N11157, N11155, N3849);
buf BUF1 (N11158, N11151);
or OR3 (N11159, N11157, N9414, N866);
and AND4 (N11160, N11158, N3856, N8890, N11098);
and AND4 (N11161, N11154, N5577, N9088, N4406);
nor NOR4 (N11162, N11161, N11144, N9375, N7265);
nand NAND2 (N11163, N913, N8170);
and AND2 (N11164, N11149, N8329);
or OR3 (N11165, N11156, N6343, N2675);
not NOT1 (N11166, N11145);
xor XOR2 (N11167, N11160, N4051);
and AND4 (N11168, N11167, N7046, N494, N5225);
or OR2 (N11169, N11166, N5893);
buf BUF1 (N11170, N11159);
or OR4 (N11171, N11168, N3324, N4132, N5705);
nand NAND3 (N11172, N11162, N6306, N5888);
and AND4 (N11173, N11170, N1329, N9090, N4795);
nor NOR2 (N11174, N11164, N4217);
xor XOR2 (N11175, N11171, N1283);
and AND4 (N11176, N11174, N10625, N6476, N5823);
not NOT1 (N11177, N11165);
not NOT1 (N11178, N11143);
nor NOR3 (N11179, N11152, N3339, N6249);
and AND2 (N11180, N11178, N6566);
nor NOR3 (N11181, N11180, N10672, N5129);
nand NAND4 (N11182, N11169, N8234, N4699, N6833);
and AND3 (N11183, N11173, N7101, N6844);
xor XOR2 (N11184, N11176, N8835);
nor NOR4 (N11185, N11183, N5271, N6311, N5441);
xor XOR2 (N11186, N11182, N1022);
xor XOR2 (N11187, N11177, N6676);
or OR3 (N11188, N11185, N7906, N5217);
and AND2 (N11189, N11150, N1678);
buf BUF1 (N11190, N11172);
or OR2 (N11191, N11190, N1967);
xor XOR2 (N11192, N11184, N10838);
buf BUF1 (N11193, N11189);
xor XOR2 (N11194, N11175, N3658);
not NOT1 (N11195, N11181);
and AND4 (N11196, N11193, N10873, N2093, N2701);
nand NAND2 (N11197, N11192, N9900);
not NOT1 (N11198, N11191);
or OR4 (N11199, N11188, N9216, N1262, N2476);
nor NOR3 (N11200, N11199, N595, N5997);
or OR3 (N11201, N11198, N7501, N9547);
nor NOR4 (N11202, N11179, N9175, N4424, N5904);
and AND2 (N11203, N11195, N7943);
xor XOR2 (N11204, N11200, N2231);
buf BUF1 (N11205, N11201);
nor NOR2 (N11206, N11204, N8603);
and AND3 (N11207, N11205, N9412, N9247);
nand NAND3 (N11208, N11197, N196, N6670);
not NOT1 (N11209, N11187);
xor XOR2 (N11210, N11208, N2212);
or OR2 (N11211, N11196, N909);
buf BUF1 (N11212, N11163);
not NOT1 (N11213, N11186);
nor NOR4 (N11214, N11212, N9799, N5290, N3324);
nand NAND2 (N11215, N11194, N6952);
not NOT1 (N11216, N11215);
nor NOR4 (N11217, N11207, N5027, N7111, N5531);
nand NAND4 (N11218, N11202, N9431, N6430, N3988);
or OR3 (N11219, N11211, N2638, N3470);
xor XOR2 (N11220, N11218, N2900);
and AND4 (N11221, N11213, N7664, N5757, N4378);
nand NAND4 (N11222, N11206, N3527, N7861, N1628);
xor XOR2 (N11223, N11216, N10875);
nor NOR4 (N11224, N11209, N8071, N3196, N7475);
and AND2 (N11225, N11223, N1821);
and AND4 (N11226, N11221, N2448, N4178, N307);
nand NAND2 (N11227, N11224, N5684);
not NOT1 (N11228, N11220);
buf BUF1 (N11229, N11217);
nor NOR3 (N11230, N11227, N2, N5397);
and AND2 (N11231, N11228, N11174);
not NOT1 (N11232, N11210);
xor XOR2 (N11233, N11219, N231);
and AND4 (N11234, N11231, N2537, N10405, N1658);
not NOT1 (N11235, N11226);
xor XOR2 (N11236, N11232, N4591);
xor XOR2 (N11237, N11230, N1813);
and AND3 (N11238, N11236, N1774, N6645);
or OR4 (N11239, N11235, N8904, N2579, N9735);
or OR4 (N11240, N11234, N823, N1029, N9082);
buf BUF1 (N11241, N11239);
and AND4 (N11242, N11233, N9030, N7985, N4686);
nor NOR2 (N11243, N11225, N4902);
or OR2 (N11244, N11240, N4966);
and AND2 (N11245, N11222, N189);
nor NOR4 (N11246, N11229, N8024, N1043, N745);
or OR4 (N11247, N11242, N4865, N7182, N671);
and AND2 (N11248, N11244, N6582);
or OR2 (N11249, N11237, N1819);
nand NAND3 (N11250, N11243, N3612, N8018);
and AND3 (N11251, N11238, N8783, N6310);
not NOT1 (N11252, N11249);
or OR4 (N11253, N11251, N8608, N1308, N8943);
nor NOR4 (N11254, N11248, N6557, N2038, N9822);
not NOT1 (N11255, N11246);
and AND2 (N11256, N11250, N5916);
nor NOR4 (N11257, N11245, N7784, N7178, N10343);
nand NAND2 (N11258, N11252, N3057);
nor NOR4 (N11259, N11247, N1964, N11051, N4853);
and AND3 (N11260, N11253, N2841, N1335);
xor XOR2 (N11261, N11203, N11226);
nor NOR2 (N11262, N11256, N212);
nor NOR4 (N11263, N11258, N8077, N7426, N7718);
not NOT1 (N11264, N11214);
and AND3 (N11265, N11257, N731, N5689);
not NOT1 (N11266, N11265);
not NOT1 (N11267, N11264);
or OR4 (N11268, N11266, N6651, N8576, N10233);
or OR4 (N11269, N11268, N2099, N1854, N8413);
xor XOR2 (N11270, N11254, N10736);
not NOT1 (N11271, N11263);
nor NOR2 (N11272, N11255, N1162);
xor XOR2 (N11273, N11269, N10637);
buf BUF1 (N11274, N11272);
or OR3 (N11275, N11273, N9983, N1260);
xor XOR2 (N11276, N11241, N4368);
and AND2 (N11277, N11270, N2606);
nand NAND3 (N11278, N11260, N9472, N2417);
xor XOR2 (N11279, N11271, N10790);
and AND3 (N11280, N11279, N5994, N5119);
nor NOR2 (N11281, N11267, N335);
nand NAND4 (N11282, N11277, N3955, N6495, N10289);
nand NAND3 (N11283, N11276, N2216, N6835);
buf BUF1 (N11284, N11278);
xor XOR2 (N11285, N11259, N2226);
xor XOR2 (N11286, N11283, N9340);
xor XOR2 (N11287, N11275, N157);
and AND3 (N11288, N11274, N2094, N1602);
nand NAND3 (N11289, N11262, N2008, N9354);
or OR3 (N11290, N11284, N1812, N6756);
nand NAND4 (N11291, N11280, N3019, N5493, N1118);
nand NAND4 (N11292, N11281, N9746, N7242, N6431);
and AND3 (N11293, N11282, N286, N628);
nand NAND3 (N11294, N11292, N8442, N5656);
buf BUF1 (N11295, N11288);
or OR2 (N11296, N11289, N7229);
not NOT1 (N11297, N11261);
and AND2 (N11298, N11297, N10883);
or OR3 (N11299, N11287, N6454, N6205);
buf BUF1 (N11300, N11296);
xor XOR2 (N11301, N11293, N353);
not NOT1 (N11302, N11299);
and AND3 (N11303, N11298, N7953, N8249);
or OR2 (N11304, N11290, N10639);
nand NAND4 (N11305, N11295, N476, N4243, N5733);
nor NOR2 (N11306, N11305, N6384);
nand NAND2 (N11307, N11303, N8374);
nor NOR2 (N11308, N11306, N10528);
nor NOR3 (N11309, N11300, N9967, N8541);
nor NOR2 (N11310, N11294, N2295);
nor NOR2 (N11311, N11310, N4461);
nor NOR2 (N11312, N11301, N5162);
xor XOR2 (N11313, N11286, N10221);
not NOT1 (N11314, N11312);
xor XOR2 (N11315, N11313, N934);
nor NOR2 (N11316, N11302, N9019);
buf BUF1 (N11317, N11304);
nor NOR2 (N11318, N11309, N3145);
buf BUF1 (N11319, N11307);
nor NOR3 (N11320, N11311, N8713, N2170);
or OR4 (N11321, N11314, N6985, N5803, N1031);
and AND3 (N11322, N11291, N10952, N9338);
or OR4 (N11323, N11319, N6292, N1070, N9463);
xor XOR2 (N11324, N11322, N10229);
or OR2 (N11325, N11316, N2219);
buf BUF1 (N11326, N11315);
or OR3 (N11327, N11318, N1908, N2749);
or OR3 (N11328, N11308, N1386, N6743);
and AND4 (N11329, N11317, N528, N8467, N5257);
not NOT1 (N11330, N11285);
nor NOR3 (N11331, N11327, N10650, N3907);
or OR4 (N11332, N11331, N3583, N5168, N9040);
buf BUF1 (N11333, N11324);
nand NAND4 (N11334, N11330, N7909, N4389, N9864);
buf BUF1 (N11335, N11328);
or OR2 (N11336, N11335, N3453);
or OR2 (N11337, N11334, N3223);
nand NAND3 (N11338, N11321, N2683, N8558);
nand NAND4 (N11339, N11329, N2792, N10162, N6470);
or OR2 (N11340, N11337, N5698);
xor XOR2 (N11341, N11339, N4220);
or OR2 (N11342, N11333, N332);
or OR4 (N11343, N11332, N1391, N2441, N9695);
xor XOR2 (N11344, N11320, N2808);
or OR3 (N11345, N11336, N5992, N7857);
or OR4 (N11346, N11341, N4097, N8127, N10668);
nor NOR3 (N11347, N11338, N5208, N7067);
buf BUF1 (N11348, N11340);
or OR2 (N11349, N11325, N9107);
not NOT1 (N11350, N11345);
nor NOR3 (N11351, N11323, N1794, N11166);
buf BUF1 (N11352, N11344);
xor XOR2 (N11353, N11346, N8474);
buf BUF1 (N11354, N11348);
not NOT1 (N11355, N11354);
buf BUF1 (N11356, N11355);
buf BUF1 (N11357, N11356);
not NOT1 (N11358, N11352);
xor XOR2 (N11359, N11357, N957);
nand NAND2 (N11360, N11359, N7219);
nor NOR3 (N11361, N11347, N2125, N5691);
or OR3 (N11362, N11349, N7943, N3308);
not NOT1 (N11363, N11343);
nand NAND2 (N11364, N11358, N6448);
buf BUF1 (N11365, N11360);
nor NOR2 (N11366, N11342, N4591);
nand NAND4 (N11367, N11366, N1736, N7911, N4285);
xor XOR2 (N11368, N11351, N8074);
and AND4 (N11369, N11367, N851, N10329, N8241);
buf BUF1 (N11370, N11326);
not NOT1 (N11371, N11365);
buf BUF1 (N11372, N11368);
and AND4 (N11373, N11364, N6838, N5811, N7889);
and AND4 (N11374, N11372, N2427, N2036, N9291);
nor NOR2 (N11375, N11371, N5904);
and AND2 (N11376, N11373, N1975);
or OR3 (N11377, N11361, N2672, N7509);
not NOT1 (N11378, N11377);
buf BUF1 (N11379, N11374);
nor NOR2 (N11380, N11379, N6922);
or OR3 (N11381, N11376, N10559, N62);
nand NAND3 (N11382, N11362, N4664, N10392);
not NOT1 (N11383, N11382);
or OR2 (N11384, N11381, N8182);
or OR4 (N11385, N11353, N10773, N7742, N7395);
not NOT1 (N11386, N11385);
or OR4 (N11387, N11363, N5818, N4664, N1772);
nor NOR2 (N11388, N11384, N2810);
nor NOR2 (N11389, N11386, N10015);
buf BUF1 (N11390, N11370);
and AND2 (N11391, N11387, N10401);
not NOT1 (N11392, N11375);
not NOT1 (N11393, N11350);
nand NAND3 (N11394, N11393, N7707, N3979);
nand NAND4 (N11395, N11369, N6040, N5710, N3146);
not NOT1 (N11396, N11394);
nor NOR3 (N11397, N11389, N8017, N1944);
xor XOR2 (N11398, N11380, N7256);
xor XOR2 (N11399, N11397, N2462);
nand NAND4 (N11400, N11399, N8366, N8444, N5872);
nor NOR3 (N11401, N11395, N1020, N4433);
not NOT1 (N11402, N11383);
or OR4 (N11403, N11401, N9046, N10968, N9964);
xor XOR2 (N11404, N11388, N3424);
not NOT1 (N11405, N11403);
nor NOR2 (N11406, N11398, N2419);
nor NOR3 (N11407, N11391, N7171, N4365);
nand NAND2 (N11408, N11404, N5149);
buf BUF1 (N11409, N11407);
not NOT1 (N11410, N11396);
xor XOR2 (N11411, N11400, N310);
and AND2 (N11412, N11408, N2658);
or OR2 (N11413, N11410, N3051);
xor XOR2 (N11414, N11412, N2919);
and AND3 (N11415, N11392, N950, N8151);
not NOT1 (N11416, N11415);
buf BUF1 (N11417, N11402);
not NOT1 (N11418, N11416);
nand NAND2 (N11419, N11390, N5719);
not NOT1 (N11420, N11417);
not NOT1 (N11421, N11420);
nand NAND3 (N11422, N11413, N10426, N7126);
and AND3 (N11423, N11414, N1220, N4961);
nand NAND2 (N11424, N11418, N5225);
buf BUF1 (N11425, N11421);
or OR2 (N11426, N11409, N6268);
and AND4 (N11427, N11424, N4475, N7693, N7973);
not NOT1 (N11428, N11378);
buf BUF1 (N11429, N11428);
nor NOR2 (N11430, N11425, N7647);
nor NOR3 (N11431, N11423, N10795, N8896);
xor XOR2 (N11432, N11431, N6850);
nor NOR4 (N11433, N11419, N2072, N1140, N597);
or OR3 (N11434, N11405, N6280, N979);
not NOT1 (N11435, N11422);
xor XOR2 (N11436, N11427, N3486);
or OR4 (N11437, N11406, N1311, N5338, N8875);
and AND4 (N11438, N11411, N261, N7547, N10301);
nor NOR3 (N11439, N11430, N10142, N357);
or OR4 (N11440, N11438, N5345, N6979, N631);
buf BUF1 (N11441, N11426);
nand NAND3 (N11442, N11434, N6688, N4318);
not NOT1 (N11443, N11433);
and AND3 (N11444, N11441, N2663, N8982);
buf BUF1 (N11445, N11442);
xor XOR2 (N11446, N11432, N8595);
and AND4 (N11447, N11436, N3882, N3549, N7019);
and AND2 (N11448, N11435, N7448);
nor NOR2 (N11449, N11448, N10627);
or OR2 (N11450, N11449, N519);
xor XOR2 (N11451, N11445, N6765);
or OR2 (N11452, N11451, N3374);
buf BUF1 (N11453, N11440);
xor XOR2 (N11454, N11447, N2522);
nor NOR3 (N11455, N11453, N8939, N2983);
and AND4 (N11456, N11437, N662, N6517, N1137);
nor NOR4 (N11457, N11429, N869, N10612, N5788);
buf BUF1 (N11458, N11443);
not NOT1 (N11459, N11444);
nor NOR4 (N11460, N11455, N1786, N6780, N1145);
or OR4 (N11461, N11454, N410, N6981, N4109);
and AND4 (N11462, N11450, N3526, N7402, N10452);
or OR4 (N11463, N11460, N9057, N3500, N11394);
not NOT1 (N11464, N11461);
xor XOR2 (N11465, N11462, N10724);
nor NOR2 (N11466, N11457, N3992);
and AND2 (N11467, N11459, N1505);
nor NOR3 (N11468, N11463, N5797, N7718);
not NOT1 (N11469, N11458);
xor XOR2 (N11470, N11469, N9089);
or OR4 (N11471, N11456, N4893, N10010, N6752);
and AND2 (N11472, N11465, N9100);
nand NAND3 (N11473, N11470, N2942, N7127);
not NOT1 (N11474, N11467);
and AND3 (N11475, N11466, N8411, N8152);
and AND2 (N11476, N11474, N9830);
xor XOR2 (N11477, N11446, N7242);
not NOT1 (N11478, N11476);
buf BUF1 (N11479, N11468);
or OR2 (N11480, N11452, N3345);
buf BUF1 (N11481, N11439);
nor NOR4 (N11482, N11472, N1876, N9111, N9993);
and AND2 (N11483, N11471, N502);
or OR3 (N11484, N11481, N3485, N2250);
nor NOR2 (N11485, N11464, N4344);
and AND4 (N11486, N11484, N8476, N3893, N4727);
xor XOR2 (N11487, N11480, N8370);
xor XOR2 (N11488, N11475, N10320);
or OR3 (N11489, N11473, N5947, N1799);
nor NOR4 (N11490, N11482, N3531, N2609, N5436);
not NOT1 (N11491, N11479);
and AND2 (N11492, N11485, N6550);
nor NOR2 (N11493, N11489, N7203);
or OR2 (N11494, N11493, N8408);
nor NOR2 (N11495, N11491, N1212);
nor NOR3 (N11496, N11488, N3092, N2071);
nand NAND2 (N11497, N11490, N9402);
and AND4 (N11498, N11497, N9340, N157, N239);
nand NAND3 (N11499, N11478, N10406, N6145);
nand NAND4 (N11500, N11494, N10787, N780, N10797);
not NOT1 (N11501, N11495);
nor NOR3 (N11502, N11477, N6168, N2610);
xor XOR2 (N11503, N11492, N554);
not NOT1 (N11504, N11496);
and AND3 (N11505, N11503, N548, N10480);
xor XOR2 (N11506, N11487, N1745);
or OR2 (N11507, N11506, N5812);
or OR4 (N11508, N11502, N4219, N1564, N609);
and AND2 (N11509, N11498, N11429);
not NOT1 (N11510, N11504);
and AND2 (N11511, N11501, N917);
nor NOR2 (N11512, N11483, N10226);
buf BUF1 (N11513, N11505);
nor NOR2 (N11514, N11512, N2653);
xor XOR2 (N11515, N11509, N6013);
buf BUF1 (N11516, N11514);
xor XOR2 (N11517, N11515, N8388);
or OR3 (N11518, N11499, N910, N10454);
and AND4 (N11519, N11517, N1382, N11107, N9687);
xor XOR2 (N11520, N11508, N3623);
buf BUF1 (N11521, N11516);
xor XOR2 (N11522, N11521, N498);
not NOT1 (N11523, N11507);
nor NOR2 (N11524, N11523, N4780);
not NOT1 (N11525, N11500);
xor XOR2 (N11526, N11519, N5707);
not NOT1 (N11527, N11518);
nand NAND4 (N11528, N11527, N721, N5865, N3227);
not NOT1 (N11529, N11520);
buf BUF1 (N11530, N11511);
nand NAND3 (N11531, N11510, N6358, N9970);
buf BUF1 (N11532, N11528);
buf BUF1 (N11533, N11529);
or OR3 (N11534, N11486, N5591, N7029);
and AND4 (N11535, N11524, N6525, N10994, N9292);
nor NOR2 (N11536, N11534, N2770);
not NOT1 (N11537, N11533);
nand NAND2 (N11538, N11513, N7904);
nand NAND4 (N11539, N11530, N6597, N84, N7913);
buf BUF1 (N11540, N11539);
nand NAND4 (N11541, N11537, N1774, N7844, N7987);
or OR2 (N11542, N11536, N2424);
nor NOR3 (N11543, N11531, N516, N10020);
and AND4 (N11544, N11522, N2067, N2760, N4196);
and AND2 (N11545, N11540, N2329);
nand NAND4 (N11546, N11532, N8851, N10493, N6636);
nor NOR4 (N11547, N11525, N8794, N1499, N5903);
and AND3 (N11548, N11541, N4586, N2629);
xor XOR2 (N11549, N11526, N996);
nand NAND4 (N11550, N11549, N2892, N6488, N1404);
and AND2 (N11551, N11538, N3261);
and AND4 (N11552, N11535, N4958, N596, N3236);
or OR2 (N11553, N11550, N11246);
not NOT1 (N11554, N11543);
not NOT1 (N11555, N11552);
xor XOR2 (N11556, N11548, N3847);
buf BUF1 (N11557, N11551);
nor NOR4 (N11558, N11544, N2476, N11426, N7125);
xor XOR2 (N11559, N11556, N10149);
not NOT1 (N11560, N11553);
and AND4 (N11561, N11545, N8398, N4308, N1388);
or OR4 (N11562, N11560, N342, N3048, N382);
or OR4 (N11563, N11559, N1694, N8684, N6839);
xor XOR2 (N11564, N11546, N3547);
not NOT1 (N11565, N11554);
and AND2 (N11566, N11558, N4763);
and AND4 (N11567, N11563, N7052, N7923, N6058);
and AND3 (N11568, N11542, N3530, N10405);
and AND2 (N11569, N11565, N10387);
or OR4 (N11570, N11547, N5158, N9037, N1323);
or OR3 (N11571, N11566, N1633, N4829);
not NOT1 (N11572, N11561);
nand NAND4 (N11573, N11572, N10150, N8382, N5855);
nand NAND4 (N11574, N11562, N602, N4802, N8350);
or OR2 (N11575, N11574, N3965);
nand NAND3 (N11576, N11557, N1629, N1243);
and AND3 (N11577, N11567, N9749, N5013);
xor XOR2 (N11578, N11573, N1915);
nor NOR2 (N11579, N11576, N6849);
xor XOR2 (N11580, N11568, N1383);
nor NOR4 (N11581, N11580, N107, N335, N9984);
xor XOR2 (N11582, N11579, N4472);
or OR3 (N11583, N11578, N3123, N10271);
or OR4 (N11584, N11571, N1718, N6969, N8582);
nor NOR2 (N11585, N11577, N913);
nor NOR4 (N11586, N11575, N2639, N3821, N3858);
xor XOR2 (N11587, N11583, N10306);
and AND2 (N11588, N11587, N9198);
and AND4 (N11589, N11581, N7460, N6037, N3506);
buf BUF1 (N11590, N11569);
nand NAND4 (N11591, N11570, N5197, N6820, N7505);
xor XOR2 (N11592, N11586, N11521);
nor NOR4 (N11593, N11582, N11052, N2337, N10630);
nor NOR4 (N11594, N11564, N7694, N4833, N2921);
or OR2 (N11595, N11591, N2631);
not NOT1 (N11596, N11594);
nand NAND2 (N11597, N11584, N2765);
or OR4 (N11598, N11590, N178, N2945, N9018);
buf BUF1 (N11599, N11593);
and AND2 (N11600, N11592, N3755);
or OR4 (N11601, N11596, N11117, N8669, N10346);
nor NOR3 (N11602, N11599, N5480, N2943);
buf BUF1 (N11603, N11597);
nand NAND4 (N11604, N11603, N5807, N8768, N4957);
xor XOR2 (N11605, N11555, N9963);
nor NOR3 (N11606, N11589, N9969, N1903);
or OR3 (N11607, N11605, N5674, N7824);
xor XOR2 (N11608, N11585, N10828);
buf BUF1 (N11609, N11588);
buf BUF1 (N11610, N11604);
or OR2 (N11611, N11600, N10454);
and AND2 (N11612, N11606, N5424);
nor NOR4 (N11613, N11601, N6028, N11147, N1644);
nand NAND2 (N11614, N11607, N11552);
not NOT1 (N11615, N11595);
and AND2 (N11616, N11609, N9542);
or OR3 (N11617, N11613, N5692, N6157);
or OR2 (N11618, N11610, N8735);
not NOT1 (N11619, N11618);
or OR4 (N11620, N11614, N8743, N4266, N334);
nor NOR4 (N11621, N11615, N3096, N9050, N8028);
and AND3 (N11622, N11598, N11132, N1531);
nor NOR2 (N11623, N11617, N10937);
nand NAND2 (N11624, N11621, N2850);
buf BUF1 (N11625, N11616);
xor XOR2 (N11626, N11608, N10962);
or OR2 (N11627, N11620, N202);
not NOT1 (N11628, N11623);
xor XOR2 (N11629, N11627, N1150);
nand NAND2 (N11630, N11625, N6053);
nand NAND2 (N11631, N11611, N7945);
nand NAND3 (N11632, N11628, N2255, N10375);
xor XOR2 (N11633, N11626, N4367);
not NOT1 (N11634, N11622);
not NOT1 (N11635, N11631);
buf BUF1 (N11636, N11632);
or OR2 (N11637, N11619, N4219);
xor XOR2 (N11638, N11633, N3513);
nand NAND4 (N11639, N11602, N7346, N1004, N4212);
not NOT1 (N11640, N11629);
not NOT1 (N11641, N11639);
xor XOR2 (N11642, N11624, N6699);
not NOT1 (N11643, N11637);
not NOT1 (N11644, N11638);
nand NAND3 (N11645, N11634, N135, N2388);
xor XOR2 (N11646, N11641, N8448);
xor XOR2 (N11647, N11646, N6979);
and AND3 (N11648, N11630, N5121, N7225);
nor NOR3 (N11649, N11636, N3973, N10964);
or OR3 (N11650, N11645, N4900, N2644);
buf BUF1 (N11651, N11635);
xor XOR2 (N11652, N11612, N4225);
xor XOR2 (N11653, N11640, N2749);
xor XOR2 (N11654, N11644, N2282);
buf BUF1 (N11655, N11649);
not NOT1 (N11656, N11650);
nor NOR4 (N11657, N11656, N11491, N9509, N2325);
not NOT1 (N11658, N11657);
and AND3 (N11659, N11655, N10566, N6537);
not NOT1 (N11660, N11651);
nor NOR3 (N11661, N11642, N7311, N2103);
and AND2 (N11662, N11660, N9983);
and AND4 (N11663, N11643, N3680, N7997, N3564);
and AND3 (N11664, N11653, N764, N9121);
or OR4 (N11665, N11664, N2453, N11630, N11157);
xor XOR2 (N11666, N11663, N10529);
or OR2 (N11667, N11647, N6807);
nand NAND3 (N11668, N11662, N2527, N2050);
buf BUF1 (N11669, N11659);
or OR3 (N11670, N11665, N4750, N5643);
and AND2 (N11671, N11652, N6604);
nand NAND3 (N11672, N11671, N5256, N6266);
buf BUF1 (N11673, N11666);
nor NOR2 (N11674, N11669, N10909);
buf BUF1 (N11675, N11661);
buf BUF1 (N11676, N11654);
and AND3 (N11677, N11674, N3861, N5547);
nor NOR2 (N11678, N11673, N7056);
and AND2 (N11679, N11668, N934);
xor XOR2 (N11680, N11676, N1279);
or OR2 (N11681, N11667, N11413);
nand NAND4 (N11682, N11670, N499, N9455, N8226);
buf BUF1 (N11683, N11677);
not NOT1 (N11684, N11679);
xor XOR2 (N11685, N11658, N9292);
xor XOR2 (N11686, N11680, N6221);
not NOT1 (N11687, N11672);
and AND4 (N11688, N11648, N5641, N7573, N2827);
and AND2 (N11689, N11678, N83);
nand NAND3 (N11690, N11686, N9777, N5207);
not NOT1 (N11691, N11684);
not NOT1 (N11692, N11675);
nand NAND4 (N11693, N11688, N608, N7456, N8589);
or OR3 (N11694, N11685, N1204, N6626);
and AND2 (N11695, N11690, N104);
nor NOR3 (N11696, N11692, N802, N5980);
nand NAND4 (N11697, N11687, N8606, N2290, N1484);
nand NAND2 (N11698, N11694, N8689);
not NOT1 (N11699, N11682);
and AND3 (N11700, N11693, N3380, N8898);
xor XOR2 (N11701, N11697, N755);
and AND3 (N11702, N11701, N6699, N7666);
and AND2 (N11703, N11691, N5780);
not NOT1 (N11704, N11683);
nand NAND2 (N11705, N11698, N7920);
buf BUF1 (N11706, N11704);
buf BUF1 (N11707, N11696);
nand NAND4 (N11708, N11703, N8308, N2250, N46);
nor NOR2 (N11709, N11699, N11129);
nor NOR3 (N11710, N11709, N693, N6273);
nor NOR4 (N11711, N11695, N1940, N5756, N3027);
buf BUF1 (N11712, N11702);
buf BUF1 (N11713, N11708);
xor XOR2 (N11714, N11706, N5389);
xor XOR2 (N11715, N11681, N203);
not NOT1 (N11716, N11715);
and AND2 (N11717, N11714, N337);
and AND3 (N11718, N11712, N5230, N1322);
not NOT1 (N11719, N11716);
and AND3 (N11720, N11707, N5286, N1177);
nand NAND4 (N11721, N11718, N3773, N66, N244);
not NOT1 (N11722, N11720);
or OR4 (N11723, N11689, N7627, N4921, N8708);
nor NOR4 (N11724, N11705, N10922, N5599, N9669);
not NOT1 (N11725, N11711);
xor XOR2 (N11726, N11713, N1091);
buf BUF1 (N11727, N11710);
buf BUF1 (N11728, N11723);
and AND4 (N11729, N11728, N5860, N9609, N11093);
nand NAND2 (N11730, N11722, N6121);
xor XOR2 (N11731, N11730, N6708);
nand NAND4 (N11732, N11724, N1817, N10332, N4676);
nor NOR3 (N11733, N11727, N1926, N5621);
nor NOR2 (N11734, N11732, N9524);
and AND2 (N11735, N11719, N7490);
nand NAND2 (N11736, N11733, N3518);
nand NAND4 (N11737, N11717, N2789, N7275, N8734);
or OR2 (N11738, N11726, N6136);
not NOT1 (N11739, N11734);
nand NAND3 (N11740, N11737, N9075, N8012);
buf BUF1 (N11741, N11700);
nand NAND3 (N11742, N11736, N547, N2007);
or OR4 (N11743, N11721, N8186, N7441, N4472);
nor NOR3 (N11744, N11739, N8347, N3954);
buf BUF1 (N11745, N11735);
nand NAND3 (N11746, N11731, N9381, N9621);
not NOT1 (N11747, N11738);
or OR2 (N11748, N11747, N5063);
or OR4 (N11749, N11740, N5593, N166, N7036);
xor XOR2 (N11750, N11743, N4812);
buf BUF1 (N11751, N11750);
buf BUF1 (N11752, N11729);
xor XOR2 (N11753, N11744, N3138);
not NOT1 (N11754, N11749);
not NOT1 (N11755, N11752);
nand NAND2 (N11756, N11745, N3230);
buf BUF1 (N11757, N11753);
buf BUF1 (N11758, N11725);
buf BUF1 (N11759, N11757);
xor XOR2 (N11760, N11748, N6099);
nand NAND2 (N11761, N11756, N11631);
xor XOR2 (N11762, N11760, N1308);
and AND2 (N11763, N11755, N9659);
xor XOR2 (N11764, N11759, N9099);
or OR2 (N11765, N11763, N710);
not NOT1 (N11766, N11746);
nand NAND3 (N11767, N11761, N9663, N9591);
and AND2 (N11768, N11765, N3797);
nor NOR3 (N11769, N11742, N3992, N342);
buf BUF1 (N11770, N11768);
or OR4 (N11771, N11766, N7444, N11628, N11263);
xor XOR2 (N11772, N11754, N9170);
buf BUF1 (N11773, N11764);
and AND2 (N11774, N11758, N10655);
buf BUF1 (N11775, N11774);
or OR4 (N11776, N11741, N7597, N2662, N6741);
and AND4 (N11777, N11775, N27, N3903, N3944);
or OR4 (N11778, N11772, N11342, N3710, N765);
and AND2 (N11779, N11770, N1689);
or OR4 (N11780, N11771, N7426, N676, N8303);
not NOT1 (N11781, N11780);
nor NOR3 (N11782, N11777, N5193, N7642);
or OR3 (N11783, N11779, N6241, N8448);
and AND3 (N11784, N11773, N10968, N4001);
nand NAND3 (N11785, N11781, N8147, N8256);
xor XOR2 (N11786, N11769, N11120);
xor XOR2 (N11787, N11785, N10753);
or OR3 (N11788, N11783, N6505, N1519);
nand NAND4 (N11789, N11788, N7341, N4638, N4789);
nor NOR2 (N11790, N11778, N4375);
not NOT1 (N11791, N11784);
nor NOR2 (N11792, N11791, N10829);
not NOT1 (N11793, N11792);
nor NOR3 (N11794, N11776, N512, N253);
nor NOR3 (N11795, N11794, N345, N319);
buf BUF1 (N11796, N11782);
or OR3 (N11797, N11793, N10137, N8931);
buf BUF1 (N11798, N11786);
buf BUF1 (N11799, N11796);
xor XOR2 (N11800, N11799, N8597);
not NOT1 (N11801, N11789);
nor NOR3 (N11802, N11800, N5853, N1454);
buf BUF1 (N11803, N11787);
nand NAND3 (N11804, N11751, N1675, N6243);
nand NAND4 (N11805, N11767, N4200, N10493, N6051);
nor NOR3 (N11806, N11804, N5857, N1902);
nor NOR3 (N11807, N11801, N10066, N11301);
not NOT1 (N11808, N11798);
nor NOR3 (N11809, N11762, N9922, N2089);
nand NAND2 (N11810, N11806, N3568);
or OR3 (N11811, N11809, N11081, N2272);
xor XOR2 (N11812, N11810, N3720);
nand NAND3 (N11813, N11808, N2583, N8771);
nor NOR2 (N11814, N11813, N7881);
xor XOR2 (N11815, N11807, N9160);
nor NOR4 (N11816, N11790, N2529, N6905, N8740);
nor NOR2 (N11817, N11816, N10738);
or OR2 (N11818, N11795, N8220);
nand NAND2 (N11819, N11814, N6482);
xor XOR2 (N11820, N11811, N625);
not NOT1 (N11821, N11803);
and AND4 (N11822, N11819, N5049, N7941, N2339);
not NOT1 (N11823, N11812);
nand NAND3 (N11824, N11817, N8418, N9465);
nand NAND4 (N11825, N11805, N6126, N2843, N4549);
nand NAND2 (N11826, N11818, N4230);
or OR4 (N11827, N11824, N7737, N6524, N5227);
and AND2 (N11828, N11802, N402);
nand NAND4 (N11829, N11825, N1329, N8206, N10445);
or OR3 (N11830, N11820, N5388, N11459);
buf BUF1 (N11831, N11823);
nor NOR3 (N11832, N11797, N5546, N4952);
or OR2 (N11833, N11832, N92);
xor XOR2 (N11834, N11831, N4649);
or OR2 (N11835, N11827, N7465);
not NOT1 (N11836, N11833);
not NOT1 (N11837, N11836);
or OR2 (N11838, N11828, N902);
buf BUF1 (N11839, N11838);
not NOT1 (N11840, N11835);
or OR3 (N11841, N11829, N10388, N537);
or OR2 (N11842, N11839, N10012);
nand NAND2 (N11843, N11815, N11156);
nand NAND2 (N11844, N11837, N6865);
buf BUF1 (N11845, N11834);
nor NOR4 (N11846, N11845, N10438, N10288, N8632);
nand NAND2 (N11847, N11840, N2910);
nand NAND4 (N11848, N11846, N4874, N6902, N2338);
or OR4 (N11849, N11847, N4013, N4967, N8230);
nor NOR2 (N11850, N11821, N8075);
nand NAND3 (N11851, N11844, N5978, N3045);
nor NOR3 (N11852, N11841, N4776, N1664);
xor XOR2 (N11853, N11848, N6915);
xor XOR2 (N11854, N11822, N9531);
xor XOR2 (N11855, N11850, N1015);
or OR2 (N11856, N11855, N2868);
not NOT1 (N11857, N11852);
or OR3 (N11858, N11851, N10728, N11359);
not NOT1 (N11859, N11854);
and AND4 (N11860, N11843, N9411, N1409, N7445);
buf BUF1 (N11861, N11849);
or OR2 (N11862, N11856, N11654);
not NOT1 (N11863, N11859);
xor XOR2 (N11864, N11861, N5340);
not NOT1 (N11865, N11863);
nor NOR2 (N11866, N11864, N3952);
buf BUF1 (N11867, N11853);
or OR2 (N11868, N11865, N9699);
nor NOR4 (N11869, N11860, N627, N6867, N7755);
or OR4 (N11870, N11862, N3833, N8091, N8833);
xor XOR2 (N11871, N11869, N210);
or OR4 (N11872, N11866, N7394, N11105, N6383);
and AND4 (N11873, N11871, N7226, N4298, N7030);
and AND2 (N11874, N11870, N917);
and AND4 (N11875, N11867, N9551, N7710, N9106);
xor XOR2 (N11876, N11875, N11214);
or OR3 (N11877, N11842, N11756, N3434);
buf BUF1 (N11878, N11872);
xor XOR2 (N11879, N11874, N8808);
and AND4 (N11880, N11857, N6843, N2860, N6047);
buf BUF1 (N11881, N11830);
and AND2 (N11882, N11881, N1442);
xor XOR2 (N11883, N11879, N3955);
nor NOR3 (N11884, N11880, N1287, N10632);
and AND2 (N11885, N11858, N104);
buf BUF1 (N11886, N11884);
and AND3 (N11887, N11885, N1474, N8056);
xor XOR2 (N11888, N11886, N2952);
or OR2 (N11889, N11878, N11514);
and AND2 (N11890, N11887, N8435);
buf BUF1 (N11891, N11826);
and AND4 (N11892, N11889, N11777, N2393, N5394);
xor XOR2 (N11893, N11877, N1404);
buf BUF1 (N11894, N11892);
buf BUF1 (N11895, N11891);
xor XOR2 (N11896, N11883, N2363);
xor XOR2 (N11897, N11895, N9597);
and AND3 (N11898, N11896, N10484, N6989);
or OR2 (N11899, N11873, N5247);
or OR2 (N11900, N11898, N516);
and AND3 (N11901, N11868, N3062, N7205);
buf BUF1 (N11902, N11882);
not NOT1 (N11903, N11899);
buf BUF1 (N11904, N11890);
nand NAND4 (N11905, N11888, N8226, N9721, N1219);
nor NOR4 (N11906, N11901, N279, N3616, N232);
and AND4 (N11907, N11897, N11149, N9953, N1044);
nand NAND2 (N11908, N11894, N9989);
and AND4 (N11909, N11876, N349, N10965, N10229);
xor XOR2 (N11910, N11902, N3650);
nor NOR3 (N11911, N11900, N7965, N9909);
or OR3 (N11912, N11904, N11639, N6295);
not NOT1 (N11913, N11909);
xor XOR2 (N11914, N11911, N11517);
nor NOR4 (N11915, N11914, N1478, N2832, N6462);
buf BUF1 (N11916, N11913);
nor NOR4 (N11917, N11912, N10116, N4134, N3782);
not NOT1 (N11918, N11906);
and AND4 (N11919, N11916, N7220, N4405, N6437);
nand NAND4 (N11920, N11918, N2390, N6513, N76);
nor NOR3 (N11921, N11893, N9642, N8468);
xor XOR2 (N11922, N11907, N9458);
xor XOR2 (N11923, N11908, N6523);
nand NAND3 (N11924, N11910, N5388, N5464);
nor NOR4 (N11925, N11903, N4558, N1559, N7229);
buf BUF1 (N11926, N11917);
or OR2 (N11927, N11905, N4926);
nand NAND2 (N11928, N11927, N7824);
and AND3 (N11929, N11919, N7279, N44);
buf BUF1 (N11930, N11921);
buf BUF1 (N11931, N11920);
nor NOR2 (N11932, N11924, N8825);
xor XOR2 (N11933, N11923, N11879);
xor XOR2 (N11934, N11932, N3309);
nor NOR2 (N11935, N11931, N10920);
xor XOR2 (N11936, N11929, N4307);
nand NAND2 (N11937, N11915, N4733);
nand NAND4 (N11938, N11937, N161, N6548, N2310);
and AND3 (N11939, N11934, N8821, N7575);
nor NOR3 (N11940, N11938, N763, N4334);
and AND2 (N11941, N11930, N4560);
and AND4 (N11942, N11925, N2655, N9957, N4300);
nand NAND4 (N11943, N11936, N1242, N11318, N464);
and AND3 (N11944, N11943, N8206, N3356);
nand NAND2 (N11945, N11922, N10795);
buf BUF1 (N11946, N11935);
nand NAND4 (N11947, N11944, N2515, N10745, N5587);
or OR3 (N11948, N11946, N9221, N11041);
buf BUF1 (N11949, N11933);
nand NAND2 (N11950, N11947, N7943);
and AND3 (N11951, N11942, N10748, N9728);
buf BUF1 (N11952, N11950);
nand NAND3 (N11953, N11948, N4756, N10636);
nand NAND3 (N11954, N11941, N4398, N9295);
nor NOR4 (N11955, N11926, N4231, N5152, N987);
buf BUF1 (N11956, N11954);
nand NAND3 (N11957, N11928, N808, N10009);
not NOT1 (N11958, N11939);
nand NAND2 (N11959, N11949, N2452);
xor XOR2 (N11960, N11951, N10419);
buf BUF1 (N11961, N11959);
and AND4 (N11962, N11961, N10568, N11103, N6454);
nor NOR4 (N11963, N11953, N11294, N8202, N5830);
xor XOR2 (N11964, N11962, N6137);
buf BUF1 (N11965, N11945);
and AND4 (N11966, N11958, N4733, N10009, N11942);
and AND3 (N11967, N11940, N7128, N5108);
and AND4 (N11968, N11960, N10528, N3784, N4732);
buf BUF1 (N11969, N11963);
xor XOR2 (N11970, N11957, N4649);
xor XOR2 (N11971, N11966, N6432);
nand NAND3 (N11972, N11971, N2261, N5697);
nand NAND4 (N11973, N11967, N1308, N2400, N2562);
buf BUF1 (N11974, N11964);
nand NAND3 (N11975, N11973, N3775, N8045);
xor XOR2 (N11976, N11972, N614);
not NOT1 (N11977, N11956);
nor NOR2 (N11978, N11977, N10759);
buf BUF1 (N11979, N11978);
not NOT1 (N11980, N11965);
and AND3 (N11981, N11955, N7258, N4795);
buf BUF1 (N11982, N11974);
not NOT1 (N11983, N11970);
not NOT1 (N11984, N11981);
not NOT1 (N11985, N11982);
not NOT1 (N11986, N11952);
and AND4 (N11987, N11975, N1402, N8999, N8667);
or OR4 (N11988, N11986, N3912, N2495, N2740);
and AND4 (N11989, N11980, N2211, N4206, N2972);
nor NOR4 (N11990, N11988, N3086, N5715, N1919);
xor XOR2 (N11991, N11976, N6300);
buf BUF1 (N11992, N11983);
or OR2 (N11993, N11969, N4180);
buf BUF1 (N11994, N11990);
not NOT1 (N11995, N11987);
and AND4 (N11996, N11993, N11829, N2105, N5140);
not NOT1 (N11997, N11979);
nor NOR4 (N11998, N11984, N4288, N2759, N4063);
nand NAND4 (N11999, N11985, N5991, N146, N8813);
or OR3 (N12000, N11994, N4660, N8169);
nor NOR2 (N12001, N11989, N3918);
xor XOR2 (N12002, N12001, N5960);
not NOT1 (N12003, N12002);
nor NOR2 (N12004, N11997, N5516);
or OR4 (N12005, N11996, N11110, N1656, N9331);
or OR3 (N12006, N11992, N7021, N10846);
buf BUF1 (N12007, N11995);
xor XOR2 (N12008, N12000, N4436);
nor NOR3 (N12009, N11999, N5877, N5901);
nand NAND2 (N12010, N12004, N6146);
or OR3 (N12011, N11968, N1716, N187);
nand NAND4 (N12012, N12008, N4665, N10127, N9692);
buf BUF1 (N12013, N12010);
nor NOR3 (N12014, N12006, N10979, N10760);
not NOT1 (N12015, N12013);
nand NAND2 (N12016, N12014, N4942);
not NOT1 (N12017, N12005);
xor XOR2 (N12018, N12003, N8227);
xor XOR2 (N12019, N12012, N3667);
not NOT1 (N12020, N12019);
buf BUF1 (N12021, N12007);
buf BUF1 (N12022, N11998);
or OR4 (N12023, N12016, N7252, N4892, N2411);
not NOT1 (N12024, N12011);
nor NOR2 (N12025, N12009, N1386);
not NOT1 (N12026, N12017);
xor XOR2 (N12027, N12020, N2445);
nor NOR2 (N12028, N12026, N5204);
or OR3 (N12029, N12022, N995, N4305);
nor NOR3 (N12030, N12021, N4970, N5394);
buf BUF1 (N12031, N12028);
not NOT1 (N12032, N12015);
not NOT1 (N12033, N12025);
nand NAND2 (N12034, N12023, N5366);
buf BUF1 (N12035, N12034);
not NOT1 (N12036, N12024);
not NOT1 (N12037, N12027);
buf BUF1 (N12038, N12032);
xor XOR2 (N12039, N12036, N6410);
not NOT1 (N12040, N12039);
and AND2 (N12041, N12018, N7807);
and AND2 (N12042, N12038, N1654);
nand NAND3 (N12043, N12042, N5777, N9278);
nand NAND3 (N12044, N12029, N8810, N11560);
not NOT1 (N12045, N11991);
xor XOR2 (N12046, N12031, N11026);
or OR2 (N12047, N12035, N10924);
buf BUF1 (N12048, N12030);
not NOT1 (N12049, N12037);
nand NAND2 (N12050, N12040, N4429);
or OR4 (N12051, N12041, N4742, N1851, N669);
nand NAND2 (N12052, N12051, N3542);
nor NOR4 (N12053, N12050, N8519, N4398, N3996);
xor XOR2 (N12054, N12049, N1869);
and AND3 (N12055, N12048, N4965, N3383);
or OR2 (N12056, N12055, N8149);
or OR2 (N12057, N12046, N4610);
xor XOR2 (N12058, N12033, N1864);
nand NAND4 (N12059, N12053, N4988, N3229, N9277);
not NOT1 (N12060, N12043);
buf BUF1 (N12061, N12052);
xor XOR2 (N12062, N12044, N6930);
nor NOR2 (N12063, N12061, N5571);
xor XOR2 (N12064, N12060, N6869);
or OR3 (N12065, N12062, N3735, N9159);
or OR3 (N12066, N12063, N6823, N6391);
nor NOR3 (N12067, N12058, N4509, N1987);
nand NAND4 (N12068, N12066, N3676, N1042, N10272);
not NOT1 (N12069, N12056);
xor XOR2 (N12070, N12054, N5809);
nor NOR3 (N12071, N12067, N6212, N1973);
nand NAND4 (N12072, N12059, N1909, N4866, N5201);
not NOT1 (N12073, N12057);
or OR4 (N12074, N12069, N3838, N9844, N999);
buf BUF1 (N12075, N12047);
not NOT1 (N12076, N12045);
nand NAND4 (N12077, N12070, N5993, N3653, N2424);
xor XOR2 (N12078, N12072, N7147);
xor XOR2 (N12079, N12071, N9061);
buf BUF1 (N12080, N12077);
nand NAND3 (N12081, N12079, N221, N3879);
xor XOR2 (N12082, N12080, N2987);
or OR2 (N12083, N12074, N10570);
nor NOR4 (N12084, N12073, N3996, N5445, N11492);
buf BUF1 (N12085, N12064);
nor NOR4 (N12086, N12065, N272, N6611, N10872);
nand NAND3 (N12087, N12084, N7094, N1289);
not NOT1 (N12088, N12083);
not NOT1 (N12089, N12085);
nand NAND3 (N12090, N12082, N6078, N7679);
nand NAND2 (N12091, N12078, N9822);
nand NAND3 (N12092, N12076, N7077, N4086);
nand NAND2 (N12093, N12092, N1047);
xor XOR2 (N12094, N12090, N11329);
nor NOR3 (N12095, N12075, N509, N11253);
buf BUF1 (N12096, N12081);
and AND2 (N12097, N12091, N12004);
xor XOR2 (N12098, N12097, N6726);
nor NOR4 (N12099, N12096, N4560, N253, N6371);
xor XOR2 (N12100, N12099, N230);
xor XOR2 (N12101, N12100, N3642);
not NOT1 (N12102, N12086);
or OR2 (N12103, N12068, N6276);
or OR3 (N12104, N12098, N7454, N3504);
nor NOR4 (N12105, N12103, N628, N6139, N2468);
buf BUF1 (N12106, N12095);
not NOT1 (N12107, N12106);
xor XOR2 (N12108, N12088, N11975);
buf BUF1 (N12109, N12104);
xor XOR2 (N12110, N12108, N8913);
buf BUF1 (N12111, N12101);
or OR4 (N12112, N12105, N11003, N2315, N10215);
not NOT1 (N12113, N12089);
and AND4 (N12114, N12112, N9178, N6419, N3243);
xor XOR2 (N12115, N12109, N10035);
and AND3 (N12116, N12110, N7341, N9313);
nand NAND2 (N12117, N12094, N9076);
nor NOR2 (N12118, N12114, N10725);
nor NOR4 (N12119, N12093, N1527, N7296, N10927);
nand NAND2 (N12120, N12117, N12019);
not NOT1 (N12121, N12111);
and AND2 (N12122, N12115, N6742);
nand NAND4 (N12123, N12107, N8960, N1659, N7545);
buf BUF1 (N12124, N12122);
and AND2 (N12125, N12119, N6428);
not NOT1 (N12126, N12118);
or OR4 (N12127, N12087, N5978, N5519, N6413);
xor XOR2 (N12128, N12124, N5635);
not NOT1 (N12129, N12116);
and AND4 (N12130, N12129, N4859, N4897, N1213);
or OR3 (N12131, N12102, N1928, N7418);
nor NOR2 (N12132, N12131, N9504);
buf BUF1 (N12133, N12123);
nor NOR2 (N12134, N12130, N7516);
nand NAND3 (N12135, N12125, N2443, N928);
or OR2 (N12136, N12133, N1786);
and AND4 (N12137, N12134, N6694, N2694, N9364);
not NOT1 (N12138, N12132);
and AND4 (N12139, N12136, N6220, N10759, N4563);
and AND4 (N12140, N12127, N11310, N9504, N9583);
xor XOR2 (N12141, N12121, N10728);
buf BUF1 (N12142, N12137);
nand NAND4 (N12143, N12120, N1850, N7384, N6543);
or OR4 (N12144, N12126, N2034, N961, N6176);
not NOT1 (N12145, N12135);
nand NAND4 (N12146, N12128, N6312, N8927, N7068);
not NOT1 (N12147, N12142);
buf BUF1 (N12148, N12146);
nor NOR2 (N12149, N12138, N3699);
not NOT1 (N12150, N12148);
not NOT1 (N12151, N12139);
not NOT1 (N12152, N12113);
nand NAND2 (N12153, N12141, N9143);
not NOT1 (N12154, N12153);
not NOT1 (N12155, N12154);
buf BUF1 (N12156, N12140);
buf BUF1 (N12157, N12152);
xor XOR2 (N12158, N12149, N12115);
not NOT1 (N12159, N12150);
not NOT1 (N12160, N12155);
not NOT1 (N12161, N12145);
nand NAND3 (N12162, N12157, N2202, N11172);
xor XOR2 (N12163, N12144, N7418);
not NOT1 (N12164, N12143);
buf BUF1 (N12165, N12156);
nor NOR2 (N12166, N12160, N907);
nor NOR3 (N12167, N12159, N8912, N1265);
nand NAND4 (N12168, N12164, N3662, N11720, N8538);
not NOT1 (N12169, N12162);
and AND3 (N12170, N12168, N6568, N6436);
xor XOR2 (N12171, N12167, N10167);
not NOT1 (N12172, N12165);
xor XOR2 (N12173, N12151, N8149);
and AND3 (N12174, N12170, N8525, N10916);
or OR2 (N12175, N12169, N110);
nor NOR3 (N12176, N12158, N9695, N7555);
nor NOR2 (N12177, N12171, N6147);
or OR3 (N12178, N12175, N8018, N11085);
nor NOR2 (N12179, N12161, N6037);
nor NOR2 (N12180, N12166, N5992);
or OR2 (N12181, N12147, N1894);
buf BUF1 (N12182, N12180);
not NOT1 (N12183, N12174);
not NOT1 (N12184, N12172);
nor NOR4 (N12185, N12181, N1050, N6429, N3348);
buf BUF1 (N12186, N12183);
xor XOR2 (N12187, N12182, N11219);
buf BUF1 (N12188, N12184);
not NOT1 (N12189, N12186);
buf BUF1 (N12190, N12185);
or OR4 (N12191, N12177, N2070, N3716, N9455);
and AND2 (N12192, N12191, N2581);
not NOT1 (N12193, N12188);
or OR4 (N12194, N12163, N3586, N10869, N11515);
nor NOR4 (N12195, N12187, N8200, N6681, N725);
xor XOR2 (N12196, N12190, N8917);
not NOT1 (N12197, N12178);
nor NOR3 (N12198, N12189, N1999, N3808);
and AND4 (N12199, N12176, N4742, N6060, N9462);
nand NAND2 (N12200, N12193, N1248);
xor XOR2 (N12201, N12192, N504);
buf BUF1 (N12202, N12179);
xor XOR2 (N12203, N12197, N9623);
and AND4 (N12204, N12194, N7764, N10324, N11214);
nand NAND3 (N12205, N12198, N5863, N2607);
and AND2 (N12206, N12201, N10994);
xor XOR2 (N12207, N12173, N11628);
nor NOR2 (N12208, N12202, N7015);
nor NOR3 (N12209, N12207, N6443, N3408);
nand NAND2 (N12210, N12206, N10409);
buf BUF1 (N12211, N12210);
not NOT1 (N12212, N12195);
xor XOR2 (N12213, N12208, N9832);
nand NAND3 (N12214, N12204, N4956, N4350);
xor XOR2 (N12215, N12196, N10102);
xor XOR2 (N12216, N12215, N3997);
not NOT1 (N12217, N12209);
not NOT1 (N12218, N12205);
or OR2 (N12219, N12218, N10540);
or OR2 (N12220, N12211, N7541);
nand NAND3 (N12221, N12220, N6434, N7254);
or OR2 (N12222, N12213, N1513);
xor XOR2 (N12223, N12200, N6031);
and AND3 (N12224, N12214, N4234, N5289);
xor XOR2 (N12225, N12219, N3293);
not NOT1 (N12226, N12216);
nor NOR3 (N12227, N12203, N2207, N11334);
xor XOR2 (N12228, N12225, N5164);
xor XOR2 (N12229, N12226, N5011);
nor NOR2 (N12230, N12221, N9345);
nand NAND3 (N12231, N12230, N7578, N2747);
nand NAND3 (N12232, N12229, N5972, N7779);
buf BUF1 (N12233, N12227);
or OR2 (N12234, N12228, N99);
nand NAND2 (N12235, N12223, N4991);
and AND4 (N12236, N12222, N11724, N8340, N6489);
nand NAND4 (N12237, N12233, N11685, N3548, N8206);
or OR4 (N12238, N12236, N3082, N11964, N6619);
and AND2 (N12239, N12232, N6440);
not NOT1 (N12240, N12231);
buf BUF1 (N12241, N12239);
not NOT1 (N12242, N12199);
or OR2 (N12243, N12242, N1666);
nand NAND4 (N12244, N12217, N11944, N4144, N11697);
or OR3 (N12245, N12244, N9474, N11526);
buf BUF1 (N12246, N12235);
or OR3 (N12247, N12234, N8252, N10426);
nand NAND4 (N12248, N12246, N6803, N8312, N12099);
not NOT1 (N12249, N12241);
and AND2 (N12250, N12224, N986);
nor NOR3 (N12251, N12245, N669, N1223);
xor XOR2 (N12252, N12249, N7916);
buf BUF1 (N12253, N12250);
nand NAND3 (N12254, N12212, N9567, N11747);
and AND3 (N12255, N12253, N10346, N73);
nand NAND4 (N12256, N12255, N7524, N1412, N6336);
buf BUF1 (N12257, N12254);
and AND4 (N12258, N12237, N11203, N9530, N5265);
xor XOR2 (N12259, N12251, N7509);
xor XOR2 (N12260, N12252, N11482);
not NOT1 (N12261, N12256);
or OR3 (N12262, N12258, N2621, N7141);
not NOT1 (N12263, N12259);
not NOT1 (N12264, N12257);
not NOT1 (N12265, N12243);
or OR4 (N12266, N12248, N10589, N10644, N7686);
or OR2 (N12267, N12264, N3981);
nand NAND2 (N12268, N12265, N11567);
nand NAND4 (N12269, N12266, N9090, N8491, N3163);
nand NAND3 (N12270, N12261, N1880, N10823);
or OR4 (N12271, N12267, N10135, N847, N939);
not NOT1 (N12272, N12260);
or OR2 (N12273, N12263, N467);
not NOT1 (N12274, N12272);
nor NOR3 (N12275, N12273, N1513, N2343);
and AND2 (N12276, N12271, N4017);
nor NOR2 (N12277, N12276, N3684);
or OR4 (N12278, N12269, N2861, N9521, N4732);
and AND2 (N12279, N12275, N10506);
nor NOR2 (N12280, N12238, N657);
not NOT1 (N12281, N12278);
nand NAND2 (N12282, N12268, N7908);
not NOT1 (N12283, N12247);
nor NOR2 (N12284, N12270, N8161);
or OR2 (N12285, N12281, N5396);
buf BUF1 (N12286, N12284);
or OR3 (N12287, N12280, N1707, N8314);
nor NOR4 (N12288, N12282, N1477, N8678, N1765);
xor XOR2 (N12289, N12287, N6079);
not NOT1 (N12290, N12279);
not NOT1 (N12291, N12285);
not NOT1 (N12292, N12290);
nor NOR4 (N12293, N12283, N8892, N9186, N1641);
not NOT1 (N12294, N12288);
and AND3 (N12295, N12291, N10674, N1380);
and AND4 (N12296, N12294, N4676, N9667, N11830);
buf BUF1 (N12297, N12293);
or OR3 (N12298, N12297, N4607, N11913);
or OR3 (N12299, N12295, N7607, N8158);
nand NAND2 (N12300, N12286, N12207);
nand NAND3 (N12301, N12299, N17, N4111);
not NOT1 (N12302, N12298);
buf BUF1 (N12303, N12302);
nor NOR2 (N12304, N12301, N3608);
xor XOR2 (N12305, N12300, N2394);
and AND2 (N12306, N12296, N460);
buf BUF1 (N12307, N12303);
or OR3 (N12308, N12307, N7750, N9990);
nor NOR3 (N12309, N12277, N12032, N10038);
nand NAND3 (N12310, N12240, N11431, N3794);
nand NAND2 (N12311, N12310, N8187);
and AND3 (N12312, N12311, N9340, N2806);
xor XOR2 (N12313, N12305, N546);
buf BUF1 (N12314, N12313);
and AND4 (N12315, N12274, N3409, N427, N7921);
and AND4 (N12316, N12292, N6003, N4581, N2975);
xor XOR2 (N12317, N12306, N703);
and AND4 (N12318, N12308, N638, N7348, N2835);
nand NAND3 (N12319, N12318, N4604, N6543);
buf BUF1 (N12320, N12304);
not NOT1 (N12321, N12312);
nor NOR3 (N12322, N12315, N12043, N3836);
and AND2 (N12323, N12320, N10794);
nor NOR2 (N12324, N12316, N6677);
and AND2 (N12325, N12317, N12264);
buf BUF1 (N12326, N12262);
and AND3 (N12327, N12309, N4913, N3618);
and AND2 (N12328, N12289, N12025);
xor XOR2 (N12329, N12326, N12200);
xor XOR2 (N12330, N12325, N9238);
nor NOR3 (N12331, N12323, N2540, N5009);
nor NOR2 (N12332, N12321, N12215);
and AND2 (N12333, N12332, N2780);
nand NAND2 (N12334, N12330, N9124);
buf BUF1 (N12335, N12319);
not NOT1 (N12336, N12334);
and AND4 (N12337, N12329, N863, N9221, N8779);
xor XOR2 (N12338, N12314, N6324);
xor XOR2 (N12339, N12335, N11614);
nand NAND4 (N12340, N12337, N7972, N243, N6476);
nor NOR3 (N12341, N12328, N6271, N7883);
nor NOR3 (N12342, N12322, N7362, N6283);
and AND4 (N12343, N12340, N10214, N1209, N9446);
nor NOR4 (N12344, N12327, N12000, N6829, N10879);
and AND3 (N12345, N12341, N11156, N9055);
nor NOR3 (N12346, N12324, N6571, N9896);
and AND3 (N12347, N12333, N5004, N9413);
not NOT1 (N12348, N12346);
nand NAND3 (N12349, N12343, N5797, N4103);
not NOT1 (N12350, N12338);
or OR3 (N12351, N12342, N228, N631);
or OR2 (N12352, N12349, N7490);
not NOT1 (N12353, N12331);
xor XOR2 (N12354, N12348, N5098);
xor XOR2 (N12355, N12344, N6667);
nor NOR2 (N12356, N12354, N2098);
and AND4 (N12357, N12347, N3143, N2319, N5234);
nand NAND4 (N12358, N12351, N1433, N2163, N3547);
buf BUF1 (N12359, N12339);
xor XOR2 (N12360, N12356, N9456);
and AND2 (N12361, N12358, N6603);
nand NAND4 (N12362, N12336, N2303, N580, N8287);
or OR2 (N12363, N12352, N5527);
not NOT1 (N12364, N12362);
and AND2 (N12365, N12360, N9574);
nand NAND2 (N12366, N12364, N2134);
not NOT1 (N12367, N12363);
buf BUF1 (N12368, N12367);
and AND3 (N12369, N12345, N9159, N9278);
and AND4 (N12370, N12368, N1880, N2254, N11399);
xor XOR2 (N12371, N12359, N276);
and AND4 (N12372, N12357, N10053, N6162, N2337);
not NOT1 (N12373, N12366);
xor XOR2 (N12374, N12350, N7241);
buf BUF1 (N12375, N12372);
xor XOR2 (N12376, N12370, N3262);
or OR3 (N12377, N12374, N5597, N3689);
and AND3 (N12378, N12377, N10071, N1613);
nor NOR4 (N12379, N12353, N6805, N7182, N7718);
nand NAND2 (N12380, N12369, N7869);
and AND4 (N12381, N12355, N3800, N5344, N5623);
or OR2 (N12382, N12373, N9206);
or OR4 (N12383, N12381, N10696, N5516, N1960);
nand NAND4 (N12384, N12378, N8876, N5603, N3331);
nand NAND2 (N12385, N12379, N8277);
nand NAND3 (N12386, N12380, N9222, N2603);
and AND2 (N12387, N12375, N2140);
buf BUF1 (N12388, N12365);
and AND3 (N12389, N12361, N3036, N9898);
not NOT1 (N12390, N12384);
or OR2 (N12391, N12382, N7584);
nand NAND2 (N12392, N12387, N10741);
xor XOR2 (N12393, N12388, N1102);
nor NOR3 (N12394, N12392, N5079, N8466);
buf BUF1 (N12395, N12394);
buf BUF1 (N12396, N12383);
buf BUF1 (N12397, N12376);
not NOT1 (N12398, N12393);
and AND4 (N12399, N12386, N5866, N5699, N3316);
xor XOR2 (N12400, N12398, N9419);
nor NOR2 (N12401, N12397, N9580);
or OR2 (N12402, N12399, N10750);
nand NAND2 (N12403, N12401, N4053);
buf BUF1 (N12404, N12371);
xor XOR2 (N12405, N12400, N11544);
nand NAND4 (N12406, N12404, N9483, N11134, N12286);
and AND3 (N12407, N12406, N7874, N222);
xor XOR2 (N12408, N12407, N5352);
not NOT1 (N12409, N12391);
buf BUF1 (N12410, N12395);
not NOT1 (N12411, N12405);
not NOT1 (N12412, N12402);
not NOT1 (N12413, N12390);
buf BUF1 (N12414, N12396);
nor NOR2 (N12415, N12408, N8193);
not NOT1 (N12416, N12413);
not NOT1 (N12417, N12409);
xor XOR2 (N12418, N12417, N10992);
nand NAND4 (N12419, N12385, N1225, N5196, N8839);
xor XOR2 (N12420, N12415, N9074);
nand NAND2 (N12421, N12411, N2456);
xor XOR2 (N12422, N12416, N10501);
nand NAND4 (N12423, N12389, N1719, N7069, N618);
and AND3 (N12424, N12419, N1527, N6199);
buf BUF1 (N12425, N12412);
xor XOR2 (N12426, N12421, N5325);
not NOT1 (N12427, N12403);
or OR4 (N12428, N12422, N343, N3947, N9900);
or OR2 (N12429, N12423, N9253);
xor XOR2 (N12430, N12420, N2095);
buf BUF1 (N12431, N12425);
xor XOR2 (N12432, N12418, N10581);
or OR3 (N12433, N12410, N2880, N7538);
and AND3 (N12434, N12432, N4689, N2809);
and AND3 (N12435, N12430, N768, N2047);
nand NAND4 (N12436, N12428, N9587, N7339, N448);
xor XOR2 (N12437, N12436, N10875);
xor XOR2 (N12438, N12424, N4721);
xor XOR2 (N12439, N12426, N12245);
xor XOR2 (N12440, N12434, N6841);
or OR4 (N12441, N12439, N1451, N9290, N7387);
nor NOR2 (N12442, N12431, N10785);
nand NAND2 (N12443, N12440, N1368);
nand NAND3 (N12444, N12429, N9909, N5647);
buf BUF1 (N12445, N12437);
or OR2 (N12446, N12441, N7244);
buf BUF1 (N12447, N12443);
not NOT1 (N12448, N12444);
or OR3 (N12449, N12414, N1154, N1453);
xor XOR2 (N12450, N12445, N7020);
nor NOR2 (N12451, N12450, N7511);
nor NOR4 (N12452, N12448, N11733, N10730, N5668);
nand NAND3 (N12453, N12447, N7077, N9120);
xor XOR2 (N12454, N12442, N6606);
xor XOR2 (N12455, N12433, N8119);
not NOT1 (N12456, N12454);
xor XOR2 (N12457, N12427, N9490);
nand NAND3 (N12458, N12438, N4239, N11797);
or OR4 (N12459, N12455, N4123, N10115, N2265);
buf BUF1 (N12460, N12457);
buf BUF1 (N12461, N12451);
nand NAND4 (N12462, N12458, N11492, N7733, N12005);
xor XOR2 (N12463, N12460, N2380);
and AND3 (N12464, N12452, N9796, N6276);
nor NOR3 (N12465, N12446, N5849, N10828);
xor XOR2 (N12466, N12461, N8154);
buf BUF1 (N12467, N12462);
nand NAND4 (N12468, N12464, N12019, N9503, N11425);
xor XOR2 (N12469, N12463, N12269);
and AND3 (N12470, N12467, N10098, N1622);
buf BUF1 (N12471, N12449);
buf BUF1 (N12472, N12456);
nor NOR2 (N12473, N12466, N11015);
not NOT1 (N12474, N12469);
not NOT1 (N12475, N12470);
and AND3 (N12476, N12435, N6899, N965);
buf BUF1 (N12477, N12473);
nor NOR2 (N12478, N12471, N10153);
or OR2 (N12479, N12476, N11395);
nand NAND4 (N12480, N12465, N8251, N6557, N8771);
buf BUF1 (N12481, N12468);
or OR4 (N12482, N12459, N10439, N3926, N2554);
not NOT1 (N12483, N12479);
xor XOR2 (N12484, N12480, N1566);
and AND3 (N12485, N12453, N1607, N9129);
xor XOR2 (N12486, N12484, N10259);
nand NAND3 (N12487, N12485, N2662, N6841);
nand NAND4 (N12488, N12481, N5538, N962, N3275);
or OR3 (N12489, N12482, N8417, N7903);
or OR4 (N12490, N12489, N11069, N12111, N7422);
nand NAND3 (N12491, N12486, N2439, N12228);
nand NAND4 (N12492, N12483, N11358, N11020, N3636);
nor NOR2 (N12493, N12490, N7213);
nand NAND2 (N12494, N12472, N10722);
nor NOR4 (N12495, N12492, N9900, N12455, N652);
nand NAND3 (N12496, N12495, N6293, N5737);
xor XOR2 (N12497, N12496, N10786);
or OR4 (N12498, N12497, N10910, N7734, N1357);
xor XOR2 (N12499, N12498, N2389);
not NOT1 (N12500, N12488);
buf BUF1 (N12501, N12478);
and AND2 (N12502, N12494, N10066);
or OR3 (N12503, N12474, N4574, N10881);
nor NOR4 (N12504, N12503, N1451, N6347, N9957);
nor NOR3 (N12505, N12491, N4320, N5457);
xor XOR2 (N12506, N12475, N5283);
nand NAND2 (N12507, N12502, N4811);
nand NAND2 (N12508, N12499, N11507);
or OR3 (N12509, N12508, N5654, N8612);
xor XOR2 (N12510, N12505, N4470);
xor XOR2 (N12511, N12510, N5604);
not NOT1 (N12512, N12487);
nor NOR4 (N12513, N12493, N11896, N5149, N1674);
xor XOR2 (N12514, N12504, N6910);
nor NOR2 (N12515, N12514, N11588);
not NOT1 (N12516, N12507);
buf BUF1 (N12517, N12477);
nor NOR2 (N12518, N12512, N2853);
nand NAND3 (N12519, N12515, N6137, N9852);
nor NOR2 (N12520, N12511, N11978);
buf BUF1 (N12521, N12506);
or OR3 (N12522, N12513, N1320, N5645);
or OR4 (N12523, N12522, N3955, N2391, N11803);
xor XOR2 (N12524, N12501, N8024);
not NOT1 (N12525, N12520);
and AND4 (N12526, N12500, N6617, N65, N10715);
nand NAND3 (N12527, N12523, N2740, N5594);
or OR3 (N12528, N12509, N1668, N5);
xor XOR2 (N12529, N12525, N2735);
nor NOR2 (N12530, N12518, N6886);
or OR3 (N12531, N12517, N11562, N10201);
nand NAND4 (N12532, N12531, N2772, N85, N5796);
xor XOR2 (N12533, N12532, N6207);
nand NAND3 (N12534, N12527, N6287, N5388);
nand NAND4 (N12535, N12521, N851, N1833, N7947);
buf BUF1 (N12536, N12526);
xor XOR2 (N12537, N12534, N9649);
xor XOR2 (N12538, N12533, N8448);
nand NAND3 (N12539, N12516, N8739, N7225);
or OR2 (N12540, N12519, N10652);
nand NAND3 (N12541, N12535, N2071, N4181);
and AND3 (N12542, N12539, N9407, N10197);
not NOT1 (N12543, N12542);
xor XOR2 (N12544, N12536, N6296);
and AND3 (N12545, N12524, N5648, N8007);
and AND3 (N12546, N12544, N4077, N8578);
nor NOR3 (N12547, N12530, N11292, N5618);
nand NAND2 (N12548, N12537, N9093);
xor XOR2 (N12549, N12538, N5789);
xor XOR2 (N12550, N12529, N5536);
nand NAND3 (N12551, N12548, N8007, N2825);
or OR4 (N12552, N12550, N478, N10418, N10017);
nand NAND3 (N12553, N12546, N2680, N7295);
or OR2 (N12554, N12551, N2682);
buf BUF1 (N12555, N12545);
xor XOR2 (N12556, N12553, N1384);
nand NAND2 (N12557, N12543, N4449);
buf BUF1 (N12558, N12556);
or OR4 (N12559, N12557, N11258, N7011, N11030);
and AND4 (N12560, N12549, N1563, N8229, N6569);
buf BUF1 (N12561, N12541);
buf BUF1 (N12562, N12555);
and AND3 (N12563, N12558, N474, N8639);
nor NOR2 (N12564, N12528, N4433);
xor XOR2 (N12565, N12560, N5052);
or OR2 (N12566, N12559, N2430);
nand NAND2 (N12567, N12563, N5777);
nor NOR2 (N12568, N12554, N9543);
xor XOR2 (N12569, N12565, N11333);
buf BUF1 (N12570, N12540);
not NOT1 (N12571, N12567);
and AND4 (N12572, N12547, N4619, N1578, N10977);
and AND4 (N12573, N12566, N2569, N8039, N11847);
nor NOR2 (N12574, N12561, N1130);
buf BUF1 (N12575, N12569);
xor XOR2 (N12576, N12574, N6033);
buf BUF1 (N12577, N12576);
nand NAND4 (N12578, N12571, N6531, N11306, N3367);
xor XOR2 (N12579, N12578, N2815);
nor NOR4 (N12580, N12564, N10763, N5760, N8764);
not NOT1 (N12581, N12568);
and AND4 (N12582, N12570, N6819, N10215, N300);
not NOT1 (N12583, N12579);
or OR3 (N12584, N12575, N9095, N982);
xor XOR2 (N12585, N12584, N2225);
xor XOR2 (N12586, N12583, N9692);
nand NAND3 (N12587, N12586, N755, N3800);
buf BUF1 (N12588, N12572);
not NOT1 (N12589, N12581);
buf BUF1 (N12590, N12587);
or OR2 (N12591, N12589, N2531);
and AND4 (N12592, N12580, N4821, N10536, N11223);
nor NOR4 (N12593, N12573, N3407, N339, N7493);
xor XOR2 (N12594, N12552, N8994);
xor XOR2 (N12595, N12590, N8309);
nand NAND3 (N12596, N12577, N104, N9455);
or OR3 (N12597, N12594, N1757, N3613);
buf BUF1 (N12598, N12596);
nor NOR3 (N12599, N12595, N1065, N1415);
and AND2 (N12600, N12591, N6107);
buf BUF1 (N12601, N12598);
not NOT1 (N12602, N12601);
or OR3 (N12603, N12599, N9564, N175);
nand NAND4 (N12604, N12600, N9479, N8939, N2673);
nand NAND3 (N12605, N12604, N205, N4723);
nand NAND2 (N12606, N12605, N1761);
or OR2 (N12607, N12602, N10286);
or OR2 (N12608, N12607, N1622);
or OR2 (N12609, N12585, N7428);
or OR4 (N12610, N12609, N4423, N2010, N11891);
nor NOR4 (N12611, N12592, N9124, N2351, N12062);
or OR4 (N12612, N12593, N6351, N11471, N7567);
buf BUF1 (N12613, N12582);
or OR2 (N12614, N12606, N9595);
nor NOR4 (N12615, N12603, N8275, N9664, N7615);
nand NAND2 (N12616, N12597, N3188);
and AND4 (N12617, N12588, N5201, N6771, N3953);
or OR2 (N12618, N12562, N4499);
xor XOR2 (N12619, N12611, N3872);
and AND2 (N12620, N12613, N2500);
buf BUF1 (N12621, N12617);
not NOT1 (N12622, N12618);
not NOT1 (N12623, N12615);
or OR3 (N12624, N12614, N5882, N9725);
not NOT1 (N12625, N12620);
or OR4 (N12626, N12612, N4531, N10708, N9633);
xor XOR2 (N12627, N12619, N12521);
xor XOR2 (N12628, N12616, N804);
and AND3 (N12629, N12627, N9186, N11092);
xor XOR2 (N12630, N12623, N7761);
nor NOR3 (N12631, N12621, N12150, N10906);
buf BUF1 (N12632, N12610);
nor NOR2 (N12633, N12626, N5867);
and AND3 (N12634, N12629, N349, N8628);
not NOT1 (N12635, N12625);
or OR2 (N12636, N12632, N4912);
nand NAND2 (N12637, N12628, N3592);
or OR2 (N12638, N12636, N6990);
nor NOR3 (N12639, N12634, N4297, N4328);
nor NOR3 (N12640, N12637, N9705, N5432);
buf BUF1 (N12641, N12633);
and AND3 (N12642, N12631, N96, N3728);
xor XOR2 (N12643, N12630, N955);
nor NOR2 (N12644, N12608, N4137);
not NOT1 (N12645, N12642);
and AND4 (N12646, N12624, N4979, N7912, N5724);
xor XOR2 (N12647, N12635, N1784);
and AND3 (N12648, N12622, N1667, N12089);
buf BUF1 (N12649, N12641);
or OR4 (N12650, N12647, N8691, N2321, N5047);
nand NAND4 (N12651, N12650, N1470, N7876, N3211);
not NOT1 (N12652, N12645);
buf BUF1 (N12653, N12644);
buf BUF1 (N12654, N12640);
xor XOR2 (N12655, N12643, N7084);
nor NOR4 (N12656, N12652, N11081, N7242, N10029);
buf BUF1 (N12657, N12646);
xor XOR2 (N12658, N12651, N7183);
buf BUF1 (N12659, N12648);
nor NOR4 (N12660, N12658, N12504, N4716, N5386);
and AND3 (N12661, N12660, N11559, N12645);
or OR2 (N12662, N12659, N4281);
xor XOR2 (N12663, N12655, N7308);
xor XOR2 (N12664, N12649, N12228);
and AND2 (N12665, N12662, N2866);
or OR4 (N12666, N12661, N5324, N4543, N11039);
buf BUF1 (N12667, N12666);
not NOT1 (N12668, N12663);
or OR2 (N12669, N12667, N8509);
nor NOR4 (N12670, N12654, N7133, N11470, N11871);
nor NOR3 (N12671, N12665, N6485, N11313);
and AND4 (N12672, N12664, N448, N7831, N4847);
nand NAND4 (N12673, N12653, N6121, N9342, N87);
nor NOR3 (N12674, N12671, N6486, N2436);
and AND4 (N12675, N12656, N11179, N4745, N7917);
and AND2 (N12676, N12669, N2333);
buf BUF1 (N12677, N12673);
xor XOR2 (N12678, N12670, N6517);
and AND3 (N12679, N12676, N7345, N8656);
buf BUF1 (N12680, N12668);
or OR3 (N12681, N12638, N2485, N12530);
not NOT1 (N12682, N12657);
or OR2 (N12683, N12639, N5046);
xor XOR2 (N12684, N12675, N6989);
xor XOR2 (N12685, N12680, N9841);
not NOT1 (N12686, N12678);
nor NOR4 (N12687, N12683, N11525, N12117, N5350);
buf BUF1 (N12688, N12684);
xor XOR2 (N12689, N12686, N11930);
xor XOR2 (N12690, N12677, N8951);
not NOT1 (N12691, N12689);
nand NAND2 (N12692, N12681, N9037);
or OR2 (N12693, N12685, N2666);
buf BUF1 (N12694, N12690);
buf BUF1 (N12695, N12693);
or OR4 (N12696, N12691, N4607, N2796, N12382);
nor NOR2 (N12697, N12682, N7585);
not NOT1 (N12698, N12679);
not NOT1 (N12699, N12694);
buf BUF1 (N12700, N12695);
or OR4 (N12701, N12698, N3659, N7901, N5875);
buf BUF1 (N12702, N12696);
xor XOR2 (N12703, N12699, N828);
and AND3 (N12704, N12687, N12660, N11108);
not NOT1 (N12705, N12674);
buf BUF1 (N12706, N12672);
xor XOR2 (N12707, N12706, N9709);
buf BUF1 (N12708, N12703);
and AND2 (N12709, N12692, N4168);
nor NOR4 (N12710, N12708, N1300, N2210, N1437);
xor XOR2 (N12711, N12704, N5793);
not NOT1 (N12712, N12707);
not NOT1 (N12713, N12711);
xor XOR2 (N12714, N12697, N2618);
nor NOR4 (N12715, N12705, N4461, N4241, N7192);
buf BUF1 (N12716, N12715);
or OR3 (N12717, N12714, N8933, N868);
and AND3 (N12718, N12688, N7329, N9912);
xor XOR2 (N12719, N12712, N4246);
nand NAND2 (N12720, N12710, N4512);
nor NOR2 (N12721, N12719, N4415);
nand NAND2 (N12722, N12720, N1646);
and AND2 (N12723, N12713, N1797);
nor NOR2 (N12724, N12723, N7267);
and AND3 (N12725, N12709, N11458, N2946);
not NOT1 (N12726, N12717);
xor XOR2 (N12727, N12722, N4479);
nand NAND4 (N12728, N12718, N10102, N12663, N10091);
or OR3 (N12729, N12701, N12191, N7536);
not NOT1 (N12730, N12727);
xor XOR2 (N12731, N12729, N6829);
xor XOR2 (N12732, N12700, N10969);
nand NAND3 (N12733, N12702, N10323, N12619);
nand NAND4 (N12734, N12721, N10040, N11271, N3511);
and AND3 (N12735, N12726, N12211, N3924);
nand NAND3 (N12736, N12725, N8471, N2309);
buf BUF1 (N12737, N12732);
xor XOR2 (N12738, N12731, N1422);
buf BUF1 (N12739, N12736);
or OR4 (N12740, N12733, N3359, N6888, N6820);
buf BUF1 (N12741, N12740);
not NOT1 (N12742, N12734);
and AND3 (N12743, N12741, N9117, N4020);
nand NAND2 (N12744, N12739, N1778);
xor XOR2 (N12745, N12724, N7068);
and AND2 (N12746, N12738, N12105);
not NOT1 (N12747, N12744);
or OR4 (N12748, N12746, N7808, N1861, N11743);
and AND4 (N12749, N12743, N4, N10203, N11403);
or OR2 (N12750, N12745, N5177);
buf BUF1 (N12751, N12749);
and AND4 (N12752, N12737, N3766, N4760, N8805);
buf BUF1 (N12753, N12747);
xor XOR2 (N12754, N12752, N7068);
nor NOR2 (N12755, N12754, N6427);
not NOT1 (N12756, N12730);
nor NOR3 (N12757, N12742, N6522, N2768);
not NOT1 (N12758, N12735);
nor NOR4 (N12759, N12755, N1797, N4226, N3186);
or OR4 (N12760, N12728, N1094, N11857, N5788);
not NOT1 (N12761, N12751);
xor XOR2 (N12762, N12753, N11395);
or OR4 (N12763, N12761, N9567, N1256, N1257);
and AND3 (N12764, N12758, N12430, N7019);
buf BUF1 (N12765, N12716);
and AND3 (N12766, N12765, N7904, N12285);
nand NAND4 (N12767, N12750, N1945, N5369, N5908);
xor XOR2 (N12768, N12766, N6673);
not NOT1 (N12769, N12757);
or OR4 (N12770, N12763, N244, N6838, N10473);
nand NAND3 (N12771, N12768, N8448, N12170);
or OR2 (N12772, N12762, N11479);
xor XOR2 (N12773, N12772, N2601);
or OR3 (N12774, N12759, N6134, N889);
not NOT1 (N12775, N12756);
not NOT1 (N12776, N12764);
not NOT1 (N12777, N12748);
nand NAND2 (N12778, N12771, N3726);
not NOT1 (N12779, N12767);
buf BUF1 (N12780, N12776);
or OR2 (N12781, N12774, N11028);
not NOT1 (N12782, N12769);
buf BUF1 (N12783, N12773);
not NOT1 (N12784, N12778);
buf BUF1 (N12785, N12770);
nand NAND2 (N12786, N12783, N12222);
or OR3 (N12787, N12781, N11717, N2286);
buf BUF1 (N12788, N12785);
and AND3 (N12789, N12788, N9730, N12764);
and AND3 (N12790, N12779, N8270, N1603);
nand NAND2 (N12791, N12777, N12318);
not NOT1 (N12792, N12787);
buf BUF1 (N12793, N12791);
xor XOR2 (N12794, N12793, N10117);
buf BUF1 (N12795, N12782);
buf BUF1 (N12796, N12792);
xor XOR2 (N12797, N12789, N4890);
and AND2 (N12798, N12797, N7355);
and AND4 (N12799, N12798, N7233, N11288, N5878);
and AND4 (N12800, N12795, N6119, N2126, N10830);
not NOT1 (N12801, N12784);
and AND4 (N12802, N12786, N8496, N5634, N12332);
or OR4 (N12803, N12799, N4688, N2165, N10194);
nand NAND3 (N12804, N12790, N2024, N2906);
and AND4 (N12805, N12794, N6953, N8209, N678);
not NOT1 (N12806, N12805);
or OR3 (N12807, N12796, N6780, N9058);
or OR3 (N12808, N12760, N7027, N1896);
nor NOR3 (N12809, N12804, N1132, N8081);
nand NAND4 (N12810, N12775, N7901, N1697, N11604);
nand NAND3 (N12811, N12800, N7684, N2187);
buf BUF1 (N12812, N12801);
xor XOR2 (N12813, N12809, N399);
buf BUF1 (N12814, N12808);
buf BUF1 (N12815, N12780);
or OR2 (N12816, N12807, N11867);
buf BUF1 (N12817, N12813);
not NOT1 (N12818, N12816);
buf BUF1 (N12819, N12810);
nor NOR4 (N12820, N12806, N8966, N6989, N12436);
or OR3 (N12821, N12812, N3969, N4634);
nand NAND4 (N12822, N12818, N1135, N8838, N12359);
and AND3 (N12823, N12803, N2349, N6981);
and AND3 (N12824, N12820, N9848, N9704);
or OR3 (N12825, N12815, N578, N10114);
nor NOR2 (N12826, N12821, N8441);
nand NAND3 (N12827, N12825, N11416, N1420);
not NOT1 (N12828, N12826);
and AND2 (N12829, N12828, N10769);
xor XOR2 (N12830, N12811, N9552);
or OR2 (N12831, N12819, N7712);
xor XOR2 (N12832, N12827, N5822);
nor NOR3 (N12833, N12814, N3323, N6441);
and AND3 (N12834, N12817, N10629, N1272);
or OR2 (N12835, N12824, N1498);
or OR4 (N12836, N12802, N8907, N8741, N4425);
xor XOR2 (N12837, N12836, N1412);
and AND3 (N12838, N12830, N11817, N6983);
nand NAND3 (N12839, N12831, N6904, N6943);
or OR4 (N12840, N12829, N1988, N12198, N5141);
or OR3 (N12841, N12832, N4656, N8525);
nor NOR3 (N12842, N12834, N1837, N3848);
and AND2 (N12843, N12822, N5999);
nor NOR4 (N12844, N12835, N1311, N714, N3855);
and AND4 (N12845, N12843, N9657, N6876, N1010);
xor XOR2 (N12846, N12840, N10882);
nor NOR4 (N12847, N12845, N6137, N2232, N1490);
not NOT1 (N12848, N12844);
or OR4 (N12849, N12846, N11474, N286, N9233);
xor XOR2 (N12850, N12841, N10554);
xor XOR2 (N12851, N12849, N2343);
and AND3 (N12852, N12851, N4465, N8947);
not NOT1 (N12853, N12850);
and AND3 (N12854, N12847, N4785, N8147);
buf BUF1 (N12855, N12823);
or OR4 (N12856, N12848, N7526, N11809, N12584);
xor XOR2 (N12857, N12838, N12417);
buf BUF1 (N12858, N12855);
buf BUF1 (N12859, N12839);
nand NAND3 (N12860, N12854, N1671, N10799);
or OR3 (N12861, N12858, N11839, N4364);
or OR4 (N12862, N12842, N4967, N7820, N2290);
and AND3 (N12863, N12857, N8816, N6551);
nand NAND2 (N12864, N12859, N3644);
and AND3 (N12865, N12837, N9856, N135);
nand NAND4 (N12866, N12856, N4237, N7278, N9194);
not NOT1 (N12867, N12863);
nor NOR3 (N12868, N12864, N6782, N2858);
and AND4 (N12869, N12867, N401, N7001, N1370);
and AND3 (N12870, N12852, N3003, N2245);
and AND4 (N12871, N12869, N3872, N59, N8414);
or OR4 (N12872, N12853, N294, N2662, N3446);
xor XOR2 (N12873, N12866, N28);
not NOT1 (N12874, N12870);
nor NOR2 (N12875, N12872, N12035);
and AND4 (N12876, N12871, N8884, N11386, N10642);
xor XOR2 (N12877, N12865, N1367);
nand NAND3 (N12878, N12873, N12352, N7686);
nand NAND2 (N12879, N12877, N6635);
xor XOR2 (N12880, N12876, N1465);
and AND3 (N12881, N12874, N8949, N11049);
buf BUF1 (N12882, N12875);
or OR3 (N12883, N12868, N9949, N10068);
nand NAND3 (N12884, N12879, N4235, N12197);
nand NAND3 (N12885, N12833, N711, N7435);
nor NOR4 (N12886, N12880, N908, N3545, N7507);
or OR3 (N12887, N12886, N12870, N5897);
xor XOR2 (N12888, N12881, N575);
or OR4 (N12889, N12887, N7064, N10059, N12230);
xor XOR2 (N12890, N12885, N8758);
nor NOR3 (N12891, N12888, N8173, N4232);
xor XOR2 (N12892, N12883, N5593);
buf BUF1 (N12893, N12861);
and AND3 (N12894, N12891, N11199, N1849);
not NOT1 (N12895, N12890);
and AND3 (N12896, N12862, N4199, N4620);
nor NOR2 (N12897, N12884, N9701);
nand NAND4 (N12898, N12878, N12225, N2114, N12266);
xor XOR2 (N12899, N12898, N7821);
or OR2 (N12900, N12895, N7383);
and AND2 (N12901, N12899, N1272);
or OR3 (N12902, N12900, N7344, N4238);
and AND4 (N12903, N12892, N1531, N11358, N1120);
or OR4 (N12904, N12896, N9227, N8708, N4014);
and AND2 (N12905, N12860, N8340);
buf BUF1 (N12906, N12893);
nor NOR4 (N12907, N12904, N12616, N560, N3619);
nor NOR2 (N12908, N12897, N10210);
and AND3 (N12909, N12906, N7195, N9709);
xor XOR2 (N12910, N12903, N8392);
nand NAND2 (N12911, N12902, N9915);
not NOT1 (N12912, N12882);
xor XOR2 (N12913, N12909, N5729);
nor NOR3 (N12914, N12905, N4782, N11162);
or OR4 (N12915, N12889, N1927, N9854, N4224);
nand NAND2 (N12916, N12908, N8652);
not NOT1 (N12917, N12912);
xor XOR2 (N12918, N12915, N11280);
or OR3 (N12919, N12911, N1747, N9578);
or OR4 (N12920, N12918, N7747, N8127, N5704);
nand NAND2 (N12921, N12914, N9625);
not NOT1 (N12922, N12920);
or OR2 (N12923, N12921, N10016);
not NOT1 (N12924, N12923);
and AND3 (N12925, N12924, N10503, N6465);
nand NAND2 (N12926, N12917, N12293);
buf BUF1 (N12927, N12894);
nand NAND3 (N12928, N12919, N9122, N7835);
xor XOR2 (N12929, N12901, N8425);
nand NAND3 (N12930, N12913, N7251, N6642);
nor NOR2 (N12931, N12910, N3164);
nor NOR4 (N12932, N12907, N12102, N7477, N5373);
xor XOR2 (N12933, N12931, N2981);
not NOT1 (N12934, N12926);
nand NAND4 (N12935, N12927, N5400, N9179, N86);
and AND4 (N12936, N12925, N8370, N4527, N7240);
and AND4 (N12937, N12930, N4814, N1987, N12762);
or OR3 (N12938, N12929, N955, N774);
buf BUF1 (N12939, N12933);
xor XOR2 (N12940, N12937, N1879);
not NOT1 (N12941, N12932);
and AND2 (N12942, N12940, N4969);
nand NAND4 (N12943, N12936, N10496, N373, N7267);
xor XOR2 (N12944, N12943, N2549);
xor XOR2 (N12945, N12939, N6771);
and AND3 (N12946, N12945, N7963, N10506);
not NOT1 (N12947, N12935);
or OR2 (N12948, N12946, N6494);
xor XOR2 (N12949, N12922, N4406);
xor XOR2 (N12950, N12941, N2093);
and AND2 (N12951, N12934, N6875);
and AND4 (N12952, N12928, N6006, N1257, N1178);
nand NAND2 (N12953, N12916, N1913);
xor XOR2 (N12954, N12942, N581);
xor XOR2 (N12955, N12949, N4289);
and AND2 (N12956, N12938, N6361);
buf BUF1 (N12957, N12956);
buf BUF1 (N12958, N12952);
nand NAND2 (N12959, N12948, N4693);
nor NOR3 (N12960, N12951, N133, N7724);
not NOT1 (N12961, N12955);
and AND3 (N12962, N12950, N8110, N10562);
buf BUF1 (N12963, N12957);
and AND4 (N12964, N12954, N626, N8991, N5212);
not NOT1 (N12965, N12958);
xor XOR2 (N12966, N12964, N11813);
nor NOR4 (N12967, N12947, N4189, N2293, N6664);
or OR3 (N12968, N12944, N1446, N8556);
xor XOR2 (N12969, N12963, N1012);
nor NOR2 (N12970, N12967, N7422);
buf BUF1 (N12971, N12960);
not NOT1 (N12972, N12959);
not NOT1 (N12973, N12966);
and AND2 (N12974, N12968, N11354);
not NOT1 (N12975, N12973);
not NOT1 (N12976, N12974);
buf BUF1 (N12977, N12975);
or OR3 (N12978, N12972, N11348, N5558);
or OR2 (N12979, N12962, N9312);
and AND3 (N12980, N12976, N1385, N6736);
buf BUF1 (N12981, N12979);
nor NOR2 (N12982, N12981, N2161);
or OR3 (N12983, N12971, N5164, N12391);
and AND4 (N12984, N12961, N12872, N7032, N7920);
nand NAND2 (N12985, N12982, N10526);
not NOT1 (N12986, N12978);
or OR4 (N12987, N12985, N1105, N2937, N11733);
xor XOR2 (N12988, N12969, N7713);
xor XOR2 (N12989, N12970, N799);
and AND4 (N12990, N12984, N4899, N7060, N8433);
xor XOR2 (N12991, N12990, N6726);
and AND3 (N12992, N12965, N4461, N7317);
xor XOR2 (N12993, N12991, N6811);
or OR4 (N12994, N12992, N8460, N5024, N6519);
or OR4 (N12995, N12980, N4850, N2809, N9538);
xor XOR2 (N12996, N12993, N6697);
or OR3 (N12997, N12977, N5261, N8077);
and AND2 (N12998, N12989, N1878);
and AND3 (N12999, N12986, N4533, N7664);
buf BUF1 (N13000, N12997);
nand NAND2 (N13001, N12988, N5741);
or OR4 (N13002, N12994, N12439, N6035, N3947);
not NOT1 (N13003, N12983);
not NOT1 (N13004, N13003);
nand NAND3 (N13005, N13004, N11289, N6201);
and AND3 (N13006, N13001, N9441, N2141);
nor NOR3 (N13007, N12953, N10110, N5789);
or OR3 (N13008, N13000, N9405, N1903);
buf BUF1 (N13009, N13007);
not NOT1 (N13010, N13005);
nand NAND4 (N13011, N12996, N12922, N5074, N10017);
not NOT1 (N13012, N13002);
not NOT1 (N13013, N12987);
nor NOR2 (N13014, N13012, N43);
not NOT1 (N13015, N13010);
not NOT1 (N13016, N13009);
nand NAND4 (N13017, N12995, N11751, N2204, N12522);
or OR3 (N13018, N12998, N6981, N10774);
not NOT1 (N13019, N12999);
nor NOR2 (N13020, N13018, N2876);
nand NAND2 (N13021, N13006, N7724);
not NOT1 (N13022, N13011);
not NOT1 (N13023, N13017);
buf BUF1 (N13024, N13016);
nand NAND4 (N13025, N13023, N7438, N3099, N6389);
or OR4 (N13026, N13024, N10137, N3233, N1143);
xor XOR2 (N13027, N13013, N9294);
nand NAND4 (N13028, N13025, N8981, N1590, N4904);
xor XOR2 (N13029, N13020, N11004);
or OR4 (N13030, N13026, N12367, N3409, N5635);
and AND3 (N13031, N13015, N4227, N7098);
nor NOR2 (N13032, N13008, N111);
not NOT1 (N13033, N13019);
nor NOR3 (N13034, N13033, N10064, N2930);
and AND3 (N13035, N13030, N10873, N4760);
nor NOR4 (N13036, N13032, N2508, N6847, N5100);
or OR4 (N13037, N13031, N11593, N12513, N12254);
or OR2 (N13038, N13027, N4934);
nor NOR2 (N13039, N13022, N7067);
xor XOR2 (N13040, N13038, N3282);
nand NAND2 (N13041, N13028, N10726);
or OR4 (N13042, N13037, N375, N6543, N5704);
xor XOR2 (N13043, N13039, N12727);
nor NOR4 (N13044, N13042, N2190, N933, N3508);
xor XOR2 (N13045, N13041, N3141);
buf BUF1 (N13046, N13045);
not NOT1 (N13047, N13029);
nor NOR4 (N13048, N13043, N8487, N4705, N3742);
buf BUF1 (N13049, N13021);
and AND2 (N13050, N13046, N3083);
xor XOR2 (N13051, N13036, N4903);
nand NAND2 (N13052, N13014, N9685);
and AND3 (N13053, N13044, N3921, N8727);
not NOT1 (N13054, N13048);
buf BUF1 (N13055, N13054);
buf BUF1 (N13056, N13035);
nor NOR4 (N13057, N13055, N8424, N12223, N4341);
nor NOR3 (N13058, N13056, N8824, N12720);
buf BUF1 (N13059, N13053);
nor NOR2 (N13060, N13040, N7528);
or OR2 (N13061, N13034, N6043);
nor NOR3 (N13062, N13047, N2906, N11384);
nand NAND4 (N13063, N13050, N1825, N4696, N3828);
nor NOR4 (N13064, N13062, N7853, N2696, N8658);
not NOT1 (N13065, N13052);
nand NAND3 (N13066, N13058, N4637, N5715);
or OR2 (N13067, N13060, N9252);
or OR3 (N13068, N13066, N3819, N11090);
xor XOR2 (N13069, N13063, N11328);
nand NAND4 (N13070, N13068, N11906, N2823, N7281);
or OR3 (N13071, N13059, N5355, N3488);
nor NOR2 (N13072, N13057, N4925);
nor NOR2 (N13073, N13070, N5172);
nor NOR3 (N13074, N13049, N5029, N12277);
nor NOR3 (N13075, N13061, N8494, N5719);
buf BUF1 (N13076, N13071);
buf BUF1 (N13077, N13065);
nor NOR4 (N13078, N13076, N6402, N3327, N6563);
nor NOR2 (N13079, N13051, N1424);
xor XOR2 (N13080, N13077, N11688);
nor NOR4 (N13081, N13078, N8257, N3377, N967);
or OR2 (N13082, N13064, N1851);
nor NOR2 (N13083, N13072, N9180);
or OR3 (N13084, N13074, N9897, N1944);
buf BUF1 (N13085, N13082);
buf BUF1 (N13086, N13085);
nand NAND3 (N13087, N13084, N6938, N11127);
nand NAND4 (N13088, N13081, N11670, N49, N5406);
and AND3 (N13089, N13086, N1009, N6622);
nand NAND4 (N13090, N13089, N10744, N12568, N9606);
xor XOR2 (N13091, N13075, N2749);
and AND2 (N13092, N13087, N120);
buf BUF1 (N13093, N13092);
and AND2 (N13094, N13069, N206);
not NOT1 (N13095, N13090);
or OR4 (N13096, N13091, N1963, N7408, N3471);
nand NAND4 (N13097, N13088, N4071, N3318, N11319);
nand NAND4 (N13098, N13097, N5049, N3304, N4136);
buf BUF1 (N13099, N13083);
or OR2 (N13100, N13079, N4401);
xor XOR2 (N13101, N13080, N7592);
and AND4 (N13102, N13093, N3033, N921, N11313);
nor NOR3 (N13103, N13098, N1258, N4443);
nor NOR4 (N13104, N13096, N10699, N5358, N7154);
buf BUF1 (N13105, N13101);
nor NOR2 (N13106, N13105, N6595);
nand NAND4 (N13107, N13100, N5536, N8616, N2118);
buf BUF1 (N13108, N13102);
nand NAND4 (N13109, N13073, N3110, N12990, N6517);
or OR3 (N13110, N13099, N5956, N847);
nor NOR4 (N13111, N13104, N7375, N12860, N1381);
buf BUF1 (N13112, N13109);
nor NOR4 (N13113, N13111, N10612, N6018, N3352);
and AND2 (N13114, N13106, N2627);
nand NAND4 (N13115, N13113, N5663, N10808, N12508);
or OR2 (N13116, N13110, N7402);
buf BUF1 (N13117, N13067);
buf BUF1 (N13118, N13117);
xor XOR2 (N13119, N13115, N5865);
buf BUF1 (N13120, N13119);
nand NAND4 (N13121, N13120, N555, N11906, N4411);
xor XOR2 (N13122, N13116, N6266);
not NOT1 (N13123, N13118);
nand NAND4 (N13124, N13122, N588, N3741, N8992);
not NOT1 (N13125, N13095);
nor NOR3 (N13126, N13094, N11894, N1055);
xor XOR2 (N13127, N13107, N10778);
or OR4 (N13128, N13124, N11474, N1385, N13015);
nand NAND3 (N13129, N13128, N4650, N10509);
or OR4 (N13130, N13129, N11524, N9730, N1764);
not NOT1 (N13131, N13130);
nand NAND4 (N13132, N13112, N1934, N10616, N7328);
buf BUF1 (N13133, N13131);
and AND4 (N13134, N13103, N8547, N6674, N2355);
not NOT1 (N13135, N13126);
buf BUF1 (N13136, N13134);
nand NAND3 (N13137, N13114, N5914, N11032);
xor XOR2 (N13138, N13123, N5432);
nand NAND4 (N13139, N13138, N9300, N11735, N4607);
and AND3 (N13140, N13135, N752, N9627);
nor NOR4 (N13141, N13133, N10614, N12098, N4312);
xor XOR2 (N13142, N13137, N7893);
and AND3 (N13143, N13125, N9055, N11107);
not NOT1 (N13144, N13121);
nor NOR2 (N13145, N13140, N2665);
not NOT1 (N13146, N13132);
or OR3 (N13147, N13127, N591, N8044);
and AND4 (N13148, N13136, N7654, N6877, N2375);
or OR2 (N13149, N13142, N1331);
and AND3 (N13150, N13146, N1988, N7284);
not NOT1 (N13151, N13149);
xor XOR2 (N13152, N13108, N373);
not NOT1 (N13153, N13143);
nor NOR3 (N13154, N13141, N492, N4093);
nand NAND2 (N13155, N13151, N9277);
not NOT1 (N13156, N13154);
xor XOR2 (N13157, N13147, N8845);
and AND3 (N13158, N13156, N11665, N8598);
not NOT1 (N13159, N13139);
buf BUF1 (N13160, N13155);
not NOT1 (N13161, N13157);
xor XOR2 (N13162, N13153, N7144);
not NOT1 (N13163, N13150);
xor XOR2 (N13164, N13161, N9386);
and AND2 (N13165, N13152, N2603);
xor XOR2 (N13166, N13163, N10601);
nand NAND4 (N13167, N13148, N1202, N12713, N1733);
nand NAND4 (N13168, N13167, N12522, N2752, N12023);
and AND3 (N13169, N13144, N6475, N6208);
nand NAND2 (N13170, N13169, N2627);
or OR2 (N13171, N13160, N575);
and AND3 (N13172, N13165, N8584, N2945);
nand NAND4 (N13173, N13166, N7683, N4662, N8416);
xor XOR2 (N13174, N13170, N9785);
xor XOR2 (N13175, N13159, N7491);
not NOT1 (N13176, N13171);
nand NAND2 (N13177, N13176, N11626);
nand NAND4 (N13178, N13177, N11967, N5195, N4142);
and AND4 (N13179, N13158, N3385, N1830, N6427);
not NOT1 (N13180, N13178);
nor NOR2 (N13181, N13162, N6522);
not NOT1 (N13182, N13168);
buf BUF1 (N13183, N13182);
xor XOR2 (N13184, N13164, N9188);
xor XOR2 (N13185, N13173, N6189);
nand NAND2 (N13186, N13145, N11969);
xor XOR2 (N13187, N13174, N2074);
not NOT1 (N13188, N13184);
buf BUF1 (N13189, N13186);
and AND2 (N13190, N13189, N10904);
and AND3 (N13191, N13183, N1318, N9461);
and AND2 (N13192, N13188, N2320);
nand NAND3 (N13193, N13185, N8469, N10871);
and AND3 (N13194, N13190, N4215, N6386);
and AND3 (N13195, N13192, N6554, N5914);
nor NOR3 (N13196, N13194, N11509, N6584);
not NOT1 (N13197, N13179);
and AND3 (N13198, N13180, N7354, N10676);
nor NOR3 (N13199, N13172, N1175, N5904);
buf BUF1 (N13200, N13199);
buf BUF1 (N13201, N13198);
nand NAND2 (N13202, N13197, N12077);
nor NOR2 (N13203, N13193, N653);
or OR4 (N13204, N13191, N12342, N1441, N7569);
or OR2 (N13205, N13181, N11376);
buf BUF1 (N13206, N13201);
xor XOR2 (N13207, N13205, N9089);
xor XOR2 (N13208, N13206, N5047);
xor XOR2 (N13209, N13208, N12921);
or OR4 (N13210, N13204, N10119, N12682, N3530);
nand NAND3 (N13211, N13195, N2244, N3612);
not NOT1 (N13212, N13175);
buf BUF1 (N13213, N13187);
nor NOR4 (N13214, N13202, N3865, N11693, N6492);
nand NAND2 (N13215, N13203, N1566);
buf BUF1 (N13216, N13196);
nand NAND4 (N13217, N13210, N9137, N7906, N5573);
and AND3 (N13218, N13217, N5998, N1919);
nand NAND2 (N13219, N13214, N1858);
or OR3 (N13220, N13215, N6084, N9621);
or OR3 (N13221, N13213, N1589, N5872);
xor XOR2 (N13222, N13219, N1791);
buf BUF1 (N13223, N13212);
xor XOR2 (N13224, N13222, N3526);
or OR3 (N13225, N13211, N6605, N79);
and AND2 (N13226, N13220, N11727);
or OR4 (N13227, N13223, N4034, N6981, N6588);
nor NOR2 (N13228, N13218, N1956);
not NOT1 (N13229, N13227);
buf BUF1 (N13230, N13226);
not NOT1 (N13231, N13225);
nand NAND2 (N13232, N13221, N10712);
buf BUF1 (N13233, N13228);
and AND3 (N13234, N13231, N8125, N291);
buf BUF1 (N13235, N13234);
xor XOR2 (N13236, N13232, N8075);
nor NOR3 (N13237, N13209, N1755, N6082);
and AND4 (N13238, N13233, N9165, N2077, N10783);
nor NOR3 (N13239, N13230, N2326, N4309);
not NOT1 (N13240, N13239);
and AND2 (N13241, N13200, N9030);
or OR4 (N13242, N13229, N8247, N3804, N8511);
or OR4 (N13243, N13224, N7830, N1093, N3739);
nor NOR3 (N13244, N13235, N9677, N11341);
buf BUF1 (N13245, N13241);
xor XOR2 (N13246, N13238, N1376);
buf BUF1 (N13247, N13244);
xor XOR2 (N13248, N13240, N3104);
xor XOR2 (N13249, N13245, N8216);
nor NOR2 (N13250, N13246, N5973);
buf BUF1 (N13251, N13243);
buf BUF1 (N13252, N13216);
nor NOR3 (N13253, N13251, N7761, N327);
xor XOR2 (N13254, N13249, N12994);
buf BUF1 (N13255, N13250);
buf BUF1 (N13256, N13252);
buf BUF1 (N13257, N13253);
xor XOR2 (N13258, N13237, N7038);
or OR2 (N13259, N13254, N11832);
not NOT1 (N13260, N13259);
nand NAND2 (N13261, N13236, N6918);
nand NAND4 (N13262, N13256, N2643, N5987, N5787);
nand NAND4 (N13263, N13258, N9415, N10246, N2029);
or OR4 (N13264, N13263, N6687, N6419, N996);
and AND3 (N13265, N13207, N9169, N13262);
or OR4 (N13266, N1199, N10968, N7135, N7830);
and AND2 (N13267, N13247, N7611);
xor XOR2 (N13268, N13267, N11578);
buf BUF1 (N13269, N13266);
nand NAND4 (N13270, N13269, N7452, N12983, N9915);
xor XOR2 (N13271, N13242, N4451);
or OR4 (N13272, N13260, N714, N3096, N5653);
xor XOR2 (N13273, N13268, N11300);
xor XOR2 (N13274, N13273, N4743);
buf BUF1 (N13275, N13257);
buf BUF1 (N13276, N13265);
nor NOR4 (N13277, N13261, N3080, N1898, N5940);
or OR3 (N13278, N13276, N782, N7923);
or OR4 (N13279, N13255, N12598, N6970, N624);
nor NOR4 (N13280, N13271, N4301, N9738, N11843);
nand NAND2 (N13281, N13277, N2488);
buf BUF1 (N13282, N13248);
not NOT1 (N13283, N13280);
xor XOR2 (N13284, N13281, N9995);
not NOT1 (N13285, N13264);
nor NOR4 (N13286, N13275, N12493, N4553, N8946);
nand NAND2 (N13287, N13270, N294);
buf BUF1 (N13288, N13285);
nand NAND3 (N13289, N13282, N11012, N3077);
buf BUF1 (N13290, N13286);
buf BUF1 (N13291, N13288);
nand NAND2 (N13292, N13291, N4363);
or OR2 (N13293, N13279, N11268);
nand NAND2 (N13294, N13292, N3098);
or OR4 (N13295, N13283, N5712, N3428, N728);
xor XOR2 (N13296, N13284, N4730);
buf BUF1 (N13297, N13290);
buf BUF1 (N13298, N13296);
xor XOR2 (N13299, N13298, N921);
xor XOR2 (N13300, N13294, N5124);
not NOT1 (N13301, N13293);
or OR4 (N13302, N13300, N8854, N8780, N3896);
nor NOR2 (N13303, N13295, N3487);
nand NAND4 (N13304, N13303, N5980, N4620, N4045);
buf BUF1 (N13305, N13304);
not NOT1 (N13306, N13289);
and AND2 (N13307, N13302, N2535);
buf BUF1 (N13308, N13297);
nand NAND3 (N13309, N13305, N434, N13003);
and AND3 (N13310, N13274, N7929, N6008);
nor NOR2 (N13311, N13272, N12784);
nand NAND4 (N13312, N13287, N4216, N11681, N2430);
or OR4 (N13313, N13310, N624, N10769, N4899);
xor XOR2 (N13314, N13313, N981);
and AND3 (N13315, N13314, N11856, N1133);
nor NOR2 (N13316, N13311, N649);
not NOT1 (N13317, N13309);
not NOT1 (N13318, N13306);
not NOT1 (N13319, N13301);
nor NOR4 (N13320, N13299, N1974, N1993, N625);
and AND3 (N13321, N13318, N2098, N3461);
and AND3 (N13322, N13317, N10496, N887);
nor NOR3 (N13323, N13316, N435, N195);
buf BUF1 (N13324, N13315);
nor NOR2 (N13325, N13321, N9580);
not NOT1 (N13326, N13324);
buf BUF1 (N13327, N13322);
buf BUF1 (N13328, N13323);
and AND4 (N13329, N13320, N87, N811, N12792);
or OR4 (N13330, N13319, N6689, N10642, N5156);
nand NAND4 (N13331, N13325, N9638, N7405, N8994);
and AND2 (N13332, N13327, N9338);
nor NOR3 (N13333, N13307, N4382, N5142);
and AND3 (N13334, N13328, N4915, N5756);
and AND4 (N13335, N13329, N1648, N10393, N11996);
or OR4 (N13336, N13334, N12711, N6209, N10051);
not NOT1 (N13337, N13331);
xor XOR2 (N13338, N13336, N5728);
and AND4 (N13339, N13326, N3863, N6628, N9927);
not NOT1 (N13340, N13333);
and AND3 (N13341, N13332, N2706, N4578);
xor XOR2 (N13342, N13338, N9796);
nor NOR2 (N13343, N13335, N10031);
or OR2 (N13344, N13343, N9874);
nand NAND2 (N13345, N13340, N7348);
not NOT1 (N13346, N13345);
buf BUF1 (N13347, N13339);
nor NOR2 (N13348, N13342, N5494);
and AND2 (N13349, N13337, N12740);
buf BUF1 (N13350, N13341);
xor XOR2 (N13351, N13346, N2267);
buf BUF1 (N13352, N13308);
not NOT1 (N13353, N13348);
xor XOR2 (N13354, N13312, N10318);
buf BUF1 (N13355, N13344);
and AND3 (N13356, N13330, N3799, N10622);
nor NOR4 (N13357, N13347, N2434, N7218, N3201);
nor NOR2 (N13358, N13355, N1789);
nor NOR3 (N13359, N13349, N6334, N1725);
not NOT1 (N13360, N13357);
and AND4 (N13361, N13359, N8947, N8257, N11549);
nor NOR2 (N13362, N13361, N10388);
nand NAND4 (N13363, N13353, N8524, N6570, N2324);
xor XOR2 (N13364, N13360, N8839);
nor NOR2 (N13365, N13363, N13080);
nor NOR3 (N13366, N13351, N153, N4441);
or OR3 (N13367, N13356, N10534, N6127);
or OR2 (N13368, N13362, N6305);
or OR4 (N13369, N13358, N5032, N11355, N8084);
and AND3 (N13370, N13364, N9104, N12025);
nor NOR4 (N13371, N13370, N2938, N9959, N12516);
nand NAND3 (N13372, N13368, N7755, N8459);
or OR4 (N13373, N13371, N8703, N6091, N5014);
not NOT1 (N13374, N13278);
buf BUF1 (N13375, N13369);
or OR4 (N13376, N13375, N6275, N11117, N683);
and AND3 (N13377, N13366, N8750, N13311);
nor NOR4 (N13378, N13352, N9746, N2149, N13);
xor XOR2 (N13379, N13376, N2164);
not NOT1 (N13380, N13379);
or OR4 (N13381, N13377, N12453, N3378, N10515);
or OR2 (N13382, N13373, N11974);
nor NOR2 (N13383, N13382, N1431);
nor NOR2 (N13384, N13365, N9774);
not NOT1 (N13385, N13378);
nor NOR3 (N13386, N13381, N6503, N4857);
or OR2 (N13387, N13380, N5605);
xor XOR2 (N13388, N13374, N4520);
and AND2 (N13389, N13372, N4689);
and AND3 (N13390, N13367, N12209, N11809);
and AND3 (N13391, N13385, N8312, N10330);
nor NOR2 (N13392, N13391, N12192);
not NOT1 (N13393, N13384);
nand NAND4 (N13394, N13383, N3299, N4625, N8652);
or OR3 (N13395, N13392, N11618, N3043);
nor NOR3 (N13396, N13393, N11810, N1991);
xor XOR2 (N13397, N13390, N5142);
xor XOR2 (N13398, N13354, N3669);
or OR2 (N13399, N13389, N13254);
nor NOR3 (N13400, N13399, N6570, N7175);
nor NOR3 (N13401, N13394, N443, N5174);
nand NAND4 (N13402, N13397, N6885, N1006, N6883);
nor NOR4 (N13403, N13402, N12712, N210, N12355);
or OR2 (N13404, N13388, N5370);
buf BUF1 (N13405, N13404);
not NOT1 (N13406, N13403);
not NOT1 (N13407, N13395);
nor NOR3 (N13408, N13398, N1567, N5665);
xor XOR2 (N13409, N13350, N8133);
xor XOR2 (N13410, N13396, N7825);
nand NAND3 (N13411, N13400, N12358, N1410);
xor XOR2 (N13412, N13409, N12831);
nand NAND3 (N13413, N13410, N10496, N8836);
buf BUF1 (N13414, N13413);
or OR3 (N13415, N13407, N918, N8264);
buf BUF1 (N13416, N13386);
or OR4 (N13417, N13411, N8590, N10811, N6678);
nor NOR2 (N13418, N13408, N9171);
xor XOR2 (N13419, N13401, N2022);
nor NOR2 (N13420, N13415, N1038);
and AND3 (N13421, N13418, N6705, N5587);
buf BUF1 (N13422, N13412);
xor XOR2 (N13423, N13422, N7614);
and AND4 (N13424, N13405, N3877, N11600, N10162);
nand NAND2 (N13425, N13416, N10936);
or OR2 (N13426, N13421, N4502);
or OR2 (N13427, N13387, N8006);
buf BUF1 (N13428, N13426);
and AND2 (N13429, N13424, N1259);
not NOT1 (N13430, N13427);
or OR3 (N13431, N13414, N2527, N4341);
nor NOR4 (N13432, N13429, N8258, N5874, N12348);
nor NOR3 (N13433, N13423, N2368, N498);
not NOT1 (N13434, N13406);
nand NAND2 (N13435, N13428, N2532);
buf BUF1 (N13436, N13432);
nand NAND2 (N13437, N13435, N7051);
or OR4 (N13438, N13420, N5894, N781, N12602);
and AND2 (N13439, N13431, N12699);
or OR2 (N13440, N13430, N8762);
not NOT1 (N13441, N13440);
nand NAND2 (N13442, N13438, N11744);
xor XOR2 (N13443, N13434, N539);
nor NOR3 (N13444, N13436, N7848, N5256);
nor NOR3 (N13445, N13433, N7252, N8531);
xor XOR2 (N13446, N13441, N7962);
buf BUF1 (N13447, N13419);
xor XOR2 (N13448, N13444, N3801);
nand NAND2 (N13449, N13439, N2301);
not NOT1 (N13450, N13447);
buf BUF1 (N13451, N13449);
not NOT1 (N13452, N13437);
not NOT1 (N13453, N13445);
nor NOR4 (N13454, N13452, N7005, N13004, N12974);
buf BUF1 (N13455, N13450);
buf BUF1 (N13456, N13446);
or OR3 (N13457, N13417, N8697, N5171);
and AND3 (N13458, N13456, N9479, N10535);
nand NAND2 (N13459, N13425, N936);
not NOT1 (N13460, N13455);
and AND4 (N13461, N13442, N1099, N11509, N4115);
buf BUF1 (N13462, N13454);
not NOT1 (N13463, N13443);
buf BUF1 (N13464, N13461);
nor NOR3 (N13465, N13457, N11460, N1920);
xor XOR2 (N13466, N13458, N8129);
or OR2 (N13467, N13463, N11100);
not NOT1 (N13468, N13466);
nor NOR2 (N13469, N13451, N11679);
and AND4 (N13470, N13462, N1526, N5712, N5190);
xor XOR2 (N13471, N13467, N4813);
nor NOR4 (N13472, N13464, N7691, N7780, N13261);
buf BUF1 (N13473, N13471);
nor NOR3 (N13474, N13465, N854, N9118);
xor XOR2 (N13475, N13473, N8550);
not NOT1 (N13476, N13475);
buf BUF1 (N13477, N13472);
buf BUF1 (N13478, N13469);
buf BUF1 (N13479, N13478);
not NOT1 (N13480, N13460);
nor NOR3 (N13481, N13476, N9388, N11687);
and AND3 (N13482, N13479, N7310, N4050);
not NOT1 (N13483, N13448);
xor XOR2 (N13484, N13453, N10903);
or OR4 (N13485, N13474, N6095, N11306, N10978);
xor XOR2 (N13486, N13468, N5304);
and AND3 (N13487, N13484, N10662, N11205);
and AND4 (N13488, N13485, N2058, N8233, N13231);
nand NAND2 (N13489, N13487, N3979);
and AND3 (N13490, N13480, N10920, N8710);
xor XOR2 (N13491, N13477, N3213);
nand NAND2 (N13492, N13489, N11323);
nand NAND2 (N13493, N13488, N5929);
or OR4 (N13494, N13493, N10057, N13025, N8053);
and AND4 (N13495, N13481, N8474, N8452, N6318);
or OR2 (N13496, N13494, N115);
or OR3 (N13497, N13482, N11240, N4639);
nor NOR2 (N13498, N13490, N12614);
xor XOR2 (N13499, N13491, N2567);
buf BUF1 (N13500, N13470);
buf BUF1 (N13501, N13500);
and AND3 (N13502, N13495, N12430, N2697);
xor XOR2 (N13503, N13492, N5647);
or OR2 (N13504, N13498, N8498);
or OR2 (N13505, N13501, N4532);
nor NOR4 (N13506, N13497, N12577, N7327, N11971);
buf BUF1 (N13507, N13506);
xor XOR2 (N13508, N13504, N2584);
buf BUF1 (N13509, N13508);
or OR3 (N13510, N13503, N11480, N4137);
xor XOR2 (N13511, N13505, N5714);
and AND4 (N13512, N13459, N8476, N5206, N1718);
not NOT1 (N13513, N13483);
or OR3 (N13514, N13496, N2810, N7978);
or OR2 (N13515, N13507, N3976);
not NOT1 (N13516, N13502);
buf BUF1 (N13517, N13510);
and AND4 (N13518, N13515, N2103, N4949, N4344);
nor NOR3 (N13519, N13512, N6920, N7091);
nor NOR2 (N13520, N13514, N12580);
xor XOR2 (N13521, N13499, N7737);
xor XOR2 (N13522, N13486, N7132);
and AND2 (N13523, N13509, N1013);
nand NAND4 (N13524, N13520, N7939, N5142, N8471);
and AND2 (N13525, N13513, N3968);
buf BUF1 (N13526, N13523);
and AND3 (N13527, N13518, N13031, N6129);
not NOT1 (N13528, N13519);
not NOT1 (N13529, N13522);
and AND3 (N13530, N13526, N6760, N57);
nand NAND3 (N13531, N13525, N9602, N3717);
or OR3 (N13532, N13530, N1875, N3349);
buf BUF1 (N13533, N13516);
nor NOR4 (N13534, N13527, N10728, N4823, N1353);
not NOT1 (N13535, N13521);
not NOT1 (N13536, N13533);
or OR3 (N13537, N13517, N3016, N11727);
or OR2 (N13538, N13534, N759);
buf BUF1 (N13539, N13532);
xor XOR2 (N13540, N13531, N6085);
xor XOR2 (N13541, N13529, N7204);
and AND2 (N13542, N13539, N5971);
and AND4 (N13543, N13537, N11657, N7264, N1016);
not NOT1 (N13544, N13524);
nand NAND3 (N13545, N13540, N5191, N11237);
buf BUF1 (N13546, N13535);
xor XOR2 (N13547, N13541, N9883);
buf BUF1 (N13548, N13538);
buf BUF1 (N13549, N13542);
and AND3 (N13550, N13536, N6264, N7350);
buf BUF1 (N13551, N13544);
and AND4 (N13552, N13549, N10954, N7525, N788);
and AND2 (N13553, N13548, N11055);
nor NOR4 (N13554, N13552, N4769, N7492, N1762);
xor XOR2 (N13555, N13543, N10554);
and AND4 (N13556, N13511, N11408, N11122, N8472);
and AND4 (N13557, N13546, N8691, N8343, N3701);
nand NAND2 (N13558, N13557, N6350);
xor XOR2 (N13559, N13528, N6618);
and AND3 (N13560, N13550, N7010, N6187);
nand NAND4 (N13561, N13558, N9864, N11765, N12929);
xor XOR2 (N13562, N13553, N8905);
xor XOR2 (N13563, N13545, N12466);
xor XOR2 (N13564, N13561, N11493);
and AND4 (N13565, N13563, N9028, N12836, N12386);
xor XOR2 (N13566, N13564, N10639);
nor NOR2 (N13567, N13555, N2963);
not NOT1 (N13568, N13547);
nor NOR4 (N13569, N13566, N7399, N5109, N5561);
xor XOR2 (N13570, N13562, N2787);
nand NAND4 (N13571, N13570, N10528, N4078, N4025);
and AND2 (N13572, N13571, N6383);
and AND2 (N13573, N13559, N12586);
xor XOR2 (N13574, N13567, N6840);
not NOT1 (N13575, N13551);
nand NAND4 (N13576, N13560, N12046, N8405, N10559);
and AND2 (N13577, N13554, N9189);
and AND3 (N13578, N13573, N7751, N11636);
nor NOR3 (N13579, N13568, N6322, N11696);
xor XOR2 (N13580, N13575, N6038);
and AND2 (N13581, N13579, N7862);
nand NAND4 (N13582, N13556, N9528, N11099, N10931);
buf BUF1 (N13583, N13572);
xor XOR2 (N13584, N13580, N9006);
or OR4 (N13585, N13582, N2130, N6853, N6102);
nand NAND3 (N13586, N13577, N1535, N12925);
buf BUF1 (N13587, N13586);
and AND3 (N13588, N13574, N11273, N9728);
xor XOR2 (N13589, N13565, N3257);
nor NOR3 (N13590, N13588, N5231, N11652);
nand NAND4 (N13591, N13583, N6462, N5947, N6966);
nand NAND2 (N13592, N13589, N12916);
buf BUF1 (N13593, N13591);
not NOT1 (N13594, N13569);
nor NOR2 (N13595, N13581, N12459);
or OR3 (N13596, N13578, N342, N5086);
not NOT1 (N13597, N13594);
and AND2 (N13598, N13576, N11320);
buf BUF1 (N13599, N13597);
not NOT1 (N13600, N13584);
nand NAND3 (N13601, N13599, N13160, N11772);
or OR2 (N13602, N13593, N236);
and AND4 (N13603, N13601, N8128, N1720, N162);
buf BUF1 (N13604, N13585);
or OR2 (N13605, N13595, N3324);
nand NAND2 (N13606, N13598, N7501);
or OR3 (N13607, N13603, N13071, N4545);
or OR3 (N13608, N13606, N9065, N4486);
nor NOR2 (N13609, N13596, N11120);
not NOT1 (N13610, N13587);
or OR3 (N13611, N13590, N11558, N7051);
not NOT1 (N13612, N13605);
or OR4 (N13613, N13610, N17, N12784, N10712);
and AND3 (N13614, N13600, N9389, N1690);
nand NAND3 (N13615, N13604, N8052, N5773);
or OR4 (N13616, N13611, N10541, N995, N4551);
nand NAND4 (N13617, N13616, N4754, N4297, N10914);
and AND4 (N13618, N13607, N5836, N2330, N6719);
buf BUF1 (N13619, N13617);
buf BUF1 (N13620, N13609);
not NOT1 (N13621, N13592);
nand NAND3 (N13622, N13615, N1942, N851);
nand NAND4 (N13623, N13621, N12003, N2568, N835);
buf BUF1 (N13624, N13622);
nand NAND4 (N13625, N13624, N9644, N605, N10427);
xor XOR2 (N13626, N13618, N8374);
or OR2 (N13627, N13623, N546);
and AND2 (N13628, N13614, N3452);
and AND2 (N13629, N13628, N2026);
buf BUF1 (N13630, N13627);
or OR2 (N13631, N13619, N1939);
buf BUF1 (N13632, N13602);
not NOT1 (N13633, N13629);
nand NAND2 (N13634, N13631, N1106);
not NOT1 (N13635, N13625);
nor NOR3 (N13636, N13612, N13518, N9844);
nor NOR4 (N13637, N13613, N641, N8050, N238);
buf BUF1 (N13638, N13620);
nand NAND4 (N13639, N13626, N6911, N842, N13194);
not NOT1 (N13640, N13639);
or OR4 (N13641, N13608, N4271, N11110, N9538);
nand NAND4 (N13642, N13632, N9292, N1506, N9889);
not NOT1 (N13643, N13630);
and AND3 (N13644, N13638, N10051, N11595);
not NOT1 (N13645, N13637);
buf BUF1 (N13646, N13643);
not NOT1 (N13647, N13646);
and AND4 (N13648, N13634, N12563, N9251, N7645);
xor XOR2 (N13649, N13633, N10610);
buf BUF1 (N13650, N13641);
not NOT1 (N13651, N13644);
and AND2 (N13652, N13640, N12745);
or OR4 (N13653, N13645, N6285, N2093, N12958);
buf BUF1 (N13654, N13649);
buf BUF1 (N13655, N13636);
nand NAND3 (N13656, N13635, N7135, N7498);
nor NOR3 (N13657, N13656, N4425, N8567);
nor NOR2 (N13658, N13648, N1619);
xor XOR2 (N13659, N13650, N637);
or OR3 (N13660, N13658, N7710, N3094);
buf BUF1 (N13661, N13654);
or OR3 (N13662, N13653, N9809, N8127);
not NOT1 (N13663, N13659);
nand NAND3 (N13664, N13661, N10969, N8780);
and AND3 (N13665, N13655, N3265, N8060);
not NOT1 (N13666, N13662);
buf BUF1 (N13667, N13664);
buf BUF1 (N13668, N13651);
or OR3 (N13669, N13668, N2839, N1339);
or OR2 (N13670, N13663, N1448);
not NOT1 (N13671, N13657);
buf BUF1 (N13672, N13665);
not NOT1 (N13673, N13669);
or OR3 (N13674, N13667, N5394, N7872);
xor XOR2 (N13675, N13671, N1126);
not NOT1 (N13676, N13660);
not NOT1 (N13677, N13670);
and AND2 (N13678, N13666, N10975);
nor NOR4 (N13679, N13647, N10165, N2568, N11857);
and AND3 (N13680, N13673, N9586, N13417);
nor NOR4 (N13681, N13677, N533, N4442, N2443);
buf BUF1 (N13682, N13681);
nand NAND4 (N13683, N13652, N5393, N11585, N12032);
xor XOR2 (N13684, N13678, N6768);
not NOT1 (N13685, N13680);
or OR4 (N13686, N13672, N9337, N5428, N867);
nor NOR3 (N13687, N13642, N4328, N12803);
nand NAND3 (N13688, N13682, N5470, N6100);
buf BUF1 (N13689, N13676);
xor XOR2 (N13690, N13675, N13307);
xor XOR2 (N13691, N13690, N5476);
not NOT1 (N13692, N13683);
or OR3 (N13693, N13691, N11870, N4495);
and AND4 (N13694, N13684, N9046, N10114, N10186);
and AND4 (N13695, N13688, N6801, N857, N2086);
nand NAND2 (N13696, N13679, N8946);
nor NOR4 (N13697, N13694, N10591, N1612, N10537);
xor XOR2 (N13698, N13693, N23);
nor NOR2 (N13699, N13689, N7267);
or OR3 (N13700, N13698, N8890, N13529);
xor XOR2 (N13701, N13699, N3422);
not NOT1 (N13702, N13697);
xor XOR2 (N13703, N13686, N2616);
nand NAND4 (N13704, N13692, N5839, N11587, N1155);
nor NOR4 (N13705, N13702, N9081, N9478, N1176);
nor NOR3 (N13706, N13674, N8475, N1962);
xor XOR2 (N13707, N13700, N3769);
xor XOR2 (N13708, N13687, N10739);
not NOT1 (N13709, N13703);
and AND2 (N13710, N13709, N13158);
nand NAND2 (N13711, N13685, N9418);
buf BUF1 (N13712, N13696);
not NOT1 (N13713, N13705);
xor XOR2 (N13714, N13706, N11739);
xor XOR2 (N13715, N13707, N1645);
nand NAND4 (N13716, N13701, N34, N7751, N8361);
and AND2 (N13717, N13708, N9889);
buf BUF1 (N13718, N13714);
nand NAND3 (N13719, N13718, N10499, N12990);
not NOT1 (N13720, N13713);
nor NOR3 (N13721, N13719, N3953, N11755);
not NOT1 (N13722, N13711);
nor NOR3 (N13723, N13712, N1159, N7614);
xor XOR2 (N13724, N13695, N10777);
nor NOR4 (N13725, N13717, N12534, N2157, N10406);
buf BUF1 (N13726, N13724);
not NOT1 (N13727, N13716);
and AND3 (N13728, N13704, N10491, N10988);
not NOT1 (N13729, N13710);
not NOT1 (N13730, N13723);
and AND3 (N13731, N13725, N7353, N12347);
not NOT1 (N13732, N13731);
or OR3 (N13733, N13732, N13121, N13287);
and AND4 (N13734, N13730, N3921, N2345, N5249);
not NOT1 (N13735, N13733);
and AND3 (N13736, N13720, N13562, N4950);
and AND4 (N13737, N13721, N1547, N1430, N3390);
or OR4 (N13738, N13737, N10524, N7252, N10808);
xor XOR2 (N13739, N13722, N13193);
nor NOR3 (N13740, N13738, N9822, N5631);
not NOT1 (N13741, N13735);
not NOT1 (N13742, N13740);
and AND3 (N13743, N13728, N12357, N6471);
not NOT1 (N13744, N13734);
xor XOR2 (N13745, N13744, N8809);
nor NOR3 (N13746, N13742, N7581, N9816);
or OR4 (N13747, N13746, N8251, N9162, N10503);
or OR4 (N13748, N13739, N5322, N13521, N12141);
not NOT1 (N13749, N13736);
nor NOR3 (N13750, N13741, N1887, N13037);
buf BUF1 (N13751, N13726);
or OR3 (N13752, N13729, N9827, N927);
not NOT1 (N13753, N13743);
nand NAND4 (N13754, N13745, N7243, N998, N7163);
or OR2 (N13755, N13754, N1439);
or OR3 (N13756, N13751, N6739, N5529);
buf BUF1 (N13757, N13715);
nor NOR3 (N13758, N13756, N11254, N6729);
buf BUF1 (N13759, N13758);
and AND2 (N13760, N13727, N6356);
or OR2 (N13761, N13752, N3466);
nor NOR2 (N13762, N13748, N8206);
and AND3 (N13763, N13761, N1212, N10038);
xor XOR2 (N13764, N13755, N4334);
nand NAND3 (N13765, N13764, N8140, N1469);
or OR2 (N13766, N13750, N6388);
or OR3 (N13767, N13765, N13516, N9462);
and AND4 (N13768, N13753, N2136, N63, N2039);
xor XOR2 (N13769, N13757, N5710);
nor NOR4 (N13770, N13766, N4873, N7014, N6091);
not NOT1 (N13771, N13770);
buf BUF1 (N13772, N13747);
not NOT1 (N13773, N13759);
xor XOR2 (N13774, N13760, N12190);
and AND4 (N13775, N13749, N7441, N9535, N2525);
nand NAND2 (N13776, N13762, N5463);
xor XOR2 (N13777, N13774, N5859);
and AND3 (N13778, N13775, N13167, N6792);
nand NAND2 (N13779, N13763, N2114);
not NOT1 (N13780, N13777);
xor XOR2 (N13781, N13771, N7740);
nand NAND2 (N13782, N13778, N1051);
not NOT1 (N13783, N13776);
nand NAND2 (N13784, N13782, N12465);
not NOT1 (N13785, N13783);
nor NOR4 (N13786, N13780, N11513, N8017, N7972);
not NOT1 (N13787, N13784);
or OR3 (N13788, N13768, N1673, N590);
and AND4 (N13789, N13772, N1551, N12215, N1184);
buf BUF1 (N13790, N13767);
xor XOR2 (N13791, N13779, N13207);
and AND4 (N13792, N13791, N1300, N3229, N12694);
buf BUF1 (N13793, N13786);
nand NAND2 (N13794, N13785, N1945);
nand NAND2 (N13795, N13769, N3136);
buf BUF1 (N13796, N13790);
not NOT1 (N13797, N13781);
nor NOR3 (N13798, N13789, N12365, N1133);
buf BUF1 (N13799, N13793);
nand NAND3 (N13800, N13797, N7848, N1694);
buf BUF1 (N13801, N13795);
nand NAND3 (N13802, N13788, N3669, N3984);
nand NAND3 (N13803, N13800, N2414, N4817);
nand NAND2 (N13804, N13802, N7710);
and AND3 (N13805, N13803, N8385, N7500);
or OR3 (N13806, N13801, N13163, N350);
nor NOR2 (N13807, N13806, N12012);
not NOT1 (N13808, N13798);
buf BUF1 (N13809, N13807);
buf BUF1 (N13810, N13773);
xor XOR2 (N13811, N13808, N153);
buf BUF1 (N13812, N13792);
or OR3 (N13813, N13811, N3609, N13564);
nor NOR4 (N13814, N13805, N7373, N3746, N11875);
nand NAND3 (N13815, N13814, N11779, N5359);
or OR4 (N13816, N13804, N11186, N9002, N5778);
nand NAND3 (N13817, N13796, N4721, N4924);
buf BUF1 (N13818, N13816);
or OR3 (N13819, N13799, N2823, N6961);
nor NOR4 (N13820, N13819, N13024, N7817, N8721);
nor NOR2 (N13821, N13810, N5604);
nor NOR2 (N13822, N13815, N11978);
and AND4 (N13823, N13822, N596, N8298, N9876);
nand NAND4 (N13824, N13817, N11285, N8291, N5519);
not NOT1 (N13825, N13794);
not NOT1 (N13826, N13812);
and AND3 (N13827, N13821, N6915, N10197);
nand NAND2 (N13828, N13818, N13113);
buf BUF1 (N13829, N13809);
xor XOR2 (N13830, N13824, N386);
nand NAND4 (N13831, N13830, N11347, N1583, N8768);
or OR2 (N13832, N13787, N12081);
buf BUF1 (N13833, N13823);
xor XOR2 (N13834, N13832, N2455);
xor XOR2 (N13835, N13833, N10992);
buf BUF1 (N13836, N13829);
nor NOR3 (N13837, N13825, N3410, N13033);
and AND4 (N13838, N13820, N8946, N11460, N11414);
and AND4 (N13839, N13828, N6431, N12754, N4082);
nor NOR4 (N13840, N13835, N1506, N407, N8410);
nand NAND4 (N13841, N13836, N6367, N10404, N9301);
and AND3 (N13842, N13813, N11972, N4001);
buf BUF1 (N13843, N13839);
xor XOR2 (N13844, N13843, N4141);
nand NAND2 (N13845, N13826, N8664);
xor XOR2 (N13846, N13834, N5348);
xor XOR2 (N13847, N13837, N10825);
or OR3 (N13848, N13838, N8453, N2247);
not NOT1 (N13849, N13845);
or OR2 (N13850, N13849, N11423);
or OR3 (N13851, N13840, N7863, N13850);
nand NAND3 (N13852, N11429, N13399, N6450);
xor XOR2 (N13853, N13846, N9593);
nor NOR3 (N13854, N13853, N12194, N2043);
nor NOR2 (N13855, N13847, N8241);
or OR3 (N13856, N13831, N3016, N13199);
and AND3 (N13857, N13842, N2006, N9639);
not NOT1 (N13858, N13857);
nor NOR2 (N13859, N13856, N11698);
not NOT1 (N13860, N13855);
buf BUF1 (N13861, N13858);
or OR2 (N13862, N13861, N8377);
nor NOR4 (N13863, N13851, N6314, N4638, N10628);
and AND3 (N13864, N13844, N4909, N6626);
buf BUF1 (N13865, N13854);
not NOT1 (N13866, N13859);
nor NOR4 (N13867, N13864, N11204, N580, N10187);
buf BUF1 (N13868, N13863);
not NOT1 (N13869, N13866);
not NOT1 (N13870, N13862);
nor NOR2 (N13871, N13868, N9864);
nand NAND2 (N13872, N13865, N12161);
or OR2 (N13873, N13827, N6199);
buf BUF1 (N13874, N13872);
or OR2 (N13875, N13874, N9076);
and AND2 (N13876, N13875, N1186);
nand NAND3 (N13877, N13873, N3916, N12411);
nand NAND2 (N13878, N13877, N9313);
nor NOR2 (N13879, N13852, N5909);
buf BUF1 (N13880, N13878);
buf BUF1 (N13881, N13841);
not NOT1 (N13882, N13870);
buf BUF1 (N13883, N13871);
or OR2 (N13884, N13883, N8441);
buf BUF1 (N13885, N13869);
or OR3 (N13886, N13879, N12804, N414);
buf BUF1 (N13887, N13860);
xor XOR2 (N13888, N13882, N3416);
buf BUF1 (N13889, N13876);
not NOT1 (N13890, N13848);
xor XOR2 (N13891, N13887, N10169);
nor NOR2 (N13892, N13889, N2065);
not NOT1 (N13893, N13881);
and AND4 (N13894, N13885, N3411, N13820, N9949);
and AND2 (N13895, N13890, N2209);
nand NAND3 (N13896, N13880, N8793, N665);
buf BUF1 (N13897, N13891);
or OR4 (N13898, N13888, N5827, N13430, N5309);
and AND4 (N13899, N13886, N3717, N8578, N7588);
nor NOR2 (N13900, N13894, N3857);
xor XOR2 (N13901, N13893, N239);
xor XOR2 (N13902, N13898, N12032);
or OR2 (N13903, N13867, N229);
or OR3 (N13904, N13895, N10264, N11496);
and AND4 (N13905, N13902, N4318, N4614, N4615);
xor XOR2 (N13906, N13899, N11598);
not NOT1 (N13907, N13896);
and AND3 (N13908, N13904, N7582, N13355);
nor NOR4 (N13909, N13884, N6390, N8111, N8272);
and AND4 (N13910, N13905, N10435, N8925, N6224);
and AND2 (N13911, N13901, N13611);
buf BUF1 (N13912, N13911);
nand NAND2 (N13913, N13910, N12931);
nor NOR3 (N13914, N13892, N5967, N6010);
nand NAND4 (N13915, N13897, N6407, N5995, N3661);
or OR3 (N13916, N13914, N10919, N3878);
buf BUF1 (N13917, N13912);
or OR4 (N13918, N13913, N9817, N5622, N7631);
nor NOR3 (N13919, N13918, N10084, N6325);
nand NAND4 (N13920, N13900, N11553, N10905, N5025);
nand NAND4 (N13921, N13908, N8423, N5116, N11633);
nor NOR2 (N13922, N13919, N6320);
not NOT1 (N13923, N13906);
nand NAND4 (N13924, N13921, N10772, N11021, N55);
or OR4 (N13925, N13920, N3485, N10178, N4189);
nor NOR4 (N13926, N13903, N481, N2812, N3728);
not NOT1 (N13927, N13926);
or OR3 (N13928, N13925, N6888, N10136);
not NOT1 (N13929, N13922);
and AND3 (N13930, N13915, N5475, N5985);
nor NOR3 (N13931, N13928, N3417, N6608);
and AND2 (N13932, N13924, N9765);
buf BUF1 (N13933, N13930);
buf BUF1 (N13934, N13923);
or OR3 (N13935, N13909, N13049, N7411);
not NOT1 (N13936, N13933);
xor XOR2 (N13937, N13935, N3020);
not NOT1 (N13938, N13932);
xor XOR2 (N13939, N13934, N9983);
nor NOR3 (N13940, N13929, N5112, N3332);
nand NAND2 (N13941, N13936, N7651);
not NOT1 (N13942, N13927);
nand NAND3 (N13943, N13939, N10172, N5316);
or OR2 (N13944, N13941, N4023);
buf BUF1 (N13945, N13940);
and AND3 (N13946, N13943, N9510, N9151);
nor NOR4 (N13947, N13938, N8667, N4531, N11666);
not NOT1 (N13948, N13942);
xor XOR2 (N13949, N13917, N893);
buf BUF1 (N13950, N13949);
buf BUF1 (N13951, N13944);
nand NAND3 (N13952, N13916, N394, N689);
nand NAND4 (N13953, N13931, N11029, N2080, N2174);
nand NAND4 (N13954, N13951, N11384, N4525, N3);
or OR3 (N13955, N13946, N9149, N3691);
and AND4 (N13956, N13907, N7034, N13696, N6677);
or OR3 (N13957, N13950, N12477, N11723);
and AND4 (N13958, N13937, N2175, N1079, N5492);
and AND3 (N13959, N13956, N4658, N11312);
xor XOR2 (N13960, N13954, N6568);
not NOT1 (N13961, N13960);
nand NAND2 (N13962, N13952, N13499);
nand NAND2 (N13963, N13958, N12770);
and AND2 (N13964, N13947, N9986);
nor NOR4 (N13965, N13959, N13872, N11903, N261);
or OR4 (N13966, N13953, N5292, N897, N919);
and AND4 (N13967, N13964, N11031, N7727, N682);
or OR3 (N13968, N13963, N12830, N5897);
not NOT1 (N13969, N13962);
and AND4 (N13970, N13969, N13835, N8037, N9111);
buf BUF1 (N13971, N13967);
nand NAND3 (N13972, N13955, N4415, N12933);
or OR4 (N13973, N13948, N8389, N10624, N10488);
and AND3 (N13974, N13945, N7332, N8589);
nor NOR3 (N13975, N13968, N12998, N11035);
buf BUF1 (N13976, N13972);
not NOT1 (N13977, N13976);
or OR4 (N13978, N13970, N957, N5704, N194);
or OR4 (N13979, N13975, N12747, N2743, N6438);
nor NOR4 (N13980, N13974, N4759, N12303, N8034);
xor XOR2 (N13981, N13980, N2520);
nand NAND4 (N13982, N13965, N6398, N2519, N11267);
or OR2 (N13983, N13978, N5729);
not NOT1 (N13984, N13977);
not NOT1 (N13985, N13981);
nand NAND2 (N13986, N13984, N212);
buf BUF1 (N13987, N13961);
nand NAND4 (N13988, N13982, N21, N7778, N9730);
not NOT1 (N13989, N13983);
nand NAND2 (N13990, N13966, N5596);
not NOT1 (N13991, N13990);
nand NAND3 (N13992, N13987, N3130, N13395);
buf BUF1 (N13993, N13986);
nand NAND2 (N13994, N13971, N2851);
and AND3 (N13995, N13988, N8083, N392);
nor NOR4 (N13996, N13993, N11788, N6561, N3890);
nor NOR2 (N13997, N13996, N13797);
buf BUF1 (N13998, N13979);
buf BUF1 (N13999, N13991);
and AND2 (N14000, N13973, N1983);
buf BUF1 (N14001, N13957);
nor NOR4 (N14002, N13998, N2733, N12815, N12100);
and AND4 (N14003, N13995, N7404, N9093, N9345);
and AND4 (N14004, N13999, N305, N11496, N10539);
nor NOR2 (N14005, N13985, N2413);
nand NAND4 (N14006, N13989, N3398, N8559, N5477);
buf BUF1 (N14007, N14006);
nand NAND2 (N14008, N13994, N6963);
not NOT1 (N14009, N14001);
and AND4 (N14010, N14008, N2379, N726, N3052);
not NOT1 (N14011, N14003);
and AND3 (N14012, N14000, N12898, N3789);
buf BUF1 (N14013, N14010);
nor NOR3 (N14014, N13992, N1131, N9035);
or OR2 (N14015, N14009, N2166);
xor XOR2 (N14016, N14011, N9977);
nand NAND3 (N14017, N14016, N4087, N11574);
buf BUF1 (N14018, N14002);
buf BUF1 (N14019, N14014);
not NOT1 (N14020, N14013);
not NOT1 (N14021, N14019);
buf BUF1 (N14022, N14015);
and AND3 (N14023, N14007, N2812, N6466);
or OR4 (N14024, N14017, N10468, N7225, N1350);
buf BUF1 (N14025, N14012);
and AND2 (N14026, N14018, N8159);
nor NOR2 (N14027, N14023, N1257);
xor XOR2 (N14028, N13997, N8061);
xor XOR2 (N14029, N14026, N7606);
not NOT1 (N14030, N14028);
nand NAND2 (N14031, N14005, N11905);
or OR2 (N14032, N14025, N13186);
nor NOR4 (N14033, N14031, N3996, N13780, N8631);
or OR4 (N14034, N14004, N6136, N2289, N7364);
xor XOR2 (N14035, N14024, N9374);
xor XOR2 (N14036, N14033, N12111);
buf BUF1 (N14037, N14027);
buf BUF1 (N14038, N14030);
xor XOR2 (N14039, N14032, N9425);
buf BUF1 (N14040, N14039);
nand NAND2 (N14041, N14021, N13098);
not NOT1 (N14042, N14037);
xor XOR2 (N14043, N14036, N2729);
buf BUF1 (N14044, N14043);
not NOT1 (N14045, N14042);
nor NOR3 (N14046, N14034, N2526, N2005);
nor NOR4 (N14047, N14041, N3274, N1332, N3821);
nand NAND2 (N14048, N14040, N12905);
buf BUF1 (N14049, N14047);
and AND4 (N14050, N14038, N4344, N10826, N4723);
nand NAND2 (N14051, N14035, N12981);
buf BUF1 (N14052, N14045);
xor XOR2 (N14053, N14048, N9912);
buf BUF1 (N14054, N14051);
or OR2 (N14055, N14022, N3105);
and AND2 (N14056, N14049, N10854);
nor NOR3 (N14057, N14053, N4772, N1184);
not NOT1 (N14058, N14056);
or OR3 (N14059, N14058, N3075, N4150);
or OR3 (N14060, N14055, N1960, N12820);
or OR4 (N14061, N14060, N10177, N13499, N7271);
buf BUF1 (N14062, N14054);
or OR3 (N14063, N14061, N1223, N892);
nor NOR2 (N14064, N14029, N9986);
or OR4 (N14065, N14052, N4362, N9132, N1346);
nor NOR4 (N14066, N14050, N9492, N12073, N11714);
xor XOR2 (N14067, N14062, N5412);
not NOT1 (N14068, N14067);
not NOT1 (N14069, N14059);
or OR2 (N14070, N14064, N8851);
not NOT1 (N14071, N14057);
nand NAND3 (N14072, N14070, N1246, N10163);
xor XOR2 (N14073, N14071, N8901);
nor NOR4 (N14074, N14072, N2266, N11492, N2638);
nor NOR3 (N14075, N14065, N2981, N4073);
xor XOR2 (N14076, N14073, N12692);
nand NAND2 (N14077, N14066, N9985);
xor XOR2 (N14078, N14046, N3477);
nor NOR4 (N14079, N14069, N10027, N5797, N12259);
xor XOR2 (N14080, N14076, N5635);
buf BUF1 (N14081, N14068);
xor XOR2 (N14082, N14063, N4244);
xor XOR2 (N14083, N14081, N13250);
nand NAND2 (N14084, N14083, N10736);
and AND3 (N14085, N14044, N12849, N13892);
nor NOR3 (N14086, N14084, N12089, N11323);
nand NAND3 (N14087, N14077, N7041, N118);
buf BUF1 (N14088, N14075);
not NOT1 (N14089, N14087);
nand NAND4 (N14090, N14088, N7661, N9237, N4047);
not NOT1 (N14091, N14074);
or OR2 (N14092, N14085, N2287);
buf BUF1 (N14093, N14089);
buf BUF1 (N14094, N14090);
buf BUF1 (N14095, N14093);
xor XOR2 (N14096, N14078, N10626);
buf BUF1 (N14097, N14094);
not NOT1 (N14098, N14020);
buf BUF1 (N14099, N14095);
xor XOR2 (N14100, N14096, N12110);
not NOT1 (N14101, N14099);
buf BUF1 (N14102, N14091);
not NOT1 (N14103, N14101);
nand NAND4 (N14104, N14102, N4662, N5641, N651);
buf BUF1 (N14105, N14092);
nand NAND3 (N14106, N14097, N13788, N3959);
nand NAND4 (N14107, N14082, N10872, N8214, N4460);
and AND2 (N14108, N14106, N13746);
buf BUF1 (N14109, N14100);
nor NOR4 (N14110, N14109, N7325, N12845, N9264);
not NOT1 (N14111, N14104);
nor NOR3 (N14112, N14110, N14071, N6611);
not NOT1 (N14113, N14103);
buf BUF1 (N14114, N14079);
or OR3 (N14115, N14105, N2045, N7091);
nor NOR2 (N14116, N14098, N12365);
or OR2 (N14117, N14086, N4316);
buf BUF1 (N14118, N14111);
not NOT1 (N14119, N14118);
not NOT1 (N14120, N14107);
buf BUF1 (N14121, N14120);
not NOT1 (N14122, N14112);
nor NOR2 (N14123, N14119, N4713);
not NOT1 (N14124, N14123);
and AND4 (N14125, N14124, N8828, N6086, N2745);
or OR2 (N14126, N14122, N6715);
buf BUF1 (N14127, N14080);
or OR3 (N14128, N14108, N4813, N5791);
or OR2 (N14129, N14121, N9255);
nor NOR3 (N14130, N14113, N6180, N11724);
not NOT1 (N14131, N14130);
buf BUF1 (N14132, N14126);
or OR2 (N14133, N14114, N9158);
nand NAND4 (N14134, N14132, N10307, N4530, N1350);
and AND2 (N14135, N14127, N2105);
buf BUF1 (N14136, N14133);
nor NOR3 (N14137, N14115, N5812, N7269);
nor NOR2 (N14138, N14117, N6601);
not NOT1 (N14139, N14125);
nand NAND3 (N14140, N14116, N514, N1651);
xor XOR2 (N14141, N14134, N3429);
not NOT1 (N14142, N14139);
buf BUF1 (N14143, N14138);
xor XOR2 (N14144, N14141, N9514);
or OR2 (N14145, N14129, N9099);
nor NOR2 (N14146, N14143, N3003);
not NOT1 (N14147, N14136);
buf BUF1 (N14148, N14140);
or OR4 (N14149, N14142, N1232, N11017, N8312);
xor XOR2 (N14150, N14144, N3352);
buf BUF1 (N14151, N14146);
buf BUF1 (N14152, N14131);
nand NAND4 (N14153, N14148, N626, N13781, N13067);
nand NAND3 (N14154, N14152, N5193, N3118);
not NOT1 (N14155, N14137);
buf BUF1 (N14156, N14128);
and AND4 (N14157, N14155, N7639, N1494, N13784);
nor NOR2 (N14158, N14157, N3757);
nand NAND2 (N14159, N14147, N6279);
xor XOR2 (N14160, N14156, N8249);
nor NOR4 (N14161, N14158, N6382, N4994, N3236);
and AND3 (N14162, N14135, N3429, N3015);
or OR3 (N14163, N14162, N2203, N3020);
nor NOR3 (N14164, N14149, N7734, N6530);
and AND3 (N14165, N14161, N3145, N12650);
and AND4 (N14166, N14153, N6944, N3640, N9719);
nor NOR3 (N14167, N14150, N11533, N7724);
buf BUF1 (N14168, N14166);
nor NOR4 (N14169, N14165, N11755, N12637, N10305);
or OR2 (N14170, N14167, N11238);
nor NOR2 (N14171, N14160, N191);
or OR4 (N14172, N14164, N257, N7685, N6103);
nand NAND3 (N14173, N14159, N12777, N13968);
nor NOR4 (N14174, N14168, N9598, N5807, N5835);
and AND4 (N14175, N14173, N6844, N7805, N7291);
nand NAND3 (N14176, N14171, N13752, N2518);
nand NAND2 (N14177, N14163, N11951);
or OR3 (N14178, N14145, N8315, N3642);
buf BUF1 (N14179, N14174);
or OR3 (N14180, N14179, N11585, N13538);
or OR2 (N14181, N14180, N13544);
or OR4 (N14182, N14181, N8058, N13835, N928);
and AND2 (N14183, N14170, N3526);
buf BUF1 (N14184, N14169);
buf BUF1 (N14185, N14184);
nand NAND2 (N14186, N14182, N8186);
nor NOR3 (N14187, N14151, N9619, N12689);
xor XOR2 (N14188, N14186, N14143);
nor NOR3 (N14189, N14185, N4897, N11248);
nor NOR3 (N14190, N14188, N12610, N7694);
xor XOR2 (N14191, N14177, N13379);
and AND4 (N14192, N14190, N5518, N9728, N11058);
nand NAND3 (N14193, N14187, N8184, N2409);
not NOT1 (N14194, N14176);
not NOT1 (N14195, N14191);
xor XOR2 (N14196, N14194, N5241);
not NOT1 (N14197, N14178);
xor XOR2 (N14198, N14154, N8434);
and AND3 (N14199, N14192, N12195, N10493);
or OR2 (N14200, N14196, N4642);
nor NOR4 (N14201, N14195, N5986, N5537, N3334);
xor XOR2 (N14202, N14198, N8369);
xor XOR2 (N14203, N14172, N13689);
not NOT1 (N14204, N14201);
and AND4 (N14205, N14199, N712, N13451, N10645);
nor NOR2 (N14206, N14202, N13567);
and AND4 (N14207, N14189, N3176, N7489, N7299);
or OR2 (N14208, N14207, N9479);
nand NAND3 (N14209, N14197, N1721, N3719);
and AND4 (N14210, N14209, N21, N1441, N3613);
buf BUF1 (N14211, N14183);
buf BUF1 (N14212, N14204);
xor XOR2 (N14213, N14212, N1795);
or OR2 (N14214, N14175, N13450);
and AND4 (N14215, N14206, N9, N9685, N3098);
nand NAND2 (N14216, N14211, N7339);
nand NAND4 (N14217, N14193, N3735, N5640, N3783);
nor NOR3 (N14218, N14215, N8623, N9066);
buf BUF1 (N14219, N14213);
buf BUF1 (N14220, N14217);
not NOT1 (N14221, N14218);
nor NOR3 (N14222, N14216, N3326, N6743);
xor XOR2 (N14223, N14222, N10470);
nor NOR3 (N14224, N14220, N12181, N5907);
xor XOR2 (N14225, N14221, N13888);
and AND4 (N14226, N14214, N9871, N2669, N4037);
buf BUF1 (N14227, N14225);
nor NOR3 (N14228, N14226, N9458, N13700);
buf BUF1 (N14229, N14223);
and AND4 (N14230, N14200, N1516, N9729, N2946);
or OR3 (N14231, N14210, N9593, N5433);
or OR4 (N14232, N14227, N6847, N3021, N11489);
nand NAND2 (N14233, N14219, N5677);
and AND2 (N14234, N14233, N11700);
or OR3 (N14235, N14231, N11603, N9231);
not NOT1 (N14236, N14203);
xor XOR2 (N14237, N14208, N9031);
or OR4 (N14238, N14230, N1158, N7564, N4405);
nor NOR4 (N14239, N14205, N12934, N6729, N1895);
nand NAND2 (N14240, N14235, N3398);
and AND2 (N14241, N14238, N4630);
and AND3 (N14242, N14224, N6207, N5128);
and AND4 (N14243, N14240, N1304, N2097, N2605);
nand NAND3 (N14244, N14229, N5820, N4713);
xor XOR2 (N14245, N14228, N9311);
nand NAND3 (N14246, N14237, N9553, N5910);
xor XOR2 (N14247, N14242, N5774);
not NOT1 (N14248, N14232);
not NOT1 (N14249, N14239);
not NOT1 (N14250, N14236);
nand NAND2 (N14251, N14249, N7373);
nand NAND2 (N14252, N14245, N10389);
or OR3 (N14253, N14250, N7557, N5786);
buf BUF1 (N14254, N14241);
not NOT1 (N14255, N14251);
not NOT1 (N14256, N14248);
nor NOR3 (N14257, N14256, N14241, N11490);
not NOT1 (N14258, N14247);
not NOT1 (N14259, N14252);
buf BUF1 (N14260, N14243);
nor NOR3 (N14261, N14253, N9747, N7932);
xor XOR2 (N14262, N14246, N384);
and AND4 (N14263, N14259, N7711, N271, N13916);
nand NAND3 (N14264, N14262, N13550, N9637);
not NOT1 (N14265, N14234);
nand NAND2 (N14266, N14264, N11864);
nor NOR4 (N14267, N14265, N1856, N8199, N3549);
nor NOR2 (N14268, N14267, N13710);
or OR3 (N14269, N14263, N8676, N731);
and AND3 (N14270, N14261, N12246, N10468);
not NOT1 (N14271, N14258);
nand NAND3 (N14272, N14271, N5434, N13682);
or OR3 (N14273, N14272, N5959, N8957);
nand NAND4 (N14274, N14269, N840, N4438, N10660);
not NOT1 (N14275, N14255);
not NOT1 (N14276, N14270);
or OR2 (N14277, N14274, N4667);
or OR3 (N14278, N14254, N6063, N3065);
buf BUF1 (N14279, N14275);
or OR4 (N14280, N14276, N14231, N3289, N12997);
or OR2 (N14281, N14266, N525);
not NOT1 (N14282, N14278);
or OR4 (N14283, N14244, N5403, N1575, N7857);
and AND4 (N14284, N14260, N387, N508, N4730);
or OR3 (N14285, N14284, N6599, N2320);
buf BUF1 (N14286, N14281);
buf BUF1 (N14287, N14279);
nand NAND3 (N14288, N14268, N8351, N13497);
nor NOR2 (N14289, N14273, N11968);
xor XOR2 (N14290, N14285, N8942);
xor XOR2 (N14291, N14257, N13355);
not NOT1 (N14292, N14280);
or OR3 (N14293, N14283, N1670, N7643);
not NOT1 (N14294, N14282);
nand NAND3 (N14295, N14288, N13888, N11129);
or OR3 (N14296, N14286, N13874, N9032);
xor XOR2 (N14297, N14295, N13681);
buf BUF1 (N14298, N14293);
nor NOR3 (N14299, N14298, N7244, N6103);
not NOT1 (N14300, N14277);
and AND4 (N14301, N14291, N371, N12226, N4816);
or OR4 (N14302, N14292, N1815, N2082, N11818);
or OR3 (N14303, N14299, N10495, N12610);
not NOT1 (N14304, N14301);
buf BUF1 (N14305, N14290);
or OR4 (N14306, N14300, N9119, N5152, N7654);
nand NAND4 (N14307, N14305, N5417, N1845, N2811);
nand NAND4 (N14308, N14297, N677, N384, N13116);
and AND3 (N14309, N14306, N1287, N2814);
nor NOR3 (N14310, N14307, N7135, N10169);
not NOT1 (N14311, N14287);
not NOT1 (N14312, N14304);
nand NAND3 (N14313, N14296, N12091, N11825);
nand NAND4 (N14314, N14302, N3907, N13233, N8436);
buf BUF1 (N14315, N14314);
not NOT1 (N14316, N14311);
and AND2 (N14317, N14310, N5653);
nor NOR3 (N14318, N14313, N3887, N13355);
nor NOR2 (N14319, N14315, N9078);
xor XOR2 (N14320, N14308, N5430);
not NOT1 (N14321, N14289);
nand NAND2 (N14322, N14318, N5114);
nor NOR2 (N14323, N14294, N9666);
not NOT1 (N14324, N14322);
not NOT1 (N14325, N14320);
or OR3 (N14326, N14323, N987, N12858);
buf BUF1 (N14327, N14303);
nor NOR4 (N14328, N14316, N13348, N11493, N8046);
or OR4 (N14329, N14309, N8867, N10696, N10569);
buf BUF1 (N14330, N14326);
and AND3 (N14331, N14330, N10186, N11129);
not NOT1 (N14332, N14325);
or OR3 (N14333, N14317, N463, N4204);
nor NOR4 (N14334, N14332, N8807, N2227, N10709);
not NOT1 (N14335, N14334);
nor NOR2 (N14336, N14324, N9212);
not NOT1 (N14337, N14335);
nand NAND3 (N14338, N14321, N2920, N10399);
buf BUF1 (N14339, N14329);
buf BUF1 (N14340, N14331);
or OR2 (N14341, N14327, N7365);
and AND3 (N14342, N14333, N11802, N8993);
nor NOR2 (N14343, N14337, N11012);
and AND2 (N14344, N14341, N10372);
nand NAND3 (N14345, N14343, N1603, N1375);
xor XOR2 (N14346, N14340, N8309);
xor XOR2 (N14347, N14336, N6330);
buf BUF1 (N14348, N14342);
and AND4 (N14349, N14312, N10367, N12358, N8271);
xor XOR2 (N14350, N14347, N10368);
buf BUF1 (N14351, N14338);
nor NOR3 (N14352, N14351, N10590, N4339);
or OR4 (N14353, N14346, N8415, N7381, N10168);
or OR4 (N14354, N14328, N4892, N9991, N1766);
not NOT1 (N14355, N14352);
nand NAND4 (N14356, N14345, N14162, N2288, N1857);
xor XOR2 (N14357, N14339, N9139);
nor NOR3 (N14358, N14319, N2864, N1401);
nor NOR2 (N14359, N14348, N8480);
and AND2 (N14360, N14357, N11919);
xor XOR2 (N14361, N14353, N11006);
or OR4 (N14362, N14355, N3544, N8715, N10937);
nand NAND4 (N14363, N14360, N10356, N11044, N1812);
xor XOR2 (N14364, N14356, N12453);
buf BUF1 (N14365, N14363);
or OR4 (N14366, N14358, N13952, N2054, N2743);
and AND4 (N14367, N14362, N5068, N12506, N10481);
nand NAND2 (N14368, N14367, N858);
nor NOR3 (N14369, N14344, N5543, N3168);
buf BUF1 (N14370, N14366);
nand NAND3 (N14371, N14354, N10666, N11900);
and AND4 (N14372, N14361, N4048, N2437, N8530);
not NOT1 (N14373, N14350);
nand NAND3 (N14374, N14365, N8979, N2980);
or OR2 (N14375, N14368, N1463);
nor NOR3 (N14376, N14373, N7315, N13836);
and AND3 (N14377, N14359, N3546, N1464);
buf BUF1 (N14378, N14375);
nor NOR4 (N14379, N14369, N12516, N372, N7875);
or OR2 (N14380, N14364, N1354);
or OR2 (N14381, N14371, N6182);
xor XOR2 (N14382, N14377, N14321);
buf BUF1 (N14383, N14370);
not NOT1 (N14384, N14382);
xor XOR2 (N14385, N14374, N12242);
buf BUF1 (N14386, N14372);
xor XOR2 (N14387, N14383, N8075);
xor XOR2 (N14388, N14387, N3388);
and AND4 (N14389, N14378, N9389, N10543, N7825);
nand NAND2 (N14390, N14381, N3204);
nor NOR4 (N14391, N14380, N10023, N9319, N7576);
buf BUF1 (N14392, N14391);
nand NAND3 (N14393, N14389, N9242, N3177);
and AND3 (N14394, N14385, N14218, N2438);
xor XOR2 (N14395, N14376, N10633);
or OR4 (N14396, N14393, N10760, N2575, N2185);
buf BUF1 (N14397, N14384);
or OR3 (N14398, N14349, N5826, N1728);
not NOT1 (N14399, N14395);
xor XOR2 (N14400, N14398, N12954);
or OR3 (N14401, N14400, N5023, N11274);
or OR2 (N14402, N14388, N8218);
not NOT1 (N14403, N14397);
nand NAND2 (N14404, N14390, N2509);
nand NAND2 (N14405, N14396, N9550);
nand NAND4 (N14406, N14392, N3483, N3739, N598);
nor NOR3 (N14407, N14401, N13885, N928);
nor NOR4 (N14408, N14407, N13542, N14075, N2676);
xor XOR2 (N14409, N14406, N8196);
or OR3 (N14410, N14379, N14394, N2160);
and AND4 (N14411, N5545, N2775, N10701, N12721);
or OR3 (N14412, N14403, N1529, N5798);
and AND4 (N14413, N14412, N6957, N12111, N9886);
or OR3 (N14414, N14410, N5843, N12196);
or OR2 (N14415, N14409, N7310);
xor XOR2 (N14416, N14411, N2579);
nand NAND2 (N14417, N14413, N10939);
or OR2 (N14418, N14402, N11487);
nor NOR4 (N14419, N14404, N3478, N5147, N4107);
buf BUF1 (N14420, N14386);
not NOT1 (N14421, N14420);
and AND4 (N14422, N14405, N8521, N6533, N11235);
xor XOR2 (N14423, N14408, N8634);
nand NAND3 (N14424, N14423, N5214, N11111);
xor XOR2 (N14425, N14419, N2873);
nor NOR4 (N14426, N14418, N5819, N1674, N392);
not NOT1 (N14427, N14399);
nor NOR4 (N14428, N14415, N12303, N843, N8474);
xor XOR2 (N14429, N14426, N1848);
xor XOR2 (N14430, N14414, N10031);
nand NAND3 (N14431, N14425, N7538, N9484);
and AND2 (N14432, N14422, N12001);
not NOT1 (N14433, N14417);
nand NAND3 (N14434, N14421, N13201, N11799);
nor NOR3 (N14435, N14429, N9079, N9283);
or OR3 (N14436, N14430, N3243, N1658);
xor XOR2 (N14437, N14428, N11440);
buf BUF1 (N14438, N14432);
nand NAND3 (N14439, N14433, N5622, N7135);
and AND2 (N14440, N14431, N3969);
buf BUF1 (N14441, N14436);
nor NOR4 (N14442, N14434, N7563, N3836, N7100);
xor XOR2 (N14443, N14416, N5134);
not NOT1 (N14444, N14442);
buf BUF1 (N14445, N14435);
buf BUF1 (N14446, N14444);
nor NOR4 (N14447, N14446, N10726, N3770, N8912);
buf BUF1 (N14448, N14441);
or OR4 (N14449, N14445, N10195, N417, N13016);
nand NAND3 (N14450, N14447, N4776, N11018);
nand NAND2 (N14451, N14439, N1547);
nand NAND2 (N14452, N14440, N1088);
and AND3 (N14453, N14450, N8412, N12522);
or OR3 (N14454, N14451, N3781, N937);
nand NAND2 (N14455, N14424, N11736);
nand NAND4 (N14456, N14438, N9696, N10443, N11985);
buf BUF1 (N14457, N14448);
or OR4 (N14458, N14453, N4301, N1018, N10607);
and AND4 (N14459, N14458, N6765, N9822, N12532);
nand NAND2 (N14460, N14437, N8407);
xor XOR2 (N14461, N14454, N6392);
xor XOR2 (N14462, N14456, N11307);
and AND2 (N14463, N14449, N9896);
and AND4 (N14464, N14452, N4596, N5492, N3821);
xor XOR2 (N14465, N14464, N1562);
xor XOR2 (N14466, N14462, N12473);
nor NOR4 (N14467, N14443, N11170, N6070, N14419);
buf BUF1 (N14468, N14466);
xor XOR2 (N14469, N14457, N5693);
or OR3 (N14470, N14460, N8914, N3069);
nand NAND3 (N14471, N14455, N929, N1719);
buf BUF1 (N14472, N14463);
not NOT1 (N14473, N14459);
not NOT1 (N14474, N14461);
or OR3 (N14475, N14471, N587, N3924);
and AND3 (N14476, N14474, N10364, N5143);
and AND4 (N14477, N14465, N612, N2050, N6448);
not NOT1 (N14478, N14427);
nand NAND2 (N14479, N14472, N359);
nor NOR4 (N14480, N14476, N7358, N13587, N2423);
and AND3 (N14481, N14480, N5113, N116);
nand NAND4 (N14482, N14479, N7140, N8842, N4917);
not NOT1 (N14483, N14482);
or OR3 (N14484, N14481, N9590, N653);
not NOT1 (N14485, N14468);
xor XOR2 (N14486, N14470, N7138);
or OR2 (N14487, N14473, N13430);
xor XOR2 (N14488, N14477, N8766);
or OR2 (N14489, N14478, N13023);
buf BUF1 (N14490, N14487);
or OR4 (N14491, N14467, N11842, N11159, N10564);
nand NAND2 (N14492, N14475, N10231);
and AND3 (N14493, N14485, N3732, N3354);
not NOT1 (N14494, N14489);
xor XOR2 (N14495, N14493, N14353);
nand NAND3 (N14496, N14488, N1607, N7276);
nand NAND4 (N14497, N14494, N5236, N3715, N12543);
or OR4 (N14498, N14469, N9568, N9543, N1718);
buf BUF1 (N14499, N14497);
nand NAND2 (N14500, N14495, N8790);
and AND3 (N14501, N14496, N4512, N5532);
not NOT1 (N14502, N14491);
or OR3 (N14503, N14483, N5533, N7997);
buf BUF1 (N14504, N14486);
not NOT1 (N14505, N14503);
xor XOR2 (N14506, N14490, N8356);
not NOT1 (N14507, N14492);
buf BUF1 (N14508, N14501);
and AND3 (N14509, N14498, N11930, N915);
and AND4 (N14510, N14506, N3938, N1665, N6843);
not NOT1 (N14511, N14504);
xor XOR2 (N14512, N14499, N13009);
nor NOR2 (N14513, N14511, N8448);
or OR3 (N14514, N14510, N10030, N8192);
nor NOR4 (N14515, N14502, N14050, N4950, N3878);
or OR2 (N14516, N14512, N12721);
nand NAND2 (N14517, N14513, N2469);
and AND4 (N14518, N14515, N8610, N1869, N3364);
or OR3 (N14519, N14518, N8200, N11391);
or OR2 (N14520, N14516, N13413);
nand NAND4 (N14521, N14520, N8105, N10870, N2083);
and AND3 (N14522, N14517, N8496, N9854);
or OR2 (N14523, N14514, N355);
and AND4 (N14524, N14509, N1661, N1557, N4980);
buf BUF1 (N14525, N14521);
buf BUF1 (N14526, N14525);
buf BUF1 (N14527, N14508);
or OR4 (N14528, N14507, N13104, N1053, N12990);
buf BUF1 (N14529, N14524);
and AND2 (N14530, N14529, N372);
not NOT1 (N14531, N14522);
or OR4 (N14532, N14484, N1007, N708, N1788);
nor NOR2 (N14533, N14530, N11319);
not NOT1 (N14534, N14526);
xor XOR2 (N14535, N14500, N2109);
nor NOR2 (N14536, N14531, N12886);
nand NAND4 (N14537, N14536, N1727, N8019, N12420);
buf BUF1 (N14538, N14519);
xor XOR2 (N14539, N14534, N9050);
not NOT1 (N14540, N14533);
nand NAND2 (N14541, N14523, N1888);
xor XOR2 (N14542, N14535, N9322);
buf BUF1 (N14543, N14505);
or OR4 (N14544, N14527, N10914, N3432, N1000);
nand NAND2 (N14545, N14544, N651);
and AND4 (N14546, N14543, N7575, N2418, N12358);
or OR4 (N14547, N14542, N7774, N5794, N8165);
buf BUF1 (N14548, N14538);
not NOT1 (N14549, N14532);
nor NOR3 (N14550, N14547, N2511, N12098);
buf BUF1 (N14551, N14539);
nand NAND3 (N14552, N14537, N10808, N6921);
or OR4 (N14553, N14546, N11015, N2623, N8047);
and AND3 (N14554, N14540, N498, N5246);
and AND4 (N14555, N14548, N12755, N7998, N1522);
buf BUF1 (N14556, N14549);
xor XOR2 (N14557, N14554, N7289);
xor XOR2 (N14558, N14556, N7251);
not NOT1 (N14559, N14552);
not NOT1 (N14560, N14558);
and AND2 (N14561, N14555, N9009);
xor XOR2 (N14562, N14557, N4241);
not NOT1 (N14563, N14550);
not NOT1 (N14564, N14553);
buf BUF1 (N14565, N14551);
or OR3 (N14566, N14564, N690, N6018);
or OR4 (N14567, N14566, N6224, N12667, N1494);
not NOT1 (N14568, N14541);
not NOT1 (N14569, N14567);
or OR2 (N14570, N14568, N2810);
nor NOR2 (N14571, N14560, N4070);
not NOT1 (N14572, N14528);
nand NAND4 (N14573, N14571, N4053, N5740, N11723);
xor XOR2 (N14574, N14572, N5301);
buf BUF1 (N14575, N14570);
buf BUF1 (N14576, N14573);
or OR2 (N14577, N14563, N12310);
nand NAND4 (N14578, N14561, N9444, N3982, N8732);
and AND3 (N14579, N14569, N14200, N6867);
not NOT1 (N14580, N14559);
not NOT1 (N14581, N14579);
buf BUF1 (N14582, N14578);
and AND4 (N14583, N14576, N11547, N9410, N13888);
nor NOR3 (N14584, N14581, N10423, N6426);
not NOT1 (N14585, N14565);
and AND4 (N14586, N14580, N7254, N6521, N10873);
and AND3 (N14587, N14584, N677, N9299);
xor XOR2 (N14588, N14562, N7121);
not NOT1 (N14589, N14585);
and AND4 (N14590, N14577, N2980, N3253, N10468);
buf BUF1 (N14591, N14582);
nand NAND2 (N14592, N14545, N4651);
nor NOR4 (N14593, N14574, N12279, N9413, N1248);
and AND4 (N14594, N14590, N5447, N1069, N12950);
nor NOR4 (N14595, N14593, N8409, N8164, N4362);
nor NOR2 (N14596, N14592, N2824);
not NOT1 (N14597, N14587);
nand NAND3 (N14598, N14575, N9955, N3575);
xor XOR2 (N14599, N14583, N12835);
xor XOR2 (N14600, N14597, N3334);
xor XOR2 (N14601, N14596, N13083);
nor NOR3 (N14602, N14599, N9764, N14271);
nor NOR4 (N14603, N14601, N5012, N7584, N8770);
nand NAND3 (N14604, N14588, N4790, N814);
nand NAND4 (N14605, N14595, N1682, N8911, N3491);
nand NAND3 (N14606, N14586, N2963, N5916);
xor XOR2 (N14607, N14594, N229);
nand NAND3 (N14608, N14605, N1649, N3778);
nor NOR2 (N14609, N14604, N2075);
and AND3 (N14610, N14598, N13809, N12230);
not NOT1 (N14611, N14591);
nor NOR3 (N14612, N14611, N12396, N11408);
not NOT1 (N14613, N14602);
nand NAND4 (N14614, N14606, N3559, N6715, N1827);
xor XOR2 (N14615, N14614, N4784);
xor XOR2 (N14616, N14600, N10088);
nor NOR2 (N14617, N14603, N10902);
nand NAND4 (N14618, N14613, N648, N772, N848);
and AND3 (N14619, N14612, N1048, N7113);
and AND2 (N14620, N14618, N1836);
and AND4 (N14621, N14615, N9466, N11109, N8128);
or OR2 (N14622, N14589, N6610);
buf BUF1 (N14623, N14619);
xor XOR2 (N14624, N14620, N13314);
nand NAND3 (N14625, N14608, N4128, N11341);
or OR2 (N14626, N14625, N7473);
xor XOR2 (N14627, N14609, N10899);
and AND4 (N14628, N14607, N1787, N337, N5976);
nor NOR2 (N14629, N14622, N12744);
or OR2 (N14630, N14623, N3902);
nor NOR3 (N14631, N14617, N8568, N6913);
nor NOR3 (N14632, N14629, N2083, N6985);
xor XOR2 (N14633, N14616, N10240);
and AND2 (N14634, N14630, N12203);
xor XOR2 (N14635, N14633, N3998);
and AND4 (N14636, N14627, N12075, N2804, N7569);
nor NOR2 (N14637, N14624, N2427);
buf BUF1 (N14638, N14636);
nand NAND3 (N14639, N14634, N9596, N8689);
or OR3 (N14640, N14637, N2504, N1601);
and AND2 (N14641, N14621, N13927);
buf BUF1 (N14642, N14639);
nand NAND3 (N14643, N14638, N7229, N4793);
xor XOR2 (N14644, N14632, N7680);
xor XOR2 (N14645, N14628, N11136);
xor XOR2 (N14646, N14641, N8899);
not NOT1 (N14647, N14640);
not NOT1 (N14648, N14644);
not NOT1 (N14649, N14646);
xor XOR2 (N14650, N14648, N11468);
and AND4 (N14651, N14610, N9056, N7875, N1505);
nand NAND4 (N14652, N14649, N741, N5631, N6164);
xor XOR2 (N14653, N14647, N5808);
or OR4 (N14654, N14643, N5347, N1731, N3922);
and AND3 (N14655, N14635, N11351, N1943);
xor XOR2 (N14656, N14645, N5804);
nor NOR2 (N14657, N14650, N11021);
and AND2 (N14658, N14654, N11415);
and AND2 (N14659, N14653, N12199);
buf BUF1 (N14660, N14642);
not NOT1 (N14661, N14655);
nor NOR4 (N14662, N14661, N6105, N8274, N11446);
nand NAND3 (N14663, N14657, N6797, N14650);
xor XOR2 (N14664, N14662, N12610);
nor NOR4 (N14665, N14631, N11450, N5170, N11096);
and AND4 (N14666, N14658, N4281, N11859, N11675);
nor NOR4 (N14667, N14660, N11117, N3993, N12143);
nand NAND2 (N14668, N14656, N4796);
or OR2 (N14669, N14666, N13058);
nand NAND4 (N14670, N14669, N6574, N324, N2229);
buf BUF1 (N14671, N14659);
not NOT1 (N14672, N14670);
and AND2 (N14673, N14672, N9123);
and AND4 (N14674, N14665, N12919, N9271, N4291);
not NOT1 (N14675, N14651);
and AND3 (N14676, N14664, N12765, N12164);
or OR4 (N14677, N14671, N9665, N9108, N2419);
nor NOR2 (N14678, N14677, N6727);
xor XOR2 (N14679, N14667, N463);
buf BUF1 (N14680, N14675);
and AND4 (N14681, N14668, N13074, N3885, N3923);
buf BUF1 (N14682, N14626);
or OR3 (N14683, N14678, N1798, N14143);
or OR2 (N14684, N14680, N995);
and AND2 (N14685, N14684, N211);
and AND3 (N14686, N14663, N3893, N4237);
buf BUF1 (N14687, N14686);
nor NOR2 (N14688, N14685, N6055);
xor XOR2 (N14689, N14683, N4939);
xor XOR2 (N14690, N14682, N9784);
xor XOR2 (N14691, N14681, N11389);
xor XOR2 (N14692, N14676, N11625);
or OR2 (N14693, N14692, N11738);
or OR4 (N14694, N14687, N6388, N979, N10579);
buf BUF1 (N14695, N14688);
xor XOR2 (N14696, N14693, N4807);
nor NOR2 (N14697, N14689, N6713);
or OR2 (N14698, N14691, N4111);
nor NOR2 (N14699, N14697, N6374);
nor NOR3 (N14700, N14696, N1886, N4815);
and AND2 (N14701, N14694, N8032);
nand NAND2 (N14702, N14700, N10610);
not NOT1 (N14703, N14695);
and AND4 (N14704, N14652, N9385, N4412, N2042);
not NOT1 (N14705, N14704);
or OR2 (N14706, N14699, N12323);
and AND4 (N14707, N14690, N12180, N1109, N2332);
and AND3 (N14708, N14707, N294, N12691);
not NOT1 (N14709, N14708);
buf BUF1 (N14710, N14679);
and AND3 (N14711, N14698, N10288, N3848);
nand NAND4 (N14712, N14674, N6846, N2827, N8247);
xor XOR2 (N14713, N14710, N4691);
nand NAND3 (N14714, N14705, N5149, N4777);
not NOT1 (N14715, N14701);
or OR2 (N14716, N14673, N7015);
xor XOR2 (N14717, N14711, N6267);
or OR2 (N14718, N14714, N136);
nor NOR3 (N14719, N14709, N5723, N7944);
nand NAND2 (N14720, N14718, N12707);
nor NOR4 (N14721, N14703, N8491, N6485, N8189);
or OR3 (N14722, N14716, N8804, N13535);
and AND3 (N14723, N14722, N7894, N9150);
xor XOR2 (N14724, N14717, N14155);
nor NOR4 (N14725, N14721, N3063, N6078, N10022);
or OR2 (N14726, N14706, N12600);
nand NAND2 (N14727, N14723, N11173);
not NOT1 (N14728, N14725);
and AND3 (N14729, N14728, N12527, N4019);
and AND3 (N14730, N14712, N12583, N189);
nand NAND4 (N14731, N14730, N6259, N14463, N8129);
buf BUF1 (N14732, N14713);
nor NOR3 (N14733, N14726, N9138, N10191);
nor NOR2 (N14734, N14719, N2301);
xor XOR2 (N14735, N14724, N3181);
nor NOR3 (N14736, N14733, N7512, N11833);
buf BUF1 (N14737, N14735);
nand NAND4 (N14738, N14702, N1845, N1935, N13233);
not NOT1 (N14739, N14737);
xor XOR2 (N14740, N14739, N3698);
or OR3 (N14741, N14727, N13124, N10916);
nand NAND4 (N14742, N14741, N5586, N8327, N7554);
nor NOR3 (N14743, N14738, N8853, N10875);
nor NOR3 (N14744, N14729, N8953, N13733);
not NOT1 (N14745, N14731);
xor XOR2 (N14746, N14715, N3289);
not NOT1 (N14747, N14736);
xor XOR2 (N14748, N14732, N10234);
not NOT1 (N14749, N14734);
nand NAND2 (N14750, N14740, N5750);
xor XOR2 (N14751, N14744, N12589);
xor XOR2 (N14752, N14745, N5417);
not NOT1 (N14753, N14750);
xor XOR2 (N14754, N14746, N1230);
nor NOR3 (N14755, N14754, N4100, N5028);
not NOT1 (N14756, N14751);
or OR2 (N14757, N14742, N10760);
nand NAND2 (N14758, N14757, N10202);
nand NAND3 (N14759, N14753, N2869, N14565);
nand NAND3 (N14760, N14758, N9882, N209);
xor XOR2 (N14761, N14759, N1310);
xor XOR2 (N14762, N14720, N11484);
nand NAND2 (N14763, N14743, N3259);
buf BUF1 (N14764, N14760);
nand NAND3 (N14765, N14747, N4351, N9065);
or OR4 (N14766, N14765, N5527, N6897, N8481);
nand NAND4 (N14767, N14762, N703, N12784, N8549);
or OR3 (N14768, N14761, N13117, N383);
xor XOR2 (N14769, N14755, N4666);
and AND2 (N14770, N14749, N12778);
nand NAND3 (N14771, N14752, N5126, N11608);
nand NAND4 (N14772, N14769, N6949, N3566, N13391);
or OR2 (N14773, N14770, N10915);
and AND2 (N14774, N14767, N12422);
nand NAND2 (N14775, N14764, N13082);
nand NAND4 (N14776, N14772, N4765, N8554, N13167);
buf BUF1 (N14777, N14756);
not NOT1 (N14778, N14763);
not NOT1 (N14779, N14748);
not NOT1 (N14780, N14778);
xor XOR2 (N14781, N14771, N11736);
and AND2 (N14782, N14766, N3512);
nand NAND3 (N14783, N14776, N14317, N1933);
or OR4 (N14784, N14783, N10604, N6213, N9276);
nand NAND4 (N14785, N14780, N5499, N5212, N8668);
nand NAND3 (N14786, N14768, N9888, N14458);
buf BUF1 (N14787, N14779);
or OR4 (N14788, N14775, N2282, N5541, N1066);
nor NOR2 (N14789, N14777, N2594);
nand NAND3 (N14790, N14786, N2394, N12378);
buf BUF1 (N14791, N14790);
not NOT1 (N14792, N14787);
and AND2 (N14793, N14782, N4181);
and AND2 (N14794, N14788, N5958);
nor NOR4 (N14795, N14792, N13061, N218, N4160);
nor NOR2 (N14796, N14773, N1650);
not NOT1 (N14797, N14785);
nand NAND3 (N14798, N14794, N12866, N6101);
and AND4 (N14799, N14796, N916, N8489, N84);
buf BUF1 (N14800, N14781);
buf BUF1 (N14801, N14774);
nor NOR3 (N14802, N14795, N5108, N13166);
not NOT1 (N14803, N14784);
or OR4 (N14804, N14800, N4360, N10020, N3564);
and AND3 (N14805, N14793, N2951, N8169);
and AND4 (N14806, N14791, N6457, N11804, N6834);
nor NOR3 (N14807, N14801, N279, N9250);
nand NAND3 (N14808, N14807, N6501, N4863);
nand NAND2 (N14809, N14798, N5621);
not NOT1 (N14810, N14799);
buf BUF1 (N14811, N14802);
nor NOR4 (N14812, N14811, N559, N574, N1431);
buf BUF1 (N14813, N14803);
xor XOR2 (N14814, N14813, N2007);
buf BUF1 (N14815, N14797);
nor NOR2 (N14816, N14789, N6156);
xor XOR2 (N14817, N14806, N8187);
nand NAND3 (N14818, N14815, N1914, N7180);
not NOT1 (N14819, N14804);
nand NAND2 (N14820, N14818, N10227);
buf BUF1 (N14821, N14808);
xor XOR2 (N14822, N14817, N6141);
buf BUF1 (N14823, N14812);
buf BUF1 (N14824, N14816);
xor XOR2 (N14825, N14819, N8020);
or OR3 (N14826, N14822, N1539, N5036);
or OR3 (N14827, N14814, N14023, N7571);
or OR3 (N14828, N14824, N2170, N11382);
xor XOR2 (N14829, N14810, N5915);
or OR3 (N14830, N14826, N3203, N6212);
not NOT1 (N14831, N14809);
buf BUF1 (N14832, N14829);
buf BUF1 (N14833, N14823);
not NOT1 (N14834, N14825);
not NOT1 (N14835, N14820);
or OR2 (N14836, N14827, N1012);
buf BUF1 (N14837, N14821);
buf BUF1 (N14838, N14834);
xor XOR2 (N14839, N14837, N11604);
nand NAND3 (N14840, N14838, N13957, N6533);
and AND2 (N14841, N14839, N3822);
not NOT1 (N14842, N14830);
buf BUF1 (N14843, N14831);
nor NOR3 (N14844, N14842, N4146, N2701);
not NOT1 (N14845, N14835);
nor NOR2 (N14846, N14841, N3896);
and AND3 (N14847, N14843, N3248, N10175);
xor XOR2 (N14848, N14846, N14262);
and AND3 (N14849, N14836, N717, N12222);
not NOT1 (N14850, N14845);
nor NOR2 (N14851, N14844, N14312);
not NOT1 (N14852, N14849);
and AND4 (N14853, N14851, N7699, N7593, N9906);
not NOT1 (N14854, N14848);
xor XOR2 (N14855, N14852, N4536);
nand NAND2 (N14856, N14828, N13401);
buf BUF1 (N14857, N14840);
and AND3 (N14858, N14857, N5248, N4501);
xor XOR2 (N14859, N14854, N1123);
xor XOR2 (N14860, N14805, N6027);
and AND4 (N14861, N14833, N2804, N10243, N12321);
and AND2 (N14862, N14860, N111);
nor NOR4 (N14863, N14855, N13654, N1024, N8531);
nand NAND2 (N14864, N14858, N6442);
nor NOR3 (N14865, N14856, N10823, N11417);
xor XOR2 (N14866, N14859, N8692);
nand NAND2 (N14867, N14866, N12060);
and AND2 (N14868, N14850, N7737);
not NOT1 (N14869, N14832);
or OR2 (N14870, N14861, N688);
nor NOR3 (N14871, N14868, N13942, N5842);
and AND2 (N14872, N14862, N11647);
buf BUF1 (N14873, N14865);
buf BUF1 (N14874, N14864);
nand NAND2 (N14875, N14847, N12293);
and AND4 (N14876, N14863, N9384, N3803, N6185);
nor NOR2 (N14877, N14867, N4874);
xor XOR2 (N14878, N14872, N3017);
or OR3 (N14879, N14877, N13647, N4588);
xor XOR2 (N14880, N14874, N5708);
or OR3 (N14881, N14880, N13168, N3779);
buf BUF1 (N14882, N14869);
nor NOR4 (N14883, N14876, N4998, N7773, N14752);
not NOT1 (N14884, N14881);
buf BUF1 (N14885, N14882);
and AND3 (N14886, N14884, N2988, N6828);
nand NAND3 (N14887, N14875, N1330, N13438);
nand NAND3 (N14888, N14887, N10960, N5524);
nand NAND3 (N14889, N14873, N1566, N6989);
and AND2 (N14890, N14879, N6989);
buf BUF1 (N14891, N14888);
xor XOR2 (N14892, N14886, N880);
nor NOR2 (N14893, N14889, N8849);
not NOT1 (N14894, N14892);
nand NAND4 (N14895, N14890, N1849, N3163, N10791);
buf BUF1 (N14896, N14891);
or OR3 (N14897, N14894, N2550, N9388);
not NOT1 (N14898, N14885);
not NOT1 (N14899, N14893);
and AND4 (N14900, N14899, N8420, N7873, N12282);
nor NOR4 (N14901, N14896, N2271, N2529, N709);
not NOT1 (N14902, N14878);
nand NAND2 (N14903, N14901, N10896);
nor NOR4 (N14904, N14898, N7258, N4068, N848);
nand NAND2 (N14905, N14904, N12536);
nand NAND2 (N14906, N14903, N3013);
not NOT1 (N14907, N14897);
and AND2 (N14908, N14870, N5990);
not NOT1 (N14909, N14908);
and AND4 (N14910, N14871, N2017, N2934, N7034);
nor NOR4 (N14911, N14902, N5175, N5227, N3118);
and AND4 (N14912, N14895, N7047, N2281, N1769);
buf BUF1 (N14913, N14906);
xor XOR2 (N14914, N14883, N476);
and AND3 (N14915, N14900, N14686, N11862);
nand NAND2 (N14916, N14914, N4069);
not NOT1 (N14917, N14853);
and AND3 (N14918, N14916, N3963, N66);
xor XOR2 (N14919, N14913, N1699);
not NOT1 (N14920, N14917);
and AND3 (N14921, N14919, N836, N4337);
or OR2 (N14922, N14918, N2099);
not NOT1 (N14923, N14921);
or OR3 (N14924, N14907, N11122, N2126);
or OR3 (N14925, N14920, N824, N13969);
xor XOR2 (N14926, N14910, N12027);
or OR3 (N14927, N14909, N14806, N8989);
not NOT1 (N14928, N14926);
and AND2 (N14929, N14923, N12362);
xor XOR2 (N14930, N14911, N10719);
xor XOR2 (N14931, N14930, N14849);
xor XOR2 (N14932, N14925, N5900);
and AND4 (N14933, N14924, N2165, N10029, N11651);
not NOT1 (N14934, N14933);
nand NAND3 (N14935, N14922, N6486, N9236);
or OR2 (N14936, N14915, N11602);
or OR2 (N14937, N14912, N4488);
nand NAND2 (N14938, N14928, N13176);
buf BUF1 (N14939, N14936);
and AND3 (N14940, N14935, N1888, N12107);
buf BUF1 (N14941, N14934);
nor NOR2 (N14942, N14941, N10058);
xor XOR2 (N14943, N14905, N6971);
nor NOR4 (N14944, N14932, N1917, N3822, N951);
not NOT1 (N14945, N14937);
nand NAND3 (N14946, N14938, N8789, N4954);
nand NAND4 (N14947, N14939, N7235, N12186, N5248);
and AND4 (N14948, N14946, N10940, N4549, N3452);
buf BUF1 (N14949, N14947);
or OR2 (N14950, N14942, N14787);
or OR2 (N14951, N14949, N484);
not NOT1 (N14952, N14950);
or OR3 (N14953, N14944, N11355, N14929);
xor XOR2 (N14954, N7124, N14523);
xor XOR2 (N14955, N14948, N12122);
and AND3 (N14956, N14954, N13840, N11162);
xor XOR2 (N14957, N14940, N3432);
nor NOR3 (N14958, N14951, N4690, N1211);
buf BUF1 (N14959, N14955);
xor XOR2 (N14960, N14931, N11610);
nand NAND2 (N14961, N14927, N2212);
buf BUF1 (N14962, N14952);
buf BUF1 (N14963, N14959);
nor NOR4 (N14964, N14956, N6274, N4026, N7606);
xor XOR2 (N14965, N14953, N14004);
nor NOR3 (N14966, N14957, N9970, N13069);
or OR4 (N14967, N14961, N11171, N2483, N12862);
or OR4 (N14968, N14963, N8999, N4882, N2764);
xor XOR2 (N14969, N14960, N6281);
xor XOR2 (N14970, N14967, N6459);
or OR2 (N14971, N14943, N9726);
nand NAND4 (N14972, N14970, N5161, N8381, N10789);
or OR2 (N14973, N14969, N9331);
xor XOR2 (N14974, N14964, N2387);
not NOT1 (N14975, N14958);
nor NOR3 (N14976, N14965, N11122, N5858);
xor XOR2 (N14977, N14968, N12278);
xor XOR2 (N14978, N14977, N6137);
not NOT1 (N14979, N14978);
buf BUF1 (N14980, N14945);
xor XOR2 (N14981, N14972, N7700);
and AND3 (N14982, N14973, N10469, N3038);
not NOT1 (N14983, N14979);
and AND2 (N14984, N14971, N3469);
xor XOR2 (N14985, N14974, N7576);
and AND2 (N14986, N14985, N1275);
nand NAND2 (N14987, N14976, N11770);
buf BUF1 (N14988, N14966);
xor XOR2 (N14989, N14988, N13892);
and AND3 (N14990, N14983, N7680, N8369);
xor XOR2 (N14991, N14986, N4948);
and AND2 (N14992, N14962, N2343);
and AND2 (N14993, N14982, N10068);
nor NOR3 (N14994, N14987, N8442, N10168);
and AND4 (N14995, N14992, N5864, N10443, N11450);
and AND3 (N14996, N14980, N7429, N10069);
not NOT1 (N14997, N14981);
and AND4 (N14998, N14995, N6510, N2211, N11099);
or OR4 (N14999, N14993, N5285, N409, N2857);
nand NAND4 (N15000, N14997, N6832, N2917, N7564);
nor NOR3 (N15001, N15000, N9871, N1248);
nand NAND4 (N15002, N14991, N166, N5253, N12666);
or OR2 (N15003, N14996, N10399);
nand NAND2 (N15004, N14989, N9815);
nor NOR3 (N15005, N14994, N7092, N5449);
xor XOR2 (N15006, N14998, N1664);
nor NOR3 (N15007, N15004, N14518, N2921);
nand NAND2 (N15008, N15005, N11305);
xor XOR2 (N15009, N15008, N4259);
nor NOR2 (N15010, N14975, N8821);
xor XOR2 (N15011, N15003, N1022);
not NOT1 (N15012, N15001);
or OR4 (N15013, N15007, N13017, N8845, N5511);
and AND4 (N15014, N15009, N11777, N13207, N9281);
buf BUF1 (N15015, N14984);
nor NOR2 (N15016, N15015, N6166);
and AND2 (N15017, N15012, N13204);
or OR4 (N15018, N15017, N14102, N12708, N10887);
or OR4 (N15019, N15002, N6572, N1871, N4262);
nand NAND4 (N15020, N14990, N12146, N12424, N306);
nor NOR3 (N15021, N15006, N3247, N2250);
xor XOR2 (N15022, N15014, N8737);
nor NOR3 (N15023, N14999, N1271, N6067);
and AND2 (N15024, N15013, N7440);
xor XOR2 (N15025, N15020, N14834);
not NOT1 (N15026, N15016);
nand NAND2 (N15027, N15021, N9948);
not NOT1 (N15028, N15024);
nor NOR4 (N15029, N15019, N6978, N12567, N1247);
nand NAND4 (N15030, N15027, N1841, N12751, N8323);
buf BUF1 (N15031, N15029);
buf BUF1 (N15032, N15011);
and AND4 (N15033, N15018, N14090, N9166, N14942);
buf BUF1 (N15034, N15026);
nor NOR4 (N15035, N15025, N7455, N797, N130);
and AND4 (N15036, N15030, N9116, N843, N2529);
xor XOR2 (N15037, N15033, N7704);
not NOT1 (N15038, N15035);
nor NOR3 (N15039, N15023, N14553, N13932);
and AND4 (N15040, N15022, N11054, N1680, N289);
and AND4 (N15041, N15032, N771, N2550, N12188);
nor NOR3 (N15042, N15028, N10337, N7067);
or OR2 (N15043, N15040, N6241);
xor XOR2 (N15044, N15041, N12483);
and AND3 (N15045, N15010, N12886, N8516);
and AND3 (N15046, N15036, N13940, N10457);
buf BUF1 (N15047, N15044);
not NOT1 (N15048, N15042);
and AND4 (N15049, N15046, N5645, N7533, N12910);
buf BUF1 (N15050, N15039);
xor XOR2 (N15051, N15043, N75);
not NOT1 (N15052, N15050);
nand NAND4 (N15053, N15045, N8384, N9435, N12122);
nor NOR4 (N15054, N15034, N4060, N8004, N5897);
and AND2 (N15055, N15049, N14841);
and AND3 (N15056, N15047, N14758, N2462);
buf BUF1 (N15057, N15056);
buf BUF1 (N15058, N15053);
not NOT1 (N15059, N15038);
nor NOR2 (N15060, N15031, N1819);
nand NAND4 (N15061, N15048, N5094, N839, N9593);
xor XOR2 (N15062, N15055, N7936);
buf BUF1 (N15063, N15037);
or OR2 (N15064, N15061, N6245);
not NOT1 (N15065, N15064);
nand NAND4 (N15066, N15060, N4985, N6342, N6821);
nand NAND4 (N15067, N15052, N6189, N7270, N9959);
nand NAND4 (N15068, N15057, N3036, N8138, N10627);
not NOT1 (N15069, N15062);
nor NOR2 (N15070, N15068, N2928);
nand NAND2 (N15071, N15069, N1095);
not NOT1 (N15072, N15051);
nor NOR2 (N15073, N15063, N12794);
nand NAND4 (N15074, N15070, N12233, N11486, N513);
xor XOR2 (N15075, N15058, N4790);
nor NOR4 (N15076, N15065, N9670, N8094, N6476);
not NOT1 (N15077, N15073);
buf BUF1 (N15078, N15076);
buf BUF1 (N15079, N15072);
nor NOR4 (N15080, N15074, N9620, N12188, N11443);
not NOT1 (N15081, N15075);
xor XOR2 (N15082, N15054, N14122);
and AND4 (N15083, N15080, N3582, N7780, N4799);
not NOT1 (N15084, N15059);
not NOT1 (N15085, N15077);
nor NOR4 (N15086, N15082, N5274, N13170, N13501);
nand NAND3 (N15087, N15078, N7704, N7058);
or OR4 (N15088, N15081, N8995, N14541, N12620);
or OR3 (N15089, N15079, N14940, N1972);
nand NAND3 (N15090, N15071, N10444, N13643);
xor XOR2 (N15091, N15090, N1817);
nor NOR3 (N15092, N15086, N487, N3007);
and AND2 (N15093, N15067, N261);
xor XOR2 (N15094, N15088, N8879);
buf BUF1 (N15095, N15094);
buf BUF1 (N15096, N15087);
not NOT1 (N15097, N15095);
nor NOR3 (N15098, N15084, N6341, N6120);
not NOT1 (N15099, N15066);
buf BUF1 (N15100, N15089);
or OR3 (N15101, N15098, N257, N10093);
nor NOR3 (N15102, N15085, N9999, N10879);
nand NAND2 (N15103, N15100, N14890);
and AND2 (N15104, N15099, N14806);
nand NAND4 (N15105, N15097, N14401, N4448, N3686);
or OR3 (N15106, N15093, N3272, N9716);
xor XOR2 (N15107, N15103, N4675);
and AND3 (N15108, N15106, N4254, N699);
not NOT1 (N15109, N15092);
or OR3 (N15110, N15109, N341, N9708);
nand NAND3 (N15111, N15104, N3614, N1257);
or OR2 (N15112, N15107, N4603);
xor XOR2 (N15113, N15105, N12631);
nand NAND4 (N15114, N15108, N4680, N7733, N13741);
nand NAND2 (N15115, N15102, N7910);
not NOT1 (N15116, N15110);
or OR2 (N15117, N15111, N5372);
nor NOR4 (N15118, N15116, N9172, N10052, N9419);
xor XOR2 (N15119, N15091, N13542);
not NOT1 (N15120, N15113);
buf BUF1 (N15121, N15120);
xor XOR2 (N15122, N15096, N11995);
nor NOR4 (N15123, N15101, N6747, N11709, N10451);
or OR2 (N15124, N15114, N3298);
not NOT1 (N15125, N15115);
or OR2 (N15126, N15125, N4512);
and AND4 (N15127, N15121, N3875, N8365, N12973);
nand NAND4 (N15128, N15112, N14972, N6460, N6636);
xor XOR2 (N15129, N15118, N11187);
xor XOR2 (N15130, N15123, N4590);
xor XOR2 (N15131, N15124, N5719);
and AND4 (N15132, N15117, N3810, N12035, N4344);
nand NAND3 (N15133, N15128, N12741, N1856);
nor NOR3 (N15134, N15119, N3338, N4747);
not NOT1 (N15135, N15133);
not NOT1 (N15136, N15134);
or OR3 (N15137, N15129, N4198, N5481);
or OR3 (N15138, N15127, N4326, N7650);
buf BUF1 (N15139, N15132);
nor NOR2 (N15140, N15135, N8257);
not NOT1 (N15141, N15122);
and AND2 (N15142, N15139, N13623);
or OR3 (N15143, N15140, N6296, N9522);
xor XOR2 (N15144, N15143, N14760);
and AND2 (N15145, N15130, N8349);
and AND4 (N15146, N15131, N14262, N1374, N7086);
buf BUF1 (N15147, N15126);
not NOT1 (N15148, N15136);
nor NOR4 (N15149, N15144, N14000, N11546, N14136);
not NOT1 (N15150, N15138);
nor NOR2 (N15151, N15137, N829);
not NOT1 (N15152, N15149);
not NOT1 (N15153, N15146);
nand NAND3 (N15154, N15145, N12704, N4040);
buf BUF1 (N15155, N15142);
buf BUF1 (N15156, N15150);
not NOT1 (N15157, N15153);
not NOT1 (N15158, N15083);
or OR2 (N15159, N15152, N2839);
buf BUF1 (N15160, N15157);
nor NOR4 (N15161, N15156, N8626, N6775, N3683);
nand NAND3 (N15162, N15160, N9960, N3068);
and AND4 (N15163, N15151, N12041, N1342, N14302);
not NOT1 (N15164, N15141);
buf BUF1 (N15165, N15159);
and AND4 (N15166, N15148, N8283, N8967, N6116);
and AND3 (N15167, N15147, N3244, N6074);
buf BUF1 (N15168, N15155);
or OR4 (N15169, N15162, N5714, N1977, N13970);
buf BUF1 (N15170, N15164);
xor XOR2 (N15171, N15169, N10745);
buf BUF1 (N15172, N15154);
or OR3 (N15173, N15166, N9357, N7758);
not NOT1 (N15174, N15167);
buf BUF1 (N15175, N15172);
xor XOR2 (N15176, N15171, N5431);
or OR2 (N15177, N15176, N9721);
nand NAND4 (N15178, N15174, N7820, N8370, N8446);
not NOT1 (N15179, N15165);
nor NOR3 (N15180, N15163, N14345, N8931);
not NOT1 (N15181, N15161);
or OR3 (N15182, N15158, N13315, N7505);
xor XOR2 (N15183, N15175, N8077);
and AND4 (N15184, N15173, N3513, N9587, N11207);
or OR4 (N15185, N15170, N11670, N9380, N8322);
and AND4 (N15186, N15180, N14911, N1183, N557);
or OR4 (N15187, N15185, N2841, N12782, N6715);
and AND3 (N15188, N15168, N7688, N11524);
xor XOR2 (N15189, N15179, N5877);
nand NAND4 (N15190, N15184, N12221, N11124, N14363);
nor NOR3 (N15191, N15178, N12897, N4656);
xor XOR2 (N15192, N15187, N4061);
nor NOR2 (N15193, N15189, N12945);
buf BUF1 (N15194, N15191);
or OR3 (N15195, N15181, N1672, N1928);
nand NAND2 (N15196, N15177, N1024);
not NOT1 (N15197, N15195);
not NOT1 (N15198, N15194);
nand NAND2 (N15199, N15186, N10722);
buf BUF1 (N15200, N15188);
or OR4 (N15201, N15200, N9697, N10276, N14449);
and AND4 (N15202, N15196, N6274, N11009, N6563);
or OR3 (N15203, N15199, N1946, N9918);
or OR3 (N15204, N15198, N829, N10882);
xor XOR2 (N15205, N15197, N362);
not NOT1 (N15206, N15204);
xor XOR2 (N15207, N15190, N1327);
nor NOR3 (N15208, N15183, N15047, N6896);
xor XOR2 (N15209, N15205, N14212);
buf BUF1 (N15210, N15208);
not NOT1 (N15211, N15182);
and AND3 (N15212, N15192, N9096, N11180);
not NOT1 (N15213, N15210);
not NOT1 (N15214, N15202);
and AND4 (N15215, N15207, N3000, N5848, N5434);
xor XOR2 (N15216, N15193, N2526);
nor NOR3 (N15217, N15206, N9239, N5180);
not NOT1 (N15218, N15213);
and AND2 (N15219, N15203, N10885);
or OR3 (N15220, N15214, N12062, N12099);
or OR3 (N15221, N15209, N10397, N27);
nand NAND4 (N15222, N15212, N2833, N9970, N6213);
not NOT1 (N15223, N15219);
not NOT1 (N15224, N15215);
nand NAND4 (N15225, N15217, N10844, N5536, N3346);
xor XOR2 (N15226, N15223, N4783);
not NOT1 (N15227, N15218);
buf BUF1 (N15228, N15226);
xor XOR2 (N15229, N15201, N11028);
nor NOR4 (N15230, N15211, N2084, N13482, N3068);
not NOT1 (N15231, N15222);
and AND4 (N15232, N15227, N14756, N12751, N1626);
or OR2 (N15233, N15224, N184);
or OR3 (N15234, N15230, N3000, N4317);
buf BUF1 (N15235, N15234);
or OR2 (N15236, N15225, N30);
or OR3 (N15237, N15236, N9113, N6786);
or OR3 (N15238, N15233, N7740, N14407);
or OR2 (N15239, N15231, N11586);
and AND3 (N15240, N15220, N9682, N4622);
not NOT1 (N15241, N15216);
nor NOR3 (N15242, N15239, N8473, N683);
or OR4 (N15243, N15228, N14118, N6745, N4139);
buf BUF1 (N15244, N15242);
not NOT1 (N15245, N15240);
or OR3 (N15246, N15232, N519, N14007);
nor NOR3 (N15247, N15241, N2071, N11747);
nand NAND4 (N15248, N15247, N9061, N12735, N14628);
nand NAND2 (N15249, N15221, N10422);
nor NOR4 (N15250, N15238, N10680, N9461, N9773);
xor XOR2 (N15251, N15235, N4246);
or OR3 (N15252, N15248, N11585, N4316);
nand NAND3 (N15253, N15251, N109, N14174);
not NOT1 (N15254, N15246);
and AND4 (N15255, N15244, N3566, N7399, N9427);
nor NOR3 (N15256, N15250, N9467, N2875);
nor NOR3 (N15257, N15243, N11954, N4683);
xor XOR2 (N15258, N15252, N11124);
not NOT1 (N15259, N15254);
nor NOR4 (N15260, N15257, N6464, N711, N1536);
not NOT1 (N15261, N15260);
nand NAND4 (N15262, N15258, N8259, N8513, N11420);
nor NOR4 (N15263, N15229, N7336, N8556, N4258);
not NOT1 (N15264, N15249);
buf BUF1 (N15265, N15261);
buf BUF1 (N15266, N15245);
or OR2 (N15267, N15264, N8712);
buf BUF1 (N15268, N15253);
xor XOR2 (N15269, N15237, N3375);
xor XOR2 (N15270, N15262, N12699);
and AND3 (N15271, N15266, N15133, N3639);
nor NOR2 (N15272, N15259, N7776);
nor NOR3 (N15273, N15271, N3995, N7954);
xor XOR2 (N15274, N15265, N13497);
and AND4 (N15275, N15256, N5350, N7703, N12866);
nor NOR2 (N15276, N15275, N10823);
or OR4 (N15277, N15274, N13204, N15242, N6725);
or OR3 (N15278, N15277, N2167, N12975);
buf BUF1 (N15279, N15273);
not NOT1 (N15280, N15272);
xor XOR2 (N15281, N15268, N10119);
and AND2 (N15282, N15276, N6282);
not NOT1 (N15283, N15267);
buf BUF1 (N15284, N15255);
xor XOR2 (N15285, N15280, N14813);
not NOT1 (N15286, N15279);
and AND4 (N15287, N15285, N5479, N13460, N10159);
and AND2 (N15288, N15287, N290);
nand NAND4 (N15289, N15281, N14037, N11618, N13725);
buf BUF1 (N15290, N15263);
and AND2 (N15291, N15270, N9257);
xor XOR2 (N15292, N15291, N1590);
nand NAND4 (N15293, N15290, N2939, N6195, N364);
buf BUF1 (N15294, N15293);
nand NAND3 (N15295, N15283, N4806, N4577);
nor NOR2 (N15296, N15286, N9766);
nand NAND4 (N15297, N15296, N2627, N5250, N13303);
and AND2 (N15298, N15294, N6213);
buf BUF1 (N15299, N15278);
and AND4 (N15300, N15299, N10197, N8164, N1867);
or OR3 (N15301, N15292, N3078, N1553);
buf BUF1 (N15302, N15284);
or OR4 (N15303, N15282, N3168, N5167, N9705);
not NOT1 (N15304, N15302);
buf BUF1 (N15305, N15298);
or OR4 (N15306, N15305, N8021, N4313, N11351);
buf BUF1 (N15307, N15288);
not NOT1 (N15308, N15289);
nor NOR2 (N15309, N15301, N7873);
xor XOR2 (N15310, N15309, N11502);
or OR2 (N15311, N15297, N6753);
xor XOR2 (N15312, N15295, N8362);
xor XOR2 (N15313, N15303, N5601);
nor NOR2 (N15314, N15313, N269);
not NOT1 (N15315, N15310);
nor NOR4 (N15316, N15300, N3235, N3294, N1665);
and AND3 (N15317, N15307, N5435, N2914);
or OR2 (N15318, N15308, N1085);
buf BUF1 (N15319, N15306);
nor NOR4 (N15320, N15316, N8472, N7408, N8524);
nor NOR4 (N15321, N15315, N1969, N9981, N7510);
xor XOR2 (N15322, N15318, N440);
buf BUF1 (N15323, N15304);
or OR2 (N15324, N15312, N14660);
and AND2 (N15325, N15319, N1355);
buf BUF1 (N15326, N15325);
buf BUF1 (N15327, N15321);
not NOT1 (N15328, N15311);
nor NOR2 (N15329, N15326, N158);
nor NOR2 (N15330, N15327, N13834);
and AND2 (N15331, N15324, N8831);
nand NAND4 (N15332, N15330, N12165, N12096, N10788);
and AND3 (N15333, N15320, N14875, N9868);
or OR3 (N15334, N15331, N14543, N10191);
and AND2 (N15335, N15269, N4317);
or OR4 (N15336, N15329, N3474, N13794, N6441);
not NOT1 (N15337, N15317);
xor XOR2 (N15338, N15332, N11212);
xor XOR2 (N15339, N15323, N10716);
not NOT1 (N15340, N15338);
and AND2 (N15341, N15328, N8027);
and AND2 (N15342, N15336, N14988);
or OR4 (N15343, N15342, N10274, N5393, N5463);
nand NAND3 (N15344, N15335, N3045, N6317);
or OR4 (N15345, N15339, N4091, N9933, N14165);
or OR4 (N15346, N15337, N5537, N1336, N12944);
or OR3 (N15347, N15344, N1464, N6998);
and AND3 (N15348, N15334, N12625, N2394);
not NOT1 (N15349, N15333);
and AND4 (N15350, N15348, N11268, N11467, N12515);
not NOT1 (N15351, N15340);
or OR2 (N15352, N15351, N13581);
nor NOR2 (N15353, N15346, N7802);
buf BUF1 (N15354, N15314);
nor NOR3 (N15355, N15345, N10940, N9278);
and AND2 (N15356, N15354, N6889);
nand NAND2 (N15357, N15353, N11613);
and AND4 (N15358, N15352, N6434, N7124, N2568);
and AND4 (N15359, N15355, N9347, N8250, N6872);
nor NOR2 (N15360, N15349, N969);
xor XOR2 (N15361, N15343, N623);
not NOT1 (N15362, N15361);
buf BUF1 (N15363, N15347);
nor NOR4 (N15364, N15359, N6333, N8553, N13772);
or OR3 (N15365, N15356, N13745, N8442);
xor XOR2 (N15366, N15363, N10913);
nor NOR3 (N15367, N15360, N4799, N6777);
xor XOR2 (N15368, N15366, N2898);
or OR3 (N15369, N15365, N691, N1318);
or OR4 (N15370, N15362, N14340, N11446, N12380);
not NOT1 (N15371, N15341);
nand NAND2 (N15372, N15358, N13859);
nand NAND2 (N15373, N15371, N14355);
or OR3 (N15374, N15373, N6043, N11600);
nor NOR2 (N15375, N15357, N12152);
nor NOR4 (N15376, N15364, N12389, N12450, N12374);
not NOT1 (N15377, N15375);
nor NOR3 (N15378, N15322, N13799, N6661);
or OR3 (N15379, N15374, N861, N14660);
and AND2 (N15380, N15378, N13855);
or OR3 (N15381, N15376, N10707, N12613);
nor NOR3 (N15382, N15377, N14959, N8177);
and AND3 (N15383, N15372, N1156, N11489);
buf BUF1 (N15384, N15383);
and AND4 (N15385, N15379, N1715, N7100, N14643);
nor NOR3 (N15386, N15382, N15207, N15270);
or OR4 (N15387, N15384, N3879, N13458, N2856);
or OR4 (N15388, N15370, N6474, N2257, N4851);
xor XOR2 (N15389, N15368, N15228);
not NOT1 (N15390, N15380);
not NOT1 (N15391, N15386);
and AND4 (N15392, N15388, N3144, N2422, N4598);
or OR3 (N15393, N15381, N4187, N3926);
buf BUF1 (N15394, N15350);
nor NOR4 (N15395, N15367, N2004, N7804, N7758);
not NOT1 (N15396, N15387);
nor NOR3 (N15397, N15392, N4551, N3121);
or OR4 (N15398, N15369, N5412, N13121, N2115);
buf BUF1 (N15399, N15393);
xor XOR2 (N15400, N15396, N5399);
buf BUF1 (N15401, N15397);
nand NAND2 (N15402, N15395, N10566);
nor NOR3 (N15403, N15400, N13004, N5635);
xor XOR2 (N15404, N15398, N13996);
or OR2 (N15405, N15404, N8664);
not NOT1 (N15406, N15390);
xor XOR2 (N15407, N15406, N1598);
nor NOR2 (N15408, N15405, N6020);
buf BUF1 (N15409, N15391);
xor XOR2 (N15410, N15409, N13351);
xor XOR2 (N15411, N15401, N10691);
xor XOR2 (N15412, N15407, N5962);
xor XOR2 (N15413, N15402, N6745);
nor NOR3 (N15414, N15399, N10219, N13092);
and AND2 (N15415, N15389, N7186);
buf BUF1 (N15416, N15403);
and AND4 (N15417, N15413, N10437, N12836, N7964);
nor NOR2 (N15418, N15411, N2201);
nor NOR4 (N15419, N15415, N72, N6641, N11545);
nor NOR3 (N15420, N15410, N13569, N280);
or OR3 (N15421, N15412, N952, N2368);
buf BUF1 (N15422, N15414);
nand NAND3 (N15423, N15417, N2782, N10717);
buf BUF1 (N15424, N15421);
or OR3 (N15425, N15422, N8484, N11477);
buf BUF1 (N15426, N15420);
buf BUF1 (N15427, N15408);
nor NOR2 (N15428, N15385, N8065);
buf BUF1 (N15429, N15419);
or OR4 (N15430, N15429, N11451, N3201, N8130);
and AND4 (N15431, N15427, N3161, N15031, N831);
xor XOR2 (N15432, N15424, N2206);
nand NAND2 (N15433, N15430, N13183);
nand NAND2 (N15434, N15394, N7006);
nand NAND3 (N15435, N15423, N2653, N10743);
buf BUF1 (N15436, N15418);
or OR4 (N15437, N15428, N4817, N607, N1940);
buf BUF1 (N15438, N15426);
xor XOR2 (N15439, N15433, N4650);
nand NAND3 (N15440, N15439, N10991, N4224);
not NOT1 (N15441, N15434);
or OR3 (N15442, N15432, N13579, N10949);
nand NAND3 (N15443, N15442, N14649, N4931);
and AND4 (N15444, N15435, N11190, N12629, N8000);
not NOT1 (N15445, N15438);
xor XOR2 (N15446, N15436, N3937);
not NOT1 (N15447, N15446);
and AND2 (N15448, N15416, N6256);
xor XOR2 (N15449, N15425, N9944);
and AND2 (N15450, N15441, N12460);
not NOT1 (N15451, N15447);
not NOT1 (N15452, N15449);
not NOT1 (N15453, N15452);
nand NAND4 (N15454, N15443, N8501, N1742, N7186);
and AND4 (N15455, N15450, N1213, N13249, N1543);
nand NAND4 (N15456, N15431, N13071, N3166, N5246);
and AND3 (N15457, N15456, N8660, N9027);
xor XOR2 (N15458, N15455, N10269);
buf BUF1 (N15459, N15457);
buf BUF1 (N15460, N15440);
buf BUF1 (N15461, N15451);
xor XOR2 (N15462, N15437, N5221);
not NOT1 (N15463, N15448);
not NOT1 (N15464, N15459);
buf BUF1 (N15465, N15444);
nor NOR4 (N15466, N15453, N3515, N6362, N2200);
not NOT1 (N15467, N15465);
nor NOR3 (N15468, N15466, N6452, N9718);
and AND2 (N15469, N15468, N6717);
xor XOR2 (N15470, N15458, N399);
buf BUF1 (N15471, N15461);
nor NOR4 (N15472, N15469, N5333, N15068, N5758);
nor NOR3 (N15473, N15467, N11243, N1816);
nor NOR2 (N15474, N15473, N2794);
or OR4 (N15475, N15460, N7523, N10535, N3847);
nand NAND3 (N15476, N15475, N8353, N4551);
xor XOR2 (N15477, N15474, N12738);
nand NAND2 (N15478, N15477, N11738);
nand NAND2 (N15479, N15470, N12251);
not NOT1 (N15480, N15471);
buf BUF1 (N15481, N15445);
nand NAND3 (N15482, N15454, N13493, N6745);
nand NAND3 (N15483, N15478, N2951, N7832);
buf BUF1 (N15484, N15479);
not NOT1 (N15485, N15472);
nand NAND2 (N15486, N15483, N5501);
not NOT1 (N15487, N15462);
nor NOR2 (N15488, N15484, N5530);
or OR4 (N15489, N15486, N10025, N6440, N4589);
or OR3 (N15490, N15481, N2536, N14160);
buf BUF1 (N15491, N15490);
buf BUF1 (N15492, N15476);
xor XOR2 (N15493, N15492, N6426);
or OR2 (N15494, N15489, N6148);
buf BUF1 (N15495, N15482);
not NOT1 (N15496, N15494);
buf BUF1 (N15497, N15495);
not NOT1 (N15498, N15488);
buf BUF1 (N15499, N15487);
nand NAND4 (N15500, N15498, N12624, N11710, N3583);
xor XOR2 (N15501, N15497, N7762);
buf BUF1 (N15502, N15499);
and AND4 (N15503, N15493, N12086, N14865, N14506);
or OR2 (N15504, N15491, N5477);
nand NAND4 (N15505, N15502, N11020, N12905, N6333);
nor NOR3 (N15506, N15500, N15080, N2514);
xor XOR2 (N15507, N15503, N13263);
xor XOR2 (N15508, N15505, N9152);
and AND4 (N15509, N15508, N6339, N12366, N9477);
xor XOR2 (N15510, N15463, N9450);
or OR2 (N15511, N15506, N4082);
xor XOR2 (N15512, N15511, N3157);
nor NOR3 (N15513, N15504, N1492, N10673);
or OR3 (N15514, N15507, N13335, N13910);
not NOT1 (N15515, N15513);
xor XOR2 (N15516, N15514, N7542);
xor XOR2 (N15517, N15501, N14555);
or OR3 (N15518, N15485, N9078, N2355);
not NOT1 (N15519, N15510);
buf BUF1 (N15520, N15512);
xor XOR2 (N15521, N15509, N3410);
and AND2 (N15522, N15496, N5489);
buf BUF1 (N15523, N15464);
xor XOR2 (N15524, N15518, N1131);
nand NAND3 (N15525, N15522, N9033, N4663);
xor XOR2 (N15526, N15521, N12518);
nor NOR2 (N15527, N15520, N10364);
and AND2 (N15528, N15517, N1397);
xor XOR2 (N15529, N15527, N669);
not NOT1 (N15530, N15525);
buf BUF1 (N15531, N15529);
or OR4 (N15532, N15523, N11778, N7123, N7393);
not NOT1 (N15533, N15532);
nand NAND3 (N15534, N15528, N9490, N1161);
nand NAND2 (N15535, N15534, N13904);
nand NAND3 (N15536, N15515, N11881, N2685);
buf BUF1 (N15537, N15536);
buf BUF1 (N15538, N15535);
nand NAND3 (N15539, N15526, N6917, N2248);
and AND4 (N15540, N15480, N5023, N11139, N1562);
nand NAND4 (N15541, N15531, N11888, N3995, N11631);
xor XOR2 (N15542, N15537, N9637);
or OR4 (N15543, N15530, N10261, N10075, N2980);
or OR3 (N15544, N15538, N4220, N15413);
nor NOR3 (N15545, N15516, N10355, N1556);
nor NOR2 (N15546, N15539, N2160);
and AND3 (N15547, N15533, N10354, N1265);
nor NOR2 (N15548, N15542, N11742);
nor NOR3 (N15549, N15543, N9541, N14599);
and AND2 (N15550, N15546, N8883);
or OR3 (N15551, N15519, N9692, N2368);
or OR2 (N15552, N15551, N15117);
and AND2 (N15553, N15545, N295);
buf BUF1 (N15554, N15549);
buf BUF1 (N15555, N15524);
xor XOR2 (N15556, N15540, N14147);
buf BUF1 (N15557, N15544);
not NOT1 (N15558, N15554);
and AND2 (N15559, N15547, N6314);
xor XOR2 (N15560, N15548, N4958);
nand NAND2 (N15561, N15553, N12977);
buf BUF1 (N15562, N15555);
xor XOR2 (N15563, N15558, N4208);
nor NOR3 (N15564, N15561, N12892, N10676);
or OR3 (N15565, N15564, N10174, N8144);
and AND3 (N15566, N15556, N4529, N4084);
nand NAND3 (N15567, N15559, N295, N13759);
nor NOR4 (N15568, N15557, N11364, N13500, N13500);
nor NOR4 (N15569, N15560, N8518, N4310, N4437);
or OR2 (N15570, N15562, N14431);
xor XOR2 (N15571, N15541, N2860);
and AND3 (N15572, N15567, N5621, N1431);
xor XOR2 (N15573, N15552, N450);
nor NOR3 (N15574, N15566, N4756, N1515);
buf BUF1 (N15575, N15550);
xor XOR2 (N15576, N15572, N9603);
nor NOR4 (N15577, N15569, N13078, N158, N15311);
nand NAND2 (N15578, N15570, N13071);
nand NAND2 (N15579, N15565, N10631);
buf BUF1 (N15580, N15578);
buf BUF1 (N15581, N15580);
buf BUF1 (N15582, N15574);
not NOT1 (N15583, N15582);
not NOT1 (N15584, N15571);
nor NOR3 (N15585, N15568, N14610, N14001);
nor NOR2 (N15586, N15575, N5972);
or OR3 (N15587, N15563, N1872, N7879);
buf BUF1 (N15588, N15573);
nand NAND4 (N15589, N15576, N13652, N4032, N14219);
and AND4 (N15590, N15584, N7843, N13024, N9429);
nor NOR4 (N15591, N15589, N7922, N8828, N9555);
nand NAND2 (N15592, N15590, N1515);
xor XOR2 (N15593, N15585, N2370);
not NOT1 (N15594, N15579);
and AND2 (N15595, N15594, N993);
xor XOR2 (N15596, N15593, N7826);
buf BUF1 (N15597, N15577);
nand NAND3 (N15598, N15597, N8681, N7453);
nand NAND3 (N15599, N15596, N12513, N4865);
buf BUF1 (N15600, N15587);
nor NOR2 (N15601, N15581, N12807);
not NOT1 (N15602, N15595);
or OR3 (N15603, N15601, N13329, N10996);
not NOT1 (N15604, N15602);
xor XOR2 (N15605, N15603, N2242);
or OR3 (N15606, N15592, N5618, N6164);
not NOT1 (N15607, N15606);
and AND4 (N15608, N15600, N11775, N13977, N8584);
or OR2 (N15609, N15605, N13014);
xor XOR2 (N15610, N15604, N9337);
xor XOR2 (N15611, N15610, N11657);
not NOT1 (N15612, N15607);
xor XOR2 (N15613, N15591, N1129);
not NOT1 (N15614, N15586);
nand NAND4 (N15615, N15609, N10196, N10019, N8413);
nor NOR3 (N15616, N15612, N11331, N15386);
nor NOR2 (N15617, N15614, N1601);
buf BUF1 (N15618, N15583);
and AND3 (N15619, N15616, N2125, N5814);
buf BUF1 (N15620, N15599);
nand NAND2 (N15621, N15598, N3421);
buf BUF1 (N15622, N15617);
xor XOR2 (N15623, N15588, N3943);
and AND4 (N15624, N15613, N1880, N2996, N10403);
or OR3 (N15625, N15623, N10870, N5674);
buf BUF1 (N15626, N15618);
buf BUF1 (N15627, N15615);
nand NAND2 (N15628, N15624, N3283);
not NOT1 (N15629, N15627);
xor XOR2 (N15630, N15629, N2340);
and AND4 (N15631, N15619, N3316, N9916, N15076);
buf BUF1 (N15632, N15625);
nand NAND3 (N15633, N15621, N15360, N4395);
nand NAND2 (N15634, N15631, N7600);
and AND4 (N15635, N15633, N15487, N5408, N8856);
xor XOR2 (N15636, N15620, N15429);
not NOT1 (N15637, N15635);
or OR2 (N15638, N15634, N2812);
not NOT1 (N15639, N15630);
xor XOR2 (N15640, N15611, N994);
or OR4 (N15641, N15640, N14822, N14193, N14790);
not NOT1 (N15642, N15638);
or OR4 (N15643, N15637, N4997, N11495, N15589);
not NOT1 (N15644, N15608);
nor NOR4 (N15645, N15626, N1812, N10088, N6626);
buf BUF1 (N15646, N15643);
xor XOR2 (N15647, N15645, N12901);
and AND2 (N15648, N15636, N10831);
nor NOR2 (N15649, N15646, N9683);
nand NAND3 (N15650, N15622, N2882, N8769);
not NOT1 (N15651, N15650);
xor XOR2 (N15652, N15649, N10018);
not NOT1 (N15653, N15628);
and AND2 (N15654, N15644, N6140);
nand NAND2 (N15655, N15648, N7077);
xor XOR2 (N15656, N15651, N7997);
and AND2 (N15657, N15641, N9064);
or OR3 (N15658, N15657, N4535, N4434);
nand NAND2 (N15659, N15655, N14394);
or OR3 (N15660, N15642, N1325, N2119);
xor XOR2 (N15661, N15639, N10413);
nor NOR4 (N15662, N15647, N8854, N12285, N10264);
nor NOR3 (N15663, N15659, N14888, N4499);
and AND3 (N15664, N15652, N11463, N9852);
and AND4 (N15665, N15654, N14806, N8628, N7493);
xor XOR2 (N15666, N15664, N5551);
nor NOR3 (N15667, N15663, N14921, N640);
and AND2 (N15668, N15653, N4010);
or OR2 (N15669, N15667, N9239);
not NOT1 (N15670, N15661);
buf BUF1 (N15671, N15670);
xor XOR2 (N15672, N15660, N3224);
nand NAND4 (N15673, N15669, N6553, N12386, N9862);
buf BUF1 (N15674, N15671);
xor XOR2 (N15675, N15674, N11086);
and AND2 (N15676, N15665, N13554);
nor NOR4 (N15677, N15676, N14554, N1067, N10965);
or OR4 (N15678, N15673, N3860, N885, N7545);
or OR3 (N15679, N15656, N13951, N4491);
nor NOR2 (N15680, N15658, N14927);
or OR3 (N15681, N15672, N10416, N2474);
nor NOR4 (N15682, N15681, N10579, N4882, N7495);
and AND2 (N15683, N15632, N11619);
not NOT1 (N15684, N15682);
not NOT1 (N15685, N15683);
and AND2 (N15686, N15678, N6194);
not NOT1 (N15687, N15679);
xor XOR2 (N15688, N15675, N12783);
xor XOR2 (N15689, N15688, N11449);
and AND3 (N15690, N15685, N13928, N7626);
not NOT1 (N15691, N15666);
nor NOR4 (N15692, N15677, N13724, N14096, N656);
or OR3 (N15693, N15691, N8493, N15315);
not NOT1 (N15694, N15662);
and AND3 (N15695, N15668, N5582, N4612);
or OR4 (N15696, N15687, N6661, N2387, N13421);
buf BUF1 (N15697, N15696);
nand NAND3 (N15698, N15694, N10712, N6902);
not NOT1 (N15699, N15689);
xor XOR2 (N15700, N15684, N11566);
and AND2 (N15701, N15680, N12911);
not NOT1 (N15702, N15701);
and AND2 (N15703, N15693, N13816);
xor XOR2 (N15704, N15695, N1711);
nor NOR3 (N15705, N15700, N3035, N3029);
nand NAND3 (N15706, N15686, N4389, N7548);
xor XOR2 (N15707, N15704, N13404);
or OR3 (N15708, N15707, N2988, N2714);
buf BUF1 (N15709, N15705);
nor NOR2 (N15710, N15708, N10718);
and AND2 (N15711, N15692, N531);
or OR3 (N15712, N15690, N15287, N14720);
xor XOR2 (N15713, N15702, N168);
or OR3 (N15714, N15709, N13951, N14457);
or OR3 (N15715, N15699, N14431, N10119);
not NOT1 (N15716, N15706);
and AND2 (N15717, N15712, N8448);
xor XOR2 (N15718, N15713, N3462);
xor XOR2 (N15719, N15711, N6791);
not NOT1 (N15720, N15703);
buf BUF1 (N15721, N15710);
xor XOR2 (N15722, N15697, N2342);
not NOT1 (N15723, N15721);
or OR2 (N15724, N15723, N13628);
and AND2 (N15725, N15715, N5804);
and AND4 (N15726, N15719, N2536, N4639, N10668);
nor NOR3 (N15727, N15722, N12227, N12586);
not NOT1 (N15728, N15717);
or OR4 (N15729, N15728, N10631, N4030, N14387);
xor XOR2 (N15730, N15729, N5229);
or OR3 (N15731, N15730, N2433, N13972);
not NOT1 (N15732, N15718);
or OR3 (N15733, N15716, N4162, N3094);
xor XOR2 (N15734, N15714, N4605);
nor NOR3 (N15735, N15731, N5413, N13728);
not NOT1 (N15736, N15720);
buf BUF1 (N15737, N15735);
or OR2 (N15738, N15726, N4810);
or OR2 (N15739, N15732, N11609);
buf BUF1 (N15740, N15727);
nand NAND3 (N15741, N15736, N13144, N11168);
buf BUF1 (N15742, N15738);
not NOT1 (N15743, N15724);
and AND3 (N15744, N15742, N5153, N6195);
and AND2 (N15745, N15744, N4944);
not NOT1 (N15746, N15737);
xor XOR2 (N15747, N15741, N12370);
nor NOR4 (N15748, N15739, N6983, N344, N2254);
or OR2 (N15749, N15733, N8902);
xor XOR2 (N15750, N15734, N1123);
or OR3 (N15751, N15745, N10153, N2846);
not NOT1 (N15752, N15750);
or OR2 (N15753, N15743, N4408);
or OR2 (N15754, N15740, N3526);
nand NAND4 (N15755, N15754, N3042, N2457, N5762);
buf BUF1 (N15756, N15698);
buf BUF1 (N15757, N15748);
buf BUF1 (N15758, N15757);
buf BUF1 (N15759, N15756);
nand NAND4 (N15760, N15746, N5883, N2201, N7758);
nand NAND4 (N15761, N15747, N4771, N11673, N2846);
buf BUF1 (N15762, N15752);
nand NAND4 (N15763, N15758, N15227, N6910, N1399);
nor NOR3 (N15764, N15759, N4592, N10480);
or OR2 (N15765, N15755, N3631);
or OR3 (N15766, N15765, N10711, N11299);
nand NAND4 (N15767, N15764, N490, N6103, N10146);
buf BUF1 (N15768, N15760);
xor XOR2 (N15769, N15725, N2924);
nor NOR2 (N15770, N15763, N14606);
xor XOR2 (N15771, N15766, N13833);
or OR3 (N15772, N15771, N3447, N347);
not NOT1 (N15773, N15769);
xor XOR2 (N15774, N15768, N15580);
and AND3 (N15775, N15749, N14664, N1347);
nand NAND2 (N15776, N15767, N3828);
and AND2 (N15777, N15776, N15634);
xor XOR2 (N15778, N15751, N15101);
nand NAND3 (N15779, N15753, N6627, N12377);
or OR3 (N15780, N15778, N1791, N11380);
nand NAND2 (N15781, N15780, N8153);
nand NAND3 (N15782, N15772, N11769, N7579);
nand NAND2 (N15783, N15770, N12782);
and AND3 (N15784, N15761, N8869, N13529);
not NOT1 (N15785, N15762);
xor XOR2 (N15786, N15773, N8576);
xor XOR2 (N15787, N15777, N5104);
nor NOR2 (N15788, N15781, N4174);
xor XOR2 (N15789, N15785, N10260);
nor NOR3 (N15790, N15784, N10993, N13930);
buf BUF1 (N15791, N15775);
not NOT1 (N15792, N15779);
nand NAND4 (N15793, N15788, N6886, N2829, N7205);
and AND4 (N15794, N15782, N3337, N14958, N11496);
nand NAND2 (N15795, N15786, N9955);
buf BUF1 (N15796, N15774);
nand NAND2 (N15797, N15796, N8195);
and AND3 (N15798, N15794, N7811, N11724);
xor XOR2 (N15799, N15797, N464);
and AND3 (N15800, N15795, N8011, N3104);
nor NOR3 (N15801, N15798, N13716, N15194);
not NOT1 (N15802, N15789);
or OR2 (N15803, N15793, N12300);
nor NOR2 (N15804, N15799, N220);
and AND4 (N15805, N15783, N12682, N5033, N7175);
xor XOR2 (N15806, N15800, N4287);
buf BUF1 (N15807, N15791);
not NOT1 (N15808, N15807);
xor XOR2 (N15809, N15802, N7769);
xor XOR2 (N15810, N15809, N12764);
or OR3 (N15811, N15806, N4882, N4586);
not NOT1 (N15812, N15810);
or OR3 (N15813, N15804, N6531, N5359);
or OR4 (N15814, N15801, N4561, N9942, N4102);
nand NAND2 (N15815, N15805, N3818);
not NOT1 (N15816, N15814);
buf BUF1 (N15817, N15803);
or OR4 (N15818, N15812, N15265, N7591, N1900);
buf BUF1 (N15819, N15790);
xor XOR2 (N15820, N15808, N11276);
not NOT1 (N15821, N15813);
nor NOR2 (N15822, N15819, N6904);
not NOT1 (N15823, N15787);
xor XOR2 (N15824, N15821, N10367);
or OR4 (N15825, N15816, N6816, N5548, N14508);
buf BUF1 (N15826, N15818);
nand NAND2 (N15827, N15817, N14584);
or OR2 (N15828, N15822, N13011);
nor NOR3 (N15829, N15827, N5795, N1468);
xor XOR2 (N15830, N15792, N8842);
buf BUF1 (N15831, N15811);
xor XOR2 (N15832, N15830, N783);
or OR4 (N15833, N15826, N5372, N8491, N7896);
and AND2 (N15834, N15823, N8250);
and AND4 (N15835, N15824, N14898, N10077, N9435);
nand NAND2 (N15836, N15832, N2956);
and AND2 (N15837, N15831, N10609);
not NOT1 (N15838, N15815);
or OR3 (N15839, N15835, N11850, N10613);
and AND3 (N15840, N15820, N2355, N8305);
nand NAND3 (N15841, N15837, N10949, N11240);
xor XOR2 (N15842, N15838, N9700);
nand NAND2 (N15843, N15841, N8991);
or OR2 (N15844, N15829, N11691);
nand NAND3 (N15845, N15844, N7955, N8918);
xor XOR2 (N15846, N15839, N2262);
xor XOR2 (N15847, N15833, N14140);
not NOT1 (N15848, N15847);
nor NOR2 (N15849, N15825, N8070);
xor XOR2 (N15850, N15843, N11875);
not NOT1 (N15851, N15849);
and AND3 (N15852, N15828, N8028, N3889);
xor XOR2 (N15853, N15842, N14585);
nor NOR3 (N15854, N15840, N9323, N8805);
or OR3 (N15855, N15834, N2922, N7202);
xor XOR2 (N15856, N15836, N15493);
not NOT1 (N15857, N15848);
nand NAND3 (N15858, N15857, N15113, N15410);
xor XOR2 (N15859, N15853, N14532);
buf BUF1 (N15860, N15854);
buf BUF1 (N15861, N15855);
xor XOR2 (N15862, N15852, N3090);
buf BUF1 (N15863, N15856);
nand NAND3 (N15864, N15862, N1946, N4462);
nor NOR2 (N15865, N15863, N10162);
or OR3 (N15866, N15864, N1825, N882);
not NOT1 (N15867, N15845);
and AND4 (N15868, N15865, N1936, N12482, N14854);
not NOT1 (N15869, N15851);
and AND4 (N15870, N15850, N9544, N10718, N15863);
not NOT1 (N15871, N15868);
nand NAND3 (N15872, N15846, N3804, N12020);
nor NOR2 (N15873, N15861, N1679);
not NOT1 (N15874, N15858);
not NOT1 (N15875, N15869);
nand NAND4 (N15876, N15873, N8369, N2675, N2291);
xor XOR2 (N15877, N15876, N9934);
nor NOR3 (N15878, N15871, N8827, N5852);
nor NOR3 (N15879, N15877, N6930, N11164);
xor XOR2 (N15880, N15879, N10296);
nor NOR3 (N15881, N15859, N13786, N14201);
and AND2 (N15882, N15872, N11525);
xor XOR2 (N15883, N15867, N7291);
xor XOR2 (N15884, N15883, N10302);
or OR4 (N15885, N15870, N7403, N7480, N15426);
not NOT1 (N15886, N15884);
and AND2 (N15887, N15878, N11740);
nor NOR4 (N15888, N15887, N4349, N6066, N2733);
xor XOR2 (N15889, N15881, N11274);
buf BUF1 (N15890, N15886);
not NOT1 (N15891, N15860);
nor NOR2 (N15892, N15885, N11218);
and AND2 (N15893, N15889, N6440);
and AND4 (N15894, N15882, N13018, N11853, N12718);
or OR2 (N15895, N15880, N13010);
nor NOR4 (N15896, N15894, N5804, N3716, N14622);
nand NAND2 (N15897, N15890, N3255);
buf BUF1 (N15898, N15893);
xor XOR2 (N15899, N15895, N518);
nor NOR4 (N15900, N15896, N8256, N14792, N3279);
xor XOR2 (N15901, N15866, N1751);
not NOT1 (N15902, N15892);
nand NAND3 (N15903, N15888, N7577, N15395);
xor XOR2 (N15904, N15902, N13666);
buf BUF1 (N15905, N15874);
nor NOR4 (N15906, N15875, N5338, N13126, N10939);
not NOT1 (N15907, N15901);
or OR2 (N15908, N15899, N11649);
nor NOR2 (N15909, N15903, N1152);
xor XOR2 (N15910, N15898, N10448);
nand NAND4 (N15911, N15910, N2383, N10171, N4017);
or OR4 (N15912, N15904, N15345, N10596, N3559);
nor NOR3 (N15913, N15912, N5481, N10907);
xor XOR2 (N15914, N15906, N2061);
not NOT1 (N15915, N15905);
not NOT1 (N15916, N15907);
buf BUF1 (N15917, N15897);
or OR3 (N15918, N15911, N9747, N6763);
not NOT1 (N15919, N15918);
or OR2 (N15920, N15916, N7598);
buf BUF1 (N15921, N15920);
nor NOR2 (N15922, N15891, N3313);
not NOT1 (N15923, N15914);
and AND2 (N15924, N15915, N2628);
nor NOR2 (N15925, N15922, N3820);
nor NOR2 (N15926, N15919, N10845);
and AND4 (N15927, N15921, N2633, N13893, N993);
nand NAND2 (N15928, N15926, N7774);
not NOT1 (N15929, N15917);
or OR2 (N15930, N15913, N7639);
nor NOR2 (N15931, N15929, N9900);
or OR2 (N15932, N15925, N5390);
nor NOR4 (N15933, N15909, N8968, N778, N13401);
and AND4 (N15934, N15932, N10591, N10712, N3664);
or OR2 (N15935, N15908, N15089);
and AND4 (N15936, N15928, N3256, N12998, N5224);
not NOT1 (N15937, N15927);
or OR3 (N15938, N15900, N2269, N1174);
nor NOR3 (N15939, N15933, N10200, N14783);
nor NOR2 (N15940, N15934, N14590);
and AND2 (N15941, N15936, N14820);
not NOT1 (N15942, N15931);
nand NAND2 (N15943, N15940, N5272);
xor XOR2 (N15944, N15943, N10547);
or OR4 (N15945, N15930, N3432, N13384, N10337);
and AND4 (N15946, N15924, N2359, N11599, N14214);
xor XOR2 (N15947, N15946, N4862);
not NOT1 (N15948, N15935);
nand NAND3 (N15949, N15944, N6212, N4256);
xor XOR2 (N15950, N15923, N6204);
buf BUF1 (N15951, N15937);
nand NAND3 (N15952, N15938, N11718, N14235);
xor XOR2 (N15953, N15945, N15727);
or OR3 (N15954, N15952, N4307, N5862);
xor XOR2 (N15955, N15951, N2555);
xor XOR2 (N15956, N15955, N9886);
xor XOR2 (N15957, N15941, N5092);
or OR2 (N15958, N15954, N63);
xor XOR2 (N15959, N15957, N3249);
and AND2 (N15960, N15953, N4397);
not NOT1 (N15961, N15939);
xor XOR2 (N15962, N15942, N9166);
or OR3 (N15963, N15959, N13281, N1997);
nor NOR4 (N15964, N15960, N3129, N4186, N6890);
or OR3 (N15965, N15961, N6839, N8550);
buf BUF1 (N15966, N15965);
nor NOR3 (N15967, N15949, N12252, N2389);
and AND3 (N15968, N15962, N3378, N13399);
buf BUF1 (N15969, N15947);
nor NOR3 (N15970, N15966, N14693, N11817);
and AND2 (N15971, N15948, N11647);
nand NAND2 (N15972, N15970, N15384);
and AND2 (N15973, N15958, N14576);
buf BUF1 (N15974, N15956);
nor NOR2 (N15975, N15950, N5264);
nand NAND4 (N15976, N15975, N8289, N9794, N12453);
xor XOR2 (N15977, N15974, N12107);
not NOT1 (N15978, N15972);
buf BUF1 (N15979, N15971);
and AND3 (N15980, N15978, N12058, N1040);
nor NOR4 (N15981, N15967, N2480, N2431, N15442);
and AND2 (N15982, N15976, N5767);
nor NOR3 (N15983, N15963, N11284, N9087);
not NOT1 (N15984, N15981);
not NOT1 (N15985, N15968);
nand NAND2 (N15986, N15979, N3044);
or OR3 (N15987, N15969, N3427, N1373);
or OR2 (N15988, N15964, N5576);
not NOT1 (N15989, N15973);
xor XOR2 (N15990, N15980, N9671);
and AND4 (N15991, N15983, N8796, N12878, N15934);
nand NAND2 (N15992, N15984, N7179);
or OR3 (N15993, N15982, N14056, N10344);
xor XOR2 (N15994, N15986, N1749);
not NOT1 (N15995, N15991);
nor NOR4 (N15996, N15987, N2341, N6441, N11809);
not NOT1 (N15997, N15985);
xor XOR2 (N15998, N15994, N1600);
buf BUF1 (N15999, N15997);
nand NAND2 (N16000, N15996, N12127);
buf BUF1 (N16001, N15990);
and AND3 (N16002, N16000, N1491, N1808);
and AND4 (N16003, N15977, N8351, N15903, N11474);
and AND3 (N16004, N15993, N15929, N8260);
nor NOR4 (N16005, N15999, N7497, N8932, N11332);
nor NOR4 (N16006, N16004, N1451, N13365, N13607);
buf BUF1 (N16007, N16006);
buf BUF1 (N16008, N15995);
xor XOR2 (N16009, N16002, N3540);
nor NOR4 (N16010, N15992, N3447, N5198, N13719);
and AND3 (N16011, N16010, N2952, N2661);
buf BUF1 (N16012, N16003);
nand NAND4 (N16013, N16001, N10907, N12469, N11051);
and AND3 (N16014, N15989, N8988, N14679);
buf BUF1 (N16015, N16009);
nand NAND4 (N16016, N16011, N1785, N6199, N315);
not NOT1 (N16017, N16014);
and AND3 (N16018, N16007, N1019, N1880);
or OR3 (N16019, N16018, N7982, N13549);
buf BUF1 (N16020, N16016);
nor NOR3 (N16021, N16015, N15530, N7604);
nor NOR2 (N16022, N16013, N3647);
buf BUF1 (N16023, N16012);
or OR2 (N16024, N16023, N6776);
and AND4 (N16025, N16022, N1950, N12129, N10487);
nand NAND3 (N16026, N16020, N3853, N5325);
or OR2 (N16027, N16026, N15928);
and AND2 (N16028, N16021, N10733);
or OR2 (N16029, N16027, N3658);
buf BUF1 (N16030, N15998);
xor XOR2 (N16031, N16028, N4773);
xor XOR2 (N16032, N16025, N15875);
buf BUF1 (N16033, N16032);
xor XOR2 (N16034, N16031, N4950);
not NOT1 (N16035, N16024);
buf BUF1 (N16036, N16008);
buf BUF1 (N16037, N15988);
buf BUF1 (N16038, N16033);
nand NAND4 (N16039, N16037, N3724, N14080, N4827);
xor XOR2 (N16040, N16035, N50);
nand NAND4 (N16041, N16040, N4803, N12450, N10788);
nand NAND3 (N16042, N16038, N14812, N2652);
nor NOR4 (N16043, N16019, N14405, N5351, N11999);
nor NOR2 (N16044, N16043, N13774);
and AND3 (N16045, N16017, N2217, N7922);
nand NAND2 (N16046, N16039, N2844);
or OR2 (N16047, N16045, N4546);
xor XOR2 (N16048, N16029, N9852);
nand NAND4 (N16049, N16042, N13452, N15893, N8670);
buf BUF1 (N16050, N16046);
or OR4 (N16051, N16050, N11527, N14061, N11656);
or OR2 (N16052, N16048, N10583);
buf BUF1 (N16053, N16041);
xor XOR2 (N16054, N16051, N6703);
and AND4 (N16055, N16005, N1849, N3180, N10206);
nor NOR3 (N16056, N16047, N8231, N14105);
nor NOR4 (N16057, N16054, N8791, N3569, N431);
or OR3 (N16058, N16036, N3220, N10582);
and AND3 (N16059, N16052, N6819, N12973);
xor XOR2 (N16060, N16044, N10002);
and AND2 (N16061, N16030, N4188);
xor XOR2 (N16062, N16053, N2820);
not NOT1 (N16063, N16049);
or OR4 (N16064, N16059, N6573, N116, N13407);
buf BUF1 (N16065, N16056);
nor NOR2 (N16066, N16063, N3897);
not NOT1 (N16067, N16065);
or OR4 (N16068, N16064, N11953, N11891, N10243);
nand NAND4 (N16069, N16062, N6132, N5218, N11096);
not NOT1 (N16070, N16058);
or OR4 (N16071, N16034, N2843, N14710, N643);
nand NAND3 (N16072, N16071, N5267, N1321);
or OR2 (N16073, N16067, N7633);
nor NOR3 (N16074, N16069, N10663, N3003);
or OR2 (N16075, N16070, N8780);
buf BUF1 (N16076, N16057);
or OR3 (N16077, N16072, N6027, N1124);
or OR3 (N16078, N16077, N7610, N10776);
and AND3 (N16079, N16073, N6431, N14210);
and AND3 (N16080, N16074, N10106, N1686);
or OR2 (N16081, N16080, N4566);
and AND4 (N16082, N16081, N7561, N5504, N10566);
and AND4 (N16083, N16066, N10996, N11714, N5070);
and AND2 (N16084, N16079, N13060);
and AND2 (N16085, N16083, N2627);
nand NAND4 (N16086, N16055, N11296, N8493, N6159);
not NOT1 (N16087, N16061);
nor NOR4 (N16088, N16087, N14543, N15384, N13008);
or OR2 (N16089, N16082, N9383);
nand NAND2 (N16090, N16086, N5866);
and AND4 (N16091, N16060, N15390, N6941, N4700);
and AND2 (N16092, N16084, N11975);
or OR2 (N16093, N16075, N3456);
and AND4 (N16094, N16093, N9858, N11192, N11639);
buf BUF1 (N16095, N16091);
or OR4 (N16096, N16085, N9804, N9789, N9214);
buf BUF1 (N16097, N16094);
buf BUF1 (N16098, N16078);
and AND3 (N16099, N16076, N8054, N15822);
or OR4 (N16100, N16096, N5889, N9868, N7810);
nor NOR4 (N16101, N16092, N14441, N9502, N15101);
buf BUF1 (N16102, N16100);
not NOT1 (N16103, N16099);
and AND3 (N16104, N16103, N7779, N2688);
nand NAND3 (N16105, N16104, N12985, N1163);
xor XOR2 (N16106, N16095, N14335);
nor NOR3 (N16107, N16088, N4409, N2991);
nor NOR3 (N16108, N16101, N10229, N13674);
nor NOR2 (N16109, N16098, N3025);
and AND2 (N16110, N16109, N13250);
or OR2 (N16111, N16105, N14230);
nand NAND2 (N16112, N16068, N4268);
xor XOR2 (N16113, N16102, N841);
nand NAND3 (N16114, N16111, N15883, N7672);
or OR3 (N16115, N16112, N14199, N134);
xor XOR2 (N16116, N16108, N14820);
nor NOR2 (N16117, N16106, N15027);
buf BUF1 (N16118, N16090);
buf BUF1 (N16119, N16107);
buf BUF1 (N16120, N16114);
not NOT1 (N16121, N16115);
nand NAND3 (N16122, N16118, N15567, N5337);
nor NOR2 (N16123, N16110, N4798);
not NOT1 (N16124, N16116);
nor NOR4 (N16125, N16097, N1910, N12267, N859);
not NOT1 (N16126, N16122);
and AND4 (N16127, N16121, N4089, N12540, N13056);
or OR3 (N16128, N16124, N10046, N14181);
or OR4 (N16129, N16089, N11715, N1262, N14874);
not NOT1 (N16130, N16123);
or OR4 (N16131, N16125, N4230, N449, N8424);
and AND2 (N16132, N16113, N10123);
nand NAND2 (N16133, N16129, N5330);
nor NOR3 (N16134, N16117, N15150, N13133);
buf BUF1 (N16135, N16130);
or OR2 (N16136, N16119, N8611);
xor XOR2 (N16137, N16131, N1117);
buf BUF1 (N16138, N16134);
xor XOR2 (N16139, N16127, N2450);
nand NAND4 (N16140, N16135, N11843, N12132, N15009);
nand NAND3 (N16141, N16133, N6224, N15748);
nor NOR4 (N16142, N16138, N6064, N3995, N12169);
xor XOR2 (N16143, N16139, N294);
and AND3 (N16144, N16132, N15144, N10691);
and AND3 (N16145, N16136, N12318, N356);
and AND3 (N16146, N16142, N13405, N6628);
or OR2 (N16147, N16143, N1850);
nor NOR2 (N16148, N16144, N4396);
nor NOR2 (N16149, N16137, N5198);
nor NOR2 (N16150, N16120, N3431);
not NOT1 (N16151, N16145);
or OR2 (N16152, N16149, N2020);
xor XOR2 (N16153, N16126, N1638);
xor XOR2 (N16154, N16151, N6219);
and AND2 (N16155, N16140, N8161);
not NOT1 (N16156, N16154);
buf BUF1 (N16157, N16156);
nor NOR4 (N16158, N16155, N1757, N13315, N1241);
nor NOR2 (N16159, N16158, N13869);
nand NAND3 (N16160, N16147, N3321, N6606);
nand NAND2 (N16161, N16152, N12968);
not NOT1 (N16162, N16150);
buf BUF1 (N16163, N16162);
not NOT1 (N16164, N16148);
nand NAND3 (N16165, N16159, N3286, N9611);
xor XOR2 (N16166, N16164, N12038);
and AND2 (N16167, N16146, N4222);
nand NAND2 (N16168, N16160, N8024);
not NOT1 (N16169, N16128);
xor XOR2 (N16170, N16167, N2453);
not NOT1 (N16171, N16141);
nor NOR4 (N16172, N16169, N2292, N630, N10138);
not NOT1 (N16173, N16168);
buf BUF1 (N16174, N16170);
or OR2 (N16175, N16165, N7346);
and AND4 (N16176, N16166, N12990, N11591, N10883);
not NOT1 (N16177, N16172);
and AND2 (N16178, N16173, N4337);
nand NAND4 (N16179, N16161, N13943, N1445, N7223);
or OR4 (N16180, N16171, N3419, N681, N13481);
not NOT1 (N16181, N16163);
and AND3 (N16182, N16180, N8799, N4724);
buf BUF1 (N16183, N16177);
nand NAND3 (N16184, N16157, N10075, N7436);
nand NAND3 (N16185, N16174, N6803, N15042);
nand NAND2 (N16186, N16176, N6706);
xor XOR2 (N16187, N16153, N16007);
nor NOR2 (N16188, N16185, N7898);
and AND4 (N16189, N16183, N1250, N13932, N10944);
not NOT1 (N16190, N16175);
not NOT1 (N16191, N16187);
and AND2 (N16192, N16188, N4554);
or OR3 (N16193, N16181, N2595, N8743);
and AND4 (N16194, N16178, N2467, N15950, N451);
nand NAND2 (N16195, N16191, N953);
or OR4 (N16196, N16182, N4323, N15320, N5089);
nor NOR3 (N16197, N16192, N4323, N7742);
xor XOR2 (N16198, N16194, N8231);
xor XOR2 (N16199, N16193, N10898);
nor NOR4 (N16200, N16189, N3058, N5100, N15569);
and AND3 (N16201, N16200, N8345, N6298);
xor XOR2 (N16202, N16184, N8541);
xor XOR2 (N16203, N16199, N5625);
or OR4 (N16204, N16203, N14, N8568, N3274);
or OR3 (N16205, N16201, N11775, N3868);
nor NOR4 (N16206, N16195, N11985, N3024, N10272);
not NOT1 (N16207, N16204);
nand NAND3 (N16208, N16202, N6344, N10214);
not NOT1 (N16209, N16206);
xor XOR2 (N16210, N16179, N6784);
and AND2 (N16211, N16196, N14068);
nor NOR4 (N16212, N16205, N15693, N13969, N5494);
xor XOR2 (N16213, N16209, N9405);
nor NOR4 (N16214, N16207, N9975, N10544, N11620);
nand NAND2 (N16215, N16214, N2655);
or OR4 (N16216, N16198, N13229, N6426, N11343);
or OR3 (N16217, N16208, N11099, N11686);
or OR3 (N16218, N16212, N13182, N2608);
not NOT1 (N16219, N16216);
xor XOR2 (N16220, N16218, N8623);
xor XOR2 (N16221, N16219, N295);
nor NOR2 (N16222, N16197, N14447);
nand NAND3 (N16223, N16186, N2398, N785);
xor XOR2 (N16224, N16213, N6071);
buf BUF1 (N16225, N16217);
nor NOR3 (N16226, N16222, N13216, N1718);
or OR3 (N16227, N16225, N14702, N8778);
or OR3 (N16228, N16223, N1408, N9206);
not NOT1 (N16229, N16210);
or OR3 (N16230, N16227, N997, N5060);
xor XOR2 (N16231, N16221, N7121);
nand NAND4 (N16232, N16226, N3449, N12919, N8460);
xor XOR2 (N16233, N16215, N14896);
not NOT1 (N16234, N16233);
not NOT1 (N16235, N16231);
xor XOR2 (N16236, N16230, N15105);
buf BUF1 (N16237, N16190);
buf BUF1 (N16238, N16224);
nor NOR3 (N16239, N16234, N12710, N3481);
buf BUF1 (N16240, N16239);
xor XOR2 (N16241, N16232, N14001);
and AND2 (N16242, N16220, N6380);
buf BUF1 (N16243, N16211);
or OR2 (N16244, N16237, N12889);
xor XOR2 (N16245, N16241, N14230);
nand NAND3 (N16246, N16243, N15587, N6041);
xor XOR2 (N16247, N16240, N15556);
nor NOR2 (N16248, N16245, N2591);
and AND3 (N16249, N16248, N4731, N4345);
or OR3 (N16250, N16228, N2262, N13907);
or OR3 (N16251, N16244, N5349, N10128);
not NOT1 (N16252, N16235);
nor NOR3 (N16253, N16247, N13529, N12778);
or OR3 (N16254, N16250, N2050, N15225);
not NOT1 (N16255, N16254);
xor XOR2 (N16256, N16252, N13427);
nand NAND4 (N16257, N16253, N12841, N3847, N10207);
nor NOR4 (N16258, N16238, N2721, N1179, N8909);
nor NOR2 (N16259, N16255, N4114);
not NOT1 (N16260, N16256);
nor NOR4 (N16261, N16260, N2182, N11693, N5419);
or OR3 (N16262, N16259, N1175, N7914);
not NOT1 (N16263, N16246);
buf BUF1 (N16264, N16263);
and AND3 (N16265, N16249, N11971, N10233);
and AND3 (N16266, N16229, N1086, N288);
nor NOR3 (N16267, N16251, N3211, N9410);
buf BUF1 (N16268, N16236);
nand NAND2 (N16269, N16262, N1302);
nand NAND3 (N16270, N16268, N16067, N9110);
buf BUF1 (N16271, N16265);
not NOT1 (N16272, N16257);
xor XOR2 (N16273, N16264, N13342);
nand NAND2 (N16274, N16271, N15231);
nor NOR3 (N16275, N16270, N4388, N10282);
nand NAND4 (N16276, N16267, N15243, N955, N5307);
nand NAND3 (N16277, N16269, N7085, N14625);
not NOT1 (N16278, N16258);
xor XOR2 (N16279, N16274, N16043);
buf BUF1 (N16280, N16266);
and AND3 (N16281, N16273, N16262, N12044);
not NOT1 (N16282, N16280);
not NOT1 (N16283, N16278);
or OR2 (N16284, N16272, N9223);
or OR2 (N16285, N16279, N2480);
and AND3 (N16286, N16276, N10568, N12183);
xor XOR2 (N16287, N16286, N1604);
buf BUF1 (N16288, N16275);
not NOT1 (N16289, N16282);
buf BUF1 (N16290, N16283);
and AND3 (N16291, N16288, N10985, N1948);
xor XOR2 (N16292, N16290, N11592);
or OR4 (N16293, N16291, N11424, N10925, N14136);
buf BUF1 (N16294, N16281);
and AND2 (N16295, N16292, N7266);
nor NOR2 (N16296, N16277, N11204);
buf BUF1 (N16297, N16289);
or OR4 (N16298, N16297, N5211, N7330, N6319);
not NOT1 (N16299, N16285);
xor XOR2 (N16300, N16298, N15406);
nor NOR2 (N16301, N16300, N2796);
nor NOR4 (N16302, N16287, N11266, N8360, N10054);
xor XOR2 (N16303, N16296, N3282);
xor XOR2 (N16304, N16293, N13606);
buf BUF1 (N16305, N16295);
not NOT1 (N16306, N16299);
xor XOR2 (N16307, N16301, N9031);
nor NOR4 (N16308, N16242, N627, N6699, N14490);
xor XOR2 (N16309, N16307, N6195);
nor NOR2 (N16310, N16261, N11821);
and AND3 (N16311, N16303, N11096, N9489);
xor XOR2 (N16312, N16305, N13608);
or OR4 (N16313, N16306, N16114, N14558, N4188);
buf BUF1 (N16314, N16302);
xor XOR2 (N16315, N16284, N10965);
and AND3 (N16316, N16310, N1961, N9613);
or OR2 (N16317, N16316, N944);
buf BUF1 (N16318, N16314);
not NOT1 (N16319, N16313);
xor XOR2 (N16320, N16308, N533);
nand NAND2 (N16321, N16304, N1077);
not NOT1 (N16322, N16318);
or OR4 (N16323, N16315, N13328, N2500, N1867);
not NOT1 (N16324, N16317);
not NOT1 (N16325, N16322);
nor NOR4 (N16326, N16311, N16258, N3816, N14873);
or OR3 (N16327, N16325, N3070, N16310);
not NOT1 (N16328, N16326);
or OR2 (N16329, N16294, N4591);
and AND4 (N16330, N16329, N10286, N9047, N11096);
xor XOR2 (N16331, N16309, N9554);
nand NAND4 (N16332, N16330, N9546, N2551, N7793);
and AND2 (N16333, N16332, N8849);
nand NAND2 (N16334, N16331, N782);
nor NOR4 (N16335, N16324, N10178, N13704, N7159);
nand NAND2 (N16336, N16320, N4141);
buf BUF1 (N16337, N16323);
nand NAND2 (N16338, N16328, N9424);
nor NOR2 (N16339, N16321, N11353);
and AND3 (N16340, N16335, N6589, N13354);
nor NOR4 (N16341, N16327, N5490, N10831, N12796);
and AND4 (N16342, N16338, N14653, N2996, N11112);
not NOT1 (N16343, N16337);
nand NAND4 (N16344, N16312, N3995, N327, N7488);
and AND2 (N16345, N16342, N12802);
xor XOR2 (N16346, N16336, N2377);
nand NAND2 (N16347, N16319, N6110);
not NOT1 (N16348, N16345);
nor NOR3 (N16349, N16341, N5069, N11500);
or OR2 (N16350, N16343, N14098);
xor XOR2 (N16351, N16333, N1631);
or OR2 (N16352, N16350, N12167);
nand NAND3 (N16353, N16348, N9021, N1988);
buf BUF1 (N16354, N16351);
or OR2 (N16355, N16354, N14793);
or OR4 (N16356, N16340, N10014, N3637, N3459);
xor XOR2 (N16357, N16346, N2394);
or OR4 (N16358, N16347, N15814, N15516, N5611);
nor NOR4 (N16359, N16356, N7666, N10541, N5806);
or OR3 (N16360, N16349, N8900, N11644);
buf BUF1 (N16361, N16344);
or OR4 (N16362, N16358, N700, N8032, N15245);
or OR3 (N16363, N16355, N1199, N8811);
not NOT1 (N16364, N16361);
nand NAND2 (N16365, N16352, N6155);
xor XOR2 (N16366, N16339, N6279);
or OR4 (N16367, N16353, N10887, N5169, N4316);
xor XOR2 (N16368, N16365, N15636);
xor XOR2 (N16369, N16366, N388);
or OR2 (N16370, N16363, N5813);
and AND4 (N16371, N16364, N9124, N4410, N13482);
and AND3 (N16372, N16370, N6500, N7148);
buf BUF1 (N16373, N16372);
and AND2 (N16374, N16359, N6403);
nor NOR4 (N16375, N16374, N671, N8815, N11848);
or OR3 (N16376, N16371, N7940, N457);
buf BUF1 (N16377, N16367);
xor XOR2 (N16378, N16360, N2532);
or OR2 (N16379, N16368, N3900);
xor XOR2 (N16380, N16362, N10707);
xor XOR2 (N16381, N16379, N1531);
nor NOR4 (N16382, N16378, N14596, N9390, N985);
xor XOR2 (N16383, N16381, N2016);
or OR2 (N16384, N16334, N10498);
nor NOR2 (N16385, N16384, N14859);
nand NAND4 (N16386, N16380, N12026, N534, N6712);
xor XOR2 (N16387, N16373, N16069);
and AND4 (N16388, N16377, N6941, N15148, N469);
nor NOR3 (N16389, N16369, N16380, N11938);
nor NOR3 (N16390, N16375, N10916, N7760);
or OR2 (N16391, N16390, N14231);
or OR2 (N16392, N16386, N6330);
and AND2 (N16393, N16388, N8014);
or OR4 (N16394, N16393, N7014, N15366, N5356);
and AND4 (N16395, N16383, N11651, N5991, N3442);
xor XOR2 (N16396, N16385, N7962);
nor NOR4 (N16397, N16389, N7501, N8804, N3313);
nand NAND4 (N16398, N16391, N13283, N691, N2050);
nand NAND3 (N16399, N16394, N9339, N9579);
not NOT1 (N16400, N16397);
nor NOR4 (N16401, N16357, N10651, N16001, N9173);
and AND3 (N16402, N16382, N2196, N2104);
xor XOR2 (N16403, N16392, N10009);
and AND3 (N16404, N16403, N3526, N13156);
not NOT1 (N16405, N16399);
buf BUF1 (N16406, N16402);
xor XOR2 (N16407, N16404, N14254);
not NOT1 (N16408, N16387);
xor XOR2 (N16409, N16400, N10746);
not NOT1 (N16410, N16409);
xor XOR2 (N16411, N16396, N3326);
xor XOR2 (N16412, N16406, N506);
nor NOR3 (N16413, N16408, N20, N8311);
nand NAND2 (N16414, N16395, N2919);
or OR3 (N16415, N16376, N3157, N1814);
or OR4 (N16416, N16401, N6313, N7007, N7095);
and AND3 (N16417, N16407, N9775, N13117);
buf BUF1 (N16418, N16413);
and AND4 (N16419, N16418, N5547, N5755, N12253);
nand NAND2 (N16420, N16419, N7330);
xor XOR2 (N16421, N16405, N6699);
not NOT1 (N16422, N16421);
not NOT1 (N16423, N16398);
not NOT1 (N16424, N16422);
buf BUF1 (N16425, N16424);
not NOT1 (N16426, N16420);
and AND2 (N16427, N16414, N603);
nand NAND4 (N16428, N16423, N5170, N6400, N10961);
buf BUF1 (N16429, N16412);
and AND4 (N16430, N16427, N768, N5910, N9984);
and AND3 (N16431, N16415, N249, N1130);
or OR4 (N16432, N16426, N9618, N10102, N5404);
nor NOR2 (N16433, N16428, N11888);
nor NOR3 (N16434, N16430, N12938, N8361);
buf BUF1 (N16435, N16416);
not NOT1 (N16436, N16433);
nor NOR3 (N16437, N16432, N14520, N14611);
nor NOR4 (N16438, N16417, N2655, N7534, N7621);
buf BUF1 (N16439, N16410);
and AND2 (N16440, N16436, N9461);
and AND2 (N16441, N16438, N15431);
and AND2 (N16442, N16431, N4293);
buf BUF1 (N16443, N16440);
xor XOR2 (N16444, N16435, N10595);
buf BUF1 (N16445, N16444);
and AND3 (N16446, N16442, N14863, N635);
xor XOR2 (N16447, N16411, N9960);
nand NAND4 (N16448, N16439, N15562, N9582, N12061);
xor XOR2 (N16449, N16445, N9399);
not NOT1 (N16450, N16429);
and AND4 (N16451, N16443, N8333, N4997, N2558);
not NOT1 (N16452, N16446);
nand NAND3 (N16453, N16441, N12357, N5472);
nand NAND4 (N16454, N16453, N3710, N10920, N11138);
not NOT1 (N16455, N16452);
and AND2 (N16456, N16451, N2288);
and AND3 (N16457, N16449, N14901, N11984);
or OR2 (N16458, N16434, N13352);
nor NOR3 (N16459, N16425, N13132, N14676);
buf BUF1 (N16460, N16448);
and AND4 (N16461, N16437, N8321, N11305, N217);
xor XOR2 (N16462, N16450, N15566);
xor XOR2 (N16463, N16461, N13293);
nand NAND3 (N16464, N16460, N5641, N8641);
or OR2 (N16465, N16459, N13393);
nor NOR3 (N16466, N16456, N3783, N2277);
xor XOR2 (N16467, N16455, N8051);
not NOT1 (N16468, N16465);
buf BUF1 (N16469, N16468);
or OR3 (N16470, N16463, N14565, N585);
nor NOR4 (N16471, N16469, N13209, N6475, N182);
buf BUF1 (N16472, N16462);
nor NOR2 (N16473, N16467, N5271);
or OR4 (N16474, N16470, N14972, N11156, N2128);
and AND2 (N16475, N16466, N9873);
nor NOR4 (N16476, N16471, N9908, N7684, N2886);
nor NOR4 (N16477, N16457, N7981, N15777, N10194);
not NOT1 (N16478, N16475);
buf BUF1 (N16479, N16464);
nor NOR3 (N16480, N16477, N8379, N8618);
and AND3 (N16481, N16479, N1009, N1851);
nor NOR3 (N16482, N16473, N10938, N5571);
nor NOR3 (N16483, N16478, N11671, N1211);
buf BUF1 (N16484, N16474);
nor NOR4 (N16485, N16454, N15113, N13236, N3807);
xor XOR2 (N16486, N16483, N15249);
nor NOR2 (N16487, N16447, N6910);
and AND3 (N16488, N16484, N337, N8239);
and AND4 (N16489, N16488, N1208, N10813, N15456);
or OR2 (N16490, N16480, N5940);
or OR4 (N16491, N16472, N10110, N13644, N11233);
and AND3 (N16492, N16486, N12664, N8372);
or OR2 (N16493, N16485, N4861);
not NOT1 (N16494, N16487);
xor XOR2 (N16495, N16476, N4264);
not NOT1 (N16496, N16494);
nor NOR2 (N16497, N16493, N3371);
and AND2 (N16498, N16481, N15945);
buf BUF1 (N16499, N16489);
xor XOR2 (N16500, N16458, N11525);
or OR3 (N16501, N16492, N3625, N5185);
nor NOR4 (N16502, N16501, N15967, N16356, N8571);
nor NOR3 (N16503, N16495, N5923, N885);
and AND2 (N16504, N16496, N6163);
or OR3 (N16505, N16482, N5534, N327);
nor NOR4 (N16506, N16491, N3148, N2256, N11090);
xor XOR2 (N16507, N16502, N817);
nand NAND3 (N16508, N16497, N10510, N2330);
or OR4 (N16509, N16503, N11092, N15493, N9588);
xor XOR2 (N16510, N16505, N13872);
nand NAND4 (N16511, N16490, N7099, N15545, N9426);
nand NAND3 (N16512, N16499, N3822, N8510);
nor NOR4 (N16513, N16511, N8127, N6973, N6095);
xor XOR2 (N16514, N16512, N1266);
or OR4 (N16515, N16498, N6786, N11073, N10064);
xor XOR2 (N16516, N16504, N12960);
xor XOR2 (N16517, N16507, N11365);
xor XOR2 (N16518, N16506, N11251);
or OR3 (N16519, N16515, N11760, N9000);
nand NAND2 (N16520, N16509, N4716);
or OR2 (N16521, N16500, N1049);
buf BUF1 (N16522, N16510);
not NOT1 (N16523, N16516);
nor NOR4 (N16524, N16517, N13641, N8182, N12166);
not NOT1 (N16525, N16518);
nor NOR3 (N16526, N16523, N5145, N14230);
nor NOR2 (N16527, N16526, N11735);
nand NAND2 (N16528, N16522, N15956);
nor NOR4 (N16529, N16519, N9928, N6457, N2830);
not NOT1 (N16530, N16520);
buf BUF1 (N16531, N16527);
nand NAND4 (N16532, N16508, N8241, N11746, N5238);
nor NOR4 (N16533, N16528, N2670, N8552, N4771);
xor XOR2 (N16534, N16525, N5698);
nand NAND3 (N16535, N16534, N12183, N4788);
nor NOR3 (N16536, N16531, N2874, N13903);
nand NAND4 (N16537, N16514, N12941, N12884, N2083);
xor XOR2 (N16538, N16513, N14182);
nand NAND4 (N16539, N16524, N4328, N4644, N12847);
xor XOR2 (N16540, N16532, N12751);
buf BUF1 (N16541, N16530);
nor NOR3 (N16542, N16529, N5091, N4856);
xor XOR2 (N16543, N16538, N15931);
or OR3 (N16544, N16539, N11662, N16531);
not NOT1 (N16545, N16541);
and AND4 (N16546, N16542, N5463, N10758, N1921);
not NOT1 (N16547, N16535);
or OR3 (N16548, N16521, N12334, N10706);
or OR4 (N16549, N16548, N758, N12262, N4124);
nor NOR4 (N16550, N16536, N8758, N3704, N2004);
nor NOR3 (N16551, N16546, N16341, N1012);
buf BUF1 (N16552, N16550);
or OR4 (N16553, N16552, N10186, N6490, N10883);
nor NOR3 (N16554, N16540, N1907, N7743);
buf BUF1 (N16555, N16547);
nor NOR2 (N16556, N16545, N949);
not NOT1 (N16557, N16544);
buf BUF1 (N16558, N16553);
and AND3 (N16559, N16549, N16086, N15789);
not NOT1 (N16560, N16533);
and AND4 (N16561, N16560, N13176, N14598, N6353);
nor NOR3 (N16562, N16556, N7269, N2738);
xor XOR2 (N16563, N16555, N6953);
and AND3 (N16564, N16562, N5553, N10311);
nand NAND4 (N16565, N16564, N4554, N548, N9148);
xor XOR2 (N16566, N16551, N10913);
nand NAND4 (N16567, N16561, N6985, N2295, N13162);
nor NOR2 (N16568, N16565, N12071);
or OR3 (N16569, N16537, N15250, N8874);
not NOT1 (N16570, N16568);
nand NAND3 (N16571, N16566, N11339, N13829);
and AND3 (N16572, N16543, N8727, N10234);
nand NAND2 (N16573, N16554, N13666);
nand NAND3 (N16574, N16563, N4286, N1056);
nand NAND4 (N16575, N16557, N15598, N1759, N12786);
and AND4 (N16576, N16571, N13411, N10989, N1210);
nand NAND2 (N16577, N16574, N9381);
and AND3 (N16578, N16559, N11609, N13608);
and AND4 (N16579, N16572, N7239, N15551, N5208);
buf BUF1 (N16580, N16558);
xor XOR2 (N16581, N16576, N15496);
buf BUF1 (N16582, N16575);
buf BUF1 (N16583, N16577);
buf BUF1 (N16584, N16573);
and AND4 (N16585, N16569, N10467, N13881, N12791);
xor XOR2 (N16586, N16570, N7637);
buf BUF1 (N16587, N16582);
or OR3 (N16588, N16578, N3058, N16307);
xor XOR2 (N16589, N16585, N12389);
buf BUF1 (N16590, N16579);
nand NAND4 (N16591, N16581, N2419, N12089, N4949);
buf BUF1 (N16592, N16591);
nand NAND4 (N16593, N16567, N3186, N7567, N700);
xor XOR2 (N16594, N16586, N15417);
or OR3 (N16595, N16589, N8281, N10127);
not NOT1 (N16596, N16580);
or OR2 (N16597, N16595, N4144);
or OR2 (N16598, N16592, N884);
or OR4 (N16599, N16588, N11098, N4182, N8614);
nor NOR3 (N16600, N16598, N5705, N4024);
xor XOR2 (N16601, N16599, N8929);
or OR3 (N16602, N16601, N5918, N9352);
buf BUF1 (N16603, N16602);
and AND3 (N16604, N16596, N1886, N2130);
buf BUF1 (N16605, N16587);
and AND4 (N16606, N16584, N3230, N11900, N12938);
nand NAND2 (N16607, N16583, N15598);
not NOT1 (N16608, N16603);
or OR2 (N16609, N16606, N2491);
nor NOR3 (N16610, N16607, N11911, N4366);
and AND4 (N16611, N16597, N7860, N4809, N8138);
buf BUF1 (N16612, N16610);
xor XOR2 (N16613, N16594, N1480);
buf BUF1 (N16614, N16609);
not NOT1 (N16615, N16613);
nand NAND3 (N16616, N16590, N8763, N12633);
xor XOR2 (N16617, N16605, N9611);
xor XOR2 (N16618, N16600, N13909);
not NOT1 (N16619, N16614);
and AND3 (N16620, N16616, N15210, N4359);
not NOT1 (N16621, N16620);
buf BUF1 (N16622, N16618);
xor XOR2 (N16623, N16593, N3660);
nand NAND3 (N16624, N16612, N3963, N12856);
and AND3 (N16625, N16623, N9100, N536);
or OR4 (N16626, N16619, N4869, N8909, N11715);
not NOT1 (N16627, N16626);
and AND2 (N16628, N16617, N14176);
buf BUF1 (N16629, N16608);
buf BUF1 (N16630, N16621);
not NOT1 (N16631, N16628);
xor XOR2 (N16632, N16629, N14730);
buf BUF1 (N16633, N16630);
buf BUF1 (N16634, N16611);
nor NOR4 (N16635, N16633, N10964, N2321, N14856);
xor XOR2 (N16636, N16604, N10788);
nand NAND4 (N16637, N16635, N13961, N11644, N12825);
buf BUF1 (N16638, N16625);
nor NOR2 (N16639, N16636, N10224);
nor NOR3 (N16640, N16631, N2913, N2642);
buf BUF1 (N16641, N16638);
and AND3 (N16642, N16639, N15626, N5708);
not NOT1 (N16643, N16642);
nor NOR4 (N16644, N16637, N11096, N5237, N13119);
buf BUF1 (N16645, N16624);
nand NAND2 (N16646, N16640, N6576);
xor XOR2 (N16647, N16645, N2965);
buf BUF1 (N16648, N16647);
buf BUF1 (N16649, N16646);
buf BUF1 (N16650, N16644);
nand NAND2 (N16651, N16648, N7513);
or OR3 (N16652, N16643, N8110, N9237);
or OR3 (N16653, N16652, N5343, N13361);
nand NAND2 (N16654, N16650, N1358);
or OR3 (N16655, N16654, N10231, N14663);
and AND2 (N16656, N16622, N6419);
or OR3 (N16657, N16656, N3567, N10043);
or OR4 (N16658, N16649, N15581, N444, N15035);
nand NAND3 (N16659, N16655, N3241, N10398);
or OR3 (N16660, N16627, N11140, N2711);
not NOT1 (N16661, N16641);
nor NOR4 (N16662, N16634, N2729, N5871, N8825);
nand NAND2 (N16663, N16662, N12197);
xor XOR2 (N16664, N16632, N9817);
not NOT1 (N16665, N16661);
not NOT1 (N16666, N16658);
or OR3 (N16667, N16665, N11646, N3174);
buf BUF1 (N16668, N16657);
nand NAND3 (N16669, N16659, N1672, N2654);
not NOT1 (N16670, N16615);
and AND3 (N16671, N16653, N3830, N10685);
nor NOR3 (N16672, N16667, N7982, N8421);
not NOT1 (N16673, N16660);
xor XOR2 (N16674, N16664, N1803);
or OR2 (N16675, N16674, N14964);
nor NOR3 (N16676, N16669, N13102, N13299);
and AND4 (N16677, N16663, N12411, N9815, N9874);
xor XOR2 (N16678, N16671, N13326);
buf BUF1 (N16679, N16668);
nor NOR2 (N16680, N16666, N4391);
xor XOR2 (N16681, N16651, N7027);
buf BUF1 (N16682, N16680);
and AND4 (N16683, N16670, N9501, N850, N695);
buf BUF1 (N16684, N16676);
buf BUF1 (N16685, N16673);
not NOT1 (N16686, N16678);
nor NOR4 (N16687, N16684, N6498, N10893, N8778);
not NOT1 (N16688, N16687);
and AND4 (N16689, N16686, N6735, N8895, N2529);
nor NOR2 (N16690, N16688, N12619);
or OR3 (N16691, N16675, N13919, N15693);
nand NAND4 (N16692, N16689, N14814, N10906, N14178);
xor XOR2 (N16693, N16682, N8534);
nand NAND2 (N16694, N16683, N2607);
not NOT1 (N16695, N16692);
nor NOR3 (N16696, N16681, N16572, N9677);
nand NAND3 (N16697, N16693, N9661, N6141);
not NOT1 (N16698, N16691);
nor NOR3 (N16699, N16685, N3637, N1757);
and AND3 (N16700, N16694, N9746, N9085);
nor NOR3 (N16701, N16679, N12473, N3553);
xor XOR2 (N16702, N16696, N647);
nor NOR3 (N16703, N16690, N2282, N88);
buf BUF1 (N16704, N16697);
nand NAND2 (N16705, N16698, N3725);
nand NAND4 (N16706, N16700, N3616, N15070, N10152);
nand NAND2 (N16707, N16703, N5623);
and AND2 (N16708, N16705, N7184);
xor XOR2 (N16709, N16707, N1688);
nor NOR2 (N16710, N16701, N6768);
xor XOR2 (N16711, N16677, N1667);
or OR3 (N16712, N16702, N14650, N2667);
nand NAND3 (N16713, N16711, N6193, N8521);
not NOT1 (N16714, N16713);
nor NOR4 (N16715, N16709, N15261, N3715, N13204);
nand NAND3 (N16716, N16704, N10726, N14072);
nand NAND4 (N16717, N16712, N9758, N8421, N2597);
xor XOR2 (N16718, N16715, N89);
buf BUF1 (N16719, N16718);
and AND3 (N16720, N16716, N13897, N5101);
not NOT1 (N16721, N16708);
and AND2 (N16722, N16672, N15556);
nor NOR2 (N16723, N16706, N556);
buf BUF1 (N16724, N16699);
nand NAND4 (N16725, N16723, N3622, N12821, N7423);
or OR4 (N16726, N16719, N2339, N6284, N11008);
nand NAND4 (N16727, N16717, N4630, N8245, N7382);
xor XOR2 (N16728, N16714, N13353);
not NOT1 (N16729, N16720);
and AND3 (N16730, N16721, N14443, N8315);
xor XOR2 (N16731, N16725, N6199);
not NOT1 (N16732, N16729);
buf BUF1 (N16733, N16724);
and AND2 (N16734, N16710, N6293);
nand NAND4 (N16735, N16734, N11683, N6487, N1039);
nor NOR2 (N16736, N16732, N6909);
nand NAND4 (N16737, N16695, N756, N13495, N2480);
and AND2 (N16738, N16730, N12613);
nor NOR4 (N16739, N16735, N391, N9642, N8980);
or OR3 (N16740, N16731, N7350, N413);
not NOT1 (N16741, N16727);
or OR3 (N16742, N16740, N481, N1367);
not NOT1 (N16743, N16728);
buf BUF1 (N16744, N16722);
not NOT1 (N16745, N16738);
nor NOR2 (N16746, N16737, N12092);
or OR3 (N16747, N16726, N2588, N2683);
and AND4 (N16748, N16745, N14953, N2796, N5550);
and AND2 (N16749, N16741, N8065);
xor XOR2 (N16750, N16746, N12204);
and AND3 (N16751, N16747, N5400, N15141);
nor NOR3 (N16752, N16744, N13141, N6475);
xor XOR2 (N16753, N16742, N9422);
and AND3 (N16754, N16749, N10737, N7241);
xor XOR2 (N16755, N16736, N14270);
xor XOR2 (N16756, N16748, N8457);
and AND3 (N16757, N16753, N13907, N14215);
nand NAND2 (N16758, N16754, N11964);
or OR2 (N16759, N16757, N2753);
or OR3 (N16760, N16733, N9280, N4301);
nand NAND4 (N16761, N16752, N9858, N3339, N14238);
or OR2 (N16762, N16761, N8739);
or OR4 (N16763, N16755, N7356, N15320, N8971);
buf BUF1 (N16764, N16759);
buf BUF1 (N16765, N16739);
nand NAND3 (N16766, N16758, N2167, N2971);
buf BUF1 (N16767, N16760);
xor XOR2 (N16768, N16765, N5261);
xor XOR2 (N16769, N16743, N8860);
buf BUF1 (N16770, N16767);
xor XOR2 (N16771, N16750, N13724);
and AND2 (N16772, N16762, N5891);
nand NAND3 (N16773, N16764, N6282, N4983);
nand NAND3 (N16774, N16770, N16687, N6017);
not NOT1 (N16775, N16773);
xor XOR2 (N16776, N16756, N5758);
and AND2 (N16777, N16771, N5700);
nand NAND3 (N16778, N16766, N503, N12529);
not NOT1 (N16779, N16777);
or OR4 (N16780, N16776, N12952, N8509, N10285);
or OR3 (N16781, N16769, N3110, N4453);
and AND2 (N16782, N16768, N6365);
and AND4 (N16783, N16751, N12967, N15177, N200);
nand NAND2 (N16784, N16763, N13377);
and AND2 (N16785, N16772, N5426);
nand NAND2 (N16786, N16782, N5721);
nand NAND4 (N16787, N16778, N4036, N4694, N7441);
nand NAND3 (N16788, N16785, N6552, N35);
nor NOR2 (N16789, N16788, N15313);
nor NOR3 (N16790, N16774, N11010, N10031);
nor NOR2 (N16791, N16779, N16772);
buf BUF1 (N16792, N16790);
xor XOR2 (N16793, N16784, N12187);
or OR2 (N16794, N16792, N2697);
buf BUF1 (N16795, N16783);
nand NAND3 (N16796, N16789, N504, N8498);
and AND4 (N16797, N16795, N6865, N13546, N10840);
nor NOR3 (N16798, N16775, N8405, N9670);
buf BUF1 (N16799, N16793);
nor NOR4 (N16800, N16787, N5313, N3026, N8805);
and AND4 (N16801, N16781, N4335, N9126, N11721);
nor NOR2 (N16802, N16780, N5507);
buf BUF1 (N16803, N16798);
nand NAND4 (N16804, N16801, N3563, N1831, N3249);
xor XOR2 (N16805, N16803, N5159);
buf BUF1 (N16806, N16802);
and AND3 (N16807, N16800, N13270, N15380);
xor XOR2 (N16808, N16807, N6332);
and AND3 (N16809, N16805, N7813, N8825);
and AND4 (N16810, N16806, N2983, N13942, N3292);
nor NOR2 (N16811, N16810, N5254);
nor NOR2 (N16812, N16794, N4167);
nor NOR2 (N16813, N16799, N5853);
xor XOR2 (N16814, N16786, N8544);
buf BUF1 (N16815, N16804);
nor NOR3 (N16816, N16797, N2510, N2244);
xor XOR2 (N16817, N16816, N3861);
not NOT1 (N16818, N16808);
buf BUF1 (N16819, N16818);
or OR2 (N16820, N16791, N3132);
or OR4 (N16821, N16815, N14263, N3478, N5774);
xor XOR2 (N16822, N16811, N4664);
and AND2 (N16823, N16809, N5377);
not NOT1 (N16824, N16819);
nor NOR2 (N16825, N16796, N6151);
xor XOR2 (N16826, N16817, N4608);
not NOT1 (N16827, N16822);
and AND2 (N16828, N16825, N14753);
xor XOR2 (N16829, N16813, N15993);
nand NAND3 (N16830, N16829, N4997, N14981);
nor NOR2 (N16831, N16814, N1066);
nand NAND4 (N16832, N16821, N15387, N9665, N13239);
not NOT1 (N16833, N16827);
nand NAND3 (N16834, N16831, N1539, N875);
or OR3 (N16835, N16830, N14797, N5056);
nand NAND3 (N16836, N16823, N12599, N15372);
xor XOR2 (N16837, N16828, N4927);
buf BUF1 (N16838, N16833);
nand NAND2 (N16839, N16820, N14422);
not NOT1 (N16840, N16835);
or OR3 (N16841, N16812, N263, N16691);
or OR2 (N16842, N16841, N3042);
not NOT1 (N16843, N16842);
nor NOR2 (N16844, N16843, N9422);
buf BUF1 (N16845, N16834);
not NOT1 (N16846, N16826);
or OR4 (N16847, N16838, N845, N11311, N2944);
nor NOR2 (N16848, N16832, N13120);
not NOT1 (N16849, N16845);
nor NOR3 (N16850, N16848, N14960, N3717);
nand NAND2 (N16851, N16836, N6872);
or OR4 (N16852, N16846, N11969, N13634, N15534);
buf BUF1 (N16853, N16852);
or OR4 (N16854, N16851, N2142, N1724, N11277);
nand NAND2 (N16855, N16840, N15486);
xor XOR2 (N16856, N16853, N13080);
not NOT1 (N16857, N16847);
nand NAND4 (N16858, N16854, N12847, N6326, N5385);
or OR2 (N16859, N16837, N16787);
buf BUF1 (N16860, N16844);
and AND3 (N16861, N16849, N11967, N10762);
buf BUF1 (N16862, N16859);
and AND3 (N16863, N16861, N7740, N1721);
or OR4 (N16864, N16850, N4233, N8538, N13470);
not NOT1 (N16865, N16855);
nor NOR3 (N16866, N16858, N12539, N12063);
and AND3 (N16867, N16862, N4192, N13511);
not NOT1 (N16868, N16857);
buf BUF1 (N16869, N16824);
not NOT1 (N16870, N16868);
xor XOR2 (N16871, N16864, N2493);
and AND2 (N16872, N16865, N16076);
or OR3 (N16873, N16871, N7662, N11242);
and AND4 (N16874, N16870, N15043, N14835, N14343);
buf BUF1 (N16875, N16873);
not NOT1 (N16876, N16874);
nor NOR4 (N16877, N16839, N9885, N2113, N5268);
not NOT1 (N16878, N16867);
and AND3 (N16879, N16872, N4166, N1637);
nor NOR4 (N16880, N16878, N10377, N8453, N5203);
nor NOR3 (N16881, N16880, N2796, N14708);
xor XOR2 (N16882, N16876, N13966);
buf BUF1 (N16883, N16856);
xor XOR2 (N16884, N16883, N10673);
not NOT1 (N16885, N16881);
not NOT1 (N16886, N16869);
xor XOR2 (N16887, N16866, N13465);
nor NOR4 (N16888, N16879, N12690, N2249, N1986);
xor XOR2 (N16889, N16888, N791);
and AND4 (N16890, N16889, N9340, N12201, N4589);
and AND2 (N16891, N16890, N16274);
nand NAND4 (N16892, N16863, N9595, N1952, N13824);
nor NOR2 (N16893, N16891, N980);
nand NAND2 (N16894, N16860, N5775);
buf BUF1 (N16895, N16887);
nor NOR2 (N16896, N16884, N11081);
not NOT1 (N16897, N16875);
nand NAND2 (N16898, N16885, N6058);
nand NAND4 (N16899, N16895, N5805, N7997, N3220);
nor NOR4 (N16900, N16896, N5510, N465, N5965);
or OR4 (N16901, N16882, N4159, N10208, N2800);
nand NAND3 (N16902, N16893, N2096, N12790);
not NOT1 (N16903, N16886);
not NOT1 (N16904, N16900);
xor XOR2 (N16905, N16899, N15975);
xor XOR2 (N16906, N16892, N12952);
not NOT1 (N16907, N16877);
nor NOR3 (N16908, N16897, N6609, N16581);
not NOT1 (N16909, N16903);
not NOT1 (N16910, N16898);
nor NOR2 (N16911, N16904, N10516);
nand NAND4 (N16912, N16909, N13839, N8496, N16904);
and AND3 (N16913, N16908, N2862, N2870);
xor XOR2 (N16914, N16907, N6498);
nand NAND2 (N16915, N16902, N7787);
xor XOR2 (N16916, N16911, N14255);
buf BUF1 (N16917, N16906);
not NOT1 (N16918, N16905);
nor NOR3 (N16919, N16894, N15918, N8428);
nor NOR4 (N16920, N16912, N13270, N9893, N9093);
nor NOR4 (N16921, N16918, N5948, N11290, N15441);
buf BUF1 (N16922, N16913);
nor NOR3 (N16923, N16916, N2754, N2909);
buf BUF1 (N16924, N16915);
nor NOR4 (N16925, N16922, N12184, N3084, N4516);
or OR4 (N16926, N16920, N12892, N5293, N12002);
xor XOR2 (N16927, N16924, N2405);
or OR3 (N16928, N16923, N2896, N1003);
buf BUF1 (N16929, N16928);
or OR3 (N16930, N16914, N12740, N13145);
xor XOR2 (N16931, N16921, N14286);
nand NAND2 (N16932, N16930, N8081);
xor XOR2 (N16933, N16919, N2982);
xor XOR2 (N16934, N16929, N1136);
nand NAND4 (N16935, N16910, N13325, N12078, N1791);
xor XOR2 (N16936, N16917, N9702);
nor NOR3 (N16937, N16927, N10279, N8000);
buf BUF1 (N16938, N16936);
xor XOR2 (N16939, N16937, N7584);
xor XOR2 (N16940, N16901, N13457);
nor NOR2 (N16941, N16935, N2651);
or OR4 (N16942, N16933, N780, N4672, N15591);
buf BUF1 (N16943, N16940);
xor XOR2 (N16944, N16942, N13850);
nand NAND2 (N16945, N16926, N7612);
buf BUF1 (N16946, N16945);
buf BUF1 (N16947, N16934);
xor XOR2 (N16948, N16939, N9658);
buf BUF1 (N16949, N16931);
and AND4 (N16950, N16938, N1964, N1545, N4213);
and AND4 (N16951, N16947, N5677, N16858, N16048);
nand NAND2 (N16952, N16949, N1027);
not NOT1 (N16953, N16948);
buf BUF1 (N16954, N16925);
nand NAND2 (N16955, N16941, N12162);
xor XOR2 (N16956, N16955, N6038);
buf BUF1 (N16957, N16950);
and AND4 (N16958, N16943, N16855, N6932, N3235);
nand NAND4 (N16959, N16946, N3896, N13477, N10609);
nand NAND4 (N16960, N16954, N12005, N5604, N4650);
buf BUF1 (N16961, N16953);
buf BUF1 (N16962, N16944);
xor XOR2 (N16963, N16958, N618);
not NOT1 (N16964, N16962);
and AND4 (N16965, N16957, N8765, N3084, N4719);
nand NAND4 (N16966, N16964, N11782, N13052, N9671);
and AND2 (N16967, N16951, N3255);
and AND3 (N16968, N16952, N6988, N4660);
buf BUF1 (N16969, N16959);
or OR3 (N16970, N16966, N2351, N13065);
buf BUF1 (N16971, N16965);
and AND4 (N16972, N16969, N12452, N54, N11320);
or OR3 (N16973, N16967, N2903, N14105);
and AND4 (N16974, N16972, N15311, N11199, N12842);
nor NOR2 (N16975, N16968, N9325);
buf BUF1 (N16976, N16961);
xor XOR2 (N16977, N16971, N12989);
not NOT1 (N16978, N16963);
nor NOR2 (N16979, N16978, N4228);
and AND4 (N16980, N16973, N10423, N7689, N2994);
buf BUF1 (N16981, N16974);
and AND4 (N16982, N16960, N7909, N14062, N107);
nand NAND3 (N16983, N16981, N13044, N9393);
buf BUF1 (N16984, N16980);
nand NAND4 (N16985, N16977, N16718, N16546, N9579);
xor XOR2 (N16986, N16985, N1992);
nand NAND3 (N16987, N16984, N3639, N9813);
and AND2 (N16988, N16976, N15799);
xor XOR2 (N16989, N16987, N1902);
not NOT1 (N16990, N16988);
or OR4 (N16991, N16956, N3365, N9289, N11774);
xor XOR2 (N16992, N16932, N9569);
or OR3 (N16993, N16989, N10145, N7376);
xor XOR2 (N16994, N16979, N5784);
buf BUF1 (N16995, N16983);
not NOT1 (N16996, N16975);
not NOT1 (N16997, N16996);
nor NOR4 (N16998, N16995, N248, N10869, N2327);
nor NOR4 (N16999, N16986, N14237, N11377, N14449);
or OR3 (N17000, N16993, N4970, N6383);
xor XOR2 (N17001, N17000, N13702);
and AND4 (N17002, N16992, N4808, N252, N7114);
nand NAND2 (N17003, N16999, N10073);
and AND3 (N17004, N16970, N9333, N10055);
buf BUF1 (N17005, N16994);
xor XOR2 (N17006, N17001, N14996);
and AND2 (N17007, N16997, N12497);
buf BUF1 (N17008, N17006);
or OR3 (N17009, N16998, N2719, N11370);
and AND2 (N17010, N17007, N7190);
buf BUF1 (N17011, N16991);
nand NAND3 (N17012, N17002, N1527, N13316);
buf BUF1 (N17013, N17003);
or OR2 (N17014, N16982, N11664);
or OR2 (N17015, N17005, N8755);
nand NAND4 (N17016, N17004, N4427, N9946, N5866);
nand NAND4 (N17017, N17009, N5039, N3749, N4724);
not NOT1 (N17018, N17013);
xor XOR2 (N17019, N16990, N16412);
and AND4 (N17020, N17016, N8535, N82, N5408);
or OR4 (N17021, N17012, N12427, N10589, N7842);
nand NAND3 (N17022, N17019, N10669, N2851);
and AND4 (N17023, N17015, N5684, N11150, N13847);
not NOT1 (N17024, N17010);
xor XOR2 (N17025, N17021, N12491);
nand NAND2 (N17026, N17024, N15783);
xor XOR2 (N17027, N17023, N4590);
and AND3 (N17028, N17025, N8935, N10171);
not NOT1 (N17029, N17017);
buf BUF1 (N17030, N17027);
and AND3 (N17031, N17026, N2549, N2911);
xor XOR2 (N17032, N17014, N6862);
buf BUF1 (N17033, N17030);
nor NOR2 (N17034, N17018, N11396);
nor NOR3 (N17035, N17011, N11226, N1573);
nor NOR3 (N17036, N17022, N8372, N13240);
nand NAND3 (N17037, N17031, N11678, N10997);
and AND4 (N17038, N17036, N11520, N12976, N816);
xor XOR2 (N17039, N17035, N11313);
nand NAND4 (N17040, N17039, N9559, N12810, N10313);
not NOT1 (N17041, N17033);
xor XOR2 (N17042, N17008, N16334);
nor NOR4 (N17043, N17028, N15974, N16988, N13887);
not NOT1 (N17044, N17034);
not NOT1 (N17045, N17043);
nand NAND2 (N17046, N17038, N13481);
and AND2 (N17047, N17020, N742);
and AND3 (N17048, N17041, N3135, N16940);
xor XOR2 (N17049, N17048, N2327);
and AND2 (N17050, N17049, N3126);
buf BUF1 (N17051, N17050);
or OR4 (N17052, N17040, N3821, N9436, N1871);
xor XOR2 (N17053, N17044, N12551);
not NOT1 (N17054, N17051);
or OR4 (N17055, N17046, N10409, N15241, N9848);
not NOT1 (N17056, N17032);
and AND4 (N17057, N17037, N7156, N10873, N5037);
or OR4 (N17058, N17057, N14465, N4449, N7243);
or OR2 (N17059, N17053, N1444);
or OR2 (N17060, N17029, N16746);
xor XOR2 (N17061, N17055, N14755);
or OR4 (N17062, N17052, N13931, N12456, N13857);
nor NOR3 (N17063, N17062, N9271, N3679);
nand NAND3 (N17064, N17058, N10543, N2461);
nor NOR2 (N17065, N17054, N7637);
and AND2 (N17066, N17065, N5319);
and AND3 (N17067, N17047, N1550, N2035);
not NOT1 (N17068, N17060);
buf BUF1 (N17069, N17045);
and AND2 (N17070, N17063, N16086);
or OR4 (N17071, N17070, N13319, N4700, N9627);
buf BUF1 (N17072, N17059);
and AND4 (N17073, N17066, N3163, N9228, N268);
nor NOR2 (N17074, N17067, N8170);
not NOT1 (N17075, N17071);
not NOT1 (N17076, N17061);
buf BUF1 (N17077, N17069);
buf BUF1 (N17078, N17075);
nor NOR4 (N17079, N17077, N11663, N7303, N353);
or OR3 (N17080, N17079, N13242, N12303);
and AND4 (N17081, N17068, N11780, N3643, N15532);
and AND3 (N17082, N17042, N5534, N364);
nand NAND4 (N17083, N17056, N7800, N16118, N13822);
xor XOR2 (N17084, N17082, N958);
not NOT1 (N17085, N17078);
or OR3 (N17086, N17083, N9371, N16544);
nand NAND4 (N17087, N17086, N4591, N7722, N14559);
xor XOR2 (N17088, N17080, N12354);
xor XOR2 (N17089, N17085, N7573);
nand NAND4 (N17090, N17064, N4628, N7353, N1777);
nor NOR2 (N17091, N17074, N11829);
not NOT1 (N17092, N17089);
or OR4 (N17093, N17092, N15028, N15376, N8106);
and AND4 (N17094, N17073, N15498, N9414, N13510);
xor XOR2 (N17095, N17088, N3766);
or OR2 (N17096, N17087, N14049);
nor NOR2 (N17097, N17090, N16076);
xor XOR2 (N17098, N17096, N15050);
xor XOR2 (N17099, N17091, N15041);
nand NAND4 (N17100, N17072, N13093, N13240, N15330);
buf BUF1 (N17101, N17081);
or OR3 (N17102, N17093, N722, N15626);
and AND3 (N17103, N17102, N14315, N9822);
buf BUF1 (N17104, N17094);
nor NOR2 (N17105, N17084, N6263);
or OR4 (N17106, N17103, N452, N539, N5069);
and AND3 (N17107, N17076, N4601, N1487);
buf BUF1 (N17108, N17100);
not NOT1 (N17109, N17099);
nand NAND3 (N17110, N17105, N4237, N2058);
and AND4 (N17111, N17108, N6970, N734, N2234);
not NOT1 (N17112, N17111);
and AND2 (N17113, N17098, N2646);
buf BUF1 (N17114, N17101);
or OR4 (N17115, N17106, N4324, N2193, N7999);
buf BUF1 (N17116, N17112);
and AND4 (N17117, N17095, N13438, N14068, N15608);
buf BUF1 (N17118, N17113);
nor NOR4 (N17119, N17117, N25, N8091, N11059);
or OR4 (N17120, N17119, N5343, N8883, N15142);
nand NAND2 (N17121, N17110, N6731);
xor XOR2 (N17122, N17104, N4358);
and AND4 (N17123, N17114, N3089, N8781, N10657);
buf BUF1 (N17124, N17121);
xor XOR2 (N17125, N17122, N6465);
nor NOR3 (N17126, N17123, N10234, N10749);
not NOT1 (N17127, N17124);
or OR3 (N17128, N17115, N10935, N9506);
nand NAND2 (N17129, N17127, N8247);
or OR4 (N17130, N17118, N9959, N1513, N329);
nand NAND4 (N17131, N17129, N8596, N13610, N2112);
xor XOR2 (N17132, N17116, N3479);
and AND2 (N17133, N17132, N3347);
or OR4 (N17134, N17126, N1302, N14351, N3628);
xor XOR2 (N17135, N17134, N14573);
or OR3 (N17136, N17130, N15281, N11642);
nor NOR2 (N17137, N17131, N9987);
and AND3 (N17138, N17136, N13161, N11890);
nor NOR4 (N17139, N17125, N16857, N13665, N6323);
buf BUF1 (N17140, N17128);
buf BUF1 (N17141, N17097);
and AND3 (N17142, N17135, N16812, N12747);
xor XOR2 (N17143, N17133, N8096);
not NOT1 (N17144, N17142);
or OR3 (N17145, N17120, N3870, N4349);
xor XOR2 (N17146, N17140, N431);
or OR2 (N17147, N17139, N11176);
not NOT1 (N17148, N17109);
xor XOR2 (N17149, N17144, N16625);
or OR4 (N17150, N17137, N3000, N5821, N8196);
xor XOR2 (N17151, N17148, N2752);
or OR2 (N17152, N17107, N4687);
and AND4 (N17153, N17147, N5790, N7183, N9944);
not NOT1 (N17154, N17149);
xor XOR2 (N17155, N17141, N11202);
xor XOR2 (N17156, N17151, N8810);
nand NAND4 (N17157, N17145, N2973, N15702, N7180);
not NOT1 (N17158, N17143);
or OR2 (N17159, N17150, N5208);
and AND4 (N17160, N17156, N5912, N13541, N10671);
not NOT1 (N17161, N17159);
xor XOR2 (N17162, N17152, N10915);
or OR3 (N17163, N17153, N12108, N15781);
not NOT1 (N17164, N17163);
nor NOR4 (N17165, N17155, N12697, N12814, N8310);
buf BUF1 (N17166, N17157);
and AND4 (N17167, N17146, N15578, N6515, N2633);
xor XOR2 (N17168, N17138, N7737);
buf BUF1 (N17169, N17167);
nand NAND2 (N17170, N17162, N14153);
or OR4 (N17171, N17158, N8078, N2859, N6644);
and AND3 (N17172, N17154, N10728, N10202);
and AND2 (N17173, N17164, N1568);
and AND4 (N17174, N17171, N1020, N14339, N1552);
buf BUF1 (N17175, N17169);
nand NAND4 (N17176, N17174, N451, N4390, N8927);
nand NAND3 (N17177, N17160, N12423, N4479);
nor NOR2 (N17178, N17170, N607);
and AND3 (N17179, N17173, N5347, N4650);
xor XOR2 (N17180, N17178, N15649);
buf BUF1 (N17181, N17172);
nand NAND4 (N17182, N17177, N4671, N4021, N8021);
nand NAND3 (N17183, N17165, N7342, N6372);
or OR2 (N17184, N17168, N214);
or OR2 (N17185, N17166, N4699);
not NOT1 (N17186, N17180);
nor NOR2 (N17187, N17161, N4729);
or OR3 (N17188, N17184, N7558, N9763);
nor NOR2 (N17189, N17181, N13818);
buf BUF1 (N17190, N17186);
or OR3 (N17191, N17175, N8641, N7884);
xor XOR2 (N17192, N17188, N13577);
nor NOR2 (N17193, N17191, N10652);
xor XOR2 (N17194, N17192, N14385);
buf BUF1 (N17195, N17193);
buf BUF1 (N17196, N17195);
nand NAND3 (N17197, N17182, N14787, N6561);
buf BUF1 (N17198, N17179);
or OR3 (N17199, N17187, N16314, N7036);
not NOT1 (N17200, N17196);
and AND4 (N17201, N17199, N1926, N13876, N3461);
xor XOR2 (N17202, N17176, N9690);
or OR4 (N17203, N17189, N16865, N10115, N1119);
nor NOR2 (N17204, N17190, N15816);
and AND3 (N17205, N17183, N9480, N16296);
buf BUF1 (N17206, N17201);
or OR3 (N17207, N17198, N6525, N9202);
buf BUF1 (N17208, N17185);
nand NAND4 (N17209, N17200, N12273, N8397, N6262);
or OR4 (N17210, N17206, N5407, N15011, N8367);
xor XOR2 (N17211, N17210, N12673);
buf BUF1 (N17212, N17194);
nand NAND3 (N17213, N17204, N15837, N7591);
nand NAND2 (N17214, N17207, N2077);
not NOT1 (N17215, N17209);
xor XOR2 (N17216, N17215, N16999);
xor XOR2 (N17217, N17212, N13411);
xor XOR2 (N17218, N17213, N15505);
nand NAND4 (N17219, N17217, N684, N12100, N17025);
xor XOR2 (N17220, N17211, N3137);
nor NOR3 (N17221, N17219, N1316, N10143);
xor XOR2 (N17222, N17205, N4720);
buf BUF1 (N17223, N17221);
or OR4 (N17224, N17216, N10649, N1106, N9149);
nor NOR2 (N17225, N17197, N667);
buf BUF1 (N17226, N17218);
or OR3 (N17227, N17226, N10058, N758);
nand NAND3 (N17228, N17214, N13444, N11162);
not NOT1 (N17229, N17222);
not NOT1 (N17230, N17208);
nand NAND2 (N17231, N17225, N3473);
xor XOR2 (N17232, N17220, N2656);
and AND2 (N17233, N17224, N11688);
or OR4 (N17234, N17233, N3113, N2220, N3221);
nand NAND3 (N17235, N17229, N13505, N16260);
and AND4 (N17236, N17234, N8156, N7985, N4085);
buf BUF1 (N17237, N17236);
not NOT1 (N17238, N17202);
buf BUF1 (N17239, N17231);
or OR3 (N17240, N17235, N6522, N17177);
and AND2 (N17241, N17230, N6646);
xor XOR2 (N17242, N17227, N4876);
buf BUF1 (N17243, N17223);
and AND2 (N17244, N17238, N15153);
not NOT1 (N17245, N17241);
or OR2 (N17246, N17242, N6357);
buf BUF1 (N17247, N17232);
nand NAND4 (N17248, N17240, N6412, N822, N13783);
and AND4 (N17249, N17239, N4617, N3236, N10906);
nand NAND4 (N17250, N17247, N11433, N15715, N6713);
not NOT1 (N17251, N17228);
and AND2 (N17252, N17243, N9847);
and AND2 (N17253, N17249, N15435);
nor NOR4 (N17254, N17237, N15198, N2506, N9427);
and AND4 (N17255, N17244, N13827, N353, N5352);
buf BUF1 (N17256, N17252);
nand NAND3 (N17257, N17248, N9963, N1490);
or OR4 (N17258, N17253, N2882, N11603, N1131);
nand NAND2 (N17259, N17257, N8997);
nor NOR3 (N17260, N17246, N3553, N1179);
and AND2 (N17261, N17255, N11427);
nand NAND2 (N17262, N17261, N7361);
or OR3 (N17263, N17258, N2891, N16012);
buf BUF1 (N17264, N17260);
nand NAND3 (N17265, N17263, N5743, N16109);
and AND4 (N17266, N17265, N946, N8102, N3261);
buf BUF1 (N17267, N17203);
and AND2 (N17268, N17259, N3987);
and AND4 (N17269, N17245, N9372, N9594, N12085);
not NOT1 (N17270, N17266);
not NOT1 (N17271, N17264);
nor NOR3 (N17272, N17254, N5300, N11119);
and AND4 (N17273, N17250, N16735, N11255, N9004);
and AND3 (N17274, N17256, N15041, N4538);
and AND2 (N17275, N17272, N7267);
or OR4 (N17276, N17267, N7007, N11613, N5386);
xor XOR2 (N17277, N17251, N8463);
and AND4 (N17278, N17273, N7856, N14574, N1261);
nor NOR4 (N17279, N17275, N17169, N6850, N11782);
nor NOR2 (N17280, N17278, N923);
and AND4 (N17281, N17270, N13146, N6786, N10997);
nand NAND2 (N17282, N17276, N11432);
and AND4 (N17283, N17281, N2733, N9218, N3232);
xor XOR2 (N17284, N17268, N6582);
buf BUF1 (N17285, N17274);
xor XOR2 (N17286, N17277, N9308);
nand NAND4 (N17287, N17262, N13484, N13176, N15018);
buf BUF1 (N17288, N17282);
nor NOR2 (N17289, N17285, N5082);
or OR3 (N17290, N17271, N16550, N9146);
xor XOR2 (N17291, N17286, N1984);
nand NAND2 (N17292, N17280, N1178);
buf BUF1 (N17293, N17283);
nand NAND3 (N17294, N17287, N17160, N7098);
nand NAND2 (N17295, N17292, N16092);
nor NOR4 (N17296, N17288, N17051, N6982, N10037);
or OR4 (N17297, N17284, N2325, N4017, N15277);
buf BUF1 (N17298, N17291);
nand NAND3 (N17299, N17296, N6945, N3921);
not NOT1 (N17300, N17293);
or OR2 (N17301, N17298, N2498);
and AND2 (N17302, N17279, N15597);
nor NOR4 (N17303, N17300, N13294, N6954, N1798);
nor NOR4 (N17304, N17289, N12832, N15122, N6705);
or OR3 (N17305, N17302, N5874, N8424);
nor NOR3 (N17306, N17301, N2143, N2399);
buf BUF1 (N17307, N17299);
xor XOR2 (N17308, N17303, N1855);
xor XOR2 (N17309, N17297, N9853);
nand NAND4 (N17310, N17290, N10437, N14041, N643);
and AND2 (N17311, N17309, N6248);
or OR2 (N17312, N17307, N3001);
nor NOR2 (N17313, N17311, N13396);
nor NOR2 (N17314, N17313, N1335);
not NOT1 (N17315, N17314);
buf BUF1 (N17316, N17294);
and AND3 (N17317, N17305, N11916, N11513);
and AND4 (N17318, N17308, N1572, N16780, N10936);
not NOT1 (N17319, N17304);
nand NAND2 (N17320, N17295, N9896);
buf BUF1 (N17321, N17316);
not NOT1 (N17322, N17319);
not NOT1 (N17323, N17306);
nor NOR2 (N17324, N17312, N3029);
and AND4 (N17325, N17323, N4010, N8275, N11868);
and AND2 (N17326, N17310, N1923);
or OR4 (N17327, N17320, N11988, N13299, N3328);
nand NAND3 (N17328, N17327, N10067, N9861);
nand NAND4 (N17329, N17325, N1366, N6674, N14001);
and AND3 (N17330, N17318, N10786, N5428);
nand NAND3 (N17331, N17315, N876, N17171);
buf BUF1 (N17332, N17329);
xor XOR2 (N17333, N17330, N5124);
not NOT1 (N17334, N17324);
nor NOR4 (N17335, N17269, N15263, N13356, N11258);
buf BUF1 (N17336, N17333);
or OR2 (N17337, N17332, N804);
or OR4 (N17338, N17326, N11856, N16637, N16459);
nor NOR2 (N17339, N17334, N2096);
or OR3 (N17340, N17337, N5072, N9901);
nand NAND4 (N17341, N17336, N3781, N16658, N1988);
not NOT1 (N17342, N17338);
and AND2 (N17343, N17339, N1379);
and AND4 (N17344, N17340, N738, N10728, N10670);
buf BUF1 (N17345, N17317);
nor NOR2 (N17346, N17328, N11848);
nor NOR2 (N17347, N17335, N15278);
xor XOR2 (N17348, N17321, N571);
nand NAND3 (N17349, N17345, N1264, N9613);
or OR4 (N17350, N17342, N12991, N3494, N146);
nand NAND4 (N17351, N17322, N4100, N5318, N8364);
nand NAND2 (N17352, N17350, N16820);
buf BUF1 (N17353, N17351);
not NOT1 (N17354, N17353);
nand NAND2 (N17355, N17349, N12281);
nand NAND4 (N17356, N17346, N13894, N2222, N1730);
not NOT1 (N17357, N17347);
not NOT1 (N17358, N17354);
xor XOR2 (N17359, N17356, N8312);
nor NOR4 (N17360, N17331, N642, N4914, N12619);
nand NAND2 (N17361, N17343, N9533);
nand NAND2 (N17362, N17355, N3130);
and AND2 (N17363, N17360, N719);
buf BUF1 (N17364, N17363);
and AND3 (N17365, N17341, N8970, N12648);
or OR2 (N17366, N17358, N1371);
nand NAND2 (N17367, N17359, N3687);
not NOT1 (N17368, N17367);
nor NOR2 (N17369, N17366, N9222);
and AND3 (N17370, N17368, N7420, N3170);
xor XOR2 (N17371, N17365, N10843);
not NOT1 (N17372, N17362);
xor XOR2 (N17373, N17369, N2175);
nand NAND4 (N17374, N17348, N12531, N1377, N7980);
buf BUF1 (N17375, N17374);
not NOT1 (N17376, N17372);
nor NOR3 (N17377, N17364, N13778, N14539);
xor XOR2 (N17378, N17376, N16924);
xor XOR2 (N17379, N17370, N2541);
xor XOR2 (N17380, N17344, N9777);
and AND3 (N17381, N17380, N12400, N113);
buf BUF1 (N17382, N17379);
buf BUF1 (N17383, N17381);
nor NOR4 (N17384, N17352, N4571, N15350, N6174);
xor XOR2 (N17385, N17377, N7487);
nand NAND4 (N17386, N17375, N8485, N10429, N3450);
or OR2 (N17387, N17386, N3119);
buf BUF1 (N17388, N17371);
xor XOR2 (N17389, N17382, N13057);
nor NOR4 (N17390, N17361, N15560, N7739, N10691);
not NOT1 (N17391, N17388);
not NOT1 (N17392, N17389);
not NOT1 (N17393, N17392);
nor NOR3 (N17394, N17387, N2042, N13889);
and AND3 (N17395, N17391, N12671, N4942);
and AND4 (N17396, N17357, N5725, N4755, N14530);
nand NAND4 (N17397, N17383, N4017, N5298, N10961);
nor NOR2 (N17398, N17378, N17235);
xor XOR2 (N17399, N17390, N13120);
and AND4 (N17400, N17384, N6969, N9465, N7051);
and AND3 (N17401, N17397, N13505, N17230);
buf BUF1 (N17402, N17393);
not NOT1 (N17403, N17373);
not NOT1 (N17404, N17385);
nand NAND3 (N17405, N17404, N14925, N890);
nor NOR4 (N17406, N17399, N8940, N14828, N6877);
nand NAND3 (N17407, N17402, N470, N10304);
or OR3 (N17408, N17403, N13908, N4243);
nand NAND4 (N17409, N17395, N3248, N7251, N14861);
or OR3 (N17410, N17408, N10233, N16131);
buf BUF1 (N17411, N17394);
buf BUF1 (N17412, N17411);
nor NOR4 (N17413, N17407, N8900, N10888, N16553);
and AND3 (N17414, N17398, N569, N2922);
buf BUF1 (N17415, N17414);
nand NAND4 (N17416, N17410, N13598, N13725, N6427);
and AND4 (N17417, N17396, N649, N2529, N7477);
buf BUF1 (N17418, N17409);
and AND4 (N17419, N17405, N10655, N13304, N11618);
buf BUF1 (N17420, N17416);
xor XOR2 (N17421, N17420, N12951);
and AND2 (N17422, N17406, N7366);
and AND4 (N17423, N17401, N7654, N9488, N9226);
nor NOR3 (N17424, N17421, N15661, N4884);
nand NAND2 (N17425, N17419, N13762);
buf BUF1 (N17426, N17413);
not NOT1 (N17427, N17412);
nand NAND2 (N17428, N17422, N2640);
not NOT1 (N17429, N17417);
nand NAND2 (N17430, N17423, N6505);
buf BUF1 (N17431, N17429);
and AND2 (N17432, N17427, N11421);
buf BUF1 (N17433, N17424);
xor XOR2 (N17434, N17432, N5038);
buf BUF1 (N17435, N17428);
nand NAND2 (N17436, N17434, N14376);
or OR2 (N17437, N17431, N14120);
not NOT1 (N17438, N17437);
buf BUF1 (N17439, N17430);
not NOT1 (N17440, N17433);
or OR2 (N17441, N17435, N12379);
and AND3 (N17442, N17436, N8850, N3444);
buf BUF1 (N17443, N17441);
not NOT1 (N17444, N17400);
nor NOR2 (N17445, N17442, N8035);
not NOT1 (N17446, N17418);
or OR2 (N17447, N17425, N12379);
or OR4 (N17448, N17426, N11014, N3023, N13836);
and AND3 (N17449, N17439, N12355, N7545);
xor XOR2 (N17450, N17446, N13090);
nand NAND3 (N17451, N17415, N5692, N3308);
nor NOR2 (N17452, N17445, N3697);
or OR2 (N17453, N17448, N15559);
nand NAND3 (N17454, N17450, N10239, N6099);
and AND4 (N17455, N17453, N12656, N3813, N12411);
nand NAND3 (N17456, N17454, N3529, N12387);
and AND3 (N17457, N17438, N11903, N2131);
nand NAND2 (N17458, N17444, N7292);
not NOT1 (N17459, N17457);
xor XOR2 (N17460, N17447, N6507);
buf BUF1 (N17461, N17443);
buf BUF1 (N17462, N17460);
xor XOR2 (N17463, N17449, N10091);
not NOT1 (N17464, N17462);
buf BUF1 (N17465, N17461);
nand NAND2 (N17466, N17459, N14586);
or OR2 (N17467, N17451, N9966);
nor NOR3 (N17468, N17464, N17092, N4560);
and AND2 (N17469, N17465, N6540);
xor XOR2 (N17470, N17456, N13673);
nor NOR2 (N17471, N17458, N6300);
and AND3 (N17472, N17467, N4914, N3739);
not NOT1 (N17473, N17471);
and AND2 (N17474, N17455, N1525);
nand NAND4 (N17475, N17468, N13573, N3736, N17050);
and AND4 (N17476, N17472, N10058, N14119, N1677);
or OR3 (N17477, N17452, N6934, N1618);
or OR3 (N17478, N17477, N5142, N17199);
buf BUF1 (N17479, N17470);
nor NOR4 (N17480, N17475, N16162, N5066, N11683);
nor NOR3 (N17481, N17476, N7134, N17174);
not NOT1 (N17482, N17463);
not NOT1 (N17483, N17481);
and AND3 (N17484, N17480, N6499, N2667);
not NOT1 (N17485, N17466);
nand NAND4 (N17486, N17482, N17075, N11459, N5074);
not NOT1 (N17487, N17469);
xor XOR2 (N17488, N17483, N4325);
xor XOR2 (N17489, N17440, N2244);
nand NAND4 (N17490, N17474, N16888, N3999, N609);
not NOT1 (N17491, N17487);
or OR3 (N17492, N17491, N16932, N15655);
nor NOR4 (N17493, N17489, N7931, N8226, N3884);
nor NOR2 (N17494, N17484, N12965);
or OR3 (N17495, N17473, N16747, N13461);
nand NAND4 (N17496, N17478, N1109, N15015, N11115);
not NOT1 (N17497, N17479);
xor XOR2 (N17498, N17494, N13131);
not NOT1 (N17499, N17496);
xor XOR2 (N17500, N17499, N7308);
buf BUF1 (N17501, N17493);
buf BUF1 (N17502, N17500);
xor XOR2 (N17503, N17497, N4169);
buf BUF1 (N17504, N17503);
buf BUF1 (N17505, N17485);
nor NOR3 (N17506, N17504, N5989, N15584);
nor NOR3 (N17507, N17486, N16920, N14784);
nand NAND2 (N17508, N17490, N3527);
nand NAND4 (N17509, N17501, N12488, N7706, N14888);
buf BUF1 (N17510, N17502);
buf BUF1 (N17511, N17488);
or OR3 (N17512, N17495, N492, N12489);
buf BUF1 (N17513, N17506);
nor NOR2 (N17514, N17512, N13626);
xor XOR2 (N17515, N17514, N2739);
nor NOR2 (N17516, N17510, N9701);
or OR3 (N17517, N17492, N16834, N7775);
or OR2 (N17518, N17509, N14220);
nor NOR4 (N17519, N17505, N1093, N2070, N3483);
not NOT1 (N17520, N17511);
xor XOR2 (N17521, N17516, N14433);
xor XOR2 (N17522, N17513, N1609);
nand NAND2 (N17523, N17520, N6012);
xor XOR2 (N17524, N17522, N11622);
nand NAND4 (N17525, N17508, N15816, N15358, N4750);
xor XOR2 (N17526, N17521, N11818);
nor NOR2 (N17527, N17523, N15965);
not NOT1 (N17528, N17527);
buf BUF1 (N17529, N17515);
xor XOR2 (N17530, N17528, N7188);
xor XOR2 (N17531, N17526, N9964);
not NOT1 (N17532, N17529);
nand NAND4 (N17533, N17518, N4725, N9266, N17107);
buf BUF1 (N17534, N17519);
and AND2 (N17535, N17524, N14836);
not NOT1 (N17536, N17531);
xor XOR2 (N17537, N17498, N1344);
or OR2 (N17538, N17533, N5478);
nand NAND3 (N17539, N17517, N3804, N8448);
nor NOR3 (N17540, N17525, N1022, N7409);
not NOT1 (N17541, N17534);
xor XOR2 (N17542, N17541, N15689);
xor XOR2 (N17543, N17542, N14889);
not NOT1 (N17544, N17540);
or OR3 (N17545, N17535, N8450, N6604);
xor XOR2 (N17546, N17539, N4103);
or OR4 (N17547, N17546, N14264, N15967, N6737);
not NOT1 (N17548, N17545);
xor XOR2 (N17549, N17548, N6458);
nor NOR2 (N17550, N17544, N222);
xor XOR2 (N17551, N17530, N6402);
nand NAND3 (N17552, N17538, N2944, N2520);
and AND2 (N17553, N17547, N6258);
xor XOR2 (N17554, N17553, N6844);
not NOT1 (N17555, N17543);
not NOT1 (N17556, N17550);
buf BUF1 (N17557, N17551);
xor XOR2 (N17558, N17532, N16207);
and AND4 (N17559, N17556, N733, N10777, N11382);
nor NOR3 (N17560, N17507, N13226, N15882);
nand NAND2 (N17561, N17537, N56);
or OR3 (N17562, N17559, N191, N5043);
xor XOR2 (N17563, N17552, N296);
nand NAND2 (N17564, N17554, N15005);
and AND2 (N17565, N17558, N15365);
and AND2 (N17566, N17536, N3538);
or OR2 (N17567, N17566, N9431);
nand NAND3 (N17568, N17557, N16437, N3669);
or OR2 (N17569, N17568, N12089);
xor XOR2 (N17570, N17567, N2692);
nor NOR3 (N17571, N17563, N14590, N14847);
not NOT1 (N17572, N17561);
nor NOR3 (N17573, N17572, N7860, N14238);
or OR4 (N17574, N17573, N2583, N12527, N1410);
or OR2 (N17575, N17574, N12297);
not NOT1 (N17576, N17549);
xor XOR2 (N17577, N17571, N14030);
and AND2 (N17578, N17575, N4318);
buf BUF1 (N17579, N17565);
or OR3 (N17580, N17579, N9581, N4039);
nor NOR2 (N17581, N17577, N15084);
nor NOR2 (N17582, N17569, N16650);
or OR3 (N17583, N17570, N36, N14040);
nand NAND4 (N17584, N17578, N14365, N8830, N14584);
and AND3 (N17585, N17582, N5548, N6606);
or OR4 (N17586, N17581, N16476, N6687, N1058);
nor NOR2 (N17587, N17560, N9452);
xor XOR2 (N17588, N17580, N14175);
buf BUF1 (N17589, N17564);
and AND4 (N17590, N17584, N3352, N10987, N9778);
nand NAND3 (N17591, N17589, N11763, N5608);
xor XOR2 (N17592, N17555, N11421);
nor NOR2 (N17593, N17591, N7436);
nand NAND3 (N17594, N17592, N14213, N557);
and AND2 (N17595, N17594, N16440);
buf BUF1 (N17596, N17583);
buf BUF1 (N17597, N17590);
and AND4 (N17598, N17587, N3835, N15137, N5878);
xor XOR2 (N17599, N17562, N10299);
not NOT1 (N17600, N17595);
nor NOR2 (N17601, N17593, N10190);
xor XOR2 (N17602, N17586, N1529);
xor XOR2 (N17603, N17601, N12608);
nor NOR4 (N17604, N17603, N10299, N1760, N691);
or OR4 (N17605, N17588, N1943, N267, N12436);
xor XOR2 (N17606, N17604, N5569);
or OR4 (N17607, N17600, N5768, N14920, N1872);
not NOT1 (N17608, N17596);
nand NAND2 (N17609, N17606, N14917);
nand NAND3 (N17610, N17599, N3672, N5463);
and AND2 (N17611, N17605, N1282);
or OR4 (N17612, N17611, N3719, N5816, N10538);
buf BUF1 (N17613, N17585);
not NOT1 (N17614, N17612);
nor NOR3 (N17615, N17613, N10183, N3858);
nor NOR4 (N17616, N17615, N2724, N13135, N1628);
or OR3 (N17617, N17610, N13366, N11869);
not NOT1 (N17618, N17598);
nand NAND4 (N17619, N17616, N14259, N16724, N13960);
not NOT1 (N17620, N17602);
or OR3 (N17621, N17614, N6878, N3124);
or OR3 (N17622, N17607, N9000, N11264);
and AND4 (N17623, N17618, N1456, N5694, N12389);
and AND2 (N17624, N17620, N13454);
nor NOR2 (N17625, N17576, N9899);
or OR2 (N17626, N17617, N3164);
or OR2 (N17627, N17608, N11741);
xor XOR2 (N17628, N17597, N15253);
xor XOR2 (N17629, N17623, N5142);
or OR4 (N17630, N17627, N2841, N2775, N485);
and AND3 (N17631, N17624, N7882, N7182);
or OR4 (N17632, N17631, N4017, N4704, N7020);
or OR4 (N17633, N17630, N16028, N10836, N3873);
xor XOR2 (N17634, N17628, N6840);
buf BUF1 (N17635, N17632);
nand NAND4 (N17636, N17619, N4333, N9210, N1989);
nor NOR3 (N17637, N17625, N16327, N2924);
or OR4 (N17638, N17622, N13019, N8436, N15786);
and AND2 (N17639, N17629, N444);
xor XOR2 (N17640, N17635, N14289);
not NOT1 (N17641, N17621);
and AND4 (N17642, N17637, N11613, N3849, N2976);
or OR4 (N17643, N17642, N12566, N6664, N17469);
or OR4 (N17644, N17639, N8504, N1123, N10983);
xor XOR2 (N17645, N17644, N8259);
and AND4 (N17646, N17634, N718, N2732, N15234);
nor NOR3 (N17647, N17646, N2351, N3740);
and AND2 (N17648, N17647, N9665);
buf BUF1 (N17649, N17640);
or OR2 (N17650, N17609, N10129);
not NOT1 (N17651, N17649);
and AND3 (N17652, N17645, N13485, N6888);
buf BUF1 (N17653, N17652);
not NOT1 (N17654, N17636);
xor XOR2 (N17655, N17633, N4791);
or OR2 (N17656, N17653, N6020);
buf BUF1 (N17657, N17656);
buf BUF1 (N17658, N17655);
nor NOR2 (N17659, N17641, N10472);
xor XOR2 (N17660, N17659, N4232);
buf BUF1 (N17661, N17658);
xor XOR2 (N17662, N17638, N14605);
nand NAND2 (N17663, N17662, N12630);
nand NAND4 (N17664, N17626, N10950, N13538, N892);
not NOT1 (N17665, N17663);
xor XOR2 (N17666, N17650, N12140);
nor NOR3 (N17667, N17648, N12004, N2169);
or OR3 (N17668, N17657, N6112, N10839);
nand NAND3 (N17669, N17664, N8470, N8610);
not NOT1 (N17670, N17669);
nand NAND3 (N17671, N17665, N16916, N14078);
or OR2 (N17672, N17660, N16620);
and AND2 (N17673, N17671, N1081);
not NOT1 (N17674, N17643);
or OR4 (N17675, N17674, N11755, N7861, N15749);
xor XOR2 (N17676, N17661, N1458);
or OR3 (N17677, N17672, N7383, N7951);
not NOT1 (N17678, N17651);
buf BUF1 (N17679, N17678);
not NOT1 (N17680, N17677);
not NOT1 (N17681, N17670);
nor NOR2 (N17682, N17654, N10169);
xor XOR2 (N17683, N17680, N6891);
not NOT1 (N17684, N17666);
buf BUF1 (N17685, N17679);
nand NAND4 (N17686, N17675, N11736, N8657, N7728);
xor XOR2 (N17687, N17686, N428);
nand NAND3 (N17688, N17667, N16218, N7431);
nor NOR2 (N17689, N17676, N14408);
buf BUF1 (N17690, N17688);
nor NOR2 (N17691, N17673, N14736);
nor NOR4 (N17692, N17690, N4855, N12597, N379);
not NOT1 (N17693, N17689);
nor NOR3 (N17694, N17668, N5065, N13416);
nor NOR3 (N17695, N17681, N14462, N6642);
nand NAND3 (N17696, N17684, N11708, N7786);
xor XOR2 (N17697, N17696, N9849);
nor NOR2 (N17698, N17682, N7783);
or OR4 (N17699, N17695, N9754, N15611, N5691);
and AND2 (N17700, N17692, N15024);
buf BUF1 (N17701, N17697);
or OR4 (N17702, N17687, N15614, N17073, N9829);
xor XOR2 (N17703, N17698, N14488);
not NOT1 (N17704, N17685);
buf BUF1 (N17705, N17699);
and AND3 (N17706, N17705, N1323, N14551);
not NOT1 (N17707, N17693);
and AND2 (N17708, N17694, N6308);
not NOT1 (N17709, N17703);
or OR2 (N17710, N17702, N2588);
buf BUF1 (N17711, N17710);
and AND4 (N17712, N17706, N12847, N6725, N4992);
not NOT1 (N17713, N17708);
nand NAND3 (N17714, N17713, N413, N3623);
xor XOR2 (N17715, N17704, N16202);
or OR3 (N17716, N17711, N6087, N2780);
or OR3 (N17717, N17701, N8025, N6958);
nand NAND4 (N17718, N17709, N1672, N1337, N10613);
not NOT1 (N17719, N17715);
not NOT1 (N17720, N17691);
and AND2 (N17721, N17718, N3766);
nor NOR4 (N17722, N17683, N881, N11221, N17566);
buf BUF1 (N17723, N17707);
not NOT1 (N17724, N17712);
xor XOR2 (N17725, N17721, N1091);
buf BUF1 (N17726, N17717);
not NOT1 (N17727, N17722);
nand NAND4 (N17728, N17720, N4148, N4745, N17098);
not NOT1 (N17729, N17725);
nor NOR3 (N17730, N17716, N9223, N8379);
not NOT1 (N17731, N17724);
xor XOR2 (N17732, N17727, N12239);
xor XOR2 (N17733, N17714, N5437);
xor XOR2 (N17734, N17729, N11094);
nor NOR3 (N17735, N17731, N7900, N15216);
and AND2 (N17736, N17726, N2052);
and AND4 (N17737, N17733, N13694, N5445, N13310);
and AND4 (N17738, N17734, N4389, N9274, N8320);
nand NAND2 (N17739, N17719, N15348);
xor XOR2 (N17740, N17728, N8172);
nor NOR2 (N17741, N17738, N7263);
and AND3 (N17742, N17739, N9790, N13992);
not NOT1 (N17743, N17741);
nor NOR4 (N17744, N17735, N10919, N10932, N4540);
nand NAND4 (N17745, N17700, N13259, N14299, N6537);
and AND2 (N17746, N17730, N1804);
buf BUF1 (N17747, N17736);
buf BUF1 (N17748, N17744);
buf BUF1 (N17749, N17740);
nor NOR4 (N17750, N17723, N1782, N7836, N10819);
nand NAND4 (N17751, N17745, N14750, N1707, N8918);
buf BUF1 (N17752, N17743);
nand NAND3 (N17753, N17749, N8731, N14184);
nor NOR4 (N17754, N17753, N380, N15434, N12056);
buf BUF1 (N17755, N17752);
nand NAND3 (N17756, N17754, N5914, N668);
nor NOR2 (N17757, N17748, N5513);
and AND4 (N17758, N17732, N1099, N4675, N9290);
nand NAND4 (N17759, N17750, N3853, N7866, N13422);
not NOT1 (N17760, N17737);
not NOT1 (N17761, N17746);
and AND4 (N17762, N17751, N11834, N2838, N4458);
and AND3 (N17763, N17756, N1620, N4653);
not NOT1 (N17764, N17763);
nand NAND2 (N17765, N17760, N15604);
or OR4 (N17766, N17759, N7956, N2417, N3229);
and AND3 (N17767, N17766, N8682, N6892);
xor XOR2 (N17768, N17765, N779);
nor NOR3 (N17769, N17768, N12262, N13026);
nand NAND2 (N17770, N17764, N15096);
nand NAND4 (N17771, N17770, N3508, N9133, N4886);
buf BUF1 (N17772, N17767);
or OR4 (N17773, N17742, N12971, N1407, N17548);
xor XOR2 (N17774, N17755, N13580);
buf BUF1 (N17775, N17769);
or OR2 (N17776, N17762, N2379);
nor NOR4 (N17777, N17761, N12501, N2958, N6739);
or OR3 (N17778, N17773, N13555, N992);
not NOT1 (N17779, N17771);
or OR2 (N17780, N17757, N10861);
and AND4 (N17781, N17778, N2127, N9298, N14308);
not NOT1 (N17782, N17747);
xor XOR2 (N17783, N17780, N699);
not NOT1 (N17784, N17772);
not NOT1 (N17785, N17758);
buf BUF1 (N17786, N17777);
xor XOR2 (N17787, N17786, N1854);
or OR3 (N17788, N17775, N10515, N1974);
xor XOR2 (N17789, N17785, N6596);
xor XOR2 (N17790, N17781, N13576);
nand NAND3 (N17791, N17783, N5432, N10828);
buf BUF1 (N17792, N17776);
or OR3 (N17793, N17788, N3636, N6307);
and AND4 (N17794, N17791, N11100, N5702, N17271);
or OR4 (N17795, N17793, N11882, N3987, N2698);
buf BUF1 (N17796, N17789);
not NOT1 (N17797, N17796);
nor NOR2 (N17798, N17794, N16465);
not NOT1 (N17799, N17792);
or OR3 (N17800, N17787, N11992, N7073);
and AND3 (N17801, N17797, N9418, N8168);
xor XOR2 (N17802, N17801, N2897);
nand NAND2 (N17803, N17799, N9300);
not NOT1 (N17804, N17800);
buf BUF1 (N17805, N17802);
nand NAND4 (N17806, N17803, N5556, N6631, N3028);
or OR4 (N17807, N17784, N3662, N279, N4838);
nor NOR4 (N17808, N17782, N6469, N17365, N13962);
or OR3 (N17809, N17790, N8503, N12991);
xor XOR2 (N17810, N17779, N3271);
nor NOR4 (N17811, N17805, N16468, N4911, N9447);
xor XOR2 (N17812, N17808, N9933);
and AND4 (N17813, N17810, N15680, N11806, N9135);
xor XOR2 (N17814, N17813, N1832);
nand NAND3 (N17815, N17798, N14813, N2039);
buf BUF1 (N17816, N17795);
nand NAND4 (N17817, N17774, N2574, N2066, N2227);
nor NOR4 (N17818, N17807, N16015, N4838, N13601);
and AND2 (N17819, N17815, N12727);
not NOT1 (N17820, N17809);
not NOT1 (N17821, N17811);
and AND2 (N17822, N17819, N9524);
xor XOR2 (N17823, N17820, N4360);
xor XOR2 (N17824, N17812, N14709);
or OR3 (N17825, N17817, N9990, N8310);
buf BUF1 (N17826, N17823);
buf BUF1 (N17827, N17818);
nand NAND2 (N17828, N17816, N8565);
or OR3 (N17829, N17828, N16210, N13116);
not NOT1 (N17830, N17822);
buf BUF1 (N17831, N17826);
or OR4 (N17832, N17831, N12103, N15665, N17657);
and AND3 (N17833, N17821, N10154, N6775);
nor NOR4 (N17834, N17806, N6292, N1116, N14148);
buf BUF1 (N17835, N17834);
and AND3 (N17836, N17833, N8953, N17316);
xor XOR2 (N17837, N17804, N92);
and AND4 (N17838, N17837, N14849, N3653, N2555);
and AND3 (N17839, N17829, N5965, N751);
or OR2 (N17840, N17832, N1213);
not NOT1 (N17841, N17827);
nor NOR4 (N17842, N17841, N5144, N11490, N8004);
nand NAND4 (N17843, N17836, N14768, N4885, N5580);
nor NOR3 (N17844, N17839, N4255, N11419);
or OR4 (N17845, N17830, N1677, N2819, N7860);
nor NOR4 (N17846, N17814, N12586, N10575, N11264);
and AND2 (N17847, N17844, N10952);
xor XOR2 (N17848, N17824, N15380);
nor NOR4 (N17849, N17843, N3241, N753, N2166);
xor XOR2 (N17850, N17846, N9132);
buf BUF1 (N17851, N17848);
not NOT1 (N17852, N17842);
not NOT1 (N17853, N17847);
buf BUF1 (N17854, N17852);
or OR4 (N17855, N17849, N16290, N3250, N2768);
xor XOR2 (N17856, N17838, N6000);
nand NAND4 (N17857, N17850, N13927, N16196, N2040);
nand NAND3 (N17858, N17851, N13907, N16497);
nand NAND3 (N17859, N17854, N17798, N2973);
not NOT1 (N17860, N17853);
nand NAND4 (N17861, N17855, N7008, N14512, N8856);
not NOT1 (N17862, N17825);
buf BUF1 (N17863, N17857);
and AND2 (N17864, N17861, N243);
buf BUF1 (N17865, N17840);
or OR3 (N17866, N17845, N4640, N17771);
and AND3 (N17867, N17865, N11432, N8341);
or OR3 (N17868, N17858, N9697, N15060);
and AND4 (N17869, N17835, N17088, N4844, N4974);
xor XOR2 (N17870, N17868, N2410);
buf BUF1 (N17871, N17866);
buf BUF1 (N17872, N17869);
or OR2 (N17873, N17871, N901);
xor XOR2 (N17874, N17864, N3066);
or OR4 (N17875, N17859, N10796, N5770, N17081);
buf BUF1 (N17876, N17872);
xor XOR2 (N17877, N17856, N119);
nor NOR3 (N17878, N17862, N363, N7074);
nor NOR2 (N17879, N17874, N12260);
or OR2 (N17880, N17876, N7422);
nor NOR2 (N17881, N17875, N1691);
nor NOR3 (N17882, N17877, N4372, N12112);
buf BUF1 (N17883, N17860);
nand NAND4 (N17884, N17883, N5037, N17267, N4923);
nand NAND2 (N17885, N17880, N17175);
not NOT1 (N17886, N17879);
buf BUF1 (N17887, N17881);
not NOT1 (N17888, N17873);
not NOT1 (N17889, N17884);
and AND3 (N17890, N17886, N17888, N3376);
not NOT1 (N17891, N3047);
nand NAND4 (N17892, N17889, N13847, N5588, N9949);
buf BUF1 (N17893, N17878);
nor NOR2 (N17894, N17891, N3933);
and AND2 (N17895, N17890, N16219);
xor XOR2 (N17896, N17867, N231);
nor NOR3 (N17897, N17896, N6847, N8745);
nor NOR4 (N17898, N17897, N16916, N255, N3131);
and AND3 (N17899, N17870, N15555, N6601);
not NOT1 (N17900, N17899);
or OR3 (N17901, N17898, N13893, N5966);
nand NAND2 (N17902, N17863, N10244);
nor NOR2 (N17903, N17893, N12967);
or OR3 (N17904, N17901, N7428, N13174);
not NOT1 (N17905, N17902);
nor NOR2 (N17906, N17895, N16387);
nor NOR3 (N17907, N17903, N5301, N13606);
and AND2 (N17908, N17905, N2389);
and AND2 (N17909, N17907, N14455);
nor NOR4 (N17910, N17906, N13020, N3831, N6996);
and AND2 (N17911, N17900, N1454);
xor XOR2 (N17912, N17882, N17316);
nand NAND2 (N17913, N17894, N15211);
buf BUF1 (N17914, N17885);
buf BUF1 (N17915, N17908);
xor XOR2 (N17916, N17913, N8842);
xor XOR2 (N17917, N17912, N5423);
nor NOR4 (N17918, N17916, N1024, N2998, N16048);
nand NAND4 (N17919, N17892, N13935, N3191, N14490);
and AND4 (N17920, N17914, N17162, N12847, N14302);
nor NOR2 (N17921, N17917, N9700);
nor NOR3 (N17922, N17910, N285, N7700);
nand NAND2 (N17923, N17911, N5265);
xor XOR2 (N17924, N17920, N13147);
or OR4 (N17925, N17923, N15889, N4231, N16133);
not NOT1 (N17926, N17918);
not NOT1 (N17927, N17926);
buf BUF1 (N17928, N17915);
buf BUF1 (N17929, N17924);
buf BUF1 (N17930, N17925);
or OR4 (N17931, N17929, N9403, N8689, N9380);
or OR2 (N17932, N17921, N14526);
or OR2 (N17933, N17928, N10454);
and AND2 (N17934, N17922, N15014);
nand NAND4 (N17935, N17934, N3531, N3622, N5635);
not NOT1 (N17936, N17887);
buf BUF1 (N17937, N17931);
xor XOR2 (N17938, N17930, N11465);
not NOT1 (N17939, N17937);
and AND4 (N17940, N17932, N17900, N4352, N8960);
nand NAND3 (N17941, N17904, N949, N2124);
or OR4 (N17942, N17935, N10083, N1567, N1710);
nor NOR4 (N17943, N17933, N7589, N14984, N8783);
buf BUF1 (N17944, N17940);
nor NOR2 (N17945, N17941, N2211);
nor NOR2 (N17946, N17944, N12803);
or OR3 (N17947, N17927, N11113, N6029);
nand NAND2 (N17948, N17936, N15815);
not NOT1 (N17949, N17943);
nor NOR3 (N17950, N17938, N7, N9769);
nand NAND4 (N17951, N17945, N14444, N10433, N4687);
or OR2 (N17952, N17919, N14780);
not NOT1 (N17953, N17939);
and AND4 (N17954, N17950, N2349, N10575, N5298);
xor XOR2 (N17955, N17948, N10706);
and AND4 (N17956, N17955, N13251, N14662, N12977);
nor NOR3 (N17957, N17947, N13033, N9991);
nand NAND3 (N17958, N17952, N15210, N3146);
buf BUF1 (N17959, N17953);
buf BUF1 (N17960, N17942);
and AND3 (N17961, N17949, N489, N467);
buf BUF1 (N17962, N17946);
and AND2 (N17963, N17954, N8503);
nor NOR2 (N17964, N17951, N866);
or OR3 (N17965, N17957, N17876, N15442);
and AND2 (N17966, N17964, N4234);
nor NOR4 (N17967, N17959, N565, N8106, N2039);
and AND2 (N17968, N17909, N16464);
xor XOR2 (N17969, N17956, N7578);
buf BUF1 (N17970, N17966);
and AND2 (N17971, N17958, N10519);
and AND4 (N17972, N17963, N17650, N8821, N3717);
not NOT1 (N17973, N17962);
and AND3 (N17974, N17961, N9439, N14531);
xor XOR2 (N17975, N17974, N5458);
or OR4 (N17976, N17967, N7458, N9191, N8277);
xor XOR2 (N17977, N17973, N13000);
xor XOR2 (N17978, N17972, N3775);
not NOT1 (N17979, N17965);
xor XOR2 (N17980, N17977, N16840);
buf BUF1 (N17981, N17960);
buf BUF1 (N17982, N17980);
or OR3 (N17983, N17979, N6974, N4165);
or OR2 (N17984, N17981, N14797);
or OR4 (N17985, N17976, N196, N8861, N7388);
nand NAND4 (N17986, N17985, N8986, N11454, N859);
not NOT1 (N17987, N17971);
and AND2 (N17988, N17984, N5600);
not NOT1 (N17989, N17983);
and AND2 (N17990, N17982, N15416);
xor XOR2 (N17991, N17989, N13369);
xor XOR2 (N17992, N17988, N2779);
buf BUF1 (N17993, N17987);
buf BUF1 (N17994, N17970);
xor XOR2 (N17995, N17990, N12057);
xor XOR2 (N17996, N17993, N8623);
nand NAND3 (N17997, N17995, N8664, N13324);
nand NAND3 (N17998, N17969, N4158, N4264);
buf BUF1 (N17999, N17986);
nor NOR2 (N18000, N17978, N2607);
not NOT1 (N18001, N17968);
nor NOR2 (N18002, N17996, N16610);
nor NOR3 (N18003, N17975, N10168, N7295);
xor XOR2 (N18004, N17991, N13998);
and AND4 (N18005, N18004, N11792, N9642, N8952);
nand NAND3 (N18006, N17998, N10999, N12396);
not NOT1 (N18007, N17997);
and AND2 (N18008, N18005, N2856);
and AND2 (N18009, N18003, N361);
or OR3 (N18010, N18007, N16468, N2719);
buf BUF1 (N18011, N18000);
and AND3 (N18012, N17992, N11279, N7712);
xor XOR2 (N18013, N18002, N8247);
nand NAND2 (N18014, N18011, N16550);
nand NAND3 (N18015, N17999, N325, N2802);
nand NAND2 (N18016, N18009, N8303);
nor NOR3 (N18017, N17994, N15543, N14309);
nor NOR2 (N18018, N18014, N824);
nor NOR2 (N18019, N18017, N16450);
not NOT1 (N18020, N18001);
nand NAND2 (N18021, N18020, N5138);
nor NOR2 (N18022, N18016, N2838);
buf BUF1 (N18023, N18015);
or OR3 (N18024, N18021, N5231, N16656);
or OR2 (N18025, N18024, N7150);
not NOT1 (N18026, N18013);
or OR4 (N18027, N18025, N3848, N7820, N6814);
nand NAND4 (N18028, N18019, N17800, N13769, N5258);
buf BUF1 (N18029, N18023);
and AND3 (N18030, N18026, N10032, N6901);
xor XOR2 (N18031, N18029, N13812);
and AND2 (N18032, N18008, N10250);
xor XOR2 (N18033, N18028, N688);
xor XOR2 (N18034, N18031, N14513);
xor XOR2 (N18035, N18030, N11976);
not NOT1 (N18036, N18027);
nand NAND4 (N18037, N18010, N2255, N10082, N12994);
and AND2 (N18038, N18037, N2603);
xor XOR2 (N18039, N18036, N14818);
or OR2 (N18040, N18018, N11838);
or OR4 (N18041, N18033, N16847, N683, N16024);
nor NOR3 (N18042, N18034, N8587, N7577);
not NOT1 (N18043, N18040);
or OR3 (N18044, N18032, N14981, N4194);
nor NOR3 (N18045, N18041, N14655, N15453);
xor XOR2 (N18046, N18012, N881);
or OR4 (N18047, N18038, N14633, N6680, N2567);
not NOT1 (N18048, N18045);
xor XOR2 (N18049, N18022, N16952);
buf BUF1 (N18050, N18042);
nand NAND2 (N18051, N18044, N9131);
xor XOR2 (N18052, N18047, N10821);
nor NOR4 (N18053, N18050, N10170, N15403, N6670);
nor NOR4 (N18054, N18046, N8971, N15025, N13693);
xor XOR2 (N18055, N18049, N3150);
xor XOR2 (N18056, N18035, N15117);
xor XOR2 (N18057, N18054, N3299);
xor XOR2 (N18058, N18048, N14200);
xor XOR2 (N18059, N18052, N16257);
and AND4 (N18060, N18055, N1318, N7584, N5737);
nor NOR2 (N18061, N18057, N1766);
buf BUF1 (N18062, N18058);
or OR2 (N18063, N18060, N1960);
xor XOR2 (N18064, N18053, N6273);
nand NAND4 (N18065, N18061, N8431, N459, N332);
not NOT1 (N18066, N18051);
nor NOR2 (N18067, N18063, N2885);
or OR2 (N18068, N18062, N18055);
nand NAND2 (N18069, N18066, N11529);
xor XOR2 (N18070, N18056, N13739);
nand NAND2 (N18071, N18006, N15368);
nor NOR3 (N18072, N18039, N2780, N740);
buf BUF1 (N18073, N18072);
nand NAND3 (N18074, N18069, N16443, N5526);
nand NAND4 (N18075, N18065, N17554, N17601, N8645);
not NOT1 (N18076, N18073);
nor NOR3 (N18077, N18064, N4958, N7601);
or OR3 (N18078, N18043, N5718, N4623);
not NOT1 (N18079, N18068);
or OR4 (N18080, N18077, N15659, N3743, N6678);
xor XOR2 (N18081, N18075, N9048);
nand NAND4 (N18082, N18059, N12454, N3105, N14967);
nand NAND4 (N18083, N18079, N4751, N10284, N12987);
or OR2 (N18084, N18078, N6871);
nand NAND3 (N18085, N18071, N2260, N11466);
not NOT1 (N18086, N18076);
buf BUF1 (N18087, N18082);
buf BUF1 (N18088, N18067);
nor NOR3 (N18089, N18070, N11824, N14420);
or OR2 (N18090, N18080, N16676);
xor XOR2 (N18091, N18090, N16782);
and AND4 (N18092, N18083, N14292, N17164, N12256);
xor XOR2 (N18093, N18081, N16561);
nor NOR3 (N18094, N18085, N9752, N5382);
buf BUF1 (N18095, N18087);
or OR4 (N18096, N18095, N4226, N10558, N9858);
xor XOR2 (N18097, N18074, N3365);
or OR3 (N18098, N18091, N13765, N7453);
nand NAND4 (N18099, N18092, N378, N9869, N8395);
xor XOR2 (N18100, N18098, N15955);
nand NAND4 (N18101, N18089, N3807, N15302, N11160);
buf BUF1 (N18102, N18099);
or OR3 (N18103, N18101, N10446, N14660);
nor NOR4 (N18104, N18103, N7076, N7318, N4455);
or OR4 (N18105, N18093, N2147, N3505, N9571);
and AND2 (N18106, N18094, N10858);
nor NOR2 (N18107, N18106, N933);
nand NAND4 (N18108, N18107, N12776, N16343, N16770);
xor XOR2 (N18109, N18088, N13921);
and AND3 (N18110, N18105, N8979, N14194);
nand NAND4 (N18111, N18108, N14382, N965, N7042);
nand NAND2 (N18112, N18100, N17961);
nand NAND2 (N18113, N18102, N7902);
nand NAND2 (N18114, N18109, N6424);
and AND2 (N18115, N18113, N10319);
nand NAND3 (N18116, N18084, N7349, N16573);
buf BUF1 (N18117, N18116);
buf BUF1 (N18118, N18104);
nor NOR2 (N18119, N18097, N3057);
or OR2 (N18120, N18117, N10075);
nor NOR4 (N18121, N18111, N9880, N3746, N3660);
nor NOR2 (N18122, N18096, N13945);
xor XOR2 (N18123, N18122, N2242);
buf BUF1 (N18124, N18114);
and AND2 (N18125, N18124, N5664);
xor XOR2 (N18126, N18121, N16991);
and AND2 (N18127, N18110, N11400);
or OR2 (N18128, N18126, N12363);
nor NOR4 (N18129, N18119, N7977, N8259, N14918);
nor NOR4 (N18130, N18086, N9214, N6819, N9233);
nand NAND2 (N18131, N18123, N14446);
not NOT1 (N18132, N18112);
nand NAND2 (N18133, N18129, N8084);
buf BUF1 (N18134, N18125);
not NOT1 (N18135, N18118);
nor NOR2 (N18136, N18115, N3086);
or OR2 (N18137, N18127, N10247);
nor NOR2 (N18138, N18134, N13309);
nand NAND4 (N18139, N18128, N17286, N14802, N2270);
nand NAND3 (N18140, N18139, N10139, N10768);
or OR3 (N18141, N18133, N12682, N8492);
nor NOR2 (N18142, N18132, N1200);
nor NOR2 (N18143, N18135, N9154);
and AND4 (N18144, N18138, N5255, N8242, N5518);
xor XOR2 (N18145, N18131, N3169);
buf BUF1 (N18146, N18143);
not NOT1 (N18147, N18120);
nor NOR3 (N18148, N18136, N8422, N661);
and AND2 (N18149, N18140, N10133);
buf BUF1 (N18150, N18137);
buf BUF1 (N18151, N18147);
not NOT1 (N18152, N18148);
buf BUF1 (N18153, N18150);
buf BUF1 (N18154, N18145);
nor NOR4 (N18155, N18153, N2104, N212, N4586);
xor XOR2 (N18156, N18141, N957);
nand NAND3 (N18157, N18155, N17239, N11365);
buf BUF1 (N18158, N18157);
nor NOR3 (N18159, N18158, N14779, N15942);
nor NOR2 (N18160, N18142, N10835);
xor XOR2 (N18161, N18154, N3419);
and AND4 (N18162, N18144, N15870, N2165, N6102);
or OR4 (N18163, N18146, N15695, N17676, N16064);
or OR4 (N18164, N18161, N9358, N11320, N5685);
or OR4 (N18165, N18156, N6598, N3463, N2684);
or OR3 (N18166, N18163, N12475, N3369);
not NOT1 (N18167, N18159);
xor XOR2 (N18168, N18165, N16364);
nor NOR4 (N18169, N18152, N4439, N17846, N944);
and AND3 (N18170, N18169, N6935, N17959);
or OR3 (N18171, N18166, N2431, N10522);
xor XOR2 (N18172, N18170, N4916);
or OR2 (N18173, N18171, N15454);
buf BUF1 (N18174, N18149);
xor XOR2 (N18175, N18164, N9741);
not NOT1 (N18176, N18172);
xor XOR2 (N18177, N18173, N12069);
nand NAND3 (N18178, N18176, N17721, N13550);
buf BUF1 (N18179, N18160);
buf BUF1 (N18180, N18177);
xor XOR2 (N18181, N18175, N8943);
or OR3 (N18182, N18179, N2383, N5536);
xor XOR2 (N18183, N18174, N6657);
or OR3 (N18184, N18130, N18153, N9709);
buf BUF1 (N18185, N18178);
xor XOR2 (N18186, N18183, N13508);
not NOT1 (N18187, N18151);
nor NOR3 (N18188, N18186, N15494, N8110);
xor XOR2 (N18189, N18180, N14512);
nand NAND4 (N18190, N18187, N7975, N5939, N15702);
xor XOR2 (N18191, N18167, N8110);
not NOT1 (N18192, N18188);
not NOT1 (N18193, N18191);
and AND3 (N18194, N18184, N9429, N3189);
xor XOR2 (N18195, N18168, N5956);
nor NOR2 (N18196, N18193, N9560);
nand NAND2 (N18197, N18192, N1561);
and AND2 (N18198, N18195, N17054);
and AND4 (N18199, N18181, N5682, N11418, N220);
buf BUF1 (N18200, N18189);
not NOT1 (N18201, N18185);
buf BUF1 (N18202, N18200);
or OR2 (N18203, N18162, N17713);
nand NAND3 (N18204, N18194, N2316, N2521);
not NOT1 (N18205, N18198);
or OR3 (N18206, N18190, N888, N16613);
xor XOR2 (N18207, N18204, N12204);
buf BUF1 (N18208, N18203);
not NOT1 (N18209, N18205);
xor XOR2 (N18210, N18209, N17620);
and AND3 (N18211, N18202, N1292, N8232);
or OR4 (N18212, N18208, N15680, N16226, N6398);
or OR4 (N18213, N18182, N5667, N6331, N17734);
buf BUF1 (N18214, N18207);
or OR4 (N18215, N18199, N12378, N10595, N12286);
and AND3 (N18216, N18210, N5008, N15714);
buf BUF1 (N18217, N18214);
and AND4 (N18218, N18213, N9871, N17929, N9281);
or OR4 (N18219, N18216, N4445, N12195, N14201);
buf BUF1 (N18220, N18212);
xor XOR2 (N18221, N18197, N14306);
nor NOR2 (N18222, N18219, N4671);
buf BUF1 (N18223, N18215);
and AND2 (N18224, N18201, N15401);
and AND3 (N18225, N18206, N3835, N3343);
xor XOR2 (N18226, N18217, N2548);
buf BUF1 (N18227, N18218);
and AND2 (N18228, N18227, N6931);
buf BUF1 (N18229, N18196);
nor NOR4 (N18230, N18226, N8764, N15532, N4169);
and AND3 (N18231, N18221, N6063, N15690);
or OR3 (N18232, N18222, N15353, N5959);
nand NAND3 (N18233, N18224, N9146, N4271);
nand NAND3 (N18234, N18223, N8623, N2725);
xor XOR2 (N18235, N18228, N15752);
nor NOR2 (N18236, N18231, N466);
buf BUF1 (N18237, N18235);
or OR2 (N18238, N18233, N4972);
nand NAND3 (N18239, N18236, N1834, N3705);
buf BUF1 (N18240, N18232);
xor XOR2 (N18241, N18240, N3322);
not NOT1 (N18242, N18229);
nor NOR4 (N18243, N18238, N8635, N9548, N17451);
and AND4 (N18244, N18220, N11771, N328, N8306);
and AND4 (N18245, N18239, N10066, N11432, N9989);
xor XOR2 (N18246, N18225, N7965);
or OR4 (N18247, N18242, N1949, N4292, N4711);
xor XOR2 (N18248, N18230, N15412);
nor NOR3 (N18249, N18247, N16859, N9482);
nand NAND4 (N18250, N18237, N14125, N12095, N17436);
nand NAND2 (N18251, N18250, N3504);
or OR2 (N18252, N18244, N4186);
xor XOR2 (N18253, N18241, N17376);
not NOT1 (N18254, N18248);
nand NAND3 (N18255, N18211, N12152, N8112);
buf BUF1 (N18256, N18253);
buf BUF1 (N18257, N18254);
xor XOR2 (N18258, N18257, N17996);
or OR4 (N18259, N18258, N8509, N3690, N2373);
xor XOR2 (N18260, N18246, N14011);
or OR4 (N18261, N18245, N9119, N15511, N7608);
or OR4 (N18262, N18260, N9707, N672, N6106);
nand NAND4 (N18263, N18252, N3752, N8979, N6100);
buf BUF1 (N18264, N18251);
buf BUF1 (N18265, N18264);
or OR2 (N18266, N18263, N6892);
buf BUF1 (N18267, N18265);
xor XOR2 (N18268, N18267, N13546);
nor NOR2 (N18269, N18268, N6052);
buf BUF1 (N18270, N18266);
nor NOR4 (N18271, N18262, N10112, N5913, N17878);
nor NOR2 (N18272, N18261, N4577);
or OR3 (N18273, N18243, N13308, N4154);
buf BUF1 (N18274, N18255);
nor NOR4 (N18275, N18269, N3991, N8216, N561);
nor NOR2 (N18276, N18274, N12764);
not NOT1 (N18277, N18271);
nand NAND4 (N18278, N18270, N4626, N2755, N10971);
or OR3 (N18279, N18256, N12177, N7841);
or OR2 (N18280, N18259, N17910);
xor XOR2 (N18281, N18279, N14880);
not NOT1 (N18282, N18275);
not NOT1 (N18283, N18281);
buf BUF1 (N18284, N18249);
xor XOR2 (N18285, N18273, N10330);
buf BUF1 (N18286, N18272);
or OR3 (N18287, N18278, N5846, N3929);
nor NOR2 (N18288, N18234, N3245);
not NOT1 (N18289, N18285);
nand NAND2 (N18290, N18277, N8973);
xor XOR2 (N18291, N18290, N17035);
xor XOR2 (N18292, N18284, N17902);
buf BUF1 (N18293, N18286);
not NOT1 (N18294, N18289);
and AND3 (N18295, N18294, N11674, N11290);
not NOT1 (N18296, N18295);
nand NAND2 (N18297, N18291, N13654);
or OR4 (N18298, N18276, N1621, N7359, N4413);
and AND4 (N18299, N18287, N10351, N10997, N4497);
nor NOR3 (N18300, N18298, N12676, N15908);
and AND2 (N18301, N18293, N15754);
and AND3 (N18302, N18280, N12677, N6724);
buf BUF1 (N18303, N18282);
not NOT1 (N18304, N18299);
or OR4 (N18305, N18292, N17554, N5164, N10014);
xor XOR2 (N18306, N18300, N17591);
buf BUF1 (N18307, N18283);
buf BUF1 (N18308, N18305);
buf BUF1 (N18309, N18303);
nor NOR3 (N18310, N18306, N3969, N15486);
buf BUF1 (N18311, N18308);
or OR2 (N18312, N18296, N2511);
buf BUF1 (N18313, N18297);
not NOT1 (N18314, N18304);
or OR2 (N18315, N18307, N6164);
nor NOR4 (N18316, N18310, N982, N12686, N17852);
nor NOR3 (N18317, N18311, N15715, N8190);
nor NOR3 (N18318, N18315, N9213, N10196);
not NOT1 (N18319, N18313);
and AND4 (N18320, N18301, N7645, N13987, N11956);
or OR3 (N18321, N18312, N6544, N1100);
or OR3 (N18322, N18314, N7781, N13976);
nor NOR4 (N18323, N18318, N8278, N12166, N6066);
xor XOR2 (N18324, N18317, N14831);
nand NAND2 (N18325, N18288, N490);
nand NAND2 (N18326, N18316, N7027);
nand NAND3 (N18327, N18321, N14675, N15672);
buf BUF1 (N18328, N18319);
not NOT1 (N18329, N18320);
or OR2 (N18330, N18326, N14820);
xor XOR2 (N18331, N18323, N13410);
not NOT1 (N18332, N18329);
and AND4 (N18333, N18302, N8767, N9488, N9831);
xor XOR2 (N18334, N18324, N3809);
xor XOR2 (N18335, N18334, N10414);
nor NOR2 (N18336, N18322, N15140);
nor NOR2 (N18337, N18327, N15250);
buf BUF1 (N18338, N18330);
nand NAND3 (N18339, N18336, N16276, N378);
xor XOR2 (N18340, N18335, N382);
buf BUF1 (N18341, N18309);
or OR2 (N18342, N18338, N16034);
and AND4 (N18343, N18325, N8544, N6442, N9504);
not NOT1 (N18344, N18332);
not NOT1 (N18345, N18341);
nand NAND2 (N18346, N18333, N11936);
xor XOR2 (N18347, N18343, N5115);
or OR4 (N18348, N18331, N4223, N1446, N13770);
nor NOR2 (N18349, N18340, N16268);
nand NAND2 (N18350, N18346, N3375);
xor XOR2 (N18351, N18347, N9128);
and AND2 (N18352, N18339, N8140);
nor NOR2 (N18353, N18345, N3934);
not NOT1 (N18354, N18337);
nor NOR3 (N18355, N18352, N15676, N5519);
and AND4 (N18356, N18350, N11378, N2512, N12190);
xor XOR2 (N18357, N18351, N11619);
buf BUF1 (N18358, N18355);
xor XOR2 (N18359, N18353, N9959);
or OR2 (N18360, N18357, N4122);
nor NOR4 (N18361, N18359, N5061, N6178, N13129);
nand NAND4 (N18362, N18328, N13446, N11641, N9808);
or OR3 (N18363, N18360, N7597, N5914);
nand NAND3 (N18364, N18342, N14729, N627);
not NOT1 (N18365, N18344);
xor XOR2 (N18366, N18364, N10074);
or OR3 (N18367, N18348, N16729, N15692);
nand NAND4 (N18368, N18365, N8030, N15149, N2509);
buf BUF1 (N18369, N18368);
nand NAND3 (N18370, N18362, N14612, N5665);
nand NAND2 (N18371, N18370, N3805);
buf BUF1 (N18372, N18356);
xor XOR2 (N18373, N18363, N616);
xor XOR2 (N18374, N18366, N14189);
or OR4 (N18375, N18367, N562, N13701, N5527);
not NOT1 (N18376, N18372);
nor NOR4 (N18377, N18376, N11523, N2065, N12409);
nand NAND2 (N18378, N18349, N10475);
xor XOR2 (N18379, N18375, N8538);
nor NOR4 (N18380, N18354, N3678, N15035, N11561);
buf BUF1 (N18381, N18361);
nor NOR3 (N18382, N18380, N18112, N10745);
or OR2 (N18383, N18371, N344);
nor NOR2 (N18384, N18377, N10340);
nor NOR3 (N18385, N18382, N12870, N8004);
not NOT1 (N18386, N18378);
and AND3 (N18387, N18373, N5716, N13790);
and AND4 (N18388, N18384, N649, N8566, N8613);
buf BUF1 (N18389, N18385);
or OR3 (N18390, N18381, N12963, N6499);
xor XOR2 (N18391, N18386, N12405);
buf BUF1 (N18392, N18391);
xor XOR2 (N18393, N18390, N14040);
nand NAND2 (N18394, N18393, N13207);
and AND2 (N18395, N18369, N13641);
or OR3 (N18396, N18395, N9171, N5062);
nor NOR2 (N18397, N18379, N8245);
xor XOR2 (N18398, N18383, N1205);
xor XOR2 (N18399, N18396, N1600);
not NOT1 (N18400, N18388);
and AND2 (N18401, N18392, N4113);
or OR2 (N18402, N18389, N135);
nor NOR3 (N18403, N18401, N11401, N13756);
xor XOR2 (N18404, N18398, N5178);
not NOT1 (N18405, N18403);
nand NAND2 (N18406, N18404, N13511);
not NOT1 (N18407, N18394);
not NOT1 (N18408, N18400);
not NOT1 (N18409, N18407);
nand NAND4 (N18410, N18409, N4991, N10877, N2381);
buf BUF1 (N18411, N18358);
buf BUF1 (N18412, N18374);
nor NOR4 (N18413, N18397, N15944, N1316, N8978);
and AND4 (N18414, N18410, N1449, N3838, N7612);
xor XOR2 (N18415, N18402, N12918);
nor NOR3 (N18416, N18405, N9271, N16357);
nand NAND2 (N18417, N18406, N1427);
buf BUF1 (N18418, N18413);
nor NOR4 (N18419, N18418, N3734, N3674, N591);
xor XOR2 (N18420, N18417, N9710);
buf BUF1 (N18421, N18415);
nor NOR2 (N18422, N18419, N11571);
buf BUF1 (N18423, N18416);
xor XOR2 (N18424, N18423, N6706);
nor NOR3 (N18425, N18399, N3129, N5997);
nand NAND2 (N18426, N18425, N7595);
nand NAND4 (N18427, N18426, N8485, N9018, N8641);
buf BUF1 (N18428, N18424);
nand NAND4 (N18429, N18412, N3961, N2771, N8083);
nor NOR2 (N18430, N18421, N4359);
or OR2 (N18431, N18420, N10118);
or OR3 (N18432, N18430, N7220, N5526);
xor XOR2 (N18433, N18422, N9811);
nand NAND3 (N18434, N18387, N14945, N9811);
buf BUF1 (N18435, N18428);
nand NAND2 (N18436, N18434, N7481);
not NOT1 (N18437, N18427);
xor XOR2 (N18438, N18432, N14217);
xor XOR2 (N18439, N18408, N16404);
nand NAND4 (N18440, N18411, N9506, N16262, N7985);
and AND4 (N18441, N18433, N9762, N3965, N18237);
buf BUF1 (N18442, N18438);
nand NAND4 (N18443, N18414, N17415, N806, N2200);
and AND3 (N18444, N18437, N5830, N9247);
nand NAND2 (N18445, N18439, N15992);
nor NOR4 (N18446, N18443, N4052, N4833, N8386);
xor XOR2 (N18447, N18441, N5222);
xor XOR2 (N18448, N18445, N17903);
not NOT1 (N18449, N18436);
nor NOR4 (N18450, N18448, N5803, N11505, N12061);
buf BUF1 (N18451, N18447);
buf BUF1 (N18452, N18450);
buf BUF1 (N18453, N18452);
and AND3 (N18454, N18446, N17227, N13504);
buf BUF1 (N18455, N18431);
buf BUF1 (N18456, N18444);
or OR3 (N18457, N18442, N8576, N9619);
and AND3 (N18458, N18455, N5105, N36);
nand NAND3 (N18459, N18449, N190, N14428);
xor XOR2 (N18460, N18458, N5357);
nand NAND3 (N18461, N18451, N3867, N18436);
nand NAND3 (N18462, N18429, N15717, N15963);
nor NOR3 (N18463, N18453, N16446, N4023);
not NOT1 (N18464, N18435);
nor NOR3 (N18465, N18456, N15641, N453);
and AND4 (N18466, N18462, N2758, N6443, N16155);
nor NOR2 (N18467, N18461, N4921);
nor NOR4 (N18468, N18457, N2988, N5759, N15488);
xor XOR2 (N18469, N18463, N4292);
buf BUF1 (N18470, N18459);
xor XOR2 (N18471, N18470, N11484);
xor XOR2 (N18472, N18468, N113);
xor XOR2 (N18473, N18460, N8837);
not NOT1 (N18474, N18464);
nand NAND4 (N18475, N18465, N5911, N809, N13047);
xor XOR2 (N18476, N18469, N16644);
and AND3 (N18477, N18472, N327, N16246);
nand NAND2 (N18478, N18477, N17424);
nand NAND4 (N18479, N18454, N11464, N862, N13714);
nand NAND3 (N18480, N18478, N6550, N11537);
buf BUF1 (N18481, N18466);
xor XOR2 (N18482, N18474, N56);
xor XOR2 (N18483, N18475, N15304);
nand NAND2 (N18484, N18473, N6890);
xor XOR2 (N18485, N18484, N17430);
buf BUF1 (N18486, N18467);
nor NOR4 (N18487, N18476, N13230, N687, N11553);
and AND3 (N18488, N18482, N10276, N3162);
buf BUF1 (N18489, N18471);
xor XOR2 (N18490, N18485, N16866);
nor NOR4 (N18491, N18487, N15435, N12123, N7125);
buf BUF1 (N18492, N18491);
and AND3 (N18493, N18486, N8446, N10616);
xor XOR2 (N18494, N18483, N16004);
nand NAND2 (N18495, N18488, N143);
nor NOR2 (N18496, N18481, N15288);
buf BUF1 (N18497, N18480);
or OR3 (N18498, N18489, N18262, N5119);
nand NAND2 (N18499, N18497, N16848);
buf BUF1 (N18500, N18498);
nor NOR2 (N18501, N18493, N13941);
not NOT1 (N18502, N18495);
or OR4 (N18503, N18492, N13434, N2034, N12002);
and AND4 (N18504, N18490, N13236, N6056, N7487);
nor NOR3 (N18505, N18504, N3649, N17748);
or OR4 (N18506, N18496, N6380, N16976, N9089);
not NOT1 (N18507, N18502);
not NOT1 (N18508, N18503);
nand NAND4 (N18509, N18499, N4298, N357, N10134);
not NOT1 (N18510, N18505);
buf BUF1 (N18511, N18494);
or OR4 (N18512, N18506, N16622, N3626, N17178);
nor NOR4 (N18513, N18512, N4546, N963, N14977);
nor NOR3 (N18514, N18501, N14271, N273);
xor XOR2 (N18515, N18514, N14375);
xor XOR2 (N18516, N18507, N6846);
buf BUF1 (N18517, N18500);
buf BUF1 (N18518, N18509);
nor NOR4 (N18519, N18510, N2748, N1675, N5600);
and AND3 (N18520, N18511, N9202, N5393);
nor NOR2 (N18521, N18516, N307);
and AND2 (N18522, N18515, N17889);
nor NOR4 (N18523, N18513, N1479, N17209, N8305);
buf BUF1 (N18524, N18519);
or OR4 (N18525, N18524, N11576, N674, N618);
not NOT1 (N18526, N18523);
not NOT1 (N18527, N18508);
xor XOR2 (N18528, N18520, N12909);
xor XOR2 (N18529, N18528, N6477);
and AND3 (N18530, N18525, N8680, N6996);
xor XOR2 (N18531, N18529, N17977);
and AND3 (N18532, N18531, N31, N15440);
and AND4 (N18533, N18517, N6850, N3992, N3320);
xor XOR2 (N18534, N18526, N16426);
not NOT1 (N18535, N18534);
nor NOR3 (N18536, N18532, N1829, N11847);
or OR2 (N18537, N18518, N12400);
and AND2 (N18538, N18533, N9818);
not NOT1 (N18539, N18527);
nor NOR3 (N18540, N18537, N13105, N15733);
nor NOR2 (N18541, N18522, N4885);
nor NOR2 (N18542, N18538, N6545);
buf BUF1 (N18543, N18542);
nor NOR2 (N18544, N18521, N11805);
nand NAND2 (N18545, N18539, N16843);
not NOT1 (N18546, N18544);
not NOT1 (N18547, N18530);
and AND3 (N18548, N18540, N452, N303);
xor XOR2 (N18549, N18543, N4652);
and AND3 (N18550, N18546, N17823, N4701);
buf BUF1 (N18551, N18549);
and AND3 (N18552, N18545, N5346, N17578);
and AND4 (N18553, N18550, N6463, N8912, N2130);
nand NAND3 (N18554, N18553, N7469, N3177);
not NOT1 (N18555, N18440);
xor XOR2 (N18556, N18555, N8191);
not NOT1 (N18557, N18535);
and AND4 (N18558, N18547, N7049, N3983, N17263);
not NOT1 (N18559, N18557);
nand NAND4 (N18560, N18554, N2098, N3726, N15155);
not NOT1 (N18561, N18558);
and AND2 (N18562, N18479, N16603);
not NOT1 (N18563, N18536);
nand NAND2 (N18564, N18562, N17164);
buf BUF1 (N18565, N18560);
and AND3 (N18566, N18551, N11784, N3813);
and AND4 (N18567, N18541, N1293, N2930, N17058);
nand NAND2 (N18568, N18567, N8152);
xor XOR2 (N18569, N18563, N8224);
buf BUF1 (N18570, N18552);
nand NAND4 (N18571, N18556, N3853, N14385, N12823);
xor XOR2 (N18572, N18569, N11105);
buf BUF1 (N18573, N18572);
buf BUF1 (N18574, N18564);
nor NOR2 (N18575, N18574, N12796);
nor NOR4 (N18576, N18571, N13979, N14819, N15494);
not NOT1 (N18577, N18575);
and AND2 (N18578, N18573, N16685);
xor XOR2 (N18579, N18559, N9693);
or OR2 (N18580, N18565, N4236);
nand NAND2 (N18581, N18579, N9665);
and AND4 (N18582, N18548, N13640, N14153, N12941);
buf BUF1 (N18583, N18561);
or OR3 (N18584, N18583, N11813, N18206);
xor XOR2 (N18585, N18584, N15143);
not NOT1 (N18586, N18576);
xor XOR2 (N18587, N18585, N7074);
not NOT1 (N18588, N18587);
nor NOR2 (N18589, N18568, N15314);
and AND4 (N18590, N18566, N15249, N11704, N2812);
xor XOR2 (N18591, N18581, N10256);
not NOT1 (N18592, N18582);
xor XOR2 (N18593, N18586, N11614);
or OR2 (N18594, N18578, N9818);
xor XOR2 (N18595, N18592, N7413);
not NOT1 (N18596, N18580);
nand NAND4 (N18597, N18570, N9107, N397, N16115);
nand NAND2 (N18598, N18590, N16745);
xor XOR2 (N18599, N18588, N4889);
not NOT1 (N18600, N18577);
buf BUF1 (N18601, N18589);
nand NAND3 (N18602, N18598, N17776, N15012);
nand NAND4 (N18603, N18593, N1575, N6513, N8820);
xor XOR2 (N18604, N18597, N6893);
and AND4 (N18605, N18599, N15997, N13178, N2196);
not NOT1 (N18606, N18595);
or OR4 (N18607, N18602, N8672, N4710, N6053);
not NOT1 (N18608, N18603);
buf BUF1 (N18609, N18596);
not NOT1 (N18610, N18601);
nor NOR2 (N18611, N18607, N10891);
nand NAND3 (N18612, N18600, N9843, N16559);
nand NAND3 (N18613, N18606, N12803, N12632);
not NOT1 (N18614, N18613);
nand NAND2 (N18615, N18610, N23);
not NOT1 (N18616, N18591);
and AND4 (N18617, N18612, N5200, N14361, N2924);
not NOT1 (N18618, N18617);
and AND3 (N18619, N18609, N15628, N7380);
or OR4 (N18620, N18614, N8816, N10592, N7869);
buf BUF1 (N18621, N18620);
nand NAND4 (N18622, N18618, N18509, N6997, N11055);
not NOT1 (N18623, N18616);
nand NAND2 (N18624, N18605, N3736);
nor NOR3 (N18625, N18594, N59, N12267);
and AND4 (N18626, N18615, N13556, N17334, N14867);
buf BUF1 (N18627, N18608);
nor NOR2 (N18628, N18611, N16455);
and AND2 (N18629, N18619, N3287);
not NOT1 (N18630, N18621);
nand NAND4 (N18631, N18623, N4487, N15892, N17201);
xor XOR2 (N18632, N18631, N14776);
or OR3 (N18633, N18627, N8321, N14403);
xor XOR2 (N18634, N18633, N14932);
and AND2 (N18635, N18604, N6161);
buf BUF1 (N18636, N18632);
nor NOR4 (N18637, N18636, N16079, N426, N10046);
nand NAND2 (N18638, N18622, N6444);
nand NAND2 (N18639, N18628, N2836);
and AND4 (N18640, N18638, N12336, N18263, N4601);
nand NAND3 (N18641, N18639, N8517, N11516);
or OR4 (N18642, N18625, N3944, N14768, N10623);
not NOT1 (N18643, N18637);
and AND4 (N18644, N18642, N17271, N6704, N5076);
or OR2 (N18645, N18635, N17094);
not NOT1 (N18646, N18626);
buf BUF1 (N18647, N18624);
not NOT1 (N18648, N18641);
or OR4 (N18649, N18630, N7403, N16834, N10596);
nand NAND3 (N18650, N18649, N6398, N3961);
xor XOR2 (N18651, N18629, N11178);
not NOT1 (N18652, N18647);
not NOT1 (N18653, N18640);
and AND3 (N18654, N18646, N12694, N17837);
buf BUF1 (N18655, N18652);
not NOT1 (N18656, N18655);
xor XOR2 (N18657, N18651, N5199);
not NOT1 (N18658, N18648);
xor XOR2 (N18659, N18657, N3923);
nand NAND2 (N18660, N18643, N10784);
buf BUF1 (N18661, N18658);
nand NAND2 (N18662, N18659, N1048);
nor NOR4 (N18663, N18661, N13828, N13489, N3759);
nand NAND4 (N18664, N18654, N7160, N16500, N17682);
buf BUF1 (N18665, N18656);
buf BUF1 (N18666, N18663);
nor NOR2 (N18667, N18662, N4774);
or OR3 (N18668, N18644, N14404, N9620);
or OR3 (N18669, N18653, N8920, N8298);
not NOT1 (N18670, N18668);
xor XOR2 (N18671, N18645, N7479);
and AND3 (N18672, N18671, N18557, N4440);
not NOT1 (N18673, N18634);
or OR4 (N18674, N18673, N1487, N9045, N10585);
and AND4 (N18675, N18669, N6788, N11813, N18199);
xor XOR2 (N18676, N18667, N2723);
buf BUF1 (N18677, N18666);
buf BUF1 (N18678, N18676);
nand NAND3 (N18679, N18664, N9606, N871);
nor NOR4 (N18680, N18660, N5628, N18280, N15238);
and AND2 (N18681, N18680, N15075);
xor XOR2 (N18682, N18650, N9496);
xor XOR2 (N18683, N18665, N9415);
nor NOR2 (N18684, N18672, N9443);
and AND3 (N18685, N18670, N16346, N515);
nor NOR4 (N18686, N18685, N11428, N14379, N14842);
buf BUF1 (N18687, N18678);
not NOT1 (N18688, N18687);
nor NOR2 (N18689, N18684, N16498);
and AND3 (N18690, N18686, N14043, N3047);
and AND2 (N18691, N18675, N3344);
and AND2 (N18692, N18690, N13107);
and AND3 (N18693, N18688, N13981, N269);
and AND4 (N18694, N18693, N13188, N3341, N8086);
and AND4 (N18695, N18692, N12347, N6430, N13339);
nand NAND3 (N18696, N18681, N11870, N13195);
nand NAND2 (N18697, N18696, N9281);
nand NAND2 (N18698, N18683, N7853);
buf BUF1 (N18699, N18677);
or OR3 (N18700, N18682, N7482, N377);
and AND3 (N18701, N18700, N9193, N2095);
and AND4 (N18702, N18674, N18435, N16910, N13415);
and AND2 (N18703, N18697, N6436);
or OR3 (N18704, N18699, N3000, N14615);
nand NAND4 (N18705, N18691, N6110, N4067, N6347);
not NOT1 (N18706, N18703);
buf BUF1 (N18707, N18694);
or OR4 (N18708, N18707, N11298, N4033, N16455);
not NOT1 (N18709, N18706);
buf BUF1 (N18710, N18702);
nor NOR4 (N18711, N18704, N14471, N18189, N864);
buf BUF1 (N18712, N18708);
not NOT1 (N18713, N18701);
buf BUF1 (N18714, N18712);
not NOT1 (N18715, N18705);
and AND4 (N18716, N18709, N16126, N15568, N6523);
and AND2 (N18717, N18695, N207);
nor NOR2 (N18718, N18698, N17726);
nor NOR2 (N18719, N18716, N6210);
not NOT1 (N18720, N18710);
nand NAND3 (N18721, N18720, N5172, N14213);
or OR3 (N18722, N18719, N7782, N4458);
nand NAND4 (N18723, N18715, N18005, N11157, N2846);
buf BUF1 (N18724, N18722);
or OR4 (N18725, N18713, N7111, N4137, N2942);
or OR4 (N18726, N18718, N6530, N1725, N11243);
nor NOR2 (N18727, N18714, N11060);
nand NAND4 (N18728, N18721, N8985, N17683, N5113);
nor NOR4 (N18729, N18726, N15600, N13820, N18462);
xor XOR2 (N18730, N18727, N16067);
buf BUF1 (N18731, N18730);
nand NAND4 (N18732, N18689, N9995, N18062, N1216);
nor NOR4 (N18733, N18717, N8087, N7958, N15187);
or OR3 (N18734, N18679, N3507, N2629);
buf BUF1 (N18735, N18729);
and AND3 (N18736, N18711, N6992, N16581);
nor NOR4 (N18737, N18735, N11890, N8708, N6316);
buf BUF1 (N18738, N18723);
and AND3 (N18739, N18725, N9415, N468);
buf BUF1 (N18740, N18734);
xor XOR2 (N18741, N18732, N18008);
xor XOR2 (N18742, N18724, N1513);
or OR3 (N18743, N18739, N181, N7659);
buf BUF1 (N18744, N18728);
buf BUF1 (N18745, N18743);
or OR2 (N18746, N18745, N1404);
nor NOR3 (N18747, N18733, N11370, N18031);
or OR2 (N18748, N18738, N14025);
not NOT1 (N18749, N18747);
buf BUF1 (N18750, N18746);
or OR3 (N18751, N18748, N7857, N4639);
xor XOR2 (N18752, N18741, N7998);
and AND4 (N18753, N18737, N16013, N15938, N8968);
nor NOR3 (N18754, N18731, N6843, N14611);
nand NAND2 (N18755, N18742, N1800);
nand NAND2 (N18756, N18755, N5038);
not NOT1 (N18757, N18752);
xor XOR2 (N18758, N18754, N7086);
and AND2 (N18759, N18749, N18000);
xor XOR2 (N18760, N18756, N11609);
not NOT1 (N18761, N18750);
or OR2 (N18762, N18740, N10866);
not NOT1 (N18763, N18753);
or OR3 (N18764, N18763, N3754, N11206);
buf BUF1 (N18765, N18744);
nor NOR3 (N18766, N18751, N13198, N11774);
and AND2 (N18767, N18759, N15064);
nor NOR4 (N18768, N18766, N6525, N8066, N11205);
and AND4 (N18769, N18764, N6068, N6544, N3620);
nand NAND4 (N18770, N18768, N15282, N3962, N17092);
nor NOR4 (N18771, N18765, N1634, N6890, N16975);
or OR3 (N18772, N18767, N12224, N15822);
nand NAND4 (N18773, N18761, N12820, N9094, N14179);
nor NOR4 (N18774, N18758, N1836, N9787, N13280);
nor NOR3 (N18775, N18762, N7440, N12584);
nand NAND4 (N18776, N18774, N10709, N13152, N1054);
buf BUF1 (N18777, N18769);
xor XOR2 (N18778, N18776, N5270);
nand NAND2 (N18779, N18777, N11578);
not NOT1 (N18780, N18770);
nor NOR2 (N18781, N18772, N3266);
or OR2 (N18782, N18781, N14395);
and AND2 (N18783, N18778, N4080);
buf BUF1 (N18784, N18780);
buf BUF1 (N18785, N18779);
not NOT1 (N18786, N18785);
nor NOR4 (N18787, N18786, N13901, N4615, N9520);
nor NOR3 (N18788, N18784, N17658, N6117);
nand NAND2 (N18789, N18782, N6280);
and AND4 (N18790, N18787, N12517, N367, N2797);
xor XOR2 (N18791, N18757, N14284);
xor XOR2 (N18792, N18771, N18190);
or OR2 (N18793, N18773, N11900);
not NOT1 (N18794, N18783);
xor XOR2 (N18795, N18792, N14509);
nand NAND4 (N18796, N18795, N12533, N8606, N9411);
not NOT1 (N18797, N18788);
or OR4 (N18798, N18790, N13082, N4856, N2444);
or OR3 (N18799, N18796, N3079, N919);
xor XOR2 (N18800, N18775, N14195);
not NOT1 (N18801, N18760);
nor NOR4 (N18802, N18801, N6836, N18167, N15822);
not NOT1 (N18803, N18789);
not NOT1 (N18804, N18794);
or OR3 (N18805, N18803, N10791, N10343);
xor XOR2 (N18806, N18736, N15209);
nor NOR2 (N18807, N18804, N16853);
nand NAND2 (N18808, N18807, N9681);
or OR4 (N18809, N18797, N5899, N8348, N16170);
xor XOR2 (N18810, N18809, N12906);
and AND3 (N18811, N18810, N154, N5551);
not NOT1 (N18812, N18793);
or OR4 (N18813, N18806, N18142, N16513, N10543);
nor NOR4 (N18814, N18808, N15997, N6973, N2236);
or OR2 (N18815, N18813, N9738);
buf BUF1 (N18816, N18814);
nor NOR2 (N18817, N18815, N3618);
and AND3 (N18818, N18811, N3901, N3976);
buf BUF1 (N18819, N18800);
buf BUF1 (N18820, N18799);
and AND3 (N18821, N18805, N4992, N14977);
not NOT1 (N18822, N18821);
buf BUF1 (N18823, N18819);
not NOT1 (N18824, N18791);
not NOT1 (N18825, N18820);
nor NOR4 (N18826, N18822, N14370, N15009, N4705);
xor XOR2 (N18827, N18818, N2340);
xor XOR2 (N18828, N18817, N16686);
not NOT1 (N18829, N18827);
not NOT1 (N18830, N18812);
nor NOR4 (N18831, N18802, N12435, N16535, N10204);
buf BUF1 (N18832, N18831);
and AND3 (N18833, N18825, N5391, N6184);
buf BUF1 (N18834, N18816);
nor NOR2 (N18835, N18833, N3989);
or OR3 (N18836, N18824, N16083, N15594);
not NOT1 (N18837, N18828);
nand NAND4 (N18838, N18836, N14450, N15450, N6086);
and AND2 (N18839, N18832, N4059);
xor XOR2 (N18840, N18834, N15109);
xor XOR2 (N18841, N18839, N8926);
nand NAND4 (N18842, N18837, N10043, N8664, N6235);
xor XOR2 (N18843, N18830, N4609);
nor NOR2 (N18844, N18798, N8928);
nand NAND4 (N18845, N18829, N18521, N17891, N13402);
buf BUF1 (N18846, N18826);
or OR2 (N18847, N18835, N4212);
not NOT1 (N18848, N18843);
and AND3 (N18849, N18848, N14513, N12425);
nand NAND3 (N18850, N18849, N7464, N16534);
not NOT1 (N18851, N18838);
nor NOR4 (N18852, N18842, N15851, N16756, N17283);
xor XOR2 (N18853, N18845, N16600);
nand NAND3 (N18854, N18846, N13322, N14537);
nor NOR3 (N18855, N18823, N8231, N17352);
and AND3 (N18856, N18841, N10558, N10543);
nor NOR2 (N18857, N18854, N2123);
buf BUF1 (N18858, N18852);
xor XOR2 (N18859, N18853, N620);
xor XOR2 (N18860, N18858, N8984);
or OR2 (N18861, N18860, N15646);
nor NOR2 (N18862, N18859, N7135);
and AND3 (N18863, N18857, N4627, N5283);
nand NAND3 (N18864, N18863, N1463, N3844);
nor NOR3 (N18865, N18847, N16178, N1427);
or OR4 (N18866, N18851, N14181, N9948, N16856);
not NOT1 (N18867, N18865);
not NOT1 (N18868, N18861);
not NOT1 (N18869, N18868);
nor NOR3 (N18870, N18856, N1424, N5309);
buf BUF1 (N18871, N18864);
not NOT1 (N18872, N18866);
nand NAND3 (N18873, N18855, N2785, N16396);
nand NAND2 (N18874, N18873, N1662);
buf BUF1 (N18875, N18869);
not NOT1 (N18876, N18870);
nor NOR4 (N18877, N18872, N8734, N16468, N5581);
not NOT1 (N18878, N18850);
buf BUF1 (N18879, N18840);
nor NOR3 (N18880, N18874, N9993, N10383);
nand NAND4 (N18881, N18876, N9637, N8107, N8484);
and AND3 (N18882, N18878, N12104, N6798);
buf BUF1 (N18883, N18880);
not NOT1 (N18884, N18882);
buf BUF1 (N18885, N18867);
nand NAND3 (N18886, N18844, N2058, N9098);
buf BUF1 (N18887, N18884);
and AND3 (N18888, N18881, N16782, N992);
not NOT1 (N18889, N18871);
not NOT1 (N18890, N18889);
nor NOR2 (N18891, N18886, N10760);
nor NOR2 (N18892, N18862, N11655);
and AND3 (N18893, N18883, N9323, N18148);
buf BUF1 (N18894, N18891);
not NOT1 (N18895, N18875);
not NOT1 (N18896, N18877);
buf BUF1 (N18897, N18879);
or OR2 (N18898, N18893, N6920);
nor NOR3 (N18899, N18895, N8881, N11854);
nor NOR4 (N18900, N18887, N16359, N1758, N72);
nor NOR3 (N18901, N18888, N17615, N3355);
buf BUF1 (N18902, N18890);
nand NAND3 (N18903, N18900, N7767, N3019);
nor NOR3 (N18904, N18897, N1863, N11894);
nand NAND4 (N18905, N18902, N9864, N4636, N2004);
nand NAND3 (N18906, N18892, N10153, N5961);
and AND2 (N18907, N18896, N15719);
not NOT1 (N18908, N18901);
buf BUF1 (N18909, N18907);
nand NAND2 (N18910, N18898, N3859);
nor NOR2 (N18911, N18885, N17481);
not NOT1 (N18912, N18899);
nor NOR4 (N18913, N18904, N7047, N6059, N15253);
xor XOR2 (N18914, N18905, N9733);
not NOT1 (N18915, N18908);
and AND2 (N18916, N18911, N17982);
xor XOR2 (N18917, N18903, N11819);
xor XOR2 (N18918, N18913, N18310);
buf BUF1 (N18919, N18906);
nor NOR2 (N18920, N18915, N12264);
xor XOR2 (N18921, N18912, N2210);
buf BUF1 (N18922, N18916);
not NOT1 (N18923, N18919);
or OR4 (N18924, N18922, N7720, N4478, N17711);
xor XOR2 (N18925, N18917, N11430);
xor XOR2 (N18926, N18894, N16100);
not NOT1 (N18927, N18925);
buf BUF1 (N18928, N18914);
or OR4 (N18929, N18926, N1164, N5567, N9585);
or OR3 (N18930, N18920, N18254, N15325);
buf BUF1 (N18931, N18910);
xor XOR2 (N18932, N18927, N17407);
xor XOR2 (N18933, N18932, N6687);
or OR2 (N18934, N18921, N16082);
buf BUF1 (N18935, N18918);
and AND4 (N18936, N18928, N7958, N9928, N18282);
buf BUF1 (N18937, N18924);
buf BUF1 (N18938, N18937);
or OR2 (N18939, N18923, N5258);
not NOT1 (N18940, N18933);
not NOT1 (N18941, N18936);
not NOT1 (N18942, N18929);
buf BUF1 (N18943, N18934);
buf BUF1 (N18944, N18909);
and AND4 (N18945, N18940, N12985, N8070, N1886);
buf BUF1 (N18946, N18939);
and AND4 (N18947, N18931, N11583, N3605, N3160);
and AND4 (N18948, N18930, N5284, N2134, N17906);
and AND4 (N18949, N18944, N14588, N3261, N7662);
buf BUF1 (N18950, N18938);
not NOT1 (N18951, N18942);
xor XOR2 (N18952, N18945, N1637);
xor XOR2 (N18953, N18952, N9461);
xor XOR2 (N18954, N18950, N18891);
and AND4 (N18955, N18946, N15388, N11553, N7206);
buf BUF1 (N18956, N18948);
not NOT1 (N18957, N18941);
xor XOR2 (N18958, N18947, N17153);
and AND3 (N18959, N18949, N6659, N1098);
nand NAND4 (N18960, N18957, N7120, N7555, N4300);
not NOT1 (N18961, N18943);
or OR4 (N18962, N18954, N15041, N14905, N10879);
not NOT1 (N18963, N18951);
or OR4 (N18964, N18956, N16773, N11128, N4507);
not NOT1 (N18965, N18964);
xor XOR2 (N18966, N18963, N9827);
nand NAND3 (N18967, N18960, N15375, N25);
or OR3 (N18968, N18935, N10471, N16174);
not NOT1 (N18969, N18961);
xor XOR2 (N18970, N18965, N8896);
xor XOR2 (N18971, N18955, N18555);
nor NOR3 (N18972, N18953, N17742, N12533);
and AND3 (N18973, N18958, N15061, N13830);
nor NOR3 (N18974, N18969, N7229, N5052);
not NOT1 (N18975, N18959);
xor XOR2 (N18976, N18973, N11512);
not NOT1 (N18977, N18970);
nand NAND4 (N18978, N18971, N7729, N12921, N14681);
buf BUF1 (N18979, N18967);
or OR2 (N18980, N18976, N5971);
not NOT1 (N18981, N18974);
nand NAND2 (N18982, N18972, N5892);
xor XOR2 (N18983, N18981, N17037);
xor XOR2 (N18984, N18977, N3405);
not NOT1 (N18985, N18982);
nand NAND3 (N18986, N18985, N13476, N11872);
buf BUF1 (N18987, N18986);
and AND4 (N18988, N18978, N15977, N9943, N12252);
buf BUF1 (N18989, N18975);
not NOT1 (N18990, N18989);
and AND3 (N18991, N18979, N15618, N9272);
or OR2 (N18992, N18988, N2409);
nand NAND3 (N18993, N18968, N10073, N6727);
not NOT1 (N18994, N18966);
buf BUF1 (N18995, N18987);
and AND3 (N18996, N18984, N2264, N14050);
nor NOR2 (N18997, N18991, N13259);
buf BUF1 (N18998, N18992);
buf BUF1 (N18999, N18995);
nor NOR3 (N19000, N18980, N18750, N15016);
and AND4 (N19001, N18990, N6826, N18773, N6417);
or OR2 (N19002, N19000, N11273);
or OR2 (N19003, N19001, N7309);
nand NAND3 (N19004, N18993, N13438, N18364);
nor NOR4 (N19005, N18994, N3987, N6237, N6715);
xor XOR2 (N19006, N18962, N8832);
and AND3 (N19007, N19006, N9104, N1395);
xor XOR2 (N19008, N19004, N13689);
not NOT1 (N19009, N18999);
not NOT1 (N19010, N19009);
not NOT1 (N19011, N18997);
or OR3 (N19012, N19008, N3525, N15333);
nand NAND2 (N19013, N18998, N4460);
xor XOR2 (N19014, N19012, N5412);
nor NOR2 (N19015, N19005, N3013);
not NOT1 (N19016, N19013);
or OR2 (N19017, N19014, N13847);
xor XOR2 (N19018, N19011, N12493);
nand NAND3 (N19019, N19017, N13190, N9081);
or OR4 (N19020, N19003, N15106, N14531, N11514);
nor NOR3 (N19021, N19018, N5798, N7254);
buf BUF1 (N19022, N18996);
not NOT1 (N19023, N19015);
nor NOR3 (N19024, N18983, N16265, N6380);
xor XOR2 (N19025, N19007, N10715);
nor NOR2 (N19026, N19016, N3589);
and AND3 (N19027, N19025, N11688, N12353);
not NOT1 (N19028, N19002);
xor XOR2 (N19029, N19021, N11453);
not NOT1 (N19030, N19024);
and AND2 (N19031, N19019, N7879);
nor NOR4 (N19032, N19010, N8673, N15750, N8903);
or OR2 (N19033, N19032, N5003);
nor NOR4 (N19034, N19031, N10607, N98, N8097);
nor NOR4 (N19035, N19026, N16283, N11323, N12478);
xor XOR2 (N19036, N19023, N3188);
nor NOR3 (N19037, N19030, N697, N12553);
nand NAND2 (N19038, N19027, N18795);
and AND3 (N19039, N19035, N18366, N16256);
nor NOR2 (N19040, N19029, N554);
nor NOR2 (N19041, N19037, N14855);
xor XOR2 (N19042, N19022, N15793);
nor NOR3 (N19043, N19034, N3031, N9401);
nor NOR2 (N19044, N19033, N12773);
and AND3 (N19045, N19039, N11015, N14617);
or OR3 (N19046, N19020, N10719, N11458);
xor XOR2 (N19047, N19040, N17657);
xor XOR2 (N19048, N19047, N7138);
not NOT1 (N19049, N19044);
or OR4 (N19050, N19043, N16213, N17525, N3206);
and AND4 (N19051, N19049, N10547, N12944, N11822);
buf BUF1 (N19052, N19036);
nor NOR2 (N19053, N19028, N18072);
and AND4 (N19054, N19052, N3028, N3650, N725);
nor NOR4 (N19055, N19046, N1110, N2169, N3135);
buf BUF1 (N19056, N19045);
buf BUF1 (N19057, N19053);
nand NAND3 (N19058, N19055, N14737, N2888);
buf BUF1 (N19059, N19057);
and AND3 (N19060, N19050, N2265, N15538);
nand NAND2 (N19061, N19038, N5390);
and AND3 (N19062, N19042, N14992, N1117);
or OR2 (N19063, N19061, N8027);
and AND3 (N19064, N19051, N1742, N892);
xor XOR2 (N19065, N19041, N400);
or OR4 (N19066, N19060, N9471, N3975, N16868);
xor XOR2 (N19067, N19064, N14827);
nand NAND4 (N19068, N19056, N7473, N1644, N12419);
or OR2 (N19069, N19063, N3838);
or OR4 (N19070, N19048, N17267, N6077, N15204);
buf BUF1 (N19071, N19066);
nand NAND3 (N19072, N19068, N2362, N6661);
xor XOR2 (N19073, N19069, N17724);
and AND2 (N19074, N19072, N9488);
nand NAND2 (N19075, N19059, N7507);
or OR4 (N19076, N19065, N7471, N13980, N3444);
buf BUF1 (N19077, N19074);
xor XOR2 (N19078, N19054, N18963);
nor NOR4 (N19079, N19078, N5408, N17831, N14236);
nor NOR2 (N19080, N19058, N15726);
xor XOR2 (N19081, N19067, N7308);
buf BUF1 (N19082, N19080);
and AND2 (N19083, N19070, N15877);
and AND4 (N19084, N19073, N13738, N2645, N4445);
nand NAND4 (N19085, N19071, N5172, N17877, N13210);
nor NOR3 (N19086, N19081, N7194, N12845);
not NOT1 (N19087, N19075);
buf BUF1 (N19088, N19062);
buf BUF1 (N19089, N19077);
xor XOR2 (N19090, N19088, N2870);
xor XOR2 (N19091, N19087, N15271);
nand NAND2 (N19092, N19091, N6831);
buf BUF1 (N19093, N19079);
and AND2 (N19094, N19083, N15886);
not NOT1 (N19095, N19089);
not NOT1 (N19096, N19076);
nand NAND3 (N19097, N19086, N15289, N1446);
or OR4 (N19098, N19094, N3383, N17333, N13129);
and AND2 (N19099, N19085, N3455);
nand NAND3 (N19100, N19095, N19071, N1817);
or OR4 (N19101, N19100, N4669, N12515, N10875);
xor XOR2 (N19102, N19097, N4683);
nand NAND3 (N19103, N19098, N10381, N13805);
nand NAND4 (N19104, N19103, N11134, N2398, N18421);
nand NAND2 (N19105, N19102, N16834);
buf BUF1 (N19106, N19084);
xor XOR2 (N19107, N19090, N15103);
not NOT1 (N19108, N19107);
buf BUF1 (N19109, N19093);
or OR3 (N19110, N19106, N18777, N2182);
xor XOR2 (N19111, N19110, N12368);
buf BUF1 (N19112, N19101);
or OR4 (N19113, N19108, N16047, N8216, N13829);
or OR2 (N19114, N19112, N19090);
buf BUF1 (N19115, N19111);
and AND3 (N19116, N19104, N13470, N830);
or OR4 (N19117, N19115, N1566, N1177, N16270);
and AND4 (N19118, N19109, N3728, N5373, N2530);
nor NOR3 (N19119, N19092, N1179, N18939);
nor NOR2 (N19120, N19082, N3919);
xor XOR2 (N19121, N19105, N4109);
nor NOR4 (N19122, N19099, N3971, N1956, N4022);
nand NAND3 (N19123, N19119, N4528, N7947);
or OR4 (N19124, N19096, N16281, N14474, N15709);
buf BUF1 (N19125, N19114);
xor XOR2 (N19126, N19123, N2508);
buf BUF1 (N19127, N19126);
xor XOR2 (N19128, N19122, N4425);
or OR2 (N19129, N19117, N2758);
not NOT1 (N19130, N19118);
not NOT1 (N19131, N19116);
nor NOR4 (N19132, N19131, N2277, N2963, N4703);
xor XOR2 (N19133, N19132, N7435);
buf BUF1 (N19134, N19129);
buf BUF1 (N19135, N19113);
buf BUF1 (N19136, N19130);
or OR2 (N19137, N19128, N13741);
not NOT1 (N19138, N19127);
nor NOR4 (N19139, N19120, N16478, N5904, N6136);
buf BUF1 (N19140, N19121);
and AND2 (N19141, N19138, N19134);
not NOT1 (N19142, N13993);
buf BUF1 (N19143, N19139);
buf BUF1 (N19144, N19124);
or OR3 (N19145, N19144, N4536, N13601);
nor NOR3 (N19146, N19137, N10342, N6650);
xor XOR2 (N19147, N19142, N12440);
and AND2 (N19148, N19125, N13713);
buf BUF1 (N19149, N19141);
nor NOR4 (N19150, N19143, N10235, N11873, N2632);
buf BUF1 (N19151, N19140);
or OR4 (N19152, N19149, N8498, N5128, N6544);
not NOT1 (N19153, N19150);
buf BUF1 (N19154, N19153);
nand NAND4 (N19155, N19136, N15636, N11976, N2826);
xor XOR2 (N19156, N19145, N934);
and AND3 (N19157, N19148, N14162, N6497);
and AND2 (N19158, N19147, N13073);
or OR4 (N19159, N19151, N4507, N1200, N14871);
nor NOR4 (N19160, N19152, N18706, N2337, N12736);
nor NOR2 (N19161, N19133, N11657);
not NOT1 (N19162, N19155);
and AND4 (N19163, N19157, N6644, N343, N19066);
or OR3 (N19164, N19146, N18343, N1696);
buf BUF1 (N19165, N19160);
xor XOR2 (N19166, N19135, N10196);
buf BUF1 (N19167, N19162);
buf BUF1 (N19168, N19165);
and AND2 (N19169, N19168, N18352);
nand NAND2 (N19170, N19156, N3102);
buf BUF1 (N19171, N19163);
buf BUF1 (N19172, N19158);
nand NAND2 (N19173, N19166, N6178);
nor NOR4 (N19174, N19159, N8003, N18843, N13888);
not NOT1 (N19175, N19161);
buf BUF1 (N19176, N19174);
nor NOR3 (N19177, N19173, N7992, N10858);
nand NAND3 (N19178, N19175, N18547, N13825);
and AND3 (N19179, N19167, N3167, N4771);
nor NOR4 (N19180, N19164, N16004, N14502, N11277);
nand NAND3 (N19181, N19171, N1961, N17987);
or OR4 (N19182, N19178, N11592, N4931, N1715);
xor XOR2 (N19183, N19169, N16136);
and AND3 (N19184, N19172, N10218, N18474);
buf BUF1 (N19185, N19177);
buf BUF1 (N19186, N19183);
xor XOR2 (N19187, N19185, N17673);
nor NOR4 (N19188, N19187, N3821, N16650, N12783);
buf BUF1 (N19189, N19188);
buf BUF1 (N19190, N19179);
buf BUF1 (N19191, N19186);
buf BUF1 (N19192, N19181);
or OR2 (N19193, N19180, N18813);
and AND2 (N19194, N19193, N8727);
or OR2 (N19195, N19170, N17823);
not NOT1 (N19196, N19189);
buf BUF1 (N19197, N19190);
nand NAND4 (N19198, N19192, N11377, N11619, N17138);
xor XOR2 (N19199, N19154, N13966);
xor XOR2 (N19200, N19197, N3433);
not NOT1 (N19201, N19194);
nor NOR4 (N19202, N19198, N14252, N13858, N8124);
nor NOR2 (N19203, N19201, N14579);
and AND3 (N19204, N19176, N8449, N18434);
not NOT1 (N19205, N19184);
buf BUF1 (N19206, N19199);
xor XOR2 (N19207, N19205, N12050);
xor XOR2 (N19208, N19191, N291);
nor NOR4 (N19209, N19207, N2035, N4873, N8193);
buf BUF1 (N19210, N19195);
xor XOR2 (N19211, N19200, N2762);
nor NOR3 (N19212, N19203, N4012, N7699);
buf BUF1 (N19213, N19196);
or OR4 (N19214, N19211, N6953, N14517, N8130);
or OR2 (N19215, N19208, N4345);
and AND3 (N19216, N19213, N7690, N8857);
not NOT1 (N19217, N19202);
xor XOR2 (N19218, N19209, N18430);
not NOT1 (N19219, N19218);
xor XOR2 (N19220, N19206, N8938);
nor NOR4 (N19221, N19204, N534, N18879, N12729);
buf BUF1 (N19222, N19221);
and AND4 (N19223, N19215, N12974, N12933, N3362);
or OR4 (N19224, N19223, N2726, N10960, N37);
or OR4 (N19225, N19214, N10342, N6713, N1106);
buf BUF1 (N19226, N19219);
xor XOR2 (N19227, N19224, N14051);
xor XOR2 (N19228, N19217, N8220);
or OR3 (N19229, N19226, N12832, N10041);
xor XOR2 (N19230, N19225, N11079);
nor NOR3 (N19231, N19220, N17045, N17773);
or OR3 (N19232, N19212, N8449, N1050);
or OR4 (N19233, N19222, N3885, N3620, N8838);
nand NAND2 (N19234, N19232, N3919);
and AND3 (N19235, N19229, N14165, N273);
or OR4 (N19236, N19235, N19152, N11115, N12927);
or OR3 (N19237, N19182, N9143, N11885);
nor NOR3 (N19238, N19237, N14342, N3436);
or OR4 (N19239, N19227, N9739, N13055, N4444);
and AND2 (N19240, N19238, N3930);
buf BUF1 (N19241, N19231);
nor NOR2 (N19242, N19233, N14793);
not NOT1 (N19243, N19239);
not NOT1 (N19244, N19210);
nand NAND3 (N19245, N19230, N9482, N15785);
buf BUF1 (N19246, N19244);
xor XOR2 (N19247, N19242, N18302);
not NOT1 (N19248, N19240);
nand NAND2 (N19249, N19248, N5905);
not NOT1 (N19250, N19228);
or OR3 (N19251, N19216, N17216, N13943);
xor XOR2 (N19252, N19236, N9978);
nor NOR3 (N19253, N19250, N17663, N11284);
or OR3 (N19254, N19246, N2269, N155);
buf BUF1 (N19255, N19243);
buf BUF1 (N19256, N19241);
nand NAND3 (N19257, N19252, N13684, N5126);
buf BUF1 (N19258, N19255);
nor NOR3 (N19259, N19258, N6606, N15819);
not NOT1 (N19260, N19247);
xor XOR2 (N19261, N19259, N7052);
nand NAND4 (N19262, N19261, N14526, N15372, N6850);
not NOT1 (N19263, N19256);
nand NAND3 (N19264, N19260, N4257, N11425);
nand NAND2 (N19265, N19254, N16726);
nand NAND3 (N19266, N19262, N15104, N1454);
nor NOR3 (N19267, N19264, N11447, N16);
xor XOR2 (N19268, N19266, N12805);
not NOT1 (N19269, N19251);
or OR3 (N19270, N19263, N1369, N15485);
xor XOR2 (N19271, N19253, N1068);
nor NOR4 (N19272, N19267, N308, N5236, N18451);
nor NOR2 (N19273, N19268, N12477);
nor NOR3 (N19274, N19272, N13709, N18739);
nor NOR2 (N19275, N19234, N8412);
or OR2 (N19276, N19270, N7193);
nor NOR3 (N19277, N19257, N8538, N12914);
buf BUF1 (N19278, N19269);
or OR2 (N19279, N19249, N574);
nand NAND2 (N19280, N19245, N4538);
not NOT1 (N19281, N19265);
and AND4 (N19282, N19274, N10744, N17639, N5147);
buf BUF1 (N19283, N19279);
not NOT1 (N19284, N19281);
nand NAND2 (N19285, N19278, N1277);
not NOT1 (N19286, N19273);
not NOT1 (N19287, N19275);
or OR4 (N19288, N19284, N1965, N19038, N2032);
buf BUF1 (N19289, N19277);
xor XOR2 (N19290, N19280, N8831);
not NOT1 (N19291, N19288);
or OR2 (N19292, N19276, N6967);
and AND2 (N19293, N19283, N6851);
or OR3 (N19294, N19290, N2209, N8714);
buf BUF1 (N19295, N19282);
and AND2 (N19296, N19285, N11823);
or OR2 (N19297, N19289, N11029);
and AND3 (N19298, N19291, N11607, N10950);
or OR4 (N19299, N19294, N15209, N1788, N365);
not NOT1 (N19300, N19271);
buf BUF1 (N19301, N19295);
nor NOR4 (N19302, N19292, N6284, N14009, N9832);
not NOT1 (N19303, N19297);
not NOT1 (N19304, N19298);
and AND4 (N19305, N19301, N3402, N1913, N17105);
buf BUF1 (N19306, N19303);
nor NOR2 (N19307, N19305, N3354);
xor XOR2 (N19308, N19299, N9394);
not NOT1 (N19309, N19300);
nand NAND2 (N19310, N19308, N9114);
xor XOR2 (N19311, N19286, N15448);
or OR4 (N19312, N19304, N6725, N4251, N9286);
or OR2 (N19313, N19296, N18684);
nand NAND2 (N19314, N19312, N1141);
not NOT1 (N19315, N19306);
or OR3 (N19316, N19315, N6493, N2325);
buf BUF1 (N19317, N19309);
xor XOR2 (N19318, N19302, N1166);
nand NAND4 (N19319, N19318, N8069, N18117, N1904);
nand NAND4 (N19320, N19313, N6402, N6448, N1477);
and AND4 (N19321, N19310, N10104, N11825, N9756);
and AND4 (N19322, N19321, N1694, N18416, N9125);
xor XOR2 (N19323, N19293, N8461);
not NOT1 (N19324, N19322);
not NOT1 (N19325, N19311);
nand NAND3 (N19326, N19320, N6928, N2652);
nand NAND2 (N19327, N19287, N5473);
nor NOR4 (N19328, N19319, N1666, N5705, N9379);
and AND4 (N19329, N19323, N15396, N5963, N11361);
nor NOR4 (N19330, N19326, N134, N6240, N15266);
buf BUF1 (N19331, N19307);
nand NAND3 (N19332, N19328, N12335, N17172);
xor XOR2 (N19333, N19329, N18111);
nand NAND3 (N19334, N19332, N4961, N15752);
and AND2 (N19335, N19327, N13296);
nor NOR4 (N19336, N19314, N13711, N9030, N1659);
xor XOR2 (N19337, N19316, N13523);
not NOT1 (N19338, N19334);
buf BUF1 (N19339, N19324);
and AND3 (N19340, N19330, N4943, N5155);
not NOT1 (N19341, N19338);
xor XOR2 (N19342, N19325, N4134);
or OR4 (N19343, N19339, N5344, N14035, N18955);
buf BUF1 (N19344, N19337);
nor NOR4 (N19345, N19341, N15998, N12341, N9314);
nor NOR2 (N19346, N19335, N8941);
not NOT1 (N19347, N19317);
nor NOR2 (N19348, N19342, N10693);
xor XOR2 (N19349, N19344, N3613);
or OR4 (N19350, N19348, N14422, N13925, N10232);
nand NAND2 (N19351, N19350, N12213);
buf BUF1 (N19352, N19331);
nor NOR4 (N19353, N19333, N16016, N17368, N13722);
nor NOR3 (N19354, N19351, N1261, N8924);
and AND4 (N19355, N19347, N18903, N1949, N218);
nand NAND2 (N19356, N19345, N6838);
buf BUF1 (N19357, N19352);
nor NOR4 (N19358, N19354, N5076, N7817, N11294);
buf BUF1 (N19359, N19353);
and AND4 (N19360, N19349, N2884, N13194, N1976);
and AND3 (N19361, N19360, N9268, N13557);
or OR2 (N19362, N19340, N5806);
and AND4 (N19363, N19336, N18257, N4678, N6605);
xor XOR2 (N19364, N19356, N18737);
and AND4 (N19365, N19363, N1749, N7562, N10591);
xor XOR2 (N19366, N19359, N813);
and AND3 (N19367, N19355, N3559, N1630);
nor NOR3 (N19368, N19366, N8178, N7921);
xor XOR2 (N19369, N19362, N11742);
buf BUF1 (N19370, N19365);
and AND2 (N19371, N19364, N4752);
nor NOR4 (N19372, N19343, N15681, N15443, N7168);
buf BUF1 (N19373, N19358);
xor XOR2 (N19374, N19373, N3777);
and AND4 (N19375, N19357, N18642, N13850, N16241);
or OR3 (N19376, N19367, N3288, N7120);
nand NAND2 (N19377, N19346, N15828);
buf BUF1 (N19378, N19369);
buf BUF1 (N19379, N19368);
not NOT1 (N19380, N19378);
nor NOR4 (N19381, N19376, N3394, N14376, N2755);
nand NAND3 (N19382, N19371, N6742, N18915);
buf BUF1 (N19383, N19382);
or OR2 (N19384, N19374, N7787);
buf BUF1 (N19385, N19361);
xor XOR2 (N19386, N19372, N15024);
not NOT1 (N19387, N19383);
and AND2 (N19388, N19380, N2405);
nor NOR2 (N19389, N19385, N2030);
buf BUF1 (N19390, N19388);
or OR2 (N19391, N19381, N3347);
xor XOR2 (N19392, N19390, N11978);
or OR2 (N19393, N19392, N8375);
buf BUF1 (N19394, N19387);
or OR4 (N19395, N19384, N1226, N4851, N7208);
buf BUF1 (N19396, N19377);
buf BUF1 (N19397, N19394);
and AND3 (N19398, N19379, N5448, N2798);
or OR4 (N19399, N19397, N16672, N10876, N5030);
buf BUF1 (N19400, N19399);
nand NAND4 (N19401, N19370, N1184, N7997, N18933);
and AND4 (N19402, N19386, N16066, N9157, N13431);
and AND3 (N19403, N19396, N5153, N2030);
nand NAND4 (N19404, N19402, N8525, N18512, N8028);
nand NAND2 (N19405, N19391, N9910);
buf BUF1 (N19406, N19389);
not NOT1 (N19407, N19404);
nand NAND2 (N19408, N19400, N11257);
xor XOR2 (N19409, N19401, N18383);
nand NAND2 (N19410, N19398, N16542);
xor XOR2 (N19411, N19407, N18635);
and AND4 (N19412, N19393, N14509, N16796, N15714);
nor NOR3 (N19413, N19405, N16929, N2734);
or OR2 (N19414, N19410, N7495);
or OR3 (N19415, N19412, N4713, N3528);
or OR2 (N19416, N19409, N3439);
nand NAND3 (N19417, N19375, N5334, N7966);
and AND4 (N19418, N19411, N3355, N4203, N5005);
and AND2 (N19419, N19413, N271);
nor NOR3 (N19420, N19395, N5363, N7265);
buf BUF1 (N19421, N19406);
nor NOR2 (N19422, N19421, N6734);
or OR4 (N19423, N19416, N2833, N3013, N10098);
or OR4 (N19424, N19415, N5630, N3402, N7412);
xor XOR2 (N19425, N19408, N2653);
buf BUF1 (N19426, N19424);
nand NAND3 (N19427, N19418, N9199, N9867);
xor XOR2 (N19428, N19414, N142);
not NOT1 (N19429, N19417);
buf BUF1 (N19430, N19419);
nand NAND2 (N19431, N19425, N16069);
xor XOR2 (N19432, N19422, N10525);
buf BUF1 (N19433, N19431);
buf BUF1 (N19434, N19433);
xor XOR2 (N19435, N19427, N8648);
buf BUF1 (N19436, N19420);
or OR3 (N19437, N19423, N681, N12084);
not NOT1 (N19438, N19436);
and AND3 (N19439, N19438, N4329, N17051);
xor XOR2 (N19440, N19429, N4986);
or OR4 (N19441, N19430, N7463, N13272, N14751);
not NOT1 (N19442, N19434);
xor XOR2 (N19443, N19437, N13930);
nand NAND2 (N19444, N19443, N16470);
or OR3 (N19445, N19442, N7350, N2245);
nand NAND2 (N19446, N19439, N3094);
and AND2 (N19447, N19441, N15518);
nand NAND2 (N19448, N19435, N3609);
not NOT1 (N19449, N19428);
buf BUF1 (N19450, N19426);
xor XOR2 (N19451, N19450, N14370);
nor NOR4 (N19452, N19449, N4262, N11110, N13507);
xor XOR2 (N19453, N19446, N16130);
or OR4 (N19454, N19440, N14913, N15195, N18207);
nor NOR3 (N19455, N19453, N6091, N3938);
buf BUF1 (N19456, N19445);
nor NOR2 (N19457, N19444, N12598);
or OR2 (N19458, N19447, N14225);
nand NAND3 (N19459, N19448, N18126, N16703);
not NOT1 (N19460, N19432);
nand NAND3 (N19461, N19403, N6153, N2019);
buf BUF1 (N19462, N19460);
buf BUF1 (N19463, N19462);
not NOT1 (N19464, N19459);
nor NOR2 (N19465, N19464, N9477);
and AND3 (N19466, N19451, N15056, N4542);
and AND2 (N19467, N19463, N18824);
buf BUF1 (N19468, N19458);
and AND4 (N19469, N19461, N16083, N4653, N1587);
and AND4 (N19470, N19465, N5918, N14090, N15899);
and AND2 (N19471, N19456, N2633);
or OR2 (N19472, N19468, N5119);
buf BUF1 (N19473, N19457);
nand NAND3 (N19474, N19471, N15574, N6376);
not NOT1 (N19475, N19474);
nor NOR3 (N19476, N19473, N18801, N15930);
nor NOR4 (N19477, N19466, N4178, N17848, N11083);
not NOT1 (N19478, N19455);
nor NOR3 (N19479, N19454, N6502, N14261);
nor NOR3 (N19480, N19478, N8548, N13322);
not NOT1 (N19481, N19480);
nor NOR3 (N19482, N19481, N12322, N14254);
and AND3 (N19483, N19467, N12263, N18233);
nor NOR3 (N19484, N19472, N12965, N6394);
buf BUF1 (N19485, N19477);
or OR2 (N19486, N19483, N16593);
buf BUF1 (N19487, N19469);
not NOT1 (N19488, N19485);
nor NOR2 (N19489, N19487, N12498);
and AND4 (N19490, N19486, N6225, N5232, N15575);
buf BUF1 (N19491, N19470);
not NOT1 (N19492, N19488);
nand NAND4 (N19493, N19484, N8762, N16974, N16288);
or OR3 (N19494, N19475, N10356, N12685);
not NOT1 (N19495, N19493);
nand NAND4 (N19496, N19489, N5724, N5548, N16599);
or OR2 (N19497, N19494, N6951);
xor XOR2 (N19498, N19482, N19490);
nand NAND2 (N19499, N7868, N1496);
xor XOR2 (N19500, N19497, N3633);
xor XOR2 (N19501, N19492, N11112);
nand NAND3 (N19502, N19500, N14638, N16703);
not NOT1 (N19503, N19452);
buf BUF1 (N19504, N19476);
and AND2 (N19505, N19498, N17920);
nand NAND4 (N19506, N19503, N2868, N2010, N16871);
and AND2 (N19507, N19496, N12926);
and AND3 (N19508, N19506, N15279, N19239);
xor XOR2 (N19509, N19501, N2591);
nor NOR2 (N19510, N19507, N15055);
xor XOR2 (N19511, N19479, N7802);
buf BUF1 (N19512, N19510);
nor NOR3 (N19513, N19491, N11368, N8010);
or OR4 (N19514, N19509, N9531, N3322, N7859);
or OR4 (N19515, N19502, N10758, N11500, N2219);
nor NOR2 (N19516, N19513, N8921);
xor XOR2 (N19517, N19505, N15698);
xor XOR2 (N19518, N19516, N14022);
nor NOR4 (N19519, N19504, N18805, N11334, N13926);
nor NOR2 (N19520, N19514, N6064);
nand NAND2 (N19521, N19520, N15863);
or OR2 (N19522, N19515, N9632);
not NOT1 (N19523, N19512);
or OR4 (N19524, N19508, N9387, N8273, N12069);
and AND4 (N19525, N19523, N4890, N677, N10008);
not NOT1 (N19526, N19511);
buf BUF1 (N19527, N19525);
xor XOR2 (N19528, N19517, N6275);
buf BUF1 (N19529, N19524);
nand NAND2 (N19530, N19527, N1765);
not NOT1 (N19531, N19528);
buf BUF1 (N19532, N19531);
and AND2 (N19533, N19529, N11415);
xor XOR2 (N19534, N19521, N12146);
and AND3 (N19535, N19526, N11832, N3197);
or OR4 (N19536, N19535, N5392, N15074, N17144);
buf BUF1 (N19537, N19518);
and AND3 (N19538, N19530, N17264, N5930);
nor NOR4 (N19539, N19538, N12404, N15019, N9863);
xor XOR2 (N19540, N19533, N12781);
buf BUF1 (N19541, N19537);
nand NAND4 (N19542, N19532, N16764, N11886, N1191);
and AND3 (N19543, N19539, N1431, N11117);
nand NAND4 (N19544, N19519, N8779, N7762, N12371);
buf BUF1 (N19545, N19534);
xor XOR2 (N19546, N19536, N11357);
xor XOR2 (N19547, N19522, N729);
buf BUF1 (N19548, N19541);
nand NAND2 (N19549, N19543, N1425);
xor XOR2 (N19550, N19542, N8357);
xor XOR2 (N19551, N19550, N16305);
buf BUF1 (N19552, N19549);
nand NAND2 (N19553, N19548, N15379);
nor NOR3 (N19554, N19546, N13881, N11317);
xor XOR2 (N19555, N19540, N15246);
nor NOR2 (N19556, N19545, N4475);
or OR4 (N19557, N19544, N12251, N12117, N15591);
nand NAND4 (N19558, N19495, N7777, N2902, N3227);
nand NAND4 (N19559, N19499, N2489, N2080, N17887);
or OR2 (N19560, N19555, N12998);
buf BUF1 (N19561, N19560);
xor XOR2 (N19562, N19554, N10529);
buf BUF1 (N19563, N19561);
nand NAND2 (N19564, N19547, N15283);
not NOT1 (N19565, N19562);
buf BUF1 (N19566, N19552);
buf BUF1 (N19567, N19564);
and AND2 (N19568, N19559, N12752);
xor XOR2 (N19569, N19568, N6267);
nor NOR4 (N19570, N19551, N14807, N899, N12946);
xor XOR2 (N19571, N19570, N836);
and AND3 (N19572, N19571, N14429, N7214);
xor XOR2 (N19573, N19556, N18802);
buf BUF1 (N19574, N19569);
nor NOR2 (N19575, N19567, N3114);
xor XOR2 (N19576, N19563, N421);
or OR3 (N19577, N19566, N18803, N6352);
not NOT1 (N19578, N19572);
not NOT1 (N19579, N19578);
buf BUF1 (N19580, N19553);
nor NOR3 (N19581, N19576, N6775, N10572);
nor NOR4 (N19582, N19577, N17234, N14585, N484);
buf BUF1 (N19583, N19557);
not NOT1 (N19584, N19575);
nor NOR2 (N19585, N19579, N304);
and AND4 (N19586, N19580, N493, N14005, N1269);
buf BUF1 (N19587, N19573);
xor XOR2 (N19588, N19574, N5088);
xor XOR2 (N19589, N19584, N18106);
xor XOR2 (N19590, N19589, N3363);
and AND4 (N19591, N19558, N16820, N9489, N12841);
or OR2 (N19592, N19582, N13951);
and AND4 (N19593, N19592, N19504, N19131, N1101);
nand NAND3 (N19594, N19590, N8304, N3534);
nand NAND2 (N19595, N19583, N3617);
xor XOR2 (N19596, N19585, N15587);
not NOT1 (N19597, N19565);
nor NOR4 (N19598, N19597, N6415, N7492, N4810);
nand NAND3 (N19599, N19594, N2184, N6656);
nand NAND3 (N19600, N19599, N10552, N5662);
xor XOR2 (N19601, N19593, N14891);
or OR2 (N19602, N19600, N12263);
not NOT1 (N19603, N19598);
and AND2 (N19604, N19601, N15519);
not NOT1 (N19605, N19586);
and AND2 (N19606, N19596, N4427);
or OR4 (N19607, N19587, N6621, N8312, N10560);
xor XOR2 (N19608, N19606, N5819);
and AND2 (N19609, N19607, N8586);
buf BUF1 (N19610, N19603);
xor XOR2 (N19611, N19591, N11278);
and AND2 (N19612, N19595, N11695);
and AND4 (N19613, N19610, N9276, N18895, N18698);
buf BUF1 (N19614, N19608);
or OR2 (N19615, N19604, N2586);
nor NOR3 (N19616, N19614, N5238, N9069);
and AND4 (N19617, N19615, N14012, N16636, N2017);
xor XOR2 (N19618, N19612, N12695);
and AND3 (N19619, N19588, N6743, N2105);
nand NAND2 (N19620, N19619, N16943);
not NOT1 (N19621, N19605);
buf BUF1 (N19622, N19621);
nand NAND3 (N19623, N19581, N14497, N1899);
buf BUF1 (N19624, N19622);
buf BUF1 (N19625, N19616);
nor NOR3 (N19626, N19609, N1187, N16258);
nand NAND2 (N19627, N19617, N3706);
nand NAND4 (N19628, N19620, N11094, N16972, N13396);
not NOT1 (N19629, N19627);
nand NAND2 (N19630, N19618, N16269);
or OR3 (N19631, N19623, N4153, N2967);
xor XOR2 (N19632, N19630, N7388);
xor XOR2 (N19633, N19613, N5935);
and AND2 (N19634, N19631, N19099);
or OR2 (N19635, N19629, N18636);
and AND2 (N19636, N19602, N1572);
nand NAND4 (N19637, N19628, N861, N3487, N17310);
not NOT1 (N19638, N19635);
and AND4 (N19639, N19611, N5739, N8927, N16193);
not NOT1 (N19640, N19626);
or OR4 (N19641, N19625, N10185, N3419, N14921);
nor NOR4 (N19642, N19633, N16097, N6003, N2814);
not NOT1 (N19643, N19636);
or OR4 (N19644, N19641, N9267, N10936, N9199);
nand NAND4 (N19645, N19638, N12124, N8853, N15013);
nand NAND4 (N19646, N19637, N968, N7561, N16338);
and AND2 (N19647, N19645, N12751);
and AND2 (N19648, N19640, N15399);
and AND4 (N19649, N19639, N4957, N14210, N9030);
buf BUF1 (N19650, N19624);
nand NAND3 (N19651, N19648, N4646, N12918);
buf BUF1 (N19652, N19632);
nor NOR3 (N19653, N19646, N6632, N2812);
xor XOR2 (N19654, N19651, N3255);
buf BUF1 (N19655, N19644);
or OR4 (N19656, N19647, N11277, N4720, N2789);
xor XOR2 (N19657, N19653, N5214);
nand NAND2 (N19658, N19656, N4935);
or OR4 (N19659, N19657, N7280, N14058, N11990);
nand NAND4 (N19660, N19634, N4621, N4366, N8992);
not NOT1 (N19661, N19655);
nand NAND2 (N19662, N19660, N17950);
nand NAND4 (N19663, N19649, N1461, N16239, N13782);
nand NAND2 (N19664, N19643, N4155);
not NOT1 (N19665, N19652);
nor NOR4 (N19666, N19658, N16722, N16420, N3448);
or OR2 (N19667, N19664, N8624);
or OR3 (N19668, N19662, N16532, N1754);
and AND2 (N19669, N19659, N7419);
nand NAND3 (N19670, N19661, N4376, N6261);
nor NOR4 (N19671, N19668, N10351, N210, N15188);
nor NOR4 (N19672, N19650, N8450, N10511, N9899);
or OR3 (N19673, N19672, N10857, N10039);
not NOT1 (N19674, N19642);
nor NOR4 (N19675, N19665, N14490, N473, N6720);
nand NAND3 (N19676, N19674, N3880, N720);
nor NOR2 (N19677, N19676, N7963);
nor NOR2 (N19678, N19666, N13988);
and AND3 (N19679, N19675, N10291, N16620);
buf BUF1 (N19680, N19667);
buf BUF1 (N19681, N19663);
not NOT1 (N19682, N19678);
nor NOR3 (N19683, N19670, N10159, N9566);
xor XOR2 (N19684, N19683, N19236);
and AND4 (N19685, N19673, N727, N15821, N13534);
xor XOR2 (N19686, N19680, N2614);
and AND4 (N19687, N19677, N12381, N7964, N15770);
xor XOR2 (N19688, N19671, N9593);
xor XOR2 (N19689, N19654, N13141);
nor NOR2 (N19690, N19684, N472);
not NOT1 (N19691, N19682);
and AND3 (N19692, N19681, N4516, N9834);
xor XOR2 (N19693, N19679, N5116);
xor XOR2 (N19694, N19686, N16058);
nand NAND3 (N19695, N19694, N7207, N4942);
or OR3 (N19696, N19685, N7537, N981);
and AND2 (N19697, N19690, N19243);
nor NOR3 (N19698, N19689, N1040, N18284);
and AND2 (N19699, N19692, N16208);
and AND3 (N19700, N19699, N7893, N12079);
xor XOR2 (N19701, N19688, N2376);
nand NAND3 (N19702, N19687, N1754, N13696);
and AND2 (N19703, N19698, N2455);
xor XOR2 (N19704, N19696, N6415);
nor NOR3 (N19705, N19691, N12504, N15592);
not NOT1 (N19706, N19697);
buf BUF1 (N19707, N19702);
buf BUF1 (N19708, N19700);
xor XOR2 (N19709, N19705, N18629);
nand NAND4 (N19710, N19704, N12864, N18685, N17749);
not NOT1 (N19711, N19669);
buf BUF1 (N19712, N19707);
nor NOR4 (N19713, N19695, N15255, N5029, N9718);
xor XOR2 (N19714, N19701, N8754);
and AND4 (N19715, N19710, N15780, N14909, N9987);
or OR4 (N19716, N19708, N15979, N15917, N4388);
nand NAND3 (N19717, N19716, N4936, N18277);
xor XOR2 (N19718, N19711, N826);
not NOT1 (N19719, N19717);
xor XOR2 (N19720, N19713, N5902);
buf BUF1 (N19721, N19720);
xor XOR2 (N19722, N19709, N19620);
not NOT1 (N19723, N19722);
xor XOR2 (N19724, N19719, N3723);
buf BUF1 (N19725, N19714);
nand NAND2 (N19726, N19718, N10369);
xor XOR2 (N19727, N19715, N17503);
nand NAND2 (N19728, N19712, N19648);
and AND3 (N19729, N19693, N6562, N4976);
not NOT1 (N19730, N19729);
xor XOR2 (N19731, N19727, N19294);
xor XOR2 (N19732, N19725, N9000);
nor NOR4 (N19733, N19728, N9272, N4352, N14752);
buf BUF1 (N19734, N19703);
nor NOR2 (N19735, N19732, N16961);
not NOT1 (N19736, N19724);
nor NOR2 (N19737, N19723, N4969);
and AND3 (N19738, N19733, N15595, N3583);
not NOT1 (N19739, N19738);
not NOT1 (N19740, N19737);
not NOT1 (N19741, N19731);
nand NAND2 (N19742, N19721, N2411);
or OR2 (N19743, N19739, N12643);
nor NOR4 (N19744, N19736, N11152, N3197, N8009);
xor XOR2 (N19745, N19730, N3053);
buf BUF1 (N19746, N19745);
not NOT1 (N19747, N19743);
and AND4 (N19748, N19741, N678, N208, N3262);
or OR2 (N19749, N19747, N274);
nor NOR2 (N19750, N19749, N12730);
buf BUF1 (N19751, N19740);
and AND2 (N19752, N19735, N9955);
nor NOR2 (N19753, N19726, N18139);
nor NOR3 (N19754, N19748, N8345, N14226);
nand NAND3 (N19755, N19742, N19298, N8671);
nor NOR4 (N19756, N19752, N17993, N4833, N10622);
nand NAND4 (N19757, N19750, N18022, N18202, N9963);
xor XOR2 (N19758, N19751, N14786);
not NOT1 (N19759, N19753);
xor XOR2 (N19760, N19754, N5442);
nand NAND3 (N19761, N19759, N2255, N6647);
or OR3 (N19762, N19734, N4146, N8364);
xor XOR2 (N19763, N19760, N13440);
nand NAND4 (N19764, N19744, N18565, N3664, N5351);
buf BUF1 (N19765, N19756);
nor NOR3 (N19766, N19764, N2323, N13269);
buf BUF1 (N19767, N19762);
nor NOR3 (N19768, N19766, N1564, N1496);
buf BUF1 (N19769, N19768);
not NOT1 (N19770, N19755);
not NOT1 (N19771, N19761);
nand NAND4 (N19772, N19770, N156, N16292, N11565);
or OR2 (N19773, N19771, N9616);
xor XOR2 (N19774, N19746, N3639);
or OR2 (N19775, N19767, N10899);
xor XOR2 (N19776, N19773, N12744);
xor XOR2 (N19777, N19772, N18033);
or OR4 (N19778, N19775, N152, N18098, N229);
xor XOR2 (N19779, N19776, N1869);
nand NAND2 (N19780, N19777, N16144);
xor XOR2 (N19781, N19774, N5616);
nand NAND4 (N19782, N19781, N3958, N17289, N3035);
or OR2 (N19783, N19779, N15765);
or OR4 (N19784, N19782, N294, N12563, N8967);
or OR3 (N19785, N19758, N6548, N8134);
and AND4 (N19786, N19769, N13140, N2583, N67);
or OR3 (N19787, N19778, N235, N11809);
nand NAND3 (N19788, N19783, N12176, N10833);
and AND3 (N19789, N19788, N7385, N9525);
not NOT1 (N19790, N19787);
not NOT1 (N19791, N19785);
and AND2 (N19792, N19757, N14905);
nand NAND4 (N19793, N19780, N5294, N17382, N9613);
xor XOR2 (N19794, N19792, N3987);
and AND2 (N19795, N19763, N11281);
and AND4 (N19796, N19793, N8985, N6946, N14731);
and AND3 (N19797, N19784, N5254, N8654);
xor XOR2 (N19798, N19795, N4253);
nand NAND4 (N19799, N19797, N11831, N11238, N15489);
and AND3 (N19800, N19706, N1106, N212);
buf BUF1 (N19801, N19789);
and AND3 (N19802, N19765, N12294, N5247);
or OR2 (N19803, N19790, N3858);
buf BUF1 (N19804, N19801);
nand NAND4 (N19805, N19794, N3246, N19275, N12447);
xor XOR2 (N19806, N19802, N16808);
or OR3 (N19807, N19791, N16305, N18659);
buf BUF1 (N19808, N19786);
buf BUF1 (N19809, N19803);
buf BUF1 (N19810, N19805);
not NOT1 (N19811, N19810);
nand NAND2 (N19812, N19804, N14743);
not NOT1 (N19813, N19807);
buf BUF1 (N19814, N19813);
nor NOR3 (N19815, N19806, N19070, N7214);
nor NOR4 (N19816, N19814, N9650, N5938, N13871);
and AND4 (N19817, N19799, N2546, N1517, N5324);
and AND2 (N19818, N19798, N18887);
nor NOR3 (N19819, N19812, N8341, N7331);
nand NAND2 (N19820, N19819, N17941);
and AND2 (N19821, N19815, N10224);
nor NOR3 (N19822, N19800, N4766, N7580);
nor NOR3 (N19823, N19817, N11879, N15523);
nor NOR3 (N19824, N19808, N13645, N9602);
nor NOR4 (N19825, N19822, N17514, N7778, N14658);
nand NAND3 (N19826, N19818, N13496, N143);
not NOT1 (N19827, N19811);
or OR4 (N19828, N19820, N7805, N14200, N14281);
or OR4 (N19829, N19821, N19588, N4731, N18663);
buf BUF1 (N19830, N19796);
and AND3 (N19831, N19829, N18355, N5989);
or OR2 (N19832, N19828, N18270);
buf BUF1 (N19833, N19809);
not NOT1 (N19834, N19823);
xor XOR2 (N19835, N19816, N3529);
nand NAND3 (N19836, N19833, N3934, N6083);
or OR3 (N19837, N19827, N4026, N4731);
and AND4 (N19838, N19837, N400, N18488, N17735);
buf BUF1 (N19839, N19835);
or OR4 (N19840, N19832, N15322, N8402, N12396);
nor NOR4 (N19841, N19830, N1484, N1752, N7042);
nor NOR2 (N19842, N19834, N13947);
or OR3 (N19843, N19831, N11714, N3912);
buf BUF1 (N19844, N19826);
buf BUF1 (N19845, N19825);
not NOT1 (N19846, N19844);
or OR4 (N19847, N19839, N15688, N9869, N15956);
not NOT1 (N19848, N19838);
not NOT1 (N19849, N19836);
and AND3 (N19850, N19848, N11833, N19693);
xor XOR2 (N19851, N19841, N18011);
xor XOR2 (N19852, N19845, N18484);
or OR3 (N19853, N19851, N1318, N12910);
buf BUF1 (N19854, N19849);
buf BUF1 (N19855, N19847);
nor NOR4 (N19856, N19843, N10390, N18967, N12138);
or OR3 (N19857, N19852, N12619, N540);
and AND3 (N19858, N19824, N1876, N13039);
nor NOR2 (N19859, N19853, N5323);
nor NOR2 (N19860, N19842, N1369);
buf BUF1 (N19861, N19857);
not NOT1 (N19862, N19854);
or OR3 (N19863, N19861, N9135, N4528);
buf BUF1 (N19864, N19850);
and AND2 (N19865, N19864, N11822);
nor NOR4 (N19866, N19865, N7883, N12404, N18536);
nor NOR3 (N19867, N19866, N10427, N7050);
not NOT1 (N19868, N19856);
or OR2 (N19869, N19860, N7436);
nor NOR3 (N19870, N19858, N4511, N10163);
nand NAND3 (N19871, N19867, N19671, N3157);
not NOT1 (N19872, N19868);
xor XOR2 (N19873, N19863, N3992);
nand NAND2 (N19874, N19840, N894);
buf BUF1 (N19875, N19871);
and AND3 (N19876, N19875, N14529, N16851);
not NOT1 (N19877, N19876);
and AND4 (N19878, N19862, N4864, N17928, N1001);
nand NAND4 (N19879, N19859, N10203, N11156, N1478);
or OR3 (N19880, N19846, N3634, N986);
nor NOR3 (N19881, N19879, N9027, N12211);
xor XOR2 (N19882, N19880, N7779);
buf BUF1 (N19883, N19881);
buf BUF1 (N19884, N19874);
xor XOR2 (N19885, N19872, N1263);
xor XOR2 (N19886, N19877, N5632);
nand NAND3 (N19887, N19886, N6557, N3991);
xor XOR2 (N19888, N19869, N11065);
nand NAND3 (N19889, N19884, N11979, N8146);
nand NAND2 (N19890, N19888, N10506);
and AND3 (N19891, N19883, N13077, N8556);
nor NOR4 (N19892, N19870, N2568, N19465, N17745);
nor NOR2 (N19893, N19885, N13346);
buf BUF1 (N19894, N19887);
nand NAND4 (N19895, N19878, N3760, N4336, N5834);
nor NOR4 (N19896, N19855, N14765, N10107, N17165);
nor NOR3 (N19897, N19895, N10324, N9970);
and AND2 (N19898, N19891, N18634);
not NOT1 (N19899, N19897);
xor XOR2 (N19900, N19889, N4859);
not NOT1 (N19901, N19896);
nand NAND4 (N19902, N19898, N16367, N5583, N5576);
not NOT1 (N19903, N19890);
buf BUF1 (N19904, N19882);
not NOT1 (N19905, N19899);
buf BUF1 (N19906, N19904);
xor XOR2 (N19907, N19894, N3976);
buf BUF1 (N19908, N19901);
and AND4 (N19909, N19902, N9222, N1529, N7991);
nor NOR2 (N19910, N19907, N8518);
nand NAND3 (N19911, N19893, N6431, N1141);
nand NAND2 (N19912, N19909, N17616);
nand NAND3 (N19913, N19873, N6286, N1003);
nand NAND3 (N19914, N19911, N6207, N13808);
nand NAND3 (N19915, N19908, N19607, N11976);
xor XOR2 (N19916, N19913, N4136);
or OR3 (N19917, N19915, N9963, N11718);
nor NOR4 (N19918, N19905, N8073, N9895, N12039);
buf BUF1 (N19919, N19906);
or OR2 (N19920, N19916, N16260);
or OR2 (N19921, N19910, N4499);
nor NOR3 (N19922, N19903, N15078, N891);
buf BUF1 (N19923, N19922);
and AND3 (N19924, N19912, N8030, N10732);
not NOT1 (N19925, N19918);
or OR4 (N19926, N19923, N8101, N1624, N919);
nand NAND4 (N19927, N19925, N9114, N15720, N8743);
nand NAND3 (N19928, N19921, N2413, N7539);
nor NOR4 (N19929, N19928, N19817, N8961, N11974);
and AND2 (N19930, N19892, N17351);
nor NOR4 (N19931, N19927, N11811, N11009, N7512);
nor NOR2 (N19932, N19920, N8167);
xor XOR2 (N19933, N19900, N11776);
nor NOR4 (N19934, N19926, N16120, N13501, N16941);
nor NOR3 (N19935, N19932, N3498, N1545);
or OR4 (N19936, N19929, N11808, N1436, N18860);
and AND4 (N19937, N19914, N16692, N4341, N1837);
xor XOR2 (N19938, N19936, N15508);
and AND3 (N19939, N19938, N12996, N8111);
and AND3 (N19940, N19919, N16118, N8966);
nand NAND2 (N19941, N19917, N12116);
nor NOR4 (N19942, N19930, N9664, N2636, N2151);
nor NOR3 (N19943, N19924, N1663, N7664);
nand NAND3 (N19944, N19934, N19287, N8668);
nor NOR4 (N19945, N19935, N1261, N10761, N16598);
xor XOR2 (N19946, N19937, N3726);
and AND2 (N19947, N19943, N12209);
not NOT1 (N19948, N19931);
buf BUF1 (N19949, N19939);
nand NAND4 (N19950, N19947, N10668, N4061, N2625);
or OR3 (N19951, N19944, N934, N15308);
and AND3 (N19952, N19950, N10391, N19665);
xor XOR2 (N19953, N19942, N9844);
and AND3 (N19954, N19949, N17512, N12881);
nor NOR4 (N19955, N19941, N5153, N11688, N12925);
nor NOR4 (N19956, N19953, N19699, N7123, N4960);
nor NOR4 (N19957, N19954, N3163, N19677, N6311);
or OR2 (N19958, N19945, N11353);
or OR2 (N19959, N19958, N7186);
nand NAND3 (N19960, N19948, N2451, N4706);
nand NAND4 (N19961, N19957, N6376, N19392, N6516);
xor XOR2 (N19962, N19940, N10468);
nand NAND2 (N19963, N19959, N6054);
nor NOR2 (N19964, N19955, N11506);
not NOT1 (N19965, N19962);
not NOT1 (N19966, N19946);
not NOT1 (N19967, N19961);
nor NOR2 (N19968, N19956, N2119);
nor NOR4 (N19969, N19933, N7217, N15384, N7500);
xor XOR2 (N19970, N19960, N6674);
not NOT1 (N19971, N19951);
buf BUF1 (N19972, N19969);
and AND2 (N19973, N19968, N7007);
nor NOR4 (N19974, N19967, N13622, N6986, N509);
nand NAND2 (N19975, N19972, N11274);
or OR4 (N19976, N19964, N8822, N13734, N14188);
or OR4 (N19977, N19976, N14546, N7303, N3124);
xor XOR2 (N19978, N19966, N3569);
nand NAND3 (N19979, N19978, N11679, N19173);
nand NAND2 (N19980, N19973, N10205);
nor NOR4 (N19981, N19965, N13243, N8987, N6675);
buf BUF1 (N19982, N19971);
xor XOR2 (N19983, N19977, N3797);
nor NOR2 (N19984, N19952, N10216);
nor NOR2 (N19985, N19975, N14109);
buf BUF1 (N19986, N19970);
buf BUF1 (N19987, N19983);
buf BUF1 (N19988, N19981);
and AND3 (N19989, N19982, N6441, N6363);
or OR2 (N19990, N19987, N19481);
xor XOR2 (N19991, N19988, N18827);
nor NOR3 (N19992, N19989, N19769, N11963);
xor XOR2 (N19993, N19979, N11138);
nand NAND2 (N19994, N19992, N8825);
nor NOR3 (N19995, N19994, N8232, N11718);
or OR4 (N19996, N19993, N18314, N2149, N5291);
nor NOR2 (N19997, N19985, N11276);
xor XOR2 (N19998, N19997, N19547);
or OR4 (N19999, N19974, N12240, N18826, N15150);
and AND3 (N20000, N19980, N10915, N14730);
buf BUF1 (N20001, N19998);
buf BUF1 (N20002, N19990);
and AND3 (N20003, N19986, N7159, N16405);
nor NOR2 (N20004, N19984, N9896);
buf BUF1 (N20005, N20000);
or OR2 (N20006, N19963, N17357);
not NOT1 (N20007, N19999);
and AND2 (N20008, N19991, N995);
buf BUF1 (N20009, N20004);
xor XOR2 (N20010, N19995, N15425);
and AND3 (N20011, N20003, N4502, N505);
or OR3 (N20012, N20005, N19710, N3298);
xor XOR2 (N20013, N20008, N12252);
nor NOR4 (N20014, N20011, N238, N4491, N3141);
or OR3 (N20015, N20012, N15239, N9874);
and AND4 (N20016, N20009, N13155, N919, N719);
nand NAND4 (N20017, N20014, N16640, N12373, N4818);
not NOT1 (N20018, N20013);
xor XOR2 (N20019, N20001, N6746);
buf BUF1 (N20020, N19996);
not NOT1 (N20021, N20006);
buf BUF1 (N20022, N20007);
nand NAND2 (N20023, N20016, N12971);
and AND2 (N20024, N20015, N1649);
and AND4 (N20025, N20022, N16, N15945, N8796);
nand NAND4 (N20026, N20019, N17654, N15874, N17169);
xor XOR2 (N20027, N20018, N3789);
xor XOR2 (N20028, N20020, N17547);
and AND2 (N20029, N20017, N10636);
or OR2 (N20030, N20024, N7496);
nand NAND2 (N20031, N20028, N1784);
and AND3 (N20032, N20021, N4057, N2463);
buf BUF1 (N20033, N20030);
buf BUF1 (N20034, N20023);
or OR3 (N20035, N20010, N15180, N17759);
not NOT1 (N20036, N20032);
not NOT1 (N20037, N20035);
xor XOR2 (N20038, N20037, N9205);
nand NAND3 (N20039, N20038, N4273, N11909);
not NOT1 (N20040, N20039);
nor NOR3 (N20041, N20036, N10442, N12390);
nand NAND3 (N20042, N20027, N9334, N10504);
or OR2 (N20043, N20041, N3009);
nor NOR4 (N20044, N20033, N5116, N15069, N3847);
nand NAND2 (N20045, N20025, N7994);
xor XOR2 (N20046, N20045, N2407);
or OR4 (N20047, N20043, N3715, N14215, N7354);
nand NAND2 (N20048, N20040, N3464);
or OR3 (N20049, N20048, N15192, N18794);
nor NOR4 (N20050, N20049, N468, N9400, N12234);
not NOT1 (N20051, N20044);
or OR4 (N20052, N20042, N15072, N1068, N16205);
nand NAND2 (N20053, N20026, N8173);
nor NOR3 (N20054, N20029, N5614, N16625);
buf BUF1 (N20055, N20053);
not NOT1 (N20056, N20054);
not NOT1 (N20057, N20034);
and AND2 (N20058, N20055, N3483);
not NOT1 (N20059, N20056);
nand NAND2 (N20060, N20050, N13278);
nand NAND4 (N20061, N20058, N8762, N2735, N9502);
and AND2 (N20062, N20031, N1317);
and AND3 (N20063, N20051, N15686, N17508);
buf BUF1 (N20064, N20052);
or OR2 (N20065, N20002, N14313);
not NOT1 (N20066, N20059);
nor NOR3 (N20067, N20047, N15513, N313);
buf BUF1 (N20068, N20062);
nand NAND2 (N20069, N20057, N9159);
or OR2 (N20070, N20068, N14740);
and AND4 (N20071, N20046, N14740, N18512, N14527);
buf BUF1 (N20072, N20061);
nor NOR3 (N20073, N20065, N4662, N6105);
not NOT1 (N20074, N20064);
nand NAND3 (N20075, N20060, N6683, N8517);
and AND2 (N20076, N20066, N1766);
buf BUF1 (N20077, N20067);
nor NOR3 (N20078, N20073, N3928, N12808);
nand NAND3 (N20079, N20063, N13112, N4900);
not NOT1 (N20080, N20078);
and AND4 (N20081, N20071, N12086, N2228, N952);
nand NAND4 (N20082, N20075, N8175, N906, N16348);
nor NOR2 (N20083, N20069, N16309);
nor NOR2 (N20084, N20081, N12553);
not NOT1 (N20085, N20076);
nor NOR3 (N20086, N20082, N6219, N257);
xor XOR2 (N20087, N20077, N3422);
not NOT1 (N20088, N20086);
buf BUF1 (N20089, N20079);
and AND3 (N20090, N20088, N13036, N10171);
nor NOR4 (N20091, N20090, N4665, N13518, N1755);
nor NOR2 (N20092, N20074, N1040);
and AND2 (N20093, N20080, N18421);
buf BUF1 (N20094, N20091);
not NOT1 (N20095, N20085);
xor XOR2 (N20096, N20084, N11443);
and AND4 (N20097, N20070, N333, N9976, N19794);
or OR2 (N20098, N20083, N10728);
nor NOR2 (N20099, N20095, N6969);
buf BUF1 (N20100, N20072);
or OR4 (N20101, N20100, N6520, N3024, N18448);
xor XOR2 (N20102, N20087, N12244);
not NOT1 (N20103, N20093);
buf BUF1 (N20104, N20099);
buf BUF1 (N20105, N20098);
xor XOR2 (N20106, N20102, N19275);
or OR4 (N20107, N20103, N9876, N17556, N9827);
nand NAND2 (N20108, N20104, N14056);
or OR3 (N20109, N20105, N11814, N2925);
nand NAND4 (N20110, N20092, N11341, N6772, N11937);
nand NAND4 (N20111, N20101, N15298, N15032, N3921);
and AND4 (N20112, N20108, N11079, N6097, N6110);
not NOT1 (N20113, N20110);
and AND3 (N20114, N20112, N173, N2345);
xor XOR2 (N20115, N20114, N9400);
xor XOR2 (N20116, N20097, N1839);
and AND4 (N20117, N20096, N1976, N3967, N11619);
xor XOR2 (N20118, N20089, N6440);
or OR2 (N20119, N20094, N4572);
not NOT1 (N20120, N20117);
nand NAND4 (N20121, N20113, N10493, N16039, N8601);
or OR2 (N20122, N20115, N18016);
and AND2 (N20123, N20107, N17555);
nor NOR2 (N20124, N20109, N17661);
xor XOR2 (N20125, N20106, N2548);
not NOT1 (N20126, N20111);
buf BUF1 (N20127, N20120);
buf BUF1 (N20128, N20121);
xor XOR2 (N20129, N20127, N14667);
and AND3 (N20130, N20129, N1871, N9811);
nor NOR3 (N20131, N20126, N1327, N11032);
buf BUF1 (N20132, N20116);
or OR2 (N20133, N20118, N11040);
and AND3 (N20134, N20133, N16877, N14562);
xor XOR2 (N20135, N20131, N8673);
nand NAND3 (N20136, N20135, N18935, N5902);
nor NOR4 (N20137, N20134, N1484, N13842, N7074);
and AND4 (N20138, N20124, N6245, N7295, N10366);
buf BUF1 (N20139, N20138);
buf BUF1 (N20140, N20132);
not NOT1 (N20141, N20125);
xor XOR2 (N20142, N20119, N18040);
and AND3 (N20143, N20123, N11701, N2198);
xor XOR2 (N20144, N20122, N18277);
nor NOR4 (N20145, N20130, N798, N17691, N8810);
or OR2 (N20146, N20136, N4061);
and AND3 (N20147, N20139, N15557, N17024);
and AND4 (N20148, N20140, N8775, N5116, N13442);
buf BUF1 (N20149, N20143);
buf BUF1 (N20150, N20144);
and AND4 (N20151, N20128, N14481, N5788, N7107);
nand NAND4 (N20152, N20146, N11719, N18953, N3634);
buf BUF1 (N20153, N20148);
and AND4 (N20154, N20147, N5974, N7752, N4502);
not NOT1 (N20155, N20153);
not NOT1 (N20156, N20149);
nand NAND4 (N20157, N20155, N4422, N326, N9084);
not NOT1 (N20158, N20150);
nand NAND2 (N20159, N20157, N2157);
not NOT1 (N20160, N20151);
buf BUF1 (N20161, N20145);
buf BUF1 (N20162, N20158);
and AND4 (N20163, N20159, N20116, N1714, N3142);
or OR3 (N20164, N20161, N10590, N15269);
or OR2 (N20165, N20152, N5987);
and AND4 (N20166, N20141, N8335, N9290, N5459);
buf BUF1 (N20167, N20154);
buf BUF1 (N20168, N20137);
nand NAND4 (N20169, N20163, N1580, N1557, N12083);
nor NOR2 (N20170, N20165, N7527);
nand NAND3 (N20171, N20164, N18366, N11953);
not NOT1 (N20172, N20168);
nand NAND4 (N20173, N20142, N18012, N4037, N7513);
or OR4 (N20174, N20156, N1609, N14073, N17868);
not NOT1 (N20175, N20160);
nand NAND4 (N20176, N20173, N14972, N18006, N3620);
and AND3 (N20177, N20169, N15711, N17033);
not NOT1 (N20178, N20177);
buf BUF1 (N20179, N20174);
nand NAND2 (N20180, N20162, N116);
buf BUF1 (N20181, N20175);
buf BUF1 (N20182, N20176);
nor NOR2 (N20183, N20166, N10540);
nor NOR3 (N20184, N20170, N14769, N11880);
xor XOR2 (N20185, N20178, N14202);
not NOT1 (N20186, N20179);
nor NOR4 (N20187, N20181, N17597, N9066, N12363);
or OR4 (N20188, N20186, N17393, N11339, N12070);
not NOT1 (N20189, N20187);
or OR2 (N20190, N20185, N9617);
not NOT1 (N20191, N20171);
and AND2 (N20192, N20191, N13232);
and AND3 (N20193, N20180, N12903, N18656);
not NOT1 (N20194, N20192);
buf BUF1 (N20195, N20182);
buf BUF1 (N20196, N20195);
or OR3 (N20197, N20194, N3790, N20002);
nor NOR2 (N20198, N20193, N18114);
nor NOR3 (N20199, N20188, N15612, N3927);
buf BUF1 (N20200, N20167);
buf BUF1 (N20201, N20198);
xor XOR2 (N20202, N20184, N20188);
or OR3 (N20203, N20189, N18736, N928);
buf BUF1 (N20204, N20190);
and AND4 (N20205, N20202, N23, N2232, N101);
nor NOR4 (N20206, N20199, N7424, N3947, N3721);
buf BUF1 (N20207, N20204);
nand NAND2 (N20208, N20206, N864);
and AND4 (N20209, N20205, N18364, N13853, N8204);
and AND3 (N20210, N20172, N7130, N11622);
or OR3 (N20211, N20197, N383, N1493);
buf BUF1 (N20212, N20210);
or OR4 (N20213, N20207, N13056, N7597, N3965);
nor NOR2 (N20214, N20209, N1190);
buf BUF1 (N20215, N20196);
not NOT1 (N20216, N20213);
nor NOR3 (N20217, N20203, N11356, N4239);
and AND3 (N20218, N20216, N2658, N10783);
or OR3 (N20219, N20218, N11071, N14508);
and AND2 (N20220, N20183, N13937);
or OR4 (N20221, N20217, N2232, N5704, N14838);
xor XOR2 (N20222, N20219, N19955);
nand NAND4 (N20223, N20221, N5740, N8569, N1370);
not NOT1 (N20224, N20222);
and AND2 (N20225, N20223, N3756);
not NOT1 (N20226, N20212);
xor XOR2 (N20227, N20220, N18471);
or OR2 (N20228, N20215, N17199);
nor NOR3 (N20229, N20225, N1521, N17160);
xor XOR2 (N20230, N20227, N17954);
xor XOR2 (N20231, N20214, N19635);
xor XOR2 (N20232, N20201, N19561);
nor NOR3 (N20233, N20211, N19755, N7049);
buf BUF1 (N20234, N20200);
xor XOR2 (N20235, N20224, N11314);
or OR2 (N20236, N20235, N14917);
nor NOR2 (N20237, N20230, N10293);
buf BUF1 (N20238, N20208);
buf BUF1 (N20239, N20228);
or OR2 (N20240, N20226, N16845);
buf BUF1 (N20241, N20240);
not NOT1 (N20242, N20239);
nand NAND2 (N20243, N20236, N19169);
buf BUF1 (N20244, N20234);
and AND4 (N20245, N20238, N6444, N13495, N19020);
xor XOR2 (N20246, N20244, N7930);
not NOT1 (N20247, N20245);
not NOT1 (N20248, N20242);
or OR4 (N20249, N20232, N8533, N6569, N10288);
or OR3 (N20250, N20243, N6252, N16002);
xor XOR2 (N20251, N20248, N19658);
xor XOR2 (N20252, N20231, N3434);
xor XOR2 (N20253, N20229, N17959);
nand NAND2 (N20254, N20246, N8206);
nor NOR3 (N20255, N20252, N19908, N2088);
and AND3 (N20256, N20247, N2486, N10815);
buf BUF1 (N20257, N20250);
not NOT1 (N20258, N20233);
or OR4 (N20259, N20255, N16222, N19616, N9307);
and AND2 (N20260, N20251, N13339);
not NOT1 (N20261, N20254);
nor NOR4 (N20262, N20261, N10132, N16789, N5379);
or OR4 (N20263, N20256, N8600, N8937, N17360);
not NOT1 (N20264, N20263);
or OR3 (N20265, N20249, N8166, N3533);
nand NAND2 (N20266, N20259, N9471);
nand NAND2 (N20267, N20265, N19521);
and AND3 (N20268, N20264, N16406, N19652);
not NOT1 (N20269, N20260);
and AND4 (N20270, N20267, N4200, N10322, N7035);
buf BUF1 (N20271, N20257);
nand NAND2 (N20272, N20269, N16);
not NOT1 (N20273, N20258);
or OR3 (N20274, N20262, N1932, N3310);
nor NOR4 (N20275, N20270, N2600, N8006, N16048);
nand NAND2 (N20276, N20268, N18108);
buf BUF1 (N20277, N20271);
nor NOR3 (N20278, N20276, N4982, N13180);
and AND2 (N20279, N20278, N17607);
not NOT1 (N20280, N20279);
xor XOR2 (N20281, N20237, N5429);
and AND2 (N20282, N20275, N1310);
nand NAND3 (N20283, N20272, N12818, N4632);
not NOT1 (N20284, N20277);
xor XOR2 (N20285, N20283, N451);
buf BUF1 (N20286, N20280);
nor NOR2 (N20287, N20241, N2837);
buf BUF1 (N20288, N20274);
not NOT1 (N20289, N20286);
nor NOR3 (N20290, N20287, N19870, N7874);
xor XOR2 (N20291, N20266, N18957);
buf BUF1 (N20292, N20281);
or OR4 (N20293, N20284, N17600, N1325, N7368);
or OR4 (N20294, N20285, N18432, N11627, N14599);
nor NOR2 (N20295, N20289, N14700);
or OR3 (N20296, N20288, N8682, N18069);
buf BUF1 (N20297, N20253);
not NOT1 (N20298, N20292);
xor XOR2 (N20299, N20293, N6323);
nor NOR3 (N20300, N20297, N1066, N14158);
nor NOR2 (N20301, N20290, N18293);
not NOT1 (N20302, N20282);
buf BUF1 (N20303, N20294);
buf BUF1 (N20304, N20301);
buf BUF1 (N20305, N20304);
buf BUF1 (N20306, N20295);
nand NAND2 (N20307, N20298, N9155);
nand NAND3 (N20308, N20303, N3935, N1082);
nand NAND2 (N20309, N20299, N7118);
and AND2 (N20310, N20273, N5569);
nor NOR4 (N20311, N20307, N12043, N2066, N10582);
or OR3 (N20312, N20309, N7057, N13788);
buf BUF1 (N20313, N20305);
or OR3 (N20314, N20311, N6063, N13757);
not NOT1 (N20315, N20291);
or OR3 (N20316, N20306, N16790, N802);
nor NOR2 (N20317, N20310, N6484);
nor NOR2 (N20318, N20312, N16868);
and AND2 (N20319, N20313, N7990);
or OR4 (N20320, N20318, N17995, N8461, N5540);
xor XOR2 (N20321, N20320, N4751);
and AND2 (N20322, N20314, N8143);
or OR2 (N20323, N20300, N5538);
nand NAND2 (N20324, N20322, N1087);
or OR3 (N20325, N20308, N11934, N5683);
or OR3 (N20326, N20302, N20259, N3131);
nor NOR4 (N20327, N20324, N3402, N2744, N11722);
or OR4 (N20328, N20315, N18562, N13163, N2684);
nand NAND3 (N20329, N20317, N17747, N19009);
nor NOR2 (N20330, N20321, N12071);
nand NAND4 (N20331, N20326, N13913, N13904, N11003);
not NOT1 (N20332, N20327);
buf BUF1 (N20333, N20328);
not NOT1 (N20334, N20319);
buf BUF1 (N20335, N20325);
buf BUF1 (N20336, N20323);
buf BUF1 (N20337, N20335);
buf BUF1 (N20338, N20316);
and AND4 (N20339, N20333, N16518, N2309, N10910);
and AND4 (N20340, N20338, N7137, N4790, N15045);
nor NOR4 (N20341, N20332, N4111, N2588, N5445);
or OR4 (N20342, N20334, N10676, N16609, N19579);
and AND2 (N20343, N20342, N11484);
nand NAND3 (N20344, N20331, N3116, N6964);
buf BUF1 (N20345, N20341);
nand NAND3 (N20346, N20344, N14872, N2866);
or OR3 (N20347, N20337, N15888, N11650);
not NOT1 (N20348, N20330);
nand NAND2 (N20349, N20339, N2331);
nand NAND2 (N20350, N20340, N8521);
nor NOR3 (N20351, N20348, N5731, N2588);
not NOT1 (N20352, N20329);
or OR2 (N20353, N20347, N18665);
not NOT1 (N20354, N20353);
xor XOR2 (N20355, N20343, N8685);
buf BUF1 (N20356, N20336);
nand NAND4 (N20357, N20355, N5106, N10287, N4753);
nor NOR3 (N20358, N20352, N16087, N12325);
or OR4 (N20359, N20351, N17899, N8432, N7769);
and AND4 (N20360, N20345, N197, N3939, N3105);
or OR4 (N20361, N20360, N2733, N13108, N5777);
not NOT1 (N20362, N20349);
buf BUF1 (N20363, N20358);
buf BUF1 (N20364, N20346);
and AND2 (N20365, N20356, N16209);
or OR3 (N20366, N20354, N7343, N20059);
not NOT1 (N20367, N20350);
buf BUF1 (N20368, N20366);
or OR2 (N20369, N20365, N11856);
or OR4 (N20370, N20359, N17499, N10382, N5136);
buf BUF1 (N20371, N20296);
not NOT1 (N20372, N20368);
nand NAND2 (N20373, N20369, N636);
nand NAND4 (N20374, N20362, N10972, N19039, N19524);
not NOT1 (N20375, N20370);
xor XOR2 (N20376, N20371, N17597);
nor NOR4 (N20377, N20367, N5545, N14877, N7562);
nand NAND3 (N20378, N20375, N12031, N6936);
not NOT1 (N20379, N20374);
and AND4 (N20380, N20373, N9247, N7918, N20272);
xor XOR2 (N20381, N20379, N15517);
nor NOR4 (N20382, N20364, N19681, N14787, N3191);
nor NOR2 (N20383, N20380, N11366);
or OR3 (N20384, N20372, N841, N76);
nand NAND3 (N20385, N20382, N1779, N10984);
or OR4 (N20386, N20377, N13850, N13074, N3837);
or OR2 (N20387, N20384, N102);
nor NOR2 (N20388, N20381, N12287);
nor NOR4 (N20389, N20388, N20339, N39, N3497);
and AND3 (N20390, N20361, N5401, N3143);
nand NAND3 (N20391, N20363, N1318, N13616);
xor XOR2 (N20392, N20383, N12491);
xor XOR2 (N20393, N20376, N18056);
or OR3 (N20394, N20393, N9069, N14226);
not NOT1 (N20395, N20357);
and AND4 (N20396, N20387, N15648, N19298, N7891);
and AND4 (N20397, N20396, N5160, N14398, N4958);
nand NAND4 (N20398, N20378, N243, N19727, N12870);
and AND2 (N20399, N20394, N579);
and AND3 (N20400, N20398, N17448, N8659);
not NOT1 (N20401, N20385);
xor XOR2 (N20402, N20399, N1588);
buf BUF1 (N20403, N20386);
xor XOR2 (N20404, N20390, N17559);
nand NAND3 (N20405, N20403, N2579, N9358);
not NOT1 (N20406, N20400);
and AND2 (N20407, N20392, N386);
nand NAND2 (N20408, N20407, N15785);
not NOT1 (N20409, N20406);
nor NOR3 (N20410, N20405, N17574, N1830);
nor NOR4 (N20411, N20409, N3086, N16485, N19331);
nand NAND4 (N20412, N20401, N16522, N17964, N1190);
or OR2 (N20413, N20404, N13226);
not NOT1 (N20414, N20389);
and AND2 (N20415, N20412, N19303);
and AND2 (N20416, N20413, N17529);
xor XOR2 (N20417, N20402, N6120);
nor NOR4 (N20418, N20410, N8407, N9637, N6081);
and AND2 (N20419, N20416, N14620);
xor XOR2 (N20420, N20395, N9821);
or OR2 (N20421, N20397, N11422);
or OR3 (N20422, N20418, N10616, N3409);
or OR3 (N20423, N20417, N8716, N3377);
nand NAND3 (N20424, N20411, N1929, N20059);
xor XOR2 (N20425, N20422, N11365);
not NOT1 (N20426, N20414);
not NOT1 (N20427, N20425);
nand NAND2 (N20428, N20420, N14404);
buf BUF1 (N20429, N20428);
xor XOR2 (N20430, N20424, N13341);
not NOT1 (N20431, N20421);
xor XOR2 (N20432, N20419, N9296);
buf BUF1 (N20433, N20426);
buf BUF1 (N20434, N20427);
nor NOR3 (N20435, N20434, N19321, N12223);
and AND3 (N20436, N20415, N5799, N13328);
buf BUF1 (N20437, N20435);
nand NAND2 (N20438, N20423, N18766);
nor NOR2 (N20439, N20391, N5059);
or OR3 (N20440, N20436, N15523, N18092);
or OR3 (N20441, N20438, N8096, N5182);
or OR3 (N20442, N20431, N19698, N12781);
buf BUF1 (N20443, N20433);
and AND4 (N20444, N20441, N15220, N16351, N1821);
buf BUF1 (N20445, N20429);
buf BUF1 (N20446, N20442);
and AND2 (N20447, N20437, N10395);
and AND2 (N20448, N20432, N3893);
and AND3 (N20449, N20408, N726, N7595);
and AND2 (N20450, N20449, N12379);
or OR4 (N20451, N20445, N20208, N316, N19035);
or OR3 (N20452, N20440, N17102, N14846);
not NOT1 (N20453, N20430);
buf BUF1 (N20454, N20450);
buf BUF1 (N20455, N20448);
nand NAND3 (N20456, N20443, N1480, N20378);
not NOT1 (N20457, N20453);
and AND4 (N20458, N20451, N3518, N3940, N10627);
or OR2 (N20459, N20455, N1318);
and AND2 (N20460, N20439, N13782);
buf BUF1 (N20461, N20460);
xor XOR2 (N20462, N20458, N1121);
nand NAND2 (N20463, N20456, N6590);
nor NOR4 (N20464, N20461, N6570, N18618, N11140);
xor XOR2 (N20465, N20457, N7599);
and AND4 (N20466, N20462, N1566, N8343, N9334);
or OR3 (N20467, N20454, N1426, N18075);
not NOT1 (N20468, N20446);
not NOT1 (N20469, N20467);
not NOT1 (N20470, N20452);
and AND3 (N20471, N20465, N13043, N13653);
and AND3 (N20472, N20463, N16427, N9606);
not NOT1 (N20473, N20464);
buf BUF1 (N20474, N20469);
not NOT1 (N20475, N20459);
xor XOR2 (N20476, N20444, N206);
or OR4 (N20477, N20468, N8890, N9768, N5208);
or OR4 (N20478, N20475, N9577, N4644, N437);
nand NAND2 (N20479, N20472, N13507);
buf BUF1 (N20480, N20466);
or OR3 (N20481, N20474, N11101, N16127);
nand NAND2 (N20482, N20470, N20401);
nand NAND3 (N20483, N20447, N2945, N10920);
nand NAND3 (N20484, N20471, N13539, N16031);
or OR4 (N20485, N20479, N19823, N9013, N4221);
buf BUF1 (N20486, N20477);
nor NOR2 (N20487, N20481, N4289);
and AND4 (N20488, N20487, N10228, N8220, N11673);
or OR3 (N20489, N20476, N1662, N5051);
buf BUF1 (N20490, N20478);
and AND2 (N20491, N20484, N12812);
or OR2 (N20492, N20488, N471);
not NOT1 (N20493, N20486);
or OR2 (N20494, N20492, N16451);
nand NAND2 (N20495, N20493, N18107);
or OR4 (N20496, N20494, N13360, N16671, N10806);
or OR4 (N20497, N20491, N13518, N7106, N11243);
or OR3 (N20498, N20497, N8133, N12261);
xor XOR2 (N20499, N20482, N19235);
xor XOR2 (N20500, N20496, N13070);
nor NOR2 (N20501, N20499, N7711);
buf BUF1 (N20502, N20495);
xor XOR2 (N20503, N20501, N13437);
or OR2 (N20504, N20473, N8149);
nand NAND3 (N20505, N20485, N9738, N16802);
or OR4 (N20506, N20498, N968, N7628, N11507);
buf BUF1 (N20507, N20502);
nand NAND3 (N20508, N20503, N9840, N14059);
not NOT1 (N20509, N20505);
or OR4 (N20510, N20506, N7371, N10548, N13657);
nand NAND3 (N20511, N20500, N18382, N16307);
nand NAND3 (N20512, N20509, N5745, N15513);
buf BUF1 (N20513, N20512);
xor XOR2 (N20514, N20490, N6590);
and AND4 (N20515, N20483, N9350, N16702, N8366);
buf BUF1 (N20516, N20507);
nand NAND4 (N20517, N20516, N11454, N15042, N18441);
nor NOR3 (N20518, N20504, N12396, N18420);
not NOT1 (N20519, N20515);
and AND4 (N20520, N20480, N9206, N7465, N5466);
and AND4 (N20521, N20508, N3277, N10962, N7281);
and AND3 (N20522, N20518, N11192, N2347);
nor NOR4 (N20523, N20519, N3068, N6841, N20478);
nand NAND4 (N20524, N20511, N11677, N13882, N3572);
nor NOR2 (N20525, N20523, N987);
and AND4 (N20526, N20522, N17069, N18279, N11633);
not NOT1 (N20527, N20514);
buf BUF1 (N20528, N20520);
nor NOR3 (N20529, N20510, N19764, N3910);
nand NAND2 (N20530, N20526, N15748);
and AND2 (N20531, N20530, N1515);
xor XOR2 (N20532, N20521, N14308);
buf BUF1 (N20533, N20524);
nor NOR3 (N20534, N20525, N19435, N1588);
xor XOR2 (N20535, N20517, N5939);
and AND2 (N20536, N20532, N19206);
or OR3 (N20537, N20489, N1128, N9565);
nor NOR3 (N20538, N20531, N15687, N1188);
not NOT1 (N20539, N20537);
xor XOR2 (N20540, N20529, N10716);
xor XOR2 (N20541, N20536, N14720);
xor XOR2 (N20542, N20528, N13871);
xor XOR2 (N20543, N20538, N6833);
nand NAND3 (N20544, N20527, N9140, N8161);
and AND3 (N20545, N20533, N9367, N20321);
and AND3 (N20546, N20544, N19797, N9629);
not NOT1 (N20547, N20535);
nand NAND2 (N20548, N20539, N1298);
or OR2 (N20549, N20545, N14063);
and AND4 (N20550, N20542, N19423, N264, N13665);
or OR4 (N20551, N20548, N17063, N13861, N16713);
xor XOR2 (N20552, N20540, N11657);
nand NAND2 (N20553, N20552, N12805);
nor NOR4 (N20554, N20546, N1616, N14004, N4978);
xor XOR2 (N20555, N20550, N15688);
and AND2 (N20556, N20554, N172);
nand NAND2 (N20557, N20547, N8624);
and AND4 (N20558, N20534, N3137, N8990, N8689);
or OR2 (N20559, N20556, N6524);
xor XOR2 (N20560, N20558, N9888);
nand NAND3 (N20561, N20549, N15688, N3129);
or OR4 (N20562, N20513, N16855, N690, N4832);
and AND3 (N20563, N20561, N9903, N5894);
not NOT1 (N20564, N20563);
not NOT1 (N20565, N20543);
not NOT1 (N20566, N20551);
not NOT1 (N20567, N20557);
buf BUF1 (N20568, N20559);
or OR2 (N20569, N20568, N15734);
nand NAND3 (N20570, N20562, N3362, N20318);
or OR2 (N20571, N20567, N19526);
nand NAND3 (N20572, N20566, N5412, N10850);
nor NOR4 (N20573, N20564, N5352, N10057, N6853);
nor NOR2 (N20574, N20541, N18887);
xor XOR2 (N20575, N20574, N12605);
not NOT1 (N20576, N20572);
xor XOR2 (N20577, N20571, N6663);
xor XOR2 (N20578, N20553, N7332);
buf BUF1 (N20579, N20576);
not NOT1 (N20580, N20565);
not NOT1 (N20581, N20577);
xor XOR2 (N20582, N20555, N8508);
nand NAND2 (N20583, N20579, N16992);
not NOT1 (N20584, N20581);
xor XOR2 (N20585, N20573, N7259);
buf BUF1 (N20586, N20585);
or OR2 (N20587, N20586, N7301);
not NOT1 (N20588, N20584);
nor NOR3 (N20589, N20587, N10390, N20154);
not NOT1 (N20590, N20570);
not NOT1 (N20591, N20590);
not NOT1 (N20592, N20583);
or OR4 (N20593, N20560, N8347, N18865, N13715);
not NOT1 (N20594, N20582);
xor XOR2 (N20595, N20588, N3673);
buf BUF1 (N20596, N20595);
nor NOR4 (N20597, N20592, N9949, N19521, N541);
not NOT1 (N20598, N20594);
nand NAND4 (N20599, N20589, N11170, N10877, N3124);
buf BUF1 (N20600, N20575);
buf BUF1 (N20601, N20599);
nand NAND4 (N20602, N20569, N18162, N2778, N19086);
nand NAND2 (N20603, N20598, N10061);
and AND4 (N20604, N20601, N17465, N849, N386);
nand NAND3 (N20605, N20578, N1738, N11191);
nand NAND3 (N20606, N20591, N15316, N18301);
or OR4 (N20607, N20602, N16470, N20298, N221);
not NOT1 (N20608, N20605);
or OR2 (N20609, N20607, N5444);
nor NOR2 (N20610, N20596, N2924);
or OR4 (N20611, N20609, N4997, N13318, N18691);
nand NAND3 (N20612, N20611, N12851, N6586);
and AND3 (N20613, N20597, N9462, N13830);
or OR3 (N20614, N20603, N5709, N2603);
nand NAND2 (N20615, N20613, N12567);
xor XOR2 (N20616, N20593, N13864);
and AND2 (N20617, N20608, N2306);
nor NOR3 (N20618, N20616, N13006, N14747);
buf BUF1 (N20619, N20615);
nor NOR2 (N20620, N20600, N8757);
nor NOR3 (N20621, N20618, N1066, N13948);
not NOT1 (N20622, N20606);
nor NOR4 (N20623, N20612, N15933, N4257, N1497);
nand NAND3 (N20624, N20614, N1473, N1402);
buf BUF1 (N20625, N20610);
xor XOR2 (N20626, N20624, N7297);
nand NAND2 (N20627, N20623, N16881);
not NOT1 (N20628, N20617);
or OR3 (N20629, N20621, N14233, N9540);
nor NOR4 (N20630, N20627, N16542, N14274, N2765);
xor XOR2 (N20631, N20626, N5419);
and AND4 (N20632, N20580, N14285, N9609, N12375);
or OR2 (N20633, N20631, N161);
nor NOR2 (N20634, N20620, N5641);
xor XOR2 (N20635, N20628, N8773);
not NOT1 (N20636, N20634);
and AND2 (N20637, N20625, N12757);
or OR4 (N20638, N20632, N17987, N7268, N12822);
and AND2 (N20639, N20637, N19979);
or OR4 (N20640, N20604, N20364, N11992, N17958);
nor NOR4 (N20641, N20630, N8772, N11878, N9140);
nand NAND2 (N20642, N20622, N14876);
nor NOR2 (N20643, N20639, N2205);
and AND3 (N20644, N20641, N4097, N6500);
nor NOR3 (N20645, N20629, N18026, N14506);
or OR2 (N20646, N20619, N6136);
or OR4 (N20647, N20643, N14204, N7501, N7950);
nor NOR4 (N20648, N20642, N8139, N4077, N7271);
buf BUF1 (N20649, N20635);
or OR2 (N20650, N20647, N13368);
not NOT1 (N20651, N20638);
buf BUF1 (N20652, N20646);
and AND4 (N20653, N20644, N4442, N17707, N532);
nor NOR3 (N20654, N20651, N7335, N14930);
buf BUF1 (N20655, N20636);
nand NAND4 (N20656, N20648, N6858, N16281, N4894);
or OR2 (N20657, N20645, N6406);
or OR3 (N20658, N20655, N1261, N19371);
nand NAND2 (N20659, N20649, N11518);
xor XOR2 (N20660, N20657, N2041);
nand NAND2 (N20661, N20656, N890);
not NOT1 (N20662, N20658);
or OR3 (N20663, N20661, N19704, N7025);
buf BUF1 (N20664, N20640);
buf BUF1 (N20665, N20659);
and AND3 (N20666, N20662, N7322, N3479);
buf BUF1 (N20667, N20654);
xor XOR2 (N20668, N20633, N12814);
not NOT1 (N20669, N20668);
or OR2 (N20670, N20666, N1369);
or OR4 (N20671, N20664, N12299, N6798, N20096);
nand NAND4 (N20672, N20671, N19737, N4400, N426);
and AND3 (N20673, N20669, N468, N13072);
or OR3 (N20674, N20653, N11349, N12585);
nand NAND2 (N20675, N20660, N4415);
xor XOR2 (N20676, N20665, N112);
nand NAND2 (N20677, N20674, N12356);
nor NOR4 (N20678, N20650, N19073, N6027, N12620);
and AND4 (N20679, N20652, N16942, N14110, N14035);
buf BUF1 (N20680, N20677);
nor NOR2 (N20681, N20673, N20317);
not NOT1 (N20682, N20681);
or OR3 (N20683, N20679, N15265, N10436);
or OR2 (N20684, N20678, N11351);
xor XOR2 (N20685, N20683, N14293);
nor NOR2 (N20686, N20670, N17423);
buf BUF1 (N20687, N20682);
or OR2 (N20688, N20686, N19787);
nor NOR3 (N20689, N20672, N3007, N5242);
nor NOR4 (N20690, N20689, N19534, N4241, N1152);
and AND2 (N20691, N20684, N18015);
and AND2 (N20692, N20663, N19416);
buf BUF1 (N20693, N20690);
not NOT1 (N20694, N20688);
xor XOR2 (N20695, N20687, N1632);
xor XOR2 (N20696, N20675, N13726);
and AND4 (N20697, N20692, N2559, N3146, N16144);
xor XOR2 (N20698, N20676, N14189);
or OR4 (N20699, N20697, N7480, N11589, N15374);
or OR2 (N20700, N20680, N6097);
xor XOR2 (N20701, N20667, N220);
and AND2 (N20702, N20693, N1697);
and AND3 (N20703, N20696, N16589, N8864);
or OR3 (N20704, N20695, N11240, N100);
nor NOR2 (N20705, N20704, N19761);
nor NOR2 (N20706, N20700, N20166);
buf BUF1 (N20707, N20691);
nor NOR2 (N20708, N20705, N15314);
not NOT1 (N20709, N20685);
nor NOR3 (N20710, N20703, N10612, N8547);
not NOT1 (N20711, N20698);
and AND2 (N20712, N20709, N15343);
or OR3 (N20713, N20701, N3528, N5682);
nor NOR4 (N20714, N20710, N13605, N12539, N20681);
and AND4 (N20715, N20699, N19549, N10166, N7088);
not NOT1 (N20716, N20711);
buf BUF1 (N20717, N20694);
nand NAND4 (N20718, N20706, N2176, N1427, N14139);
buf BUF1 (N20719, N20708);
not NOT1 (N20720, N20714);
not NOT1 (N20721, N20718);
buf BUF1 (N20722, N20717);
nand NAND4 (N20723, N20702, N13862, N6597, N16116);
nor NOR4 (N20724, N20713, N10565, N9571, N19223);
nand NAND3 (N20725, N20716, N10363, N4415);
buf BUF1 (N20726, N20725);
or OR2 (N20727, N20723, N11214);
xor XOR2 (N20728, N20720, N14814);
buf BUF1 (N20729, N20724);
or OR4 (N20730, N20712, N170, N14056, N4077);
nand NAND4 (N20731, N20715, N9820, N16160, N15587);
not NOT1 (N20732, N20719);
not NOT1 (N20733, N20726);
nand NAND2 (N20734, N20728, N6906);
or OR3 (N20735, N20730, N438, N19456);
or OR4 (N20736, N20729, N13821, N5596, N15828);
not NOT1 (N20737, N20735);
buf BUF1 (N20738, N20722);
xor XOR2 (N20739, N20733, N19315);
nor NOR4 (N20740, N20727, N7306, N8155, N14957);
buf BUF1 (N20741, N20739);
xor XOR2 (N20742, N20740, N11982);
xor XOR2 (N20743, N20738, N8190);
nor NOR4 (N20744, N20737, N14157, N2933, N15496);
nor NOR3 (N20745, N20732, N7815, N17998);
not NOT1 (N20746, N20742);
or OR4 (N20747, N20736, N10778, N6711, N17406);
not NOT1 (N20748, N20746);
not NOT1 (N20749, N20707);
xor XOR2 (N20750, N20748, N14817);
nand NAND2 (N20751, N20745, N17210);
or OR4 (N20752, N20743, N8325, N18061, N9329);
or OR2 (N20753, N20741, N10194);
buf BUF1 (N20754, N20747);
not NOT1 (N20755, N20750);
or OR3 (N20756, N20749, N8853, N17718);
and AND4 (N20757, N20756, N11212, N1064, N7657);
xor XOR2 (N20758, N20751, N19345);
nand NAND4 (N20759, N20757, N7731, N7968, N15401);
nand NAND3 (N20760, N20754, N1299, N11397);
not NOT1 (N20761, N20744);
not NOT1 (N20762, N20755);
or OR2 (N20763, N20753, N4713);
buf BUF1 (N20764, N20721);
buf BUF1 (N20765, N20758);
buf BUF1 (N20766, N20765);
or OR2 (N20767, N20734, N10578);
xor XOR2 (N20768, N20767, N3680);
and AND2 (N20769, N20761, N8290);
and AND3 (N20770, N20763, N11825, N8634);
not NOT1 (N20771, N20769);
or OR4 (N20772, N20764, N7834, N7999, N15201);
nand NAND4 (N20773, N20762, N3152, N10927, N3037);
xor XOR2 (N20774, N20768, N15033);
buf BUF1 (N20775, N20759);
or OR2 (N20776, N20774, N5430);
xor XOR2 (N20777, N20776, N5325);
or OR2 (N20778, N20772, N2858);
buf BUF1 (N20779, N20773);
or OR3 (N20780, N20775, N6327, N6810);
nor NOR3 (N20781, N20777, N3118, N267);
nor NOR3 (N20782, N20752, N37, N17382);
or OR4 (N20783, N20781, N10861, N19569, N3157);
and AND3 (N20784, N20731, N11503, N5653);
buf BUF1 (N20785, N20780);
xor XOR2 (N20786, N20783, N13202);
nor NOR2 (N20787, N20771, N18408);
not NOT1 (N20788, N20787);
not NOT1 (N20789, N20788);
nor NOR4 (N20790, N20789, N9226, N11860, N4830);
nand NAND3 (N20791, N20760, N15535, N17997);
xor XOR2 (N20792, N20779, N18647);
not NOT1 (N20793, N20785);
buf BUF1 (N20794, N20792);
or OR2 (N20795, N20770, N11182);
not NOT1 (N20796, N20782);
nand NAND3 (N20797, N20794, N10070, N3246);
or OR2 (N20798, N20790, N19675);
not NOT1 (N20799, N20796);
nand NAND4 (N20800, N20778, N1931, N2631, N73);
or OR4 (N20801, N20797, N4861, N18694, N10104);
and AND4 (N20802, N20766, N3946, N6253, N8326);
nor NOR2 (N20803, N20784, N10698);
xor XOR2 (N20804, N20793, N1848);
and AND2 (N20805, N20804, N10542);
nand NAND4 (N20806, N20803, N4048, N10720, N10552);
xor XOR2 (N20807, N20802, N2533);
or OR2 (N20808, N20806, N14909);
nand NAND2 (N20809, N20800, N935);
and AND3 (N20810, N20786, N8407, N6347);
not NOT1 (N20811, N20809);
not NOT1 (N20812, N20801);
nor NOR2 (N20813, N20791, N4868);
buf BUF1 (N20814, N20799);
xor XOR2 (N20815, N20805, N5132);
not NOT1 (N20816, N20814);
or OR3 (N20817, N20808, N2965, N1231);
and AND3 (N20818, N20817, N6204, N14395);
nand NAND4 (N20819, N20811, N13794, N9414, N18073);
not NOT1 (N20820, N20795);
not NOT1 (N20821, N20815);
nor NOR3 (N20822, N20816, N3276, N11150);
buf BUF1 (N20823, N20822);
buf BUF1 (N20824, N20798);
buf BUF1 (N20825, N20819);
not NOT1 (N20826, N20823);
nor NOR3 (N20827, N20825, N10953, N14781);
xor XOR2 (N20828, N20818, N16122);
or OR3 (N20829, N20810, N14792, N16106);
not NOT1 (N20830, N20824);
not NOT1 (N20831, N20830);
not NOT1 (N20832, N20812);
and AND4 (N20833, N20807, N1995, N17670, N19148);
nor NOR4 (N20834, N20827, N11759, N4558, N7821);
xor XOR2 (N20835, N20820, N18277);
and AND3 (N20836, N20826, N2203, N20358);
xor XOR2 (N20837, N20828, N6560);
and AND3 (N20838, N20813, N6924, N5732);
xor XOR2 (N20839, N20821, N6687);
xor XOR2 (N20840, N20833, N2584);
buf BUF1 (N20841, N20837);
nor NOR3 (N20842, N20832, N1778, N10503);
or OR3 (N20843, N20842, N3489, N3155);
or OR2 (N20844, N20829, N327);
or OR2 (N20845, N20839, N4028);
buf BUF1 (N20846, N20841);
and AND3 (N20847, N20834, N12586, N18429);
and AND2 (N20848, N20831, N6981);
nor NOR3 (N20849, N20848, N3367, N12275);
buf BUF1 (N20850, N20843);
xor XOR2 (N20851, N20836, N1764);
buf BUF1 (N20852, N20846);
nor NOR2 (N20853, N20850, N2833);
buf BUF1 (N20854, N20838);
or OR4 (N20855, N20852, N14171, N7812, N17443);
buf BUF1 (N20856, N20840);
nand NAND3 (N20857, N20844, N15781, N15102);
not NOT1 (N20858, N20835);
buf BUF1 (N20859, N20855);
or OR4 (N20860, N20847, N10437, N17694, N9531);
or OR3 (N20861, N20860, N11238, N5942);
nor NOR4 (N20862, N20856, N10037, N1781, N18644);
buf BUF1 (N20863, N20845);
not NOT1 (N20864, N20854);
xor XOR2 (N20865, N20849, N3368);
xor XOR2 (N20866, N20859, N16820);
or OR4 (N20867, N20857, N8453, N20777, N8275);
buf BUF1 (N20868, N20864);
nand NAND4 (N20869, N20865, N7424, N16906, N18027);
xor XOR2 (N20870, N20867, N15672);
nor NOR2 (N20871, N20863, N16607);
xor XOR2 (N20872, N20870, N5353);
xor XOR2 (N20873, N20869, N701);
not NOT1 (N20874, N20868);
nand NAND3 (N20875, N20853, N6895, N1597);
and AND4 (N20876, N20861, N9803, N4965, N1960);
and AND2 (N20877, N20851, N2858);
not NOT1 (N20878, N20876);
or OR3 (N20879, N20872, N6002, N11042);
or OR3 (N20880, N20871, N10050, N17920);
xor XOR2 (N20881, N20866, N7682);
nor NOR4 (N20882, N20877, N3658, N5644, N613);
not NOT1 (N20883, N20874);
not NOT1 (N20884, N20858);
or OR2 (N20885, N20880, N15298);
nand NAND2 (N20886, N20878, N15304);
or OR2 (N20887, N20886, N2086);
or OR3 (N20888, N20879, N17391, N16975);
or OR4 (N20889, N20883, N12839, N19550, N5638);
buf BUF1 (N20890, N20885);
or OR4 (N20891, N20884, N530, N13993, N14525);
not NOT1 (N20892, N20881);
xor XOR2 (N20893, N20889, N12339);
and AND2 (N20894, N20875, N4952);
or OR3 (N20895, N20873, N17297, N2844);
nand NAND2 (N20896, N20894, N17818);
or OR3 (N20897, N20892, N17583, N6304);
buf BUF1 (N20898, N20893);
nand NAND3 (N20899, N20898, N14701, N20848);
not NOT1 (N20900, N20899);
or OR4 (N20901, N20896, N4675, N3158, N13939);
not NOT1 (N20902, N20862);
or OR2 (N20903, N20891, N8196);
nor NOR3 (N20904, N20882, N18063, N4742);
and AND2 (N20905, N20897, N11224);
xor XOR2 (N20906, N20888, N1342);
not NOT1 (N20907, N20887);
nand NAND4 (N20908, N20905, N4271, N848, N4641);
nor NOR2 (N20909, N20903, N16075);
and AND4 (N20910, N20901, N7981, N3757, N3304);
nor NOR2 (N20911, N20904, N3190);
xor XOR2 (N20912, N20907, N10311);
or OR4 (N20913, N20902, N4790, N4124, N6039);
or OR2 (N20914, N20900, N18683);
and AND3 (N20915, N20895, N7919, N7240);
nand NAND4 (N20916, N20906, N10743, N3535, N11764);
and AND3 (N20917, N20908, N2124, N13270);
and AND3 (N20918, N20911, N10929, N11431);
nor NOR3 (N20919, N20914, N14676, N17584);
not NOT1 (N20920, N20910);
not NOT1 (N20921, N20917);
nand NAND2 (N20922, N20921, N17797);
nor NOR4 (N20923, N20915, N8882, N17944, N15398);
or OR3 (N20924, N20916, N12910, N9570);
not NOT1 (N20925, N20909);
xor XOR2 (N20926, N20925, N14764);
not NOT1 (N20927, N20919);
or OR2 (N20928, N20890, N2118);
buf BUF1 (N20929, N20924);
xor XOR2 (N20930, N20923, N8044);
nor NOR4 (N20931, N20912, N16532, N9449, N12576);
buf BUF1 (N20932, N20913);
or OR3 (N20933, N20928, N14994, N300);
not NOT1 (N20934, N20933);
and AND2 (N20935, N20929, N18135);
and AND3 (N20936, N20927, N16547, N12671);
buf BUF1 (N20937, N20920);
nand NAND4 (N20938, N20922, N5500, N15019, N8236);
and AND3 (N20939, N20937, N10671, N9470);
not NOT1 (N20940, N20918);
nand NAND2 (N20941, N20934, N15167);
xor XOR2 (N20942, N20940, N20922);
or OR4 (N20943, N20938, N19867, N10695, N12112);
or OR4 (N20944, N20943, N4826, N3561, N8522);
nor NOR4 (N20945, N20932, N3181, N20114, N17590);
nand NAND3 (N20946, N20945, N8468, N12364);
and AND3 (N20947, N20936, N11094, N20119);
not NOT1 (N20948, N20944);
or OR3 (N20949, N20939, N6199, N11282);
nor NOR4 (N20950, N20942, N14448, N10541, N1088);
and AND4 (N20951, N20926, N17649, N11292, N8057);
not NOT1 (N20952, N20946);
not NOT1 (N20953, N20935);
not NOT1 (N20954, N20947);
not NOT1 (N20955, N20953);
nor NOR3 (N20956, N20952, N9080, N6260);
xor XOR2 (N20957, N20950, N4339);
nand NAND3 (N20958, N20948, N14257, N14475);
and AND4 (N20959, N20955, N20242, N558, N12352);
nor NOR3 (N20960, N20959, N17938, N13575);
buf BUF1 (N20961, N20956);
not NOT1 (N20962, N20949);
and AND3 (N20963, N20962, N8605, N4904);
nand NAND3 (N20964, N20930, N5311, N13759);
not NOT1 (N20965, N20954);
buf BUF1 (N20966, N20941);
and AND4 (N20967, N20966, N270, N10049, N5704);
xor XOR2 (N20968, N20961, N4239);
nor NOR3 (N20969, N20967, N20954, N447);
or OR2 (N20970, N20963, N19485);
not NOT1 (N20971, N20969);
buf BUF1 (N20972, N20957);
nand NAND3 (N20973, N20931, N17160, N11680);
buf BUF1 (N20974, N20965);
or OR2 (N20975, N20968, N8753);
xor XOR2 (N20976, N20973, N3700);
nor NOR3 (N20977, N20970, N4018, N6165);
nor NOR2 (N20978, N20964, N6080);
or OR2 (N20979, N20958, N6965);
nand NAND4 (N20980, N20975, N18485, N6366, N19167);
not NOT1 (N20981, N20974);
nor NOR2 (N20982, N20951, N3761);
nor NOR3 (N20983, N20978, N14671, N13086);
and AND4 (N20984, N20983, N20113, N18858, N16471);
xor XOR2 (N20985, N20977, N10009);
or OR4 (N20986, N20971, N10847, N18708, N5903);
or OR3 (N20987, N20986, N6116, N8367);
and AND4 (N20988, N20982, N2075, N14930, N12578);
nor NOR3 (N20989, N20972, N16232, N15075);
nor NOR3 (N20990, N20988, N16439, N20744);
or OR3 (N20991, N20976, N2759, N9044);
or OR3 (N20992, N20960, N629, N18812);
buf BUF1 (N20993, N20984);
nor NOR2 (N20994, N20987, N5229);
buf BUF1 (N20995, N20980);
not NOT1 (N20996, N20989);
not NOT1 (N20997, N20993);
xor XOR2 (N20998, N20996, N3899);
or OR4 (N20999, N20994, N14769, N8658, N16188);
xor XOR2 (N21000, N20981, N2639);
not NOT1 (N21001, N20992);
buf BUF1 (N21002, N20979);
and AND3 (N21003, N21001, N300, N12749);
nand NAND2 (N21004, N20999, N1638);
not NOT1 (N21005, N20998);
or OR3 (N21006, N20991, N7994, N19217);
buf BUF1 (N21007, N20990);
buf BUF1 (N21008, N21003);
nor NOR4 (N21009, N21002, N685, N17728, N17111);
buf BUF1 (N21010, N20985);
not NOT1 (N21011, N20995);
not NOT1 (N21012, N21011);
or OR3 (N21013, N21010, N5902, N4636);
or OR4 (N21014, N21000, N875, N19665, N11930);
nor NOR3 (N21015, N21013, N3226, N10698);
not NOT1 (N21016, N21014);
nand NAND3 (N21017, N21012, N14446, N10177);
nor NOR3 (N21018, N21004, N499, N6591);
not NOT1 (N21019, N21018);
and AND4 (N21020, N21016, N8093, N11051, N10852);
nor NOR3 (N21021, N21017, N6956, N17625);
nor NOR4 (N21022, N21020, N9209, N7291, N10395);
nor NOR3 (N21023, N21022, N14311, N14901);
xor XOR2 (N21024, N21006, N16675);
buf BUF1 (N21025, N21009);
not NOT1 (N21026, N21007);
nor NOR3 (N21027, N20997, N18811, N11444);
nand NAND3 (N21028, N21005, N19298, N712);
nand NAND2 (N21029, N21025, N14621);
nand NAND3 (N21030, N21019, N16231, N4097);
buf BUF1 (N21031, N21027);
nor NOR4 (N21032, N21026, N20068, N15812, N5387);
not NOT1 (N21033, N21028);
buf BUF1 (N21034, N21032);
buf BUF1 (N21035, N21023);
or OR3 (N21036, N21034, N7288, N10472);
or OR2 (N21037, N21030, N5023);
nand NAND4 (N21038, N21033, N20098, N14242, N10894);
buf BUF1 (N21039, N21037);
buf BUF1 (N21040, N21008);
or OR4 (N21041, N21038, N20361, N3839, N10518);
nor NOR3 (N21042, N21024, N6405, N9234);
nand NAND2 (N21043, N21036, N5823);
nand NAND2 (N21044, N21031, N13820);
or OR4 (N21045, N21035, N13665, N15199, N20024);
buf BUF1 (N21046, N21015);
not NOT1 (N21047, N21039);
buf BUF1 (N21048, N21045);
buf BUF1 (N21049, N21040);
or OR3 (N21050, N21041, N2269, N10986);
buf BUF1 (N21051, N21029);
nand NAND3 (N21052, N21050, N19279, N15214);
or OR2 (N21053, N21042, N18232);
and AND3 (N21054, N21049, N17343, N13576);
nand NAND4 (N21055, N21043, N17458, N7636, N5744);
nor NOR4 (N21056, N21053, N5280, N18653, N14313);
xor XOR2 (N21057, N21052, N19228);
nor NOR4 (N21058, N21054, N9722, N12397, N9093);
xor XOR2 (N21059, N21046, N8417);
xor XOR2 (N21060, N21051, N4710);
nor NOR2 (N21061, N21055, N7265);
nand NAND4 (N21062, N21048, N16941, N8609, N12462);
xor XOR2 (N21063, N21061, N20466);
nor NOR3 (N21064, N21062, N16630, N18648);
not NOT1 (N21065, N21057);
buf BUF1 (N21066, N21063);
nand NAND2 (N21067, N21064, N17482);
buf BUF1 (N21068, N21059);
not NOT1 (N21069, N21058);
nand NAND3 (N21070, N21066, N10510, N4971);
or OR3 (N21071, N21060, N17356, N17615);
not NOT1 (N21072, N21065);
and AND4 (N21073, N21067, N2788, N8001, N9174);
xor XOR2 (N21074, N21044, N9111);
nor NOR3 (N21075, N21072, N11832, N1912);
nor NOR4 (N21076, N21071, N2057, N14532, N4632);
and AND3 (N21077, N21073, N2710, N259);
buf BUF1 (N21078, N21069);
not NOT1 (N21079, N21056);
xor XOR2 (N21080, N21077, N141);
not NOT1 (N21081, N21021);
nor NOR3 (N21082, N21075, N18859, N13308);
buf BUF1 (N21083, N21074);
buf BUF1 (N21084, N21079);
buf BUF1 (N21085, N21082);
and AND4 (N21086, N21047, N329, N12862, N6933);
or OR4 (N21087, N21081, N17381, N13634, N16822);
or OR3 (N21088, N21084, N18523, N20145);
and AND3 (N21089, N21083, N5068, N3955);
not NOT1 (N21090, N21080);
buf BUF1 (N21091, N21078);
nor NOR4 (N21092, N21086, N16248, N927, N13576);
and AND2 (N21093, N21087, N2052);
buf BUF1 (N21094, N21093);
nand NAND2 (N21095, N21085, N16171);
and AND3 (N21096, N21092, N10225, N12669);
and AND3 (N21097, N21068, N15078, N113);
xor XOR2 (N21098, N21070, N11528);
buf BUF1 (N21099, N21098);
and AND4 (N21100, N21091, N3167, N14071, N5451);
or OR2 (N21101, N21094, N11514);
or OR2 (N21102, N21101, N9588);
xor XOR2 (N21103, N21096, N14555);
xor XOR2 (N21104, N21100, N9236);
buf BUF1 (N21105, N21102);
not NOT1 (N21106, N21089);
buf BUF1 (N21107, N21103);
nor NOR4 (N21108, N21076, N5851, N13949, N20313);
nor NOR2 (N21109, N21088, N9717);
or OR3 (N21110, N21108, N11610, N15292);
nand NAND2 (N21111, N21099, N14278);
nand NAND2 (N21112, N21090, N9798);
and AND3 (N21113, N21109, N2868, N10695);
and AND4 (N21114, N21106, N13162, N3442, N16512);
buf BUF1 (N21115, N21105);
nor NOR4 (N21116, N21115, N10780, N3524, N11825);
xor XOR2 (N21117, N21097, N15173);
not NOT1 (N21118, N21111);
buf BUF1 (N21119, N21107);
nor NOR2 (N21120, N21118, N12899);
xor XOR2 (N21121, N21095, N454);
or OR2 (N21122, N21119, N4432);
xor XOR2 (N21123, N21117, N2965);
and AND3 (N21124, N21114, N17936, N18669);
not NOT1 (N21125, N21124);
nor NOR3 (N21126, N21123, N18221, N2760);
nor NOR4 (N21127, N21110, N4867, N13240, N15100);
buf BUF1 (N21128, N21113);
buf BUF1 (N21129, N21128);
not NOT1 (N21130, N21126);
not NOT1 (N21131, N21120);
or OR4 (N21132, N21125, N20457, N5182, N14783);
nor NOR4 (N21133, N21127, N773, N6342, N13021);
or OR2 (N21134, N21133, N9616);
nor NOR2 (N21135, N21130, N1077);
not NOT1 (N21136, N21129);
or OR2 (N21137, N21116, N12425);
xor XOR2 (N21138, N21122, N6401);
not NOT1 (N21139, N21135);
not NOT1 (N21140, N21112);
not NOT1 (N21141, N21137);
and AND2 (N21142, N21132, N15741);
not NOT1 (N21143, N21141);
nand NAND3 (N21144, N21140, N16758, N20129);
nor NOR2 (N21145, N21144, N19361);
not NOT1 (N21146, N21134);
nand NAND4 (N21147, N21146, N15699, N1865, N7903);
xor XOR2 (N21148, N21142, N14749);
or OR4 (N21149, N21145, N1640, N5047, N7712);
not NOT1 (N21150, N21136);
nand NAND4 (N21151, N21138, N6629, N10012, N5082);
and AND3 (N21152, N21139, N20624, N5050);
or OR2 (N21153, N21131, N10882);
or OR3 (N21154, N21152, N20011, N9190);
xor XOR2 (N21155, N21148, N13791);
and AND4 (N21156, N21149, N15579, N19833, N2479);
nand NAND2 (N21157, N21104, N13550);
nor NOR3 (N21158, N21150, N11658, N14564);
not NOT1 (N21159, N21158);
xor XOR2 (N21160, N21157, N12679);
nand NAND2 (N21161, N21143, N10322);
buf BUF1 (N21162, N21154);
xor XOR2 (N21163, N21159, N13664);
buf BUF1 (N21164, N21147);
buf BUF1 (N21165, N21155);
buf BUF1 (N21166, N21121);
not NOT1 (N21167, N21161);
or OR4 (N21168, N21160, N6925, N7363, N5699);
buf BUF1 (N21169, N21164);
and AND4 (N21170, N21163, N15736, N13344, N14986);
or OR2 (N21171, N21162, N18919);
nor NOR4 (N21172, N21168, N4084, N19396, N19411);
not NOT1 (N21173, N21153);
nor NOR3 (N21174, N21166, N12001, N416);
or OR2 (N21175, N21167, N15550);
or OR3 (N21176, N21174, N1984, N11675);
nor NOR4 (N21177, N21173, N14353, N5677, N10350);
not NOT1 (N21178, N21170);
buf BUF1 (N21179, N21169);
and AND2 (N21180, N21175, N20835);
or OR4 (N21181, N21178, N1924, N10950, N8652);
and AND4 (N21182, N21179, N20232, N826, N6237);
or OR3 (N21183, N21151, N2291, N11171);
not NOT1 (N21184, N21182);
not NOT1 (N21185, N21177);
buf BUF1 (N21186, N21183);
nand NAND3 (N21187, N21171, N3312, N16741);
nor NOR2 (N21188, N21185, N17905);
nor NOR3 (N21189, N21184, N313, N8136);
xor XOR2 (N21190, N21165, N11030);
or OR2 (N21191, N21181, N14443);
nand NAND2 (N21192, N21190, N12962);
or OR2 (N21193, N21186, N18939);
nand NAND4 (N21194, N21192, N9031, N18946, N16362);
or OR3 (N21195, N21172, N18207, N6321);
not NOT1 (N21196, N21180);
nand NAND4 (N21197, N21195, N16533, N13386, N13131);
not NOT1 (N21198, N21188);
not NOT1 (N21199, N21193);
buf BUF1 (N21200, N21199);
nand NAND2 (N21201, N21187, N6334);
buf BUF1 (N21202, N21191);
buf BUF1 (N21203, N21202);
not NOT1 (N21204, N21201);
xor XOR2 (N21205, N21196, N11644);
not NOT1 (N21206, N21204);
and AND2 (N21207, N21189, N7115);
not NOT1 (N21208, N21205);
not NOT1 (N21209, N21156);
nor NOR2 (N21210, N21208, N15848);
xor XOR2 (N21211, N21198, N6506);
xor XOR2 (N21212, N21210, N13140);
not NOT1 (N21213, N21197);
xor XOR2 (N21214, N21203, N17215);
nor NOR4 (N21215, N21212, N6933, N18759, N12328);
or OR2 (N21216, N21206, N10665);
and AND2 (N21217, N21215, N13229);
nor NOR4 (N21218, N21213, N5723, N3896, N15357);
nor NOR2 (N21219, N21216, N16991);
nor NOR2 (N21220, N21176, N20287);
not NOT1 (N21221, N21200);
or OR3 (N21222, N21194, N7346, N16077);
or OR3 (N21223, N21220, N15492, N1748);
and AND2 (N21224, N21207, N8077);
or OR4 (N21225, N21219, N19738, N4211, N9420);
nor NOR4 (N21226, N21221, N4793, N5785, N2175);
or OR2 (N21227, N21211, N19378);
or OR3 (N21228, N21218, N21049, N20515);
not NOT1 (N21229, N21222);
nor NOR3 (N21230, N21224, N14810, N880);
and AND4 (N21231, N21227, N8793, N2856, N17398);
and AND3 (N21232, N21230, N7277, N13432);
nand NAND4 (N21233, N21229, N9145, N4140, N4818);
or OR2 (N21234, N21214, N12730);
nor NOR2 (N21235, N21209, N18551);
xor XOR2 (N21236, N21225, N10737);
not NOT1 (N21237, N21234);
nor NOR4 (N21238, N21217, N13881, N2935, N6534);
xor XOR2 (N21239, N21238, N13226);
xor XOR2 (N21240, N21237, N20743);
xor XOR2 (N21241, N21236, N15850);
xor XOR2 (N21242, N21231, N9262);
buf BUF1 (N21243, N21232);
and AND2 (N21244, N21233, N12075);
xor XOR2 (N21245, N21223, N9688);
not NOT1 (N21246, N21235);
xor XOR2 (N21247, N21246, N13167);
xor XOR2 (N21248, N21245, N12042);
nor NOR2 (N21249, N21241, N9815);
or OR2 (N21250, N21226, N12146);
or OR4 (N21251, N21228, N3243, N4939, N7771);
nor NOR2 (N21252, N21243, N19699);
not NOT1 (N21253, N21252);
nand NAND4 (N21254, N21239, N14049, N12131, N20617);
nand NAND3 (N21255, N21253, N7244, N18071);
buf BUF1 (N21256, N21248);
and AND3 (N21257, N21251, N16656, N4588);
xor XOR2 (N21258, N21256, N15522);
xor XOR2 (N21259, N21250, N11182);
xor XOR2 (N21260, N21254, N13599);
nand NAND3 (N21261, N21247, N6781, N2012);
not NOT1 (N21262, N21255);
buf BUF1 (N21263, N21249);
nor NOR4 (N21264, N21261, N13987, N19496, N620);
or OR3 (N21265, N21259, N9958, N13566);
not NOT1 (N21266, N21264);
nor NOR3 (N21267, N21265, N2732, N6043);
buf BUF1 (N21268, N21244);
nor NOR2 (N21269, N21257, N7241);
nand NAND2 (N21270, N21263, N20737);
xor XOR2 (N21271, N21267, N957);
or OR3 (N21272, N21269, N16808, N3585);
xor XOR2 (N21273, N21262, N9853);
buf BUF1 (N21274, N21266);
nor NOR3 (N21275, N21268, N10385, N8760);
not NOT1 (N21276, N21258);
nand NAND4 (N21277, N21273, N12244, N5467, N8842);
not NOT1 (N21278, N21260);
or OR4 (N21279, N21276, N14999, N7568, N17225);
buf BUF1 (N21280, N21274);
not NOT1 (N21281, N21278);
xor XOR2 (N21282, N21279, N1780);
nor NOR2 (N21283, N21282, N16063);
nor NOR4 (N21284, N21283, N8126, N2833, N18147);
and AND4 (N21285, N21280, N1389, N3445, N18013);
and AND2 (N21286, N21281, N2507);
and AND4 (N21287, N21271, N3086, N14281, N14383);
not NOT1 (N21288, N21286);
xor XOR2 (N21289, N21272, N16972);
buf BUF1 (N21290, N21277);
nand NAND3 (N21291, N21284, N5078, N10521);
nor NOR4 (N21292, N21287, N181, N17692, N8376);
or OR2 (N21293, N21242, N6454);
nor NOR3 (N21294, N21285, N20591, N18441);
buf BUF1 (N21295, N21275);
buf BUF1 (N21296, N21288);
buf BUF1 (N21297, N21294);
buf BUF1 (N21298, N21293);
and AND2 (N21299, N21240, N7623);
xor XOR2 (N21300, N21297, N2821);
or OR2 (N21301, N21291, N10774);
or OR4 (N21302, N21270, N2304, N10873, N3011);
and AND2 (N21303, N21289, N11509);
nor NOR4 (N21304, N21303, N18277, N9566, N6027);
or OR4 (N21305, N21296, N6803, N2883, N19270);
or OR3 (N21306, N21298, N16483, N2025);
not NOT1 (N21307, N21299);
nor NOR3 (N21308, N21301, N1452, N15953);
or OR4 (N21309, N21305, N13052, N15565, N20073);
nor NOR2 (N21310, N21302, N20364);
nand NAND2 (N21311, N21308, N15177);
buf BUF1 (N21312, N21311);
xor XOR2 (N21313, N21295, N16111);
buf BUF1 (N21314, N21300);
nand NAND4 (N21315, N21306, N2272, N21256, N18318);
or OR3 (N21316, N21313, N18669, N9507);
nand NAND3 (N21317, N21315, N12377, N8753);
nand NAND2 (N21318, N21310, N11145);
nor NOR4 (N21319, N21316, N9917, N14483, N2177);
xor XOR2 (N21320, N21304, N18200);
nor NOR3 (N21321, N21314, N17130, N21113);
xor XOR2 (N21322, N21312, N18124);
or OR2 (N21323, N21318, N18381);
nand NAND3 (N21324, N21317, N8303, N9863);
nand NAND4 (N21325, N21290, N8548, N16483, N4137);
or OR4 (N21326, N21324, N20081, N5752, N2677);
not NOT1 (N21327, N21309);
buf BUF1 (N21328, N21326);
nor NOR4 (N21329, N21320, N6739, N12686, N7418);
xor XOR2 (N21330, N21323, N16276);
nor NOR4 (N21331, N21325, N19197, N1987, N5989);
or OR3 (N21332, N21322, N6992, N483);
buf BUF1 (N21333, N21319);
xor XOR2 (N21334, N21330, N10111);
buf BUF1 (N21335, N21332);
nor NOR4 (N21336, N21333, N4211, N15457, N8192);
xor XOR2 (N21337, N21307, N1709);
nand NAND2 (N21338, N21331, N13709);
or OR4 (N21339, N21338, N2936, N5647, N16233);
or OR3 (N21340, N21336, N9828, N6460);
xor XOR2 (N21341, N21321, N214);
xor XOR2 (N21342, N21329, N13665);
nor NOR3 (N21343, N21342, N18412, N4109);
buf BUF1 (N21344, N21335);
buf BUF1 (N21345, N21328);
nand NAND2 (N21346, N21343, N8496);
buf BUF1 (N21347, N21337);
and AND2 (N21348, N21346, N12249);
or OR3 (N21349, N21340, N13940, N7874);
xor XOR2 (N21350, N21339, N15404);
buf BUF1 (N21351, N21349);
not NOT1 (N21352, N21292);
nor NOR2 (N21353, N21352, N14364);
and AND3 (N21354, N21334, N755, N11300);
buf BUF1 (N21355, N21341);
or OR3 (N21356, N21354, N2789, N6418);
and AND3 (N21357, N21344, N17392, N12652);
not NOT1 (N21358, N21351);
nand NAND2 (N21359, N21327, N807);
and AND2 (N21360, N21350, N762);
not NOT1 (N21361, N21355);
or OR4 (N21362, N21353, N12156, N17387, N10759);
buf BUF1 (N21363, N21345);
buf BUF1 (N21364, N21348);
or OR2 (N21365, N21359, N4375);
nand NAND4 (N21366, N21357, N10928, N13403, N12016);
nand NAND4 (N21367, N21364, N12501, N17349, N19183);
or OR2 (N21368, N21360, N419);
nor NOR4 (N21369, N21356, N14375, N500, N19267);
nand NAND2 (N21370, N21366, N11069);
nand NAND3 (N21371, N21365, N9643, N318);
nand NAND3 (N21372, N21347, N1636, N11351);
buf BUF1 (N21373, N21362);
xor XOR2 (N21374, N21373, N10130);
or OR3 (N21375, N21369, N18456, N3307);
not NOT1 (N21376, N21361);
not NOT1 (N21377, N21370);
nand NAND3 (N21378, N21376, N5954, N17596);
buf BUF1 (N21379, N21377);
nor NOR3 (N21380, N21378, N18224, N9024);
or OR2 (N21381, N21358, N15594);
or OR3 (N21382, N21379, N10578, N12823);
or OR3 (N21383, N21371, N165, N4406);
nor NOR2 (N21384, N21374, N18891);
nor NOR2 (N21385, N21384, N9971);
nand NAND2 (N21386, N21375, N5375);
not NOT1 (N21387, N21383);
not NOT1 (N21388, N21363);
and AND2 (N21389, N21381, N6370);
nor NOR3 (N21390, N21385, N4515, N11245);
nand NAND4 (N21391, N21390, N15349, N20253, N7092);
nor NOR3 (N21392, N21380, N7459, N11375);
buf BUF1 (N21393, N21372);
nor NOR4 (N21394, N21368, N436, N10847, N12002);
buf BUF1 (N21395, N21388);
and AND2 (N21396, N21393, N9191);
and AND3 (N21397, N21396, N3681, N10107);
nor NOR4 (N21398, N21395, N17553, N8475, N19496);
xor XOR2 (N21399, N21367, N15791);
not NOT1 (N21400, N21387);
and AND3 (N21401, N21382, N344, N11406);
or OR4 (N21402, N21391, N1195, N13972, N16187);
buf BUF1 (N21403, N21397);
and AND4 (N21404, N21399, N12069, N13451, N13528);
nand NAND2 (N21405, N21401, N4379);
buf BUF1 (N21406, N21394);
or OR2 (N21407, N21403, N15692);
nand NAND4 (N21408, N21386, N10917, N20977, N20860);
not NOT1 (N21409, N21405);
buf BUF1 (N21410, N21400);
not NOT1 (N21411, N21409);
xor XOR2 (N21412, N21398, N2703);
nand NAND2 (N21413, N21402, N13156);
not NOT1 (N21414, N21404);
not NOT1 (N21415, N21413);
and AND2 (N21416, N21406, N11648);
buf BUF1 (N21417, N21410);
nor NOR3 (N21418, N21416, N15363, N17343);
buf BUF1 (N21419, N21407);
not NOT1 (N21420, N21418);
and AND2 (N21421, N21419, N14199);
nor NOR2 (N21422, N21408, N17646);
or OR3 (N21423, N21414, N12785, N4555);
not NOT1 (N21424, N21412);
nand NAND3 (N21425, N21415, N11693, N19537);
nand NAND4 (N21426, N21389, N19404, N9453, N754);
and AND3 (N21427, N21420, N17767, N7537);
xor XOR2 (N21428, N21422, N14920);
nand NAND2 (N21429, N21421, N17046);
or OR2 (N21430, N21417, N18731);
xor XOR2 (N21431, N21424, N154);
nand NAND2 (N21432, N21431, N10943);
or OR3 (N21433, N21425, N3200, N3317);
nand NAND2 (N21434, N21429, N13237);
xor XOR2 (N21435, N21411, N14316);
buf BUF1 (N21436, N21423);
and AND3 (N21437, N21434, N17456, N20216);
and AND2 (N21438, N21392, N10428);
nand NAND4 (N21439, N21433, N181, N18845, N10569);
and AND2 (N21440, N21427, N18745);
nand NAND2 (N21441, N21428, N8155);
nor NOR4 (N21442, N21440, N15628, N2125, N13584);
not NOT1 (N21443, N21439);
nand NAND2 (N21444, N21442, N12688);
nor NOR3 (N21445, N21444, N6704, N5037);
nand NAND2 (N21446, N21441, N15371);
not NOT1 (N21447, N21435);
xor XOR2 (N21448, N21443, N1990);
xor XOR2 (N21449, N21438, N9880);
not NOT1 (N21450, N21449);
and AND2 (N21451, N21445, N17309);
buf BUF1 (N21452, N21436);
nand NAND2 (N21453, N21451, N15234);
xor XOR2 (N21454, N21432, N16670);
and AND3 (N21455, N21450, N1394, N6759);
and AND4 (N21456, N21454, N4888, N2759, N14052);
nand NAND2 (N21457, N21447, N21438);
nand NAND2 (N21458, N21452, N16768);
and AND3 (N21459, N21458, N4129, N12336);
xor XOR2 (N21460, N21437, N14878);
not NOT1 (N21461, N21459);
nor NOR4 (N21462, N21426, N13032, N13207, N14623);
xor XOR2 (N21463, N21461, N15604);
buf BUF1 (N21464, N21463);
nor NOR2 (N21465, N21464, N18349);
nor NOR4 (N21466, N21448, N13114, N11722, N12916);
not NOT1 (N21467, N21446);
xor XOR2 (N21468, N21467, N4182);
nand NAND3 (N21469, N21462, N15620, N2544);
or OR4 (N21470, N21465, N1648, N182, N5669);
nand NAND4 (N21471, N21468, N6815, N3725, N12266);
nor NOR2 (N21472, N21455, N16455);
nor NOR4 (N21473, N21457, N20514, N3463, N10578);
xor XOR2 (N21474, N21456, N7953);
nand NAND3 (N21475, N21473, N12873, N3432);
nand NAND2 (N21476, N21466, N5942);
xor XOR2 (N21477, N21476, N6081);
buf BUF1 (N21478, N21430);
and AND2 (N21479, N21469, N17830);
nor NOR3 (N21480, N21460, N1539, N15134);
and AND4 (N21481, N21472, N16238, N14940, N12110);
not NOT1 (N21482, N21475);
xor XOR2 (N21483, N21453, N9320);
or OR2 (N21484, N21483, N585);
or OR2 (N21485, N21479, N16144);
or OR4 (N21486, N21478, N13414, N8520, N20325);
nor NOR3 (N21487, N21470, N7490, N7963);
not NOT1 (N21488, N21480);
or OR2 (N21489, N21485, N2004);
nor NOR2 (N21490, N21482, N15364);
and AND4 (N21491, N21487, N15151, N14162, N18534);
or OR2 (N21492, N21486, N18242);
or OR4 (N21493, N21490, N13250, N112, N17191);
nand NAND4 (N21494, N21489, N17525, N4862, N10168);
not NOT1 (N21495, N21493);
buf BUF1 (N21496, N21494);
nor NOR4 (N21497, N21484, N20665, N2496, N13590);
and AND3 (N21498, N21497, N13270, N20720);
nand NAND3 (N21499, N21491, N9599, N15120);
nand NAND3 (N21500, N21492, N2945, N11473);
not NOT1 (N21501, N21481);
not NOT1 (N21502, N21488);
nand NAND3 (N21503, N21502, N16169, N8475);
nand NAND4 (N21504, N21503, N21105, N11332, N16141);
buf BUF1 (N21505, N21504);
not NOT1 (N21506, N21471);
buf BUF1 (N21507, N21500);
nor NOR2 (N21508, N21498, N20507);
xor XOR2 (N21509, N21505, N9300);
xor XOR2 (N21510, N21477, N17704);
nand NAND2 (N21511, N21510, N14007);
xor XOR2 (N21512, N21507, N15535);
or OR3 (N21513, N21495, N15291, N17794);
or OR3 (N21514, N21511, N13137, N7065);
nand NAND4 (N21515, N21514, N20600, N19838, N8502);
not NOT1 (N21516, N21515);
nand NAND2 (N21517, N21506, N2836);
buf BUF1 (N21518, N21496);
nor NOR2 (N21519, N21518, N17696);
and AND4 (N21520, N21499, N3473, N11396, N12708);
and AND2 (N21521, N21512, N6349);
not NOT1 (N21522, N21517);
buf BUF1 (N21523, N21474);
nand NAND2 (N21524, N21516, N14043);
buf BUF1 (N21525, N21508);
nor NOR4 (N21526, N21522, N5397, N10961, N19410);
xor XOR2 (N21527, N21523, N1941);
not NOT1 (N21528, N21509);
or OR2 (N21529, N21526, N15296);
and AND4 (N21530, N21528, N742, N1657, N762);
or OR2 (N21531, N21521, N7075);
xor XOR2 (N21532, N21519, N8331);
nor NOR3 (N21533, N21531, N11403, N15400);
and AND4 (N21534, N21525, N17394, N3362, N12779);
buf BUF1 (N21535, N21527);
and AND2 (N21536, N21534, N16485);
not NOT1 (N21537, N21532);
and AND2 (N21538, N21535, N21162);
not NOT1 (N21539, N21513);
or OR4 (N21540, N21533, N11723, N3757, N3709);
buf BUF1 (N21541, N21530);
and AND4 (N21542, N21501, N8268, N14103, N20235);
xor XOR2 (N21543, N21539, N15898);
xor XOR2 (N21544, N21520, N8647);
nand NAND4 (N21545, N21537, N15181, N15225, N16962);
buf BUF1 (N21546, N21538);
nand NAND3 (N21547, N21529, N4354, N10824);
nand NAND2 (N21548, N21546, N1764);
and AND4 (N21549, N21541, N15737, N7072, N14307);
or OR2 (N21550, N21543, N18747);
and AND3 (N21551, N21547, N8870, N20451);
nand NAND3 (N21552, N21548, N20914, N15251);
not NOT1 (N21553, N21524);
not NOT1 (N21554, N21549);
or OR3 (N21555, N21542, N5843, N6944);
or OR4 (N21556, N21545, N4051, N478, N17662);
or OR2 (N21557, N21556, N2538);
and AND4 (N21558, N21554, N9313, N21297, N3419);
nand NAND2 (N21559, N21555, N17531);
and AND2 (N21560, N21551, N4923);
nor NOR4 (N21561, N21536, N10636, N8425, N12387);
and AND3 (N21562, N21561, N11188, N14057);
and AND4 (N21563, N21562, N2105, N17638, N16154);
and AND3 (N21564, N21544, N17128, N17433);
and AND3 (N21565, N21550, N7184, N6541);
or OR2 (N21566, N21564, N607);
and AND4 (N21567, N21559, N5706, N17725, N16719);
or OR4 (N21568, N21553, N11569, N452, N5753);
or OR2 (N21569, N21558, N6052);
buf BUF1 (N21570, N21557);
or OR2 (N21571, N21567, N7824);
nor NOR4 (N21572, N21540, N18763, N9523, N58);
xor XOR2 (N21573, N21552, N10074);
or OR4 (N21574, N21573, N9468, N21251, N15099);
or OR3 (N21575, N21571, N13343, N20703);
buf BUF1 (N21576, N21569);
buf BUF1 (N21577, N21576);
and AND4 (N21578, N21570, N19726, N2075, N4830);
nor NOR2 (N21579, N21574, N3856);
not NOT1 (N21580, N21565);
not NOT1 (N21581, N21578);
xor XOR2 (N21582, N21575, N7687);
buf BUF1 (N21583, N21563);
nor NOR3 (N21584, N21560, N19205, N6712);
buf BUF1 (N21585, N21572);
buf BUF1 (N21586, N21584);
or OR3 (N21587, N21581, N21179, N19204);
or OR3 (N21588, N21586, N16318, N2575);
nor NOR2 (N21589, N21580, N20405);
or OR2 (N21590, N21589, N1847);
buf BUF1 (N21591, N21587);
xor XOR2 (N21592, N21582, N2912);
nand NAND3 (N21593, N21592, N12273, N13567);
nand NAND2 (N21594, N21579, N15837);
not NOT1 (N21595, N21577);
and AND2 (N21596, N21591, N4820);
and AND4 (N21597, N21596, N11259, N16, N15761);
and AND2 (N21598, N21568, N21142);
buf BUF1 (N21599, N21593);
nand NAND3 (N21600, N21594, N11463, N19021);
buf BUF1 (N21601, N21595);
nor NOR4 (N21602, N21566, N12699, N2934, N17805);
buf BUF1 (N21603, N21599);
buf BUF1 (N21604, N21603);
xor XOR2 (N21605, N21583, N794);
and AND2 (N21606, N21590, N18152);
nor NOR4 (N21607, N21598, N3775, N21162, N10541);
buf BUF1 (N21608, N21600);
xor XOR2 (N21609, N21602, N18799);
not NOT1 (N21610, N21607);
buf BUF1 (N21611, N21605);
xor XOR2 (N21612, N21606, N21071);
buf BUF1 (N21613, N21597);
nand NAND4 (N21614, N21601, N19319, N7786, N11842);
not NOT1 (N21615, N21612);
and AND4 (N21616, N21610, N21467, N6941, N16440);
buf BUF1 (N21617, N21609);
or OR3 (N21618, N21614, N16445, N20758);
and AND3 (N21619, N21616, N8807, N13574);
and AND3 (N21620, N21617, N3465, N7449);
xor XOR2 (N21621, N21585, N7827);
xor XOR2 (N21622, N21588, N3490);
and AND2 (N21623, N21611, N4975);
or OR3 (N21624, N21613, N21252, N20124);
not NOT1 (N21625, N21604);
xor XOR2 (N21626, N21624, N18769);
xor XOR2 (N21627, N21625, N13231);
or OR4 (N21628, N21618, N4766, N6026, N1859);
buf BUF1 (N21629, N21619);
or OR3 (N21630, N21615, N8585, N16778);
and AND3 (N21631, N21628, N5234, N18787);
nor NOR2 (N21632, N21608, N15516);
or OR3 (N21633, N21622, N14647, N16987);
xor XOR2 (N21634, N21630, N14693);
nor NOR3 (N21635, N21631, N13549, N16686);
nor NOR2 (N21636, N21620, N14759);
buf BUF1 (N21637, N21629);
not NOT1 (N21638, N21627);
or OR3 (N21639, N21636, N7861, N19438);
nor NOR2 (N21640, N21621, N1194);
nand NAND4 (N21641, N21639, N21344, N20415, N15901);
or OR2 (N21642, N21635, N21257);
buf BUF1 (N21643, N21632);
buf BUF1 (N21644, N21633);
and AND4 (N21645, N21641, N7380, N7892, N2145);
and AND3 (N21646, N21637, N12562, N18347);
not NOT1 (N21647, N21634);
buf BUF1 (N21648, N21642);
buf BUF1 (N21649, N21644);
and AND4 (N21650, N21648, N296, N10319, N17183);
buf BUF1 (N21651, N21650);
xor XOR2 (N21652, N21651, N14299);
buf BUF1 (N21653, N21626);
not NOT1 (N21654, N21623);
nand NAND2 (N21655, N21649, N14177);
nor NOR4 (N21656, N21653, N18948, N12975, N3962);
nand NAND3 (N21657, N21656, N16779, N15887);
or OR2 (N21658, N21638, N8056);
buf BUF1 (N21659, N21646);
and AND2 (N21660, N21647, N3849);
xor XOR2 (N21661, N21658, N1717);
and AND4 (N21662, N21645, N15986, N4441, N9742);
or OR2 (N21663, N21662, N17530);
nor NOR4 (N21664, N21660, N6014, N20930, N5835);
and AND2 (N21665, N21663, N1682);
xor XOR2 (N21666, N21654, N286);
or OR2 (N21667, N21664, N13497);
buf BUF1 (N21668, N21666);
xor XOR2 (N21669, N21659, N20966);
nor NOR2 (N21670, N21661, N2328);
buf BUF1 (N21671, N21665);
and AND2 (N21672, N21657, N8584);
nor NOR4 (N21673, N21672, N8203, N1892, N662);
nand NAND2 (N21674, N21652, N11742);
xor XOR2 (N21675, N21670, N9752);
not NOT1 (N21676, N21673);
xor XOR2 (N21677, N21668, N20974);
not NOT1 (N21678, N21667);
and AND2 (N21679, N21674, N5224);
not NOT1 (N21680, N21677);
buf BUF1 (N21681, N21679);
nand NAND4 (N21682, N21671, N752, N7848, N20219);
nand NAND4 (N21683, N21675, N18249, N817, N4695);
buf BUF1 (N21684, N21683);
nor NOR4 (N21685, N21643, N975, N3739, N13411);
nand NAND3 (N21686, N21685, N15542, N9316);
xor XOR2 (N21687, N21682, N13336);
buf BUF1 (N21688, N21676);
or OR4 (N21689, N21684, N5108, N18601, N11984);
not NOT1 (N21690, N21688);
buf BUF1 (N21691, N21680);
nand NAND4 (N21692, N21655, N16668, N20903, N15931);
nor NOR2 (N21693, N21678, N3285);
or OR2 (N21694, N21692, N2821);
buf BUF1 (N21695, N21687);
buf BUF1 (N21696, N21669);
not NOT1 (N21697, N21686);
and AND4 (N21698, N21681, N16331, N19256, N11424);
and AND2 (N21699, N21696, N9586);
not NOT1 (N21700, N21699);
or OR3 (N21701, N21694, N1933, N13711);
or OR2 (N21702, N21701, N11346);
not NOT1 (N21703, N21693);
xor XOR2 (N21704, N21695, N13912);
xor XOR2 (N21705, N21690, N7064);
and AND2 (N21706, N21702, N14057);
xor XOR2 (N21707, N21704, N4844);
or OR2 (N21708, N21689, N15435);
buf BUF1 (N21709, N21691);
buf BUF1 (N21710, N21698);
not NOT1 (N21711, N21707);
and AND3 (N21712, N21711, N17290, N5702);
xor XOR2 (N21713, N21708, N7619);
or OR4 (N21714, N21710, N213, N7784, N9099);
and AND2 (N21715, N21700, N10717);
not NOT1 (N21716, N21640);
buf BUF1 (N21717, N21703);
nand NAND4 (N21718, N21713, N7144, N17575, N15012);
nor NOR3 (N21719, N21718, N4758, N13056);
and AND2 (N21720, N21712, N13019);
nor NOR4 (N21721, N21719, N10199, N869, N436);
and AND4 (N21722, N21720, N87, N16226, N21182);
buf BUF1 (N21723, N21697);
nand NAND2 (N21724, N21706, N4041);
not NOT1 (N21725, N21721);
nor NOR4 (N21726, N21716, N17246, N12020, N3726);
nor NOR3 (N21727, N21725, N10709, N9047);
not NOT1 (N21728, N21714);
nand NAND4 (N21729, N21728, N11775, N15264, N17558);
xor XOR2 (N21730, N21709, N16747);
or OR3 (N21731, N21729, N9317, N563);
nand NAND2 (N21732, N21730, N535);
nor NOR3 (N21733, N21732, N7919, N9475);
xor XOR2 (N21734, N21733, N4412);
buf BUF1 (N21735, N21715);
buf BUF1 (N21736, N21735);
not NOT1 (N21737, N21705);
not NOT1 (N21738, N21734);
nand NAND2 (N21739, N21723, N5441);
buf BUF1 (N21740, N21739);
xor XOR2 (N21741, N21724, N15570);
and AND2 (N21742, N21717, N9127);
nor NOR2 (N21743, N21737, N19635);
buf BUF1 (N21744, N21742);
nor NOR2 (N21745, N21722, N19454);
not NOT1 (N21746, N21744);
and AND3 (N21747, N21726, N517, N10501);
xor XOR2 (N21748, N21741, N2735);
xor XOR2 (N21749, N21748, N5592);
or OR4 (N21750, N21736, N14225, N18563, N10394);
and AND3 (N21751, N21749, N20837, N16602);
nand NAND3 (N21752, N21750, N5487, N6832);
not NOT1 (N21753, N21745);
nand NAND4 (N21754, N21753, N3744, N10649, N3652);
xor XOR2 (N21755, N21727, N10311);
not NOT1 (N21756, N21738);
xor XOR2 (N21757, N21751, N20084);
xor XOR2 (N21758, N21752, N18168);
and AND4 (N21759, N21731, N4737, N503, N1001);
buf BUF1 (N21760, N21755);
or OR4 (N21761, N21746, N15836, N8612, N13408);
and AND3 (N21762, N21759, N9611, N7836);
nor NOR4 (N21763, N21757, N17970, N5880, N12223);
and AND2 (N21764, N21756, N12976);
or OR3 (N21765, N21762, N13828, N1033);
and AND2 (N21766, N21760, N18017);
and AND2 (N21767, N21743, N13508);
buf BUF1 (N21768, N21747);
nand NAND3 (N21769, N21767, N9001, N11827);
nand NAND4 (N21770, N21769, N5746, N1840, N5341);
nand NAND4 (N21771, N21763, N9475, N20319, N2624);
not NOT1 (N21772, N21768);
nor NOR2 (N21773, N21770, N6300);
xor XOR2 (N21774, N21772, N9544);
or OR2 (N21775, N21765, N3584);
buf BUF1 (N21776, N21764);
or OR4 (N21777, N21771, N13128, N10538, N4294);
or OR4 (N21778, N21761, N7478, N18119, N10935);
xor XOR2 (N21779, N21776, N3236);
xor XOR2 (N21780, N21775, N3178);
xor XOR2 (N21781, N21740, N10101);
and AND2 (N21782, N21781, N3548);
and AND4 (N21783, N21778, N1005, N19933, N7624);
nand NAND2 (N21784, N21754, N2485);
not NOT1 (N21785, N21766);
and AND3 (N21786, N21780, N1910, N20003);
buf BUF1 (N21787, N21784);
nand NAND2 (N21788, N21782, N3187);
or OR4 (N21789, N21758, N5880, N19420, N2181);
buf BUF1 (N21790, N21787);
buf BUF1 (N21791, N21779);
or OR4 (N21792, N21789, N10650, N4531, N11436);
and AND3 (N21793, N21791, N21257, N21257);
or OR2 (N21794, N21773, N18400);
not NOT1 (N21795, N21788);
or OR2 (N21796, N21774, N716);
or OR4 (N21797, N21794, N3466, N7697, N7019);
not NOT1 (N21798, N21790);
not NOT1 (N21799, N21798);
nand NAND2 (N21800, N21785, N8669);
buf BUF1 (N21801, N21796);
nor NOR3 (N21802, N21792, N1545, N4018);
buf BUF1 (N21803, N21800);
nor NOR3 (N21804, N21801, N10557, N66);
not NOT1 (N21805, N21777);
nand NAND3 (N21806, N21803, N11969, N18120);
or OR4 (N21807, N21786, N14507, N11967, N12956);
nand NAND2 (N21808, N21807, N7469);
xor XOR2 (N21809, N21805, N19421);
buf BUF1 (N21810, N21795);
xor XOR2 (N21811, N21802, N11058);
and AND3 (N21812, N21793, N403, N10446);
not NOT1 (N21813, N21808);
xor XOR2 (N21814, N21783, N12373);
nor NOR4 (N21815, N21804, N1532, N2329, N3595);
nand NAND3 (N21816, N21810, N16595, N20366);
nor NOR2 (N21817, N21815, N6895);
nand NAND2 (N21818, N21813, N7222);
buf BUF1 (N21819, N21818);
buf BUF1 (N21820, N21799);
buf BUF1 (N21821, N21812);
buf BUF1 (N21822, N21814);
and AND4 (N21823, N21819, N10857, N12939, N264);
nor NOR2 (N21824, N21806, N12250);
buf BUF1 (N21825, N21797);
buf BUF1 (N21826, N21824);
nor NOR4 (N21827, N21823, N4209, N21171, N9172);
xor XOR2 (N21828, N21825, N2865);
not NOT1 (N21829, N21827);
not NOT1 (N21830, N21829);
nand NAND4 (N21831, N21817, N12075, N12735, N17900);
not NOT1 (N21832, N21826);
or OR4 (N21833, N21828, N4565, N879, N3940);
buf BUF1 (N21834, N21832);
xor XOR2 (N21835, N21830, N3157);
nand NAND4 (N21836, N21831, N3146, N10182, N16130);
not NOT1 (N21837, N21833);
not NOT1 (N21838, N21835);
or OR2 (N21839, N21836, N5245);
nor NOR2 (N21840, N21821, N9713);
nand NAND3 (N21841, N21837, N13082, N9005);
not NOT1 (N21842, N21841);
or OR2 (N21843, N21842, N21336);
xor XOR2 (N21844, N21816, N15619);
buf BUF1 (N21845, N21839);
nor NOR3 (N21846, N21811, N8454, N10575);
nor NOR4 (N21847, N21844, N1785, N3362, N10349);
buf BUF1 (N21848, N21834);
xor XOR2 (N21849, N21847, N11862);
buf BUF1 (N21850, N21845);
xor XOR2 (N21851, N21820, N10682);
nor NOR2 (N21852, N21822, N21734);
nor NOR4 (N21853, N21846, N17320, N623, N6584);
nor NOR2 (N21854, N21853, N21799);
nor NOR4 (N21855, N21851, N2859, N5266, N10070);
buf BUF1 (N21856, N21840);
or OR4 (N21857, N21850, N21567, N3879, N20761);
xor XOR2 (N21858, N21843, N11580);
and AND3 (N21859, N21858, N16716, N20207);
buf BUF1 (N21860, N21855);
and AND2 (N21861, N21849, N17812);
and AND2 (N21862, N21859, N6663);
nor NOR4 (N21863, N21860, N4878, N13025, N17323);
not NOT1 (N21864, N21861);
nor NOR3 (N21865, N21864, N5810, N10436);
xor XOR2 (N21866, N21865, N1618);
or OR2 (N21867, N21857, N20971);
nor NOR4 (N21868, N21854, N14062, N16950, N14895);
nand NAND3 (N21869, N21838, N3940, N2244);
and AND4 (N21870, N21863, N11349, N14049, N16068);
xor XOR2 (N21871, N21868, N16048);
xor XOR2 (N21872, N21866, N19020);
xor XOR2 (N21873, N21809, N20565);
or OR4 (N21874, N21871, N19384, N1119, N17456);
and AND4 (N21875, N21872, N10065, N13720, N17571);
nand NAND4 (N21876, N21870, N2121, N19760, N8218);
or OR4 (N21877, N21856, N1609, N14392, N3977);
nand NAND3 (N21878, N21875, N20521, N4435);
not NOT1 (N21879, N21862);
buf BUF1 (N21880, N21848);
or OR3 (N21881, N21878, N231, N3225);
xor XOR2 (N21882, N21876, N13469);
nand NAND3 (N21883, N21877, N2188, N8614);
nor NOR3 (N21884, N21867, N13487, N6579);
buf BUF1 (N21885, N21874);
nor NOR3 (N21886, N21880, N6801, N16285);
nor NOR4 (N21887, N21883, N17332, N1703, N21811);
xor XOR2 (N21888, N21869, N1525);
not NOT1 (N21889, N21884);
xor XOR2 (N21890, N21882, N1210);
xor XOR2 (N21891, N21879, N17010);
or OR4 (N21892, N21888, N1032, N12271, N15768);
or OR2 (N21893, N21873, N4113);
nand NAND4 (N21894, N21852, N15854, N1211, N19337);
nand NAND3 (N21895, N21890, N1665, N8585);
buf BUF1 (N21896, N21892);
xor XOR2 (N21897, N21895, N1647);
xor XOR2 (N21898, N21897, N11118);
xor XOR2 (N21899, N21896, N20271);
xor XOR2 (N21900, N21886, N19500);
or OR4 (N21901, N21887, N13031, N19615, N14869);
nand NAND3 (N21902, N21893, N21022, N5246);
or OR4 (N21903, N21891, N12579, N17695, N1494);
nor NOR2 (N21904, N21903, N19957);
and AND3 (N21905, N21902, N1908, N7621);
not NOT1 (N21906, N21899);
or OR3 (N21907, N21885, N9145, N19190);
nor NOR4 (N21908, N21894, N2087, N12266, N21577);
nor NOR4 (N21909, N21908, N8296, N8629, N8248);
nand NAND2 (N21910, N21905, N18893);
xor XOR2 (N21911, N21898, N12351);
buf BUF1 (N21912, N21907);
nor NOR3 (N21913, N21911, N11917, N3089);
nor NOR2 (N21914, N21904, N7568);
xor XOR2 (N21915, N21913, N7103);
xor XOR2 (N21916, N21881, N9403);
nand NAND4 (N21917, N21915, N4979, N21799, N16862);
nor NOR2 (N21918, N21889, N1169);
or OR3 (N21919, N21912, N19439, N790);
or OR2 (N21920, N21909, N7436);
or OR4 (N21921, N21900, N11572, N887, N5428);
nor NOR2 (N21922, N21910, N20634);
buf BUF1 (N21923, N21901);
xor XOR2 (N21924, N21918, N1363);
nor NOR3 (N21925, N21906, N16266, N11945);
nand NAND2 (N21926, N21924, N19380);
nor NOR2 (N21927, N21926, N1670);
buf BUF1 (N21928, N21921);
buf BUF1 (N21929, N21923);
nand NAND2 (N21930, N21928, N17210);
or OR4 (N21931, N21929, N21773, N16537, N4852);
nand NAND2 (N21932, N21922, N18586);
nand NAND3 (N21933, N21919, N15311, N15291);
nand NAND4 (N21934, N21916, N4241, N10075, N21206);
xor XOR2 (N21935, N21914, N6281);
or OR2 (N21936, N21935, N132);
and AND3 (N21937, N21933, N18423, N13808);
not NOT1 (N21938, N21917);
and AND4 (N21939, N21927, N15632, N2326, N16832);
and AND3 (N21940, N21930, N8177, N17384);
buf BUF1 (N21941, N21936);
not NOT1 (N21942, N21932);
or OR2 (N21943, N21931, N12829);
nand NAND2 (N21944, N21939, N7977);
and AND3 (N21945, N21934, N10715, N6845);
and AND3 (N21946, N21937, N8757, N7992);
nand NAND4 (N21947, N21940, N20674, N19586, N13244);
buf BUF1 (N21948, N21920);
nand NAND4 (N21949, N21938, N12109, N11906, N11126);
xor XOR2 (N21950, N21944, N15095);
nor NOR4 (N21951, N21942, N18793, N14803, N1991);
nor NOR3 (N21952, N21951, N1906, N10554);
xor XOR2 (N21953, N21941, N9431);
and AND3 (N21954, N21949, N8140, N18649);
xor XOR2 (N21955, N21947, N15193);
not NOT1 (N21956, N21950);
buf BUF1 (N21957, N21925);
nand NAND2 (N21958, N21956, N17925);
nor NOR3 (N21959, N21945, N6034, N15026);
and AND4 (N21960, N21948, N14270, N16677, N21669);
not NOT1 (N21961, N21946);
and AND3 (N21962, N21960, N19926, N1150);
nor NOR3 (N21963, N21962, N2296, N15164);
nand NAND2 (N21964, N21963, N16382);
and AND4 (N21965, N21953, N4140, N15805, N7248);
not NOT1 (N21966, N21943);
xor XOR2 (N21967, N21966, N6877);
xor XOR2 (N21968, N21967, N10954);
nor NOR2 (N21969, N21961, N1881);
or OR2 (N21970, N21955, N6314);
nor NOR4 (N21971, N21954, N13492, N2485, N19667);
or OR3 (N21972, N21958, N17563, N10076);
nand NAND4 (N21973, N21965, N16833, N18611, N11354);
not NOT1 (N21974, N21968);
nor NOR2 (N21975, N21952, N4724);
not NOT1 (N21976, N21964);
or OR2 (N21977, N21969, N6537);
and AND3 (N21978, N21971, N2418, N14211);
or OR4 (N21979, N21974, N8181, N388, N4791);
buf BUF1 (N21980, N21970);
and AND3 (N21981, N21977, N7065, N14612);
or OR4 (N21982, N21980, N2392, N16404, N18590);
buf BUF1 (N21983, N21957);
nor NOR2 (N21984, N21982, N13051);
or OR2 (N21985, N21975, N663);
and AND4 (N21986, N21973, N5727, N2195, N12974);
nor NOR3 (N21987, N21981, N11754, N3373);
buf BUF1 (N21988, N21984);
buf BUF1 (N21989, N21972);
nor NOR3 (N21990, N21976, N5145, N9538);
nand NAND3 (N21991, N21989, N1952, N19110);
nor NOR4 (N21992, N21991, N13707, N6168, N33);
and AND2 (N21993, N21987, N5674);
and AND4 (N21994, N21978, N13351, N13114, N11407);
buf BUF1 (N21995, N21986);
xor XOR2 (N21996, N21993, N2674);
or OR2 (N21997, N21995, N1287);
or OR3 (N21998, N21992, N3938, N16150);
buf BUF1 (N21999, N21959);
not NOT1 (N22000, N21985);
nor NOR2 (N22001, N21998, N5869);
buf BUF1 (N22002, N21979);
and AND3 (N22003, N22000, N970, N12199);
xor XOR2 (N22004, N21999, N4084);
or OR2 (N22005, N21988, N21796);
or OR3 (N22006, N21990, N19480, N6898);
nor NOR3 (N22007, N21983, N19765, N7872);
and AND2 (N22008, N22007, N11379);
and AND2 (N22009, N22008, N20093);
not NOT1 (N22010, N21997);
xor XOR2 (N22011, N21994, N20142);
nor NOR4 (N22012, N21996, N3488, N3669, N19514);
nor NOR3 (N22013, N22005, N15555, N9850);
nor NOR3 (N22014, N22002, N7351, N9831);
nand NAND2 (N22015, N22009, N3251);
nand NAND2 (N22016, N22004, N8342);
or OR4 (N22017, N22011, N2296, N15993, N17840);
and AND4 (N22018, N22017, N17710, N19642, N13256);
or OR3 (N22019, N22018, N2079, N6646);
buf BUF1 (N22020, N22012);
not NOT1 (N22021, N22003);
nor NOR4 (N22022, N22001, N2063, N15639, N7709);
nor NOR3 (N22023, N22019, N18030, N1357);
nor NOR4 (N22024, N22023, N10511, N15366, N2952);
xor XOR2 (N22025, N22016, N9005);
or OR2 (N22026, N22024, N1698);
nand NAND3 (N22027, N22020, N18879, N12027);
xor XOR2 (N22028, N22026, N8619);
and AND4 (N22029, N22006, N6630, N17369, N5130);
buf BUF1 (N22030, N22013);
buf BUF1 (N22031, N22025);
xor XOR2 (N22032, N22022, N4619);
and AND4 (N22033, N22030, N19388, N1109, N2288);
or OR4 (N22034, N22010, N16941, N2552, N4589);
or OR3 (N22035, N22028, N14129, N17161);
xor XOR2 (N22036, N22021, N14682);
and AND3 (N22037, N22035, N18955, N20510);
nor NOR2 (N22038, N22037, N2047);
and AND3 (N22039, N22034, N2242, N5624);
nor NOR4 (N22040, N22033, N15535, N20487, N7967);
nand NAND4 (N22041, N22027, N5892, N3700, N8093);
nor NOR4 (N22042, N22038, N5258, N15959, N3238);
and AND2 (N22043, N22014, N17485);
nand NAND4 (N22044, N22042, N16138, N6697, N4842);
nand NAND4 (N22045, N22036, N20458, N14774, N17691);
nand NAND4 (N22046, N22015, N10453, N2157, N16748);
or OR2 (N22047, N22040, N20124);
not NOT1 (N22048, N22046);
or OR3 (N22049, N22047, N7324, N12546);
nor NOR2 (N22050, N22049, N244);
nor NOR3 (N22051, N22039, N8410, N14231);
and AND3 (N22052, N22041, N16706, N9748);
xor XOR2 (N22053, N22044, N18517);
not NOT1 (N22054, N22043);
nor NOR4 (N22055, N22052, N3366, N9594, N4672);
not NOT1 (N22056, N22032);
and AND2 (N22057, N22054, N12848);
nor NOR4 (N22058, N22055, N21129, N7842, N15055);
not NOT1 (N22059, N22053);
nor NOR4 (N22060, N22051, N20478, N15427, N21210);
nor NOR4 (N22061, N22060, N13465, N5760, N19447);
and AND2 (N22062, N22058, N9955);
or OR3 (N22063, N22062, N16953, N4441);
nor NOR3 (N22064, N22057, N4036, N15340);
not NOT1 (N22065, N22029);
not NOT1 (N22066, N22048);
nor NOR4 (N22067, N22045, N16817, N18401, N7645);
or OR4 (N22068, N22064, N4273, N12493, N16243);
not NOT1 (N22069, N22050);
and AND3 (N22070, N22066, N1064, N17877);
not NOT1 (N22071, N22031);
not NOT1 (N22072, N22070);
and AND2 (N22073, N22065, N5308);
and AND4 (N22074, N22073, N21024, N12443, N10522);
or OR3 (N22075, N22069, N19332, N21861);
and AND2 (N22076, N22059, N10078);
or OR4 (N22077, N22061, N20504, N152, N14320);
nor NOR3 (N22078, N22068, N16910, N18211);
nor NOR4 (N22079, N22076, N11142, N10733, N20474);
xor XOR2 (N22080, N22074, N20884);
or OR3 (N22081, N22079, N17895, N4222);
not NOT1 (N22082, N22075);
nand NAND3 (N22083, N22078, N14254, N3338);
and AND3 (N22084, N22080, N7751, N10046);
xor XOR2 (N22085, N22082, N10208);
and AND3 (N22086, N22085, N19485, N9814);
and AND4 (N22087, N22083, N14024, N14239, N8990);
nand NAND3 (N22088, N22056, N1366, N7587);
or OR4 (N22089, N22071, N1507, N410, N14263);
buf BUF1 (N22090, N22077);
nand NAND3 (N22091, N22089, N11021, N16616);
nand NAND4 (N22092, N22086, N12642, N17055, N5038);
or OR3 (N22093, N22063, N20086, N20845);
not NOT1 (N22094, N22084);
and AND3 (N22095, N22094, N10018, N3281);
buf BUF1 (N22096, N22088);
nand NAND4 (N22097, N22081, N16174, N19340, N11657);
or OR3 (N22098, N22093, N8919, N3015);
buf BUF1 (N22099, N22097);
buf BUF1 (N22100, N22098);
buf BUF1 (N22101, N22087);
xor XOR2 (N22102, N22092, N18514);
or OR2 (N22103, N22067, N11973);
and AND3 (N22104, N22096, N18324, N16340);
nand NAND3 (N22105, N22091, N19818, N19753);
nand NAND2 (N22106, N22101, N15551);
nand NAND2 (N22107, N22103, N7337);
not NOT1 (N22108, N22099);
and AND4 (N22109, N22095, N4030, N16114, N21923);
buf BUF1 (N22110, N22109);
buf BUF1 (N22111, N22104);
nand NAND3 (N22112, N22102, N7465, N14861);
and AND3 (N22113, N22100, N19319, N2465);
not NOT1 (N22114, N22090);
not NOT1 (N22115, N22072);
buf BUF1 (N22116, N22111);
not NOT1 (N22117, N22112);
nand NAND2 (N22118, N22115, N8540);
and AND2 (N22119, N22110, N13554);
buf BUF1 (N22120, N22113);
or OR2 (N22121, N22119, N17019);
nor NOR3 (N22122, N22118, N153, N21254);
nor NOR4 (N22123, N22105, N14259, N4495, N3304);
or OR2 (N22124, N22122, N7376);
nand NAND3 (N22125, N22107, N656, N5030);
and AND2 (N22126, N22114, N1195);
and AND2 (N22127, N22117, N22003);
and AND3 (N22128, N22123, N4236, N11486);
or OR4 (N22129, N22124, N16047, N13695, N21440);
nor NOR4 (N22130, N22106, N13233, N5052, N9254);
not NOT1 (N22131, N22125);
or OR4 (N22132, N22131, N22122, N17378, N4723);
not NOT1 (N22133, N22132);
nand NAND3 (N22134, N22108, N6938, N20446);
or OR3 (N22135, N22126, N5382, N1193);
and AND3 (N22136, N22133, N3259, N7005);
nand NAND3 (N22137, N22121, N18167, N7935);
xor XOR2 (N22138, N22136, N5759);
and AND4 (N22139, N22130, N11051, N12996, N10616);
nor NOR3 (N22140, N22137, N16135, N15675);
xor XOR2 (N22141, N22135, N1942);
or OR2 (N22142, N22138, N4582);
buf BUF1 (N22143, N22129);
buf BUF1 (N22144, N22143);
or OR3 (N22145, N22141, N21834, N4737);
and AND2 (N22146, N22128, N13443);
and AND4 (N22147, N22145, N2130, N8710, N12356);
or OR2 (N22148, N22127, N5530);
xor XOR2 (N22149, N22142, N555);
xor XOR2 (N22150, N22116, N10378);
nor NOR3 (N22151, N22149, N15686, N16984);
nor NOR3 (N22152, N22140, N14529, N9840);
and AND2 (N22153, N22150, N14928);
buf BUF1 (N22154, N22134);
xor XOR2 (N22155, N22144, N12080);
xor XOR2 (N22156, N22155, N17638);
buf BUF1 (N22157, N22154);
not NOT1 (N22158, N22147);
and AND2 (N22159, N22148, N21203);
nor NOR3 (N22160, N22159, N2904, N2486);
nand NAND3 (N22161, N22152, N1568, N12480);
not NOT1 (N22162, N22160);
not NOT1 (N22163, N22157);
buf BUF1 (N22164, N22151);
nor NOR3 (N22165, N22158, N14800, N8824);
buf BUF1 (N22166, N22165);
not NOT1 (N22167, N22120);
xor XOR2 (N22168, N22161, N7384);
nor NOR2 (N22169, N22156, N15166);
xor XOR2 (N22170, N22139, N17938);
buf BUF1 (N22171, N22164);
buf BUF1 (N22172, N22169);
not NOT1 (N22173, N22153);
nor NOR4 (N22174, N22173, N15315, N13599, N9454);
nand NAND2 (N22175, N22163, N12591);
and AND3 (N22176, N22174, N10225, N8145);
and AND3 (N22177, N22176, N10288, N4850);
nor NOR2 (N22178, N22175, N398);
xor XOR2 (N22179, N22170, N10347);
nor NOR2 (N22180, N22166, N21513);
not NOT1 (N22181, N22180);
xor XOR2 (N22182, N22172, N15258);
buf BUF1 (N22183, N22182);
nor NOR4 (N22184, N22146, N6073, N2157, N15160);
not NOT1 (N22185, N22178);
xor XOR2 (N22186, N22184, N7104);
and AND4 (N22187, N22168, N11255, N9815, N20902);
not NOT1 (N22188, N22179);
not NOT1 (N22189, N22185);
nand NAND2 (N22190, N22177, N7850);
or OR2 (N22191, N22187, N15734);
xor XOR2 (N22192, N22183, N7380);
and AND3 (N22193, N22189, N17991, N12891);
nand NAND3 (N22194, N22181, N20522, N6496);
and AND3 (N22195, N22191, N7416, N7491);
xor XOR2 (N22196, N22167, N4971);
not NOT1 (N22197, N22195);
or OR4 (N22198, N22188, N2691, N13075, N16089);
or OR3 (N22199, N22197, N1979, N21940);
and AND2 (N22200, N22198, N11224);
nor NOR3 (N22201, N22190, N11374, N6631);
not NOT1 (N22202, N22192);
nand NAND4 (N22203, N22196, N785, N7444, N612);
or OR3 (N22204, N22200, N13001, N17241);
not NOT1 (N22205, N22201);
nand NAND2 (N22206, N22193, N18370);
xor XOR2 (N22207, N22205, N19170);
and AND3 (N22208, N22194, N16406, N21920);
nand NAND2 (N22209, N22199, N4086);
xor XOR2 (N22210, N22171, N15060);
nand NAND3 (N22211, N22210, N12438, N14029);
and AND2 (N22212, N22203, N7355);
nand NAND4 (N22213, N22206, N3777, N8938, N6725);
buf BUF1 (N22214, N22213);
and AND3 (N22215, N22209, N15091, N13354);
nor NOR4 (N22216, N22207, N17525, N19475, N1987);
not NOT1 (N22217, N22216);
xor XOR2 (N22218, N22214, N3186);
xor XOR2 (N22219, N22208, N3950);
buf BUF1 (N22220, N22219);
or OR2 (N22221, N22204, N2970);
or OR2 (N22222, N22202, N17082);
buf BUF1 (N22223, N22220);
nand NAND3 (N22224, N22186, N4387, N12651);
nor NOR2 (N22225, N22162, N17996);
xor XOR2 (N22226, N22217, N9334);
and AND3 (N22227, N22222, N21565, N783);
nand NAND2 (N22228, N22223, N2662);
buf BUF1 (N22229, N22212);
not NOT1 (N22230, N22218);
nand NAND2 (N22231, N22229, N14077);
buf BUF1 (N22232, N22215);
nand NAND4 (N22233, N22221, N5428, N15076, N14587);
or OR3 (N22234, N22226, N7140, N16436);
nor NOR2 (N22235, N22234, N2962);
buf BUF1 (N22236, N22225);
not NOT1 (N22237, N22230);
xor XOR2 (N22238, N22232, N7148);
not NOT1 (N22239, N22227);
nand NAND4 (N22240, N22231, N8388, N19791, N11746);
and AND4 (N22241, N22224, N8605, N14976, N4899);
nor NOR2 (N22242, N22228, N11806);
buf BUF1 (N22243, N22211);
not NOT1 (N22244, N22242);
and AND3 (N22245, N22233, N18002, N13954);
or OR3 (N22246, N22238, N4609, N18225);
buf BUF1 (N22247, N22244);
or OR2 (N22248, N22245, N13183);
and AND3 (N22249, N22246, N1831, N16859);
nand NAND3 (N22250, N22235, N9330, N10320);
nor NOR3 (N22251, N22236, N15817, N11079);
not NOT1 (N22252, N22241);
nor NOR3 (N22253, N22243, N10104, N12835);
nor NOR3 (N22254, N22237, N6323, N17365);
xor XOR2 (N22255, N22253, N17077);
or OR4 (N22256, N22254, N10636, N4621, N5759);
buf BUF1 (N22257, N22249);
not NOT1 (N22258, N22257);
or OR3 (N22259, N22251, N3600, N11389);
nand NAND4 (N22260, N22248, N894, N4929, N15221);
and AND3 (N22261, N22250, N17613, N17791);
nand NAND3 (N22262, N22258, N21289, N3138);
or OR4 (N22263, N22255, N14573, N13631, N282);
xor XOR2 (N22264, N22256, N5897);
and AND3 (N22265, N22259, N15466, N10994);
buf BUF1 (N22266, N22263);
nor NOR2 (N22267, N22239, N14087);
and AND2 (N22268, N22267, N15252);
and AND2 (N22269, N22260, N5783);
and AND2 (N22270, N22252, N5471);
nand NAND2 (N22271, N22247, N18625);
buf BUF1 (N22272, N22264);
nor NOR4 (N22273, N22262, N7330, N15177, N22105);
nor NOR2 (N22274, N22240, N14587);
not NOT1 (N22275, N22261);
nand NAND3 (N22276, N22271, N8465, N4601);
nand NAND4 (N22277, N22272, N20791, N4521, N9998);
not NOT1 (N22278, N22273);
and AND4 (N22279, N22278, N3648, N9756, N7946);
xor XOR2 (N22280, N22269, N9282);
nor NOR4 (N22281, N22274, N21714, N7010, N2824);
nor NOR2 (N22282, N22266, N7856);
xor XOR2 (N22283, N22281, N20958);
nand NAND3 (N22284, N22283, N6726, N4493);
nand NAND2 (N22285, N22282, N5502);
or OR2 (N22286, N22268, N6221);
nand NAND4 (N22287, N22275, N12346, N20866, N10326);
nand NAND2 (N22288, N22287, N6831);
or OR4 (N22289, N22285, N16225, N16810, N11047);
buf BUF1 (N22290, N22279);
and AND4 (N22291, N22286, N1514, N7095, N15485);
nand NAND4 (N22292, N22280, N355, N20, N9430);
not NOT1 (N22293, N22288);
nor NOR2 (N22294, N22284, N16656);
buf BUF1 (N22295, N22291);
nor NOR3 (N22296, N22293, N7848, N16903);
xor XOR2 (N22297, N22276, N8856);
nand NAND2 (N22298, N22294, N19515);
not NOT1 (N22299, N22265);
not NOT1 (N22300, N22270);
nor NOR2 (N22301, N22295, N2795);
buf BUF1 (N22302, N22298);
nor NOR2 (N22303, N22292, N10196);
xor XOR2 (N22304, N22277, N21910);
buf BUF1 (N22305, N22289);
xor XOR2 (N22306, N22297, N6201);
not NOT1 (N22307, N22303);
xor XOR2 (N22308, N22296, N19173);
nand NAND2 (N22309, N22306, N18457);
nand NAND2 (N22310, N22307, N3462);
buf BUF1 (N22311, N22300);
not NOT1 (N22312, N22305);
buf BUF1 (N22313, N22301);
nand NAND2 (N22314, N22313, N5472);
xor XOR2 (N22315, N22309, N19067);
nand NAND2 (N22316, N22314, N4409);
nand NAND4 (N22317, N22308, N11206, N8385, N6321);
xor XOR2 (N22318, N22311, N21955);
nand NAND3 (N22319, N22304, N13191, N21375);
buf BUF1 (N22320, N22319);
and AND2 (N22321, N22316, N17827);
or OR2 (N22322, N22302, N13460);
buf BUF1 (N22323, N22310);
not NOT1 (N22324, N22321);
not NOT1 (N22325, N22323);
nor NOR3 (N22326, N22325, N12879, N13096);
xor XOR2 (N22327, N22299, N20272);
xor XOR2 (N22328, N22320, N686);
nand NAND4 (N22329, N22317, N10626, N20191, N6347);
not NOT1 (N22330, N22290);
not NOT1 (N22331, N22312);
and AND2 (N22332, N22315, N10496);
and AND2 (N22333, N22324, N2590);
not NOT1 (N22334, N22327);
nor NOR2 (N22335, N22328, N17985);
buf BUF1 (N22336, N22332);
not NOT1 (N22337, N22322);
or OR3 (N22338, N22331, N18702, N18850);
buf BUF1 (N22339, N22318);
and AND4 (N22340, N22334, N5498, N6706, N14544);
and AND4 (N22341, N22340, N8775, N8448, N13641);
nand NAND4 (N22342, N22338, N17380, N7440, N3367);
nor NOR3 (N22343, N22337, N229, N18666);
nand NAND3 (N22344, N22341, N7150, N15096);
nor NOR2 (N22345, N22342, N20163);
or OR3 (N22346, N22333, N12271, N9351);
and AND2 (N22347, N22345, N1435);
or OR2 (N22348, N22326, N12739);
not NOT1 (N22349, N22346);
and AND3 (N22350, N22335, N3201, N19933);
nand NAND2 (N22351, N22349, N11274);
nor NOR3 (N22352, N22344, N14924, N14323);
nor NOR4 (N22353, N22352, N14076, N21925, N4686);
nor NOR4 (N22354, N22348, N3759, N14007, N21761);
and AND4 (N22355, N22347, N7558, N3664, N10136);
buf BUF1 (N22356, N22343);
buf BUF1 (N22357, N22353);
xor XOR2 (N22358, N22350, N11443);
or OR2 (N22359, N22354, N2112);
or OR2 (N22360, N22329, N13376);
nand NAND4 (N22361, N22359, N7652, N316, N4340);
not NOT1 (N22362, N22361);
nor NOR2 (N22363, N22330, N12394);
xor XOR2 (N22364, N22363, N6142);
nor NOR4 (N22365, N22360, N17897, N16844, N19381);
xor XOR2 (N22366, N22364, N8106);
and AND2 (N22367, N22356, N964);
or OR4 (N22368, N22336, N19856, N2739, N19056);
buf BUF1 (N22369, N22355);
buf BUF1 (N22370, N22367);
buf BUF1 (N22371, N22362);
nand NAND2 (N22372, N22365, N734);
or OR4 (N22373, N22368, N13208, N19146, N15687);
nor NOR2 (N22374, N22371, N8971);
not NOT1 (N22375, N22369);
nand NAND2 (N22376, N22358, N6821);
xor XOR2 (N22377, N22372, N17913);
nor NOR2 (N22378, N22370, N13522);
or OR2 (N22379, N22375, N7471);
and AND3 (N22380, N22351, N5070, N10177);
nand NAND3 (N22381, N22366, N20045, N5533);
or OR3 (N22382, N22377, N16237, N2986);
not NOT1 (N22383, N22379);
not NOT1 (N22384, N22383);
or OR2 (N22385, N22381, N8362);
xor XOR2 (N22386, N22373, N2280);
and AND3 (N22387, N22386, N2463, N3084);
not NOT1 (N22388, N22378);
xor XOR2 (N22389, N22387, N6171);
nand NAND4 (N22390, N22376, N15412, N14520, N15336);
not NOT1 (N22391, N22382);
xor XOR2 (N22392, N22339, N20614);
xor XOR2 (N22393, N22388, N15334);
and AND3 (N22394, N22385, N333, N13653);
buf BUF1 (N22395, N22384);
and AND3 (N22396, N22391, N19529, N5529);
and AND4 (N22397, N22357, N13171, N3677, N5964);
buf BUF1 (N22398, N22393);
buf BUF1 (N22399, N22396);
nor NOR2 (N22400, N22389, N19071);
and AND3 (N22401, N22374, N11867, N3687);
and AND4 (N22402, N22400, N9181, N1889, N3759);
nand NAND4 (N22403, N22392, N9649, N15269, N16055);
xor XOR2 (N22404, N22401, N6919);
xor XOR2 (N22405, N22404, N11929);
buf BUF1 (N22406, N22395);
and AND3 (N22407, N22398, N16528, N8161);
or OR3 (N22408, N22405, N12686, N20194);
nand NAND3 (N22409, N22399, N3562, N15384);
buf BUF1 (N22410, N22380);
buf BUF1 (N22411, N22410);
buf BUF1 (N22412, N22403);
or OR3 (N22413, N22409, N309, N15036);
nor NOR4 (N22414, N22394, N10327, N13798, N12644);
or OR3 (N22415, N22414, N17337, N2739);
nand NAND3 (N22416, N22411, N11270, N19139);
buf BUF1 (N22417, N22413);
not NOT1 (N22418, N22408);
buf BUF1 (N22419, N22415);
buf BUF1 (N22420, N22407);
not NOT1 (N22421, N22417);
or OR4 (N22422, N22397, N2776, N16880, N9018);
and AND3 (N22423, N22402, N3392, N16845);
xor XOR2 (N22424, N22419, N18780);
buf BUF1 (N22425, N22420);
and AND3 (N22426, N22424, N9443, N19992);
buf BUF1 (N22427, N22390);
xor XOR2 (N22428, N22418, N20109);
xor XOR2 (N22429, N22412, N6716);
and AND4 (N22430, N22406, N18194, N11262, N3132);
nand NAND2 (N22431, N22429, N21975);
or OR4 (N22432, N22428, N13110, N14999, N884);
nor NOR4 (N22433, N22431, N8441, N5197, N10510);
nand NAND2 (N22434, N22416, N16941);
xor XOR2 (N22435, N22427, N18527);
nor NOR2 (N22436, N22432, N21073);
or OR4 (N22437, N22423, N16508, N17945, N16120);
not NOT1 (N22438, N22422);
and AND3 (N22439, N22435, N18215, N5804);
not NOT1 (N22440, N22425);
and AND4 (N22441, N22437, N22344, N4132, N8781);
nand NAND4 (N22442, N22433, N1635, N1626, N10231);
xor XOR2 (N22443, N22442, N8012);
or OR3 (N22444, N22443, N16414, N21489);
nor NOR4 (N22445, N22441, N19155, N2267, N582);
xor XOR2 (N22446, N22426, N16745);
nor NOR3 (N22447, N22421, N9431, N14294);
buf BUF1 (N22448, N22446);
nand NAND2 (N22449, N22438, N12593);
xor XOR2 (N22450, N22445, N1673);
and AND4 (N22451, N22439, N17049, N1276, N4186);
buf BUF1 (N22452, N22444);
or OR3 (N22453, N22447, N3804, N15722);
buf BUF1 (N22454, N22448);
buf BUF1 (N22455, N22454);
xor XOR2 (N22456, N22449, N12533);
not NOT1 (N22457, N22430);
and AND2 (N22458, N22440, N13653);
or OR2 (N22459, N22455, N21317);
or OR3 (N22460, N22436, N6818, N1198);
not NOT1 (N22461, N22456);
buf BUF1 (N22462, N22451);
not NOT1 (N22463, N22460);
and AND2 (N22464, N22434, N12954);
nand NAND2 (N22465, N22463, N21790);
or OR2 (N22466, N22457, N12582);
and AND3 (N22467, N22450, N5531, N2770);
and AND3 (N22468, N22465, N17439, N11720);
or OR4 (N22469, N22462, N7644, N11022, N665);
buf BUF1 (N22470, N22459);
buf BUF1 (N22471, N22458);
not NOT1 (N22472, N22453);
xor XOR2 (N22473, N22468, N15117);
nand NAND2 (N22474, N22452, N6495);
buf BUF1 (N22475, N22471);
xor XOR2 (N22476, N22473, N21921);
and AND4 (N22477, N22474, N18339, N9835, N19431);
nor NOR2 (N22478, N22470, N20504);
buf BUF1 (N22479, N22464);
and AND4 (N22480, N22472, N16945, N11995, N9808);
xor XOR2 (N22481, N22478, N8144);
xor XOR2 (N22482, N22461, N14051);
nand NAND3 (N22483, N22477, N18672, N1188);
or OR2 (N22484, N22481, N17751);
buf BUF1 (N22485, N22469);
not NOT1 (N22486, N22484);
or OR2 (N22487, N22480, N17685);
nor NOR3 (N22488, N22487, N14900, N17973);
not NOT1 (N22489, N22467);
nand NAND4 (N22490, N22482, N16279, N11207, N17810);
and AND2 (N22491, N22476, N17583);
not NOT1 (N22492, N22489);
or OR2 (N22493, N22491, N15285);
not NOT1 (N22494, N22466);
and AND3 (N22495, N22485, N10349, N8938);
nand NAND3 (N22496, N22486, N4705, N20811);
nor NOR3 (N22497, N22494, N21338, N5782);
not NOT1 (N22498, N22493);
and AND3 (N22499, N22483, N16360, N12054);
and AND2 (N22500, N22475, N14361);
buf BUF1 (N22501, N22490);
and AND4 (N22502, N22501, N5774, N10079, N2619);
xor XOR2 (N22503, N22488, N2462);
not NOT1 (N22504, N22503);
nor NOR2 (N22505, N22498, N15580);
buf BUF1 (N22506, N22499);
nor NOR2 (N22507, N22496, N11852);
nor NOR2 (N22508, N22502, N11786);
and AND2 (N22509, N22504, N6709);
xor XOR2 (N22510, N22507, N10941);
not NOT1 (N22511, N22506);
not NOT1 (N22512, N22497);
not NOT1 (N22513, N22479);
not NOT1 (N22514, N22492);
xor XOR2 (N22515, N22500, N20017);
and AND2 (N22516, N22495, N2386);
buf BUF1 (N22517, N22514);
xor XOR2 (N22518, N22511, N21871);
nand NAND2 (N22519, N22512, N8958);
xor XOR2 (N22520, N22519, N5727);
or OR4 (N22521, N22520, N15442, N5676, N11490);
not NOT1 (N22522, N22518);
nor NOR3 (N22523, N22521, N9664, N11825);
or OR2 (N22524, N22510, N7792);
xor XOR2 (N22525, N22516, N5651);
buf BUF1 (N22526, N22525);
buf BUF1 (N22527, N22509);
buf BUF1 (N22528, N22527);
buf BUF1 (N22529, N22515);
not NOT1 (N22530, N22524);
nand NAND3 (N22531, N22522, N18985, N13520);
nand NAND2 (N22532, N22505, N21679);
and AND3 (N22533, N22531, N3708, N18941);
not NOT1 (N22534, N22513);
nand NAND3 (N22535, N22523, N10832, N5193);
nand NAND3 (N22536, N22508, N21998, N17923);
nor NOR2 (N22537, N22535, N9906);
nand NAND3 (N22538, N22528, N21676, N2757);
not NOT1 (N22539, N22530);
buf BUF1 (N22540, N22539);
buf BUF1 (N22541, N22517);
and AND2 (N22542, N22540, N10477);
not NOT1 (N22543, N22534);
xor XOR2 (N22544, N22536, N19236);
nand NAND3 (N22545, N22532, N12356, N7595);
or OR3 (N22546, N22542, N2411, N17211);
nor NOR2 (N22547, N22526, N289);
xor XOR2 (N22548, N22544, N6774);
buf BUF1 (N22549, N22533);
and AND3 (N22550, N22529, N18231, N8276);
or OR3 (N22551, N22549, N5447, N12394);
xor XOR2 (N22552, N22541, N10874);
nor NOR2 (N22553, N22538, N20405);
xor XOR2 (N22554, N22537, N17482);
xor XOR2 (N22555, N22552, N69);
nor NOR2 (N22556, N22547, N4674);
not NOT1 (N22557, N22551);
xor XOR2 (N22558, N22546, N1908);
nor NOR2 (N22559, N22555, N17169);
and AND2 (N22560, N22559, N10546);
nor NOR3 (N22561, N22548, N2883, N19796);
nor NOR3 (N22562, N22550, N20363, N22501);
and AND4 (N22563, N22562, N21258, N12206, N16646);
buf BUF1 (N22564, N22558);
xor XOR2 (N22565, N22563, N20665);
nand NAND2 (N22566, N22561, N13703);
buf BUF1 (N22567, N22557);
and AND3 (N22568, N22554, N18053, N13154);
and AND4 (N22569, N22553, N292, N16512, N10730);
or OR4 (N22570, N22565, N14085, N20563, N21701);
buf BUF1 (N22571, N22570);
nand NAND4 (N22572, N22545, N14999, N21988, N11979);
not NOT1 (N22573, N22571);
buf BUF1 (N22574, N22560);
or OR4 (N22575, N22573, N10238, N14951, N20228);
and AND2 (N22576, N22543, N9957);
nor NOR4 (N22577, N22564, N7897, N8732, N22157);
buf BUF1 (N22578, N22577);
and AND2 (N22579, N22578, N13145);
nor NOR4 (N22580, N22568, N630, N15395, N13443);
xor XOR2 (N22581, N22567, N12986);
nand NAND3 (N22582, N22581, N9801, N16848);
and AND3 (N22583, N22575, N15459, N7589);
nand NAND2 (N22584, N22580, N19168);
nand NAND3 (N22585, N22574, N21, N15493);
xor XOR2 (N22586, N22582, N1887);
buf BUF1 (N22587, N22556);
nor NOR2 (N22588, N22586, N18817);
and AND4 (N22589, N22587, N21939, N18144, N17719);
not NOT1 (N22590, N22579);
nor NOR2 (N22591, N22583, N8510);
nand NAND3 (N22592, N22584, N8821, N13958);
and AND4 (N22593, N22589, N11436, N21716, N12532);
and AND2 (N22594, N22576, N7937);
not NOT1 (N22595, N22590);
not NOT1 (N22596, N22588);
and AND4 (N22597, N22593, N19221, N9466, N18773);
and AND4 (N22598, N22566, N4083, N5223, N15462);
or OR2 (N22599, N22598, N19356);
nand NAND3 (N22600, N22599, N10989, N18633);
xor XOR2 (N22601, N22569, N20868);
xor XOR2 (N22602, N22601, N12753);
nand NAND4 (N22603, N22595, N10259, N11864, N3552);
xor XOR2 (N22604, N22591, N608);
nor NOR3 (N22605, N22597, N162, N19095);
xor XOR2 (N22606, N22572, N96);
or OR4 (N22607, N22603, N12118, N22182, N18440);
or OR2 (N22608, N22585, N20200);
buf BUF1 (N22609, N22600);
buf BUF1 (N22610, N22604);
and AND4 (N22611, N22602, N15793, N8901, N5106);
and AND3 (N22612, N22605, N20272, N17177);
or OR2 (N22613, N22609, N13604);
not NOT1 (N22614, N22611);
xor XOR2 (N22615, N22610, N8332);
and AND3 (N22616, N22614, N16527, N821);
and AND3 (N22617, N22612, N21257, N22343);
or OR2 (N22618, N22606, N1974);
not NOT1 (N22619, N22608);
and AND3 (N22620, N22592, N10714, N4300);
buf BUF1 (N22621, N22617);
buf BUF1 (N22622, N22621);
xor XOR2 (N22623, N22616, N1176);
nor NOR4 (N22624, N22607, N5486, N16376, N16545);
buf BUF1 (N22625, N22624);
nor NOR2 (N22626, N22623, N14187);
or OR3 (N22627, N22618, N1933, N1320);
buf BUF1 (N22628, N22626);
or OR2 (N22629, N22620, N12533);
xor XOR2 (N22630, N22629, N21047);
not NOT1 (N22631, N22613);
buf BUF1 (N22632, N22631);
nand NAND2 (N22633, N22630, N4047);
xor XOR2 (N22634, N22615, N14631);
and AND2 (N22635, N22634, N6681);
and AND3 (N22636, N22625, N8274, N2329);
not NOT1 (N22637, N22596);
xor XOR2 (N22638, N22628, N10472);
not NOT1 (N22639, N22619);
xor XOR2 (N22640, N22638, N13543);
and AND4 (N22641, N22627, N4488, N1438, N18653);
buf BUF1 (N22642, N22637);
xor XOR2 (N22643, N22594, N4348);
nor NOR4 (N22644, N22622, N10207, N7788, N14624);
xor XOR2 (N22645, N22643, N6232);
nand NAND2 (N22646, N22636, N10406);
xor XOR2 (N22647, N22633, N22239);
buf BUF1 (N22648, N22632);
nor NOR4 (N22649, N22647, N16230, N5227, N15207);
or OR2 (N22650, N22639, N21115);
or OR3 (N22651, N22645, N13483, N7849);
or OR2 (N22652, N22650, N18911);
and AND4 (N22653, N22644, N21389, N20332, N12071);
or OR3 (N22654, N22642, N760, N12681);
buf BUF1 (N22655, N22651);
xor XOR2 (N22656, N22648, N20897);
xor XOR2 (N22657, N22646, N2415);
or OR4 (N22658, N22654, N15297, N7339, N21914);
nand NAND2 (N22659, N22656, N20831);
buf BUF1 (N22660, N22655);
nor NOR3 (N22661, N22649, N15037, N13360);
buf BUF1 (N22662, N22653);
nand NAND4 (N22663, N22662, N13274, N3861, N6669);
nand NAND3 (N22664, N22641, N16030, N17542);
or OR4 (N22665, N22652, N17255, N19042, N15794);
nor NOR3 (N22666, N22640, N2635, N12654);
buf BUF1 (N22667, N22665);
or OR2 (N22668, N22667, N17601);
and AND4 (N22669, N22668, N22317, N8263, N16851);
nand NAND4 (N22670, N22663, N10801, N5693, N12583);
nand NAND2 (N22671, N22657, N4279);
and AND3 (N22672, N22669, N19508, N8477);
not NOT1 (N22673, N22666);
or OR2 (N22674, N22661, N20486);
and AND4 (N22675, N22671, N5804, N9908, N10199);
or OR2 (N22676, N22670, N1450);
nand NAND2 (N22677, N22674, N15366);
xor XOR2 (N22678, N22660, N10612);
xor XOR2 (N22679, N22635, N5961);
and AND2 (N22680, N22679, N11357);
xor XOR2 (N22681, N22673, N20857);
nor NOR3 (N22682, N22675, N17472, N11899);
not NOT1 (N22683, N22659);
not NOT1 (N22684, N22678);
nor NOR3 (N22685, N22683, N9457, N9531);
nand NAND3 (N22686, N22680, N22019, N7238);
buf BUF1 (N22687, N22676);
xor XOR2 (N22688, N22685, N14021);
buf BUF1 (N22689, N22664);
buf BUF1 (N22690, N22687);
nand NAND2 (N22691, N22681, N2047);
xor XOR2 (N22692, N22684, N1621);
xor XOR2 (N22693, N22692, N596);
not NOT1 (N22694, N22658);
nand NAND4 (N22695, N22677, N4638, N9689, N6627);
buf BUF1 (N22696, N22690);
not NOT1 (N22697, N22672);
and AND4 (N22698, N22694, N3756, N10144, N14332);
not NOT1 (N22699, N22686);
not NOT1 (N22700, N22699);
nand NAND4 (N22701, N22693, N3691, N1907, N10756);
nor NOR3 (N22702, N22691, N20151, N8087);
and AND4 (N22703, N22698, N16080, N16427, N16410);
not NOT1 (N22704, N22700);
not NOT1 (N22705, N22701);
not NOT1 (N22706, N22705);
xor XOR2 (N22707, N22706, N2402);
nand NAND3 (N22708, N22688, N11975, N21535);
not NOT1 (N22709, N22695);
or OR2 (N22710, N22708, N6981);
buf BUF1 (N22711, N22689);
or OR2 (N22712, N22704, N12695);
not NOT1 (N22713, N22697);
xor XOR2 (N22714, N22711, N10437);
nor NOR2 (N22715, N22702, N8241);
or OR3 (N22716, N22713, N2285, N14228);
and AND3 (N22717, N22715, N5510, N1199);
or OR2 (N22718, N22696, N7219);
nor NOR4 (N22719, N22718, N19016, N10866, N18058);
or OR3 (N22720, N22714, N9894, N1090);
and AND3 (N22721, N22710, N9268, N4175);
xor XOR2 (N22722, N22712, N4077);
nand NAND3 (N22723, N22722, N4131, N11098);
or OR3 (N22724, N22720, N7194, N17637);
nand NAND4 (N22725, N22716, N851, N19922, N13270);
buf BUF1 (N22726, N22724);
nor NOR3 (N22727, N22703, N9136, N8680);
and AND4 (N22728, N22726, N15227, N5860, N13493);
or OR4 (N22729, N22682, N10184, N11650, N22585);
or OR4 (N22730, N22723, N10361, N4943, N14064);
or OR3 (N22731, N22729, N13944, N16061);
and AND3 (N22732, N22717, N7584, N11584);
and AND4 (N22733, N22707, N760, N6327, N21340);
buf BUF1 (N22734, N22728);
nand NAND3 (N22735, N22725, N13870, N20014);
and AND3 (N22736, N22719, N5522, N12022);
or OR3 (N22737, N22731, N9292, N11233);
buf BUF1 (N22738, N22736);
not NOT1 (N22739, N22732);
buf BUF1 (N22740, N22709);
buf BUF1 (N22741, N22739);
and AND3 (N22742, N22727, N6115, N8326);
nand NAND4 (N22743, N22730, N4994, N22178, N13313);
nor NOR3 (N22744, N22721, N21043, N10362);
and AND4 (N22745, N22735, N7993, N13854, N7631);
nand NAND3 (N22746, N22734, N20769, N2893);
and AND4 (N22747, N22745, N20393, N4122, N18837);
nor NOR2 (N22748, N22747, N20164);
nand NAND2 (N22749, N22743, N673);
nand NAND3 (N22750, N22741, N11696, N19234);
nor NOR2 (N22751, N22746, N11289);
xor XOR2 (N22752, N22751, N14883);
nor NOR2 (N22753, N22749, N4003);
xor XOR2 (N22754, N22750, N6083);
or OR3 (N22755, N22733, N8963, N493);
not NOT1 (N22756, N22754);
or OR3 (N22757, N22740, N16564, N14993);
xor XOR2 (N22758, N22756, N6030);
buf BUF1 (N22759, N22737);
nand NAND3 (N22760, N22752, N5318, N872);
nor NOR4 (N22761, N22755, N10202, N4863, N1912);
not NOT1 (N22762, N22761);
xor XOR2 (N22763, N22742, N9440);
nor NOR3 (N22764, N22760, N21814, N10151);
nand NAND2 (N22765, N22759, N18772);
buf BUF1 (N22766, N22758);
nand NAND3 (N22767, N22763, N9939, N21193);
nor NOR4 (N22768, N22762, N18151, N1295, N2744);
not NOT1 (N22769, N22767);
or OR3 (N22770, N22738, N2287, N9468);
nand NAND2 (N22771, N22753, N11305);
or OR3 (N22772, N22744, N18308, N197);
nand NAND2 (N22773, N22765, N16080);
nand NAND4 (N22774, N22768, N9456, N3716, N17483);
nand NAND4 (N22775, N22748, N5559, N14331, N8358);
nor NOR2 (N22776, N22766, N12309);
xor XOR2 (N22777, N22772, N15365);
nor NOR3 (N22778, N22769, N14529, N17443);
and AND2 (N22779, N22774, N22628);
or OR4 (N22780, N22757, N5530, N7768, N20321);
and AND4 (N22781, N22775, N6229, N13255, N18964);
xor XOR2 (N22782, N22771, N14840);
nand NAND2 (N22783, N22778, N20059);
nand NAND4 (N22784, N22773, N6562, N12646, N16627);
and AND4 (N22785, N22783, N14289, N19920, N15676);
nand NAND2 (N22786, N22782, N22276);
nand NAND2 (N22787, N22786, N5785);
not NOT1 (N22788, N22776);
and AND2 (N22789, N22788, N14958);
nor NOR3 (N22790, N22785, N3114, N15183);
or OR3 (N22791, N22789, N9691, N5282);
and AND3 (N22792, N22780, N18658, N424);
nand NAND3 (N22793, N22777, N1549, N10746);
and AND4 (N22794, N22770, N11561, N9518, N3094);
and AND4 (N22795, N22784, N22658, N22235, N14988);
nand NAND3 (N22796, N22781, N1065, N21996);
nor NOR4 (N22797, N22793, N20324, N2192, N12672);
not NOT1 (N22798, N22791);
not NOT1 (N22799, N22796);
buf BUF1 (N22800, N22764);
not NOT1 (N22801, N22800);
and AND3 (N22802, N22797, N8999, N13189);
not NOT1 (N22803, N22779);
nand NAND2 (N22804, N22787, N11774);
nor NOR2 (N22805, N22804, N20033);
buf BUF1 (N22806, N22801);
buf BUF1 (N22807, N22792);
nand NAND3 (N22808, N22790, N4716, N731);
buf BUF1 (N22809, N22802);
xor XOR2 (N22810, N22808, N13314);
not NOT1 (N22811, N22803);
nand NAND2 (N22812, N22805, N14991);
xor XOR2 (N22813, N22809, N11859);
nor NOR2 (N22814, N22812, N12875);
nand NAND2 (N22815, N22795, N19002);
or OR4 (N22816, N22798, N19021, N1182, N4335);
or OR3 (N22817, N22814, N9493, N16871);
nor NOR3 (N22818, N22799, N7409, N6173);
nand NAND2 (N22819, N22813, N20747);
not NOT1 (N22820, N22818);
xor XOR2 (N22821, N22807, N3140);
and AND2 (N22822, N22816, N9071);
nor NOR3 (N22823, N22815, N10446, N9327);
nor NOR3 (N22824, N22810, N10192, N6453);
or OR4 (N22825, N22806, N17801, N17556, N19443);
or OR3 (N22826, N22824, N14380, N11261);
nor NOR3 (N22827, N22817, N8655, N702);
nor NOR2 (N22828, N22794, N13780);
xor XOR2 (N22829, N22826, N8022);
and AND2 (N22830, N22820, N8389);
and AND3 (N22831, N22821, N17107, N13154);
and AND3 (N22832, N22827, N13765, N1076);
not NOT1 (N22833, N22831);
nand NAND2 (N22834, N22822, N14991);
not NOT1 (N22835, N22825);
nor NOR4 (N22836, N22811, N10766, N12528, N13909);
buf BUF1 (N22837, N22833);
and AND4 (N22838, N22823, N8917, N247, N355);
or OR4 (N22839, N22830, N1197, N461, N13492);
not NOT1 (N22840, N22832);
nor NOR4 (N22841, N22836, N8272, N21503, N17685);
xor XOR2 (N22842, N22841, N15821);
nand NAND4 (N22843, N22819, N6231, N15239, N12166);
xor XOR2 (N22844, N22842, N20980);
nor NOR3 (N22845, N22843, N11152, N14830);
nor NOR4 (N22846, N22834, N658, N12949, N1225);
nand NAND3 (N22847, N22840, N1711, N14888);
nand NAND3 (N22848, N22847, N20493, N5068);
xor XOR2 (N22849, N22835, N10581);
not NOT1 (N22850, N22848);
nand NAND2 (N22851, N22846, N18408);
and AND3 (N22852, N22845, N15934, N16498);
and AND3 (N22853, N22844, N10383, N15453);
xor XOR2 (N22854, N22850, N8517);
xor XOR2 (N22855, N22829, N14430);
nand NAND3 (N22856, N22837, N10190, N20666);
not NOT1 (N22857, N22828);
or OR2 (N22858, N22855, N3147);
nor NOR2 (N22859, N22853, N15404);
and AND2 (N22860, N22859, N3400);
or OR3 (N22861, N22839, N13734, N732);
xor XOR2 (N22862, N22856, N14975);
not NOT1 (N22863, N22854);
buf BUF1 (N22864, N22838);
and AND3 (N22865, N22860, N7729, N8827);
or OR2 (N22866, N22863, N17757);
nand NAND4 (N22867, N22858, N10458, N3523, N14981);
not NOT1 (N22868, N22857);
not NOT1 (N22869, N22849);
xor XOR2 (N22870, N22867, N19695);
nor NOR2 (N22871, N22865, N14262);
xor XOR2 (N22872, N22870, N13793);
or OR2 (N22873, N22866, N17032);
not NOT1 (N22874, N22861);
buf BUF1 (N22875, N22869);
nor NOR4 (N22876, N22862, N22364, N11763, N17269);
nand NAND4 (N22877, N22851, N15080, N11993, N20725);
xor XOR2 (N22878, N22873, N14579);
xor XOR2 (N22879, N22876, N19641);
not NOT1 (N22880, N22868);
nor NOR4 (N22881, N22872, N10644, N5937, N18457);
and AND2 (N22882, N22880, N11426);
and AND2 (N22883, N22874, N7810);
nand NAND3 (N22884, N22879, N10688, N21461);
nor NOR3 (N22885, N22883, N17265, N6270);
buf BUF1 (N22886, N22871);
nor NOR4 (N22887, N22852, N22837, N4056, N9993);
nor NOR2 (N22888, N22881, N18612);
nand NAND4 (N22889, N22885, N21363, N21719, N18639);
and AND2 (N22890, N22864, N17082);
not NOT1 (N22891, N22889);
and AND2 (N22892, N22888, N17174);
xor XOR2 (N22893, N22875, N8327);
nand NAND2 (N22894, N22878, N221);
nor NOR2 (N22895, N22893, N14995);
xor XOR2 (N22896, N22887, N6808);
nor NOR4 (N22897, N22884, N13933, N9738, N6754);
or OR2 (N22898, N22877, N1852);
nor NOR2 (N22899, N22890, N20739);
buf BUF1 (N22900, N22898);
not NOT1 (N22901, N22894);
buf BUF1 (N22902, N22891);
buf BUF1 (N22903, N22892);
xor XOR2 (N22904, N22895, N15028);
buf BUF1 (N22905, N22900);
not NOT1 (N22906, N22901);
or OR2 (N22907, N22896, N13996);
not NOT1 (N22908, N22904);
buf BUF1 (N22909, N22905);
not NOT1 (N22910, N22902);
not NOT1 (N22911, N22907);
nand NAND2 (N22912, N22908, N9659);
and AND4 (N22913, N22910, N21627, N4175, N5286);
and AND3 (N22914, N22903, N8731, N5985);
xor XOR2 (N22915, N22914, N16907);
nand NAND3 (N22916, N22906, N889, N16474);
not NOT1 (N22917, N22913);
not NOT1 (N22918, N22912);
not NOT1 (N22919, N22897);
not NOT1 (N22920, N22886);
buf BUF1 (N22921, N22882);
buf BUF1 (N22922, N22921);
nor NOR4 (N22923, N22920, N11146, N1517, N3486);
buf BUF1 (N22924, N22915);
not NOT1 (N22925, N22909);
nor NOR2 (N22926, N22911, N2794);
and AND3 (N22927, N22924, N12312, N6146);
or OR4 (N22928, N22899, N1012, N17430, N21748);
buf BUF1 (N22929, N22916);
buf BUF1 (N22930, N22918);
or OR4 (N22931, N22930, N6971, N1547, N20614);
xor XOR2 (N22932, N22928, N17219);
or OR3 (N22933, N22925, N1044, N868);
and AND2 (N22934, N22932, N17899);
buf BUF1 (N22935, N22927);
not NOT1 (N22936, N22922);
or OR4 (N22937, N22923, N11787, N10873, N22155);
buf BUF1 (N22938, N22931);
buf BUF1 (N22939, N22935);
and AND3 (N22940, N22933, N13578, N22164);
buf BUF1 (N22941, N22939);
nand NAND2 (N22942, N22926, N7756);
nand NAND4 (N22943, N22917, N14083, N7113, N22480);
or OR3 (N22944, N22936, N13656, N17351);
and AND2 (N22945, N22919, N672);
xor XOR2 (N22946, N22929, N5563);
buf BUF1 (N22947, N22938);
and AND4 (N22948, N22940, N17585, N22236, N20750);
or OR3 (N22949, N22942, N12871, N9373);
nand NAND3 (N22950, N22941, N3478, N19736);
not NOT1 (N22951, N22947);
nand NAND3 (N22952, N22948, N9722, N16763);
nand NAND4 (N22953, N22951, N2336, N14060, N16190);
nand NAND4 (N22954, N22944, N2093, N15914, N6702);
nand NAND3 (N22955, N22943, N5764, N13820);
nand NAND3 (N22956, N22934, N16967, N14948);
nor NOR2 (N22957, N22949, N17240);
xor XOR2 (N22958, N22946, N6696);
buf BUF1 (N22959, N22956);
buf BUF1 (N22960, N22952);
nand NAND4 (N22961, N22958, N17898, N18282, N3914);
buf BUF1 (N22962, N22953);
or OR4 (N22963, N22961, N19547, N19332, N16745);
nand NAND4 (N22964, N22954, N5698, N13071, N1383);
xor XOR2 (N22965, N22959, N13990);
xor XOR2 (N22966, N22960, N22059);
buf BUF1 (N22967, N22963);
nand NAND2 (N22968, N22945, N15083);
xor XOR2 (N22969, N22957, N3180);
xor XOR2 (N22970, N22955, N18985);
and AND4 (N22971, N22968, N5492, N20139, N6949);
xor XOR2 (N22972, N22950, N7833);
not NOT1 (N22973, N22964);
and AND4 (N22974, N22970, N22736, N8473, N19188);
or OR2 (N22975, N22972, N15497);
nand NAND3 (N22976, N22975, N10649, N21582);
xor XOR2 (N22977, N22966, N1683);
and AND2 (N22978, N22969, N10525);
not NOT1 (N22979, N22971);
nor NOR3 (N22980, N22977, N2973, N8582);
nand NAND4 (N22981, N22980, N11248, N22662, N2831);
not NOT1 (N22982, N22973);
xor XOR2 (N22983, N22974, N20326);
or OR3 (N22984, N22976, N18971, N13684);
and AND4 (N22985, N22984, N18753, N21748, N4379);
and AND4 (N22986, N22937, N13045, N727, N10618);
nor NOR3 (N22987, N22986, N8465, N22177);
xor XOR2 (N22988, N22981, N166);
buf BUF1 (N22989, N22987);
buf BUF1 (N22990, N22962);
nor NOR3 (N22991, N22979, N9545, N14698);
xor XOR2 (N22992, N22985, N132);
nor NOR4 (N22993, N22978, N10689, N18733, N7640);
buf BUF1 (N22994, N22990);
buf BUF1 (N22995, N22965);
xor XOR2 (N22996, N22992, N8645);
xor XOR2 (N22997, N22994, N4766);
buf BUF1 (N22998, N22993);
not NOT1 (N22999, N22995);
not NOT1 (N23000, N22967);
xor XOR2 (N23001, N22983, N16783);
xor XOR2 (N23002, N22989, N5273);
and AND3 (N23003, N23001, N18794, N20119);
xor XOR2 (N23004, N23000, N13835);
or OR2 (N23005, N22996, N1632);
xor XOR2 (N23006, N22991, N17432);
nand NAND4 (N23007, N23006, N20865, N9399, N1483);
or OR3 (N23008, N22988, N7739, N12911);
not NOT1 (N23009, N22998);
nor NOR2 (N23010, N23004, N837);
or OR3 (N23011, N23010, N13277, N6207);
nor NOR4 (N23012, N23007, N6512, N18939, N22802);
nand NAND2 (N23013, N23005, N19288);
not NOT1 (N23014, N22982);
not NOT1 (N23015, N23009);
nor NOR2 (N23016, N23011, N14034);
not NOT1 (N23017, N23002);
and AND2 (N23018, N23017, N15383);
or OR4 (N23019, N23014, N20877, N443, N11772);
xor XOR2 (N23020, N23018, N7045);
buf BUF1 (N23021, N23008);
xor XOR2 (N23022, N23015, N20431);
not NOT1 (N23023, N23019);
not NOT1 (N23024, N22999);
buf BUF1 (N23025, N23016);
or OR2 (N23026, N23021, N12520);
or OR3 (N23027, N23013, N5688, N1385);
buf BUF1 (N23028, N23020);
buf BUF1 (N23029, N23023);
or OR4 (N23030, N23003, N21693, N9673, N20842);
not NOT1 (N23031, N22997);
nand NAND3 (N23032, N23030, N20797, N19584);
nor NOR4 (N23033, N23012, N7332, N17672, N898);
nor NOR2 (N23034, N23024, N1849);
and AND2 (N23035, N23026, N22557);
and AND3 (N23036, N23032, N12538, N14336);
not NOT1 (N23037, N23022);
and AND3 (N23038, N23031, N14880, N18490);
nand NAND2 (N23039, N23033, N13887);
buf BUF1 (N23040, N23036);
or OR4 (N23041, N23028, N18317, N16718, N15311);
not NOT1 (N23042, N23034);
nor NOR4 (N23043, N23037, N13876, N855, N8415);
not NOT1 (N23044, N23038);
nor NOR4 (N23045, N23029, N12385, N5808, N22915);
nor NOR2 (N23046, N23025, N1834);
xor XOR2 (N23047, N23045, N195);
or OR3 (N23048, N23043, N10475, N1372);
buf BUF1 (N23049, N23027);
nand NAND2 (N23050, N23040, N11562);
and AND4 (N23051, N23041, N9276, N13603, N15740);
not NOT1 (N23052, N23042);
not NOT1 (N23053, N23047);
or OR3 (N23054, N23035, N706, N10167);
nand NAND3 (N23055, N23054, N3520, N16495);
nor NOR4 (N23056, N23055, N17481, N12851, N16138);
buf BUF1 (N23057, N23049);
and AND3 (N23058, N23052, N5844, N22447);
not NOT1 (N23059, N23057);
buf BUF1 (N23060, N23044);
not NOT1 (N23061, N23059);
nand NAND2 (N23062, N23061, N6508);
nand NAND3 (N23063, N23060, N5926, N2044);
nand NAND3 (N23064, N23039, N13096, N12981);
and AND4 (N23065, N23053, N237, N14580, N1254);
nor NOR2 (N23066, N23062, N17553);
nand NAND2 (N23067, N23064, N13946);
and AND4 (N23068, N23065, N20258, N15142, N8769);
nor NOR3 (N23069, N23063, N19223, N152);
nor NOR4 (N23070, N23069, N12758, N13752, N9899);
nand NAND3 (N23071, N23050, N3456, N6269);
nor NOR3 (N23072, N23058, N14069, N7758);
buf BUF1 (N23073, N23068);
nand NAND2 (N23074, N23072, N10215);
not NOT1 (N23075, N23051);
xor XOR2 (N23076, N23046, N11917);
nand NAND4 (N23077, N23070, N12629, N4997, N22465);
nor NOR3 (N23078, N23071, N5590, N20188);
nor NOR4 (N23079, N23056, N4952, N6579, N11252);
buf BUF1 (N23080, N23078);
not NOT1 (N23081, N23048);
and AND2 (N23082, N23066, N4478);
not NOT1 (N23083, N23077);
not NOT1 (N23084, N23076);
or OR4 (N23085, N23073, N6780, N15159, N71);
and AND2 (N23086, N23067, N22585);
nand NAND3 (N23087, N23083, N12759, N9951);
or OR3 (N23088, N23079, N13022, N22657);
and AND4 (N23089, N23088, N20460, N16407, N7400);
or OR3 (N23090, N23075, N17207, N20312);
or OR4 (N23091, N23089, N10573, N14193, N16537);
nand NAND2 (N23092, N23074, N13274);
and AND3 (N23093, N23085, N15702, N11320);
nor NOR3 (N23094, N23081, N10442, N21420);
nand NAND3 (N23095, N23086, N12543, N21043);
nor NOR2 (N23096, N23094, N14422);
xor XOR2 (N23097, N23091, N14279);
and AND3 (N23098, N23093, N10334, N4234);
buf BUF1 (N23099, N23097);
xor XOR2 (N23100, N23090, N3629);
buf BUF1 (N23101, N23080);
not NOT1 (N23102, N23082);
not NOT1 (N23103, N23100);
buf BUF1 (N23104, N23103);
and AND2 (N23105, N23102, N1394);
buf BUF1 (N23106, N23087);
nand NAND3 (N23107, N23101, N9248, N19266);
nand NAND3 (N23108, N23096, N2563, N2259);
nor NOR2 (N23109, N23104, N11148);
xor XOR2 (N23110, N23098, N22311);
or OR3 (N23111, N23099, N20973, N6014);
xor XOR2 (N23112, N23108, N22223);
and AND2 (N23113, N23110, N2849);
buf BUF1 (N23114, N23111);
and AND2 (N23115, N23092, N17815);
nand NAND3 (N23116, N23095, N11488, N16975);
nand NAND4 (N23117, N23107, N9971, N14359, N7279);
not NOT1 (N23118, N23113);
buf BUF1 (N23119, N23118);
not NOT1 (N23120, N23114);
nor NOR3 (N23121, N23119, N15497, N599);
xor XOR2 (N23122, N23106, N22401);
and AND3 (N23123, N23109, N4407, N19931);
buf BUF1 (N23124, N23115);
buf BUF1 (N23125, N23105);
or OR4 (N23126, N23116, N20776, N13172, N8015);
not NOT1 (N23127, N23126);
nor NOR4 (N23128, N23127, N9667, N13509, N10675);
nor NOR2 (N23129, N23122, N12390);
nand NAND4 (N23130, N23084, N21212, N7323, N16194);
and AND4 (N23131, N23117, N8728, N19491, N13155);
nor NOR3 (N23132, N23124, N3398, N14396);
xor XOR2 (N23133, N23130, N16417);
xor XOR2 (N23134, N23128, N2250);
or OR2 (N23135, N23129, N1213);
nor NOR2 (N23136, N23121, N19845);
nand NAND2 (N23137, N23135, N562);
buf BUF1 (N23138, N23133);
nand NAND2 (N23139, N23138, N9512);
or OR3 (N23140, N23123, N8261, N21060);
or OR2 (N23141, N23120, N20898);
buf BUF1 (N23142, N23132);
not NOT1 (N23143, N23139);
buf BUF1 (N23144, N23141);
nor NOR2 (N23145, N23144, N5365);
or OR3 (N23146, N23145, N18658, N15026);
not NOT1 (N23147, N23137);
and AND4 (N23148, N23125, N6091, N6124, N12637);
buf BUF1 (N23149, N23112);
xor XOR2 (N23150, N23146, N9111);
nor NOR4 (N23151, N23142, N7703, N12272, N13866);
nand NAND3 (N23152, N23134, N8916, N5848);
nand NAND4 (N23153, N23147, N14086, N21524, N19436);
and AND4 (N23154, N23140, N15238, N7934, N16209);
nor NOR2 (N23155, N23154, N16373);
and AND2 (N23156, N23151, N4759);
and AND2 (N23157, N23152, N15412);
xor XOR2 (N23158, N23157, N15858);
or OR2 (N23159, N23150, N22209);
not NOT1 (N23160, N23155);
xor XOR2 (N23161, N23131, N7237);
nor NOR2 (N23162, N23158, N19095);
or OR2 (N23163, N23148, N11481);
xor XOR2 (N23164, N23159, N3550);
buf BUF1 (N23165, N23136);
not NOT1 (N23166, N23161);
buf BUF1 (N23167, N23166);
and AND3 (N23168, N23167, N13093, N3743);
buf BUF1 (N23169, N23165);
buf BUF1 (N23170, N23160);
xor XOR2 (N23171, N23164, N375);
not NOT1 (N23172, N23168);
and AND3 (N23173, N23149, N12420, N19265);
buf BUF1 (N23174, N23169);
or OR3 (N23175, N23143, N23065, N11639);
xor XOR2 (N23176, N23172, N16377);
and AND2 (N23177, N23162, N15606);
and AND3 (N23178, N23171, N5217, N20483);
xor XOR2 (N23179, N23178, N21510);
xor XOR2 (N23180, N23163, N9350);
nand NAND2 (N23181, N23156, N7035);
buf BUF1 (N23182, N23175);
xor XOR2 (N23183, N23180, N17008);
nand NAND3 (N23184, N23176, N5861, N16381);
nor NOR4 (N23185, N23179, N21506, N21853, N21532);
nor NOR2 (N23186, N23185, N21976);
and AND3 (N23187, N23174, N15615, N15292);
nand NAND3 (N23188, N23183, N22226, N355);
not NOT1 (N23189, N23177);
nand NAND4 (N23190, N23170, N5636, N3552, N4820);
nor NOR3 (N23191, N23186, N20076, N5632);
and AND4 (N23192, N23181, N20200, N5167, N15922);
xor XOR2 (N23193, N23189, N19803);
xor XOR2 (N23194, N23153, N51);
nand NAND4 (N23195, N23187, N14292, N117, N4864);
buf BUF1 (N23196, N23184);
xor XOR2 (N23197, N23192, N19900);
not NOT1 (N23198, N23182);
xor XOR2 (N23199, N23198, N18649);
nand NAND2 (N23200, N23196, N20223);
or OR4 (N23201, N23190, N11736, N2179, N13485);
and AND4 (N23202, N23193, N7701, N15427, N5352);
nor NOR3 (N23203, N23191, N7041, N5377);
and AND3 (N23204, N23173, N21241, N3418);
not NOT1 (N23205, N23194);
or OR2 (N23206, N23205, N15145);
xor XOR2 (N23207, N23204, N10601);
nand NAND4 (N23208, N23197, N12478, N437, N8344);
and AND2 (N23209, N23207, N15966);
xor XOR2 (N23210, N23206, N16592);
not NOT1 (N23211, N23202);
and AND3 (N23212, N23201, N22102, N13691);
and AND2 (N23213, N23210, N8403);
nand NAND4 (N23214, N23211, N10795, N20082, N21687);
nand NAND2 (N23215, N23199, N15805);
nand NAND4 (N23216, N23200, N19431, N21277, N14466);
buf BUF1 (N23217, N23213);
and AND4 (N23218, N23216, N23107, N1741, N1982);
or OR3 (N23219, N23217, N18241, N14453);
not NOT1 (N23220, N23208);
or OR2 (N23221, N23203, N10106);
not NOT1 (N23222, N23221);
not NOT1 (N23223, N23212);
buf BUF1 (N23224, N23220);
nor NOR2 (N23225, N23214, N19336);
nor NOR2 (N23226, N23222, N6209);
nor NOR2 (N23227, N23215, N12291);
buf BUF1 (N23228, N23218);
nand NAND4 (N23229, N23219, N11801, N22124, N16235);
or OR4 (N23230, N23226, N17724, N908, N20817);
and AND2 (N23231, N23230, N2261);
not NOT1 (N23232, N23223);
nand NAND2 (N23233, N23225, N6428);
nand NAND2 (N23234, N23232, N10495);
xor XOR2 (N23235, N23231, N7646);
not NOT1 (N23236, N23227);
nand NAND3 (N23237, N23235, N3029, N19359);
or OR4 (N23238, N23195, N10496, N9192, N18572);
or OR4 (N23239, N23188, N5598, N9486, N5361);
not NOT1 (N23240, N23228);
nor NOR4 (N23241, N23234, N11977, N5085, N14493);
nor NOR4 (N23242, N23239, N3399, N9889, N26);
nor NOR3 (N23243, N23224, N22628, N7247);
or OR2 (N23244, N23238, N15017);
and AND2 (N23245, N23242, N14585);
xor XOR2 (N23246, N23236, N8119);
nor NOR4 (N23247, N23246, N15794, N615, N3701);
not NOT1 (N23248, N23245);
buf BUF1 (N23249, N23229);
nor NOR2 (N23250, N23249, N11953);
not NOT1 (N23251, N23237);
xor XOR2 (N23252, N23241, N6384);
not NOT1 (N23253, N23244);
and AND4 (N23254, N23250, N2391, N71, N10095);
buf BUF1 (N23255, N23251);
nor NOR2 (N23256, N23255, N12980);
buf BUF1 (N23257, N23233);
not NOT1 (N23258, N23252);
or OR4 (N23259, N23248, N7738, N16553, N22627);
buf BUF1 (N23260, N23254);
not NOT1 (N23261, N23253);
xor XOR2 (N23262, N23257, N12845);
nand NAND3 (N23263, N23262, N22566, N8985);
not NOT1 (N23264, N23247);
or OR2 (N23265, N23209, N11387);
xor XOR2 (N23266, N23258, N19262);
not NOT1 (N23267, N23264);
nand NAND4 (N23268, N23266, N3752, N888, N1606);
not NOT1 (N23269, N23265);
not NOT1 (N23270, N23240);
buf BUF1 (N23271, N23268);
or OR2 (N23272, N23267, N23078);
xor XOR2 (N23273, N23270, N20519);
nand NAND2 (N23274, N23269, N13532);
not NOT1 (N23275, N23243);
or OR3 (N23276, N23271, N2587, N21891);
nand NAND2 (N23277, N23260, N4679);
xor XOR2 (N23278, N23256, N7708);
buf BUF1 (N23279, N23276);
nand NAND2 (N23280, N23261, N14590);
buf BUF1 (N23281, N23278);
nor NOR3 (N23282, N23274, N8898, N14686);
not NOT1 (N23283, N23273);
buf BUF1 (N23284, N23272);
nand NAND3 (N23285, N23259, N4893, N20610);
or OR3 (N23286, N23281, N22456, N18219);
xor XOR2 (N23287, N23280, N16569);
nand NAND4 (N23288, N23286, N4917, N9948, N1130);
buf BUF1 (N23289, N23263);
not NOT1 (N23290, N23289);
buf BUF1 (N23291, N23283);
buf BUF1 (N23292, N23279);
or OR2 (N23293, N23291, N2840);
or OR3 (N23294, N23275, N14221, N15217);
nor NOR4 (N23295, N23293, N2015, N11496, N8223);
xor XOR2 (N23296, N23290, N9188);
or OR3 (N23297, N23292, N987, N13101);
or OR4 (N23298, N23296, N11119, N6917, N5999);
nand NAND3 (N23299, N23294, N14412, N9088);
nor NOR3 (N23300, N23285, N15385, N15319);
xor XOR2 (N23301, N23284, N14487);
not NOT1 (N23302, N23287);
xor XOR2 (N23303, N23277, N20261);
buf BUF1 (N23304, N23302);
not NOT1 (N23305, N23301);
buf BUF1 (N23306, N23299);
not NOT1 (N23307, N23300);
xor XOR2 (N23308, N23304, N13174);
and AND2 (N23309, N23297, N6743);
nor NOR3 (N23310, N23305, N7932, N20415);
nand NAND2 (N23311, N23306, N16919);
buf BUF1 (N23312, N23309);
or OR2 (N23313, N23310, N2900);
buf BUF1 (N23314, N23288);
buf BUF1 (N23315, N23312);
or OR3 (N23316, N23313, N15088, N13848);
xor XOR2 (N23317, N23308, N14986);
nor NOR4 (N23318, N23282, N12535, N6679, N1230);
nor NOR3 (N23319, N23315, N18256, N22025);
nand NAND3 (N23320, N23307, N13566, N21183);
nor NOR3 (N23321, N23314, N2428, N15100);
and AND4 (N23322, N23319, N18919, N12859, N12276);
not NOT1 (N23323, N23316);
nor NOR2 (N23324, N23311, N21646);
or OR2 (N23325, N23295, N11059);
and AND2 (N23326, N23298, N14785);
or OR3 (N23327, N23303, N9071, N7190);
not NOT1 (N23328, N23323);
nand NAND4 (N23329, N23325, N15894, N12679, N12363);
and AND3 (N23330, N23318, N10631, N4469);
nor NOR3 (N23331, N23329, N20003, N15878);
not NOT1 (N23332, N23317);
and AND4 (N23333, N23332, N11192, N6244, N18500);
xor XOR2 (N23334, N23331, N7803);
or OR2 (N23335, N23326, N12696);
nor NOR2 (N23336, N23334, N14239);
xor XOR2 (N23337, N23335, N544);
or OR2 (N23338, N23322, N14344);
and AND3 (N23339, N23324, N7121, N22075);
or OR3 (N23340, N23333, N3664, N2385);
nand NAND3 (N23341, N23321, N21090, N16046);
nand NAND4 (N23342, N23320, N2, N13, N11663);
and AND3 (N23343, N23337, N4253, N7206);
buf BUF1 (N23344, N23328);
xor XOR2 (N23345, N23342, N22589);
not NOT1 (N23346, N23341);
not NOT1 (N23347, N23340);
buf BUF1 (N23348, N23327);
nor NOR4 (N23349, N23344, N13661, N21157, N12420);
nand NAND4 (N23350, N23336, N601, N20993, N8291);
and AND4 (N23351, N23338, N7488, N1580, N9159);
nor NOR4 (N23352, N23348, N3847, N4743, N20543);
nand NAND4 (N23353, N23339, N21242, N22801, N8786);
nor NOR2 (N23354, N23347, N15626);
nand NAND3 (N23355, N23352, N2289, N9842);
or OR2 (N23356, N23346, N6485);
or OR4 (N23357, N23343, N12225, N15452, N12906);
or OR4 (N23358, N23356, N5417, N7839, N4576);
buf BUF1 (N23359, N23351);
xor XOR2 (N23360, N23354, N12262);
nand NAND3 (N23361, N23330, N15945, N17037);
and AND3 (N23362, N23353, N18004, N7132);
nor NOR2 (N23363, N23349, N1839);
xor XOR2 (N23364, N23345, N295);
nor NOR4 (N23365, N23355, N6474, N13989, N682);
xor XOR2 (N23366, N23360, N4050);
and AND2 (N23367, N23357, N20850);
xor XOR2 (N23368, N23367, N10519);
nor NOR4 (N23369, N23358, N2436, N8541, N155);
nor NOR4 (N23370, N23366, N19162, N3472, N12079);
or OR3 (N23371, N23363, N17403, N15133);
nor NOR3 (N23372, N23368, N13757, N14030);
not NOT1 (N23373, N23362);
xor XOR2 (N23374, N23350, N22982);
not NOT1 (N23375, N23374);
nand NAND3 (N23376, N23365, N14668, N20790);
nand NAND2 (N23377, N23359, N9562);
xor XOR2 (N23378, N23370, N8819);
not NOT1 (N23379, N23377);
nand NAND3 (N23380, N23361, N12210, N3793);
or OR4 (N23381, N23372, N11977, N15881, N11001);
not NOT1 (N23382, N23378);
or OR3 (N23383, N23371, N22815, N19615);
not NOT1 (N23384, N23375);
nor NOR2 (N23385, N23380, N19854);
buf BUF1 (N23386, N23381);
and AND4 (N23387, N23364, N17408, N8775, N6753);
nor NOR3 (N23388, N23386, N22778, N19931);
buf BUF1 (N23389, N23387);
xor XOR2 (N23390, N23382, N21949);
nor NOR3 (N23391, N23390, N13731, N289);
buf BUF1 (N23392, N23385);
not NOT1 (N23393, N23379);
nor NOR4 (N23394, N23376, N16124, N4555, N14029);
xor XOR2 (N23395, N23388, N12650);
or OR3 (N23396, N23389, N11477, N2686);
buf BUF1 (N23397, N23395);
buf BUF1 (N23398, N23373);
nand NAND4 (N23399, N23393, N22286, N20948, N9645);
nor NOR4 (N23400, N23396, N9875, N19044, N22116);
buf BUF1 (N23401, N23369);
not NOT1 (N23402, N23398);
buf BUF1 (N23403, N23401);
nor NOR3 (N23404, N23397, N3489, N1660);
buf BUF1 (N23405, N23383);
buf BUF1 (N23406, N23391);
not NOT1 (N23407, N23384);
xor XOR2 (N23408, N23404, N16145);
buf BUF1 (N23409, N23408);
nand NAND2 (N23410, N23399, N10787);
not NOT1 (N23411, N23405);
not NOT1 (N23412, N23402);
nand NAND4 (N23413, N23406, N6850, N305, N1030);
buf BUF1 (N23414, N23409);
xor XOR2 (N23415, N23410, N248);
nor NOR4 (N23416, N23413, N15554, N16501, N6842);
and AND2 (N23417, N23403, N12495);
xor XOR2 (N23418, N23407, N13418);
buf BUF1 (N23419, N23392);
nor NOR4 (N23420, N23415, N19573, N18038, N20782);
buf BUF1 (N23421, N23400);
nand NAND2 (N23422, N23394, N12832);
nor NOR3 (N23423, N23422, N1438, N4290);
buf BUF1 (N23424, N23423);
nor NOR2 (N23425, N23420, N21191);
or OR2 (N23426, N23424, N11629);
buf BUF1 (N23427, N23426);
xor XOR2 (N23428, N23412, N1489);
xor XOR2 (N23429, N23414, N14688);
or OR3 (N23430, N23411, N1174, N11004);
or OR2 (N23431, N23419, N10919);
and AND3 (N23432, N23421, N1535, N14552);
nor NOR3 (N23433, N23432, N22117, N8073);
or OR3 (N23434, N23427, N9887, N6455);
nand NAND3 (N23435, N23430, N19189, N20481);
or OR3 (N23436, N23431, N5874, N18411);
nor NOR4 (N23437, N23417, N2983, N7106, N1717);
not NOT1 (N23438, N23436);
not NOT1 (N23439, N23418);
buf BUF1 (N23440, N23435);
xor XOR2 (N23441, N23428, N14800);
nand NAND4 (N23442, N23433, N6789, N12674, N3292);
nand NAND4 (N23443, N23438, N3652, N10774, N22188);
and AND4 (N23444, N23442, N931, N19806, N12912);
xor XOR2 (N23445, N23439, N22556);
xor XOR2 (N23446, N23443, N7339);
xor XOR2 (N23447, N23425, N22143);
and AND2 (N23448, N23437, N4603);
nand NAND4 (N23449, N23446, N13736, N9567, N7286);
or OR4 (N23450, N23416, N2902, N22130, N5952);
not NOT1 (N23451, N23450);
not NOT1 (N23452, N23445);
and AND3 (N23453, N23447, N19111, N11021);
buf BUF1 (N23454, N23449);
not NOT1 (N23455, N23454);
xor XOR2 (N23456, N23451, N11432);
xor XOR2 (N23457, N23440, N22324);
nand NAND4 (N23458, N23456, N5876, N5019, N6556);
buf BUF1 (N23459, N23444);
xor XOR2 (N23460, N23458, N3515);
not NOT1 (N23461, N23460);
buf BUF1 (N23462, N23457);
buf BUF1 (N23463, N23459);
xor XOR2 (N23464, N23448, N18623);
not NOT1 (N23465, N23453);
not NOT1 (N23466, N23455);
nor NOR3 (N23467, N23452, N6780, N21883);
or OR2 (N23468, N23463, N16234);
buf BUF1 (N23469, N23441);
nor NOR3 (N23470, N23429, N23336, N7039);
xor XOR2 (N23471, N23470, N10714);
not NOT1 (N23472, N23471);
not NOT1 (N23473, N23462);
not NOT1 (N23474, N23468);
buf BUF1 (N23475, N23473);
not NOT1 (N23476, N23465);
buf BUF1 (N23477, N23467);
not NOT1 (N23478, N23472);
or OR4 (N23479, N23464, N20887, N15566, N21563);
nand NAND3 (N23480, N23475, N16045, N23288);
nor NOR3 (N23481, N23478, N11576, N8688);
or OR4 (N23482, N23479, N5377, N23298, N1072);
and AND4 (N23483, N23477, N10950, N23375, N12307);
not NOT1 (N23484, N23483);
buf BUF1 (N23485, N23484);
nand NAND3 (N23486, N23482, N2230, N10774);
or OR4 (N23487, N23486, N15536, N6600, N7680);
or OR4 (N23488, N23480, N8574, N23412, N12409);
or OR2 (N23489, N23481, N13487);
nand NAND3 (N23490, N23469, N16766, N4914);
and AND3 (N23491, N23476, N18594, N13509);
nand NAND2 (N23492, N23474, N14048);
buf BUF1 (N23493, N23492);
and AND3 (N23494, N23491, N21684, N1537);
xor XOR2 (N23495, N23489, N21461);
nand NAND4 (N23496, N23490, N8571, N21194, N7352);
xor XOR2 (N23497, N23495, N9332);
xor XOR2 (N23498, N23493, N3627);
nand NAND2 (N23499, N23434, N8529);
not NOT1 (N23500, N23485);
xor XOR2 (N23501, N23498, N7188);
buf BUF1 (N23502, N23461);
or OR4 (N23503, N23494, N9985, N2276, N17886);
nor NOR3 (N23504, N23488, N19127, N12144);
not NOT1 (N23505, N23497);
nand NAND2 (N23506, N23505, N1487);
nor NOR3 (N23507, N23506, N20518, N731);
nor NOR3 (N23508, N23504, N20372, N6857);
not NOT1 (N23509, N23508);
and AND4 (N23510, N23496, N8572, N20859, N6725);
buf BUF1 (N23511, N23466);
and AND4 (N23512, N23500, N7475, N19601, N10561);
nand NAND4 (N23513, N23510, N8185, N21056, N20437);
nand NAND4 (N23514, N23501, N16962, N9787, N7295);
and AND3 (N23515, N23503, N11955, N11106);
and AND2 (N23516, N23502, N14144);
buf BUF1 (N23517, N23487);
nand NAND4 (N23518, N23517, N14122, N3889, N9292);
not NOT1 (N23519, N23507);
buf BUF1 (N23520, N23515);
xor XOR2 (N23521, N23520, N17001);
nor NOR4 (N23522, N23518, N7079, N4996, N15777);
nor NOR4 (N23523, N23521, N15373, N9058, N2661);
not NOT1 (N23524, N23514);
and AND3 (N23525, N23519, N10830, N1885);
xor XOR2 (N23526, N23524, N8396);
nor NOR3 (N23527, N23522, N10874, N22764);
nor NOR4 (N23528, N23511, N7804, N9252, N9993);
not NOT1 (N23529, N23516);
and AND2 (N23530, N23523, N18478);
not NOT1 (N23531, N23526);
xor XOR2 (N23532, N23499, N8750);
or OR4 (N23533, N23532, N22680, N2303, N15897);
nor NOR2 (N23534, N23528, N21476);
nand NAND3 (N23535, N23513, N22969, N20196);
xor XOR2 (N23536, N23533, N12572);
nand NAND2 (N23537, N23525, N6494);
and AND3 (N23538, N23534, N4042, N18647);
not NOT1 (N23539, N23509);
nand NAND2 (N23540, N23529, N17795);
not NOT1 (N23541, N23538);
not NOT1 (N23542, N23541);
and AND3 (N23543, N23512, N2624, N13777);
nor NOR3 (N23544, N23535, N8986, N17372);
not NOT1 (N23545, N23544);
nand NAND3 (N23546, N23536, N13691, N19182);
or OR3 (N23547, N23531, N15090, N1120);
nand NAND2 (N23548, N23527, N6989);
nand NAND3 (N23549, N23542, N12343, N19833);
buf BUF1 (N23550, N23548);
and AND3 (N23551, N23549, N8064, N19517);
buf BUF1 (N23552, N23546);
nor NOR2 (N23553, N23539, N17845);
nand NAND3 (N23554, N23553, N21023, N16736);
not NOT1 (N23555, N23537);
nor NOR2 (N23556, N23550, N19881);
nand NAND2 (N23557, N23530, N2846);
nand NAND3 (N23558, N23543, N71, N16504);
not NOT1 (N23559, N23555);
nand NAND4 (N23560, N23556, N14508, N10030, N4877);
xor XOR2 (N23561, N23547, N3466);
buf BUF1 (N23562, N23560);
nand NAND2 (N23563, N23540, N22615);
nor NOR4 (N23564, N23552, N5697, N20763, N5669);
buf BUF1 (N23565, N23554);
and AND2 (N23566, N23561, N12359);
xor XOR2 (N23567, N23562, N10536);
xor XOR2 (N23568, N23557, N5161);
xor XOR2 (N23569, N23551, N2645);
nor NOR4 (N23570, N23569, N5884, N5715, N14312);
or OR4 (N23571, N23565, N22951, N16891, N19189);
nor NOR4 (N23572, N23558, N11523, N20556, N20227);
nor NOR2 (N23573, N23570, N2318);
and AND3 (N23574, N23545, N1856, N5287);
xor XOR2 (N23575, N23566, N225);
buf BUF1 (N23576, N23559);
nand NAND3 (N23577, N23575, N18660, N23008);
nand NAND4 (N23578, N23564, N21294, N22237, N13979);
nand NAND3 (N23579, N23577, N12457, N8521);
and AND4 (N23580, N23578, N2688, N833, N119);
or OR3 (N23581, N23571, N12890, N15472);
and AND4 (N23582, N23579, N20654, N11545, N10797);
or OR4 (N23583, N23582, N5366, N7268, N22969);
nand NAND2 (N23584, N23567, N16443);
and AND2 (N23585, N23576, N12260);
not NOT1 (N23586, N23581);
xor XOR2 (N23587, N23584, N20412);
nand NAND2 (N23588, N23563, N16840);
buf BUF1 (N23589, N23574);
nor NOR3 (N23590, N23588, N17611, N16356);
or OR4 (N23591, N23585, N23406, N22300, N7604);
nor NOR3 (N23592, N23590, N7190, N12681);
or OR3 (N23593, N23573, N4324, N8818);
nor NOR4 (N23594, N23592, N13772, N12807, N7867);
buf BUF1 (N23595, N23583);
or OR4 (N23596, N23568, N8988, N10360, N14866);
buf BUF1 (N23597, N23595);
or OR2 (N23598, N23596, N21274);
buf BUF1 (N23599, N23587);
or OR2 (N23600, N23598, N10910);
buf BUF1 (N23601, N23589);
and AND3 (N23602, N23586, N22041, N4565);
or OR2 (N23603, N23602, N10980);
nor NOR2 (N23604, N23593, N15163);
and AND4 (N23605, N23572, N17844, N20992, N5233);
xor XOR2 (N23606, N23604, N3951);
and AND4 (N23607, N23597, N18133, N16740, N4580);
nand NAND3 (N23608, N23603, N17269, N9009);
not NOT1 (N23609, N23594);
not NOT1 (N23610, N23601);
nand NAND2 (N23611, N23606, N2218);
buf BUF1 (N23612, N23611);
or OR4 (N23613, N23599, N10165, N7160, N6162);
xor XOR2 (N23614, N23609, N13460);
and AND2 (N23615, N23605, N11535);
buf BUF1 (N23616, N23614);
xor XOR2 (N23617, N23580, N17945);
or OR4 (N23618, N23615, N21230, N14283, N7937);
and AND2 (N23619, N23610, N5557);
xor XOR2 (N23620, N23618, N14528);
not NOT1 (N23621, N23600);
nand NAND4 (N23622, N23617, N2201, N11396, N19837);
nand NAND3 (N23623, N23608, N11211, N12757);
or OR2 (N23624, N23619, N10087);
not NOT1 (N23625, N23622);
or OR4 (N23626, N23621, N1345, N3154, N15615);
xor XOR2 (N23627, N23620, N13137);
nand NAND2 (N23628, N23625, N12409);
xor XOR2 (N23629, N23623, N8121);
not NOT1 (N23630, N23624);
nand NAND3 (N23631, N23607, N9484, N21507);
buf BUF1 (N23632, N23612);
or OR2 (N23633, N23591, N9175);
nor NOR3 (N23634, N23631, N12126, N21628);
or OR3 (N23635, N23632, N9326, N21446);
or OR3 (N23636, N23613, N2861, N19837);
nand NAND2 (N23637, N23628, N13926);
not NOT1 (N23638, N23636);
nand NAND3 (N23639, N23629, N15073, N22590);
nand NAND2 (N23640, N23627, N5873);
or OR2 (N23641, N23640, N14030);
xor XOR2 (N23642, N23635, N20342);
not NOT1 (N23643, N23638);
xor XOR2 (N23644, N23641, N19688);
buf BUF1 (N23645, N23633);
buf BUF1 (N23646, N23645);
nand NAND4 (N23647, N23630, N11669, N16980, N2664);
or OR2 (N23648, N23626, N7546);
nor NOR3 (N23649, N23639, N17246, N3106);
or OR3 (N23650, N23648, N15154, N8241);
or OR3 (N23651, N23646, N22053, N6704);
nor NOR4 (N23652, N23637, N14396, N23461, N22296);
buf BUF1 (N23653, N23634);
buf BUF1 (N23654, N23650);
and AND3 (N23655, N23616, N13302, N21882);
buf BUF1 (N23656, N23647);
nand NAND3 (N23657, N23643, N11487, N23530);
or OR4 (N23658, N23642, N1873, N17269, N5425);
and AND4 (N23659, N23649, N14824, N3436, N15297);
not NOT1 (N23660, N23656);
xor XOR2 (N23661, N23658, N21486);
or OR2 (N23662, N23661, N17716);
buf BUF1 (N23663, N23655);
xor XOR2 (N23664, N23644, N6030);
xor XOR2 (N23665, N23664, N13180);
nand NAND3 (N23666, N23657, N12011, N10294);
buf BUF1 (N23667, N23665);
or OR3 (N23668, N23651, N12656, N281);
not NOT1 (N23669, N23662);
and AND2 (N23670, N23663, N19352);
not NOT1 (N23671, N23670);
buf BUF1 (N23672, N23652);
nor NOR4 (N23673, N23668, N7526, N18168, N18335);
nand NAND3 (N23674, N23660, N2059, N20151);
buf BUF1 (N23675, N23673);
nand NAND2 (N23676, N23672, N454);
nor NOR3 (N23677, N23674, N16314, N18216);
xor XOR2 (N23678, N23675, N8683);
nand NAND3 (N23679, N23671, N9481, N18983);
buf BUF1 (N23680, N23659);
nand NAND2 (N23681, N23679, N9270);
and AND3 (N23682, N23676, N6270, N18351);
xor XOR2 (N23683, N23666, N21184);
buf BUF1 (N23684, N23654);
or OR4 (N23685, N23678, N22985, N7540, N8299);
xor XOR2 (N23686, N23667, N19753);
nand NAND2 (N23687, N23669, N17617);
buf BUF1 (N23688, N23653);
not NOT1 (N23689, N23684);
buf BUF1 (N23690, N23685);
and AND4 (N23691, N23690, N20542, N4243, N4129);
nand NAND4 (N23692, N23686, N19604, N1486, N16119);
not NOT1 (N23693, N23682);
buf BUF1 (N23694, N23687);
xor XOR2 (N23695, N23691, N21428);
not NOT1 (N23696, N23695);
buf BUF1 (N23697, N23696);
nor NOR2 (N23698, N23680, N9382);
not NOT1 (N23699, N23698);
nand NAND2 (N23700, N23693, N10794);
not NOT1 (N23701, N23689);
buf BUF1 (N23702, N23697);
nand NAND4 (N23703, N23700, N16427, N20455, N6652);
xor XOR2 (N23704, N23694, N4801);
nand NAND3 (N23705, N23699, N8493, N22543);
buf BUF1 (N23706, N23681);
buf BUF1 (N23707, N23702);
not NOT1 (N23708, N23701);
and AND4 (N23709, N23677, N16446, N15763, N13000);
not NOT1 (N23710, N23705);
not NOT1 (N23711, N23704);
buf BUF1 (N23712, N23692);
or OR2 (N23713, N23688, N9778);
or OR3 (N23714, N23706, N10396, N15057);
xor XOR2 (N23715, N23712, N15462);
nand NAND3 (N23716, N23709, N20503, N23237);
buf BUF1 (N23717, N23716);
or OR3 (N23718, N23717, N14318, N16540);
buf BUF1 (N23719, N23707);
and AND3 (N23720, N23683, N11483, N15803);
buf BUF1 (N23721, N23715);
buf BUF1 (N23722, N23714);
or OR4 (N23723, N23711, N18383, N6832, N11293);
nor NOR2 (N23724, N23721, N19842);
nand NAND2 (N23725, N23718, N3437);
buf BUF1 (N23726, N23723);
or OR3 (N23727, N23708, N21510, N11468);
nand NAND4 (N23728, N23713, N818, N12783, N23540);
not NOT1 (N23729, N23703);
nand NAND4 (N23730, N23729, N15381, N10043, N1351);
or OR4 (N23731, N23710, N4878, N309, N963);
nor NOR4 (N23732, N23730, N7576, N22266, N13719);
buf BUF1 (N23733, N23722);
or OR3 (N23734, N23728, N21156, N14889);
buf BUF1 (N23735, N23727);
nor NOR4 (N23736, N23724, N16664, N21698, N16680);
and AND3 (N23737, N23733, N22330, N15804);
not NOT1 (N23738, N23735);
not NOT1 (N23739, N23725);
or OR4 (N23740, N23737, N4727, N7208, N3127);
nor NOR3 (N23741, N23726, N6737, N20432);
and AND3 (N23742, N23734, N18447, N10108);
or OR4 (N23743, N23738, N14853, N20298, N7984);
nand NAND2 (N23744, N23743, N5448);
nor NOR2 (N23745, N23744, N14804);
buf BUF1 (N23746, N23736);
nand NAND4 (N23747, N23746, N19162, N2970, N14871);
buf BUF1 (N23748, N23741);
nor NOR4 (N23749, N23720, N12283, N16184, N18238);
xor XOR2 (N23750, N23731, N13139);
or OR2 (N23751, N23750, N13958);
and AND3 (N23752, N23749, N19580, N5402);
buf BUF1 (N23753, N23745);
nand NAND2 (N23754, N23739, N8042);
nand NAND4 (N23755, N23740, N2668, N16847, N18512);
nor NOR2 (N23756, N23732, N10640);
xor XOR2 (N23757, N23751, N4001);
xor XOR2 (N23758, N23755, N4053);
or OR2 (N23759, N23747, N9383);
nand NAND3 (N23760, N23758, N20943, N13301);
buf BUF1 (N23761, N23752);
nor NOR3 (N23762, N23754, N604, N18850);
nor NOR2 (N23763, N23756, N20798);
nor NOR3 (N23764, N23760, N11531, N2321);
xor XOR2 (N23765, N23757, N16456);
and AND2 (N23766, N23765, N21487);
nor NOR2 (N23767, N23761, N16446);
buf BUF1 (N23768, N23764);
and AND4 (N23769, N23753, N6614, N4524, N3386);
nor NOR3 (N23770, N23767, N12144, N1512);
and AND2 (N23771, N23763, N16528);
nor NOR3 (N23772, N23762, N19605, N12040);
not NOT1 (N23773, N23769);
nand NAND3 (N23774, N23719, N21629, N17163);
and AND3 (N23775, N23773, N8737, N6378);
nor NOR4 (N23776, N23775, N3261, N539, N14677);
xor XOR2 (N23777, N23768, N7652);
nor NOR2 (N23778, N23774, N15793);
nor NOR2 (N23779, N23772, N22107);
buf BUF1 (N23780, N23776);
nor NOR2 (N23781, N23748, N15787);
or OR4 (N23782, N23766, N15715, N4708, N19494);
nand NAND3 (N23783, N23781, N11138, N17067);
or OR2 (N23784, N23742, N2921);
nor NOR3 (N23785, N23784, N14429, N6899);
nand NAND3 (N23786, N23778, N15421, N12917);
xor XOR2 (N23787, N23779, N4328);
nor NOR2 (N23788, N23759, N1382);
or OR2 (N23789, N23786, N15365);
nor NOR3 (N23790, N23782, N1899, N12992);
and AND3 (N23791, N23789, N3752, N13348);
or OR2 (N23792, N23790, N212);
buf BUF1 (N23793, N23792);
not NOT1 (N23794, N23777);
and AND2 (N23795, N23793, N19242);
buf BUF1 (N23796, N23783);
or OR4 (N23797, N23788, N10756, N16255, N4166);
xor XOR2 (N23798, N23794, N17041);
not NOT1 (N23799, N23770);
xor XOR2 (N23800, N23795, N16055);
nand NAND2 (N23801, N23787, N1723);
nor NOR4 (N23802, N23796, N9213, N2722, N1146);
and AND3 (N23803, N23802, N3942, N21006);
or OR3 (N23804, N23800, N2119, N4182);
and AND2 (N23805, N23799, N17138);
not NOT1 (N23806, N23801);
not NOT1 (N23807, N23785);
not NOT1 (N23808, N23805);
nand NAND3 (N23809, N23806, N17796, N11596);
not NOT1 (N23810, N23803);
buf BUF1 (N23811, N23804);
and AND2 (N23812, N23780, N22555);
not NOT1 (N23813, N23810);
nor NOR2 (N23814, N23791, N23069);
or OR2 (N23815, N23811, N2049);
xor XOR2 (N23816, N23808, N8781);
xor XOR2 (N23817, N23812, N10316);
or OR3 (N23818, N23815, N11993, N1801);
not NOT1 (N23819, N23814);
buf BUF1 (N23820, N23818);
not NOT1 (N23821, N23817);
xor XOR2 (N23822, N23813, N2657);
buf BUF1 (N23823, N23816);
buf BUF1 (N23824, N23821);
nor NOR2 (N23825, N23823, N2558);
and AND3 (N23826, N23822, N9860, N19670);
nand NAND2 (N23827, N23797, N8555);
or OR3 (N23828, N23809, N17942, N18543);
xor XOR2 (N23829, N23826, N13314);
and AND2 (N23830, N23825, N18178);
xor XOR2 (N23831, N23807, N13603);
or OR3 (N23832, N23798, N16459, N1306);
nand NAND3 (N23833, N23820, N16191, N7354);
nor NOR2 (N23834, N23819, N16485);
buf BUF1 (N23835, N23833);
xor XOR2 (N23836, N23828, N14487);
or OR4 (N23837, N23835, N15955, N12544, N23544);
not NOT1 (N23838, N23837);
nand NAND3 (N23839, N23824, N8679, N20405);
buf BUF1 (N23840, N23839);
or OR2 (N23841, N23838, N5543);
xor XOR2 (N23842, N23841, N12200);
nand NAND3 (N23843, N23831, N1857, N3295);
and AND2 (N23844, N23836, N10442);
or OR4 (N23845, N23832, N2426, N20793, N8665);
and AND3 (N23846, N23829, N20825, N6914);
buf BUF1 (N23847, N23843);
or OR2 (N23848, N23847, N21668);
and AND2 (N23849, N23846, N7525);
nand NAND3 (N23850, N23834, N4061, N3506);
buf BUF1 (N23851, N23771);
nand NAND2 (N23852, N23849, N13643);
or OR2 (N23853, N23840, N7779);
and AND3 (N23854, N23842, N3654, N1456);
nor NOR2 (N23855, N23827, N21284);
xor XOR2 (N23856, N23851, N12222);
buf BUF1 (N23857, N23853);
or OR3 (N23858, N23844, N9188, N6906);
not NOT1 (N23859, N23848);
or OR2 (N23860, N23858, N10478);
nor NOR4 (N23861, N23859, N17187, N21911, N19006);
buf BUF1 (N23862, N23850);
buf BUF1 (N23863, N23856);
xor XOR2 (N23864, N23857, N1773);
not NOT1 (N23865, N23855);
nor NOR4 (N23866, N23862, N23474, N12333, N1661);
xor XOR2 (N23867, N23854, N4188);
xor XOR2 (N23868, N23860, N23867);
nand NAND4 (N23869, N2883, N20186, N3587, N11907);
not NOT1 (N23870, N23863);
or OR4 (N23871, N23864, N16557, N7102, N5735);
not NOT1 (N23872, N23866);
nand NAND2 (N23873, N23865, N22584);
and AND4 (N23874, N23852, N8673, N9928, N18209);
buf BUF1 (N23875, N23830);
or OR3 (N23876, N23869, N20164, N18958);
xor XOR2 (N23877, N23861, N17939);
nand NAND2 (N23878, N23870, N12341);
xor XOR2 (N23879, N23875, N10340);
nand NAND4 (N23880, N23871, N9873, N17795, N712);
not NOT1 (N23881, N23872);
nor NOR2 (N23882, N23878, N5564);
nand NAND3 (N23883, N23881, N3034, N6864);
nand NAND2 (N23884, N23845, N10621);
nor NOR2 (N23885, N23876, N14837);
nand NAND3 (N23886, N23884, N11368, N9463);
xor XOR2 (N23887, N23886, N5006);
xor XOR2 (N23888, N23882, N11166);
or OR2 (N23889, N23887, N4057);
nor NOR4 (N23890, N23885, N14259, N18971, N14029);
not NOT1 (N23891, N23873);
nand NAND3 (N23892, N23888, N22459, N9199);
and AND3 (N23893, N23883, N21564, N21309);
buf BUF1 (N23894, N23874);
buf BUF1 (N23895, N23879);
not NOT1 (N23896, N23880);
xor XOR2 (N23897, N23893, N12248);
buf BUF1 (N23898, N23892);
not NOT1 (N23899, N23895);
buf BUF1 (N23900, N23890);
or OR4 (N23901, N23897, N10165, N1012, N18265);
or OR4 (N23902, N23889, N13899, N7357, N7032);
not NOT1 (N23903, N23877);
xor XOR2 (N23904, N23896, N18532);
xor XOR2 (N23905, N23901, N17003);
xor XOR2 (N23906, N23868, N12153);
xor XOR2 (N23907, N23900, N1667);
xor XOR2 (N23908, N23891, N6760);
and AND4 (N23909, N23899, N13073, N1439, N20370);
nand NAND2 (N23910, N23903, N22124);
nor NOR3 (N23911, N23898, N7744, N22499);
not NOT1 (N23912, N23911);
and AND2 (N23913, N23908, N1186);
xor XOR2 (N23914, N23904, N22997);
xor XOR2 (N23915, N23914, N12265);
buf BUF1 (N23916, N23915);
nand NAND4 (N23917, N23910, N6826, N13248, N18309);
buf BUF1 (N23918, N23917);
nand NAND2 (N23919, N23894, N11619);
xor XOR2 (N23920, N23916, N2988);
buf BUF1 (N23921, N23909);
or OR3 (N23922, N23921, N14802, N10629);
nand NAND2 (N23923, N23905, N12021);
or OR2 (N23924, N23919, N8424);
xor XOR2 (N23925, N23906, N16342);
nor NOR4 (N23926, N23918, N301, N14786, N22582);
and AND2 (N23927, N23913, N12858);
nor NOR3 (N23928, N23927, N3447, N7212);
not NOT1 (N23929, N23923);
or OR4 (N23930, N23912, N23787, N19088, N6525);
or OR3 (N23931, N23926, N4402, N23909);
nand NAND4 (N23932, N23930, N3544, N1276, N502);
nor NOR3 (N23933, N23928, N20299, N512);
and AND4 (N23934, N23929, N21695, N9459, N2337);
and AND3 (N23935, N23924, N11517, N22576);
or OR2 (N23936, N23922, N20751);
nand NAND3 (N23937, N23931, N11989, N14603);
buf BUF1 (N23938, N23902);
buf BUF1 (N23939, N23934);
not NOT1 (N23940, N23925);
and AND4 (N23941, N23933, N15694, N19385, N11363);
nand NAND4 (N23942, N23941, N18865, N18087, N6894);
not NOT1 (N23943, N23938);
xor XOR2 (N23944, N23937, N425);
nand NAND3 (N23945, N23944, N6300, N11114);
nor NOR2 (N23946, N23935, N16725);
xor XOR2 (N23947, N23920, N19532);
nand NAND2 (N23948, N23936, N16581);
or OR2 (N23949, N23947, N4801);
nand NAND2 (N23950, N23942, N22956);
buf BUF1 (N23951, N23948);
xor XOR2 (N23952, N23932, N7576);
nand NAND3 (N23953, N23940, N10176, N11620);
not NOT1 (N23954, N23943);
nand NAND2 (N23955, N23939, N2534);
xor XOR2 (N23956, N23951, N21861);
xor XOR2 (N23957, N23956, N18162);
not NOT1 (N23958, N23957);
not NOT1 (N23959, N23954);
nand NAND4 (N23960, N23958, N7511, N18996, N3031);
and AND4 (N23961, N23952, N18172, N19443, N23236);
buf BUF1 (N23962, N23959);
nor NOR4 (N23963, N23949, N21441, N18485, N7087);
or OR2 (N23964, N23962, N5421);
buf BUF1 (N23965, N23945);
nand NAND4 (N23966, N23946, N10752, N13135, N13568);
xor XOR2 (N23967, N23907, N12848);
xor XOR2 (N23968, N23961, N5879);
buf BUF1 (N23969, N23965);
or OR2 (N23970, N23963, N18335);
and AND4 (N23971, N23967, N19267, N18381, N15928);
nor NOR2 (N23972, N23964, N1197);
buf BUF1 (N23973, N23960);
nand NAND3 (N23974, N23953, N18644, N3906);
nor NOR4 (N23975, N23970, N11058, N18170, N23071);
nand NAND2 (N23976, N23969, N20984);
buf BUF1 (N23977, N23974);
xor XOR2 (N23978, N23955, N19018);
and AND3 (N23979, N23977, N6308, N14);
nand NAND4 (N23980, N23968, N1283, N16822, N15222);
not NOT1 (N23981, N23950);
buf BUF1 (N23982, N23981);
buf BUF1 (N23983, N23966);
not NOT1 (N23984, N23971);
not NOT1 (N23985, N23973);
not NOT1 (N23986, N23975);
not NOT1 (N23987, N23978);
not NOT1 (N23988, N23976);
buf BUF1 (N23989, N23984);
nand NAND3 (N23990, N23983, N9881, N3891);
nor NOR2 (N23991, N23990, N3151);
or OR2 (N23992, N23982, N5430);
not NOT1 (N23993, N23986);
and AND4 (N23994, N23987, N725, N19859, N23837);
nand NAND4 (N23995, N23989, N1508, N13600, N18212);
xor XOR2 (N23996, N23991, N10137);
and AND2 (N23997, N23985, N17129);
or OR3 (N23998, N23992, N1619, N23445);
buf BUF1 (N23999, N23993);
buf BUF1 (N24000, N23972);
xor XOR2 (N24001, N23995, N3574);
and AND4 (N24002, N23979, N293, N7477, N2770);
and AND4 (N24003, N24001, N4657, N7091, N6882);
xor XOR2 (N24004, N24003, N3189);
nor NOR4 (N24005, N23999, N10287, N9143, N5250);
nor NOR4 (N24006, N23988, N3102, N4893, N9157);
not NOT1 (N24007, N24002);
and AND2 (N24008, N23997, N3710);
nand NAND2 (N24009, N23994, N6317);
buf BUF1 (N24010, N23980);
buf BUF1 (N24011, N24009);
buf BUF1 (N24012, N24007);
nor NOR2 (N24013, N23998, N17880);
buf BUF1 (N24014, N24004);
and AND3 (N24015, N24000, N14481, N72);
and AND4 (N24016, N24012, N20130, N13752, N19379);
and AND3 (N24017, N24005, N17175, N14628);
or OR2 (N24018, N24011, N1738);
xor XOR2 (N24019, N24010, N13631);
nor NOR3 (N24020, N24016, N5807, N7645);
and AND2 (N24021, N24018, N10313);
nand NAND3 (N24022, N24020, N3878, N601);
xor XOR2 (N24023, N24021, N14983);
or OR2 (N24024, N24006, N10269);
xor XOR2 (N24025, N24024, N11004);
or OR2 (N24026, N24019, N11915);
not NOT1 (N24027, N24013);
and AND2 (N24028, N24017, N10002);
nor NOR4 (N24029, N24025, N3174, N426, N18412);
buf BUF1 (N24030, N24027);
buf BUF1 (N24031, N24030);
or OR3 (N24032, N24028, N258, N8184);
buf BUF1 (N24033, N24015);
buf BUF1 (N24034, N24031);
and AND2 (N24035, N24032, N5403);
or OR3 (N24036, N23996, N13255, N8808);
not NOT1 (N24037, N24029);
not NOT1 (N24038, N24034);
nand NAND4 (N24039, N24036, N13730, N4333, N17375);
nor NOR4 (N24040, N24033, N13475, N23582, N12006);
buf BUF1 (N24041, N24038);
xor XOR2 (N24042, N24041, N4547);
xor XOR2 (N24043, N24026, N6006);
nand NAND3 (N24044, N24042, N5563, N16735);
and AND2 (N24045, N24040, N14095);
and AND4 (N24046, N24045, N16229, N19293, N14966);
xor XOR2 (N24047, N24043, N19409);
buf BUF1 (N24048, N24047);
or OR2 (N24049, N24037, N3818);
and AND2 (N24050, N24014, N7339);
nor NOR4 (N24051, N24039, N11128, N22449, N5045);
nor NOR3 (N24052, N24050, N2470, N5578);
or OR2 (N24053, N24023, N19747);
and AND3 (N24054, N24052, N5148, N8976);
not NOT1 (N24055, N24054);
xor XOR2 (N24056, N24053, N11452);
buf BUF1 (N24057, N24044);
or OR2 (N24058, N24056, N5069);
and AND2 (N24059, N24051, N21413);
and AND2 (N24060, N24055, N15993);
nor NOR4 (N24061, N24059, N13234, N12149, N8757);
buf BUF1 (N24062, N24060);
nand NAND2 (N24063, N24046, N22724);
nand NAND3 (N24064, N24063, N613, N20609);
nor NOR2 (N24065, N24049, N12204);
buf BUF1 (N24066, N24022);
buf BUF1 (N24067, N24065);
xor XOR2 (N24068, N24061, N8787);
buf BUF1 (N24069, N24008);
and AND3 (N24070, N24066, N10043, N9195);
nand NAND4 (N24071, N24057, N2074, N13386, N15539);
and AND2 (N24072, N24062, N4050);
not NOT1 (N24073, N24071);
buf BUF1 (N24074, N24058);
buf BUF1 (N24075, N24070);
buf BUF1 (N24076, N24035);
and AND3 (N24077, N24073, N2544, N5080);
not NOT1 (N24078, N24069);
and AND4 (N24079, N24048, N3284, N4770, N24055);
or OR4 (N24080, N24075, N15738, N11598, N18655);
nand NAND3 (N24081, N24072, N3829, N4680);
nand NAND4 (N24082, N24076, N17641, N20286, N11752);
not NOT1 (N24083, N24080);
nand NAND4 (N24084, N24077, N5254, N15883, N16834);
buf BUF1 (N24085, N24078);
and AND3 (N24086, N24067, N11847, N7326);
xor XOR2 (N24087, N24083, N18764);
xor XOR2 (N24088, N24074, N5167);
xor XOR2 (N24089, N24088, N2164);
not NOT1 (N24090, N24068);
xor XOR2 (N24091, N24064, N8704);
and AND2 (N24092, N24091, N20778);
buf BUF1 (N24093, N24089);
and AND3 (N24094, N24081, N9147, N1921);
xor XOR2 (N24095, N24087, N18421);
buf BUF1 (N24096, N24090);
or OR4 (N24097, N24096, N4777, N10770, N19335);
nor NOR2 (N24098, N24095, N9809);
or OR2 (N24099, N24094, N17956);
nand NAND2 (N24100, N24093, N14119);
buf BUF1 (N24101, N24099);
nor NOR4 (N24102, N24084, N10485, N12266, N3099);
or OR4 (N24103, N24082, N13117, N21158, N6715);
or OR2 (N24104, N24098, N3167);
nand NAND3 (N24105, N24079, N3950, N14876);
not NOT1 (N24106, N24105);
nor NOR3 (N24107, N24104, N2950, N21256);
xor XOR2 (N24108, N24100, N9651);
nand NAND3 (N24109, N24097, N18454, N12760);
buf BUF1 (N24110, N24086);
nand NAND2 (N24111, N24102, N6252);
or OR4 (N24112, N24111, N9164, N11057, N23295);
and AND2 (N24113, N24107, N4535);
buf BUF1 (N24114, N24110);
buf BUF1 (N24115, N24085);
or OR2 (N24116, N24103, N23520);
xor XOR2 (N24117, N24115, N20184);
or OR2 (N24118, N24101, N21489);
nand NAND2 (N24119, N24114, N21784);
or OR2 (N24120, N24116, N6163);
and AND4 (N24121, N24109, N3227, N21264, N900);
nand NAND2 (N24122, N24106, N17331);
nor NOR4 (N24123, N24122, N10423, N23647, N18364);
and AND3 (N24124, N24117, N16597, N17080);
and AND2 (N24125, N24123, N8866);
xor XOR2 (N24126, N24118, N23492);
or OR2 (N24127, N24121, N6321);
xor XOR2 (N24128, N24112, N7955);
not NOT1 (N24129, N24127);
not NOT1 (N24130, N24125);
buf BUF1 (N24131, N24119);
or OR4 (N24132, N24092, N10364, N9130, N16717);
nor NOR2 (N24133, N24113, N23474);
nor NOR4 (N24134, N24132, N11435, N12052, N4873);
xor XOR2 (N24135, N24130, N20860);
buf BUF1 (N24136, N24126);
buf BUF1 (N24137, N24129);
buf BUF1 (N24138, N24128);
not NOT1 (N24139, N24134);
buf BUF1 (N24140, N24139);
or OR4 (N24141, N24120, N6222, N11076, N840);
or OR3 (N24142, N24131, N12573, N5745);
not NOT1 (N24143, N24133);
buf BUF1 (N24144, N24124);
or OR2 (N24145, N24140, N11991);
xor XOR2 (N24146, N24137, N15141);
and AND3 (N24147, N24145, N22784, N13563);
or OR4 (N24148, N24143, N3607, N20958, N22623);
nor NOR3 (N24149, N24135, N10928, N7333);
nand NAND2 (N24150, N24141, N3063);
or OR4 (N24151, N24149, N8214, N22535, N18967);
nand NAND3 (N24152, N24146, N21396, N1265);
xor XOR2 (N24153, N24138, N22296);
xor XOR2 (N24154, N24142, N15509);
xor XOR2 (N24155, N24144, N20028);
not NOT1 (N24156, N24147);
nor NOR4 (N24157, N24136, N10863, N14854, N2858);
buf BUF1 (N24158, N24150);
nor NOR4 (N24159, N24158, N19210, N9084, N10385);
or OR2 (N24160, N24108, N19168);
or OR2 (N24161, N24160, N5296);
or OR2 (N24162, N24148, N3759);
buf BUF1 (N24163, N24152);
nor NOR2 (N24164, N24153, N7045);
and AND4 (N24165, N24159, N11714, N2277, N16255);
nor NOR3 (N24166, N24165, N7385, N9827);
xor XOR2 (N24167, N24156, N6498);
buf BUF1 (N24168, N24167);
xor XOR2 (N24169, N24161, N16192);
nor NOR4 (N24170, N24155, N11737, N6787, N17266);
nor NOR2 (N24171, N24163, N9430);
buf BUF1 (N24172, N24164);
xor XOR2 (N24173, N24151, N5585);
and AND4 (N24174, N24169, N18918, N1703, N7649);
buf BUF1 (N24175, N24171);
or OR3 (N24176, N24168, N652, N18895);
nor NOR4 (N24177, N24174, N9529, N23022, N14044);
or OR3 (N24178, N24170, N3727, N3399);
nand NAND3 (N24179, N24178, N4379, N3427);
not NOT1 (N24180, N24162);
nand NAND3 (N24181, N24154, N23025, N20845);
nand NAND4 (N24182, N24181, N21549, N20571, N4602);
and AND2 (N24183, N24166, N18914);
xor XOR2 (N24184, N24157, N19107);
or OR4 (N24185, N24172, N4557, N22646, N13657);
nand NAND2 (N24186, N24179, N2428);
xor XOR2 (N24187, N24173, N16684);
or OR3 (N24188, N24187, N12071, N7213);
xor XOR2 (N24189, N24182, N5028);
and AND4 (N24190, N24184, N802, N12618, N9269);
xor XOR2 (N24191, N24175, N332);
and AND3 (N24192, N24189, N3467, N19130);
and AND4 (N24193, N24183, N7038, N41, N3512);
buf BUF1 (N24194, N24193);
nand NAND2 (N24195, N24188, N19115);
nor NOR3 (N24196, N24191, N5666, N12532);
not NOT1 (N24197, N24194);
nand NAND2 (N24198, N24185, N2916);
nand NAND4 (N24199, N24198, N5747, N19770, N2016);
and AND2 (N24200, N24197, N5647);
or OR2 (N24201, N24176, N19858);
buf BUF1 (N24202, N24177);
or OR3 (N24203, N24180, N19703, N12338);
or OR2 (N24204, N24203, N6300);
buf BUF1 (N24205, N24195);
nand NAND2 (N24206, N24205, N23652);
nor NOR4 (N24207, N24186, N17306, N18263, N21424);
or OR3 (N24208, N24204, N13352, N16739);
nor NOR3 (N24209, N24207, N19385, N8233);
nand NAND2 (N24210, N24190, N16517);
xor XOR2 (N24211, N24202, N17760);
or OR4 (N24212, N24196, N13532, N23540, N7045);
nor NOR4 (N24213, N24212, N9908, N17740, N2876);
not NOT1 (N24214, N24209);
nand NAND3 (N24215, N24201, N17212, N11965);
and AND2 (N24216, N24211, N16339);
nor NOR4 (N24217, N24206, N13991, N4087, N503);
and AND3 (N24218, N24215, N21637, N22933);
or OR4 (N24219, N24210, N9069, N1048, N12839);
xor XOR2 (N24220, N24208, N14394);
xor XOR2 (N24221, N24192, N13730);
or OR4 (N24222, N24199, N13747, N22265, N22224);
not NOT1 (N24223, N24218);
nand NAND2 (N24224, N24213, N14864);
not NOT1 (N24225, N24217);
nand NAND4 (N24226, N24224, N7449, N19671, N16982);
buf BUF1 (N24227, N24216);
buf BUF1 (N24228, N24200);
buf BUF1 (N24229, N24222);
or OR2 (N24230, N24223, N24183);
nor NOR4 (N24231, N24214, N14288, N877, N16964);
not NOT1 (N24232, N24231);
nand NAND3 (N24233, N24225, N9243, N9926);
nand NAND3 (N24234, N24228, N22049, N22132);
not NOT1 (N24235, N24234);
xor XOR2 (N24236, N24233, N17056);
xor XOR2 (N24237, N24227, N14103);
nand NAND2 (N24238, N24219, N16833);
xor XOR2 (N24239, N24220, N10458);
and AND2 (N24240, N24226, N10920);
or OR2 (N24241, N24232, N15112);
or OR3 (N24242, N24235, N6520, N106);
nand NAND4 (N24243, N24236, N24037, N366, N22551);
and AND3 (N24244, N24239, N14796, N22421);
not NOT1 (N24245, N24230);
nand NAND4 (N24246, N24241, N10121, N8036, N6149);
nand NAND3 (N24247, N24245, N4745, N1920);
nor NOR4 (N24248, N24221, N7150, N1862, N4262);
buf BUF1 (N24249, N24229);
not NOT1 (N24250, N24240);
or OR3 (N24251, N24247, N901, N22286);
or OR2 (N24252, N24238, N6325);
and AND4 (N24253, N24250, N14534, N2980, N11288);
buf BUF1 (N24254, N24237);
not NOT1 (N24255, N24244);
buf BUF1 (N24256, N24251);
nand NAND3 (N24257, N24256, N14674, N22125);
nor NOR3 (N24258, N24242, N16323, N11744);
or OR4 (N24259, N24243, N15565, N9270, N20852);
nor NOR4 (N24260, N24248, N3748, N8660, N6621);
xor XOR2 (N24261, N24260, N955);
buf BUF1 (N24262, N24254);
not NOT1 (N24263, N24261);
nand NAND3 (N24264, N24253, N1035, N2957);
and AND4 (N24265, N24246, N17194, N3481, N21304);
or OR2 (N24266, N24259, N21708);
not NOT1 (N24267, N24249);
not NOT1 (N24268, N24258);
and AND3 (N24269, N24255, N17828, N7833);
and AND2 (N24270, N24268, N15657);
and AND3 (N24271, N24264, N14687, N10565);
buf BUF1 (N24272, N24257);
nor NOR4 (N24273, N24266, N22135, N16106, N10721);
nor NOR2 (N24274, N24273, N13914);
xor XOR2 (N24275, N24270, N16961);
xor XOR2 (N24276, N24272, N23826);
xor XOR2 (N24277, N24252, N13318);
nand NAND2 (N24278, N24277, N23557);
nor NOR3 (N24279, N24278, N18456, N23738);
nand NAND2 (N24280, N24275, N22840);
not NOT1 (N24281, N24269);
xor XOR2 (N24282, N24281, N11928);
buf BUF1 (N24283, N24262);
or OR4 (N24284, N24276, N6446, N2114, N16316);
buf BUF1 (N24285, N24280);
or OR2 (N24286, N24283, N20332);
nor NOR4 (N24287, N24286, N14084, N6737, N2640);
not NOT1 (N24288, N24284);
not NOT1 (N24289, N24285);
xor XOR2 (N24290, N24289, N24269);
and AND3 (N24291, N24274, N10189, N21719);
nor NOR4 (N24292, N24287, N23756, N17384, N571);
or OR4 (N24293, N24279, N21230, N10318, N15066);
buf BUF1 (N24294, N24288);
and AND4 (N24295, N24290, N6235, N16917, N3381);
xor XOR2 (N24296, N24282, N23881);
and AND2 (N24297, N24295, N14899);
nand NAND3 (N24298, N24267, N7833, N16774);
not NOT1 (N24299, N24265);
buf BUF1 (N24300, N24271);
xor XOR2 (N24301, N24298, N21561);
not NOT1 (N24302, N24263);
not NOT1 (N24303, N24299);
xor XOR2 (N24304, N24302, N8383);
buf BUF1 (N24305, N24297);
or OR2 (N24306, N24294, N14179);
or OR2 (N24307, N24292, N19886);
buf BUF1 (N24308, N24293);
or OR2 (N24309, N24301, N4895);
or OR3 (N24310, N24308, N14426, N12540);
xor XOR2 (N24311, N24296, N5970);
nand NAND2 (N24312, N24304, N10241);
buf BUF1 (N24313, N24300);
buf BUF1 (N24314, N24291);
buf BUF1 (N24315, N24311);
nor NOR2 (N24316, N24306, N20750);
not NOT1 (N24317, N24312);
nor NOR2 (N24318, N24317, N12425);
nand NAND2 (N24319, N24318, N3840);
nand NAND2 (N24320, N24310, N10978);
buf BUF1 (N24321, N24305);
and AND2 (N24322, N24309, N7681);
not NOT1 (N24323, N24303);
and AND4 (N24324, N24307, N20139, N11156, N15486);
buf BUF1 (N24325, N24316);
nand NAND4 (N24326, N24313, N13785, N15554, N15949);
not NOT1 (N24327, N24324);
buf BUF1 (N24328, N24322);
or OR3 (N24329, N24323, N2879, N22642);
or OR4 (N24330, N24328, N18711, N7059, N6512);
buf BUF1 (N24331, N24321);
or OR2 (N24332, N24330, N9667);
or OR4 (N24333, N24320, N13617, N15500, N7226);
buf BUF1 (N24334, N24333);
not NOT1 (N24335, N24329);
nand NAND2 (N24336, N24327, N981);
buf BUF1 (N24337, N24319);
xor XOR2 (N24338, N24315, N1376);
nand NAND3 (N24339, N24325, N20782, N15563);
not NOT1 (N24340, N24331);
buf BUF1 (N24341, N24332);
and AND3 (N24342, N24339, N24134, N2729);
not NOT1 (N24343, N24335);
nor NOR2 (N24344, N24326, N18700);
and AND2 (N24345, N24336, N4320);
nor NOR4 (N24346, N24338, N12997, N20734, N6953);
or OR3 (N24347, N24343, N23100, N15836);
not NOT1 (N24348, N24340);
nand NAND4 (N24349, N24341, N2344, N22885, N18904);
xor XOR2 (N24350, N24342, N1464);
nor NOR4 (N24351, N24345, N8891, N6781, N24144);
buf BUF1 (N24352, N24334);
nor NOR3 (N24353, N24314, N2695, N14269);
nor NOR4 (N24354, N24344, N123, N105, N2173);
nor NOR2 (N24355, N24351, N908);
xor XOR2 (N24356, N24352, N1524);
xor XOR2 (N24357, N24355, N19595);
not NOT1 (N24358, N24357);
buf BUF1 (N24359, N24346);
or OR2 (N24360, N24337, N21529);
and AND2 (N24361, N24353, N9245);
xor XOR2 (N24362, N24347, N13498);
xor XOR2 (N24363, N24361, N23964);
nand NAND3 (N24364, N24354, N5013, N18095);
and AND2 (N24365, N24349, N4475);
buf BUF1 (N24366, N24360);
or OR2 (N24367, N24364, N3258);
and AND4 (N24368, N24366, N14098, N23717, N900);
and AND2 (N24369, N24348, N10748);
nand NAND3 (N24370, N24368, N23835, N19853);
and AND2 (N24371, N24356, N1544);
and AND2 (N24372, N24358, N2080);
and AND2 (N24373, N24363, N12350);
and AND3 (N24374, N24372, N412, N22684);
and AND4 (N24375, N24350, N21706, N2827, N6807);
nand NAND2 (N24376, N24369, N9418);
nand NAND3 (N24377, N24359, N19586, N10807);
or OR4 (N24378, N24375, N16098, N9726, N8745);
nand NAND3 (N24379, N24365, N10100, N21112);
buf BUF1 (N24380, N24376);
buf BUF1 (N24381, N24367);
not NOT1 (N24382, N24379);
xor XOR2 (N24383, N24380, N2017);
buf BUF1 (N24384, N24373);
buf BUF1 (N24385, N24378);
or OR2 (N24386, N24377, N3542);
or OR2 (N24387, N24383, N20838);
xor XOR2 (N24388, N24362, N15792);
not NOT1 (N24389, N24384);
or OR4 (N24390, N24382, N23599, N16410, N5433);
or OR4 (N24391, N24385, N18921, N20163, N11019);
and AND3 (N24392, N24387, N9859, N12028);
buf BUF1 (N24393, N24392);
or OR3 (N24394, N24386, N2353, N18934);
nand NAND2 (N24395, N24390, N15297);
xor XOR2 (N24396, N24389, N15408);
not NOT1 (N24397, N24388);
not NOT1 (N24398, N24381);
nand NAND4 (N24399, N24395, N3032, N21769, N16501);
nor NOR4 (N24400, N24394, N12406, N22120, N11363);
not NOT1 (N24401, N24400);
not NOT1 (N24402, N24396);
buf BUF1 (N24403, N24374);
xor XOR2 (N24404, N24393, N11174);
and AND2 (N24405, N24399, N15664);
xor XOR2 (N24406, N24401, N22259);
buf BUF1 (N24407, N24370);
nand NAND4 (N24408, N24404, N7219, N4854, N20408);
xor XOR2 (N24409, N24397, N7323);
nor NOR4 (N24410, N24402, N9307, N15453, N22498);
not NOT1 (N24411, N24405);
nand NAND2 (N24412, N24409, N16949);
or OR4 (N24413, N24412, N107, N10664, N21823);
nand NAND3 (N24414, N24413, N2062, N11763);
nor NOR4 (N24415, N24406, N8599, N16615, N18112);
xor XOR2 (N24416, N24411, N12845);
buf BUF1 (N24417, N24403);
nor NOR4 (N24418, N24416, N6511, N2600, N3988);
or OR2 (N24419, N24407, N8514);
not NOT1 (N24420, N24415);
or OR3 (N24421, N24417, N4722, N8940);
buf BUF1 (N24422, N24419);
or OR2 (N24423, N24418, N385);
xor XOR2 (N24424, N24398, N19454);
not NOT1 (N24425, N24424);
nor NOR2 (N24426, N24423, N9285);
nand NAND3 (N24427, N24391, N20454, N2649);
xor XOR2 (N24428, N24410, N17086);
nand NAND3 (N24429, N24425, N4976, N8162);
buf BUF1 (N24430, N24428);
xor XOR2 (N24431, N24414, N8247);
xor XOR2 (N24432, N24429, N9787);
or OR2 (N24433, N24420, N3140);
nor NOR4 (N24434, N24431, N4943, N14765, N24196);
nand NAND3 (N24435, N24371, N10102, N14033);
nor NOR4 (N24436, N24435, N12971, N10822, N979);
nand NAND4 (N24437, N24436, N10826, N6239, N10382);
not NOT1 (N24438, N24421);
nor NOR3 (N24439, N24408, N16222, N24043);
xor XOR2 (N24440, N24426, N19214);
or OR2 (N24441, N24434, N5408);
nand NAND4 (N24442, N24440, N12635, N10196, N17892);
and AND2 (N24443, N24433, N17506);
buf BUF1 (N24444, N24437);
nor NOR3 (N24445, N24430, N18232, N10818);
nand NAND3 (N24446, N24443, N1509, N19242);
and AND3 (N24447, N24438, N12488, N11086);
nand NAND3 (N24448, N24439, N13975, N20029);
nor NOR2 (N24449, N24422, N16156);
not NOT1 (N24450, N24448);
buf BUF1 (N24451, N24442);
not NOT1 (N24452, N24445);
nor NOR3 (N24453, N24447, N7600, N16453);
or OR3 (N24454, N24444, N19915, N22967);
nand NAND4 (N24455, N24446, N1668, N6259, N18753);
and AND2 (N24456, N24453, N19705);
and AND3 (N24457, N24451, N11495, N2850);
buf BUF1 (N24458, N24427);
xor XOR2 (N24459, N24441, N9187);
buf BUF1 (N24460, N24454);
nor NOR4 (N24461, N24450, N13180, N22117, N18717);
nand NAND4 (N24462, N24455, N15949, N3821, N2337);
nor NOR2 (N24463, N24457, N16575);
and AND4 (N24464, N24432, N14232, N18093, N3621);
buf BUF1 (N24465, N24462);
not NOT1 (N24466, N24456);
and AND2 (N24467, N24461, N16949);
nor NOR4 (N24468, N24466, N21605, N6709, N19878);
nand NAND4 (N24469, N24464, N16263, N21814, N12352);
buf BUF1 (N24470, N24449);
not NOT1 (N24471, N24469);
buf BUF1 (N24472, N24460);
nor NOR4 (N24473, N24463, N20130, N22596, N15866);
not NOT1 (N24474, N24468);
and AND2 (N24475, N24465, N8300);
buf BUF1 (N24476, N24470);
buf BUF1 (N24477, N24458);
and AND3 (N24478, N24472, N20419, N4370);
and AND4 (N24479, N24477, N12039, N5969, N7240);
buf BUF1 (N24480, N24475);
xor XOR2 (N24481, N24459, N23758);
nor NOR4 (N24482, N24471, N5561, N9970, N7559);
and AND3 (N24483, N24473, N13591, N20266);
and AND2 (N24484, N24482, N23186);
buf BUF1 (N24485, N24484);
not NOT1 (N24486, N24476);
buf BUF1 (N24487, N24479);
nor NOR4 (N24488, N24481, N6599, N11806, N924);
buf BUF1 (N24489, N24486);
or OR2 (N24490, N24478, N529);
xor XOR2 (N24491, N24474, N23684);
xor XOR2 (N24492, N24490, N4917);
xor XOR2 (N24493, N24487, N23718);
not NOT1 (N24494, N24488);
nor NOR2 (N24495, N24493, N15060);
buf BUF1 (N24496, N24489);
xor XOR2 (N24497, N24494, N20380);
nand NAND4 (N24498, N24495, N7635, N10186, N240);
and AND3 (N24499, N24491, N13051, N8379);
nand NAND4 (N24500, N24483, N24454, N5111, N4837);
or OR4 (N24501, N24499, N8846, N17376, N10203);
not NOT1 (N24502, N24501);
or OR3 (N24503, N24452, N4839, N1225);
nand NAND3 (N24504, N24485, N20297, N5859);
buf BUF1 (N24505, N24503);
or OR3 (N24506, N24496, N21345, N17452);
nand NAND2 (N24507, N24467, N24506);
not NOT1 (N24508, N12192);
and AND3 (N24509, N24508, N19782, N12735);
not NOT1 (N24510, N24500);
xor XOR2 (N24511, N24492, N8260);
nor NOR4 (N24512, N24480, N3521, N3834, N10461);
buf BUF1 (N24513, N24504);
or OR2 (N24514, N24498, N12711);
buf BUF1 (N24515, N24514);
xor XOR2 (N24516, N24515, N6751);
and AND2 (N24517, N24511, N20185);
buf BUF1 (N24518, N24502);
and AND3 (N24519, N24513, N22415, N23006);
and AND4 (N24520, N24519, N12506, N13267, N8490);
not NOT1 (N24521, N24497);
xor XOR2 (N24522, N24518, N16173);
and AND4 (N24523, N24510, N20626, N18369, N19182);
nor NOR2 (N24524, N24505, N12823);
xor XOR2 (N24525, N24524, N15884);
nor NOR4 (N24526, N24520, N10252, N5507, N18679);
not NOT1 (N24527, N24526);
nand NAND4 (N24528, N24522, N18651, N17045, N21157);
buf BUF1 (N24529, N24525);
nor NOR4 (N24530, N24528, N904, N7666, N13509);
nand NAND3 (N24531, N24530, N13649, N4359);
or OR3 (N24532, N24517, N11759, N228);
and AND3 (N24533, N24532, N9324, N11224);
nor NOR4 (N24534, N24509, N21882, N14216, N11327);
and AND2 (N24535, N24521, N20384);
buf BUF1 (N24536, N24527);
or OR4 (N24537, N24529, N18422, N13730, N12681);
nand NAND2 (N24538, N24516, N10331);
not NOT1 (N24539, N24537);
nand NAND3 (N24540, N24523, N12751, N14830);
or OR2 (N24541, N24533, N23637);
and AND2 (N24542, N24540, N1958);
xor XOR2 (N24543, N24531, N8460);
xor XOR2 (N24544, N24535, N13098);
and AND2 (N24545, N24542, N24053);
nor NOR4 (N24546, N24536, N6138, N2720, N17969);
xor XOR2 (N24547, N24507, N12037);
buf BUF1 (N24548, N24539);
not NOT1 (N24549, N24545);
or OR3 (N24550, N24512, N18238, N21001);
nor NOR4 (N24551, N24534, N3855, N15524, N23027);
nor NOR2 (N24552, N24549, N5049);
nand NAND3 (N24553, N24546, N6095, N15818);
nor NOR3 (N24554, N24544, N2343, N7938);
xor XOR2 (N24555, N24550, N19223);
not NOT1 (N24556, N24552);
not NOT1 (N24557, N24551);
nand NAND3 (N24558, N24555, N12534, N17767);
nor NOR3 (N24559, N24548, N1781, N16903);
nand NAND4 (N24560, N24538, N18862, N9074, N19623);
not NOT1 (N24561, N24543);
and AND2 (N24562, N24547, N5135);
nand NAND2 (N24563, N24541, N11113);
buf BUF1 (N24564, N24562);
nor NOR3 (N24565, N24564, N10088, N17904);
nor NOR2 (N24566, N24557, N23837);
nor NOR3 (N24567, N24566, N24203, N20668);
or OR3 (N24568, N24563, N8682, N18631);
not NOT1 (N24569, N24567);
or OR4 (N24570, N24569, N24331, N18553, N6193);
nand NAND4 (N24571, N24560, N615, N10593, N23954);
nand NAND3 (N24572, N24558, N23052, N780);
xor XOR2 (N24573, N24556, N5712);
buf BUF1 (N24574, N24553);
nand NAND3 (N24575, N24574, N18887, N19101);
not NOT1 (N24576, N24575);
and AND4 (N24577, N24554, N5282, N10030, N14992);
buf BUF1 (N24578, N24568);
nand NAND2 (N24579, N24572, N360);
buf BUF1 (N24580, N24559);
or OR2 (N24581, N24579, N7581);
nand NAND2 (N24582, N24576, N19721);
nor NOR4 (N24583, N24580, N6780, N3430, N5845);
and AND2 (N24584, N24578, N537);
and AND2 (N24585, N24582, N16648);
buf BUF1 (N24586, N24583);
xor XOR2 (N24587, N24586, N17397);
xor XOR2 (N24588, N24571, N8117);
or OR2 (N24589, N24585, N19233);
not NOT1 (N24590, N24587);
nor NOR4 (N24591, N24589, N21750, N24448, N21390);
and AND2 (N24592, N24570, N9815);
nand NAND4 (N24593, N24573, N3923, N5294, N4427);
not NOT1 (N24594, N24590);
xor XOR2 (N24595, N24588, N8889);
nand NAND2 (N24596, N24584, N6075);
nand NAND2 (N24597, N24592, N21624);
or OR4 (N24598, N24581, N7751, N620, N7295);
not NOT1 (N24599, N24596);
not NOT1 (N24600, N24599);
buf BUF1 (N24601, N24593);
xor XOR2 (N24602, N24600, N11822);
xor XOR2 (N24603, N24597, N711);
xor XOR2 (N24604, N24598, N9607);
nand NAND3 (N24605, N24595, N541, N10106);
and AND4 (N24606, N24601, N8006, N4451, N3557);
nand NAND3 (N24607, N24604, N20448, N23905);
and AND2 (N24608, N24603, N12923);
buf BUF1 (N24609, N24602);
not NOT1 (N24610, N24565);
buf BUF1 (N24611, N24605);
xor XOR2 (N24612, N24608, N12824);
nor NOR3 (N24613, N24612, N19122, N2924);
xor XOR2 (N24614, N24613, N14102);
and AND2 (N24615, N24561, N2185);
nand NAND4 (N24616, N24610, N3742, N6148, N19455);
buf BUF1 (N24617, N24577);
or OR4 (N24618, N24617, N21072, N18158, N1653);
and AND2 (N24619, N24594, N6869);
and AND2 (N24620, N24591, N11453);
and AND3 (N24621, N24611, N23283, N5915);
or OR4 (N24622, N24606, N18158, N17156, N13992);
not NOT1 (N24623, N24622);
or OR2 (N24624, N24614, N14244);
or OR4 (N24625, N24623, N21493, N17032, N2163);
xor XOR2 (N24626, N24619, N9089);
or OR3 (N24627, N24626, N2607, N8347);
and AND2 (N24628, N24625, N3702);
nor NOR2 (N24629, N24616, N14555);
buf BUF1 (N24630, N24629);
xor XOR2 (N24631, N24621, N6524);
buf BUF1 (N24632, N24618);
buf BUF1 (N24633, N24609);
nand NAND3 (N24634, N24607, N4121, N17866);
nand NAND2 (N24635, N24627, N10914);
and AND3 (N24636, N24631, N584, N13831);
or OR2 (N24637, N24624, N23307);
buf BUF1 (N24638, N24615);
nor NOR4 (N24639, N24620, N14654, N9268, N21030);
not NOT1 (N24640, N24632);
buf BUF1 (N24641, N24628);
and AND2 (N24642, N24636, N5041);
nor NOR4 (N24643, N24638, N6076, N6053, N11066);
xor XOR2 (N24644, N24634, N21409);
buf BUF1 (N24645, N24643);
nand NAND2 (N24646, N24633, N4737);
nand NAND3 (N24647, N24637, N468, N15176);
not NOT1 (N24648, N24645);
xor XOR2 (N24649, N24642, N8358);
nor NOR4 (N24650, N24646, N6316, N5433, N4479);
nand NAND2 (N24651, N24647, N2790);
and AND4 (N24652, N24630, N9676, N1118, N9428);
nor NOR3 (N24653, N24650, N19795, N1468);
nor NOR4 (N24654, N24635, N11620, N18913, N24582);
not NOT1 (N24655, N24639);
not NOT1 (N24656, N24652);
buf BUF1 (N24657, N24653);
xor XOR2 (N24658, N24656, N16362);
or OR3 (N24659, N24640, N21081, N18965);
nand NAND2 (N24660, N24659, N18832);
and AND4 (N24661, N24660, N214, N14693, N13401);
nand NAND4 (N24662, N24644, N5228, N3112, N3711);
nor NOR4 (N24663, N24655, N20730, N1101, N12432);
not NOT1 (N24664, N24648);
not NOT1 (N24665, N24641);
nand NAND4 (N24666, N24661, N1951, N9271, N2151);
nor NOR3 (N24667, N24664, N20198, N20926);
nand NAND3 (N24668, N24651, N767, N11874);
buf BUF1 (N24669, N24657);
nand NAND4 (N24670, N24662, N10338, N2145, N23266);
nor NOR2 (N24671, N24663, N16201);
not NOT1 (N24672, N24670);
nand NAND2 (N24673, N24669, N24442);
nand NAND4 (N24674, N24667, N7623, N13511, N9462);
buf BUF1 (N24675, N24672);
xor XOR2 (N24676, N24666, N10823);
buf BUF1 (N24677, N24668);
not NOT1 (N24678, N24675);
xor XOR2 (N24679, N24676, N6738);
not NOT1 (N24680, N24674);
buf BUF1 (N24681, N24673);
buf BUF1 (N24682, N24680);
buf BUF1 (N24683, N24681);
nand NAND2 (N24684, N24649, N4259);
nor NOR3 (N24685, N24682, N7477, N18765);
nor NOR3 (N24686, N24658, N7292, N22580);
nor NOR3 (N24687, N24677, N300, N114);
nand NAND4 (N24688, N24671, N22431, N16783, N19534);
and AND2 (N24689, N24685, N9358);
or OR2 (N24690, N24687, N9540);
xor XOR2 (N24691, N24689, N215);
buf BUF1 (N24692, N24683);
nand NAND4 (N24693, N24654, N8007, N5331, N3159);
and AND4 (N24694, N24688, N12704, N11494, N24296);
buf BUF1 (N24695, N24678);
nand NAND3 (N24696, N24691, N18904, N7046);
xor XOR2 (N24697, N24684, N20415);
or OR2 (N24698, N24696, N5174);
and AND2 (N24699, N24697, N10815);
buf BUF1 (N24700, N24698);
buf BUF1 (N24701, N24690);
not NOT1 (N24702, N24692);
nand NAND4 (N24703, N24693, N6140, N3399, N18730);
xor XOR2 (N24704, N24694, N4427);
xor XOR2 (N24705, N24700, N12728);
not NOT1 (N24706, N24665);
buf BUF1 (N24707, N24686);
nand NAND4 (N24708, N24707, N22253, N6400, N15293);
buf BUF1 (N24709, N24699);
not NOT1 (N24710, N24702);
not NOT1 (N24711, N24695);
and AND3 (N24712, N24701, N16209, N16402);
xor XOR2 (N24713, N24709, N6667);
xor XOR2 (N24714, N24710, N11549);
not NOT1 (N24715, N24714);
not NOT1 (N24716, N24679);
and AND3 (N24717, N24712, N18171, N2270);
or OR3 (N24718, N24703, N14617, N3309);
and AND3 (N24719, N24711, N4517, N15253);
nand NAND2 (N24720, N24706, N3285);
or OR4 (N24721, N24705, N15710, N23793, N22841);
nand NAND2 (N24722, N24713, N4415);
or OR3 (N24723, N24716, N8281, N19659);
not NOT1 (N24724, N24708);
and AND4 (N24725, N24717, N4615, N16140, N8849);
not NOT1 (N24726, N24721);
xor XOR2 (N24727, N24720, N16404);
nand NAND2 (N24728, N24726, N1999);
or OR4 (N24729, N24724, N11590, N10068, N6227);
nor NOR4 (N24730, N24704, N5347, N12042, N18926);
or OR3 (N24731, N24725, N20707, N23338);
buf BUF1 (N24732, N24728);
nand NAND4 (N24733, N24729, N5542, N5973, N21662);
and AND3 (N24734, N24722, N14178, N12897);
nand NAND4 (N24735, N24733, N2885, N11470, N1256);
buf BUF1 (N24736, N24719);
nor NOR4 (N24737, N24730, N13279, N4895, N21439);
or OR3 (N24738, N24731, N22873, N15405);
nand NAND4 (N24739, N24727, N7140, N11747, N23975);
nand NAND4 (N24740, N24715, N651, N3287, N3983);
not NOT1 (N24741, N24718);
nand NAND3 (N24742, N24740, N5032, N3558);
xor XOR2 (N24743, N24739, N21960);
nor NOR3 (N24744, N24738, N17680, N630);
not NOT1 (N24745, N24735);
and AND4 (N24746, N24734, N10866, N17957, N13616);
and AND4 (N24747, N24744, N2864, N12176, N11347);
buf BUF1 (N24748, N24742);
buf BUF1 (N24749, N24736);
or OR4 (N24750, N24747, N19793, N22140, N9527);
buf BUF1 (N24751, N24741);
and AND3 (N24752, N24748, N24595, N13052);
xor XOR2 (N24753, N24746, N16119);
xor XOR2 (N24754, N24743, N2744);
not NOT1 (N24755, N24754);
nand NAND2 (N24756, N24755, N16115);
or OR3 (N24757, N24750, N2411, N17197);
buf BUF1 (N24758, N24732);
not NOT1 (N24759, N24756);
or OR2 (N24760, N24753, N14374);
and AND3 (N24761, N24758, N17798, N8628);
buf BUF1 (N24762, N24751);
buf BUF1 (N24763, N24762);
xor XOR2 (N24764, N24723, N3);
not NOT1 (N24765, N24737);
nand NAND2 (N24766, N24764, N6644);
buf BUF1 (N24767, N24745);
nor NOR3 (N24768, N24766, N3817, N16704);
or OR3 (N24769, N24759, N8459, N6139);
xor XOR2 (N24770, N24760, N7020);
nor NOR4 (N24771, N24757, N12753, N18129, N15054);
xor XOR2 (N24772, N24768, N23005);
xor XOR2 (N24773, N24770, N8089);
and AND2 (N24774, N24769, N14476);
not NOT1 (N24775, N24774);
xor XOR2 (N24776, N24752, N6053);
nand NAND2 (N24777, N24761, N2119);
nor NOR3 (N24778, N24767, N2807, N9554);
xor XOR2 (N24779, N24776, N22718);
nor NOR2 (N24780, N24779, N18150);
nor NOR4 (N24781, N24773, N24280, N4758, N19773);
buf BUF1 (N24782, N24765);
and AND4 (N24783, N24749, N20590, N18833, N7988);
or OR3 (N24784, N24777, N18886, N8773);
nor NOR3 (N24785, N24778, N3556, N21201);
or OR3 (N24786, N24775, N14951, N1156);
xor XOR2 (N24787, N24783, N19790);
and AND3 (N24788, N24772, N24293, N6874);
buf BUF1 (N24789, N24787);
buf BUF1 (N24790, N24789);
nor NOR3 (N24791, N24763, N1988, N15969);
not NOT1 (N24792, N24784);
nor NOR3 (N24793, N24782, N14042, N22472);
and AND3 (N24794, N24793, N8151, N3230);
xor XOR2 (N24795, N24790, N14678);
nor NOR2 (N24796, N24780, N21029);
nor NOR3 (N24797, N24791, N19892, N1951);
and AND4 (N24798, N24781, N3801, N18322, N4961);
xor XOR2 (N24799, N24792, N24594);
or OR3 (N24800, N24796, N6104, N10924);
nand NAND3 (N24801, N24800, N7781, N21163);
not NOT1 (N24802, N24771);
nor NOR2 (N24803, N24788, N15151);
buf BUF1 (N24804, N24799);
or OR3 (N24805, N24794, N14927, N3663);
nor NOR3 (N24806, N24805, N8014, N20719);
nor NOR3 (N24807, N24806, N4697, N12541);
nand NAND4 (N24808, N24785, N781, N7961, N24161);
nand NAND3 (N24809, N24798, N17907, N13396);
not NOT1 (N24810, N24797);
nor NOR2 (N24811, N24810, N22897);
nand NAND4 (N24812, N24803, N21414, N3918, N18191);
nand NAND4 (N24813, N24801, N15304, N7807, N13915);
nand NAND3 (N24814, N24811, N10673, N18533);
or OR3 (N24815, N24807, N19081, N20658);
xor XOR2 (N24816, N24813, N1179);
nand NAND4 (N24817, N24802, N23676, N4282, N22238);
or OR3 (N24818, N24808, N20647, N428);
nor NOR2 (N24819, N24795, N4618);
or OR3 (N24820, N24812, N14570, N14969);
nor NOR4 (N24821, N24815, N22732, N15537, N22153);
nor NOR2 (N24822, N24819, N10627);
and AND3 (N24823, N24821, N10524, N12413);
buf BUF1 (N24824, N24823);
not NOT1 (N24825, N24824);
nand NAND3 (N24826, N24822, N21765, N24179);
and AND4 (N24827, N24820, N19620, N12752, N17394);
or OR2 (N24828, N24827, N21797);
nand NAND3 (N24829, N24817, N11933, N12942);
nand NAND4 (N24830, N24818, N6278, N14925, N16791);
or OR3 (N24831, N24814, N23495, N19264);
buf BUF1 (N24832, N24786);
nand NAND4 (N24833, N24826, N11299, N14821, N14635);
buf BUF1 (N24834, N24832);
and AND2 (N24835, N24831, N19717);
and AND4 (N24836, N24834, N7552, N3324, N9829);
and AND4 (N24837, N24828, N14105, N5715, N3306);
buf BUF1 (N24838, N24833);
nor NOR4 (N24839, N24838, N7777, N7272, N9371);
nand NAND2 (N24840, N24829, N4162);
nand NAND4 (N24841, N24804, N18481, N16996, N23471);
not NOT1 (N24842, N24830);
or OR4 (N24843, N24825, N4671, N14675, N11289);
and AND4 (N24844, N24842, N5651, N4195, N7665);
nor NOR4 (N24845, N24839, N6459, N11215, N9602);
not NOT1 (N24846, N24835);
buf BUF1 (N24847, N24837);
not NOT1 (N24848, N24816);
nand NAND2 (N24849, N24843, N20693);
buf BUF1 (N24850, N24840);
and AND4 (N24851, N24846, N15328, N2040, N373);
and AND3 (N24852, N24836, N1762, N6170);
or OR4 (N24853, N24847, N3407, N13505, N15818);
buf BUF1 (N24854, N24841);
not NOT1 (N24855, N24844);
xor XOR2 (N24856, N24852, N24078);
not NOT1 (N24857, N24850);
buf BUF1 (N24858, N24845);
nand NAND2 (N24859, N24855, N18899);
nor NOR3 (N24860, N24809, N2785, N15836);
and AND2 (N24861, N24848, N1953);
buf BUF1 (N24862, N24859);
or OR2 (N24863, N24857, N1355);
or OR2 (N24864, N24860, N9880);
or OR3 (N24865, N24858, N326, N1857);
xor XOR2 (N24866, N24849, N3994);
nor NOR3 (N24867, N24861, N9505, N22743);
and AND3 (N24868, N24866, N2632, N9727);
nand NAND4 (N24869, N24862, N15751, N8526, N3037);
buf BUF1 (N24870, N24851);
nor NOR3 (N24871, N24867, N9071, N23642);
xor XOR2 (N24872, N24871, N37);
not NOT1 (N24873, N24869);
not NOT1 (N24874, N24873);
xor XOR2 (N24875, N24864, N21620);
and AND3 (N24876, N24853, N15547, N12774);
or OR2 (N24877, N24856, N17803);
xor XOR2 (N24878, N24854, N13326);
and AND3 (N24879, N24863, N8264, N15042);
nor NOR2 (N24880, N24875, N13850);
or OR2 (N24881, N24880, N22824);
buf BUF1 (N24882, N24870);
or OR4 (N24883, N24882, N20714, N12250, N8056);
and AND4 (N24884, N24872, N12391, N3738, N10152);
not NOT1 (N24885, N24865);
nand NAND2 (N24886, N24879, N9543);
xor XOR2 (N24887, N24883, N238);
or OR3 (N24888, N24884, N2280, N21299);
xor XOR2 (N24889, N24887, N23471);
nand NAND3 (N24890, N24877, N17354, N19048);
or OR3 (N24891, N24868, N3285, N15435);
nor NOR3 (N24892, N24890, N132, N17792);
xor XOR2 (N24893, N24888, N22794);
nor NOR2 (N24894, N24874, N1514);
nand NAND4 (N24895, N24886, N10897, N7231, N1977);
nand NAND2 (N24896, N24894, N3803);
xor XOR2 (N24897, N24893, N7782);
not NOT1 (N24898, N24889);
and AND4 (N24899, N24896, N3388, N20058, N9039);
and AND3 (N24900, N24878, N4101, N19009);
xor XOR2 (N24901, N24895, N7470);
xor XOR2 (N24902, N24892, N14415);
not NOT1 (N24903, N24897);
xor XOR2 (N24904, N24881, N10741);
not NOT1 (N24905, N24901);
or OR2 (N24906, N24900, N23587);
nor NOR3 (N24907, N24899, N22890, N13568);
nand NAND2 (N24908, N24906, N11148);
not NOT1 (N24909, N24908);
and AND2 (N24910, N24905, N14805);
not NOT1 (N24911, N24898);
buf BUF1 (N24912, N24904);
nand NAND4 (N24913, N24907, N2417, N17198, N4568);
nand NAND3 (N24914, N24912, N9613, N21388);
and AND3 (N24915, N24902, N13834, N9984);
or OR3 (N24916, N24911, N24774, N4203);
buf BUF1 (N24917, N24914);
buf BUF1 (N24918, N24916);
xor XOR2 (N24919, N24885, N22186);
nand NAND3 (N24920, N24915, N20832, N17631);
not NOT1 (N24921, N24917);
buf BUF1 (N24922, N24921);
and AND2 (N24923, N24891, N8074);
xor XOR2 (N24924, N24909, N18270);
nor NOR3 (N24925, N24913, N10056, N526);
not NOT1 (N24926, N24876);
or OR4 (N24927, N24926, N23906, N22063, N11968);
not NOT1 (N24928, N24910);
and AND2 (N24929, N24919, N19110);
not NOT1 (N24930, N24925);
and AND3 (N24931, N24929, N9908, N19981);
not NOT1 (N24932, N24918);
xor XOR2 (N24933, N24924, N16570);
xor XOR2 (N24934, N24933, N19871);
and AND2 (N24935, N24932, N21128);
not NOT1 (N24936, N24931);
nor NOR2 (N24937, N24922, N5980);
and AND4 (N24938, N24934, N23544, N10247, N19012);
and AND4 (N24939, N24923, N17822, N5338, N17984);
and AND4 (N24940, N24939, N4116, N2987, N6247);
or OR3 (N24941, N24936, N14585, N18033);
nor NOR3 (N24942, N24941, N22429, N11716);
nor NOR2 (N24943, N24920, N7563);
or OR4 (N24944, N24903, N4133, N14868, N2325);
not NOT1 (N24945, N24935);
buf BUF1 (N24946, N24927);
buf BUF1 (N24947, N24928);
xor XOR2 (N24948, N24940, N8132);
and AND2 (N24949, N24944, N4462);
nor NOR2 (N24950, N24942, N23484);
or OR4 (N24951, N24937, N16027, N4105, N78);
buf BUF1 (N24952, N24930);
or OR3 (N24953, N24950, N23426, N586);
nand NAND3 (N24954, N24945, N9274, N7880);
nor NOR4 (N24955, N24946, N5985, N19089, N13473);
buf BUF1 (N24956, N24947);
nand NAND4 (N24957, N24938, N21, N16970, N12827);
nand NAND2 (N24958, N24955, N16965);
xor XOR2 (N24959, N24948, N22371);
buf BUF1 (N24960, N24949);
nor NOR2 (N24961, N24951, N21862);
not NOT1 (N24962, N24957);
xor XOR2 (N24963, N24960, N6416);
and AND2 (N24964, N24952, N16521);
buf BUF1 (N24965, N24962);
buf BUF1 (N24966, N24953);
or OR2 (N24967, N24964, N10196);
xor XOR2 (N24968, N24954, N19427);
nor NOR2 (N24969, N24965, N17791);
nor NOR3 (N24970, N24968, N13425, N11901);
nor NOR2 (N24971, N24956, N14247);
xor XOR2 (N24972, N24967, N7788);
or OR2 (N24973, N24972, N16412);
and AND3 (N24974, N24971, N5056, N6293);
or OR4 (N24975, N24958, N18011, N16609, N2763);
nor NOR4 (N24976, N24961, N6788, N7687, N16520);
nor NOR2 (N24977, N24966, N11743);
not NOT1 (N24978, N24943);
nand NAND4 (N24979, N24975, N617, N14231, N11279);
or OR2 (N24980, N24979, N5574);
nand NAND3 (N24981, N24976, N11370, N2841);
xor XOR2 (N24982, N24978, N2461);
buf BUF1 (N24983, N24963);
nand NAND4 (N24984, N24974, N8400, N5842, N9255);
xor XOR2 (N24985, N24982, N4395);
and AND4 (N24986, N24984, N12778, N5097, N10081);
and AND3 (N24987, N24977, N12591, N4677);
buf BUF1 (N24988, N24980);
nor NOR4 (N24989, N24985, N4634, N21623, N590);
or OR4 (N24990, N24969, N13326, N7890, N12697);
or OR4 (N24991, N24986, N22482, N14217, N4779);
buf BUF1 (N24992, N24983);
nor NOR3 (N24993, N24987, N15309, N12555);
buf BUF1 (N24994, N24992);
buf BUF1 (N24995, N24988);
or OR3 (N24996, N24995, N15818, N9664);
nand NAND4 (N24997, N24959, N1794, N10790, N23492);
and AND2 (N24998, N24973, N4466);
nor NOR3 (N24999, N24997, N10987, N17807);
and AND2 (N25000, N24998, N14121);
or OR2 (N25001, N24989, N24808);
xor XOR2 (N25002, N24981, N9522);
xor XOR2 (N25003, N24994, N6279);
and AND4 (N25004, N24999, N24913, N4685, N18789);
and AND3 (N25005, N24991, N10012, N8783);
buf BUF1 (N25006, N25000);
not NOT1 (N25007, N24990);
nor NOR3 (N25008, N25004, N6477, N11722);
xor XOR2 (N25009, N24993, N4379);
and AND2 (N25010, N24996, N10921);
xor XOR2 (N25011, N24970, N21657);
not NOT1 (N25012, N25008);
nor NOR3 (N25013, N25003, N5623, N17898);
and AND2 (N25014, N25005, N18210);
xor XOR2 (N25015, N25007, N19725);
or OR3 (N25016, N25009, N13904, N16866);
or OR4 (N25017, N25016, N9561, N2395, N23275);
or OR4 (N25018, N25010, N22081, N8743, N9690);
or OR2 (N25019, N25006, N10287);
buf BUF1 (N25020, N25019);
not NOT1 (N25021, N25013);
nand NAND2 (N25022, N25012, N8706);
not NOT1 (N25023, N25014);
nor NOR3 (N25024, N25011, N21822, N19015);
xor XOR2 (N25025, N25017, N8772);
nor NOR2 (N25026, N25001, N13185);
and AND2 (N25027, N25015, N6071);
nand NAND4 (N25028, N25002, N5926, N8730, N11810);
nand NAND3 (N25029, N25018, N650, N1015);
or OR3 (N25030, N25022, N18254, N11359);
nor NOR4 (N25031, N25023, N5808, N12139, N14448);
nand NAND4 (N25032, N25028, N18763, N12149, N24279);
nor NOR3 (N25033, N25027, N23235, N24357);
and AND4 (N25034, N25031, N11551, N17843, N9592);
nand NAND2 (N25035, N25029, N2338);
nor NOR2 (N25036, N25030, N9890);
nor NOR2 (N25037, N25032, N22723);
not NOT1 (N25038, N25026);
and AND3 (N25039, N25024, N21450, N24520);
not NOT1 (N25040, N25037);
xor XOR2 (N25041, N25036, N23915);
or OR3 (N25042, N25041, N2803, N8356);
nand NAND2 (N25043, N25040, N14580);
nor NOR2 (N25044, N25039, N19387);
buf BUF1 (N25045, N25038);
or OR4 (N25046, N25033, N8804, N10809, N14625);
nand NAND2 (N25047, N25042, N15665);
buf BUF1 (N25048, N25046);
not NOT1 (N25049, N25048);
nor NOR2 (N25050, N25020, N2676);
or OR4 (N25051, N25044, N22379, N22212, N10328);
buf BUF1 (N25052, N25045);
nor NOR3 (N25053, N25025, N14007, N18720);
xor XOR2 (N25054, N25050, N10537);
nand NAND4 (N25055, N25051, N16129, N3500, N7241);
and AND4 (N25056, N25034, N22849, N3170, N3461);
or OR2 (N25057, N25043, N11675);
not NOT1 (N25058, N25057);
or OR4 (N25059, N25021, N132, N7722, N22629);
nand NAND3 (N25060, N25035, N9869, N7667);
nand NAND3 (N25061, N25049, N6359, N20804);
xor XOR2 (N25062, N25053, N1343);
or OR2 (N25063, N25047, N4782);
not NOT1 (N25064, N25056);
xor XOR2 (N25065, N25052, N8772);
not NOT1 (N25066, N25055);
or OR2 (N25067, N25063, N3601);
not NOT1 (N25068, N25054);
not NOT1 (N25069, N25064);
not NOT1 (N25070, N25060);
or OR3 (N25071, N25061, N1108, N24112);
or OR2 (N25072, N25066, N23233);
buf BUF1 (N25073, N25058);
xor XOR2 (N25074, N25072, N16392);
and AND2 (N25075, N25059, N15744);
nor NOR2 (N25076, N25068, N2868);
or OR4 (N25077, N25062, N21144, N472, N22210);
buf BUF1 (N25078, N25071);
or OR4 (N25079, N25074, N10150, N4072, N21392);
or OR2 (N25080, N25079, N19466);
not NOT1 (N25081, N25078);
xor XOR2 (N25082, N25069, N11876);
or OR2 (N25083, N25080, N17068);
nand NAND4 (N25084, N25073, N17869, N21262, N16014);
buf BUF1 (N25085, N25076);
or OR4 (N25086, N25075, N9454, N12503, N1886);
nor NOR4 (N25087, N25077, N4091, N15276, N4741);
nor NOR2 (N25088, N25085, N18037);
nand NAND4 (N25089, N25083, N17096, N24414, N4490);
and AND2 (N25090, N25065, N6408);
or OR4 (N25091, N25084, N11240, N23870, N3618);
buf BUF1 (N25092, N25070);
nor NOR4 (N25093, N25082, N11837, N22312, N18334);
or OR4 (N25094, N25067, N19615, N7626, N5407);
xor XOR2 (N25095, N25092, N2278);
not NOT1 (N25096, N25089);
nand NAND4 (N25097, N25094, N4982, N19434, N23925);
nand NAND3 (N25098, N25096, N18276, N499);
buf BUF1 (N25099, N25081);
or OR4 (N25100, N25095, N2128, N1111, N17716);
not NOT1 (N25101, N25100);
not NOT1 (N25102, N25098);
xor XOR2 (N25103, N25091, N8173);
and AND4 (N25104, N25099, N16256, N15554, N20813);
and AND2 (N25105, N25097, N9444);
or OR4 (N25106, N25086, N19712, N17761, N23578);
or OR2 (N25107, N25102, N1114);
or OR4 (N25108, N25093, N15504, N1407, N3052);
nand NAND3 (N25109, N25103, N55, N5716);
and AND4 (N25110, N25087, N3176, N1560, N20880);
nand NAND3 (N25111, N25107, N24944, N9989);
nor NOR2 (N25112, N25106, N9570);
buf BUF1 (N25113, N25111);
and AND3 (N25114, N25112, N8850, N24892);
nand NAND2 (N25115, N25108, N12669);
nor NOR2 (N25116, N25105, N3908);
and AND3 (N25117, N25115, N9972, N1191);
nand NAND4 (N25118, N25116, N14956, N16559, N1576);
buf BUF1 (N25119, N25088);
not NOT1 (N25120, N25101);
not NOT1 (N25121, N25110);
or OR3 (N25122, N25117, N9711, N14619);
xor XOR2 (N25123, N25109, N24766);
and AND2 (N25124, N25122, N15458);
nand NAND4 (N25125, N25124, N2949, N7725, N8220);
nor NOR2 (N25126, N25121, N16509);
nand NAND2 (N25127, N25126, N4660);
nor NOR3 (N25128, N25127, N2641, N14132);
or OR4 (N25129, N25114, N3553, N14375, N22443);
and AND3 (N25130, N25128, N20741, N6253);
not NOT1 (N25131, N25129);
xor XOR2 (N25132, N25125, N16453);
and AND4 (N25133, N25130, N14709, N12290, N10514);
nor NOR3 (N25134, N25120, N23449, N1033);
or OR2 (N25135, N25119, N13441);
and AND2 (N25136, N25133, N19503);
nor NOR4 (N25137, N25134, N4018, N13972, N4293);
buf BUF1 (N25138, N25131);
nor NOR2 (N25139, N25090, N16760);
xor XOR2 (N25140, N25137, N9641);
or OR3 (N25141, N25113, N7056, N15565);
and AND4 (N25142, N25135, N21866, N1545, N12378);
or OR3 (N25143, N25123, N5494, N19419);
nand NAND3 (N25144, N25136, N14758, N18499);
nor NOR3 (N25145, N25143, N18403, N6946);
nor NOR2 (N25146, N25140, N19686);
and AND4 (N25147, N25142, N11923, N2862, N17259);
xor XOR2 (N25148, N25139, N21350);
buf BUF1 (N25149, N25148);
or OR4 (N25150, N25132, N21419, N22385, N6635);
or OR3 (N25151, N25149, N10137, N20138);
not NOT1 (N25152, N25141);
not NOT1 (N25153, N25147);
and AND3 (N25154, N25144, N15776, N10572);
or OR4 (N25155, N25153, N23013, N16540, N9224);
and AND4 (N25156, N25145, N1005, N2916, N22212);
nand NAND3 (N25157, N25156, N11068, N13409);
buf BUF1 (N25158, N25150);
nand NAND4 (N25159, N25154, N3117, N18157, N10662);
nand NAND3 (N25160, N25138, N3161, N1975);
buf BUF1 (N25161, N25146);
nor NOR4 (N25162, N25157, N2871, N15693, N9515);
xor XOR2 (N25163, N25161, N5775);
or OR4 (N25164, N25160, N18791, N4681, N19555);
xor XOR2 (N25165, N25158, N14538);
buf BUF1 (N25166, N25155);
and AND2 (N25167, N25152, N24724);
buf BUF1 (N25168, N25164);
or OR4 (N25169, N25167, N4545, N9994, N17055);
xor XOR2 (N25170, N25166, N8023);
buf BUF1 (N25171, N25169);
and AND4 (N25172, N25162, N20716, N19301, N9032);
xor XOR2 (N25173, N25159, N7241);
buf BUF1 (N25174, N25171);
nor NOR3 (N25175, N25174, N21348, N12010);
and AND4 (N25176, N25163, N8550, N1838, N7329);
not NOT1 (N25177, N25104);
or OR4 (N25178, N25173, N3108, N24922, N22312);
or OR4 (N25179, N25118, N22146, N10173, N14918);
buf BUF1 (N25180, N25177);
or OR2 (N25181, N25151, N9782);
and AND3 (N25182, N25165, N24515, N12772);
nor NOR2 (N25183, N25181, N25012);
or OR2 (N25184, N25178, N1217);
nor NOR3 (N25185, N25179, N12073, N22900);
and AND2 (N25186, N25172, N2217);
nand NAND3 (N25187, N25186, N4092, N7582);
nor NOR2 (N25188, N25176, N12162);
buf BUF1 (N25189, N25168);
xor XOR2 (N25190, N25183, N21364);
not NOT1 (N25191, N25185);
buf BUF1 (N25192, N25180);
and AND2 (N25193, N25170, N22394);
and AND2 (N25194, N25189, N11232);
buf BUF1 (N25195, N25190);
or OR2 (N25196, N25191, N16901);
or OR2 (N25197, N25187, N18791);
nor NOR3 (N25198, N25196, N17586, N19726);
nand NAND4 (N25199, N25197, N14339, N5098, N18636);
not NOT1 (N25200, N25192);
or OR2 (N25201, N25194, N5453);
or OR2 (N25202, N25182, N21300);
buf BUF1 (N25203, N25200);
nor NOR3 (N25204, N25188, N10763, N6515);
not NOT1 (N25205, N25198);
and AND2 (N25206, N25199, N20446);
and AND2 (N25207, N25206, N14889);
not NOT1 (N25208, N25202);
xor XOR2 (N25209, N25195, N8489);
nor NOR2 (N25210, N25193, N17503);
or OR2 (N25211, N25210, N5904);
xor XOR2 (N25212, N25211, N23062);
xor XOR2 (N25213, N25175, N19877);
or OR3 (N25214, N25203, N21407, N1058);
and AND4 (N25215, N25204, N7343, N9020, N20646);
or OR2 (N25216, N25205, N10735);
nand NAND2 (N25217, N25216, N16335);
nand NAND4 (N25218, N25213, N12567, N7184, N14238);
not NOT1 (N25219, N25217);
nor NOR4 (N25220, N25214, N11172, N5057, N12768);
xor XOR2 (N25221, N25208, N961);
or OR2 (N25222, N25212, N1284);
xor XOR2 (N25223, N25221, N2471);
buf BUF1 (N25224, N25215);
xor XOR2 (N25225, N25222, N20135);
not NOT1 (N25226, N25224);
or OR2 (N25227, N25207, N24592);
not NOT1 (N25228, N25201);
or OR2 (N25229, N25218, N18997);
xor XOR2 (N25230, N25228, N22400);
or OR2 (N25231, N25227, N8537);
nand NAND2 (N25232, N25220, N24780);
not NOT1 (N25233, N25184);
xor XOR2 (N25234, N25232, N2940);
buf BUF1 (N25235, N25226);
buf BUF1 (N25236, N25234);
not NOT1 (N25237, N25231);
xor XOR2 (N25238, N25235, N6338);
buf BUF1 (N25239, N25223);
xor XOR2 (N25240, N25238, N6586);
or OR2 (N25241, N25225, N17337);
nor NOR2 (N25242, N25233, N18101);
and AND2 (N25243, N25240, N23339);
not NOT1 (N25244, N25230);
xor XOR2 (N25245, N25241, N6758);
nor NOR2 (N25246, N25219, N12422);
xor XOR2 (N25247, N25246, N11212);
and AND3 (N25248, N25209, N1805, N2741);
nor NOR3 (N25249, N25247, N14523, N11088);
nand NAND2 (N25250, N25249, N16015);
xor XOR2 (N25251, N25236, N10768);
and AND3 (N25252, N25242, N4988, N2118);
nor NOR4 (N25253, N25237, N12531, N24610, N8600);
nor NOR4 (N25254, N25250, N18109, N3359, N11397);
nand NAND2 (N25255, N25239, N13315);
xor XOR2 (N25256, N25229, N21223);
not NOT1 (N25257, N25248);
or OR4 (N25258, N25252, N24506, N12920, N2464);
or OR3 (N25259, N25245, N12906, N9367);
not NOT1 (N25260, N25244);
nor NOR3 (N25261, N25254, N20202, N15263);
buf BUF1 (N25262, N25257);
xor XOR2 (N25263, N25255, N14785);
nor NOR3 (N25264, N25258, N8101, N3187);
buf BUF1 (N25265, N25260);
nor NOR4 (N25266, N25253, N16258, N11336, N10927);
buf BUF1 (N25267, N25263);
nand NAND3 (N25268, N25259, N11985, N1063);
nand NAND2 (N25269, N25251, N25205);
buf BUF1 (N25270, N25269);
and AND3 (N25271, N25256, N23380, N14383);
not NOT1 (N25272, N25270);
buf BUF1 (N25273, N25264);
and AND3 (N25274, N25272, N9849, N14200);
or OR4 (N25275, N25273, N11176, N9155, N23834);
buf BUF1 (N25276, N25243);
nor NOR4 (N25277, N25265, N17453, N23591, N21557);
and AND4 (N25278, N25274, N6205, N9212, N3265);
and AND2 (N25279, N25276, N10469);
not NOT1 (N25280, N25261);
xor XOR2 (N25281, N25267, N16495);
buf BUF1 (N25282, N25280);
nand NAND4 (N25283, N25266, N2919, N6287, N18400);
or OR3 (N25284, N25279, N5081, N9514);
or OR4 (N25285, N25275, N19794, N3537, N9412);
not NOT1 (N25286, N25278);
buf BUF1 (N25287, N25271);
not NOT1 (N25288, N25287);
xor XOR2 (N25289, N25277, N23740);
nand NAND3 (N25290, N25282, N14761, N12402);
or OR4 (N25291, N25283, N8034, N2959, N13070);
or OR3 (N25292, N25289, N20508, N15187);
buf BUF1 (N25293, N25284);
not NOT1 (N25294, N25290);
not NOT1 (N25295, N25291);
buf BUF1 (N25296, N25262);
or OR2 (N25297, N25286, N21273);
or OR3 (N25298, N25295, N8891, N4842);
not NOT1 (N25299, N25293);
nor NOR3 (N25300, N25294, N18189, N6781);
buf BUF1 (N25301, N25285);
not NOT1 (N25302, N25296);
xor XOR2 (N25303, N25298, N16116);
buf BUF1 (N25304, N25303);
nand NAND2 (N25305, N25288, N20489);
or OR4 (N25306, N25281, N7136, N22170, N17953);
or OR3 (N25307, N25301, N4534, N20647);
xor XOR2 (N25308, N25304, N7527);
and AND3 (N25309, N25268, N23194, N7268);
nor NOR3 (N25310, N25300, N12021, N25274);
and AND4 (N25311, N25309, N4665, N1384, N4138);
not NOT1 (N25312, N25306);
xor XOR2 (N25313, N25292, N9879);
nand NAND3 (N25314, N25308, N24549, N22382);
buf BUF1 (N25315, N25314);
or OR4 (N25316, N25299, N5246, N9644, N5491);
and AND2 (N25317, N25297, N20047);
buf BUF1 (N25318, N25310);
or OR2 (N25319, N25307, N17318);
nand NAND3 (N25320, N25312, N12513, N23213);
not NOT1 (N25321, N25316);
nor NOR2 (N25322, N25319, N1827);
and AND2 (N25323, N25302, N19212);
buf BUF1 (N25324, N25305);
and AND2 (N25325, N25311, N1290);
nand NAND4 (N25326, N25320, N4974, N19489, N6888);
not NOT1 (N25327, N25322);
buf BUF1 (N25328, N25318);
or OR3 (N25329, N25325, N306, N11177);
and AND3 (N25330, N25329, N932, N25324);
nand NAND3 (N25331, N15517, N7894, N4194);
buf BUF1 (N25332, N25328);
or OR2 (N25333, N25332, N19632);
not NOT1 (N25334, N25315);
buf BUF1 (N25335, N25327);
not NOT1 (N25336, N25334);
not NOT1 (N25337, N25333);
nand NAND4 (N25338, N25317, N21293, N4842, N24548);
xor XOR2 (N25339, N25313, N2272);
or OR4 (N25340, N25337, N14908, N19048, N329);
or OR4 (N25341, N25335, N14911, N11992, N5603);
not NOT1 (N25342, N25338);
nor NOR4 (N25343, N25340, N23448, N10824, N12472);
not NOT1 (N25344, N25330);
and AND4 (N25345, N25342, N18104, N9880, N11914);
nor NOR4 (N25346, N25321, N20776, N7800, N6288);
nor NOR4 (N25347, N25336, N15971, N25043, N7036);
nand NAND4 (N25348, N25346, N16403, N23815, N7915);
buf BUF1 (N25349, N25331);
not NOT1 (N25350, N25347);
xor XOR2 (N25351, N25350, N19444);
buf BUF1 (N25352, N25343);
nor NOR3 (N25353, N25345, N2855, N14004);
nor NOR3 (N25354, N25351, N10356, N19771);
nor NOR4 (N25355, N25341, N24496, N15775, N4791);
and AND2 (N25356, N25348, N8185);
not NOT1 (N25357, N25356);
and AND2 (N25358, N25354, N23070);
nand NAND2 (N25359, N25355, N7749);
not NOT1 (N25360, N25349);
not NOT1 (N25361, N25344);
nor NOR4 (N25362, N25360, N21037, N16691, N7556);
xor XOR2 (N25363, N25352, N22235);
buf BUF1 (N25364, N25363);
xor XOR2 (N25365, N25326, N10365);
buf BUF1 (N25366, N25365);
and AND2 (N25367, N25358, N21028);
and AND2 (N25368, N25367, N19352);
nor NOR3 (N25369, N25368, N11004, N1297);
nor NOR3 (N25370, N25362, N8317, N22134);
buf BUF1 (N25371, N25366);
nor NOR4 (N25372, N25357, N19478, N20059, N12062);
and AND2 (N25373, N25339, N13048);
nor NOR2 (N25374, N25370, N22048);
buf BUF1 (N25375, N25323);
or OR4 (N25376, N25359, N15463, N23578, N16191);
or OR2 (N25377, N25374, N14021);
xor XOR2 (N25378, N25377, N1546);
nor NOR3 (N25379, N25373, N22606, N4424);
nor NOR3 (N25380, N25364, N11931, N13325);
nand NAND4 (N25381, N25376, N18226, N11936, N12319);
not NOT1 (N25382, N25379);
buf BUF1 (N25383, N25380);
nor NOR2 (N25384, N25372, N606);
or OR4 (N25385, N25375, N24552, N16804, N13453);
nand NAND4 (N25386, N25384, N6674, N24407, N13341);
buf BUF1 (N25387, N25378);
buf BUF1 (N25388, N25361);
or OR4 (N25389, N25386, N22712, N10930, N24058);
buf BUF1 (N25390, N25383);
nor NOR3 (N25391, N25390, N1550, N194);
and AND4 (N25392, N25369, N11724, N14372, N2618);
not NOT1 (N25393, N25381);
nor NOR4 (N25394, N25392, N20354, N15201, N22612);
and AND3 (N25395, N25387, N10967, N15787);
xor XOR2 (N25396, N25395, N16013);
xor XOR2 (N25397, N25389, N23150);
xor XOR2 (N25398, N25394, N1484);
xor XOR2 (N25399, N25391, N19413);
or OR2 (N25400, N25353, N8505);
and AND4 (N25401, N25398, N25326, N14109, N18126);
xor XOR2 (N25402, N25385, N20033);
not NOT1 (N25403, N25396);
nor NOR2 (N25404, N25382, N4146);
buf BUF1 (N25405, N25400);
xor XOR2 (N25406, N25401, N16591);
nor NOR3 (N25407, N25399, N16879, N21528);
not NOT1 (N25408, N25404);
nor NOR4 (N25409, N25402, N9950, N16605, N24381);
and AND3 (N25410, N25406, N14146, N17506);
or OR2 (N25411, N25409, N3236);
nand NAND2 (N25412, N25397, N8157);
nand NAND2 (N25413, N25393, N23235);
buf BUF1 (N25414, N25410);
or OR2 (N25415, N25408, N15947);
nor NOR3 (N25416, N25415, N3215, N19527);
or OR2 (N25417, N25411, N22810);
nand NAND4 (N25418, N25412, N20515, N25388, N7754);
nor NOR3 (N25419, N8506, N21208, N19656);
and AND4 (N25420, N25417, N10064, N10706, N19142);
nor NOR2 (N25421, N25420, N23445);
not NOT1 (N25422, N25416);
and AND3 (N25423, N25405, N10382, N4636);
or OR4 (N25424, N25403, N7117, N20952, N8697);
nor NOR3 (N25425, N25423, N20372, N2849);
nor NOR3 (N25426, N25421, N12454, N665);
nor NOR3 (N25427, N25426, N1634, N4364);
xor XOR2 (N25428, N25414, N3162);
or OR3 (N25429, N25371, N3201, N12498);
buf BUF1 (N25430, N25407);
nor NOR3 (N25431, N25424, N7876, N310);
nand NAND4 (N25432, N25413, N14238, N14911, N6550);
buf BUF1 (N25433, N25419);
not NOT1 (N25434, N25425);
or OR4 (N25435, N25427, N867, N13829, N21240);
xor XOR2 (N25436, N25434, N14026);
buf BUF1 (N25437, N25430);
nand NAND4 (N25438, N25429, N10675, N19401, N13992);
not NOT1 (N25439, N25436);
buf BUF1 (N25440, N25433);
and AND2 (N25441, N25437, N22601);
nand NAND3 (N25442, N25418, N16633, N103);
nor NOR2 (N25443, N25440, N21477);
not NOT1 (N25444, N25443);
xor XOR2 (N25445, N25435, N22085);
xor XOR2 (N25446, N25438, N19762);
buf BUF1 (N25447, N25439);
nor NOR2 (N25448, N25431, N7080);
not NOT1 (N25449, N25444);
buf BUF1 (N25450, N25447);
not NOT1 (N25451, N25448);
or OR4 (N25452, N25442, N14139, N18926, N1211);
not NOT1 (N25453, N25422);
xor XOR2 (N25454, N25446, N16445);
nor NOR4 (N25455, N25451, N17183, N9560, N12413);
not NOT1 (N25456, N25445);
xor XOR2 (N25457, N25441, N21409);
xor XOR2 (N25458, N25452, N15549);
nor NOR3 (N25459, N25428, N25034, N3178);
xor XOR2 (N25460, N25459, N17796);
and AND2 (N25461, N25453, N14662);
nand NAND2 (N25462, N25454, N20560);
nor NOR4 (N25463, N25457, N18182, N13767, N5584);
nor NOR2 (N25464, N25432, N620);
or OR3 (N25465, N25458, N16892, N6401);
buf BUF1 (N25466, N25461);
xor XOR2 (N25467, N25460, N10622);
buf BUF1 (N25468, N25464);
or OR4 (N25469, N25450, N9017, N22129, N8565);
nor NOR3 (N25470, N25463, N182, N7050);
not NOT1 (N25471, N25467);
nor NOR3 (N25472, N25462, N5423, N2350);
or OR2 (N25473, N25469, N15884);
buf BUF1 (N25474, N25468);
not NOT1 (N25475, N25472);
buf BUF1 (N25476, N25466);
and AND3 (N25477, N25456, N18706, N1334);
nand NAND3 (N25478, N25449, N3698, N23628);
nor NOR3 (N25479, N25470, N22734, N24677);
nor NOR2 (N25480, N25471, N8201);
buf BUF1 (N25481, N25478);
buf BUF1 (N25482, N25465);
and AND4 (N25483, N25477, N18163, N8540, N14209);
nor NOR3 (N25484, N25455, N4018, N24193);
nand NAND3 (N25485, N25482, N6376, N13091);
buf BUF1 (N25486, N25481);
nor NOR2 (N25487, N25484, N18691);
nor NOR3 (N25488, N25483, N22346, N21521);
or OR4 (N25489, N25479, N2313, N23758, N11871);
or OR3 (N25490, N25485, N10732, N3027);
xor XOR2 (N25491, N25489, N9462);
xor XOR2 (N25492, N25473, N6028);
nor NOR3 (N25493, N25475, N3455, N19118);
not NOT1 (N25494, N25493);
and AND2 (N25495, N25490, N13772);
xor XOR2 (N25496, N25480, N25155);
and AND2 (N25497, N25495, N19403);
and AND2 (N25498, N25476, N16439);
buf BUF1 (N25499, N25494);
nand NAND4 (N25500, N25497, N13101, N18772, N16541);
and AND2 (N25501, N25498, N4709);
and AND2 (N25502, N25488, N12655);
not NOT1 (N25503, N25499);
and AND4 (N25504, N25474, N7597, N23676, N13718);
nand NAND4 (N25505, N25504, N4860, N22142, N16114);
nor NOR4 (N25506, N25505, N5037, N2114, N7437);
nand NAND4 (N25507, N25501, N12926, N6725, N25334);
xor XOR2 (N25508, N25502, N1690);
and AND4 (N25509, N25496, N19057, N1612, N20642);
nor NOR2 (N25510, N25491, N22080);
or OR4 (N25511, N25510, N19056, N7297, N17369);
nand NAND3 (N25512, N25500, N14168, N19458);
nand NAND2 (N25513, N25511, N2430);
and AND3 (N25514, N25486, N4786, N15048);
not NOT1 (N25515, N25487);
or OR3 (N25516, N25513, N414, N18836);
and AND3 (N25517, N25515, N23032, N20730);
buf BUF1 (N25518, N25508);
xor XOR2 (N25519, N25492, N4646);
xor XOR2 (N25520, N25509, N14174);
nor NOR2 (N25521, N25512, N1688);
or OR4 (N25522, N25506, N8784, N12422, N10622);
nor NOR2 (N25523, N25521, N20661);
not NOT1 (N25524, N25522);
and AND4 (N25525, N25523, N22703, N21358, N9483);
and AND3 (N25526, N25517, N22981, N17161);
and AND4 (N25527, N25514, N13921, N22228, N21930);
nor NOR2 (N25528, N25507, N9820);
buf BUF1 (N25529, N25525);
and AND4 (N25530, N25529, N7606, N17569, N8345);
buf BUF1 (N25531, N25524);
xor XOR2 (N25532, N25531, N3857);
nand NAND3 (N25533, N25519, N4995, N25122);
not NOT1 (N25534, N25526);
not NOT1 (N25535, N25520);
not NOT1 (N25536, N25503);
and AND3 (N25537, N25527, N1533, N20384);
and AND2 (N25538, N25537, N22715);
or OR4 (N25539, N25530, N1622, N1900, N4857);
xor XOR2 (N25540, N25539, N14257);
xor XOR2 (N25541, N25535, N1374);
xor XOR2 (N25542, N25518, N10563);
nand NAND4 (N25543, N25540, N22193, N24407, N3968);
nor NOR3 (N25544, N25542, N16062, N22699);
buf BUF1 (N25545, N25528);
or OR2 (N25546, N25536, N10941);
not NOT1 (N25547, N25541);
nor NOR2 (N25548, N25544, N17964);
nand NAND2 (N25549, N25545, N1340);
or OR2 (N25550, N25532, N17416);
or OR4 (N25551, N25550, N22834, N22434, N22697);
and AND2 (N25552, N25543, N19180);
xor XOR2 (N25553, N25549, N22680);
and AND2 (N25554, N25534, N1122);
nand NAND2 (N25555, N25533, N9784);
buf BUF1 (N25556, N25553);
not NOT1 (N25557, N25551);
nand NAND3 (N25558, N25538, N5615, N22228);
nor NOR3 (N25559, N25552, N25046, N6745);
and AND4 (N25560, N25546, N1435, N19383, N4217);
nand NAND3 (N25561, N25557, N14728, N11659);
or OR2 (N25562, N25560, N24127);
and AND3 (N25563, N25548, N12294, N942);
and AND3 (N25564, N25556, N19784, N21261);
nor NOR4 (N25565, N25561, N8166, N1858, N13126);
and AND3 (N25566, N25554, N16426, N7979);
and AND2 (N25567, N25563, N9180);
not NOT1 (N25568, N25565);
nor NOR3 (N25569, N25516, N24209, N5891);
and AND2 (N25570, N25559, N8170);
not NOT1 (N25571, N25558);
nand NAND2 (N25572, N25547, N21823);
nand NAND3 (N25573, N25570, N8902, N24837);
not NOT1 (N25574, N25567);
not NOT1 (N25575, N25562);
buf BUF1 (N25576, N25564);
and AND4 (N25577, N25573, N17527, N3643, N19166);
nand NAND4 (N25578, N25577, N23324, N6194, N14805);
and AND4 (N25579, N25568, N12436, N9536, N14297);
nor NOR3 (N25580, N25574, N15976, N14283);
xor XOR2 (N25581, N25555, N15509);
xor XOR2 (N25582, N25576, N8834);
not NOT1 (N25583, N25572);
or OR2 (N25584, N25582, N18202);
xor XOR2 (N25585, N25575, N22578);
or OR4 (N25586, N25580, N1948, N20512, N1586);
not NOT1 (N25587, N25566);
and AND3 (N25588, N25583, N4802, N6687);
nand NAND2 (N25589, N25585, N24337);
not NOT1 (N25590, N25587);
xor XOR2 (N25591, N25581, N9308);
buf BUF1 (N25592, N25588);
buf BUF1 (N25593, N25571);
buf BUF1 (N25594, N25590);
or OR4 (N25595, N25592, N10139, N14329, N461);
nor NOR2 (N25596, N25589, N18191);
and AND4 (N25597, N25584, N10389, N7259, N25101);
or OR3 (N25598, N25578, N18091, N17421);
not NOT1 (N25599, N25597);
and AND4 (N25600, N25595, N6950, N12802, N13709);
nor NOR2 (N25601, N25598, N14252);
nor NOR3 (N25602, N25591, N9399, N22158);
buf BUF1 (N25603, N25594);
xor XOR2 (N25604, N25600, N4735);
nor NOR3 (N25605, N25602, N24139, N14652);
xor XOR2 (N25606, N25603, N4554);
and AND4 (N25607, N25605, N18370, N15605, N1686);
not NOT1 (N25608, N25593);
nand NAND2 (N25609, N25596, N9485);
nor NOR2 (N25610, N25579, N4267);
nor NOR3 (N25611, N25586, N13138, N10464);
nor NOR2 (N25612, N25608, N5219);
nand NAND3 (N25613, N25610, N12902, N25219);
or OR4 (N25614, N25609, N12065, N23501, N13066);
or OR4 (N25615, N25599, N14678, N11227, N21291);
not NOT1 (N25616, N25606);
buf BUF1 (N25617, N25604);
xor XOR2 (N25618, N25607, N8789);
xor XOR2 (N25619, N25616, N25603);
endmodule