// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19;

output N380,N415,N403,N407,N405,N412,N411,N389,N418,N419;

buf BUF1 (N20, N9);
xor XOR2 (N21, N19, N3);
nand NAND4 (N22, N16, N17, N3, N18);
and AND2 (N23, N9, N21);
and AND2 (N24, N4, N7);
not NOT1 (N25, N17);
and AND4 (N26, N4, N19, N1, N22);
or OR4 (N27, N24, N6, N11, N22);
nand NAND4 (N28, N7, N16, N14, N8);
buf BUF1 (N29, N1);
nor NOR2 (N30, N26, N9);
buf BUF1 (N31, N26);
nand NAND2 (N32, N2, N10);
not NOT1 (N33, N18);
nand NAND4 (N34, N33, N1, N33, N30);
buf BUF1 (N35, N26);
not NOT1 (N36, N32);
xor XOR2 (N37, N25, N17);
buf BUF1 (N38, N35);
nand NAND2 (N39, N20, N33);
nand NAND3 (N40, N38, N11, N20);
not NOT1 (N41, N37);
or OR4 (N42, N31, N32, N11, N39);
nor NOR4 (N43, N6, N32, N21, N38);
xor XOR2 (N44, N28, N3);
nor NOR2 (N45, N41, N3);
xor XOR2 (N46, N27, N8);
xor XOR2 (N47, N23, N21);
xor XOR2 (N48, N40, N42);
nand NAND2 (N49, N34, N33);
buf BUF1 (N50, N22);
or OR3 (N51, N50, N44, N22);
not NOT1 (N52, N49);
or OR2 (N53, N6, N44);
buf BUF1 (N54, N46);
and AND4 (N55, N53, N36, N52, N17);
nand NAND4 (N56, N3, N13, N3, N41);
nor NOR2 (N57, N48, N24);
nor NOR4 (N58, N4, N1, N26, N28);
not NOT1 (N59, N55);
nor NOR3 (N60, N47, N42, N21);
nor NOR3 (N61, N43, N15, N25);
not NOT1 (N62, N59);
not NOT1 (N63, N29);
not NOT1 (N64, N62);
buf BUF1 (N65, N51);
nand NAND4 (N66, N64, N3, N63, N49);
nand NAND4 (N67, N39, N42, N20, N10);
not NOT1 (N68, N66);
not NOT1 (N69, N58);
not NOT1 (N70, N68);
and AND3 (N71, N61, N25, N32);
and AND3 (N72, N45, N51, N28);
not NOT1 (N73, N56);
not NOT1 (N74, N57);
buf BUF1 (N75, N72);
nand NAND3 (N76, N54, N1, N50);
nor NOR3 (N77, N75, N17, N35);
and AND3 (N78, N70, N42, N42);
xor XOR2 (N79, N77, N55);
and AND3 (N80, N74, N19, N74);
and AND2 (N81, N80, N23);
not NOT1 (N82, N69);
nand NAND2 (N83, N78, N35);
not NOT1 (N84, N82);
not NOT1 (N85, N60);
xor XOR2 (N86, N76, N30);
buf BUF1 (N87, N73);
nand NAND4 (N88, N79, N46, N75, N23);
xor XOR2 (N89, N85, N11);
not NOT1 (N90, N71);
nand NAND2 (N91, N90, N49);
xor XOR2 (N92, N86, N56);
xor XOR2 (N93, N84, N38);
nand NAND3 (N94, N92, N30, N2);
nand NAND2 (N95, N89, N82);
or OR4 (N96, N95, N85, N86, N38);
buf BUF1 (N97, N91);
or OR3 (N98, N96, N28, N18);
not NOT1 (N99, N81);
not NOT1 (N100, N83);
or OR4 (N101, N65, N30, N69, N22);
nor NOR4 (N102, N101, N46, N41, N6);
not NOT1 (N103, N88);
not NOT1 (N104, N94);
not NOT1 (N105, N87);
nor NOR2 (N106, N97, N93);
xor XOR2 (N107, N94, N104);
nand NAND3 (N108, N96, N95, N97);
nand NAND2 (N109, N102, N106);
or OR3 (N110, N67, N52, N60);
nand NAND2 (N111, N23, N30);
or OR2 (N112, N100, N70);
xor XOR2 (N113, N111, N69);
not NOT1 (N114, N105);
xor XOR2 (N115, N98, N89);
not NOT1 (N116, N110);
or OR2 (N117, N115, N82);
buf BUF1 (N118, N109);
or OR3 (N119, N99, N101, N59);
and AND4 (N120, N118, N119, N99, N113);
and AND2 (N121, N21, N96);
not NOT1 (N122, N107);
xor XOR2 (N123, N35, N28);
nand NAND2 (N124, N114, N63);
and AND4 (N125, N112, N63, N17, N88);
nand NAND4 (N126, N116, N12, N117, N20);
nand NAND3 (N127, N77, N113, N5);
buf BUF1 (N128, N121);
nand NAND4 (N129, N123, N37, N26, N68);
and AND2 (N130, N129, N22);
or OR4 (N131, N124, N11, N107, N3);
and AND2 (N132, N122, N112);
buf BUF1 (N133, N126);
not NOT1 (N134, N103);
buf BUF1 (N135, N130);
or OR2 (N136, N125, N114);
xor XOR2 (N137, N136, N101);
buf BUF1 (N138, N108);
and AND3 (N139, N137, N115, N69);
nor NOR2 (N140, N133, N34);
buf BUF1 (N141, N138);
nand NAND2 (N142, N128, N82);
xor XOR2 (N143, N127, N32);
not NOT1 (N144, N139);
or OR3 (N145, N131, N50, N47);
buf BUF1 (N146, N132);
and AND2 (N147, N144, N68);
and AND4 (N148, N135, N50, N50, N19);
and AND4 (N149, N147, N118, N143, N4);
buf BUF1 (N150, N60);
nor NOR4 (N151, N141, N147, N145, N91);
nand NAND3 (N152, N78, N7, N140);
nand NAND4 (N153, N35, N133, N73, N78);
and AND3 (N154, N149, N132, N77);
and AND2 (N155, N151, N66);
nor NOR3 (N156, N154, N38, N62);
buf BUF1 (N157, N156);
not NOT1 (N158, N155);
xor XOR2 (N159, N148, N151);
and AND2 (N160, N152, N137);
nor NOR4 (N161, N153, N14, N66, N107);
and AND3 (N162, N158, N80, N5);
or OR4 (N163, N161, N156, N71, N60);
nor NOR2 (N164, N134, N36);
and AND2 (N165, N142, N140);
xor XOR2 (N166, N150, N132);
or OR2 (N167, N157, N146);
nand NAND3 (N168, N26, N71, N129);
not NOT1 (N169, N160);
not NOT1 (N170, N163);
or OR4 (N171, N165, N94, N62, N152);
or OR4 (N172, N168, N4, N24, N25);
nor NOR4 (N173, N167, N117, N141, N160);
nor NOR3 (N174, N162, N146, N128);
xor XOR2 (N175, N120, N48);
and AND3 (N176, N172, N114, N70);
xor XOR2 (N177, N159, N133);
buf BUF1 (N178, N166);
or OR4 (N179, N169, N101, N98, N160);
buf BUF1 (N180, N174);
and AND3 (N181, N175, N126, N41);
nand NAND4 (N182, N176, N158, N14, N80);
and AND2 (N183, N179, N142);
nand NAND2 (N184, N173, N139);
and AND2 (N185, N164, N133);
or OR3 (N186, N171, N16, N58);
buf BUF1 (N187, N178);
nor NOR4 (N188, N177, N98, N4, N117);
nor NOR3 (N189, N186, N154, N33);
xor XOR2 (N190, N180, N164);
not NOT1 (N191, N170);
not NOT1 (N192, N181);
buf BUF1 (N193, N190);
and AND3 (N194, N185, N65, N90);
xor XOR2 (N195, N184, N138);
buf BUF1 (N196, N182);
nand NAND2 (N197, N193, N52);
nand NAND3 (N198, N191, N66, N189);
and AND2 (N199, N190, N85);
xor XOR2 (N200, N198, N90);
not NOT1 (N201, N195);
or OR4 (N202, N201, N74, N110, N133);
nand NAND3 (N203, N200, N100, N48);
nand NAND4 (N204, N183, N119, N144, N101);
buf BUF1 (N205, N204);
and AND4 (N206, N203, N50, N17, N201);
not NOT1 (N207, N194);
or OR3 (N208, N192, N52, N30);
nand NAND4 (N209, N187, N131, N90, N203);
nand NAND3 (N210, N188, N130, N83);
or OR2 (N211, N209, N64);
xor XOR2 (N212, N205, N78);
not NOT1 (N213, N208);
nand NAND4 (N214, N206, N98, N116, N167);
and AND4 (N215, N213, N189, N183, N210);
buf BUF1 (N216, N53);
xor XOR2 (N217, N211, N7);
nand NAND2 (N218, N197, N131);
buf BUF1 (N219, N217);
not NOT1 (N220, N196);
xor XOR2 (N221, N214, N32);
buf BUF1 (N222, N212);
nor NOR2 (N223, N215, N106);
or OR4 (N224, N219, N69, N178, N146);
or OR3 (N225, N222, N127, N170);
buf BUF1 (N226, N220);
and AND4 (N227, N226, N39, N217, N124);
nor NOR4 (N228, N199, N193, N12, N130);
not NOT1 (N229, N207);
not NOT1 (N230, N228);
nor NOR4 (N231, N227, N2, N69, N148);
and AND4 (N232, N229, N109, N64, N63);
nand NAND3 (N233, N221, N147, N128);
nand NAND4 (N234, N224, N60, N100, N92);
or OR3 (N235, N225, N68, N214);
and AND4 (N236, N235, N120, N176, N49);
xor XOR2 (N237, N218, N93);
buf BUF1 (N238, N223);
nor NOR2 (N239, N232, N105);
not NOT1 (N240, N239);
buf BUF1 (N241, N237);
nor NOR4 (N242, N216, N226, N197, N51);
or OR4 (N243, N242, N77, N135, N234);
and AND4 (N244, N89, N74, N93, N144);
not NOT1 (N245, N231);
nand NAND2 (N246, N230, N15);
nor NOR2 (N247, N240, N20);
xor XOR2 (N248, N241, N44);
and AND4 (N249, N245, N190, N75, N1);
xor XOR2 (N250, N247, N248);
buf BUF1 (N251, N187);
nand NAND4 (N252, N246, N223, N83, N246);
not NOT1 (N253, N250);
and AND4 (N254, N202, N82, N171, N200);
and AND3 (N255, N253, N93, N67);
nor NOR2 (N256, N254, N84);
buf BUF1 (N257, N233);
xor XOR2 (N258, N256, N126);
nand NAND4 (N259, N244, N228, N206, N31);
nand NAND2 (N260, N259, N191);
nor NOR3 (N261, N243, N133, N216);
or OR3 (N262, N258, N207, N135);
not NOT1 (N263, N260);
nand NAND2 (N264, N261, N204);
buf BUF1 (N265, N249);
nand NAND4 (N266, N255, N134, N260, N152);
or OR2 (N267, N262, N180);
not NOT1 (N268, N257);
or OR4 (N269, N266, N225, N115, N31);
buf BUF1 (N270, N264);
nand NAND2 (N271, N270, N163);
and AND4 (N272, N269, N67, N182, N74);
and AND2 (N273, N265, N140);
nand NAND4 (N274, N268, N270, N69, N228);
not NOT1 (N275, N272);
or OR3 (N276, N263, N262, N124);
nand NAND2 (N277, N276, N179);
nor NOR4 (N278, N252, N260, N47, N103);
xor XOR2 (N279, N267, N5);
xor XOR2 (N280, N279, N225);
buf BUF1 (N281, N251);
not NOT1 (N282, N238);
not NOT1 (N283, N278);
buf BUF1 (N284, N280);
nor NOR3 (N285, N284, N178, N276);
nand NAND3 (N286, N275, N20, N102);
or OR2 (N287, N273, N169);
buf BUF1 (N288, N287);
xor XOR2 (N289, N281, N29);
xor XOR2 (N290, N236, N271);
buf BUF1 (N291, N38);
xor XOR2 (N292, N282, N230);
and AND2 (N293, N283, N131);
not NOT1 (N294, N285);
nor NOR4 (N295, N294, N137, N263, N141);
not NOT1 (N296, N289);
or OR4 (N297, N290, N245, N123, N295);
buf BUF1 (N298, N287);
nor NOR4 (N299, N292, N212, N126, N89);
xor XOR2 (N300, N286, N11);
and AND2 (N301, N297, N43);
and AND4 (N302, N296, N146, N301, N88);
xor XOR2 (N303, N293, N247);
buf BUF1 (N304, N21);
and AND3 (N305, N291, N166, N177);
not NOT1 (N306, N298);
or OR3 (N307, N288, N127, N44);
and AND2 (N308, N300, N88);
and AND2 (N309, N299, N135);
buf BUF1 (N310, N303);
xor XOR2 (N311, N274, N271);
xor XOR2 (N312, N306, N233);
and AND2 (N313, N307, N148);
not NOT1 (N314, N309);
nor NOR4 (N315, N312, N3, N121, N255);
nand NAND3 (N316, N277, N116, N222);
buf BUF1 (N317, N305);
and AND3 (N318, N304, N34, N155);
nand NAND2 (N319, N317, N174);
nor NOR2 (N320, N319, N6);
and AND2 (N321, N315, N211);
buf BUF1 (N322, N316);
or OR4 (N323, N308, N187, N41, N310);
or OR2 (N324, N140, N108);
buf BUF1 (N325, N322);
nor NOR3 (N326, N320, N28, N110);
or OR4 (N327, N318, N198, N30, N118);
not NOT1 (N328, N302);
buf BUF1 (N329, N327);
nand NAND4 (N330, N311, N247, N2, N107);
xor XOR2 (N331, N324, N229);
nand NAND3 (N332, N326, N7, N204);
nor NOR2 (N333, N323, N118);
or OR4 (N334, N321, N65, N296, N105);
not NOT1 (N335, N333);
nand NAND2 (N336, N314, N292);
xor XOR2 (N337, N328, N151);
nor NOR3 (N338, N330, N146, N279);
xor XOR2 (N339, N337, N242);
xor XOR2 (N340, N331, N146);
or OR2 (N341, N336, N61);
nand NAND3 (N342, N338, N288, N190);
nor NOR4 (N343, N335, N35, N216, N212);
and AND2 (N344, N339, N255);
nor NOR4 (N345, N341, N334, N146, N200);
buf BUF1 (N346, N138);
nor NOR3 (N347, N342, N65, N10);
buf BUF1 (N348, N345);
xor XOR2 (N349, N340, N280);
and AND4 (N350, N313, N83, N99, N66);
nor NOR4 (N351, N344, N93, N61, N193);
buf BUF1 (N352, N349);
and AND4 (N353, N347, N240, N263, N144);
or OR2 (N354, N352, N335);
nor NOR3 (N355, N348, N43, N212);
xor XOR2 (N356, N350, N232);
or OR2 (N357, N329, N80);
not NOT1 (N358, N353);
nor NOR2 (N359, N355, N62);
buf BUF1 (N360, N325);
or OR2 (N361, N343, N260);
not NOT1 (N362, N360);
nor NOR2 (N363, N361, N152);
nand NAND4 (N364, N358, N121, N287, N339);
or OR3 (N365, N356, N124, N103);
nand NAND3 (N366, N365, N18, N220);
xor XOR2 (N367, N364, N92);
nor NOR2 (N368, N359, N78);
xor XOR2 (N369, N368, N164);
nor NOR2 (N370, N363, N98);
xor XOR2 (N371, N332, N144);
nand NAND2 (N372, N346, N23);
or OR2 (N373, N357, N109);
not NOT1 (N374, N351);
xor XOR2 (N375, N367, N225);
nand NAND2 (N376, N354, N50);
nand NAND4 (N377, N374, N2, N21, N126);
or OR2 (N378, N376, N290);
or OR4 (N379, N371, N87, N216, N336);
nand NAND2 (N380, N377, N362);
buf BUF1 (N381, N108);
nand NAND3 (N382, N375, N14, N67);
nor NOR2 (N383, N370, N226);
nor NOR3 (N384, N373, N292, N92);
nor NOR3 (N385, N384, N109, N258);
xor XOR2 (N386, N379, N312);
nor NOR2 (N387, N381, N324);
not NOT1 (N388, N387);
or OR4 (N389, N388, N37, N35, N282);
or OR4 (N390, N386, N371, N295, N62);
nor NOR4 (N391, N390, N317, N194, N115);
or OR3 (N392, N369, N245, N68);
and AND2 (N393, N383, N219);
buf BUF1 (N394, N378);
or OR2 (N395, N382, N33);
xor XOR2 (N396, N385, N115);
xor XOR2 (N397, N391, N363);
buf BUF1 (N398, N396);
nor NOR4 (N399, N398, N146, N136, N175);
nor NOR4 (N400, N393, N186, N340, N227);
not NOT1 (N401, N372);
buf BUF1 (N402, N401);
not NOT1 (N403, N399);
not NOT1 (N404, N402);
xor XOR2 (N405, N400, N280);
and AND3 (N406, N366, N58, N231);
xor XOR2 (N407, N406, N143);
not NOT1 (N408, N395);
nand NAND4 (N409, N397, N307, N283, N352);
or OR4 (N410, N409, N58, N193, N106);
not NOT1 (N411, N404);
or OR4 (N412, N392, N31, N410, N171);
xor XOR2 (N413, N317, N31);
nand NAND2 (N414, N413, N291);
nand NAND4 (N415, N414, N160, N278, N123);
xor XOR2 (N416, N394, N259);
not NOT1 (N417, N408);
nor NOR3 (N418, N417, N67, N77);
buf BUF1 (N419, N416);
endmodule