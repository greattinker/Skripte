// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10;

output N2001,N1996,N2008,N2004,N1990,N1999,N2006,N2003,N2007,N2010;

nand NAND2 (N11, N9, N1);
buf BUF1 (N12, N6);
buf BUF1 (N13, N12);
nor NOR4 (N14, N3, N10, N7, N3);
nand NAND2 (N15, N11, N3);
xor XOR2 (N16, N1, N9);
and AND3 (N17, N9, N11, N10);
not NOT1 (N18, N3);
not NOT1 (N19, N1);
nor NOR2 (N20, N9, N19);
not NOT1 (N21, N2);
xor XOR2 (N22, N15, N4);
nor NOR3 (N23, N3, N3, N13);
or OR3 (N24, N16, N10, N9);
xor XOR2 (N25, N17, N22);
or OR2 (N26, N20, N8);
nand NAND3 (N27, N12, N19, N2);
not NOT1 (N28, N14);
xor XOR2 (N29, N26, N11);
and AND3 (N30, N12, N29, N14);
nor NOR2 (N31, N7, N15);
xor XOR2 (N32, N24, N20);
and AND3 (N33, N3, N8, N23);
xor XOR2 (N34, N14, N6);
xor XOR2 (N35, N27, N29);
xor XOR2 (N36, N33, N6);
not NOT1 (N37, N28);
and AND4 (N38, N30, N27, N19, N20);
not NOT1 (N39, N37);
nor NOR2 (N40, N39, N11);
xor XOR2 (N41, N38, N26);
xor XOR2 (N42, N21, N29);
xor XOR2 (N43, N32, N8);
or OR4 (N44, N42, N14, N18, N9);
and AND4 (N45, N2, N18, N39, N40);
not NOT1 (N46, N29);
not NOT1 (N47, N25);
and AND3 (N48, N34, N18, N13);
xor XOR2 (N49, N47, N34);
not NOT1 (N50, N44);
not NOT1 (N51, N45);
nor NOR3 (N52, N43, N15, N5);
or OR2 (N53, N48, N49);
not NOT1 (N54, N50);
nand NAND4 (N55, N1, N19, N14, N13);
nor NOR3 (N56, N55, N54, N1);
and AND3 (N57, N31, N47, N4);
nor NOR2 (N58, N21, N40);
or OR4 (N59, N46, N44, N3, N27);
or OR2 (N60, N35, N11);
buf BUF1 (N61, N52);
nor NOR2 (N62, N61, N30);
and AND4 (N63, N59, N51, N3, N61);
nand NAND3 (N64, N22, N1, N33);
nor NOR2 (N65, N56, N8);
xor XOR2 (N66, N41, N29);
buf BUF1 (N67, N60);
xor XOR2 (N68, N67, N27);
not NOT1 (N69, N64);
buf BUF1 (N70, N53);
and AND3 (N71, N63, N1, N6);
xor XOR2 (N72, N58, N25);
nor NOR4 (N73, N62, N57, N13, N10);
xor XOR2 (N74, N64, N31);
nand NAND2 (N75, N70, N31);
buf BUF1 (N76, N66);
and AND3 (N77, N75, N11, N33);
buf BUF1 (N78, N71);
or OR4 (N79, N68, N41, N54, N78);
or OR2 (N80, N62, N58);
xor XOR2 (N81, N36, N61);
nand NAND4 (N82, N79, N56, N31, N22);
nor NOR3 (N83, N80, N26, N47);
or OR2 (N84, N74, N71);
and AND4 (N85, N72, N73, N77, N48);
not NOT1 (N86, N9);
not NOT1 (N87, N19);
and AND4 (N88, N69, N25, N67, N10);
nor NOR3 (N89, N84, N88, N20);
not NOT1 (N90, N40);
not NOT1 (N91, N83);
or OR3 (N92, N91, N56, N71);
not NOT1 (N93, N81);
and AND4 (N94, N85, N49, N14, N14);
xor XOR2 (N95, N65, N44);
and AND2 (N96, N82, N60);
and AND3 (N97, N86, N80, N94);
nand NAND3 (N98, N46, N2, N46);
xor XOR2 (N99, N97, N90);
buf BUF1 (N100, N51);
or OR4 (N101, N89, N33, N40, N88);
and AND2 (N102, N92, N70);
buf BUF1 (N103, N100);
buf BUF1 (N104, N93);
and AND3 (N105, N103, N80, N71);
not NOT1 (N106, N96);
or OR2 (N107, N95, N7);
nor NOR2 (N108, N101, N66);
not NOT1 (N109, N99);
nor NOR3 (N110, N106, N89, N52);
not NOT1 (N111, N98);
and AND4 (N112, N108, N45, N59, N25);
xor XOR2 (N113, N109, N112);
buf BUF1 (N114, N107);
or OR3 (N115, N93, N5, N26);
not NOT1 (N116, N102);
or OR4 (N117, N110, N73, N48, N52);
nor NOR2 (N118, N116, N38);
buf BUF1 (N119, N105);
or OR2 (N120, N119, N106);
not NOT1 (N121, N111);
not NOT1 (N122, N115);
nand NAND4 (N123, N76, N73, N68, N16);
xor XOR2 (N124, N118, N54);
nand NAND3 (N125, N87, N38, N117);
and AND3 (N126, N104, N58, N38);
nor NOR2 (N127, N126, N89);
or OR3 (N128, N63, N67, N50);
nor NOR2 (N129, N114, N39);
nand NAND3 (N130, N120, N94, N77);
not NOT1 (N131, N122);
or OR2 (N132, N129, N2);
not NOT1 (N133, N130);
and AND4 (N134, N132, N36, N48, N45);
nand NAND2 (N135, N127, N101);
xor XOR2 (N136, N123, N20);
buf BUF1 (N137, N134);
not NOT1 (N138, N131);
nand NAND2 (N139, N138, N110);
buf BUF1 (N140, N121);
nand NAND2 (N141, N136, N102);
and AND3 (N142, N124, N15, N110);
nor NOR4 (N143, N137, N77, N125, N76);
and AND3 (N144, N42, N54, N20);
or OR2 (N145, N141, N10);
not NOT1 (N146, N133);
not NOT1 (N147, N144);
nor NOR4 (N148, N145, N8, N84, N41);
nand NAND2 (N149, N143, N16);
buf BUF1 (N150, N142);
or OR3 (N151, N139, N8, N91);
xor XOR2 (N152, N135, N119);
and AND2 (N153, N149, N46);
nand NAND2 (N154, N146, N47);
nor NOR3 (N155, N150, N20, N18);
or OR4 (N156, N113, N82, N140, N25);
or OR3 (N157, N19, N131, N26);
buf BUF1 (N158, N151);
nor NOR3 (N159, N155, N31, N29);
xor XOR2 (N160, N154, N118);
nand NAND3 (N161, N160, N42, N51);
nor NOR4 (N162, N147, N73, N159, N157);
buf BUF1 (N163, N4);
xor XOR2 (N164, N88, N63);
and AND3 (N165, N163, N135, N70);
not NOT1 (N166, N128);
and AND4 (N167, N161, N1, N9, N103);
and AND4 (N168, N158, N134, N125, N4);
and AND2 (N169, N152, N37);
xor XOR2 (N170, N167, N38);
or OR2 (N171, N156, N56);
nand NAND3 (N172, N165, N156, N111);
xor XOR2 (N173, N169, N113);
or OR4 (N174, N162, N163, N102, N45);
nor NOR4 (N175, N173, N122, N87, N10);
buf BUF1 (N176, N153);
nand NAND4 (N177, N174, N168, N68, N24);
xor XOR2 (N178, N170, N51);
or OR2 (N179, N113, N84);
nand NAND2 (N180, N166, N141);
buf BUF1 (N181, N176);
not NOT1 (N182, N172);
and AND4 (N183, N175, N32, N145, N39);
or OR2 (N184, N178, N87);
nand NAND3 (N185, N182, N150, N134);
and AND3 (N186, N171, N24, N60);
or OR4 (N187, N185, N180, N85, N72);
or OR3 (N188, N136, N52, N42);
or OR3 (N189, N184, N46, N129);
nand NAND4 (N190, N188, N29, N101, N106);
buf BUF1 (N191, N187);
buf BUF1 (N192, N181);
xor XOR2 (N193, N177, N19);
xor XOR2 (N194, N192, N187);
buf BUF1 (N195, N191);
nand NAND4 (N196, N179, N12, N57, N103);
xor XOR2 (N197, N193, N130);
nand NAND2 (N198, N194, N129);
not NOT1 (N199, N148);
buf BUF1 (N200, N190);
not NOT1 (N201, N199);
xor XOR2 (N202, N195, N56);
xor XOR2 (N203, N202, N129);
or OR3 (N204, N198, N114, N7);
not NOT1 (N205, N196);
not NOT1 (N206, N204);
xor XOR2 (N207, N186, N150);
nand NAND2 (N208, N183, N189);
not NOT1 (N209, N61);
and AND2 (N210, N206, N30);
nand NAND2 (N211, N208, N144);
or OR4 (N212, N200, N135, N128, N115);
or OR4 (N213, N201, N203, N162, N95);
nor NOR4 (N214, N44, N2, N59, N75);
and AND4 (N215, N214, N131, N46, N26);
xor XOR2 (N216, N197, N83);
nor NOR2 (N217, N212, N174);
not NOT1 (N218, N205);
nand NAND4 (N219, N217, N119, N21, N199);
or OR4 (N220, N210, N207, N89, N104);
xor XOR2 (N221, N50, N214);
nand NAND3 (N222, N164, N150, N86);
or OR2 (N223, N222, N187);
buf BUF1 (N224, N221);
xor XOR2 (N225, N213, N183);
and AND4 (N226, N224, N25, N111, N5);
buf BUF1 (N227, N226);
or OR3 (N228, N211, N114, N31);
xor XOR2 (N229, N219, N32);
nor NOR4 (N230, N225, N68, N16, N46);
or OR2 (N231, N209, N210);
buf BUF1 (N232, N220);
and AND4 (N233, N231, N74, N215, N55);
xor XOR2 (N234, N144, N13);
or OR3 (N235, N227, N197, N32);
nor NOR2 (N236, N230, N136);
buf BUF1 (N237, N223);
or OR2 (N238, N237, N71);
or OR3 (N239, N218, N36, N30);
or OR2 (N240, N216, N15);
xor XOR2 (N241, N233, N164);
buf BUF1 (N242, N234);
not NOT1 (N243, N236);
xor XOR2 (N244, N243, N53);
not NOT1 (N245, N241);
nand NAND4 (N246, N229, N218, N121, N239);
buf BUF1 (N247, N140);
not NOT1 (N248, N240);
nand NAND3 (N249, N244, N240, N105);
nand NAND4 (N250, N232, N43, N120, N136);
or OR4 (N251, N246, N183, N22, N180);
xor XOR2 (N252, N228, N115);
and AND3 (N253, N242, N178, N104);
buf BUF1 (N254, N249);
or OR2 (N255, N238, N64);
or OR2 (N256, N250, N150);
or OR4 (N257, N248, N82, N69, N234);
xor XOR2 (N258, N247, N81);
nand NAND3 (N259, N254, N117, N86);
and AND4 (N260, N256, N88, N216, N114);
nor NOR2 (N261, N252, N194);
or OR3 (N262, N245, N26, N45);
nand NAND4 (N263, N262, N239, N222, N205);
buf BUF1 (N264, N263);
buf BUF1 (N265, N258);
not NOT1 (N266, N264);
xor XOR2 (N267, N265, N95);
not NOT1 (N268, N259);
or OR2 (N269, N257, N138);
buf BUF1 (N270, N235);
and AND2 (N271, N270, N99);
nand NAND3 (N272, N255, N119, N205);
not NOT1 (N273, N260);
not NOT1 (N274, N272);
xor XOR2 (N275, N261, N139);
nand NAND3 (N276, N271, N48, N215);
or OR3 (N277, N268, N189, N60);
nor NOR2 (N278, N267, N66);
or OR3 (N279, N269, N59, N248);
buf BUF1 (N280, N273);
nand NAND3 (N281, N251, N177, N204);
nor NOR2 (N282, N274, N242);
xor XOR2 (N283, N282, N211);
nand NAND2 (N284, N275, N56);
nand NAND4 (N285, N284, N8, N126, N213);
xor XOR2 (N286, N276, N27);
xor XOR2 (N287, N278, N59);
and AND3 (N288, N283, N204, N21);
and AND4 (N289, N286, N179, N270, N165);
nor NOR4 (N290, N277, N3, N113, N266);
and AND2 (N291, N8, N196);
not NOT1 (N292, N280);
and AND2 (N293, N292, N280);
nor NOR4 (N294, N288, N197, N40, N200);
or OR2 (N295, N253, N131);
or OR4 (N296, N281, N54, N287, N99);
not NOT1 (N297, N239);
buf BUF1 (N298, N285);
buf BUF1 (N299, N296);
nand NAND3 (N300, N295, N16, N150);
and AND4 (N301, N294, N231, N226, N94);
not NOT1 (N302, N293);
not NOT1 (N303, N297);
nor NOR2 (N304, N299, N123);
or OR3 (N305, N303, N234, N84);
not NOT1 (N306, N298);
nand NAND3 (N307, N302, N121, N43);
xor XOR2 (N308, N300, N53);
nor NOR3 (N309, N305, N106, N85);
buf BUF1 (N310, N308);
or OR2 (N311, N309, N99);
nor NOR3 (N312, N311, N209, N131);
nand NAND3 (N313, N312, N66, N176);
not NOT1 (N314, N306);
not NOT1 (N315, N291);
or OR3 (N316, N301, N71, N129);
xor XOR2 (N317, N310, N26);
not NOT1 (N318, N307);
nor NOR4 (N319, N289, N22, N57, N169);
and AND3 (N320, N279, N18, N270);
xor XOR2 (N321, N313, N214);
nand NAND3 (N322, N314, N234, N257);
nand NAND4 (N323, N319, N237, N210, N281);
buf BUF1 (N324, N316);
not NOT1 (N325, N318);
nor NOR2 (N326, N324, N235);
nand NAND4 (N327, N325, N40, N53, N165);
or OR4 (N328, N322, N222, N170, N73);
or OR2 (N329, N326, N311);
xor XOR2 (N330, N290, N77);
xor XOR2 (N331, N323, N205);
or OR2 (N332, N315, N293);
and AND3 (N333, N320, N85, N207);
nand NAND2 (N334, N317, N54);
not NOT1 (N335, N334);
xor XOR2 (N336, N333, N80);
buf BUF1 (N337, N336);
not NOT1 (N338, N332);
buf BUF1 (N339, N328);
xor XOR2 (N340, N337, N316);
nand NAND4 (N341, N340, N294, N210, N206);
buf BUF1 (N342, N327);
nor NOR2 (N343, N341, N169);
nor NOR2 (N344, N343, N274);
nand NAND2 (N345, N321, N190);
and AND3 (N346, N339, N15, N184);
buf BUF1 (N347, N342);
nand NAND2 (N348, N346, N112);
nand NAND2 (N349, N347, N193);
nor NOR3 (N350, N345, N97, N118);
and AND2 (N351, N349, N271);
xor XOR2 (N352, N350, N340);
nand NAND3 (N353, N352, N163, N11);
or OR4 (N354, N344, N110, N125, N198);
not NOT1 (N355, N338);
buf BUF1 (N356, N335);
xor XOR2 (N357, N354, N183);
nand NAND2 (N358, N353, N122);
or OR4 (N359, N357, N355, N81, N213);
buf BUF1 (N360, N11);
nor NOR2 (N361, N329, N343);
and AND2 (N362, N358, N21);
not NOT1 (N363, N351);
nand NAND3 (N364, N360, N270, N185);
or OR2 (N365, N363, N279);
nand NAND2 (N366, N359, N74);
nor NOR4 (N367, N365, N307, N258, N207);
or OR2 (N368, N366, N216);
not NOT1 (N369, N368);
xor XOR2 (N370, N348, N204);
nor NOR4 (N371, N331, N170, N67, N25);
not NOT1 (N372, N304);
buf BUF1 (N373, N330);
xor XOR2 (N374, N364, N223);
nand NAND4 (N375, N374, N322, N337, N40);
nor NOR3 (N376, N372, N237, N65);
buf BUF1 (N377, N370);
xor XOR2 (N378, N356, N338);
nand NAND4 (N379, N378, N163, N243, N308);
or OR4 (N380, N379, N376, N164, N284);
not NOT1 (N381, N347);
nand NAND2 (N382, N367, N47);
nor NOR3 (N383, N375, N176, N36);
and AND3 (N384, N373, N147, N258);
xor XOR2 (N385, N382, N246);
xor XOR2 (N386, N381, N344);
nand NAND4 (N387, N369, N285, N11, N336);
and AND3 (N388, N361, N362, N349);
and AND3 (N389, N382, N305, N293);
and AND4 (N390, N386, N323, N318, N299);
xor XOR2 (N391, N389, N236);
nor NOR3 (N392, N384, N112, N332);
xor XOR2 (N393, N377, N192);
buf BUF1 (N394, N371);
or OR3 (N395, N390, N218, N95);
not NOT1 (N396, N392);
not NOT1 (N397, N387);
nand NAND2 (N398, N397, N19);
xor XOR2 (N399, N396, N354);
nor NOR2 (N400, N388, N165);
nand NAND2 (N401, N400, N370);
nor NOR3 (N402, N380, N35, N105);
and AND4 (N403, N385, N122, N89, N214);
buf BUF1 (N404, N394);
not NOT1 (N405, N398);
not NOT1 (N406, N393);
xor XOR2 (N407, N391, N398);
nand NAND3 (N408, N403, N40, N258);
or OR3 (N409, N402, N376, N271);
or OR2 (N410, N399, N363);
buf BUF1 (N411, N410);
or OR2 (N412, N411, N106);
xor XOR2 (N413, N395, N62);
nor NOR3 (N414, N406, N253, N214);
nor NOR4 (N415, N405, N148, N18, N198);
or OR3 (N416, N404, N125, N153);
or OR3 (N417, N408, N378, N413);
nand NAND3 (N418, N119, N52, N166);
buf BUF1 (N419, N401);
and AND2 (N420, N417, N43);
nand NAND3 (N421, N419, N61, N183);
or OR3 (N422, N420, N83, N384);
buf BUF1 (N423, N383);
or OR4 (N424, N416, N397, N241, N34);
not NOT1 (N425, N424);
buf BUF1 (N426, N422);
buf BUF1 (N427, N412);
not NOT1 (N428, N425);
not NOT1 (N429, N415);
nor NOR3 (N430, N418, N201, N81);
buf BUF1 (N431, N430);
nor NOR4 (N432, N421, N387, N118, N190);
buf BUF1 (N433, N426);
nor NOR2 (N434, N423, N277);
nor NOR4 (N435, N433, N388, N381, N63);
nor NOR2 (N436, N435, N45);
nor NOR4 (N437, N429, N290, N407, N377);
buf BUF1 (N438, N157);
buf BUF1 (N439, N428);
xor XOR2 (N440, N431, N69);
and AND3 (N441, N434, N306, N268);
buf BUF1 (N442, N427);
nand NAND2 (N443, N432, N214);
nand NAND2 (N444, N414, N361);
not NOT1 (N445, N443);
xor XOR2 (N446, N440, N190);
not NOT1 (N447, N409);
xor XOR2 (N448, N436, N357);
xor XOR2 (N449, N448, N389);
or OR3 (N450, N447, N207, N116);
buf BUF1 (N451, N445);
nor NOR3 (N452, N451, N206, N143);
and AND3 (N453, N444, N83, N194);
not NOT1 (N454, N437);
nand NAND3 (N455, N453, N25, N321);
buf BUF1 (N456, N438);
or OR4 (N457, N454, N208, N255, N415);
xor XOR2 (N458, N456, N240);
nor NOR3 (N459, N458, N409, N336);
buf BUF1 (N460, N441);
nand NAND3 (N461, N449, N138, N43);
nor NOR2 (N462, N455, N173);
or OR2 (N463, N450, N25);
buf BUF1 (N464, N442);
xor XOR2 (N465, N457, N456);
not NOT1 (N466, N462);
not NOT1 (N467, N465);
nor NOR4 (N468, N459, N134, N377, N114);
or OR3 (N469, N452, N317, N205);
buf BUF1 (N470, N468);
nor NOR2 (N471, N461, N240);
and AND3 (N472, N469, N342, N49);
buf BUF1 (N473, N466);
nor NOR4 (N474, N463, N115, N391, N10);
nand NAND3 (N475, N473, N131, N146);
buf BUF1 (N476, N470);
not NOT1 (N477, N464);
not NOT1 (N478, N439);
and AND4 (N479, N472, N318, N393, N184);
nor NOR3 (N480, N475, N2, N142);
xor XOR2 (N481, N477, N239);
or OR4 (N482, N481, N416, N427, N74);
xor XOR2 (N483, N467, N3);
not NOT1 (N484, N482);
or OR4 (N485, N480, N325, N141, N153);
nand NAND4 (N486, N484, N377, N241, N141);
nor NOR2 (N487, N485, N300);
nand NAND4 (N488, N471, N75, N75, N144);
nand NAND2 (N489, N476, N262);
nand NAND2 (N490, N489, N371);
not NOT1 (N491, N460);
or OR4 (N492, N487, N313, N116, N163);
and AND3 (N493, N446, N130, N19);
and AND2 (N494, N474, N132);
nor NOR2 (N495, N478, N481);
xor XOR2 (N496, N479, N1);
and AND3 (N497, N495, N426, N436);
or OR3 (N498, N486, N44, N137);
and AND2 (N499, N491, N35);
xor XOR2 (N500, N488, N88);
and AND4 (N501, N498, N159, N161, N118);
nor NOR2 (N502, N494, N408);
and AND3 (N503, N492, N235, N381);
not NOT1 (N504, N501);
not NOT1 (N505, N504);
and AND4 (N506, N497, N277, N133, N45);
xor XOR2 (N507, N506, N232);
or OR4 (N508, N500, N250, N498, N396);
nor NOR3 (N509, N502, N123, N235);
xor XOR2 (N510, N507, N162);
nor NOR3 (N511, N510, N173, N123);
and AND2 (N512, N511, N415);
xor XOR2 (N513, N483, N127);
xor XOR2 (N514, N496, N164);
or OR4 (N515, N512, N393, N309, N405);
and AND2 (N516, N503, N84);
buf BUF1 (N517, N499);
not NOT1 (N518, N517);
and AND4 (N519, N515, N79, N300, N151);
buf BUF1 (N520, N514);
or OR3 (N521, N490, N466, N414);
or OR4 (N522, N513, N458, N230, N184);
xor XOR2 (N523, N516, N482);
nand NAND4 (N524, N519, N289, N164, N444);
buf BUF1 (N525, N522);
buf BUF1 (N526, N524);
or OR4 (N527, N525, N29, N133, N77);
not NOT1 (N528, N523);
not NOT1 (N529, N518);
or OR3 (N530, N526, N171, N191);
and AND2 (N531, N493, N206);
xor XOR2 (N532, N521, N513);
not NOT1 (N533, N508);
and AND2 (N534, N530, N91);
buf BUF1 (N535, N531);
and AND3 (N536, N533, N237, N218);
nand NAND3 (N537, N505, N480, N492);
and AND3 (N538, N536, N101, N222);
or OR3 (N539, N534, N513, N1);
nor NOR4 (N540, N539, N330, N10, N203);
and AND2 (N541, N520, N158);
and AND2 (N542, N529, N175);
nor NOR3 (N543, N537, N65, N532);
not NOT1 (N544, N493);
nor NOR3 (N545, N528, N406, N370);
nand NAND2 (N546, N527, N243);
xor XOR2 (N547, N544, N504);
nor NOR4 (N548, N540, N76, N481, N98);
nand NAND3 (N549, N546, N92, N171);
nor NOR3 (N550, N535, N391, N48);
and AND2 (N551, N543, N515);
nor NOR2 (N552, N542, N419);
nor NOR2 (N553, N545, N51);
not NOT1 (N554, N509);
or OR2 (N555, N554, N429);
buf BUF1 (N556, N538);
xor XOR2 (N557, N552, N409);
nand NAND4 (N558, N549, N352, N298, N340);
nand NAND2 (N559, N551, N361);
buf BUF1 (N560, N555);
not NOT1 (N561, N558);
nand NAND3 (N562, N557, N131, N369);
nand NAND4 (N563, N550, N127, N102, N144);
buf BUF1 (N564, N559);
nand NAND3 (N565, N553, N438, N148);
xor XOR2 (N566, N548, N509);
and AND4 (N567, N566, N270, N461, N312);
nor NOR4 (N568, N547, N234, N416, N546);
not NOT1 (N569, N560);
nor NOR2 (N570, N568, N163);
nand NAND2 (N571, N563, N139);
nand NAND2 (N572, N569, N458);
nor NOR4 (N573, N571, N546, N328, N141);
xor XOR2 (N574, N572, N151);
nor NOR2 (N575, N573, N526);
nor NOR3 (N576, N574, N483, N436);
and AND3 (N577, N561, N347, N157);
buf BUF1 (N578, N541);
nand NAND2 (N579, N578, N519);
nand NAND2 (N580, N576, N140);
not NOT1 (N581, N579);
or OR4 (N582, N577, N78, N514, N94);
and AND2 (N583, N581, N156);
buf BUF1 (N584, N562);
not NOT1 (N585, N575);
nor NOR4 (N586, N583, N522, N411, N79);
nor NOR4 (N587, N564, N154, N109, N94);
or OR4 (N588, N586, N102, N481, N533);
xor XOR2 (N589, N588, N375);
nand NAND2 (N590, N570, N553);
or OR2 (N591, N587, N284);
or OR2 (N592, N580, N458);
buf BUF1 (N593, N567);
or OR3 (N594, N590, N61, N308);
and AND3 (N595, N592, N395, N544);
not NOT1 (N596, N582);
buf BUF1 (N597, N591);
and AND2 (N598, N595, N310);
xor XOR2 (N599, N589, N225);
and AND4 (N600, N599, N379, N342, N120);
xor XOR2 (N601, N596, N309);
xor XOR2 (N602, N584, N594);
nor NOR3 (N603, N265, N562, N203);
nand NAND2 (N604, N600, N448);
xor XOR2 (N605, N556, N258);
not NOT1 (N606, N598);
nor NOR2 (N607, N606, N86);
nor NOR4 (N608, N597, N492, N596, N116);
not NOT1 (N609, N603);
nand NAND2 (N610, N593, N402);
or OR2 (N611, N585, N98);
buf BUF1 (N612, N611);
or OR2 (N613, N612, N158);
or OR4 (N614, N607, N125, N39, N86);
or OR4 (N615, N610, N231, N113, N202);
nand NAND4 (N616, N601, N468, N538, N378);
and AND3 (N617, N608, N614, N599);
and AND3 (N618, N118, N522, N509);
not NOT1 (N619, N616);
xor XOR2 (N620, N604, N152);
nor NOR3 (N621, N609, N64, N471);
and AND2 (N622, N617, N527);
buf BUF1 (N623, N565);
nand NAND4 (N624, N621, N219, N79, N202);
xor XOR2 (N625, N605, N552);
not NOT1 (N626, N622);
xor XOR2 (N627, N619, N264);
nand NAND2 (N628, N625, N613);
xor XOR2 (N629, N325, N187);
and AND4 (N630, N628, N627, N438, N550);
xor XOR2 (N631, N268, N555);
nor NOR4 (N632, N629, N363, N276, N112);
xor XOR2 (N633, N602, N468);
xor XOR2 (N634, N631, N610);
nor NOR3 (N635, N623, N228, N294);
nor NOR3 (N636, N634, N311, N165);
xor XOR2 (N637, N635, N626);
or OR4 (N638, N251, N278, N318, N100);
buf BUF1 (N639, N620);
nor NOR3 (N640, N637, N47, N137);
buf BUF1 (N641, N633);
not NOT1 (N642, N638);
buf BUF1 (N643, N624);
xor XOR2 (N644, N615, N512);
nand NAND2 (N645, N632, N326);
buf BUF1 (N646, N640);
nand NAND4 (N647, N639, N282, N94, N446);
nand NAND3 (N648, N618, N210, N24);
and AND3 (N649, N648, N423, N53);
not NOT1 (N650, N649);
xor XOR2 (N651, N641, N264);
xor XOR2 (N652, N645, N29);
nand NAND2 (N653, N651, N383);
xor XOR2 (N654, N647, N581);
buf BUF1 (N655, N646);
nor NOR2 (N656, N644, N313);
nand NAND2 (N657, N630, N487);
buf BUF1 (N658, N652);
or OR3 (N659, N643, N388, N405);
nor NOR4 (N660, N657, N461, N344, N614);
or OR2 (N661, N642, N340);
and AND3 (N662, N654, N326, N22);
nand NAND4 (N663, N661, N377, N436, N60);
buf BUF1 (N664, N659);
buf BUF1 (N665, N662);
nor NOR3 (N666, N665, N188, N123);
nor NOR2 (N667, N664, N414);
nand NAND4 (N668, N660, N92, N574, N148);
xor XOR2 (N669, N663, N317);
xor XOR2 (N670, N668, N11);
buf BUF1 (N671, N636);
and AND3 (N672, N666, N208, N364);
or OR4 (N673, N670, N391, N456, N517);
not NOT1 (N674, N653);
not NOT1 (N675, N669);
nand NAND4 (N676, N667, N69, N312, N339);
and AND3 (N677, N676, N28, N154);
not NOT1 (N678, N650);
xor XOR2 (N679, N677, N91);
and AND4 (N680, N658, N302, N176, N112);
buf BUF1 (N681, N680);
or OR3 (N682, N671, N476, N129);
and AND2 (N683, N675, N551);
buf BUF1 (N684, N655);
buf BUF1 (N685, N682);
not NOT1 (N686, N673);
xor XOR2 (N687, N656, N231);
buf BUF1 (N688, N679);
not NOT1 (N689, N686);
or OR2 (N690, N685, N553);
not NOT1 (N691, N683);
xor XOR2 (N692, N690, N183);
nor NOR4 (N693, N689, N312, N25, N266);
nor NOR3 (N694, N688, N421, N202);
buf BUF1 (N695, N687);
and AND2 (N696, N674, N86);
buf BUF1 (N697, N691);
nand NAND4 (N698, N694, N568, N531, N576);
xor XOR2 (N699, N696, N13);
buf BUF1 (N700, N699);
nand NAND4 (N701, N693, N185, N670, N687);
not NOT1 (N702, N672);
and AND4 (N703, N697, N235, N7, N11);
xor XOR2 (N704, N692, N466);
and AND4 (N705, N684, N481, N481, N28);
buf BUF1 (N706, N700);
and AND4 (N707, N706, N33, N55, N317);
or OR2 (N708, N701, N80);
nand NAND3 (N709, N708, N242, N665);
and AND3 (N710, N705, N485, N666);
buf BUF1 (N711, N710);
buf BUF1 (N712, N681);
not NOT1 (N713, N695);
nand NAND3 (N714, N702, N230, N553);
nor NOR3 (N715, N711, N342, N474);
xor XOR2 (N716, N698, N433);
or OR3 (N717, N703, N17, N22);
nand NAND2 (N718, N678, N345);
nor NOR4 (N719, N713, N47, N302, N556);
or OR4 (N720, N707, N251, N100, N477);
nand NAND2 (N721, N719, N628);
nor NOR4 (N722, N704, N714, N125, N504);
nand NAND4 (N723, N239, N324, N540, N401);
nand NAND4 (N724, N716, N488, N715, N400);
and AND4 (N725, N373, N388, N459, N558);
not NOT1 (N726, N721);
not NOT1 (N727, N725);
nand NAND2 (N728, N712, N154);
nand NAND4 (N729, N726, N693, N439, N554);
or OR3 (N730, N728, N497, N413);
or OR2 (N731, N723, N281);
nand NAND4 (N732, N718, N315, N332, N93);
xor XOR2 (N733, N722, N37);
buf BUF1 (N734, N730);
not NOT1 (N735, N732);
xor XOR2 (N736, N717, N314);
xor XOR2 (N737, N720, N420);
not NOT1 (N738, N731);
not NOT1 (N739, N733);
nand NAND3 (N740, N734, N636, N466);
buf BUF1 (N741, N740);
and AND2 (N742, N727, N639);
xor XOR2 (N743, N735, N272);
nor NOR2 (N744, N738, N141);
and AND3 (N745, N744, N287, N509);
or OR3 (N746, N724, N330, N495);
and AND4 (N747, N742, N733, N367, N272);
xor XOR2 (N748, N729, N111);
nand NAND4 (N749, N748, N650, N721, N440);
xor XOR2 (N750, N743, N671);
and AND2 (N751, N739, N505);
nor NOR3 (N752, N746, N116, N177);
and AND4 (N753, N741, N10, N427, N248);
xor XOR2 (N754, N737, N436);
xor XOR2 (N755, N754, N366);
xor XOR2 (N756, N755, N291);
not NOT1 (N757, N751);
xor XOR2 (N758, N709, N58);
nand NAND2 (N759, N758, N456);
not NOT1 (N760, N757);
nand NAND2 (N761, N759, N6);
nor NOR4 (N762, N760, N330, N298, N241);
nand NAND4 (N763, N762, N544, N100, N10);
not NOT1 (N764, N747);
not NOT1 (N765, N761);
buf BUF1 (N766, N752);
not NOT1 (N767, N753);
not NOT1 (N768, N767);
or OR2 (N769, N765, N645);
not NOT1 (N770, N764);
buf BUF1 (N771, N768);
xor XOR2 (N772, N736, N700);
or OR2 (N773, N771, N693);
buf BUF1 (N774, N763);
nor NOR2 (N775, N774, N595);
and AND4 (N776, N775, N121, N682, N151);
buf BUF1 (N777, N756);
nor NOR4 (N778, N773, N294, N677, N566);
not NOT1 (N779, N778);
not NOT1 (N780, N777);
xor XOR2 (N781, N779, N237);
buf BUF1 (N782, N766);
or OR3 (N783, N776, N488, N753);
and AND3 (N784, N781, N689, N386);
buf BUF1 (N785, N783);
and AND2 (N786, N784, N620);
not NOT1 (N787, N770);
nor NOR4 (N788, N786, N605, N230, N291);
nor NOR3 (N789, N785, N584, N775);
nor NOR2 (N790, N788, N218);
not NOT1 (N791, N789);
not NOT1 (N792, N749);
nand NAND4 (N793, N772, N526, N231, N497);
or OR4 (N794, N791, N33, N695, N544);
and AND4 (N795, N745, N82, N204, N336);
nor NOR4 (N796, N750, N216, N113, N713);
not NOT1 (N797, N796);
or OR4 (N798, N790, N566, N562, N372);
and AND4 (N799, N787, N166, N446, N498);
or OR3 (N800, N797, N414, N671);
or OR4 (N801, N780, N669, N14, N564);
nor NOR3 (N802, N799, N552, N665);
xor XOR2 (N803, N798, N722);
buf BUF1 (N804, N803);
nor NOR4 (N805, N801, N797, N506, N165);
not NOT1 (N806, N805);
nand NAND4 (N807, N793, N140, N7, N751);
not NOT1 (N808, N794);
buf BUF1 (N809, N804);
buf BUF1 (N810, N792);
nor NOR3 (N811, N810, N183, N194);
or OR3 (N812, N802, N301, N577);
and AND2 (N813, N811, N454);
not NOT1 (N814, N769);
buf BUF1 (N815, N806);
buf BUF1 (N816, N782);
or OR2 (N817, N813, N217);
nor NOR3 (N818, N809, N283, N764);
nor NOR3 (N819, N817, N401, N326);
buf BUF1 (N820, N812);
nand NAND3 (N821, N808, N251, N271);
nor NOR3 (N822, N821, N593, N631);
xor XOR2 (N823, N816, N729);
buf BUF1 (N824, N800);
nor NOR2 (N825, N824, N492);
xor XOR2 (N826, N814, N55);
nor NOR3 (N827, N818, N463, N110);
or OR2 (N828, N822, N317);
xor XOR2 (N829, N827, N477);
nand NAND3 (N830, N829, N787, N629);
not NOT1 (N831, N807);
not NOT1 (N832, N823);
or OR2 (N833, N826, N712);
buf BUF1 (N834, N833);
or OR2 (N835, N815, N443);
xor XOR2 (N836, N835, N58);
not NOT1 (N837, N828);
nor NOR4 (N838, N831, N551, N93, N797);
not NOT1 (N839, N820);
not NOT1 (N840, N832);
and AND3 (N841, N795, N212, N430);
and AND4 (N842, N834, N100, N481, N590);
xor XOR2 (N843, N839, N746);
and AND3 (N844, N840, N75, N482);
not NOT1 (N845, N841);
xor XOR2 (N846, N838, N91);
nor NOR4 (N847, N836, N204, N31, N597);
buf BUF1 (N848, N837);
not NOT1 (N849, N830);
xor XOR2 (N850, N825, N838);
nand NAND3 (N851, N849, N760, N87);
not NOT1 (N852, N845);
or OR3 (N853, N842, N726, N30);
or OR4 (N854, N843, N243, N347, N400);
buf BUF1 (N855, N819);
nor NOR3 (N856, N847, N98, N330);
buf BUF1 (N857, N851);
not NOT1 (N858, N848);
nand NAND4 (N859, N858, N77, N444, N484);
xor XOR2 (N860, N844, N199);
not NOT1 (N861, N850);
nand NAND4 (N862, N855, N187, N486, N161);
not NOT1 (N863, N846);
nor NOR3 (N864, N856, N758, N659);
nor NOR3 (N865, N852, N270, N46);
and AND4 (N866, N859, N426, N740, N659);
not NOT1 (N867, N864);
nor NOR3 (N868, N853, N216, N726);
and AND3 (N869, N868, N855, N431);
or OR2 (N870, N863, N28);
nand NAND4 (N871, N857, N724, N585, N646);
or OR2 (N872, N870, N622);
nor NOR4 (N873, N869, N726, N871, N692);
or OR4 (N874, N584, N659, N193, N581);
or OR2 (N875, N867, N223);
not NOT1 (N876, N865);
buf BUF1 (N877, N875);
or OR2 (N878, N862, N428);
xor XOR2 (N879, N877, N778);
not NOT1 (N880, N879);
and AND4 (N881, N860, N145, N123, N669);
and AND4 (N882, N866, N856, N678, N114);
and AND4 (N883, N872, N607, N192, N543);
not NOT1 (N884, N861);
not NOT1 (N885, N876);
nand NAND3 (N886, N880, N800, N144);
and AND4 (N887, N881, N687, N648, N220);
not NOT1 (N888, N882);
xor XOR2 (N889, N886, N244);
nor NOR4 (N890, N878, N470, N255, N278);
nand NAND3 (N891, N884, N354, N549);
or OR3 (N892, N890, N708, N6);
xor XOR2 (N893, N888, N298);
nand NAND4 (N894, N892, N262, N65, N395);
and AND2 (N895, N894, N502);
or OR4 (N896, N885, N567, N132, N205);
not NOT1 (N897, N873);
xor XOR2 (N898, N896, N439);
not NOT1 (N899, N898);
nand NAND4 (N900, N897, N181, N214, N375);
nor NOR3 (N901, N893, N615, N190);
or OR2 (N902, N889, N888);
or OR4 (N903, N891, N192, N302, N392);
and AND2 (N904, N902, N299);
buf BUF1 (N905, N854);
buf BUF1 (N906, N874);
buf BUF1 (N907, N883);
buf BUF1 (N908, N907);
or OR3 (N909, N899, N562, N642);
nor NOR4 (N910, N903, N685, N510, N637);
buf BUF1 (N911, N908);
nand NAND2 (N912, N904, N585);
xor XOR2 (N913, N911, N322);
and AND3 (N914, N901, N626, N344);
and AND2 (N915, N912, N11);
nand NAND3 (N916, N900, N623, N733);
xor XOR2 (N917, N914, N566);
not NOT1 (N918, N895);
or OR2 (N919, N913, N209);
nor NOR4 (N920, N915, N205, N131, N100);
not NOT1 (N921, N917);
buf BUF1 (N922, N918);
nor NOR3 (N923, N909, N655, N65);
xor XOR2 (N924, N922, N819);
not NOT1 (N925, N916);
xor XOR2 (N926, N905, N313);
not NOT1 (N927, N887);
not NOT1 (N928, N927);
not NOT1 (N929, N925);
buf BUF1 (N930, N910);
or OR2 (N931, N921, N337);
xor XOR2 (N932, N919, N128);
xor XOR2 (N933, N923, N839);
nor NOR3 (N934, N931, N856, N597);
nor NOR4 (N935, N926, N96, N118, N481);
buf BUF1 (N936, N930);
nand NAND4 (N937, N933, N876, N539, N870);
not NOT1 (N938, N932);
and AND3 (N939, N935, N324, N432);
not NOT1 (N940, N928);
not NOT1 (N941, N937);
xor XOR2 (N942, N940, N294);
nor NOR4 (N943, N906, N636, N222, N257);
nand NAND4 (N944, N924, N674, N622, N89);
not NOT1 (N945, N943);
or OR4 (N946, N939, N608, N160, N771);
xor XOR2 (N947, N920, N85);
buf BUF1 (N948, N946);
nor NOR2 (N949, N936, N915);
buf BUF1 (N950, N942);
nor NOR4 (N951, N934, N194, N69, N131);
nor NOR4 (N952, N938, N627, N837, N721);
or OR3 (N953, N941, N809, N30);
not NOT1 (N954, N949);
nand NAND3 (N955, N948, N235, N691);
or OR4 (N956, N951, N551, N949, N198);
nand NAND2 (N957, N929, N677);
and AND4 (N958, N953, N833, N621, N706);
or OR2 (N959, N952, N125);
not NOT1 (N960, N956);
nor NOR4 (N961, N945, N433, N420, N19);
not NOT1 (N962, N960);
nand NAND4 (N963, N944, N245, N276, N589);
buf BUF1 (N964, N957);
nand NAND2 (N965, N959, N266);
nand NAND2 (N966, N954, N602);
nor NOR2 (N967, N966, N665);
not NOT1 (N968, N958);
not NOT1 (N969, N965);
nor NOR4 (N970, N963, N253, N164, N451);
nor NOR3 (N971, N962, N442, N772);
nor NOR2 (N972, N969, N684);
nand NAND2 (N973, N967, N555);
nor NOR3 (N974, N968, N412, N649);
nor NOR2 (N975, N947, N329);
buf BUF1 (N976, N955);
xor XOR2 (N977, N964, N371);
or OR2 (N978, N971, N53);
or OR2 (N979, N976, N135);
not NOT1 (N980, N961);
not NOT1 (N981, N978);
not NOT1 (N982, N979);
not NOT1 (N983, N980);
and AND2 (N984, N950, N178);
nor NOR3 (N985, N973, N589, N980);
or OR2 (N986, N974, N424);
nand NAND4 (N987, N982, N807, N617, N846);
buf BUF1 (N988, N987);
or OR2 (N989, N981, N902);
nand NAND2 (N990, N983, N366);
and AND4 (N991, N975, N598, N118, N322);
xor XOR2 (N992, N972, N626);
or OR4 (N993, N989, N698, N141, N670);
nand NAND4 (N994, N970, N415, N143, N294);
xor XOR2 (N995, N992, N216);
xor XOR2 (N996, N984, N850);
nand NAND4 (N997, N988, N464, N91, N605);
nand NAND4 (N998, N996, N710, N283, N142);
nand NAND4 (N999, N997, N25, N65, N449);
not NOT1 (N1000, N990);
nor NOR4 (N1001, N1000, N908, N566, N797);
nor NOR3 (N1002, N999, N2, N290);
and AND3 (N1003, N993, N354, N770);
nor NOR4 (N1004, N1003, N155, N953, N922);
nor NOR3 (N1005, N1002, N795, N443);
or OR2 (N1006, N991, N752);
xor XOR2 (N1007, N998, N737);
or OR3 (N1008, N994, N940, N411);
or OR3 (N1009, N977, N229, N402);
and AND4 (N1010, N1006, N777, N108, N381);
or OR4 (N1011, N1008, N992, N912, N312);
nor NOR3 (N1012, N985, N309, N96);
and AND2 (N1013, N1007, N799);
xor XOR2 (N1014, N1012, N470);
and AND2 (N1015, N1005, N554);
and AND2 (N1016, N1009, N293);
or OR4 (N1017, N1016, N624, N824, N504);
xor XOR2 (N1018, N1015, N538);
nand NAND3 (N1019, N1013, N998, N403);
and AND4 (N1020, N1018, N349, N18, N263);
or OR3 (N1021, N995, N646, N378);
nor NOR3 (N1022, N1019, N792, N626);
and AND3 (N1023, N1014, N575, N883);
and AND4 (N1024, N1020, N794, N865, N543);
nor NOR2 (N1025, N1011, N320);
not NOT1 (N1026, N1023);
nor NOR4 (N1027, N1026, N915, N671, N290);
nor NOR4 (N1028, N1024, N109, N43, N467);
nand NAND3 (N1029, N1025, N1016, N825);
buf BUF1 (N1030, N1017);
nor NOR2 (N1031, N1021, N751);
nor NOR2 (N1032, N1029, N288);
and AND3 (N1033, N1030, N20, N177);
or OR4 (N1034, N1027, N466, N589, N688);
buf BUF1 (N1035, N1001);
nor NOR4 (N1036, N1034, N314, N596, N747);
nor NOR3 (N1037, N1031, N281, N289);
not NOT1 (N1038, N1037);
and AND2 (N1039, N1004, N782);
nor NOR2 (N1040, N1032, N582);
and AND4 (N1041, N1033, N186, N505, N865);
nor NOR4 (N1042, N986, N372, N65, N221);
buf BUF1 (N1043, N1040);
nor NOR3 (N1044, N1041, N676, N369);
nor NOR4 (N1045, N1035, N685, N276, N276);
buf BUF1 (N1046, N1028);
not NOT1 (N1047, N1042);
or OR3 (N1048, N1038, N455, N353);
and AND4 (N1049, N1036, N508, N308, N149);
nand NAND2 (N1050, N1022, N290);
and AND3 (N1051, N1045, N301, N109);
and AND4 (N1052, N1051, N224, N642, N687);
nor NOR3 (N1053, N1044, N807, N147);
nor NOR2 (N1054, N1052, N468);
and AND4 (N1055, N1048, N714, N342, N543);
nand NAND4 (N1056, N1055, N705, N1038, N169);
nor NOR4 (N1057, N1039, N749, N736, N443);
buf BUF1 (N1058, N1057);
not NOT1 (N1059, N1058);
and AND4 (N1060, N1010, N553, N348, N405);
nor NOR3 (N1061, N1047, N799, N714);
not NOT1 (N1062, N1061);
xor XOR2 (N1063, N1059, N132);
not NOT1 (N1064, N1043);
and AND2 (N1065, N1060, N474);
xor XOR2 (N1066, N1065, N576);
xor XOR2 (N1067, N1050, N85);
not NOT1 (N1068, N1056);
nor NOR4 (N1069, N1068, N773, N10, N18);
nor NOR4 (N1070, N1054, N134, N407, N746);
nor NOR3 (N1071, N1046, N806, N895);
not NOT1 (N1072, N1053);
nor NOR2 (N1073, N1063, N46);
and AND3 (N1074, N1064, N407, N62);
or OR2 (N1075, N1070, N708);
and AND3 (N1076, N1074, N281, N427);
and AND4 (N1077, N1069, N658, N661, N648);
xor XOR2 (N1078, N1062, N548);
or OR3 (N1079, N1049, N765, N155);
not NOT1 (N1080, N1073);
and AND3 (N1081, N1076, N43, N370);
buf BUF1 (N1082, N1072);
buf BUF1 (N1083, N1080);
buf BUF1 (N1084, N1077);
and AND2 (N1085, N1082, N480);
and AND3 (N1086, N1084, N841, N911);
or OR2 (N1087, N1075, N657);
nor NOR2 (N1088, N1071, N1013);
nand NAND3 (N1089, N1087, N887, N736);
not NOT1 (N1090, N1089);
and AND4 (N1091, N1079, N714, N92, N106);
nand NAND4 (N1092, N1086, N187, N944, N761);
xor XOR2 (N1093, N1078, N369);
or OR4 (N1094, N1081, N912, N590, N630);
or OR3 (N1095, N1091, N556, N1016);
buf BUF1 (N1096, N1094);
and AND3 (N1097, N1085, N853, N593);
buf BUF1 (N1098, N1097);
nor NOR4 (N1099, N1067, N797, N582, N260);
xor XOR2 (N1100, N1099, N451);
buf BUF1 (N1101, N1095);
nand NAND3 (N1102, N1083, N40, N945);
and AND4 (N1103, N1096, N770, N510, N952);
not NOT1 (N1104, N1101);
xor XOR2 (N1105, N1104, N741);
nand NAND3 (N1106, N1092, N594, N389);
not NOT1 (N1107, N1093);
xor XOR2 (N1108, N1107, N140);
xor XOR2 (N1109, N1098, N891);
buf BUF1 (N1110, N1100);
xor XOR2 (N1111, N1103, N529);
buf BUF1 (N1112, N1111);
or OR2 (N1113, N1090, N733);
or OR4 (N1114, N1105, N723, N836, N739);
and AND3 (N1115, N1102, N251, N362);
nand NAND3 (N1116, N1112, N362, N207);
xor XOR2 (N1117, N1109, N489);
xor XOR2 (N1118, N1117, N500);
buf BUF1 (N1119, N1118);
nand NAND2 (N1120, N1114, N722);
buf BUF1 (N1121, N1088);
not NOT1 (N1122, N1121);
not NOT1 (N1123, N1066);
nand NAND4 (N1124, N1122, N1113, N192, N619);
buf BUF1 (N1125, N796);
not NOT1 (N1126, N1119);
buf BUF1 (N1127, N1106);
or OR3 (N1128, N1127, N454, N323);
nand NAND3 (N1129, N1123, N587, N102);
xor XOR2 (N1130, N1128, N735);
or OR2 (N1131, N1115, N903);
buf BUF1 (N1132, N1116);
not NOT1 (N1133, N1124);
and AND3 (N1134, N1108, N597, N945);
not NOT1 (N1135, N1110);
xor XOR2 (N1136, N1133, N129);
xor XOR2 (N1137, N1129, N915);
and AND2 (N1138, N1131, N200);
buf BUF1 (N1139, N1134);
or OR2 (N1140, N1136, N37);
buf BUF1 (N1141, N1137);
nor NOR4 (N1142, N1140, N444, N498, N418);
xor XOR2 (N1143, N1142, N649);
not NOT1 (N1144, N1120);
nor NOR2 (N1145, N1130, N717);
nand NAND2 (N1146, N1135, N196);
nor NOR2 (N1147, N1138, N154);
not NOT1 (N1148, N1143);
nor NOR4 (N1149, N1145, N401, N308, N116);
and AND3 (N1150, N1141, N112, N300);
xor XOR2 (N1151, N1150, N149);
and AND4 (N1152, N1125, N911, N395, N364);
nor NOR2 (N1153, N1149, N417);
and AND2 (N1154, N1126, N66);
or OR3 (N1155, N1132, N960, N38);
xor XOR2 (N1156, N1154, N332);
nand NAND2 (N1157, N1155, N121);
buf BUF1 (N1158, N1148);
or OR2 (N1159, N1146, N74);
not NOT1 (N1160, N1139);
nand NAND3 (N1161, N1159, N1089, N519);
xor XOR2 (N1162, N1158, N73);
xor XOR2 (N1163, N1160, N942);
nor NOR2 (N1164, N1147, N452);
and AND2 (N1165, N1163, N476);
or OR2 (N1166, N1151, N675);
or OR3 (N1167, N1164, N310, N543);
and AND3 (N1168, N1161, N756, N189);
or OR2 (N1169, N1166, N580);
not NOT1 (N1170, N1168);
nand NAND4 (N1171, N1156, N1106, N462, N635);
xor XOR2 (N1172, N1152, N852);
buf BUF1 (N1173, N1153);
and AND2 (N1174, N1162, N224);
and AND3 (N1175, N1167, N1126, N493);
nand NAND2 (N1176, N1170, N743);
and AND2 (N1177, N1173, N74);
not NOT1 (N1178, N1172);
buf BUF1 (N1179, N1169);
not NOT1 (N1180, N1177);
buf BUF1 (N1181, N1180);
xor XOR2 (N1182, N1144, N801);
or OR4 (N1183, N1174, N94, N196, N201);
not NOT1 (N1184, N1165);
not NOT1 (N1185, N1182);
not NOT1 (N1186, N1184);
or OR3 (N1187, N1183, N700, N265);
nand NAND2 (N1188, N1186, N435);
buf BUF1 (N1189, N1181);
nor NOR3 (N1190, N1178, N529, N272);
or OR2 (N1191, N1175, N15);
nand NAND4 (N1192, N1179, N193, N856, N862);
buf BUF1 (N1193, N1192);
xor XOR2 (N1194, N1187, N920);
nand NAND3 (N1195, N1188, N793, N567);
and AND2 (N1196, N1185, N861);
nor NOR3 (N1197, N1194, N401, N540);
nand NAND3 (N1198, N1190, N351, N1028);
not NOT1 (N1199, N1171);
xor XOR2 (N1200, N1157, N5);
nor NOR3 (N1201, N1197, N247, N47);
or OR4 (N1202, N1201, N214, N1201, N226);
and AND3 (N1203, N1199, N874, N52);
nand NAND2 (N1204, N1191, N1160);
nor NOR2 (N1205, N1196, N109);
nor NOR3 (N1206, N1205, N255, N745);
xor XOR2 (N1207, N1200, N508);
nor NOR2 (N1208, N1193, N657);
not NOT1 (N1209, N1202);
buf BUF1 (N1210, N1203);
nor NOR2 (N1211, N1176, N1063);
and AND4 (N1212, N1195, N24, N612, N1164);
nor NOR2 (N1213, N1207, N667);
and AND4 (N1214, N1206, N392, N347, N916);
not NOT1 (N1215, N1212);
buf BUF1 (N1216, N1213);
nand NAND3 (N1217, N1211, N138, N843);
buf BUF1 (N1218, N1204);
xor XOR2 (N1219, N1189, N1064);
nand NAND2 (N1220, N1214, N889);
nor NOR2 (N1221, N1215, N432);
or OR3 (N1222, N1209, N803, N1043);
not NOT1 (N1223, N1216);
buf BUF1 (N1224, N1218);
xor XOR2 (N1225, N1222, N187);
or OR4 (N1226, N1224, N74, N459, N751);
or OR2 (N1227, N1208, N703);
xor XOR2 (N1228, N1225, N242);
not NOT1 (N1229, N1220);
or OR4 (N1230, N1219, N210, N308, N540);
xor XOR2 (N1231, N1223, N866);
not NOT1 (N1232, N1226);
nor NOR4 (N1233, N1227, N394, N536, N738);
and AND2 (N1234, N1221, N1186);
nand NAND3 (N1235, N1210, N945, N116);
and AND3 (N1236, N1230, N1005, N789);
xor XOR2 (N1237, N1233, N780);
xor XOR2 (N1238, N1236, N650);
or OR4 (N1239, N1235, N234, N1031, N1040);
nand NAND2 (N1240, N1232, N1020);
or OR2 (N1241, N1238, N234);
and AND3 (N1242, N1231, N392, N1088);
nor NOR3 (N1243, N1242, N242, N407);
nor NOR3 (N1244, N1198, N71, N835);
and AND4 (N1245, N1229, N304, N1107, N614);
or OR3 (N1246, N1217, N233, N44);
and AND2 (N1247, N1228, N496);
not NOT1 (N1248, N1244);
not NOT1 (N1249, N1248);
buf BUF1 (N1250, N1243);
buf BUF1 (N1251, N1246);
and AND2 (N1252, N1234, N339);
nand NAND4 (N1253, N1245, N420, N653, N725);
and AND2 (N1254, N1250, N347);
nand NAND2 (N1255, N1252, N818);
nor NOR4 (N1256, N1249, N1045, N293, N199);
nor NOR2 (N1257, N1254, N599);
xor XOR2 (N1258, N1247, N454);
or OR4 (N1259, N1257, N758, N172, N163);
or OR4 (N1260, N1255, N206, N434, N1117);
nand NAND3 (N1261, N1240, N1140, N1088);
and AND3 (N1262, N1239, N175, N50);
and AND3 (N1263, N1253, N28, N761);
and AND4 (N1264, N1251, N564, N554, N549);
not NOT1 (N1265, N1260);
nor NOR2 (N1266, N1259, N283);
or OR3 (N1267, N1266, N300, N610);
not NOT1 (N1268, N1241);
not NOT1 (N1269, N1258);
nand NAND3 (N1270, N1265, N1042, N57);
or OR4 (N1271, N1264, N1053, N660, N393);
nand NAND3 (N1272, N1268, N419, N2);
nand NAND4 (N1273, N1271, N354, N662, N211);
and AND2 (N1274, N1273, N8);
nand NAND3 (N1275, N1262, N222, N72);
buf BUF1 (N1276, N1269);
nor NOR2 (N1277, N1270, N371);
not NOT1 (N1278, N1263);
nand NAND4 (N1279, N1277, N1143, N1187, N441);
xor XOR2 (N1280, N1237, N686);
nand NAND2 (N1281, N1279, N624);
buf BUF1 (N1282, N1278);
or OR3 (N1283, N1281, N745, N1227);
nand NAND4 (N1284, N1256, N1218, N1077, N946);
or OR4 (N1285, N1261, N129, N837, N957);
xor XOR2 (N1286, N1267, N626);
or OR4 (N1287, N1284, N586, N715, N515);
or OR4 (N1288, N1286, N413, N738, N160);
xor XOR2 (N1289, N1287, N1271);
and AND4 (N1290, N1288, N373, N288, N931);
or OR2 (N1291, N1275, N670);
not NOT1 (N1292, N1283);
not NOT1 (N1293, N1292);
buf BUF1 (N1294, N1274);
and AND2 (N1295, N1294, N757);
or OR4 (N1296, N1272, N1204, N240, N391);
or OR4 (N1297, N1290, N618, N337, N264);
or OR2 (N1298, N1296, N708);
not NOT1 (N1299, N1285);
not NOT1 (N1300, N1298);
and AND2 (N1301, N1291, N959);
not NOT1 (N1302, N1297);
or OR2 (N1303, N1301, N612);
buf BUF1 (N1304, N1280);
nor NOR4 (N1305, N1282, N885, N481, N1300);
or OR4 (N1306, N361, N449, N64, N1147);
buf BUF1 (N1307, N1289);
and AND2 (N1308, N1305, N780);
nand NAND4 (N1309, N1307, N68, N312, N974);
and AND2 (N1310, N1276, N491);
xor XOR2 (N1311, N1306, N586);
and AND3 (N1312, N1303, N37, N472);
and AND4 (N1313, N1312, N1046, N753, N679);
and AND2 (N1314, N1311, N174);
xor XOR2 (N1315, N1293, N532);
not NOT1 (N1316, N1299);
xor XOR2 (N1317, N1310, N67);
xor XOR2 (N1318, N1302, N886);
or OR2 (N1319, N1295, N938);
nor NOR2 (N1320, N1314, N523);
xor XOR2 (N1321, N1319, N785);
or OR2 (N1322, N1304, N314);
nor NOR2 (N1323, N1321, N578);
buf BUF1 (N1324, N1318);
and AND3 (N1325, N1308, N132, N917);
nor NOR3 (N1326, N1316, N1208, N788);
buf BUF1 (N1327, N1313);
or OR4 (N1328, N1315, N1280, N752, N271);
or OR2 (N1329, N1328, N612);
nor NOR4 (N1330, N1323, N691, N268, N58);
nand NAND2 (N1331, N1320, N601);
nand NAND4 (N1332, N1330, N139, N1287, N939);
or OR3 (N1333, N1325, N554, N1043);
xor XOR2 (N1334, N1324, N749);
not NOT1 (N1335, N1331);
and AND2 (N1336, N1309, N379);
or OR2 (N1337, N1317, N1008);
xor XOR2 (N1338, N1337, N1052);
nand NAND4 (N1339, N1332, N2, N633, N296);
buf BUF1 (N1340, N1339);
or OR2 (N1341, N1334, N664);
xor XOR2 (N1342, N1340, N430);
nand NAND4 (N1343, N1322, N653, N365, N31);
xor XOR2 (N1344, N1326, N865);
and AND2 (N1345, N1342, N858);
not NOT1 (N1346, N1336);
nor NOR2 (N1347, N1344, N294);
buf BUF1 (N1348, N1341);
not NOT1 (N1349, N1345);
buf BUF1 (N1350, N1348);
nor NOR4 (N1351, N1350, N788, N432, N1085);
nor NOR4 (N1352, N1338, N47, N1127, N1061);
nor NOR2 (N1353, N1346, N994);
xor XOR2 (N1354, N1343, N863);
buf BUF1 (N1355, N1347);
xor XOR2 (N1356, N1351, N331);
xor XOR2 (N1357, N1356, N1199);
nor NOR4 (N1358, N1333, N289, N855, N30);
not NOT1 (N1359, N1354);
nand NAND4 (N1360, N1353, N116, N207, N900);
and AND3 (N1361, N1352, N200, N925);
xor XOR2 (N1362, N1329, N173);
and AND4 (N1363, N1362, N356, N1013, N555);
or OR4 (N1364, N1355, N34, N503, N1128);
and AND4 (N1365, N1327, N80, N856, N486);
and AND3 (N1366, N1358, N782, N553);
not NOT1 (N1367, N1359);
buf BUF1 (N1368, N1357);
not NOT1 (N1369, N1367);
nor NOR4 (N1370, N1363, N454, N292, N556);
xor XOR2 (N1371, N1349, N192);
nand NAND3 (N1372, N1364, N112, N861);
xor XOR2 (N1373, N1335, N900);
nor NOR3 (N1374, N1361, N449, N582);
and AND4 (N1375, N1366, N1201, N1111, N1126);
nor NOR3 (N1376, N1360, N503, N1067);
buf BUF1 (N1377, N1370);
nand NAND2 (N1378, N1371, N379);
or OR2 (N1379, N1375, N1139);
not NOT1 (N1380, N1372);
not NOT1 (N1381, N1379);
nor NOR2 (N1382, N1380, N750);
buf BUF1 (N1383, N1377);
and AND4 (N1384, N1369, N628, N1371, N1250);
and AND3 (N1385, N1368, N420, N952);
buf BUF1 (N1386, N1383);
or OR4 (N1387, N1382, N954, N195, N840);
not NOT1 (N1388, N1385);
nor NOR3 (N1389, N1381, N1031, N655);
nand NAND3 (N1390, N1365, N667, N983);
not NOT1 (N1391, N1389);
xor XOR2 (N1392, N1387, N485);
not NOT1 (N1393, N1390);
buf BUF1 (N1394, N1392);
buf BUF1 (N1395, N1376);
nand NAND4 (N1396, N1386, N690, N830, N1340);
or OR2 (N1397, N1396, N307);
or OR3 (N1398, N1397, N162, N1060);
nand NAND4 (N1399, N1388, N1011, N1040, N843);
or OR3 (N1400, N1391, N220, N837);
not NOT1 (N1401, N1374);
nor NOR2 (N1402, N1399, N1071);
or OR3 (N1403, N1402, N1366, N372);
xor XOR2 (N1404, N1393, N735);
and AND4 (N1405, N1394, N9, N1319, N372);
nand NAND4 (N1406, N1384, N1357, N440, N1357);
buf BUF1 (N1407, N1403);
buf BUF1 (N1408, N1395);
not NOT1 (N1409, N1398);
or OR2 (N1410, N1378, N952);
nand NAND4 (N1411, N1400, N652, N56, N1317);
not NOT1 (N1412, N1405);
not NOT1 (N1413, N1407);
nor NOR2 (N1414, N1412, N524);
or OR3 (N1415, N1406, N676, N89);
or OR3 (N1416, N1413, N362, N1327);
xor XOR2 (N1417, N1404, N395);
nand NAND4 (N1418, N1414, N258, N345, N697);
xor XOR2 (N1419, N1411, N747);
and AND2 (N1420, N1410, N817);
and AND2 (N1421, N1419, N489);
and AND4 (N1422, N1408, N671, N806, N614);
not NOT1 (N1423, N1422);
nand NAND4 (N1424, N1421, N791, N1215, N514);
xor XOR2 (N1425, N1418, N250);
nor NOR2 (N1426, N1373, N453);
and AND3 (N1427, N1426, N1293, N834);
or OR3 (N1428, N1417, N482, N1303);
or OR2 (N1429, N1427, N1132);
nor NOR4 (N1430, N1416, N1220, N485, N67);
nor NOR4 (N1431, N1425, N494, N1426, N135);
xor XOR2 (N1432, N1424, N13);
not NOT1 (N1433, N1431);
not NOT1 (N1434, N1430);
and AND2 (N1435, N1401, N944);
nand NAND4 (N1436, N1432, N737, N571, N1097);
buf BUF1 (N1437, N1423);
not NOT1 (N1438, N1435);
buf BUF1 (N1439, N1434);
buf BUF1 (N1440, N1429);
xor XOR2 (N1441, N1415, N326);
not NOT1 (N1442, N1441);
xor XOR2 (N1443, N1409, N971);
nor NOR3 (N1444, N1440, N960, N913);
or OR2 (N1445, N1428, N239);
xor XOR2 (N1446, N1437, N769);
not NOT1 (N1447, N1443);
nand NAND3 (N1448, N1445, N7, N917);
nand NAND2 (N1449, N1433, N895);
buf BUF1 (N1450, N1438);
buf BUF1 (N1451, N1449);
xor XOR2 (N1452, N1451, N1350);
buf BUF1 (N1453, N1439);
nand NAND2 (N1454, N1444, N890);
nor NOR3 (N1455, N1453, N1061, N74);
not NOT1 (N1456, N1446);
xor XOR2 (N1457, N1448, N823);
nor NOR2 (N1458, N1452, N135);
nor NOR3 (N1459, N1457, N1405, N1292);
and AND3 (N1460, N1420, N1367, N1384);
and AND3 (N1461, N1447, N1401, N426);
xor XOR2 (N1462, N1461, N470);
buf BUF1 (N1463, N1442);
nor NOR3 (N1464, N1460, N1009, N505);
or OR2 (N1465, N1462, N236);
not NOT1 (N1466, N1459);
and AND4 (N1467, N1458, N439, N198, N767);
nor NOR2 (N1468, N1463, N560);
xor XOR2 (N1469, N1465, N607);
not NOT1 (N1470, N1466);
not NOT1 (N1471, N1454);
buf BUF1 (N1472, N1456);
nand NAND4 (N1473, N1467, N409, N1143, N998);
and AND3 (N1474, N1472, N1426, N204);
buf BUF1 (N1475, N1468);
not NOT1 (N1476, N1473);
nor NOR2 (N1477, N1450, N197);
buf BUF1 (N1478, N1455);
nor NOR3 (N1479, N1474, N1128, N241);
xor XOR2 (N1480, N1479, N848);
or OR3 (N1481, N1469, N852, N353);
nand NAND4 (N1482, N1436, N214, N195, N90);
xor XOR2 (N1483, N1464, N1205);
not NOT1 (N1484, N1475);
buf BUF1 (N1485, N1483);
nor NOR3 (N1486, N1480, N287, N1259);
not NOT1 (N1487, N1482);
not NOT1 (N1488, N1481);
xor XOR2 (N1489, N1485, N1087);
xor XOR2 (N1490, N1478, N531);
and AND4 (N1491, N1470, N1010, N526, N1440);
or OR2 (N1492, N1490, N1289);
nand NAND2 (N1493, N1492, N1358);
xor XOR2 (N1494, N1489, N1064);
xor XOR2 (N1495, N1484, N1014);
not NOT1 (N1496, N1471);
nand NAND3 (N1497, N1488, N1302, N1022);
and AND2 (N1498, N1493, N480);
buf BUF1 (N1499, N1476);
buf BUF1 (N1500, N1498);
and AND3 (N1501, N1500, N372, N368);
or OR3 (N1502, N1496, N931, N753);
nand NAND4 (N1503, N1494, N450, N1327, N776);
nor NOR3 (N1504, N1495, N247, N165);
or OR3 (N1505, N1487, N635, N282);
or OR3 (N1506, N1486, N1489, N1325);
not NOT1 (N1507, N1491);
not NOT1 (N1508, N1505);
not NOT1 (N1509, N1503);
or OR2 (N1510, N1508, N1504);
buf BUF1 (N1511, N10);
or OR2 (N1512, N1477, N568);
and AND3 (N1513, N1511, N1106, N563);
buf BUF1 (N1514, N1512);
not NOT1 (N1515, N1499);
xor XOR2 (N1516, N1510, N435);
nand NAND2 (N1517, N1497, N1456);
nand NAND2 (N1518, N1516, N1370);
and AND2 (N1519, N1507, N41);
not NOT1 (N1520, N1506);
nor NOR3 (N1521, N1501, N672, N1213);
buf BUF1 (N1522, N1502);
nand NAND4 (N1523, N1509, N37, N59, N550);
and AND2 (N1524, N1522, N55);
and AND3 (N1525, N1515, N914, N1347);
not NOT1 (N1526, N1524);
or OR2 (N1527, N1526, N419);
xor XOR2 (N1528, N1520, N1487);
or OR3 (N1529, N1528, N477, N462);
nand NAND2 (N1530, N1527, N472);
or OR2 (N1531, N1518, N431);
xor XOR2 (N1532, N1523, N1140);
nor NOR3 (N1533, N1514, N1433, N1134);
xor XOR2 (N1534, N1530, N138);
xor XOR2 (N1535, N1531, N88);
nand NAND3 (N1536, N1513, N1460, N213);
nand NAND3 (N1537, N1535, N1166, N1357);
nor NOR2 (N1538, N1533, N1074);
xor XOR2 (N1539, N1529, N635);
and AND2 (N1540, N1538, N966);
or OR2 (N1541, N1532, N1345);
nand NAND4 (N1542, N1534, N820, N1308, N65);
xor XOR2 (N1543, N1521, N237);
nand NAND2 (N1544, N1519, N62);
buf BUF1 (N1545, N1536);
not NOT1 (N1546, N1539);
buf BUF1 (N1547, N1542);
or OR2 (N1548, N1525, N19);
xor XOR2 (N1549, N1537, N1372);
xor XOR2 (N1550, N1517, N73);
or OR3 (N1551, N1546, N1048, N642);
not NOT1 (N1552, N1550);
nand NAND4 (N1553, N1549, N701, N1464, N152);
and AND3 (N1554, N1551, N1149, N1507);
and AND3 (N1555, N1543, N354, N1395);
not NOT1 (N1556, N1541);
or OR4 (N1557, N1540, N359, N721, N1556);
nor NOR2 (N1558, N1145, N81);
not NOT1 (N1559, N1544);
buf BUF1 (N1560, N1548);
buf BUF1 (N1561, N1558);
nand NAND3 (N1562, N1552, N331, N524);
nor NOR3 (N1563, N1555, N45, N1067);
nor NOR3 (N1564, N1562, N986, N1304);
or OR2 (N1565, N1563, N1363);
buf BUF1 (N1566, N1565);
nor NOR2 (N1567, N1561, N900);
not NOT1 (N1568, N1566);
nor NOR4 (N1569, N1545, N578, N672, N569);
not NOT1 (N1570, N1553);
or OR3 (N1571, N1570, N670, N1312);
or OR3 (N1572, N1568, N253, N241);
buf BUF1 (N1573, N1560);
nor NOR4 (N1574, N1564, N183, N1214, N157);
not NOT1 (N1575, N1559);
nand NAND3 (N1576, N1547, N1364, N404);
nand NAND4 (N1577, N1557, N871, N705, N668);
or OR2 (N1578, N1571, N1273);
nor NOR2 (N1579, N1567, N1067);
nand NAND4 (N1580, N1577, N1425, N636, N203);
nor NOR3 (N1581, N1580, N1293, N625);
xor XOR2 (N1582, N1579, N1523);
and AND3 (N1583, N1554, N1341, N1216);
nand NAND4 (N1584, N1578, N394, N57, N1178);
buf BUF1 (N1585, N1569);
and AND4 (N1586, N1574, N567, N456, N683);
or OR3 (N1587, N1585, N988, N623);
nand NAND4 (N1588, N1587, N1210, N1492, N918);
buf BUF1 (N1589, N1588);
not NOT1 (N1590, N1582);
nand NAND2 (N1591, N1583, N741);
not NOT1 (N1592, N1572);
nor NOR3 (N1593, N1576, N950, N555);
nor NOR4 (N1594, N1592, N1467, N1216, N7);
nor NOR3 (N1595, N1584, N993, N642);
or OR3 (N1596, N1581, N445, N670);
not NOT1 (N1597, N1593);
xor XOR2 (N1598, N1590, N1569);
xor XOR2 (N1599, N1575, N132);
xor XOR2 (N1600, N1586, N74);
or OR4 (N1601, N1600, N301, N718, N489);
xor XOR2 (N1602, N1594, N1497);
nor NOR2 (N1603, N1601, N842);
nor NOR2 (N1604, N1591, N48);
or OR2 (N1605, N1595, N641);
nand NAND3 (N1606, N1589, N942, N131);
buf BUF1 (N1607, N1573);
nor NOR2 (N1608, N1602, N317);
nor NOR4 (N1609, N1605, N78, N1582, N1333);
nand NAND4 (N1610, N1598, N1010, N58, N723);
xor XOR2 (N1611, N1603, N656);
nor NOR2 (N1612, N1597, N46);
buf BUF1 (N1613, N1606);
xor XOR2 (N1614, N1612, N997);
not NOT1 (N1615, N1607);
buf BUF1 (N1616, N1614);
and AND4 (N1617, N1609, N207, N240, N507);
or OR3 (N1618, N1611, N27, N455);
not NOT1 (N1619, N1616);
xor XOR2 (N1620, N1608, N78);
buf BUF1 (N1621, N1613);
buf BUF1 (N1622, N1617);
not NOT1 (N1623, N1615);
not NOT1 (N1624, N1610);
not NOT1 (N1625, N1620);
buf BUF1 (N1626, N1623);
xor XOR2 (N1627, N1618, N844);
or OR3 (N1628, N1627, N1374, N1337);
nor NOR4 (N1629, N1622, N1013, N771, N863);
or OR2 (N1630, N1629, N1402);
not NOT1 (N1631, N1624);
buf BUF1 (N1632, N1596);
and AND2 (N1633, N1626, N810);
not NOT1 (N1634, N1632);
xor XOR2 (N1635, N1633, N169);
nand NAND3 (N1636, N1631, N667, N432);
nor NOR3 (N1637, N1635, N744, N859);
and AND3 (N1638, N1621, N1091, N563);
xor XOR2 (N1639, N1628, N917);
buf BUF1 (N1640, N1630);
not NOT1 (N1641, N1637);
nand NAND3 (N1642, N1619, N1334, N1538);
buf BUF1 (N1643, N1625);
or OR4 (N1644, N1643, N1625, N583, N713);
buf BUF1 (N1645, N1644);
nor NOR2 (N1646, N1639, N735);
buf BUF1 (N1647, N1638);
and AND3 (N1648, N1641, N698, N146);
not NOT1 (N1649, N1634);
nand NAND4 (N1650, N1640, N1462, N1011, N1407);
buf BUF1 (N1651, N1636);
nand NAND4 (N1652, N1604, N763, N1230, N636);
xor XOR2 (N1653, N1650, N344);
and AND4 (N1654, N1647, N400, N1606, N746);
nand NAND2 (N1655, N1648, N1499);
buf BUF1 (N1656, N1654);
buf BUF1 (N1657, N1642);
and AND2 (N1658, N1599, N1330);
xor XOR2 (N1659, N1657, N993);
xor XOR2 (N1660, N1649, N97);
xor XOR2 (N1661, N1656, N570);
or OR2 (N1662, N1655, N311);
xor XOR2 (N1663, N1646, N580);
or OR3 (N1664, N1659, N415, N1341);
nor NOR2 (N1665, N1645, N1375);
xor XOR2 (N1666, N1652, N1312);
buf BUF1 (N1667, N1666);
nand NAND2 (N1668, N1660, N321);
xor XOR2 (N1669, N1662, N745);
nor NOR2 (N1670, N1668, N1594);
xor XOR2 (N1671, N1653, N1080);
nor NOR2 (N1672, N1658, N489);
and AND2 (N1673, N1671, N617);
not NOT1 (N1674, N1667);
not NOT1 (N1675, N1672);
nor NOR3 (N1676, N1674, N1412, N747);
not NOT1 (N1677, N1661);
or OR2 (N1678, N1664, N1156);
buf BUF1 (N1679, N1678);
xor XOR2 (N1680, N1675, N1169);
nor NOR2 (N1681, N1663, N1632);
buf BUF1 (N1682, N1680);
not NOT1 (N1683, N1677);
not NOT1 (N1684, N1669);
nor NOR3 (N1685, N1683, N499, N1574);
or OR2 (N1686, N1670, N1193);
nand NAND2 (N1687, N1676, N1065);
xor XOR2 (N1688, N1687, N1236);
xor XOR2 (N1689, N1684, N1135);
xor XOR2 (N1690, N1686, N709);
nor NOR2 (N1691, N1688, N148);
nor NOR3 (N1692, N1685, N576, N1589);
nand NAND3 (N1693, N1651, N1188, N415);
and AND4 (N1694, N1692, N1035, N1544, N1595);
nand NAND3 (N1695, N1673, N1258, N1074);
nand NAND4 (N1696, N1693, N597, N1214, N1038);
nand NAND2 (N1697, N1691, N438);
or OR3 (N1698, N1681, N495, N221);
and AND3 (N1699, N1696, N495, N1149);
or OR3 (N1700, N1697, N965, N1588);
or OR2 (N1701, N1695, N599);
not NOT1 (N1702, N1689);
xor XOR2 (N1703, N1702, N1171);
nand NAND3 (N1704, N1690, N841, N588);
buf BUF1 (N1705, N1704);
buf BUF1 (N1706, N1700);
or OR4 (N1707, N1699, N495, N979, N500);
not NOT1 (N1708, N1701);
nand NAND4 (N1709, N1706, N1157, N409, N695);
xor XOR2 (N1710, N1698, N412);
nand NAND4 (N1711, N1665, N442, N1329, N1402);
buf BUF1 (N1712, N1709);
nor NOR2 (N1713, N1707, N548);
nand NAND3 (N1714, N1705, N1498, N878);
and AND3 (N1715, N1713, N1703, N1294);
buf BUF1 (N1716, N1408);
nand NAND2 (N1717, N1716, N8);
xor XOR2 (N1718, N1712, N1450);
buf BUF1 (N1719, N1711);
nor NOR3 (N1720, N1694, N1543, N388);
not NOT1 (N1721, N1715);
xor XOR2 (N1722, N1718, N996);
or OR3 (N1723, N1679, N529, N363);
xor XOR2 (N1724, N1714, N665);
not NOT1 (N1725, N1717);
not NOT1 (N1726, N1721);
or OR3 (N1727, N1682, N989, N1397);
not NOT1 (N1728, N1724);
not NOT1 (N1729, N1722);
nor NOR2 (N1730, N1708, N702);
nor NOR3 (N1731, N1719, N629, N840);
xor XOR2 (N1732, N1723, N1534);
buf BUF1 (N1733, N1728);
and AND2 (N1734, N1733, N1523);
not NOT1 (N1735, N1731);
not NOT1 (N1736, N1727);
or OR2 (N1737, N1732, N1266);
nand NAND3 (N1738, N1736, N1164, N684);
buf BUF1 (N1739, N1720);
buf BUF1 (N1740, N1726);
or OR3 (N1741, N1730, N216, N712);
buf BUF1 (N1742, N1739);
nand NAND4 (N1743, N1737, N313, N862, N796);
and AND3 (N1744, N1738, N660, N1286);
nand NAND3 (N1745, N1710, N705, N601);
not NOT1 (N1746, N1735);
nor NOR3 (N1747, N1729, N1076, N1501);
buf BUF1 (N1748, N1734);
nor NOR3 (N1749, N1748, N1047, N444);
xor XOR2 (N1750, N1749, N764);
and AND3 (N1751, N1741, N41, N1130);
buf BUF1 (N1752, N1740);
nand NAND4 (N1753, N1746, N1603, N337, N1122);
not NOT1 (N1754, N1743);
buf BUF1 (N1755, N1751);
nand NAND2 (N1756, N1745, N70);
nand NAND4 (N1757, N1744, N1624, N1359, N1348);
nor NOR2 (N1758, N1756, N942);
nor NOR2 (N1759, N1753, N872);
and AND4 (N1760, N1758, N1031, N1399, N1108);
nand NAND2 (N1761, N1747, N208);
xor XOR2 (N1762, N1759, N855);
and AND4 (N1763, N1725, N1488, N825, N997);
not NOT1 (N1764, N1752);
nand NAND4 (N1765, N1762, N393, N5, N1557);
and AND4 (N1766, N1750, N1190, N414, N834);
buf BUF1 (N1767, N1765);
nand NAND3 (N1768, N1761, N103, N612);
or OR2 (N1769, N1767, N199);
nand NAND4 (N1770, N1757, N608, N657, N1597);
or OR4 (N1771, N1770, N751, N267, N1056);
buf BUF1 (N1772, N1763);
buf BUF1 (N1773, N1769);
nor NOR4 (N1774, N1742, N397, N1647, N916);
or OR3 (N1775, N1764, N796, N158);
and AND3 (N1776, N1768, N1408, N348);
not NOT1 (N1777, N1771);
not NOT1 (N1778, N1760);
nand NAND4 (N1779, N1777, N35, N1426, N1086);
nand NAND2 (N1780, N1772, N1677);
or OR2 (N1781, N1778, N1493);
nor NOR2 (N1782, N1780, N1525);
xor XOR2 (N1783, N1775, N175);
xor XOR2 (N1784, N1782, N76);
buf BUF1 (N1785, N1783);
nand NAND4 (N1786, N1754, N81, N1757, N1345);
not NOT1 (N1787, N1776);
xor XOR2 (N1788, N1774, N1520);
buf BUF1 (N1789, N1785);
and AND4 (N1790, N1784, N1062, N576, N1435);
and AND2 (N1791, N1766, N786);
not NOT1 (N1792, N1789);
not NOT1 (N1793, N1790);
nor NOR4 (N1794, N1755, N901, N945, N81);
nand NAND3 (N1795, N1779, N1769, N41);
or OR2 (N1796, N1788, N1176);
buf BUF1 (N1797, N1791);
or OR2 (N1798, N1793, N74);
xor XOR2 (N1799, N1798, N1138);
not NOT1 (N1800, N1786);
and AND2 (N1801, N1796, N876);
xor XOR2 (N1802, N1799, N930);
nand NAND3 (N1803, N1787, N1477, N259);
not NOT1 (N1804, N1801);
not NOT1 (N1805, N1804);
buf BUF1 (N1806, N1792);
buf BUF1 (N1807, N1806);
or OR2 (N1808, N1797, N1157);
and AND2 (N1809, N1794, N1186);
nor NOR2 (N1810, N1807, N977);
xor XOR2 (N1811, N1795, N335);
xor XOR2 (N1812, N1810, N948);
or OR3 (N1813, N1781, N1024, N1105);
xor XOR2 (N1814, N1773, N821);
xor XOR2 (N1815, N1811, N245);
buf BUF1 (N1816, N1812);
nor NOR3 (N1817, N1808, N1597, N1729);
nand NAND2 (N1818, N1815, N1569);
xor XOR2 (N1819, N1817, N1022);
buf BUF1 (N1820, N1800);
or OR2 (N1821, N1809, N1195);
nand NAND3 (N1822, N1805, N818, N41);
nor NOR2 (N1823, N1814, N1265);
buf BUF1 (N1824, N1822);
nand NAND2 (N1825, N1823, N1524);
nor NOR4 (N1826, N1821, N399, N59, N1382);
buf BUF1 (N1827, N1824);
xor XOR2 (N1828, N1825, N1281);
and AND4 (N1829, N1827, N427, N1126, N248);
nor NOR2 (N1830, N1816, N1215);
nand NAND4 (N1831, N1826, N784, N222, N447);
buf BUF1 (N1832, N1813);
nand NAND3 (N1833, N1832, N1140, N825);
or OR2 (N1834, N1819, N614);
or OR2 (N1835, N1831, N1385);
or OR4 (N1836, N1829, N1305, N1483, N329);
buf BUF1 (N1837, N1802);
or OR2 (N1838, N1834, N1051);
not NOT1 (N1839, N1838);
and AND2 (N1840, N1818, N1748);
or OR3 (N1841, N1820, N1045, N1562);
nand NAND2 (N1842, N1833, N1124);
not NOT1 (N1843, N1836);
and AND4 (N1844, N1840, N944, N1272, N554);
or OR2 (N1845, N1830, N470);
not NOT1 (N1846, N1841);
or OR3 (N1847, N1842, N1661, N933);
not NOT1 (N1848, N1828);
xor XOR2 (N1849, N1845, N618);
nor NOR3 (N1850, N1844, N1239, N911);
nor NOR4 (N1851, N1850, N1235, N195, N1582);
nand NAND4 (N1852, N1803, N1766, N1796, N1438);
buf BUF1 (N1853, N1847);
buf BUF1 (N1854, N1851);
not NOT1 (N1855, N1849);
nand NAND2 (N1856, N1855, N552);
not NOT1 (N1857, N1854);
and AND3 (N1858, N1839, N302, N1367);
and AND2 (N1859, N1857, N1070);
xor XOR2 (N1860, N1852, N810);
buf BUF1 (N1861, N1837);
or OR4 (N1862, N1848, N1860, N249, N1335);
buf BUF1 (N1863, N1330);
nand NAND3 (N1864, N1863, N42, N922);
or OR2 (N1865, N1862, N1858);
or OR3 (N1866, N1240, N778, N386);
not NOT1 (N1867, N1856);
buf BUF1 (N1868, N1864);
nor NOR3 (N1869, N1846, N1567, N430);
not NOT1 (N1870, N1843);
and AND2 (N1871, N1870, N1099);
not NOT1 (N1872, N1859);
and AND2 (N1873, N1872, N618);
nor NOR4 (N1874, N1835, N1804, N1374, N1188);
not NOT1 (N1875, N1874);
nand NAND4 (N1876, N1865, N985, N1840, N1310);
and AND2 (N1877, N1875, N542);
nor NOR2 (N1878, N1867, N505);
nor NOR4 (N1879, N1869, N80, N602, N706);
or OR2 (N1880, N1866, N444);
or OR3 (N1881, N1877, N1012, N297);
and AND2 (N1882, N1876, N1292);
nand NAND4 (N1883, N1868, N655, N687, N464);
xor XOR2 (N1884, N1882, N127);
nand NAND4 (N1885, N1861, N552, N1671, N782);
not NOT1 (N1886, N1883);
or OR4 (N1887, N1880, N474, N882, N1285);
nor NOR3 (N1888, N1886, N30, N1553);
buf BUF1 (N1889, N1887);
xor XOR2 (N1890, N1853, N1367);
xor XOR2 (N1891, N1879, N655);
not NOT1 (N1892, N1881);
nand NAND3 (N1893, N1878, N1742, N967);
buf BUF1 (N1894, N1888);
nor NOR2 (N1895, N1892, N1140);
not NOT1 (N1896, N1884);
xor XOR2 (N1897, N1890, N379);
xor XOR2 (N1898, N1891, N1);
buf BUF1 (N1899, N1871);
and AND3 (N1900, N1898, N1130, N537);
and AND2 (N1901, N1900, N1103);
nor NOR4 (N1902, N1901, N33, N1636, N645);
buf BUF1 (N1903, N1895);
xor XOR2 (N1904, N1903, N1560);
nand NAND3 (N1905, N1889, N1226, N1445);
xor XOR2 (N1906, N1885, N937);
or OR2 (N1907, N1896, N879);
xor XOR2 (N1908, N1897, N1124);
and AND4 (N1909, N1894, N1679, N6, N212);
or OR4 (N1910, N1908, N69, N169, N1219);
or OR3 (N1911, N1906, N673, N1816);
not NOT1 (N1912, N1911);
nor NOR2 (N1913, N1907, N1527);
not NOT1 (N1914, N1905);
nor NOR3 (N1915, N1914, N562, N2);
buf BUF1 (N1916, N1909);
or OR3 (N1917, N1912, N136, N755);
nor NOR3 (N1918, N1917, N1546, N1795);
nand NAND3 (N1919, N1893, N991, N653);
buf BUF1 (N1920, N1873);
or OR2 (N1921, N1919, N1445);
not NOT1 (N1922, N1913);
nand NAND4 (N1923, N1902, N170, N641, N894);
nand NAND2 (N1924, N1916, N1130);
not NOT1 (N1925, N1915);
nor NOR3 (N1926, N1899, N1375, N277);
and AND4 (N1927, N1926, N162, N1407, N1514);
nor NOR4 (N1928, N1921, N1627, N1631, N197);
buf BUF1 (N1929, N1910);
and AND3 (N1930, N1924, N85, N1587);
buf BUF1 (N1931, N1930);
and AND3 (N1932, N1925, N1648, N1299);
buf BUF1 (N1933, N1931);
nor NOR4 (N1934, N1904, N1871, N135, N275);
not NOT1 (N1935, N1918);
nand NAND2 (N1936, N1935, N1825);
buf BUF1 (N1937, N1932);
and AND2 (N1938, N1933, N202);
buf BUF1 (N1939, N1928);
or OR4 (N1940, N1934, N1634, N519, N1922);
not NOT1 (N1941, N870);
or OR2 (N1942, N1929, N1796);
buf BUF1 (N1943, N1937);
or OR2 (N1944, N1941, N1184);
xor XOR2 (N1945, N1940, N1128);
and AND3 (N1946, N1939, N565, N1768);
buf BUF1 (N1947, N1946);
xor XOR2 (N1948, N1923, N1924);
buf BUF1 (N1949, N1947);
and AND3 (N1950, N1936, N1469, N1899);
not NOT1 (N1951, N1950);
or OR3 (N1952, N1951, N1727, N581);
xor XOR2 (N1953, N1927, N1884);
nand NAND3 (N1954, N1949, N102, N1784);
xor XOR2 (N1955, N1948, N364);
not NOT1 (N1956, N1938);
buf BUF1 (N1957, N1954);
and AND4 (N1958, N1956, N1678, N454, N1399);
nor NOR3 (N1959, N1953, N1291, N561);
or OR3 (N1960, N1944, N496, N650);
buf BUF1 (N1961, N1960);
or OR4 (N1962, N1957, N88, N1180, N800);
xor XOR2 (N1963, N1920, N1619);
nor NOR2 (N1964, N1961, N1378);
xor XOR2 (N1965, N1945, N459);
or OR2 (N1966, N1955, N595);
xor XOR2 (N1967, N1966, N1031);
xor XOR2 (N1968, N1963, N1260);
nor NOR2 (N1969, N1962, N106);
xor XOR2 (N1970, N1967, N1501);
xor XOR2 (N1971, N1959, N509);
and AND2 (N1972, N1971, N287);
and AND2 (N1973, N1952, N682);
not NOT1 (N1974, N1969);
and AND2 (N1975, N1958, N1268);
or OR4 (N1976, N1965, N1421, N1726, N338);
buf BUF1 (N1977, N1968);
buf BUF1 (N1978, N1976);
xor XOR2 (N1979, N1974, N654);
and AND4 (N1980, N1977, N1370, N1261, N1672);
not NOT1 (N1981, N1979);
nor NOR3 (N1982, N1978, N833, N47);
nor NOR4 (N1983, N1982, N159, N667, N1184);
not NOT1 (N1984, N1980);
nand NAND3 (N1985, N1981, N693, N1116);
and AND3 (N1986, N1972, N231, N601);
not NOT1 (N1987, N1986);
nor NOR3 (N1988, N1983, N40, N780);
buf BUF1 (N1989, N1943);
nand NAND2 (N1990, N1970, N1283);
nand NAND2 (N1991, N1987, N71);
or OR2 (N1992, N1988, N1572);
or OR4 (N1993, N1989, N955, N1486, N1260);
and AND4 (N1994, N1984, N129, N1306, N506);
or OR2 (N1995, N1992, N1706);
nor NOR4 (N1996, N1985, N433, N1861, N306);
not NOT1 (N1997, N1993);
nand NAND2 (N1998, N1995, N124);
nor NOR4 (N1999, N1942, N1782, N885, N293);
nand NAND3 (N2000, N1973, N1198, N181);
xor XOR2 (N2001, N1975, N1557);
nor NOR3 (N2002, N1964, N777, N1022);
nor NOR2 (N2003, N1997, N1550);
buf BUF1 (N2004, N1998);
buf BUF1 (N2005, N2000);
or OR2 (N2006, N1991, N1975);
xor XOR2 (N2007, N2005, N470);
not NOT1 (N2008, N2002);
buf BUF1 (N2009, N1994);
and AND2 (N2010, N2009, N1792);
endmodule