// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13;

output N512,N507,N506,N500,N492,N489,N511,N510,N509,N513;

and AND4 (N14, N7, N12, N10, N4);
xor XOR2 (N15, N11, N3);
nand NAND3 (N16, N10, N15, N7);
buf BUF1 (N17, N16);
or OR4 (N18, N9, N16, N3, N16);
xor XOR2 (N19, N15, N11);
or OR4 (N20, N17, N9, N15, N13);
nor NOR2 (N21, N7, N11);
xor XOR2 (N22, N21, N1);
buf BUF1 (N23, N8);
not NOT1 (N24, N17);
nor NOR3 (N25, N21, N19, N1);
nand NAND2 (N26, N15, N23);
or OR3 (N27, N16, N26, N6);
nor NOR4 (N28, N4, N19, N8, N17);
and AND4 (N29, N2, N4, N11, N20);
buf BUF1 (N30, N17);
and AND4 (N31, N22, N26, N2, N9);
buf BUF1 (N32, N7);
buf BUF1 (N33, N28);
and AND3 (N34, N25, N4, N20);
nand NAND2 (N35, N14, N8);
not NOT1 (N36, N34);
and AND3 (N37, N35, N5, N24);
nand NAND3 (N38, N14, N4, N32);
not NOT1 (N39, N2);
buf BUF1 (N40, N38);
nand NAND3 (N41, N27, N11, N32);
and AND3 (N42, N37, N22, N32);
xor XOR2 (N43, N31, N9);
or OR4 (N44, N42, N31, N1, N6);
buf BUF1 (N45, N36);
xor XOR2 (N46, N39, N37);
buf BUF1 (N47, N44);
nor NOR2 (N48, N41, N4);
buf BUF1 (N49, N29);
nand NAND2 (N50, N40, N26);
nor NOR3 (N51, N30, N31, N30);
and AND3 (N52, N45, N20, N38);
or OR2 (N53, N47, N18);
and AND2 (N54, N49, N8);
nor NOR3 (N55, N2, N27, N25);
nor NOR2 (N56, N53, N47);
buf BUF1 (N57, N43);
buf BUF1 (N58, N33);
nor NOR4 (N59, N51, N57, N7, N32);
not NOT1 (N60, N41);
not NOT1 (N61, N56);
buf BUF1 (N62, N52);
not NOT1 (N63, N58);
and AND3 (N64, N59, N59, N4);
xor XOR2 (N65, N46, N42);
or OR2 (N66, N64, N55);
nand NAND4 (N67, N33, N35, N12, N22);
not NOT1 (N68, N48);
xor XOR2 (N69, N63, N61);
not NOT1 (N70, N12);
nand NAND4 (N71, N62, N61, N58, N11);
not NOT1 (N72, N65);
buf BUF1 (N73, N70);
not NOT1 (N74, N60);
not NOT1 (N75, N67);
nor NOR3 (N76, N72, N70, N34);
nand NAND2 (N77, N75, N16);
nand NAND4 (N78, N71, N8, N15, N24);
buf BUF1 (N79, N77);
and AND4 (N80, N76, N19, N9, N16);
or OR2 (N81, N79, N22);
or OR2 (N82, N74, N76);
buf BUF1 (N83, N54);
xor XOR2 (N84, N50, N69);
not NOT1 (N85, N4);
and AND4 (N86, N80, N84, N53, N30);
and AND2 (N87, N70, N51);
buf BUF1 (N88, N73);
xor XOR2 (N89, N81, N4);
xor XOR2 (N90, N68, N44);
nor NOR3 (N91, N88, N2, N22);
not NOT1 (N92, N82);
nor NOR3 (N93, N92, N89, N47);
and AND4 (N94, N25, N75, N48, N36);
buf BUF1 (N95, N66);
xor XOR2 (N96, N91, N40);
xor XOR2 (N97, N83, N49);
buf BUF1 (N98, N96);
not NOT1 (N99, N85);
not NOT1 (N100, N78);
xor XOR2 (N101, N90, N55);
nand NAND4 (N102, N97, N12, N48, N101);
xor XOR2 (N103, N27, N74);
buf BUF1 (N104, N93);
and AND2 (N105, N95, N50);
xor XOR2 (N106, N86, N63);
nand NAND3 (N107, N105, N36, N2);
or OR4 (N108, N98, N55, N63, N30);
xor XOR2 (N109, N94, N105);
and AND3 (N110, N87, N36, N12);
and AND2 (N111, N103, N105);
nor NOR2 (N112, N108, N12);
or OR4 (N113, N99, N76, N17, N107);
xor XOR2 (N114, N63, N21);
and AND2 (N115, N113, N50);
xor XOR2 (N116, N102, N64);
nand NAND2 (N117, N115, N21);
or OR3 (N118, N112, N57, N4);
nand NAND2 (N119, N117, N60);
xor XOR2 (N120, N118, N116);
and AND4 (N121, N64, N57, N27, N60);
xor XOR2 (N122, N121, N70);
buf BUF1 (N123, N109);
xor XOR2 (N124, N106, N21);
xor XOR2 (N125, N111, N30);
buf BUF1 (N126, N110);
and AND4 (N127, N104, N30, N94, N26);
buf BUF1 (N128, N120);
nand NAND4 (N129, N127, N17, N59, N114);
nand NAND2 (N130, N22, N86);
xor XOR2 (N131, N130, N5);
not NOT1 (N132, N125);
not NOT1 (N133, N132);
nor NOR3 (N134, N129, N121, N1);
nand NAND2 (N135, N119, N70);
and AND4 (N136, N131, N51, N93, N113);
buf BUF1 (N137, N134);
nor NOR2 (N138, N133, N14);
xor XOR2 (N139, N124, N98);
or OR3 (N140, N137, N139, N58);
and AND4 (N141, N48, N7, N77, N37);
or OR4 (N142, N135, N101, N93, N28);
and AND2 (N143, N138, N88);
nor NOR4 (N144, N123, N39, N56, N72);
nor NOR2 (N145, N144, N123);
not NOT1 (N146, N128);
nand NAND2 (N147, N141, N71);
xor XOR2 (N148, N136, N140);
nand NAND4 (N149, N120, N97, N37, N112);
and AND2 (N150, N122, N3);
xor XOR2 (N151, N145, N89);
not NOT1 (N152, N100);
or OR2 (N153, N149, N122);
and AND2 (N154, N148, N36);
or OR2 (N155, N146, N55);
or OR2 (N156, N126, N26);
or OR2 (N157, N152, N75);
and AND4 (N158, N155, N85, N26, N124);
and AND4 (N159, N156, N25, N48, N99);
buf BUF1 (N160, N151);
not NOT1 (N161, N142);
nand NAND2 (N162, N143, N124);
buf BUF1 (N163, N159);
and AND4 (N164, N163, N3, N159, N19);
xor XOR2 (N165, N164, N78);
buf BUF1 (N166, N150);
nor NOR3 (N167, N165, N19, N18);
buf BUF1 (N168, N153);
buf BUF1 (N169, N166);
and AND3 (N170, N168, N130, N95);
or OR2 (N171, N154, N72);
nand NAND3 (N172, N147, N142, N151);
and AND2 (N173, N172, N45);
not NOT1 (N174, N173);
and AND4 (N175, N169, N164, N118, N9);
nand NAND2 (N176, N175, N157);
xor XOR2 (N177, N37, N6);
nor NOR2 (N178, N176, N167);
nor NOR2 (N179, N141, N54);
not NOT1 (N180, N158);
or OR4 (N181, N177, N32, N44, N160);
and AND2 (N182, N7, N113);
or OR3 (N183, N179, N88, N45);
or OR3 (N184, N170, N147, N70);
or OR4 (N185, N171, N7, N104, N12);
not NOT1 (N186, N183);
nor NOR2 (N187, N182, N2);
nor NOR3 (N188, N161, N1, N24);
and AND3 (N189, N162, N184, N1);
or OR4 (N190, N68, N148, N81, N41);
buf BUF1 (N191, N181);
nor NOR4 (N192, N190, N43, N85, N96);
nor NOR3 (N193, N192, N78, N113);
nor NOR2 (N194, N188, N108);
or OR3 (N195, N185, N86, N64);
xor XOR2 (N196, N195, N92);
nor NOR3 (N197, N193, N148, N82);
xor XOR2 (N198, N189, N27);
or OR4 (N199, N187, N147, N34, N186);
not NOT1 (N200, N68);
nor NOR3 (N201, N174, N126, N75);
xor XOR2 (N202, N198, N50);
xor XOR2 (N203, N178, N18);
and AND4 (N204, N197, N45, N177, N151);
or OR4 (N205, N199, N106, N70, N79);
nand NAND3 (N206, N196, N165, N76);
nand NAND4 (N207, N204, N11, N102, N45);
not NOT1 (N208, N202);
nor NOR4 (N209, N180, N200, N42, N172);
xor XOR2 (N210, N8, N195);
or OR4 (N211, N209, N34, N56, N5);
not NOT1 (N212, N207);
nand NAND3 (N213, N212, N99, N114);
and AND3 (N214, N203, N135, N118);
nand NAND4 (N215, N208, N177, N214, N46);
not NOT1 (N216, N31);
xor XOR2 (N217, N201, N131);
and AND2 (N218, N216, N111);
nor NOR4 (N219, N218, N55, N218, N29);
nand NAND3 (N220, N194, N160, N177);
xor XOR2 (N221, N191, N166);
not NOT1 (N222, N210);
nor NOR3 (N223, N221, N55, N19);
nor NOR2 (N224, N215, N101);
nand NAND4 (N225, N213, N154, N135, N81);
or OR4 (N226, N206, N141, N51, N220);
or OR4 (N227, N43, N89, N127, N118);
and AND2 (N228, N211, N194);
nor NOR3 (N229, N217, N199, N37);
xor XOR2 (N230, N222, N67);
buf BUF1 (N231, N229);
and AND2 (N232, N227, N164);
and AND3 (N233, N225, N222, N17);
nand NAND3 (N234, N232, N86, N7);
or OR3 (N235, N228, N136, N68);
nand NAND3 (N236, N219, N46, N111);
buf BUF1 (N237, N226);
nor NOR4 (N238, N223, N131, N20, N71);
xor XOR2 (N239, N237, N123);
not NOT1 (N240, N239);
and AND2 (N241, N224, N104);
not NOT1 (N242, N238);
nand NAND2 (N243, N233, N115);
not NOT1 (N244, N236);
or OR4 (N245, N244, N69, N225, N167);
nor NOR3 (N246, N240, N129, N87);
buf BUF1 (N247, N231);
and AND4 (N248, N234, N119, N40, N70);
or OR2 (N249, N230, N161);
and AND4 (N250, N235, N119, N54, N151);
and AND3 (N251, N247, N173, N45);
xor XOR2 (N252, N205, N130);
nor NOR4 (N253, N246, N43, N68, N160);
buf BUF1 (N254, N243);
and AND3 (N255, N248, N133, N199);
and AND4 (N256, N245, N55, N23, N128);
xor XOR2 (N257, N252, N202);
xor XOR2 (N258, N249, N77);
or OR3 (N259, N258, N211, N188);
not NOT1 (N260, N259);
nor NOR3 (N261, N253, N234, N60);
xor XOR2 (N262, N254, N259);
and AND3 (N263, N256, N38, N92);
nor NOR3 (N264, N262, N80, N257);
xor XOR2 (N265, N54, N201);
nand NAND2 (N266, N250, N60);
or OR2 (N267, N241, N169);
xor XOR2 (N268, N264, N11);
not NOT1 (N269, N255);
xor XOR2 (N270, N251, N12);
buf BUF1 (N271, N260);
nor NOR3 (N272, N242, N228, N67);
and AND4 (N273, N269, N206, N216, N65);
and AND2 (N274, N266, N261);
xor XOR2 (N275, N219, N229);
nand NAND2 (N276, N263, N181);
nand NAND3 (N277, N273, N246, N174);
or OR4 (N278, N274, N144, N210, N24);
nand NAND4 (N279, N277, N177, N247, N10);
not NOT1 (N280, N267);
nand NAND4 (N281, N275, N144, N20, N24);
nor NOR4 (N282, N271, N54, N89, N191);
not NOT1 (N283, N272);
nand NAND2 (N284, N265, N53);
and AND3 (N285, N270, N14, N165);
xor XOR2 (N286, N283, N109);
not NOT1 (N287, N268);
nor NOR3 (N288, N276, N98, N133);
not NOT1 (N289, N285);
buf BUF1 (N290, N282);
or OR2 (N291, N279, N53);
and AND3 (N292, N288, N110, N86);
nor NOR2 (N293, N278, N33);
not NOT1 (N294, N291);
or OR4 (N295, N287, N258, N220, N172);
buf BUF1 (N296, N286);
nand NAND4 (N297, N294, N88, N129, N126);
nor NOR4 (N298, N297, N21, N178, N34);
buf BUF1 (N299, N284);
xor XOR2 (N300, N292, N83);
and AND2 (N301, N296, N61);
and AND3 (N302, N281, N146, N253);
nand NAND4 (N303, N301, N136, N25, N20);
or OR3 (N304, N295, N52, N248);
nand NAND2 (N305, N298, N210);
or OR2 (N306, N280, N218);
buf BUF1 (N307, N302);
or OR3 (N308, N303, N203, N41);
buf BUF1 (N309, N307);
nor NOR4 (N310, N309, N77, N88, N241);
xor XOR2 (N311, N305, N192);
nor NOR4 (N312, N293, N126, N311, N66);
not NOT1 (N313, N210);
nor NOR2 (N314, N299, N211);
nor NOR2 (N315, N306, N210);
xor XOR2 (N316, N290, N267);
xor XOR2 (N317, N300, N213);
nor NOR4 (N318, N308, N298, N191, N186);
not NOT1 (N319, N310);
and AND3 (N320, N317, N289, N90);
or OR2 (N321, N249, N304);
xor XOR2 (N322, N117, N306);
nand NAND3 (N323, N316, N146, N9);
or OR3 (N324, N318, N267, N106);
xor XOR2 (N325, N322, N99);
not NOT1 (N326, N319);
not NOT1 (N327, N324);
nor NOR4 (N328, N325, N157, N193, N25);
not NOT1 (N329, N326);
buf BUF1 (N330, N314);
or OR4 (N331, N330, N137, N113, N52);
nand NAND4 (N332, N327, N273, N6, N86);
xor XOR2 (N333, N312, N254);
nor NOR2 (N334, N320, N38);
buf BUF1 (N335, N321);
buf BUF1 (N336, N329);
or OR4 (N337, N315, N101, N21, N311);
nor NOR2 (N338, N334, N310);
or OR3 (N339, N332, N203, N147);
and AND2 (N340, N313, N277);
xor XOR2 (N341, N323, N152);
nand NAND2 (N342, N339, N327);
or OR2 (N343, N338, N45);
nor NOR3 (N344, N341, N76, N210);
nor NOR3 (N345, N331, N78, N3);
nand NAND2 (N346, N333, N78);
or OR4 (N347, N337, N335, N24, N117);
not NOT1 (N348, N20);
and AND3 (N349, N328, N1, N313);
xor XOR2 (N350, N342, N173);
not NOT1 (N351, N346);
and AND2 (N352, N348, N135);
nand NAND2 (N353, N349, N37);
nor NOR2 (N354, N347, N231);
or OR3 (N355, N343, N151, N158);
xor XOR2 (N356, N353, N46);
xor XOR2 (N357, N355, N269);
xor XOR2 (N358, N354, N92);
xor XOR2 (N359, N356, N110);
and AND3 (N360, N357, N336, N159);
buf BUF1 (N361, N76);
and AND4 (N362, N359, N148, N274, N333);
buf BUF1 (N363, N350);
nand NAND3 (N364, N340, N141, N28);
or OR3 (N365, N358, N8, N341);
nand NAND4 (N366, N344, N361, N18, N128);
nor NOR2 (N367, N186, N16);
nand NAND4 (N368, N351, N42, N124, N73);
nand NAND4 (N369, N365, N303, N128, N77);
nand NAND3 (N370, N366, N233, N204);
xor XOR2 (N371, N370, N208);
or OR4 (N372, N364, N187, N257, N205);
buf BUF1 (N373, N352);
nor NOR2 (N374, N362, N355);
or OR4 (N375, N345, N183, N370, N316);
not NOT1 (N376, N360);
not NOT1 (N377, N374);
xor XOR2 (N378, N368, N202);
nor NOR4 (N379, N369, N84, N23, N99);
xor XOR2 (N380, N375, N150);
or OR3 (N381, N380, N205, N63);
and AND2 (N382, N376, N42);
nor NOR3 (N383, N382, N366, N243);
xor XOR2 (N384, N378, N368);
nor NOR2 (N385, N372, N84);
xor XOR2 (N386, N363, N18);
or OR3 (N387, N373, N238, N11);
and AND4 (N388, N385, N337, N154, N317);
buf BUF1 (N389, N383);
not NOT1 (N390, N386);
or OR2 (N391, N381, N285);
xor XOR2 (N392, N377, N184);
not NOT1 (N393, N391);
not NOT1 (N394, N367);
and AND4 (N395, N389, N276, N88, N66);
buf BUF1 (N396, N384);
and AND2 (N397, N371, N382);
nand NAND3 (N398, N396, N57, N186);
xor XOR2 (N399, N395, N389);
nor NOR3 (N400, N394, N206, N159);
not NOT1 (N401, N397);
or OR2 (N402, N393, N17);
or OR2 (N403, N398, N44);
nand NAND2 (N404, N387, N227);
or OR4 (N405, N400, N252, N322, N93);
xor XOR2 (N406, N403, N132);
and AND3 (N407, N379, N244, N194);
xor XOR2 (N408, N399, N1);
or OR4 (N409, N392, N135, N233, N245);
and AND3 (N410, N388, N262, N61);
or OR3 (N411, N404, N271, N256);
buf BUF1 (N412, N407);
and AND3 (N413, N411, N4, N406);
not NOT1 (N414, N349);
buf BUF1 (N415, N412);
not NOT1 (N416, N405);
nand NAND2 (N417, N408, N145);
nor NOR4 (N418, N401, N284, N242, N311);
buf BUF1 (N419, N418);
or OR4 (N420, N414, N135, N120, N252);
buf BUF1 (N421, N390);
not NOT1 (N422, N416);
or OR3 (N423, N417, N174, N323);
nand NAND4 (N424, N422, N262, N403, N93);
or OR3 (N425, N421, N377, N337);
nand NAND4 (N426, N419, N139, N174, N66);
nor NOR3 (N427, N409, N360, N28);
xor XOR2 (N428, N413, N378);
or OR3 (N429, N410, N139, N249);
not NOT1 (N430, N428);
nor NOR4 (N431, N415, N28, N275, N236);
nand NAND3 (N432, N420, N374, N63);
not NOT1 (N433, N430);
and AND4 (N434, N425, N321, N287, N217);
xor XOR2 (N435, N432, N276);
and AND4 (N436, N429, N187, N42, N268);
xor XOR2 (N437, N431, N388);
buf BUF1 (N438, N402);
or OR2 (N439, N424, N44);
nor NOR2 (N440, N433, N168);
or OR3 (N441, N437, N249, N160);
buf BUF1 (N442, N436);
nand NAND4 (N443, N439, N96, N15, N382);
nor NOR2 (N444, N434, N414);
nor NOR2 (N445, N440, N301);
nor NOR3 (N446, N443, N182, N147);
nor NOR2 (N447, N446, N135);
nand NAND2 (N448, N444, N138);
and AND4 (N449, N448, N85, N304, N326);
nand NAND3 (N450, N426, N395, N381);
nor NOR4 (N451, N427, N388, N63, N309);
not NOT1 (N452, N423);
and AND2 (N453, N447, N177);
buf BUF1 (N454, N450);
nor NOR2 (N455, N449, N126);
nand NAND2 (N456, N442, N186);
and AND4 (N457, N454, N184, N50, N280);
nor NOR2 (N458, N457, N240);
and AND3 (N459, N452, N150, N439);
buf BUF1 (N460, N455);
nor NOR3 (N461, N458, N190, N70);
xor XOR2 (N462, N451, N49);
buf BUF1 (N463, N438);
not NOT1 (N464, N462);
xor XOR2 (N465, N445, N19);
or OR2 (N466, N456, N206);
xor XOR2 (N467, N453, N384);
not NOT1 (N468, N460);
or OR2 (N469, N461, N389);
xor XOR2 (N470, N435, N103);
nand NAND4 (N471, N464, N362, N158, N336);
and AND4 (N472, N466, N123, N266, N315);
xor XOR2 (N473, N470, N267);
nand NAND2 (N474, N468, N72);
xor XOR2 (N475, N463, N204);
nand NAND4 (N476, N441, N81, N267, N217);
not NOT1 (N477, N475);
not NOT1 (N478, N465);
nor NOR2 (N479, N478, N238);
nand NAND2 (N480, N467, N92);
and AND2 (N481, N472, N448);
and AND2 (N482, N477, N333);
not NOT1 (N483, N476);
xor XOR2 (N484, N479, N70);
buf BUF1 (N485, N481);
nand NAND2 (N486, N471, N329);
or OR3 (N487, N485, N82, N91);
and AND3 (N488, N459, N338, N454);
buf BUF1 (N489, N484);
nor NOR2 (N490, N487, N243);
or OR4 (N491, N474, N34, N223, N236);
not NOT1 (N492, N482);
nor NOR2 (N493, N490, N335);
or OR4 (N494, N493, N410, N115, N198);
xor XOR2 (N495, N488, N51);
nand NAND4 (N496, N483, N37, N272, N274);
not NOT1 (N497, N480);
or OR3 (N498, N469, N106, N3);
nand NAND2 (N499, N491, N428);
nor NOR2 (N500, N499, N99);
buf BUF1 (N501, N495);
or OR3 (N502, N501, N191, N486);
xor XOR2 (N503, N154, N241);
or OR4 (N504, N503, N449, N20, N430);
buf BUF1 (N505, N502);
or OR2 (N506, N498, N288);
or OR2 (N507, N473, N50);
nor NOR3 (N508, N494, N83, N357);
and AND3 (N509, N504, N189, N97);
and AND2 (N510, N505, N353);
xor XOR2 (N511, N496, N479);
not NOT1 (N512, N508);
nor NOR2 (N513, N497, N323);
endmodule