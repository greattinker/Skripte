// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12;

output N8005,N8004,N7999,N8008,N8011,N8006,N7994,N8010,N7996,N8012;

nor NOR4 (N13, N6, N2, N10, N12);
and AND4 (N14, N5, N5, N8, N5);
nor NOR2 (N15, N2, N5);
and AND2 (N16, N9, N5);
buf BUF1 (N17, N11);
xor XOR2 (N18, N13, N17);
buf BUF1 (N19, N17);
buf BUF1 (N20, N1);
xor XOR2 (N21, N8, N15);
and AND4 (N22, N16, N2, N11, N8);
nand NAND3 (N23, N22, N6, N12);
nand NAND2 (N24, N16, N3);
not NOT1 (N25, N22);
nand NAND3 (N26, N15, N12, N25);
not NOT1 (N27, N15);
buf BUF1 (N28, N10);
nor NOR3 (N29, N28, N8, N17);
xor XOR2 (N30, N14, N10);
nand NAND2 (N31, N27, N24);
or OR4 (N32, N10, N1, N19, N18);
not NOT1 (N33, N3);
not NOT1 (N34, N33);
or OR4 (N35, N31, N27, N6, N3);
or OR2 (N36, N9, N9);
xor XOR2 (N37, N21, N22);
buf BUF1 (N38, N32);
not NOT1 (N39, N35);
buf BUF1 (N40, N20);
not NOT1 (N41, N36);
not NOT1 (N42, N39);
nand NAND2 (N43, N41, N2);
nand NAND2 (N44, N43, N13);
nor NOR4 (N45, N30, N34, N37, N42);
and AND2 (N46, N3, N15);
nor NOR2 (N47, N5, N37);
or OR2 (N48, N18, N19);
xor XOR2 (N49, N23, N9);
nor NOR3 (N50, N45, N28, N6);
not NOT1 (N51, N40);
not NOT1 (N52, N46);
nand NAND2 (N53, N50, N23);
buf BUF1 (N54, N29);
and AND4 (N55, N38, N10, N37, N2);
buf BUF1 (N56, N49);
buf BUF1 (N57, N44);
not NOT1 (N58, N57);
nand NAND2 (N59, N56, N56);
nand NAND2 (N60, N52, N22);
xor XOR2 (N61, N59, N34);
or OR2 (N62, N58, N12);
and AND4 (N63, N51, N29, N13, N12);
not NOT1 (N64, N53);
and AND2 (N65, N60, N30);
or OR4 (N66, N26, N4, N34, N3);
nand NAND4 (N67, N64, N10, N33, N58);
xor XOR2 (N68, N63, N30);
and AND4 (N69, N54, N65, N15, N22);
or OR3 (N70, N20, N26, N21);
not NOT1 (N71, N61);
or OR2 (N72, N70, N52);
not NOT1 (N73, N48);
not NOT1 (N74, N73);
or OR3 (N75, N71, N6, N32);
and AND3 (N76, N55, N51, N38);
and AND2 (N77, N68, N64);
nor NOR3 (N78, N75, N52, N26);
not NOT1 (N79, N72);
nor NOR2 (N80, N69, N51);
or OR4 (N81, N67, N74, N5, N8);
not NOT1 (N82, N29);
nor NOR2 (N83, N76, N77);
or OR2 (N84, N29, N59);
and AND3 (N85, N47, N60, N58);
nand NAND3 (N86, N79, N73, N83);
nor NOR2 (N87, N32, N40);
buf BUF1 (N88, N85);
nor NOR4 (N89, N88, N64, N55, N22);
nor NOR2 (N90, N84, N11);
nor NOR4 (N91, N82, N19, N38, N30);
not NOT1 (N92, N81);
nand NAND4 (N93, N86, N15, N84, N6);
not NOT1 (N94, N92);
or OR4 (N95, N87, N5, N8, N62);
not NOT1 (N96, N17);
xor XOR2 (N97, N80, N40);
nand NAND3 (N98, N95, N34, N10);
buf BUF1 (N99, N93);
nor NOR2 (N100, N94, N1);
not NOT1 (N101, N97);
not NOT1 (N102, N98);
not NOT1 (N103, N100);
buf BUF1 (N104, N96);
nand NAND2 (N105, N101, N46);
or OR2 (N106, N89, N23);
xor XOR2 (N107, N106, N43);
not NOT1 (N108, N102);
xor XOR2 (N109, N105, N15);
nand NAND4 (N110, N109, N65, N87, N79);
buf BUF1 (N111, N78);
not NOT1 (N112, N104);
xor XOR2 (N113, N108, N1);
or OR3 (N114, N90, N76, N13);
and AND2 (N115, N66, N78);
buf BUF1 (N116, N114);
xor XOR2 (N117, N110, N30);
and AND3 (N118, N113, N114, N112);
or OR2 (N119, N19, N62);
nand NAND4 (N120, N118, N37, N94, N96);
buf BUF1 (N121, N107);
nor NOR4 (N122, N116, N47, N79, N48);
and AND4 (N123, N117, N3, N21, N56);
and AND3 (N124, N103, N1, N73);
nor NOR4 (N125, N115, N124, N28, N105);
nand NAND3 (N126, N46, N12, N71);
not NOT1 (N127, N125);
buf BUF1 (N128, N99);
not NOT1 (N129, N128);
and AND3 (N130, N126, N92, N91);
and AND2 (N131, N26, N13);
and AND2 (N132, N130, N104);
not NOT1 (N133, N127);
and AND2 (N134, N133, N4);
and AND4 (N135, N134, N109, N109, N81);
nor NOR4 (N136, N121, N128, N10, N106);
nor NOR4 (N137, N135, N104, N97, N49);
nor NOR4 (N138, N131, N131, N106, N61);
xor XOR2 (N139, N129, N14);
buf BUF1 (N140, N111);
nor NOR3 (N141, N119, N77, N16);
nor NOR3 (N142, N141, N118, N78);
nand NAND3 (N143, N123, N78, N58);
xor XOR2 (N144, N140, N104);
nor NOR4 (N145, N138, N135, N34, N5);
nor NOR2 (N146, N132, N104);
nor NOR4 (N147, N142, N4, N24, N135);
or OR3 (N148, N143, N44, N146);
nand NAND4 (N149, N42, N100, N110, N123);
nand NAND4 (N150, N122, N2, N7, N68);
not NOT1 (N151, N120);
buf BUF1 (N152, N148);
and AND3 (N153, N136, N91, N110);
nand NAND3 (N154, N144, N12, N64);
buf BUF1 (N155, N145);
and AND4 (N156, N151, N126, N106, N93);
or OR2 (N157, N155, N119);
nor NOR4 (N158, N157, N53, N26, N109);
buf BUF1 (N159, N153);
and AND4 (N160, N150, N73, N145, N123);
and AND2 (N161, N159, N53);
xor XOR2 (N162, N161, N92);
nand NAND4 (N163, N156, N55, N134, N67);
nand NAND3 (N164, N163, N19, N1);
nand NAND2 (N165, N149, N90);
nor NOR4 (N166, N147, N57, N20, N150);
nor NOR3 (N167, N152, N36, N61);
buf BUF1 (N168, N154);
not NOT1 (N169, N164);
nor NOR3 (N170, N162, N25, N73);
not NOT1 (N171, N170);
not NOT1 (N172, N139);
and AND3 (N173, N160, N123, N143);
buf BUF1 (N174, N166);
xor XOR2 (N175, N169, N172);
or OR4 (N176, N28, N149, N11, N98);
or OR2 (N177, N137, N74);
and AND2 (N178, N176, N147);
nand NAND3 (N179, N173, N14, N58);
not NOT1 (N180, N174);
nor NOR4 (N181, N167, N76, N66, N63);
not NOT1 (N182, N165);
or OR4 (N183, N158, N129, N131, N80);
xor XOR2 (N184, N178, N107);
xor XOR2 (N185, N183, N171);
or OR3 (N186, N28, N41, N121);
nor NOR2 (N187, N179, N35);
or OR4 (N188, N181, N71, N70, N137);
nor NOR3 (N189, N186, N5, N71);
buf BUF1 (N190, N180);
and AND2 (N191, N187, N60);
nand NAND2 (N192, N190, N150);
xor XOR2 (N193, N182, N82);
buf BUF1 (N194, N192);
xor XOR2 (N195, N177, N133);
and AND2 (N196, N168, N37);
and AND4 (N197, N191, N65, N82, N191);
nand NAND4 (N198, N193, N98, N102, N146);
nand NAND3 (N199, N189, N8, N165);
xor XOR2 (N200, N196, N122);
xor XOR2 (N201, N185, N105);
or OR3 (N202, N201, N175, N131);
nand NAND2 (N203, N180, N191);
not NOT1 (N204, N184);
not NOT1 (N205, N195);
not NOT1 (N206, N188);
or OR2 (N207, N203, N134);
xor XOR2 (N208, N205, N33);
nor NOR2 (N209, N199, N51);
buf BUF1 (N210, N200);
nor NOR2 (N211, N210, N204);
not NOT1 (N212, N61);
nor NOR3 (N213, N202, N160, N89);
xor XOR2 (N214, N208, N58);
not NOT1 (N215, N206);
buf BUF1 (N216, N215);
or OR3 (N217, N213, N46, N166);
buf BUF1 (N218, N194);
or OR3 (N219, N217, N119, N149);
xor XOR2 (N220, N216, N118);
nand NAND4 (N221, N197, N71, N196, N31);
not NOT1 (N222, N198);
buf BUF1 (N223, N219);
and AND3 (N224, N212, N80, N14);
xor XOR2 (N225, N207, N93);
and AND4 (N226, N214, N128, N185, N119);
or OR4 (N227, N223, N168, N185, N134);
buf BUF1 (N228, N225);
nor NOR2 (N229, N209, N129);
buf BUF1 (N230, N222);
xor XOR2 (N231, N218, N133);
buf BUF1 (N232, N231);
buf BUF1 (N233, N224);
or OR2 (N234, N233, N179);
not NOT1 (N235, N221);
buf BUF1 (N236, N234);
nand NAND3 (N237, N227, N76, N39);
nand NAND4 (N238, N236, N85, N214, N64);
buf BUF1 (N239, N232);
buf BUF1 (N240, N238);
xor XOR2 (N241, N235, N2);
nor NOR3 (N242, N229, N222, N91);
not NOT1 (N243, N242);
and AND2 (N244, N230, N109);
not NOT1 (N245, N211);
xor XOR2 (N246, N240, N211);
not NOT1 (N247, N226);
xor XOR2 (N248, N237, N178);
nor NOR4 (N249, N248, N114, N201, N151);
buf BUF1 (N250, N247);
and AND3 (N251, N243, N54, N95);
not NOT1 (N252, N228);
nand NAND4 (N253, N244, N95, N207, N62);
or OR2 (N254, N245, N244);
or OR4 (N255, N246, N142, N200, N151);
buf BUF1 (N256, N241);
or OR4 (N257, N250, N86, N148, N116);
buf BUF1 (N258, N251);
not NOT1 (N259, N220);
and AND4 (N260, N255, N7, N254, N83);
nand NAND2 (N261, N78, N66);
buf BUF1 (N262, N256);
and AND4 (N263, N261, N160, N211, N253);
or OR3 (N264, N262, N198, N184);
xor XOR2 (N265, N147, N220);
nand NAND3 (N266, N249, N3, N31);
buf BUF1 (N267, N258);
buf BUF1 (N268, N266);
nor NOR3 (N269, N257, N15, N208);
not NOT1 (N270, N259);
xor XOR2 (N271, N239, N260);
buf BUF1 (N272, N188);
nand NAND2 (N273, N270, N138);
and AND4 (N274, N252, N89, N178, N135);
xor XOR2 (N275, N265, N206);
buf BUF1 (N276, N269);
nor NOR3 (N277, N275, N2, N193);
not NOT1 (N278, N272);
not NOT1 (N279, N274);
buf BUF1 (N280, N273);
not NOT1 (N281, N276);
or OR3 (N282, N280, N212, N74);
buf BUF1 (N283, N268);
nand NAND2 (N284, N263, N74);
nor NOR3 (N285, N264, N59, N52);
or OR3 (N286, N277, N241, N110);
nor NOR2 (N287, N286, N71);
and AND2 (N288, N279, N193);
or OR4 (N289, N283, N86, N265, N58);
and AND4 (N290, N287, N272, N36, N156);
or OR2 (N291, N288, N52);
not NOT1 (N292, N290);
xor XOR2 (N293, N282, N22);
nor NOR4 (N294, N267, N85, N160, N209);
nand NAND4 (N295, N281, N247, N196, N45);
not NOT1 (N296, N293);
not NOT1 (N297, N294);
nand NAND3 (N298, N292, N186, N192);
nor NOR2 (N299, N284, N96);
not NOT1 (N300, N291);
not NOT1 (N301, N298);
nor NOR4 (N302, N295, N164, N209, N290);
not NOT1 (N303, N271);
nor NOR2 (N304, N285, N34);
and AND2 (N305, N278, N277);
xor XOR2 (N306, N296, N176);
nand NAND3 (N307, N303, N195, N108);
not NOT1 (N308, N307);
nand NAND2 (N309, N304, N81);
not NOT1 (N310, N297);
nand NAND3 (N311, N308, N37, N161);
and AND4 (N312, N305, N265, N135, N196);
or OR2 (N313, N289, N113);
xor XOR2 (N314, N311, N259);
or OR2 (N315, N306, N272);
buf BUF1 (N316, N310);
xor XOR2 (N317, N299, N35);
xor XOR2 (N318, N313, N226);
nor NOR2 (N319, N300, N152);
and AND4 (N320, N314, N61, N268, N31);
or OR4 (N321, N319, N50, N97, N76);
and AND2 (N322, N316, N36);
or OR2 (N323, N321, N96);
or OR2 (N324, N318, N89);
nand NAND2 (N325, N315, N159);
not NOT1 (N326, N317);
nor NOR3 (N327, N326, N305, N221);
not NOT1 (N328, N301);
not NOT1 (N329, N322);
or OR3 (N330, N325, N258, N273);
not NOT1 (N331, N327);
buf BUF1 (N332, N320);
xor XOR2 (N333, N312, N217);
not NOT1 (N334, N331);
buf BUF1 (N335, N329);
not NOT1 (N336, N330);
or OR4 (N337, N302, N209, N1, N271);
nor NOR4 (N338, N334, N17, N264, N10);
buf BUF1 (N339, N309);
xor XOR2 (N340, N336, N74);
not NOT1 (N341, N332);
and AND4 (N342, N333, N220, N235, N14);
nor NOR4 (N343, N335, N124, N217, N233);
nand NAND4 (N344, N324, N135, N314, N269);
nor NOR4 (N345, N337, N277, N337, N18);
not NOT1 (N346, N340);
and AND3 (N347, N342, N11, N339);
not NOT1 (N348, N56);
or OR2 (N349, N346, N83);
or OR2 (N350, N349, N23);
and AND4 (N351, N350, N238, N158, N12);
nor NOR2 (N352, N351, N299);
or OR3 (N353, N341, N43, N131);
buf BUF1 (N354, N347);
buf BUF1 (N355, N348);
not NOT1 (N356, N343);
xor XOR2 (N357, N344, N323);
not NOT1 (N358, N81);
buf BUF1 (N359, N328);
and AND3 (N360, N354, N235, N235);
nor NOR4 (N361, N358, N192, N248, N309);
or OR4 (N362, N355, N263, N57, N124);
nand NAND2 (N363, N338, N190);
not NOT1 (N364, N362);
nand NAND2 (N365, N360, N53);
xor XOR2 (N366, N363, N57);
nand NAND4 (N367, N364, N354, N67, N30);
xor XOR2 (N368, N357, N192);
xor XOR2 (N369, N368, N245);
not NOT1 (N370, N366);
nand NAND4 (N371, N370, N300, N177, N118);
not NOT1 (N372, N352);
buf BUF1 (N373, N361);
buf BUF1 (N374, N373);
buf BUF1 (N375, N353);
nand NAND4 (N376, N371, N353, N317, N9);
xor XOR2 (N377, N372, N306);
buf BUF1 (N378, N345);
and AND3 (N379, N359, N25, N20);
nor NOR3 (N380, N375, N116, N85);
xor XOR2 (N381, N356, N88);
xor XOR2 (N382, N374, N19);
and AND2 (N383, N382, N232);
not NOT1 (N384, N378);
nor NOR2 (N385, N369, N224);
or OR2 (N386, N381, N71);
nand NAND4 (N387, N367, N258, N346, N12);
or OR4 (N388, N379, N316, N67, N374);
nor NOR2 (N389, N383, N312);
or OR4 (N390, N377, N220, N300, N11);
or OR4 (N391, N389, N121, N390, N26);
nor NOR2 (N392, N101, N378);
xor XOR2 (N393, N391, N201);
xor XOR2 (N394, N386, N20);
not NOT1 (N395, N376);
or OR2 (N396, N385, N290);
or OR2 (N397, N365, N30);
xor XOR2 (N398, N395, N114);
nand NAND2 (N399, N380, N167);
and AND3 (N400, N392, N398, N336);
nor NOR4 (N401, N284, N267, N30, N148);
nor NOR2 (N402, N396, N49);
not NOT1 (N403, N388);
nor NOR4 (N404, N387, N337, N87, N119);
xor XOR2 (N405, N384, N204);
nand NAND3 (N406, N404, N263, N26);
nand NAND2 (N407, N399, N14);
nand NAND3 (N408, N393, N329, N199);
nor NOR3 (N409, N403, N31, N243);
xor XOR2 (N410, N406, N37);
nand NAND4 (N411, N394, N117, N121, N302);
buf BUF1 (N412, N409);
and AND2 (N413, N408, N368);
and AND4 (N414, N405, N36, N240, N355);
or OR3 (N415, N413, N82, N226);
not NOT1 (N416, N397);
xor XOR2 (N417, N407, N155);
not NOT1 (N418, N410);
not NOT1 (N419, N411);
and AND4 (N420, N418, N321, N355, N297);
or OR4 (N421, N400, N243, N314, N192);
nor NOR4 (N422, N414, N66, N347, N244);
nand NAND3 (N423, N417, N98, N340);
xor XOR2 (N424, N421, N22);
and AND4 (N425, N423, N389, N143, N164);
nor NOR3 (N426, N425, N139, N280);
nor NOR3 (N427, N424, N273, N426);
or OR2 (N428, N377, N140);
nand NAND4 (N429, N422, N89, N173, N381);
nor NOR3 (N430, N419, N378, N32);
or OR4 (N431, N401, N347, N374, N243);
nand NAND2 (N432, N428, N108);
or OR2 (N433, N429, N249);
nand NAND4 (N434, N433, N84, N93, N391);
and AND3 (N435, N427, N42, N417);
xor XOR2 (N436, N402, N161);
buf BUF1 (N437, N420);
and AND3 (N438, N416, N435, N85);
and AND4 (N439, N163, N17, N376, N111);
nand NAND2 (N440, N412, N188);
buf BUF1 (N441, N431);
not NOT1 (N442, N432);
not NOT1 (N443, N440);
buf BUF1 (N444, N415);
and AND4 (N445, N439, N90, N186, N172);
or OR2 (N446, N436, N325);
nor NOR3 (N447, N434, N159, N68);
nand NAND4 (N448, N442, N362, N225, N162);
or OR2 (N449, N441, N257);
not NOT1 (N450, N437);
or OR2 (N451, N438, N362);
nand NAND3 (N452, N446, N267, N441);
or OR4 (N453, N447, N130, N27, N333);
and AND3 (N454, N448, N405, N322);
xor XOR2 (N455, N443, N194);
or OR2 (N456, N449, N98);
not NOT1 (N457, N450);
buf BUF1 (N458, N457);
buf BUF1 (N459, N430);
nor NOR3 (N460, N444, N56, N360);
or OR4 (N461, N455, N147, N299, N174);
nand NAND3 (N462, N445, N451, N385);
or OR4 (N463, N353, N45, N62, N137);
buf BUF1 (N464, N456);
nor NOR4 (N465, N461, N71, N255, N192);
and AND3 (N466, N454, N443, N279);
nor NOR3 (N467, N463, N380, N65);
or OR3 (N468, N462, N442, N355);
nand NAND4 (N469, N467, N323, N117, N315);
not NOT1 (N470, N453);
buf BUF1 (N471, N459);
nand NAND2 (N472, N464, N70);
or OR3 (N473, N471, N346, N13);
nand NAND2 (N474, N472, N121);
nand NAND3 (N475, N458, N427, N323);
nor NOR3 (N476, N469, N199, N384);
buf BUF1 (N477, N452);
and AND4 (N478, N476, N326, N286, N403);
nor NOR3 (N479, N460, N111, N415);
buf BUF1 (N480, N466);
nor NOR3 (N481, N475, N373, N326);
buf BUF1 (N482, N477);
or OR4 (N483, N465, N379, N446, N404);
buf BUF1 (N484, N478);
nor NOR3 (N485, N481, N145, N351);
or OR2 (N486, N474, N286);
xor XOR2 (N487, N468, N319);
nor NOR3 (N488, N470, N176, N160);
nor NOR4 (N489, N488, N87, N427, N284);
nand NAND2 (N490, N489, N250);
or OR4 (N491, N479, N183, N388, N148);
nand NAND4 (N492, N490, N227, N137, N1);
not NOT1 (N493, N483);
nor NOR3 (N494, N492, N366, N486);
nor NOR2 (N495, N320, N220);
xor XOR2 (N496, N495, N206);
buf BUF1 (N497, N487);
and AND3 (N498, N480, N39, N314);
and AND3 (N499, N494, N206, N379);
xor XOR2 (N500, N484, N34);
nand NAND4 (N501, N485, N181, N465, N201);
not NOT1 (N502, N500);
xor XOR2 (N503, N482, N500);
or OR3 (N504, N501, N93, N151);
nand NAND2 (N505, N503, N15);
or OR2 (N506, N502, N203);
nor NOR4 (N507, N497, N273, N427, N106);
buf BUF1 (N508, N499);
and AND4 (N509, N491, N399, N222, N9);
or OR2 (N510, N498, N11);
buf BUF1 (N511, N504);
and AND4 (N512, N496, N217, N412, N190);
buf BUF1 (N513, N507);
and AND2 (N514, N508, N45);
or OR3 (N515, N506, N260, N431);
buf BUF1 (N516, N505);
nand NAND3 (N517, N509, N446, N339);
not NOT1 (N518, N516);
nor NOR2 (N519, N517, N512);
and AND4 (N520, N198, N224, N456, N472);
or OR2 (N521, N514, N188);
xor XOR2 (N522, N515, N453);
xor XOR2 (N523, N518, N21);
not NOT1 (N524, N473);
buf BUF1 (N525, N522);
nand NAND2 (N526, N510, N291);
not NOT1 (N527, N519);
and AND3 (N528, N493, N486, N335);
and AND4 (N529, N525, N483, N299, N493);
buf BUF1 (N530, N523);
and AND4 (N531, N511, N208, N214, N320);
xor XOR2 (N532, N524, N187);
nor NOR3 (N533, N526, N498, N222);
and AND4 (N534, N530, N129, N339, N68);
and AND3 (N535, N521, N302, N383);
nor NOR4 (N536, N527, N374, N405, N88);
and AND3 (N537, N536, N411, N420);
or OR2 (N538, N528, N144);
and AND4 (N539, N533, N158, N402, N148);
xor XOR2 (N540, N534, N195);
or OR4 (N541, N538, N326, N232, N399);
and AND4 (N542, N541, N414, N494, N24);
not NOT1 (N543, N539);
or OR2 (N544, N513, N327);
or OR3 (N545, N531, N456, N216);
nor NOR2 (N546, N545, N542);
not NOT1 (N547, N333);
xor XOR2 (N548, N546, N148);
buf BUF1 (N549, N547);
nor NOR2 (N550, N520, N112);
and AND3 (N551, N529, N445, N509);
nor NOR3 (N552, N551, N445, N86);
nand NAND3 (N553, N549, N282, N17);
not NOT1 (N554, N535);
or OR2 (N555, N552, N397);
not NOT1 (N556, N543);
nand NAND3 (N557, N532, N341, N220);
nand NAND2 (N558, N554, N150);
nor NOR4 (N559, N548, N210, N37, N399);
or OR4 (N560, N553, N520, N467, N559);
and AND4 (N561, N34, N319, N151, N442);
and AND4 (N562, N561, N242, N486, N34);
xor XOR2 (N563, N556, N185);
and AND3 (N564, N550, N126, N463);
nor NOR4 (N565, N540, N79, N210, N532);
or OR3 (N566, N562, N541, N468);
and AND2 (N567, N564, N51);
not NOT1 (N568, N560);
and AND3 (N569, N567, N82, N333);
nand NAND3 (N570, N565, N433, N466);
not NOT1 (N571, N557);
or OR3 (N572, N558, N349, N504);
nand NAND4 (N573, N537, N323, N74, N113);
and AND3 (N574, N570, N327, N155);
xor XOR2 (N575, N571, N369);
not NOT1 (N576, N555);
nor NOR3 (N577, N572, N92, N295);
or OR3 (N578, N575, N539, N406);
and AND3 (N579, N578, N498, N256);
and AND3 (N580, N568, N343, N6);
or OR2 (N581, N573, N301);
and AND4 (N582, N576, N219, N30, N441);
and AND3 (N583, N574, N238, N451);
xor XOR2 (N584, N582, N408);
and AND4 (N585, N579, N412, N74, N465);
or OR3 (N586, N580, N531, N52);
buf BUF1 (N587, N563);
nand NAND4 (N588, N586, N528, N219, N137);
buf BUF1 (N589, N544);
nor NOR2 (N590, N587, N190);
buf BUF1 (N591, N585);
nor NOR4 (N592, N577, N278, N176, N544);
buf BUF1 (N593, N590);
buf BUF1 (N594, N592);
nand NAND3 (N595, N594, N482, N368);
buf BUF1 (N596, N593);
not NOT1 (N597, N595);
xor XOR2 (N598, N584, N496);
xor XOR2 (N599, N583, N335);
not NOT1 (N600, N591);
nor NOR2 (N601, N566, N563);
and AND4 (N602, N589, N257, N126, N533);
nor NOR2 (N603, N599, N332);
and AND3 (N604, N597, N134, N129);
buf BUF1 (N605, N569);
and AND2 (N606, N581, N454);
buf BUF1 (N607, N605);
and AND2 (N608, N598, N261);
not NOT1 (N609, N608);
or OR2 (N610, N607, N87);
xor XOR2 (N611, N609, N397);
nor NOR3 (N612, N603, N410, N65);
or OR2 (N613, N601, N326);
not NOT1 (N614, N610);
nand NAND4 (N615, N613, N85, N193, N366);
nor NOR3 (N616, N604, N422, N232);
not NOT1 (N617, N596);
nor NOR2 (N618, N588, N67);
and AND2 (N619, N615, N42);
not NOT1 (N620, N617);
and AND4 (N621, N612, N374, N520, N152);
nor NOR4 (N622, N611, N150, N201, N478);
nand NAND3 (N623, N620, N323, N549);
xor XOR2 (N624, N621, N134);
or OR2 (N625, N616, N171);
buf BUF1 (N626, N625);
or OR4 (N627, N602, N378, N218, N367);
nor NOR3 (N628, N626, N625, N396);
xor XOR2 (N629, N614, N258);
nor NOR3 (N630, N627, N144, N237);
nor NOR4 (N631, N618, N399, N182, N487);
nor NOR3 (N632, N629, N521, N29);
nand NAND4 (N633, N622, N504, N513, N572);
buf BUF1 (N634, N628);
and AND4 (N635, N631, N608, N218, N243);
not NOT1 (N636, N630);
nand NAND3 (N637, N619, N215, N328);
or OR2 (N638, N624, N80);
and AND2 (N639, N623, N564);
nand NAND2 (N640, N637, N91);
or OR4 (N641, N639, N321, N506, N532);
not NOT1 (N642, N633);
nor NOR4 (N643, N600, N342, N291, N520);
buf BUF1 (N644, N634);
xor XOR2 (N645, N641, N256);
nand NAND2 (N646, N644, N244);
or OR2 (N647, N643, N426);
not NOT1 (N648, N645);
buf BUF1 (N649, N642);
and AND3 (N650, N636, N559, N264);
xor XOR2 (N651, N638, N468);
nor NOR2 (N652, N648, N488);
nor NOR4 (N653, N651, N362, N295, N342);
xor XOR2 (N654, N635, N207);
nand NAND3 (N655, N653, N151, N196);
nor NOR4 (N656, N654, N640, N29, N280);
nand NAND4 (N657, N71, N607, N78, N580);
not NOT1 (N658, N650);
not NOT1 (N659, N655);
not NOT1 (N660, N657);
xor XOR2 (N661, N659, N618);
not NOT1 (N662, N647);
not NOT1 (N663, N656);
buf BUF1 (N664, N646);
and AND4 (N665, N661, N462, N471, N420);
nor NOR4 (N666, N606, N238, N308, N218);
not NOT1 (N667, N658);
xor XOR2 (N668, N663, N419);
xor XOR2 (N669, N649, N388);
buf BUF1 (N670, N667);
nor NOR2 (N671, N665, N276);
nand NAND4 (N672, N664, N11, N81, N262);
or OR2 (N673, N666, N137);
buf BUF1 (N674, N662);
buf BUF1 (N675, N669);
and AND3 (N676, N671, N591, N119);
buf BUF1 (N677, N668);
not NOT1 (N678, N673);
or OR4 (N679, N674, N336, N214, N209);
not NOT1 (N680, N632);
nand NAND2 (N681, N677, N248);
xor XOR2 (N682, N681, N197);
nand NAND4 (N683, N682, N297, N315, N266);
nor NOR3 (N684, N652, N639, N566);
buf BUF1 (N685, N678);
nor NOR3 (N686, N683, N38, N458);
or OR3 (N687, N660, N99, N461);
nor NOR3 (N688, N680, N617, N257);
nor NOR3 (N689, N675, N263, N656);
or OR4 (N690, N686, N629, N177, N447);
buf BUF1 (N691, N688);
nor NOR3 (N692, N676, N182, N93);
and AND3 (N693, N670, N266, N90);
buf BUF1 (N694, N679);
nand NAND3 (N695, N692, N524, N214);
or OR2 (N696, N672, N133);
not NOT1 (N697, N693);
and AND2 (N698, N685, N335);
and AND3 (N699, N687, N13, N676);
xor XOR2 (N700, N696, N532);
nor NOR2 (N701, N699, N539);
nor NOR3 (N702, N700, N324, N434);
buf BUF1 (N703, N697);
xor XOR2 (N704, N690, N90);
or OR2 (N705, N684, N270);
nor NOR3 (N706, N705, N374, N202);
xor XOR2 (N707, N689, N292);
buf BUF1 (N708, N706);
xor XOR2 (N709, N702, N236);
buf BUF1 (N710, N708);
nor NOR3 (N711, N694, N217, N239);
not NOT1 (N712, N710);
buf BUF1 (N713, N703);
not NOT1 (N714, N695);
and AND4 (N715, N704, N657, N513, N607);
nand NAND3 (N716, N713, N353, N708);
or OR4 (N717, N711, N182, N555, N461);
or OR3 (N718, N691, N591, N345);
and AND2 (N719, N707, N439);
nand NAND4 (N720, N717, N271, N401, N99);
or OR3 (N721, N716, N472, N473);
or OR4 (N722, N698, N410, N146, N362);
or OR2 (N723, N722, N325);
or OR2 (N724, N721, N500);
nor NOR4 (N725, N714, N487, N377, N204);
or OR2 (N726, N701, N81);
nor NOR4 (N727, N709, N47, N427, N242);
buf BUF1 (N728, N719);
xor XOR2 (N729, N720, N22);
and AND4 (N730, N712, N234, N447, N368);
or OR4 (N731, N715, N191, N694, N610);
nor NOR2 (N732, N728, N469);
xor XOR2 (N733, N724, N692);
and AND4 (N734, N718, N108, N271, N346);
and AND3 (N735, N734, N273, N473);
not NOT1 (N736, N733);
nor NOR3 (N737, N736, N444, N13);
or OR4 (N738, N732, N436, N147, N335);
nand NAND2 (N739, N723, N612);
nand NAND4 (N740, N731, N434, N9, N485);
and AND2 (N741, N739, N165);
buf BUF1 (N742, N740);
buf BUF1 (N743, N729);
nand NAND4 (N744, N735, N199, N251, N617);
nand NAND3 (N745, N744, N113, N15);
buf BUF1 (N746, N742);
and AND4 (N747, N737, N221, N331, N265);
and AND2 (N748, N747, N235);
nand NAND3 (N749, N738, N217, N127);
nand NAND3 (N750, N743, N522, N653);
and AND2 (N751, N745, N592);
buf BUF1 (N752, N730);
and AND2 (N753, N726, N539);
nor NOR2 (N754, N749, N203);
nand NAND4 (N755, N741, N626, N525, N216);
nand NAND4 (N756, N755, N350, N30, N87);
buf BUF1 (N757, N727);
buf BUF1 (N758, N757);
or OR2 (N759, N751, N682);
not NOT1 (N760, N746);
and AND3 (N761, N750, N129, N35);
and AND3 (N762, N759, N175, N544);
xor XOR2 (N763, N758, N611);
or OR2 (N764, N761, N610);
not NOT1 (N765, N764);
buf BUF1 (N766, N756);
xor XOR2 (N767, N748, N145);
xor XOR2 (N768, N765, N748);
and AND4 (N769, N754, N421, N33, N275);
not NOT1 (N770, N769);
or OR2 (N771, N760, N651);
nor NOR3 (N772, N767, N162, N613);
nor NOR3 (N773, N753, N637, N716);
and AND4 (N774, N763, N679, N244, N437);
buf BUF1 (N775, N752);
nor NOR4 (N776, N768, N653, N765, N492);
or OR3 (N777, N771, N454, N198);
or OR2 (N778, N762, N194);
buf BUF1 (N779, N778);
nor NOR4 (N780, N773, N775, N401, N778);
or OR2 (N781, N335, N605);
and AND2 (N782, N779, N193);
nor NOR2 (N783, N774, N321);
nor NOR2 (N784, N777, N138);
xor XOR2 (N785, N725, N654);
or OR3 (N786, N782, N663, N730);
nand NAND3 (N787, N772, N16, N47);
not NOT1 (N788, N785);
xor XOR2 (N789, N770, N343);
not NOT1 (N790, N786);
buf BUF1 (N791, N784);
xor XOR2 (N792, N787, N338);
buf BUF1 (N793, N792);
buf BUF1 (N794, N793);
nand NAND4 (N795, N766, N109, N527, N688);
buf BUF1 (N796, N791);
or OR4 (N797, N795, N631, N93, N745);
and AND3 (N798, N790, N221, N134);
buf BUF1 (N799, N783);
not NOT1 (N800, N794);
not NOT1 (N801, N780);
buf BUF1 (N802, N788);
buf BUF1 (N803, N796);
nor NOR4 (N804, N799, N210, N770, N33);
nor NOR3 (N805, N776, N351, N355);
and AND3 (N806, N804, N443, N708);
nor NOR3 (N807, N789, N754, N787);
and AND2 (N808, N781, N153);
or OR4 (N809, N807, N39, N187, N469);
buf BUF1 (N810, N808);
xor XOR2 (N811, N802, N402);
xor XOR2 (N812, N798, N792);
nor NOR2 (N813, N797, N81);
buf BUF1 (N814, N813);
nand NAND2 (N815, N809, N553);
nand NAND4 (N816, N814, N704, N134, N513);
not NOT1 (N817, N816);
nor NOR3 (N818, N801, N717, N707);
nor NOR3 (N819, N800, N320, N595);
not NOT1 (N820, N811);
xor XOR2 (N821, N818, N292);
nand NAND3 (N822, N820, N60, N572);
nor NOR2 (N823, N812, N420);
buf BUF1 (N824, N823);
buf BUF1 (N825, N803);
buf BUF1 (N826, N825);
xor XOR2 (N827, N821, N194);
nor NOR3 (N828, N826, N26, N373);
nand NAND2 (N829, N815, N53);
xor XOR2 (N830, N817, N15);
xor XOR2 (N831, N824, N378);
or OR2 (N832, N827, N723);
or OR4 (N833, N830, N830, N510, N498);
not NOT1 (N834, N833);
buf BUF1 (N835, N834);
and AND4 (N836, N819, N436, N262, N302);
nor NOR3 (N837, N806, N133, N696);
and AND3 (N838, N829, N253, N370);
not NOT1 (N839, N838);
not NOT1 (N840, N832);
or OR3 (N841, N837, N813, N403);
not NOT1 (N842, N839);
xor XOR2 (N843, N842, N509);
and AND4 (N844, N828, N253, N284, N38);
or OR3 (N845, N841, N369, N512);
xor XOR2 (N846, N822, N161);
not NOT1 (N847, N835);
buf BUF1 (N848, N845);
or OR3 (N849, N848, N187, N248);
xor XOR2 (N850, N847, N805);
nor NOR4 (N851, N769, N4, N441, N643);
nor NOR4 (N852, N831, N177, N87, N427);
not NOT1 (N853, N851);
or OR4 (N854, N840, N758, N209, N230);
or OR4 (N855, N843, N738, N229, N195);
or OR3 (N856, N852, N297, N247);
buf BUF1 (N857, N850);
and AND4 (N858, N857, N307, N55, N482);
nand NAND4 (N859, N836, N475, N406, N848);
or OR3 (N860, N844, N305, N549);
nand NAND3 (N861, N858, N727, N108);
or OR2 (N862, N860, N92);
nor NOR3 (N863, N846, N377, N701);
nor NOR2 (N864, N810, N760);
or OR4 (N865, N859, N79, N407, N347);
or OR2 (N866, N856, N643);
and AND2 (N867, N849, N824);
and AND4 (N868, N864, N846, N301, N287);
and AND2 (N869, N854, N282);
not NOT1 (N870, N869);
xor XOR2 (N871, N862, N553);
buf BUF1 (N872, N855);
buf BUF1 (N873, N872);
and AND3 (N874, N870, N58, N403);
or OR3 (N875, N853, N636, N525);
or OR3 (N876, N873, N622, N390);
buf BUF1 (N877, N871);
xor XOR2 (N878, N865, N115);
nand NAND2 (N879, N867, N155);
nand NAND4 (N880, N876, N309, N827, N281);
or OR2 (N881, N878, N742);
nand NAND3 (N882, N880, N163, N457);
and AND2 (N883, N868, N452);
nor NOR4 (N884, N882, N293, N824, N298);
buf BUF1 (N885, N874);
and AND4 (N886, N861, N787, N586, N208);
not NOT1 (N887, N877);
xor XOR2 (N888, N884, N704);
buf BUF1 (N889, N875);
nand NAND3 (N890, N887, N447, N454);
and AND4 (N891, N866, N23, N337, N368);
and AND2 (N892, N885, N438);
and AND3 (N893, N889, N484, N825);
and AND4 (N894, N891, N195, N109, N836);
nand NAND2 (N895, N888, N541);
nand NAND4 (N896, N886, N309, N183, N735);
buf BUF1 (N897, N883);
or OR2 (N898, N863, N252);
buf BUF1 (N899, N895);
and AND2 (N900, N897, N45);
not NOT1 (N901, N890);
not NOT1 (N902, N900);
not NOT1 (N903, N899);
buf BUF1 (N904, N896);
buf BUF1 (N905, N893);
xor XOR2 (N906, N903, N744);
nor NOR3 (N907, N904, N331, N718);
nand NAND3 (N908, N901, N189, N181);
buf BUF1 (N909, N898);
nand NAND2 (N910, N909, N263);
xor XOR2 (N911, N894, N145);
not NOT1 (N912, N907);
and AND3 (N913, N908, N216, N197);
and AND4 (N914, N881, N19, N561, N359);
xor XOR2 (N915, N906, N691);
buf BUF1 (N916, N892);
or OR3 (N917, N915, N230, N856);
nand NAND3 (N918, N910, N40, N501);
xor XOR2 (N919, N917, N207);
buf BUF1 (N920, N911);
not NOT1 (N921, N905);
and AND2 (N922, N918, N748);
and AND3 (N923, N913, N441, N797);
nand NAND2 (N924, N920, N658);
nand NAND4 (N925, N912, N691, N822, N529);
and AND3 (N926, N916, N267, N621);
buf BUF1 (N927, N922);
not NOT1 (N928, N927);
not NOT1 (N929, N914);
xor XOR2 (N930, N928, N362);
or OR2 (N931, N879, N617);
xor XOR2 (N932, N919, N254);
nor NOR2 (N933, N932, N64);
nand NAND4 (N934, N902, N345, N443, N707);
or OR3 (N935, N931, N415, N600);
not NOT1 (N936, N934);
or OR4 (N937, N936, N409, N646, N317);
xor XOR2 (N938, N930, N876);
nand NAND3 (N939, N937, N113, N529);
not NOT1 (N940, N933);
or OR2 (N941, N938, N434);
nor NOR2 (N942, N940, N350);
or OR4 (N943, N941, N709, N620, N314);
and AND3 (N944, N923, N237, N939);
not NOT1 (N945, N797);
xor XOR2 (N946, N945, N151);
xor XOR2 (N947, N926, N237);
or OR3 (N948, N947, N637, N803);
nor NOR2 (N949, N929, N740);
not NOT1 (N950, N949);
nand NAND3 (N951, N950, N877, N467);
nand NAND2 (N952, N943, N714);
and AND3 (N953, N944, N629, N201);
not NOT1 (N954, N924);
and AND3 (N955, N954, N842, N615);
xor XOR2 (N956, N951, N377);
nor NOR3 (N957, N921, N77, N81);
nand NAND2 (N958, N946, N449);
nor NOR3 (N959, N942, N699, N229);
nand NAND3 (N960, N956, N592, N632);
nand NAND3 (N961, N957, N503, N691);
buf BUF1 (N962, N961);
buf BUF1 (N963, N955);
and AND2 (N964, N958, N299);
xor XOR2 (N965, N948, N590);
and AND4 (N966, N960, N311, N650, N892);
and AND2 (N967, N925, N646);
and AND4 (N968, N953, N956, N961, N397);
xor XOR2 (N969, N959, N720);
not NOT1 (N970, N964);
or OR2 (N971, N968, N749);
and AND4 (N972, N967, N629, N269, N842);
nor NOR2 (N973, N935, N748);
nor NOR3 (N974, N965, N770, N66);
nor NOR2 (N975, N971, N73);
xor XOR2 (N976, N952, N969);
and AND2 (N977, N213, N433);
xor XOR2 (N978, N975, N631);
nand NAND2 (N979, N970, N170);
and AND4 (N980, N979, N55, N404, N95);
buf BUF1 (N981, N980);
and AND4 (N982, N966, N622, N264, N134);
not NOT1 (N983, N963);
nor NOR3 (N984, N983, N266, N347);
nand NAND2 (N985, N978, N655);
nor NOR2 (N986, N984, N260);
nor NOR2 (N987, N981, N668);
buf BUF1 (N988, N982);
not NOT1 (N989, N985);
buf BUF1 (N990, N972);
nor NOR3 (N991, N989, N208, N259);
xor XOR2 (N992, N986, N895);
and AND3 (N993, N987, N331, N201);
buf BUF1 (N994, N976);
and AND4 (N995, N973, N197, N259, N464);
and AND2 (N996, N962, N57);
not NOT1 (N997, N993);
nand NAND3 (N998, N994, N927, N163);
buf BUF1 (N999, N992);
nor NOR2 (N1000, N990, N597);
nand NAND4 (N1001, N997, N753, N241, N669);
buf BUF1 (N1002, N1000);
not NOT1 (N1003, N977);
buf BUF1 (N1004, N999);
buf BUF1 (N1005, N998);
and AND4 (N1006, N991, N970, N556, N491);
buf BUF1 (N1007, N974);
and AND2 (N1008, N1001, N761);
xor XOR2 (N1009, N1008, N288);
not NOT1 (N1010, N995);
buf BUF1 (N1011, N988);
or OR2 (N1012, N1007, N994);
xor XOR2 (N1013, N1005, N833);
nor NOR4 (N1014, N1012, N835, N505, N918);
nor NOR3 (N1015, N1002, N744, N166);
xor XOR2 (N1016, N1006, N463);
or OR4 (N1017, N1013, N338, N573, N803);
or OR2 (N1018, N1003, N703);
or OR2 (N1019, N1018, N295);
buf BUF1 (N1020, N1016);
xor XOR2 (N1021, N1019, N761);
or OR2 (N1022, N996, N741);
or OR4 (N1023, N1017, N675, N886, N552);
xor XOR2 (N1024, N1022, N1022);
and AND4 (N1025, N1015, N375, N521, N95);
and AND4 (N1026, N1010, N642, N780, N393);
not NOT1 (N1027, N1026);
not NOT1 (N1028, N1004);
nand NAND2 (N1029, N1009, N318);
not NOT1 (N1030, N1023);
not NOT1 (N1031, N1027);
xor XOR2 (N1032, N1021, N210);
nor NOR4 (N1033, N1029, N653, N80, N228);
and AND3 (N1034, N1028, N789, N904);
xor XOR2 (N1035, N1033, N211);
xor XOR2 (N1036, N1030, N683);
nand NAND3 (N1037, N1036, N242, N909);
buf BUF1 (N1038, N1014);
buf BUF1 (N1039, N1024);
buf BUF1 (N1040, N1031);
buf BUF1 (N1041, N1032);
buf BUF1 (N1042, N1041);
not NOT1 (N1043, N1039);
nor NOR4 (N1044, N1042, N47, N1041, N715);
buf BUF1 (N1045, N1040);
or OR2 (N1046, N1020, N893);
buf BUF1 (N1047, N1037);
not NOT1 (N1048, N1044);
xor XOR2 (N1049, N1011, N960);
buf BUF1 (N1050, N1043);
not NOT1 (N1051, N1045);
nor NOR2 (N1052, N1049, N302);
nand NAND3 (N1053, N1046, N292, N956);
nor NOR3 (N1054, N1025, N671, N849);
xor XOR2 (N1055, N1047, N180);
buf BUF1 (N1056, N1053);
not NOT1 (N1057, N1035);
nor NOR2 (N1058, N1034, N989);
and AND4 (N1059, N1056, N851, N996, N971);
nor NOR2 (N1060, N1048, N703);
nor NOR2 (N1061, N1052, N126);
nand NAND3 (N1062, N1050, N148, N790);
buf BUF1 (N1063, N1057);
or OR2 (N1064, N1051, N219);
buf BUF1 (N1065, N1038);
and AND4 (N1066, N1055, N240, N836, N894);
nor NOR3 (N1067, N1058, N313, N303);
buf BUF1 (N1068, N1064);
or OR3 (N1069, N1068, N774, N1009);
xor XOR2 (N1070, N1067, N530);
and AND2 (N1071, N1059, N388);
not NOT1 (N1072, N1066);
xor XOR2 (N1073, N1070, N611);
nor NOR3 (N1074, N1069, N47, N740);
xor XOR2 (N1075, N1063, N877);
nor NOR2 (N1076, N1071, N238);
xor XOR2 (N1077, N1060, N1015);
not NOT1 (N1078, N1061);
nor NOR4 (N1079, N1078, N553, N341, N647);
buf BUF1 (N1080, N1072);
or OR3 (N1081, N1080, N644, N501);
or OR3 (N1082, N1079, N7, N71);
not NOT1 (N1083, N1081);
not NOT1 (N1084, N1076);
not NOT1 (N1085, N1062);
or OR3 (N1086, N1074, N994, N840);
not NOT1 (N1087, N1075);
buf BUF1 (N1088, N1082);
and AND4 (N1089, N1073, N599, N484, N264);
nand NAND3 (N1090, N1077, N88, N1062);
nand NAND4 (N1091, N1089, N447, N81, N619);
nor NOR3 (N1092, N1086, N215, N99);
nand NAND4 (N1093, N1054, N104, N142, N645);
or OR4 (N1094, N1085, N860, N639, N17);
xor XOR2 (N1095, N1090, N1026);
not NOT1 (N1096, N1091);
xor XOR2 (N1097, N1084, N561);
not NOT1 (N1098, N1096);
xor XOR2 (N1099, N1065, N4);
buf BUF1 (N1100, N1087);
not NOT1 (N1101, N1095);
and AND2 (N1102, N1088, N952);
nand NAND4 (N1103, N1097, N806, N650, N727);
xor XOR2 (N1104, N1093, N902);
and AND3 (N1105, N1083, N947, N638);
not NOT1 (N1106, N1105);
not NOT1 (N1107, N1102);
buf BUF1 (N1108, N1092);
not NOT1 (N1109, N1094);
not NOT1 (N1110, N1106);
nor NOR2 (N1111, N1109, N511);
buf BUF1 (N1112, N1098);
not NOT1 (N1113, N1110);
buf BUF1 (N1114, N1103);
buf BUF1 (N1115, N1101);
nand NAND4 (N1116, N1115, N451, N856, N296);
xor XOR2 (N1117, N1104, N818);
not NOT1 (N1118, N1113);
and AND3 (N1119, N1116, N28, N177);
nor NOR4 (N1120, N1117, N33, N410, N1084);
nor NOR3 (N1121, N1100, N744, N800);
not NOT1 (N1122, N1120);
not NOT1 (N1123, N1118);
buf BUF1 (N1124, N1111);
or OR4 (N1125, N1107, N1035, N392, N364);
xor XOR2 (N1126, N1108, N145);
xor XOR2 (N1127, N1124, N223);
or OR2 (N1128, N1121, N451);
or OR3 (N1129, N1099, N869, N60);
nor NOR4 (N1130, N1123, N43, N1008, N176);
xor XOR2 (N1131, N1127, N243);
nand NAND3 (N1132, N1119, N203, N161);
and AND2 (N1133, N1114, N413);
nor NOR4 (N1134, N1132, N206, N96, N791);
buf BUF1 (N1135, N1122);
buf BUF1 (N1136, N1128);
xor XOR2 (N1137, N1112, N137);
and AND2 (N1138, N1129, N958);
buf BUF1 (N1139, N1125);
or OR2 (N1140, N1126, N644);
buf BUF1 (N1141, N1140);
nand NAND3 (N1142, N1137, N960, N1013);
nor NOR3 (N1143, N1135, N306, N725);
not NOT1 (N1144, N1134);
buf BUF1 (N1145, N1136);
buf BUF1 (N1146, N1145);
nor NOR3 (N1147, N1131, N370, N342);
or OR3 (N1148, N1130, N175, N680);
nor NOR2 (N1149, N1133, N1044);
buf BUF1 (N1150, N1141);
or OR2 (N1151, N1150, N505);
xor XOR2 (N1152, N1142, N381);
and AND2 (N1153, N1149, N341);
nor NOR4 (N1154, N1152, N317, N746, N74);
nor NOR4 (N1155, N1144, N1141, N476, N31);
buf BUF1 (N1156, N1138);
nand NAND4 (N1157, N1148, N95, N880, N875);
and AND4 (N1158, N1147, N184, N326, N856);
xor XOR2 (N1159, N1158, N1151);
buf BUF1 (N1160, N489);
nor NOR2 (N1161, N1157, N277);
buf BUF1 (N1162, N1156);
not NOT1 (N1163, N1159);
nand NAND3 (N1164, N1143, N505, N329);
and AND2 (N1165, N1163, N299);
nand NAND3 (N1166, N1153, N384, N651);
nor NOR2 (N1167, N1161, N773);
nand NAND3 (N1168, N1154, N1143, N963);
nor NOR4 (N1169, N1160, N102, N334, N1023);
or OR3 (N1170, N1165, N686, N506);
and AND2 (N1171, N1164, N919);
nand NAND2 (N1172, N1170, N815);
or OR2 (N1173, N1168, N897);
buf BUF1 (N1174, N1173);
or OR3 (N1175, N1155, N743, N406);
xor XOR2 (N1176, N1146, N528);
xor XOR2 (N1177, N1139, N718);
not NOT1 (N1178, N1166);
buf BUF1 (N1179, N1174);
xor XOR2 (N1180, N1175, N683);
xor XOR2 (N1181, N1172, N777);
and AND3 (N1182, N1180, N808, N714);
buf BUF1 (N1183, N1182);
nand NAND2 (N1184, N1169, N1152);
and AND2 (N1185, N1183, N1020);
xor XOR2 (N1186, N1171, N606);
not NOT1 (N1187, N1186);
xor XOR2 (N1188, N1162, N342);
and AND4 (N1189, N1176, N274, N679, N299);
and AND2 (N1190, N1177, N713);
xor XOR2 (N1191, N1187, N340);
not NOT1 (N1192, N1191);
or OR4 (N1193, N1188, N326, N888, N405);
buf BUF1 (N1194, N1178);
nand NAND4 (N1195, N1194, N516, N201, N121);
buf BUF1 (N1196, N1192);
or OR4 (N1197, N1181, N734, N403, N1040);
and AND2 (N1198, N1190, N1143);
and AND2 (N1199, N1197, N578);
not NOT1 (N1200, N1196);
xor XOR2 (N1201, N1195, N805);
nand NAND4 (N1202, N1198, N906, N979, N25);
buf BUF1 (N1203, N1179);
buf BUF1 (N1204, N1167);
or OR3 (N1205, N1202, N49, N94);
nand NAND4 (N1206, N1189, N699, N440, N855);
nor NOR3 (N1207, N1206, N822, N477);
nand NAND2 (N1208, N1205, N971);
not NOT1 (N1209, N1201);
and AND4 (N1210, N1203, N828, N47, N188);
nor NOR2 (N1211, N1207, N517);
or OR4 (N1212, N1210, N1105, N210, N345);
xor XOR2 (N1213, N1185, N814);
nor NOR4 (N1214, N1199, N173, N846, N117);
not NOT1 (N1215, N1212);
buf BUF1 (N1216, N1209);
xor XOR2 (N1217, N1193, N588);
nand NAND3 (N1218, N1213, N362, N954);
buf BUF1 (N1219, N1184);
buf BUF1 (N1220, N1217);
and AND2 (N1221, N1218, N1142);
or OR3 (N1222, N1204, N771, N531);
buf BUF1 (N1223, N1220);
or OR3 (N1224, N1208, N151, N648);
nand NAND3 (N1225, N1216, N1152, N1194);
xor XOR2 (N1226, N1222, N875);
buf BUF1 (N1227, N1225);
buf BUF1 (N1228, N1223);
buf BUF1 (N1229, N1215);
buf BUF1 (N1230, N1224);
xor XOR2 (N1231, N1228, N712);
nand NAND2 (N1232, N1231, N354);
nand NAND3 (N1233, N1226, N435, N930);
or OR4 (N1234, N1232, N618, N642, N570);
nor NOR3 (N1235, N1211, N47, N1134);
buf BUF1 (N1236, N1234);
xor XOR2 (N1237, N1214, N199);
or OR4 (N1238, N1219, N56, N515, N991);
not NOT1 (N1239, N1227);
and AND4 (N1240, N1200, N660, N798, N625);
xor XOR2 (N1241, N1233, N449);
nand NAND3 (N1242, N1229, N1179, N7);
not NOT1 (N1243, N1241);
nor NOR2 (N1244, N1242, N951);
buf BUF1 (N1245, N1237);
xor XOR2 (N1246, N1238, N344);
nand NAND3 (N1247, N1239, N993, N139);
nand NAND2 (N1248, N1240, N153);
not NOT1 (N1249, N1245);
and AND2 (N1250, N1244, N91);
or OR2 (N1251, N1247, N423);
xor XOR2 (N1252, N1236, N810);
not NOT1 (N1253, N1243);
xor XOR2 (N1254, N1248, N38);
nand NAND3 (N1255, N1235, N472, N1244);
or OR3 (N1256, N1249, N26, N538);
or OR4 (N1257, N1254, N433, N965, N673);
or OR4 (N1258, N1252, N159, N240, N139);
nor NOR4 (N1259, N1246, N831, N442, N465);
nand NAND4 (N1260, N1257, N740, N1244, N514);
nand NAND3 (N1261, N1260, N850, N243);
nand NAND3 (N1262, N1259, N336, N537);
nand NAND3 (N1263, N1255, N813, N239);
buf BUF1 (N1264, N1251);
xor XOR2 (N1265, N1230, N918);
nor NOR3 (N1266, N1261, N1088, N617);
or OR4 (N1267, N1263, N1221, N787, N977);
not NOT1 (N1268, N143);
not NOT1 (N1269, N1266);
and AND4 (N1270, N1268, N1051, N737, N906);
nor NOR2 (N1271, N1264, N1213);
and AND4 (N1272, N1258, N607, N100, N1045);
nor NOR2 (N1273, N1256, N383);
nand NAND3 (N1274, N1265, N809, N1138);
nand NAND4 (N1275, N1274, N778, N1033, N59);
not NOT1 (N1276, N1271);
xor XOR2 (N1277, N1267, N822);
buf BUF1 (N1278, N1269);
buf BUF1 (N1279, N1276);
or OR4 (N1280, N1253, N784, N1001, N249);
buf BUF1 (N1281, N1273);
nor NOR2 (N1282, N1281, N30);
or OR4 (N1283, N1278, N576, N60, N312);
xor XOR2 (N1284, N1280, N277);
not NOT1 (N1285, N1277);
or OR3 (N1286, N1279, N259, N1091);
xor XOR2 (N1287, N1270, N426);
not NOT1 (N1288, N1284);
and AND4 (N1289, N1287, N941, N228, N757);
nor NOR2 (N1290, N1275, N597);
and AND2 (N1291, N1286, N943);
and AND4 (N1292, N1291, N914, N97, N607);
or OR3 (N1293, N1289, N408, N880);
xor XOR2 (N1294, N1282, N1048);
xor XOR2 (N1295, N1288, N1083);
xor XOR2 (N1296, N1293, N266);
xor XOR2 (N1297, N1295, N244);
not NOT1 (N1298, N1290);
not NOT1 (N1299, N1285);
not NOT1 (N1300, N1250);
buf BUF1 (N1301, N1296);
xor XOR2 (N1302, N1297, N699);
buf BUF1 (N1303, N1301);
nand NAND4 (N1304, N1298, N859, N889, N390);
xor XOR2 (N1305, N1262, N1183);
buf BUF1 (N1306, N1294);
nand NAND4 (N1307, N1292, N771, N793, N406);
not NOT1 (N1308, N1299);
nand NAND4 (N1309, N1303, N1136, N767, N1210);
not NOT1 (N1310, N1304);
and AND4 (N1311, N1308, N406, N665, N723);
nand NAND4 (N1312, N1306, N751, N258, N329);
xor XOR2 (N1313, N1302, N223);
or OR2 (N1314, N1309, N341);
and AND2 (N1315, N1307, N1168);
xor XOR2 (N1316, N1311, N386);
nor NOR2 (N1317, N1283, N816);
and AND2 (N1318, N1300, N1254);
not NOT1 (N1319, N1310);
buf BUF1 (N1320, N1272);
nand NAND3 (N1321, N1319, N630, N524);
nand NAND4 (N1322, N1313, N617, N1198, N659);
not NOT1 (N1323, N1318);
buf BUF1 (N1324, N1316);
xor XOR2 (N1325, N1312, N940);
nand NAND2 (N1326, N1322, N937);
not NOT1 (N1327, N1315);
or OR4 (N1328, N1323, N370, N343, N1195);
not NOT1 (N1329, N1328);
xor XOR2 (N1330, N1327, N367);
not NOT1 (N1331, N1320);
or OR3 (N1332, N1325, N843, N219);
nand NAND3 (N1333, N1330, N1115, N584);
not NOT1 (N1334, N1321);
buf BUF1 (N1335, N1326);
or OR2 (N1336, N1331, N1282);
buf BUF1 (N1337, N1335);
nor NOR3 (N1338, N1334, N80, N186);
or OR2 (N1339, N1314, N462);
and AND4 (N1340, N1333, N505, N167, N869);
or OR4 (N1341, N1340, N71, N266, N427);
and AND4 (N1342, N1341, N228, N375, N1239);
buf BUF1 (N1343, N1317);
xor XOR2 (N1344, N1338, N1124);
and AND3 (N1345, N1339, N653, N1010);
not NOT1 (N1346, N1336);
and AND3 (N1347, N1345, N18, N75);
nor NOR4 (N1348, N1347, N326, N491, N52);
or OR4 (N1349, N1329, N727, N948, N427);
xor XOR2 (N1350, N1305, N351);
and AND4 (N1351, N1324, N265, N1341, N994);
buf BUF1 (N1352, N1342);
nor NOR2 (N1353, N1343, N1066);
nor NOR4 (N1354, N1353, N234, N864, N160);
not NOT1 (N1355, N1344);
not NOT1 (N1356, N1354);
nand NAND4 (N1357, N1348, N272, N601, N473);
xor XOR2 (N1358, N1349, N767);
not NOT1 (N1359, N1352);
buf BUF1 (N1360, N1357);
not NOT1 (N1361, N1359);
xor XOR2 (N1362, N1332, N719);
nand NAND3 (N1363, N1337, N811, N47);
buf BUF1 (N1364, N1355);
not NOT1 (N1365, N1364);
and AND3 (N1366, N1351, N804, N997);
and AND4 (N1367, N1356, N1043, N737, N1259);
or OR3 (N1368, N1367, N1061, N475);
not NOT1 (N1369, N1360);
xor XOR2 (N1370, N1369, N1296);
and AND2 (N1371, N1363, N910);
xor XOR2 (N1372, N1370, N1014);
xor XOR2 (N1373, N1358, N616);
or OR3 (N1374, N1372, N702, N406);
nand NAND3 (N1375, N1350, N751, N881);
or OR2 (N1376, N1375, N108);
buf BUF1 (N1377, N1376);
and AND4 (N1378, N1373, N1249, N1018, N458);
or OR3 (N1379, N1362, N934, N1258);
nand NAND2 (N1380, N1346, N1310);
xor XOR2 (N1381, N1377, N25);
xor XOR2 (N1382, N1381, N221);
buf BUF1 (N1383, N1371);
buf BUF1 (N1384, N1365);
not NOT1 (N1385, N1382);
or OR2 (N1386, N1379, N755);
buf BUF1 (N1387, N1361);
nor NOR4 (N1388, N1380, N217, N149, N1074);
and AND2 (N1389, N1388, N649);
buf BUF1 (N1390, N1389);
or OR3 (N1391, N1374, N641, N307);
not NOT1 (N1392, N1366);
nand NAND3 (N1393, N1385, N1352, N554);
nand NAND2 (N1394, N1378, N465);
not NOT1 (N1395, N1393);
and AND4 (N1396, N1383, N1252, N502, N1115);
nand NAND4 (N1397, N1384, N7, N228, N1054);
xor XOR2 (N1398, N1386, N702);
nand NAND4 (N1399, N1395, N432, N1315, N517);
xor XOR2 (N1400, N1398, N651);
or OR4 (N1401, N1392, N758, N1179, N601);
nand NAND2 (N1402, N1368, N379);
and AND4 (N1403, N1394, N297, N644, N1261);
not NOT1 (N1404, N1397);
xor XOR2 (N1405, N1402, N499);
nor NOR2 (N1406, N1403, N79);
buf BUF1 (N1407, N1396);
buf BUF1 (N1408, N1390);
nor NOR4 (N1409, N1406, N1092, N296, N223);
or OR3 (N1410, N1387, N752, N528);
or OR4 (N1411, N1391, N1339, N1369, N1257);
nor NOR4 (N1412, N1410, N1363, N724, N367);
nor NOR2 (N1413, N1408, N163);
nor NOR3 (N1414, N1401, N173, N59);
or OR4 (N1415, N1399, N239, N968, N1241);
buf BUF1 (N1416, N1409);
not NOT1 (N1417, N1414);
buf BUF1 (N1418, N1417);
and AND3 (N1419, N1404, N184, N1275);
xor XOR2 (N1420, N1419, N1062);
buf BUF1 (N1421, N1405);
buf BUF1 (N1422, N1418);
nand NAND3 (N1423, N1420, N459, N1233);
not NOT1 (N1424, N1407);
not NOT1 (N1425, N1423);
nor NOR3 (N1426, N1411, N1029, N755);
buf BUF1 (N1427, N1424);
nor NOR2 (N1428, N1413, N85);
nor NOR4 (N1429, N1421, N1011, N620, N1328);
nor NOR2 (N1430, N1412, N854);
or OR3 (N1431, N1426, N11, N855);
not NOT1 (N1432, N1430);
not NOT1 (N1433, N1428);
and AND2 (N1434, N1432, N1429);
nand NAND4 (N1435, N1250, N452, N409, N1292);
buf BUF1 (N1436, N1427);
xor XOR2 (N1437, N1434, N366);
xor XOR2 (N1438, N1433, N616);
and AND4 (N1439, N1437, N1173, N1436, N694);
buf BUF1 (N1440, N1114);
nor NOR4 (N1441, N1435, N220, N507, N603);
nand NAND2 (N1442, N1416, N635);
not NOT1 (N1443, N1442);
not NOT1 (N1444, N1415);
nor NOR2 (N1445, N1422, N652);
nor NOR2 (N1446, N1431, N993);
buf BUF1 (N1447, N1445);
xor XOR2 (N1448, N1447, N1166);
nand NAND2 (N1449, N1446, N1126);
not NOT1 (N1450, N1449);
and AND2 (N1451, N1400, N151);
not NOT1 (N1452, N1450);
and AND3 (N1453, N1451, N41, N478);
or OR4 (N1454, N1444, N79, N1402, N1119);
xor XOR2 (N1455, N1439, N635);
nor NOR3 (N1456, N1440, N1141, N987);
nor NOR2 (N1457, N1441, N275);
xor XOR2 (N1458, N1454, N335);
and AND3 (N1459, N1455, N1450, N918);
not NOT1 (N1460, N1457);
nand NAND4 (N1461, N1452, N828, N571, N543);
buf BUF1 (N1462, N1453);
buf BUF1 (N1463, N1461);
xor XOR2 (N1464, N1425, N1096);
nor NOR4 (N1465, N1438, N169, N1221, N690);
not NOT1 (N1466, N1458);
xor XOR2 (N1467, N1465, N1095);
or OR4 (N1468, N1467, N503, N1230, N224);
xor XOR2 (N1469, N1463, N801);
nand NAND2 (N1470, N1464, N2);
nor NOR2 (N1471, N1466, N493);
or OR4 (N1472, N1443, N355, N324, N553);
buf BUF1 (N1473, N1460);
nor NOR2 (N1474, N1470, N358);
and AND2 (N1475, N1473, N1354);
nand NAND3 (N1476, N1475, N1143, N1330);
and AND3 (N1477, N1472, N1242, N266);
nor NOR3 (N1478, N1474, N952, N164);
and AND3 (N1479, N1459, N1392, N1190);
nand NAND2 (N1480, N1456, N769);
or OR2 (N1481, N1462, N909);
nor NOR2 (N1482, N1480, N1410);
and AND2 (N1483, N1477, N315);
or OR4 (N1484, N1479, N111, N1214, N323);
buf BUF1 (N1485, N1469);
nand NAND4 (N1486, N1468, N788, N28, N797);
buf BUF1 (N1487, N1481);
xor XOR2 (N1488, N1487, N1008);
nand NAND2 (N1489, N1476, N251);
nand NAND2 (N1490, N1484, N595);
not NOT1 (N1491, N1482);
nand NAND2 (N1492, N1478, N1035);
nor NOR2 (N1493, N1490, N1020);
nand NAND3 (N1494, N1491, N866, N329);
not NOT1 (N1495, N1494);
and AND3 (N1496, N1486, N493, N375);
nand NAND2 (N1497, N1448, N974);
and AND4 (N1498, N1483, N1137, N43, N1201);
or OR2 (N1499, N1488, N503);
and AND2 (N1500, N1496, N14);
buf BUF1 (N1501, N1499);
and AND4 (N1502, N1471, N753, N472, N744);
and AND4 (N1503, N1493, N301, N1220, N1456);
not NOT1 (N1504, N1501);
not NOT1 (N1505, N1485);
not NOT1 (N1506, N1489);
not NOT1 (N1507, N1502);
not NOT1 (N1508, N1498);
not NOT1 (N1509, N1508);
and AND2 (N1510, N1509, N577);
xor XOR2 (N1511, N1504, N859);
nor NOR2 (N1512, N1507, N173);
buf BUF1 (N1513, N1500);
nand NAND3 (N1514, N1503, N364, N584);
xor XOR2 (N1515, N1505, N1274);
nand NAND4 (N1516, N1511, N286, N1115, N1161);
and AND2 (N1517, N1497, N557);
not NOT1 (N1518, N1495);
or OR4 (N1519, N1516, N1408, N274, N1129);
buf BUF1 (N1520, N1515);
buf BUF1 (N1521, N1506);
not NOT1 (N1522, N1521);
nor NOR3 (N1523, N1522, N517, N1323);
or OR4 (N1524, N1517, N1318, N929, N330);
nor NOR2 (N1525, N1492, N462);
nand NAND2 (N1526, N1512, N499);
nand NAND2 (N1527, N1514, N472);
nor NOR4 (N1528, N1519, N701, N800, N1403);
and AND2 (N1529, N1510, N91);
nand NAND2 (N1530, N1518, N1496);
nand NAND2 (N1531, N1525, N1267);
xor XOR2 (N1532, N1527, N505);
nand NAND3 (N1533, N1523, N901, N313);
xor XOR2 (N1534, N1530, N88);
buf BUF1 (N1535, N1531);
and AND2 (N1536, N1513, N1476);
nor NOR2 (N1537, N1534, N1447);
nand NAND4 (N1538, N1532, N584, N1242, N966);
xor XOR2 (N1539, N1538, N508);
nor NOR3 (N1540, N1529, N1019, N1284);
or OR2 (N1541, N1524, N873);
or OR2 (N1542, N1520, N1267);
buf BUF1 (N1543, N1536);
not NOT1 (N1544, N1526);
buf BUF1 (N1545, N1533);
or OR3 (N1546, N1540, N832, N798);
or OR4 (N1547, N1541, N1347, N1199, N210);
or OR3 (N1548, N1542, N596, N264);
and AND3 (N1549, N1543, N1372, N846);
nor NOR2 (N1550, N1548, N1177);
nand NAND3 (N1551, N1535, N221, N848);
and AND3 (N1552, N1528, N273, N901);
buf BUF1 (N1553, N1551);
nand NAND3 (N1554, N1544, N327, N902);
and AND4 (N1555, N1547, N802, N615, N1148);
nor NOR3 (N1556, N1549, N929, N665);
not NOT1 (N1557, N1545);
nor NOR2 (N1558, N1537, N118);
nor NOR4 (N1559, N1557, N691, N1277, N238);
not NOT1 (N1560, N1556);
not NOT1 (N1561, N1546);
nor NOR2 (N1562, N1558, N852);
xor XOR2 (N1563, N1552, N1172);
nand NAND4 (N1564, N1553, N151, N1052, N1450);
buf BUF1 (N1565, N1563);
nand NAND2 (N1566, N1565, N1523);
not NOT1 (N1567, N1539);
buf BUF1 (N1568, N1560);
nand NAND2 (N1569, N1564, N356);
and AND4 (N1570, N1569, N192, N613, N851);
and AND4 (N1571, N1559, N589, N1175, N464);
not NOT1 (N1572, N1555);
nand NAND2 (N1573, N1561, N1085);
and AND3 (N1574, N1573, N216, N612);
or OR3 (N1575, N1554, N294, N1118);
xor XOR2 (N1576, N1575, N601);
buf BUF1 (N1577, N1576);
buf BUF1 (N1578, N1574);
xor XOR2 (N1579, N1567, N1190);
or OR3 (N1580, N1550, N1218, N1300);
buf BUF1 (N1581, N1566);
nor NOR2 (N1582, N1580, N29);
not NOT1 (N1583, N1571);
nor NOR3 (N1584, N1578, N1231, N371);
buf BUF1 (N1585, N1584);
not NOT1 (N1586, N1577);
and AND3 (N1587, N1586, N547, N1366);
or OR3 (N1588, N1587, N872, N357);
nand NAND4 (N1589, N1568, N1147, N266, N381);
xor XOR2 (N1590, N1579, N238);
or OR4 (N1591, N1589, N798, N311, N1247);
not NOT1 (N1592, N1591);
nand NAND4 (N1593, N1570, N739, N1172, N1283);
or OR2 (N1594, N1562, N971);
nor NOR4 (N1595, N1594, N1498, N253, N35);
buf BUF1 (N1596, N1588);
xor XOR2 (N1597, N1595, N66);
nor NOR2 (N1598, N1592, N1153);
buf BUF1 (N1599, N1582);
nor NOR2 (N1600, N1598, N613);
not NOT1 (N1601, N1590);
or OR2 (N1602, N1596, N897);
and AND2 (N1603, N1599, N926);
buf BUF1 (N1604, N1600);
buf BUF1 (N1605, N1585);
xor XOR2 (N1606, N1602, N630);
nand NAND4 (N1607, N1603, N504, N717, N485);
xor XOR2 (N1608, N1593, N685);
or OR2 (N1609, N1583, N899);
and AND4 (N1610, N1607, N753, N1033, N243);
buf BUF1 (N1611, N1610);
nor NOR3 (N1612, N1581, N343, N130);
xor XOR2 (N1613, N1604, N135);
not NOT1 (N1614, N1605);
and AND4 (N1615, N1572, N544, N1311, N1007);
nor NOR3 (N1616, N1597, N1234, N126);
nand NAND4 (N1617, N1612, N381, N1054, N445);
and AND3 (N1618, N1606, N804, N1501);
xor XOR2 (N1619, N1611, N1558);
nand NAND2 (N1620, N1619, N774);
nand NAND3 (N1621, N1620, N1481, N791);
buf BUF1 (N1622, N1616);
xor XOR2 (N1623, N1613, N1121);
buf BUF1 (N1624, N1617);
buf BUF1 (N1625, N1615);
buf BUF1 (N1626, N1622);
and AND4 (N1627, N1621, N919, N456, N1209);
or OR3 (N1628, N1614, N787, N373);
and AND3 (N1629, N1623, N1120, N404);
nor NOR4 (N1630, N1626, N934, N1191, N225);
nand NAND3 (N1631, N1624, N1085, N303);
xor XOR2 (N1632, N1608, N188);
and AND2 (N1633, N1601, N1357);
and AND3 (N1634, N1628, N996, N1411);
and AND3 (N1635, N1631, N879, N1007);
nor NOR2 (N1636, N1635, N244);
and AND4 (N1637, N1632, N1001, N804, N635);
buf BUF1 (N1638, N1633);
xor XOR2 (N1639, N1638, N444);
or OR3 (N1640, N1639, N809, N126);
and AND4 (N1641, N1636, N1534, N1473, N1056);
xor XOR2 (N1642, N1641, N1001);
nand NAND3 (N1643, N1625, N267, N758);
nand NAND4 (N1644, N1629, N1465, N753, N277);
not NOT1 (N1645, N1637);
not NOT1 (N1646, N1640);
and AND3 (N1647, N1642, N1506, N1157);
xor XOR2 (N1648, N1647, N1358);
or OR2 (N1649, N1643, N640);
buf BUF1 (N1650, N1646);
nand NAND4 (N1651, N1644, N1191, N184, N1443);
not NOT1 (N1652, N1650);
buf BUF1 (N1653, N1609);
nand NAND2 (N1654, N1651, N1536);
xor XOR2 (N1655, N1652, N1137);
nand NAND2 (N1656, N1630, N612);
nor NOR2 (N1657, N1634, N216);
nand NAND2 (N1658, N1649, N1363);
or OR4 (N1659, N1654, N609, N878, N270);
nor NOR3 (N1660, N1645, N1165, N181);
or OR3 (N1661, N1655, N1650, N737);
and AND2 (N1662, N1627, N144);
nor NOR4 (N1663, N1659, N1528, N1586, N433);
xor XOR2 (N1664, N1653, N1254);
nor NOR2 (N1665, N1660, N695);
xor XOR2 (N1666, N1665, N1128);
and AND3 (N1667, N1664, N1608, N410);
or OR3 (N1668, N1656, N86, N1212);
nand NAND2 (N1669, N1662, N652);
xor XOR2 (N1670, N1618, N547);
buf BUF1 (N1671, N1670);
buf BUF1 (N1672, N1667);
nand NAND3 (N1673, N1671, N1035, N804);
not NOT1 (N1674, N1669);
xor XOR2 (N1675, N1661, N92);
buf BUF1 (N1676, N1668);
buf BUF1 (N1677, N1674);
and AND3 (N1678, N1673, N289, N423);
buf BUF1 (N1679, N1676);
or OR4 (N1680, N1658, N25, N322, N17);
nand NAND2 (N1681, N1678, N700);
nand NAND3 (N1682, N1672, N876, N953);
xor XOR2 (N1683, N1677, N937);
not NOT1 (N1684, N1683);
or OR2 (N1685, N1657, N902);
xor XOR2 (N1686, N1648, N600);
not NOT1 (N1687, N1680);
nand NAND4 (N1688, N1666, N1581, N646, N1338);
not NOT1 (N1689, N1681);
and AND3 (N1690, N1675, N1517, N240);
nand NAND2 (N1691, N1684, N237);
nor NOR4 (N1692, N1686, N1398, N1199, N540);
not NOT1 (N1693, N1691);
nand NAND2 (N1694, N1693, N1637);
or OR4 (N1695, N1679, N1625, N893, N1179);
xor XOR2 (N1696, N1690, N200);
or OR4 (N1697, N1682, N233, N1294, N76);
nor NOR2 (N1698, N1663, N1209);
and AND4 (N1699, N1698, N673, N1575, N1035);
not NOT1 (N1700, N1688);
and AND2 (N1701, N1699, N246);
and AND3 (N1702, N1687, N1381, N416);
and AND3 (N1703, N1694, N1186, N1620);
or OR3 (N1704, N1685, N60, N1670);
not NOT1 (N1705, N1696);
and AND2 (N1706, N1701, N1188);
buf BUF1 (N1707, N1705);
nor NOR3 (N1708, N1704, N790, N115);
nor NOR3 (N1709, N1689, N1491, N232);
nand NAND3 (N1710, N1708, N1118, N1444);
not NOT1 (N1711, N1700);
and AND3 (N1712, N1703, N1489, N356);
or OR3 (N1713, N1707, N732, N1557);
xor XOR2 (N1714, N1697, N1454);
nor NOR3 (N1715, N1692, N294, N293);
xor XOR2 (N1716, N1711, N559);
not NOT1 (N1717, N1713);
or OR2 (N1718, N1702, N172);
xor XOR2 (N1719, N1716, N434);
nor NOR2 (N1720, N1719, N773);
xor XOR2 (N1721, N1706, N668);
nand NAND3 (N1722, N1709, N764, N1624);
or OR3 (N1723, N1714, N397, N1665);
xor XOR2 (N1724, N1723, N1142);
nor NOR4 (N1725, N1717, N260, N1631, N278);
and AND2 (N1726, N1720, N1218);
buf BUF1 (N1727, N1724);
and AND3 (N1728, N1722, N1326, N66);
and AND3 (N1729, N1712, N1593, N1277);
and AND3 (N1730, N1727, N1628, N1131);
nand NAND4 (N1731, N1695, N944, N1725, N1049);
and AND2 (N1732, N1020, N993);
buf BUF1 (N1733, N1729);
xor XOR2 (N1734, N1721, N714);
not NOT1 (N1735, N1710);
buf BUF1 (N1736, N1715);
not NOT1 (N1737, N1734);
nand NAND4 (N1738, N1730, N1669, N622, N1402);
or OR2 (N1739, N1735, N506);
and AND4 (N1740, N1728, N1358, N797, N607);
nand NAND4 (N1741, N1737, N1738, N1467, N1073);
nand NAND3 (N1742, N1447, N832, N1423);
or OR2 (N1743, N1740, N1612);
and AND2 (N1744, N1742, N1495);
not NOT1 (N1745, N1731);
buf BUF1 (N1746, N1726);
not NOT1 (N1747, N1744);
xor XOR2 (N1748, N1743, N1483);
or OR2 (N1749, N1718, N1507);
nor NOR2 (N1750, N1749, N1613);
nand NAND2 (N1751, N1748, N568);
or OR3 (N1752, N1745, N467, N1427);
buf BUF1 (N1753, N1736);
nor NOR2 (N1754, N1752, N41);
and AND4 (N1755, N1733, N927, N214, N1157);
nor NOR4 (N1756, N1750, N945, N675, N167);
nor NOR2 (N1757, N1754, N1192);
xor XOR2 (N1758, N1747, N1273);
buf BUF1 (N1759, N1741);
not NOT1 (N1760, N1756);
and AND2 (N1761, N1753, N1496);
and AND4 (N1762, N1732, N77, N1095, N729);
not NOT1 (N1763, N1758);
and AND4 (N1764, N1739, N160, N569, N997);
nand NAND4 (N1765, N1755, N875, N1274, N1312);
not NOT1 (N1766, N1764);
not NOT1 (N1767, N1762);
not NOT1 (N1768, N1767);
nand NAND4 (N1769, N1759, N511, N1006, N288);
buf BUF1 (N1770, N1768);
nand NAND3 (N1771, N1766, N1670, N1064);
not NOT1 (N1772, N1761);
not NOT1 (N1773, N1765);
buf BUF1 (N1774, N1770);
and AND3 (N1775, N1751, N1367, N379);
nor NOR4 (N1776, N1772, N289, N1721, N1459);
nand NAND3 (N1777, N1757, N1647, N212);
or OR2 (N1778, N1746, N401);
or OR3 (N1779, N1774, N1285, N908);
xor XOR2 (N1780, N1779, N1200);
xor XOR2 (N1781, N1771, N1014);
and AND2 (N1782, N1777, N227);
xor XOR2 (N1783, N1781, N1183);
nor NOR3 (N1784, N1780, N485, N1623);
not NOT1 (N1785, N1760);
xor XOR2 (N1786, N1763, N1751);
not NOT1 (N1787, N1778);
and AND4 (N1788, N1776, N49, N928, N780);
or OR3 (N1789, N1784, N267, N23);
or OR3 (N1790, N1775, N59, N259);
or OR4 (N1791, N1788, N1285, N1449, N1556);
nand NAND4 (N1792, N1790, N1175, N959, N225);
and AND3 (N1793, N1792, N532, N896);
nor NOR4 (N1794, N1789, N1466, N879, N653);
nand NAND2 (N1795, N1794, N1039);
nand NAND2 (N1796, N1782, N1492);
and AND4 (N1797, N1791, N1623, N794, N12);
not NOT1 (N1798, N1785);
not NOT1 (N1799, N1773);
or OR4 (N1800, N1799, N1429, N863, N1770);
and AND2 (N1801, N1795, N1547);
buf BUF1 (N1802, N1783);
or OR3 (N1803, N1797, N1277, N1127);
and AND3 (N1804, N1796, N1000, N1127);
xor XOR2 (N1805, N1793, N889);
or OR2 (N1806, N1786, N1520);
or OR2 (N1807, N1800, N1805);
nand NAND3 (N1808, N1497, N1188, N432);
or OR4 (N1809, N1787, N1398, N1302, N559);
or OR2 (N1810, N1809, N1693);
buf BUF1 (N1811, N1769);
and AND3 (N1812, N1803, N994, N1135);
nor NOR3 (N1813, N1806, N881, N1641);
not NOT1 (N1814, N1798);
buf BUF1 (N1815, N1808);
nor NOR2 (N1816, N1812, N1027);
not NOT1 (N1817, N1816);
or OR4 (N1818, N1810, N1246, N505, N1476);
nand NAND4 (N1819, N1801, N1069, N1406, N1436);
and AND2 (N1820, N1813, N1109);
or OR4 (N1821, N1815, N316, N1599, N69);
nor NOR4 (N1822, N1818, N541, N487, N920);
or OR3 (N1823, N1811, N504, N141);
nor NOR4 (N1824, N1802, N1359, N1047, N1283);
nand NAND2 (N1825, N1821, N326);
xor XOR2 (N1826, N1817, N1117);
nor NOR3 (N1827, N1823, N1776, N145);
not NOT1 (N1828, N1826);
buf BUF1 (N1829, N1804);
nand NAND3 (N1830, N1822, N93, N1487);
and AND4 (N1831, N1814, N1743, N116, N1267);
and AND2 (N1832, N1825, N1549);
or OR4 (N1833, N1827, N1133, N1282, N1450);
not NOT1 (N1834, N1829);
or OR3 (N1835, N1833, N1063, N543);
and AND3 (N1836, N1824, N1055, N70);
or OR4 (N1837, N1820, N778, N1047, N95);
not NOT1 (N1838, N1807);
nand NAND2 (N1839, N1832, N144);
buf BUF1 (N1840, N1830);
or OR3 (N1841, N1828, N49, N1547);
not NOT1 (N1842, N1819);
not NOT1 (N1843, N1836);
buf BUF1 (N1844, N1838);
nor NOR2 (N1845, N1841, N1306);
nand NAND4 (N1846, N1834, N1615, N564, N476);
xor XOR2 (N1847, N1842, N1023);
and AND3 (N1848, N1847, N1439, N1786);
buf BUF1 (N1849, N1837);
not NOT1 (N1850, N1840);
not NOT1 (N1851, N1848);
not NOT1 (N1852, N1849);
or OR4 (N1853, N1844, N1274, N353, N1068);
xor XOR2 (N1854, N1835, N1415);
and AND2 (N1855, N1850, N966);
buf BUF1 (N1856, N1846);
nand NAND4 (N1857, N1839, N938, N585, N847);
and AND3 (N1858, N1845, N1720, N636);
and AND2 (N1859, N1855, N1024);
buf BUF1 (N1860, N1852);
nand NAND2 (N1861, N1857, N357);
xor XOR2 (N1862, N1831, N1650);
buf BUF1 (N1863, N1856);
not NOT1 (N1864, N1863);
or OR4 (N1865, N1860, N418, N724, N1855);
and AND2 (N1866, N1859, N384);
not NOT1 (N1867, N1862);
buf BUF1 (N1868, N1851);
or OR3 (N1869, N1864, N1725, N1305);
nor NOR2 (N1870, N1843, N1575);
xor XOR2 (N1871, N1869, N1332);
and AND2 (N1872, N1858, N1773);
or OR2 (N1873, N1870, N1858);
xor XOR2 (N1874, N1854, N67);
nand NAND2 (N1875, N1865, N659);
nor NOR3 (N1876, N1873, N1031, N1511);
buf BUF1 (N1877, N1876);
xor XOR2 (N1878, N1853, N142);
or OR2 (N1879, N1867, N824);
or OR4 (N1880, N1868, N388, N1232, N664);
nand NAND4 (N1881, N1880, N1148, N820, N1136);
buf BUF1 (N1882, N1866);
or OR2 (N1883, N1861, N44);
nand NAND3 (N1884, N1882, N944, N1572);
buf BUF1 (N1885, N1878);
and AND2 (N1886, N1872, N1568);
xor XOR2 (N1887, N1886, N267);
nor NOR4 (N1888, N1884, N77, N835, N1828);
and AND2 (N1889, N1881, N272);
xor XOR2 (N1890, N1885, N1317);
not NOT1 (N1891, N1889);
not NOT1 (N1892, N1874);
xor XOR2 (N1893, N1875, N469);
or OR4 (N1894, N1890, N190, N791, N41);
and AND3 (N1895, N1877, N1636, N452);
or OR2 (N1896, N1893, N1837);
not NOT1 (N1897, N1894);
or OR2 (N1898, N1879, N272);
nand NAND2 (N1899, N1891, N1472);
not NOT1 (N1900, N1897);
or OR4 (N1901, N1898, N1680, N1399, N1230);
not NOT1 (N1902, N1901);
xor XOR2 (N1903, N1896, N808);
buf BUF1 (N1904, N1883);
nand NAND2 (N1905, N1899, N809);
nand NAND4 (N1906, N1904, N700, N1425, N633);
nor NOR3 (N1907, N1895, N366, N1280);
buf BUF1 (N1908, N1892);
nor NOR2 (N1909, N1900, N1484);
or OR4 (N1910, N1888, N268, N1007, N1144);
and AND2 (N1911, N1909, N457);
or OR4 (N1912, N1907, N1197, N160, N1066);
or OR3 (N1913, N1910, N574, N1809);
and AND4 (N1914, N1905, N1653, N691, N439);
and AND2 (N1915, N1911, N1583);
nand NAND2 (N1916, N1903, N217);
nand NAND2 (N1917, N1916, N1215);
and AND4 (N1918, N1914, N363, N802, N12);
xor XOR2 (N1919, N1912, N1359);
or OR3 (N1920, N1902, N1752, N67);
buf BUF1 (N1921, N1919);
and AND4 (N1922, N1913, N1390, N335, N55);
nand NAND2 (N1923, N1906, N1848);
nand NAND2 (N1924, N1908, N894);
or OR3 (N1925, N1915, N922, N1751);
nand NAND3 (N1926, N1923, N39, N74);
xor XOR2 (N1927, N1922, N1708);
buf BUF1 (N1928, N1926);
xor XOR2 (N1929, N1918, N1692);
nor NOR3 (N1930, N1928, N650, N213);
or OR3 (N1931, N1871, N213, N1349);
xor XOR2 (N1932, N1924, N656);
nand NAND3 (N1933, N1887, N1627, N1138);
not NOT1 (N1934, N1933);
not NOT1 (N1935, N1929);
nor NOR3 (N1936, N1932, N338, N29);
xor XOR2 (N1937, N1931, N937);
not NOT1 (N1938, N1921);
buf BUF1 (N1939, N1920);
xor XOR2 (N1940, N1939, N937);
xor XOR2 (N1941, N1930, N1658);
or OR3 (N1942, N1934, N1302, N1872);
nand NAND2 (N1943, N1936, N180);
buf BUF1 (N1944, N1935);
not NOT1 (N1945, N1938);
xor XOR2 (N1946, N1944, N613);
nor NOR2 (N1947, N1943, N659);
or OR4 (N1948, N1946, N1625, N505, N1831);
and AND3 (N1949, N1947, N458, N382);
xor XOR2 (N1950, N1925, N1702);
not NOT1 (N1951, N1948);
nor NOR4 (N1952, N1937, N1352, N745, N1543);
or OR3 (N1953, N1951, N610, N1665);
buf BUF1 (N1954, N1953);
buf BUF1 (N1955, N1950);
nor NOR2 (N1956, N1949, N403);
nor NOR2 (N1957, N1952, N1768);
not NOT1 (N1958, N1954);
buf BUF1 (N1959, N1945);
or OR3 (N1960, N1917, N629, N1285);
nand NAND3 (N1961, N1956, N284, N992);
or OR4 (N1962, N1927, N1217, N1202, N689);
xor XOR2 (N1963, N1958, N964);
nand NAND4 (N1964, N1960, N59, N873, N678);
and AND3 (N1965, N1963, N365, N1547);
xor XOR2 (N1966, N1957, N172);
buf BUF1 (N1967, N1961);
or OR4 (N1968, N1966, N933, N1003, N897);
nand NAND2 (N1969, N1942, N633);
or OR4 (N1970, N1967, N279, N616, N1379);
nor NOR4 (N1971, N1962, N1527, N1612, N358);
nand NAND3 (N1972, N1955, N1580, N1007);
buf BUF1 (N1973, N1959);
not NOT1 (N1974, N1970);
xor XOR2 (N1975, N1941, N777);
not NOT1 (N1976, N1972);
xor XOR2 (N1977, N1965, N371);
buf BUF1 (N1978, N1964);
nor NOR2 (N1979, N1968, N565);
or OR4 (N1980, N1971, N1764, N1546, N1146);
not NOT1 (N1981, N1974);
and AND2 (N1982, N1969, N252);
xor XOR2 (N1983, N1982, N134);
and AND4 (N1984, N1980, N1249, N674, N1693);
xor XOR2 (N1985, N1976, N1943);
not NOT1 (N1986, N1985);
nand NAND3 (N1987, N1977, N1762, N1222);
buf BUF1 (N1988, N1981);
xor XOR2 (N1989, N1940, N616);
nor NOR4 (N1990, N1984, N783, N661, N1871);
nor NOR4 (N1991, N1978, N1950, N1009, N258);
nor NOR4 (N1992, N1990, N1349, N1638, N1440);
nor NOR2 (N1993, N1987, N1500);
buf BUF1 (N1994, N1991);
not NOT1 (N1995, N1988);
not NOT1 (N1996, N1994);
or OR2 (N1997, N1995, N275);
buf BUF1 (N1998, N1975);
buf BUF1 (N1999, N1992);
or OR2 (N2000, N1989, N1918);
nor NOR3 (N2001, N1986, N1985, N1409);
buf BUF1 (N2002, N1979);
not NOT1 (N2003, N2000);
xor XOR2 (N2004, N1993, N1028);
xor XOR2 (N2005, N1973, N1732);
buf BUF1 (N2006, N2001);
buf BUF1 (N2007, N1999);
xor XOR2 (N2008, N1997, N1066);
nor NOR2 (N2009, N1998, N1596);
or OR4 (N2010, N2009, N1670, N1906, N441);
nor NOR3 (N2011, N2003, N1686, N1280);
nand NAND2 (N2012, N1983, N351);
and AND4 (N2013, N2006, N751, N1859, N939);
or OR2 (N2014, N2013, N633);
xor XOR2 (N2015, N2004, N942);
not NOT1 (N2016, N2015);
and AND2 (N2017, N2008, N1077);
nand NAND3 (N2018, N2011, N1440, N931);
buf BUF1 (N2019, N2005);
nor NOR4 (N2020, N2016, N1292, N1347, N1672);
or OR4 (N2021, N2012, N451, N1692, N1173);
not NOT1 (N2022, N2020);
nand NAND2 (N2023, N2022, N1331);
not NOT1 (N2024, N2019);
buf BUF1 (N2025, N2010);
nand NAND4 (N2026, N2007, N190, N253, N444);
or OR3 (N2027, N2021, N709, N481);
nor NOR3 (N2028, N2024, N839, N875);
nor NOR4 (N2029, N2027, N1992, N82, N521);
nor NOR4 (N2030, N2023, N625, N1176, N1375);
nor NOR3 (N2031, N2014, N671, N1969);
buf BUF1 (N2032, N2002);
and AND4 (N2033, N2029, N369, N447, N596);
nor NOR2 (N2034, N2017, N1905);
nor NOR4 (N2035, N2033, N1874, N1565, N260);
not NOT1 (N2036, N2028);
xor XOR2 (N2037, N2031, N1869);
not NOT1 (N2038, N2025);
nand NAND4 (N2039, N2034, N397, N2014, N281);
or OR3 (N2040, N2018, N1269, N1494);
not NOT1 (N2041, N2026);
or OR3 (N2042, N2030, N975, N473);
nand NAND2 (N2043, N2035, N176);
or OR2 (N2044, N2041, N797);
nor NOR3 (N2045, N2044, N422, N1963);
nand NAND4 (N2046, N2042, N1564, N862, N1125);
and AND2 (N2047, N2039, N1864);
not NOT1 (N2048, N2037);
nor NOR3 (N2049, N2036, N631, N1981);
nor NOR4 (N2050, N2047, N327, N1405, N1277);
not NOT1 (N2051, N2048);
not NOT1 (N2052, N2050);
and AND2 (N2053, N2043, N112);
xor XOR2 (N2054, N2046, N1872);
xor XOR2 (N2055, N2032, N826);
nor NOR2 (N2056, N2055, N1504);
nor NOR3 (N2057, N2056, N1203, N1818);
nor NOR2 (N2058, N2053, N2032);
nand NAND2 (N2059, N2051, N116);
buf BUF1 (N2060, N2038);
not NOT1 (N2061, N2054);
not NOT1 (N2062, N2059);
not NOT1 (N2063, N2049);
nand NAND3 (N2064, N2040, N62, N1183);
nor NOR2 (N2065, N2063, N1672);
buf BUF1 (N2066, N1996);
and AND4 (N2067, N2045, N1596, N806, N1557);
nor NOR3 (N2068, N2052, N710, N1954);
buf BUF1 (N2069, N2066);
nor NOR2 (N2070, N2065, N307);
and AND4 (N2071, N2062, N1437, N1204, N1048);
buf BUF1 (N2072, N2058);
buf BUF1 (N2073, N2060);
nor NOR4 (N2074, N2067, N296, N67, N563);
buf BUF1 (N2075, N2057);
nand NAND2 (N2076, N2070, N1996);
and AND3 (N2077, N2061, N1873, N910);
buf BUF1 (N2078, N2072);
xor XOR2 (N2079, N2073, N1811);
and AND2 (N2080, N2078, N1300);
buf BUF1 (N2081, N2077);
nand NAND2 (N2082, N2076, N1423);
not NOT1 (N2083, N2069);
not NOT1 (N2084, N2071);
and AND2 (N2085, N2079, N1249);
nor NOR4 (N2086, N2075, N826, N1598, N1677);
buf BUF1 (N2087, N2080);
buf BUF1 (N2088, N2083);
buf BUF1 (N2089, N2068);
not NOT1 (N2090, N2064);
nor NOR3 (N2091, N2074, N1812, N260);
or OR4 (N2092, N2084, N1642, N871, N339);
or OR3 (N2093, N2088, N1750, N2037);
xor XOR2 (N2094, N2093, N1167);
xor XOR2 (N2095, N2086, N683);
nand NAND3 (N2096, N2081, N737, N1957);
nand NAND2 (N2097, N2096, N1427);
xor XOR2 (N2098, N2091, N1508);
or OR2 (N2099, N2082, N216);
or OR2 (N2100, N2098, N1831);
or OR4 (N2101, N2085, N1332, N567, N875);
and AND3 (N2102, N2101, N1116, N925);
or OR3 (N2103, N2089, N735, N625);
not NOT1 (N2104, N2095);
not NOT1 (N2105, N2099);
nand NAND2 (N2106, N2105, N1527);
xor XOR2 (N2107, N2097, N625);
buf BUF1 (N2108, N2094);
buf BUF1 (N2109, N2104);
buf BUF1 (N2110, N2087);
and AND3 (N2111, N2109, N1050, N2009);
nor NOR4 (N2112, N2103, N484, N1149, N759);
xor XOR2 (N2113, N2102, N126);
xor XOR2 (N2114, N2107, N1798);
or OR3 (N2115, N2110, N175, N1513);
buf BUF1 (N2116, N2113);
nand NAND3 (N2117, N2111, N1783, N2099);
or OR2 (N2118, N2106, N523);
and AND2 (N2119, N2112, N836);
nor NOR4 (N2120, N2108, N1036, N1087, N599);
and AND4 (N2121, N2118, N1746, N634, N1423);
nor NOR2 (N2122, N2121, N186);
or OR2 (N2123, N2115, N724);
nand NAND4 (N2124, N2120, N528, N1796, N1351);
nor NOR4 (N2125, N2119, N1513, N1349, N1341);
buf BUF1 (N2126, N2116);
not NOT1 (N2127, N2123);
not NOT1 (N2128, N2092);
nor NOR2 (N2129, N2114, N2019);
xor XOR2 (N2130, N2122, N1690);
and AND4 (N2131, N2128, N75, N1632, N1185);
buf BUF1 (N2132, N2129);
or OR3 (N2133, N2100, N794, N549);
buf BUF1 (N2134, N2127);
not NOT1 (N2135, N2117);
not NOT1 (N2136, N2090);
not NOT1 (N2137, N2132);
and AND2 (N2138, N2137, N1823);
or OR4 (N2139, N2138, N1595, N1572, N964);
xor XOR2 (N2140, N2125, N1734);
nand NAND3 (N2141, N2139, N1852, N929);
nand NAND2 (N2142, N2124, N1391);
or OR4 (N2143, N2136, N530, N1281, N70);
and AND2 (N2144, N2134, N902);
nor NOR3 (N2145, N2130, N1681, N45);
nor NOR4 (N2146, N2141, N1601, N889, N625);
nor NOR2 (N2147, N2126, N2134);
xor XOR2 (N2148, N2133, N1127);
nor NOR4 (N2149, N2145, N577, N1537, N128);
not NOT1 (N2150, N2143);
or OR2 (N2151, N2147, N414);
nor NOR2 (N2152, N2135, N51);
and AND4 (N2153, N2142, N1505, N163, N2141);
xor XOR2 (N2154, N2146, N364);
xor XOR2 (N2155, N2150, N349);
nor NOR3 (N2156, N2155, N753, N1597);
buf BUF1 (N2157, N2149);
buf BUF1 (N2158, N2144);
and AND4 (N2159, N2131, N1236, N1161, N1553);
and AND2 (N2160, N2148, N1926);
xor XOR2 (N2161, N2158, N680);
nor NOR4 (N2162, N2156, N142, N189, N75);
xor XOR2 (N2163, N2157, N485);
nor NOR4 (N2164, N2154, N205, N1459, N223);
nor NOR4 (N2165, N2151, N1687, N898, N1254);
nand NAND4 (N2166, N2165, N916, N1697, N1366);
nor NOR4 (N2167, N2159, N180, N999, N324);
nand NAND2 (N2168, N2140, N289);
nor NOR4 (N2169, N2162, N307, N108, N1311);
not NOT1 (N2170, N2169);
xor XOR2 (N2171, N2152, N910);
not NOT1 (N2172, N2168);
and AND3 (N2173, N2167, N329, N7);
nand NAND4 (N2174, N2173, N1727, N692, N736);
nand NAND4 (N2175, N2170, N1080, N1463, N1554);
nor NOR2 (N2176, N2153, N534);
and AND2 (N2177, N2164, N149);
and AND4 (N2178, N2172, N1518, N1640, N2166);
buf BUF1 (N2179, N602);
and AND3 (N2180, N2175, N1454, N537);
or OR4 (N2181, N2176, N2136, N1608, N1695);
xor XOR2 (N2182, N2177, N666);
buf BUF1 (N2183, N2160);
not NOT1 (N2184, N2183);
buf BUF1 (N2185, N2184);
not NOT1 (N2186, N2174);
not NOT1 (N2187, N2163);
or OR2 (N2188, N2181, N23);
buf BUF1 (N2189, N2179);
buf BUF1 (N2190, N2185);
not NOT1 (N2191, N2188);
nor NOR4 (N2192, N2171, N242, N1204, N310);
or OR4 (N2193, N2178, N405, N813, N1134);
nand NAND2 (N2194, N2186, N1780);
xor XOR2 (N2195, N2193, N1562);
nor NOR4 (N2196, N2180, N937, N1941, N1180);
nand NAND2 (N2197, N2192, N560);
xor XOR2 (N2198, N2189, N838);
and AND3 (N2199, N2197, N1007, N864);
xor XOR2 (N2200, N2191, N1008);
buf BUF1 (N2201, N2198);
not NOT1 (N2202, N2195);
not NOT1 (N2203, N2194);
buf BUF1 (N2204, N2187);
buf BUF1 (N2205, N2201);
not NOT1 (N2206, N2161);
buf BUF1 (N2207, N2206);
xor XOR2 (N2208, N2190, N1848);
not NOT1 (N2209, N2205);
xor XOR2 (N2210, N2207, N835);
and AND2 (N2211, N2200, N1250);
or OR4 (N2212, N2210, N1272, N1403, N423);
and AND3 (N2213, N2209, N1793, N315);
nor NOR4 (N2214, N2203, N1191, N1690, N1894);
xor XOR2 (N2215, N2213, N862);
not NOT1 (N2216, N2208);
xor XOR2 (N2217, N2215, N1781);
and AND2 (N2218, N2217, N572);
xor XOR2 (N2219, N2202, N28);
or OR2 (N2220, N2216, N285);
or OR3 (N2221, N2219, N1735, N1484);
not NOT1 (N2222, N2220);
xor XOR2 (N2223, N2196, N762);
xor XOR2 (N2224, N2222, N1355);
or OR2 (N2225, N2199, N1040);
buf BUF1 (N2226, N2182);
xor XOR2 (N2227, N2211, N678);
not NOT1 (N2228, N2204);
and AND2 (N2229, N2228, N400);
nand NAND2 (N2230, N2221, N727);
not NOT1 (N2231, N2227);
xor XOR2 (N2232, N2224, N1401);
nand NAND4 (N2233, N2212, N2002, N1066, N148);
buf BUF1 (N2234, N2229);
or OR2 (N2235, N2231, N162);
nand NAND4 (N2236, N2235, N36, N884, N470);
xor XOR2 (N2237, N2226, N2210);
nand NAND2 (N2238, N2236, N1271);
xor XOR2 (N2239, N2232, N1208);
nand NAND2 (N2240, N2238, N1505);
buf BUF1 (N2241, N2240);
and AND2 (N2242, N2230, N1584);
buf BUF1 (N2243, N2241);
and AND2 (N2244, N2234, N140);
buf BUF1 (N2245, N2225);
nand NAND4 (N2246, N2214, N1088, N1513, N1851);
not NOT1 (N2247, N2242);
buf BUF1 (N2248, N2223);
and AND2 (N2249, N2239, N1298);
nand NAND3 (N2250, N2246, N595, N1560);
nor NOR2 (N2251, N2237, N2223);
nor NOR3 (N2252, N2244, N1754, N310);
or OR3 (N2253, N2247, N1010, N903);
nor NOR3 (N2254, N2252, N1198, N1723);
xor XOR2 (N2255, N2250, N2168);
nor NOR4 (N2256, N2253, N594, N1500, N2243);
xor XOR2 (N2257, N1534, N2236);
and AND2 (N2258, N2257, N1978);
not NOT1 (N2259, N2258);
not NOT1 (N2260, N2259);
nor NOR3 (N2261, N2251, N2177, N329);
xor XOR2 (N2262, N2261, N1092);
or OR2 (N2263, N2255, N149);
nand NAND2 (N2264, N2254, N969);
or OR4 (N2265, N2260, N31, N736, N1154);
xor XOR2 (N2266, N2264, N1714);
xor XOR2 (N2267, N2249, N2216);
and AND2 (N2268, N2256, N412);
nand NAND2 (N2269, N2245, N984);
nor NOR3 (N2270, N2263, N1808, N128);
xor XOR2 (N2271, N2265, N2175);
and AND2 (N2272, N2269, N1534);
not NOT1 (N2273, N2233);
nor NOR3 (N2274, N2248, N346, N663);
nor NOR3 (N2275, N2271, N399, N739);
not NOT1 (N2276, N2272);
and AND2 (N2277, N2275, N634);
and AND4 (N2278, N2262, N2207, N234, N1319);
xor XOR2 (N2279, N2277, N2102);
not NOT1 (N2280, N2267);
not NOT1 (N2281, N2273);
nor NOR4 (N2282, N2266, N1457, N445, N1931);
buf BUF1 (N2283, N2274);
xor XOR2 (N2284, N2280, N1777);
xor XOR2 (N2285, N2276, N1740);
nor NOR2 (N2286, N2282, N2124);
not NOT1 (N2287, N2268);
xor XOR2 (N2288, N2278, N1978);
not NOT1 (N2289, N2286);
buf BUF1 (N2290, N2270);
not NOT1 (N2291, N2289);
nor NOR4 (N2292, N2285, N1239, N2054, N751);
nor NOR2 (N2293, N2290, N1913);
nand NAND2 (N2294, N2292, N2210);
not NOT1 (N2295, N2279);
buf BUF1 (N2296, N2284);
xor XOR2 (N2297, N2287, N358);
xor XOR2 (N2298, N2291, N411);
or OR2 (N2299, N2293, N2276);
buf BUF1 (N2300, N2294);
nor NOR3 (N2301, N2281, N842, N1679);
and AND3 (N2302, N2297, N142, N321);
xor XOR2 (N2303, N2299, N329);
buf BUF1 (N2304, N2295);
xor XOR2 (N2305, N2302, N1803);
not NOT1 (N2306, N2303);
and AND4 (N2307, N2218, N487, N59, N1155);
or OR3 (N2308, N2307, N519, N380);
nand NAND4 (N2309, N2296, N213, N1054, N1326);
and AND3 (N2310, N2298, N861, N855);
nand NAND3 (N2311, N2306, N2024, N2085);
nor NOR3 (N2312, N2310, N1106, N1197);
xor XOR2 (N2313, N2311, N1811);
or OR4 (N2314, N2308, N1068, N909, N597);
or OR4 (N2315, N2313, N995, N898, N2267);
and AND4 (N2316, N2314, N1648, N1898, N230);
not NOT1 (N2317, N2312);
buf BUF1 (N2318, N2301);
xor XOR2 (N2319, N2304, N350);
not NOT1 (N2320, N2315);
and AND4 (N2321, N2288, N833, N60, N1627);
xor XOR2 (N2322, N2300, N2161);
xor XOR2 (N2323, N2322, N1166);
buf BUF1 (N2324, N2319);
not NOT1 (N2325, N2324);
or OR4 (N2326, N2321, N421, N431, N876);
nand NAND2 (N2327, N2316, N2053);
xor XOR2 (N2328, N2309, N628);
and AND3 (N2329, N2325, N2267, N1417);
and AND2 (N2330, N2317, N724);
and AND4 (N2331, N2330, N917, N1575, N2153);
not NOT1 (N2332, N2329);
not NOT1 (N2333, N2327);
buf BUF1 (N2334, N2318);
or OR4 (N2335, N2331, N2248, N1812, N469);
nand NAND4 (N2336, N2326, N2161, N670, N832);
not NOT1 (N2337, N2283);
or OR3 (N2338, N2334, N2260, N1455);
and AND3 (N2339, N2328, N569, N367);
nand NAND4 (N2340, N2338, N631, N1525, N2052);
or OR2 (N2341, N2340, N544);
or OR2 (N2342, N2305, N93);
or OR4 (N2343, N2341, N857, N1812, N150);
and AND3 (N2344, N2339, N2010, N487);
and AND2 (N2345, N2333, N1574);
and AND4 (N2346, N2332, N1077, N2138, N892);
not NOT1 (N2347, N2342);
nor NOR4 (N2348, N2347, N427, N1335, N1868);
nor NOR2 (N2349, N2346, N617);
buf BUF1 (N2350, N2345);
not NOT1 (N2351, N2348);
nand NAND3 (N2352, N2350, N1513, N2004);
nand NAND2 (N2353, N2336, N1447);
and AND4 (N2354, N2352, N289, N1641, N1153);
and AND2 (N2355, N2337, N2132);
buf BUF1 (N2356, N2323);
nand NAND2 (N2357, N2344, N1251);
xor XOR2 (N2358, N2351, N708);
nand NAND3 (N2359, N2349, N2024, N412);
or OR2 (N2360, N2356, N2044);
xor XOR2 (N2361, N2359, N1494);
or OR4 (N2362, N2335, N1345, N721, N973);
or OR4 (N2363, N2320, N334, N790, N91);
nor NOR3 (N2364, N2363, N2204, N53);
not NOT1 (N2365, N2358);
xor XOR2 (N2366, N2360, N2271);
xor XOR2 (N2367, N2353, N710);
or OR3 (N2368, N2365, N1087, N196);
not NOT1 (N2369, N2364);
nor NOR3 (N2370, N2369, N800, N625);
or OR2 (N2371, N2367, N2311);
and AND2 (N2372, N2361, N959);
and AND3 (N2373, N2362, N2213, N208);
nor NOR2 (N2374, N2354, N389);
nor NOR2 (N2375, N2368, N1354);
nor NOR2 (N2376, N2373, N275);
buf BUF1 (N2377, N2376);
or OR3 (N2378, N2355, N1643, N1513);
nor NOR3 (N2379, N2343, N1213, N1979);
nand NAND3 (N2380, N2366, N660, N1279);
nand NAND2 (N2381, N2374, N1893);
buf BUF1 (N2382, N2357);
buf BUF1 (N2383, N2382);
nor NOR4 (N2384, N2370, N510, N543, N2061);
xor XOR2 (N2385, N2377, N1998);
xor XOR2 (N2386, N2379, N1627);
not NOT1 (N2387, N2380);
xor XOR2 (N2388, N2372, N1893);
nand NAND4 (N2389, N2385, N692, N1871, N526);
buf BUF1 (N2390, N2386);
not NOT1 (N2391, N2390);
or OR4 (N2392, N2375, N1046, N57, N767);
nor NOR2 (N2393, N2387, N616);
and AND2 (N2394, N2384, N2108);
xor XOR2 (N2395, N2394, N1363);
xor XOR2 (N2396, N2392, N1485);
xor XOR2 (N2397, N2383, N1500);
xor XOR2 (N2398, N2393, N793);
and AND2 (N2399, N2391, N309);
not NOT1 (N2400, N2371);
xor XOR2 (N2401, N2395, N1933);
nor NOR4 (N2402, N2400, N919, N2237, N84);
and AND2 (N2403, N2401, N1637);
nor NOR3 (N2404, N2389, N1309, N1418);
and AND4 (N2405, N2378, N1237, N518, N1593);
or OR4 (N2406, N2396, N564, N1422, N947);
or OR3 (N2407, N2404, N1711, N468);
not NOT1 (N2408, N2403);
nor NOR2 (N2409, N2406, N1755);
nand NAND4 (N2410, N2397, N1959, N1715, N117);
buf BUF1 (N2411, N2405);
xor XOR2 (N2412, N2399, N88);
or OR4 (N2413, N2398, N1111, N324, N536);
buf BUF1 (N2414, N2388);
nand NAND3 (N2415, N2413, N1738, N1509);
xor XOR2 (N2416, N2414, N170);
not NOT1 (N2417, N2416);
nor NOR2 (N2418, N2410, N1675);
or OR2 (N2419, N2402, N914);
or OR4 (N2420, N2415, N656, N739, N976);
buf BUF1 (N2421, N2407);
nor NOR3 (N2422, N2418, N1368, N1081);
and AND2 (N2423, N2419, N978);
nor NOR3 (N2424, N2420, N2127, N992);
and AND2 (N2425, N2409, N1887);
and AND3 (N2426, N2423, N906, N2315);
xor XOR2 (N2427, N2426, N1441);
not NOT1 (N2428, N2425);
not NOT1 (N2429, N2412);
not NOT1 (N2430, N2429);
buf BUF1 (N2431, N2408);
not NOT1 (N2432, N2381);
nor NOR3 (N2433, N2422, N1309, N2406);
buf BUF1 (N2434, N2430);
and AND4 (N2435, N2427, N1422, N139, N485);
xor XOR2 (N2436, N2411, N1200);
or OR3 (N2437, N2436, N52, N1001);
nor NOR3 (N2438, N2433, N123, N1833);
not NOT1 (N2439, N2424);
xor XOR2 (N2440, N2434, N558);
not NOT1 (N2441, N2440);
not NOT1 (N2442, N2417);
not NOT1 (N2443, N2435);
and AND3 (N2444, N2438, N203, N317);
xor XOR2 (N2445, N2444, N1008);
or OR3 (N2446, N2441, N1470, N745);
nor NOR3 (N2447, N2432, N946, N2013);
not NOT1 (N2448, N2445);
and AND4 (N2449, N2447, N1011, N600, N220);
not NOT1 (N2450, N2431);
buf BUF1 (N2451, N2442);
not NOT1 (N2452, N2428);
nand NAND4 (N2453, N2421, N308, N1446, N1474);
xor XOR2 (N2454, N2452, N517);
xor XOR2 (N2455, N2451, N558);
or OR4 (N2456, N2439, N1165, N1928, N1172);
nand NAND3 (N2457, N2454, N1205, N2370);
nand NAND3 (N2458, N2446, N1710, N1138);
not NOT1 (N2459, N2448);
and AND2 (N2460, N2458, N897);
xor XOR2 (N2461, N2457, N1426);
nor NOR3 (N2462, N2450, N704, N1019);
buf BUF1 (N2463, N2459);
buf BUF1 (N2464, N2453);
not NOT1 (N2465, N2443);
nand NAND2 (N2466, N2465, N1230);
buf BUF1 (N2467, N2437);
xor XOR2 (N2468, N2467, N2150);
nand NAND3 (N2469, N2468, N1300, N2283);
not NOT1 (N2470, N2456);
not NOT1 (N2471, N2466);
not NOT1 (N2472, N2469);
nand NAND4 (N2473, N2470, N1028, N985, N1168);
and AND4 (N2474, N2472, N2383, N410, N848);
xor XOR2 (N2475, N2449, N1272);
nor NOR2 (N2476, N2474, N2379);
or OR4 (N2477, N2461, N1939, N896, N1447);
and AND2 (N2478, N2462, N52);
or OR3 (N2479, N2478, N1810, N1909);
and AND2 (N2480, N2464, N940);
xor XOR2 (N2481, N2479, N2241);
nand NAND3 (N2482, N2455, N1000, N414);
nor NOR4 (N2483, N2460, N514, N1151, N521);
nand NAND2 (N2484, N2481, N2212);
xor XOR2 (N2485, N2476, N398);
xor XOR2 (N2486, N2482, N1227);
not NOT1 (N2487, N2483);
buf BUF1 (N2488, N2477);
and AND2 (N2489, N2471, N788);
and AND3 (N2490, N2463, N1706, N1643);
xor XOR2 (N2491, N2480, N2387);
or OR2 (N2492, N2488, N2046);
not NOT1 (N2493, N2475);
or OR2 (N2494, N2489, N2062);
nand NAND3 (N2495, N2490, N2408, N326);
nand NAND3 (N2496, N2484, N2348, N1063);
nand NAND2 (N2497, N2491, N1933);
and AND3 (N2498, N2493, N372, N286);
not NOT1 (N2499, N2492);
buf BUF1 (N2500, N2495);
or OR3 (N2501, N2496, N1182, N595);
nand NAND3 (N2502, N2500, N247, N1590);
or OR3 (N2503, N2497, N427, N1359);
or OR2 (N2504, N2487, N1437);
or OR4 (N2505, N2504, N1733, N2208, N952);
buf BUF1 (N2506, N2485);
and AND3 (N2507, N2486, N177, N466);
buf BUF1 (N2508, N2498);
or OR4 (N2509, N2499, N88, N1445, N2411);
xor XOR2 (N2510, N2501, N1425);
nand NAND3 (N2511, N2506, N1153, N2027);
xor XOR2 (N2512, N2508, N637);
xor XOR2 (N2513, N2507, N216);
xor XOR2 (N2514, N2505, N2220);
and AND4 (N2515, N2511, N1154, N513, N1684);
nor NOR2 (N2516, N2514, N1893);
not NOT1 (N2517, N2513);
nand NAND2 (N2518, N2502, N1726);
or OR4 (N2519, N2518, N2193, N2050, N1841);
or OR4 (N2520, N2494, N1704, N863, N990);
nor NOR2 (N2521, N2473, N452);
not NOT1 (N2522, N2512);
xor XOR2 (N2523, N2515, N409);
or OR4 (N2524, N2517, N81, N1570, N1330);
buf BUF1 (N2525, N2520);
nor NOR2 (N2526, N2503, N771);
buf BUF1 (N2527, N2519);
not NOT1 (N2528, N2523);
nand NAND2 (N2529, N2516, N1089);
or OR3 (N2530, N2528, N641, N2178);
xor XOR2 (N2531, N2526, N2513);
or OR3 (N2532, N2521, N1372, N647);
and AND4 (N2533, N2530, N2187, N1329, N564);
and AND3 (N2534, N2522, N1757, N1261);
xor XOR2 (N2535, N2510, N985);
buf BUF1 (N2536, N2527);
or OR4 (N2537, N2531, N218, N2203, N2433);
not NOT1 (N2538, N2535);
buf BUF1 (N2539, N2532);
and AND2 (N2540, N2534, N915);
not NOT1 (N2541, N2538);
nand NAND2 (N2542, N2539, N801);
or OR2 (N2543, N2509, N1098);
not NOT1 (N2544, N2537);
buf BUF1 (N2545, N2529);
or OR4 (N2546, N2533, N1496, N683, N1796);
xor XOR2 (N2547, N2544, N328);
not NOT1 (N2548, N2524);
nor NOR3 (N2549, N2547, N2200, N1481);
and AND2 (N2550, N2541, N1996);
or OR3 (N2551, N2542, N1624, N2091);
or OR3 (N2552, N2545, N1797, N718);
nand NAND3 (N2553, N2551, N169, N708);
or OR4 (N2554, N2550, N2342, N313, N1557);
not NOT1 (N2555, N2553);
nor NOR4 (N2556, N2555, N2435, N574, N2007);
not NOT1 (N2557, N2552);
buf BUF1 (N2558, N2546);
nand NAND4 (N2559, N2549, N1434, N395, N1513);
not NOT1 (N2560, N2554);
and AND3 (N2561, N2560, N93, N248);
or OR3 (N2562, N2557, N1286, N669);
and AND4 (N2563, N2548, N1111, N1112, N872);
and AND2 (N2564, N2536, N1911);
nor NOR3 (N2565, N2525, N1181, N341);
buf BUF1 (N2566, N2558);
not NOT1 (N2567, N2562);
nor NOR2 (N2568, N2561, N1487);
or OR3 (N2569, N2564, N367, N1415);
or OR4 (N2570, N2569, N1040, N2546, N1404);
xor XOR2 (N2571, N2540, N1373);
xor XOR2 (N2572, N2568, N1010);
and AND2 (N2573, N2566, N351);
xor XOR2 (N2574, N2563, N1943);
or OR3 (N2575, N2574, N2030, N765);
or OR2 (N2576, N2570, N1846);
nand NAND2 (N2577, N2573, N1770);
nor NOR4 (N2578, N2576, N644, N1513, N227);
nand NAND2 (N2579, N2556, N2465);
nand NAND4 (N2580, N2571, N2579, N1825, N664);
buf BUF1 (N2581, N934);
nor NOR3 (N2582, N2567, N1628, N2163);
xor XOR2 (N2583, N2565, N2155);
and AND2 (N2584, N2580, N29);
or OR3 (N2585, N2577, N32, N922);
and AND4 (N2586, N2572, N516, N1052, N1292);
xor XOR2 (N2587, N2586, N2272);
nand NAND2 (N2588, N2578, N42);
nand NAND2 (N2589, N2581, N2271);
buf BUF1 (N2590, N2584);
and AND4 (N2591, N2588, N1522, N1301, N2276);
and AND3 (N2592, N2543, N1454, N296);
and AND2 (N2593, N2589, N499);
nor NOR4 (N2594, N2585, N1133, N725, N2593);
not NOT1 (N2595, N488);
xor XOR2 (N2596, N2582, N1222);
buf BUF1 (N2597, N2583);
nor NOR4 (N2598, N2595, N914, N394, N1267);
xor XOR2 (N2599, N2591, N779);
xor XOR2 (N2600, N2559, N703);
buf BUF1 (N2601, N2596);
nand NAND2 (N2602, N2599, N1452);
and AND2 (N2603, N2600, N1794);
xor XOR2 (N2604, N2603, N33);
xor XOR2 (N2605, N2604, N625);
buf BUF1 (N2606, N2601);
buf BUF1 (N2607, N2587);
and AND2 (N2608, N2590, N972);
xor XOR2 (N2609, N2607, N695);
buf BUF1 (N2610, N2609);
buf BUF1 (N2611, N2594);
xor XOR2 (N2612, N2605, N194);
buf BUF1 (N2613, N2611);
xor XOR2 (N2614, N2606, N2261);
or OR2 (N2615, N2608, N617);
xor XOR2 (N2616, N2597, N506);
nor NOR2 (N2617, N2602, N1457);
buf BUF1 (N2618, N2598);
nand NAND3 (N2619, N2592, N112, N1098);
xor XOR2 (N2620, N2575, N648);
and AND2 (N2621, N2616, N1038);
or OR2 (N2622, N2617, N1432);
nor NOR3 (N2623, N2610, N1747, N1689);
nor NOR3 (N2624, N2613, N1593, N1136);
nand NAND2 (N2625, N2623, N1637);
and AND3 (N2626, N2619, N1019, N694);
not NOT1 (N2627, N2626);
nand NAND4 (N2628, N2625, N580, N1056, N2163);
nand NAND4 (N2629, N2614, N2180, N1108, N967);
and AND3 (N2630, N2612, N1606, N1207);
nand NAND2 (N2631, N2621, N545);
nand NAND3 (N2632, N2615, N318, N2341);
not NOT1 (N2633, N2628);
buf BUF1 (N2634, N2620);
not NOT1 (N2635, N2622);
buf BUF1 (N2636, N2627);
xor XOR2 (N2637, N2632, N740);
not NOT1 (N2638, N2631);
buf BUF1 (N2639, N2636);
xor XOR2 (N2640, N2635, N2484);
xor XOR2 (N2641, N2638, N2300);
not NOT1 (N2642, N2629);
not NOT1 (N2643, N2624);
buf BUF1 (N2644, N2640);
xor XOR2 (N2645, N2644, N279);
not NOT1 (N2646, N2630);
or OR2 (N2647, N2642, N2455);
nand NAND3 (N2648, N2643, N1271, N2526);
nor NOR3 (N2649, N2634, N1465, N832);
xor XOR2 (N2650, N2645, N1232);
nand NAND3 (N2651, N2650, N1472, N2424);
nand NAND3 (N2652, N2648, N2136, N1113);
or OR4 (N2653, N2646, N2036, N1574, N22);
nor NOR4 (N2654, N2653, N1444, N2127, N1753);
xor XOR2 (N2655, N2639, N439);
or OR3 (N2656, N2655, N1887, N92);
buf BUF1 (N2657, N2637);
not NOT1 (N2658, N2649);
not NOT1 (N2659, N2618);
not NOT1 (N2660, N2651);
buf BUF1 (N2661, N2660);
not NOT1 (N2662, N2661);
and AND3 (N2663, N2652, N2387, N1088);
and AND2 (N2664, N2633, N2291);
or OR4 (N2665, N2658, N1714, N2023, N2373);
nor NOR2 (N2666, N2647, N1500);
or OR3 (N2667, N2659, N814, N534);
buf BUF1 (N2668, N2641);
buf BUF1 (N2669, N2668);
nand NAND4 (N2670, N2654, N1693, N2255, N1467);
not NOT1 (N2671, N2669);
buf BUF1 (N2672, N2667);
nand NAND3 (N2673, N2657, N2564, N2310);
xor XOR2 (N2674, N2665, N2418);
xor XOR2 (N2675, N2672, N503);
buf BUF1 (N2676, N2666);
or OR3 (N2677, N2673, N968, N243);
xor XOR2 (N2678, N2677, N2156);
or OR3 (N2679, N2676, N710, N1018);
xor XOR2 (N2680, N2675, N1287);
xor XOR2 (N2681, N2674, N1497);
buf BUF1 (N2682, N2681);
nand NAND2 (N2683, N2678, N2256);
nand NAND3 (N2684, N2682, N915, N1559);
nand NAND2 (N2685, N2670, N1604);
nand NAND3 (N2686, N2679, N609, N2431);
buf BUF1 (N2687, N2684);
not NOT1 (N2688, N2687);
and AND2 (N2689, N2671, N2169);
buf BUF1 (N2690, N2683);
and AND3 (N2691, N2690, N1816, N744);
nor NOR2 (N2692, N2663, N1046);
not NOT1 (N2693, N2656);
buf BUF1 (N2694, N2686);
nand NAND4 (N2695, N2680, N17, N912, N1672);
or OR2 (N2696, N2694, N1725);
or OR3 (N2697, N2692, N779, N2284);
buf BUF1 (N2698, N2689);
not NOT1 (N2699, N2693);
xor XOR2 (N2700, N2695, N2546);
xor XOR2 (N2701, N2662, N822);
xor XOR2 (N2702, N2698, N1872);
or OR2 (N2703, N2691, N1525);
nor NOR3 (N2704, N2664, N2654, N531);
or OR4 (N2705, N2696, N2446, N612, N2435);
nand NAND3 (N2706, N2688, N1799, N264);
nor NOR4 (N2707, N2700, N1461, N2455, N1486);
and AND4 (N2708, N2685, N1058, N1746, N1045);
and AND3 (N2709, N2699, N2260, N137);
buf BUF1 (N2710, N2702);
and AND4 (N2711, N2710, N2044, N1502, N2076);
nor NOR3 (N2712, N2704, N1000, N1349);
and AND3 (N2713, N2697, N120, N1377);
or OR3 (N2714, N2713, N1573, N1143);
xor XOR2 (N2715, N2708, N1559);
and AND2 (N2716, N2706, N1960);
buf BUF1 (N2717, N2716);
xor XOR2 (N2718, N2714, N59);
buf BUF1 (N2719, N2711);
and AND2 (N2720, N2703, N1868);
not NOT1 (N2721, N2720);
nor NOR4 (N2722, N2715, N1174, N1961, N2014);
xor XOR2 (N2723, N2719, N838);
not NOT1 (N2724, N2722);
buf BUF1 (N2725, N2724);
and AND4 (N2726, N2707, N1666, N1107, N323);
nor NOR4 (N2727, N2723, N2562, N1376, N1430);
and AND4 (N2728, N2725, N459, N2489, N639);
or OR3 (N2729, N2712, N261, N299);
and AND2 (N2730, N2721, N1842);
and AND2 (N2731, N2717, N2722);
or OR4 (N2732, N2727, N969, N1572, N138);
not NOT1 (N2733, N2732);
or OR2 (N2734, N2718, N47);
xor XOR2 (N2735, N2731, N1523);
and AND3 (N2736, N2735, N1132, N2195);
not NOT1 (N2737, N2733);
nand NAND2 (N2738, N2726, N528);
or OR3 (N2739, N2730, N2259, N1978);
not NOT1 (N2740, N2734);
or OR3 (N2741, N2709, N1193, N713);
nand NAND4 (N2742, N2705, N2330, N2655, N1458);
not NOT1 (N2743, N2742);
xor XOR2 (N2744, N2743, N1414);
not NOT1 (N2745, N2737);
not NOT1 (N2746, N2745);
xor XOR2 (N2747, N2740, N1853);
or OR3 (N2748, N2728, N126, N207);
buf BUF1 (N2749, N2738);
nor NOR2 (N2750, N2739, N1320);
and AND3 (N2751, N2748, N2013, N1538);
buf BUF1 (N2752, N2744);
nor NOR4 (N2753, N2736, N2348, N1248, N304);
not NOT1 (N2754, N2751);
xor XOR2 (N2755, N2741, N1227);
not NOT1 (N2756, N2749);
xor XOR2 (N2757, N2746, N2738);
buf BUF1 (N2758, N2757);
and AND3 (N2759, N2729, N554, N892);
and AND4 (N2760, N2747, N2619, N2357, N2513);
not NOT1 (N2761, N2754);
buf BUF1 (N2762, N2750);
xor XOR2 (N2763, N2752, N1415);
not NOT1 (N2764, N2756);
and AND2 (N2765, N2764, N211);
or OR4 (N2766, N2763, N1690, N2522, N2041);
nand NAND2 (N2767, N2753, N754);
nor NOR4 (N2768, N2766, N1833, N1324, N1383);
or OR2 (N2769, N2759, N594);
buf BUF1 (N2770, N2767);
nor NOR4 (N2771, N2770, N2699, N1099, N1922);
and AND4 (N2772, N2755, N41, N901, N446);
nor NOR4 (N2773, N2765, N1706, N280, N529);
not NOT1 (N2774, N2761);
buf BUF1 (N2775, N2771);
xor XOR2 (N2776, N2768, N1099);
or OR3 (N2777, N2775, N1096, N2683);
and AND4 (N2778, N2769, N2126, N896, N2277);
xor XOR2 (N2779, N2776, N1864);
nand NAND3 (N2780, N2774, N1087, N500);
not NOT1 (N2781, N2760);
buf BUF1 (N2782, N2779);
nand NAND3 (N2783, N2762, N2685, N78);
or OR3 (N2784, N2777, N625, N1841);
or OR4 (N2785, N2701, N854, N1253, N2493);
nor NOR2 (N2786, N2784, N2330);
or OR2 (N2787, N2786, N186);
and AND2 (N2788, N2778, N2592);
nor NOR4 (N2789, N2772, N2039, N2016, N1870);
nor NOR3 (N2790, N2781, N2167, N4);
or OR3 (N2791, N2790, N913, N823);
nand NAND3 (N2792, N2782, N2367, N2363);
not NOT1 (N2793, N2792);
nand NAND3 (N2794, N2783, N540, N1834);
xor XOR2 (N2795, N2780, N750);
nor NOR2 (N2796, N2794, N482);
or OR4 (N2797, N2793, N1147, N339, N1608);
xor XOR2 (N2798, N2796, N891);
or OR4 (N2799, N2758, N596, N1965, N13);
not NOT1 (N2800, N2773);
not NOT1 (N2801, N2785);
nand NAND2 (N2802, N2797, N412);
not NOT1 (N2803, N2799);
or OR2 (N2804, N2787, N1922);
nor NOR4 (N2805, N2795, N1165, N776, N2121);
nor NOR2 (N2806, N2791, N1152);
xor XOR2 (N2807, N2789, N1628);
nand NAND2 (N2808, N2801, N2032);
or OR2 (N2809, N2798, N1420);
nor NOR3 (N2810, N2806, N93, N878);
nand NAND3 (N2811, N2804, N663, N999);
buf BUF1 (N2812, N2807);
nor NOR3 (N2813, N2805, N795, N1154);
buf BUF1 (N2814, N2808);
not NOT1 (N2815, N2813);
nor NOR4 (N2816, N2800, N1032, N1193, N2005);
nand NAND3 (N2817, N2788, N1743, N1106);
or OR3 (N2818, N2812, N1051, N1438);
buf BUF1 (N2819, N2816);
nor NOR2 (N2820, N2817, N678);
or OR4 (N2821, N2809, N1229, N759, N1532);
xor XOR2 (N2822, N2802, N430);
or OR4 (N2823, N2819, N2320, N624, N2810);
buf BUF1 (N2824, N1666);
not NOT1 (N2825, N2803);
nor NOR3 (N2826, N2822, N349, N699);
buf BUF1 (N2827, N2824);
not NOT1 (N2828, N2815);
xor XOR2 (N2829, N2814, N304);
nor NOR3 (N2830, N2821, N2186, N856);
not NOT1 (N2831, N2818);
or OR4 (N2832, N2811, N1498, N1842, N1539);
buf BUF1 (N2833, N2831);
nor NOR2 (N2834, N2828, N2734);
buf BUF1 (N2835, N2826);
and AND2 (N2836, N2823, N2541);
or OR3 (N2837, N2834, N2263, N1055);
xor XOR2 (N2838, N2837, N534);
or OR4 (N2839, N2838, N585, N2459, N2833);
xor XOR2 (N2840, N536, N1738);
nor NOR3 (N2841, N2829, N1640, N2755);
nor NOR3 (N2842, N2830, N1928, N2053);
buf BUF1 (N2843, N2839);
or OR4 (N2844, N2843, N1600, N1487, N1062);
or OR4 (N2845, N2835, N1488, N1960, N532);
nand NAND2 (N2846, N2836, N1107);
xor XOR2 (N2847, N2832, N2816);
and AND2 (N2848, N2845, N640);
nor NOR2 (N2849, N2820, N547);
nand NAND4 (N2850, N2840, N2655, N646, N2839);
xor XOR2 (N2851, N2827, N1334);
buf BUF1 (N2852, N2848);
and AND3 (N2853, N2847, N2100, N114);
xor XOR2 (N2854, N2850, N2061);
or OR4 (N2855, N2851, N2581, N1429, N2171);
xor XOR2 (N2856, N2853, N1811);
not NOT1 (N2857, N2852);
not NOT1 (N2858, N2854);
xor XOR2 (N2859, N2856, N2039);
nor NOR3 (N2860, N2858, N1335, N2139);
buf BUF1 (N2861, N2849);
and AND2 (N2862, N2859, N2057);
buf BUF1 (N2863, N2857);
xor XOR2 (N2864, N2841, N1227);
nor NOR3 (N2865, N2864, N212, N1800);
xor XOR2 (N2866, N2825, N2220);
nor NOR3 (N2867, N2865, N1381, N1185);
xor XOR2 (N2868, N2867, N1144);
buf BUF1 (N2869, N2862);
and AND4 (N2870, N2860, N2742, N468, N1604);
nor NOR3 (N2871, N2868, N2416, N358);
nor NOR3 (N2872, N2866, N1858, N2165);
nor NOR4 (N2873, N2870, N176, N1331, N1567);
nand NAND2 (N2874, N2872, N368);
or OR3 (N2875, N2844, N1790, N1042);
nand NAND4 (N2876, N2874, N2772, N126, N953);
not NOT1 (N2877, N2855);
xor XOR2 (N2878, N2873, N1594);
xor XOR2 (N2879, N2869, N2407);
or OR2 (N2880, N2877, N271);
and AND2 (N2881, N2861, N707);
or OR2 (N2882, N2846, N2626);
not NOT1 (N2883, N2863);
not NOT1 (N2884, N2871);
nand NAND2 (N2885, N2879, N273);
and AND2 (N2886, N2880, N1340);
and AND4 (N2887, N2886, N2802, N1811, N2021);
and AND2 (N2888, N2842, N2762);
and AND3 (N2889, N2882, N2234, N2496);
not NOT1 (N2890, N2878);
or OR4 (N2891, N2890, N2322, N789, N2221);
xor XOR2 (N2892, N2887, N587);
nor NOR4 (N2893, N2876, N1368, N513, N778);
not NOT1 (N2894, N2884);
nor NOR2 (N2895, N2892, N542);
nand NAND2 (N2896, N2894, N1575);
nor NOR3 (N2897, N2896, N1173, N2393);
nor NOR4 (N2898, N2885, N1591, N1277, N1887);
xor XOR2 (N2899, N2897, N1791);
buf BUF1 (N2900, N2888);
buf BUF1 (N2901, N2883);
nor NOR4 (N2902, N2889, N1908, N1779, N1604);
xor XOR2 (N2903, N2900, N1413);
not NOT1 (N2904, N2901);
nor NOR4 (N2905, N2898, N2651, N1321, N2747);
nor NOR3 (N2906, N2902, N1158, N1271);
xor XOR2 (N2907, N2893, N2212);
nor NOR2 (N2908, N2903, N66);
xor XOR2 (N2909, N2895, N2696);
xor XOR2 (N2910, N2905, N1478);
or OR2 (N2911, N2875, N2556);
nor NOR4 (N2912, N2910, N1762, N2861, N2699);
not NOT1 (N2913, N2891);
nand NAND3 (N2914, N2904, N2389, N986);
nand NAND4 (N2915, N2907, N1178, N2773, N2712);
buf BUF1 (N2916, N2906);
not NOT1 (N2917, N2899);
buf BUF1 (N2918, N2908);
and AND3 (N2919, N2913, N1491, N311);
not NOT1 (N2920, N2881);
or OR3 (N2921, N2909, N152, N1340);
nor NOR2 (N2922, N2915, N2569);
nor NOR2 (N2923, N2912, N56);
and AND2 (N2924, N2919, N2826);
nand NAND2 (N2925, N2923, N1991);
nor NOR3 (N2926, N2921, N1878, N426);
nand NAND2 (N2927, N2914, N1356);
nor NOR3 (N2928, N2926, N2411, N1268);
or OR4 (N2929, N2920, N2066, N1050, N1540);
nor NOR4 (N2930, N2928, N787, N2825, N2813);
xor XOR2 (N2931, N2925, N572);
and AND2 (N2932, N2916, N1352);
or OR2 (N2933, N2924, N1380);
and AND2 (N2934, N2929, N365);
or OR4 (N2935, N2918, N1624, N2530, N2925);
xor XOR2 (N2936, N2934, N426);
or OR2 (N2937, N2933, N1052);
xor XOR2 (N2938, N2911, N2836);
and AND2 (N2939, N2922, N2005);
nand NAND2 (N2940, N2939, N418);
not NOT1 (N2941, N2932);
nand NAND3 (N2942, N2937, N1887, N1579);
nor NOR4 (N2943, N2941, N2024, N1750, N2755);
and AND4 (N2944, N2940, N2513, N1447, N2642);
nor NOR3 (N2945, N2927, N1162, N789);
xor XOR2 (N2946, N2930, N2069);
or OR4 (N2947, N2943, N207, N403, N1180);
not NOT1 (N2948, N2935);
and AND4 (N2949, N2936, N1228, N498, N325);
or OR3 (N2950, N2938, N2041, N1001);
or OR4 (N2951, N2917, N1088, N2280, N254);
nand NAND3 (N2952, N2948, N110, N2020);
xor XOR2 (N2953, N2949, N287);
nor NOR4 (N2954, N2931, N1862, N1949, N2647);
buf BUF1 (N2955, N2950);
and AND4 (N2956, N2952, N2875, N1072, N2306);
buf BUF1 (N2957, N2945);
and AND4 (N2958, N2957, N1861, N1214, N875);
nor NOR4 (N2959, N2946, N1953, N2770, N2116);
or OR4 (N2960, N2944, N1884, N2569, N2450);
nand NAND4 (N2961, N2942, N2062, N667, N1527);
and AND4 (N2962, N2953, N296, N823, N2434);
not NOT1 (N2963, N2962);
not NOT1 (N2964, N2947);
nand NAND3 (N2965, N2956, N437, N666);
buf BUF1 (N2966, N2955);
xor XOR2 (N2967, N2964, N1276);
nand NAND2 (N2968, N2966, N1155);
xor XOR2 (N2969, N2951, N2339);
xor XOR2 (N2970, N2954, N2820);
buf BUF1 (N2971, N2959);
and AND2 (N2972, N2969, N935);
nor NOR2 (N2973, N2960, N1517);
buf BUF1 (N2974, N2968);
nand NAND4 (N2975, N2961, N1586, N2224, N321);
nor NOR2 (N2976, N2974, N627);
nand NAND2 (N2977, N2976, N1598);
or OR3 (N2978, N2973, N2290, N1562);
xor XOR2 (N2979, N2972, N225);
nor NOR2 (N2980, N2965, N2896);
not NOT1 (N2981, N2975);
nor NOR2 (N2982, N2979, N1019);
xor XOR2 (N2983, N2970, N938);
buf BUF1 (N2984, N2967);
buf BUF1 (N2985, N2971);
buf BUF1 (N2986, N2980);
buf BUF1 (N2987, N2978);
and AND3 (N2988, N2958, N1411, N1470);
xor XOR2 (N2989, N2982, N524);
buf BUF1 (N2990, N2988);
not NOT1 (N2991, N2990);
and AND4 (N2992, N2963, N1109, N865, N976);
xor XOR2 (N2993, N2977, N138);
and AND2 (N2994, N2981, N2470);
nand NAND3 (N2995, N2993, N1858, N1479);
or OR2 (N2996, N2987, N2357);
and AND3 (N2997, N2983, N1137, N40);
nand NAND4 (N2998, N2984, N1896, N1722, N2880);
buf BUF1 (N2999, N2992);
nand NAND2 (N3000, N2986, N1809);
xor XOR2 (N3001, N2998, N245);
nand NAND2 (N3002, N2997, N736);
xor XOR2 (N3003, N3001, N1182);
xor XOR2 (N3004, N2985, N1759);
nor NOR2 (N3005, N2994, N2372);
nand NAND4 (N3006, N3002, N289, N1996, N532);
nand NAND4 (N3007, N3004, N2518, N559, N2852);
nor NOR2 (N3008, N2996, N322);
buf BUF1 (N3009, N3007);
nor NOR3 (N3010, N3006, N2086, N1095);
buf BUF1 (N3011, N2991);
or OR2 (N3012, N3000, N1665);
or OR4 (N3013, N2989, N2051, N2405, N1725);
xor XOR2 (N3014, N3011, N2755);
not NOT1 (N3015, N3008);
not NOT1 (N3016, N3009);
not NOT1 (N3017, N3005);
nand NAND3 (N3018, N3014, N2962, N1011);
not NOT1 (N3019, N3015);
and AND3 (N3020, N3003, N2284, N3006);
nor NOR4 (N3021, N3010, N947, N1473, N737);
xor XOR2 (N3022, N3018, N1834);
nand NAND3 (N3023, N2995, N2947, N2287);
buf BUF1 (N3024, N3016);
xor XOR2 (N3025, N3017, N367);
nor NOR3 (N3026, N3012, N1349, N2675);
not NOT1 (N3027, N3013);
nor NOR2 (N3028, N2999, N2845);
buf BUF1 (N3029, N3023);
nand NAND3 (N3030, N3021, N1103, N1315);
or OR3 (N3031, N3026, N2696, N2538);
xor XOR2 (N3032, N3025, N2705);
not NOT1 (N3033, N3022);
or OR4 (N3034, N3028, N1981, N1334, N946);
or OR4 (N3035, N3032, N3031, N98, N2440);
buf BUF1 (N3036, N2290);
buf BUF1 (N3037, N3030);
not NOT1 (N3038, N3034);
xor XOR2 (N3039, N3038, N1882);
nor NOR4 (N3040, N3036, N1731, N1468, N981);
not NOT1 (N3041, N3040);
xor XOR2 (N3042, N3019, N2277);
not NOT1 (N3043, N3020);
xor XOR2 (N3044, N3035, N2236);
nand NAND4 (N3045, N3027, N340, N2097, N2350);
buf BUF1 (N3046, N3024);
nand NAND2 (N3047, N3044, N1094);
or OR2 (N3048, N3033, N1586);
not NOT1 (N3049, N3041);
xor XOR2 (N3050, N3046, N1249);
not NOT1 (N3051, N3049);
or OR4 (N3052, N3051, N146, N588, N372);
nor NOR4 (N3053, N3029, N2941, N2530, N2104);
xor XOR2 (N3054, N3052, N1842);
xor XOR2 (N3055, N3047, N2123);
or OR4 (N3056, N3042, N3004, N1978, N2667);
nand NAND4 (N3057, N3045, N1911, N967, N1349);
nor NOR3 (N3058, N3056, N1575, N2923);
xor XOR2 (N3059, N3058, N1962);
buf BUF1 (N3060, N3057);
buf BUF1 (N3061, N3059);
nand NAND3 (N3062, N3055, N1849, N1053);
or OR4 (N3063, N3060, N1464, N622, N518);
not NOT1 (N3064, N3037);
or OR4 (N3065, N3061, N1512, N2362, N1679);
or OR4 (N3066, N3062, N319, N727, N1831);
and AND4 (N3067, N3065, N2086, N218, N2783);
nor NOR3 (N3068, N3067, N53, N695);
buf BUF1 (N3069, N3039);
or OR4 (N3070, N3054, N2965, N2307, N1362);
or OR2 (N3071, N3068, N1665);
and AND2 (N3072, N3063, N909);
buf BUF1 (N3073, N3048);
and AND2 (N3074, N3073, N508);
or OR3 (N3075, N3069, N1630, N1328);
not NOT1 (N3076, N3043);
or OR3 (N3077, N3070, N1605, N2059);
nor NOR2 (N3078, N3076, N3029);
nand NAND3 (N3079, N3074, N1251, N1296);
buf BUF1 (N3080, N3072);
buf BUF1 (N3081, N3053);
and AND4 (N3082, N3080, N1157, N771, N395);
and AND3 (N3083, N3064, N2062, N887);
nand NAND3 (N3084, N3050, N3044, N2487);
xor XOR2 (N3085, N3082, N686);
buf BUF1 (N3086, N3081);
nand NAND4 (N3087, N3079, N1612, N40, N1686);
nor NOR2 (N3088, N3071, N1260);
not NOT1 (N3089, N3086);
buf BUF1 (N3090, N3089);
not NOT1 (N3091, N3083);
nand NAND4 (N3092, N3078, N1242, N1311, N2395);
buf BUF1 (N3093, N3085);
xor XOR2 (N3094, N3077, N2470);
or OR2 (N3095, N3075, N520);
buf BUF1 (N3096, N3094);
and AND3 (N3097, N3090, N2022, N320);
nor NOR2 (N3098, N3088, N2923);
buf BUF1 (N3099, N3096);
and AND2 (N3100, N3099, N1829);
nor NOR4 (N3101, N3092, N1573, N2681, N1554);
not NOT1 (N3102, N3098);
or OR4 (N3103, N3084, N87, N2580, N2842);
xor XOR2 (N3104, N3066, N760);
nand NAND3 (N3105, N3095, N1708, N1617);
buf BUF1 (N3106, N3091);
xor XOR2 (N3107, N3102, N297);
nand NAND2 (N3108, N3100, N2842);
nor NOR2 (N3109, N3093, N2866);
or OR2 (N3110, N3097, N132);
not NOT1 (N3111, N3105);
not NOT1 (N3112, N3107);
nor NOR2 (N3113, N3106, N2158);
xor XOR2 (N3114, N3110, N762);
buf BUF1 (N3115, N3112);
and AND4 (N3116, N3104, N3043, N1692, N2559);
and AND3 (N3117, N3116, N1018, N2132);
nor NOR4 (N3118, N3117, N862, N1529, N251);
or OR2 (N3119, N3103, N1430);
and AND2 (N3120, N3115, N3112);
buf BUF1 (N3121, N3108);
nand NAND2 (N3122, N3101, N2142);
nor NOR4 (N3123, N3087, N2550, N715, N1337);
nand NAND2 (N3124, N3118, N1860);
and AND2 (N3125, N3122, N2126);
nand NAND4 (N3126, N3113, N1845, N1447, N1478);
nand NAND2 (N3127, N3126, N1756);
nand NAND4 (N3128, N3125, N1816, N890, N1157);
buf BUF1 (N3129, N3120);
nand NAND4 (N3130, N3128, N1758, N1026, N2956);
nand NAND2 (N3131, N3130, N2501);
nand NAND4 (N3132, N3119, N1583, N2312, N1144);
or OR2 (N3133, N3121, N2961);
xor XOR2 (N3134, N3132, N2982);
nor NOR3 (N3135, N3124, N425, N2915);
xor XOR2 (N3136, N3127, N83);
xor XOR2 (N3137, N3133, N2475);
and AND4 (N3138, N3134, N1560, N1345, N2124);
xor XOR2 (N3139, N3138, N2270);
xor XOR2 (N3140, N3129, N772);
or OR2 (N3141, N3140, N2152);
xor XOR2 (N3142, N3131, N256);
nand NAND2 (N3143, N3141, N969);
xor XOR2 (N3144, N3137, N2798);
or OR2 (N3145, N3111, N2884);
buf BUF1 (N3146, N3136);
nand NAND3 (N3147, N3135, N830, N1071);
nor NOR2 (N3148, N3139, N1274);
xor XOR2 (N3149, N3109, N1196);
nand NAND2 (N3150, N3147, N834);
nor NOR4 (N3151, N3149, N651, N2941, N1667);
and AND3 (N3152, N3114, N1279, N2054);
and AND3 (N3153, N3148, N3136, N2972);
nor NOR2 (N3154, N3146, N1349);
nor NOR4 (N3155, N3123, N2502, N2829, N2749);
nor NOR2 (N3156, N3151, N2693);
and AND3 (N3157, N3150, N1103, N3044);
xor XOR2 (N3158, N3145, N155);
buf BUF1 (N3159, N3153);
nor NOR4 (N3160, N3154, N2509, N2266, N931);
nand NAND4 (N3161, N3156, N1326, N1923, N1827);
nor NOR2 (N3162, N3144, N667);
and AND2 (N3163, N3152, N2600);
nor NOR2 (N3164, N3163, N2279);
and AND4 (N3165, N3155, N1738, N513, N929);
or OR4 (N3166, N3158, N2024, N1704, N355);
buf BUF1 (N3167, N3166);
xor XOR2 (N3168, N3159, N2228);
nand NAND2 (N3169, N3165, N338);
or OR4 (N3170, N3167, N651, N2733, N2133);
and AND2 (N3171, N3160, N1502);
or OR2 (N3172, N3157, N227);
and AND4 (N3173, N3161, N1490, N2280, N865);
nor NOR2 (N3174, N3168, N2701);
not NOT1 (N3175, N3174);
nand NAND4 (N3176, N3175, N481, N1226, N2073);
buf BUF1 (N3177, N3176);
nand NAND2 (N3178, N3177, N64);
or OR3 (N3179, N3173, N2841, N2228);
nor NOR4 (N3180, N3178, N2168, N119, N1933);
xor XOR2 (N3181, N3172, N2089);
and AND3 (N3182, N3179, N1257, N237);
or OR2 (N3183, N3162, N2014);
nor NOR4 (N3184, N3182, N164, N589, N2027);
buf BUF1 (N3185, N3184);
buf BUF1 (N3186, N3171);
not NOT1 (N3187, N3185);
buf BUF1 (N3188, N3142);
nand NAND2 (N3189, N3183, N1318);
and AND3 (N3190, N3164, N2329, N2987);
or OR3 (N3191, N3143, N1906, N1285);
or OR2 (N3192, N3187, N1220);
or OR4 (N3193, N3188, N2904, N1622, N2780);
or OR4 (N3194, N3189, N2829, N2127, N2967);
not NOT1 (N3195, N3170);
and AND4 (N3196, N3194, N166, N1809, N2308);
buf BUF1 (N3197, N3191);
not NOT1 (N3198, N3197);
buf BUF1 (N3199, N3186);
and AND2 (N3200, N3196, N2441);
not NOT1 (N3201, N3199);
buf BUF1 (N3202, N3195);
not NOT1 (N3203, N3192);
or OR3 (N3204, N3193, N406, N2080);
nor NOR3 (N3205, N3181, N1991, N1913);
or OR2 (N3206, N3169, N95);
not NOT1 (N3207, N3204);
nor NOR3 (N3208, N3198, N1443, N54);
not NOT1 (N3209, N3201);
nand NAND4 (N3210, N3205, N158, N909, N760);
xor XOR2 (N3211, N3180, N2882);
nor NOR3 (N3212, N3211, N845, N1871);
nand NAND3 (N3213, N3208, N742, N1928);
and AND4 (N3214, N3200, N241, N484, N3163);
nand NAND2 (N3215, N3214, N763);
not NOT1 (N3216, N3202);
and AND4 (N3217, N3206, N3007, N265, N1318);
or OR3 (N3218, N3212, N1690, N1532);
nor NOR3 (N3219, N3218, N2574, N3204);
buf BUF1 (N3220, N3217);
nand NAND3 (N3221, N3203, N1955, N1246);
nand NAND4 (N3222, N3221, N682, N724, N3142);
and AND4 (N3223, N3216, N1561, N2725, N2887);
or OR4 (N3224, N3222, N1487, N1857, N2770);
nor NOR3 (N3225, N3224, N1046, N1254);
or OR3 (N3226, N3207, N1248, N1559);
buf BUF1 (N3227, N3219);
nand NAND3 (N3228, N3213, N687, N2793);
nand NAND2 (N3229, N3225, N1294);
not NOT1 (N3230, N3226);
xor XOR2 (N3231, N3228, N1755);
nand NAND3 (N3232, N3215, N2770, N1895);
xor XOR2 (N3233, N3229, N3198);
nor NOR2 (N3234, N3231, N2149);
buf BUF1 (N3235, N3233);
buf BUF1 (N3236, N3230);
nor NOR3 (N3237, N3232, N2194, N1924);
buf BUF1 (N3238, N3210);
buf BUF1 (N3239, N3209);
nor NOR3 (N3240, N3227, N373, N2574);
nor NOR4 (N3241, N3190, N1796, N534, N803);
not NOT1 (N3242, N3235);
buf BUF1 (N3243, N3238);
buf BUF1 (N3244, N3243);
nand NAND2 (N3245, N3244, N239);
or OR4 (N3246, N3240, N3231, N3177, N1481);
xor XOR2 (N3247, N3223, N3226);
nor NOR4 (N3248, N3237, N259, N1636, N1523);
or OR2 (N3249, N3248, N1526);
nand NAND3 (N3250, N3220, N1578, N2173);
and AND3 (N3251, N3250, N617, N3141);
nor NOR4 (N3252, N3234, N446, N3041, N2170);
and AND2 (N3253, N3249, N2522);
buf BUF1 (N3254, N3252);
nand NAND3 (N3255, N3254, N2588, N2007);
xor XOR2 (N3256, N3253, N1374);
not NOT1 (N3257, N3245);
nor NOR3 (N3258, N3236, N1157, N153);
and AND4 (N3259, N3246, N3249, N646, N604);
nor NOR4 (N3260, N3255, N2834, N1230, N49);
xor XOR2 (N3261, N3256, N636);
not NOT1 (N3262, N3261);
nand NAND4 (N3263, N3239, N1862, N1257, N450);
not NOT1 (N3264, N3241);
nand NAND2 (N3265, N3262, N1250);
nand NAND4 (N3266, N3259, N1199, N1779, N1749);
xor XOR2 (N3267, N3264, N2250);
or OR3 (N3268, N3247, N56, N2511);
xor XOR2 (N3269, N3266, N1364);
not NOT1 (N3270, N3268);
nor NOR4 (N3271, N3251, N898, N593, N20);
buf BUF1 (N3272, N3263);
nor NOR2 (N3273, N3269, N3011);
and AND4 (N3274, N3242, N833, N1435, N432);
buf BUF1 (N3275, N3273);
nand NAND4 (N3276, N3258, N3148, N2418, N586);
and AND2 (N3277, N3271, N2805);
nand NAND3 (N3278, N3260, N1896, N1432);
xor XOR2 (N3279, N3276, N1426);
nand NAND2 (N3280, N3265, N3245);
or OR4 (N3281, N3272, N1835, N300, N3256);
and AND3 (N3282, N3280, N2838, N2265);
xor XOR2 (N3283, N3278, N341);
and AND3 (N3284, N3274, N976, N1668);
buf BUF1 (N3285, N3277);
xor XOR2 (N3286, N3282, N1789);
or OR4 (N3287, N3275, N877, N3179, N1644);
and AND2 (N3288, N3267, N2740);
xor XOR2 (N3289, N3257, N2031);
or OR2 (N3290, N3270, N377);
xor XOR2 (N3291, N3284, N1430);
or OR2 (N3292, N3285, N2944);
nand NAND3 (N3293, N3290, N2975, N3217);
not NOT1 (N3294, N3292);
or OR2 (N3295, N3288, N1643);
nor NOR4 (N3296, N3295, N2583, N2279, N130);
not NOT1 (N3297, N3291);
buf BUF1 (N3298, N3281);
xor XOR2 (N3299, N3297, N2567);
not NOT1 (N3300, N3299);
not NOT1 (N3301, N3279);
not NOT1 (N3302, N3301);
nor NOR4 (N3303, N3287, N2767, N1161, N2782);
or OR3 (N3304, N3286, N2112, N141);
xor XOR2 (N3305, N3303, N991);
xor XOR2 (N3306, N3304, N157);
and AND2 (N3307, N3283, N1644);
xor XOR2 (N3308, N3294, N380);
xor XOR2 (N3309, N3296, N2709);
not NOT1 (N3310, N3300);
nand NAND4 (N3311, N3289, N1502, N713, N1873);
xor XOR2 (N3312, N3307, N997);
buf BUF1 (N3313, N3302);
not NOT1 (N3314, N3293);
not NOT1 (N3315, N3308);
xor XOR2 (N3316, N3315, N391);
or OR4 (N3317, N3305, N2053, N27, N2934);
or OR3 (N3318, N3314, N94, N2283);
buf BUF1 (N3319, N3298);
nand NAND3 (N3320, N3311, N609, N1849);
or OR2 (N3321, N3309, N147);
buf BUF1 (N3322, N3312);
nor NOR2 (N3323, N3321, N1038);
nor NOR2 (N3324, N3306, N205);
nor NOR2 (N3325, N3310, N48);
xor XOR2 (N3326, N3318, N2090);
nor NOR4 (N3327, N3324, N1833, N1546, N3194);
and AND4 (N3328, N3327, N1540, N2370, N1445);
nand NAND2 (N3329, N3326, N2438);
not NOT1 (N3330, N3313);
or OR3 (N3331, N3317, N443, N2720);
or OR2 (N3332, N3331, N2808);
and AND2 (N3333, N3319, N196);
not NOT1 (N3334, N3322);
xor XOR2 (N3335, N3334, N3090);
xor XOR2 (N3336, N3333, N1164);
xor XOR2 (N3337, N3328, N2449);
or OR2 (N3338, N3323, N378);
or OR3 (N3339, N3330, N1666, N2276);
nand NAND4 (N3340, N3338, N1902, N2879, N2864);
nor NOR4 (N3341, N3332, N2277, N3053, N1068);
or OR2 (N3342, N3325, N398);
xor XOR2 (N3343, N3316, N2634);
buf BUF1 (N3344, N3320);
not NOT1 (N3345, N3341);
or OR4 (N3346, N3345, N137, N1298, N2280);
nand NAND2 (N3347, N3342, N3265);
xor XOR2 (N3348, N3329, N2047);
and AND4 (N3349, N3339, N2831, N1705, N2594);
nor NOR2 (N3350, N3349, N687);
and AND4 (N3351, N3348, N3297, N1013, N1379);
not NOT1 (N3352, N3346);
not NOT1 (N3353, N3336);
xor XOR2 (N3354, N3347, N2668);
not NOT1 (N3355, N3335);
xor XOR2 (N3356, N3354, N857);
nor NOR3 (N3357, N3352, N2465, N2134);
or OR3 (N3358, N3343, N267, N127);
xor XOR2 (N3359, N3358, N416);
buf BUF1 (N3360, N3353);
nor NOR3 (N3361, N3350, N135, N2680);
and AND3 (N3362, N3355, N5, N193);
xor XOR2 (N3363, N3340, N1724);
not NOT1 (N3364, N3356);
buf BUF1 (N3365, N3364);
or OR4 (N3366, N3365, N3029, N2786, N2437);
and AND3 (N3367, N3366, N2512, N597);
nor NOR3 (N3368, N3337, N3359, N1023);
nand NAND2 (N3369, N841, N464);
not NOT1 (N3370, N3357);
xor XOR2 (N3371, N3369, N3054);
nor NOR2 (N3372, N3360, N12);
nand NAND3 (N3373, N3362, N397, N522);
nor NOR2 (N3374, N3371, N508);
or OR4 (N3375, N3351, N2053, N2754, N1530);
and AND3 (N3376, N3370, N2731, N2928);
nand NAND3 (N3377, N3374, N2337, N2296);
not NOT1 (N3378, N3367);
and AND2 (N3379, N3378, N3246);
or OR2 (N3380, N3376, N3143);
nand NAND2 (N3381, N3344, N2858);
buf BUF1 (N3382, N3380);
or OR4 (N3383, N3379, N2680, N523, N2674);
or OR2 (N3384, N3382, N112);
xor XOR2 (N3385, N3372, N2189);
and AND3 (N3386, N3373, N419, N1939);
xor XOR2 (N3387, N3384, N1974);
and AND2 (N3388, N3387, N220);
or OR4 (N3389, N3386, N609, N466, N1248);
nand NAND2 (N3390, N3377, N970);
buf BUF1 (N3391, N3383);
or OR4 (N3392, N3390, N153, N1352, N3087);
not NOT1 (N3393, N3381);
not NOT1 (N3394, N3385);
not NOT1 (N3395, N3391);
or OR2 (N3396, N3388, N718);
and AND2 (N3397, N3394, N3046);
nor NOR4 (N3398, N3368, N355, N1687, N3289);
and AND4 (N3399, N3393, N220, N1776, N3022);
nand NAND2 (N3400, N3363, N504);
not NOT1 (N3401, N3399);
buf BUF1 (N3402, N3392);
or OR2 (N3403, N3389, N704);
xor XOR2 (N3404, N3395, N411);
not NOT1 (N3405, N3361);
nor NOR4 (N3406, N3401, N231, N1501, N317);
or OR2 (N3407, N3403, N1223);
not NOT1 (N3408, N3405);
buf BUF1 (N3409, N3404);
buf BUF1 (N3410, N3375);
nor NOR3 (N3411, N3398, N116, N3337);
buf BUF1 (N3412, N3400);
nor NOR4 (N3413, N3396, N1307, N138, N571);
buf BUF1 (N3414, N3408);
or OR3 (N3415, N3407, N3224, N776);
nor NOR4 (N3416, N3415, N2558, N267, N1562);
and AND4 (N3417, N3412, N2160, N2369, N786);
nand NAND2 (N3418, N3411, N3365);
not NOT1 (N3419, N3402);
or OR3 (N3420, N3418, N1564, N1770);
nor NOR4 (N3421, N3419, N2668, N1827, N647);
xor XOR2 (N3422, N3406, N2877);
nand NAND4 (N3423, N3420, N1154, N2418, N2425);
xor XOR2 (N3424, N3422, N1634);
nand NAND4 (N3425, N3416, N2482, N1253, N230);
not NOT1 (N3426, N3397);
or OR2 (N3427, N3423, N3385);
not NOT1 (N3428, N3425);
and AND2 (N3429, N3428, N2138);
xor XOR2 (N3430, N3426, N2991);
buf BUF1 (N3431, N3409);
and AND3 (N3432, N3431, N1170, N148);
buf BUF1 (N3433, N3413);
not NOT1 (N3434, N3410);
not NOT1 (N3435, N3432);
and AND3 (N3436, N3414, N3399, N3048);
xor XOR2 (N3437, N3434, N867);
nand NAND2 (N3438, N3433, N1429);
nor NOR3 (N3439, N3427, N752, N802);
or OR4 (N3440, N3424, N3068, N2311, N1514);
or OR2 (N3441, N3438, N1313);
not NOT1 (N3442, N3421);
and AND2 (N3443, N3437, N347);
xor XOR2 (N3444, N3440, N234);
nand NAND4 (N3445, N3439, N474, N1174, N1669);
xor XOR2 (N3446, N3430, N1798);
nand NAND3 (N3447, N3444, N873, N983);
nor NOR2 (N3448, N3441, N2048);
nor NOR3 (N3449, N3448, N2819, N2494);
not NOT1 (N3450, N3435);
and AND3 (N3451, N3449, N2612, N992);
not NOT1 (N3452, N3450);
not NOT1 (N3453, N3451);
nor NOR3 (N3454, N3445, N2825, N1323);
xor XOR2 (N3455, N3453, N781);
nand NAND2 (N3456, N3417, N1682);
xor XOR2 (N3457, N3447, N1686);
buf BUF1 (N3458, N3442);
xor XOR2 (N3459, N3436, N1674);
nor NOR3 (N3460, N3458, N2456, N352);
buf BUF1 (N3461, N3443);
buf BUF1 (N3462, N3457);
or OR4 (N3463, N3446, N1694, N569, N3374);
not NOT1 (N3464, N3461);
or OR4 (N3465, N3464, N643, N2114, N2849);
nor NOR3 (N3466, N3456, N2700, N2235);
xor XOR2 (N3467, N3462, N876);
buf BUF1 (N3468, N3454);
nand NAND2 (N3469, N3467, N2217);
nor NOR4 (N3470, N3429, N144, N874, N1953);
or OR3 (N3471, N3452, N3061, N3225);
buf BUF1 (N3472, N3465);
xor XOR2 (N3473, N3472, N708);
and AND2 (N3474, N3473, N261);
or OR4 (N3475, N3455, N153, N3261, N1074);
not NOT1 (N3476, N3463);
buf BUF1 (N3477, N3469);
xor XOR2 (N3478, N3460, N1289);
xor XOR2 (N3479, N3475, N81);
xor XOR2 (N3480, N3479, N3164);
not NOT1 (N3481, N3466);
nand NAND2 (N3482, N3474, N1924);
and AND2 (N3483, N3459, N1188);
not NOT1 (N3484, N3480);
buf BUF1 (N3485, N3483);
nand NAND4 (N3486, N3468, N105, N2057, N473);
nor NOR4 (N3487, N3484, N2918, N306, N1769);
and AND4 (N3488, N3471, N569, N2173, N2279);
nor NOR2 (N3489, N3485, N3405);
xor XOR2 (N3490, N3488, N119);
not NOT1 (N3491, N3490);
nand NAND4 (N3492, N3476, N2356, N40, N1739);
buf BUF1 (N3493, N3470);
buf BUF1 (N3494, N3491);
not NOT1 (N3495, N3481);
buf BUF1 (N3496, N3495);
and AND3 (N3497, N3482, N1639, N1540);
not NOT1 (N3498, N3478);
nand NAND3 (N3499, N3494, N2853, N2553);
not NOT1 (N3500, N3498);
not NOT1 (N3501, N3499);
and AND3 (N3502, N3489, N42, N2602);
nor NOR3 (N3503, N3496, N1619, N191);
nor NOR2 (N3504, N3500, N1829);
and AND2 (N3505, N3487, N2169);
nor NOR4 (N3506, N3505, N924, N3196, N3421);
buf BUF1 (N3507, N3493);
buf BUF1 (N3508, N3503);
or OR3 (N3509, N3497, N2566, N3459);
or OR3 (N3510, N3492, N2898, N693);
nand NAND4 (N3511, N3486, N169, N607, N2851);
or OR4 (N3512, N3508, N1313, N1564, N2220);
buf BUF1 (N3513, N3512);
nand NAND2 (N3514, N3504, N2095);
and AND4 (N3515, N3510, N862, N315, N492);
not NOT1 (N3516, N3501);
not NOT1 (N3517, N3506);
buf BUF1 (N3518, N3514);
nor NOR4 (N3519, N3515, N2118, N1134, N3344);
or OR3 (N3520, N3516, N3061, N3178);
nand NAND2 (N3521, N3507, N2624);
not NOT1 (N3522, N3513);
and AND4 (N3523, N3511, N21, N305, N2599);
xor XOR2 (N3524, N3520, N254);
and AND2 (N3525, N3517, N2891);
nor NOR2 (N3526, N3524, N3215);
and AND2 (N3527, N3509, N1153);
buf BUF1 (N3528, N3477);
buf BUF1 (N3529, N3525);
nand NAND4 (N3530, N3528, N1958, N1179, N1693);
nand NAND4 (N3531, N3519, N1851, N2611, N1864);
not NOT1 (N3532, N3529);
not NOT1 (N3533, N3518);
and AND4 (N3534, N3532, N2486, N1797, N196);
nor NOR3 (N3535, N3526, N468, N3289);
or OR3 (N3536, N3534, N3149, N73);
or OR3 (N3537, N3533, N2106, N441);
buf BUF1 (N3538, N3531);
not NOT1 (N3539, N3502);
xor XOR2 (N3540, N3538, N939);
or OR3 (N3541, N3536, N3059, N1016);
nor NOR2 (N3542, N3540, N980);
nand NAND4 (N3543, N3521, N2154, N1690, N895);
nand NAND3 (N3544, N3530, N453, N3055);
or OR2 (N3545, N3535, N1346);
not NOT1 (N3546, N3523);
nand NAND2 (N3547, N3537, N508);
buf BUF1 (N3548, N3539);
nor NOR4 (N3549, N3527, N1963, N1139, N2029);
nand NAND3 (N3550, N3546, N3518, N211);
or OR3 (N3551, N3543, N928, N2323);
not NOT1 (N3552, N3545);
or OR3 (N3553, N3542, N379, N392);
nand NAND2 (N3554, N3548, N170);
not NOT1 (N3555, N3552);
or OR4 (N3556, N3547, N1427, N2917, N2582);
nor NOR3 (N3557, N3556, N923, N1203);
buf BUF1 (N3558, N3555);
xor XOR2 (N3559, N3541, N2853);
xor XOR2 (N3560, N3550, N1908);
xor XOR2 (N3561, N3522, N228);
xor XOR2 (N3562, N3553, N160);
and AND4 (N3563, N3549, N2834, N1676, N3465);
nand NAND3 (N3564, N3554, N2560, N910);
and AND4 (N3565, N3551, N3489, N391, N1093);
not NOT1 (N3566, N3565);
nand NAND4 (N3567, N3564, N2581, N923, N2969);
xor XOR2 (N3568, N3561, N1219);
buf BUF1 (N3569, N3568);
and AND2 (N3570, N3559, N1694);
xor XOR2 (N3571, N3570, N2906);
or OR4 (N3572, N3571, N562, N2310, N251);
or OR2 (N3573, N3544, N1040);
buf BUF1 (N3574, N3560);
nor NOR4 (N3575, N3563, N893, N468, N2918);
nand NAND3 (N3576, N3573, N1024, N1194);
nand NAND3 (N3577, N3575, N3020, N1712);
or OR3 (N3578, N3572, N2137, N2723);
not NOT1 (N3579, N3577);
buf BUF1 (N3580, N3557);
not NOT1 (N3581, N3578);
xor XOR2 (N3582, N3567, N2019);
not NOT1 (N3583, N3580);
or OR4 (N3584, N3581, N2015, N956, N2051);
nor NOR2 (N3585, N3566, N500);
or OR2 (N3586, N3569, N2335);
and AND2 (N3587, N3586, N1347);
or OR3 (N3588, N3562, N1815, N283);
or OR4 (N3589, N3579, N3117, N411, N3374);
buf BUF1 (N3590, N3558);
nand NAND3 (N3591, N3588, N985, N1868);
and AND3 (N3592, N3591, N2568, N2629);
nor NOR3 (N3593, N3592, N3439, N3065);
nand NAND3 (N3594, N3585, N2506, N3005);
nor NOR3 (N3595, N3593, N282, N3097);
nor NOR4 (N3596, N3576, N933, N493, N417);
or OR4 (N3597, N3574, N3150, N560, N1824);
or OR4 (N3598, N3584, N3045, N557, N554);
and AND4 (N3599, N3589, N378, N436, N2472);
nand NAND4 (N3600, N3587, N2891, N1678, N2365);
not NOT1 (N3601, N3594);
not NOT1 (N3602, N3601);
or OR3 (N3603, N3600, N2274, N157);
xor XOR2 (N3604, N3603, N1121);
buf BUF1 (N3605, N3590);
or OR4 (N3606, N3602, N2924, N3025, N3324);
or OR3 (N3607, N3582, N1897, N3494);
and AND3 (N3608, N3596, N170, N1538);
nor NOR2 (N3609, N3598, N2955);
nor NOR4 (N3610, N3609, N2126, N675, N1556);
or OR4 (N3611, N3608, N2511, N990, N548);
xor XOR2 (N3612, N3610, N1455);
not NOT1 (N3613, N3605);
nor NOR2 (N3614, N3604, N624);
or OR3 (N3615, N3612, N606, N986);
or OR4 (N3616, N3614, N2735, N2512, N3167);
and AND4 (N3617, N3606, N1677, N1260, N2609);
nand NAND4 (N3618, N3615, N2324, N2334, N2471);
or OR4 (N3619, N3613, N153, N1293, N1417);
buf BUF1 (N3620, N3616);
and AND4 (N3621, N3611, N3566, N2120, N346);
nand NAND4 (N3622, N3618, N1505, N3297, N1945);
and AND4 (N3623, N3622, N1721, N323, N2276);
buf BUF1 (N3624, N3597);
or OR3 (N3625, N3620, N2664, N986);
and AND2 (N3626, N3625, N1974);
nor NOR4 (N3627, N3617, N347, N2780, N1711);
nor NOR3 (N3628, N3619, N2473, N1598);
or OR3 (N3629, N3607, N1612, N706);
nor NOR2 (N3630, N3621, N986);
nand NAND2 (N3631, N3627, N1753);
xor XOR2 (N3632, N3629, N880);
or OR4 (N3633, N3599, N2269, N801, N2873);
and AND4 (N3634, N3632, N2466, N2048, N1226);
nand NAND4 (N3635, N3633, N941, N3132, N3542);
and AND3 (N3636, N3630, N2408, N2188);
nand NAND4 (N3637, N3635, N1243, N2299, N1083);
and AND2 (N3638, N3583, N1899);
not NOT1 (N3639, N3623);
and AND2 (N3640, N3634, N673);
and AND2 (N3641, N3595, N1246);
xor XOR2 (N3642, N3637, N183);
nand NAND2 (N3643, N3631, N3009);
and AND3 (N3644, N3639, N2663, N192);
buf BUF1 (N3645, N3628);
or OR4 (N3646, N3645, N390, N852, N1910);
buf BUF1 (N3647, N3646);
not NOT1 (N3648, N3638);
and AND3 (N3649, N3624, N529, N2718);
nor NOR2 (N3650, N3648, N3214);
nor NOR4 (N3651, N3647, N2224, N3571, N2592);
not NOT1 (N3652, N3626);
buf BUF1 (N3653, N3651);
xor XOR2 (N3654, N3650, N2070);
nand NAND4 (N3655, N3641, N777, N2010, N3251);
nand NAND4 (N3656, N3652, N3583, N3630, N1482);
buf BUF1 (N3657, N3654);
xor XOR2 (N3658, N3655, N399);
buf BUF1 (N3659, N3642);
and AND4 (N3660, N3656, N1260, N1767, N2790);
nand NAND4 (N3661, N3658, N2811, N2693, N2446);
nand NAND4 (N3662, N3649, N937, N1159, N934);
nor NOR4 (N3663, N3661, N3157, N1156, N1283);
not NOT1 (N3664, N3659);
buf BUF1 (N3665, N3663);
not NOT1 (N3666, N3665);
not NOT1 (N3667, N3643);
nand NAND2 (N3668, N3664, N2126);
xor XOR2 (N3669, N3662, N3643);
not NOT1 (N3670, N3668);
buf BUF1 (N3671, N3640);
not NOT1 (N3672, N3666);
buf BUF1 (N3673, N3670);
nor NOR3 (N3674, N3671, N653, N1884);
nor NOR3 (N3675, N3669, N3316, N1303);
and AND2 (N3676, N3653, N1472);
nand NAND4 (N3677, N3676, N2753, N2619, N2764);
or OR3 (N3678, N3672, N1861, N1229);
nand NAND3 (N3679, N3660, N873, N132);
and AND3 (N3680, N3673, N458, N3206);
and AND3 (N3681, N3680, N1773, N1272);
nor NOR2 (N3682, N3667, N3494);
buf BUF1 (N3683, N3682);
not NOT1 (N3684, N3678);
or OR4 (N3685, N3657, N2055, N3471, N2573);
xor XOR2 (N3686, N3674, N161);
nand NAND4 (N3687, N3686, N776, N2576, N1330);
and AND3 (N3688, N3685, N1162, N1373);
xor XOR2 (N3689, N3636, N2182);
xor XOR2 (N3690, N3684, N3295);
nor NOR2 (N3691, N3679, N97);
not NOT1 (N3692, N3677);
nor NOR2 (N3693, N3689, N3418);
not NOT1 (N3694, N3687);
nor NOR2 (N3695, N3692, N665);
buf BUF1 (N3696, N3693);
nand NAND2 (N3697, N3695, N3448);
not NOT1 (N3698, N3694);
buf BUF1 (N3699, N3644);
nand NAND4 (N3700, N3691, N706, N3153, N1111);
buf BUF1 (N3701, N3697);
not NOT1 (N3702, N3701);
or OR3 (N3703, N3700, N3022, N1190);
or OR4 (N3704, N3683, N768, N3319, N3250);
xor XOR2 (N3705, N3703, N966);
nand NAND4 (N3706, N3699, N939, N3601, N2631);
or OR2 (N3707, N3705, N3570);
nand NAND4 (N3708, N3681, N2741, N3690, N1165);
and AND3 (N3709, N459, N1572, N769);
xor XOR2 (N3710, N3675, N932);
buf BUF1 (N3711, N3706);
buf BUF1 (N3712, N3711);
or OR3 (N3713, N3709, N821, N1674);
and AND4 (N3714, N3707, N3337, N2722, N1150);
and AND3 (N3715, N3702, N104, N2044);
nor NOR4 (N3716, N3696, N544, N1810, N857);
not NOT1 (N3717, N3712);
nor NOR4 (N3718, N3710, N3511, N2117, N1340);
not NOT1 (N3719, N3717);
nand NAND3 (N3720, N3708, N1384, N733);
nor NOR4 (N3721, N3719, N2747, N2884, N1502);
nor NOR2 (N3722, N3716, N2811);
xor XOR2 (N3723, N3714, N2521);
xor XOR2 (N3724, N3723, N2621);
or OR2 (N3725, N3722, N3602);
or OR2 (N3726, N3721, N3096);
or OR2 (N3727, N3704, N481);
and AND2 (N3728, N3724, N1275);
nand NAND4 (N3729, N3725, N2299, N3266, N2325);
nand NAND4 (N3730, N3720, N611, N2181, N2373);
nand NAND3 (N3731, N3718, N2911, N1435);
or OR2 (N3732, N3728, N1363);
or OR2 (N3733, N3731, N1);
or OR3 (N3734, N3730, N3155, N2664);
nor NOR2 (N3735, N3688, N3001);
xor XOR2 (N3736, N3735, N703);
xor XOR2 (N3737, N3734, N2727);
and AND4 (N3738, N3736, N1201, N1920, N2519);
and AND2 (N3739, N3733, N2497);
buf BUF1 (N3740, N3727);
nor NOR2 (N3741, N3740, N2168);
nor NOR2 (N3742, N3713, N1129);
nor NOR3 (N3743, N3742, N2041, N247);
nand NAND2 (N3744, N3738, N1120);
not NOT1 (N3745, N3732);
buf BUF1 (N3746, N3744);
nand NAND4 (N3747, N3698, N2550, N3097, N3264);
xor XOR2 (N3748, N3747, N2349);
buf BUF1 (N3749, N3739);
buf BUF1 (N3750, N3748);
buf BUF1 (N3751, N3741);
and AND3 (N3752, N3715, N917, N2211);
xor XOR2 (N3753, N3745, N934);
nor NOR4 (N3754, N3753, N469, N1280, N416);
or OR3 (N3755, N3729, N3085, N911);
not NOT1 (N3756, N3751);
buf BUF1 (N3757, N3752);
buf BUF1 (N3758, N3749);
xor XOR2 (N3759, N3726, N1645);
nand NAND3 (N3760, N3754, N1427, N3505);
buf BUF1 (N3761, N3760);
nand NAND2 (N3762, N3759, N2074);
and AND3 (N3763, N3746, N2385, N1138);
or OR2 (N3764, N3756, N2664);
nand NAND2 (N3765, N3743, N1674);
or OR3 (N3766, N3757, N2233, N11);
nand NAND3 (N3767, N3737, N405, N2452);
xor XOR2 (N3768, N3761, N3400);
and AND2 (N3769, N3767, N2855);
not NOT1 (N3770, N3762);
xor XOR2 (N3771, N3766, N1361);
nand NAND2 (N3772, N3763, N94);
and AND3 (N3773, N3755, N247, N1305);
buf BUF1 (N3774, N3771);
buf BUF1 (N3775, N3758);
xor XOR2 (N3776, N3775, N1830);
not NOT1 (N3777, N3773);
and AND4 (N3778, N3764, N1509, N3124, N401);
nor NOR2 (N3779, N3750, N2532);
buf BUF1 (N3780, N3769);
buf BUF1 (N3781, N3765);
buf BUF1 (N3782, N3776);
nand NAND3 (N3783, N3770, N353, N365);
and AND4 (N3784, N3777, N705, N3370, N2380);
nor NOR4 (N3785, N3781, N1752, N1279, N1382);
nand NAND2 (N3786, N3784, N2658);
not NOT1 (N3787, N3780);
not NOT1 (N3788, N3787);
nor NOR2 (N3789, N3779, N3541);
nor NOR4 (N3790, N3786, N1515, N2893, N3147);
nand NAND4 (N3791, N3778, N3301, N1293, N1685);
buf BUF1 (N3792, N3790);
and AND2 (N3793, N3792, N564);
buf BUF1 (N3794, N3782);
buf BUF1 (N3795, N3772);
nand NAND4 (N3796, N3794, N247, N1432, N824);
nor NOR3 (N3797, N3789, N3671, N1209);
buf BUF1 (N3798, N3797);
and AND4 (N3799, N3774, N2978, N2951, N754);
not NOT1 (N3800, N3791);
buf BUF1 (N3801, N3788);
not NOT1 (N3802, N3801);
not NOT1 (N3803, N3768);
nand NAND4 (N3804, N3783, N10, N3423, N1163);
nor NOR3 (N3805, N3799, N3369, N170);
or OR2 (N3806, N3793, N3275);
xor XOR2 (N3807, N3796, N289);
nor NOR2 (N3808, N3800, N3721);
or OR4 (N3809, N3785, N3104, N980, N3280);
nand NAND4 (N3810, N3808, N2945, N600, N340);
nand NAND2 (N3811, N3802, N2090);
not NOT1 (N3812, N3806);
not NOT1 (N3813, N3810);
nor NOR2 (N3814, N3807, N275);
not NOT1 (N3815, N3798);
nor NOR4 (N3816, N3805, N862, N3235, N850);
not NOT1 (N3817, N3803);
nand NAND4 (N3818, N3795, N2657, N2941, N330);
xor XOR2 (N3819, N3818, N2463);
and AND3 (N3820, N3812, N1231, N3800);
nand NAND3 (N3821, N3804, N591, N1996);
xor XOR2 (N3822, N3819, N2251);
buf BUF1 (N3823, N3821);
xor XOR2 (N3824, N3811, N3442);
xor XOR2 (N3825, N3814, N2268);
xor XOR2 (N3826, N3823, N69);
nor NOR3 (N3827, N3820, N2518, N3370);
nor NOR2 (N3828, N3826, N3153);
nor NOR3 (N3829, N3824, N89, N2233);
nand NAND4 (N3830, N3828, N1695, N2012, N1071);
or OR3 (N3831, N3816, N2558, N2279);
xor XOR2 (N3832, N3822, N500);
not NOT1 (N3833, N3813);
buf BUF1 (N3834, N3829);
nand NAND2 (N3835, N3834, N2549);
not NOT1 (N3836, N3815);
xor XOR2 (N3837, N3836, N1758);
xor XOR2 (N3838, N3835, N1107);
and AND3 (N3839, N3809, N1681, N2921);
and AND3 (N3840, N3837, N609, N1913);
and AND3 (N3841, N3839, N3453, N1218);
or OR2 (N3842, N3817, N3291);
xor XOR2 (N3843, N3831, N3061);
not NOT1 (N3844, N3825);
xor XOR2 (N3845, N3827, N1446);
xor XOR2 (N3846, N3842, N3604);
or OR4 (N3847, N3838, N890, N3717, N1230);
not NOT1 (N3848, N3844);
and AND4 (N3849, N3833, N168, N1076, N3043);
nor NOR3 (N3850, N3849, N2336, N1635);
and AND2 (N3851, N3848, N2517);
not NOT1 (N3852, N3847);
and AND3 (N3853, N3840, N922, N3802);
buf BUF1 (N3854, N3851);
buf BUF1 (N3855, N3845);
nand NAND3 (N3856, N3852, N971, N2554);
not NOT1 (N3857, N3841);
xor XOR2 (N3858, N3854, N2252);
nand NAND3 (N3859, N3846, N2161, N3354);
and AND4 (N3860, N3843, N1643, N1702, N1550);
buf BUF1 (N3861, N3857);
xor XOR2 (N3862, N3830, N350);
nand NAND2 (N3863, N3861, N1890);
buf BUF1 (N3864, N3855);
and AND2 (N3865, N3856, N1456);
and AND2 (N3866, N3865, N3234);
nor NOR4 (N3867, N3863, N3173, N1071, N1252);
not NOT1 (N3868, N3867);
xor XOR2 (N3869, N3864, N338);
nor NOR3 (N3870, N3868, N3020, N3825);
nor NOR3 (N3871, N3866, N3295, N80);
xor XOR2 (N3872, N3832, N89);
or OR3 (N3873, N3871, N3821, N3261);
nand NAND2 (N3874, N3853, N2811);
and AND2 (N3875, N3859, N1273);
nor NOR4 (N3876, N3874, N3030, N3383, N2365);
and AND4 (N3877, N3869, N553, N2998, N2847);
xor XOR2 (N3878, N3860, N1397);
and AND2 (N3879, N3875, N2882);
nand NAND3 (N3880, N3878, N923, N895);
xor XOR2 (N3881, N3880, N2924);
xor XOR2 (N3882, N3879, N2028);
nand NAND4 (N3883, N3877, N3077, N2320, N1230);
buf BUF1 (N3884, N3873);
buf BUF1 (N3885, N3862);
and AND3 (N3886, N3883, N1299, N824);
nand NAND2 (N3887, N3885, N3483);
nand NAND2 (N3888, N3850, N2945);
xor XOR2 (N3889, N3872, N2806);
or OR3 (N3890, N3858, N2896, N1120);
nand NAND2 (N3891, N3890, N2494);
xor XOR2 (N3892, N3888, N158);
buf BUF1 (N3893, N3876);
xor XOR2 (N3894, N3889, N3209);
buf BUF1 (N3895, N3881);
nor NOR3 (N3896, N3893, N3435, N1562);
and AND3 (N3897, N3892, N1130, N1639);
nand NAND2 (N3898, N3897, N2283);
nand NAND4 (N3899, N3884, N2444, N3267, N3278);
buf BUF1 (N3900, N3894);
and AND2 (N3901, N3891, N2931);
buf BUF1 (N3902, N3895);
nand NAND3 (N3903, N3887, N3577, N471);
not NOT1 (N3904, N3901);
buf BUF1 (N3905, N3882);
or OR4 (N3906, N3902, N2816, N670, N746);
and AND4 (N3907, N3886, N826, N132, N160);
and AND4 (N3908, N3896, N3549, N897, N2278);
buf BUF1 (N3909, N3904);
and AND4 (N3910, N3898, N3144, N181, N498);
xor XOR2 (N3911, N3903, N2537);
nand NAND3 (N3912, N3899, N2594, N2536);
nand NAND4 (N3913, N3910, N949, N1828, N3194);
or OR4 (N3914, N3912, N3006, N251, N861);
and AND3 (N3915, N3911, N2545, N2099);
nand NAND4 (N3916, N3913, N2840, N1629, N1371);
or OR4 (N3917, N3908, N1630, N613, N1335);
not NOT1 (N3918, N3907);
buf BUF1 (N3919, N3915);
nand NAND2 (N3920, N3914, N3044);
nand NAND2 (N3921, N3919, N1674);
not NOT1 (N3922, N3870);
not NOT1 (N3923, N3909);
nand NAND3 (N3924, N3900, N857, N3895);
not NOT1 (N3925, N3924);
nor NOR2 (N3926, N3905, N2701);
or OR3 (N3927, N3906, N825, N2787);
nor NOR3 (N3928, N3920, N32, N12);
nand NAND3 (N3929, N3916, N418, N1733);
not NOT1 (N3930, N3926);
not NOT1 (N3931, N3921);
and AND4 (N3932, N3931, N1566, N3454, N853);
xor XOR2 (N3933, N3932, N1316);
nand NAND4 (N3934, N3917, N1535, N1621, N2783);
buf BUF1 (N3935, N3930);
buf BUF1 (N3936, N3935);
or OR4 (N3937, N3933, N1173, N470, N3097);
xor XOR2 (N3938, N3918, N3744);
xor XOR2 (N3939, N3934, N1105);
or OR3 (N3940, N3927, N1537, N3277);
or OR3 (N3941, N3938, N292, N1944);
or OR2 (N3942, N3941, N3719);
nand NAND4 (N3943, N3936, N3583, N1590, N3071);
nor NOR2 (N3944, N3939, N1614);
xor XOR2 (N3945, N3928, N115);
nor NOR4 (N3946, N3922, N1068, N273, N2368);
and AND4 (N3947, N3940, N2769, N2365, N2906);
or OR3 (N3948, N3925, N1691, N2707);
nand NAND2 (N3949, N3945, N2410);
nand NAND2 (N3950, N3942, N2637);
xor XOR2 (N3951, N3948, N546);
not NOT1 (N3952, N3943);
or OR4 (N3953, N3944, N910, N965, N18);
or OR2 (N3954, N3953, N3279);
nand NAND4 (N3955, N3952, N3954, N2634, N1552);
nor NOR2 (N3956, N593, N2552);
xor XOR2 (N3957, N3955, N1861);
and AND4 (N3958, N3947, N112, N240, N1519);
nor NOR4 (N3959, N3923, N111, N854, N3232);
and AND4 (N3960, N3959, N1740, N425, N700);
not NOT1 (N3961, N3951);
xor XOR2 (N3962, N3961, N1627);
nand NAND4 (N3963, N3956, N1314, N1228, N2301);
xor XOR2 (N3964, N3957, N785);
nand NAND2 (N3965, N3962, N1687);
buf BUF1 (N3966, N3965);
xor XOR2 (N3967, N3966, N127);
buf BUF1 (N3968, N3960);
nor NOR2 (N3969, N3937, N1759);
nand NAND3 (N3970, N3949, N937, N1824);
xor XOR2 (N3971, N3958, N2115);
xor XOR2 (N3972, N3929, N813);
nor NOR3 (N3973, N3969, N1340, N940);
buf BUF1 (N3974, N3963);
buf BUF1 (N3975, N3968);
nand NAND2 (N3976, N3964, N2745);
not NOT1 (N3977, N3972);
nor NOR2 (N3978, N3975, N1289);
not NOT1 (N3979, N3973);
or OR4 (N3980, N3970, N3541, N1623, N104);
buf BUF1 (N3981, N3946);
or OR3 (N3982, N3981, N311, N1442);
xor XOR2 (N3983, N3980, N2360);
xor XOR2 (N3984, N3979, N2696);
or OR3 (N3985, N3976, N957, N1768);
or OR3 (N3986, N3974, N1788, N3469);
and AND2 (N3987, N3971, N2859);
not NOT1 (N3988, N3977);
xor XOR2 (N3989, N3967, N517);
and AND4 (N3990, N3986, N945, N2998, N3796);
buf BUF1 (N3991, N3987);
xor XOR2 (N3992, N3988, N3072);
or OR4 (N3993, N3985, N2235, N3378, N1273);
buf BUF1 (N3994, N3978);
or OR4 (N3995, N3994, N2076, N3836, N641);
nor NOR4 (N3996, N3992, N3385, N900, N687);
buf BUF1 (N3997, N3995);
buf BUF1 (N3998, N3996);
not NOT1 (N3999, N3983);
nand NAND4 (N4000, N3998, N1359, N1945, N175);
buf BUF1 (N4001, N3990);
and AND4 (N4002, N3989, N1264, N1323, N2446);
and AND2 (N4003, N3991, N3596);
xor XOR2 (N4004, N4003, N1703);
buf BUF1 (N4005, N4002);
or OR4 (N4006, N4001, N2507, N3801, N715);
not NOT1 (N4007, N4006);
and AND2 (N4008, N4007, N3325);
xor XOR2 (N4009, N3982, N3211);
nor NOR2 (N4010, N4004, N2136);
nor NOR4 (N4011, N4010, N2103, N2855, N882);
nor NOR4 (N4012, N3950, N767, N1908, N2701);
nor NOR4 (N4013, N4012, N2464, N300, N3999);
and AND2 (N4014, N15, N2944);
and AND2 (N4015, N4000, N2477);
not NOT1 (N4016, N4005);
not NOT1 (N4017, N3997);
xor XOR2 (N4018, N4013, N1244);
and AND3 (N4019, N3993, N3423, N3921);
not NOT1 (N4020, N4014);
xor XOR2 (N4021, N4015, N2604);
nand NAND3 (N4022, N4009, N3641, N2596);
nor NOR3 (N4023, N4016, N2585, N2520);
and AND3 (N4024, N4020, N3087, N2557);
and AND4 (N4025, N4008, N455, N1567, N6);
or OR4 (N4026, N4019, N1575, N729, N2916);
nand NAND2 (N4027, N4011, N2822);
or OR4 (N4028, N4024, N1302, N3091, N1948);
xor XOR2 (N4029, N4025, N383);
not NOT1 (N4030, N4018);
nand NAND2 (N4031, N4027, N1272);
not NOT1 (N4032, N4029);
nand NAND2 (N4033, N4030, N1001);
buf BUF1 (N4034, N4031);
xor XOR2 (N4035, N4033, N1145);
not NOT1 (N4036, N4022);
or OR4 (N4037, N4021, N2564, N3269, N3646);
and AND4 (N4038, N4017, N3347, N739, N213);
xor XOR2 (N4039, N4026, N182);
or OR4 (N4040, N4028, N1969, N1958, N2275);
nand NAND3 (N4041, N3984, N1899, N2059);
xor XOR2 (N4042, N4034, N1767);
and AND4 (N4043, N4041, N288, N1493, N3865);
not NOT1 (N4044, N4043);
nor NOR4 (N4045, N4035, N3559, N186, N1587);
nand NAND2 (N4046, N4044, N3076);
buf BUF1 (N4047, N4036);
nor NOR4 (N4048, N4032, N2077, N88, N732);
nor NOR3 (N4049, N4038, N4001, N3078);
nor NOR4 (N4050, N4040, N1301, N3273, N2100);
and AND4 (N4051, N4045, N1620, N986, N2426);
xor XOR2 (N4052, N4050, N671);
and AND2 (N4053, N4046, N3576);
not NOT1 (N4054, N4047);
and AND2 (N4055, N4039, N2117);
xor XOR2 (N4056, N4053, N3656);
nor NOR4 (N4057, N4048, N1771, N1235, N1341);
buf BUF1 (N4058, N4051);
nand NAND3 (N4059, N4023, N2162, N1927);
not NOT1 (N4060, N4059);
nor NOR2 (N4061, N4060, N1194);
buf BUF1 (N4062, N4061);
xor XOR2 (N4063, N4037, N3098);
and AND4 (N4064, N4062, N604, N3571, N2970);
not NOT1 (N4065, N4052);
buf BUF1 (N4066, N4056);
nand NAND2 (N4067, N4049, N1337);
and AND2 (N4068, N4065, N3016);
xor XOR2 (N4069, N4058, N1333);
buf BUF1 (N4070, N4069);
xor XOR2 (N4071, N4055, N1155);
nand NAND3 (N4072, N4066, N2775, N319);
and AND4 (N4073, N4063, N1285, N2125, N122);
not NOT1 (N4074, N4057);
xor XOR2 (N4075, N4068, N2942);
and AND2 (N4076, N4067, N3041);
buf BUF1 (N4077, N4074);
xor XOR2 (N4078, N4077, N539);
nand NAND3 (N4079, N4078, N681, N3333);
not NOT1 (N4080, N4076);
buf BUF1 (N4081, N4070);
buf BUF1 (N4082, N4081);
and AND2 (N4083, N4064, N3165);
or OR2 (N4084, N4082, N2311);
or OR4 (N4085, N4080, N743, N3649, N1633);
and AND2 (N4086, N4075, N2076);
or OR4 (N4087, N4073, N1201, N1350, N1430);
buf BUF1 (N4088, N4086);
nor NOR3 (N4089, N4088, N986, N2830);
and AND2 (N4090, N4085, N3827);
nor NOR3 (N4091, N4089, N534, N1710);
buf BUF1 (N4092, N4084);
or OR3 (N4093, N4083, N2830, N2292);
buf BUF1 (N4094, N4054);
or OR4 (N4095, N4093, N2565, N3585, N3048);
nand NAND4 (N4096, N4090, N3069, N3946, N2899);
not NOT1 (N4097, N4091);
and AND2 (N4098, N4079, N3706);
nor NOR3 (N4099, N4098, N2153, N1567);
and AND2 (N4100, N4071, N1195);
nor NOR3 (N4101, N4097, N2993, N3355);
and AND2 (N4102, N4042, N2431);
or OR3 (N4103, N4099, N1388, N3575);
not NOT1 (N4104, N4094);
or OR3 (N4105, N4095, N3069, N2388);
xor XOR2 (N4106, N4105, N3200);
buf BUF1 (N4107, N4087);
or OR4 (N4108, N4107, N3037, N1680, N635);
buf BUF1 (N4109, N4100);
buf BUF1 (N4110, N4101);
nand NAND3 (N4111, N4102, N2594, N3435);
nand NAND4 (N4112, N4109, N1440, N2271, N1216);
xor XOR2 (N4113, N4092, N4112);
or OR2 (N4114, N2077, N3176);
and AND2 (N4115, N4104, N684);
and AND3 (N4116, N4115, N756, N3320);
or OR4 (N4117, N4111, N3582, N1720, N149);
and AND3 (N4118, N4096, N2854, N558);
not NOT1 (N4119, N4116);
nor NOR4 (N4120, N4119, N3376, N3909, N1024);
buf BUF1 (N4121, N4108);
nor NOR2 (N4122, N4118, N3451);
xor XOR2 (N4123, N4121, N2514);
xor XOR2 (N4124, N4114, N293);
not NOT1 (N4125, N4120);
and AND2 (N4126, N4072, N1136);
or OR3 (N4127, N4126, N2316, N3836);
and AND4 (N4128, N4122, N2492, N1656, N4046);
and AND4 (N4129, N4128, N1183, N3651, N3747);
nand NAND2 (N4130, N4106, N2783);
buf BUF1 (N4131, N4125);
xor XOR2 (N4132, N4117, N502);
or OR3 (N4133, N4127, N3457, N3410);
not NOT1 (N4134, N4113);
not NOT1 (N4135, N4123);
nand NAND3 (N4136, N4134, N1555, N2818);
and AND2 (N4137, N4124, N1703);
xor XOR2 (N4138, N4136, N2442);
xor XOR2 (N4139, N4135, N1322);
buf BUF1 (N4140, N4133);
buf BUF1 (N4141, N4129);
not NOT1 (N4142, N4103);
and AND4 (N4143, N4130, N465, N3663, N3713);
nand NAND2 (N4144, N4139, N605);
and AND2 (N4145, N4144, N3732);
and AND3 (N4146, N4131, N3310, N2535);
not NOT1 (N4147, N4138);
xor XOR2 (N4148, N4137, N679);
nor NOR3 (N4149, N4140, N3629, N192);
and AND2 (N4150, N4142, N2800);
not NOT1 (N4151, N4110);
buf BUF1 (N4152, N4145);
and AND2 (N4153, N4152, N3445);
nand NAND3 (N4154, N4153, N413, N3722);
not NOT1 (N4155, N4154);
nor NOR4 (N4156, N4141, N265, N2382, N3242);
and AND3 (N4157, N4143, N2728, N1786);
or OR4 (N4158, N4150, N3563, N755, N3654);
buf BUF1 (N4159, N4149);
and AND3 (N4160, N4132, N4059, N1383);
not NOT1 (N4161, N4147);
buf BUF1 (N4162, N4155);
not NOT1 (N4163, N4157);
not NOT1 (N4164, N4160);
nor NOR4 (N4165, N4159, N2086, N641, N1068);
not NOT1 (N4166, N4164);
and AND2 (N4167, N4166, N564);
and AND2 (N4168, N4146, N440);
nor NOR2 (N4169, N4168, N4073);
and AND3 (N4170, N4148, N3305, N141);
buf BUF1 (N4171, N4151);
nand NAND4 (N4172, N4167, N3394, N1623, N2704);
nor NOR2 (N4173, N4162, N3244);
or OR4 (N4174, N4169, N4064, N1517, N1840);
and AND4 (N4175, N4163, N1091, N2768, N2800);
buf BUF1 (N4176, N4165);
and AND4 (N4177, N4170, N3402, N1800, N427);
or OR4 (N4178, N4156, N716, N229, N2241);
nand NAND4 (N4179, N4171, N2377, N3179, N1130);
or OR2 (N4180, N4158, N2339);
xor XOR2 (N4181, N4172, N2536);
nand NAND3 (N4182, N4180, N1490, N4153);
nand NAND4 (N4183, N4177, N3036, N4053, N1329);
nor NOR3 (N4184, N4175, N859, N2563);
not NOT1 (N4185, N4182);
buf BUF1 (N4186, N4174);
not NOT1 (N4187, N4179);
and AND4 (N4188, N4184, N1771, N3545, N2002);
nor NOR4 (N4189, N4176, N2277, N1815, N4044);
nor NOR3 (N4190, N4187, N3128, N1280);
not NOT1 (N4191, N4186);
and AND2 (N4192, N4183, N1033);
buf BUF1 (N4193, N4191);
nor NOR3 (N4194, N4161, N3226, N574);
nor NOR3 (N4195, N4188, N1751, N1405);
nand NAND3 (N4196, N4173, N156, N3669);
nand NAND4 (N4197, N4192, N4137, N450, N845);
nand NAND4 (N4198, N4181, N3333, N2111, N1534);
or OR4 (N4199, N4194, N4038, N1154, N1476);
xor XOR2 (N4200, N4196, N3941);
not NOT1 (N4201, N4189);
and AND2 (N4202, N4185, N150);
or OR4 (N4203, N4201, N810, N4162, N2943);
and AND2 (N4204, N4197, N48);
buf BUF1 (N4205, N4199);
not NOT1 (N4206, N4193);
buf BUF1 (N4207, N4205);
xor XOR2 (N4208, N4203, N1273);
nor NOR4 (N4209, N4202, N2406, N305, N2380);
or OR2 (N4210, N4190, N1404);
or OR3 (N4211, N4195, N526, N2162);
buf BUF1 (N4212, N4208);
or OR3 (N4213, N4210, N1503, N2493);
or OR2 (N4214, N4213, N911);
nand NAND4 (N4215, N4206, N1459, N2034, N3738);
and AND4 (N4216, N4198, N42, N835, N2978);
buf BUF1 (N4217, N4209);
xor XOR2 (N4218, N4215, N3598);
not NOT1 (N4219, N4200);
nor NOR4 (N4220, N4216, N2871, N2126, N2331);
buf BUF1 (N4221, N4207);
not NOT1 (N4222, N4212);
buf BUF1 (N4223, N4222);
not NOT1 (N4224, N4178);
buf BUF1 (N4225, N4224);
xor XOR2 (N4226, N4221, N419);
xor XOR2 (N4227, N4218, N438);
or OR4 (N4228, N4219, N1358, N3242, N3483);
and AND2 (N4229, N4217, N3225);
buf BUF1 (N4230, N4214);
not NOT1 (N4231, N4230);
nand NAND3 (N4232, N4211, N1775, N1584);
and AND4 (N4233, N4223, N2918, N752, N850);
or OR3 (N4234, N4231, N3207, N1105);
xor XOR2 (N4235, N4226, N503);
buf BUF1 (N4236, N4228);
and AND2 (N4237, N4220, N548);
and AND2 (N4238, N4235, N570);
and AND2 (N4239, N4238, N984);
nand NAND4 (N4240, N4225, N1355, N1999, N2237);
nor NOR4 (N4241, N4227, N1655, N1170, N4034);
not NOT1 (N4242, N4241);
not NOT1 (N4243, N4240);
nor NOR3 (N4244, N4236, N3791, N917);
xor XOR2 (N4245, N4229, N530);
nand NAND3 (N4246, N4232, N1051, N2743);
nand NAND2 (N4247, N4246, N2182);
xor XOR2 (N4248, N4244, N2700);
xor XOR2 (N4249, N4239, N1062);
and AND4 (N4250, N4248, N2638, N2951, N3651);
and AND4 (N4251, N4250, N1431, N56, N2056);
buf BUF1 (N4252, N4251);
not NOT1 (N4253, N4247);
not NOT1 (N4254, N4253);
or OR4 (N4255, N4252, N656, N3686, N2478);
or OR4 (N4256, N4234, N832, N3273, N2542);
xor XOR2 (N4257, N4242, N2542);
nor NOR2 (N4258, N4255, N3005);
nor NOR2 (N4259, N4243, N260);
nand NAND4 (N4260, N4237, N1504, N2276, N4120);
and AND4 (N4261, N4260, N1753, N1112, N403);
not NOT1 (N4262, N4245);
not NOT1 (N4263, N4261);
nor NOR4 (N4264, N4249, N2052, N4045, N1415);
or OR4 (N4265, N4262, N428, N193, N393);
or OR3 (N4266, N4264, N3305, N1443);
nand NAND3 (N4267, N4263, N2345, N516);
nor NOR2 (N4268, N4257, N3006);
xor XOR2 (N4269, N4268, N1125);
nand NAND2 (N4270, N4204, N3133);
and AND2 (N4271, N4256, N2641);
buf BUF1 (N4272, N4270);
not NOT1 (N4273, N4258);
and AND3 (N4274, N4269, N1919, N950);
not NOT1 (N4275, N4271);
buf BUF1 (N4276, N4266);
nor NOR2 (N4277, N4267, N455);
nand NAND2 (N4278, N4254, N285);
or OR4 (N4279, N4272, N1191, N639, N716);
nand NAND3 (N4280, N4274, N2244, N3258);
buf BUF1 (N4281, N4259);
not NOT1 (N4282, N4280);
or OR2 (N4283, N4233, N1958);
nand NAND2 (N4284, N4265, N3456);
nand NAND4 (N4285, N4276, N1101, N4153, N2267);
xor XOR2 (N4286, N4275, N2234);
buf BUF1 (N4287, N4283);
and AND2 (N4288, N4273, N1870);
buf BUF1 (N4289, N4284);
nand NAND4 (N4290, N4282, N1740, N160, N2436);
or OR3 (N4291, N4285, N1405, N2304);
or OR3 (N4292, N4289, N2582, N2067);
not NOT1 (N4293, N4278);
buf BUF1 (N4294, N4281);
xor XOR2 (N4295, N4294, N719);
nand NAND3 (N4296, N4295, N3302, N1426);
or OR2 (N4297, N4296, N4186);
and AND3 (N4298, N4292, N487, N1312);
not NOT1 (N4299, N4290);
or OR3 (N4300, N4279, N3898, N3778);
nor NOR3 (N4301, N4293, N1802, N2520);
nand NAND3 (N4302, N4286, N2808, N196);
xor XOR2 (N4303, N4298, N1234);
nand NAND3 (N4304, N4287, N2923, N1122);
and AND4 (N4305, N4304, N2844, N942, N4275);
and AND4 (N4306, N4297, N4299, N1832, N2203);
xor XOR2 (N4307, N4257, N2112);
or OR4 (N4308, N4277, N2501, N3718, N1482);
and AND3 (N4309, N4300, N2401, N3795);
nand NAND4 (N4310, N4306, N1525, N216, N1355);
buf BUF1 (N4311, N4301);
or OR3 (N4312, N4308, N2848, N3584);
nor NOR2 (N4313, N4305, N3770);
nor NOR2 (N4314, N4313, N2293);
and AND2 (N4315, N4302, N3981);
nor NOR4 (N4316, N4314, N737, N373, N1385);
not NOT1 (N4317, N4291);
nand NAND4 (N4318, N4288, N2735, N1761, N3288);
nor NOR3 (N4319, N4310, N3871, N79);
nor NOR4 (N4320, N4317, N3355, N2468, N3781);
nand NAND4 (N4321, N4303, N1741, N854, N185);
and AND3 (N4322, N4321, N218, N2741);
xor XOR2 (N4323, N4309, N1290);
nand NAND2 (N4324, N4316, N866);
nand NAND3 (N4325, N4311, N137, N2543);
buf BUF1 (N4326, N4312);
nor NOR4 (N4327, N4325, N3472, N2543, N715);
and AND3 (N4328, N4320, N292, N2783);
nand NAND3 (N4329, N4324, N3568, N2033);
not NOT1 (N4330, N4319);
not NOT1 (N4331, N4307);
nand NAND3 (N4332, N4315, N245, N4274);
and AND2 (N4333, N4322, N135);
buf BUF1 (N4334, N4328);
or OR2 (N4335, N4331, N1109);
or OR3 (N4336, N4333, N4174, N3191);
and AND3 (N4337, N4318, N308, N1016);
xor XOR2 (N4338, N4332, N1576);
and AND4 (N4339, N4323, N1544, N4155, N1098);
or OR3 (N4340, N4335, N1503, N3620);
not NOT1 (N4341, N4326);
or OR4 (N4342, N4336, N30, N25, N2794);
buf BUF1 (N4343, N4340);
nor NOR4 (N4344, N4334, N861, N3418, N2952);
buf BUF1 (N4345, N4329);
buf BUF1 (N4346, N4338);
not NOT1 (N4347, N4344);
xor XOR2 (N4348, N4346, N2565);
nor NOR3 (N4349, N4327, N1833, N924);
nor NOR4 (N4350, N4345, N1478, N3767, N2057);
buf BUF1 (N4351, N4342);
not NOT1 (N4352, N4330);
buf BUF1 (N4353, N4350);
nand NAND3 (N4354, N4347, N41, N2657);
buf BUF1 (N4355, N4351);
xor XOR2 (N4356, N4353, N194);
xor XOR2 (N4357, N4337, N3443);
buf BUF1 (N4358, N4357);
xor XOR2 (N4359, N4341, N1886);
buf BUF1 (N4360, N4356);
not NOT1 (N4361, N4354);
not NOT1 (N4362, N4359);
or OR4 (N4363, N4360, N1814, N1851, N193);
nor NOR2 (N4364, N4358, N480);
nand NAND4 (N4365, N4362, N896, N1160, N2596);
and AND2 (N4366, N4363, N2534);
xor XOR2 (N4367, N4366, N2012);
nand NAND2 (N4368, N4365, N3203);
or OR3 (N4369, N4348, N2032, N662);
buf BUF1 (N4370, N4361);
and AND2 (N4371, N4369, N94);
nor NOR3 (N4372, N4370, N3285, N1013);
and AND3 (N4373, N4367, N3028, N3533);
nand NAND3 (N4374, N4352, N1914, N3798);
nor NOR3 (N4375, N4368, N3561, N212);
buf BUF1 (N4376, N4364);
xor XOR2 (N4377, N4349, N4311);
nor NOR4 (N4378, N4371, N3458, N2245, N2410);
xor XOR2 (N4379, N4374, N3719);
not NOT1 (N4380, N4339);
nand NAND4 (N4381, N4378, N2861, N1888, N1851);
and AND4 (N4382, N4377, N4015, N993, N326);
and AND4 (N4383, N4381, N2613, N3269, N3484);
xor XOR2 (N4384, N4376, N1766);
or OR2 (N4385, N4343, N917);
buf BUF1 (N4386, N4383);
xor XOR2 (N4387, N4373, N3370);
not NOT1 (N4388, N4386);
xor XOR2 (N4389, N4387, N896);
not NOT1 (N4390, N4384);
and AND3 (N4391, N4375, N1364, N3109);
xor XOR2 (N4392, N4385, N1626);
and AND4 (N4393, N4392, N1846, N3410, N2156);
nand NAND4 (N4394, N4393, N907, N255, N4393);
buf BUF1 (N4395, N4372);
or OR2 (N4396, N4389, N1982);
buf BUF1 (N4397, N4388);
not NOT1 (N4398, N4390);
and AND4 (N4399, N4397, N541, N1730, N3260);
nand NAND4 (N4400, N4379, N2111, N769, N958);
nand NAND3 (N4401, N4398, N546, N4146);
and AND3 (N4402, N4395, N2260, N2801);
buf BUF1 (N4403, N4382);
nand NAND2 (N4404, N4399, N147);
nor NOR4 (N4405, N4402, N3881, N2650, N3078);
nand NAND3 (N4406, N4401, N1320, N2354);
not NOT1 (N4407, N4391);
and AND3 (N4408, N4400, N2635, N1810);
not NOT1 (N4409, N4355);
nand NAND3 (N4410, N4404, N3563, N3223);
and AND3 (N4411, N4405, N404, N663);
or OR3 (N4412, N4406, N1496, N3445);
xor XOR2 (N4413, N4412, N3513);
nand NAND4 (N4414, N4413, N4204, N3978, N2426);
and AND3 (N4415, N4394, N2719, N308);
buf BUF1 (N4416, N4407);
nor NOR3 (N4417, N4396, N49, N696);
xor XOR2 (N4418, N4417, N1351);
and AND3 (N4419, N4409, N581, N833);
xor XOR2 (N4420, N4380, N4245);
not NOT1 (N4421, N4408);
or OR4 (N4422, N4410, N2839, N3706, N705);
xor XOR2 (N4423, N4418, N2332);
nand NAND2 (N4424, N4422, N1729);
buf BUF1 (N4425, N4423);
buf BUF1 (N4426, N4419);
not NOT1 (N4427, N4411);
and AND4 (N4428, N4426, N1566, N509, N4160);
nor NOR4 (N4429, N4421, N2950, N2949, N1813);
nand NAND3 (N4430, N4429, N1434, N3592);
buf BUF1 (N4431, N4430);
nand NAND4 (N4432, N4420, N3547, N765, N2491);
buf BUF1 (N4433, N4414);
nor NOR4 (N4434, N4416, N2233, N3906, N1469);
nand NAND4 (N4435, N4432, N3400, N3767, N992);
not NOT1 (N4436, N4435);
or OR2 (N4437, N4403, N2061);
nor NOR2 (N4438, N4424, N3125);
not NOT1 (N4439, N4438);
nand NAND3 (N4440, N4428, N3253, N255);
nor NOR2 (N4441, N4425, N3918);
not NOT1 (N4442, N4439);
xor XOR2 (N4443, N4415, N1590);
buf BUF1 (N4444, N4443);
nor NOR4 (N4445, N4437, N567, N1960, N3003);
not NOT1 (N4446, N4444);
and AND4 (N4447, N4436, N2542, N2247, N84);
and AND2 (N4448, N4433, N782);
xor XOR2 (N4449, N4446, N3009);
and AND3 (N4450, N4434, N475, N2309);
nor NOR4 (N4451, N4440, N1665, N703, N273);
or OR3 (N4452, N4441, N4272, N2229);
or OR4 (N4453, N4448, N3397, N2078, N3906);
nand NAND3 (N4454, N4450, N654, N3070);
or OR2 (N4455, N4453, N1925);
nor NOR3 (N4456, N4454, N584, N779);
not NOT1 (N4457, N4451);
xor XOR2 (N4458, N4455, N3942);
not NOT1 (N4459, N4458);
nand NAND2 (N4460, N4456, N3900);
nand NAND4 (N4461, N4449, N2168, N2586, N1691);
xor XOR2 (N4462, N4447, N3933);
buf BUF1 (N4463, N4461);
xor XOR2 (N4464, N4462, N1384);
nor NOR4 (N4465, N4452, N2749, N2708, N1907);
buf BUF1 (N4466, N4442);
and AND2 (N4467, N4459, N951);
or OR4 (N4468, N4464, N3076, N528, N2332);
nand NAND4 (N4469, N4467, N3075, N291, N2367);
nor NOR4 (N4470, N4457, N3829, N2665, N4469);
buf BUF1 (N4471, N2139);
or OR4 (N4472, N4465, N2244, N3479, N3512);
and AND4 (N4473, N4431, N2494, N2180, N2169);
xor XOR2 (N4474, N4472, N3709);
or OR3 (N4475, N4460, N3789, N2726);
or OR3 (N4476, N4427, N3121, N2742);
not NOT1 (N4477, N4445);
nand NAND2 (N4478, N4468, N221);
nor NOR2 (N4479, N4463, N3900);
buf BUF1 (N4480, N4473);
xor XOR2 (N4481, N4478, N3691);
xor XOR2 (N4482, N4475, N3141);
xor XOR2 (N4483, N4480, N91);
nor NOR3 (N4484, N4466, N1094, N4057);
not NOT1 (N4485, N4482);
not NOT1 (N4486, N4479);
xor XOR2 (N4487, N4481, N1397);
and AND4 (N4488, N4476, N1642, N287, N2693);
or OR4 (N4489, N4484, N371, N1837, N2482);
xor XOR2 (N4490, N4477, N3224);
nand NAND3 (N4491, N4490, N423, N4298);
nand NAND4 (N4492, N4471, N684, N1817, N21);
or OR2 (N4493, N4491, N4479);
or OR4 (N4494, N4474, N47, N2467, N1651);
nand NAND4 (N4495, N4493, N4032, N897, N913);
buf BUF1 (N4496, N4470);
and AND3 (N4497, N4489, N2508, N1787);
buf BUF1 (N4498, N4486);
not NOT1 (N4499, N4483);
and AND2 (N4500, N4485, N689);
buf BUF1 (N4501, N4487);
not NOT1 (N4502, N4497);
nor NOR2 (N4503, N4496, N3519);
not NOT1 (N4504, N4498);
or OR4 (N4505, N4503, N2235, N3308, N1495);
not NOT1 (N4506, N4500);
nand NAND4 (N4507, N4506, N906, N2144, N250);
not NOT1 (N4508, N4495);
or OR3 (N4509, N4488, N2204, N4350);
nand NAND4 (N4510, N4492, N1668, N2417, N1916);
and AND3 (N4511, N4499, N2348, N600);
nor NOR3 (N4512, N4504, N3953, N3283);
nor NOR3 (N4513, N4502, N3563, N3431);
and AND3 (N4514, N4505, N342, N156);
nor NOR4 (N4515, N4511, N734, N506, N3266);
nor NOR3 (N4516, N4508, N1270, N1100);
buf BUF1 (N4517, N4510);
nand NAND2 (N4518, N4517, N1153);
nor NOR4 (N4519, N4501, N3990, N3428, N2160);
nor NOR2 (N4520, N4494, N2057);
not NOT1 (N4521, N4507);
xor XOR2 (N4522, N4516, N3200);
xor XOR2 (N4523, N4520, N1644);
not NOT1 (N4524, N4515);
and AND2 (N4525, N4512, N3181);
nand NAND4 (N4526, N4521, N2480, N827, N3173);
xor XOR2 (N4527, N4526, N3868);
buf BUF1 (N4528, N4514);
xor XOR2 (N4529, N4523, N1520);
nand NAND4 (N4530, N4528, N3624, N4373, N32);
nor NOR2 (N4531, N4524, N1813);
and AND4 (N4532, N4525, N496, N4314, N1532);
xor XOR2 (N4533, N4509, N4279);
nor NOR2 (N4534, N4530, N370);
xor XOR2 (N4535, N4527, N2876);
or OR3 (N4536, N4532, N2574, N2352);
nand NAND2 (N4537, N4534, N2158);
nor NOR3 (N4538, N4535, N3724, N3351);
or OR3 (N4539, N4529, N1966, N3989);
not NOT1 (N4540, N4522);
not NOT1 (N4541, N4533);
and AND4 (N4542, N4537, N1017, N734, N55);
not NOT1 (N4543, N4513);
or OR3 (N4544, N4540, N3177, N3883);
nand NAND4 (N4545, N4536, N4252, N4428, N858);
and AND3 (N4546, N4543, N1239, N88);
and AND3 (N4547, N4545, N2618, N2610);
xor XOR2 (N4548, N4546, N1243);
not NOT1 (N4549, N4547);
xor XOR2 (N4550, N4541, N70);
xor XOR2 (N4551, N4519, N2642);
not NOT1 (N4552, N4531);
or OR2 (N4553, N4552, N2861);
xor XOR2 (N4554, N4549, N4075);
not NOT1 (N4555, N4548);
not NOT1 (N4556, N4544);
not NOT1 (N4557, N4550);
and AND2 (N4558, N4542, N687);
and AND2 (N4559, N4554, N1884);
and AND4 (N4560, N4551, N3263, N4348, N3816);
nand NAND3 (N4561, N4553, N1891, N953);
buf BUF1 (N4562, N4556);
or OR3 (N4563, N4559, N2065, N884);
and AND4 (N4564, N4539, N539, N1617, N181);
and AND2 (N4565, N4561, N2975);
buf BUF1 (N4566, N4557);
not NOT1 (N4567, N4558);
or OR4 (N4568, N4560, N4504, N3865, N3105);
or OR2 (N4569, N4538, N750);
not NOT1 (N4570, N4563);
nand NAND2 (N4571, N4518, N4130);
and AND2 (N4572, N4567, N4);
or OR2 (N4573, N4572, N3371);
not NOT1 (N4574, N4568);
buf BUF1 (N4575, N4566);
xor XOR2 (N4576, N4555, N1884);
xor XOR2 (N4577, N4576, N1256);
and AND2 (N4578, N4570, N1069);
buf BUF1 (N4579, N4571);
nand NAND4 (N4580, N4573, N1518, N1257, N76);
xor XOR2 (N4581, N4578, N2445);
or OR2 (N4582, N4569, N4440);
not NOT1 (N4583, N4579);
buf BUF1 (N4584, N4575);
buf BUF1 (N4585, N4584);
xor XOR2 (N4586, N4564, N46);
and AND4 (N4587, N4565, N3085, N3686, N1619);
and AND2 (N4588, N4586, N2407);
buf BUF1 (N4589, N4562);
or OR3 (N4590, N4574, N4298, N4256);
and AND4 (N4591, N4581, N2475, N2686, N1383);
and AND3 (N4592, N4582, N1019, N2136);
xor XOR2 (N4593, N4585, N4263);
buf BUF1 (N4594, N4591);
not NOT1 (N4595, N4580);
not NOT1 (N4596, N4588);
buf BUF1 (N4597, N4595);
and AND2 (N4598, N4587, N4461);
xor XOR2 (N4599, N4596, N1339);
or OR3 (N4600, N4593, N1772, N885);
nor NOR2 (N4601, N4599, N2776);
or OR4 (N4602, N4601, N2083, N3957, N4184);
buf BUF1 (N4603, N4577);
nand NAND4 (N4604, N4602, N4542, N2887, N1273);
nor NOR2 (N4605, N4600, N2660);
or OR3 (N4606, N4598, N2758, N2388);
nand NAND3 (N4607, N4606, N1310, N1997);
not NOT1 (N4608, N4583);
not NOT1 (N4609, N4589);
nor NOR4 (N4610, N4605, N2691, N142, N167);
nor NOR4 (N4611, N4603, N4109, N900, N1755);
and AND2 (N4612, N4611, N1472);
nand NAND2 (N4613, N4607, N4110);
xor XOR2 (N4614, N4609, N691);
nand NAND3 (N4615, N4604, N578, N216);
or OR2 (N4616, N4592, N4047);
or OR4 (N4617, N4597, N1261, N4596, N550);
nand NAND2 (N4618, N4610, N520);
and AND2 (N4619, N4613, N1477);
xor XOR2 (N4620, N4616, N1339);
not NOT1 (N4621, N4590);
xor XOR2 (N4622, N4615, N3920);
nand NAND2 (N4623, N4608, N277);
and AND4 (N4624, N4617, N4573, N689, N2551);
not NOT1 (N4625, N4624);
nand NAND4 (N4626, N4614, N418, N1157, N4135);
buf BUF1 (N4627, N4622);
buf BUF1 (N4628, N4626);
not NOT1 (N4629, N4625);
nand NAND2 (N4630, N4623, N432);
and AND3 (N4631, N4627, N1692, N3067);
xor XOR2 (N4632, N4630, N3726);
nand NAND4 (N4633, N4619, N4566, N1927, N3330);
and AND3 (N4634, N4629, N2864, N3615);
nor NOR3 (N4635, N4618, N3571, N3847);
nor NOR4 (N4636, N4631, N1991, N1571, N3937);
or OR2 (N4637, N4620, N4229);
nand NAND4 (N4638, N4621, N3169, N4403, N2250);
not NOT1 (N4639, N4634);
buf BUF1 (N4640, N4637);
xor XOR2 (N4641, N4628, N4302);
buf BUF1 (N4642, N4612);
or OR3 (N4643, N4633, N2796, N512);
not NOT1 (N4644, N4639);
nor NOR4 (N4645, N4644, N213, N416, N4308);
or OR3 (N4646, N4632, N1719, N1357);
not NOT1 (N4647, N4643);
nand NAND4 (N4648, N4645, N4427, N1537, N1228);
nand NAND4 (N4649, N4642, N3474, N2186, N1897);
not NOT1 (N4650, N4636);
xor XOR2 (N4651, N4650, N1790);
and AND3 (N4652, N4635, N4469, N217);
nand NAND4 (N4653, N4638, N1095, N2058, N2383);
xor XOR2 (N4654, N4653, N3716);
xor XOR2 (N4655, N4640, N529);
nand NAND4 (N4656, N4655, N3539, N4255, N4208);
not NOT1 (N4657, N4654);
nand NAND4 (N4658, N4648, N3990, N4493, N4188);
xor XOR2 (N4659, N4656, N1261);
or OR4 (N4660, N4652, N2475, N3642, N4129);
xor XOR2 (N4661, N4646, N1539);
not NOT1 (N4662, N4651);
xor XOR2 (N4663, N4660, N2877);
xor XOR2 (N4664, N4594, N586);
or OR3 (N4665, N4664, N2038, N1210);
not NOT1 (N4666, N4647);
nor NOR2 (N4667, N4663, N1591);
nor NOR3 (N4668, N4657, N2073, N3587);
or OR4 (N4669, N4661, N4422, N2685, N2237);
or OR4 (N4670, N4641, N3035, N3275, N3816);
nand NAND2 (N4671, N4667, N4026);
or OR2 (N4672, N4671, N2554);
nor NOR4 (N4673, N4669, N2670, N2282, N1767);
nor NOR4 (N4674, N4668, N4472, N2788, N4492);
or OR4 (N4675, N4662, N1785, N4310, N4218);
or OR3 (N4676, N4672, N2543, N1906);
nor NOR3 (N4677, N4670, N1829, N3447);
or OR4 (N4678, N4666, N4274, N3154, N2232);
buf BUF1 (N4679, N4675);
and AND4 (N4680, N4678, N779, N2455, N1778);
buf BUF1 (N4681, N4676);
nand NAND2 (N4682, N4681, N1834);
not NOT1 (N4683, N4679);
nor NOR2 (N4684, N4649, N3917);
not NOT1 (N4685, N4665);
xor XOR2 (N4686, N4684, N1976);
or OR4 (N4687, N4683, N769, N4242, N1039);
or OR3 (N4688, N4680, N1396, N2276);
nor NOR2 (N4689, N4686, N2381);
and AND3 (N4690, N4685, N2171, N786);
nor NOR3 (N4691, N4673, N2395, N1305);
nand NAND3 (N4692, N4688, N3368, N435);
or OR2 (N4693, N4674, N2);
not NOT1 (N4694, N4691);
xor XOR2 (N4695, N4693, N2171);
nor NOR3 (N4696, N4695, N4550, N390);
and AND2 (N4697, N4677, N411);
not NOT1 (N4698, N4694);
nand NAND2 (N4699, N4698, N2187);
nor NOR2 (N4700, N4697, N4220);
and AND2 (N4701, N4690, N3236);
xor XOR2 (N4702, N4701, N4046);
and AND4 (N4703, N4700, N3211, N764, N2372);
nand NAND3 (N4704, N4699, N4423, N343);
or OR2 (N4705, N4704, N1761);
buf BUF1 (N4706, N4659);
and AND4 (N4707, N4703, N3007, N1943, N577);
xor XOR2 (N4708, N4705, N3374);
or OR4 (N4709, N4687, N289, N3572, N2524);
and AND2 (N4710, N4702, N4163);
and AND2 (N4711, N4709, N4077);
nor NOR4 (N4712, N4711, N362, N2457, N1273);
not NOT1 (N4713, N4707);
xor XOR2 (N4714, N4710, N3100);
and AND3 (N4715, N4682, N1336, N3558);
not NOT1 (N4716, N4713);
nor NOR3 (N4717, N4658, N188, N2932);
nand NAND2 (N4718, N4715, N2865);
not NOT1 (N4719, N4708);
nand NAND2 (N4720, N4689, N3234);
nor NOR3 (N4721, N4720, N3975, N2411);
nor NOR3 (N4722, N4717, N4303, N2989);
nand NAND2 (N4723, N4716, N2204);
buf BUF1 (N4724, N4692);
xor XOR2 (N4725, N4696, N3787);
buf BUF1 (N4726, N4712);
not NOT1 (N4727, N4706);
or OR4 (N4728, N4718, N514, N2308, N3111);
or OR3 (N4729, N4719, N1172, N4274);
buf BUF1 (N4730, N4725);
and AND2 (N4731, N4723, N223);
not NOT1 (N4732, N4729);
nand NAND3 (N4733, N4730, N3479, N1788);
nor NOR4 (N4734, N4714, N869, N1471, N2662);
nand NAND4 (N4735, N4734, N373, N1575, N3362);
nand NAND2 (N4736, N4722, N1976);
and AND2 (N4737, N4735, N2791);
xor XOR2 (N4738, N4727, N3241);
nor NOR2 (N4739, N4733, N3387);
xor XOR2 (N4740, N4731, N967);
nand NAND4 (N4741, N4732, N446, N4611, N1090);
or OR2 (N4742, N4724, N128);
and AND4 (N4743, N4728, N231, N99, N2611);
and AND3 (N4744, N4741, N3185, N4364);
or OR4 (N4745, N4736, N1580, N1891, N2907);
buf BUF1 (N4746, N4739);
or OR3 (N4747, N4742, N202, N3009);
nand NAND3 (N4748, N4747, N2184, N1506);
not NOT1 (N4749, N4721);
nor NOR3 (N4750, N4737, N2027, N36);
and AND3 (N4751, N4726, N637, N1332);
and AND2 (N4752, N4740, N198);
nor NOR3 (N4753, N4745, N3294, N1181);
and AND4 (N4754, N4751, N850, N1196, N2805);
xor XOR2 (N4755, N4744, N1077);
buf BUF1 (N4756, N4755);
buf BUF1 (N4757, N4750);
nor NOR4 (N4758, N4748, N3222, N4368, N3462);
nor NOR4 (N4759, N4738, N1074, N3720, N3694);
buf BUF1 (N4760, N4746);
nand NAND4 (N4761, N4749, N2506, N1664, N24);
nor NOR2 (N4762, N4757, N4503);
not NOT1 (N4763, N4756);
buf BUF1 (N4764, N4758);
nor NOR2 (N4765, N4759, N2093);
nand NAND2 (N4766, N4764, N1814);
not NOT1 (N4767, N4763);
not NOT1 (N4768, N4762);
xor XOR2 (N4769, N4765, N2969);
nor NOR3 (N4770, N4768, N39, N1156);
nand NAND4 (N4771, N4766, N758, N580, N871);
nor NOR4 (N4772, N4754, N1851, N4204, N1585);
not NOT1 (N4773, N4760);
nand NAND3 (N4774, N4771, N3845, N3002);
or OR4 (N4775, N4774, N1438, N2665, N1311);
and AND2 (N4776, N4775, N2243);
nor NOR4 (N4777, N4767, N671, N820, N4609);
or OR2 (N4778, N4752, N1366);
not NOT1 (N4779, N4777);
nand NAND4 (N4780, N4776, N4600, N2674, N838);
not NOT1 (N4781, N4743);
buf BUF1 (N4782, N4770);
buf BUF1 (N4783, N4761);
nand NAND3 (N4784, N4783, N4187, N2186);
xor XOR2 (N4785, N4778, N4360);
and AND2 (N4786, N4784, N4259);
or OR3 (N4787, N4769, N719, N4333);
and AND3 (N4788, N4780, N4241, N2925);
not NOT1 (N4789, N4782);
not NOT1 (N4790, N4781);
nor NOR3 (N4791, N4785, N102, N3910);
or OR2 (N4792, N4773, N2312);
nor NOR3 (N4793, N4789, N260, N679);
buf BUF1 (N4794, N4772);
not NOT1 (N4795, N4787);
or OR4 (N4796, N4792, N2389, N3763, N2274);
nor NOR2 (N4797, N4779, N2663);
or OR2 (N4798, N4791, N809);
and AND2 (N4799, N4793, N4167);
nand NAND4 (N4800, N4786, N4310, N858, N3694);
buf BUF1 (N4801, N4794);
nor NOR2 (N4802, N4800, N931);
nor NOR4 (N4803, N4788, N812, N2369, N4593);
not NOT1 (N4804, N4753);
and AND3 (N4805, N4795, N2542, N3305);
buf BUF1 (N4806, N4805);
and AND3 (N4807, N4804, N3669, N4147);
nand NAND3 (N4808, N4790, N1421, N4167);
nand NAND3 (N4809, N4806, N3710, N2283);
xor XOR2 (N4810, N4796, N630);
and AND2 (N4811, N4809, N3058);
xor XOR2 (N4812, N4801, N476);
and AND3 (N4813, N4802, N2339, N2409);
and AND2 (N4814, N4797, N4070);
nor NOR3 (N4815, N4814, N729, N3196);
not NOT1 (N4816, N4799);
buf BUF1 (N4817, N4813);
not NOT1 (N4818, N4807);
or OR2 (N4819, N4798, N4665);
or OR3 (N4820, N4810, N3275, N1617);
or OR4 (N4821, N4815, N3424, N2861, N1837);
not NOT1 (N4822, N4803);
or OR2 (N4823, N4820, N4281);
and AND2 (N4824, N4816, N3121);
not NOT1 (N4825, N4824);
buf BUF1 (N4826, N4812);
nand NAND4 (N4827, N4808, N2609, N3066, N669);
or OR3 (N4828, N4811, N441, N4470);
buf BUF1 (N4829, N4817);
nor NOR3 (N4830, N4823, N2463, N1273);
and AND2 (N4831, N4828, N3354);
nand NAND4 (N4832, N4818, N1818, N2028, N1227);
not NOT1 (N4833, N4827);
buf BUF1 (N4834, N4821);
buf BUF1 (N4835, N4825);
xor XOR2 (N4836, N4831, N4580);
xor XOR2 (N4837, N4819, N1192);
nand NAND4 (N4838, N4834, N2411, N1888, N3221);
and AND3 (N4839, N4835, N3512, N1410);
buf BUF1 (N4840, N4826);
or OR4 (N4841, N4829, N2588, N2394, N3697);
and AND2 (N4842, N4833, N425);
not NOT1 (N4843, N4838);
nand NAND4 (N4844, N4843, N2491, N1754, N407);
nand NAND2 (N4845, N4832, N262);
xor XOR2 (N4846, N4836, N694);
or OR4 (N4847, N4841, N412, N4091, N2667);
nand NAND3 (N4848, N4830, N378, N3299);
not NOT1 (N4849, N4840);
not NOT1 (N4850, N4847);
and AND2 (N4851, N4837, N3607);
or OR3 (N4852, N4842, N4200, N311);
not NOT1 (N4853, N4839);
not NOT1 (N4854, N4848);
xor XOR2 (N4855, N4845, N1244);
nand NAND3 (N4856, N4853, N4731, N1425);
nor NOR3 (N4857, N4849, N133, N1831);
nand NAND2 (N4858, N4857, N2757);
nor NOR4 (N4859, N4858, N4172, N1873, N2843);
nor NOR3 (N4860, N4859, N2736, N1987);
and AND3 (N4861, N4860, N913, N2655);
buf BUF1 (N4862, N4861);
xor XOR2 (N4863, N4844, N3768);
nor NOR4 (N4864, N4854, N4828, N2798, N3778);
nand NAND3 (N4865, N4822, N3173, N2380);
not NOT1 (N4866, N4863);
and AND2 (N4867, N4862, N2530);
or OR2 (N4868, N4846, N4367);
xor XOR2 (N4869, N4867, N4311);
and AND2 (N4870, N4864, N1720);
nand NAND2 (N4871, N4850, N132);
or OR4 (N4872, N4865, N793, N2139, N3697);
nand NAND3 (N4873, N4870, N1320, N1135);
nand NAND3 (N4874, N4872, N3909, N1620);
or OR2 (N4875, N4851, N409);
nand NAND4 (N4876, N4874, N1913, N3373, N363);
buf BUF1 (N4877, N4871);
not NOT1 (N4878, N4876);
not NOT1 (N4879, N4878);
or OR3 (N4880, N4877, N1142, N4077);
nor NOR3 (N4881, N4875, N2757, N3195);
buf BUF1 (N4882, N4866);
xor XOR2 (N4883, N4852, N654);
xor XOR2 (N4884, N4883, N3815);
and AND3 (N4885, N4855, N3320, N1187);
buf BUF1 (N4886, N4884);
xor XOR2 (N4887, N4856, N1788);
xor XOR2 (N4888, N4881, N973);
or OR2 (N4889, N4868, N2607);
and AND2 (N4890, N4885, N690);
or OR4 (N4891, N4890, N801, N240, N4859);
buf BUF1 (N4892, N4891);
not NOT1 (N4893, N4886);
not NOT1 (N4894, N4889);
and AND2 (N4895, N4873, N1507);
and AND2 (N4896, N4892, N4516);
buf BUF1 (N4897, N4895);
nand NAND2 (N4898, N4894, N2781);
nand NAND4 (N4899, N4880, N2360, N912, N2014);
nand NAND3 (N4900, N4897, N415, N4214);
or OR4 (N4901, N4900, N2621, N3418, N430);
nor NOR2 (N4902, N4899, N1833);
nor NOR4 (N4903, N4882, N1617, N3749, N3862);
nand NAND4 (N4904, N4903, N1553, N2236, N1968);
and AND4 (N4905, N4896, N1375, N1533, N85);
nor NOR3 (N4906, N4905, N2559, N3075);
not NOT1 (N4907, N4902);
buf BUF1 (N4908, N4906);
and AND2 (N4909, N4904, N4825);
and AND4 (N4910, N4888, N2957, N3839, N1297);
or OR2 (N4911, N4887, N157);
nand NAND3 (N4912, N4879, N4832, N295);
and AND3 (N4913, N4893, N2751, N4508);
and AND3 (N4914, N4869, N502, N1858);
not NOT1 (N4915, N4901);
nor NOR3 (N4916, N4915, N3021, N4083);
nor NOR3 (N4917, N4907, N2447, N2664);
and AND4 (N4918, N4910, N4506, N3074, N4064);
buf BUF1 (N4919, N4918);
nor NOR3 (N4920, N4913, N3349, N4658);
nor NOR2 (N4921, N4914, N368);
and AND2 (N4922, N4921, N3976);
not NOT1 (N4923, N4920);
nor NOR3 (N4924, N4909, N1086, N4082);
not NOT1 (N4925, N4912);
nand NAND3 (N4926, N4925, N1983, N4350);
not NOT1 (N4927, N4916);
not NOT1 (N4928, N4898);
buf BUF1 (N4929, N4924);
and AND3 (N4930, N4927, N4290, N1262);
nor NOR3 (N4931, N4911, N2125, N3567);
not NOT1 (N4932, N4923);
buf BUF1 (N4933, N4932);
xor XOR2 (N4934, N4926, N344);
not NOT1 (N4935, N4922);
buf BUF1 (N4936, N4935);
nor NOR2 (N4937, N4933, N4279);
nand NAND4 (N4938, N4908, N157, N3276, N918);
buf BUF1 (N4939, N4937);
or OR2 (N4940, N4938, N392);
buf BUF1 (N4941, N4928);
nor NOR2 (N4942, N4934, N613);
nor NOR4 (N4943, N4930, N2302, N2949, N4032);
nand NAND2 (N4944, N4941, N2006);
buf BUF1 (N4945, N4919);
buf BUF1 (N4946, N4936);
xor XOR2 (N4947, N4944, N1835);
nor NOR2 (N4948, N4939, N4352);
and AND4 (N4949, N4948, N552, N1340, N3269);
nor NOR4 (N4950, N4931, N4613, N3244, N3112);
or OR2 (N4951, N4943, N2182);
or OR4 (N4952, N4945, N172, N3760, N2620);
nor NOR3 (N4953, N4929, N2418, N1749);
nor NOR3 (N4954, N4946, N4775, N4682);
or OR2 (N4955, N4952, N4072);
and AND2 (N4956, N4940, N4652);
nand NAND2 (N4957, N4949, N1536);
buf BUF1 (N4958, N4950);
or OR4 (N4959, N4917, N3010, N2520, N3984);
not NOT1 (N4960, N4957);
nor NOR2 (N4961, N4958, N729);
not NOT1 (N4962, N4942);
nor NOR2 (N4963, N4962, N3095);
or OR4 (N4964, N4953, N4686, N1426, N1918);
xor XOR2 (N4965, N4951, N3725);
buf BUF1 (N4966, N4960);
or OR3 (N4967, N4961, N2717, N2435);
or OR3 (N4968, N4964, N4337, N403);
and AND2 (N4969, N4965, N3760);
nor NOR4 (N4970, N4967, N3383, N3508, N2199);
nor NOR3 (N4971, N4970, N2935, N2322);
nor NOR3 (N4972, N4947, N4856, N3009);
and AND2 (N4973, N4956, N91);
buf BUF1 (N4974, N4955);
and AND2 (N4975, N4966, N2175);
buf BUF1 (N4976, N4954);
nor NOR4 (N4977, N4959, N2902, N4519, N2043);
and AND4 (N4978, N4975, N3788, N1812, N3495);
nor NOR4 (N4979, N4969, N4027, N1595, N4513);
buf BUF1 (N4980, N4978);
or OR3 (N4981, N4963, N1245, N1096);
not NOT1 (N4982, N4979);
nand NAND3 (N4983, N4972, N4543, N4266);
nor NOR3 (N4984, N4982, N2164, N2916);
nor NOR4 (N4985, N4981, N2194, N4047, N2016);
not NOT1 (N4986, N4976);
nor NOR2 (N4987, N4985, N2126);
nand NAND2 (N4988, N4968, N2919);
buf BUF1 (N4989, N4980);
and AND3 (N4990, N4977, N145, N549);
buf BUF1 (N4991, N4990);
xor XOR2 (N4992, N4989, N3237);
xor XOR2 (N4993, N4992, N2786);
nand NAND3 (N4994, N4991, N328, N775);
or OR2 (N4995, N4988, N4681);
and AND4 (N4996, N4994, N4504, N4444, N2200);
xor XOR2 (N4997, N4995, N269);
nand NAND2 (N4998, N4971, N2231);
nand NAND4 (N4999, N4997, N1208, N2097, N4112);
nand NAND4 (N5000, N4986, N4240, N108, N2229);
not NOT1 (N5001, N4974);
xor XOR2 (N5002, N5001, N1960);
not NOT1 (N5003, N5002);
and AND2 (N5004, N4983, N4983);
buf BUF1 (N5005, N5003);
xor XOR2 (N5006, N4973, N3959);
not NOT1 (N5007, N4987);
buf BUF1 (N5008, N5000);
nor NOR2 (N5009, N5005, N1338);
nand NAND2 (N5010, N5007, N2250);
not NOT1 (N5011, N4993);
and AND2 (N5012, N5006, N4348);
or OR3 (N5013, N5009, N4981, N995);
nand NAND2 (N5014, N4998, N1890);
not NOT1 (N5015, N5008);
xor XOR2 (N5016, N5012, N2234);
not NOT1 (N5017, N5004);
nor NOR2 (N5018, N5017, N3987);
nand NAND2 (N5019, N5018, N1156);
nor NOR4 (N5020, N5015, N3929, N1575, N2785);
nand NAND2 (N5021, N4996, N3468);
and AND4 (N5022, N5016, N65, N1195, N1275);
buf BUF1 (N5023, N5020);
buf BUF1 (N5024, N5022);
nand NAND4 (N5025, N5021, N4097, N3614, N3441);
nor NOR3 (N5026, N5013, N849, N2791);
and AND3 (N5027, N4984, N149, N4428);
nor NOR2 (N5028, N5025, N4883);
or OR2 (N5029, N5010, N1230);
nor NOR2 (N5030, N5023, N107);
nand NAND4 (N5031, N4999, N4060, N4507, N4012);
buf BUF1 (N5032, N5031);
nand NAND4 (N5033, N5029, N4848, N2243, N2839);
buf BUF1 (N5034, N5024);
xor XOR2 (N5035, N5033, N4578);
nor NOR4 (N5036, N5032, N2563, N2362, N1913);
not NOT1 (N5037, N5026);
nor NOR3 (N5038, N5011, N4143, N2862);
nor NOR3 (N5039, N5036, N1228, N4347);
and AND3 (N5040, N5034, N93, N3706);
xor XOR2 (N5041, N5038, N1557);
not NOT1 (N5042, N5040);
nand NAND3 (N5043, N5039, N3985, N1331);
nor NOR4 (N5044, N5042, N3067, N4083, N603);
and AND2 (N5045, N5037, N611);
nor NOR2 (N5046, N5030, N4645);
nor NOR3 (N5047, N5041, N3879, N4024);
not NOT1 (N5048, N5035);
or OR3 (N5049, N5028, N1986, N2979);
not NOT1 (N5050, N5044);
not NOT1 (N5051, N5049);
nand NAND4 (N5052, N5047, N3158, N774, N957);
and AND4 (N5053, N5043, N1162, N720, N4476);
and AND4 (N5054, N5048, N4113, N4128, N4697);
not NOT1 (N5055, N5046);
or OR4 (N5056, N5051, N43, N48, N526);
buf BUF1 (N5057, N5045);
and AND2 (N5058, N5054, N917);
buf BUF1 (N5059, N5053);
or OR3 (N5060, N5014, N876, N47);
or OR3 (N5061, N5056, N745, N1924);
nand NAND2 (N5062, N5052, N4349);
and AND4 (N5063, N5057, N3371, N2203, N1461);
not NOT1 (N5064, N5061);
and AND2 (N5065, N5060, N5006);
nor NOR3 (N5066, N5055, N1781, N3498);
buf BUF1 (N5067, N5050);
xor XOR2 (N5068, N5027, N4758);
and AND3 (N5069, N5058, N3281, N2375);
nor NOR2 (N5070, N5069, N769);
nand NAND3 (N5071, N5066, N3008, N2007);
and AND4 (N5072, N5019, N180, N2962, N1252);
and AND2 (N5073, N5071, N2309);
not NOT1 (N5074, N5068);
xor XOR2 (N5075, N5063, N1678);
xor XOR2 (N5076, N5072, N3004);
not NOT1 (N5077, N5062);
buf BUF1 (N5078, N5076);
xor XOR2 (N5079, N5067, N2348);
buf BUF1 (N5080, N5074);
not NOT1 (N5081, N5064);
nand NAND3 (N5082, N5078, N3491, N3659);
not NOT1 (N5083, N5081);
nor NOR4 (N5084, N5082, N111, N1971, N1459);
nor NOR3 (N5085, N5075, N3550, N4302);
buf BUF1 (N5086, N5079);
buf BUF1 (N5087, N5059);
buf BUF1 (N5088, N5083);
or OR3 (N5089, N5080, N4024, N3397);
buf BUF1 (N5090, N5089);
or OR3 (N5091, N5087, N3533, N3553);
xor XOR2 (N5092, N5091, N4139);
nor NOR3 (N5093, N5085, N4837, N4703);
xor XOR2 (N5094, N5093, N3918);
not NOT1 (N5095, N5094);
xor XOR2 (N5096, N5086, N352);
nor NOR4 (N5097, N5065, N4605, N2442, N321);
nand NAND4 (N5098, N5088, N3080, N1568, N4424);
not NOT1 (N5099, N5098);
nor NOR2 (N5100, N5097, N4393);
nand NAND4 (N5101, N5100, N4357, N2398, N2695);
and AND4 (N5102, N5096, N4654, N4381, N4485);
nor NOR3 (N5103, N5073, N4737, N3705);
or OR2 (N5104, N5095, N3512);
and AND2 (N5105, N5104, N3675);
nor NOR2 (N5106, N5099, N4077);
or OR2 (N5107, N5106, N445);
or OR4 (N5108, N5102, N811, N4486, N3159);
nor NOR2 (N5109, N5103, N2126);
nor NOR2 (N5110, N5105, N2544);
not NOT1 (N5111, N5108);
xor XOR2 (N5112, N5084, N1101);
buf BUF1 (N5113, N5110);
nor NOR2 (N5114, N5111, N3403);
and AND4 (N5115, N5092, N2629, N2813, N1071);
xor XOR2 (N5116, N5112, N2564);
nand NAND3 (N5117, N5090, N2713, N2194);
not NOT1 (N5118, N5107);
nor NOR2 (N5119, N5113, N3064);
xor XOR2 (N5120, N5101, N4544);
nand NAND4 (N5121, N5070, N74, N1441, N1141);
or OR2 (N5122, N5118, N4394);
nor NOR2 (N5123, N5122, N4836);
or OR3 (N5124, N5115, N4450, N1252);
or OR2 (N5125, N5123, N4138);
nor NOR3 (N5126, N5125, N936, N3024);
nor NOR3 (N5127, N5126, N2490, N4735);
or OR3 (N5128, N5117, N4411, N1509);
buf BUF1 (N5129, N5128);
buf BUF1 (N5130, N5114);
not NOT1 (N5131, N5130);
nor NOR2 (N5132, N5129, N4131);
and AND4 (N5133, N5121, N3993, N4599, N1463);
buf BUF1 (N5134, N5131);
and AND2 (N5135, N5133, N4349);
not NOT1 (N5136, N5132);
xor XOR2 (N5137, N5120, N1766);
buf BUF1 (N5138, N5136);
xor XOR2 (N5139, N5124, N2777);
or OR2 (N5140, N5119, N1358);
buf BUF1 (N5141, N5135);
nand NAND2 (N5142, N5137, N1216);
or OR3 (N5143, N5134, N4950, N2259);
and AND3 (N5144, N5143, N4455, N3772);
or OR4 (N5145, N5116, N2087, N3344, N1098);
or OR4 (N5146, N5077, N1753, N4947, N4567);
and AND2 (N5147, N5138, N188);
buf BUF1 (N5148, N5141);
not NOT1 (N5149, N5109);
not NOT1 (N5150, N5139);
nand NAND4 (N5151, N5140, N3851, N2598, N1331);
buf BUF1 (N5152, N5147);
and AND4 (N5153, N5145, N1049, N2470, N3794);
and AND3 (N5154, N5127, N358, N4177);
or OR2 (N5155, N5144, N2887);
buf BUF1 (N5156, N5153);
buf BUF1 (N5157, N5142);
nor NOR4 (N5158, N5156, N270, N4179, N1703);
and AND2 (N5159, N5157, N542);
and AND4 (N5160, N5149, N4353, N1440, N4210);
nand NAND3 (N5161, N5150, N2446, N854);
nand NAND2 (N5162, N5160, N2504);
nor NOR4 (N5163, N5155, N1244, N2440, N760);
or OR4 (N5164, N5163, N5119, N1292, N3903);
xor XOR2 (N5165, N5162, N2680);
nor NOR4 (N5166, N5154, N2214, N3052, N4240);
and AND4 (N5167, N5164, N212, N4466, N2127);
nor NOR2 (N5168, N5151, N186);
nand NAND2 (N5169, N5168, N616);
nor NOR3 (N5170, N5166, N2382, N2738);
xor XOR2 (N5171, N5152, N1306);
nand NAND2 (N5172, N5167, N4537);
nor NOR2 (N5173, N5169, N1972);
nor NOR4 (N5174, N5159, N2067, N4707, N4518);
not NOT1 (N5175, N5172);
nor NOR4 (N5176, N5170, N4093, N2801, N3249);
xor XOR2 (N5177, N5158, N1322);
not NOT1 (N5178, N5165);
not NOT1 (N5179, N5176);
xor XOR2 (N5180, N5173, N2375);
not NOT1 (N5181, N5180);
not NOT1 (N5182, N5181);
or OR3 (N5183, N5161, N3918, N3423);
or OR3 (N5184, N5177, N1310, N1665);
buf BUF1 (N5185, N5178);
not NOT1 (N5186, N5182);
nand NAND4 (N5187, N5186, N1256, N2449, N3345);
nand NAND3 (N5188, N5183, N3974, N602);
buf BUF1 (N5189, N5188);
nand NAND2 (N5190, N5187, N2935);
and AND2 (N5191, N5190, N4118);
nand NAND2 (N5192, N5184, N2732);
buf BUF1 (N5193, N5192);
nor NOR4 (N5194, N5148, N1173, N3774, N1154);
buf BUF1 (N5195, N5175);
nand NAND2 (N5196, N5185, N2651);
and AND3 (N5197, N5194, N2116, N171);
not NOT1 (N5198, N5193);
nor NOR3 (N5199, N5171, N4373, N831);
nor NOR3 (N5200, N5179, N4137, N1313);
nor NOR3 (N5201, N5199, N2678, N2799);
xor XOR2 (N5202, N5200, N2397);
nor NOR3 (N5203, N5191, N2791, N2047);
buf BUF1 (N5204, N5203);
or OR4 (N5205, N5189, N2179, N1686, N3508);
buf BUF1 (N5206, N5205);
nand NAND3 (N5207, N5201, N394, N1880);
xor XOR2 (N5208, N5202, N4740);
buf BUF1 (N5209, N5206);
buf BUF1 (N5210, N5195);
xor XOR2 (N5211, N5204, N4605);
nor NOR2 (N5212, N5211, N2941);
and AND3 (N5213, N5174, N413, N4179);
nor NOR4 (N5214, N5208, N4239, N1325, N2525);
not NOT1 (N5215, N5196);
and AND3 (N5216, N5212, N2911, N2435);
xor XOR2 (N5217, N5215, N1513);
not NOT1 (N5218, N5197);
nand NAND2 (N5219, N5210, N3079);
buf BUF1 (N5220, N5213);
nand NAND2 (N5221, N5146, N3643);
or OR4 (N5222, N5216, N2868, N3990, N4600);
xor XOR2 (N5223, N5222, N2710);
xor XOR2 (N5224, N5220, N1526);
nand NAND3 (N5225, N5217, N374, N1717);
and AND2 (N5226, N5219, N768);
xor XOR2 (N5227, N5224, N3626);
not NOT1 (N5228, N5198);
nor NOR3 (N5229, N5221, N3169, N4714);
and AND2 (N5230, N5226, N5103);
xor XOR2 (N5231, N5225, N4711);
not NOT1 (N5232, N5209);
or OR3 (N5233, N5223, N1119, N3565);
and AND3 (N5234, N5218, N100, N3410);
and AND4 (N5235, N5228, N3019, N4561, N291);
and AND4 (N5236, N5232, N2640, N128, N857);
xor XOR2 (N5237, N5229, N2187);
and AND2 (N5238, N5234, N2413);
or OR4 (N5239, N5238, N3784, N4289, N1975);
not NOT1 (N5240, N5207);
xor XOR2 (N5241, N5231, N5146);
nor NOR2 (N5242, N5235, N4810);
xor XOR2 (N5243, N5240, N3910);
xor XOR2 (N5244, N5230, N4877);
nand NAND2 (N5245, N5237, N602);
and AND3 (N5246, N5241, N3188, N1000);
xor XOR2 (N5247, N5239, N3728);
nor NOR2 (N5248, N5244, N2239);
and AND4 (N5249, N5246, N3266, N2408, N2464);
buf BUF1 (N5250, N5247);
not NOT1 (N5251, N5236);
or OR3 (N5252, N5251, N2878, N428);
or OR2 (N5253, N5242, N256);
or OR4 (N5254, N5248, N2331, N2189, N4602);
not NOT1 (N5255, N5254);
buf BUF1 (N5256, N5214);
nor NOR2 (N5257, N5227, N3335);
and AND4 (N5258, N5257, N5244, N2649, N1386);
or OR4 (N5259, N5258, N1620, N2769, N5174);
buf BUF1 (N5260, N5243);
nand NAND2 (N5261, N5256, N3204);
and AND3 (N5262, N5259, N4067, N730);
buf BUF1 (N5263, N5262);
nand NAND2 (N5264, N5260, N3234);
nor NOR3 (N5265, N5249, N3940, N4081);
buf BUF1 (N5266, N5255);
or OR3 (N5267, N5263, N274, N4582);
xor XOR2 (N5268, N5245, N4273);
nor NOR4 (N5269, N5252, N2794, N4781, N393);
xor XOR2 (N5270, N5268, N3109);
and AND3 (N5271, N5267, N880, N56);
or OR3 (N5272, N5250, N1002, N1858);
xor XOR2 (N5273, N5271, N801);
not NOT1 (N5274, N5270);
xor XOR2 (N5275, N5266, N2993);
xor XOR2 (N5276, N5233, N80);
and AND2 (N5277, N5274, N2358);
or OR3 (N5278, N5269, N1920, N4342);
not NOT1 (N5279, N5273);
nand NAND2 (N5280, N5253, N4795);
or OR3 (N5281, N5277, N2841, N1013);
not NOT1 (N5282, N5276);
and AND2 (N5283, N5281, N3121);
not NOT1 (N5284, N5265);
nor NOR4 (N5285, N5283, N368, N2318, N3680);
and AND2 (N5286, N5261, N1464);
xor XOR2 (N5287, N5286, N4235);
nand NAND3 (N5288, N5285, N2787, N649);
buf BUF1 (N5289, N5279);
and AND3 (N5290, N5275, N3370, N2838);
xor XOR2 (N5291, N5280, N2725);
buf BUF1 (N5292, N5287);
and AND3 (N5293, N5292, N2081, N4583);
or OR4 (N5294, N5278, N2131, N4488, N803);
and AND4 (N5295, N5282, N2036, N5071, N2329);
and AND2 (N5296, N5294, N5108);
nor NOR4 (N5297, N5290, N1942, N2013, N2007);
nand NAND4 (N5298, N5297, N3562, N1115, N1657);
and AND3 (N5299, N5272, N1627, N196);
nor NOR3 (N5300, N5295, N1747, N4558);
not NOT1 (N5301, N5299);
xor XOR2 (N5302, N5288, N3159);
not NOT1 (N5303, N5284);
or OR3 (N5304, N5302, N2285, N4057);
xor XOR2 (N5305, N5304, N3017);
xor XOR2 (N5306, N5298, N173);
nor NOR4 (N5307, N5303, N4706, N1653, N2914);
not NOT1 (N5308, N5296);
or OR3 (N5309, N5301, N3505, N4439);
nor NOR3 (N5310, N5293, N2872, N4192);
or OR4 (N5311, N5305, N4085, N4082, N1905);
nand NAND2 (N5312, N5289, N1457);
xor XOR2 (N5313, N5264, N5291);
xor XOR2 (N5314, N5275, N4840);
not NOT1 (N5315, N5306);
xor XOR2 (N5316, N5309, N5006);
or OR2 (N5317, N5308, N4889);
nor NOR4 (N5318, N5300, N3026, N327, N3553);
nor NOR3 (N5319, N5307, N4008, N240);
not NOT1 (N5320, N5313);
buf BUF1 (N5321, N5319);
xor XOR2 (N5322, N5321, N1705);
nand NAND3 (N5323, N5320, N4452, N1617);
and AND4 (N5324, N5310, N96, N75, N4926);
and AND3 (N5325, N5322, N5171, N2844);
nand NAND3 (N5326, N5312, N2052, N892);
nor NOR4 (N5327, N5326, N1277, N4996, N5319);
and AND2 (N5328, N5311, N2366);
xor XOR2 (N5329, N5316, N4577);
or OR3 (N5330, N5328, N449, N4528);
not NOT1 (N5331, N5330);
xor XOR2 (N5332, N5323, N2124);
nor NOR4 (N5333, N5332, N141, N2221, N2768);
xor XOR2 (N5334, N5329, N1620);
not NOT1 (N5335, N5317);
nand NAND2 (N5336, N5315, N5197);
xor XOR2 (N5337, N5333, N3540);
nor NOR4 (N5338, N5336, N4989, N1396, N3192);
or OR2 (N5339, N5331, N3428);
or OR4 (N5340, N5337, N460, N153, N1506);
not NOT1 (N5341, N5334);
nand NAND4 (N5342, N5324, N3101, N1394, N4023);
not NOT1 (N5343, N5341);
nand NAND2 (N5344, N5338, N4433);
and AND3 (N5345, N5342, N2178, N3953);
nor NOR2 (N5346, N5343, N2937);
nor NOR2 (N5347, N5314, N4521);
xor XOR2 (N5348, N5344, N3953);
nand NAND4 (N5349, N5348, N3854, N2437, N1700);
or OR4 (N5350, N5340, N2867, N4399, N841);
and AND4 (N5351, N5350, N1097, N764, N5090);
or OR4 (N5352, N5325, N2897, N4564, N2788);
nand NAND4 (N5353, N5347, N4672, N726, N734);
nor NOR4 (N5354, N5339, N5012, N1769, N3119);
nand NAND2 (N5355, N5327, N3199);
nand NAND2 (N5356, N5352, N4540);
not NOT1 (N5357, N5335);
nand NAND3 (N5358, N5351, N2133, N3648);
or OR3 (N5359, N5356, N435, N3768);
nand NAND4 (N5360, N5355, N1373, N4865, N849);
nand NAND4 (N5361, N5360, N3276, N2639, N4376);
and AND4 (N5362, N5318, N5090, N4900, N2179);
and AND2 (N5363, N5358, N659);
and AND4 (N5364, N5357, N4125, N4590, N3948);
xor XOR2 (N5365, N5346, N4099);
or OR4 (N5366, N5345, N1105, N4233, N1132);
buf BUF1 (N5367, N5349);
or OR3 (N5368, N5353, N3371, N1103);
not NOT1 (N5369, N5364);
xor XOR2 (N5370, N5365, N381);
nor NOR3 (N5371, N5366, N1977, N5245);
or OR4 (N5372, N5354, N4440, N2781, N3201);
and AND4 (N5373, N5368, N5330, N2240, N1513);
buf BUF1 (N5374, N5370);
not NOT1 (N5375, N5369);
buf BUF1 (N5376, N5371);
nor NOR4 (N5377, N5367, N3440, N1959, N4421);
buf BUF1 (N5378, N5372);
and AND4 (N5379, N5363, N424, N1110, N4429);
or OR3 (N5380, N5374, N5256, N4133);
and AND3 (N5381, N5379, N3548, N150);
not NOT1 (N5382, N5373);
or OR4 (N5383, N5359, N2709, N3738, N2510);
or OR4 (N5384, N5378, N3334, N3508, N320);
nor NOR2 (N5385, N5375, N2477);
not NOT1 (N5386, N5380);
and AND2 (N5387, N5383, N5159);
buf BUF1 (N5388, N5377);
nand NAND2 (N5389, N5361, N1234);
xor XOR2 (N5390, N5362, N261);
buf BUF1 (N5391, N5376);
nor NOR3 (N5392, N5387, N2661, N4058);
and AND3 (N5393, N5382, N309, N4101);
or OR4 (N5394, N5386, N261, N2885, N5061);
nor NOR2 (N5395, N5384, N4361);
not NOT1 (N5396, N5391);
nand NAND3 (N5397, N5393, N1900, N1880);
not NOT1 (N5398, N5395);
or OR3 (N5399, N5381, N4521, N1282);
nor NOR2 (N5400, N5396, N1602);
and AND4 (N5401, N5394, N2932, N3150, N635);
or OR4 (N5402, N5385, N3647, N2298, N3665);
nor NOR2 (N5403, N5392, N1227);
not NOT1 (N5404, N5390);
buf BUF1 (N5405, N5399);
or OR4 (N5406, N5404, N2503, N4546, N1339);
nor NOR2 (N5407, N5402, N1741);
buf BUF1 (N5408, N5401);
buf BUF1 (N5409, N5405);
buf BUF1 (N5410, N5397);
and AND2 (N5411, N5388, N1159);
nor NOR4 (N5412, N5408, N657, N800, N970);
or OR2 (N5413, N5412, N5364);
xor XOR2 (N5414, N5407, N1904);
nor NOR4 (N5415, N5400, N3331, N1998, N3569);
and AND3 (N5416, N5389, N149, N5174);
not NOT1 (N5417, N5415);
not NOT1 (N5418, N5413);
not NOT1 (N5419, N5418);
or OR3 (N5420, N5410, N2224, N3084);
or OR3 (N5421, N5419, N1653, N2419);
or OR4 (N5422, N5414, N406, N1835, N3724);
nor NOR2 (N5423, N5411, N3997);
buf BUF1 (N5424, N5422);
and AND3 (N5425, N5423, N3243, N4974);
nand NAND3 (N5426, N5409, N642, N1764);
and AND2 (N5427, N5426, N3859);
and AND3 (N5428, N5403, N941, N1707);
nor NOR4 (N5429, N5427, N1288, N3971, N960);
nor NOR2 (N5430, N5406, N5415);
and AND4 (N5431, N5424, N2919, N3272, N4320);
xor XOR2 (N5432, N5429, N784);
nand NAND3 (N5433, N5430, N4226, N3255);
and AND4 (N5434, N5417, N646, N535, N1854);
or OR4 (N5435, N5398, N3449, N5042, N5045);
nand NAND4 (N5436, N5421, N3045, N1590, N1294);
nor NOR2 (N5437, N5428, N649);
or OR3 (N5438, N5434, N778, N4021);
xor XOR2 (N5439, N5431, N1269);
nor NOR4 (N5440, N5435, N2273, N1458, N3464);
nor NOR3 (N5441, N5432, N2543, N2538);
not NOT1 (N5442, N5416);
nand NAND2 (N5443, N5438, N4349);
nand NAND2 (N5444, N5440, N3540);
xor XOR2 (N5445, N5444, N651);
and AND2 (N5446, N5436, N2157);
not NOT1 (N5447, N5443);
and AND2 (N5448, N5446, N2323);
buf BUF1 (N5449, N5447);
and AND2 (N5450, N5433, N1023);
not NOT1 (N5451, N5445);
and AND2 (N5452, N5450, N1674);
nor NOR3 (N5453, N5448, N3913, N355);
not NOT1 (N5454, N5420);
and AND4 (N5455, N5442, N5395, N3018, N4428);
nor NOR4 (N5456, N5454, N1119, N24, N1959);
xor XOR2 (N5457, N5453, N5294);
buf BUF1 (N5458, N5441);
not NOT1 (N5459, N5455);
buf BUF1 (N5460, N5425);
not NOT1 (N5461, N5458);
not NOT1 (N5462, N5461);
nand NAND3 (N5463, N5451, N4814, N3933);
not NOT1 (N5464, N5437);
not NOT1 (N5465, N5460);
or OR2 (N5466, N5463, N4380);
and AND2 (N5467, N5462, N3623);
or OR2 (N5468, N5457, N568);
xor XOR2 (N5469, N5459, N1203);
not NOT1 (N5470, N5468);
xor XOR2 (N5471, N5466, N111);
nor NOR4 (N5472, N5467, N4158, N473, N1225);
buf BUF1 (N5473, N5449);
buf BUF1 (N5474, N5439);
not NOT1 (N5475, N5472);
nor NOR3 (N5476, N5470, N4189, N2914);
nand NAND3 (N5477, N5475, N5028, N2240);
xor XOR2 (N5478, N5471, N177);
buf BUF1 (N5479, N5452);
buf BUF1 (N5480, N5476);
nor NOR2 (N5481, N5478, N3274);
nor NOR4 (N5482, N5464, N4260, N4833, N4383);
and AND3 (N5483, N5473, N2677, N2100);
and AND3 (N5484, N5477, N4482, N5217);
or OR2 (N5485, N5481, N4161);
and AND3 (N5486, N5484, N3891, N1980);
xor XOR2 (N5487, N5483, N5391);
not NOT1 (N5488, N5482);
buf BUF1 (N5489, N5465);
buf BUF1 (N5490, N5456);
not NOT1 (N5491, N5480);
or OR3 (N5492, N5469, N1016, N5138);
and AND3 (N5493, N5487, N5267, N2777);
or OR4 (N5494, N5474, N4124, N2353, N937);
nand NAND3 (N5495, N5488, N5058, N2289);
not NOT1 (N5496, N5485);
or OR3 (N5497, N5496, N3403, N5209);
nor NOR4 (N5498, N5490, N4589, N5149, N2483);
nand NAND4 (N5499, N5479, N4589, N5154, N1333);
nor NOR2 (N5500, N5499, N921);
or OR2 (N5501, N5486, N1780);
xor XOR2 (N5502, N5491, N51);
nor NOR3 (N5503, N5492, N669, N307);
xor XOR2 (N5504, N5497, N2790);
nand NAND3 (N5505, N5502, N3241, N2672);
nand NAND2 (N5506, N5494, N3099);
or OR2 (N5507, N5503, N633);
or OR2 (N5508, N5495, N713);
nand NAND4 (N5509, N5504, N1838, N4592, N2742);
buf BUF1 (N5510, N5505);
buf BUF1 (N5511, N5508);
nor NOR2 (N5512, N5506, N263);
and AND4 (N5513, N5493, N2667, N2934, N3577);
nor NOR3 (N5514, N5513, N4784, N1897);
and AND4 (N5515, N5511, N1181, N4430, N3000);
nand NAND4 (N5516, N5510, N5066, N383, N4016);
xor XOR2 (N5517, N5515, N5315);
not NOT1 (N5518, N5512);
nand NAND4 (N5519, N5500, N346, N884, N4163);
buf BUF1 (N5520, N5514);
not NOT1 (N5521, N5516);
nand NAND4 (N5522, N5519, N4946, N4337, N1870);
and AND3 (N5523, N5509, N1467, N4657);
buf BUF1 (N5524, N5498);
xor XOR2 (N5525, N5522, N4021);
buf BUF1 (N5526, N5524);
nor NOR3 (N5527, N5501, N2814, N4322);
buf BUF1 (N5528, N5523);
xor XOR2 (N5529, N5507, N704);
xor XOR2 (N5530, N5521, N4685);
xor XOR2 (N5531, N5520, N2969);
nand NAND3 (N5532, N5531, N2060, N3157);
not NOT1 (N5533, N5532);
nand NAND4 (N5534, N5530, N5325, N3582, N1639);
not NOT1 (N5535, N5528);
not NOT1 (N5536, N5517);
nand NAND3 (N5537, N5525, N2471, N4886);
buf BUF1 (N5538, N5535);
and AND3 (N5539, N5529, N5227, N3264);
buf BUF1 (N5540, N5539);
not NOT1 (N5541, N5526);
and AND4 (N5542, N5534, N2899, N1867, N3014);
xor XOR2 (N5543, N5537, N1159);
nor NOR2 (N5544, N5536, N2181);
nand NAND4 (N5545, N5533, N3602, N4241, N3911);
or OR4 (N5546, N5544, N911, N367, N4863);
buf BUF1 (N5547, N5489);
and AND3 (N5548, N5518, N765, N1310);
or OR4 (N5549, N5541, N2551, N1984, N986);
xor XOR2 (N5550, N5527, N161);
or OR3 (N5551, N5547, N210, N3058);
nor NOR3 (N5552, N5550, N2103, N2846);
not NOT1 (N5553, N5538);
and AND2 (N5554, N5548, N5395);
and AND2 (N5555, N5553, N3253);
or OR2 (N5556, N5554, N213);
xor XOR2 (N5557, N5552, N2416);
and AND3 (N5558, N5551, N3636, N1702);
xor XOR2 (N5559, N5558, N3993);
or OR3 (N5560, N5546, N1925, N3855);
or OR3 (N5561, N5556, N3274, N5546);
or OR4 (N5562, N5542, N12, N182, N3160);
or OR2 (N5563, N5561, N4083);
and AND2 (N5564, N5540, N3734);
buf BUF1 (N5565, N5563);
and AND2 (N5566, N5549, N3108);
buf BUF1 (N5567, N5560);
nand NAND3 (N5568, N5545, N1786, N4036);
nand NAND3 (N5569, N5564, N3243, N3229);
and AND3 (N5570, N5567, N3849, N5117);
nor NOR4 (N5571, N5559, N4290, N4571, N2367);
not NOT1 (N5572, N5566);
nand NAND2 (N5573, N5571, N5272);
not NOT1 (N5574, N5557);
buf BUF1 (N5575, N5555);
buf BUF1 (N5576, N5574);
xor XOR2 (N5577, N5565, N3479);
nand NAND3 (N5578, N5572, N2790, N2078);
not NOT1 (N5579, N5573);
xor XOR2 (N5580, N5568, N4006);
xor XOR2 (N5581, N5569, N287);
xor XOR2 (N5582, N5543, N4677);
and AND4 (N5583, N5581, N2183, N5133, N3194);
nor NOR2 (N5584, N5577, N4705);
and AND3 (N5585, N5578, N4504, N654);
buf BUF1 (N5586, N5579);
xor XOR2 (N5587, N5586, N2179);
not NOT1 (N5588, N5570);
nand NAND2 (N5589, N5582, N4350);
buf BUF1 (N5590, N5589);
or OR2 (N5591, N5580, N3544);
and AND3 (N5592, N5575, N2653, N2990);
and AND4 (N5593, N5591, N1094, N3464, N5210);
or OR4 (N5594, N5587, N4960, N4662, N2189);
xor XOR2 (N5595, N5588, N2736);
and AND4 (N5596, N5585, N3759, N465, N1013);
nor NOR4 (N5597, N5562, N5458, N2059, N2120);
not NOT1 (N5598, N5594);
nor NOR2 (N5599, N5584, N2830);
or OR2 (N5600, N5599, N4410);
and AND3 (N5601, N5592, N3865, N2932);
buf BUF1 (N5602, N5590);
not NOT1 (N5603, N5595);
or OR3 (N5604, N5601, N4590, N2769);
buf BUF1 (N5605, N5576);
not NOT1 (N5606, N5593);
not NOT1 (N5607, N5604);
not NOT1 (N5608, N5603);
nand NAND4 (N5609, N5608, N4557, N3858, N4608);
xor XOR2 (N5610, N5596, N2610);
not NOT1 (N5611, N5605);
or OR3 (N5612, N5609, N4197, N4426);
xor XOR2 (N5613, N5598, N3169);
nand NAND4 (N5614, N5602, N5045, N472, N2940);
nand NAND2 (N5615, N5600, N3903);
nor NOR4 (N5616, N5612, N493, N4181, N815);
nor NOR4 (N5617, N5616, N3446, N1359, N914);
nand NAND3 (N5618, N5613, N3104, N3140);
buf BUF1 (N5619, N5606);
or OR2 (N5620, N5597, N1341);
nand NAND4 (N5621, N5614, N2250, N135, N4237);
xor XOR2 (N5622, N5620, N3818);
buf BUF1 (N5623, N5617);
not NOT1 (N5624, N5583);
nor NOR2 (N5625, N5611, N4121);
or OR2 (N5626, N5624, N33);
buf BUF1 (N5627, N5615);
nand NAND4 (N5628, N5627, N1998, N62, N2338);
xor XOR2 (N5629, N5607, N1879);
nor NOR4 (N5630, N5626, N5245, N251, N621);
and AND3 (N5631, N5610, N282, N1586);
not NOT1 (N5632, N5625);
or OR3 (N5633, N5619, N1952, N558);
nor NOR3 (N5634, N5631, N4270, N865);
nor NOR3 (N5635, N5621, N3391, N1747);
xor XOR2 (N5636, N5634, N1530);
nand NAND3 (N5637, N5636, N3442, N2879);
xor XOR2 (N5638, N5618, N862);
not NOT1 (N5639, N5629);
and AND2 (N5640, N5639, N2543);
buf BUF1 (N5641, N5628);
nand NAND4 (N5642, N5635, N4456, N4183, N1518);
nor NOR2 (N5643, N5622, N3537);
nor NOR4 (N5644, N5623, N863, N1589, N3527);
buf BUF1 (N5645, N5643);
nand NAND3 (N5646, N5641, N4989, N5209);
nand NAND4 (N5647, N5642, N2738, N5018, N3453);
not NOT1 (N5648, N5630);
xor XOR2 (N5649, N5640, N3566);
xor XOR2 (N5650, N5649, N2595);
nor NOR4 (N5651, N5645, N549, N209, N186);
or OR4 (N5652, N5651, N4253, N4623, N371);
not NOT1 (N5653, N5647);
nor NOR3 (N5654, N5644, N96, N3254);
or OR4 (N5655, N5632, N5249, N3998, N270);
nor NOR3 (N5656, N5650, N5071, N43);
nand NAND3 (N5657, N5637, N3593, N3422);
nor NOR3 (N5658, N5656, N2552, N3879);
buf BUF1 (N5659, N5648);
nor NOR3 (N5660, N5638, N5090, N2400);
and AND4 (N5661, N5653, N5359, N3727, N4513);
not NOT1 (N5662, N5655);
xor XOR2 (N5663, N5661, N1148);
nand NAND3 (N5664, N5659, N4081, N743);
not NOT1 (N5665, N5654);
xor XOR2 (N5666, N5665, N1516);
xor XOR2 (N5667, N5658, N3894);
nor NOR4 (N5668, N5660, N2880, N1821, N383);
not NOT1 (N5669, N5668);
nor NOR2 (N5670, N5657, N3058);
nand NAND2 (N5671, N5666, N171);
nor NOR3 (N5672, N5662, N5061, N1888);
and AND2 (N5673, N5633, N5285);
or OR4 (N5674, N5671, N3869, N4207, N4920);
nand NAND4 (N5675, N5669, N1209, N5144, N3307);
not NOT1 (N5676, N5675);
not NOT1 (N5677, N5672);
or OR2 (N5678, N5667, N232);
nand NAND4 (N5679, N5646, N1944, N1483, N4797);
nand NAND4 (N5680, N5670, N641, N4909, N1338);
nand NAND4 (N5681, N5679, N2963, N4580, N1246);
xor XOR2 (N5682, N5673, N1017);
nor NOR2 (N5683, N5681, N3042);
not NOT1 (N5684, N5678);
xor XOR2 (N5685, N5674, N1303);
or OR3 (N5686, N5684, N3437, N1825);
xor XOR2 (N5687, N5680, N2354);
nor NOR4 (N5688, N5686, N761, N1483, N1837);
not NOT1 (N5689, N5683);
nor NOR2 (N5690, N5682, N26);
xor XOR2 (N5691, N5688, N4204);
xor XOR2 (N5692, N5652, N3696);
xor XOR2 (N5693, N5664, N171);
or OR2 (N5694, N5687, N5487);
xor XOR2 (N5695, N5663, N2168);
buf BUF1 (N5696, N5677);
nand NAND2 (N5697, N5692, N334);
buf BUF1 (N5698, N5685);
xor XOR2 (N5699, N5690, N5417);
and AND4 (N5700, N5693, N1909, N3718, N1728);
nand NAND4 (N5701, N5694, N3138, N5152, N5444);
buf BUF1 (N5702, N5697);
and AND3 (N5703, N5676, N981, N3171);
nand NAND2 (N5704, N5703, N3578);
or OR2 (N5705, N5695, N4879);
xor XOR2 (N5706, N5689, N3034);
nor NOR4 (N5707, N5704, N7, N5031, N4343);
not NOT1 (N5708, N5707);
nand NAND4 (N5709, N5701, N1139, N3195, N2626);
xor XOR2 (N5710, N5691, N972);
nand NAND4 (N5711, N5700, N582, N4038, N3392);
buf BUF1 (N5712, N5705);
or OR2 (N5713, N5698, N4917);
nor NOR3 (N5714, N5712, N5180, N3057);
or OR3 (N5715, N5699, N1398, N1770);
nand NAND2 (N5716, N5708, N517);
buf BUF1 (N5717, N5709);
nand NAND2 (N5718, N5706, N3155);
xor XOR2 (N5719, N5710, N3179);
or OR4 (N5720, N5713, N666, N3049, N3625);
nand NAND4 (N5721, N5696, N199, N723, N830);
xor XOR2 (N5722, N5714, N5660);
and AND2 (N5723, N5722, N2803);
xor XOR2 (N5724, N5715, N5255);
buf BUF1 (N5725, N5716);
xor XOR2 (N5726, N5724, N395);
and AND3 (N5727, N5726, N1181, N2153);
nand NAND3 (N5728, N5719, N3908, N5145);
and AND3 (N5729, N5725, N1746, N5576);
or OR4 (N5730, N5721, N5642, N2427, N5553);
buf BUF1 (N5731, N5730);
or OR2 (N5732, N5728, N2690);
nand NAND2 (N5733, N5729, N2675);
nor NOR4 (N5734, N5718, N1391, N4775, N3391);
or OR3 (N5735, N5727, N3616, N5465);
and AND4 (N5736, N5733, N674, N5662, N2855);
or OR4 (N5737, N5702, N4837, N1939, N3968);
nor NOR2 (N5738, N5717, N1384);
or OR3 (N5739, N5734, N3858, N1660);
xor XOR2 (N5740, N5736, N398);
nand NAND3 (N5741, N5732, N2960, N2484);
xor XOR2 (N5742, N5740, N5483);
xor XOR2 (N5743, N5723, N4896);
xor XOR2 (N5744, N5711, N4888);
not NOT1 (N5745, N5731);
nand NAND2 (N5746, N5744, N1440);
nand NAND2 (N5747, N5720, N590);
nor NOR4 (N5748, N5742, N5259, N3675, N3365);
buf BUF1 (N5749, N5743);
buf BUF1 (N5750, N5741);
xor XOR2 (N5751, N5738, N3525);
nor NOR2 (N5752, N5749, N476);
nand NAND2 (N5753, N5752, N5092);
buf BUF1 (N5754, N5735);
not NOT1 (N5755, N5751);
buf BUF1 (N5756, N5737);
and AND2 (N5757, N5739, N2684);
and AND3 (N5758, N5750, N993, N4522);
xor XOR2 (N5759, N5745, N3267);
not NOT1 (N5760, N5757);
nand NAND2 (N5761, N5758, N3307);
xor XOR2 (N5762, N5753, N2798);
not NOT1 (N5763, N5755);
not NOT1 (N5764, N5756);
xor XOR2 (N5765, N5747, N686);
buf BUF1 (N5766, N5765);
or OR2 (N5767, N5764, N4353);
xor XOR2 (N5768, N5760, N1055);
or OR4 (N5769, N5759, N2672, N2027, N624);
xor XOR2 (N5770, N5746, N4065);
nand NAND3 (N5771, N5761, N1985, N5357);
and AND4 (N5772, N5762, N2007, N3131, N4287);
buf BUF1 (N5773, N5754);
or OR3 (N5774, N5772, N2087, N3565);
nor NOR2 (N5775, N5771, N1000);
and AND4 (N5776, N5769, N3996, N2411, N1608);
not NOT1 (N5777, N5774);
nand NAND2 (N5778, N5763, N697);
xor XOR2 (N5779, N5768, N1081);
nor NOR2 (N5780, N5776, N1452);
xor XOR2 (N5781, N5766, N5448);
or OR2 (N5782, N5767, N2425);
or OR2 (N5783, N5780, N2820);
nor NOR4 (N5784, N5773, N2114, N4347, N420);
or OR2 (N5785, N5770, N4811);
nor NOR3 (N5786, N5784, N4247, N1430);
or OR2 (N5787, N5778, N404);
buf BUF1 (N5788, N5786);
xor XOR2 (N5789, N5787, N1815);
nand NAND4 (N5790, N5781, N1162, N4706, N4944);
and AND3 (N5791, N5777, N5343, N3904);
xor XOR2 (N5792, N5779, N4413);
buf BUF1 (N5793, N5789);
buf BUF1 (N5794, N5748);
or OR3 (N5795, N5794, N2899, N3573);
not NOT1 (N5796, N5791);
nand NAND2 (N5797, N5782, N2544);
not NOT1 (N5798, N5792);
xor XOR2 (N5799, N5795, N5143);
buf BUF1 (N5800, N5797);
nor NOR3 (N5801, N5788, N2942, N1428);
nand NAND2 (N5802, N5800, N881);
nor NOR3 (N5803, N5796, N1009, N2779);
nand NAND3 (N5804, N5799, N2165, N5051);
not NOT1 (N5805, N5804);
buf BUF1 (N5806, N5793);
and AND4 (N5807, N5775, N5695, N2593, N784);
buf BUF1 (N5808, N5806);
xor XOR2 (N5809, N5803, N4417);
or OR3 (N5810, N5807, N2691, N3464);
not NOT1 (N5811, N5790);
nor NOR4 (N5812, N5785, N5066, N4321, N2835);
nand NAND3 (N5813, N5802, N1231, N1286);
nand NAND3 (N5814, N5813, N4062, N1342);
buf BUF1 (N5815, N5783);
or OR4 (N5816, N5798, N3742, N2682, N820);
xor XOR2 (N5817, N5810, N4602);
nor NOR3 (N5818, N5812, N4075, N4017);
xor XOR2 (N5819, N5817, N1971);
or OR2 (N5820, N5805, N3038);
not NOT1 (N5821, N5816);
nor NOR4 (N5822, N5815, N691, N3244, N1653);
xor XOR2 (N5823, N5821, N2212);
xor XOR2 (N5824, N5822, N2555);
nor NOR2 (N5825, N5823, N5021);
nor NOR3 (N5826, N5820, N3683, N1498);
not NOT1 (N5827, N5801);
nor NOR2 (N5828, N5826, N4776);
not NOT1 (N5829, N5808);
and AND2 (N5830, N5818, N1104);
or OR3 (N5831, N5825, N5528, N1137);
buf BUF1 (N5832, N5824);
or OR4 (N5833, N5832, N1645, N3478, N5069);
nor NOR2 (N5834, N5830, N2989);
not NOT1 (N5835, N5814);
not NOT1 (N5836, N5835);
nand NAND3 (N5837, N5833, N2059, N723);
buf BUF1 (N5838, N5819);
nand NAND2 (N5839, N5827, N5204);
nand NAND3 (N5840, N5836, N1495, N1365);
and AND4 (N5841, N5829, N30, N160, N4753);
nor NOR4 (N5842, N5834, N547, N1145, N1403);
not NOT1 (N5843, N5842);
buf BUF1 (N5844, N5828);
and AND2 (N5845, N5838, N4389);
nor NOR3 (N5846, N5840, N2326, N504);
xor XOR2 (N5847, N5837, N3138);
buf BUF1 (N5848, N5831);
nor NOR2 (N5849, N5848, N2498);
buf BUF1 (N5850, N5849);
or OR4 (N5851, N5845, N1183, N4503, N5095);
or OR4 (N5852, N5850, N5628, N23, N5620);
nor NOR3 (N5853, N5809, N5210, N3252);
not NOT1 (N5854, N5811);
and AND3 (N5855, N5851, N5854, N4244);
or OR4 (N5856, N1898, N2011, N185, N2069);
xor XOR2 (N5857, N5852, N4144);
nand NAND2 (N5858, N5847, N560);
buf BUF1 (N5859, N5846);
nand NAND3 (N5860, N5853, N1482, N5064);
or OR3 (N5861, N5839, N4851, N3095);
or OR4 (N5862, N5859, N2081, N3104, N2230);
not NOT1 (N5863, N5860);
not NOT1 (N5864, N5862);
not NOT1 (N5865, N5844);
nor NOR2 (N5866, N5857, N4087);
nand NAND2 (N5867, N5856, N5698);
or OR4 (N5868, N5843, N1025, N927, N4214);
buf BUF1 (N5869, N5841);
xor XOR2 (N5870, N5866, N3397);
not NOT1 (N5871, N5863);
nand NAND2 (N5872, N5864, N5677);
xor XOR2 (N5873, N5861, N5832);
and AND4 (N5874, N5865, N989, N1447, N1076);
and AND4 (N5875, N5868, N3543, N5544, N2634);
xor XOR2 (N5876, N5873, N5351);
nand NAND2 (N5877, N5872, N1239);
nor NOR3 (N5878, N5870, N1560, N544);
nor NOR3 (N5879, N5877, N5280, N3023);
and AND2 (N5880, N5878, N2111);
nor NOR4 (N5881, N5874, N4028, N2971, N3922);
buf BUF1 (N5882, N5881);
nor NOR2 (N5883, N5880, N4493);
and AND2 (N5884, N5876, N5010);
xor XOR2 (N5885, N5855, N913);
buf BUF1 (N5886, N5871);
not NOT1 (N5887, N5858);
not NOT1 (N5888, N5884);
not NOT1 (N5889, N5888);
not NOT1 (N5890, N5885);
nor NOR4 (N5891, N5887, N4902, N5072, N5404);
nor NOR2 (N5892, N5890, N4487);
nor NOR2 (N5893, N5879, N1655);
nand NAND4 (N5894, N5891, N3986, N1095, N2818);
buf BUF1 (N5895, N5893);
nor NOR4 (N5896, N5894, N4, N4785, N5515);
or OR4 (N5897, N5869, N107, N2941, N2442);
not NOT1 (N5898, N5882);
nor NOR4 (N5899, N5897, N1990, N5092, N5699);
nor NOR3 (N5900, N5883, N3252, N5731);
or OR4 (N5901, N5889, N4582, N370, N2291);
and AND4 (N5902, N5899, N2976, N4288, N1173);
and AND2 (N5903, N5895, N4740);
buf BUF1 (N5904, N5901);
not NOT1 (N5905, N5902);
or OR3 (N5906, N5886, N1893, N3011);
xor XOR2 (N5907, N5904, N2494);
or OR2 (N5908, N5905, N5577);
and AND2 (N5909, N5898, N2961);
nand NAND3 (N5910, N5908, N4231, N1049);
xor XOR2 (N5911, N5892, N1425);
and AND4 (N5912, N5906, N5562, N1700, N3314);
xor XOR2 (N5913, N5903, N2683);
xor XOR2 (N5914, N5907, N2653);
buf BUF1 (N5915, N5914);
buf BUF1 (N5916, N5909);
and AND2 (N5917, N5875, N3421);
not NOT1 (N5918, N5896);
or OR2 (N5919, N5917, N1902);
nor NOR4 (N5920, N5918, N2404, N3950, N2304);
nand NAND2 (N5921, N5911, N3804);
and AND4 (N5922, N5916, N5098, N2429, N3845);
not NOT1 (N5923, N5910);
xor XOR2 (N5924, N5919, N2987);
nand NAND2 (N5925, N5920, N2510);
not NOT1 (N5926, N5922);
xor XOR2 (N5927, N5900, N4582);
xor XOR2 (N5928, N5925, N2466);
xor XOR2 (N5929, N5928, N2289);
xor XOR2 (N5930, N5912, N3006);
nor NOR3 (N5931, N5915, N4442, N3967);
buf BUF1 (N5932, N5927);
buf BUF1 (N5933, N5924);
or OR2 (N5934, N5867, N2882);
or OR2 (N5935, N5930, N2991);
or OR4 (N5936, N5934, N460, N785, N5024);
and AND4 (N5937, N5913, N1941, N1694, N2650);
buf BUF1 (N5938, N5921);
nor NOR2 (N5939, N5932, N5150);
xor XOR2 (N5940, N5936, N2358);
xor XOR2 (N5941, N5926, N3854);
nand NAND4 (N5942, N5940, N3985, N2188, N4229);
not NOT1 (N5943, N5923);
not NOT1 (N5944, N5937);
nor NOR2 (N5945, N5943, N3939);
nor NOR4 (N5946, N5944, N2834, N4702, N5367);
not NOT1 (N5947, N5946);
or OR4 (N5948, N5931, N2188, N4551, N3726);
and AND4 (N5949, N5929, N220, N551, N120);
nor NOR3 (N5950, N5947, N2066, N62);
nor NOR4 (N5951, N5941, N2950, N2930, N1192);
nand NAND3 (N5952, N5935, N5412, N5101);
nand NAND2 (N5953, N5938, N165);
or OR4 (N5954, N5945, N3822, N1236, N1070);
nor NOR2 (N5955, N5953, N5058);
nor NOR2 (N5956, N5942, N4699);
nor NOR3 (N5957, N5933, N5463, N1152);
nor NOR2 (N5958, N5952, N1594);
buf BUF1 (N5959, N5956);
nor NOR4 (N5960, N5957, N1700, N5931, N5490);
buf BUF1 (N5961, N5959);
not NOT1 (N5962, N5960);
nand NAND3 (N5963, N5955, N4307, N4762);
nand NAND3 (N5964, N5962, N5312, N1882);
not NOT1 (N5965, N5963);
and AND3 (N5966, N5964, N1428, N2770);
buf BUF1 (N5967, N5948);
xor XOR2 (N5968, N5961, N5047);
xor XOR2 (N5969, N5967, N2450);
and AND3 (N5970, N5968, N62, N2666);
and AND2 (N5971, N5958, N3112);
not NOT1 (N5972, N5950);
or OR4 (N5973, N5951, N2923, N5501, N4038);
and AND3 (N5974, N5973, N1883, N1306);
not NOT1 (N5975, N5949);
or OR2 (N5976, N5939, N4061);
and AND4 (N5977, N5972, N5300, N2230, N3733);
not NOT1 (N5978, N5966);
buf BUF1 (N5979, N5971);
or OR2 (N5980, N5954, N382);
nand NAND2 (N5981, N5976, N1036);
nand NAND3 (N5982, N5978, N5804, N4372);
not NOT1 (N5983, N5979);
xor XOR2 (N5984, N5965, N5009);
nand NAND2 (N5985, N5982, N4945);
xor XOR2 (N5986, N5980, N4376);
not NOT1 (N5987, N5981);
not NOT1 (N5988, N5969);
not NOT1 (N5989, N5974);
nand NAND4 (N5990, N5985, N3936, N3865, N4041);
or OR2 (N5991, N5987, N2203);
xor XOR2 (N5992, N5977, N3646);
nand NAND3 (N5993, N5990, N1783, N1335);
buf BUF1 (N5994, N5984);
not NOT1 (N5995, N5993);
nand NAND4 (N5996, N5994, N2510, N1817, N529);
xor XOR2 (N5997, N5983, N1024);
buf BUF1 (N5998, N5992);
nor NOR4 (N5999, N5970, N685, N5495, N5515);
and AND4 (N6000, N5998, N4894, N1725, N4719);
xor XOR2 (N6001, N5996, N4141);
xor XOR2 (N6002, N6000, N5581);
and AND3 (N6003, N5999, N263, N3530);
or OR4 (N6004, N5997, N3895, N4020, N6000);
nor NOR3 (N6005, N6001, N4699, N5403);
nand NAND3 (N6006, N6004, N62, N1401);
not NOT1 (N6007, N5988);
buf BUF1 (N6008, N6006);
or OR2 (N6009, N5991, N4468);
or OR4 (N6010, N5975, N3201, N4773, N2795);
buf BUF1 (N6011, N5989);
nand NAND3 (N6012, N6007, N263, N1051);
nor NOR3 (N6013, N5995, N64, N1889);
nor NOR3 (N6014, N6012, N3737, N145);
xor XOR2 (N6015, N6002, N1558);
nand NAND4 (N6016, N6015, N2836, N3853, N1425);
and AND4 (N6017, N6013, N2927, N665, N4752);
xor XOR2 (N6018, N6016, N5821);
and AND2 (N6019, N6003, N2411);
nand NAND2 (N6020, N6011, N5549);
and AND3 (N6021, N6017, N4091, N1112);
or OR3 (N6022, N6005, N5418, N851);
nand NAND2 (N6023, N6010, N3172);
or OR2 (N6024, N6008, N5184);
or OR4 (N6025, N6009, N3685, N5108, N4445);
buf BUF1 (N6026, N6024);
nor NOR4 (N6027, N6018, N712, N386, N4329);
nand NAND4 (N6028, N6022, N4456, N1795, N38);
or OR2 (N6029, N6025, N1251);
buf BUF1 (N6030, N6029);
buf BUF1 (N6031, N6020);
nand NAND3 (N6032, N6014, N4264, N2102);
or OR4 (N6033, N6023, N2469, N30, N5848);
or OR2 (N6034, N6033, N5091);
and AND3 (N6035, N6031, N3303, N1977);
xor XOR2 (N6036, N6021, N493);
nand NAND2 (N6037, N5986, N2634);
buf BUF1 (N6038, N6032);
nor NOR4 (N6039, N6019, N2180, N3276, N657);
and AND3 (N6040, N6039, N1377, N1453);
not NOT1 (N6041, N6027);
nor NOR2 (N6042, N6028, N1732);
or OR3 (N6043, N6035, N2471, N72);
or OR4 (N6044, N6030, N3293, N1507, N911);
nand NAND3 (N6045, N6044, N1778, N1307);
not NOT1 (N6046, N6038);
and AND4 (N6047, N6046, N2370, N1535, N2721);
buf BUF1 (N6048, N6047);
xor XOR2 (N6049, N6036, N5609);
not NOT1 (N6050, N6042);
and AND3 (N6051, N6034, N2345, N1000);
buf BUF1 (N6052, N6049);
or OR4 (N6053, N6040, N77, N1577, N4196);
not NOT1 (N6054, N6037);
buf BUF1 (N6055, N6054);
buf BUF1 (N6056, N6055);
nand NAND2 (N6057, N6051, N5242);
or OR2 (N6058, N6026, N3262);
nor NOR2 (N6059, N6050, N4906);
xor XOR2 (N6060, N6059, N2677);
xor XOR2 (N6061, N6045, N1368);
not NOT1 (N6062, N6061);
or OR4 (N6063, N6060, N4911, N4841, N3010);
nor NOR2 (N6064, N6062, N2672);
buf BUF1 (N6065, N6057);
nand NAND4 (N6066, N6064, N2731, N2141, N5555);
buf BUF1 (N6067, N6058);
nor NOR2 (N6068, N6041, N1587);
and AND3 (N6069, N6043, N3580, N1190);
or OR4 (N6070, N6056, N4309, N45, N1904);
nor NOR3 (N6071, N6067, N2409, N1159);
or OR3 (N6072, N6065, N5098, N2228);
nor NOR4 (N6073, N6052, N620, N1934, N2390);
buf BUF1 (N6074, N6072);
nor NOR3 (N6075, N6073, N5202, N5792);
buf BUF1 (N6076, N6071);
or OR4 (N6077, N6053, N819, N2003, N3175);
and AND2 (N6078, N6076, N1927);
and AND4 (N6079, N6069, N2182, N540, N5608);
nor NOR2 (N6080, N6077, N1500);
not NOT1 (N6081, N6063);
or OR3 (N6082, N6074, N2731, N496);
not NOT1 (N6083, N6082);
xor XOR2 (N6084, N6068, N3767);
not NOT1 (N6085, N6080);
or OR2 (N6086, N6048, N4430);
nor NOR4 (N6087, N6084, N1825, N1196, N5765);
or OR4 (N6088, N6085, N3037, N5691, N3602);
or OR4 (N6089, N6081, N4241, N4051, N5709);
xor XOR2 (N6090, N6086, N2447);
xor XOR2 (N6091, N6070, N5564);
nand NAND3 (N6092, N6090, N3603, N243);
xor XOR2 (N6093, N6088, N1670);
or OR3 (N6094, N6066, N3573, N5351);
or OR3 (N6095, N6083, N501, N1263);
nand NAND2 (N6096, N6093, N4997);
nor NOR3 (N6097, N6095, N1119, N2597);
nor NOR4 (N6098, N6087, N5046, N5492, N645);
nor NOR3 (N6099, N6096, N2325, N4447);
or OR3 (N6100, N6075, N4407, N3214);
buf BUF1 (N6101, N6094);
buf BUF1 (N6102, N6092);
and AND2 (N6103, N6078, N560);
nand NAND2 (N6104, N6097, N3263);
or OR4 (N6105, N6101, N1179, N2700, N4240);
nor NOR2 (N6106, N6098, N1056);
nor NOR4 (N6107, N6099, N2659, N4166, N4280);
buf BUF1 (N6108, N6105);
not NOT1 (N6109, N6104);
nor NOR2 (N6110, N6089, N2444);
nor NOR3 (N6111, N6110, N284, N3134);
buf BUF1 (N6112, N6108);
buf BUF1 (N6113, N6079);
xor XOR2 (N6114, N6103, N696);
nand NAND3 (N6115, N6112, N1171, N2547);
buf BUF1 (N6116, N6114);
xor XOR2 (N6117, N6109, N667);
or OR4 (N6118, N6113, N2561, N6102, N5727);
nor NOR4 (N6119, N3463, N496, N1169, N83);
buf BUF1 (N6120, N6111);
xor XOR2 (N6121, N6118, N2529);
xor XOR2 (N6122, N6115, N5734);
and AND2 (N6123, N6119, N358);
not NOT1 (N6124, N6106);
xor XOR2 (N6125, N6120, N4606);
buf BUF1 (N6126, N6123);
xor XOR2 (N6127, N6121, N4444);
nor NOR2 (N6128, N6127, N2965);
not NOT1 (N6129, N6117);
and AND4 (N6130, N6124, N675, N107, N534);
nand NAND3 (N6131, N6100, N4203, N4466);
xor XOR2 (N6132, N6122, N5420);
not NOT1 (N6133, N6130);
and AND3 (N6134, N6107, N5668, N5811);
and AND3 (N6135, N6116, N4917, N651);
buf BUF1 (N6136, N6132);
xor XOR2 (N6137, N6128, N2865);
nor NOR3 (N6138, N6137, N31, N1749);
nand NAND2 (N6139, N6136, N2077);
not NOT1 (N6140, N6131);
nand NAND2 (N6141, N6134, N312);
nor NOR3 (N6142, N6135, N2753, N386);
xor XOR2 (N6143, N6125, N1497);
nor NOR2 (N6144, N6138, N5303);
xor XOR2 (N6145, N6091, N3720);
or OR2 (N6146, N6143, N3687);
and AND3 (N6147, N6141, N37, N2491);
or OR3 (N6148, N6133, N5714, N5148);
buf BUF1 (N6149, N6148);
xor XOR2 (N6150, N6145, N3140);
nor NOR2 (N6151, N6144, N2861);
not NOT1 (N6152, N6139);
xor XOR2 (N6153, N6149, N331);
and AND2 (N6154, N6147, N5580);
or OR4 (N6155, N6153, N260, N4592, N4229);
nand NAND2 (N6156, N6151, N2049);
xor XOR2 (N6157, N6140, N3121);
nand NAND2 (N6158, N6155, N5076);
buf BUF1 (N6159, N6157);
or OR4 (N6160, N6152, N1538, N984, N5423);
buf BUF1 (N6161, N6126);
xor XOR2 (N6162, N6142, N2370);
nor NOR3 (N6163, N6162, N526, N550);
and AND2 (N6164, N6150, N2570);
nor NOR3 (N6165, N6159, N3875, N4881);
nand NAND2 (N6166, N6165, N4397);
not NOT1 (N6167, N6166);
not NOT1 (N6168, N6167);
xor XOR2 (N6169, N6168, N3691);
xor XOR2 (N6170, N6154, N4044);
xor XOR2 (N6171, N6170, N1966);
nor NOR3 (N6172, N6129, N5520, N4798);
nor NOR4 (N6173, N6146, N947, N5097, N4292);
nor NOR3 (N6174, N6169, N116, N6060);
and AND3 (N6175, N6161, N5571, N6095);
nand NAND2 (N6176, N6174, N306);
nand NAND3 (N6177, N6164, N3218, N1997);
not NOT1 (N6178, N6175);
nand NAND3 (N6179, N6176, N1875, N251);
nand NAND4 (N6180, N6171, N1007, N3751, N5415);
or OR2 (N6181, N6156, N5090);
nor NOR2 (N6182, N6163, N4724);
buf BUF1 (N6183, N6180);
nor NOR4 (N6184, N6183, N1080, N3437, N1316);
buf BUF1 (N6185, N6158);
not NOT1 (N6186, N6173);
not NOT1 (N6187, N6160);
or OR3 (N6188, N6185, N1519, N4500);
buf BUF1 (N6189, N6177);
not NOT1 (N6190, N6186);
or OR3 (N6191, N6184, N1431, N3467);
xor XOR2 (N6192, N6190, N62);
buf BUF1 (N6193, N6189);
xor XOR2 (N6194, N6187, N5541);
nor NOR4 (N6195, N6188, N5712, N2572, N654);
buf BUF1 (N6196, N6192);
not NOT1 (N6197, N6191);
or OR3 (N6198, N6195, N1668, N955);
and AND3 (N6199, N6197, N1269, N5599);
nor NOR3 (N6200, N6179, N1822, N3509);
buf BUF1 (N6201, N6181);
or OR4 (N6202, N6199, N3737, N5077, N839);
nand NAND3 (N6203, N6200, N440, N5865);
buf BUF1 (N6204, N6172);
nand NAND4 (N6205, N6182, N1395, N2115, N2965);
nor NOR3 (N6206, N6204, N5129, N893);
and AND2 (N6207, N6203, N680);
or OR4 (N6208, N6201, N743, N3976, N2565);
and AND2 (N6209, N6206, N5758);
nand NAND4 (N6210, N6209, N6037, N989, N1352);
nor NOR2 (N6211, N6193, N407);
buf BUF1 (N6212, N6198);
nand NAND4 (N6213, N6196, N4895, N1398, N1450);
not NOT1 (N6214, N6208);
nor NOR2 (N6215, N6205, N2004);
or OR4 (N6216, N6214, N2277, N3420, N5673);
not NOT1 (N6217, N6207);
or OR3 (N6218, N6202, N495, N5245);
or OR2 (N6219, N6211, N3386);
buf BUF1 (N6220, N6217);
buf BUF1 (N6221, N6220);
buf BUF1 (N6222, N6215);
nand NAND4 (N6223, N6212, N5019, N1609, N483);
nand NAND4 (N6224, N6218, N3070, N1180, N2025);
nor NOR3 (N6225, N6178, N4864, N6071);
nand NAND4 (N6226, N6223, N5659, N4683, N4322);
or OR4 (N6227, N6221, N4042, N5870, N4713);
and AND4 (N6228, N6225, N5988, N641, N2280);
or OR2 (N6229, N6226, N5414);
nor NOR2 (N6230, N6227, N4356);
xor XOR2 (N6231, N6228, N395);
and AND3 (N6232, N6229, N584, N2768);
xor XOR2 (N6233, N6224, N2958);
buf BUF1 (N6234, N6230);
or OR3 (N6235, N6233, N470, N6172);
not NOT1 (N6236, N6219);
or OR2 (N6237, N6236, N2409);
buf BUF1 (N6238, N6216);
nand NAND3 (N6239, N6238, N1793, N4461);
not NOT1 (N6240, N6210);
buf BUF1 (N6241, N6239);
nand NAND4 (N6242, N6231, N4921, N2078, N4920);
not NOT1 (N6243, N6237);
nor NOR4 (N6244, N6234, N5565, N3131, N2593);
xor XOR2 (N6245, N6194, N3914);
not NOT1 (N6246, N6222);
buf BUF1 (N6247, N6235);
and AND3 (N6248, N6241, N1753, N4048);
not NOT1 (N6249, N6240);
nand NAND2 (N6250, N6242, N3394);
or OR4 (N6251, N6250, N4433, N5670, N2050);
xor XOR2 (N6252, N6232, N2647);
or OR4 (N6253, N6249, N3319, N1752, N5207);
and AND2 (N6254, N6213, N3038);
nand NAND2 (N6255, N6251, N4970);
nor NOR3 (N6256, N6243, N3859, N1109);
and AND2 (N6257, N6255, N388);
xor XOR2 (N6258, N6253, N3968);
not NOT1 (N6259, N6246);
and AND4 (N6260, N6256, N3047, N3685, N4619);
nor NOR3 (N6261, N6252, N1818, N4157);
xor XOR2 (N6262, N6261, N305);
and AND4 (N6263, N6245, N5804, N2368, N4605);
nand NAND3 (N6264, N6247, N1865, N2757);
not NOT1 (N6265, N6264);
nand NAND4 (N6266, N6257, N3110, N3746, N1276);
and AND3 (N6267, N6248, N3579, N6109);
and AND3 (N6268, N6254, N2053, N4712);
nor NOR3 (N6269, N6262, N4257, N5801);
buf BUF1 (N6270, N6259);
xor XOR2 (N6271, N6267, N4680);
not NOT1 (N6272, N6266);
xor XOR2 (N6273, N6272, N3460);
buf BUF1 (N6274, N6244);
nand NAND4 (N6275, N6270, N4902, N6107, N4101);
not NOT1 (N6276, N6271);
and AND4 (N6277, N6274, N4293, N1812, N1379);
nor NOR3 (N6278, N6276, N825, N2722);
nand NAND4 (N6279, N6269, N2446, N5202, N5027);
and AND3 (N6280, N6277, N3822, N2822);
not NOT1 (N6281, N6258);
nand NAND4 (N6282, N6281, N308, N3066, N660);
buf BUF1 (N6283, N6263);
nor NOR2 (N6284, N6280, N5872);
xor XOR2 (N6285, N6265, N2089);
nor NOR2 (N6286, N6260, N5191);
not NOT1 (N6287, N6279);
and AND2 (N6288, N6284, N3906);
nand NAND3 (N6289, N6287, N4104, N4418);
and AND3 (N6290, N6288, N3835, N814);
nor NOR4 (N6291, N6275, N74, N4867, N4734);
not NOT1 (N6292, N6273);
and AND2 (N6293, N6283, N1870);
and AND4 (N6294, N6278, N1622, N4109, N939);
nand NAND3 (N6295, N6285, N3597, N829);
not NOT1 (N6296, N6289);
nor NOR4 (N6297, N6292, N366, N2057, N4516);
nor NOR3 (N6298, N6286, N3490, N1453);
buf BUF1 (N6299, N6296);
nand NAND4 (N6300, N6299, N6251, N3715, N1378);
not NOT1 (N6301, N6291);
buf BUF1 (N6302, N6290);
xor XOR2 (N6303, N6297, N5186);
nor NOR4 (N6304, N6298, N6083, N3183, N1200);
xor XOR2 (N6305, N6294, N3947);
xor XOR2 (N6306, N6305, N4112);
and AND3 (N6307, N6303, N3545, N4424);
nor NOR4 (N6308, N6307, N167, N5123, N1933);
and AND2 (N6309, N6295, N4665);
nand NAND3 (N6310, N6302, N2685, N1219);
nand NAND2 (N6311, N6268, N2517);
nand NAND3 (N6312, N6306, N4855, N2059);
xor XOR2 (N6313, N6308, N1482);
not NOT1 (N6314, N6301);
xor XOR2 (N6315, N6282, N566);
nor NOR4 (N6316, N6309, N542, N1585, N2468);
nand NAND2 (N6317, N6304, N3889);
xor XOR2 (N6318, N6315, N5029);
nor NOR4 (N6319, N6313, N5383, N2202, N2050);
nand NAND4 (N6320, N6311, N2337, N258, N3346);
buf BUF1 (N6321, N6293);
not NOT1 (N6322, N6319);
nor NOR2 (N6323, N6322, N3882);
not NOT1 (N6324, N6310);
xor XOR2 (N6325, N6318, N1151);
and AND4 (N6326, N6325, N3478, N143, N3001);
nand NAND2 (N6327, N6316, N157);
and AND3 (N6328, N6314, N2220, N5278);
or OR2 (N6329, N6328, N5364);
or OR3 (N6330, N6320, N5279, N5501);
nand NAND2 (N6331, N6326, N1551);
nor NOR4 (N6332, N6317, N5161, N1733, N522);
nand NAND3 (N6333, N6330, N4577, N4561);
nand NAND2 (N6334, N6332, N3338);
and AND3 (N6335, N6324, N5328, N1788);
nand NAND4 (N6336, N6300, N5661, N5420, N2658);
not NOT1 (N6337, N6331);
and AND3 (N6338, N6336, N2420, N1737);
and AND4 (N6339, N6335, N5338, N2948, N12);
buf BUF1 (N6340, N6337);
nor NOR4 (N6341, N6327, N4388, N3507, N5172);
nor NOR3 (N6342, N6339, N2364, N1646);
and AND4 (N6343, N6340, N1264, N6167, N5220);
nor NOR4 (N6344, N6312, N1417, N3485, N5907);
nor NOR4 (N6345, N6344, N2949, N52, N3343);
nand NAND3 (N6346, N6334, N5469, N4214);
not NOT1 (N6347, N6323);
xor XOR2 (N6348, N6342, N2529);
and AND4 (N6349, N6341, N575, N4206, N3229);
or OR4 (N6350, N6349, N1805, N3772, N3917);
nor NOR2 (N6351, N6345, N4293);
nand NAND2 (N6352, N6350, N1310);
or OR2 (N6353, N6352, N3860);
buf BUF1 (N6354, N6343);
nand NAND3 (N6355, N6346, N239, N1604);
and AND3 (N6356, N6353, N6080, N4143);
xor XOR2 (N6357, N6338, N1063);
xor XOR2 (N6358, N6356, N2587);
or OR3 (N6359, N6321, N1314, N599);
nor NOR2 (N6360, N6347, N1212);
xor XOR2 (N6361, N6351, N5808);
or OR3 (N6362, N6348, N1581, N445);
nor NOR3 (N6363, N6358, N5278, N3891);
buf BUF1 (N6364, N6359);
xor XOR2 (N6365, N6355, N2723);
and AND2 (N6366, N6357, N2829);
not NOT1 (N6367, N6363);
and AND2 (N6368, N6365, N2951);
not NOT1 (N6369, N6362);
xor XOR2 (N6370, N6367, N5083);
nor NOR4 (N6371, N6329, N1979, N776, N4779);
xor XOR2 (N6372, N6360, N1839);
nor NOR2 (N6373, N6370, N1141);
not NOT1 (N6374, N6372);
and AND2 (N6375, N6374, N2587);
xor XOR2 (N6376, N6354, N3742);
nor NOR4 (N6377, N6371, N5594, N4540, N3694);
xor XOR2 (N6378, N6376, N2356);
nand NAND2 (N6379, N6373, N5476);
buf BUF1 (N6380, N6369);
or OR3 (N6381, N6379, N637, N2427);
not NOT1 (N6382, N6364);
buf BUF1 (N6383, N6381);
and AND3 (N6384, N6366, N1387, N824);
or OR3 (N6385, N6383, N416, N383);
nand NAND2 (N6386, N6368, N1607);
nand NAND2 (N6387, N6377, N4614);
nand NAND2 (N6388, N6386, N394);
and AND3 (N6389, N6333, N3162, N5440);
and AND4 (N6390, N6385, N5597, N5867, N1346);
nor NOR3 (N6391, N6388, N4732, N5107);
nor NOR2 (N6392, N6387, N6292);
nor NOR4 (N6393, N6392, N5845, N2956, N4153);
xor XOR2 (N6394, N6384, N2729);
buf BUF1 (N6395, N6390);
buf BUF1 (N6396, N6393);
buf BUF1 (N6397, N6389);
xor XOR2 (N6398, N6391, N4845);
and AND3 (N6399, N6396, N3952, N5379);
nor NOR2 (N6400, N6378, N5856);
buf BUF1 (N6401, N6394);
and AND3 (N6402, N6361, N3069, N3061);
or OR3 (N6403, N6397, N2844, N4792);
xor XOR2 (N6404, N6403, N1047);
buf BUF1 (N6405, N6382);
nor NOR2 (N6406, N6395, N4757);
buf BUF1 (N6407, N6375);
not NOT1 (N6408, N6400);
xor XOR2 (N6409, N6407, N4387);
nand NAND3 (N6410, N6404, N2559, N5167);
nor NOR3 (N6411, N6401, N859, N3475);
nand NAND3 (N6412, N6380, N467, N4668);
or OR2 (N6413, N6410, N6190);
not NOT1 (N6414, N6398);
nand NAND4 (N6415, N6405, N5963, N4583, N4294);
nor NOR4 (N6416, N6408, N649, N573, N285);
nand NAND3 (N6417, N6406, N2655, N2917);
nand NAND4 (N6418, N6411, N5534, N1017, N6093);
not NOT1 (N6419, N6415);
or OR2 (N6420, N6399, N5423);
not NOT1 (N6421, N6418);
or OR4 (N6422, N6420, N6007, N1611, N1293);
and AND3 (N6423, N6419, N3107, N1785);
xor XOR2 (N6424, N6413, N1548);
nand NAND3 (N6425, N6423, N638, N2295);
nor NOR2 (N6426, N6402, N853);
xor XOR2 (N6427, N6424, N307);
nand NAND4 (N6428, N6421, N3198, N2962, N4834);
or OR2 (N6429, N6422, N2221);
not NOT1 (N6430, N6417);
or OR4 (N6431, N6414, N856, N816, N1758);
not NOT1 (N6432, N6416);
not NOT1 (N6433, N6429);
and AND3 (N6434, N6428, N1512, N650);
nor NOR3 (N6435, N6432, N5226, N2286);
xor XOR2 (N6436, N6426, N2918);
nor NOR2 (N6437, N6433, N2348);
nand NAND2 (N6438, N6436, N4525);
nand NAND2 (N6439, N6412, N2197);
not NOT1 (N6440, N6439);
and AND3 (N6441, N6425, N96, N3512);
nand NAND4 (N6442, N6434, N413, N2371, N6392);
or OR2 (N6443, N6440, N220);
not NOT1 (N6444, N6431);
buf BUF1 (N6445, N6435);
xor XOR2 (N6446, N6442, N1836);
nand NAND4 (N6447, N6438, N5198, N1047, N3958);
or OR4 (N6448, N6430, N1850, N5087, N1883);
or OR3 (N6449, N6446, N950, N3440);
or OR3 (N6450, N6443, N5979, N5241);
xor XOR2 (N6451, N6409, N2917);
or OR2 (N6452, N6449, N3960);
xor XOR2 (N6453, N6452, N2453);
xor XOR2 (N6454, N6437, N2618);
and AND2 (N6455, N6448, N2544);
buf BUF1 (N6456, N6450);
xor XOR2 (N6457, N6445, N1977);
nor NOR2 (N6458, N6441, N6142);
nor NOR2 (N6459, N6455, N5378);
buf BUF1 (N6460, N6427);
buf BUF1 (N6461, N6453);
nor NOR4 (N6462, N6454, N2929, N2605, N2620);
buf BUF1 (N6463, N6451);
buf BUF1 (N6464, N6461);
nand NAND4 (N6465, N6456, N5226, N2377, N2431);
not NOT1 (N6466, N6457);
buf BUF1 (N6467, N6464);
nor NOR2 (N6468, N6465, N4838);
not NOT1 (N6469, N6463);
or OR3 (N6470, N6468, N1397, N2279);
xor XOR2 (N6471, N6462, N2032);
xor XOR2 (N6472, N6467, N2160);
buf BUF1 (N6473, N6466);
and AND2 (N6474, N6472, N5272);
or OR3 (N6475, N6444, N2068, N4644);
and AND4 (N6476, N6459, N4549, N1193, N1817);
xor XOR2 (N6477, N6469, N1969);
xor XOR2 (N6478, N6471, N6268);
and AND3 (N6479, N6447, N3340, N1702);
or OR3 (N6480, N6474, N3234, N3308);
buf BUF1 (N6481, N6460);
and AND2 (N6482, N6473, N5821);
nand NAND2 (N6483, N6458, N1699);
not NOT1 (N6484, N6470);
nand NAND2 (N6485, N6483, N2796);
xor XOR2 (N6486, N6480, N4118);
or OR2 (N6487, N6475, N2332);
buf BUF1 (N6488, N6484);
xor XOR2 (N6489, N6485, N1211);
or OR4 (N6490, N6481, N1470, N869, N714);
and AND4 (N6491, N6476, N545, N6163, N5215);
not NOT1 (N6492, N6490);
not NOT1 (N6493, N6486);
and AND3 (N6494, N6493, N1017, N3671);
or OR4 (N6495, N6489, N5344, N517, N485);
or OR2 (N6496, N6477, N2153);
not NOT1 (N6497, N6491);
not NOT1 (N6498, N6488);
or OR2 (N6499, N6482, N5804);
and AND2 (N6500, N6494, N2967);
xor XOR2 (N6501, N6492, N4292);
nand NAND2 (N6502, N6495, N4741);
or OR2 (N6503, N6500, N3022);
nand NAND3 (N6504, N6497, N5349, N1988);
not NOT1 (N6505, N6503);
and AND2 (N6506, N6498, N3043);
not NOT1 (N6507, N6502);
and AND2 (N6508, N6507, N32);
or OR2 (N6509, N6505, N1353);
not NOT1 (N6510, N6478);
buf BUF1 (N6511, N6496);
buf BUF1 (N6512, N6508);
or OR2 (N6513, N6487, N5945);
nand NAND3 (N6514, N6513, N446, N2385);
or OR2 (N6515, N6506, N3694);
nor NOR2 (N6516, N6512, N1736);
nor NOR4 (N6517, N6499, N3652, N686, N4244);
nand NAND4 (N6518, N6509, N1096, N2551, N2712);
xor XOR2 (N6519, N6515, N224);
or OR3 (N6520, N6511, N30, N5114);
or OR2 (N6521, N6479, N3619);
nor NOR3 (N6522, N6517, N5307, N1828);
nor NOR2 (N6523, N6516, N1770);
xor XOR2 (N6524, N6523, N4824);
and AND3 (N6525, N6514, N1313, N1906);
nor NOR3 (N6526, N6521, N1461, N4030);
not NOT1 (N6527, N6522);
nor NOR4 (N6528, N6510, N4620, N499, N2199);
nand NAND4 (N6529, N6524, N5991, N3013, N5171);
and AND4 (N6530, N6527, N1820, N650, N4093);
not NOT1 (N6531, N6501);
or OR3 (N6532, N6520, N1788, N6060);
not NOT1 (N6533, N6529);
or OR2 (N6534, N6518, N2490);
and AND2 (N6535, N6519, N250);
xor XOR2 (N6536, N6533, N5439);
buf BUF1 (N6537, N6528);
buf BUF1 (N6538, N6526);
xor XOR2 (N6539, N6525, N5649);
nand NAND3 (N6540, N6530, N865, N3462);
and AND4 (N6541, N6531, N4570, N4914, N5350);
nor NOR4 (N6542, N6538, N3024, N3861, N2123);
not NOT1 (N6543, N6536);
not NOT1 (N6544, N6504);
nor NOR3 (N6545, N6544, N4136, N5023);
nand NAND4 (N6546, N6535, N146, N536, N641);
nand NAND2 (N6547, N6542, N6166);
nand NAND3 (N6548, N6540, N2715, N1668);
nor NOR3 (N6549, N6545, N6203, N2712);
and AND2 (N6550, N6546, N6390);
and AND3 (N6551, N6548, N354, N1998);
xor XOR2 (N6552, N6534, N5746);
and AND3 (N6553, N6541, N2567, N3761);
or OR2 (N6554, N6532, N259);
buf BUF1 (N6555, N6543);
nor NOR2 (N6556, N6554, N6215);
and AND3 (N6557, N6537, N2540, N5219);
nor NOR4 (N6558, N6553, N4618, N5237, N3226);
or OR2 (N6559, N6552, N848);
xor XOR2 (N6560, N6551, N6246);
or OR4 (N6561, N6547, N821, N2604, N5565);
nor NOR4 (N6562, N6558, N4948, N4425, N4412);
nor NOR3 (N6563, N6559, N2865, N4861);
xor XOR2 (N6564, N6560, N1346);
or OR4 (N6565, N6557, N5168, N5297, N3941);
nor NOR4 (N6566, N6555, N4703, N1707, N6031);
buf BUF1 (N6567, N6556);
nand NAND3 (N6568, N6567, N5234, N6094);
buf BUF1 (N6569, N6539);
xor XOR2 (N6570, N6549, N3303);
xor XOR2 (N6571, N6561, N4840);
or OR4 (N6572, N6550, N3680, N4937, N3445);
not NOT1 (N6573, N6562);
not NOT1 (N6574, N6569);
not NOT1 (N6575, N6570);
not NOT1 (N6576, N6564);
buf BUF1 (N6577, N6572);
and AND4 (N6578, N6568, N783, N5619, N2878);
and AND3 (N6579, N6573, N2258, N1261);
and AND2 (N6580, N6579, N2648);
and AND3 (N6581, N6577, N6302, N5992);
xor XOR2 (N6582, N6563, N1573);
buf BUF1 (N6583, N6576);
not NOT1 (N6584, N6565);
nor NOR3 (N6585, N6584, N6213, N298);
or OR3 (N6586, N6566, N2121, N2617);
not NOT1 (N6587, N6580);
not NOT1 (N6588, N6574);
nand NAND2 (N6589, N6586, N3545);
and AND3 (N6590, N6578, N6551, N615);
or OR4 (N6591, N6585, N2058, N201, N531);
xor XOR2 (N6592, N6587, N4576);
or OR2 (N6593, N6571, N5063);
buf BUF1 (N6594, N6588);
nor NOR4 (N6595, N6591, N5327, N4028, N3845);
buf BUF1 (N6596, N6595);
nand NAND2 (N6597, N6590, N3166);
buf BUF1 (N6598, N6582);
nand NAND4 (N6599, N6596, N959, N1843, N5491);
nor NOR2 (N6600, N6592, N4122);
xor XOR2 (N6601, N6598, N3288);
or OR4 (N6602, N6593, N2205, N1115, N4198);
buf BUF1 (N6603, N6599);
nand NAND2 (N6604, N6583, N1222);
buf BUF1 (N6605, N6594);
and AND2 (N6606, N6589, N1219);
or OR2 (N6607, N6575, N1626);
buf BUF1 (N6608, N6581);
not NOT1 (N6609, N6602);
nand NAND3 (N6610, N6597, N5539, N2738);
and AND3 (N6611, N6608, N4131, N290);
or OR3 (N6612, N6610, N1559, N1574);
not NOT1 (N6613, N6609);
not NOT1 (N6614, N6600);
or OR3 (N6615, N6605, N1238, N1962);
nand NAND2 (N6616, N6612, N2148);
or OR3 (N6617, N6615, N5071, N5133);
nor NOR2 (N6618, N6606, N6437);
and AND4 (N6619, N6601, N5925, N591, N5266);
xor XOR2 (N6620, N6603, N481);
buf BUF1 (N6621, N6613);
xor XOR2 (N6622, N6619, N5329);
xor XOR2 (N6623, N6621, N2251);
and AND2 (N6624, N6620, N5666);
not NOT1 (N6625, N6622);
nor NOR2 (N6626, N6623, N5083);
or OR3 (N6627, N6624, N4424, N4190);
not NOT1 (N6628, N6618);
not NOT1 (N6629, N6616);
nand NAND2 (N6630, N6604, N3104);
nand NAND4 (N6631, N6617, N4804, N2595, N5818);
nand NAND3 (N6632, N6625, N5472, N6477);
nand NAND4 (N6633, N6611, N5062, N93, N3867);
buf BUF1 (N6634, N6633);
nand NAND2 (N6635, N6607, N5354);
and AND3 (N6636, N6626, N2755, N4403);
or OR3 (N6637, N6629, N6576, N3031);
buf BUF1 (N6638, N6631);
nand NAND2 (N6639, N6638, N2864);
not NOT1 (N6640, N6628);
not NOT1 (N6641, N6627);
not NOT1 (N6642, N6636);
not NOT1 (N6643, N6632);
nor NOR3 (N6644, N6614, N6400, N2293);
not NOT1 (N6645, N6630);
or OR3 (N6646, N6645, N2806, N1310);
nand NAND2 (N6647, N6641, N6368);
xor XOR2 (N6648, N6647, N5190);
not NOT1 (N6649, N6643);
buf BUF1 (N6650, N6646);
nor NOR3 (N6651, N6637, N1136, N3156);
nor NOR3 (N6652, N6648, N4538, N1929);
xor XOR2 (N6653, N6639, N1987);
nor NOR2 (N6654, N6652, N2689);
nor NOR2 (N6655, N6653, N2959);
not NOT1 (N6656, N6651);
nand NAND2 (N6657, N6634, N2099);
and AND4 (N6658, N6635, N5410, N5838, N4823);
buf BUF1 (N6659, N6640);
nand NAND3 (N6660, N6649, N3528, N4721);
nand NAND2 (N6661, N6644, N940);
and AND4 (N6662, N6658, N2619, N4753, N4238);
nand NAND2 (N6663, N6656, N3427);
xor XOR2 (N6664, N6663, N2088);
or OR3 (N6665, N6660, N5481, N209);
not NOT1 (N6666, N6657);
xor XOR2 (N6667, N6666, N1502);
nor NOR3 (N6668, N6659, N2529, N4504);
and AND3 (N6669, N6662, N5992, N6342);
not NOT1 (N6670, N6664);
or OR4 (N6671, N6642, N1359, N6008, N2271);
and AND4 (N6672, N6655, N4045, N6591, N6062);
buf BUF1 (N6673, N6650);
buf BUF1 (N6674, N6661);
or OR4 (N6675, N6665, N2457, N346, N1702);
or OR2 (N6676, N6668, N1612);
xor XOR2 (N6677, N6674, N715);
nor NOR4 (N6678, N6677, N5922, N3827, N2812);
nor NOR3 (N6679, N6669, N1981, N2320);
not NOT1 (N6680, N6678);
xor XOR2 (N6681, N6654, N169);
or OR4 (N6682, N6670, N4320, N5562, N2617);
xor XOR2 (N6683, N6671, N1443);
or OR2 (N6684, N6681, N6273);
nor NOR3 (N6685, N6676, N4981, N3271);
buf BUF1 (N6686, N6673);
nor NOR4 (N6687, N6679, N4416, N2619, N6278);
buf BUF1 (N6688, N6667);
or OR3 (N6689, N6687, N2115, N1288);
not NOT1 (N6690, N6682);
nor NOR2 (N6691, N6675, N216);
buf BUF1 (N6692, N6683);
not NOT1 (N6693, N6686);
buf BUF1 (N6694, N6688);
or OR2 (N6695, N6672, N4954);
nand NAND3 (N6696, N6690, N6099, N5146);
nor NOR4 (N6697, N6684, N2063, N5647, N308);
buf BUF1 (N6698, N6689);
and AND4 (N6699, N6694, N4094, N3842, N3024);
and AND2 (N6700, N6680, N5552);
nor NOR2 (N6701, N6700, N881);
nor NOR2 (N6702, N6699, N6288);
buf BUF1 (N6703, N6695);
nand NAND4 (N6704, N6698, N3202, N1314, N5564);
xor XOR2 (N6705, N6685, N1497);
nand NAND2 (N6706, N6697, N2684);
buf BUF1 (N6707, N6703);
buf BUF1 (N6708, N6701);
not NOT1 (N6709, N6691);
buf BUF1 (N6710, N6705);
not NOT1 (N6711, N6707);
nand NAND4 (N6712, N6704, N3628, N6703, N4783);
buf BUF1 (N6713, N6710);
nand NAND2 (N6714, N6706, N3012);
buf BUF1 (N6715, N6693);
xor XOR2 (N6716, N6714, N5070);
nor NOR4 (N6717, N6712, N1648, N6052, N5494);
buf BUF1 (N6718, N6716);
xor XOR2 (N6719, N6713, N4311);
or OR3 (N6720, N6715, N1670, N2067);
or OR2 (N6721, N6696, N1973);
nand NAND4 (N6722, N6709, N4410, N186, N312);
buf BUF1 (N6723, N6721);
xor XOR2 (N6724, N6692, N4188);
not NOT1 (N6725, N6718);
and AND2 (N6726, N6722, N5042);
and AND3 (N6727, N6719, N224, N3605);
nor NOR4 (N6728, N6708, N3968, N159, N2687);
nand NAND3 (N6729, N6725, N3036, N6487);
xor XOR2 (N6730, N6717, N4212);
xor XOR2 (N6731, N6711, N5655);
buf BUF1 (N6732, N6729);
xor XOR2 (N6733, N6702, N5176);
or OR3 (N6734, N6732, N1080, N6459);
and AND2 (N6735, N6730, N5478);
buf BUF1 (N6736, N6731);
nand NAND2 (N6737, N6734, N4226);
xor XOR2 (N6738, N6727, N2488);
buf BUF1 (N6739, N6720);
and AND4 (N6740, N6737, N5739, N1384, N2370);
not NOT1 (N6741, N6738);
nand NAND3 (N6742, N6741, N4789, N1832);
nand NAND2 (N6743, N6742, N4441);
nor NOR2 (N6744, N6733, N5928);
or OR3 (N6745, N6739, N2487, N2665);
or OR2 (N6746, N6745, N5837);
buf BUF1 (N6747, N6736);
nand NAND4 (N6748, N6723, N1033, N5865, N5130);
or OR2 (N6749, N6748, N1469);
nand NAND2 (N6750, N6735, N2401);
buf BUF1 (N6751, N6747);
not NOT1 (N6752, N6746);
nor NOR3 (N6753, N6743, N378, N3152);
and AND4 (N6754, N6744, N3478, N416, N5561);
not NOT1 (N6755, N6749);
nor NOR3 (N6756, N6740, N4630, N734);
nand NAND3 (N6757, N6755, N6300, N6143);
or OR2 (N6758, N6754, N1723);
nand NAND3 (N6759, N6728, N4266, N6223);
not NOT1 (N6760, N6757);
nor NOR2 (N6761, N6760, N4684);
or OR2 (N6762, N6750, N6337);
xor XOR2 (N6763, N6759, N2884);
buf BUF1 (N6764, N6724);
and AND2 (N6765, N6751, N4807);
nor NOR2 (N6766, N6763, N5582);
and AND2 (N6767, N6766, N546);
nor NOR2 (N6768, N6767, N6403);
buf BUF1 (N6769, N6756);
and AND4 (N6770, N6768, N290, N2656, N4411);
or OR2 (N6771, N6764, N965);
nor NOR2 (N6772, N6765, N4978);
and AND4 (N6773, N6726, N285, N5384, N609);
nor NOR4 (N6774, N6758, N5852, N6466, N4134);
nand NAND4 (N6775, N6769, N841, N4591, N879);
xor XOR2 (N6776, N6773, N910);
buf BUF1 (N6777, N6752);
nor NOR2 (N6778, N6777, N5478);
buf BUF1 (N6779, N6762);
or OR2 (N6780, N6779, N675);
nor NOR2 (N6781, N6775, N5159);
buf BUF1 (N6782, N6761);
nand NAND2 (N6783, N6782, N6616);
xor XOR2 (N6784, N6778, N454);
or OR3 (N6785, N6783, N5998, N456);
and AND4 (N6786, N6776, N3353, N2049, N4141);
nand NAND2 (N6787, N6781, N6272);
and AND2 (N6788, N6771, N301);
and AND3 (N6789, N6774, N5798, N5741);
nand NAND3 (N6790, N6780, N3182, N4740);
buf BUF1 (N6791, N6784);
buf BUF1 (N6792, N6770);
nor NOR4 (N6793, N6785, N498, N3628, N3782);
xor XOR2 (N6794, N6791, N4390);
nand NAND2 (N6795, N6753, N1740);
and AND2 (N6796, N6792, N3525);
not NOT1 (N6797, N6789);
nand NAND2 (N6798, N6788, N3192);
nor NOR3 (N6799, N6790, N224, N4911);
and AND2 (N6800, N6797, N202);
not NOT1 (N6801, N6786);
xor XOR2 (N6802, N6795, N2687);
or OR3 (N6803, N6798, N4113, N553);
buf BUF1 (N6804, N6799);
nand NAND4 (N6805, N6804, N4360, N5603, N5373);
nand NAND3 (N6806, N6796, N4698, N2988);
nand NAND3 (N6807, N6803, N5180, N4364);
or OR2 (N6808, N6787, N3473);
nor NOR3 (N6809, N6805, N6757, N622);
buf BUF1 (N6810, N6806);
xor XOR2 (N6811, N6800, N6208);
not NOT1 (N6812, N6801);
not NOT1 (N6813, N6807);
buf BUF1 (N6814, N6809);
xor XOR2 (N6815, N6793, N2707);
or OR2 (N6816, N6810, N5577);
buf BUF1 (N6817, N6815);
nor NOR4 (N6818, N6808, N4128, N4735, N5895);
or OR4 (N6819, N6814, N2542, N2271, N2629);
nand NAND3 (N6820, N6794, N3694, N1335);
buf BUF1 (N6821, N6812);
and AND2 (N6822, N6819, N4475);
not NOT1 (N6823, N6821);
not NOT1 (N6824, N6817);
and AND2 (N6825, N6811, N2934);
or OR3 (N6826, N6822, N2080, N4738);
nand NAND2 (N6827, N6802, N841);
buf BUF1 (N6828, N6772);
and AND2 (N6829, N6818, N6378);
nor NOR3 (N6830, N6820, N4833, N5416);
nand NAND2 (N6831, N6830, N225);
or OR2 (N6832, N6826, N391);
nor NOR2 (N6833, N6832, N2137);
nand NAND4 (N6834, N6813, N4724, N4876, N3125);
buf BUF1 (N6835, N6825);
and AND3 (N6836, N6823, N4521, N6429);
buf BUF1 (N6837, N6834);
or OR2 (N6838, N6827, N6524);
and AND3 (N6839, N6838, N4994, N1719);
or OR2 (N6840, N6836, N2327);
nor NOR3 (N6841, N6835, N6542, N3730);
or OR3 (N6842, N6828, N5170, N1663);
or OR4 (N6843, N6833, N5561, N4001, N2753);
buf BUF1 (N6844, N6831);
nor NOR3 (N6845, N6829, N5660, N3987);
xor XOR2 (N6846, N6844, N2344);
buf BUF1 (N6847, N6845);
nand NAND3 (N6848, N6846, N2163, N3930);
buf BUF1 (N6849, N6816);
buf BUF1 (N6850, N6842);
or OR2 (N6851, N6824, N1609);
buf BUF1 (N6852, N6843);
not NOT1 (N6853, N6848);
nand NAND3 (N6854, N6837, N4939, N2553);
nor NOR4 (N6855, N6850, N4978, N2257, N4067);
or OR4 (N6856, N6854, N6828, N3224, N6796);
xor XOR2 (N6857, N6847, N2144);
nand NAND2 (N6858, N6857, N5315);
and AND3 (N6859, N6853, N5593, N6243);
nor NOR2 (N6860, N6859, N5332);
xor XOR2 (N6861, N6840, N6363);
nor NOR3 (N6862, N6849, N4005, N2579);
or OR3 (N6863, N6851, N845, N721);
xor XOR2 (N6864, N6855, N4253);
xor XOR2 (N6865, N6863, N2005);
or OR2 (N6866, N6839, N2740);
not NOT1 (N6867, N6852);
or OR3 (N6868, N6841, N2311, N663);
not NOT1 (N6869, N6864);
xor XOR2 (N6870, N6861, N2691);
not NOT1 (N6871, N6866);
and AND4 (N6872, N6869, N52, N5206, N5166);
nor NOR4 (N6873, N6865, N3855, N1674, N5710);
nand NAND4 (N6874, N6873, N6594, N4019, N2041);
nor NOR2 (N6875, N6868, N2405);
buf BUF1 (N6876, N6872);
xor XOR2 (N6877, N6870, N5032);
buf BUF1 (N6878, N6875);
and AND4 (N6879, N6871, N24, N2130, N973);
nor NOR4 (N6880, N6867, N919, N6608, N213);
not NOT1 (N6881, N6862);
buf BUF1 (N6882, N6876);
xor XOR2 (N6883, N6858, N4044);
nand NAND4 (N6884, N6883, N4581, N6614, N3541);
nor NOR4 (N6885, N6882, N173, N1077, N4086);
buf BUF1 (N6886, N6879);
nor NOR4 (N6887, N6860, N3267, N3306, N6647);
not NOT1 (N6888, N6887);
and AND4 (N6889, N6888, N4254, N1567, N5917);
nor NOR2 (N6890, N6877, N4137);
nor NOR4 (N6891, N6885, N3543, N1689, N2618);
nor NOR2 (N6892, N6891, N1457);
or OR4 (N6893, N6892, N3681, N5408, N5700);
not NOT1 (N6894, N6874);
nor NOR3 (N6895, N6884, N3302, N6286);
xor XOR2 (N6896, N6893, N1012);
buf BUF1 (N6897, N6889);
xor XOR2 (N6898, N6890, N6373);
and AND2 (N6899, N6880, N5501);
not NOT1 (N6900, N6881);
not NOT1 (N6901, N6894);
xor XOR2 (N6902, N6897, N4903);
nand NAND3 (N6903, N6899, N2121, N1281);
not NOT1 (N6904, N6895);
buf BUF1 (N6905, N6903);
and AND3 (N6906, N6896, N3599, N2515);
nand NAND4 (N6907, N6856, N6474, N3412, N6722);
buf BUF1 (N6908, N6898);
and AND2 (N6909, N6907, N778);
nor NOR2 (N6910, N6902, N923);
xor XOR2 (N6911, N6908, N3730);
not NOT1 (N6912, N6906);
buf BUF1 (N6913, N6905);
and AND2 (N6914, N6901, N2938);
not NOT1 (N6915, N6886);
nand NAND4 (N6916, N6909, N3564, N5314, N2432);
nor NOR2 (N6917, N6900, N5327);
nor NOR2 (N6918, N6910, N3794);
nand NAND3 (N6919, N6918, N61, N5042);
xor XOR2 (N6920, N6919, N6471);
xor XOR2 (N6921, N6920, N674);
or OR2 (N6922, N6912, N3789);
buf BUF1 (N6923, N6914);
nor NOR3 (N6924, N6921, N5849, N5419);
xor XOR2 (N6925, N6904, N6069);
xor XOR2 (N6926, N6924, N6520);
xor XOR2 (N6927, N6916, N613);
nor NOR3 (N6928, N6911, N2534, N558);
nand NAND3 (N6929, N6922, N2055, N1908);
not NOT1 (N6930, N6915);
buf BUF1 (N6931, N6927);
nor NOR4 (N6932, N6923, N2952, N6127, N4421);
buf BUF1 (N6933, N6913);
nand NAND3 (N6934, N6878, N5370, N1660);
buf BUF1 (N6935, N6933);
not NOT1 (N6936, N6931);
xor XOR2 (N6937, N6930, N1641);
or OR2 (N6938, N6926, N1099);
nand NAND3 (N6939, N6932, N4676, N3759);
xor XOR2 (N6940, N6938, N3474);
xor XOR2 (N6941, N6917, N4859);
buf BUF1 (N6942, N6934);
buf BUF1 (N6943, N6936);
nor NOR2 (N6944, N6928, N3961);
and AND4 (N6945, N6941, N54, N237, N2318);
nand NAND2 (N6946, N6940, N79);
nor NOR4 (N6947, N6929, N905, N1736, N307);
buf BUF1 (N6948, N6935);
buf BUF1 (N6949, N6925);
or OR2 (N6950, N6944, N5729);
nor NOR4 (N6951, N6942, N4920, N1473, N825);
and AND4 (N6952, N6943, N2690, N4610, N6006);
not NOT1 (N6953, N6949);
buf BUF1 (N6954, N6939);
xor XOR2 (N6955, N6954, N1175);
not NOT1 (N6956, N6951);
or OR4 (N6957, N6952, N6219, N3445, N546);
buf BUF1 (N6958, N6945);
nand NAND2 (N6959, N6955, N2865);
and AND3 (N6960, N6946, N5209, N2524);
or OR3 (N6961, N6950, N4170, N1950);
nor NOR4 (N6962, N6961, N2580, N5718, N880);
not NOT1 (N6963, N6953);
nand NAND2 (N6964, N6957, N3523);
and AND2 (N6965, N6960, N4550);
nand NAND4 (N6966, N6947, N3628, N6119, N1608);
xor XOR2 (N6967, N6937, N2014);
or OR2 (N6968, N6964, N6276);
xor XOR2 (N6969, N6958, N5897);
nor NOR2 (N6970, N6968, N563);
not NOT1 (N6971, N6970);
buf BUF1 (N6972, N6965);
nand NAND3 (N6973, N6962, N3594, N1704);
not NOT1 (N6974, N6969);
nor NOR4 (N6975, N6974, N5702, N6086, N4436);
and AND3 (N6976, N6959, N101, N557);
xor XOR2 (N6977, N6973, N2254);
nor NOR3 (N6978, N6971, N3173, N4956);
or OR4 (N6979, N6975, N523, N4900, N939);
buf BUF1 (N6980, N6956);
and AND4 (N6981, N6978, N4272, N5180, N4106);
not NOT1 (N6982, N6977);
and AND4 (N6983, N6979, N3390, N3269, N1091);
buf BUF1 (N6984, N6981);
not NOT1 (N6985, N6980);
buf BUF1 (N6986, N6966);
nand NAND3 (N6987, N6976, N2044, N5135);
not NOT1 (N6988, N6982);
and AND2 (N6989, N6986, N3554);
nand NAND4 (N6990, N6984, N6948, N4113, N2410);
not NOT1 (N6991, N1534);
nor NOR4 (N6992, N6963, N3975, N482, N3459);
nor NOR3 (N6993, N6972, N1450, N5486);
buf BUF1 (N6994, N6992);
xor XOR2 (N6995, N6989, N1009);
nor NOR4 (N6996, N6983, N4103, N3, N1734);
not NOT1 (N6997, N6995);
not NOT1 (N6998, N6997);
or OR4 (N6999, N6996, N1471, N2064, N3685);
nor NOR2 (N7000, N6987, N794);
buf BUF1 (N7001, N6990);
nand NAND2 (N7002, N7000, N4267);
nand NAND4 (N7003, N6967, N4446, N6727, N1294);
not NOT1 (N7004, N6985);
and AND3 (N7005, N6998, N5639, N1994);
not NOT1 (N7006, N6991);
not NOT1 (N7007, N7006);
xor XOR2 (N7008, N7002, N3436);
nand NAND2 (N7009, N7005, N962);
or OR4 (N7010, N7009, N5167, N4699, N5404);
nand NAND3 (N7011, N6999, N1566, N5053);
nor NOR4 (N7012, N6993, N2060, N634, N3793);
not NOT1 (N7013, N6988);
not NOT1 (N7014, N7007);
and AND2 (N7015, N7001, N1505);
buf BUF1 (N7016, N7008);
and AND4 (N7017, N7016, N5317, N452, N5894);
xor XOR2 (N7018, N7011, N3936);
not NOT1 (N7019, N7014);
buf BUF1 (N7020, N7018);
and AND4 (N7021, N7012, N288, N547, N3658);
not NOT1 (N7022, N7021);
xor XOR2 (N7023, N7010, N4314);
nand NAND4 (N7024, N7003, N6959, N6188, N170);
or OR2 (N7025, N7004, N5916);
buf BUF1 (N7026, N7025);
nor NOR2 (N7027, N6994, N4224);
not NOT1 (N7028, N7020);
or OR4 (N7029, N7019, N1226, N3116, N5374);
or OR3 (N7030, N7028, N1442, N1566);
xor XOR2 (N7031, N7024, N2516);
or OR2 (N7032, N7017, N2396);
xor XOR2 (N7033, N7023, N3598);
nand NAND3 (N7034, N7032, N365, N1762);
nand NAND3 (N7035, N7015, N6652, N7000);
buf BUF1 (N7036, N7029);
or OR4 (N7037, N7036, N6608, N4885, N3166);
not NOT1 (N7038, N7026);
and AND2 (N7039, N7033, N3292);
or OR3 (N7040, N7039, N2912, N1257);
buf BUF1 (N7041, N7030);
nand NAND3 (N7042, N7037, N2130, N6729);
not NOT1 (N7043, N7040);
or OR3 (N7044, N7043, N3674, N4711);
nand NAND3 (N7045, N7041, N3095, N4127);
buf BUF1 (N7046, N7031);
and AND4 (N7047, N7034, N3465, N1681, N3149);
xor XOR2 (N7048, N7035, N3747);
xor XOR2 (N7049, N7047, N1661);
not NOT1 (N7050, N7044);
or OR4 (N7051, N7045, N4601, N6131, N6455);
and AND2 (N7052, N7027, N4076);
nor NOR3 (N7053, N7046, N5943, N920);
nand NAND3 (N7054, N7050, N5513, N5600);
or OR2 (N7055, N7052, N5582);
or OR2 (N7056, N7042, N4243);
or OR4 (N7057, N7054, N3321, N4901, N1490);
nor NOR2 (N7058, N7057, N1386);
nand NAND4 (N7059, N7022, N5681, N6554, N130);
and AND2 (N7060, N7059, N6628);
not NOT1 (N7061, N7058);
buf BUF1 (N7062, N7013);
buf BUF1 (N7063, N7055);
buf BUF1 (N7064, N7060);
or OR3 (N7065, N7051, N2896, N5099);
and AND3 (N7066, N7038, N4355, N6077);
xor XOR2 (N7067, N7048, N1795);
nand NAND3 (N7068, N7053, N259, N6332);
and AND3 (N7069, N7065, N1117, N2005);
nor NOR2 (N7070, N7068, N3556);
not NOT1 (N7071, N7069);
buf BUF1 (N7072, N7064);
xor XOR2 (N7073, N7056, N1553);
not NOT1 (N7074, N7073);
buf BUF1 (N7075, N7071);
nor NOR2 (N7076, N7063, N5960);
xor XOR2 (N7077, N7049, N899);
nand NAND4 (N7078, N7075, N1187, N1916, N1415);
not NOT1 (N7079, N7062);
nor NOR2 (N7080, N7066, N2558);
xor XOR2 (N7081, N7074, N2335);
nor NOR3 (N7082, N7077, N5658, N4830);
xor XOR2 (N7083, N7078, N742);
xor XOR2 (N7084, N7083, N4313);
nor NOR3 (N7085, N7079, N4247, N2607);
or OR4 (N7086, N7072, N3175, N4814, N5260);
not NOT1 (N7087, N7082);
nor NOR2 (N7088, N7061, N2436);
not NOT1 (N7089, N7087);
nor NOR3 (N7090, N7084, N4488, N4860);
and AND2 (N7091, N7076, N2826);
xor XOR2 (N7092, N7088, N115);
nand NAND2 (N7093, N7067, N3995);
xor XOR2 (N7094, N7093, N6530);
nor NOR4 (N7095, N7086, N704, N390, N3934);
buf BUF1 (N7096, N7095);
nor NOR2 (N7097, N7091, N6703);
nor NOR2 (N7098, N7097, N4285);
or OR2 (N7099, N7090, N1641);
and AND4 (N7100, N7092, N815, N1896, N6326);
buf BUF1 (N7101, N7089);
xor XOR2 (N7102, N7098, N4871);
buf BUF1 (N7103, N7070);
buf BUF1 (N7104, N7094);
nand NAND4 (N7105, N7081, N5029, N3939, N514);
not NOT1 (N7106, N7101);
or OR2 (N7107, N7104, N186);
and AND3 (N7108, N7102, N6400, N4870);
and AND3 (N7109, N7108, N766, N2153);
nor NOR2 (N7110, N7103, N5536);
nor NOR4 (N7111, N7100, N5913, N3940, N2358);
xor XOR2 (N7112, N7099, N3840);
xor XOR2 (N7113, N7085, N6342);
buf BUF1 (N7114, N7111);
and AND4 (N7115, N7080, N4781, N6866, N1574);
nor NOR2 (N7116, N7110, N6718);
and AND2 (N7117, N7116, N326);
or OR2 (N7118, N7106, N6667);
or OR4 (N7119, N7117, N1762, N2819, N2426);
or OR2 (N7120, N7119, N1305);
nor NOR2 (N7121, N7107, N5639);
nor NOR2 (N7122, N7114, N307);
not NOT1 (N7123, N7096);
or OR4 (N7124, N7122, N1170, N2961, N5627);
or OR3 (N7125, N7105, N544, N1696);
not NOT1 (N7126, N7115);
nor NOR4 (N7127, N7113, N323, N1000, N4997);
nor NOR4 (N7128, N7109, N4074, N885, N5967);
or OR4 (N7129, N7128, N3508, N2937, N2873);
not NOT1 (N7130, N7118);
nand NAND4 (N7131, N7127, N661, N477, N2924);
or OR2 (N7132, N7130, N3646);
nand NAND4 (N7133, N7121, N1520, N4635, N6716);
nor NOR4 (N7134, N7120, N2907, N2522, N3758);
nand NAND2 (N7135, N7131, N3981);
nor NOR3 (N7136, N7133, N1254, N6224);
or OR3 (N7137, N7136, N1552, N4145);
xor XOR2 (N7138, N7134, N1250);
nor NOR2 (N7139, N7129, N2183);
or OR3 (N7140, N7132, N5678, N202);
and AND2 (N7141, N7123, N7006);
nor NOR4 (N7142, N7139, N1909, N5009, N700);
buf BUF1 (N7143, N7138);
buf BUF1 (N7144, N7126);
not NOT1 (N7145, N7140);
nand NAND4 (N7146, N7142, N3623, N1337, N3273);
xor XOR2 (N7147, N7143, N6260);
or OR4 (N7148, N7137, N6103, N4143, N2187);
or OR3 (N7149, N7135, N4829, N6927);
nand NAND2 (N7150, N7112, N4981);
or OR2 (N7151, N7144, N5988);
not NOT1 (N7152, N7147);
buf BUF1 (N7153, N7152);
buf BUF1 (N7154, N7145);
not NOT1 (N7155, N7151);
nand NAND3 (N7156, N7155, N1303, N3748);
buf BUF1 (N7157, N7156);
nand NAND3 (N7158, N7148, N256, N2556);
buf BUF1 (N7159, N7146);
nand NAND2 (N7160, N7141, N6896);
and AND3 (N7161, N7154, N5466, N5988);
and AND4 (N7162, N7153, N3053, N589, N2684);
buf BUF1 (N7163, N7150);
or OR4 (N7164, N7125, N5414, N83, N3082);
nand NAND4 (N7165, N7161, N2062, N4525, N6028);
buf BUF1 (N7166, N7157);
buf BUF1 (N7167, N7166);
xor XOR2 (N7168, N7124, N3262);
xor XOR2 (N7169, N7165, N1603);
buf BUF1 (N7170, N7149);
nand NAND3 (N7171, N7167, N2800, N6809);
or OR4 (N7172, N7159, N7131, N7082, N6405);
nor NOR3 (N7173, N7160, N5181, N1553);
nand NAND3 (N7174, N7162, N5926, N799);
nand NAND2 (N7175, N7163, N4026);
not NOT1 (N7176, N7170);
not NOT1 (N7177, N7176);
xor XOR2 (N7178, N7173, N1000);
and AND2 (N7179, N7168, N5630);
buf BUF1 (N7180, N7158);
buf BUF1 (N7181, N7164);
buf BUF1 (N7182, N7171);
nand NAND4 (N7183, N7175, N6746, N3037, N6216);
or OR2 (N7184, N7182, N1906);
or OR3 (N7185, N7180, N6576, N804);
or OR3 (N7186, N7174, N2631, N2932);
or OR4 (N7187, N7169, N3516, N521, N4675);
and AND4 (N7188, N7181, N1290, N6465, N59);
buf BUF1 (N7189, N7186);
or OR4 (N7190, N7177, N4190, N6143, N6191);
buf BUF1 (N7191, N7178);
nand NAND3 (N7192, N7185, N6336, N3311);
xor XOR2 (N7193, N7190, N3726);
or OR4 (N7194, N7183, N1284, N3005, N6677);
xor XOR2 (N7195, N7189, N4714);
nand NAND4 (N7196, N7184, N6175, N1421, N3499);
xor XOR2 (N7197, N7195, N6);
not NOT1 (N7198, N7188);
or OR2 (N7199, N7198, N3797);
or OR4 (N7200, N7194, N1320, N2111, N96);
not NOT1 (N7201, N7200);
nor NOR4 (N7202, N7201, N2759, N1607, N3771);
buf BUF1 (N7203, N7196);
and AND4 (N7204, N7203, N1232, N5210, N2194);
nor NOR3 (N7205, N7202, N4229, N7087);
buf BUF1 (N7206, N7193);
or OR3 (N7207, N7205, N4464, N1614);
buf BUF1 (N7208, N7187);
xor XOR2 (N7209, N7199, N290);
or OR4 (N7210, N7206, N5751, N1671, N2415);
xor XOR2 (N7211, N7204, N3722);
and AND2 (N7212, N7210, N1570);
xor XOR2 (N7213, N7191, N3319);
nor NOR4 (N7214, N7211, N3595, N4121, N3894);
buf BUF1 (N7215, N7214);
and AND3 (N7216, N7192, N7054, N6731);
and AND2 (N7217, N7213, N3666);
not NOT1 (N7218, N7215);
xor XOR2 (N7219, N7218, N4833);
xor XOR2 (N7220, N7217, N3176);
nand NAND3 (N7221, N7197, N3691, N1120);
nand NAND3 (N7222, N7212, N2751, N4449);
and AND3 (N7223, N7220, N5369, N1899);
nor NOR4 (N7224, N7216, N7174, N2497, N1344);
buf BUF1 (N7225, N7219);
and AND2 (N7226, N7225, N689);
and AND2 (N7227, N7221, N1065);
buf BUF1 (N7228, N7227);
nand NAND4 (N7229, N7224, N4282, N6798, N4432);
or OR3 (N7230, N7228, N3131, N2791);
xor XOR2 (N7231, N7226, N5652);
xor XOR2 (N7232, N7209, N5757);
buf BUF1 (N7233, N7172);
nand NAND2 (N7234, N7223, N3983);
not NOT1 (N7235, N7229);
buf BUF1 (N7236, N7222);
not NOT1 (N7237, N7235);
and AND4 (N7238, N7233, N2873, N6070, N5293);
xor XOR2 (N7239, N7236, N3323);
nor NOR4 (N7240, N7230, N5850, N7194, N3680);
not NOT1 (N7241, N7179);
not NOT1 (N7242, N7240);
buf BUF1 (N7243, N7242);
or OR2 (N7244, N7241, N6715);
nor NOR4 (N7245, N7234, N1060, N4614, N3817);
or OR4 (N7246, N7231, N4708, N2862, N1696);
nor NOR3 (N7247, N7208, N1176, N656);
and AND2 (N7248, N7246, N2822);
and AND3 (N7249, N7243, N4894, N4813);
buf BUF1 (N7250, N7245);
not NOT1 (N7251, N7237);
xor XOR2 (N7252, N7207, N1799);
and AND2 (N7253, N7250, N288);
not NOT1 (N7254, N7248);
or OR3 (N7255, N7239, N4937, N4675);
and AND4 (N7256, N7254, N5804, N3943, N3354);
nor NOR4 (N7257, N7249, N6038, N4174, N2002);
xor XOR2 (N7258, N7232, N1090);
nor NOR4 (N7259, N7255, N6136, N223, N5690);
nor NOR4 (N7260, N7257, N6647, N4466, N1545);
not NOT1 (N7261, N7244);
nand NAND3 (N7262, N7261, N3949, N4874);
buf BUF1 (N7263, N7259);
nor NOR3 (N7264, N7262, N4402, N5398);
not NOT1 (N7265, N7238);
nor NOR4 (N7266, N7251, N6408, N5203, N3725);
and AND2 (N7267, N7247, N6353);
xor XOR2 (N7268, N7260, N1325);
nand NAND4 (N7269, N7268, N5218, N503, N3902);
or OR2 (N7270, N7252, N2761);
nand NAND4 (N7271, N7263, N566, N1766, N836);
xor XOR2 (N7272, N7253, N6657);
nor NOR2 (N7273, N7256, N2271);
nand NAND2 (N7274, N7270, N1445);
buf BUF1 (N7275, N7271);
nand NAND3 (N7276, N7265, N397, N5475);
nand NAND3 (N7277, N7258, N6800, N3919);
and AND4 (N7278, N7274, N4151, N6449, N6288);
and AND2 (N7279, N7272, N6483);
or OR2 (N7280, N7279, N432);
xor XOR2 (N7281, N7267, N2396);
buf BUF1 (N7282, N7275);
buf BUF1 (N7283, N7273);
not NOT1 (N7284, N7277);
buf BUF1 (N7285, N7283);
nand NAND2 (N7286, N7278, N6893);
not NOT1 (N7287, N7281);
buf BUF1 (N7288, N7280);
nand NAND3 (N7289, N7285, N4090, N4806);
or OR2 (N7290, N7269, N3969);
not NOT1 (N7291, N7289);
xor XOR2 (N7292, N7282, N472);
or OR4 (N7293, N7284, N5281, N1936, N5960);
buf BUF1 (N7294, N7288);
xor XOR2 (N7295, N7276, N159);
buf BUF1 (N7296, N7294);
not NOT1 (N7297, N7286);
and AND3 (N7298, N7295, N952, N4541);
or OR3 (N7299, N7297, N869, N554);
not NOT1 (N7300, N7290);
nor NOR3 (N7301, N7292, N4779, N153);
and AND3 (N7302, N7293, N2961, N5846);
xor XOR2 (N7303, N7298, N1246);
xor XOR2 (N7304, N7301, N5457);
and AND3 (N7305, N7266, N5307, N1506);
not NOT1 (N7306, N7305);
xor XOR2 (N7307, N7291, N2077);
nand NAND3 (N7308, N7287, N6430, N235);
nand NAND3 (N7309, N7306, N4666, N4999);
not NOT1 (N7310, N7304);
buf BUF1 (N7311, N7309);
buf BUF1 (N7312, N7296);
not NOT1 (N7313, N7302);
or OR4 (N7314, N7311, N3116, N4849, N1637);
or OR4 (N7315, N7314, N178, N1378, N5192);
not NOT1 (N7316, N7315);
nor NOR3 (N7317, N7299, N4125, N5691);
buf BUF1 (N7318, N7310);
nand NAND2 (N7319, N7317, N709);
xor XOR2 (N7320, N7312, N842);
or OR2 (N7321, N7264, N2920);
nand NAND2 (N7322, N7300, N3614);
xor XOR2 (N7323, N7316, N59);
buf BUF1 (N7324, N7322);
and AND3 (N7325, N7319, N6484, N6732);
nor NOR4 (N7326, N7320, N965, N1875, N6067);
nand NAND4 (N7327, N7325, N6095, N456, N4595);
nor NOR2 (N7328, N7318, N2508);
or OR2 (N7329, N7308, N1969);
and AND3 (N7330, N7324, N522, N2081);
xor XOR2 (N7331, N7326, N2544);
nor NOR4 (N7332, N7331, N6419, N4975, N474);
xor XOR2 (N7333, N7327, N4717);
nand NAND2 (N7334, N7328, N6629);
nor NOR3 (N7335, N7303, N2935, N3830);
buf BUF1 (N7336, N7335);
xor XOR2 (N7337, N7334, N3647);
xor XOR2 (N7338, N7329, N6858);
or OR2 (N7339, N7337, N6588);
nor NOR4 (N7340, N7332, N6100, N2272, N953);
xor XOR2 (N7341, N7336, N408);
and AND3 (N7342, N7333, N5391, N5774);
and AND4 (N7343, N7341, N926, N6791, N6746);
nand NAND2 (N7344, N7339, N397);
nor NOR4 (N7345, N7313, N1598, N461, N6915);
or OR2 (N7346, N7330, N1833);
buf BUF1 (N7347, N7346);
not NOT1 (N7348, N7345);
not NOT1 (N7349, N7344);
nor NOR2 (N7350, N7349, N2795);
nor NOR2 (N7351, N7348, N4864);
nor NOR4 (N7352, N7323, N2452, N2456, N1124);
and AND3 (N7353, N7350, N5721, N2430);
nand NAND3 (N7354, N7343, N6389, N2690);
nor NOR3 (N7355, N7347, N3001, N5561);
nand NAND3 (N7356, N7307, N6351, N3149);
nand NAND3 (N7357, N7321, N5335, N1192);
nand NAND3 (N7358, N7354, N1309, N3798);
not NOT1 (N7359, N7356);
not NOT1 (N7360, N7342);
nor NOR3 (N7361, N7360, N4286, N2880);
not NOT1 (N7362, N7340);
nand NAND3 (N7363, N7362, N7077, N2139);
nor NOR4 (N7364, N7351, N3030, N7302, N2100);
buf BUF1 (N7365, N7357);
not NOT1 (N7366, N7363);
nand NAND4 (N7367, N7361, N1326, N355, N6586);
buf BUF1 (N7368, N7367);
xor XOR2 (N7369, N7364, N721);
not NOT1 (N7370, N7368);
not NOT1 (N7371, N7365);
buf BUF1 (N7372, N7369);
nor NOR4 (N7373, N7338, N3588, N6433, N254);
or OR4 (N7374, N7352, N3871, N1278, N1476);
nor NOR3 (N7375, N7353, N2842, N6835);
xor XOR2 (N7376, N7374, N3825);
buf BUF1 (N7377, N7366);
nor NOR2 (N7378, N7377, N6247);
not NOT1 (N7379, N7372);
not NOT1 (N7380, N7358);
or OR4 (N7381, N7380, N1293, N129, N5681);
xor XOR2 (N7382, N7379, N4769);
or OR4 (N7383, N7359, N2865, N5196, N4581);
nor NOR4 (N7384, N7355, N6188, N5855, N4540);
buf BUF1 (N7385, N7381);
and AND4 (N7386, N7383, N7220, N2130, N1636);
and AND4 (N7387, N7384, N4235, N1801, N2766);
nand NAND4 (N7388, N7375, N666, N3911, N23);
not NOT1 (N7389, N7385);
nand NAND3 (N7390, N7382, N4824, N4923);
and AND2 (N7391, N7371, N298);
and AND3 (N7392, N7387, N1918, N586);
buf BUF1 (N7393, N7386);
xor XOR2 (N7394, N7391, N560);
buf BUF1 (N7395, N7394);
and AND2 (N7396, N7378, N20);
xor XOR2 (N7397, N7395, N948);
buf BUF1 (N7398, N7393);
and AND3 (N7399, N7373, N6123, N4906);
buf BUF1 (N7400, N7389);
xor XOR2 (N7401, N7396, N4768);
xor XOR2 (N7402, N7390, N5860);
not NOT1 (N7403, N7398);
nand NAND3 (N7404, N7388, N5033, N5975);
not NOT1 (N7405, N7401);
buf BUF1 (N7406, N7404);
nor NOR3 (N7407, N7400, N5665, N422);
or OR3 (N7408, N7397, N4761, N4496);
buf BUF1 (N7409, N7392);
nand NAND4 (N7410, N7406, N1892, N1846, N6801);
nand NAND3 (N7411, N7405, N5749, N4912);
nand NAND3 (N7412, N7410, N1326, N2035);
nor NOR3 (N7413, N7402, N39, N274);
buf BUF1 (N7414, N7409);
or OR4 (N7415, N7408, N6671, N1334, N7325);
and AND2 (N7416, N7414, N3230);
not NOT1 (N7417, N7416);
xor XOR2 (N7418, N7399, N401);
nand NAND2 (N7419, N7376, N1226);
xor XOR2 (N7420, N7417, N2397);
buf BUF1 (N7421, N7411);
buf BUF1 (N7422, N7421);
not NOT1 (N7423, N7403);
not NOT1 (N7424, N7419);
buf BUF1 (N7425, N7415);
nor NOR2 (N7426, N7407, N3772);
and AND3 (N7427, N7412, N3509, N3059);
or OR3 (N7428, N7427, N6713, N639);
nor NOR3 (N7429, N7423, N6959, N7256);
or OR2 (N7430, N7428, N5777);
xor XOR2 (N7431, N7426, N1979);
xor XOR2 (N7432, N7420, N5318);
buf BUF1 (N7433, N7430);
nor NOR3 (N7434, N7424, N921, N551);
xor XOR2 (N7435, N7413, N5701);
or OR4 (N7436, N7435, N7124, N3645, N397);
and AND3 (N7437, N7432, N5345, N1985);
or OR4 (N7438, N7370, N1417, N194, N7065);
not NOT1 (N7439, N7422);
and AND3 (N7440, N7439, N1399, N4616);
nand NAND2 (N7441, N7440, N2016);
or OR4 (N7442, N7437, N808, N663, N4681);
xor XOR2 (N7443, N7442, N144);
nand NAND2 (N7444, N7443, N2762);
nand NAND4 (N7445, N7418, N6238, N353, N3821);
nand NAND4 (N7446, N7436, N6879, N5603, N6477);
xor XOR2 (N7447, N7441, N7003);
nor NOR2 (N7448, N7438, N7357);
or OR3 (N7449, N7429, N4618, N7352);
and AND3 (N7450, N7447, N6433, N7400);
nor NOR3 (N7451, N7434, N231, N1827);
nand NAND4 (N7452, N7431, N1890, N106, N6256);
buf BUF1 (N7453, N7444);
xor XOR2 (N7454, N7453, N6606);
not NOT1 (N7455, N7448);
or OR2 (N7456, N7445, N5794);
nand NAND4 (N7457, N7450, N1471, N1936, N3772);
nor NOR2 (N7458, N7452, N4116);
not NOT1 (N7459, N7457);
nor NOR2 (N7460, N7425, N376);
buf BUF1 (N7461, N7456);
and AND3 (N7462, N7446, N3586, N3996);
or OR4 (N7463, N7460, N4837, N5487, N6696);
xor XOR2 (N7464, N7458, N6682);
nand NAND3 (N7465, N7463, N3546, N677);
buf BUF1 (N7466, N7465);
or OR4 (N7467, N7433, N2311, N3147, N645);
and AND2 (N7468, N7462, N5768);
xor XOR2 (N7469, N7467, N2307);
xor XOR2 (N7470, N7454, N3926);
and AND3 (N7471, N7466, N1892, N6939);
or OR3 (N7472, N7469, N2451, N2435);
and AND4 (N7473, N7464, N4497, N672, N452);
and AND4 (N7474, N7473, N3941, N3683, N6869);
nor NOR4 (N7475, N7461, N3597, N6426, N6052);
nor NOR4 (N7476, N7451, N2497, N748, N7373);
xor XOR2 (N7477, N7459, N738);
or OR4 (N7478, N7471, N5989, N2848, N2323);
and AND3 (N7479, N7449, N4550, N1653);
nor NOR4 (N7480, N7472, N2633, N1373, N2920);
and AND4 (N7481, N7455, N3165, N2296, N4157);
and AND2 (N7482, N7481, N4308);
xor XOR2 (N7483, N7477, N1294);
nand NAND2 (N7484, N7468, N2020);
xor XOR2 (N7485, N7484, N6328);
buf BUF1 (N7486, N7470);
not NOT1 (N7487, N7478);
not NOT1 (N7488, N7485);
nor NOR2 (N7489, N7480, N5589);
buf BUF1 (N7490, N7474);
or OR3 (N7491, N7486, N2955, N4926);
buf BUF1 (N7492, N7482);
not NOT1 (N7493, N7491);
not NOT1 (N7494, N7476);
xor XOR2 (N7495, N7479, N7286);
nor NOR4 (N7496, N7488, N3239, N7043, N7018);
buf BUF1 (N7497, N7494);
nand NAND4 (N7498, N7489, N391, N3050, N3235);
nor NOR4 (N7499, N7495, N2642, N5822, N4617);
nor NOR2 (N7500, N7483, N3281);
not NOT1 (N7501, N7497);
or OR4 (N7502, N7500, N4945, N5203, N2479);
not NOT1 (N7503, N7487);
not NOT1 (N7504, N7498);
buf BUF1 (N7505, N7501);
nor NOR2 (N7506, N7490, N5558);
not NOT1 (N7507, N7475);
nor NOR4 (N7508, N7493, N5757, N5366, N5101);
or OR2 (N7509, N7507, N6221);
nand NAND3 (N7510, N7506, N7299, N7265);
xor XOR2 (N7511, N7502, N739);
buf BUF1 (N7512, N7508);
buf BUF1 (N7513, N7503);
and AND3 (N7514, N7499, N4793, N2453);
buf BUF1 (N7515, N7492);
and AND3 (N7516, N7505, N3179, N1464);
nand NAND2 (N7517, N7511, N331);
nor NOR2 (N7518, N7504, N3533);
and AND4 (N7519, N7515, N3071, N5047, N1372);
and AND2 (N7520, N7496, N6903);
xor XOR2 (N7521, N7520, N3807);
and AND4 (N7522, N7513, N2800, N5255, N218);
xor XOR2 (N7523, N7522, N160);
or OR3 (N7524, N7519, N361, N6548);
not NOT1 (N7525, N7514);
or OR4 (N7526, N7516, N581, N4129, N6678);
buf BUF1 (N7527, N7518);
xor XOR2 (N7528, N7521, N120);
xor XOR2 (N7529, N7528, N6490);
or OR2 (N7530, N7529, N6743);
nand NAND2 (N7531, N7524, N17);
buf BUF1 (N7532, N7510);
nand NAND4 (N7533, N7525, N3827, N2803, N4789);
or OR4 (N7534, N7531, N744, N4091, N1671);
nand NAND4 (N7535, N7527, N3492, N4299, N5943);
nand NAND3 (N7536, N7530, N1472, N4569);
xor XOR2 (N7537, N7535, N2269);
and AND3 (N7538, N7523, N4353, N3164);
not NOT1 (N7539, N7517);
buf BUF1 (N7540, N7534);
not NOT1 (N7541, N7532);
buf BUF1 (N7542, N7536);
nand NAND4 (N7543, N7539, N4036, N7102, N5780);
or OR3 (N7544, N7538, N3476, N5753);
xor XOR2 (N7545, N7544, N3870);
xor XOR2 (N7546, N7542, N7148);
nor NOR2 (N7547, N7540, N6000);
buf BUF1 (N7548, N7546);
xor XOR2 (N7549, N7512, N1833);
xor XOR2 (N7550, N7537, N4092);
nand NAND3 (N7551, N7547, N6141, N1340);
nand NAND2 (N7552, N7541, N319);
buf BUF1 (N7553, N7526);
nand NAND3 (N7554, N7552, N3716, N5380);
not NOT1 (N7555, N7554);
nor NOR2 (N7556, N7555, N4558);
nand NAND3 (N7557, N7533, N5285, N5844);
xor XOR2 (N7558, N7548, N5804);
nand NAND3 (N7559, N7543, N7439, N4362);
nand NAND4 (N7560, N7550, N3434, N716, N1026);
not NOT1 (N7561, N7556);
xor XOR2 (N7562, N7545, N6801);
xor XOR2 (N7563, N7559, N5620);
not NOT1 (N7564, N7509);
xor XOR2 (N7565, N7560, N2337);
not NOT1 (N7566, N7565);
and AND2 (N7567, N7566, N6395);
nand NAND2 (N7568, N7567, N3419);
xor XOR2 (N7569, N7564, N2417);
or OR4 (N7570, N7558, N2591, N303, N3636);
not NOT1 (N7571, N7563);
buf BUF1 (N7572, N7570);
not NOT1 (N7573, N7549);
xor XOR2 (N7574, N7572, N7245);
or OR4 (N7575, N7561, N5725, N7083, N6101);
not NOT1 (N7576, N7571);
nor NOR3 (N7577, N7573, N5780, N6154);
or OR3 (N7578, N7576, N3577, N5810);
or OR3 (N7579, N7551, N2832, N7327);
xor XOR2 (N7580, N7568, N1156);
nand NAND2 (N7581, N7579, N1595);
nand NAND4 (N7582, N7553, N5306, N1912, N1946);
xor XOR2 (N7583, N7569, N5738);
nor NOR2 (N7584, N7578, N2929);
xor XOR2 (N7585, N7575, N6369);
nor NOR3 (N7586, N7581, N4240, N1547);
or OR4 (N7587, N7583, N5780, N3000, N2158);
buf BUF1 (N7588, N7584);
xor XOR2 (N7589, N7557, N7532);
not NOT1 (N7590, N7582);
nand NAND3 (N7591, N7587, N5502, N4737);
nand NAND4 (N7592, N7588, N3839, N5661, N2919);
xor XOR2 (N7593, N7574, N2450);
nor NOR4 (N7594, N7593, N3918, N4784, N7039);
nor NOR3 (N7595, N7590, N7309, N656);
nor NOR4 (N7596, N7585, N7246, N6235, N4580);
or OR3 (N7597, N7592, N678, N5113);
nand NAND2 (N7598, N7580, N2390);
or OR4 (N7599, N7589, N75, N4716, N5547);
or OR2 (N7600, N7562, N1296);
nand NAND3 (N7601, N7595, N2913, N3183);
xor XOR2 (N7602, N7600, N4400);
xor XOR2 (N7603, N7601, N6599);
xor XOR2 (N7604, N7598, N4044);
or OR3 (N7605, N7597, N5612, N7074);
not NOT1 (N7606, N7594);
and AND4 (N7607, N7596, N5967, N6237, N1461);
nor NOR3 (N7608, N7607, N3088, N7572);
nand NAND2 (N7609, N7605, N1152);
and AND2 (N7610, N7577, N3434);
nor NOR2 (N7611, N7591, N1967);
not NOT1 (N7612, N7606);
not NOT1 (N7613, N7602);
or OR3 (N7614, N7612, N7167, N6960);
buf BUF1 (N7615, N7609);
or OR2 (N7616, N7604, N3680);
buf BUF1 (N7617, N7616);
nand NAND3 (N7618, N7608, N3372, N2786);
and AND3 (N7619, N7603, N7415, N942);
or OR3 (N7620, N7586, N1003, N1849);
and AND2 (N7621, N7620, N6890);
xor XOR2 (N7622, N7610, N1004);
not NOT1 (N7623, N7613);
xor XOR2 (N7624, N7621, N2886);
nand NAND3 (N7625, N7622, N2555, N1983);
not NOT1 (N7626, N7617);
or OR3 (N7627, N7619, N6696, N2280);
or OR2 (N7628, N7624, N4877);
or OR4 (N7629, N7599, N4497, N1041, N7501);
or OR4 (N7630, N7627, N7210, N1295, N6337);
xor XOR2 (N7631, N7611, N5147);
or OR3 (N7632, N7625, N1848, N2074);
xor XOR2 (N7633, N7618, N342);
and AND3 (N7634, N7632, N1019, N400);
nor NOR4 (N7635, N7634, N4657, N6276, N2540);
and AND4 (N7636, N7631, N5798, N4775, N5039);
xor XOR2 (N7637, N7615, N156);
nand NAND2 (N7638, N7636, N3568);
buf BUF1 (N7639, N7635);
nor NOR2 (N7640, N7614, N4602);
nor NOR4 (N7641, N7639, N1771, N3770, N2377);
nor NOR4 (N7642, N7623, N4430, N4456, N871);
or OR4 (N7643, N7637, N7526, N6872, N6310);
not NOT1 (N7644, N7628);
nand NAND4 (N7645, N7640, N466, N6502, N458);
not NOT1 (N7646, N7630);
buf BUF1 (N7647, N7642);
buf BUF1 (N7648, N7646);
nand NAND2 (N7649, N7647, N2117);
not NOT1 (N7650, N7626);
buf BUF1 (N7651, N7645);
or OR3 (N7652, N7629, N5839, N4238);
buf BUF1 (N7653, N7651);
nor NOR4 (N7654, N7649, N4616, N5325, N6621);
or OR4 (N7655, N7650, N547, N5960, N904);
and AND2 (N7656, N7641, N884);
nor NOR4 (N7657, N7656, N6413, N4223, N5067);
nand NAND4 (N7658, N7655, N6512, N2520, N6008);
not NOT1 (N7659, N7653);
and AND3 (N7660, N7654, N5032, N6190);
buf BUF1 (N7661, N7643);
or OR4 (N7662, N7652, N1484, N3993, N3489);
nand NAND3 (N7663, N7662, N3371, N1975);
buf BUF1 (N7664, N7633);
or OR2 (N7665, N7657, N5853);
xor XOR2 (N7666, N7661, N2503);
or OR3 (N7667, N7663, N7083, N2689);
and AND3 (N7668, N7659, N5195, N6106);
buf BUF1 (N7669, N7668);
xor XOR2 (N7670, N7660, N2619);
not NOT1 (N7671, N7666);
not NOT1 (N7672, N7667);
not NOT1 (N7673, N7665);
buf BUF1 (N7674, N7673);
buf BUF1 (N7675, N7648);
nor NOR2 (N7676, N7674, N2708);
not NOT1 (N7677, N7644);
xor XOR2 (N7678, N7677, N743);
xor XOR2 (N7679, N7669, N4463);
nor NOR2 (N7680, N7664, N2367);
not NOT1 (N7681, N7638);
nor NOR2 (N7682, N7658, N4412);
buf BUF1 (N7683, N7671);
not NOT1 (N7684, N7675);
xor XOR2 (N7685, N7676, N5738);
nor NOR2 (N7686, N7670, N6890);
nor NOR3 (N7687, N7679, N5778, N5071);
and AND3 (N7688, N7678, N7332, N6580);
or OR4 (N7689, N7686, N4986, N793, N203);
nor NOR2 (N7690, N7685, N3313);
xor XOR2 (N7691, N7680, N7613);
and AND3 (N7692, N7690, N4405, N253);
nand NAND2 (N7693, N7691, N5249);
xor XOR2 (N7694, N7672, N4624);
nor NOR3 (N7695, N7688, N6905, N610);
buf BUF1 (N7696, N7692);
nand NAND2 (N7697, N7695, N2460);
and AND2 (N7698, N7693, N901);
or OR2 (N7699, N7698, N2213);
or OR2 (N7700, N7681, N6054);
and AND4 (N7701, N7682, N2507, N2634, N3958);
nor NOR4 (N7702, N7683, N5751, N5305, N2755);
nor NOR3 (N7703, N7699, N3075, N2512);
not NOT1 (N7704, N7689);
xor XOR2 (N7705, N7703, N6290);
xor XOR2 (N7706, N7701, N5321);
and AND2 (N7707, N7694, N7285);
xor XOR2 (N7708, N7700, N1468);
nor NOR3 (N7709, N7697, N2327, N5509);
buf BUF1 (N7710, N7704);
nor NOR2 (N7711, N7684, N2722);
buf BUF1 (N7712, N7687);
nand NAND4 (N7713, N7711, N3503, N2316, N3942);
and AND2 (N7714, N7709, N6744);
not NOT1 (N7715, N7713);
not NOT1 (N7716, N7705);
not NOT1 (N7717, N7706);
and AND2 (N7718, N7708, N6986);
xor XOR2 (N7719, N7702, N5049);
or OR3 (N7720, N7718, N3313, N4547);
xor XOR2 (N7721, N7712, N5442);
xor XOR2 (N7722, N7720, N1458);
not NOT1 (N7723, N7714);
xor XOR2 (N7724, N7722, N1592);
xor XOR2 (N7725, N7723, N3379);
and AND4 (N7726, N7719, N5987, N4358, N1404);
nor NOR3 (N7727, N7726, N1247, N7423);
nand NAND4 (N7728, N7696, N3404, N6757, N1001);
buf BUF1 (N7729, N7725);
or OR2 (N7730, N7707, N6756);
and AND4 (N7731, N7727, N7228, N1854, N4358);
or OR2 (N7732, N7715, N2543);
or OR4 (N7733, N7710, N5067, N3249, N5032);
xor XOR2 (N7734, N7731, N4590);
and AND4 (N7735, N7717, N3272, N4173, N2860);
or OR3 (N7736, N7729, N5015, N2900);
nor NOR4 (N7737, N7716, N6117, N617, N167);
buf BUF1 (N7738, N7721);
xor XOR2 (N7739, N7736, N6890);
not NOT1 (N7740, N7738);
or OR4 (N7741, N7737, N2128, N5084, N4585);
and AND3 (N7742, N7733, N567, N5436);
nor NOR2 (N7743, N7732, N1166);
or OR3 (N7744, N7724, N4885, N3926);
or OR2 (N7745, N7743, N749);
and AND4 (N7746, N7730, N2116, N4660, N919);
nand NAND2 (N7747, N7739, N6490);
buf BUF1 (N7748, N7741);
xor XOR2 (N7749, N7744, N5556);
xor XOR2 (N7750, N7746, N3656);
buf BUF1 (N7751, N7740);
nand NAND3 (N7752, N7751, N5765, N2216);
or OR3 (N7753, N7742, N3597, N5149);
xor XOR2 (N7754, N7728, N5464);
and AND4 (N7755, N7745, N7741, N3991, N7429);
nand NAND2 (N7756, N7753, N6977);
xor XOR2 (N7757, N7754, N55);
and AND2 (N7758, N7756, N746);
and AND2 (N7759, N7750, N2123);
not NOT1 (N7760, N7757);
buf BUF1 (N7761, N7755);
nand NAND2 (N7762, N7752, N5099);
buf BUF1 (N7763, N7748);
xor XOR2 (N7764, N7747, N6857);
xor XOR2 (N7765, N7749, N7114);
nor NOR2 (N7766, N7760, N7618);
and AND3 (N7767, N7765, N628, N6897);
not NOT1 (N7768, N7759);
nor NOR4 (N7769, N7764, N4193, N93, N4370);
nor NOR4 (N7770, N7735, N4444, N4016, N1772);
and AND3 (N7771, N7761, N4140, N1285);
not NOT1 (N7772, N7771);
or OR3 (N7773, N7762, N5245, N32);
and AND4 (N7774, N7768, N357, N3504, N4754);
not NOT1 (N7775, N7772);
xor XOR2 (N7776, N7770, N6245);
xor XOR2 (N7777, N7766, N1956);
nand NAND4 (N7778, N7734, N6518, N1163, N3933);
not NOT1 (N7779, N7778);
and AND2 (N7780, N7769, N6039);
and AND2 (N7781, N7777, N2955);
not NOT1 (N7782, N7763);
and AND3 (N7783, N7776, N5899, N6582);
buf BUF1 (N7784, N7780);
or OR2 (N7785, N7775, N1930);
not NOT1 (N7786, N7781);
not NOT1 (N7787, N7785);
nor NOR4 (N7788, N7782, N7688, N6814, N4720);
or OR2 (N7789, N7788, N2935);
nand NAND3 (N7790, N7784, N682, N2052);
or OR3 (N7791, N7774, N4591, N141);
not NOT1 (N7792, N7787);
nand NAND2 (N7793, N7791, N6310);
nand NAND2 (N7794, N7786, N955);
buf BUF1 (N7795, N7792);
and AND2 (N7796, N7794, N6402);
and AND2 (N7797, N7773, N6860);
not NOT1 (N7798, N7796);
not NOT1 (N7799, N7758);
buf BUF1 (N7800, N7799);
nand NAND2 (N7801, N7789, N4681);
xor XOR2 (N7802, N7779, N5446);
buf BUF1 (N7803, N7767);
buf BUF1 (N7804, N7802);
xor XOR2 (N7805, N7797, N7545);
and AND3 (N7806, N7798, N1597, N7045);
xor XOR2 (N7807, N7790, N2553);
not NOT1 (N7808, N7804);
or OR3 (N7809, N7800, N7113, N7319);
buf BUF1 (N7810, N7803);
or OR3 (N7811, N7795, N5114, N3432);
not NOT1 (N7812, N7807);
nor NOR2 (N7813, N7806, N4048);
not NOT1 (N7814, N7811);
and AND2 (N7815, N7814, N2369);
not NOT1 (N7816, N7805);
nor NOR2 (N7817, N7813, N903);
not NOT1 (N7818, N7810);
nor NOR2 (N7819, N7809, N1160);
not NOT1 (N7820, N7812);
or OR4 (N7821, N7820, N4522, N4663, N1681);
buf BUF1 (N7822, N7818);
or OR2 (N7823, N7808, N1514);
nand NAND2 (N7824, N7819, N1484);
xor XOR2 (N7825, N7816, N3833);
xor XOR2 (N7826, N7783, N7769);
or OR2 (N7827, N7822, N1785);
buf BUF1 (N7828, N7821);
and AND2 (N7829, N7815, N701);
xor XOR2 (N7830, N7826, N6378);
nand NAND4 (N7831, N7801, N5328, N903, N930);
nor NOR3 (N7832, N7824, N361, N2406);
nor NOR3 (N7833, N7831, N7782, N3623);
or OR2 (N7834, N7817, N6582);
nand NAND4 (N7835, N7829, N2825, N5889, N2720);
or OR4 (N7836, N7830, N3742, N7162, N6854);
nor NOR3 (N7837, N7836, N4239, N4308);
or OR4 (N7838, N7834, N34, N5339, N4320);
not NOT1 (N7839, N7835);
and AND4 (N7840, N7833, N3561, N6680, N3880);
nor NOR4 (N7841, N7832, N5801, N6131, N4742);
nand NAND2 (N7842, N7837, N4647);
not NOT1 (N7843, N7825);
xor XOR2 (N7844, N7841, N2817);
and AND2 (N7845, N7838, N4182);
xor XOR2 (N7846, N7793, N3252);
buf BUF1 (N7847, N7840);
or OR3 (N7848, N7843, N7679, N1402);
or OR4 (N7849, N7848, N7001, N5586, N6674);
or OR4 (N7850, N7844, N7275, N3545, N7207);
nand NAND4 (N7851, N7842, N3487, N7192, N823);
nand NAND3 (N7852, N7846, N19, N1429);
buf BUF1 (N7853, N7828);
not NOT1 (N7854, N7852);
xor XOR2 (N7855, N7849, N7496);
buf BUF1 (N7856, N7854);
nand NAND2 (N7857, N7827, N6110);
buf BUF1 (N7858, N7839);
and AND3 (N7859, N7823, N3526, N7334);
nand NAND2 (N7860, N7857, N4332);
not NOT1 (N7861, N7856);
nand NAND2 (N7862, N7845, N3412);
nand NAND2 (N7863, N7850, N7551);
nor NOR2 (N7864, N7863, N5469);
xor XOR2 (N7865, N7862, N3090);
and AND2 (N7866, N7858, N6638);
and AND2 (N7867, N7847, N6779);
or OR4 (N7868, N7865, N5571, N1372, N6426);
xor XOR2 (N7869, N7855, N999);
or OR3 (N7870, N7868, N2398, N873);
and AND4 (N7871, N7867, N7485, N7570, N1786);
buf BUF1 (N7872, N7871);
xor XOR2 (N7873, N7853, N5129);
xor XOR2 (N7874, N7866, N4671);
or OR2 (N7875, N7864, N7866);
xor XOR2 (N7876, N7874, N6717);
not NOT1 (N7877, N7861);
not NOT1 (N7878, N7876);
xor XOR2 (N7879, N7859, N4729);
or OR2 (N7880, N7875, N7205);
nand NAND3 (N7881, N7879, N1180, N7154);
nor NOR4 (N7882, N7872, N2354, N3664, N5221);
xor XOR2 (N7883, N7877, N291);
buf BUF1 (N7884, N7880);
not NOT1 (N7885, N7882);
xor XOR2 (N7886, N7860, N6485);
nand NAND2 (N7887, N7869, N6016);
xor XOR2 (N7888, N7851, N7501);
not NOT1 (N7889, N7888);
not NOT1 (N7890, N7887);
not NOT1 (N7891, N7878);
nand NAND4 (N7892, N7883, N6238, N2069, N4784);
xor XOR2 (N7893, N7873, N3086);
or OR4 (N7894, N7889, N5787, N640, N3945);
buf BUF1 (N7895, N7894);
and AND2 (N7896, N7881, N5960);
xor XOR2 (N7897, N7891, N2009);
xor XOR2 (N7898, N7886, N6411);
and AND4 (N7899, N7890, N7694, N5445, N7390);
not NOT1 (N7900, N7898);
and AND4 (N7901, N7900, N1340, N3940, N6934);
not NOT1 (N7902, N7884);
or OR4 (N7903, N7893, N6796, N5314, N1887);
and AND4 (N7904, N7899, N1542, N2241, N6335);
not NOT1 (N7905, N7892);
and AND3 (N7906, N7897, N3754, N5438);
or OR3 (N7907, N7905, N1382, N5672);
nor NOR2 (N7908, N7907, N1212);
xor XOR2 (N7909, N7901, N5687);
not NOT1 (N7910, N7902);
buf BUF1 (N7911, N7885);
not NOT1 (N7912, N7896);
nor NOR3 (N7913, N7895, N7309, N6300);
or OR3 (N7914, N7910, N357, N1107);
xor XOR2 (N7915, N7913, N7877);
buf BUF1 (N7916, N7914);
or OR4 (N7917, N7906, N5462, N7045, N1164);
and AND2 (N7918, N7917, N1240);
or OR2 (N7919, N7916, N3972);
nand NAND4 (N7920, N7915, N4026, N326, N1452);
buf BUF1 (N7921, N7903);
xor XOR2 (N7922, N7904, N1282);
or OR4 (N7923, N7912, N4479, N2603, N2117);
not NOT1 (N7924, N7923);
buf BUF1 (N7925, N7921);
buf BUF1 (N7926, N7925);
buf BUF1 (N7927, N7908);
buf BUF1 (N7928, N7926);
xor XOR2 (N7929, N7920, N5455);
and AND3 (N7930, N7922, N6045, N3213);
or OR3 (N7931, N7930, N3408, N1699);
not NOT1 (N7932, N7928);
nand NAND2 (N7933, N7909, N2897);
and AND3 (N7934, N7931, N3317, N3448);
and AND3 (N7935, N7918, N7155, N4076);
not NOT1 (N7936, N7911);
nand NAND3 (N7937, N7919, N4266, N119);
and AND4 (N7938, N7934, N2089, N5945, N5554);
buf BUF1 (N7939, N7936);
xor XOR2 (N7940, N7935, N7428);
and AND2 (N7941, N7940, N5539);
or OR3 (N7942, N7870, N1138, N5141);
nand NAND3 (N7943, N7942, N6625, N96);
and AND4 (N7944, N7943, N1993, N5700, N2151);
nand NAND2 (N7945, N7937, N814);
nand NAND3 (N7946, N7945, N7608, N7733);
not NOT1 (N7947, N7933);
nor NOR2 (N7948, N7938, N3039);
buf BUF1 (N7949, N7924);
not NOT1 (N7950, N7948);
xor XOR2 (N7951, N7944, N6584);
nand NAND3 (N7952, N7939, N7549, N1611);
nand NAND2 (N7953, N7941, N5070);
nand NAND3 (N7954, N7953, N5997, N7248);
nor NOR2 (N7955, N7954, N7852);
nor NOR3 (N7956, N7955, N3182, N3054);
nand NAND3 (N7957, N7947, N1021, N2449);
xor XOR2 (N7958, N7932, N6406);
or OR4 (N7959, N7950, N1612, N1029, N6182);
xor XOR2 (N7960, N7949, N7596);
nor NOR3 (N7961, N7959, N1192, N6167);
xor XOR2 (N7962, N7952, N5403);
buf BUF1 (N7963, N7958);
nand NAND2 (N7964, N7956, N3174);
or OR2 (N7965, N7929, N3016);
or OR4 (N7966, N7957, N654, N7620, N1578);
and AND3 (N7967, N7927, N7547, N4714);
and AND2 (N7968, N7962, N1831);
xor XOR2 (N7969, N7961, N2255);
and AND3 (N7970, N7966, N228, N5073);
xor XOR2 (N7971, N7970, N4478);
buf BUF1 (N7972, N7965);
xor XOR2 (N7973, N7972, N4425);
buf BUF1 (N7974, N7946);
xor XOR2 (N7975, N7964, N6011);
xor XOR2 (N7976, N7971, N4513);
and AND3 (N7977, N7951, N1734, N6386);
and AND4 (N7978, N7963, N5689, N3166, N7122);
nor NOR2 (N7979, N7973, N1581);
xor XOR2 (N7980, N7968, N939);
nor NOR2 (N7981, N7978, N4699);
nor NOR4 (N7982, N7960, N1738, N2148, N2607);
and AND2 (N7983, N7969, N6978);
buf BUF1 (N7984, N7981);
xor XOR2 (N7985, N7967, N238);
and AND3 (N7986, N7974, N4496, N215);
nand NAND4 (N7987, N7983, N2218, N4724, N4219);
buf BUF1 (N7988, N7986);
xor XOR2 (N7989, N7975, N2805);
xor XOR2 (N7990, N7985, N6160);
buf BUF1 (N7991, N7987);
not NOT1 (N7992, N7977);
nor NOR2 (N7993, N7991, N2843);
and AND4 (N7994, N7976, N2399, N5621, N4374);
not NOT1 (N7995, N7982);
not NOT1 (N7996, N7990);
and AND4 (N7997, N7980, N197, N4790, N492);
xor XOR2 (N7998, N7997, N5236);
xor XOR2 (N7999, N7984, N7771);
nand NAND3 (N8000, N7998, N6653, N1707);
nor NOR3 (N8001, N7995, N5389, N6756);
xor XOR2 (N8002, N8001, N1231);
buf BUF1 (N8003, N8002);
or OR2 (N8004, N8000, N1723);
and AND3 (N8005, N8003, N5032, N1401);
xor XOR2 (N8006, N7979, N5303);
or OR4 (N8007, N7992, N1511, N1084, N6663);
nand NAND2 (N8008, N8007, N6912);
not NOT1 (N8009, N7989);
or OR3 (N8010, N7988, N7534, N1848);
and AND3 (N8011, N7993, N1890, N513);
or OR4 (N8012, N8009, N6405, N5137, N2376);
endmodule