// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16;

output N2989,N3010,N3009,N3002,N2992,N3015,N3011,N3014,N2999,N3016;

nor NOR2 (N17, N8, N16);
buf BUF1 (N18, N17);
and AND2 (N19, N6, N18);
not NOT1 (N20, N13);
nand NAND4 (N21, N20, N12, N10, N18);
and AND3 (N22, N16, N9, N21);
or OR2 (N23, N16, N16);
xor XOR2 (N24, N2, N1);
nand NAND2 (N25, N6, N8);
nand NAND4 (N26, N7, N17, N13, N15);
xor XOR2 (N27, N26, N12);
not NOT1 (N28, N4);
nor NOR2 (N29, N5, N5);
and AND2 (N30, N17, N15);
nor NOR4 (N31, N6, N3, N28, N10);
and AND4 (N32, N3, N1, N10, N13);
or OR2 (N33, N27, N10);
buf BUF1 (N34, N32);
or OR3 (N35, N23, N17, N25);
not NOT1 (N36, N19);
xor XOR2 (N37, N34, N32);
nand NAND4 (N38, N27, N3, N2, N21);
and AND4 (N39, N37, N22, N16, N13);
not NOT1 (N40, N31);
or OR3 (N41, N33, N13, N21);
xor XOR2 (N42, N4, N39);
and AND3 (N43, N32, N39, N2);
and AND4 (N44, N36, N43, N26, N25);
not NOT1 (N45, N9);
or OR4 (N46, N38, N9, N42, N19);
buf BUF1 (N47, N5);
buf BUF1 (N48, N44);
xor XOR2 (N49, N46, N14);
xor XOR2 (N50, N24, N21);
and AND2 (N51, N40, N38);
not NOT1 (N52, N35);
nor NOR3 (N53, N30, N43, N4);
or OR4 (N54, N52, N47, N19, N29);
xor XOR2 (N55, N36, N13);
or OR2 (N56, N5, N47);
nor NOR4 (N57, N41, N34, N36, N4);
and AND2 (N58, N50, N29);
and AND3 (N59, N51, N24, N28);
xor XOR2 (N60, N55, N40);
or OR2 (N61, N48, N47);
not NOT1 (N62, N54);
and AND3 (N63, N60, N11, N19);
and AND2 (N64, N61, N35);
or OR4 (N65, N56, N20, N55, N19);
xor XOR2 (N66, N59, N4);
nor NOR2 (N67, N65, N48);
xor XOR2 (N68, N57, N32);
or OR2 (N69, N66, N7);
nand NAND2 (N70, N62, N48);
nand NAND2 (N71, N64, N42);
nor NOR4 (N72, N70, N3, N23, N55);
and AND2 (N73, N63, N22);
nor NOR2 (N74, N58, N56);
and AND3 (N75, N74, N33, N14);
nor NOR3 (N76, N67, N57, N52);
buf BUF1 (N77, N71);
nand NAND4 (N78, N45, N29, N36, N42);
nand NAND3 (N79, N78, N28, N68);
or OR3 (N80, N76, N65, N39);
or OR3 (N81, N57, N55, N69);
not NOT1 (N82, N20);
or OR3 (N83, N75, N1, N49);
nor NOR2 (N84, N68, N73);
buf BUF1 (N85, N18);
not NOT1 (N86, N83);
nand NAND2 (N87, N77, N3);
nand NAND2 (N88, N80, N60);
xor XOR2 (N89, N81, N61);
and AND2 (N90, N86, N48);
nand NAND4 (N91, N53, N83, N30, N40);
nor NOR2 (N92, N91, N42);
nand NAND2 (N93, N85, N2);
and AND4 (N94, N79, N66, N76, N33);
and AND4 (N95, N92, N4, N29, N90);
or OR3 (N96, N80, N28, N94);
buf BUF1 (N97, N58);
buf BUF1 (N98, N84);
nand NAND2 (N99, N95, N25);
nand NAND2 (N100, N96, N94);
xor XOR2 (N101, N89, N77);
and AND2 (N102, N100, N60);
nor NOR2 (N103, N99, N13);
xor XOR2 (N104, N97, N37);
nor NOR3 (N105, N104, N99, N47);
and AND4 (N106, N93, N74, N33, N71);
nor NOR4 (N107, N106, N48, N3, N11);
not NOT1 (N108, N82);
not NOT1 (N109, N101);
buf BUF1 (N110, N107);
not NOT1 (N111, N72);
nand NAND2 (N112, N88, N93);
or OR2 (N113, N111, N34);
and AND2 (N114, N113, N35);
xor XOR2 (N115, N87, N12);
nand NAND4 (N116, N110, N115, N103, N19);
and AND4 (N117, N71, N32, N5, N41);
xor XOR2 (N118, N71, N55);
not NOT1 (N119, N117);
not NOT1 (N120, N118);
nor NOR3 (N121, N105, N62, N119);
nor NOR2 (N122, N1, N114);
or OR2 (N123, N115, N84);
nand NAND2 (N124, N102, N3);
nand NAND2 (N125, N108, N29);
not NOT1 (N126, N125);
or OR2 (N127, N116, N40);
nor NOR4 (N128, N120, N55, N72, N5);
nor NOR2 (N129, N128, N65);
buf BUF1 (N130, N126);
or OR3 (N131, N130, N69, N67);
or OR3 (N132, N122, N28, N124);
nand NAND4 (N133, N52, N48, N87, N56);
buf BUF1 (N134, N98);
or OR2 (N135, N131, N78);
not NOT1 (N136, N129);
and AND2 (N137, N123, N18);
buf BUF1 (N138, N109);
nor NOR4 (N139, N121, N112, N34, N49);
nor NOR4 (N140, N131, N58, N95, N24);
nor NOR2 (N141, N132, N29);
not NOT1 (N142, N127);
not NOT1 (N143, N133);
xor XOR2 (N144, N141, N25);
nor NOR4 (N145, N135, N58, N113, N102);
and AND3 (N146, N134, N79, N38);
buf BUF1 (N147, N139);
nor NOR2 (N148, N143, N125);
buf BUF1 (N149, N144);
nand NAND4 (N150, N148, N60, N20, N5);
or OR2 (N151, N147, N147);
or OR3 (N152, N150, N14, N126);
xor XOR2 (N153, N140, N23);
buf BUF1 (N154, N146);
buf BUF1 (N155, N151);
or OR2 (N156, N154, N92);
not NOT1 (N157, N153);
or OR3 (N158, N142, N133, N122);
xor XOR2 (N159, N158, N118);
or OR3 (N160, N149, N97, N2);
buf BUF1 (N161, N155);
nand NAND2 (N162, N145, N25);
buf BUF1 (N163, N161);
nor NOR2 (N164, N163, N54);
xor XOR2 (N165, N137, N81);
xor XOR2 (N166, N159, N128);
xor XOR2 (N167, N156, N23);
and AND4 (N168, N160, N137, N52, N88);
not NOT1 (N169, N164);
or OR2 (N170, N166, N75);
or OR3 (N171, N152, N4, N112);
nand NAND2 (N172, N162, N76);
or OR4 (N173, N171, N152, N25, N79);
not NOT1 (N174, N168);
nor NOR3 (N175, N167, N49, N64);
nand NAND2 (N176, N173, N94);
nand NAND2 (N177, N172, N98);
buf BUF1 (N178, N157);
buf BUF1 (N179, N178);
buf BUF1 (N180, N175);
buf BUF1 (N181, N170);
or OR2 (N182, N174, N58);
nor NOR3 (N183, N182, N91, N1);
and AND3 (N184, N180, N58, N148);
or OR2 (N185, N138, N101);
xor XOR2 (N186, N179, N26);
nand NAND3 (N187, N165, N149, N79);
nand NAND3 (N188, N136, N165, N48);
and AND4 (N189, N181, N25, N21, N56);
and AND4 (N190, N185, N49, N77, N57);
nand NAND3 (N191, N189, N5, N129);
and AND2 (N192, N176, N50);
or OR4 (N193, N183, N140, N112, N108);
nand NAND3 (N194, N193, N93, N74);
nand NAND2 (N195, N194, N174);
or OR4 (N196, N188, N84, N70, N163);
nand NAND2 (N197, N186, N104);
nor NOR4 (N198, N177, N193, N147, N121);
or OR4 (N199, N184, N68, N125, N174);
nor NOR3 (N200, N190, N133, N76);
buf BUF1 (N201, N197);
nand NAND3 (N202, N200, N188, N23);
not NOT1 (N203, N192);
xor XOR2 (N204, N202, N65);
and AND4 (N205, N196, N100, N152, N158);
xor XOR2 (N206, N203, N100);
or OR2 (N207, N201, N191);
and AND4 (N208, N12, N44, N26, N36);
not NOT1 (N209, N207);
and AND4 (N210, N169, N84, N110, N103);
nand NAND4 (N211, N206, N170, N162, N164);
nand NAND3 (N212, N205, N118, N76);
xor XOR2 (N213, N204, N20);
xor XOR2 (N214, N212, N8);
and AND3 (N215, N199, N138, N32);
and AND4 (N216, N208, N155, N5, N132);
and AND4 (N217, N198, N20, N87, N60);
and AND3 (N218, N187, N41, N143);
not NOT1 (N219, N195);
xor XOR2 (N220, N218, N149);
nand NAND3 (N221, N211, N189, N206);
nand NAND3 (N222, N209, N27, N52);
buf BUF1 (N223, N215);
not NOT1 (N224, N219);
nand NAND4 (N225, N224, N174, N175, N139);
xor XOR2 (N226, N216, N114);
and AND4 (N227, N222, N8, N178, N89);
nand NAND3 (N228, N220, N162, N212);
and AND2 (N229, N214, N97);
not NOT1 (N230, N229);
nand NAND4 (N231, N225, N205, N224, N197);
and AND4 (N232, N226, N62, N107, N14);
or OR3 (N233, N221, N110, N25);
not NOT1 (N234, N217);
buf BUF1 (N235, N231);
xor XOR2 (N236, N223, N174);
xor XOR2 (N237, N228, N17);
and AND4 (N238, N235, N175, N122, N200);
nand NAND2 (N239, N230, N110);
or OR4 (N240, N234, N58, N62, N65);
nand NAND4 (N241, N227, N226, N188, N231);
or OR3 (N242, N241, N98, N166);
and AND4 (N243, N233, N65, N125, N217);
and AND2 (N244, N213, N80);
xor XOR2 (N245, N244, N17);
and AND4 (N246, N237, N216, N5, N182);
buf BUF1 (N247, N240);
not NOT1 (N248, N210);
and AND2 (N249, N243, N173);
and AND2 (N250, N238, N237);
buf BUF1 (N251, N247);
nor NOR4 (N252, N251, N246, N12, N43);
nand NAND2 (N253, N231, N18);
not NOT1 (N254, N253);
buf BUF1 (N255, N245);
nor NOR4 (N256, N248, N43, N62, N19);
xor XOR2 (N257, N250, N66);
xor XOR2 (N258, N257, N146);
and AND2 (N259, N254, N27);
xor XOR2 (N260, N259, N60);
xor XOR2 (N261, N258, N127);
xor XOR2 (N262, N232, N125);
nand NAND2 (N263, N242, N144);
xor XOR2 (N264, N236, N114);
xor XOR2 (N265, N239, N17);
not NOT1 (N266, N255);
nand NAND4 (N267, N264, N23, N5, N86);
not NOT1 (N268, N263);
and AND3 (N269, N256, N4, N1);
xor XOR2 (N270, N266, N106);
and AND2 (N271, N260, N46);
or OR4 (N272, N267, N141, N111, N113);
nand NAND4 (N273, N261, N71, N159, N31);
not NOT1 (N274, N268);
nor NOR2 (N275, N252, N60);
or OR2 (N276, N269, N61);
nor NOR4 (N277, N249, N267, N58, N102);
xor XOR2 (N278, N265, N47);
buf BUF1 (N279, N272);
xor XOR2 (N280, N273, N199);
or OR2 (N281, N274, N154);
not NOT1 (N282, N280);
nand NAND2 (N283, N275, N42);
xor XOR2 (N284, N282, N146);
not NOT1 (N285, N279);
xor XOR2 (N286, N281, N105);
not NOT1 (N287, N283);
not NOT1 (N288, N287);
buf BUF1 (N289, N277);
not NOT1 (N290, N271);
nor NOR3 (N291, N284, N208, N198);
and AND4 (N292, N276, N32, N12, N246);
buf BUF1 (N293, N291);
nor NOR4 (N294, N293, N188, N25, N231);
nor NOR4 (N295, N286, N249, N203, N208);
nor NOR2 (N296, N262, N213);
nand NAND3 (N297, N289, N59, N48);
or OR4 (N298, N292, N152, N166, N157);
buf BUF1 (N299, N278);
nor NOR2 (N300, N296, N133);
and AND4 (N301, N299, N72, N198, N253);
xor XOR2 (N302, N301, N245);
and AND4 (N303, N295, N260, N171, N37);
and AND3 (N304, N300, N77, N229);
nand NAND4 (N305, N285, N213, N87, N10);
nand NAND3 (N306, N297, N141, N303);
xor XOR2 (N307, N253, N133);
or OR2 (N308, N307, N119);
and AND2 (N309, N288, N275);
not NOT1 (N310, N302);
buf BUF1 (N311, N290);
nand NAND3 (N312, N311, N43, N148);
nor NOR3 (N313, N270, N82, N140);
or OR3 (N314, N313, N60, N126);
and AND4 (N315, N304, N167, N255, N126);
nand NAND2 (N316, N310, N260);
nand NAND4 (N317, N314, N24, N254, N27);
buf BUF1 (N318, N315);
xor XOR2 (N319, N298, N188);
nor NOR3 (N320, N312, N149, N18);
buf BUF1 (N321, N318);
and AND2 (N322, N319, N232);
xor XOR2 (N323, N321, N166);
and AND2 (N324, N317, N54);
or OR4 (N325, N323, N287, N232, N104);
nand NAND3 (N326, N309, N316, N276);
not NOT1 (N327, N62);
xor XOR2 (N328, N325, N129);
nand NAND3 (N329, N305, N260, N84);
or OR2 (N330, N306, N116);
nand NAND4 (N331, N322, N321, N216, N177);
xor XOR2 (N332, N331, N291);
nand NAND3 (N333, N330, N315, N62);
nand NAND3 (N334, N320, N35, N326);
not NOT1 (N335, N50);
buf BUF1 (N336, N332);
or OR4 (N337, N333, N253, N115, N330);
not NOT1 (N338, N336);
and AND2 (N339, N294, N274);
nand NAND2 (N340, N334, N246);
xor XOR2 (N341, N337, N329);
not NOT1 (N342, N35);
buf BUF1 (N343, N308);
or OR3 (N344, N338, N208, N171);
nor NOR2 (N345, N344, N40);
nor NOR4 (N346, N324, N161, N258, N133);
nor NOR3 (N347, N335, N37, N20);
buf BUF1 (N348, N346);
nor NOR4 (N349, N342, N288, N107, N218);
nand NAND4 (N350, N340, N89, N122, N56);
and AND4 (N351, N345, N347, N39, N275);
and AND4 (N352, N314, N137, N241, N350);
or OR4 (N353, N217, N181, N346, N342);
not NOT1 (N354, N349);
not NOT1 (N355, N348);
not NOT1 (N356, N354);
or OR4 (N357, N353, N110, N56, N145);
nor NOR4 (N358, N356, N296, N350, N279);
buf BUF1 (N359, N341);
and AND2 (N360, N351, N340);
nor NOR2 (N361, N358, N109);
buf BUF1 (N362, N361);
xor XOR2 (N363, N360, N268);
or OR2 (N364, N362, N341);
not NOT1 (N365, N359);
xor XOR2 (N366, N328, N217);
nor NOR2 (N367, N357, N97);
buf BUF1 (N368, N339);
nand NAND2 (N369, N367, N363);
or OR2 (N370, N191, N178);
and AND4 (N371, N343, N79, N82, N33);
or OR3 (N372, N366, N180, N340);
nor NOR4 (N373, N352, N252, N145, N309);
buf BUF1 (N374, N373);
buf BUF1 (N375, N374);
buf BUF1 (N376, N355);
not NOT1 (N377, N364);
xor XOR2 (N378, N365, N27);
buf BUF1 (N379, N369);
xor XOR2 (N380, N371, N156);
and AND2 (N381, N327, N142);
or OR4 (N382, N378, N6, N207, N221);
and AND3 (N383, N379, N68, N100);
nand NAND4 (N384, N377, N133, N170, N279);
and AND3 (N385, N370, N77, N342);
or OR4 (N386, N381, N33, N339, N307);
xor XOR2 (N387, N383, N171);
not NOT1 (N388, N384);
buf BUF1 (N389, N368);
and AND3 (N390, N380, N388, N235);
nand NAND2 (N391, N298, N80);
buf BUF1 (N392, N390);
xor XOR2 (N393, N391, N123);
or OR4 (N394, N386, N338, N106, N299);
xor XOR2 (N395, N385, N153);
not NOT1 (N396, N394);
nor NOR4 (N397, N387, N310, N383, N139);
nor NOR2 (N398, N389, N160);
and AND4 (N399, N395, N103, N266, N63);
xor XOR2 (N400, N372, N160);
nand NAND3 (N401, N375, N161, N8);
buf BUF1 (N402, N392);
nand NAND4 (N403, N401, N163, N243, N302);
or OR3 (N404, N382, N244, N95);
nor NOR2 (N405, N400, N372);
nor NOR4 (N406, N403, N151, N198, N355);
nand NAND2 (N407, N396, N172);
and AND4 (N408, N402, N314, N7, N185);
or OR3 (N409, N404, N71, N228);
nor NOR3 (N410, N376, N40, N317);
nand NAND4 (N411, N397, N250, N405, N296);
not NOT1 (N412, N107);
nand NAND3 (N413, N399, N338, N278);
xor XOR2 (N414, N411, N45);
not NOT1 (N415, N412);
or OR3 (N416, N393, N388, N337);
or OR3 (N417, N407, N404, N316);
or OR4 (N418, N408, N205, N92, N50);
buf BUF1 (N419, N398);
not NOT1 (N420, N406);
and AND3 (N421, N416, N12, N337);
not NOT1 (N422, N421);
xor XOR2 (N423, N410, N26);
xor XOR2 (N424, N420, N91);
and AND2 (N425, N424, N247);
buf BUF1 (N426, N409);
or OR3 (N427, N417, N301, N210);
buf BUF1 (N428, N414);
and AND2 (N429, N425, N177);
and AND2 (N430, N419, N269);
or OR2 (N431, N423, N339);
buf BUF1 (N432, N426);
nand NAND4 (N433, N428, N62, N118, N390);
nand NAND4 (N434, N429, N201, N61, N256);
and AND3 (N435, N433, N202, N261);
xor XOR2 (N436, N422, N395);
not NOT1 (N437, N434);
not NOT1 (N438, N427);
xor XOR2 (N439, N431, N298);
or OR3 (N440, N438, N212, N411);
nand NAND2 (N441, N440, N353);
or OR3 (N442, N430, N101, N72);
or OR3 (N443, N439, N298, N204);
and AND3 (N444, N413, N109, N164);
and AND4 (N445, N435, N371, N350, N318);
or OR4 (N446, N415, N201, N18, N368);
or OR3 (N447, N446, N11, N346);
nand NAND2 (N448, N444, N68);
xor XOR2 (N449, N418, N222);
and AND3 (N450, N436, N153, N449);
or OR2 (N451, N101, N42);
not NOT1 (N452, N432);
nand NAND2 (N453, N450, N66);
nand NAND2 (N454, N445, N259);
nor NOR3 (N455, N443, N86, N274);
and AND4 (N456, N447, N36, N392, N338);
and AND4 (N457, N448, N350, N150, N82);
or OR3 (N458, N451, N225, N430);
or OR4 (N459, N441, N104, N7, N103);
not NOT1 (N460, N459);
not NOT1 (N461, N458);
and AND2 (N462, N437, N314);
nor NOR4 (N463, N461, N399, N329, N442);
or OR3 (N464, N390, N209, N34);
and AND3 (N465, N454, N220, N408);
nand NAND3 (N466, N460, N225, N351);
or OR3 (N467, N463, N283, N37);
and AND3 (N468, N464, N244, N367);
not NOT1 (N469, N467);
and AND2 (N470, N453, N184);
buf BUF1 (N471, N470);
nor NOR2 (N472, N468, N35);
xor XOR2 (N473, N469, N361);
buf BUF1 (N474, N462);
and AND3 (N475, N457, N46, N429);
and AND3 (N476, N466, N206, N232);
buf BUF1 (N477, N465);
nor NOR3 (N478, N472, N352, N386);
nand NAND4 (N479, N452, N168, N471, N436);
nand NAND2 (N480, N90, N425);
buf BUF1 (N481, N476);
nor NOR4 (N482, N475, N178, N65, N251);
and AND3 (N483, N481, N292, N291);
xor XOR2 (N484, N474, N310);
or OR3 (N485, N479, N401, N157);
not NOT1 (N486, N478);
or OR4 (N487, N455, N57, N197, N149);
xor XOR2 (N488, N477, N139);
buf BUF1 (N489, N485);
buf BUF1 (N490, N473);
or OR3 (N491, N482, N42, N288);
or OR4 (N492, N486, N197, N367, N160);
buf BUF1 (N493, N484);
xor XOR2 (N494, N456, N420);
and AND3 (N495, N488, N263, N213);
and AND2 (N496, N489, N337);
nor NOR4 (N497, N483, N234, N74, N319);
and AND2 (N498, N496, N25);
nor NOR4 (N499, N497, N471, N109, N239);
and AND2 (N500, N480, N294);
buf BUF1 (N501, N495);
nor NOR3 (N502, N492, N460, N464);
and AND2 (N503, N501, N200);
and AND4 (N504, N499, N477, N61, N164);
and AND2 (N505, N502, N33);
or OR2 (N506, N505, N408);
nand NAND3 (N507, N494, N57, N306);
xor XOR2 (N508, N504, N445);
or OR2 (N509, N507, N366);
and AND2 (N510, N509, N94);
and AND2 (N511, N500, N328);
or OR2 (N512, N511, N427);
or OR3 (N513, N490, N10, N108);
and AND4 (N514, N513, N100, N67, N256);
buf BUF1 (N515, N498);
xor XOR2 (N516, N491, N495);
buf BUF1 (N517, N487);
nand NAND4 (N518, N514, N378, N228, N313);
and AND3 (N519, N506, N189, N51);
nor NOR2 (N520, N510, N155);
or OR3 (N521, N508, N433, N516);
or OR3 (N522, N1, N381, N166);
and AND3 (N523, N503, N56, N211);
xor XOR2 (N524, N521, N445);
xor XOR2 (N525, N493, N378);
nand NAND2 (N526, N523, N260);
xor XOR2 (N527, N522, N455);
xor XOR2 (N528, N525, N379);
nand NAND2 (N529, N518, N322);
nand NAND4 (N530, N527, N357, N107, N254);
nand NAND2 (N531, N524, N82);
nor NOR3 (N532, N517, N330, N94);
buf BUF1 (N533, N528);
buf BUF1 (N534, N512);
and AND3 (N535, N533, N392, N352);
and AND3 (N536, N530, N530, N259);
nand NAND3 (N537, N531, N147, N399);
not NOT1 (N538, N519);
xor XOR2 (N539, N536, N196);
xor XOR2 (N540, N529, N55);
buf BUF1 (N541, N535);
nand NAND4 (N542, N520, N235, N381, N325);
nand NAND2 (N543, N537, N174);
or OR3 (N544, N540, N314, N215);
nor NOR3 (N545, N544, N182, N528);
or OR2 (N546, N515, N7);
or OR4 (N547, N538, N418, N375, N443);
xor XOR2 (N548, N546, N392);
nor NOR4 (N549, N545, N453, N416, N128);
or OR4 (N550, N547, N259, N40, N128);
buf BUF1 (N551, N526);
nand NAND4 (N552, N548, N38, N458, N6);
nand NAND3 (N553, N543, N117, N155);
nor NOR2 (N554, N553, N513);
buf BUF1 (N555, N541);
xor XOR2 (N556, N542, N179);
not NOT1 (N557, N549);
and AND4 (N558, N557, N502, N320, N156);
or OR4 (N559, N532, N463, N97, N118);
nor NOR2 (N560, N558, N326);
or OR4 (N561, N554, N229, N260, N32);
and AND4 (N562, N552, N174, N352, N523);
nand NAND4 (N563, N556, N510, N142, N547);
xor XOR2 (N564, N551, N478);
buf BUF1 (N565, N534);
nor NOR3 (N566, N555, N100, N524);
buf BUF1 (N567, N539);
not NOT1 (N568, N561);
buf BUF1 (N569, N559);
buf BUF1 (N570, N550);
xor XOR2 (N571, N564, N428);
nand NAND3 (N572, N560, N552, N235);
and AND2 (N573, N568, N285);
not NOT1 (N574, N566);
and AND4 (N575, N570, N417, N197, N532);
nand NAND4 (N576, N572, N306, N187, N254);
buf BUF1 (N577, N576);
nand NAND3 (N578, N574, N161, N172);
nor NOR4 (N579, N571, N203, N258, N280);
and AND3 (N580, N577, N4, N321);
not NOT1 (N581, N565);
or OR4 (N582, N581, N439, N423, N278);
nor NOR3 (N583, N562, N305, N16);
xor XOR2 (N584, N578, N467);
or OR3 (N585, N575, N140, N193);
or OR3 (N586, N579, N186, N68);
buf BUF1 (N587, N573);
not NOT1 (N588, N587);
and AND4 (N589, N585, N394, N583, N481);
and AND4 (N590, N566, N167, N107, N352);
xor XOR2 (N591, N590, N139);
and AND4 (N592, N563, N32, N24, N88);
or OR3 (N593, N567, N364, N312);
nand NAND4 (N594, N591, N297, N54, N63);
buf BUF1 (N595, N592);
not NOT1 (N596, N589);
nand NAND2 (N597, N580, N22);
nand NAND2 (N598, N586, N350);
or OR3 (N599, N569, N88, N158);
or OR4 (N600, N582, N319, N382, N226);
buf BUF1 (N601, N596);
and AND2 (N602, N597, N297);
not NOT1 (N603, N600);
and AND2 (N604, N598, N599);
nor NOR2 (N605, N434, N174);
or OR2 (N606, N588, N265);
or OR2 (N607, N603, N346);
not NOT1 (N608, N604);
xor XOR2 (N609, N584, N570);
xor XOR2 (N610, N601, N258);
nor NOR2 (N611, N609, N241);
and AND4 (N612, N607, N325, N420, N180);
and AND3 (N613, N608, N9, N244);
xor XOR2 (N614, N595, N196);
not NOT1 (N615, N611);
not NOT1 (N616, N606);
not NOT1 (N617, N605);
buf BUF1 (N618, N614);
or OR3 (N619, N617, N322, N201);
nand NAND3 (N620, N602, N28, N6);
xor XOR2 (N621, N620, N77);
buf BUF1 (N622, N613);
nand NAND2 (N623, N593, N54);
xor XOR2 (N624, N618, N359);
not NOT1 (N625, N619);
xor XOR2 (N626, N612, N535);
or OR3 (N627, N594, N358, N426);
nor NOR2 (N628, N610, N125);
nand NAND4 (N629, N621, N191, N510, N108);
xor XOR2 (N630, N627, N471);
or OR4 (N631, N615, N523, N262, N112);
and AND4 (N632, N628, N18, N586, N145);
and AND3 (N633, N632, N435, N480);
not NOT1 (N634, N625);
not NOT1 (N635, N629);
nor NOR3 (N636, N616, N120, N608);
or OR3 (N637, N630, N185, N263);
or OR3 (N638, N634, N493, N441);
buf BUF1 (N639, N638);
nor NOR4 (N640, N624, N464, N562, N272);
xor XOR2 (N641, N636, N348);
buf BUF1 (N642, N635);
nand NAND2 (N643, N623, N552);
nor NOR2 (N644, N631, N82);
or OR2 (N645, N644, N129);
xor XOR2 (N646, N633, N603);
nand NAND3 (N647, N642, N61, N417);
and AND4 (N648, N639, N534, N377, N405);
xor XOR2 (N649, N626, N167);
xor XOR2 (N650, N640, N350);
not NOT1 (N651, N643);
buf BUF1 (N652, N622);
xor XOR2 (N653, N645, N56);
xor XOR2 (N654, N646, N41);
nor NOR2 (N655, N652, N373);
or OR2 (N656, N655, N513);
or OR3 (N657, N637, N441, N363);
nand NAND3 (N658, N656, N221, N632);
and AND4 (N659, N651, N525, N144, N444);
and AND2 (N660, N654, N88);
nor NOR4 (N661, N653, N440, N296, N327);
not NOT1 (N662, N648);
buf BUF1 (N663, N658);
nor NOR4 (N664, N641, N119, N389, N153);
or OR4 (N665, N647, N260, N264, N287);
or OR3 (N666, N659, N332, N15);
xor XOR2 (N667, N664, N398);
not NOT1 (N668, N662);
and AND3 (N669, N660, N567, N371);
not NOT1 (N670, N661);
not NOT1 (N671, N670);
or OR2 (N672, N650, N57);
xor XOR2 (N673, N668, N589);
or OR3 (N674, N669, N578, N244);
and AND3 (N675, N674, N267, N650);
xor XOR2 (N676, N649, N347);
nor NOR4 (N677, N667, N38, N275, N347);
and AND3 (N678, N665, N589, N625);
buf BUF1 (N679, N673);
not NOT1 (N680, N675);
buf BUF1 (N681, N676);
nor NOR2 (N682, N672, N321);
buf BUF1 (N683, N657);
or OR2 (N684, N682, N609);
nand NAND2 (N685, N680, N260);
nor NOR4 (N686, N677, N58, N660, N661);
or OR4 (N687, N686, N183, N357, N69);
not NOT1 (N688, N687);
buf BUF1 (N689, N684);
or OR4 (N690, N678, N367, N126, N237);
xor XOR2 (N691, N671, N244);
nand NAND2 (N692, N679, N596);
and AND3 (N693, N685, N252, N74);
nor NOR2 (N694, N663, N623);
nand NAND2 (N695, N683, N320);
nor NOR3 (N696, N666, N223, N456);
xor XOR2 (N697, N690, N568);
and AND2 (N698, N694, N624);
xor XOR2 (N699, N698, N479);
nor NOR3 (N700, N689, N191, N3);
xor XOR2 (N701, N697, N512);
or OR4 (N702, N695, N230, N420, N184);
nand NAND3 (N703, N688, N613, N578);
nor NOR4 (N704, N692, N228, N669, N110);
not NOT1 (N705, N704);
and AND3 (N706, N681, N173, N484);
buf BUF1 (N707, N706);
xor XOR2 (N708, N700, N635);
buf BUF1 (N709, N699);
buf BUF1 (N710, N702);
or OR4 (N711, N705, N456, N687, N417);
and AND2 (N712, N693, N551);
xor XOR2 (N713, N691, N424);
nand NAND2 (N714, N710, N127);
or OR2 (N715, N707, N658);
or OR3 (N716, N712, N588, N557);
and AND3 (N717, N714, N158, N159);
not NOT1 (N718, N703);
or OR4 (N719, N711, N276, N686, N671);
and AND4 (N720, N701, N6, N455, N182);
xor XOR2 (N721, N718, N195);
xor XOR2 (N722, N719, N378);
and AND2 (N723, N713, N47);
or OR4 (N724, N715, N715, N93, N21);
nand NAND3 (N725, N716, N547, N82);
xor XOR2 (N726, N721, N410);
nor NOR3 (N727, N724, N540, N218);
and AND3 (N728, N717, N621, N706);
nor NOR2 (N729, N722, N724);
nand NAND4 (N730, N708, N686, N602, N121);
buf BUF1 (N731, N723);
not NOT1 (N732, N696);
xor XOR2 (N733, N729, N658);
or OR4 (N734, N726, N233, N439, N156);
nand NAND2 (N735, N725, N180);
buf BUF1 (N736, N720);
xor XOR2 (N737, N734, N694);
nand NAND3 (N738, N727, N527, N408);
and AND2 (N739, N732, N515);
nand NAND4 (N740, N709, N726, N554, N262);
xor XOR2 (N741, N739, N347);
buf BUF1 (N742, N731);
or OR2 (N743, N742, N486);
nor NOR3 (N744, N738, N206, N264);
nand NAND2 (N745, N744, N294);
buf BUF1 (N746, N728);
or OR3 (N747, N743, N737, N46);
nor NOR4 (N748, N649, N124, N659, N206);
nor NOR3 (N749, N740, N559, N78);
nand NAND2 (N750, N746, N148);
xor XOR2 (N751, N733, N736);
or OR3 (N752, N520, N518, N36);
nand NAND4 (N753, N730, N719, N294, N642);
not NOT1 (N754, N747);
buf BUF1 (N755, N745);
not NOT1 (N756, N752);
xor XOR2 (N757, N756, N132);
buf BUF1 (N758, N751);
nor NOR3 (N759, N750, N402, N420);
nor NOR4 (N760, N748, N471, N199, N457);
buf BUF1 (N761, N735);
or OR3 (N762, N759, N567, N338);
buf BUF1 (N763, N762);
and AND3 (N764, N749, N395, N566);
not NOT1 (N765, N760);
buf BUF1 (N766, N758);
and AND4 (N767, N763, N149, N275, N161);
nand NAND4 (N768, N765, N452, N419, N378);
nor NOR4 (N769, N741, N355, N36, N223);
or OR4 (N770, N757, N690, N440, N202);
buf BUF1 (N771, N753);
or OR2 (N772, N754, N478);
xor XOR2 (N773, N768, N591);
xor XOR2 (N774, N761, N130);
nor NOR3 (N775, N772, N497, N18);
nor NOR2 (N776, N755, N446);
xor XOR2 (N777, N770, N81);
buf BUF1 (N778, N767);
not NOT1 (N779, N769);
not NOT1 (N780, N779);
and AND2 (N781, N775, N167);
nor NOR3 (N782, N764, N529, N423);
not NOT1 (N783, N776);
xor XOR2 (N784, N781, N247);
and AND4 (N785, N782, N151, N583, N178);
nand NAND2 (N786, N780, N742);
xor XOR2 (N787, N783, N734);
nand NAND4 (N788, N786, N390, N196, N673);
nand NAND2 (N789, N778, N229);
not NOT1 (N790, N774);
not NOT1 (N791, N790);
buf BUF1 (N792, N789);
not NOT1 (N793, N785);
not NOT1 (N794, N766);
nor NOR4 (N795, N784, N642, N514, N184);
and AND4 (N796, N793, N28, N644, N201);
xor XOR2 (N797, N788, N152);
nor NOR3 (N798, N795, N313, N319);
xor XOR2 (N799, N787, N659);
buf BUF1 (N800, N777);
nor NOR4 (N801, N799, N666, N602, N525);
nor NOR2 (N802, N797, N327);
buf BUF1 (N803, N800);
nand NAND3 (N804, N773, N732, N404);
nor NOR3 (N805, N792, N707, N392);
nand NAND3 (N806, N791, N552, N497);
nor NOR2 (N807, N803, N536);
not NOT1 (N808, N804);
not NOT1 (N809, N806);
or OR4 (N810, N807, N516, N540, N214);
and AND3 (N811, N810, N90, N155);
not NOT1 (N812, N796);
buf BUF1 (N813, N801);
or OR4 (N814, N809, N2, N521, N82);
xor XOR2 (N815, N798, N440);
and AND2 (N816, N771, N462);
nand NAND4 (N817, N815, N316, N205, N190);
and AND2 (N818, N805, N252);
xor XOR2 (N819, N816, N91);
xor XOR2 (N820, N814, N671);
xor XOR2 (N821, N819, N413);
not NOT1 (N822, N812);
buf BUF1 (N823, N811);
xor XOR2 (N824, N820, N761);
buf BUF1 (N825, N824);
or OR3 (N826, N822, N254, N121);
buf BUF1 (N827, N808);
buf BUF1 (N828, N813);
nor NOR4 (N829, N821, N747, N139, N575);
and AND2 (N830, N802, N449);
buf BUF1 (N831, N817);
not NOT1 (N832, N827);
not NOT1 (N833, N831);
buf BUF1 (N834, N818);
and AND4 (N835, N833, N681, N804, N610);
nor NOR3 (N836, N829, N459, N376);
nand NAND4 (N837, N794, N247, N468, N689);
and AND2 (N838, N825, N468);
buf BUF1 (N839, N834);
or OR2 (N840, N837, N264);
nor NOR4 (N841, N838, N224, N52, N369);
nand NAND2 (N842, N841, N309);
nor NOR3 (N843, N830, N539, N353);
not NOT1 (N844, N839);
not NOT1 (N845, N842);
and AND2 (N846, N845, N817);
or OR3 (N847, N835, N742, N442);
or OR4 (N848, N840, N612, N153, N811);
buf BUF1 (N849, N826);
not NOT1 (N850, N846);
nor NOR4 (N851, N832, N265, N793, N704);
nor NOR4 (N852, N849, N122, N712, N713);
nor NOR4 (N853, N850, N836, N54, N756);
nand NAND4 (N854, N27, N644, N513, N239);
nor NOR3 (N855, N853, N310, N817);
or OR2 (N856, N823, N53);
xor XOR2 (N857, N851, N358);
nand NAND4 (N858, N847, N715, N434, N767);
xor XOR2 (N859, N852, N473);
or OR2 (N860, N843, N688);
buf BUF1 (N861, N844);
nor NOR4 (N862, N848, N24, N34, N606);
nor NOR2 (N863, N855, N404);
nand NAND4 (N864, N854, N650, N434, N58);
or OR2 (N865, N856, N183);
or OR2 (N866, N862, N69);
buf BUF1 (N867, N859);
nand NAND2 (N868, N864, N774);
or OR2 (N869, N863, N400);
and AND2 (N870, N828, N263);
buf BUF1 (N871, N869);
xor XOR2 (N872, N868, N643);
not NOT1 (N873, N861);
nand NAND2 (N874, N857, N95);
buf BUF1 (N875, N866);
or OR3 (N876, N867, N627, N333);
nor NOR2 (N877, N875, N562);
nor NOR2 (N878, N870, N371);
nand NAND3 (N879, N873, N770, N405);
nor NOR2 (N880, N858, N9);
buf BUF1 (N881, N880);
not NOT1 (N882, N872);
and AND4 (N883, N878, N788, N382, N718);
and AND4 (N884, N871, N778, N408, N44);
or OR4 (N885, N879, N248, N267, N72);
not NOT1 (N886, N865);
xor XOR2 (N887, N884, N815);
not NOT1 (N888, N874);
nand NAND3 (N889, N877, N870, N6);
not NOT1 (N890, N876);
or OR3 (N891, N860, N685, N406);
buf BUF1 (N892, N891);
nor NOR3 (N893, N883, N581, N780);
nand NAND4 (N894, N881, N742, N36, N806);
buf BUF1 (N895, N888);
or OR2 (N896, N886, N159);
or OR4 (N897, N885, N477, N829, N36);
nor NOR3 (N898, N887, N69, N391);
not NOT1 (N899, N894);
and AND4 (N900, N882, N833, N152, N780);
nor NOR2 (N901, N896, N646);
nand NAND4 (N902, N898, N457, N450, N621);
or OR4 (N903, N897, N466, N306, N3);
buf BUF1 (N904, N902);
xor XOR2 (N905, N890, N857);
xor XOR2 (N906, N893, N164);
and AND2 (N907, N900, N425);
nand NAND4 (N908, N905, N129, N863, N141);
xor XOR2 (N909, N903, N794);
not NOT1 (N910, N895);
and AND2 (N911, N910, N681);
xor XOR2 (N912, N892, N812);
and AND4 (N913, N901, N72, N890, N136);
or OR3 (N914, N907, N672, N590);
or OR3 (N915, N909, N464, N78);
nor NOR2 (N916, N904, N873);
and AND4 (N917, N916, N808, N511, N839);
nand NAND3 (N918, N908, N193, N537);
nor NOR2 (N919, N906, N9);
or OR4 (N920, N919, N795, N460, N129);
not NOT1 (N921, N912);
nand NAND2 (N922, N899, N711);
nand NAND3 (N923, N921, N46, N130);
buf BUF1 (N924, N889);
xor XOR2 (N925, N924, N74);
and AND2 (N926, N914, N744);
not NOT1 (N927, N923);
nand NAND2 (N928, N915, N780);
and AND3 (N929, N918, N883, N262);
buf BUF1 (N930, N922);
and AND4 (N931, N930, N752, N601, N127);
nand NAND2 (N932, N928, N707);
nand NAND4 (N933, N925, N113, N443, N599);
nor NOR2 (N934, N911, N548);
nor NOR4 (N935, N913, N170, N417, N904);
not NOT1 (N936, N933);
xor XOR2 (N937, N929, N207);
or OR3 (N938, N936, N724, N889);
nor NOR2 (N939, N934, N120);
nand NAND4 (N940, N937, N395, N643, N675);
buf BUF1 (N941, N935);
or OR3 (N942, N920, N149, N828);
and AND4 (N943, N917, N498, N343, N579);
nand NAND2 (N944, N941, N490);
xor XOR2 (N945, N938, N414);
xor XOR2 (N946, N931, N834);
and AND3 (N947, N932, N494, N214);
and AND3 (N948, N947, N486, N801);
not NOT1 (N949, N948);
and AND4 (N950, N949, N530, N776, N179);
and AND2 (N951, N927, N772);
buf BUF1 (N952, N945);
xor XOR2 (N953, N944, N775);
buf BUF1 (N954, N946);
xor XOR2 (N955, N950, N415);
nor NOR2 (N956, N943, N320);
and AND2 (N957, N926, N559);
xor XOR2 (N958, N942, N364);
xor XOR2 (N959, N951, N302);
buf BUF1 (N960, N959);
nand NAND2 (N961, N957, N467);
buf BUF1 (N962, N953);
or OR4 (N963, N954, N689, N424, N239);
buf BUF1 (N964, N952);
nor NOR4 (N965, N939, N74, N393, N524);
not NOT1 (N966, N961);
not NOT1 (N967, N964);
not NOT1 (N968, N940);
xor XOR2 (N969, N965, N897);
nand NAND4 (N970, N963, N45, N305, N272);
or OR2 (N971, N969, N778);
not NOT1 (N972, N968);
nand NAND4 (N973, N958, N90, N212, N545);
buf BUF1 (N974, N960);
not NOT1 (N975, N962);
nor NOR2 (N976, N975, N431);
and AND4 (N977, N956, N127, N103, N149);
and AND2 (N978, N977, N919);
nor NOR4 (N979, N973, N241, N925, N215);
nand NAND4 (N980, N970, N81, N551, N23);
nand NAND4 (N981, N974, N448, N255, N871);
buf BUF1 (N982, N955);
buf BUF1 (N983, N981);
nand NAND3 (N984, N983, N193, N316);
nand NAND2 (N985, N982, N586);
nor NOR3 (N986, N984, N25, N21);
and AND4 (N987, N986, N952, N879, N753);
xor XOR2 (N988, N972, N787);
xor XOR2 (N989, N966, N504);
or OR4 (N990, N979, N138, N195, N223);
nor NOR3 (N991, N967, N723, N777);
nor NOR3 (N992, N989, N507, N608);
nor NOR3 (N993, N987, N587, N456);
not NOT1 (N994, N971);
nor NOR3 (N995, N992, N173, N947);
nand NAND2 (N996, N991, N104);
or OR4 (N997, N993, N743, N836, N801);
nand NAND2 (N998, N997, N537);
nand NAND4 (N999, N988, N172, N339, N190);
buf BUF1 (N1000, N980);
and AND2 (N1001, N999, N589);
buf BUF1 (N1002, N996);
xor XOR2 (N1003, N1000, N466);
xor XOR2 (N1004, N990, N451);
buf BUF1 (N1005, N1004);
and AND2 (N1006, N976, N34);
or OR4 (N1007, N1005, N254, N363, N684);
nor NOR3 (N1008, N1006, N755, N192);
not NOT1 (N1009, N1002);
and AND4 (N1010, N1008, N448, N4, N305);
nor NOR3 (N1011, N995, N367, N165);
nor NOR3 (N1012, N985, N379, N756);
buf BUF1 (N1013, N978);
buf BUF1 (N1014, N1001);
xor XOR2 (N1015, N1003, N508);
xor XOR2 (N1016, N998, N522);
not NOT1 (N1017, N1015);
buf BUF1 (N1018, N1009);
xor XOR2 (N1019, N1007, N6);
nor NOR3 (N1020, N1010, N740, N743);
buf BUF1 (N1021, N1020);
and AND3 (N1022, N1018, N425, N438);
not NOT1 (N1023, N1016);
xor XOR2 (N1024, N1013, N997);
buf BUF1 (N1025, N1017);
buf BUF1 (N1026, N1023);
and AND3 (N1027, N994, N719, N42);
nor NOR4 (N1028, N1024, N323, N221, N652);
not NOT1 (N1029, N1027);
buf BUF1 (N1030, N1025);
not NOT1 (N1031, N1022);
buf BUF1 (N1032, N1028);
xor XOR2 (N1033, N1030, N3);
nand NAND4 (N1034, N1029, N412, N526, N950);
not NOT1 (N1035, N1034);
nand NAND4 (N1036, N1012, N304, N304, N753);
and AND3 (N1037, N1033, N967, N593);
xor XOR2 (N1038, N1036, N552);
nor NOR2 (N1039, N1032, N159);
nor NOR4 (N1040, N1037, N306, N148, N798);
buf BUF1 (N1041, N1040);
nand NAND3 (N1042, N1011, N478, N276);
nor NOR2 (N1043, N1026, N905);
nand NAND4 (N1044, N1031, N449, N508, N808);
not NOT1 (N1045, N1019);
xor XOR2 (N1046, N1043, N652);
nand NAND4 (N1047, N1045, N921, N433, N75);
buf BUF1 (N1048, N1021);
nor NOR4 (N1049, N1041, N517, N440, N673);
buf BUF1 (N1050, N1039);
buf BUF1 (N1051, N1049);
and AND3 (N1052, N1051, N760, N606);
buf BUF1 (N1053, N1047);
and AND2 (N1054, N1050, N679);
or OR4 (N1055, N1035, N1015, N84, N591);
or OR4 (N1056, N1044, N750, N401, N362);
not NOT1 (N1057, N1014);
nand NAND2 (N1058, N1056, N510);
and AND3 (N1059, N1052, N113, N946);
nor NOR3 (N1060, N1058, N339, N585);
nand NAND4 (N1061, N1054, N909, N476, N93);
xor XOR2 (N1062, N1046, N917);
nand NAND3 (N1063, N1055, N660, N823);
and AND2 (N1064, N1048, N948);
xor XOR2 (N1065, N1042, N136);
or OR4 (N1066, N1038, N651, N681, N671);
nor NOR3 (N1067, N1066, N22, N859);
xor XOR2 (N1068, N1062, N1008);
or OR2 (N1069, N1059, N656);
buf BUF1 (N1070, N1063);
buf BUF1 (N1071, N1053);
and AND4 (N1072, N1065, N936, N1069, N501);
or OR4 (N1073, N877, N277, N590, N911);
or OR3 (N1074, N1057, N380, N332);
xor XOR2 (N1075, N1073, N443);
and AND4 (N1076, N1068, N888, N451, N988);
not NOT1 (N1077, N1067);
nor NOR4 (N1078, N1074, N970, N28, N435);
and AND2 (N1079, N1070, N700);
and AND3 (N1080, N1076, N166, N509);
or OR3 (N1081, N1077, N161, N220);
and AND2 (N1082, N1078, N144);
and AND3 (N1083, N1079, N297, N728);
xor XOR2 (N1084, N1083, N171);
or OR3 (N1085, N1064, N539, N769);
and AND2 (N1086, N1084, N573);
nor NOR3 (N1087, N1085, N41, N946);
buf BUF1 (N1088, N1071);
nor NOR2 (N1089, N1086, N137);
and AND4 (N1090, N1082, N543, N1010, N951);
buf BUF1 (N1091, N1060);
buf BUF1 (N1092, N1075);
nand NAND4 (N1093, N1090, N284, N877, N824);
nor NOR2 (N1094, N1088, N818);
or OR2 (N1095, N1072, N1035);
nand NAND4 (N1096, N1061, N904, N957, N740);
nand NAND3 (N1097, N1080, N783, N340);
buf BUF1 (N1098, N1089);
xor XOR2 (N1099, N1092, N837);
nand NAND2 (N1100, N1081, N417);
or OR4 (N1101, N1096, N1093, N52, N635);
buf BUF1 (N1102, N964);
xor XOR2 (N1103, N1102, N960);
nor NOR3 (N1104, N1100, N132, N214);
nor NOR4 (N1105, N1097, N408, N647, N691);
buf BUF1 (N1106, N1098);
nand NAND2 (N1107, N1099, N998);
buf BUF1 (N1108, N1104);
or OR3 (N1109, N1094, N103, N517);
or OR3 (N1110, N1087, N197, N119);
and AND3 (N1111, N1107, N1099, N362);
xor XOR2 (N1112, N1101, N590);
and AND2 (N1113, N1106, N688);
nor NOR3 (N1114, N1110, N261, N368);
nand NAND2 (N1115, N1111, N942);
and AND2 (N1116, N1105, N889);
and AND3 (N1117, N1109, N998, N895);
or OR3 (N1118, N1103, N291, N235);
and AND3 (N1119, N1108, N876, N1075);
nor NOR3 (N1120, N1117, N849, N802);
nor NOR2 (N1121, N1112, N951);
not NOT1 (N1122, N1116);
buf BUF1 (N1123, N1119);
buf BUF1 (N1124, N1122);
xor XOR2 (N1125, N1120, N16);
or OR4 (N1126, N1091, N944, N59, N231);
nor NOR4 (N1127, N1118, N1057, N535, N908);
nand NAND3 (N1128, N1124, N2, N246);
xor XOR2 (N1129, N1126, N843);
and AND3 (N1130, N1121, N690, N618);
nor NOR3 (N1131, N1127, N648, N978);
nor NOR2 (N1132, N1129, N848);
nor NOR4 (N1133, N1095, N830, N366, N1003);
or OR4 (N1134, N1114, N26, N659, N793);
xor XOR2 (N1135, N1131, N423);
buf BUF1 (N1136, N1123);
or OR2 (N1137, N1134, N601);
buf BUF1 (N1138, N1115);
buf BUF1 (N1139, N1128);
buf BUF1 (N1140, N1135);
not NOT1 (N1141, N1132);
nor NOR4 (N1142, N1113, N595, N1058, N499);
nor NOR4 (N1143, N1141, N791, N789, N235);
and AND3 (N1144, N1133, N709, N795);
nor NOR4 (N1145, N1125, N767, N544, N1100);
nand NAND2 (N1146, N1138, N773);
not NOT1 (N1147, N1130);
or OR2 (N1148, N1136, N95);
nand NAND2 (N1149, N1147, N243);
nand NAND3 (N1150, N1144, N935, N532);
nor NOR4 (N1151, N1140, N730, N963, N1134);
and AND2 (N1152, N1145, N654);
or OR2 (N1153, N1149, N38);
buf BUF1 (N1154, N1142);
and AND4 (N1155, N1146, N613, N275, N772);
buf BUF1 (N1156, N1153);
buf BUF1 (N1157, N1139);
xor XOR2 (N1158, N1151, N349);
or OR2 (N1159, N1155, N196);
not NOT1 (N1160, N1158);
buf BUF1 (N1161, N1152);
not NOT1 (N1162, N1161);
and AND2 (N1163, N1156, N213);
or OR2 (N1164, N1163, N911);
nor NOR2 (N1165, N1157, N65);
xor XOR2 (N1166, N1148, N205);
or OR2 (N1167, N1159, N506);
nor NOR2 (N1168, N1166, N1017);
nor NOR2 (N1169, N1143, N645);
xor XOR2 (N1170, N1168, N437);
and AND3 (N1171, N1167, N281, N1063);
xor XOR2 (N1172, N1170, N221);
and AND4 (N1173, N1137, N339, N15, N731);
xor XOR2 (N1174, N1169, N778);
not NOT1 (N1175, N1165);
and AND2 (N1176, N1160, N477);
buf BUF1 (N1177, N1154);
or OR4 (N1178, N1164, N523, N403, N1131);
nand NAND3 (N1179, N1175, N248, N954);
buf BUF1 (N1180, N1179);
or OR3 (N1181, N1178, N911, N912);
xor XOR2 (N1182, N1177, N43);
nand NAND2 (N1183, N1174, N1090);
nor NOR4 (N1184, N1172, N139, N820, N100);
buf BUF1 (N1185, N1171);
nand NAND4 (N1186, N1181, N731, N584, N210);
buf BUF1 (N1187, N1184);
xor XOR2 (N1188, N1185, N1051);
nor NOR3 (N1189, N1186, N459, N823);
buf BUF1 (N1190, N1173);
xor XOR2 (N1191, N1189, N482);
xor XOR2 (N1192, N1187, N742);
or OR4 (N1193, N1180, N1161, N318, N59);
xor XOR2 (N1194, N1188, N1185);
xor XOR2 (N1195, N1162, N293);
or OR2 (N1196, N1182, N626);
and AND2 (N1197, N1192, N727);
not NOT1 (N1198, N1190);
not NOT1 (N1199, N1195);
nand NAND4 (N1200, N1197, N782, N820, N1102);
and AND2 (N1201, N1200, N947);
or OR3 (N1202, N1176, N129, N1179);
not NOT1 (N1203, N1194);
nand NAND3 (N1204, N1202, N964, N1023);
not NOT1 (N1205, N1150);
and AND2 (N1206, N1204, N808);
buf BUF1 (N1207, N1196);
buf BUF1 (N1208, N1207);
buf BUF1 (N1209, N1193);
not NOT1 (N1210, N1183);
nand NAND3 (N1211, N1201, N732, N304);
buf BUF1 (N1212, N1203);
xor XOR2 (N1213, N1211, N227);
and AND4 (N1214, N1205, N846, N448, N1070);
and AND3 (N1215, N1208, N844, N109);
nor NOR3 (N1216, N1215, N206, N1008);
nand NAND2 (N1217, N1213, N1164);
xor XOR2 (N1218, N1216, N532);
nor NOR4 (N1219, N1212, N64, N150, N1065);
not NOT1 (N1220, N1191);
nand NAND3 (N1221, N1198, N43, N766);
nand NAND2 (N1222, N1214, N711);
not NOT1 (N1223, N1199);
buf BUF1 (N1224, N1218);
xor XOR2 (N1225, N1219, N693);
or OR3 (N1226, N1206, N483, N356);
buf BUF1 (N1227, N1217);
buf BUF1 (N1228, N1220);
not NOT1 (N1229, N1221);
or OR4 (N1230, N1222, N212, N838, N54);
nor NOR4 (N1231, N1230, N822, N262, N406);
nand NAND2 (N1232, N1229, N628);
nor NOR3 (N1233, N1232, N501, N688);
xor XOR2 (N1234, N1226, N849);
xor XOR2 (N1235, N1209, N703);
buf BUF1 (N1236, N1235);
not NOT1 (N1237, N1233);
xor XOR2 (N1238, N1231, N1095);
not NOT1 (N1239, N1223);
or OR4 (N1240, N1239, N651, N603, N476);
xor XOR2 (N1241, N1234, N776);
buf BUF1 (N1242, N1236);
nor NOR4 (N1243, N1228, N552, N169, N696);
and AND4 (N1244, N1224, N682, N154, N812);
and AND4 (N1245, N1238, N22, N387, N1115);
xor XOR2 (N1246, N1245, N187);
xor XOR2 (N1247, N1242, N360);
buf BUF1 (N1248, N1246);
or OR2 (N1249, N1225, N422);
or OR4 (N1250, N1244, N709, N848, N708);
xor XOR2 (N1251, N1249, N57);
and AND2 (N1252, N1241, N564);
and AND4 (N1253, N1243, N149, N473, N785);
and AND2 (N1254, N1250, N1049);
and AND3 (N1255, N1252, N1029, N497);
or OR2 (N1256, N1254, N929);
nand NAND3 (N1257, N1248, N167, N133);
buf BUF1 (N1258, N1247);
not NOT1 (N1259, N1227);
xor XOR2 (N1260, N1257, N927);
buf BUF1 (N1261, N1255);
xor XOR2 (N1262, N1256, N828);
not NOT1 (N1263, N1251);
not NOT1 (N1264, N1259);
and AND2 (N1265, N1262, N1262);
nand NAND4 (N1266, N1237, N502, N1170, N1210);
not NOT1 (N1267, N89);
nor NOR2 (N1268, N1264, N577);
xor XOR2 (N1269, N1258, N28);
nand NAND3 (N1270, N1268, N631, N890);
xor XOR2 (N1271, N1269, N1124);
not NOT1 (N1272, N1266);
nand NAND3 (N1273, N1265, N1154, N451);
nor NOR2 (N1274, N1240, N215);
buf BUF1 (N1275, N1253);
and AND2 (N1276, N1267, N902);
buf BUF1 (N1277, N1272);
or OR3 (N1278, N1276, N559, N815);
nor NOR3 (N1279, N1275, N367, N353);
nor NOR2 (N1280, N1277, N455);
or OR2 (N1281, N1273, N105);
nand NAND3 (N1282, N1271, N309, N817);
buf BUF1 (N1283, N1263);
nor NOR4 (N1284, N1260, N529, N235, N1072);
nand NAND4 (N1285, N1280, N730, N244, N1156);
nand NAND3 (N1286, N1284, N6, N880);
and AND2 (N1287, N1270, N245);
not NOT1 (N1288, N1287);
not NOT1 (N1289, N1282);
or OR2 (N1290, N1278, N640);
buf BUF1 (N1291, N1290);
xor XOR2 (N1292, N1285, N604);
not NOT1 (N1293, N1289);
not NOT1 (N1294, N1291);
nand NAND2 (N1295, N1261, N118);
or OR2 (N1296, N1286, N383);
not NOT1 (N1297, N1296);
not NOT1 (N1298, N1297);
or OR3 (N1299, N1288, N938, N705);
and AND3 (N1300, N1293, N616, N67);
and AND3 (N1301, N1292, N548, N1094);
not NOT1 (N1302, N1274);
not NOT1 (N1303, N1299);
not NOT1 (N1304, N1301);
and AND2 (N1305, N1300, N103);
and AND2 (N1306, N1283, N1246);
or OR2 (N1307, N1306, N689);
and AND4 (N1308, N1295, N619, N11, N539);
buf BUF1 (N1309, N1298);
and AND2 (N1310, N1303, N1271);
xor XOR2 (N1311, N1304, N653);
nand NAND4 (N1312, N1294, N484, N276, N1151);
buf BUF1 (N1313, N1305);
nor NOR3 (N1314, N1281, N946, N929);
buf BUF1 (N1315, N1308);
or OR3 (N1316, N1314, N376, N337);
nor NOR2 (N1317, N1312, N1120);
and AND2 (N1318, N1309, N824);
nor NOR2 (N1319, N1310, N598);
nor NOR2 (N1320, N1316, N673);
and AND3 (N1321, N1319, N102, N471);
not NOT1 (N1322, N1279);
not NOT1 (N1323, N1315);
or OR2 (N1324, N1323, N773);
nor NOR4 (N1325, N1322, N901, N343, N67);
xor XOR2 (N1326, N1321, N748);
buf BUF1 (N1327, N1318);
nor NOR3 (N1328, N1327, N55, N1063);
nor NOR3 (N1329, N1326, N1140, N739);
and AND3 (N1330, N1313, N269, N672);
nand NAND3 (N1331, N1311, N350, N860);
buf BUF1 (N1332, N1307);
nand NAND4 (N1333, N1328, N1006, N435, N979);
and AND4 (N1334, N1332, N1045, N814, N818);
and AND2 (N1335, N1320, N276);
not NOT1 (N1336, N1302);
nand NAND2 (N1337, N1324, N361);
and AND4 (N1338, N1334, N1232, N100, N1309);
or OR3 (N1339, N1335, N231, N447);
nor NOR4 (N1340, N1325, N73, N969, N1114);
nor NOR3 (N1341, N1338, N92, N515);
not NOT1 (N1342, N1317);
and AND3 (N1343, N1340, N145, N1061);
nand NAND2 (N1344, N1339, N488);
xor XOR2 (N1345, N1329, N1031);
nor NOR2 (N1346, N1343, N674);
and AND2 (N1347, N1345, N78);
and AND3 (N1348, N1336, N492, N333);
and AND3 (N1349, N1344, N741, N928);
buf BUF1 (N1350, N1347);
or OR4 (N1351, N1337, N365, N1052, N862);
nor NOR3 (N1352, N1333, N545, N1034);
nand NAND2 (N1353, N1342, N750);
buf BUF1 (N1354, N1351);
and AND4 (N1355, N1330, N729, N1187, N1122);
not NOT1 (N1356, N1353);
and AND3 (N1357, N1356, N32, N478);
nor NOR3 (N1358, N1348, N866, N1226);
nor NOR2 (N1359, N1346, N1168);
xor XOR2 (N1360, N1350, N1032);
and AND3 (N1361, N1354, N776, N1143);
or OR3 (N1362, N1349, N1292, N704);
buf BUF1 (N1363, N1355);
nand NAND3 (N1364, N1361, N168, N1022);
and AND4 (N1365, N1352, N102, N1144, N191);
nor NOR3 (N1366, N1364, N424, N1238);
xor XOR2 (N1367, N1359, N712);
not NOT1 (N1368, N1358);
nand NAND2 (N1369, N1368, N158);
nor NOR3 (N1370, N1362, N785, N804);
nor NOR4 (N1371, N1366, N699, N823, N280);
nor NOR4 (N1372, N1369, N12, N405, N1275);
nand NAND3 (N1373, N1331, N1084, N64);
buf BUF1 (N1374, N1372);
nor NOR2 (N1375, N1373, N1138);
not NOT1 (N1376, N1341);
xor XOR2 (N1377, N1376, N839);
nand NAND2 (N1378, N1374, N964);
buf BUF1 (N1379, N1363);
xor XOR2 (N1380, N1367, N301);
not NOT1 (N1381, N1365);
nor NOR3 (N1382, N1370, N1343, N1295);
buf BUF1 (N1383, N1357);
buf BUF1 (N1384, N1378);
and AND3 (N1385, N1380, N885, N657);
and AND4 (N1386, N1383, N321, N1275, N122);
and AND3 (N1387, N1371, N978, N291);
or OR4 (N1388, N1377, N1198, N350, N1052);
buf BUF1 (N1389, N1384);
nor NOR3 (N1390, N1381, N749, N334);
and AND3 (N1391, N1379, N139, N1255);
nor NOR3 (N1392, N1390, N118, N994);
xor XOR2 (N1393, N1391, N1178);
or OR2 (N1394, N1392, N429);
nand NAND3 (N1395, N1394, N302, N757);
nor NOR4 (N1396, N1386, N711, N578, N1288);
xor XOR2 (N1397, N1393, N886);
not NOT1 (N1398, N1388);
nor NOR4 (N1399, N1360, N923, N1067, N62);
or OR4 (N1400, N1387, N40, N614, N450);
and AND2 (N1401, N1385, N849);
or OR3 (N1402, N1400, N541, N479);
buf BUF1 (N1403, N1402);
or OR4 (N1404, N1399, N454, N1134, N428);
nand NAND3 (N1405, N1397, N489, N789);
nor NOR4 (N1406, N1396, N474, N757, N299);
nor NOR3 (N1407, N1389, N662, N1087);
not NOT1 (N1408, N1398);
nor NOR3 (N1409, N1382, N877, N268);
not NOT1 (N1410, N1375);
buf BUF1 (N1411, N1405);
and AND2 (N1412, N1401, N320);
and AND3 (N1413, N1410, N1038, N475);
not NOT1 (N1414, N1411);
nor NOR2 (N1415, N1414, N1276);
nand NAND2 (N1416, N1407, N662);
nand NAND2 (N1417, N1415, N770);
nand NAND2 (N1418, N1413, N399);
nand NAND2 (N1419, N1416, N147);
nand NAND3 (N1420, N1403, N1176, N1047);
buf BUF1 (N1421, N1409);
nor NOR4 (N1422, N1395, N1306, N655, N858);
and AND2 (N1423, N1419, N990);
or OR3 (N1424, N1408, N624, N1126);
nand NAND4 (N1425, N1422, N817, N42, N670);
or OR3 (N1426, N1412, N77, N1380);
not NOT1 (N1427, N1426);
or OR4 (N1428, N1417, N1081, N447, N791);
or OR3 (N1429, N1404, N1393, N1185);
not NOT1 (N1430, N1420);
buf BUF1 (N1431, N1421);
nand NAND4 (N1432, N1425, N1294, N656, N731);
nand NAND2 (N1433, N1423, N1244);
not NOT1 (N1434, N1424);
nor NOR2 (N1435, N1418, N33);
buf BUF1 (N1436, N1429);
buf BUF1 (N1437, N1431);
or OR4 (N1438, N1434, N782, N855, N684);
xor XOR2 (N1439, N1406, N1032);
xor XOR2 (N1440, N1432, N372);
buf BUF1 (N1441, N1440);
nand NAND2 (N1442, N1441, N951);
and AND2 (N1443, N1430, N886);
and AND2 (N1444, N1435, N918);
xor XOR2 (N1445, N1428, N210);
xor XOR2 (N1446, N1427, N464);
and AND4 (N1447, N1437, N243, N701, N171);
xor XOR2 (N1448, N1445, N645);
not NOT1 (N1449, N1443);
xor XOR2 (N1450, N1444, N685);
or OR2 (N1451, N1436, N1360);
or OR3 (N1452, N1451, N1035, N52);
and AND3 (N1453, N1452, N1243, N878);
and AND3 (N1454, N1453, N771, N1064);
not NOT1 (N1455, N1454);
not NOT1 (N1456, N1447);
nand NAND4 (N1457, N1456, N311, N322, N445);
xor XOR2 (N1458, N1442, N239);
or OR4 (N1459, N1449, N68, N624, N1237);
nor NOR2 (N1460, N1438, N575);
buf BUF1 (N1461, N1446);
buf BUF1 (N1462, N1457);
or OR3 (N1463, N1460, N755, N131);
or OR4 (N1464, N1433, N1297, N299, N757);
buf BUF1 (N1465, N1463);
buf BUF1 (N1466, N1465);
nand NAND4 (N1467, N1464, N649, N447, N1074);
and AND3 (N1468, N1467, N118, N827);
xor XOR2 (N1469, N1458, N1453);
nor NOR2 (N1470, N1466, N1366);
or OR2 (N1471, N1462, N679);
and AND2 (N1472, N1469, N864);
nand NAND3 (N1473, N1472, N503, N203);
and AND2 (N1474, N1461, N1129);
nand NAND4 (N1475, N1470, N539, N595, N1043);
or OR4 (N1476, N1473, N257, N848, N1351);
xor XOR2 (N1477, N1455, N378);
nand NAND4 (N1478, N1459, N1236, N413, N298);
buf BUF1 (N1479, N1477);
not NOT1 (N1480, N1448);
buf BUF1 (N1481, N1476);
xor XOR2 (N1482, N1481, N576);
not NOT1 (N1483, N1482);
nand NAND3 (N1484, N1480, N1148, N1291);
nor NOR2 (N1485, N1471, N138);
not NOT1 (N1486, N1484);
and AND2 (N1487, N1485, N443);
not NOT1 (N1488, N1487);
nand NAND2 (N1489, N1478, N585);
or OR3 (N1490, N1479, N53, N691);
nor NOR2 (N1491, N1468, N1389);
not NOT1 (N1492, N1474);
nor NOR2 (N1493, N1475, N35);
and AND3 (N1494, N1483, N1083, N977);
nor NOR3 (N1495, N1493, N266, N1078);
buf BUF1 (N1496, N1495);
nand NAND2 (N1497, N1492, N500);
not NOT1 (N1498, N1497);
or OR3 (N1499, N1450, N56, N59);
nand NAND4 (N1500, N1488, N299, N852, N1288);
not NOT1 (N1501, N1499);
nand NAND4 (N1502, N1486, N1191, N1119, N958);
nand NAND3 (N1503, N1496, N1281, N605);
and AND2 (N1504, N1502, N197);
nand NAND4 (N1505, N1500, N555, N667, N102);
xor XOR2 (N1506, N1505, N817);
buf BUF1 (N1507, N1491);
not NOT1 (N1508, N1501);
nor NOR2 (N1509, N1494, N1288);
xor XOR2 (N1510, N1506, N937);
xor XOR2 (N1511, N1490, N652);
buf BUF1 (N1512, N1504);
nor NOR3 (N1513, N1439, N503, N101);
and AND2 (N1514, N1489, N1362);
buf BUF1 (N1515, N1514);
xor XOR2 (N1516, N1512, N1067);
xor XOR2 (N1517, N1508, N170);
buf BUF1 (N1518, N1516);
buf BUF1 (N1519, N1511);
xor XOR2 (N1520, N1517, N476);
or OR3 (N1521, N1498, N329, N882);
and AND2 (N1522, N1507, N355);
xor XOR2 (N1523, N1522, N844);
xor XOR2 (N1524, N1521, N1106);
or OR2 (N1525, N1524, N1222);
xor XOR2 (N1526, N1515, N117);
buf BUF1 (N1527, N1503);
nor NOR3 (N1528, N1510, N952, N570);
buf BUF1 (N1529, N1527);
nor NOR4 (N1530, N1509, N1144, N1210, N170);
and AND3 (N1531, N1529, N351, N297);
not NOT1 (N1532, N1531);
xor XOR2 (N1533, N1523, N468);
buf BUF1 (N1534, N1519);
nor NOR2 (N1535, N1530, N691);
not NOT1 (N1536, N1513);
or OR4 (N1537, N1534, N1376, N898, N693);
not NOT1 (N1538, N1536);
nor NOR2 (N1539, N1528, N1411);
nand NAND2 (N1540, N1537, N794);
not NOT1 (N1541, N1532);
nand NAND3 (N1542, N1518, N36, N1388);
not NOT1 (N1543, N1540);
not NOT1 (N1544, N1535);
and AND3 (N1545, N1526, N1256, N1329);
nor NOR3 (N1546, N1543, N585, N170);
nand NAND4 (N1547, N1542, N1391, N85, N1212);
or OR2 (N1548, N1547, N968);
buf BUF1 (N1549, N1525);
or OR3 (N1550, N1541, N648, N94);
buf BUF1 (N1551, N1549);
nor NOR2 (N1552, N1544, N183);
nor NOR3 (N1553, N1548, N960, N1471);
nand NAND3 (N1554, N1539, N875, N90);
xor XOR2 (N1555, N1520, N771);
nand NAND2 (N1556, N1550, N890);
nor NOR3 (N1557, N1553, N1213, N1240);
or OR4 (N1558, N1545, N220, N335, N712);
xor XOR2 (N1559, N1555, N1347);
buf BUF1 (N1560, N1552);
or OR2 (N1561, N1538, N176);
nand NAND3 (N1562, N1559, N958, N272);
buf BUF1 (N1563, N1558);
not NOT1 (N1564, N1560);
and AND4 (N1565, N1561, N1364, N972, N1167);
xor XOR2 (N1566, N1557, N498);
not NOT1 (N1567, N1556);
nand NAND4 (N1568, N1563, N265, N949, N1096);
xor XOR2 (N1569, N1564, N470);
nand NAND2 (N1570, N1554, N1412);
nand NAND4 (N1571, N1551, N1397, N964, N1427);
buf BUF1 (N1572, N1566);
not NOT1 (N1573, N1568);
nor NOR3 (N1574, N1533, N620, N1467);
xor XOR2 (N1575, N1570, N1313);
or OR2 (N1576, N1562, N1356);
and AND2 (N1577, N1575, N160);
or OR4 (N1578, N1576, N569, N446, N565);
nand NAND4 (N1579, N1572, N886, N213, N1526);
and AND2 (N1580, N1577, N151);
xor XOR2 (N1581, N1546, N946);
xor XOR2 (N1582, N1565, N44);
nor NOR4 (N1583, N1581, N1239, N1561, N293);
nor NOR3 (N1584, N1578, N917, N130);
and AND4 (N1585, N1579, N265, N863, N275);
and AND4 (N1586, N1569, N662, N1368, N1321);
buf BUF1 (N1587, N1586);
or OR2 (N1588, N1582, N1099);
not NOT1 (N1589, N1580);
buf BUF1 (N1590, N1573);
not NOT1 (N1591, N1583);
not NOT1 (N1592, N1589);
or OR3 (N1593, N1585, N1505, N1106);
and AND4 (N1594, N1571, N448, N1314, N744);
not NOT1 (N1595, N1591);
nand NAND3 (N1596, N1574, N1584, N240);
nor NOR3 (N1597, N898, N424, N1288);
or OR3 (N1598, N1597, N1569, N398);
nand NAND3 (N1599, N1587, N936, N550);
nand NAND3 (N1600, N1567, N868, N1100);
buf BUF1 (N1601, N1600);
and AND2 (N1602, N1590, N31);
buf BUF1 (N1603, N1595);
xor XOR2 (N1604, N1603, N106);
nor NOR2 (N1605, N1593, N1533);
not NOT1 (N1606, N1594);
buf BUF1 (N1607, N1602);
or OR3 (N1608, N1605, N479, N869);
nor NOR3 (N1609, N1608, N196, N1071);
nand NAND2 (N1610, N1609, N609);
nor NOR4 (N1611, N1592, N1188, N1078, N1582);
not NOT1 (N1612, N1610);
nand NAND2 (N1613, N1599, N328);
buf BUF1 (N1614, N1612);
not NOT1 (N1615, N1588);
xor XOR2 (N1616, N1607, N118);
nand NAND4 (N1617, N1615, N1505, N486, N774);
xor XOR2 (N1618, N1613, N790);
or OR4 (N1619, N1604, N1398, N1390, N386);
and AND4 (N1620, N1596, N472, N1538, N194);
not NOT1 (N1621, N1616);
and AND2 (N1622, N1598, N213);
xor XOR2 (N1623, N1617, N687);
buf BUF1 (N1624, N1606);
or OR4 (N1625, N1622, N75, N540, N24);
nand NAND2 (N1626, N1623, N813);
nand NAND4 (N1627, N1624, N148, N1129, N127);
xor XOR2 (N1628, N1620, N1004);
nand NAND3 (N1629, N1627, N849, N1322);
not NOT1 (N1630, N1618);
buf BUF1 (N1631, N1625);
xor XOR2 (N1632, N1628, N1168);
xor XOR2 (N1633, N1611, N70);
xor XOR2 (N1634, N1630, N449);
xor XOR2 (N1635, N1631, N1254);
or OR2 (N1636, N1621, N155);
buf BUF1 (N1637, N1632);
or OR3 (N1638, N1636, N786, N88);
nor NOR3 (N1639, N1634, N927, N1603);
or OR2 (N1640, N1635, N1443);
or OR4 (N1641, N1601, N1447, N817, N1281);
buf BUF1 (N1642, N1626);
buf BUF1 (N1643, N1639);
nor NOR2 (N1644, N1619, N1414);
and AND4 (N1645, N1614, N1190, N527, N2);
buf BUF1 (N1646, N1645);
not NOT1 (N1647, N1629);
and AND2 (N1648, N1642, N504);
nor NOR2 (N1649, N1647, N1460);
xor XOR2 (N1650, N1648, N186);
nand NAND3 (N1651, N1638, N688, N848);
nand NAND2 (N1652, N1633, N976);
nand NAND4 (N1653, N1650, N717, N1083, N1206);
or OR2 (N1654, N1640, N766);
not NOT1 (N1655, N1652);
and AND2 (N1656, N1641, N774);
buf BUF1 (N1657, N1643);
and AND3 (N1658, N1657, N177, N962);
buf BUF1 (N1659, N1654);
not NOT1 (N1660, N1658);
buf BUF1 (N1661, N1656);
not NOT1 (N1662, N1644);
nor NOR2 (N1663, N1661, N939);
or OR3 (N1664, N1662, N521, N1039);
not NOT1 (N1665, N1664);
and AND2 (N1666, N1653, N62);
nor NOR3 (N1667, N1665, N1132, N1468);
nor NOR2 (N1668, N1651, N1466);
and AND4 (N1669, N1649, N2, N265, N784);
or OR3 (N1670, N1663, N1119, N980);
nand NAND3 (N1671, N1655, N675, N521);
not NOT1 (N1672, N1668);
xor XOR2 (N1673, N1669, N699);
xor XOR2 (N1674, N1637, N1408);
nand NAND3 (N1675, N1646, N72, N750);
and AND3 (N1676, N1660, N796, N717);
buf BUF1 (N1677, N1675);
and AND2 (N1678, N1672, N1206);
nor NOR3 (N1679, N1673, N939, N1249);
and AND2 (N1680, N1666, N595);
and AND4 (N1681, N1674, N1671, N1389, N485);
xor XOR2 (N1682, N14, N328);
not NOT1 (N1683, N1659);
xor XOR2 (N1684, N1670, N566);
nor NOR2 (N1685, N1678, N979);
buf BUF1 (N1686, N1685);
not NOT1 (N1687, N1677);
not NOT1 (N1688, N1676);
nor NOR3 (N1689, N1687, N1243, N288);
xor XOR2 (N1690, N1680, N767);
or OR2 (N1691, N1688, N916);
nor NOR2 (N1692, N1686, N938);
or OR2 (N1693, N1692, N156);
or OR2 (N1694, N1682, N448);
buf BUF1 (N1695, N1679);
or OR4 (N1696, N1689, N225, N1341, N1404);
nand NAND3 (N1697, N1684, N711, N7);
nand NAND3 (N1698, N1693, N1625, N462);
and AND3 (N1699, N1681, N849, N1368);
or OR4 (N1700, N1683, N230, N676, N157);
or OR3 (N1701, N1694, N1386, N965);
and AND3 (N1702, N1690, N1612, N832);
or OR3 (N1703, N1699, N867, N1124);
and AND3 (N1704, N1701, N876, N1078);
buf BUF1 (N1705, N1704);
nand NAND3 (N1706, N1703, N476, N1397);
buf BUF1 (N1707, N1700);
or OR3 (N1708, N1705, N1500, N355);
nand NAND2 (N1709, N1698, N661);
nand NAND4 (N1710, N1708, N734, N387, N1112);
or OR4 (N1711, N1695, N874, N1618, N1027);
buf BUF1 (N1712, N1691);
and AND2 (N1713, N1707, N1242);
xor XOR2 (N1714, N1710, N120);
or OR3 (N1715, N1706, N677, N1555);
nor NOR2 (N1716, N1697, N721);
or OR3 (N1717, N1709, N953, N163);
and AND2 (N1718, N1716, N1594);
or OR2 (N1719, N1712, N81);
nor NOR2 (N1720, N1667, N949);
nor NOR3 (N1721, N1696, N1505, N657);
buf BUF1 (N1722, N1714);
or OR3 (N1723, N1702, N869, N538);
nand NAND2 (N1724, N1717, N997);
buf BUF1 (N1725, N1713);
nand NAND4 (N1726, N1722, N1638, N815, N1158);
not NOT1 (N1727, N1726);
and AND2 (N1728, N1721, N1650);
or OR2 (N1729, N1727, N357);
buf BUF1 (N1730, N1724);
and AND4 (N1731, N1720, N1395, N1240, N1032);
nand NAND3 (N1732, N1718, N344, N1038);
and AND2 (N1733, N1728, N250);
and AND4 (N1734, N1725, N1690, N786, N1654);
nor NOR2 (N1735, N1711, N593);
nor NOR2 (N1736, N1730, N869);
and AND2 (N1737, N1719, N332);
nor NOR2 (N1738, N1734, N1581);
nor NOR4 (N1739, N1737, N1502, N458, N1439);
not NOT1 (N1740, N1723);
not NOT1 (N1741, N1735);
or OR2 (N1742, N1729, N1110);
buf BUF1 (N1743, N1738);
not NOT1 (N1744, N1732);
nor NOR4 (N1745, N1743, N633, N904, N111);
and AND2 (N1746, N1744, N921);
nor NOR3 (N1747, N1745, N575, N797);
nand NAND3 (N1748, N1742, N91, N144);
buf BUF1 (N1749, N1747);
buf BUF1 (N1750, N1739);
or OR3 (N1751, N1748, N1392, N1082);
nand NAND3 (N1752, N1750, N495, N1257);
and AND3 (N1753, N1746, N1263, N515);
not NOT1 (N1754, N1752);
nor NOR3 (N1755, N1731, N903, N1285);
nand NAND2 (N1756, N1751, N154);
or OR4 (N1757, N1736, N1481, N430, N89);
buf BUF1 (N1758, N1740);
nor NOR2 (N1759, N1715, N520);
or OR3 (N1760, N1741, N646, N194);
buf BUF1 (N1761, N1756);
or OR3 (N1762, N1757, N1096, N1028);
buf BUF1 (N1763, N1733);
nand NAND2 (N1764, N1758, N293);
nor NOR2 (N1765, N1753, N1008);
nand NAND3 (N1766, N1749, N612, N211);
nor NOR2 (N1767, N1764, N85);
buf BUF1 (N1768, N1754);
or OR2 (N1769, N1759, N1014);
or OR3 (N1770, N1762, N1338, N909);
xor XOR2 (N1771, N1761, N994);
not NOT1 (N1772, N1771);
nor NOR4 (N1773, N1767, N1072, N1069, N467);
or OR4 (N1774, N1765, N912, N1328, N1322);
nand NAND2 (N1775, N1768, N1360);
buf BUF1 (N1776, N1760);
nand NAND2 (N1777, N1770, N361);
nand NAND4 (N1778, N1777, N1039, N898, N675);
nor NOR2 (N1779, N1776, N392);
not NOT1 (N1780, N1774);
nor NOR2 (N1781, N1769, N513);
nand NAND3 (N1782, N1773, N348, N724);
nor NOR3 (N1783, N1772, N1631, N1001);
not NOT1 (N1784, N1780);
not NOT1 (N1785, N1781);
nor NOR3 (N1786, N1782, N687, N74);
buf BUF1 (N1787, N1785);
or OR2 (N1788, N1766, N781);
and AND4 (N1789, N1783, N926, N1221, N291);
nand NAND4 (N1790, N1779, N261, N74, N665);
nand NAND4 (N1791, N1790, N1451, N1258, N703);
not NOT1 (N1792, N1787);
buf BUF1 (N1793, N1786);
xor XOR2 (N1794, N1775, N810);
not NOT1 (N1795, N1794);
and AND4 (N1796, N1788, N155, N1710, N1578);
not NOT1 (N1797, N1795);
nor NOR3 (N1798, N1778, N1304, N1678);
not NOT1 (N1799, N1798);
nor NOR2 (N1800, N1797, N362);
buf BUF1 (N1801, N1792);
or OR2 (N1802, N1755, N1185);
buf BUF1 (N1803, N1802);
xor XOR2 (N1804, N1796, N832);
not NOT1 (N1805, N1800);
not NOT1 (N1806, N1763);
nand NAND3 (N1807, N1784, N1563, N1371);
not NOT1 (N1808, N1793);
and AND2 (N1809, N1806, N892);
or OR4 (N1810, N1789, N1236, N662, N659);
or OR2 (N1811, N1808, N163);
buf BUF1 (N1812, N1811);
and AND3 (N1813, N1804, N874, N523);
nand NAND3 (N1814, N1791, N1694, N284);
not NOT1 (N1815, N1812);
nor NOR4 (N1816, N1810, N1235, N628, N887);
xor XOR2 (N1817, N1809, N327);
nor NOR2 (N1818, N1813, N464);
nand NAND3 (N1819, N1803, N1406, N1177);
or OR3 (N1820, N1819, N1563, N692);
xor XOR2 (N1821, N1816, N34);
nor NOR3 (N1822, N1820, N94, N807);
and AND2 (N1823, N1801, N629);
nor NOR2 (N1824, N1799, N1431);
not NOT1 (N1825, N1817);
buf BUF1 (N1826, N1822);
buf BUF1 (N1827, N1807);
nand NAND3 (N1828, N1818, N420, N322);
not NOT1 (N1829, N1827);
nor NOR2 (N1830, N1814, N1140);
buf BUF1 (N1831, N1824);
and AND3 (N1832, N1826, N1170, N807);
and AND2 (N1833, N1828, N398);
or OR2 (N1834, N1821, N877);
nor NOR4 (N1835, N1825, N1108, N1197, N1123);
not NOT1 (N1836, N1833);
not NOT1 (N1837, N1835);
xor XOR2 (N1838, N1829, N1033);
nand NAND2 (N1839, N1815, N1118);
not NOT1 (N1840, N1832);
and AND2 (N1841, N1831, N990);
buf BUF1 (N1842, N1839);
or OR3 (N1843, N1840, N352, N1589);
nor NOR4 (N1844, N1836, N1667, N501, N889);
and AND3 (N1845, N1844, N1011, N282);
buf BUF1 (N1846, N1830);
xor XOR2 (N1847, N1842, N1351);
xor XOR2 (N1848, N1805, N513);
and AND2 (N1849, N1848, N89);
and AND3 (N1850, N1841, N1574, N119);
and AND4 (N1851, N1837, N12, N291, N1027);
or OR4 (N1852, N1823, N1045, N1092, N18);
or OR2 (N1853, N1851, N1153);
or OR3 (N1854, N1847, N1523, N1546);
not NOT1 (N1855, N1853);
xor XOR2 (N1856, N1852, N73);
buf BUF1 (N1857, N1849);
nand NAND3 (N1858, N1846, N318, N807);
or OR3 (N1859, N1854, N377, N581);
buf BUF1 (N1860, N1858);
nand NAND4 (N1861, N1834, N987, N69, N42);
buf BUF1 (N1862, N1856);
buf BUF1 (N1863, N1855);
or OR4 (N1864, N1862, N715, N989, N723);
and AND3 (N1865, N1845, N1258, N1678);
or OR4 (N1866, N1860, N1345, N1098, N370);
and AND2 (N1867, N1857, N1262);
xor XOR2 (N1868, N1861, N268);
buf BUF1 (N1869, N1866);
nand NAND2 (N1870, N1868, N601);
and AND3 (N1871, N1869, N1424, N1099);
buf BUF1 (N1872, N1864);
xor XOR2 (N1873, N1870, N1057);
nor NOR2 (N1874, N1850, N359);
and AND3 (N1875, N1867, N515, N1684);
not NOT1 (N1876, N1871);
nand NAND4 (N1877, N1865, N1836, N1545, N1125);
nor NOR2 (N1878, N1859, N1573);
xor XOR2 (N1879, N1838, N866);
nor NOR3 (N1880, N1877, N1866, N1042);
nand NAND3 (N1881, N1872, N1348, N250);
nor NOR2 (N1882, N1878, N1300);
and AND4 (N1883, N1879, N112, N1235, N45);
nor NOR3 (N1884, N1843, N918, N1140);
xor XOR2 (N1885, N1874, N607);
or OR2 (N1886, N1863, N1361);
buf BUF1 (N1887, N1876);
xor XOR2 (N1888, N1875, N1252);
and AND2 (N1889, N1882, N692);
xor XOR2 (N1890, N1887, N1508);
nand NAND4 (N1891, N1885, N1038, N133, N727);
buf BUF1 (N1892, N1888);
or OR4 (N1893, N1886, N116, N753, N814);
or OR4 (N1894, N1892, N1616, N219, N274);
xor XOR2 (N1895, N1880, N1080);
buf BUF1 (N1896, N1889);
and AND4 (N1897, N1891, N1137, N922, N1099);
or OR3 (N1898, N1873, N1780, N308);
and AND3 (N1899, N1895, N120, N948);
and AND3 (N1900, N1881, N1515, N1440);
buf BUF1 (N1901, N1883);
or OR4 (N1902, N1897, N1851, N751, N65);
xor XOR2 (N1903, N1898, N1665);
not NOT1 (N1904, N1890);
xor XOR2 (N1905, N1894, N1654);
or OR4 (N1906, N1902, N1193, N322, N387);
buf BUF1 (N1907, N1900);
nand NAND4 (N1908, N1905, N403, N155, N1031);
buf BUF1 (N1909, N1904);
nand NAND4 (N1910, N1899, N217, N453, N1615);
nand NAND3 (N1911, N1903, N1481, N152);
or OR3 (N1912, N1909, N244, N1768);
xor XOR2 (N1913, N1912, N578);
or OR2 (N1914, N1884, N510);
not NOT1 (N1915, N1893);
buf BUF1 (N1916, N1896);
xor XOR2 (N1917, N1914, N1349);
nand NAND2 (N1918, N1907, N1386);
not NOT1 (N1919, N1908);
not NOT1 (N1920, N1917);
or OR3 (N1921, N1913, N449, N1124);
nand NAND4 (N1922, N1919, N827, N997, N1842);
nand NAND3 (N1923, N1922, N36, N338);
xor XOR2 (N1924, N1921, N965);
not NOT1 (N1925, N1910);
buf BUF1 (N1926, N1925);
not NOT1 (N1927, N1911);
nor NOR4 (N1928, N1906, N1800, N1048, N1422);
not NOT1 (N1929, N1927);
nor NOR4 (N1930, N1918, N1386, N435, N1424);
xor XOR2 (N1931, N1923, N157);
buf BUF1 (N1932, N1915);
or OR3 (N1933, N1932, N1801, N169);
nor NOR4 (N1934, N1901, N1801, N182, N300);
nand NAND3 (N1935, N1931, N18, N64);
not NOT1 (N1936, N1935);
or OR2 (N1937, N1916, N1221);
and AND3 (N1938, N1924, N1614, N1797);
nor NOR2 (N1939, N1936, N825);
buf BUF1 (N1940, N1920);
nand NAND3 (N1941, N1940, N366, N1867);
buf BUF1 (N1942, N1928);
nor NOR4 (N1943, N1926, N1829, N946, N1549);
or OR3 (N1944, N1937, N816, N437);
buf BUF1 (N1945, N1943);
not NOT1 (N1946, N1930);
and AND3 (N1947, N1934, N216, N1307);
and AND3 (N1948, N1942, N1698, N704);
not NOT1 (N1949, N1947);
not NOT1 (N1950, N1949);
and AND2 (N1951, N1939, N854);
nor NOR3 (N1952, N1945, N1063, N1301);
nor NOR3 (N1953, N1948, N1006, N1816);
nor NOR2 (N1954, N1933, N231);
or OR2 (N1955, N1938, N1120);
nor NOR3 (N1956, N1953, N1795, N1765);
or OR2 (N1957, N1951, N981);
buf BUF1 (N1958, N1929);
buf BUF1 (N1959, N1941);
xor XOR2 (N1960, N1946, N127);
or OR4 (N1961, N1960, N551, N1404, N1641);
xor XOR2 (N1962, N1955, N1230);
and AND2 (N1963, N1961, N787);
not NOT1 (N1964, N1950);
and AND4 (N1965, N1952, N191, N645, N1765);
or OR4 (N1966, N1944, N371, N836, N290);
buf BUF1 (N1967, N1958);
and AND2 (N1968, N1954, N403);
nand NAND4 (N1969, N1957, N406, N762, N1908);
nand NAND4 (N1970, N1963, N1564, N1741, N314);
xor XOR2 (N1971, N1956, N93);
xor XOR2 (N1972, N1962, N461);
and AND4 (N1973, N1965, N328, N440, N42);
and AND2 (N1974, N1970, N1225);
nand NAND3 (N1975, N1959, N1295, N814);
nor NOR4 (N1976, N1971, N1241, N818, N870);
xor XOR2 (N1977, N1969, N1079);
or OR4 (N1978, N1975, N381, N1158, N1953);
nand NAND3 (N1979, N1968, N1751, N1531);
nand NAND3 (N1980, N1974, N1280, N1267);
and AND3 (N1981, N1979, N1184, N136);
nand NAND3 (N1982, N1966, N1113, N252);
buf BUF1 (N1983, N1972);
not NOT1 (N1984, N1973);
nor NOR4 (N1985, N1983, N1521, N1358, N1691);
and AND2 (N1986, N1984, N725);
nor NOR2 (N1987, N1964, N863);
nor NOR3 (N1988, N1978, N1143, N568);
buf BUF1 (N1989, N1980);
nand NAND3 (N1990, N1967, N85, N1241);
buf BUF1 (N1991, N1985);
or OR3 (N1992, N1986, N1959, N406);
or OR4 (N1993, N1988, N1936, N1864, N1428);
or OR2 (N1994, N1989, N1220);
and AND2 (N1995, N1976, N1293);
nor NOR4 (N1996, N1977, N1647, N359, N953);
buf BUF1 (N1997, N1995);
nand NAND3 (N1998, N1994, N1820, N1075);
or OR3 (N1999, N1987, N1531, N1180);
nor NOR3 (N2000, N1990, N1400, N86);
not NOT1 (N2001, N1997);
not NOT1 (N2002, N1999);
nor NOR3 (N2003, N1981, N1130, N1569);
or OR3 (N2004, N1992, N1382, N259);
xor XOR2 (N2005, N2000, N871);
nor NOR3 (N2006, N1982, N838, N710);
and AND3 (N2007, N2001, N443, N598);
not NOT1 (N2008, N2004);
and AND4 (N2009, N2008, N1590, N235, N757);
not NOT1 (N2010, N2002);
nand NAND2 (N2011, N2010, N1684);
nand NAND2 (N2012, N2005, N50);
buf BUF1 (N2013, N2003);
not NOT1 (N2014, N2013);
not NOT1 (N2015, N2009);
nand NAND3 (N2016, N2015, N564, N286);
not NOT1 (N2017, N2011);
or OR2 (N2018, N2014, N1918);
not NOT1 (N2019, N1993);
buf BUF1 (N2020, N2017);
buf BUF1 (N2021, N2018);
not NOT1 (N2022, N2007);
or OR2 (N2023, N2016, N1206);
xor XOR2 (N2024, N2020, N66);
nand NAND2 (N2025, N1998, N1733);
not NOT1 (N2026, N2022);
not NOT1 (N2027, N2025);
not NOT1 (N2028, N2027);
and AND3 (N2029, N2006, N1424, N1337);
nor NOR4 (N2030, N1996, N1139, N1905, N1828);
xor XOR2 (N2031, N2024, N929);
and AND3 (N2032, N2030, N1848, N105);
buf BUF1 (N2033, N2021);
and AND4 (N2034, N2023, N933, N1093, N1364);
buf BUF1 (N2035, N2026);
xor XOR2 (N2036, N2019, N1071);
and AND4 (N2037, N2036, N750, N1469, N726);
and AND4 (N2038, N2035, N15, N2012, N1692);
xor XOR2 (N2039, N641, N1278);
not NOT1 (N2040, N2037);
nand NAND4 (N2041, N2028, N29, N176, N1726);
nor NOR3 (N2042, N2039, N1430, N1195);
buf BUF1 (N2043, N2038);
nor NOR2 (N2044, N2029, N1196);
or OR2 (N2045, N2033, N1830);
or OR4 (N2046, N2031, N202, N1447, N361);
nand NAND4 (N2047, N2045, N1207, N1934, N554);
and AND3 (N2048, N2041, N1979, N1045);
buf BUF1 (N2049, N2044);
xor XOR2 (N2050, N2049, N1803);
and AND2 (N2051, N1991, N1219);
xor XOR2 (N2052, N2046, N1562);
xor XOR2 (N2053, N2032, N943);
buf BUF1 (N2054, N2052);
or OR4 (N2055, N2054, N766, N821, N915);
not NOT1 (N2056, N2048);
nor NOR2 (N2057, N2043, N1462);
buf BUF1 (N2058, N2034);
and AND4 (N2059, N2055, N1075, N943, N527);
buf BUF1 (N2060, N2040);
xor XOR2 (N2061, N2050, N1273);
nor NOR3 (N2062, N2053, N1435, N508);
nand NAND3 (N2063, N2059, N45, N1012);
and AND2 (N2064, N2063, N976);
nor NOR3 (N2065, N2042, N1416, N266);
nand NAND3 (N2066, N2056, N348, N2054);
nand NAND2 (N2067, N2062, N1437);
and AND3 (N2068, N2057, N1168, N401);
or OR3 (N2069, N2067, N1043, N185);
buf BUF1 (N2070, N2066);
not NOT1 (N2071, N2069);
and AND2 (N2072, N2047, N659);
xor XOR2 (N2073, N2071, N1108);
buf BUF1 (N2074, N2072);
or OR2 (N2075, N2064, N434);
or OR2 (N2076, N2075, N767);
or OR4 (N2077, N2061, N129, N1315, N1518);
not NOT1 (N2078, N2060);
buf BUF1 (N2079, N2058);
not NOT1 (N2080, N2068);
nor NOR4 (N2081, N2073, N427, N4, N1963);
xor XOR2 (N2082, N2076, N1767);
xor XOR2 (N2083, N2079, N580);
and AND2 (N2084, N2065, N651);
nand NAND2 (N2085, N2080, N394);
buf BUF1 (N2086, N2082);
nor NOR2 (N2087, N2070, N992);
or OR3 (N2088, N2077, N1747, N113);
nor NOR2 (N2089, N2084, N1517);
nor NOR3 (N2090, N2085, N1531, N217);
and AND4 (N2091, N2088, N1675, N377, N775);
or OR4 (N2092, N2081, N714, N544, N2024);
nor NOR2 (N2093, N2091, N354);
buf BUF1 (N2094, N2086);
buf BUF1 (N2095, N2083);
not NOT1 (N2096, N2094);
buf BUF1 (N2097, N2051);
or OR2 (N2098, N2093, N1325);
buf BUF1 (N2099, N2087);
buf BUF1 (N2100, N2089);
and AND2 (N2101, N2090, N699);
xor XOR2 (N2102, N2099, N463);
and AND4 (N2103, N2102, N867, N1876, N86);
not NOT1 (N2104, N2097);
or OR3 (N2105, N2098, N662, N1569);
not NOT1 (N2106, N2105);
nor NOR4 (N2107, N2092, N300, N842, N2076);
and AND3 (N2108, N2096, N2039, N774);
not NOT1 (N2109, N2095);
nand NAND4 (N2110, N2107, N2012, N1150, N455);
nand NAND3 (N2111, N2110, N1182, N662);
or OR4 (N2112, N2104, N1754, N235, N1059);
nand NAND4 (N2113, N2100, N653, N1200, N653);
and AND2 (N2114, N2106, N609);
buf BUF1 (N2115, N2114);
nand NAND3 (N2116, N2078, N828, N542);
nor NOR2 (N2117, N2101, N1819);
nor NOR2 (N2118, N2116, N1288);
and AND4 (N2119, N2113, N1696, N1364, N289);
buf BUF1 (N2120, N2117);
buf BUF1 (N2121, N2074);
nand NAND2 (N2122, N2118, N23);
xor XOR2 (N2123, N2115, N536);
and AND2 (N2124, N2122, N1016);
not NOT1 (N2125, N2108);
nor NOR2 (N2126, N2112, N1298);
not NOT1 (N2127, N2123);
nand NAND2 (N2128, N2109, N1393);
nor NOR4 (N2129, N2126, N692, N979, N37);
nand NAND3 (N2130, N2111, N1953, N1139);
nor NOR4 (N2131, N2119, N405, N826, N1206);
buf BUF1 (N2132, N2103);
nand NAND2 (N2133, N2125, N489);
xor XOR2 (N2134, N2120, N1922);
and AND4 (N2135, N2127, N2057, N1181, N1729);
not NOT1 (N2136, N2124);
xor XOR2 (N2137, N2130, N232);
or OR4 (N2138, N2133, N842, N388, N485);
buf BUF1 (N2139, N2131);
and AND4 (N2140, N2138, N980, N162, N333);
xor XOR2 (N2141, N2137, N1828);
buf BUF1 (N2142, N2121);
xor XOR2 (N2143, N2128, N441);
nand NAND2 (N2144, N2143, N1270);
nor NOR4 (N2145, N2140, N1035, N1453, N392);
not NOT1 (N2146, N2134);
nand NAND4 (N2147, N2141, N878, N64, N1826);
nand NAND2 (N2148, N2132, N1369);
nand NAND2 (N2149, N2148, N1568);
xor XOR2 (N2150, N2144, N466);
not NOT1 (N2151, N2147);
nand NAND3 (N2152, N2139, N625, N818);
and AND3 (N2153, N2151, N1320, N549);
xor XOR2 (N2154, N2152, N27);
and AND3 (N2155, N2129, N1026, N1082);
buf BUF1 (N2156, N2150);
xor XOR2 (N2157, N2142, N539);
xor XOR2 (N2158, N2157, N1747);
xor XOR2 (N2159, N2136, N1476);
xor XOR2 (N2160, N2145, N1972);
nand NAND2 (N2161, N2158, N1785);
not NOT1 (N2162, N2149);
nor NOR2 (N2163, N2153, N1312);
not NOT1 (N2164, N2156);
nor NOR2 (N2165, N2161, N693);
not NOT1 (N2166, N2160);
or OR4 (N2167, N2146, N1937, N1352, N1784);
nand NAND3 (N2168, N2154, N1194, N1188);
nand NAND2 (N2169, N2168, N49);
xor XOR2 (N2170, N2159, N1783);
xor XOR2 (N2171, N2170, N1328);
nand NAND3 (N2172, N2167, N393, N997);
or OR3 (N2173, N2162, N2168, N1269);
xor XOR2 (N2174, N2135, N1730);
buf BUF1 (N2175, N2165);
xor XOR2 (N2176, N2166, N1630);
nor NOR3 (N2177, N2172, N570, N1693);
and AND3 (N2178, N2155, N1785, N1940);
buf BUF1 (N2179, N2171);
and AND4 (N2180, N2164, N225, N186, N739);
xor XOR2 (N2181, N2180, N75);
and AND4 (N2182, N2179, N883, N1358, N1659);
or OR2 (N2183, N2178, N2028);
buf BUF1 (N2184, N2177);
and AND2 (N2185, N2163, N1140);
and AND3 (N2186, N2184, N930, N1138);
nor NOR2 (N2187, N2185, N1334);
and AND3 (N2188, N2183, N1845, N821);
not NOT1 (N2189, N2186);
or OR4 (N2190, N2176, N1463, N221, N1479);
or OR3 (N2191, N2174, N2182, N1234);
not NOT1 (N2192, N978);
buf BUF1 (N2193, N2189);
and AND2 (N2194, N2190, N2116);
xor XOR2 (N2195, N2173, N150);
not NOT1 (N2196, N2194);
not NOT1 (N2197, N2188);
buf BUF1 (N2198, N2197);
xor XOR2 (N2199, N2195, N2010);
nand NAND2 (N2200, N2181, N299);
xor XOR2 (N2201, N2196, N1507);
xor XOR2 (N2202, N2200, N1842);
or OR2 (N2203, N2192, N2201);
buf BUF1 (N2204, N392);
nand NAND4 (N2205, N2198, N2110, N263, N263);
or OR4 (N2206, N2202, N36, N366, N222);
not NOT1 (N2207, N2203);
or OR2 (N2208, N2175, N915);
nand NAND4 (N2209, N2193, N644, N1392, N911);
nand NAND2 (N2210, N2169, N358);
and AND4 (N2211, N2210, N855, N955, N1169);
not NOT1 (N2212, N2199);
and AND3 (N2213, N2191, N1294, N872);
nor NOR3 (N2214, N2212, N410, N392);
buf BUF1 (N2215, N2206);
nand NAND2 (N2216, N2215, N1396);
xor XOR2 (N2217, N2208, N2182);
buf BUF1 (N2218, N2216);
xor XOR2 (N2219, N2217, N1567);
or OR2 (N2220, N2205, N729);
or OR3 (N2221, N2213, N2010, N1641);
and AND2 (N2222, N2209, N436);
and AND2 (N2223, N2222, N833);
xor XOR2 (N2224, N2220, N613);
nor NOR2 (N2225, N2211, N413);
buf BUF1 (N2226, N2225);
or OR3 (N2227, N2223, N2069, N1121);
xor XOR2 (N2228, N2187, N682);
xor XOR2 (N2229, N2228, N1294);
not NOT1 (N2230, N2227);
nor NOR3 (N2231, N2230, N2165, N492);
buf BUF1 (N2232, N2226);
buf BUF1 (N2233, N2221);
nor NOR2 (N2234, N2207, N58);
not NOT1 (N2235, N2224);
xor XOR2 (N2236, N2235, N1260);
or OR4 (N2237, N2204, N2158, N318, N1869);
nor NOR2 (N2238, N2233, N420);
or OR4 (N2239, N2236, N2233, N131, N1906);
nor NOR2 (N2240, N2218, N73);
not NOT1 (N2241, N2219);
nand NAND3 (N2242, N2238, N176, N1517);
nor NOR2 (N2243, N2232, N1775);
nor NOR2 (N2244, N2243, N2159);
and AND2 (N2245, N2234, N1191);
not NOT1 (N2246, N2241);
buf BUF1 (N2247, N2239);
or OR4 (N2248, N2242, N1006, N2064, N915);
and AND3 (N2249, N2237, N828, N863);
nand NAND2 (N2250, N2246, N323);
and AND2 (N2251, N2249, N152);
buf BUF1 (N2252, N2214);
xor XOR2 (N2253, N2248, N395);
xor XOR2 (N2254, N2231, N602);
and AND2 (N2255, N2229, N1259);
xor XOR2 (N2256, N2247, N60);
and AND3 (N2257, N2252, N1802, N1382);
or OR2 (N2258, N2253, N726);
nor NOR2 (N2259, N2257, N96);
and AND2 (N2260, N2250, N323);
and AND4 (N2261, N2256, N1787, N1528, N1443);
or OR3 (N2262, N2261, N56, N2248);
nand NAND2 (N2263, N2262, N2172);
or OR3 (N2264, N2259, N1977, N1831);
not NOT1 (N2265, N2264);
nand NAND4 (N2266, N2258, N901, N1965, N215);
buf BUF1 (N2267, N2244);
not NOT1 (N2268, N2251);
not NOT1 (N2269, N2255);
buf BUF1 (N2270, N2263);
nand NAND3 (N2271, N2245, N533, N407);
buf BUF1 (N2272, N2269);
nor NOR2 (N2273, N2240, N613);
or OR3 (N2274, N2254, N315, N1648);
not NOT1 (N2275, N2265);
or OR2 (N2276, N2268, N1142);
and AND3 (N2277, N2276, N1393, N649);
nand NAND3 (N2278, N2273, N1454, N2247);
nor NOR2 (N2279, N2272, N1011);
buf BUF1 (N2280, N2278);
not NOT1 (N2281, N2270);
nand NAND2 (N2282, N2281, N104);
or OR2 (N2283, N2267, N1508);
xor XOR2 (N2284, N2275, N47);
buf BUF1 (N2285, N2280);
or OR4 (N2286, N2282, N637, N562, N181);
nand NAND4 (N2287, N2279, N918, N2092, N196);
and AND2 (N2288, N2285, N1881);
buf BUF1 (N2289, N2277);
buf BUF1 (N2290, N2260);
buf BUF1 (N2291, N2266);
nor NOR2 (N2292, N2291, N183);
buf BUF1 (N2293, N2284);
not NOT1 (N2294, N2271);
not NOT1 (N2295, N2287);
xor XOR2 (N2296, N2290, N1459);
xor XOR2 (N2297, N2283, N6);
xor XOR2 (N2298, N2286, N189);
buf BUF1 (N2299, N2298);
not NOT1 (N2300, N2299);
nor NOR3 (N2301, N2292, N592, N1534);
buf BUF1 (N2302, N2301);
and AND4 (N2303, N2297, N1814, N924, N389);
or OR2 (N2304, N2303, N844);
xor XOR2 (N2305, N2304, N1437);
buf BUF1 (N2306, N2294);
nand NAND3 (N2307, N2293, N1386, N619);
or OR2 (N2308, N2306, N1136);
xor XOR2 (N2309, N2305, N1161);
nor NOR4 (N2310, N2308, N1122, N1974, N1328);
not NOT1 (N2311, N2309);
nand NAND4 (N2312, N2288, N647, N1069, N820);
nand NAND2 (N2313, N2274, N77);
or OR4 (N2314, N2296, N501, N1350, N1357);
not NOT1 (N2315, N2312);
or OR3 (N2316, N2310, N1493, N577);
xor XOR2 (N2317, N2316, N274);
and AND4 (N2318, N2313, N2031, N838, N1545);
nor NOR4 (N2319, N2315, N1940, N588, N6);
and AND3 (N2320, N2307, N764, N1036);
nand NAND4 (N2321, N2320, N1748, N1180, N1306);
nor NOR4 (N2322, N2318, N1878, N1566, N1193);
buf BUF1 (N2323, N2321);
buf BUF1 (N2324, N2300);
or OR2 (N2325, N2295, N997);
nor NOR4 (N2326, N2302, N2190, N53, N853);
not NOT1 (N2327, N2322);
not NOT1 (N2328, N2326);
buf BUF1 (N2329, N2323);
nand NAND3 (N2330, N2329, N952, N2034);
buf BUF1 (N2331, N2330);
and AND4 (N2332, N2327, N945, N616, N124);
not NOT1 (N2333, N2311);
or OR4 (N2334, N2314, N2026, N72, N1805);
nand NAND2 (N2335, N2328, N133);
and AND2 (N2336, N2332, N1649);
and AND3 (N2337, N2335, N279, N425);
buf BUF1 (N2338, N2331);
not NOT1 (N2339, N2334);
not NOT1 (N2340, N2338);
xor XOR2 (N2341, N2333, N993);
and AND2 (N2342, N2319, N277);
and AND3 (N2343, N2342, N948, N1162);
buf BUF1 (N2344, N2336);
buf BUF1 (N2345, N2343);
not NOT1 (N2346, N2344);
xor XOR2 (N2347, N2346, N241);
nor NOR3 (N2348, N2341, N1617, N836);
nor NOR4 (N2349, N2324, N1476, N1699, N1211);
and AND4 (N2350, N2339, N1942, N1948, N483);
nor NOR4 (N2351, N2348, N1545, N591, N1834);
nor NOR4 (N2352, N2349, N2062, N1893, N257);
and AND4 (N2353, N2340, N1731, N462, N373);
nor NOR2 (N2354, N2325, N829);
not NOT1 (N2355, N2317);
nor NOR4 (N2356, N2345, N152, N1492, N1592);
nand NAND2 (N2357, N2347, N1356);
buf BUF1 (N2358, N2350);
or OR4 (N2359, N2356, N470, N1915, N627);
nor NOR4 (N2360, N2351, N1334, N2306, N1440);
buf BUF1 (N2361, N2357);
nand NAND3 (N2362, N2360, N1097, N2290);
not NOT1 (N2363, N2359);
nor NOR3 (N2364, N2361, N1757, N1918);
and AND3 (N2365, N2354, N1466, N2194);
or OR4 (N2366, N2337, N1231, N346, N2294);
xor XOR2 (N2367, N2358, N1495);
not NOT1 (N2368, N2366);
and AND4 (N2369, N2355, N856, N1865, N1045);
nand NAND4 (N2370, N2369, N369, N1185, N531);
nand NAND4 (N2371, N2363, N1454, N1789, N519);
or OR4 (N2372, N2365, N620, N211, N80);
or OR4 (N2373, N2289, N554, N2213, N1035);
nand NAND3 (N2374, N2352, N1402, N2290);
nor NOR3 (N2375, N2353, N718, N1457);
nand NAND4 (N2376, N2375, N2325, N1685, N2085);
buf BUF1 (N2377, N2372);
buf BUF1 (N2378, N2377);
xor XOR2 (N2379, N2370, N1949);
not NOT1 (N2380, N2373);
nand NAND2 (N2381, N2380, N607);
xor XOR2 (N2382, N2367, N789);
nor NOR2 (N2383, N2381, N2311);
or OR2 (N2384, N2376, N2105);
xor XOR2 (N2385, N2378, N141);
not NOT1 (N2386, N2371);
and AND2 (N2387, N2383, N1393);
not NOT1 (N2388, N2364);
buf BUF1 (N2389, N2374);
xor XOR2 (N2390, N2384, N391);
xor XOR2 (N2391, N2387, N971);
nor NOR2 (N2392, N2389, N789);
or OR4 (N2393, N2391, N165, N853, N1231);
or OR3 (N2394, N2382, N1438, N257);
not NOT1 (N2395, N2368);
not NOT1 (N2396, N2390);
nand NAND4 (N2397, N2396, N2240, N1606, N1228);
or OR3 (N2398, N2394, N1994, N1171);
or OR4 (N2399, N2392, N639, N1724, N1950);
nor NOR3 (N2400, N2397, N1288, N1939);
or OR4 (N2401, N2398, N773, N139, N1107);
buf BUF1 (N2402, N2386);
not NOT1 (N2403, N2362);
not NOT1 (N2404, N2379);
buf BUF1 (N2405, N2385);
xor XOR2 (N2406, N2404, N1778);
and AND3 (N2407, N2400, N602, N82);
xor XOR2 (N2408, N2405, N1661);
nand NAND2 (N2409, N2401, N332);
xor XOR2 (N2410, N2395, N657);
buf BUF1 (N2411, N2393);
not NOT1 (N2412, N2399);
not NOT1 (N2413, N2412);
not NOT1 (N2414, N2407);
buf BUF1 (N2415, N2402);
nand NAND2 (N2416, N2413, N385);
nand NAND4 (N2417, N2416, N1740, N1372, N2191);
nor NOR3 (N2418, N2406, N2240, N828);
not NOT1 (N2419, N2414);
xor XOR2 (N2420, N2417, N229);
buf BUF1 (N2421, N2419);
or OR4 (N2422, N2415, N1203, N148, N1113);
nand NAND4 (N2423, N2418, N530, N1230, N875);
or OR4 (N2424, N2403, N1703, N981, N134);
nand NAND4 (N2425, N2420, N2297, N2076, N1165);
buf BUF1 (N2426, N2422);
and AND3 (N2427, N2388, N1157, N1229);
not NOT1 (N2428, N2425);
buf BUF1 (N2429, N2427);
and AND2 (N2430, N2428, N1222);
not NOT1 (N2431, N2411);
or OR2 (N2432, N2431, N943);
or OR3 (N2433, N2424, N2387, N1648);
not NOT1 (N2434, N2423);
xor XOR2 (N2435, N2421, N12);
buf BUF1 (N2436, N2426);
nor NOR3 (N2437, N2408, N2219, N2385);
nor NOR3 (N2438, N2432, N2225, N2404);
nor NOR4 (N2439, N2437, N972, N1946, N1638);
nor NOR3 (N2440, N2436, N1449, N1536);
nand NAND2 (N2441, N2409, N2193);
buf BUF1 (N2442, N2429);
and AND2 (N2443, N2442, N605);
and AND3 (N2444, N2440, N1518, N1570);
not NOT1 (N2445, N2438);
xor XOR2 (N2446, N2410, N1837);
nand NAND2 (N2447, N2445, N93);
or OR4 (N2448, N2446, N1353, N268, N8);
not NOT1 (N2449, N2435);
nor NOR2 (N2450, N2447, N433);
nand NAND3 (N2451, N2430, N2128, N1855);
not NOT1 (N2452, N2441);
xor XOR2 (N2453, N2452, N131);
buf BUF1 (N2454, N2443);
xor XOR2 (N2455, N2439, N841);
buf BUF1 (N2456, N2454);
xor XOR2 (N2457, N2455, N651);
buf BUF1 (N2458, N2456);
buf BUF1 (N2459, N2453);
nor NOR2 (N2460, N2459, N1368);
xor XOR2 (N2461, N2458, N780);
or OR4 (N2462, N2451, N1648, N1894, N795);
buf BUF1 (N2463, N2448);
xor XOR2 (N2464, N2434, N2430);
not NOT1 (N2465, N2462);
nor NOR2 (N2466, N2433, N1584);
nand NAND4 (N2467, N2450, N1560, N1110, N511);
and AND2 (N2468, N2461, N1629);
not NOT1 (N2469, N2465);
nand NAND3 (N2470, N2460, N984, N712);
xor XOR2 (N2471, N2449, N418);
buf BUF1 (N2472, N2468);
not NOT1 (N2473, N2467);
or OR4 (N2474, N2444, N217, N478, N2361);
xor XOR2 (N2475, N2469, N2473);
and AND4 (N2476, N2318, N783, N564, N468);
nor NOR3 (N2477, N2476, N2281, N263);
or OR4 (N2478, N2457, N791, N1132, N1547);
nand NAND4 (N2479, N2474, N430, N313, N356);
buf BUF1 (N2480, N2475);
nor NOR3 (N2481, N2480, N166, N972);
xor XOR2 (N2482, N2481, N213);
nand NAND2 (N2483, N2477, N560);
nand NAND4 (N2484, N2478, N904, N128, N2021);
not NOT1 (N2485, N2484);
buf BUF1 (N2486, N2463);
and AND4 (N2487, N2485, N479, N2186, N58);
xor XOR2 (N2488, N2487, N2402);
xor XOR2 (N2489, N2482, N1629);
and AND2 (N2490, N2466, N807);
nand NAND3 (N2491, N2471, N690, N1593);
not NOT1 (N2492, N2464);
xor XOR2 (N2493, N2492, N1315);
nor NOR2 (N2494, N2493, N2481);
xor XOR2 (N2495, N2490, N1345);
nand NAND3 (N2496, N2479, N2042, N1339);
xor XOR2 (N2497, N2483, N813);
or OR2 (N2498, N2486, N785);
or OR4 (N2499, N2495, N63, N2332, N1066);
or OR4 (N2500, N2489, N1822, N1639, N1534);
buf BUF1 (N2501, N2491);
or OR3 (N2502, N2500, N1843, N1225);
not NOT1 (N2503, N2488);
buf BUF1 (N2504, N2501);
buf BUF1 (N2505, N2503);
nor NOR4 (N2506, N2496, N170, N1098, N1555);
nor NOR2 (N2507, N2470, N1711);
buf BUF1 (N2508, N2498);
xor XOR2 (N2509, N2494, N141);
nand NAND3 (N2510, N2499, N1400, N368);
xor XOR2 (N2511, N2510, N1215);
xor XOR2 (N2512, N2509, N799);
buf BUF1 (N2513, N2502);
nand NAND2 (N2514, N2508, N983);
and AND2 (N2515, N2472, N1366);
and AND2 (N2516, N2507, N46);
nor NOR2 (N2517, N2506, N2054);
xor XOR2 (N2518, N2516, N794);
not NOT1 (N2519, N2515);
and AND2 (N2520, N2497, N1145);
nand NAND3 (N2521, N2520, N756, N1809);
buf BUF1 (N2522, N2521);
nor NOR4 (N2523, N2512, N1028, N511, N1388);
and AND4 (N2524, N2517, N676, N973, N1791);
xor XOR2 (N2525, N2523, N2503);
not NOT1 (N2526, N2518);
not NOT1 (N2527, N2524);
or OR3 (N2528, N2527, N2523, N564);
or OR2 (N2529, N2514, N971);
nor NOR2 (N2530, N2505, N1233);
and AND4 (N2531, N2522, N948, N1075, N2138);
and AND4 (N2532, N2504, N1625, N471, N554);
buf BUF1 (N2533, N2526);
or OR2 (N2534, N2513, N782);
buf BUF1 (N2535, N2533);
not NOT1 (N2536, N2529);
buf BUF1 (N2537, N2530);
nor NOR2 (N2538, N2536, N260);
nor NOR2 (N2539, N2532, N1981);
buf BUF1 (N2540, N2534);
and AND3 (N2541, N2525, N1632, N503);
or OR3 (N2542, N2519, N1691, N1129);
not NOT1 (N2543, N2540);
nor NOR4 (N2544, N2539, N1893, N665, N2421);
and AND4 (N2545, N2535, N1488, N21, N2102);
not NOT1 (N2546, N2528);
buf BUF1 (N2547, N2546);
or OR4 (N2548, N2511, N2477, N1238, N1568);
nor NOR3 (N2549, N2537, N1264, N777);
not NOT1 (N2550, N2542);
and AND2 (N2551, N2548, N1284);
or OR4 (N2552, N2531, N256, N2331, N737);
nor NOR2 (N2553, N2552, N1673);
and AND2 (N2554, N2547, N1423);
or OR2 (N2555, N2551, N1670);
and AND2 (N2556, N2541, N1208);
or OR2 (N2557, N2543, N1134);
or OR4 (N2558, N2550, N1364, N2070, N326);
or OR2 (N2559, N2549, N24);
nand NAND3 (N2560, N2545, N44, N669);
not NOT1 (N2561, N2544);
not NOT1 (N2562, N2553);
nor NOR4 (N2563, N2559, N1434, N1753, N2175);
nand NAND2 (N2564, N2538, N1196);
buf BUF1 (N2565, N2556);
xor XOR2 (N2566, N2563, N999);
buf BUF1 (N2567, N2564);
and AND4 (N2568, N2566, N983, N2560, N2192);
buf BUF1 (N2569, N2303);
buf BUF1 (N2570, N2568);
nor NOR2 (N2571, N2561, N1480);
not NOT1 (N2572, N2558);
buf BUF1 (N2573, N2565);
nand NAND3 (N2574, N2567, N813, N171);
nor NOR3 (N2575, N2557, N697, N1874);
not NOT1 (N2576, N2569);
nand NAND4 (N2577, N2576, N492, N76, N1514);
xor XOR2 (N2578, N2572, N108);
nor NOR4 (N2579, N2554, N242, N2215, N717);
or OR4 (N2580, N2575, N369, N461, N1497);
nand NAND3 (N2581, N2577, N2201, N2229);
xor XOR2 (N2582, N2578, N306);
buf BUF1 (N2583, N2574);
buf BUF1 (N2584, N2582);
xor XOR2 (N2585, N2555, N1284);
nor NOR3 (N2586, N2573, N1922, N582);
and AND2 (N2587, N2570, N1288);
not NOT1 (N2588, N2579);
buf BUF1 (N2589, N2571);
not NOT1 (N2590, N2584);
xor XOR2 (N2591, N2588, N950);
buf BUF1 (N2592, N2587);
or OR2 (N2593, N2591, N603);
and AND2 (N2594, N2590, N2034);
or OR2 (N2595, N2580, N2022);
or OR4 (N2596, N2586, N2358, N1317, N2472);
xor XOR2 (N2597, N2581, N922);
or OR3 (N2598, N2593, N111, N2347);
nor NOR4 (N2599, N2595, N448, N1015, N1500);
nor NOR2 (N2600, N2583, N1257);
not NOT1 (N2601, N2598);
nand NAND4 (N2602, N2596, N2447, N1290, N1035);
xor XOR2 (N2603, N2599, N886);
and AND2 (N2604, N2603, N243);
xor XOR2 (N2605, N2592, N1557);
or OR2 (N2606, N2597, N1393);
nor NOR2 (N2607, N2601, N1197);
buf BUF1 (N2608, N2600);
and AND2 (N2609, N2594, N1579);
xor XOR2 (N2610, N2562, N1033);
xor XOR2 (N2611, N2602, N14);
buf BUF1 (N2612, N2589);
not NOT1 (N2613, N2585);
not NOT1 (N2614, N2607);
nor NOR3 (N2615, N2614, N2181, N2156);
and AND3 (N2616, N2608, N645, N1596);
and AND4 (N2617, N2606, N1762, N1035, N2406);
xor XOR2 (N2618, N2610, N1900);
xor XOR2 (N2619, N2605, N1421);
and AND2 (N2620, N2615, N166);
buf BUF1 (N2621, N2611);
not NOT1 (N2622, N2621);
or OR2 (N2623, N2612, N45);
not NOT1 (N2624, N2618);
nor NOR4 (N2625, N2620, N614, N1417, N937);
and AND3 (N2626, N2619, N462, N549);
or OR2 (N2627, N2623, N1865);
and AND3 (N2628, N2609, N1474, N1652);
buf BUF1 (N2629, N2627);
or OR3 (N2630, N2604, N1132, N2036);
nand NAND2 (N2631, N2626, N2279);
buf BUF1 (N2632, N2617);
buf BUF1 (N2633, N2624);
buf BUF1 (N2634, N2631);
not NOT1 (N2635, N2628);
or OR4 (N2636, N2616, N2127, N23, N1375);
or OR4 (N2637, N2622, N2001, N1694, N1582);
and AND3 (N2638, N2613, N2569, N1061);
buf BUF1 (N2639, N2636);
or OR4 (N2640, N2637, N1806, N2607, N835);
not NOT1 (N2641, N2629);
or OR3 (N2642, N2640, N991, N1013);
nand NAND2 (N2643, N2641, N794);
nor NOR2 (N2644, N2638, N2217);
buf BUF1 (N2645, N2639);
nand NAND3 (N2646, N2643, N1275, N876);
nand NAND2 (N2647, N2632, N1024);
buf BUF1 (N2648, N2647);
xor XOR2 (N2649, N2642, N2075);
nor NOR3 (N2650, N2649, N976, N1935);
nand NAND4 (N2651, N2644, N667, N1917, N1388);
nor NOR4 (N2652, N2634, N1182, N1114, N1490);
buf BUF1 (N2653, N2650);
buf BUF1 (N2654, N2652);
or OR4 (N2655, N2648, N1997, N2183, N1975);
or OR2 (N2656, N2655, N2474);
xor XOR2 (N2657, N2656, N2492);
nand NAND4 (N2658, N2657, N2482, N1732, N1965);
xor XOR2 (N2659, N2630, N893);
buf BUF1 (N2660, N2658);
nor NOR3 (N2661, N2654, N1022, N1024);
nand NAND4 (N2662, N2635, N1796, N1625, N54);
not NOT1 (N2663, N2645);
buf BUF1 (N2664, N2661);
nor NOR3 (N2665, N2646, N128, N840);
nor NOR2 (N2666, N2665, N1839);
buf BUF1 (N2667, N2659);
xor XOR2 (N2668, N2664, N2664);
or OR4 (N2669, N2633, N97, N2532, N599);
not NOT1 (N2670, N2669);
not NOT1 (N2671, N2651);
and AND2 (N2672, N2625, N2083);
buf BUF1 (N2673, N2653);
and AND4 (N2674, N2672, N1686, N1225, N778);
and AND2 (N2675, N2673, N892);
or OR4 (N2676, N2675, N1502, N1487, N2018);
xor XOR2 (N2677, N2671, N296);
or OR3 (N2678, N2670, N656, N2609);
not NOT1 (N2679, N2677);
not NOT1 (N2680, N2668);
xor XOR2 (N2681, N2667, N2168);
xor XOR2 (N2682, N2676, N1054);
xor XOR2 (N2683, N2674, N777);
xor XOR2 (N2684, N2662, N412);
nor NOR2 (N2685, N2683, N2640);
nand NAND3 (N2686, N2681, N2527, N99);
nand NAND3 (N2687, N2686, N1073, N163);
nand NAND3 (N2688, N2679, N1484, N1367);
nand NAND4 (N2689, N2663, N2147, N1532, N2539);
and AND4 (N2690, N2680, N502, N1512, N834);
buf BUF1 (N2691, N2666);
or OR2 (N2692, N2690, N2338);
not NOT1 (N2693, N2678);
xor XOR2 (N2694, N2684, N2560);
not NOT1 (N2695, N2689);
buf BUF1 (N2696, N2682);
not NOT1 (N2697, N2660);
or OR4 (N2698, N2694, N2017, N747, N1574);
and AND3 (N2699, N2696, N2363, N41);
xor XOR2 (N2700, N2685, N2103);
or OR3 (N2701, N2693, N2243, N43);
nand NAND3 (N2702, N2687, N1842, N937);
and AND2 (N2703, N2701, N1510);
nor NOR3 (N2704, N2700, N2585, N106);
xor XOR2 (N2705, N2702, N2245);
nor NOR2 (N2706, N2697, N2443);
xor XOR2 (N2707, N2688, N2133);
buf BUF1 (N2708, N2698);
and AND4 (N2709, N2705, N2292, N1611, N1936);
xor XOR2 (N2710, N2707, N1422);
nand NAND3 (N2711, N2703, N1822, N2609);
nand NAND4 (N2712, N2704, N1851, N1314, N1961);
or OR3 (N2713, N2691, N2005, N1434);
nor NOR2 (N2714, N2695, N477);
and AND3 (N2715, N2692, N2435, N1057);
buf BUF1 (N2716, N2709);
and AND4 (N2717, N2711, N1761, N1698, N1401);
nand NAND3 (N2718, N2712, N1642, N325);
not NOT1 (N2719, N2708);
not NOT1 (N2720, N2699);
not NOT1 (N2721, N2717);
not NOT1 (N2722, N2706);
not NOT1 (N2723, N2716);
and AND4 (N2724, N2722, N331, N2492, N2424);
buf BUF1 (N2725, N2721);
buf BUF1 (N2726, N2715);
xor XOR2 (N2727, N2719, N753);
nor NOR2 (N2728, N2726, N1490);
or OR4 (N2729, N2713, N1022, N2361, N1649);
buf BUF1 (N2730, N2714);
nand NAND2 (N2731, N2727, N1738);
and AND4 (N2732, N2724, N1440, N1250, N2239);
xor XOR2 (N2733, N2723, N520);
xor XOR2 (N2734, N2720, N1243);
or OR2 (N2735, N2733, N816);
buf BUF1 (N2736, N2732);
and AND4 (N2737, N2734, N1754, N564, N1427);
or OR3 (N2738, N2710, N1205, N2430);
xor XOR2 (N2739, N2735, N1724);
nor NOR4 (N2740, N2737, N205, N1845, N2728);
xor XOR2 (N2741, N2709, N2352);
not NOT1 (N2742, N2725);
buf BUF1 (N2743, N2739);
xor XOR2 (N2744, N2742, N1761);
buf BUF1 (N2745, N2730);
buf BUF1 (N2746, N2729);
not NOT1 (N2747, N2738);
or OR3 (N2748, N2747, N668, N1031);
nand NAND3 (N2749, N2744, N2041, N2626);
or OR2 (N2750, N2743, N1514);
xor XOR2 (N2751, N2740, N2123);
xor XOR2 (N2752, N2748, N2377);
nand NAND3 (N2753, N2731, N1952, N1124);
and AND4 (N2754, N2718, N591, N103, N17);
xor XOR2 (N2755, N2753, N2492);
buf BUF1 (N2756, N2755);
xor XOR2 (N2757, N2754, N1120);
buf BUF1 (N2758, N2749);
or OR4 (N2759, N2756, N2122, N393, N234);
or OR2 (N2760, N2758, N1950);
or OR3 (N2761, N2759, N627, N1155);
nand NAND2 (N2762, N2736, N1539);
nor NOR4 (N2763, N2761, N995, N1136, N1374);
or OR3 (N2764, N2752, N1748, N2339);
nand NAND2 (N2765, N2751, N1083);
or OR4 (N2766, N2765, N2066, N244, N1165);
xor XOR2 (N2767, N2766, N1524);
not NOT1 (N2768, N2763);
nand NAND4 (N2769, N2741, N1903, N2293, N23);
and AND2 (N2770, N2745, N956);
and AND4 (N2771, N2769, N1377, N477, N1922);
and AND3 (N2772, N2768, N1521, N1566);
buf BUF1 (N2773, N2764);
xor XOR2 (N2774, N2760, N2726);
not NOT1 (N2775, N2757);
not NOT1 (N2776, N2770);
and AND3 (N2777, N2774, N1741, N461);
nand NAND4 (N2778, N2762, N217, N2617, N658);
xor XOR2 (N2779, N2777, N2084);
or OR2 (N2780, N2776, N2282);
or OR3 (N2781, N2775, N2735, N1694);
and AND3 (N2782, N2779, N1899, N1535);
and AND2 (N2783, N2782, N1256);
not NOT1 (N2784, N2767);
nand NAND4 (N2785, N2781, N2523, N2423, N646);
or OR4 (N2786, N2780, N1135, N1741, N2178);
xor XOR2 (N2787, N2783, N230);
xor XOR2 (N2788, N2784, N608);
nand NAND4 (N2789, N2778, N2216, N2049, N1130);
and AND3 (N2790, N2787, N1177, N987);
buf BUF1 (N2791, N2772);
nand NAND2 (N2792, N2788, N889);
buf BUF1 (N2793, N2750);
buf BUF1 (N2794, N2746);
nand NAND4 (N2795, N2792, N2682, N2437, N662);
or OR3 (N2796, N2789, N2539, N2302);
xor XOR2 (N2797, N2786, N2315);
or OR3 (N2798, N2797, N1019, N289);
xor XOR2 (N2799, N2793, N2180);
nor NOR3 (N2800, N2791, N29, N535);
not NOT1 (N2801, N2796);
nor NOR2 (N2802, N2801, N72);
buf BUF1 (N2803, N2795);
not NOT1 (N2804, N2773);
nand NAND4 (N2805, N2799, N2604, N942, N109);
nor NOR4 (N2806, N2785, N1571, N1255, N2405);
xor XOR2 (N2807, N2800, N1562);
nor NOR2 (N2808, N2806, N1993);
nand NAND4 (N2809, N2798, N1839, N1312, N939);
or OR3 (N2810, N2790, N5, N1051);
buf BUF1 (N2811, N2810);
nand NAND2 (N2812, N2808, N2649);
nor NOR4 (N2813, N2794, N1920, N1703, N353);
and AND2 (N2814, N2811, N2037);
not NOT1 (N2815, N2813);
not NOT1 (N2816, N2812);
nand NAND2 (N2817, N2815, N812);
xor XOR2 (N2818, N2802, N1357);
xor XOR2 (N2819, N2804, N510);
xor XOR2 (N2820, N2809, N1431);
nor NOR3 (N2821, N2820, N1962, N2450);
nor NOR3 (N2822, N2821, N1431, N2625);
nand NAND4 (N2823, N2803, N2032, N751, N2433);
nand NAND2 (N2824, N2807, N985);
and AND2 (N2825, N2824, N1499);
nand NAND2 (N2826, N2771, N2203);
or OR4 (N2827, N2817, N1040, N2095, N1863);
not NOT1 (N2828, N2825);
xor XOR2 (N2829, N2826, N283);
nor NOR4 (N2830, N2822, N243, N1514, N2690);
nand NAND2 (N2831, N2818, N2504);
and AND2 (N2832, N2819, N2510);
not NOT1 (N2833, N2831);
and AND2 (N2834, N2829, N2526);
xor XOR2 (N2835, N2827, N2614);
and AND4 (N2836, N2828, N2446, N2524, N202);
xor XOR2 (N2837, N2834, N261);
or OR4 (N2838, N2805, N2729, N1282, N2830);
or OR3 (N2839, N1228, N2835, N1929);
xor XOR2 (N2840, N1437, N2729);
and AND2 (N2841, N2833, N2522);
nor NOR3 (N2842, N2841, N1695, N1635);
and AND3 (N2843, N2816, N2308, N400);
xor XOR2 (N2844, N2832, N2620);
xor XOR2 (N2845, N2844, N415);
xor XOR2 (N2846, N2839, N2315);
nor NOR2 (N2847, N2842, N410);
nor NOR3 (N2848, N2836, N123, N619);
or OR3 (N2849, N2837, N1780, N127);
not NOT1 (N2850, N2843);
xor XOR2 (N2851, N2823, N772);
or OR2 (N2852, N2846, N2391);
nor NOR4 (N2853, N2851, N2449, N281, N1904);
or OR4 (N2854, N2853, N2023, N2735, N2735);
nor NOR2 (N2855, N2849, N2366);
or OR4 (N2856, N2850, N2679, N15, N2002);
not NOT1 (N2857, N2840);
buf BUF1 (N2858, N2838);
xor XOR2 (N2859, N2852, N2772);
nand NAND2 (N2860, N2856, N1439);
or OR4 (N2861, N2859, N1271, N332, N1487);
nor NOR2 (N2862, N2845, N1410);
and AND3 (N2863, N2814, N2224, N23);
xor XOR2 (N2864, N2861, N2465);
xor XOR2 (N2865, N2860, N811);
and AND4 (N2866, N2847, N1129, N2475, N1155);
nand NAND2 (N2867, N2865, N801);
nor NOR2 (N2868, N2857, N1837);
not NOT1 (N2869, N2864);
nor NOR2 (N2870, N2867, N1238);
nand NAND4 (N2871, N2848, N1797, N510, N1228);
xor XOR2 (N2872, N2855, N2673);
nand NAND3 (N2873, N2870, N2800, N2072);
buf BUF1 (N2874, N2868);
or OR2 (N2875, N2866, N1378);
nor NOR4 (N2876, N2873, N2184, N1811, N476);
or OR2 (N2877, N2875, N880);
not NOT1 (N2878, N2854);
nand NAND2 (N2879, N2858, N1177);
buf BUF1 (N2880, N2872);
buf BUF1 (N2881, N2869);
and AND4 (N2882, N2878, N853, N612, N1962);
or OR2 (N2883, N2879, N330);
and AND4 (N2884, N2882, N873, N2652, N2878);
not NOT1 (N2885, N2880);
or OR3 (N2886, N2863, N297, N2849);
or OR4 (N2887, N2886, N1750, N1793, N2034);
and AND2 (N2888, N2871, N1407);
and AND4 (N2889, N2885, N1012, N1723, N865);
xor XOR2 (N2890, N2862, N692);
xor XOR2 (N2891, N2874, N641);
or OR3 (N2892, N2876, N1477, N2343);
buf BUF1 (N2893, N2891);
not NOT1 (N2894, N2888);
nand NAND3 (N2895, N2884, N1119, N2346);
not NOT1 (N2896, N2893);
not NOT1 (N2897, N2894);
nor NOR3 (N2898, N2883, N925, N2135);
or OR2 (N2899, N2895, N2356);
nor NOR4 (N2900, N2898, N2068, N473, N1141);
not NOT1 (N2901, N2877);
not NOT1 (N2902, N2890);
xor XOR2 (N2903, N2892, N2124);
and AND2 (N2904, N2903, N1100);
or OR4 (N2905, N2902, N2601, N709, N1948);
not NOT1 (N2906, N2899);
buf BUF1 (N2907, N2905);
nor NOR4 (N2908, N2881, N966, N1297, N273);
nor NOR3 (N2909, N2906, N2373, N969);
not NOT1 (N2910, N2897);
and AND2 (N2911, N2887, N2901);
nor NOR4 (N2912, N1586, N2816, N1409, N657);
buf BUF1 (N2913, N2910);
and AND2 (N2914, N2896, N837);
nor NOR4 (N2915, N2913, N2913, N2642, N958);
xor XOR2 (N2916, N2908, N559);
not NOT1 (N2917, N2900);
xor XOR2 (N2918, N2917, N1064);
or OR4 (N2919, N2911, N586, N2658, N66);
not NOT1 (N2920, N2916);
xor XOR2 (N2921, N2915, N2416);
not NOT1 (N2922, N2904);
buf BUF1 (N2923, N2909);
and AND3 (N2924, N2920, N2379, N594);
nand NAND4 (N2925, N2907, N1682, N330, N759);
not NOT1 (N2926, N2924);
or OR3 (N2927, N2921, N1675, N1587);
and AND3 (N2928, N2927, N1057, N945);
or OR3 (N2929, N2919, N349, N309);
nor NOR2 (N2930, N2929, N1823);
and AND3 (N2931, N2925, N1089, N1686);
buf BUF1 (N2932, N2923);
and AND2 (N2933, N2930, N1057);
nand NAND4 (N2934, N2926, N1896, N478, N2616);
not NOT1 (N2935, N2912);
xor XOR2 (N2936, N2922, N2336);
or OR2 (N2937, N2934, N1125);
and AND2 (N2938, N2936, N2332);
xor XOR2 (N2939, N2931, N2873);
nor NOR2 (N2940, N2935, N1306);
nor NOR3 (N2941, N2933, N1520, N2595);
not NOT1 (N2942, N2939);
nand NAND3 (N2943, N2932, N2211, N2129);
nand NAND4 (N2944, N2918, N1554, N2199, N13);
nor NOR3 (N2945, N2942, N2180, N965);
xor XOR2 (N2946, N2928, N2283);
not NOT1 (N2947, N2945);
or OR3 (N2948, N2943, N2479, N2219);
not NOT1 (N2949, N2947);
and AND4 (N2950, N2940, N2406, N2072, N2043);
not NOT1 (N2951, N2949);
buf BUF1 (N2952, N2937);
not NOT1 (N2953, N2941);
xor XOR2 (N2954, N2951, N2211);
nand NAND3 (N2955, N2952, N892, N630);
xor XOR2 (N2956, N2889, N2349);
nand NAND2 (N2957, N2954, N1402);
xor XOR2 (N2958, N2956, N764);
not NOT1 (N2959, N2948);
buf BUF1 (N2960, N2958);
and AND3 (N2961, N2960, N270, N2438);
and AND2 (N2962, N2946, N942);
nand NAND2 (N2963, N2950, N1601);
not NOT1 (N2964, N2957);
xor XOR2 (N2965, N2959, N1837);
not NOT1 (N2966, N2964);
or OR4 (N2967, N2965, N2331, N1013, N912);
and AND2 (N2968, N2953, N1421);
not NOT1 (N2969, N2961);
or OR2 (N2970, N2966, N518);
buf BUF1 (N2971, N2970);
nor NOR2 (N2972, N2968, N1132);
nand NAND4 (N2973, N2963, N2389, N2468, N522);
and AND3 (N2974, N2914, N1144, N1811);
nand NAND4 (N2975, N2971, N1230, N2672, N1168);
nand NAND2 (N2976, N2944, N690);
or OR4 (N2977, N2975, N2195, N844, N1239);
xor XOR2 (N2978, N2967, N252);
nand NAND2 (N2979, N2972, N1814);
and AND3 (N2980, N2977, N2684, N1221);
buf BUF1 (N2981, N2962);
nor NOR2 (N2982, N2976, N695);
buf BUF1 (N2983, N2955);
not NOT1 (N2984, N2974);
nor NOR3 (N2985, N2979, N2226, N1691);
buf BUF1 (N2986, N2973);
nor NOR4 (N2987, N2969, N435, N2534, N373);
not NOT1 (N2988, N2978);
or OR4 (N2989, N2985, N438, N1087, N1519);
nor NOR3 (N2990, N2986, N228, N800);
xor XOR2 (N2991, N2981, N2491);
nor NOR3 (N2992, N2938, N2828, N1591);
not NOT1 (N2993, N2982);
or OR4 (N2994, N2983, N2405, N1592, N44);
buf BUF1 (N2995, N2980);
nand NAND2 (N2996, N2984, N328);
xor XOR2 (N2997, N2993, N903);
or OR3 (N2998, N2996, N2061, N1828);
nor NOR3 (N2999, N2988, N420, N621);
xor XOR2 (N3000, N2990, N1771);
nand NAND3 (N3001, N2991, N2779, N298);
not NOT1 (N3002, N3001);
nor NOR2 (N3003, N2998, N511);
and AND2 (N3004, N2987, N86);
or OR2 (N3005, N3003, N320);
xor XOR2 (N3006, N3005, N2855);
or OR4 (N3007, N2995, N1438, N916, N1544);
buf BUF1 (N3008, N3006);
not NOT1 (N3009, N3000);
nand NAND4 (N3010, N2997, N222, N1791, N302);
or OR3 (N3011, N3008, N1457, N2507);
xor XOR2 (N3012, N3004, N1480);
nand NAND4 (N3013, N2994, N2802, N1267, N585);
not NOT1 (N3014, N3013);
or OR4 (N3015, N3012, N1445, N2887, N12);
and AND4 (N3016, N3007, N2010, N1368, N1100);
endmodule