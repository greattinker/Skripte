// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15;

output N613,N610,N608,N604,N614,N609,N597,N607,N602,N615;

buf BUF1 (N16, N1);
not NOT1 (N17, N9);
nor NOR2 (N18, N10, N5);
and AND3 (N19, N17, N13, N14);
nor NOR3 (N20, N18, N16, N4);
and AND4 (N21, N8, N15, N11, N4);
and AND2 (N22, N16, N11);
or OR3 (N23, N20, N3, N16);
or OR2 (N24, N15, N5);
nand NAND4 (N25, N10, N4, N5, N10);
nor NOR4 (N26, N22, N5, N2, N11);
buf BUF1 (N27, N1);
buf BUF1 (N28, N20);
or OR3 (N29, N22, N16, N10);
and AND2 (N30, N12, N9);
or OR3 (N31, N27, N27, N16);
not NOT1 (N32, N23);
not NOT1 (N33, N32);
buf BUF1 (N34, N30);
or OR4 (N35, N24, N20, N31, N26);
or OR2 (N36, N13, N33);
xor XOR2 (N37, N25, N11);
not NOT1 (N38, N3);
nor NOR2 (N39, N33, N25);
nor NOR3 (N40, N35, N26, N25);
buf BUF1 (N41, N38);
xor XOR2 (N42, N37, N9);
nand NAND3 (N43, N36, N19, N2);
not NOT1 (N44, N1);
buf BUF1 (N45, N28);
nor NOR2 (N46, N43, N13);
nand NAND4 (N47, N41, N34, N36, N25);
or OR4 (N48, N29, N1, N40, N40);
nor NOR3 (N49, N3, N14, N18);
buf BUF1 (N50, N4);
xor XOR2 (N51, N45, N27);
nand NAND4 (N52, N21, N48, N35, N1);
or OR2 (N53, N27, N9);
nor NOR3 (N54, N53, N28, N46);
or OR2 (N55, N15, N3);
nor NOR3 (N56, N39, N38, N15);
xor XOR2 (N57, N55, N1);
nand NAND4 (N58, N47, N17, N21, N38);
buf BUF1 (N59, N57);
and AND2 (N60, N54, N6);
not NOT1 (N61, N51);
buf BUF1 (N62, N50);
xor XOR2 (N63, N56, N24);
buf BUF1 (N64, N62);
buf BUF1 (N65, N64);
nand NAND2 (N66, N49, N23);
and AND4 (N67, N61, N27, N19, N49);
or OR3 (N68, N60, N4, N1);
nand NAND4 (N69, N58, N60, N64, N45);
nand NAND3 (N70, N52, N43, N44);
nand NAND3 (N71, N70, N67, N26);
or OR2 (N72, N59, N63);
xor XOR2 (N73, N33, N14);
not NOT1 (N74, N20);
xor XOR2 (N75, N67, N33);
nor NOR3 (N76, N73, N3, N40);
not NOT1 (N77, N69);
not NOT1 (N78, N68);
not NOT1 (N79, N72);
xor XOR2 (N80, N78, N60);
xor XOR2 (N81, N71, N26);
or OR4 (N82, N42, N47, N55, N69);
or OR4 (N83, N74, N14, N46, N4);
and AND3 (N84, N80, N51, N82);
buf BUF1 (N85, N45);
xor XOR2 (N86, N66, N81);
or OR3 (N87, N10, N54, N69);
nand NAND4 (N88, N85, N69, N30, N58);
not NOT1 (N89, N75);
nor NOR4 (N90, N79, N46, N26, N47);
buf BUF1 (N91, N87);
nand NAND3 (N92, N77, N26, N84);
and AND2 (N93, N64, N48);
buf BUF1 (N94, N65);
xor XOR2 (N95, N86, N80);
nand NAND4 (N96, N93, N57, N92, N56);
and AND2 (N97, N72, N48);
or OR3 (N98, N91, N16, N54);
and AND4 (N99, N98, N95, N29, N43);
buf BUF1 (N100, N80);
xor XOR2 (N101, N94, N4);
not NOT1 (N102, N89);
nand NAND2 (N103, N101, N72);
not NOT1 (N104, N90);
and AND3 (N105, N97, N97, N83);
nand NAND3 (N106, N81, N81, N89);
xor XOR2 (N107, N103, N54);
buf BUF1 (N108, N76);
not NOT1 (N109, N102);
not NOT1 (N110, N96);
or OR3 (N111, N107, N31, N79);
buf BUF1 (N112, N109);
nand NAND3 (N113, N110, N43, N21);
and AND2 (N114, N108, N57);
not NOT1 (N115, N106);
nand NAND3 (N116, N100, N7, N7);
xor XOR2 (N117, N88, N81);
or OR3 (N118, N104, N11, N32);
or OR3 (N119, N115, N23, N102);
nand NAND4 (N120, N113, N51, N87, N13);
xor XOR2 (N121, N118, N5);
buf BUF1 (N122, N121);
or OR4 (N123, N114, N25, N6, N41);
buf BUF1 (N124, N112);
not NOT1 (N125, N123);
and AND4 (N126, N117, N117, N32, N17);
not NOT1 (N127, N125);
or OR3 (N128, N111, N19, N95);
and AND4 (N129, N124, N48, N34, N37);
or OR4 (N130, N128, N108, N27, N66);
nand NAND2 (N131, N116, N80);
nand NAND2 (N132, N130, N106);
xor XOR2 (N133, N105, N122);
nor NOR2 (N134, N78, N119);
or OR2 (N135, N67, N129);
nor NOR3 (N136, N16, N31, N16);
buf BUF1 (N137, N133);
or OR3 (N138, N134, N81, N69);
or OR2 (N139, N135, N69);
and AND3 (N140, N120, N71, N106);
not NOT1 (N141, N138);
nor NOR2 (N142, N126, N35);
and AND4 (N143, N132, N14, N15, N60);
not NOT1 (N144, N140);
buf BUF1 (N145, N141);
or OR2 (N146, N131, N31);
xor XOR2 (N147, N127, N104);
nor NOR2 (N148, N145, N78);
or OR3 (N149, N147, N40, N4);
nor NOR4 (N150, N149, N54, N137, N127);
nor NOR4 (N151, N83, N33, N31, N60);
or OR2 (N152, N148, N106);
xor XOR2 (N153, N136, N128);
xor XOR2 (N154, N146, N109);
nand NAND3 (N155, N152, N29, N101);
or OR2 (N156, N155, N125);
buf BUF1 (N157, N150);
or OR4 (N158, N156, N29, N6, N102);
xor XOR2 (N159, N143, N133);
nor NOR4 (N160, N139, N145, N145, N92);
not NOT1 (N161, N160);
buf BUF1 (N162, N99);
not NOT1 (N163, N151);
nand NAND2 (N164, N157, N15);
and AND4 (N165, N154, N83, N159, N91);
or OR4 (N166, N22, N42, N128, N150);
and AND2 (N167, N158, N131);
nor NOR3 (N168, N163, N124, N29);
nor NOR2 (N169, N168, N123);
xor XOR2 (N170, N169, N35);
not NOT1 (N171, N161);
nor NOR3 (N172, N171, N90, N70);
xor XOR2 (N173, N142, N126);
and AND2 (N174, N164, N68);
nor NOR4 (N175, N166, N5, N147, N84);
and AND4 (N176, N162, N165, N122, N151);
xor XOR2 (N177, N88, N60);
and AND2 (N178, N170, N25);
nor NOR3 (N179, N178, N95, N95);
nand NAND4 (N180, N167, N68, N9, N20);
or OR2 (N181, N174, N15);
nand NAND4 (N182, N180, N169, N23, N75);
nand NAND2 (N183, N176, N62);
buf BUF1 (N184, N175);
and AND2 (N185, N172, N81);
nand NAND4 (N186, N173, N42, N1, N150);
buf BUF1 (N187, N153);
not NOT1 (N188, N186);
xor XOR2 (N189, N177, N123);
not NOT1 (N190, N188);
and AND2 (N191, N184, N10);
not NOT1 (N192, N183);
xor XOR2 (N193, N187, N173);
and AND2 (N194, N185, N12);
xor XOR2 (N195, N182, N181);
xor XOR2 (N196, N53, N119);
buf BUF1 (N197, N189);
buf BUF1 (N198, N144);
or OR4 (N199, N190, N144, N81, N195);
and AND3 (N200, N52, N8, N52);
or OR2 (N201, N191, N145);
nand NAND4 (N202, N179, N155, N101, N164);
not NOT1 (N203, N199);
and AND4 (N204, N200, N183, N90, N183);
nor NOR3 (N205, N197, N202, N159);
xor XOR2 (N206, N46, N98);
xor XOR2 (N207, N205, N138);
not NOT1 (N208, N193);
not NOT1 (N209, N192);
xor XOR2 (N210, N208, N133);
not NOT1 (N211, N198);
or OR2 (N212, N210, N77);
buf BUF1 (N213, N211);
buf BUF1 (N214, N206);
not NOT1 (N215, N196);
buf BUF1 (N216, N212);
xor XOR2 (N217, N207, N157);
buf BUF1 (N218, N214);
buf BUF1 (N219, N203);
or OR4 (N220, N204, N156, N70, N1);
or OR3 (N221, N216, N63, N171);
and AND4 (N222, N194, N180, N128, N214);
xor XOR2 (N223, N213, N29);
or OR2 (N224, N220, N72);
xor XOR2 (N225, N219, N68);
buf BUF1 (N226, N221);
not NOT1 (N227, N215);
nand NAND4 (N228, N209, N152, N123, N31);
nand NAND4 (N229, N225, N14, N211, N111);
and AND2 (N230, N228, N134);
nand NAND4 (N231, N227, N41, N112, N59);
or OR2 (N232, N222, N212);
nor NOR3 (N233, N224, N7, N186);
or OR2 (N234, N201, N44);
buf BUF1 (N235, N230);
nand NAND4 (N236, N218, N229, N216, N224);
and AND2 (N237, N13, N96);
buf BUF1 (N238, N231);
nand NAND4 (N239, N232, N139, N204, N109);
not NOT1 (N240, N239);
xor XOR2 (N241, N240, N132);
or OR4 (N242, N223, N158, N7, N193);
not NOT1 (N243, N241);
nand NAND3 (N244, N217, N150, N184);
and AND4 (N245, N226, N72, N239, N198);
and AND2 (N246, N236, N126);
or OR3 (N247, N245, N176, N185);
or OR2 (N248, N244, N93);
xor XOR2 (N249, N237, N84);
nor NOR3 (N250, N249, N160, N216);
and AND2 (N251, N246, N68);
nor NOR4 (N252, N242, N95, N101, N224);
xor XOR2 (N253, N250, N56);
or OR4 (N254, N252, N147, N96, N178);
or OR4 (N255, N251, N163, N212, N217);
xor XOR2 (N256, N247, N109);
not NOT1 (N257, N256);
xor XOR2 (N258, N257, N56);
not NOT1 (N259, N235);
xor XOR2 (N260, N254, N89);
nor NOR2 (N261, N233, N229);
or OR4 (N262, N253, N83, N159, N233);
or OR4 (N263, N255, N256, N158, N243);
nor NOR4 (N264, N218, N134, N171, N133);
xor XOR2 (N265, N234, N105);
nand NAND4 (N266, N263, N34, N92, N240);
or OR4 (N267, N259, N113, N81, N105);
xor XOR2 (N268, N262, N203);
not NOT1 (N269, N260);
and AND3 (N270, N268, N260, N66);
and AND3 (N271, N266, N110, N255);
or OR2 (N272, N269, N113);
xor XOR2 (N273, N272, N111);
buf BUF1 (N274, N265);
or OR2 (N275, N274, N14);
nor NOR4 (N276, N264, N12, N25, N180);
buf BUF1 (N277, N270);
xor XOR2 (N278, N273, N227);
or OR3 (N279, N278, N221, N268);
nor NOR3 (N280, N238, N269, N205);
nand NAND3 (N281, N279, N43, N243);
xor XOR2 (N282, N276, N204);
nor NOR2 (N283, N280, N146);
and AND4 (N284, N275, N270, N78, N97);
and AND4 (N285, N282, N227, N196, N65);
nand NAND2 (N286, N261, N160);
xor XOR2 (N287, N248, N253);
or OR3 (N288, N286, N53, N280);
xor XOR2 (N289, N284, N275);
nand NAND4 (N290, N258, N99, N169, N83);
not NOT1 (N291, N285);
not NOT1 (N292, N290);
not NOT1 (N293, N271);
buf BUF1 (N294, N287);
nand NAND3 (N295, N292, N74, N101);
or OR2 (N296, N293, N70);
buf BUF1 (N297, N281);
or OR3 (N298, N297, N176, N171);
xor XOR2 (N299, N289, N10);
nor NOR2 (N300, N288, N157);
not NOT1 (N301, N267);
not NOT1 (N302, N294);
buf BUF1 (N303, N300);
nor NOR2 (N304, N299, N122);
buf BUF1 (N305, N296);
xor XOR2 (N306, N295, N234);
or OR2 (N307, N306, N196);
not NOT1 (N308, N303);
buf BUF1 (N309, N301);
buf BUF1 (N310, N291);
xor XOR2 (N311, N309, N99);
not NOT1 (N312, N305);
or OR3 (N313, N304, N168, N153);
nand NAND3 (N314, N277, N260, N22);
nand NAND3 (N315, N298, N195, N14);
buf BUF1 (N316, N307);
not NOT1 (N317, N311);
xor XOR2 (N318, N283, N1);
nand NAND4 (N319, N314, N162, N187, N192);
not NOT1 (N320, N319);
xor XOR2 (N321, N317, N43);
xor XOR2 (N322, N318, N87);
nor NOR4 (N323, N313, N46, N162, N322);
buf BUF1 (N324, N122);
nand NAND2 (N325, N316, N60);
or OR2 (N326, N312, N171);
nor NOR3 (N327, N321, N20, N286);
nand NAND4 (N328, N324, N56, N54, N150);
xor XOR2 (N329, N315, N12);
nor NOR4 (N330, N302, N212, N147, N16);
nand NAND4 (N331, N320, N147, N185, N274);
or OR4 (N332, N330, N250, N309, N100);
or OR2 (N333, N329, N255);
nor NOR2 (N334, N332, N170);
buf BUF1 (N335, N327);
xor XOR2 (N336, N334, N293);
or OR3 (N337, N333, N237, N322);
xor XOR2 (N338, N326, N166);
or OR3 (N339, N325, N113, N215);
and AND2 (N340, N308, N168);
not NOT1 (N341, N331);
nor NOR4 (N342, N328, N280, N92, N23);
or OR2 (N343, N337, N177);
or OR2 (N344, N342, N31);
buf BUF1 (N345, N338);
and AND4 (N346, N339, N127, N234, N31);
not NOT1 (N347, N335);
nor NOR2 (N348, N310, N14);
nor NOR4 (N349, N348, N333, N97, N160);
not NOT1 (N350, N336);
not NOT1 (N351, N343);
nand NAND4 (N352, N350, N64, N48, N167);
or OR3 (N353, N349, N96, N275);
xor XOR2 (N354, N346, N209);
not NOT1 (N355, N351);
xor XOR2 (N356, N344, N308);
nand NAND4 (N357, N356, N5, N57, N335);
not NOT1 (N358, N353);
nand NAND2 (N359, N355, N177);
nand NAND2 (N360, N345, N53);
nand NAND2 (N361, N347, N35);
xor XOR2 (N362, N359, N155);
buf BUF1 (N363, N340);
nand NAND3 (N364, N323, N188, N133);
buf BUF1 (N365, N364);
xor XOR2 (N366, N352, N133);
or OR3 (N367, N361, N330, N194);
buf BUF1 (N368, N366);
nor NOR4 (N369, N363, N130, N318, N120);
xor XOR2 (N370, N365, N93);
xor XOR2 (N371, N341, N104);
not NOT1 (N372, N370);
xor XOR2 (N373, N372, N334);
xor XOR2 (N374, N369, N261);
buf BUF1 (N375, N374);
and AND3 (N376, N373, N165, N286);
or OR4 (N377, N376, N374, N376, N261);
nor NOR3 (N378, N362, N117, N312);
not NOT1 (N379, N358);
xor XOR2 (N380, N371, N328);
nand NAND3 (N381, N377, N156, N78);
buf BUF1 (N382, N375);
buf BUF1 (N383, N354);
not NOT1 (N384, N382);
xor XOR2 (N385, N368, N179);
or OR4 (N386, N381, N329, N133, N364);
xor XOR2 (N387, N378, N156);
or OR3 (N388, N379, N263, N204);
buf BUF1 (N389, N360);
buf BUF1 (N390, N387);
and AND3 (N391, N383, N69, N299);
buf BUF1 (N392, N388);
or OR3 (N393, N386, N224, N204);
nor NOR4 (N394, N393, N368, N284, N115);
buf BUF1 (N395, N385);
or OR4 (N396, N390, N39, N128, N107);
or OR4 (N397, N357, N35, N391, N265);
xor XOR2 (N398, N82, N188);
and AND2 (N399, N367, N300);
and AND3 (N400, N395, N295, N142);
nor NOR2 (N401, N380, N205);
and AND3 (N402, N389, N183, N163);
buf BUF1 (N403, N401);
buf BUF1 (N404, N403);
and AND2 (N405, N402, N80);
not NOT1 (N406, N397);
and AND3 (N407, N405, N22, N261);
and AND4 (N408, N394, N213, N137, N381);
and AND4 (N409, N404, N212, N174, N36);
nand NAND3 (N410, N409, N108, N69);
or OR3 (N411, N410, N222, N6);
nand NAND3 (N412, N406, N1, N148);
and AND3 (N413, N399, N412, N82);
or OR2 (N414, N60, N173);
buf BUF1 (N415, N413);
and AND2 (N416, N392, N307);
xor XOR2 (N417, N411, N37);
nand NAND4 (N418, N417, N349, N13, N406);
nand NAND2 (N419, N407, N38);
xor XOR2 (N420, N419, N359);
not NOT1 (N421, N415);
buf BUF1 (N422, N408);
buf BUF1 (N423, N384);
buf BUF1 (N424, N418);
xor XOR2 (N425, N416, N174);
buf BUF1 (N426, N422);
xor XOR2 (N427, N396, N425);
not NOT1 (N428, N388);
nor NOR4 (N429, N400, N373, N41, N22);
or OR2 (N430, N424, N147);
nor NOR2 (N431, N430, N309);
xor XOR2 (N432, N429, N349);
or OR3 (N433, N421, N150, N66);
nor NOR3 (N434, N427, N180, N322);
not NOT1 (N435, N428);
nor NOR2 (N436, N398, N361);
xor XOR2 (N437, N423, N203);
or OR3 (N438, N431, N68, N204);
xor XOR2 (N439, N434, N72);
buf BUF1 (N440, N435);
nor NOR3 (N441, N436, N122, N270);
or OR4 (N442, N420, N287, N263, N439);
xor XOR2 (N443, N30, N352);
nand NAND4 (N444, N414, N148, N129, N380);
and AND3 (N445, N433, N183, N392);
or OR2 (N446, N440, N274);
and AND3 (N447, N438, N2, N283);
or OR2 (N448, N445, N328);
or OR3 (N449, N432, N448, N252);
nand NAND4 (N450, N118, N402, N77, N95);
xor XOR2 (N451, N446, N315);
or OR3 (N452, N447, N72, N369);
nand NAND4 (N453, N437, N448, N246, N323);
xor XOR2 (N454, N451, N365);
and AND4 (N455, N443, N20, N22, N156);
or OR2 (N456, N441, N182);
and AND4 (N457, N449, N226, N81, N80);
buf BUF1 (N458, N444);
nand NAND4 (N459, N442, N95, N52, N159);
and AND3 (N460, N452, N165, N190);
or OR4 (N461, N456, N296, N232, N181);
xor XOR2 (N462, N453, N170);
buf BUF1 (N463, N462);
xor XOR2 (N464, N460, N186);
not NOT1 (N465, N454);
buf BUF1 (N466, N461);
nor NOR2 (N467, N450, N106);
xor XOR2 (N468, N463, N290);
nor NOR4 (N469, N459, N449, N250, N170);
nand NAND2 (N470, N457, N115);
buf BUF1 (N471, N470);
or OR2 (N472, N466, N274);
or OR3 (N473, N467, N17, N272);
or OR4 (N474, N465, N250, N146, N294);
nand NAND4 (N475, N473, N296, N75, N205);
xor XOR2 (N476, N475, N293);
xor XOR2 (N477, N472, N15);
xor XOR2 (N478, N476, N125);
buf BUF1 (N479, N455);
not NOT1 (N480, N478);
not NOT1 (N481, N474);
nand NAND4 (N482, N479, N364, N111, N458);
xor XOR2 (N483, N242, N414);
xor XOR2 (N484, N471, N186);
not NOT1 (N485, N480);
nor NOR3 (N486, N481, N229, N333);
nand NAND2 (N487, N477, N31);
xor XOR2 (N488, N468, N230);
xor XOR2 (N489, N483, N458);
buf BUF1 (N490, N482);
nor NOR2 (N491, N426, N442);
not NOT1 (N492, N489);
and AND4 (N493, N484, N230, N325, N365);
buf BUF1 (N494, N486);
buf BUF1 (N495, N469);
not NOT1 (N496, N487);
nand NAND4 (N497, N464, N451, N431, N298);
xor XOR2 (N498, N496, N201);
nor NOR2 (N499, N494, N145);
or OR4 (N500, N488, N68, N432, N8);
xor XOR2 (N501, N498, N324);
nor NOR2 (N502, N500, N285);
buf BUF1 (N503, N497);
buf BUF1 (N504, N495);
or OR2 (N505, N499, N72);
nand NAND4 (N506, N491, N471, N254, N275);
nand NAND3 (N507, N505, N438, N487);
nand NAND2 (N508, N503, N327);
or OR3 (N509, N507, N403, N121);
nor NOR2 (N510, N504, N79);
buf BUF1 (N511, N508);
nand NAND2 (N512, N501, N492);
nand NAND3 (N513, N109, N140, N412);
nand NAND4 (N514, N493, N428, N269, N444);
not NOT1 (N515, N511);
nand NAND2 (N516, N485, N96);
buf BUF1 (N517, N490);
xor XOR2 (N518, N509, N142);
and AND4 (N519, N510, N75, N82, N124);
nand NAND2 (N520, N513, N496);
and AND2 (N521, N519, N240);
nand NAND3 (N522, N516, N505, N367);
nor NOR2 (N523, N518, N290);
nand NAND4 (N524, N517, N409, N325, N490);
xor XOR2 (N525, N523, N473);
xor XOR2 (N526, N520, N407);
nand NAND4 (N527, N502, N300, N236, N234);
nand NAND4 (N528, N524, N463, N284, N143);
or OR4 (N529, N512, N358, N377, N320);
buf BUF1 (N530, N526);
buf BUF1 (N531, N506);
nor NOR3 (N532, N529, N424, N210);
nand NAND2 (N533, N514, N399);
xor XOR2 (N534, N528, N161);
not NOT1 (N535, N533);
nor NOR3 (N536, N522, N237, N524);
buf BUF1 (N537, N515);
or OR3 (N538, N530, N229, N194);
or OR3 (N539, N532, N261, N511);
xor XOR2 (N540, N535, N214);
buf BUF1 (N541, N538);
not NOT1 (N542, N525);
or OR2 (N543, N537, N511);
or OR2 (N544, N527, N496);
or OR2 (N545, N540, N526);
nor NOR4 (N546, N542, N35, N427, N483);
or OR2 (N547, N541, N255);
not NOT1 (N548, N521);
nor NOR4 (N549, N548, N328, N251, N208);
or OR4 (N550, N543, N64, N323, N372);
nand NAND4 (N551, N550, N203, N341, N308);
xor XOR2 (N552, N546, N37);
nor NOR4 (N553, N545, N402, N435, N111);
xor XOR2 (N554, N536, N335);
and AND4 (N555, N551, N155, N139, N16);
buf BUF1 (N556, N531);
not NOT1 (N557, N534);
nor NOR2 (N558, N539, N56);
nor NOR3 (N559, N555, N143, N308);
not NOT1 (N560, N558);
and AND3 (N561, N557, N347, N66);
xor XOR2 (N562, N552, N455);
and AND2 (N563, N549, N235);
nor NOR4 (N564, N544, N479, N560, N399);
xor XOR2 (N565, N520, N533);
buf BUF1 (N566, N563);
and AND3 (N567, N547, N267, N522);
nand NAND3 (N568, N565, N161, N385);
and AND2 (N569, N561, N28);
nor NOR3 (N570, N562, N569, N342);
xor XOR2 (N571, N16, N182);
or OR4 (N572, N559, N455, N179, N119);
and AND2 (N573, N572, N449);
buf BUF1 (N574, N570);
xor XOR2 (N575, N574, N560);
xor XOR2 (N576, N571, N172);
buf BUF1 (N577, N566);
nand NAND4 (N578, N568, N551, N219, N358);
nand NAND2 (N579, N573, N319);
and AND3 (N580, N576, N346, N477);
xor XOR2 (N581, N564, N361);
xor XOR2 (N582, N581, N196);
nor NOR3 (N583, N554, N18, N486);
nand NAND3 (N584, N579, N238, N259);
or OR4 (N585, N578, N139, N28, N414);
nor NOR2 (N586, N580, N164);
nand NAND4 (N587, N582, N539, N331, N172);
nand NAND3 (N588, N585, N156, N420);
or OR4 (N589, N577, N445, N114, N154);
nor NOR3 (N590, N567, N158, N45);
not NOT1 (N591, N583);
nor NOR3 (N592, N591, N532, N4);
xor XOR2 (N593, N586, N70);
nand NAND3 (N594, N575, N328, N356);
nand NAND3 (N595, N588, N36, N586);
nor NOR4 (N596, N595, N526, N524, N393);
xor XOR2 (N597, N553, N477);
xor XOR2 (N598, N590, N35);
nor NOR3 (N599, N592, N51, N496);
xor XOR2 (N600, N589, N131);
not NOT1 (N601, N593);
and AND4 (N602, N601, N98, N167, N557);
and AND2 (N603, N584, N497);
not NOT1 (N604, N598);
nor NOR3 (N605, N594, N499, N519);
buf BUF1 (N606, N587);
nand NAND3 (N607, N599, N398, N435);
nand NAND4 (N608, N596, N106, N228, N75);
xor XOR2 (N609, N556, N96);
not NOT1 (N610, N600);
nor NOR2 (N611, N603, N541);
or OR3 (N612, N606, N472, N533);
and AND4 (N613, N605, N37, N543, N13);
buf BUF1 (N614, N612);
nor NOR3 (N615, N611, N28, N517);
endmodule