// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22;

output N3516,N3518,N3514,N3520,N3511,N3519,N3483,N3521,N3515,N3522;

buf BUF1 (N23, N19);
nor NOR4 (N24, N4, N10, N6, N8);
nand NAND4 (N25, N4, N24, N19, N11);
and AND4 (N26, N16, N8, N6, N20);
xor XOR2 (N27, N10, N14);
buf BUF1 (N28, N9);
nand NAND4 (N29, N23, N3, N24, N11);
xor XOR2 (N30, N23, N24);
not NOT1 (N31, N20);
nor NOR2 (N32, N19, N17);
and AND3 (N33, N4, N4, N9);
xor XOR2 (N34, N27, N18);
nor NOR3 (N35, N22, N18, N19);
nand NAND2 (N36, N25, N16);
and AND3 (N37, N26, N17, N24);
nor NOR4 (N38, N28, N34, N14, N19);
and AND4 (N39, N4, N35, N16, N14);
xor XOR2 (N40, N4, N33);
and AND2 (N41, N24, N18);
nand NAND2 (N42, N37, N28);
xor XOR2 (N43, N36, N7);
nor NOR2 (N44, N40, N26);
nor NOR2 (N45, N44, N4);
and AND4 (N46, N32, N45, N31, N40);
not NOT1 (N47, N43);
nor NOR4 (N48, N28, N2, N32, N18);
or OR2 (N49, N9, N6);
xor XOR2 (N50, N39, N31);
not NOT1 (N51, N47);
not NOT1 (N52, N48);
xor XOR2 (N53, N46, N5);
nor NOR4 (N54, N38, N53, N50, N2);
nand NAND3 (N55, N6, N18, N45);
xor XOR2 (N56, N52, N47);
nor NOR4 (N57, N6, N6, N28, N44);
buf BUF1 (N58, N57);
and AND3 (N59, N49, N4, N17);
and AND3 (N60, N54, N13, N1);
or OR2 (N61, N56, N40);
buf BUF1 (N62, N61);
and AND2 (N63, N30, N32);
buf BUF1 (N64, N62);
nand NAND3 (N65, N29, N14, N55);
or OR2 (N66, N60, N13);
xor XOR2 (N67, N49, N45);
nand NAND3 (N68, N59, N41, N4);
xor XOR2 (N69, N9, N50);
xor XOR2 (N70, N42, N29);
buf BUF1 (N71, N70);
and AND2 (N72, N64, N13);
xor XOR2 (N73, N51, N49);
nor NOR3 (N74, N69, N34, N61);
nand NAND4 (N75, N68, N36, N34, N16);
or OR3 (N76, N71, N19, N47);
xor XOR2 (N77, N72, N2);
not NOT1 (N78, N65);
nand NAND2 (N79, N58, N39);
or OR3 (N80, N76, N73, N7);
nor NOR4 (N81, N22, N10, N26, N74);
buf BUF1 (N82, N8);
and AND3 (N83, N77, N63, N21);
not NOT1 (N84, N1);
not NOT1 (N85, N83);
not NOT1 (N86, N67);
xor XOR2 (N87, N86, N21);
or OR3 (N88, N75, N52, N85);
nor NOR2 (N89, N22, N78);
xor XOR2 (N90, N59, N70);
buf BUF1 (N91, N80);
or OR2 (N92, N66, N72);
xor XOR2 (N93, N87, N31);
xor XOR2 (N94, N88, N90);
nand NAND2 (N95, N39, N94);
nand NAND3 (N96, N51, N9, N42);
nand NAND4 (N97, N95, N25, N1, N12);
nor NOR3 (N98, N92, N55, N29);
and AND4 (N99, N82, N14, N4, N45);
nor NOR3 (N100, N81, N94, N59);
or OR3 (N101, N93, N95, N71);
buf BUF1 (N102, N100);
or OR4 (N103, N91, N40, N47, N32);
nor NOR4 (N104, N97, N20, N8, N85);
nor NOR4 (N105, N96, N50, N64, N96);
nor NOR2 (N106, N101, N93);
buf BUF1 (N107, N102);
buf BUF1 (N108, N98);
or OR2 (N109, N79, N42);
buf BUF1 (N110, N106);
or OR4 (N111, N89, N26, N101, N60);
and AND3 (N112, N103, N63, N21);
nor NOR3 (N113, N104, N55, N95);
or OR4 (N114, N110, N11, N75, N17);
buf BUF1 (N115, N99);
buf BUF1 (N116, N111);
not NOT1 (N117, N112);
nand NAND4 (N118, N109, N74, N14, N79);
nor NOR2 (N119, N118, N35);
and AND4 (N120, N114, N93, N95, N85);
not NOT1 (N121, N84);
nand NAND4 (N122, N105, N37, N62, N88);
nor NOR3 (N123, N116, N73, N12);
nand NAND4 (N124, N119, N92, N25, N102);
xor XOR2 (N125, N122, N54);
or OR4 (N126, N117, N71, N70, N68);
not NOT1 (N127, N125);
buf BUF1 (N128, N107);
xor XOR2 (N129, N128, N95);
buf BUF1 (N130, N129);
or OR2 (N131, N121, N19);
nor NOR4 (N132, N126, N1, N57, N78);
buf BUF1 (N133, N108);
nor NOR3 (N134, N127, N124, N120);
nor NOR3 (N135, N129, N132, N88);
xor XOR2 (N136, N66, N93);
not NOT1 (N137, N72);
not NOT1 (N138, N134);
nand NAND2 (N139, N113, N137);
and AND4 (N140, N81, N34, N75, N84);
nor NOR2 (N141, N140, N129);
nand NAND2 (N142, N141, N33);
buf BUF1 (N143, N135);
buf BUF1 (N144, N143);
nor NOR2 (N145, N144, N88);
and AND3 (N146, N136, N111, N83);
nor NOR2 (N147, N138, N5);
nand NAND4 (N148, N146, N13, N109, N144);
buf BUF1 (N149, N123);
buf BUF1 (N150, N149);
xor XOR2 (N151, N150, N40);
or OR4 (N152, N133, N75, N17, N2);
not NOT1 (N153, N139);
nand NAND4 (N154, N115, N77, N136, N139);
xor XOR2 (N155, N142, N31);
nand NAND4 (N156, N147, N125, N141, N57);
or OR3 (N157, N148, N79, N134);
and AND4 (N158, N153, N47, N126, N61);
or OR4 (N159, N130, N128, N150, N157);
and AND3 (N160, N132, N39, N71);
or OR4 (N161, N155, N44, N76, N67);
and AND3 (N162, N154, N99, N80);
not NOT1 (N163, N160);
and AND4 (N164, N163, N112, N52, N69);
nor NOR4 (N165, N151, N140, N20, N25);
nor NOR3 (N166, N158, N10, N111);
xor XOR2 (N167, N156, N73);
and AND2 (N168, N145, N119);
not NOT1 (N169, N152);
xor XOR2 (N170, N159, N152);
buf BUF1 (N171, N167);
buf BUF1 (N172, N169);
or OR4 (N173, N172, N128, N129, N126);
or OR3 (N174, N161, N76, N144);
buf BUF1 (N175, N173);
buf BUF1 (N176, N164);
and AND3 (N177, N162, N113, N53);
buf BUF1 (N178, N168);
not NOT1 (N179, N131);
or OR3 (N180, N175, N148, N30);
not NOT1 (N181, N166);
nand NAND2 (N182, N179, N77);
nor NOR4 (N183, N170, N106, N86, N96);
nor NOR3 (N184, N174, N17, N48);
nand NAND2 (N185, N178, N31);
nor NOR3 (N186, N181, N101, N25);
nand NAND4 (N187, N177, N147, N125, N64);
or OR3 (N188, N185, N110, N59);
and AND3 (N189, N183, N81, N24);
not NOT1 (N190, N187);
not NOT1 (N191, N188);
xor XOR2 (N192, N182, N147);
not NOT1 (N193, N165);
buf BUF1 (N194, N171);
nor NOR4 (N195, N193, N188, N61, N181);
nand NAND3 (N196, N191, N15, N129);
nand NAND2 (N197, N194, N70);
not NOT1 (N198, N196);
not NOT1 (N199, N186);
nor NOR3 (N200, N195, N90, N39);
nand NAND4 (N201, N192, N81, N166, N75);
buf BUF1 (N202, N200);
nand NAND2 (N203, N197, N164);
xor XOR2 (N204, N184, N159);
xor XOR2 (N205, N189, N111);
nor NOR4 (N206, N205, N110, N155, N199);
nor NOR2 (N207, N67, N193);
buf BUF1 (N208, N201);
nor NOR4 (N209, N207, N135, N47, N204);
xor XOR2 (N210, N78, N30);
xor XOR2 (N211, N190, N86);
or OR3 (N212, N202, N72, N98);
not NOT1 (N213, N206);
nor NOR2 (N214, N203, N183);
xor XOR2 (N215, N214, N64);
nor NOR4 (N216, N180, N143, N178, N43);
nand NAND2 (N217, N208, N181);
or OR3 (N218, N213, N64, N164);
xor XOR2 (N219, N209, N192);
and AND2 (N220, N211, N45);
not NOT1 (N221, N215);
nor NOR4 (N222, N210, N177, N33, N56);
or OR3 (N223, N217, N193, N77);
or OR2 (N224, N218, N140);
buf BUF1 (N225, N222);
nor NOR4 (N226, N224, N42, N101, N41);
and AND3 (N227, N221, N130, N188);
or OR2 (N228, N220, N28);
and AND2 (N229, N198, N13);
or OR4 (N230, N212, N2, N117, N18);
and AND4 (N231, N227, N145, N83, N188);
not NOT1 (N232, N230);
or OR3 (N233, N219, N178, N89);
nor NOR2 (N234, N228, N102);
or OR4 (N235, N231, N130, N43, N125);
nand NAND3 (N236, N229, N97, N122);
and AND3 (N237, N236, N142, N96);
nor NOR2 (N238, N237, N58);
not NOT1 (N239, N176);
nor NOR3 (N240, N239, N206, N228);
and AND3 (N241, N225, N104, N26);
nand NAND4 (N242, N232, N220, N213, N132);
buf BUF1 (N243, N238);
and AND2 (N244, N243, N127);
buf BUF1 (N245, N235);
not NOT1 (N246, N242);
and AND2 (N247, N246, N197);
not NOT1 (N248, N240);
nand NAND4 (N249, N226, N191, N146, N248);
xor XOR2 (N250, N212, N42);
xor XOR2 (N251, N241, N133);
not NOT1 (N252, N249);
and AND2 (N253, N252, N45);
not NOT1 (N254, N216);
nor NOR4 (N255, N254, N122, N207, N6);
xor XOR2 (N256, N223, N26);
not NOT1 (N257, N245);
buf BUF1 (N258, N251);
nand NAND3 (N259, N257, N106, N185);
nand NAND3 (N260, N256, N194, N7);
or OR4 (N261, N234, N88, N214, N65);
and AND4 (N262, N250, N125, N252, N10);
nor NOR2 (N263, N261, N111);
buf BUF1 (N264, N255);
nand NAND3 (N265, N253, N143, N85);
not NOT1 (N266, N244);
and AND3 (N267, N247, N197, N228);
nor NOR3 (N268, N259, N196, N252);
xor XOR2 (N269, N233, N259);
not NOT1 (N270, N264);
nor NOR2 (N271, N262, N94);
or OR3 (N272, N268, N95, N52);
and AND3 (N273, N272, N271, N225);
or OR4 (N274, N35, N46, N142, N116);
and AND3 (N275, N267, N66, N274);
nand NAND2 (N276, N188, N51);
nor NOR4 (N277, N275, N113, N113, N105);
and AND2 (N278, N277, N262);
not NOT1 (N279, N258);
not NOT1 (N280, N260);
or OR4 (N281, N278, N209, N103, N227);
nand NAND2 (N282, N269, N210);
nand NAND4 (N283, N281, N22, N54, N133);
and AND3 (N284, N282, N51, N98);
xor XOR2 (N285, N276, N15);
or OR2 (N286, N265, N279);
and AND3 (N287, N253, N206, N245);
xor XOR2 (N288, N273, N2);
and AND4 (N289, N285, N147, N35, N21);
or OR2 (N290, N287, N37);
not NOT1 (N291, N289);
buf BUF1 (N292, N283);
nand NAND3 (N293, N280, N204, N69);
and AND2 (N294, N291, N7);
nor NOR3 (N295, N288, N280, N236);
buf BUF1 (N296, N292);
nor NOR2 (N297, N270, N2);
xor XOR2 (N298, N263, N22);
xor XOR2 (N299, N284, N282);
xor XOR2 (N300, N286, N299);
and AND4 (N301, N170, N95, N104, N85);
and AND2 (N302, N297, N242);
buf BUF1 (N303, N302);
or OR4 (N304, N296, N19, N213, N59);
xor XOR2 (N305, N301, N221);
or OR2 (N306, N305, N244);
buf BUF1 (N307, N295);
or OR4 (N308, N307, N198, N302, N147);
nand NAND4 (N309, N293, N138, N162, N161);
buf BUF1 (N310, N303);
nor NOR2 (N311, N308, N219);
and AND4 (N312, N300, N42, N12, N32);
not NOT1 (N313, N266);
xor XOR2 (N314, N311, N42);
not NOT1 (N315, N290);
xor XOR2 (N316, N312, N37);
xor XOR2 (N317, N313, N56);
buf BUF1 (N318, N304);
nor NOR2 (N319, N315, N202);
nor NOR3 (N320, N319, N194, N308);
buf BUF1 (N321, N317);
buf BUF1 (N322, N321);
nand NAND2 (N323, N294, N310);
buf BUF1 (N324, N137);
or OR3 (N325, N322, N11, N262);
xor XOR2 (N326, N320, N144);
nor NOR3 (N327, N306, N320, N228);
or OR3 (N328, N318, N134, N54);
and AND4 (N329, N325, N212, N48, N221);
nor NOR4 (N330, N327, N83, N102, N320);
xor XOR2 (N331, N324, N138);
not NOT1 (N332, N298);
nor NOR4 (N333, N328, N134, N254, N72);
buf BUF1 (N334, N331);
and AND4 (N335, N330, N125, N34, N178);
not NOT1 (N336, N316);
and AND3 (N337, N333, N28, N302);
xor XOR2 (N338, N323, N41);
nand NAND4 (N339, N335, N13, N234, N131);
nor NOR3 (N340, N309, N262, N278);
and AND4 (N341, N337, N40, N1, N253);
and AND3 (N342, N339, N187, N167);
xor XOR2 (N343, N341, N17);
buf BUF1 (N344, N336);
and AND3 (N345, N334, N337, N201);
nand NAND2 (N346, N329, N21);
nand NAND4 (N347, N314, N241, N193, N35);
nor NOR4 (N348, N338, N174, N296, N307);
or OR2 (N349, N344, N200);
nor NOR4 (N350, N348, N134, N197, N64);
buf BUF1 (N351, N326);
xor XOR2 (N352, N343, N83);
nand NAND4 (N353, N347, N194, N151, N150);
xor XOR2 (N354, N352, N281);
or OR2 (N355, N340, N133);
nand NAND4 (N356, N342, N61, N340, N26);
or OR3 (N357, N353, N236, N329);
xor XOR2 (N358, N357, N271);
xor XOR2 (N359, N355, N350);
nand NAND2 (N360, N343, N2);
nor NOR3 (N361, N359, N290, N81);
or OR4 (N362, N354, N349, N173, N151);
and AND3 (N363, N5, N31, N74);
nor NOR4 (N364, N363, N222, N229, N173);
nor NOR2 (N365, N362, N95);
nor NOR2 (N366, N356, N300);
buf BUF1 (N367, N364);
or OR4 (N368, N360, N11, N73, N49);
xor XOR2 (N369, N345, N126);
or OR4 (N370, N365, N176, N323, N42);
xor XOR2 (N371, N358, N131);
nand NAND4 (N372, N346, N173, N322, N59);
buf BUF1 (N373, N367);
or OR4 (N374, N351, N139, N6, N303);
nor NOR2 (N375, N373, N39);
xor XOR2 (N376, N375, N11);
and AND2 (N377, N332, N86);
xor XOR2 (N378, N372, N294);
nand NAND2 (N379, N378, N239);
and AND4 (N380, N377, N162, N149, N148);
nor NOR3 (N381, N369, N221, N19);
xor XOR2 (N382, N376, N288);
nand NAND2 (N383, N370, N245);
nand NAND4 (N384, N380, N80, N92, N241);
xor XOR2 (N385, N383, N187);
nor NOR3 (N386, N382, N91, N256);
nand NAND4 (N387, N366, N225, N14, N369);
nand NAND2 (N388, N386, N329);
and AND2 (N389, N381, N174);
not NOT1 (N390, N387);
or OR3 (N391, N390, N246, N12);
and AND2 (N392, N361, N116);
nor NOR3 (N393, N379, N193, N124);
or OR3 (N394, N374, N382, N249);
and AND4 (N395, N384, N385, N382, N154);
or OR2 (N396, N230, N268);
buf BUF1 (N397, N371);
and AND2 (N398, N392, N148);
xor XOR2 (N399, N368, N351);
or OR3 (N400, N397, N279, N92);
nand NAND2 (N401, N399, N162);
or OR4 (N402, N393, N136, N132, N311);
or OR3 (N403, N400, N108, N158);
buf BUF1 (N404, N402);
xor XOR2 (N405, N391, N163);
not NOT1 (N406, N405);
buf BUF1 (N407, N401);
and AND3 (N408, N406, N177, N299);
or OR4 (N409, N396, N406, N348, N20);
nor NOR2 (N410, N398, N94);
or OR3 (N411, N388, N74, N55);
nor NOR3 (N412, N411, N134, N45);
not NOT1 (N413, N403);
xor XOR2 (N414, N412, N201);
not NOT1 (N415, N409);
nand NAND3 (N416, N407, N17, N35);
or OR3 (N417, N413, N258, N343);
buf BUF1 (N418, N394);
buf BUF1 (N419, N395);
and AND2 (N420, N404, N86);
nor NOR2 (N421, N408, N416);
nand NAND3 (N422, N92, N239, N134);
not NOT1 (N423, N414);
nand NAND2 (N424, N417, N109);
not NOT1 (N425, N419);
buf BUF1 (N426, N425);
or OR4 (N427, N420, N100, N312, N117);
nor NOR4 (N428, N422, N362, N69, N198);
nand NAND4 (N429, N427, N32, N339, N91);
buf BUF1 (N430, N423);
and AND2 (N431, N424, N403);
and AND2 (N432, N389, N356);
or OR3 (N433, N430, N191, N419);
and AND4 (N434, N415, N393, N179, N323);
nand NAND4 (N435, N428, N94, N289, N274);
not NOT1 (N436, N433);
buf BUF1 (N437, N436);
not NOT1 (N438, N429);
or OR2 (N439, N421, N147);
nand NAND2 (N440, N426, N167);
nand NAND3 (N441, N431, N437, N321);
and AND4 (N442, N264, N361, N401, N201);
nor NOR3 (N443, N410, N284, N190);
and AND4 (N444, N441, N226, N318, N78);
xor XOR2 (N445, N438, N339);
or OR2 (N446, N435, N32);
buf BUF1 (N447, N434);
or OR2 (N448, N447, N349);
buf BUF1 (N449, N444);
buf BUF1 (N450, N446);
or OR4 (N451, N449, N404, N71, N150);
buf BUF1 (N452, N443);
and AND2 (N453, N451, N328);
buf BUF1 (N454, N453);
nor NOR3 (N455, N448, N333, N366);
and AND3 (N456, N432, N245, N328);
nand NAND4 (N457, N456, N118, N257, N168);
not NOT1 (N458, N418);
and AND2 (N459, N439, N411);
nor NOR3 (N460, N454, N318, N93);
buf BUF1 (N461, N455);
not NOT1 (N462, N459);
xor XOR2 (N463, N452, N368);
nand NAND3 (N464, N458, N88, N248);
not NOT1 (N465, N457);
buf BUF1 (N466, N463);
xor XOR2 (N467, N440, N339);
nor NOR4 (N468, N445, N298, N214, N205);
or OR2 (N469, N464, N51);
nor NOR4 (N470, N467, N294, N193, N46);
not NOT1 (N471, N462);
xor XOR2 (N472, N442, N237);
nor NOR2 (N473, N470, N212);
nor NOR4 (N474, N471, N399, N271, N202);
nor NOR2 (N475, N460, N231);
not NOT1 (N476, N473);
nand NAND2 (N477, N461, N47);
or OR4 (N478, N469, N302, N403, N34);
and AND4 (N479, N478, N458, N362, N32);
nand NAND3 (N480, N477, N476, N172);
and AND2 (N481, N331, N454);
nor NOR3 (N482, N480, N81, N184);
not NOT1 (N483, N481);
xor XOR2 (N484, N466, N351);
or OR3 (N485, N479, N337, N52);
nand NAND4 (N486, N482, N219, N314, N183);
buf BUF1 (N487, N483);
not NOT1 (N488, N484);
and AND3 (N489, N474, N370, N460);
xor XOR2 (N490, N489, N420);
or OR3 (N491, N468, N475, N462);
xor XOR2 (N492, N30, N477);
nand NAND4 (N493, N450, N90, N435, N83);
not NOT1 (N494, N472);
and AND2 (N495, N494, N13);
xor XOR2 (N496, N490, N130);
not NOT1 (N497, N496);
and AND3 (N498, N495, N246, N410);
or OR4 (N499, N485, N426, N83, N443);
and AND3 (N500, N493, N328, N489);
or OR3 (N501, N465, N214, N376);
not NOT1 (N502, N501);
buf BUF1 (N503, N487);
buf BUF1 (N504, N486);
nand NAND2 (N505, N498, N401);
not NOT1 (N506, N505);
buf BUF1 (N507, N488);
buf BUF1 (N508, N491);
and AND2 (N509, N499, N499);
xor XOR2 (N510, N497, N18);
buf BUF1 (N511, N503);
or OR4 (N512, N502, N364, N285, N48);
not NOT1 (N513, N506);
nand NAND4 (N514, N510, N53, N293, N230);
nand NAND2 (N515, N513, N2);
nor NOR3 (N516, N509, N30, N448);
nand NAND4 (N517, N508, N249, N138, N363);
not NOT1 (N518, N514);
and AND2 (N519, N515, N369);
buf BUF1 (N520, N500);
buf BUF1 (N521, N492);
or OR3 (N522, N512, N321, N224);
not NOT1 (N523, N511);
buf BUF1 (N524, N521);
buf BUF1 (N525, N524);
buf BUF1 (N526, N517);
or OR2 (N527, N504, N28);
buf BUF1 (N528, N522);
nand NAND3 (N529, N507, N408, N379);
xor XOR2 (N530, N523, N37);
or OR4 (N531, N519, N250, N358, N210);
nor NOR2 (N532, N526, N149);
buf BUF1 (N533, N527);
not NOT1 (N534, N529);
or OR3 (N535, N525, N191, N370);
nand NAND3 (N536, N518, N268, N73);
buf BUF1 (N537, N516);
or OR3 (N538, N537, N341, N87);
buf BUF1 (N539, N528);
buf BUF1 (N540, N533);
nand NAND3 (N541, N532, N429, N467);
nand NAND4 (N542, N536, N280, N349, N521);
not NOT1 (N543, N539);
xor XOR2 (N544, N520, N66);
nand NAND2 (N545, N544, N83);
nor NOR4 (N546, N530, N163, N414, N508);
and AND3 (N547, N535, N320, N527);
xor XOR2 (N548, N547, N541);
not NOT1 (N549, N301);
or OR3 (N550, N548, N365, N434);
xor XOR2 (N551, N550, N197);
xor XOR2 (N552, N540, N272);
nand NAND2 (N553, N551, N373);
or OR2 (N554, N553, N47);
and AND4 (N555, N554, N100, N61, N464);
xor XOR2 (N556, N545, N168);
nor NOR2 (N557, N542, N429);
nor NOR3 (N558, N534, N498, N275);
or OR2 (N559, N538, N322);
buf BUF1 (N560, N531);
xor XOR2 (N561, N555, N383);
or OR3 (N562, N552, N543, N251);
xor XOR2 (N563, N323, N234);
nand NAND2 (N564, N563, N276);
nand NAND4 (N565, N557, N399, N35, N99);
xor XOR2 (N566, N565, N558);
nor NOR2 (N567, N396, N94);
not NOT1 (N568, N546);
nor NOR2 (N569, N568, N447);
nand NAND2 (N570, N560, N240);
not NOT1 (N571, N562);
buf BUF1 (N572, N566);
nand NAND3 (N573, N561, N356, N539);
nor NOR2 (N574, N556, N503);
or OR2 (N575, N567, N455);
not NOT1 (N576, N569);
or OR4 (N577, N572, N34, N84, N329);
or OR4 (N578, N573, N375, N237, N419);
buf BUF1 (N579, N571);
nand NAND4 (N580, N549, N177, N122, N461);
xor XOR2 (N581, N575, N273);
xor XOR2 (N582, N576, N254);
not NOT1 (N583, N564);
or OR4 (N584, N579, N258, N319, N341);
nor NOR2 (N585, N584, N549);
nand NAND3 (N586, N577, N313, N334);
not NOT1 (N587, N583);
buf BUF1 (N588, N570);
nand NAND4 (N589, N587, N192, N18, N572);
xor XOR2 (N590, N589, N565);
nand NAND4 (N591, N559, N240, N174, N380);
nand NAND2 (N592, N588, N549);
nand NAND4 (N593, N582, N93, N193, N438);
nor NOR3 (N594, N580, N530, N260);
and AND4 (N595, N586, N481, N308, N444);
or OR3 (N596, N593, N312, N293);
and AND2 (N597, N574, N238);
xor XOR2 (N598, N591, N365);
xor XOR2 (N599, N594, N274);
not NOT1 (N600, N596);
and AND3 (N601, N585, N447, N158);
nand NAND2 (N602, N599, N180);
nor NOR2 (N603, N595, N394);
or OR2 (N604, N602, N295);
nand NAND3 (N605, N578, N197, N421);
and AND2 (N606, N590, N121);
and AND4 (N607, N604, N128, N56, N291);
buf BUF1 (N608, N597);
nand NAND2 (N609, N581, N407);
buf BUF1 (N610, N600);
nand NAND4 (N611, N603, N423, N379, N571);
nand NAND4 (N612, N611, N168, N171, N137);
or OR2 (N613, N598, N508);
buf BUF1 (N614, N610);
not NOT1 (N615, N614);
or OR3 (N616, N608, N58, N76);
and AND4 (N617, N615, N96, N545, N348);
buf BUF1 (N618, N606);
not NOT1 (N619, N617);
nand NAND4 (N620, N618, N269, N396, N292);
nand NAND3 (N621, N612, N121, N445);
nand NAND4 (N622, N621, N40, N401, N549);
nand NAND4 (N623, N622, N212, N119, N266);
not NOT1 (N624, N601);
not NOT1 (N625, N623);
or OR2 (N626, N624, N197);
and AND4 (N627, N620, N29, N279, N82);
not NOT1 (N628, N619);
not NOT1 (N629, N613);
not NOT1 (N630, N627);
buf BUF1 (N631, N628);
nand NAND2 (N632, N626, N336);
nor NOR4 (N633, N629, N317, N34, N5);
and AND4 (N634, N592, N281, N4, N548);
xor XOR2 (N635, N605, N18);
or OR4 (N636, N630, N581, N619, N35);
nand NAND4 (N637, N631, N129, N434, N165);
or OR4 (N638, N636, N365, N353, N150);
xor XOR2 (N639, N625, N458);
or OR4 (N640, N616, N197, N27, N288);
buf BUF1 (N641, N634);
not NOT1 (N642, N639);
buf BUF1 (N643, N638);
and AND3 (N644, N637, N297, N600);
or OR4 (N645, N643, N538, N17, N504);
and AND2 (N646, N642, N294);
buf BUF1 (N647, N640);
not NOT1 (N648, N644);
buf BUF1 (N649, N648);
nand NAND2 (N650, N649, N160);
xor XOR2 (N651, N609, N324);
buf BUF1 (N652, N635);
and AND4 (N653, N650, N388, N87, N198);
buf BUF1 (N654, N641);
nor NOR4 (N655, N633, N116, N515, N390);
nor NOR3 (N656, N632, N179, N96);
not NOT1 (N657, N607);
nor NOR4 (N658, N656, N374, N346, N448);
not NOT1 (N659, N658);
nand NAND4 (N660, N647, N217, N390, N4);
not NOT1 (N661, N653);
or OR3 (N662, N652, N561, N434);
nor NOR4 (N663, N661, N576, N522, N551);
or OR2 (N664, N662, N379);
not NOT1 (N665, N657);
nor NOR2 (N666, N646, N434);
nor NOR4 (N667, N663, N484, N598, N380);
and AND2 (N668, N645, N382);
nand NAND4 (N669, N666, N46, N223, N596);
or OR2 (N670, N659, N490);
nand NAND4 (N671, N655, N548, N452, N391);
nor NOR4 (N672, N651, N237, N150, N213);
not NOT1 (N673, N667);
xor XOR2 (N674, N660, N228);
buf BUF1 (N675, N669);
not NOT1 (N676, N654);
nand NAND3 (N677, N676, N203, N171);
and AND4 (N678, N675, N465, N513, N468);
and AND3 (N679, N670, N190, N394);
or OR2 (N680, N673, N108);
and AND3 (N681, N677, N141, N676);
not NOT1 (N682, N678);
nand NAND3 (N683, N668, N242, N620);
xor XOR2 (N684, N682, N430);
nand NAND4 (N685, N679, N148, N191, N397);
nand NAND2 (N686, N674, N311);
or OR4 (N687, N683, N544, N474, N112);
nor NOR4 (N688, N684, N378, N492, N55);
xor XOR2 (N689, N687, N678);
nand NAND3 (N690, N672, N295, N574);
nor NOR2 (N691, N690, N468);
and AND2 (N692, N671, N263);
or OR4 (N693, N685, N486, N401, N373);
or OR4 (N694, N665, N286, N14, N600);
and AND4 (N695, N686, N330, N110, N134);
and AND3 (N696, N689, N116, N158);
or OR2 (N697, N688, N672);
nand NAND3 (N698, N696, N100, N495);
nor NOR2 (N699, N695, N83);
not NOT1 (N700, N664);
xor XOR2 (N701, N700, N310);
buf BUF1 (N702, N694);
nand NAND3 (N703, N680, N639, N290);
or OR4 (N704, N701, N217, N344, N539);
nor NOR2 (N705, N698, N276);
not NOT1 (N706, N702);
nand NAND2 (N707, N699, N253);
or OR2 (N708, N706, N401);
nor NOR4 (N709, N703, N394, N104, N161);
buf BUF1 (N710, N709);
or OR4 (N711, N704, N486, N651, N23);
and AND3 (N712, N692, N535, N44);
nand NAND3 (N713, N705, N467, N116);
not NOT1 (N714, N708);
buf BUF1 (N715, N697);
or OR3 (N716, N691, N143, N25);
xor XOR2 (N717, N681, N48);
nand NAND4 (N718, N716, N547, N322, N105);
or OR4 (N719, N712, N121, N67, N122);
and AND3 (N720, N710, N665, N55);
not NOT1 (N721, N720);
and AND3 (N722, N707, N118, N690);
nor NOR4 (N723, N718, N324, N231, N531);
or OR2 (N724, N719, N286);
and AND2 (N725, N711, N221);
not NOT1 (N726, N715);
or OR3 (N727, N722, N290, N663);
buf BUF1 (N728, N723);
or OR4 (N729, N724, N208, N695, N234);
or OR2 (N730, N721, N137);
and AND4 (N731, N717, N592, N478, N166);
nand NAND3 (N732, N726, N232, N66);
xor XOR2 (N733, N727, N349);
or OR2 (N734, N731, N372);
and AND2 (N735, N732, N715);
not NOT1 (N736, N725);
buf BUF1 (N737, N733);
buf BUF1 (N738, N713);
not NOT1 (N739, N737);
not NOT1 (N740, N729);
and AND2 (N741, N736, N562);
nor NOR3 (N742, N740, N301, N696);
buf BUF1 (N743, N734);
nor NOR2 (N744, N693, N617);
nand NAND2 (N745, N735, N195);
not NOT1 (N746, N714);
buf BUF1 (N747, N741);
nor NOR3 (N748, N744, N670, N588);
nor NOR4 (N749, N728, N383, N514, N44);
not NOT1 (N750, N743);
xor XOR2 (N751, N749, N262);
and AND2 (N752, N746, N521);
and AND2 (N753, N742, N481);
and AND4 (N754, N751, N494, N65, N288);
nor NOR2 (N755, N745, N249);
not NOT1 (N756, N752);
nand NAND2 (N757, N750, N138);
nand NAND4 (N758, N747, N709, N274, N268);
or OR3 (N759, N738, N720, N164);
xor XOR2 (N760, N757, N535);
xor XOR2 (N761, N759, N259);
xor XOR2 (N762, N754, N509);
and AND2 (N763, N761, N222);
nand NAND3 (N764, N730, N555, N707);
not NOT1 (N765, N748);
nand NAND3 (N766, N764, N558, N617);
and AND4 (N767, N762, N424, N531, N239);
buf BUF1 (N768, N753);
buf BUF1 (N769, N765);
or OR2 (N770, N763, N707);
nand NAND2 (N771, N770, N348);
and AND2 (N772, N756, N441);
and AND4 (N773, N769, N214, N90, N373);
nor NOR4 (N774, N758, N648, N177, N641);
not NOT1 (N775, N760);
or OR3 (N776, N772, N644, N651);
nand NAND3 (N777, N767, N534, N383);
xor XOR2 (N778, N755, N749);
not NOT1 (N779, N766);
and AND4 (N780, N778, N470, N240, N622);
nor NOR2 (N781, N739, N67);
buf BUF1 (N782, N779);
or OR4 (N783, N780, N213, N440, N288);
or OR4 (N784, N782, N681, N129, N68);
nand NAND3 (N785, N783, N145, N23);
and AND4 (N786, N781, N501, N12, N218);
nor NOR2 (N787, N774, N694);
buf BUF1 (N788, N785);
nor NOR4 (N789, N776, N745, N465, N198);
and AND3 (N790, N771, N663, N471);
nand NAND4 (N791, N773, N248, N641, N724);
nand NAND2 (N792, N788, N267);
not NOT1 (N793, N768);
and AND3 (N794, N786, N761, N195);
or OR2 (N795, N777, N402);
buf BUF1 (N796, N793);
or OR3 (N797, N787, N146, N524);
nor NOR4 (N798, N796, N537, N623, N729);
nand NAND4 (N799, N789, N248, N657, N372);
nor NOR4 (N800, N790, N401, N470, N251);
or OR3 (N801, N792, N4, N548);
not NOT1 (N802, N791);
nor NOR3 (N803, N784, N771, N277);
nor NOR2 (N804, N798, N25);
xor XOR2 (N805, N799, N765);
and AND2 (N806, N804, N776);
buf BUF1 (N807, N797);
xor XOR2 (N808, N807, N147);
or OR3 (N809, N802, N488, N514);
not NOT1 (N810, N775);
nand NAND3 (N811, N800, N39, N131);
buf BUF1 (N812, N809);
xor XOR2 (N813, N803, N340);
xor XOR2 (N814, N813, N396);
not NOT1 (N815, N805);
xor XOR2 (N816, N808, N149);
nand NAND3 (N817, N811, N367, N260);
not NOT1 (N818, N815);
not NOT1 (N819, N816);
nor NOR4 (N820, N806, N602, N199, N557);
xor XOR2 (N821, N801, N294);
nor NOR4 (N822, N810, N788, N327, N373);
or OR4 (N823, N814, N564, N315, N444);
nand NAND4 (N824, N823, N25, N543, N815);
nand NAND3 (N825, N820, N516, N590);
xor XOR2 (N826, N794, N641);
xor XOR2 (N827, N818, N324);
xor XOR2 (N828, N826, N351);
or OR3 (N829, N827, N156, N2);
or OR4 (N830, N828, N689, N2, N483);
xor XOR2 (N831, N824, N355);
nor NOR4 (N832, N819, N782, N327, N13);
nand NAND4 (N833, N821, N284, N805, N793);
buf BUF1 (N834, N831);
buf BUF1 (N835, N829);
nor NOR3 (N836, N817, N298, N375);
and AND2 (N837, N830, N220);
or OR2 (N838, N812, N230);
and AND2 (N839, N835, N246);
buf BUF1 (N840, N834);
buf BUF1 (N841, N833);
nor NOR3 (N842, N836, N613, N601);
buf BUF1 (N843, N825);
buf BUF1 (N844, N840);
nor NOR4 (N845, N837, N257, N716, N143);
not NOT1 (N846, N841);
nand NAND2 (N847, N842, N483);
xor XOR2 (N848, N832, N799);
nand NAND2 (N849, N843, N330);
not NOT1 (N850, N844);
nor NOR2 (N851, N849, N272);
nand NAND4 (N852, N848, N250, N674, N421);
xor XOR2 (N853, N839, N542);
xor XOR2 (N854, N838, N722);
xor XOR2 (N855, N795, N446);
xor XOR2 (N856, N853, N304);
nor NOR3 (N857, N846, N702, N770);
xor XOR2 (N858, N851, N769);
or OR2 (N859, N854, N521);
and AND2 (N860, N850, N162);
nor NOR3 (N861, N860, N829, N62);
and AND2 (N862, N822, N114);
not NOT1 (N863, N845);
nand NAND4 (N864, N855, N747, N285, N720);
or OR4 (N865, N861, N64, N97, N389);
not NOT1 (N866, N859);
nor NOR4 (N867, N865, N322, N505, N55);
nor NOR4 (N868, N857, N598, N41, N808);
xor XOR2 (N869, N864, N122);
nor NOR2 (N870, N869, N695);
or OR3 (N871, N868, N53, N308);
not NOT1 (N872, N866);
and AND4 (N873, N870, N178, N748, N145);
or OR3 (N874, N863, N587, N828);
and AND4 (N875, N871, N91, N750, N214);
xor XOR2 (N876, N873, N721);
and AND4 (N877, N856, N427, N155, N769);
not NOT1 (N878, N875);
buf BUF1 (N879, N878);
xor XOR2 (N880, N879, N525);
nand NAND2 (N881, N847, N426);
nand NAND3 (N882, N876, N388, N241);
buf BUF1 (N883, N880);
and AND4 (N884, N882, N177, N555, N698);
and AND4 (N885, N883, N325, N141, N594);
nor NOR4 (N886, N862, N285, N106, N774);
not NOT1 (N887, N858);
nor NOR3 (N888, N885, N79, N175);
nand NAND4 (N889, N887, N448, N866, N765);
or OR2 (N890, N874, N139);
nor NOR3 (N891, N872, N511, N527);
nor NOR2 (N892, N888, N395);
or OR4 (N893, N891, N684, N583, N257);
or OR2 (N894, N892, N117);
and AND2 (N895, N877, N367);
buf BUF1 (N896, N884);
xor XOR2 (N897, N893, N803);
not NOT1 (N898, N881);
nand NAND2 (N899, N889, N775);
nor NOR4 (N900, N886, N416, N265, N704);
or OR3 (N901, N894, N26, N315);
xor XOR2 (N902, N901, N739);
buf BUF1 (N903, N899);
xor XOR2 (N904, N903, N81);
and AND4 (N905, N900, N887, N275, N831);
nor NOR3 (N906, N852, N2, N98);
buf BUF1 (N907, N898);
nand NAND2 (N908, N907, N361);
and AND4 (N909, N902, N734, N363, N872);
not NOT1 (N910, N906);
not NOT1 (N911, N905);
xor XOR2 (N912, N911, N580);
buf BUF1 (N913, N912);
nand NAND4 (N914, N910, N87, N397, N669);
buf BUF1 (N915, N908);
nor NOR3 (N916, N867, N64, N331);
buf BUF1 (N917, N890);
not NOT1 (N918, N913);
or OR2 (N919, N914, N529);
xor XOR2 (N920, N896, N889);
xor XOR2 (N921, N920, N270);
nand NAND4 (N922, N918, N140, N192, N1);
xor XOR2 (N923, N922, N467);
nor NOR4 (N924, N917, N775, N504, N571);
and AND2 (N925, N916, N291);
xor XOR2 (N926, N904, N148);
not NOT1 (N927, N923);
nand NAND3 (N928, N895, N477, N860);
nor NOR4 (N929, N927, N451, N7, N777);
xor XOR2 (N930, N921, N37);
or OR2 (N931, N915, N125);
nand NAND4 (N932, N925, N884, N785, N468);
buf BUF1 (N933, N929);
nor NOR2 (N934, N926, N343);
buf BUF1 (N935, N928);
xor XOR2 (N936, N897, N711);
nor NOR4 (N937, N909, N294, N470, N834);
nand NAND3 (N938, N919, N561, N678);
and AND2 (N939, N936, N515);
not NOT1 (N940, N935);
nor NOR3 (N941, N930, N928, N867);
buf BUF1 (N942, N934);
nor NOR2 (N943, N940, N193);
nand NAND2 (N944, N941, N689);
and AND4 (N945, N937, N186, N80, N683);
not NOT1 (N946, N932);
and AND4 (N947, N945, N739, N914, N887);
not NOT1 (N948, N942);
or OR2 (N949, N946, N80);
xor XOR2 (N950, N944, N542);
or OR2 (N951, N949, N685);
xor XOR2 (N952, N933, N271);
nor NOR2 (N953, N931, N535);
nor NOR4 (N954, N950, N853, N355, N121);
xor XOR2 (N955, N954, N421);
or OR3 (N956, N924, N490, N458);
nor NOR2 (N957, N952, N951);
nand NAND3 (N958, N747, N436, N103);
not NOT1 (N959, N957);
buf BUF1 (N960, N956);
nor NOR3 (N961, N953, N808, N837);
buf BUF1 (N962, N943);
buf BUF1 (N963, N959);
and AND3 (N964, N958, N71, N840);
nor NOR3 (N965, N939, N488, N512);
xor XOR2 (N966, N961, N919);
nor NOR3 (N967, N938, N444, N324);
and AND3 (N968, N964, N121, N836);
not NOT1 (N969, N965);
xor XOR2 (N970, N948, N696);
nor NOR4 (N971, N960, N496, N926, N172);
nand NAND4 (N972, N971, N177, N102, N432);
and AND3 (N973, N968, N430, N145);
nor NOR3 (N974, N962, N192, N346);
and AND4 (N975, N969, N575, N104, N264);
nor NOR3 (N976, N967, N964, N370);
nor NOR2 (N977, N970, N340);
or OR2 (N978, N977, N126);
nand NAND4 (N979, N978, N825, N468, N115);
and AND4 (N980, N979, N303, N196, N249);
nor NOR4 (N981, N980, N194, N874, N31);
nand NAND2 (N982, N972, N101);
xor XOR2 (N983, N974, N317);
buf BUF1 (N984, N975);
xor XOR2 (N985, N947, N431);
buf BUF1 (N986, N963);
nor NOR2 (N987, N985, N88);
or OR3 (N988, N982, N768, N840);
and AND3 (N989, N984, N401, N174);
nor NOR2 (N990, N983, N189);
nand NAND3 (N991, N973, N81, N173);
xor XOR2 (N992, N981, N708);
not NOT1 (N993, N988);
nand NAND2 (N994, N992, N315);
buf BUF1 (N995, N955);
nor NOR4 (N996, N987, N341, N896, N222);
not NOT1 (N997, N994);
and AND4 (N998, N966, N114, N921, N427);
nand NAND4 (N999, N976, N497, N892, N819);
and AND3 (N1000, N999, N366, N767);
and AND3 (N1001, N997, N681, N285);
nor NOR4 (N1002, N986, N663, N47, N745);
or OR4 (N1003, N989, N581, N16, N947);
nor NOR2 (N1004, N993, N889);
or OR4 (N1005, N1004, N431, N89, N254);
nand NAND4 (N1006, N1001, N637, N157, N218);
and AND2 (N1007, N1003, N808);
and AND4 (N1008, N1005, N813, N670, N321);
and AND4 (N1009, N1007, N178, N990, N968);
nand NAND3 (N1010, N884, N402, N44);
nor NOR2 (N1011, N1006, N394);
nor NOR3 (N1012, N1011, N408, N672);
xor XOR2 (N1013, N995, N6);
or OR3 (N1014, N1013, N899, N177);
xor XOR2 (N1015, N1002, N943);
nor NOR2 (N1016, N998, N558);
and AND3 (N1017, N1000, N54, N969);
or OR2 (N1018, N1016, N509);
nor NOR3 (N1019, N996, N542, N280);
or OR2 (N1020, N1014, N710);
or OR4 (N1021, N1018, N598, N912, N624);
nor NOR4 (N1022, N1015, N416, N848, N811);
or OR4 (N1023, N1010, N38, N491, N15);
or OR2 (N1024, N1023, N719);
or OR2 (N1025, N1008, N548);
xor XOR2 (N1026, N1009, N959);
buf BUF1 (N1027, N1024);
nand NAND4 (N1028, N991, N862, N7, N977);
nor NOR4 (N1029, N1025, N1004, N800, N710);
buf BUF1 (N1030, N1029);
nand NAND3 (N1031, N1012, N78, N17);
or OR4 (N1032, N1031, N109, N590, N818);
xor XOR2 (N1033, N1021, N832);
nand NAND2 (N1034, N1030, N769);
xor XOR2 (N1035, N1033, N823);
and AND4 (N1036, N1027, N22, N252, N779);
not NOT1 (N1037, N1035);
nor NOR3 (N1038, N1032, N785, N863);
nand NAND4 (N1039, N1038, N150, N232, N395);
xor XOR2 (N1040, N1026, N170);
buf BUF1 (N1041, N1036);
xor XOR2 (N1042, N1040, N582);
xor XOR2 (N1043, N1020, N455);
buf BUF1 (N1044, N1022);
or OR3 (N1045, N1028, N820, N185);
xor XOR2 (N1046, N1037, N493);
buf BUF1 (N1047, N1039);
buf BUF1 (N1048, N1047);
buf BUF1 (N1049, N1044);
buf BUF1 (N1050, N1042);
nand NAND4 (N1051, N1041, N974, N619, N786);
nand NAND3 (N1052, N1034, N685, N337);
nor NOR2 (N1053, N1043, N431);
xor XOR2 (N1054, N1052, N73);
xor XOR2 (N1055, N1049, N38);
not NOT1 (N1056, N1055);
xor XOR2 (N1057, N1056, N90);
nand NAND2 (N1058, N1053, N138);
xor XOR2 (N1059, N1017, N809);
nor NOR3 (N1060, N1019, N388, N293);
xor XOR2 (N1061, N1051, N559);
not NOT1 (N1062, N1046);
xor XOR2 (N1063, N1060, N822);
not NOT1 (N1064, N1059);
or OR4 (N1065, N1061, N630, N366, N527);
nand NAND2 (N1066, N1065, N1065);
xor XOR2 (N1067, N1050, N687);
and AND3 (N1068, N1058, N403, N98);
not NOT1 (N1069, N1057);
or OR3 (N1070, N1062, N40, N206);
xor XOR2 (N1071, N1054, N520);
buf BUF1 (N1072, N1068);
and AND4 (N1073, N1070, N942, N997, N4);
nor NOR2 (N1074, N1063, N431);
nand NAND4 (N1075, N1064, N199, N508, N198);
nand NAND2 (N1076, N1075, N110);
nor NOR4 (N1077, N1045, N992, N367, N853);
nor NOR2 (N1078, N1048, N265);
or OR3 (N1079, N1074, N31, N610);
and AND4 (N1080, N1079, N43, N678, N16);
xor XOR2 (N1081, N1069, N385);
nand NAND3 (N1082, N1077, N349, N430);
or OR3 (N1083, N1076, N628, N450);
not NOT1 (N1084, N1082);
not NOT1 (N1085, N1073);
and AND4 (N1086, N1081, N19, N136, N112);
buf BUF1 (N1087, N1086);
and AND3 (N1088, N1066, N751, N467);
nor NOR4 (N1089, N1083, N38, N123, N814);
buf BUF1 (N1090, N1085);
not NOT1 (N1091, N1084);
nor NOR4 (N1092, N1087, N150, N1009, N478);
and AND3 (N1093, N1088, N219, N120);
nand NAND4 (N1094, N1090, N1078, N379, N1006);
nor NOR2 (N1095, N478, N814);
buf BUF1 (N1096, N1092);
nand NAND2 (N1097, N1096, N556);
or OR3 (N1098, N1071, N46, N195);
and AND2 (N1099, N1093, N766);
and AND4 (N1100, N1067, N591, N326, N542);
nor NOR3 (N1101, N1094, N659, N781);
xor XOR2 (N1102, N1091, N756);
and AND3 (N1103, N1097, N685, N521);
buf BUF1 (N1104, N1100);
and AND2 (N1105, N1098, N831);
buf BUF1 (N1106, N1089);
and AND4 (N1107, N1105, N655, N674, N815);
buf BUF1 (N1108, N1101);
buf BUF1 (N1109, N1103);
buf BUF1 (N1110, N1095);
nor NOR3 (N1111, N1080, N563, N546);
and AND3 (N1112, N1111, N77, N1109);
or OR2 (N1113, N221, N366);
nor NOR4 (N1114, N1108, N456, N583, N755);
and AND4 (N1115, N1113, N421, N132, N79);
xor XOR2 (N1116, N1072, N345);
and AND3 (N1117, N1114, N615, N540);
not NOT1 (N1118, N1115);
and AND3 (N1119, N1110, N18, N43);
nand NAND3 (N1120, N1117, N572, N425);
and AND4 (N1121, N1099, N408, N645, N69);
nand NAND3 (N1122, N1112, N357, N436);
nor NOR2 (N1123, N1107, N189);
nor NOR2 (N1124, N1102, N644);
nor NOR2 (N1125, N1118, N922);
xor XOR2 (N1126, N1123, N499);
nor NOR2 (N1127, N1106, N1059);
nor NOR4 (N1128, N1116, N41, N1038, N8);
and AND2 (N1129, N1104, N1036);
xor XOR2 (N1130, N1122, N1015);
and AND4 (N1131, N1121, N779, N154, N784);
and AND4 (N1132, N1129, N907, N512, N1089);
xor XOR2 (N1133, N1131, N680);
xor XOR2 (N1134, N1119, N915);
or OR4 (N1135, N1128, N258, N192, N102);
and AND4 (N1136, N1125, N199, N627, N576);
or OR2 (N1137, N1136, N776);
nand NAND3 (N1138, N1133, N781, N49);
xor XOR2 (N1139, N1124, N802);
nor NOR4 (N1140, N1134, N360, N84, N703);
or OR4 (N1141, N1120, N969, N260, N266);
nand NAND4 (N1142, N1126, N918, N637, N1039);
nor NOR3 (N1143, N1127, N547, N838);
not NOT1 (N1144, N1132);
and AND2 (N1145, N1137, N484);
nand NAND3 (N1146, N1138, N881, N731);
and AND4 (N1147, N1130, N696, N741, N879);
nor NOR2 (N1148, N1146, N768);
buf BUF1 (N1149, N1140);
buf BUF1 (N1150, N1144);
nor NOR3 (N1151, N1148, N38, N1032);
buf BUF1 (N1152, N1147);
and AND2 (N1153, N1135, N122);
xor XOR2 (N1154, N1150, N656);
not NOT1 (N1155, N1149);
not NOT1 (N1156, N1142);
not NOT1 (N1157, N1156);
nand NAND2 (N1158, N1145, N528);
and AND2 (N1159, N1141, N1153);
and AND2 (N1160, N376, N440);
xor XOR2 (N1161, N1151, N873);
nor NOR3 (N1162, N1158, N1051, N660);
nor NOR2 (N1163, N1159, N111);
nand NAND3 (N1164, N1157, N662, N78);
not NOT1 (N1165, N1143);
buf BUF1 (N1166, N1162);
nor NOR4 (N1167, N1155, N638, N612, N790);
nor NOR4 (N1168, N1152, N300, N657, N739);
xor XOR2 (N1169, N1163, N846);
buf BUF1 (N1170, N1161);
xor XOR2 (N1171, N1165, N765);
nand NAND2 (N1172, N1154, N587);
nor NOR4 (N1173, N1164, N883, N349, N743);
nand NAND2 (N1174, N1166, N1033);
nand NAND4 (N1175, N1174, N442, N722, N997);
and AND3 (N1176, N1139, N624, N83);
nand NAND4 (N1177, N1171, N990, N1109, N1170);
not NOT1 (N1178, N934);
xor XOR2 (N1179, N1167, N1010);
and AND2 (N1180, N1176, N984);
and AND3 (N1181, N1173, N534, N67);
nor NOR4 (N1182, N1168, N552, N30, N149);
nand NAND2 (N1183, N1181, N1034);
nor NOR3 (N1184, N1179, N75, N431);
nor NOR4 (N1185, N1175, N18, N859, N847);
xor XOR2 (N1186, N1160, N226);
buf BUF1 (N1187, N1177);
or OR4 (N1188, N1178, N1055, N751, N920);
xor XOR2 (N1189, N1183, N1164);
xor XOR2 (N1190, N1185, N406);
buf BUF1 (N1191, N1188);
and AND3 (N1192, N1169, N786, N66);
buf BUF1 (N1193, N1190);
buf BUF1 (N1194, N1193);
nor NOR3 (N1195, N1184, N705, N198);
and AND3 (N1196, N1195, N404, N933);
nand NAND2 (N1197, N1172, N493);
nor NOR4 (N1198, N1194, N511, N232, N667);
xor XOR2 (N1199, N1197, N336);
xor XOR2 (N1200, N1189, N93);
nand NAND4 (N1201, N1200, N317, N206, N628);
xor XOR2 (N1202, N1187, N1013);
and AND3 (N1203, N1202, N1098, N893);
or OR4 (N1204, N1192, N902, N476, N1143);
xor XOR2 (N1205, N1203, N481);
and AND3 (N1206, N1198, N717, N839);
and AND2 (N1207, N1199, N602);
buf BUF1 (N1208, N1201);
or OR4 (N1209, N1182, N335, N520, N360);
not NOT1 (N1210, N1208);
and AND2 (N1211, N1196, N786);
buf BUF1 (N1212, N1206);
not NOT1 (N1213, N1209);
nor NOR4 (N1214, N1207, N206, N81, N852);
or OR3 (N1215, N1210, N314, N53);
not NOT1 (N1216, N1211);
nor NOR2 (N1217, N1191, N370);
or OR4 (N1218, N1216, N431, N653, N132);
nor NOR4 (N1219, N1186, N521, N307, N103);
buf BUF1 (N1220, N1180);
buf BUF1 (N1221, N1220);
nand NAND3 (N1222, N1219, N252, N76);
or OR3 (N1223, N1214, N94, N572);
xor XOR2 (N1224, N1217, N1179);
nor NOR2 (N1225, N1204, N103);
not NOT1 (N1226, N1225);
or OR2 (N1227, N1212, N482);
or OR3 (N1228, N1205, N184, N745);
buf BUF1 (N1229, N1223);
and AND4 (N1230, N1228, N711, N811, N947);
or OR4 (N1231, N1213, N1184, N699, N1055);
xor XOR2 (N1232, N1229, N471);
nor NOR3 (N1233, N1226, N1025, N657);
or OR4 (N1234, N1232, N453, N683, N558);
xor XOR2 (N1235, N1218, N810);
buf BUF1 (N1236, N1224);
buf BUF1 (N1237, N1227);
nand NAND3 (N1238, N1222, N331, N456);
buf BUF1 (N1239, N1234);
not NOT1 (N1240, N1215);
xor XOR2 (N1241, N1237, N471);
or OR3 (N1242, N1241, N406, N488);
or OR2 (N1243, N1230, N1121);
or OR4 (N1244, N1238, N290, N332, N1180);
and AND3 (N1245, N1242, N346, N396);
buf BUF1 (N1246, N1221);
or OR2 (N1247, N1245, N733);
nor NOR4 (N1248, N1236, N73, N308, N284);
nor NOR4 (N1249, N1247, N476, N613, N195);
buf BUF1 (N1250, N1243);
not NOT1 (N1251, N1246);
buf BUF1 (N1252, N1244);
and AND3 (N1253, N1251, N721, N320);
and AND3 (N1254, N1240, N752, N729);
nor NOR3 (N1255, N1252, N293, N325);
not NOT1 (N1256, N1235);
nand NAND3 (N1257, N1231, N214, N451);
nor NOR3 (N1258, N1256, N683, N211);
nand NAND4 (N1259, N1255, N237, N741, N275);
nor NOR3 (N1260, N1249, N1164, N141);
nor NOR3 (N1261, N1239, N496, N1129);
or OR4 (N1262, N1248, N1202, N372, N186);
nor NOR4 (N1263, N1250, N310, N286, N153);
buf BUF1 (N1264, N1262);
nor NOR2 (N1265, N1260, N823);
buf BUF1 (N1266, N1261);
nand NAND4 (N1267, N1264, N785, N691, N5);
xor XOR2 (N1268, N1257, N1256);
xor XOR2 (N1269, N1253, N72);
and AND2 (N1270, N1268, N785);
nand NAND3 (N1271, N1233, N1018, N1219);
and AND2 (N1272, N1258, N1083);
or OR3 (N1273, N1263, N466, N1227);
nor NOR2 (N1274, N1271, N975);
and AND4 (N1275, N1265, N717, N193, N705);
nor NOR2 (N1276, N1266, N739);
not NOT1 (N1277, N1267);
nor NOR2 (N1278, N1259, N11);
nand NAND2 (N1279, N1273, N245);
xor XOR2 (N1280, N1274, N557);
buf BUF1 (N1281, N1269);
or OR3 (N1282, N1272, N1157, N178);
nand NAND2 (N1283, N1280, N980);
or OR2 (N1284, N1279, N498);
and AND2 (N1285, N1275, N192);
xor XOR2 (N1286, N1254, N467);
not NOT1 (N1287, N1282);
nand NAND4 (N1288, N1285, N145, N1146, N631);
or OR3 (N1289, N1276, N54, N144);
and AND4 (N1290, N1284, N420, N187, N158);
not NOT1 (N1291, N1270);
nand NAND3 (N1292, N1278, N1140, N795);
or OR4 (N1293, N1289, N404, N98, N491);
xor XOR2 (N1294, N1277, N238);
buf BUF1 (N1295, N1294);
nand NAND3 (N1296, N1281, N567, N1139);
nand NAND3 (N1297, N1293, N629, N651);
nand NAND4 (N1298, N1287, N1104, N1223, N166);
xor XOR2 (N1299, N1290, N644);
xor XOR2 (N1300, N1292, N1141);
or OR2 (N1301, N1288, N845);
or OR2 (N1302, N1295, N255);
nor NOR2 (N1303, N1286, N263);
buf BUF1 (N1304, N1302);
xor XOR2 (N1305, N1296, N417);
or OR2 (N1306, N1299, N1133);
nor NOR3 (N1307, N1303, N537, N155);
not NOT1 (N1308, N1300);
nand NAND4 (N1309, N1306, N1201, N1131, N199);
and AND4 (N1310, N1309, N541, N768, N511);
or OR3 (N1311, N1301, N175, N713);
xor XOR2 (N1312, N1297, N577);
nor NOR3 (N1313, N1310, N289, N1031);
not NOT1 (N1314, N1307);
nor NOR4 (N1315, N1312, N37, N95, N540);
not NOT1 (N1316, N1315);
nor NOR2 (N1317, N1316, N134);
nor NOR3 (N1318, N1308, N1006, N908);
and AND3 (N1319, N1313, N518, N430);
not NOT1 (N1320, N1291);
and AND2 (N1321, N1319, N1229);
buf BUF1 (N1322, N1311);
and AND3 (N1323, N1314, N1224, N227);
and AND2 (N1324, N1317, N1052);
nand NAND3 (N1325, N1322, N1138, N653);
buf BUF1 (N1326, N1298);
buf BUF1 (N1327, N1320);
not NOT1 (N1328, N1324);
nand NAND3 (N1329, N1304, N582, N494);
nor NOR2 (N1330, N1326, N1096);
and AND3 (N1331, N1321, N70, N883);
or OR4 (N1332, N1328, N133, N231, N1265);
nand NAND2 (N1333, N1325, N139);
or OR3 (N1334, N1323, N385, N1152);
and AND4 (N1335, N1329, N32, N1171, N510);
nand NAND3 (N1336, N1331, N910, N345);
xor XOR2 (N1337, N1332, N455);
buf BUF1 (N1338, N1333);
nand NAND4 (N1339, N1335, N800, N608, N166);
or OR3 (N1340, N1336, N827, N1078);
nor NOR3 (N1341, N1283, N954, N705);
and AND4 (N1342, N1330, N938, N700, N1216);
or OR2 (N1343, N1305, N564);
nor NOR4 (N1344, N1342, N638, N520, N81);
buf BUF1 (N1345, N1327);
or OR4 (N1346, N1343, N1281, N1144, N1309);
and AND2 (N1347, N1337, N238);
and AND3 (N1348, N1347, N822, N1270);
or OR2 (N1349, N1344, N377);
not NOT1 (N1350, N1346);
nor NOR4 (N1351, N1341, N1267, N1244, N110);
xor XOR2 (N1352, N1318, N285);
buf BUF1 (N1353, N1352);
not NOT1 (N1354, N1353);
buf BUF1 (N1355, N1349);
buf BUF1 (N1356, N1350);
nor NOR2 (N1357, N1340, N778);
nor NOR4 (N1358, N1357, N276, N880, N504);
xor XOR2 (N1359, N1354, N42);
and AND3 (N1360, N1356, N1331, N130);
xor XOR2 (N1361, N1351, N1342);
nand NAND3 (N1362, N1338, N544, N720);
nor NOR4 (N1363, N1345, N220, N525, N132);
nor NOR3 (N1364, N1363, N985, N1096);
or OR4 (N1365, N1362, N926, N112, N890);
not NOT1 (N1366, N1359);
or OR3 (N1367, N1364, N1247, N567);
buf BUF1 (N1368, N1339);
and AND4 (N1369, N1348, N548, N115, N972);
nor NOR3 (N1370, N1369, N1181, N422);
and AND4 (N1371, N1358, N549, N1082, N516);
nor NOR2 (N1372, N1370, N108);
not NOT1 (N1373, N1334);
nor NOR3 (N1374, N1368, N749, N158);
or OR4 (N1375, N1361, N477, N1206, N1291);
nand NAND2 (N1376, N1366, N139);
xor XOR2 (N1377, N1371, N965);
xor XOR2 (N1378, N1375, N1305);
and AND2 (N1379, N1355, N45);
nand NAND3 (N1380, N1377, N179, N854);
not NOT1 (N1381, N1374);
nor NOR3 (N1382, N1380, N72, N1204);
and AND3 (N1383, N1376, N176, N282);
or OR3 (N1384, N1379, N349, N46);
buf BUF1 (N1385, N1373);
xor XOR2 (N1386, N1381, N1026);
not NOT1 (N1387, N1385);
and AND4 (N1388, N1387, N1219, N677, N253);
and AND4 (N1389, N1360, N36, N734, N307);
nand NAND4 (N1390, N1386, N289, N1355, N1320);
not NOT1 (N1391, N1389);
nor NOR4 (N1392, N1378, N352, N444, N26);
or OR2 (N1393, N1365, N455);
not NOT1 (N1394, N1393);
nor NOR2 (N1395, N1372, N1325);
not NOT1 (N1396, N1384);
xor XOR2 (N1397, N1395, N258);
nand NAND3 (N1398, N1392, N111, N274);
and AND3 (N1399, N1396, N208, N283);
nand NAND2 (N1400, N1399, N1381);
buf BUF1 (N1401, N1382);
nor NOR4 (N1402, N1383, N48, N1268, N696);
nor NOR4 (N1403, N1400, N1173, N1239, N1345);
and AND3 (N1404, N1398, N1335, N551);
nand NAND3 (N1405, N1390, N960, N759);
xor XOR2 (N1406, N1405, N68);
xor XOR2 (N1407, N1401, N798);
buf BUF1 (N1408, N1403);
or OR3 (N1409, N1394, N117, N1085);
and AND4 (N1410, N1388, N735, N94, N1302);
or OR3 (N1411, N1404, N421, N336);
nand NAND3 (N1412, N1408, N242, N1235);
and AND4 (N1413, N1402, N67, N954, N1293);
not NOT1 (N1414, N1413);
buf BUF1 (N1415, N1411);
xor XOR2 (N1416, N1412, N656);
not NOT1 (N1417, N1391);
and AND2 (N1418, N1367, N1115);
and AND3 (N1419, N1414, N158, N55);
or OR4 (N1420, N1407, N404, N52, N1258);
not NOT1 (N1421, N1406);
nor NOR4 (N1422, N1416, N460, N832, N506);
or OR2 (N1423, N1422, N921);
buf BUF1 (N1424, N1418);
nor NOR4 (N1425, N1419, N471, N1246, N979);
and AND2 (N1426, N1410, N915);
buf BUF1 (N1427, N1425);
xor XOR2 (N1428, N1409, N1232);
not NOT1 (N1429, N1415);
not NOT1 (N1430, N1397);
nor NOR4 (N1431, N1417, N820, N785, N114);
not NOT1 (N1432, N1429);
nand NAND2 (N1433, N1423, N442);
xor XOR2 (N1434, N1427, N739);
and AND4 (N1435, N1430, N1222, N1294, N736);
nand NAND2 (N1436, N1424, N940);
and AND2 (N1437, N1432, N1417);
and AND2 (N1438, N1431, N205);
not NOT1 (N1439, N1438);
nor NOR4 (N1440, N1436, N158, N784, N1033);
nand NAND3 (N1441, N1434, N332, N377);
xor XOR2 (N1442, N1428, N1376);
xor XOR2 (N1443, N1442, N250);
and AND4 (N1444, N1441, N376, N277, N1365);
buf BUF1 (N1445, N1421);
and AND2 (N1446, N1440, N802);
nor NOR4 (N1447, N1446, N680, N1212, N1358);
not NOT1 (N1448, N1447);
nor NOR3 (N1449, N1445, N1242, N1136);
buf BUF1 (N1450, N1439);
xor XOR2 (N1451, N1444, N1365);
or OR4 (N1452, N1448, N618, N388, N445);
xor XOR2 (N1453, N1437, N697);
or OR4 (N1454, N1452, N1217, N479, N599);
or OR4 (N1455, N1451, N1093, N786, N1222);
xor XOR2 (N1456, N1450, N294);
xor XOR2 (N1457, N1449, N1395);
nand NAND2 (N1458, N1443, N962);
nor NOR3 (N1459, N1458, N1123, N1424);
xor XOR2 (N1460, N1456, N1285);
nand NAND3 (N1461, N1454, N672, N274);
buf BUF1 (N1462, N1420);
nand NAND4 (N1463, N1426, N775, N555, N65);
and AND3 (N1464, N1463, N462, N520);
buf BUF1 (N1465, N1461);
and AND2 (N1466, N1465, N879);
or OR2 (N1467, N1460, N1133);
or OR4 (N1468, N1435, N854, N1437, N464);
or OR2 (N1469, N1455, N844);
buf BUF1 (N1470, N1469);
nand NAND2 (N1471, N1468, N856);
not NOT1 (N1472, N1453);
xor XOR2 (N1473, N1471, N1220);
not NOT1 (N1474, N1464);
nand NAND4 (N1475, N1467, N1436, N1193, N721);
nor NOR2 (N1476, N1466, N525);
nand NAND3 (N1477, N1459, N532, N396);
or OR2 (N1478, N1477, N827);
buf BUF1 (N1479, N1462);
nor NOR2 (N1480, N1470, N873);
not NOT1 (N1481, N1478);
nor NOR4 (N1482, N1472, N434, N114, N619);
not NOT1 (N1483, N1479);
not NOT1 (N1484, N1475);
and AND4 (N1485, N1476, N711, N1217, N831);
xor XOR2 (N1486, N1457, N907);
nand NAND4 (N1487, N1486, N1261, N1336, N743);
and AND2 (N1488, N1473, N59);
not NOT1 (N1489, N1482);
and AND3 (N1490, N1483, N705, N353);
buf BUF1 (N1491, N1484);
nand NAND4 (N1492, N1480, N641, N402, N886);
buf BUF1 (N1493, N1492);
and AND2 (N1494, N1491, N636);
xor XOR2 (N1495, N1487, N1119);
xor XOR2 (N1496, N1495, N258);
buf BUF1 (N1497, N1481);
xor XOR2 (N1498, N1490, N1053);
and AND3 (N1499, N1433, N905, N930);
and AND2 (N1500, N1496, N1131);
nand NAND3 (N1501, N1489, N1178, N445);
not NOT1 (N1502, N1499);
buf BUF1 (N1503, N1501);
nor NOR3 (N1504, N1494, N613, N1098);
buf BUF1 (N1505, N1488);
xor XOR2 (N1506, N1504, N74);
and AND2 (N1507, N1502, N1142);
xor XOR2 (N1508, N1493, N205);
nor NOR3 (N1509, N1474, N990, N31);
buf BUF1 (N1510, N1505);
or OR2 (N1511, N1508, N144);
buf BUF1 (N1512, N1500);
xor XOR2 (N1513, N1509, N350);
and AND2 (N1514, N1498, N517);
and AND3 (N1515, N1512, N441, N1030);
buf BUF1 (N1516, N1510);
and AND3 (N1517, N1506, N142, N1387);
and AND3 (N1518, N1485, N1507, N1120);
or OR4 (N1519, N1462, N261, N1360, N390);
or OR2 (N1520, N1517, N807);
nand NAND2 (N1521, N1513, N1411);
or OR2 (N1522, N1519, N1510);
nor NOR3 (N1523, N1516, N503, N1117);
not NOT1 (N1524, N1518);
buf BUF1 (N1525, N1524);
not NOT1 (N1526, N1523);
nor NOR2 (N1527, N1520, N371);
not NOT1 (N1528, N1497);
nand NAND3 (N1529, N1514, N303, N1509);
nor NOR3 (N1530, N1525, N896, N696);
or OR4 (N1531, N1522, N1186, N807, N448);
nand NAND4 (N1532, N1528, N488, N1426, N129);
or OR4 (N1533, N1526, N402, N772, N698);
xor XOR2 (N1534, N1530, N947);
and AND3 (N1535, N1521, N1108, N341);
nor NOR2 (N1536, N1511, N71);
buf BUF1 (N1537, N1535);
nand NAND2 (N1538, N1503, N216);
and AND4 (N1539, N1532, N692, N1175, N1023);
or OR4 (N1540, N1515, N20, N551, N845);
nand NAND4 (N1541, N1538, N1504, N52, N1258);
xor XOR2 (N1542, N1536, N1270);
buf BUF1 (N1543, N1529);
or OR4 (N1544, N1542, N1536, N1026, N82);
nor NOR2 (N1545, N1543, N109);
not NOT1 (N1546, N1541);
buf BUF1 (N1547, N1531);
or OR4 (N1548, N1533, N1049, N491, N1230);
not NOT1 (N1549, N1545);
nand NAND2 (N1550, N1549, N1017);
nor NOR2 (N1551, N1539, N940);
not NOT1 (N1552, N1548);
buf BUF1 (N1553, N1547);
not NOT1 (N1554, N1553);
nor NOR2 (N1555, N1552, N890);
xor XOR2 (N1556, N1527, N607);
not NOT1 (N1557, N1544);
or OR3 (N1558, N1546, N484, N583);
or OR3 (N1559, N1534, N1291, N1266);
or OR2 (N1560, N1551, N1073);
buf BUF1 (N1561, N1560);
or OR2 (N1562, N1557, N732);
xor XOR2 (N1563, N1562, N1140);
nand NAND4 (N1564, N1550, N109, N1544, N1202);
and AND2 (N1565, N1561, N203);
and AND3 (N1566, N1559, N1318, N1326);
nand NAND4 (N1567, N1555, N4, N336, N1536);
xor XOR2 (N1568, N1565, N803);
nand NAND2 (N1569, N1556, N148);
nand NAND2 (N1570, N1564, N543);
buf BUF1 (N1571, N1569);
not NOT1 (N1572, N1566);
not NOT1 (N1573, N1572);
nand NAND3 (N1574, N1558, N1498, N1191);
nand NAND4 (N1575, N1537, N766, N1258, N852);
nand NAND2 (N1576, N1563, N1557);
or OR2 (N1577, N1573, N246);
buf BUF1 (N1578, N1540);
nand NAND4 (N1579, N1574, N840, N1576, N202);
and AND2 (N1580, N450, N460);
xor XOR2 (N1581, N1575, N805);
and AND4 (N1582, N1580, N862, N886, N1381);
nor NOR4 (N1583, N1554, N561, N790, N995);
nor NOR3 (N1584, N1581, N591, N545);
xor XOR2 (N1585, N1582, N1462);
nor NOR4 (N1586, N1584, N940, N1102, N1353);
buf BUF1 (N1587, N1571);
and AND4 (N1588, N1583, N650, N1453, N1180);
not NOT1 (N1589, N1587);
and AND3 (N1590, N1589, N481, N1156);
and AND4 (N1591, N1586, N883, N1213, N714);
and AND4 (N1592, N1585, N986, N951, N389);
and AND2 (N1593, N1577, N848);
nand NAND3 (N1594, N1568, N978, N868);
nor NOR4 (N1595, N1588, N182, N784, N858);
and AND2 (N1596, N1594, N605);
xor XOR2 (N1597, N1567, N1057);
xor XOR2 (N1598, N1592, N1124);
or OR2 (N1599, N1593, N588);
xor XOR2 (N1600, N1590, N139);
or OR3 (N1601, N1579, N449, N348);
or OR3 (N1602, N1595, N1524, N785);
xor XOR2 (N1603, N1570, N55);
or OR3 (N1604, N1578, N150, N1456);
xor XOR2 (N1605, N1597, N188);
or OR2 (N1606, N1600, N315);
buf BUF1 (N1607, N1606);
or OR2 (N1608, N1601, N155);
not NOT1 (N1609, N1604);
and AND3 (N1610, N1609, N941, N840);
nand NAND4 (N1611, N1608, N65, N1471, N753);
and AND4 (N1612, N1610, N1073, N566, N728);
not NOT1 (N1613, N1612);
or OR4 (N1614, N1596, N956, N1073, N1456);
xor XOR2 (N1615, N1603, N776);
xor XOR2 (N1616, N1602, N405);
xor XOR2 (N1617, N1591, N241);
buf BUF1 (N1618, N1617);
nand NAND3 (N1619, N1616, N434, N956);
nor NOR3 (N1620, N1614, N1365, N1039);
nand NAND2 (N1621, N1613, N1296);
nand NAND3 (N1622, N1619, N906, N844);
nor NOR3 (N1623, N1622, N401, N309);
nor NOR4 (N1624, N1621, N1141, N572, N1012);
not NOT1 (N1625, N1611);
and AND3 (N1626, N1620, N42, N421);
xor XOR2 (N1627, N1598, N276);
or OR2 (N1628, N1615, N1164);
nor NOR3 (N1629, N1626, N128, N1464);
buf BUF1 (N1630, N1624);
not NOT1 (N1631, N1627);
nor NOR4 (N1632, N1628, N1543, N264, N206);
or OR2 (N1633, N1625, N440);
and AND3 (N1634, N1633, N376, N1236);
or OR3 (N1635, N1630, N60, N1129);
and AND3 (N1636, N1605, N1190, N1015);
nor NOR4 (N1637, N1634, N665, N869, N1485);
not NOT1 (N1638, N1632);
nand NAND2 (N1639, N1636, N242);
nand NAND2 (N1640, N1631, N688);
nand NAND4 (N1641, N1618, N1355, N1140, N1588);
buf BUF1 (N1642, N1639);
xor XOR2 (N1643, N1637, N557);
buf BUF1 (N1644, N1641);
nor NOR3 (N1645, N1643, N1159, N510);
nor NOR2 (N1646, N1640, N777);
and AND4 (N1647, N1599, N316, N566, N1303);
or OR2 (N1648, N1644, N279);
nand NAND2 (N1649, N1642, N1176);
and AND4 (N1650, N1648, N242, N522, N1564);
nor NOR3 (N1651, N1638, N1058, N700);
or OR3 (N1652, N1649, N596, N1642);
not NOT1 (N1653, N1645);
nor NOR2 (N1654, N1629, N250);
xor XOR2 (N1655, N1646, N52);
xor XOR2 (N1656, N1654, N231);
nand NAND3 (N1657, N1623, N1195, N1262);
xor XOR2 (N1658, N1647, N1547);
nor NOR4 (N1659, N1655, N543, N487, N735);
xor XOR2 (N1660, N1657, N1418);
xor XOR2 (N1661, N1635, N651);
nand NAND3 (N1662, N1651, N645, N427);
nor NOR2 (N1663, N1656, N489);
nand NAND4 (N1664, N1650, N1438, N1485, N849);
not NOT1 (N1665, N1658);
xor XOR2 (N1666, N1607, N170);
buf BUF1 (N1667, N1665);
or OR3 (N1668, N1664, N369, N620);
nand NAND3 (N1669, N1653, N1522, N1664);
nor NOR2 (N1670, N1669, N1258);
buf BUF1 (N1671, N1662);
or OR3 (N1672, N1652, N784, N1153);
nor NOR2 (N1673, N1670, N1586);
not NOT1 (N1674, N1672);
not NOT1 (N1675, N1666);
or OR2 (N1676, N1660, N416);
nor NOR3 (N1677, N1671, N244, N753);
or OR4 (N1678, N1668, N509, N595, N238);
buf BUF1 (N1679, N1667);
not NOT1 (N1680, N1674);
and AND4 (N1681, N1678, N1045, N693, N1592);
or OR4 (N1682, N1661, N231, N156, N192);
buf BUF1 (N1683, N1659);
nor NOR4 (N1684, N1673, N620, N209, N1430);
nor NOR3 (N1685, N1675, N1328, N1621);
or OR4 (N1686, N1676, N323, N1545, N973);
buf BUF1 (N1687, N1686);
buf BUF1 (N1688, N1683);
nor NOR2 (N1689, N1685, N521);
not NOT1 (N1690, N1689);
xor XOR2 (N1691, N1687, N1420);
not NOT1 (N1692, N1680);
or OR2 (N1693, N1663, N1176);
not NOT1 (N1694, N1679);
xor XOR2 (N1695, N1688, N1382);
or OR4 (N1696, N1677, N1205, N501, N133);
nand NAND3 (N1697, N1693, N104, N172);
xor XOR2 (N1698, N1681, N959);
buf BUF1 (N1699, N1692);
nand NAND2 (N1700, N1684, N19);
xor XOR2 (N1701, N1690, N1188);
not NOT1 (N1702, N1694);
not NOT1 (N1703, N1699);
nand NAND2 (N1704, N1697, N1071);
or OR2 (N1705, N1691, N62);
nand NAND3 (N1706, N1702, N375, N603);
xor XOR2 (N1707, N1704, N1262);
xor XOR2 (N1708, N1705, N778);
xor XOR2 (N1709, N1701, N1417);
not NOT1 (N1710, N1708);
not NOT1 (N1711, N1698);
nand NAND4 (N1712, N1703, N1532, N831, N893);
nand NAND4 (N1713, N1706, N756, N1597, N941);
and AND2 (N1714, N1695, N1355);
nor NOR3 (N1715, N1696, N1711, N1457);
nor NOR2 (N1716, N1260, N254);
buf BUF1 (N1717, N1710);
xor XOR2 (N1718, N1714, N345);
nand NAND3 (N1719, N1712, N234, N626);
and AND4 (N1720, N1715, N1311, N984, N1384);
xor XOR2 (N1721, N1700, N1585);
or OR3 (N1722, N1718, N1400, N719);
or OR4 (N1723, N1721, N349, N53, N38);
nor NOR3 (N1724, N1709, N1438, N1555);
nand NAND3 (N1725, N1682, N1102, N817);
xor XOR2 (N1726, N1719, N124);
not NOT1 (N1727, N1713);
or OR3 (N1728, N1717, N689, N844);
buf BUF1 (N1729, N1722);
not NOT1 (N1730, N1727);
not NOT1 (N1731, N1723);
nand NAND4 (N1732, N1725, N1653, N73, N127);
nor NOR2 (N1733, N1720, N74);
buf BUF1 (N1734, N1726);
xor XOR2 (N1735, N1707, N223);
nor NOR2 (N1736, N1730, N264);
and AND4 (N1737, N1736, N749, N1725, N1035);
nand NAND2 (N1738, N1724, N352);
buf BUF1 (N1739, N1716);
not NOT1 (N1740, N1738);
buf BUF1 (N1741, N1733);
not NOT1 (N1742, N1740);
not NOT1 (N1743, N1728);
buf BUF1 (N1744, N1734);
nand NAND3 (N1745, N1729, N1116, N414);
or OR2 (N1746, N1745, N255);
not NOT1 (N1747, N1737);
nor NOR4 (N1748, N1731, N721, N1634, N1529);
buf BUF1 (N1749, N1744);
nor NOR2 (N1750, N1739, N498);
or OR3 (N1751, N1749, N408, N997);
and AND4 (N1752, N1732, N901, N71, N987);
nand NAND4 (N1753, N1751, N1684, N1233, N714);
nand NAND3 (N1754, N1746, N1232, N270);
nor NOR3 (N1755, N1743, N473, N1093);
and AND3 (N1756, N1752, N555, N774);
nor NOR4 (N1757, N1741, N1322, N601, N555);
or OR2 (N1758, N1747, N813);
nor NOR4 (N1759, N1753, N1748, N1404, N275);
nand NAND3 (N1760, N1686, N202, N1051);
nand NAND3 (N1761, N1754, N219, N493);
or OR2 (N1762, N1742, N1339);
xor XOR2 (N1763, N1755, N1172);
xor XOR2 (N1764, N1763, N76);
xor XOR2 (N1765, N1762, N66);
or OR2 (N1766, N1764, N283);
xor XOR2 (N1767, N1757, N111);
not NOT1 (N1768, N1761);
xor XOR2 (N1769, N1766, N821);
nor NOR2 (N1770, N1768, N1736);
nor NOR3 (N1771, N1735, N507, N663);
not NOT1 (N1772, N1758);
nor NOR3 (N1773, N1756, N1220, N1741);
nor NOR3 (N1774, N1759, N861, N1488);
nand NAND4 (N1775, N1771, N352, N1691, N1508);
xor XOR2 (N1776, N1774, N1658);
not NOT1 (N1777, N1776);
not NOT1 (N1778, N1770);
and AND3 (N1779, N1769, N496, N334);
and AND4 (N1780, N1767, N1217, N1118, N812);
buf BUF1 (N1781, N1773);
buf BUF1 (N1782, N1778);
or OR3 (N1783, N1779, N1284, N91);
nand NAND3 (N1784, N1765, N1075, N1432);
or OR3 (N1785, N1777, N1249, N1700);
xor XOR2 (N1786, N1772, N1246);
not NOT1 (N1787, N1785);
nand NAND4 (N1788, N1784, N6, N1416, N1380);
or OR2 (N1789, N1782, N597);
not NOT1 (N1790, N1780);
nor NOR2 (N1791, N1775, N688);
and AND3 (N1792, N1783, N1401, N5);
or OR4 (N1793, N1792, N939, N1538, N1752);
nor NOR4 (N1794, N1786, N1387, N664, N743);
and AND3 (N1795, N1781, N836, N723);
buf BUF1 (N1796, N1760);
xor XOR2 (N1797, N1795, N674);
xor XOR2 (N1798, N1791, N427);
nor NOR4 (N1799, N1796, N368, N641, N411);
nand NAND3 (N1800, N1788, N1522, N313);
or OR4 (N1801, N1797, N893, N1788, N703);
or OR2 (N1802, N1800, N1679);
xor XOR2 (N1803, N1801, N1022);
xor XOR2 (N1804, N1802, N21);
not NOT1 (N1805, N1803);
xor XOR2 (N1806, N1805, N1797);
nand NAND2 (N1807, N1798, N159);
nor NOR4 (N1808, N1750, N405, N902, N1449);
nor NOR3 (N1809, N1787, N596, N1504);
not NOT1 (N1810, N1804);
or OR2 (N1811, N1794, N802);
nor NOR4 (N1812, N1790, N1529, N498, N886);
and AND3 (N1813, N1809, N1130, N624);
nor NOR2 (N1814, N1789, N1638);
and AND3 (N1815, N1814, N1157, N133);
xor XOR2 (N1816, N1813, N1136);
xor XOR2 (N1817, N1799, N1402);
not NOT1 (N1818, N1807);
and AND3 (N1819, N1793, N1294, N357);
nand NAND3 (N1820, N1819, N867, N490);
nor NOR3 (N1821, N1808, N1359, N793);
buf BUF1 (N1822, N1810);
buf BUF1 (N1823, N1818);
xor XOR2 (N1824, N1811, N1157);
and AND4 (N1825, N1822, N33, N1071, N1341);
buf BUF1 (N1826, N1816);
not NOT1 (N1827, N1806);
nand NAND3 (N1828, N1817, N1086, N1627);
and AND3 (N1829, N1820, N1120, N765);
buf BUF1 (N1830, N1827);
nor NOR2 (N1831, N1826, N983);
and AND4 (N1832, N1829, N1170, N94, N1621);
not NOT1 (N1833, N1815);
xor XOR2 (N1834, N1832, N155);
not NOT1 (N1835, N1828);
and AND3 (N1836, N1831, N521, N505);
nand NAND3 (N1837, N1835, N1595, N194);
not NOT1 (N1838, N1825);
buf BUF1 (N1839, N1821);
buf BUF1 (N1840, N1823);
and AND2 (N1841, N1812, N765);
buf BUF1 (N1842, N1841);
xor XOR2 (N1843, N1824, N1428);
and AND2 (N1844, N1836, N1826);
or OR2 (N1845, N1838, N1541);
buf BUF1 (N1846, N1842);
xor XOR2 (N1847, N1830, N1817);
nor NOR4 (N1848, N1844, N621, N393, N1798);
not NOT1 (N1849, N1833);
nor NOR3 (N1850, N1846, N3, N833);
and AND4 (N1851, N1850, N527, N1310, N1145);
and AND4 (N1852, N1840, N1623, N1161, N1129);
nor NOR3 (N1853, N1837, N534, N750);
nand NAND4 (N1854, N1851, N1019, N1104, N1434);
or OR3 (N1855, N1843, N260, N1475);
and AND4 (N1856, N1849, N1224, N1120, N1278);
nor NOR4 (N1857, N1848, N670, N311, N284);
or OR2 (N1858, N1857, N1732);
nor NOR3 (N1859, N1847, N1057, N1434);
and AND4 (N1860, N1845, N1797, N563, N169);
not NOT1 (N1861, N1855);
nand NAND2 (N1862, N1861, N425);
not NOT1 (N1863, N1854);
nor NOR2 (N1864, N1858, N498);
and AND3 (N1865, N1834, N779, N272);
or OR3 (N1866, N1856, N1696, N253);
and AND4 (N1867, N1852, N1082, N366, N221);
nor NOR2 (N1868, N1859, N801);
or OR4 (N1869, N1863, N918, N1829, N1689);
xor XOR2 (N1870, N1868, N458);
buf BUF1 (N1871, N1862);
or OR2 (N1872, N1867, N1285);
xor XOR2 (N1873, N1865, N678);
or OR4 (N1874, N1866, N384, N1227, N1522);
buf BUF1 (N1875, N1860);
buf BUF1 (N1876, N1864);
xor XOR2 (N1877, N1853, N1017);
xor XOR2 (N1878, N1871, N642);
nor NOR3 (N1879, N1869, N541, N171);
or OR3 (N1880, N1878, N1445, N664);
buf BUF1 (N1881, N1839);
nor NOR2 (N1882, N1877, N1191);
or OR2 (N1883, N1873, N1117);
xor XOR2 (N1884, N1879, N620);
nand NAND4 (N1885, N1872, N999, N1723, N1187);
xor XOR2 (N1886, N1880, N97);
xor XOR2 (N1887, N1874, N359);
nand NAND4 (N1888, N1870, N1728, N1341, N577);
xor XOR2 (N1889, N1881, N914);
nor NOR4 (N1890, N1882, N346, N924, N812);
and AND4 (N1891, N1890, N649, N414, N1312);
buf BUF1 (N1892, N1889);
or OR3 (N1893, N1884, N1008, N1606);
xor XOR2 (N1894, N1886, N1697);
buf BUF1 (N1895, N1887);
nand NAND4 (N1896, N1892, N370, N522, N1047);
and AND4 (N1897, N1876, N432, N357, N451);
buf BUF1 (N1898, N1894);
and AND3 (N1899, N1875, N937, N1100);
or OR2 (N1900, N1883, N112);
nand NAND2 (N1901, N1899, N1553);
nor NOR2 (N1902, N1891, N703);
xor XOR2 (N1903, N1885, N528);
not NOT1 (N1904, N1896);
buf BUF1 (N1905, N1904);
buf BUF1 (N1906, N1902);
buf BUF1 (N1907, N1905);
nand NAND3 (N1908, N1906, N1139, N3);
and AND3 (N1909, N1903, N459, N176);
or OR3 (N1910, N1897, N1787, N564);
not NOT1 (N1911, N1901);
xor XOR2 (N1912, N1911, N802);
and AND4 (N1913, N1907, N1882, N674, N999);
and AND2 (N1914, N1888, N1437);
nor NOR4 (N1915, N1893, N719, N1397, N1625);
or OR2 (N1916, N1895, N1088);
not NOT1 (N1917, N1913);
and AND2 (N1918, N1917, N726);
not NOT1 (N1919, N1908);
buf BUF1 (N1920, N1900);
or OR4 (N1921, N1916, N1056, N703, N1547);
buf BUF1 (N1922, N1914);
nor NOR2 (N1923, N1919, N461);
buf BUF1 (N1924, N1915);
xor XOR2 (N1925, N1922, N1316);
buf BUF1 (N1926, N1909);
not NOT1 (N1927, N1926);
or OR4 (N1928, N1924, N1609, N858, N1032);
nor NOR2 (N1929, N1921, N699);
nand NAND3 (N1930, N1927, N742, N1886);
not NOT1 (N1931, N1929);
and AND3 (N1932, N1923, N1121, N1064);
and AND2 (N1933, N1931, N1634);
buf BUF1 (N1934, N1898);
xor XOR2 (N1935, N1932, N197);
not NOT1 (N1936, N1933);
nor NOR3 (N1937, N1910, N1326, N1153);
xor XOR2 (N1938, N1920, N16);
nand NAND3 (N1939, N1925, N55, N80);
nor NOR2 (N1940, N1930, N230);
and AND3 (N1941, N1935, N1735, N1688);
not NOT1 (N1942, N1918);
nand NAND4 (N1943, N1939, N1398, N1075, N396);
xor XOR2 (N1944, N1928, N1615);
xor XOR2 (N1945, N1912, N1293);
nor NOR4 (N1946, N1945, N1501, N429, N968);
not NOT1 (N1947, N1944);
or OR4 (N1948, N1943, N51, N129, N213);
nand NAND4 (N1949, N1936, N35, N1726, N839);
buf BUF1 (N1950, N1941);
xor XOR2 (N1951, N1949, N602);
xor XOR2 (N1952, N1951, N627);
not NOT1 (N1953, N1942);
not NOT1 (N1954, N1950);
not NOT1 (N1955, N1938);
and AND4 (N1956, N1937, N1625, N1092, N1182);
buf BUF1 (N1957, N1955);
or OR3 (N1958, N1957, N1448, N1135);
xor XOR2 (N1959, N1940, N1552);
xor XOR2 (N1960, N1952, N458);
nand NAND3 (N1961, N1960, N1327, N1131);
or OR4 (N1962, N1934, N1022, N451, N830);
xor XOR2 (N1963, N1961, N519);
and AND3 (N1964, N1956, N158, N1347);
and AND4 (N1965, N1946, N1036, N263, N956);
nand NAND4 (N1966, N1954, N190, N850, N1497);
or OR4 (N1967, N1966, N803, N105, N1921);
or OR2 (N1968, N1953, N107);
nand NAND2 (N1969, N1959, N69);
or OR3 (N1970, N1948, N1962, N1674);
nor NOR3 (N1971, N274, N1601, N919);
or OR3 (N1972, N1971, N801, N665);
not NOT1 (N1973, N1947);
xor XOR2 (N1974, N1970, N1360);
nand NAND3 (N1975, N1968, N640, N1179);
xor XOR2 (N1976, N1969, N1069);
nor NOR3 (N1977, N1974, N401, N820);
xor XOR2 (N1978, N1976, N81);
or OR3 (N1979, N1978, N638, N235);
nor NOR2 (N1980, N1973, N1867);
not NOT1 (N1981, N1967);
nand NAND4 (N1982, N1963, N1948, N1558, N1926);
not NOT1 (N1983, N1982);
nand NAND3 (N1984, N1975, N1208, N948);
buf BUF1 (N1985, N1958);
buf BUF1 (N1986, N1983);
nor NOR2 (N1987, N1965, N1642);
nor NOR4 (N1988, N1986, N1213, N1933, N1550);
buf BUF1 (N1989, N1977);
not NOT1 (N1990, N1988);
buf BUF1 (N1991, N1987);
or OR3 (N1992, N1964, N1321, N1909);
nand NAND3 (N1993, N1979, N673, N1893);
xor XOR2 (N1994, N1985, N1268);
nand NAND2 (N1995, N1993, N537);
buf BUF1 (N1996, N1990);
and AND4 (N1997, N1972, N451, N119, N1565);
nor NOR3 (N1998, N1989, N995, N1677);
buf BUF1 (N1999, N1991);
xor XOR2 (N2000, N1984, N1227);
and AND4 (N2001, N1981, N1288, N365, N1773);
or OR2 (N2002, N1994, N1072);
xor XOR2 (N2003, N1996, N853);
or OR4 (N2004, N2000, N1625, N1576, N25);
not NOT1 (N2005, N2003);
not NOT1 (N2006, N1980);
nor NOR3 (N2007, N2006, N1677, N1894);
and AND2 (N2008, N2007, N459);
buf BUF1 (N2009, N1997);
xor XOR2 (N2010, N2009, N153);
and AND4 (N2011, N2010, N707, N308, N59);
nand NAND2 (N2012, N2001, N197);
nor NOR3 (N2013, N2002, N1953, N1742);
or OR2 (N2014, N1999, N1567);
buf BUF1 (N2015, N2013);
buf BUF1 (N2016, N2011);
xor XOR2 (N2017, N2016, N1419);
nor NOR4 (N2018, N2014, N181, N213, N1125);
and AND3 (N2019, N1992, N1328, N285);
or OR2 (N2020, N2017, N1535);
xor XOR2 (N2021, N2015, N976);
buf BUF1 (N2022, N1995);
buf BUF1 (N2023, N2004);
buf BUF1 (N2024, N2021);
not NOT1 (N2025, N2023);
not NOT1 (N2026, N2018);
or OR4 (N2027, N2019, N1339, N496, N1255);
nor NOR4 (N2028, N2012, N1494, N1242, N612);
buf BUF1 (N2029, N2024);
xor XOR2 (N2030, N2026, N2010);
and AND3 (N2031, N1998, N1280, N1468);
or OR3 (N2032, N2008, N686, N978);
buf BUF1 (N2033, N2020);
and AND3 (N2034, N2029, N1008, N729);
or OR4 (N2035, N2033, N243, N887, N1033);
not NOT1 (N2036, N2025);
not NOT1 (N2037, N2036);
buf BUF1 (N2038, N2037);
nand NAND4 (N2039, N2027, N1451, N620, N497);
not NOT1 (N2040, N2028);
buf BUF1 (N2041, N2038);
or OR3 (N2042, N2041, N758, N214);
nand NAND3 (N2043, N2030, N335, N1711);
or OR4 (N2044, N2042, N169, N374, N1427);
or OR4 (N2045, N2040, N45, N1610, N428);
or OR3 (N2046, N2044, N1020, N1731);
and AND4 (N2047, N2022, N691, N371, N1611);
nor NOR2 (N2048, N2045, N1770);
xor XOR2 (N2049, N2048, N1227);
not NOT1 (N2050, N2005);
or OR4 (N2051, N2034, N1701, N1859, N1501);
buf BUF1 (N2052, N2047);
and AND4 (N2053, N2051, N1577, N517, N1660);
or OR4 (N2054, N2035, N187, N1780, N976);
and AND2 (N2055, N2050, N725);
or OR4 (N2056, N2032, N1644, N1216, N280);
buf BUF1 (N2057, N2054);
xor XOR2 (N2058, N2046, N961);
buf BUF1 (N2059, N2057);
xor XOR2 (N2060, N2039, N667);
not NOT1 (N2061, N2058);
or OR4 (N2062, N2052, N977, N316, N1924);
nor NOR3 (N2063, N2053, N600, N310);
xor XOR2 (N2064, N2043, N327);
xor XOR2 (N2065, N2031, N1815);
nor NOR2 (N2066, N2062, N1699);
buf BUF1 (N2067, N2064);
and AND3 (N2068, N2061, N1933, N49);
or OR3 (N2069, N2066, N713, N555);
and AND3 (N2070, N2060, N1206, N1030);
or OR4 (N2071, N2067, N1828, N391, N1916);
or OR4 (N2072, N2068, N1332, N1318, N676);
nand NAND3 (N2073, N2063, N1638, N1017);
buf BUF1 (N2074, N2071);
nor NOR3 (N2075, N2056, N1845, N271);
and AND2 (N2076, N2075, N1148);
buf BUF1 (N2077, N2055);
and AND4 (N2078, N2069, N118, N974, N1775);
and AND3 (N2079, N2049, N838, N1372);
not NOT1 (N2080, N2070);
nand NAND4 (N2081, N2074, N907, N1991, N1671);
nand NAND2 (N2082, N2078, N1619);
xor XOR2 (N2083, N2082, N2071);
and AND4 (N2084, N2080, N1377, N364, N414);
and AND2 (N2085, N2077, N171);
or OR2 (N2086, N2072, N1823);
nand NAND3 (N2087, N2059, N1478, N429);
not NOT1 (N2088, N2087);
nor NOR3 (N2089, N2079, N1944, N915);
not NOT1 (N2090, N2084);
nor NOR3 (N2091, N2088, N1576, N1619);
nor NOR2 (N2092, N2086, N1529);
or OR3 (N2093, N2092, N1327, N2054);
or OR2 (N2094, N2073, N1252);
nor NOR4 (N2095, N2076, N554, N5, N804);
xor XOR2 (N2096, N2091, N818);
or OR2 (N2097, N2081, N25);
xor XOR2 (N2098, N2095, N1078);
xor XOR2 (N2099, N2098, N1355);
buf BUF1 (N2100, N2094);
not NOT1 (N2101, N2083);
not NOT1 (N2102, N2096);
and AND4 (N2103, N2085, N169, N267, N195);
or OR3 (N2104, N2100, N1342, N470);
nor NOR2 (N2105, N2089, N2051);
buf BUF1 (N2106, N2090);
xor XOR2 (N2107, N2104, N870);
and AND3 (N2108, N2101, N1709, N1265);
or OR2 (N2109, N2105, N1128);
buf BUF1 (N2110, N2097);
nand NAND2 (N2111, N2107, N876);
buf BUF1 (N2112, N2108);
or OR4 (N2113, N2106, N1626, N622, N158);
xor XOR2 (N2114, N2110, N1485);
not NOT1 (N2115, N2093);
and AND4 (N2116, N2111, N586, N628, N161);
xor XOR2 (N2117, N2114, N387);
buf BUF1 (N2118, N2117);
nand NAND3 (N2119, N2112, N789, N1281);
nor NOR3 (N2120, N2102, N1270, N608);
buf BUF1 (N2121, N2115);
and AND2 (N2122, N2118, N2117);
not NOT1 (N2123, N2103);
and AND4 (N2124, N2113, N1027, N2069, N553);
buf BUF1 (N2125, N2121);
and AND2 (N2126, N2099, N1009);
nor NOR4 (N2127, N2109, N945, N47, N707);
nand NAND2 (N2128, N2125, N595);
xor XOR2 (N2129, N2124, N148);
or OR3 (N2130, N2127, N1776, N463);
xor XOR2 (N2131, N2119, N36);
and AND3 (N2132, N2130, N247, N1502);
xor XOR2 (N2133, N2131, N1266);
or OR4 (N2134, N2126, N1506, N734, N715);
not NOT1 (N2135, N2132);
xor XOR2 (N2136, N2133, N945);
or OR2 (N2137, N2122, N517);
and AND3 (N2138, N2136, N133, N864);
buf BUF1 (N2139, N2116);
and AND3 (N2140, N2137, N1714, N1547);
buf BUF1 (N2141, N2135);
xor XOR2 (N2142, N2120, N1965);
nor NOR3 (N2143, N2128, N1748, N1404);
nand NAND3 (N2144, N2134, N619, N92);
and AND3 (N2145, N2140, N1586, N1833);
or OR3 (N2146, N2065, N1900, N680);
nand NAND4 (N2147, N2144, N1189, N1639, N1881);
buf BUF1 (N2148, N2129);
or OR4 (N2149, N2143, N2042, N1871, N81);
not NOT1 (N2150, N2142);
buf BUF1 (N2151, N2149);
buf BUF1 (N2152, N2139);
or OR4 (N2153, N2145, N1895, N975, N114);
xor XOR2 (N2154, N2150, N1763);
xor XOR2 (N2155, N2154, N695);
xor XOR2 (N2156, N2146, N647);
xor XOR2 (N2157, N2148, N935);
not NOT1 (N2158, N2151);
and AND4 (N2159, N2141, N1162, N1294, N97);
and AND2 (N2160, N2155, N257);
nand NAND3 (N2161, N2123, N116, N1049);
or OR3 (N2162, N2138, N557, N90);
or OR3 (N2163, N2147, N1247, N158);
not NOT1 (N2164, N2160);
not NOT1 (N2165, N2156);
buf BUF1 (N2166, N2164);
nor NOR4 (N2167, N2158, N344, N320, N1477);
buf BUF1 (N2168, N2161);
buf BUF1 (N2169, N2166);
xor XOR2 (N2170, N2159, N428);
nand NAND3 (N2171, N2162, N1731, N330);
xor XOR2 (N2172, N2153, N78);
buf BUF1 (N2173, N2172);
and AND3 (N2174, N2168, N1371, N199);
buf BUF1 (N2175, N2173);
xor XOR2 (N2176, N2167, N285);
or OR3 (N2177, N2163, N2009, N1054);
nand NAND3 (N2178, N2165, N1644, N603);
xor XOR2 (N2179, N2171, N2076);
xor XOR2 (N2180, N2157, N571);
buf BUF1 (N2181, N2175);
and AND3 (N2182, N2179, N975, N1263);
or OR2 (N2183, N2174, N721);
buf BUF1 (N2184, N2169);
nand NAND2 (N2185, N2180, N1470);
or OR2 (N2186, N2152, N1710);
nor NOR4 (N2187, N2177, N417, N908, N985);
nor NOR2 (N2188, N2182, N1073);
xor XOR2 (N2189, N2188, N1208);
xor XOR2 (N2190, N2187, N760);
not NOT1 (N2191, N2181);
not NOT1 (N2192, N2184);
xor XOR2 (N2193, N2176, N1506);
buf BUF1 (N2194, N2178);
buf BUF1 (N2195, N2192);
or OR2 (N2196, N2193, N2164);
and AND2 (N2197, N2194, N1872);
xor XOR2 (N2198, N2190, N830);
or OR2 (N2199, N2183, N904);
xor XOR2 (N2200, N2195, N108);
not NOT1 (N2201, N2191);
xor XOR2 (N2202, N2186, N959);
xor XOR2 (N2203, N2201, N1276);
not NOT1 (N2204, N2185);
xor XOR2 (N2205, N2197, N10);
nand NAND2 (N2206, N2196, N670);
nand NAND4 (N2207, N2170, N1974, N86, N146);
or OR3 (N2208, N2189, N159, N1887);
nand NAND3 (N2209, N2207, N1305, N1852);
and AND4 (N2210, N2209, N1338, N517, N414);
not NOT1 (N2211, N2200);
nand NAND3 (N2212, N2206, N832, N1234);
nand NAND4 (N2213, N2212, N1750, N1737, N40);
nand NAND4 (N2214, N2211, N1130, N1031, N916);
nor NOR2 (N2215, N2214, N106);
buf BUF1 (N2216, N2210);
xor XOR2 (N2217, N2205, N416);
buf BUF1 (N2218, N2202);
nand NAND3 (N2219, N2217, N356, N1112);
buf BUF1 (N2220, N2216);
and AND3 (N2221, N2198, N494, N451);
nand NAND2 (N2222, N2204, N124);
buf BUF1 (N2223, N2218);
or OR4 (N2224, N2199, N1667, N550, N1267);
xor XOR2 (N2225, N2222, N1871);
not NOT1 (N2226, N2224);
and AND2 (N2227, N2226, N423);
or OR3 (N2228, N2219, N480, N474);
buf BUF1 (N2229, N2228);
nor NOR4 (N2230, N2229, N1411, N1161, N1166);
buf BUF1 (N2231, N2213);
and AND2 (N2232, N2225, N178);
nand NAND2 (N2233, N2230, N1136);
buf BUF1 (N2234, N2233);
and AND4 (N2235, N2203, N2115, N2171, N1168);
xor XOR2 (N2236, N2232, N777);
buf BUF1 (N2237, N2223);
or OR3 (N2238, N2235, N91, N898);
or OR3 (N2239, N2215, N752, N404);
buf BUF1 (N2240, N2237);
and AND2 (N2241, N2231, N1729);
nand NAND3 (N2242, N2221, N1354, N1287);
and AND3 (N2243, N2227, N532, N936);
xor XOR2 (N2244, N2236, N1226);
not NOT1 (N2245, N2240);
or OR2 (N2246, N2243, N222);
nor NOR2 (N2247, N2244, N1172);
nand NAND4 (N2248, N2241, N1834, N497, N1758);
nand NAND4 (N2249, N2234, N367, N158, N2212);
buf BUF1 (N2250, N2246);
buf BUF1 (N2251, N2250);
and AND3 (N2252, N2208, N969, N1769);
not NOT1 (N2253, N2248);
xor XOR2 (N2254, N2238, N1763);
buf BUF1 (N2255, N2253);
nor NOR4 (N2256, N2245, N976, N1813, N563);
nand NAND2 (N2257, N2247, N1089);
xor XOR2 (N2258, N2255, N552);
xor XOR2 (N2259, N2239, N1415);
buf BUF1 (N2260, N2256);
nor NOR4 (N2261, N2257, N1602, N949, N2188);
not NOT1 (N2262, N2260);
nor NOR2 (N2263, N2252, N834);
xor XOR2 (N2264, N2249, N1713);
not NOT1 (N2265, N2242);
xor XOR2 (N2266, N2264, N631);
and AND3 (N2267, N2263, N945, N1620);
xor XOR2 (N2268, N2254, N887);
nor NOR4 (N2269, N2265, N1912, N967, N113);
nor NOR3 (N2270, N2267, N1564, N520);
xor XOR2 (N2271, N2258, N1936);
xor XOR2 (N2272, N2268, N1532);
and AND2 (N2273, N2251, N1159);
or OR4 (N2274, N2261, N313, N2199, N1007);
xor XOR2 (N2275, N2269, N2209);
and AND3 (N2276, N2274, N859, N872);
or OR2 (N2277, N2275, N1328);
not NOT1 (N2278, N2266);
nor NOR2 (N2279, N2270, N456);
not NOT1 (N2280, N2276);
nor NOR3 (N2281, N2279, N2129, N1585);
nand NAND3 (N2282, N2280, N42, N2275);
nand NAND4 (N2283, N2220, N1270, N917, N936);
buf BUF1 (N2284, N2272);
and AND2 (N2285, N2278, N951);
xor XOR2 (N2286, N2259, N500);
nor NOR2 (N2287, N2262, N975);
and AND4 (N2288, N2286, N1237, N14, N648);
and AND3 (N2289, N2288, N1913, N317);
buf BUF1 (N2290, N2277);
buf BUF1 (N2291, N2284);
not NOT1 (N2292, N2273);
not NOT1 (N2293, N2289);
or OR2 (N2294, N2283, N1130);
nand NAND4 (N2295, N2281, N34, N2005, N410);
xor XOR2 (N2296, N2285, N827);
nand NAND3 (N2297, N2271, N1925, N629);
xor XOR2 (N2298, N2292, N1628);
buf BUF1 (N2299, N2291);
or OR3 (N2300, N2294, N997, N503);
buf BUF1 (N2301, N2282);
nor NOR3 (N2302, N2293, N822, N302);
nand NAND4 (N2303, N2296, N1758, N875, N45);
and AND4 (N2304, N2290, N1510, N1048, N109);
nand NAND4 (N2305, N2300, N1581, N1802, N1244);
not NOT1 (N2306, N2301);
nor NOR2 (N2307, N2295, N1959);
not NOT1 (N2308, N2303);
or OR4 (N2309, N2304, N329, N1166, N951);
or OR4 (N2310, N2297, N1684, N2122, N1960);
not NOT1 (N2311, N2307);
and AND2 (N2312, N2302, N102);
or OR4 (N2313, N2306, N74, N1119, N1112);
buf BUF1 (N2314, N2299);
not NOT1 (N2315, N2298);
xor XOR2 (N2316, N2287, N589);
or OR4 (N2317, N2312, N2092, N1496, N1375);
or OR4 (N2318, N2308, N1823, N548, N2012);
buf BUF1 (N2319, N2305);
xor XOR2 (N2320, N2310, N2299);
xor XOR2 (N2321, N2316, N829);
and AND4 (N2322, N2319, N1872, N1233, N1824);
xor XOR2 (N2323, N2321, N640);
or OR2 (N2324, N2314, N2309);
and AND2 (N2325, N1200, N222);
nand NAND3 (N2326, N2320, N597, N267);
xor XOR2 (N2327, N2317, N691);
not NOT1 (N2328, N2324);
or OR2 (N2329, N2311, N688);
or OR2 (N2330, N2322, N47);
nand NAND3 (N2331, N2318, N1746, N1041);
buf BUF1 (N2332, N2315);
nor NOR2 (N2333, N2331, N664);
and AND4 (N2334, N2326, N307, N2168, N121);
buf BUF1 (N2335, N2325);
nand NAND3 (N2336, N2335, N1392, N20);
or OR3 (N2337, N2333, N205, N2045);
buf BUF1 (N2338, N2330);
not NOT1 (N2339, N2328);
nand NAND3 (N2340, N2339, N2032, N1073);
and AND2 (N2341, N2337, N1454);
xor XOR2 (N2342, N2334, N251);
nand NAND3 (N2343, N2332, N1617, N1390);
xor XOR2 (N2344, N2329, N913);
or OR2 (N2345, N2327, N542);
nor NOR3 (N2346, N2342, N718, N2094);
and AND3 (N2347, N2341, N1055, N1408);
nand NAND3 (N2348, N2336, N661, N427);
not NOT1 (N2349, N2347);
nand NAND3 (N2350, N2340, N1595, N13);
nand NAND3 (N2351, N2349, N1473, N1959);
nor NOR4 (N2352, N2338, N112, N430, N565);
nand NAND3 (N2353, N2345, N2081, N1395);
nor NOR3 (N2354, N2351, N1023, N1679);
and AND4 (N2355, N2323, N1683, N263, N1746);
nor NOR3 (N2356, N2343, N1765, N2305);
and AND2 (N2357, N2344, N1781);
not NOT1 (N2358, N2350);
nor NOR3 (N2359, N2358, N1077, N811);
not NOT1 (N2360, N2355);
not NOT1 (N2361, N2346);
nand NAND3 (N2362, N2354, N2055, N154);
nand NAND2 (N2363, N2359, N1657);
xor XOR2 (N2364, N2348, N1918);
nand NAND4 (N2365, N2360, N453, N2199, N1106);
nor NOR2 (N2366, N2363, N1733);
not NOT1 (N2367, N2356);
nand NAND4 (N2368, N2362, N262, N40, N2266);
xor XOR2 (N2369, N2313, N1473);
nor NOR2 (N2370, N2352, N968);
nand NAND2 (N2371, N2361, N2021);
and AND2 (N2372, N2364, N2325);
buf BUF1 (N2373, N2369);
xor XOR2 (N2374, N2372, N847);
and AND4 (N2375, N2367, N602, N215, N944);
nor NOR3 (N2376, N2357, N481, N902);
xor XOR2 (N2377, N2375, N1494);
xor XOR2 (N2378, N2371, N2110);
or OR2 (N2379, N2366, N125);
nand NAND2 (N2380, N2374, N140);
or OR3 (N2381, N2379, N1144, N1146);
xor XOR2 (N2382, N2368, N663);
nor NOR2 (N2383, N2378, N143);
not NOT1 (N2384, N2373);
nor NOR2 (N2385, N2381, N1578);
nand NAND3 (N2386, N2370, N2222, N1310);
xor XOR2 (N2387, N2365, N745);
buf BUF1 (N2388, N2385);
xor XOR2 (N2389, N2382, N654);
or OR3 (N2390, N2383, N883, N609);
not NOT1 (N2391, N2389);
or OR3 (N2392, N2387, N1885, N82);
or OR2 (N2393, N2390, N1715);
nor NOR3 (N2394, N2392, N646, N424);
xor XOR2 (N2395, N2394, N2286);
or OR3 (N2396, N2377, N197, N933);
not NOT1 (N2397, N2380);
not NOT1 (N2398, N2397);
or OR4 (N2399, N2386, N1556, N210, N273);
buf BUF1 (N2400, N2388);
xor XOR2 (N2401, N2353, N913);
not NOT1 (N2402, N2376);
buf BUF1 (N2403, N2399);
buf BUF1 (N2404, N2391);
nor NOR4 (N2405, N2401, N1143, N2131, N602);
not NOT1 (N2406, N2405);
xor XOR2 (N2407, N2395, N376);
or OR3 (N2408, N2402, N836, N633);
and AND3 (N2409, N2398, N70, N1651);
xor XOR2 (N2410, N2406, N546);
not NOT1 (N2411, N2400);
nand NAND3 (N2412, N2393, N432, N1065);
not NOT1 (N2413, N2411);
and AND4 (N2414, N2403, N178, N1461, N546);
xor XOR2 (N2415, N2409, N157);
nand NAND3 (N2416, N2415, N12, N1801);
not NOT1 (N2417, N2414);
or OR3 (N2418, N2384, N303, N2160);
buf BUF1 (N2419, N2396);
or OR2 (N2420, N2418, N800);
nor NOR2 (N2421, N2408, N922);
nand NAND4 (N2422, N2407, N432, N1656, N59);
buf BUF1 (N2423, N2404);
buf BUF1 (N2424, N2416);
buf BUF1 (N2425, N2422);
and AND3 (N2426, N2419, N632, N984);
nor NOR2 (N2427, N2412, N886);
buf BUF1 (N2428, N2427);
or OR2 (N2429, N2424, N2385);
buf BUF1 (N2430, N2428);
nor NOR3 (N2431, N2417, N944, N646);
buf BUF1 (N2432, N2430);
nand NAND4 (N2433, N2421, N949, N2199, N1954);
nand NAND4 (N2434, N2426, N1396, N609, N1311);
not NOT1 (N2435, N2433);
not NOT1 (N2436, N2431);
or OR3 (N2437, N2435, N1824, N882);
and AND3 (N2438, N2413, N38, N2085);
not NOT1 (N2439, N2425);
nand NAND3 (N2440, N2434, N768, N1441);
nand NAND2 (N2441, N2420, N2427);
and AND4 (N2442, N2429, N39, N312, N2110);
xor XOR2 (N2443, N2436, N47);
xor XOR2 (N2444, N2443, N1577);
nand NAND4 (N2445, N2432, N1324, N1712, N1577);
not NOT1 (N2446, N2441);
xor XOR2 (N2447, N2439, N2431);
xor XOR2 (N2448, N2437, N2422);
and AND4 (N2449, N2440, N1513, N2069, N2125);
nor NOR4 (N2450, N2446, N478, N2194, N594);
and AND3 (N2451, N2438, N1018, N1106);
and AND2 (N2452, N2447, N1619);
nand NAND4 (N2453, N2448, N1045, N1151, N301);
and AND2 (N2454, N2423, N525);
nand NAND4 (N2455, N2450, N30, N1547, N400);
or OR2 (N2456, N2455, N643);
and AND2 (N2457, N2445, N1187);
and AND4 (N2458, N2456, N119, N1675, N634);
or OR4 (N2459, N2449, N701, N1740, N1979);
nand NAND4 (N2460, N2410, N2172, N902, N1656);
nor NOR4 (N2461, N2451, N2340, N148, N320);
not NOT1 (N2462, N2452);
or OR4 (N2463, N2458, N1003, N2157, N1939);
not NOT1 (N2464, N2457);
and AND2 (N2465, N2463, N1199);
nand NAND3 (N2466, N2462, N96, N2088);
not NOT1 (N2467, N2466);
or OR3 (N2468, N2444, N1608, N843);
and AND4 (N2469, N2442, N1234, N529, N2377);
and AND4 (N2470, N2467, N989, N2096, N1929);
buf BUF1 (N2471, N2465);
and AND4 (N2472, N2460, N474, N197, N2329);
nand NAND4 (N2473, N2459, N247, N1663, N823);
buf BUF1 (N2474, N2454);
nor NOR2 (N2475, N2469, N2079);
and AND4 (N2476, N2453, N2250, N389, N960);
xor XOR2 (N2477, N2475, N442);
not NOT1 (N2478, N2472);
buf BUF1 (N2479, N2477);
buf BUF1 (N2480, N2464);
nor NOR3 (N2481, N2474, N1799, N1144);
not NOT1 (N2482, N2471);
not NOT1 (N2483, N2461);
not NOT1 (N2484, N2480);
nor NOR3 (N2485, N2476, N877, N582);
buf BUF1 (N2486, N2482);
and AND2 (N2487, N2473, N2196);
not NOT1 (N2488, N2486);
xor XOR2 (N2489, N2483, N136);
xor XOR2 (N2490, N2468, N2287);
nor NOR4 (N2491, N2481, N800, N653, N2064);
or OR4 (N2492, N2479, N1825, N445, N1226);
xor XOR2 (N2493, N2484, N2076);
nor NOR4 (N2494, N2490, N1369, N88, N1405);
xor XOR2 (N2495, N2470, N189);
xor XOR2 (N2496, N2494, N2118);
not NOT1 (N2497, N2485);
nor NOR2 (N2498, N2497, N684);
xor XOR2 (N2499, N2489, N657);
buf BUF1 (N2500, N2496);
and AND3 (N2501, N2487, N1040, N1285);
buf BUF1 (N2502, N2492);
and AND2 (N2503, N2493, N2360);
nor NOR3 (N2504, N2488, N1101, N172);
nand NAND2 (N2505, N2503, N125);
and AND3 (N2506, N2505, N384, N1644);
or OR4 (N2507, N2502, N1385, N1227, N2433);
buf BUF1 (N2508, N2507);
nor NOR2 (N2509, N2495, N2266);
nand NAND3 (N2510, N2508, N124, N2433);
and AND2 (N2511, N2501, N1030);
or OR4 (N2512, N2506, N2251, N523, N1125);
and AND4 (N2513, N2500, N1972, N1778, N1599);
buf BUF1 (N2514, N2478);
xor XOR2 (N2515, N2498, N1991);
nor NOR4 (N2516, N2509, N2170, N1094, N1206);
buf BUF1 (N2517, N2491);
or OR2 (N2518, N2499, N1092);
xor XOR2 (N2519, N2511, N456);
nor NOR3 (N2520, N2517, N1105, N1069);
not NOT1 (N2521, N2513);
and AND2 (N2522, N2504, N2155);
not NOT1 (N2523, N2519);
not NOT1 (N2524, N2518);
buf BUF1 (N2525, N2524);
nor NOR4 (N2526, N2523, N1802, N261, N349);
buf BUF1 (N2527, N2521);
xor XOR2 (N2528, N2520, N1340);
not NOT1 (N2529, N2515);
xor XOR2 (N2530, N2512, N95);
or OR3 (N2531, N2525, N971, N1543);
nor NOR3 (N2532, N2531, N995, N1613);
xor XOR2 (N2533, N2516, N384);
or OR2 (N2534, N2526, N246);
or OR4 (N2535, N2530, N2421, N1991, N1927);
xor XOR2 (N2536, N2528, N2290);
or OR2 (N2537, N2534, N860);
nor NOR4 (N2538, N2532, N1221, N1761, N1205);
not NOT1 (N2539, N2529);
buf BUF1 (N2540, N2536);
not NOT1 (N2541, N2514);
buf BUF1 (N2542, N2537);
buf BUF1 (N2543, N2535);
nand NAND4 (N2544, N2541, N1949, N995, N270);
nand NAND4 (N2545, N2527, N298, N2254, N1309);
and AND4 (N2546, N2543, N499, N1768, N373);
not NOT1 (N2547, N2538);
nor NOR3 (N2548, N2539, N1373, N1079);
xor XOR2 (N2549, N2542, N1051);
xor XOR2 (N2550, N2544, N1828);
and AND4 (N2551, N2545, N391, N325, N784);
nand NAND3 (N2552, N2547, N628, N525);
nand NAND4 (N2553, N2522, N61, N1016, N2138);
nand NAND2 (N2554, N2540, N1709);
nand NAND4 (N2555, N2549, N1945, N260, N1899);
buf BUF1 (N2556, N2551);
nor NOR2 (N2557, N2553, N638);
or OR4 (N2558, N2556, N2175, N1000, N104);
buf BUF1 (N2559, N2510);
or OR2 (N2560, N2554, N1761);
not NOT1 (N2561, N2550);
or OR4 (N2562, N2552, N1263, N2375, N2368);
xor XOR2 (N2563, N2562, N2166);
and AND4 (N2564, N2533, N565, N1042, N1001);
not NOT1 (N2565, N2563);
or OR2 (N2566, N2559, N86);
xor XOR2 (N2567, N2558, N1725);
nand NAND4 (N2568, N2561, N1290, N2184, N2177);
xor XOR2 (N2569, N2560, N1584);
and AND4 (N2570, N2548, N1105, N1008, N744);
nand NAND3 (N2571, N2569, N1067, N1738);
or OR3 (N2572, N2568, N912, N1587);
xor XOR2 (N2573, N2566, N1741);
and AND2 (N2574, N2573, N1379);
nand NAND2 (N2575, N2546, N666);
and AND4 (N2576, N2572, N1278, N1764, N1094);
not NOT1 (N2577, N2570);
nand NAND3 (N2578, N2577, N2010, N541);
nor NOR2 (N2579, N2567, N913);
nand NAND3 (N2580, N2565, N2491, N1844);
nand NAND2 (N2581, N2557, N262);
nand NAND2 (N2582, N2576, N585);
buf BUF1 (N2583, N2564);
buf BUF1 (N2584, N2583);
and AND4 (N2585, N2580, N2176, N2560, N1307);
nand NAND4 (N2586, N2575, N2509, N1860, N1063);
and AND3 (N2587, N2581, N1566, N364);
and AND2 (N2588, N2582, N1518);
buf BUF1 (N2589, N2579);
not NOT1 (N2590, N2588);
and AND4 (N2591, N2574, N2345, N501, N1358);
not NOT1 (N2592, N2555);
or OR2 (N2593, N2584, N723);
xor XOR2 (N2594, N2589, N1353);
xor XOR2 (N2595, N2585, N1652);
not NOT1 (N2596, N2571);
buf BUF1 (N2597, N2596);
nand NAND2 (N2598, N2594, N1446);
or OR2 (N2599, N2587, N1802);
or OR3 (N2600, N2595, N370, N359);
nor NOR2 (N2601, N2597, N993);
not NOT1 (N2602, N2598);
buf BUF1 (N2603, N2591);
nor NOR4 (N2604, N2603, N2287, N99, N2128);
not NOT1 (N2605, N2586);
buf BUF1 (N2606, N2592);
nor NOR3 (N2607, N2606, N738, N761);
not NOT1 (N2608, N2578);
nand NAND3 (N2609, N2599, N64, N788);
or OR4 (N2610, N2604, N2240, N2363, N2202);
or OR3 (N2611, N2593, N2234, N1036);
nand NAND4 (N2612, N2608, N1733, N1504, N2082);
buf BUF1 (N2613, N2607);
xor XOR2 (N2614, N2601, N1597);
nor NOR2 (N2615, N2609, N375);
nor NOR3 (N2616, N2605, N173, N1595);
not NOT1 (N2617, N2600);
buf BUF1 (N2618, N2617);
or OR4 (N2619, N2618, N426, N1741, N2524);
or OR4 (N2620, N2590, N2391, N533, N129);
nor NOR2 (N2621, N2616, N2599);
xor XOR2 (N2622, N2614, N1468);
nand NAND4 (N2623, N2612, N2615, N1498, N112);
and AND2 (N2624, N643, N2305);
or OR2 (N2625, N2619, N1141);
nor NOR3 (N2626, N2622, N417, N591);
nor NOR3 (N2627, N2621, N776, N2015);
or OR2 (N2628, N2625, N306);
buf BUF1 (N2629, N2620);
nand NAND2 (N2630, N2629, N1639);
buf BUF1 (N2631, N2610);
xor XOR2 (N2632, N2631, N1609);
nand NAND3 (N2633, N2626, N2067, N723);
nor NOR3 (N2634, N2613, N352, N2542);
and AND4 (N2635, N2628, N1301, N2157, N1550);
or OR3 (N2636, N2634, N397, N423);
buf BUF1 (N2637, N2635);
buf BUF1 (N2638, N2627);
xor XOR2 (N2639, N2611, N1746);
not NOT1 (N2640, N2632);
xor XOR2 (N2641, N2639, N784);
not NOT1 (N2642, N2630);
and AND3 (N2643, N2642, N1846, N2196);
and AND4 (N2644, N2624, N77, N440, N734);
xor XOR2 (N2645, N2640, N851);
buf BUF1 (N2646, N2638);
buf BUF1 (N2647, N2633);
or OR2 (N2648, N2602, N2392);
nor NOR2 (N2649, N2648, N265);
or OR2 (N2650, N2643, N940);
and AND3 (N2651, N2649, N2132, N588);
nor NOR2 (N2652, N2645, N2489);
and AND3 (N2653, N2637, N905, N1029);
nor NOR4 (N2654, N2647, N988, N219, N1042);
nand NAND2 (N2655, N2653, N1818);
nand NAND4 (N2656, N2651, N2224, N745, N1435);
xor XOR2 (N2657, N2623, N428);
or OR2 (N2658, N2644, N1494);
nand NAND4 (N2659, N2641, N509, N2105, N1404);
nand NAND2 (N2660, N2656, N431);
and AND4 (N2661, N2646, N1843, N1372, N33);
xor XOR2 (N2662, N2650, N2334);
nor NOR2 (N2663, N2654, N1897);
or OR2 (N2664, N2652, N879);
or OR4 (N2665, N2660, N303, N2076, N1050);
and AND3 (N2666, N2636, N1279, N843);
not NOT1 (N2667, N2661);
buf BUF1 (N2668, N2655);
buf BUF1 (N2669, N2657);
xor XOR2 (N2670, N2668, N1378);
and AND2 (N2671, N2664, N2408);
not NOT1 (N2672, N2670);
xor XOR2 (N2673, N2658, N2158);
nand NAND2 (N2674, N2662, N340);
and AND4 (N2675, N2667, N2084, N435, N607);
xor XOR2 (N2676, N2673, N2149);
xor XOR2 (N2677, N2674, N2547);
xor XOR2 (N2678, N2669, N208);
buf BUF1 (N2679, N2666);
and AND2 (N2680, N2671, N1747);
and AND4 (N2681, N2672, N410, N964, N1452);
buf BUF1 (N2682, N2665);
or OR4 (N2683, N2659, N2651, N378, N1467);
and AND3 (N2684, N2675, N390, N2324);
or OR2 (N2685, N2682, N1809);
nor NOR3 (N2686, N2678, N2394, N2547);
and AND2 (N2687, N2686, N2266);
and AND3 (N2688, N2677, N1062, N1780);
nor NOR4 (N2689, N2684, N208, N54, N1288);
xor XOR2 (N2690, N2679, N84);
xor XOR2 (N2691, N2663, N1480);
nand NAND2 (N2692, N2691, N1058);
or OR2 (N2693, N2680, N1956);
nor NOR3 (N2694, N2676, N2360, N2150);
nand NAND2 (N2695, N2687, N1816);
buf BUF1 (N2696, N2692);
nor NOR3 (N2697, N2683, N939, N393);
or OR3 (N2698, N2688, N1445, N295);
not NOT1 (N2699, N2694);
nor NOR3 (N2700, N2698, N2203, N2518);
nor NOR4 (N2701, N2693, N1617, N1645, N21);
nand NAND2 (N2702, N2700, N1479);
nor NOR4 (N2703, N2685, N1570, N1960, N342);
xor XOR2 (N2704, N2695, N799);
xor XOR2 (N2705, N2699, N1615);
nand NAND2 (N2706, N2697, N1772);
xor XOR2 (N2707, N2706, N1904);
or OR4 (N2708, N2681, N895, N2657, N75);
nor NOR2 (N2709, N2689, N1676);
nor NOR3 (N2710, N2704, N107, N2095);
not NOT1 (N2711, N2705);
not NOT1 (N2712, N2709);
not NOT1 (N2713, N2701);
nor NOR2 (N2714, N2711, N1650);
buf BUF1 (N2715, N2713);
xor XOR2 (N2716, N2710, N1509);
nand NAND3 (N2717, N2703, N2210, N1224);
nand NAND2 (N2718, N2707, N1119);
nor NOR2 (N2719, N2718, N1224);
and AND3 (N2720, N2708, N393, N1314);
and AND2 (N2721, N2715, N2644);
or OR3 (N2722, N2690, N2646, N685);
nand NAND2 (N2723, N2720, N1221);
not NOT1 (N2724, N2717);
nand NAND4 (N2725, N2702, N534, N2222, N1252);
or OR3 (N2726, N2712, N1257, N1113);
and AND4 (N2727, N2726, N356, N1483, N1560);
not NOT1 (N2728, N2724);
and AND3 (N2729, N2725, N2655, N1342);
xor XOR2 (N2730, N2696, N2448);
not NOT1 (N2731, N2730);
nand NAND2 (N2732, N2731, N424);
not NOT1 (N2733, N2722);
not NOT1 (N2734, N2733);
xor XOR2 (N2735, N2727, N2344);
not NOT1 (N2736, N2735);
not NOT1 (N2737, N2723);
or OR2 (N2738, N2734, N809);
not NOT1 (N2739, N2737);
xor XOR2 (N2740, N2732, N2201);
nor NOR2 (N2741, N2721, N1665);
nor NOR4 (N2742, N2740, N2237, N599, N218);
nand NAND4 (N2743, N2738, N2042, N2212, N292);
buf BUF1 (N2744, N2714);
xor XOR2 (N2745, N2744, N1384);
xor XOR2 (N2746, N2716, N397);
nor NOR2 (N2747, N2736, N2585);
xor XOR2 (N2748, N2746, N27);
buf BUF1 (N2749, N2742);
not NOT1 (N2750, N2719);
and AND3 (N2751, N2739, N601, N2409);
and AND3 (N2752, N2745, N610, N1576);
and AND4 (N2753, N2743, N824, N2109, N1577);
buf BUF1 (N2754, N2750);
or OR4 (N2755, N2752, N2177, N2148, N323);
xor XOR2 (N2756, N2747, N2019);
not NOT1 (N2757, N2754);
or OR4 (N2758, N2757, N633, N73, N332);
and AND4 (N2759, N2741, N1913, N1859, N1146);
and AND3 (N2760, N2728, N995, N1689);
and AND3 (N2761, N2760, N397, N2361);
or OR3 (N2762, N2755, N953, N662);
nand NAND2 (N2763, N2761, N1392);
nand NAND3 (N2764, N2758, N958, N2662);
buf BUF1 (N2765, N2748);
nand NAND4 (N2766, N2763, N1062, N435, N1743);
nand NAND3 (N2767, N2765, N1301, N676);
not NOT1 (N2768, N2767);
and AND3 (N2769, N2766, N1991, N1449);
not NOT1 (N2770, N2756);
nand NAND4 (N2771, N2762, N2000, N2484, N1435);
not NOT1 (N2772, N2749);
not NOT1 (N2773, N2753);
or OR4 (N2774, N2751, N864, N389, N463);
or OR2 (N2775, N2759, N599);
buf BUF1 (N2776, N2771);
or OR3 (N2777, N2769, N1142, N1786);
nand NAND2 (N2778, N2774, N1363);
and AND4 (N2779, N2768, N2598, N2424, N851);
and AND2 (N2780, N2764, N1114);
nand NAND2 (N2781, N2770, N559);
and AND3 (N2782, N2772, N2315, N1618);
and AND4 (N2783, N2776, N1306, N1560, N1515);
buf BUF1 (N2784, N2729);
nor NOR4 (N2785, N2783, N1539, N776, N1400);
buf BUF1 (N2786, N2773);
nor NOR2 (N2787, N2779, N82);
buf BUF1 (N2788, N2777);
or OR4 (N2789, N2775, N1571, N1605, N71);
nor NOR3 (N2790, N2789, N1802, N1751);
or OR3 (N2791, N2786, N567, N1304);
or OR4 (N2792, N2790, N209, N2702, N1815);
buf BUF1 (N2793, N2784);
or OR3 (N2794, N2788, N1507, N316);
nand NAND3 (N2795, N2785, N2554, N793);
and AND4 (N2796, N2781, N2559, N2092, N767);
xor XOR2 (N2797, N2795, N2744);
and AND3 (N2798, N2787, N1718, N1040);
nor NOR2 (N2799, N2794, N1503);
not NOT1 (N2800, N2797);
nor NOR4 (N2801, N2799, N633, N2449, N1782);
buf BUF1 (N2802, N2800);
or OR4 (N2803, N2796, N293, N1489, N1566);
buf BUF1 (N2804, N2792);
buf BUF1 (N2805, N2803);
and AND4 (N2806, N2798, N2293, N987, N1083);
nand NAND3 (N2807, N2793, N1449, N683);
not NOT1 (N2808, N2778);
or OR4 (N2809, N2782, N1419, N2345, N630);
nor NOR4 (N2810, N2808, N2275, N1975, N1869);
xor XOR2 (N2811, N2810, N2716);
xor XOR2 (N2812, N2805, N956);
xor XOR2 (N2813, N2807, N50);
or OR2 (N2814, N2813, N1936);
or OR2 (N2815, N2809, N363);
nor NOR3 (N2816, N2814, N1366, N1955);
not NOT1 (N2817, N2816);
not NOT1 (N2818, N2791);
not NOT1 (N2819, N2812);
buf BUF1 (N2820, N2804);
buf BUF1 (N2821, N2801);
or OR2 (N2822, N2819, N1945);
and AND3 (N2823, N2780, N76, N206);
or OR3 (N2824, N2811, N1985, N2245);
nand NAND3 (N2825, N2824, N2207, N1935);
buf BUF1 (N2826, N2821);
or OR2 (N2827, N2826, N1403);
not NOT1 (N2828, N2820);
nand NAND3 (N2829, N2815, N1439, N1562);
nand NAND2 (N2830, N2829, N2765);
nand NAND2 (N2831, N2825, N762);
nand NAND2 (N2832, N2830, N1745);
not NOT1 (N2833, N2832);
nand NAND3 (N2834, N2806, N2207, N2509);
nor NOR2 (N2835, N2822, N2457);
not NOT1 (N2836, N2818);
not NOT1 (N2837, N2817);
xor XOR2 (N2838, N2831, N654);
nor NOR3 (N2839, N2823, N1327, N2101);
not NOT1 (N2840, N2828);
nor NOR3 (N2841, N2840, N1546, N10);
buf BUF1 (N2842, N2838);
not NOT1 (N2843, N2841);
and AND3 (N2844, N2839, N1137, N1949);
or OR4 (N2845, N2835, N1499, N2048, N1450);
and AND4 (N2846, N2842, N1898, N484, N1871);
buf BUF1 (N2847, N2844);
or OR2 (N2848, N2834, N1343);
and AND2 (N2849, N2836, N910);
or OR3 (N2850, N2849, N2541, N2236);
nor NOR4 (N2851, N2833, N2142, N1356, N2614);
and AND2 (N2852, N2837, N1517);
xor XOR2 (N2853, N2848, N1141);
nand NAND4 (N2854, N2845, N2852, N2087, N280);
not NOT1 (N2855, N1233);
xor XOR2 (N2856, N2846, N369);
not NOT1 (N2857, N2854);
buf BUF1 (N2858, N2855);
or OR2 (N2859, N2847, N726);
nor NOR2 (N2860, N2802, N743);
not NOT1 (N2861, N2853);
or OR3 (N2862, N2858, N2021, N523);
and AND3 (N2863, N2859, N158, N1792);
nor NOR3 (N2864, N2860, N2527, N799);
buf BUF1 (N2865, N2843);
nor NOR2 (N2866, N2851, N808);
xor XOR2 (N2867, N2862, N2063);
nand NAND2 (N2868, N2827, N1707);
xor XOR2 (N2869, N2865, N1372);
or OR4 (N2870, N2861, N2397, N1373, N796);
nor NOR3 (N2871, N2867, N497, N667);
or OR4 (N2872, N2857, N2201, N2307, N2684);
buf BUF1 (N2873, N2871);
buf BUF1 (N2874, N2850);
not NOT1 (N2875, N2856);
or OR4 (N2876, N2863, N1077, N2103, N669);
buf BUF1 (N2877, N2874);
nor NOR2 (N2878, N2872, N806);
nand NAND3 (N2879, N2876, N868, N1741);
nor NOR3 (N2880, N2870, N1389, N872);
and AND4 (N2881, N2864, N2679, N1236, N738);
xor XOR2 (N2882, N2878, N1594);
not NOT1 (N2883, N2879);
not NOT1 (N2884, N2866);
not NOT1 (N2885, N2881);
buf BUF1 (N2886, N2868);
nand NAND2 (N2887, N2884, N2442);
or OR4 (N2888, N2885, N1547, N500, N417);
and AND2 (N2889, N2869, N884);
or OR3 (N2890, N2873, N199, N1103);
and AND3 (N2891, N2875, N908, N1517);
xor XOR2 (N2892, N2889, N418);
buf BUF1 (N2893, N2888);
nor NOR4 (N2894, N2887, N1398, N857, N2446);
buf BUF1 (N2895, N2882);
buf BUF1 (N2896, N2886);
and AND2 (N2897, N2891, N1112);
or OR4 (N2898, N2895, N1212, N24, N2482);
and AND4 (N2899, N2893, N1240, N2090, N1343);
or OR3 (N2900, N2894, N2129, N2238);
not NOT1 (N2901, N2892);
buf BUF1 (N2902, N2880);
and AND3 (N2903, N2900, N1072, N1654);
nor NOR4 (N2904, N2890, N2647, N334, N537);
and AND2 (N2905, N2903, N1837);
nor NOR4 (N2906, N2904, N1171, N622, N334);
and AND2 (N2907, N2883, N2847);
xor XOR2 (N2908, N2906, N1188);
nand NAND4 (N2909, N2901, N1504, N2700, N1207);
nand NAND3 (N2910, N2902, N1934, N2125);
or OR2 (N2911, N2909, N201);
not NOT1 (N2912, N2908);
xor XOR2 (N2913, N2905, N68);
and AND2 (N2914, N2907, N2851);
not NOT1 (N2915, N2899);
nor NOR2 (N2916, N2914, N2596);
nor NOR3 (N2917, N2915, N2466, N1934);
nor NOR3 (N2918, N2877, N2900, N2875);
not NOT1 (N2919, N2898);
and AND2 (N2920, N2910, N2282);
buf BUF1 (N2921, N2897);
and AND4 (N2922, N2920, N2385, N2076, N770);
nor NOR4 (N2923, N2919, N474, N1878, N2);
xor XOR2 (N2924, N2913, N1995);
and AND3 (N2925, N2918, N2320, N916);
buf BUF1 (N2926, N2917);
and AND4 (N2927, N2921, N2917, N767, N1758);
or OR3 (N2928, N2926, N413, N228);
not NOT1 (N2929, N2928);
and AND2 (N2930, N2916, N1594);
and AND3 (N2931, N2912, N2845, N350);
buf BUF1 (N2932, N2925);
buf BUF1 (N2933, N2931);
not NOT1 (N2934, N2911);
nand NAND4 (N2935, N2932, N1105, N1351, N2023);
and AND4 (N2936, N2922, N516, N2557, N2897);
nor NOR3 (N2937, N2929, N1548, N503);
and AND3 (N2938, N2937, N2294, N694);
nor NOR2 (N2939, N2927, N161);
buf BUF1 (N2940, N2938);
not NOT1 (N2941, N2933);
nor NOR2 (N2942, N2936, N1686);
nor NOR2 (N2943, N2923, N2121);
nand NAND3 (N2944, N2930, N230, N1151);
not NOT1 (N2945, N2934);
nand NAND3 (N2946, N2924, N400, N1146);
xor XOR2 (N2947, N2896, N2023);
xor XOR2 (N2948, N2942, N2058);
buf BUF1 (N2949, N2941);
and AND3 (N2950, N2935, N322, N229);
nand NAND3 (N2951, N2940, N1124, N2609);
buf BUF1 (N2952, N2944);
not NOT1 (N2953, N2951);
nor NOR4 (N2954, N2947, N1085, N776, N894);
nor NOR4 (N2955, N2945, N48, N2477, N1817);
xor XOR2 (N2956, N2953, N1953);
or OR3 (N2957, N2955, N2579, N1520);
xor XOR2 (N2958, N2952, N750);
nand NAND3 (N2959, N2943, N1088, N2207);
not NOT1 (N2960, N2958);
nand NAND2 (N2961, N2954, N1383);
buf BUF1 (N2962, N2959);
nor NOR3 (N2963, N2956, N2635, N2512);
buf BUF1 (N2964, N2963);
nand NAND2 (N2965, N2948, N608);
and AND3 (N2966, N2962, N671, N1125);
buf BUF1 (N2967, N2961);
xor XOR2 (N2968, N2939, N1874);
buf BUF1 (N2969, N2957);
not NOT1 (N2970, N2967);
not NOT1 (N2971, N2946);
or OR4 (N2972, N2965, N1116, N1687, N1830);
nand NAND3 (N2973, N2971, N829, N1987);
and AND2 (N2974, N2960, N2486);
or OR3 (N2975, N2972, N532, N260);
or OR2 (N2976, N2970, N2933);
or OR4 (N2977, N2949, N85, N1445, N1600);
and AND4 (N2978, N2975, N2758, N2679, N1837);
buf BUF1 (N2979, N2978);
nand NAND3 (N2980, N2964, N1303, N936);
not NOT1 (N2981, N2968);
nand NAND4 (N2982, N2969, N556, N661, N33);
and AND3 (N2983, N2950, N667, N970);
not NOT1 (N2984, N2982);
or OR3 (N2985, N2976, N1120, N2017);
nor NOR3 (N2986, N2974, N2189, N2234);
nand NAND4 (N2987, N2980, N2759, N1756, N23);
nor NOR3 (N2988, N2977, N2628, N1611);
buf BUF1 (N2989, N2973);
nand NAND3 (N2990, N2981, N1351, N414);
nand NAND3 (N2991, N2985, N431, N1570);
xor XOR2 (N2992, N2983, N2584);
buf BUF1 (N2993, N2966);
or OR4 (N2994, N2989, N1062, N1863, N134);
or OR2 (N2995, N2984, N1383);
or OR2 (N2996, N2979, N400);
nand NAND3 (N2997, N2993, N1978, N2375);
xor XOR2 (N2998, N2986, N2177);
and AND2 (N2999, N2990, N2046);
or OR4 (N3000, N2997, N1755, N1656, N2788);
not NOT1 (N3001, N2992);
nor NOR3 (N3002, N2994, N1863, N2976);
or OR3 (N3003, N2996, N2407, N492);
buf BUF1 (N3004, N3003);
and AND2 (N3005, N3001, N1872);
xor XOR2 (N3006, N2995, N688);
or OR2 (N3007, N3004, N2948);
not NOT1 (N3008, N3002);
or OR2 (N3009, N2998, N293);
or OR3 (N3010, N3007, N540, N1677);
buf BUF1 (N3011, N2999);
nor NOR3 (N3012, N3006, N1092, N465);
nor NOR4 (N3013, N3011, N1934, N2390, N2052);
nand NAND3 (N3014, N2991, N2719, N1648);
or OR2 (N3015, N3012, N1117);
xor XOR2 (N3016, N2987, N1357);
not NOT1 (N3017, N3014);
nand NAND2 (N3018, N2988, N988);
and AND3 (N3019, N3015, N2980, N988);
nand NAND3 (N3020, N3016, N2603, N2831);
buf BUF1 (N3021, N3008);
buf BUF1 (N3022, N3018);
xor XOR2 (N3023, N3005, N1910);
buf BUF1 (N3024, N3020);
nor NOR4 (N3025, N3023, N2449, N2884, N780);
xor XOR2 (N3026, N3022, N429);
or OR2 (N3027, N3025, N2829);
nor NOR4 (N3028, N3000, N978, N2889, N1252);
or OR3 (N3029, N3028, N2840, N1245);
or OR2 (N3030, N3027, N2785);
xor XOR2 (N3031, N3030, N2858);
xor XOR2 (N3032, N3029, N2497);
and AND3 (N3033, N3010, N2983, N2188);
xor XOR2 (N3034, N3017, N534);
not NOT1 (N3035, N3031);
nand NAND4 (N3036, N3021, N2730, N204, N104);
xor XOR2 (N3037, N3034, N1404);
and AND3 (N3038, N3037, N100, N855);
xor XOR2 (N3039, N3019, N1851);
buf BUF1 (N3040, N3033);
nor NOR3 (N3041, N3038, N2086, N701);
or OR2 (N3042, N3041, N773);
or OR2 (N3043, N3013, N1636);
nor NOR4 (N3044, N3009, N884, N1725, N1348);
xor XOR2 (N3045, N3044, N1544);
not NOT1 (N3046, N3036);
nand NAND4 (N3047, N3040, N933, N1481, N2937);
or OR3 (N3048, N3046, N1397, N1438);
or OR4 (N3049, N3047, N1801, N2183, N2804);
nor NOR3 (N3050, N3039, N903, N2559);
not NOT1 (N3051, N3026);
nand NAND2 (N3052, N3043, N2646);
and AND3 (N3053, N3049, N2214, N947);
not NOT1 (N3054, N3050);
buf BUF1 (N3055, N3051);
nor NOR4 (N3056, N3053, N346, N1192, N699);
buf BUF1 (N3057, N3042);
and AND2 (N3058, N3055, N1836);
buf BUF1 (N3059, N3024);
xor XOR2 (N3060, N3057, N2004);
and AND3 (N3061, N3035, N1395, N2824);
xor XOR2 (N3062, N3059, N2276);
xor XOR2 (N3063, N3061, N955);
buf BUF1 (N3064, N3056);
not NOT1 (N3065, N3063);
or OR2 (N3066, N3032, N1664);
nor NOR3 (N3067, N3060, N2590, N2099);
nand NAND2 (N3068, N3054, N1218);
nor NOR3 (N3069, N3065, N418, N111);
and AND4 (N3070, N3052, N1309, N1277, N1663);
xor XOR2 (N3071, N3066, N783);
nand NAND2 (N3072, N3069, N2446);
and AND4 (N3073, N3068, N2227, N408, N152);
buf BUF1 (N3074, N3072);
nand NAND3 (N3075, N3070, N1731, N1977);
not NOT1 (N3076, N3064);
nand NAND4 (N3077, N3076, N1177, N2894, N240);
xor XOR2 (N3078, N3071, N2330);
nand NAND3 (N3079, N3058, N999, N1947);
and AND3 (N3080, N3077, N1707, N2719);
not NOT1 (N3081, N3074);
or OR2 (N3082, N3048, N2159);
or OR3 (N3083, N3067, N1643, N785);
nand NAND4 (N3084, N3079, N2702, N2795, N2931);
nor NOR2 (N3085, N3075, N2020);
buf BUF1 (N3086, N3073);
nand NAND3 (N3087, N3082, N1660, N1655);
not NOT1 (N3088, N3085);
or OR2 (N3089, N3062, N2690);
nor NOR3 (N3090, N3084, N258, N2498);
and AND3 (N3091, N3086, N687, N20);
nand NAND4 (N3092, N3087, N2345, N524, N1755);
nand NAND4 (N3093, N3091, N2694, N2574, N1294);
and AND2 (N3094, N3093, N2311);
or OR3 (N3095, N3094, N2032, N1523);
nor NOR4 (N3096, N3095, N1964, N2148, N2434);
buf BUF1 (N3097, N3089);
xor XOR2 (N3098, N3045, N1656);
xor XOR2 (N3099, N3088, N2687);
xor XOR2 (N3100, N3097, N2167);
xor XOR2 (N3101, N3096, N747);
nor NOR4 (N3102, N3090, N400, N1672, N483);
xor XOR2 (N3103, N3101, N1543);
not NOT1 (N3104, N3098);
not NOT1 (N3105, N3100);
and AND3 (N3106, N3083, N2691, N604);
or OR3 (N3107, N3102, N1082, N829);
nand NAND2 (N3108, N3092, N855);
buf BUF1 (N3109, N3080);
or OR3 (N3110, N3099, N1706, N112);
nor NOR4 (N3111, N3108, N652, N3093, N2813);
or OR4 (N3112, N3109, N1298, N1374, N2345);
not NOT1 (N3113, N3112);
not NOT1 (N3114, N3113);
xor XOR2 (N3115, N3114, N392);
or OR4 (N3116, N3104, N2777, N2258, N947);
or OR2 (N3117, N3110, N2997);
buf BUF1 (N3118, N3105);
not NOT1 (N3119, N3117);
not NOT1 (N3120, N3081);
or OR2 (N3121, N3116, N2592);
nand NAND4 (N3122, N3106, N644, N2032, N2669);
nand NAND3 (N3123, N3115, N2883, N1620);
nor NOR2 (N3124, N3120, N1869);
nor NOR3 (N3125, N3107, N271, N2473);
buf BUF1 (N3126, N3124);
and AND3 (N3127, N3126, N2904, N1338);
and AND3 (N3128, N3119, N1452, N448);
xor XOR2 (N3129, N3118, N460);
or OR3 (N3130, N3125, N212, N1607);
buf BUF1 (N3131, N3128);
nor NOR3 (N3132, N3131, N1695, N2804);
nand NAND2 (N3133, N3078, N1118);
not NOT1 (N3134, N3130);
xor XOR2 (N3135, N3111, N2557);
or OR2 (N3136, N3103, N374);
nor NOR3 (N3137, N3132, N2180, N3131);
xor XOR2 (N3138, N3137, N2477);
xor XOR2 (N3139, N3133, N189);
not NOT1 (N3140, N3136);
and AND2 (N3141, N3122, N1046);
and AND2 (N3142, N3135, N696);
nand NAND3 (N3143, N3142, N1949, N936);
or OR3 (N3144, N3123, N2652, N1958);
buf BUF1 (N3145, N3139);
buf BUF1 (N3146, N3141);
nor NOR4 (N3147, N3121, N1241, N2394, N2874);
not NOT1 (N3148, N3147);
or OR3 (N3149, N3134, N2118, N392);
xor XOR2 (N3150, N3127, N1227);
not NOT1 (N3151, N3144);
nor NOR4 (N3152, N3151, N420, N1592, N1019);
nor NOR3 (N3153, N3143, N1034, N291);
xor XOR2 (N3154, N3146, N2376);
xor XOR2 (N3155, N3129, N3077);
xor XOR2 (N3156, N3140, N708);
nor NOR4 (N3157, N3145, N1016, N914, N822);
buf BUF1 (N3158, N3154);
or OR2 (N3159, N3158, N2739);
buf BUF1 (N3160, N3156);
or OR3 (N3161, N3159, N2707, N1266);
nor NOR4 (N3162, N3148, N1629, N238, N2898);
nand NAND2 (N3163, N3152, N1181);
or OR4 (N3164, N3161, N3081, N1329, N2908);
nand NAND4 (N3165, N3160, N711, N927, N225);
and AND2 (N3166, N3162, N2721);
not NOT1 (N3167, N3153);
nand NAND4 (N3168, N3149, N2380, N1576, N900);
buf BUF1 (N3169, N3164);
nor NOR3 (N3170, N3166, N2730, N1832);
buf BUF1 (N3171, N3163);
and AND2 (N3172, N3169, N1090);
xor XOR2 (N3173, N3165, N706);
buf BUF1 (N3174, N3170);
or OR4 (N3175, N3167, N278, N2441, N2202);
or OR2 (N3176, N3173, N746);
not NOT1 (N3177, N3171);
nor NOR2 (N3178, N3157, N2522);
nand NAND4 (N3179, N3178, N2507, N184, N1488);
xor XOR2 (N3180, N3150, N347);
or OR3 (N3181, N3168, N2413, N1583);
or OR2 (N3182, N3174, N714);
and AND2 (N3183, N3182, N2465);
or OR4 (N3184, N3177, N2331, N1248, N3065);
nand NAND4 (N3185, N3155, N2768, N2115, N1299);
nand NAND3 (N3186, N3176, N790, N1099);
or OR3 (N3187, N3184, N1161, N2725);
nand NAND2 (N3188, N3179, N2111);
buf BUF1 (N3189, N3172);
nor NOR2 (N3190, N3185, N2835);
nor NOR3 (N3191, N3190, N123, N2022);
not NOT1 (N3192, N3181);
and AND3 (N3193, N3192, N1816, N1912);
not NOT1 (N3194, N3138);
nor NOR3 (N3195, N3189, N2540, N1362);
xor XOR2 (N3196, N3194, N999);
nand NAND2 (N3197, N3196, N426);
xor XOR2 (N3198, N3191, N2335);
not NOT1 (N3199, N3197);
xor XOR2 (N3200, N3188, N2569);
not NOT1 (N3201, N3175);
xor XOR2 (N3202, N3195, N1596);
nand NAND4 (N3203, N3193, N2508, N879, N440);
buf BUF1 (N3204, N3186);
not NOT1 (N3205, N3187);
nor NOR3 (N3206, N3180, N3055, N610);
nand NAND4 (N3207, N3204, N1713, N2778, N754);
xor XOR2 (N3208, N3198, N1553);
nor NOR4 (N3209, N3201, N2586, N1356, N2151);
and AND2 (N3210, N3199, N2738);
nand NAND2 (N3211, N3200, N1683);
nand NAND2 (N3212, N3206, N453);
not NOT1 (N3213, N3183);
not NOT1 (N3214, N3209);
xor XOR2 (N3215, N3208, N2196);
not NOT1 (N3216, N3203);
nor NOR3 (N3217, N3211, N563, N502);
and AND3 (N3218, N3212, N136, N66);
nor NOR4 (N3219, N3207, N2130, N1260, N861);
or OR4 (N3220, N3214, N1013, N2789, N2360);
buf BUF1 (N3221, N3217);
and AND2 (N3222, N3210, N2643);
or OR4 (N3223, N3222, N3145, N3042, N2290);
not NOT1 (N3224, N3219);
xor XOR2 (N3225, N3216, N2644);
or OR2 (N3226, N3213, N1232);
or OR4 (N3227, N3226, N152, N3197, N2092);
and AND3 (N3228, N3224, N908, N787);
or OR3 (N3229, N3221, N226, N704);
nand NAND4 (N3230, N3225, N141, N3095, N35);
or OR3 (N3231, N3229, N1931, N2183);
buf BUF1 (N3232, N3230);
not NOT1 (N3233, N3228);
xor XOR2 (N3234, N3233, N1119);
not NOT1 (N3235, N3223);
nand NAND4 (N3236, N3215, N3105, N1501, N2989);
and AND3 (N3237, N3220, N760, N2826);
nand NAND2 (N3238, N3202, N1253);
nor NOR3 (N3239, N3227, N627, N1315);
buf BUF1 (N3240, N3218);
nor NOR2 (N3241, N3237, N1712);
nor NOR4 (N3242, N3205, N1220, N515, N220);
nand NAND4 (N3243, N3234, N306, N244, N90);
or OR3 (N3244, N3241, N663, N311);
and AND3 (N3245, N3242, N876, N2133);
not NOT1 (N3246, N3235);
nand NAND2 (N3247, N3231, N102);
nor NOR2 (N3248, N3245, N1004);
nand NAND4 (N3249, N3246, N505, N510, N423);
not NOT1 (N3250, N3236);
or OR2 (N3251, N3248, N2908);
not NOT1 (N3252, N3239);
or OR3 (N3253, N3249, N182, N1150);
xor XOR2 (N3254, N3247, N1233);
xor XOR2 (N3255, N3244, N885);
xor XOR2 (N3256, N3255, N2241);
nor NOR3 (N3257, N3254, N1628, N392);
and AND3 (N3258, N3257, N1214, N1126);
or OR4 (N3259, N3258, N2592, N1846, N1861);
xor XOR2 (N3260, N3251, N1362);
nor NOR4 (N3261, N3260, N3044, N2076, N1536);
or OR3 (N3262, N3256, N1632, N1131);
and AND4 (N3263, N3250, N1284, N2501, N2058);
nand NAND4 (N3264, N3262, N2889, N2055, N545);
nand NAND3 (N3265, N3261, N2228, N1132);
not NOT1 (N3266, N3259);
xor XOR2 (N3267, N3243, N1330);
buf BUF1 (N3268, N3238);
or OR4 (N3269, N3267, N2869, N2199, N2083);
buf BUF1 (N3270, N3266);
not NOT1 (N3271, N3270);
nand NAND2 (N3272, N3265, N2842);
and AND2 (N3273, N3268, N2266);
xor XOR2 (N3274, N3252, N908);
nand NAND2 (N3275, N3273, N567);
nor NOR2 (N3276, N3271, N950);
xor XOR2 (N3277, N3253, N550);
nor NOR4 (N3278, N3272, N2967, N2766, N2658);
and AND3 (N3279, N3274, N2970, N898);
and AND4 (N3280, N3264, N2903, N1535, N920);
nand NAND4 (N3281, N3240, N502, N17, N870);
nor NOR4 (N3282, N3280, N1397, N3079, N426);
not NOT1 (N3283, N3232);
xor XOR2 (N3284, N3283, N1671);
or OR3 (N3285, N3282, N1734, N1174);
not NOT1 (N3286, N3275);
and AND2 (N3287, N3263, N1944);
buf BUF1 (N3288, N3269);
not NOT1 (N3289, N3278);
nand NAND2 (N3290, N3287, N456);
nand NAND2 (N3291, N3279, N2852);
not NOT1 (N3292, N3286);
or OR4 (N3293, N3289, N3153, N642, N2692);
nor NOR3 (N3294, N3276, N205, N836);
xor XOR2 (N3295, N3293, N2523);
buf BUF1 (N3296, N3294);
xor XOR2 (N3297, N3290, N170);
xor XOR2 (N3298, N3285, N1539);
not NOT1 (N3299, N3298);
xor XOR2 (N3300, N3295, N3234);
not NOT1 (N3301, N3300);
not NOT1 (N3302, N3292);
buf BUF1 (N3303, N3296);
buf BUF1 (N3304, N3302);
or OR2 (N3305, N3288, N3185);
and AND4 (N3306, N3305, N2608, N833, N2120);
and AND3 (N3307, N3297, N2703, N2584);
nor NOR2 (N3308, N3291, N2853);
buf BUF1 (N3309, N3281);
and AND2 (N3310, N3284, N1460);
not NOT1 (N3311, N3307);
nor NOR2 (N3312, N3303, N2357);
not NOT1 (N3313, N3304);
or OR2 (N3314, N3306, N1015);
or OR3 (N3315, N3313, N896, N594);
or OR2 (N3316, N3310, N162);
nand NAND3 (N3317, N3311, N1255, N397);
nand NAND2 (N3318, N3315, N1633);
buf BUF1 (N3319, N3317);
and AND2 (N3320, N3277, N2064);
xor XOR2 (N3321, N3314, N2965);
nor NOR2 (N3322, N3308, N235);
buf BUF1 (N3323, N3321);
nor NOR3 (N3324, N3299, N717, N1871);
xor XOR2 (N3325, N3316, N2812);
xor XOR2 (N3326, N3322, N1678);
nand NAND3 (N3327, N3320, N2087, N151);
nand NAND3 (N3328, N3326, N2471, N2554);
xor XOR2 (N3329, N3319, N816);
nand NAND3 (N3330, N3328, N350, N1105);
xor XOR2 (N3331, N3323, N2610);
buf BUF1 (N3332, N3312);
nor NOR3 (N3333, N3324, N712, N2999);
nand NAND4 (N3334, N3332, N1758, N2242, N1608);
buf BUF1 (N3335, N3318);
and AND3 (N3336, N3335, N679, N1610);
nand NAND3 (N3337, N3309, N1012, N2006);
and AND3 (N3338, N3329, N685, N2183);
xor XOR2 (N3339, N3325, N3336);
or OR4 (N3340, N3319, N146, N553, N1779);
or OR3 (N3341, N3334, N241, N1938);
not NOT1 (N3342, N3341);
buf BUF1 (N3343, N3338);
nand NAND4 (N3344, N3343, N2722, N1397, N1833);
nand NAND4 (N3345, N3333, N1105, N2231, N858);
buf BUF1 (N3346, N3331);
nand NAND2 (N3347, N3340, N2940);
or OR2 (N3348, N3327, N45);
nand NAND4 (N3349, N3345, N54, N1800, N548);
nor NOR4 (N3350, N3337, N1564, N1029, N66);
not NOT1 (N3351, N3330);
not NOT1 (N3352, N3301);
nor NOR2 (N3353, N3339, N3115);
and AND2 (N3354, N3342, N3046);
nand NAND3 (N3355, N3349, N788, N806);
or OR4 (N3356, N3347, N2362, N1144, N1245);
not NOT1 (N3357, N3350);
or OR2 (N3358, N3355, N1021);
or OR2 (N3359, N3357, N1201);
buf BUF1 (N3360, N3359);
buf BUF1 (N3361, N3352);
and AND4 (N3362, N3346, N1996, N964, N1163);
xor XOR2 (N3363, N3358, N52);
buf BUF1 (N3364, N3353);
not NOT1 (N3365, N3344);
and AND3 (N3366, N3362, N1994, N3194);
and AND3 (N3367, N3356, N588, N541);
nor NOR4 (N3368, N3364, N2415, N1013, N947);
xor XOR2 (N3369, N3354, N3218);
buf BUF1 (N3370, N3351);
xor XOR2 (N3371, N3348, N1629);
or OR2 (N3372, N3363, N361);
nand NAND2 (N3373, N3372, N803);
or OR2 (N3374, N3370, N2154);
and AND3 (N3375, N3368, N1382, N2369);
and AND3 (N3376, N3367, N2118, N2983);
buf BUF1 (N3377, N3373);
buf BUF1 (N3378, N3366);
xor XOR2 (N3379, N3378, N2126);
nand NAND2 (N3380, N3379, N2074);
or OR2 (N3381, N3369, N670);
buf BUF1 (N3382, N3376);
nand NAND2 (N3383, N3371, N734);
xor XOR2 (N3384, N3374, N361);
buf BUF1 (N3385, N3377);
nand NAND2 (N3386, N3385, N2067);
or OR3 (N3387, N3365, N3016, N2940);
nor NOR2 (N3388, N3360, N2257);
nor NOR2 (N3389, N3387, N2047);
or OR4 (N3390, N3388, N1191, N2956, N141);
nand NAND4 (N3391, N3361, N2491, N3311, N1745);
xor XOR2 (N3392, N3390, N604);
buf BUF1 (N3393, N3375);
or OR2 (N3394, N3382, N716);
not NOT1 (N3395, N3393);
and AND3 (N3396, N3391, N1938, N38);
and AND2 (N3397, N3380, N1335);
or OR4 (N3398, N3384, N629, N2693, N2068);
nor NOR3 (N3399, N3386, N2106, N3151);
and AND3 (N3400, N3395, N1307, N2399);
buf BUF1 (N3401, N3398);
nand NAND2 (N3402, N3392, N2447);
nor NOR3 (N3403, N3389, N2115, N1982);
xor XOR2 (N3404, N3400, N3288);
xor XOR2 (N3405, N3394, N1347);
nand NAND2 (N3406, N3397, N30);
nor NOR3 (N3407, N3399, N2253, N3078);
and AND2 (N3408, N3401, N800);
or OR4 (N3409, N3403, N654, N1783, N812);
or OR2 (N3410, N3409, N2393);
nand NAND3 (N3411, N3407, N1134, N208);
buf BUF1 (N3412, N3411);
nor NOR3 (N3413, N3408, N2797, N1746);
or OR4 (N3414, N3381, N831, N516, N1728);
not NOT1 (N3415, N3383);
xor XOR2 (N3416, N3402, N2150);
nor NOR2 (N3417, N3412, N1901);
xor XOR2 (N3418, N3406, N171);
nand NAND4 (N3419, N3413, N2960, N966, N1278);
not NOT1 (N3420, N3396);
nand NAND4 (N3421, N3414, N3210, N1390, N2763);
and AND2 (N3422, N3405, N2743);
or OR4 (N3423, N3420, N551, N1850, N1297);
not NOT1 (N3424, N3416);
and AND4 (N3425, N3421, N3286, N3214, N69);
and AND3 (N3426, N3417, N3392, N2018);
and AND4 (N3427, N3415, N2998, N237, N843);
not NOT1 (N3428, N3422);
not NOT1 (N3429, N3404);
not NOT1 (N3430, N3428);
buf BUF1 (N3431, N3419);
nor NOR3 (N3432, N3430, N3326, N2696);
nor NOR4 (N3433, N3423, N366, N612, N852);
not NOT1 (N3434, N3427);
nand NAND2 (N3435, N3426, N1191);
nand NAND3 (N3436, N3434, N2103, N1348);
and AND2 (N3437, N3432, N379);
buf BUF1 (N3438, N3431);
xor XOR2 (N3439, N3429, N1763);
not NOT1 (N3440, N3433);
nor NOR4 (N3441, N3418, N3223, N2236, N345);
nand NAND3 (N3442, N3425, N1261, N943);
or OR4 (N3443, N3436, N2452, N1547, N463);
not NOT1 (N3444, N3410);
or OR4 (N3445, N3437, N1987, N2037, N3194);
xor XOR2 (N3446, N3445, N1806);
buf BUF1 (N3447, N3440);
and AND3 (N3448, N3424, N1010, N1216);
buf BUF1 (N3449, N3444);
and AND3 (N3450, N3435, N3019, N1797);
or OR3 (N3451, N3447, N3381, N45);
buf BUF1 (N3452, N3441);
buf BUF1 (N3453, N3449);
nor NOR4 (N3454, N3439, N727, N1303, N2801);
nand NAND3 (N3455, N3442, N3247, N2967);
nor NOR3 (N3456, N3455, N1817, N8);
or OR3 (N3457, N3456, N550, N2665);
and AND4 (N3458, N3454, N175, N2978, N3284);
buf BUF1 (N3459, N3453);
and AND3 (N3460, N3443, N787, N1959);
or OR2 (N3461, N3448, N2230);
and AND2 (N3462, N3458, N1653);
xor XOR2 (N3463, N3459, N357);
or OR2 (N3464, N3452, N2963);
nor NOR3 (N3465, N3438, N321, N2359);
nand NAND2 (N3466, N3446, N1811);
not NOT1 (N3467, N3466);
xor XOR2 (N3468, N3462, N3370);
and AND3 (N3469, N3451, N3212, N263);
and AND4 (N3470, N3467, N3211, N753, N2386);
nor NOR2 (N3471, N3457, N1035);
not NOT1 (N3472, N3465);
nor NOR2 (N3473, N3468, N1054);
xor XOR2 (N3474, N3461, N2898);
xor XOR2 (N3475, N3469, N3447);
or OR3 (N3476, N3450, N2860, N400);
nor NOR4 (N3477, N3476, N143, N891, N434);
not NOT1 (N3478, N3474);
nand NAND2 (N3479, N3472, N1573);
nor NOR3 (N3480, N3471, N3044, N1419);
and AND2 (N3481, N3460, N2109);
or OR3 (N3482, N3479, N2297, N3245);
buf BUF1 (N3483, N3480);
or OR4 (N3484, N3473, N316, N2339, N416);
not NOT1 (N3485, N3481);
xor XOR2 (N3486, N3484, N1738);
not NOT1 (N3487, N3470);
buf BUF1 (N3488, N3477);
buf BUF1 (N3489, N3488);
and AND2 (N3490, N3475, N565);
or OR2 (N3491, N3463, N2073);
or OR4 (N3492, N3489, N1290, N3253, N1163);
nand NAND2 (N3493, N3464, N2955);
xor XOR2 (N3494, N3486, N3310);
buf BUF1 (N3495, N3494);
nand NAND4 (N3496, N3478, N228, N596, N1110);
nor NOR3 (N3497, N3491, N1142, N1053);
buf BUF1 (N3498, N3495);
and AND3 (N3499, N3485, N2286, N2932);
not NOT1 (N3500, N3482);
nand NAND4 (N3501, N3497, N2804, N2517, N359);
not NOT1 (N3502, N3499);
xor XOR2 (N3503, N3492, N3126);
and AND4 (N3504, N3493, N946, N3319, N955);
xor XOR2 (N3505, N3498, N1757);
nor NOR4 (N3506, N3487, N1358, N254, N1396);
buf BUF1 (N3507, N3503);
nand NAND2 (N3508, N3506, N3161);
nor NOR4 (N3509, N3496, N3001, N2539, N857);
buf BUF1 (N3510, N3502);
and AND3 (N3511, N3504, N1577, N244);
and AND3 (N3512, N3510, N3075, N306);
and AND4 (N3513, N3505, N648, N851, N2820);
not NOT1 (N3514, N3508);
and AND2 (N3515, N3501, N3220);
not NOT1 (N3516, N3507);
nor NOR3 (N3517, N3513, N2496, N1657);
nand NAND2 (N3518, N3500, N2886);
buf BUF1 (N3519, N3517);
nor NOR2 (N3520, N3490, N1751);
nor NOR2 (N3521, N3512, N1320);
not NOT1 (N3522, N3509);
endmodule