// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21;

output N25620,N25619,N25615,N25616,N25607,N25614,N25613,N25617,N25618,N25621;

xor XOR2 (N22, N16, N14);
buf BUF1 (N23, N14);
and AND2 (N24, N7, N15);
nor NOR2 (N25, N21, N23);
buf BUF1 (N26, N13);
not NOT1 (N27, N25);
and AND3 (N28, N18, N1, N24);
and AND2 (N29, N2, N23);
or OR3 (N30, N24, N7, N19);
not NOT1 (N31, N2);
buf BUF1 (N32, N22);
buf BUF1 (N33, N24);
buf BUF1 (N34, N16);
nand NAND4 (N35, N24, N20, N23, N32);
buf BUF1 (N36, N18);
nor NOR2 (N37, N35, N17);
buf BUF1 (N38, N28);
xor XOR2 (N39, N34, N37);
buf BUF1 (N40, N1);
or OR3 (N41, N26, N20, N20);
or OR3 (N42, N29, N10, N17);
xor XOR2 (N43, N30, N12);
or OR4 (N44, N38, N6, N24, N12);
xor XOR2 (N45, N39, N3);
xor XOR2 (N46, N42, N19);
and AND2 (N47, N45, N9);
nand NAND2 (N48, N40, N46);
or OR2 (N49, N17, N29);
not NOT1 (N50, N47);
nand NAND3 (N51, N27, N16, N31);
nand NAND2 (N52, N2, N39);
nand NAND2 (N53, N51, N36);
and AND3 (N54, N18, N49, N17);
nand NAND2 (N55, N22, N43);
buf BUF1 (N56, N39);
xor XOR2 (N57, N55, N25);
buf BUF1 (N58, N41);
and AND2 (N59, N53, N40);
nand NAND3 (N60, N57, N2, N30);
nor NOR4 (N61, N50, N45, N53, N59);
nand NAND4 (N62, N57, N42, N17, N1);
nor NOR2 (N63, N62, N36);
and AND4 (N64, N63, N63, N21, N17);
and AND4 (N65, N48, N51, N64, N64);
or OR4 (N66, N36, N46, N64, N53);
nand NAND4 (N67, N54, N63, N17, N34);
nor NOR2 (N68, N44, N63);
nand NAND2 (N69, N68, N67);
and AND2 (N70, N63, N1);
not NOT1 (N71, N56);
buf BUF1 (N72, N70);
xor XOR2 (N73, N72, N27);
and AND2 (N74, N61, N11);
and AND2 (N75, N33, N18);
or OR2 (N76, N75, N3);
xor XOR2 (N77, N69, N47);
or OR2 (N78, N77, N43);
nand NAND2 (N79, N76, N32);
xor XOR2 (N80, N58, N35);
xor XOR2 (N81, N52, N35);
nand NAND4 (N82, N73, N39, N50, N2);
or OR4 (N83, N81, N4, N10, N57);
nand NAND4 (N84, N80, N49, N42, N23);
nand NAND2 (N85, N71, N28);
nor NOR3 (N86, N82, N12, N69);
not NOT1 (N87, N66);
not NOT1 (N88, N79);
and AND4 (N89, N85, N29, N23, N55);
and AND4 (N90, N86, N21, N3, N46);
or OR3 (N91, N88, N20, N11);
nand NAND3 (N92, N83, N22, N36);
buf BUF1 (N93, N78);
nand NAND3 (N94, N87, N41, N18);
xor XOR2 (N95, N92, N6);
xor XOR2 (N96, N89, N15);
buf BUF1 (N97, N96);
xor XOR2 (N98, N60, N83);
not NOT1 (N99, N90);
nand NAND2 (N100, N97, N6);
or OR4 (N101, N65, N87, N56, N65);
xor XOR2 (N102, N84, N8);
xor XOR2 (N103, N74, N91);
and AND3 (N104, N27, N23, N77);
xor XOR2 (N105, N98, N4);
not NOT1 (N106, N100);
buf BUF1 (N107, N104);
xor XOR2 (N108, N107, N46);
xor XOR2 (N109, N102, N67);
not NOT1 (N110, N103);
not NOT1 (N111, N105);
and AND2 (N112, N111, N17);
nor NOR3 (N113, N95, N20, N40);
nand NAND3 (N114, N113, N104, N39);
buf BUF1 (N115, N114);
xor XOR2 (N116, N99, N57);
xor XOR2 (N117, N112, N70);
and AND2 (N118, N93, N67);
nor NOR2 (N119, N110, N62);
buf BUF1 (N120, N117);
nor NOR2 (N121, N108, N16);
nand NAND3 (N122, N101, N113, N86);
xor XOR2 (N123, N115, N92);
not NOT1 (N124, N123);
xor XOR2 (N125, N121, N100);
nand NAND3 (N126, N124, N88, N116);
nor NOR2 (N127, N93, N90);
or OR4 (N128, N122, N4, N49, N51);
xor XOR2 (N129, N126, N66);
xor XOR2 (N130, N94, N113);
nor NOR3 (N131, N130, N103, N118);
and AND3 (N132, N48, N78, N25);
not NOT1 (N133, N119);
nor NOR2 (N134, N128, N84);
xor XOR2 (N135, N127, N49);
or OR3 (N136, N131, N35, N5);
nor NOR3 (N137, N129, N84, N67);
buf BUF1 (N138, N136);
nand NAND2 (N139, N138, N128);
xor XOR2 (N140, N132, N101);
nor NOR4 (N141, N137, N80, N89, N32);
or OR4 (N142, N109, N120, N95, N9);
nor NOR3 (N143, N63, N48, N117);
nor NOR3 (N144, N143, N46, N48);
xor XOR2 (N145, N142, N57);
or OR3 (N146, N106, N131, N95);
nand NAND4 (N147, N139, N23, N18, N56);
xor XOR2 (N148, N147, N89);
not NOT1 (N149, N148);
nand NAND2 (N150, N134, N102);
and AND2 (N151, N133, N134);
and AND4 (N152, N141, N50, N103, N94);
nand NAND4 (N153, N152, N70, N24, N40);
xor XOR2 (N154, N125, N27);
buf BUF1 (N155, N153);
xor XOR2 (N156, N150, N155);
and AND4 (N157, N145, N139, N150, N61);
not NOT1 (N158, N80);
xor XOR2 (N159, N135, N158);
not NOT1 (N160, N75);
nand NAND4 (N161, N160, N30, N65, N99);
not NOT1 (N162, N149);
nand NAND3 (N163, N157, N41, N69);
nor NOR4 (N164, N144, N132, N63, N125);
or OR3 (N165, N161, N48, N13);
nand NAND3 (N166, N164, N59, N125);
xor XOR2 (N167, N162, N46);
xor XOR2 (N168, N154, N73);
nand NAND2 (N169, N163, N67);
or OR3 (N170, N140, N79, N159);
and AND3 (N171, N8, N162, N11);
and AND2 (N172, N165, N137);
xor XOR2 (N173, N156, N70);
or OR3 (N174, N166, N114, N55);
nand NAND2 (N175, N171, N69);
buf BUF1 (N176, N170);
and AND2 (N177, N168, N118);
not NOT1 (N178, N169);
nor NOR3 (N179, N146, N130, N37);
not NOT1 (N180, N176);
xor XOR2 (N181, N173, N82);
and AND2 (N182, N180, N144);
or OR4 (N183, N174, N1, N140, N181);
and AND3 (N184, N13, N20, N39);
or OR4 (N185, N184, N163, N34, N163);
xor XOR2 (N186, N175, N172);
xor XOR2 (N187, N29, N53);
xor XOR2 (N188, N177, N77);
not NOT1 (N189, N179);
not NOT1 (N190, N186);
not NOT1 (N191, N187);
and AND4 (N192, N178, N138, N73, N123);
xor XOR2 (N193, N182, N52);
xor XOR2 (N194, N188, N24);
xor XOR2 (N195, N190, N108);
nor NOR3 (N196, N189, N122, N101);
buf BUF1 (N197, N193);
not NOT1 (N198, N183);
or OR3 (N199, N167, N81, N171);
and AND3 (N200, N151, N84, N130);
xor XOR2 (N201, N199, N32);
buf BUF1 (N202, N185);
xor XOR2 (N203, N200, N84);
nor NOR3 (N204, N196, N7, N148);
or OR3 (N205, N202, N11, N198);
buf BUF1 (N206, N168);
and AND4 (N207, N206, N53, N1, N36);
buf BUF1 (N208, N201);
and AND3 (N209, N207, N67, N140);
nand NAND3 (N210, N192, N144, N157);
nor NOR2 (N211, N210, N84);
not NOT1 (N212, N204);
nand NAND4 (N213, N203, N83, N136, N122);
and AND4 (N214, N213, N30, N172, N152);
and AND3 (N215, N195, N24, N24);
not NOT1 (N216, N208);
or OR4 (N217, N194, N138, N178, N210);
nand NAND3 (N218, N211, N119, N203);
nor NOR3 (N219, N205, N113, N217);
or OR4 (N220, N46, N28, N16, N101);
or OR3 (N221, N216, N150, N215);
not NOT1 (N222, N125);
xor XOR2 (N223, N214, N69);
nand NAND4 (N224, N220, N142, N198, N123);
nor NOR4 (N225, N209, N205, N140, N76);
nand NAND2 (N226, N223, N151);
or OR3 (N227, N224, N177, N165);
and AND4 (N228, N222, N217, N169, N48);
and AND4 (N229, N221, N96, N140, N78);
and AND3 (N230, N226, N100, N73);
or OR2 (N231, N212, N133);
nand NAND2 (N232, N219, N82);
nand NAND4 (N233, N225, N174, N172, N121);
buf BUF1 (N234, N232);
xor XOR2 (N235, N218, N117);
nor NOR3 (N236, N227, N120, N93);
nand NAND2 (N237, N231, N120);
not NOT1 (N238, N234);
xor XOR2 (N239, N230, N1);
not NOT1 (N240, N233);
and AND3 (N241, N240, N36, N234);
not NOT1 (N242, N238);
buf BUF1 (N243, N241);
or OR2 (N244, N236, N141);
not NOT1 (N245, N242);
buf BUF1 (N246, N228);
nor NOR4 (N247, N191, N242, N51, N73);
buf BUF1 (N248, N245);
xor XOR2 (N249, N247, N190);
nand NAND3 (N250, N229, N208, N167);
and AND4 (N251, N249, N57, N14, N172);
xor XOR2 (N252, N251, N195);
not NOT1 (N253, N248);
xor XOR2 (N254, N250, N81);
not NOT1 (N255, N246);
buf BUF1 (N256, N255);
nand NAND4 (N257, N197, N32, N218, N210);
or OR3 (N258, N239, N124, N230);
xor XOR2 (N259, N252, N173);
xor XOR2 (N260, N235, N192);
not NOT1 (N261, N257);
not NOT1 (N262, N260);
not NOT1 (N263, N258);
xor XOR2 (N264, N261, N38);
nor NOR3 (N265, N256, N173, N226);
xor XOR2 (N266, N253, N17);
and AND4 (N267, N263, N151, N20, N239);
nand NAND2 (N268, N267, N130);
buf BUF1 (N269, N266);
and AND2 (N270, N262, N260);
not NOT1 (N271, N264);
nor NOR3 (N272, N269, N31, N108);
and AND3 (N273, N244, N75, N219);
nor NOR2 (N274, N271, N26);
nand NAND4 (N275, N268, N215, N39, N216);
buf BUF1 (N276, N265);
nor NOR3 (N277, N272, N2, N204);
buf BUF1 (N278, N277);
xor XOR2 (N279, N254, N127);
not NOT1 (N280, N278);
or OR2 (N281, N276, N227);
xor XOR2 (N282, N280, N281);
buf BUF1 (N283, N245);
not NOT1 (N284, N273);
nor NOR2 (N285, N237, N189);
or OR3 (N286, N259, N223, N251);
not NOT1 (N287, N243);
not NOT1 (N288, N270);
or OR2 (N289, N288, N286);
buf BUF1 (N290, N214);
buf BUF1 (N291, N285);
buf BUF1 (N292, N289);
buf BUF1 (N293, N291);
and AND4 (N294, N293, N22, N60, N48);
or OR3 (N295, N274, N269, N138);
not NOT1 (N296, N283);
and AND2 (N297, N287, N287);
nand NAND4 (N298, N295, N175, N44, N217);
or OR4 (N299, N296, N294, N101, N213);
nand NAND2 (N300, N71, N122);
nand NAND4 (N301, N297, N56, N283, N207);
nand NAND2 (N302, N282, N163);
not NOT1 (N303, N284);
xor XOR2 (N304, N298, N149);
or OR4 (N305, N304, N37, N137, N238);
buf BUF1 (N306, N305);
buf BUF1 (N307, N302);
nand NAND3 (N308, N307, N164, N96);
and AND3 (N309, N299, N143, N96);
xor XOR2 (N310, N300, N185);
xor XOR2 (N311, N292, N107);
or OR2 (N312, N275, N14);
xor XOR2 (N313, N309, N155);
buf BUF1 (N314, N311);
xor XOR2 (N315, N314, N235);
xor XOR2 (N316, N308, N71);
nor NOR4 (N317, N303, N128, N270, N212);
and AND4 (N318, N310, N55, N246, N304);
xor XOR2 (N319, N313, N121);
nor NOR3 (N320, N279, N12, N237);
nand NAND4 (N321, N320, N35, N242, N278);
buf BUF1 (N322, N312);
nand NAND3 (N323, N290, N258, N201);
or OR2 (N324, N321, N71);
not NOT1 (N325, N315);
nor NOR2 (N326, N318, N104);
and AND2 (N327, N326, N251);
or OR2 (N328, N316, N326);
and AND3 (N329, N317, N81, N137);
not NOT1 (N330, N301);
nor NOR4 (N331, N322, N36, N263, N292);
and AND2 (N332, N327, N103);
or OR4 (N333, N324, N171, N206, N312);
not NOT1 (N334, N323);
not NOT1 (N335, N325);
buf BUF1 (N336, N306);
and AND3 (N337, N328, N51, N63);
or OR2 (N338, N333, N180);
and AND2 (N339, N330, N119);
buf BUF1 (N340, N337);
not NOT1 (N341, N334);
and AND2 (N342, N341, N340);
nand NAND2 (N343, N341, N192);
nor NOR4 (N344, N335, N110, N272, N215);
not NOT1 (N345, N342);
and AND2 (N346, N329, N90);
or OR2 (N347, N332, N68);
nor NOR2 (N348, N336, N134);
nor NOR2 (N349, N339, N273);
or OR4 (N350, N348, N137, N87, N187);
xor XOR2 (N351, N331, N314);
buf BUF1 (N352, N347);
nand NAND2 (N353, N343, N314);
xor XOR2 (N354, N346, N291);
xor XOR2 (N355, N344, N88);
and AND2 (N356, N350, N28);
and AND2 (N357, N354, N124);
not NOT1 (N358, N353);
xor XOR2 (N359, N338, N312);
nand NAND2 (N360, N351, N73);
and AND4 (N361, N359, N324, N110, N289);
or OR3 (N362, N355, N59, N344);
not NOT1 (N363, N349);
nand NAND3 (N364, N357, N189, N196);
not NOT1 (N365, N345);
buf BUF1 (N366, N363);
or OR2 (N367, N356, N146);
not NOT1 (N368, N362);
or OR2 (N369, N368, N233);
nor NOR2 (N370, N358, N322);
or OR3 (N371, N369, N308, N330);
not NOT1 (N372, N319);
or OR3 (N373, N372, N298, N245);
xor XOR2 (N374, N370, N306);
not NOT1 (N375, N373);
buf BUF1 (N376, N361);
buf BUF1 (N377, N375);
or OR4 (N378, N367, N304, N39, N183);
buf BUF1 (N379, N366);
and AND4 (N380, N360, N351, N320, N354);
nor NOR2 (N381, N365, N254);
xor XOR2 (N382, N352, N308);
and AND3 (N383, N380, N78, N225);
or OR3 (N384, N364, N250, N254);
nand NAND4 (N385, N374, N118, N158, N158);
nand NAND3 (N386, N385, N208, N297);
or OR3 (N387, N379, N31, N233);
xor XOR2 (N388, N378, N127);
and AND4 (N389, N383, N265, N221, N364);
nand NAND2 (N390, N388, N191);
nand NAND3 (N391, N390, N362, N294);
buf BUF1 (N392, N389);
buf BUF1 (N393, N376);
xor XOR2 (N394, N391, N139);
nand NAND2 (N395, N386, N341);
or OR3 (N396, N377, N137, N249);
xor XOR2 (N397, N384, N183);
or OR3 (N398, N393, N68, N374);
not NOT1 (N399, N387);
or OR3 (N400, N392, N105, N7);
not NOT1 (N401, N395);
buf BUF1 (N402, N398);
buf BUF1 (N403, N396);
not NOT1 (N404, N403);
not NOT1 (N405, N401);
and AND2 (N406, N400, N56);
not NOT1 (N407, N406);
or OR4 (N408, N399, N172, N243, N223);
xor XOR2 (N409, N402, N334);
and AND4 (N410, N405, N25, N289, N227);
and AND4 (N411, N371, N259, N245, N320);
and AND4 (N412, N408, N243, N361, N192);
not NOT1 (N413, N410);
nand NAND3 (N414, N394, N204, N55);
buf BUF1 (N415, N411);
xor XOR2 (N416, N397, N182);
and AND4 (N417, N413, N8, N300, N120);
and AND4 (N418, N407, N31, N285, N250);
buf BUF1 (N419, N382);
and AND4 (N420, N416, N75, N202, N238);
nand NAND4 (N421, N409, N288, N276, N367);
nand NAND2 (N422, N412, N345);
xor XOR2 (N423, N414, N156);
nand NAND3 (N424, N417, N20, N131);
or OR3 (N425, N423, N224, N155);
buf BUF1 (N426, N404);
not NOT1 (N427, N426);
nor NOR2 (N428, N424, N394);
not NOT1 (N429, N420);
or OR2 (N430, N381, N160);
xor XOR2 (N431, N419, N212);
and AND4 (N432, N428, N168, N12, N259);
and AND4 (N433, N422, N117, N116, N244);
nand NAND3 (N434, N425, N110, N328);
xor XOR2 (N435, N431, N259);
nand NAND4 (N436, N421, N26, N198, N80);
not NOT1 (N437, N430);
buf BUF1 (N438, N433);
or OR2 (N439, N432, N371);
nor NOR2 (N440, N418, N309);
xor XOR2 (N441, N438, N24);
nand NAND4 (N442, N440, N247, N143, N211);
nand NAND4 (N443, N437, N364, N293, N111);
or OR3 (N444, N442, N235, N106);
not NOT1 (N445, N429);
or OR3 (N446, N444, N255, N21);
xor XOR2 (N447, N439, N100);
and AND3 (N448, N443, N393, N315);
xor XOR2 (N449, N441, N164);
buf BUF1 (N450, N445);
nand NAND4 (N451, N450, N114, N85, N173);
and AND2 (N452, N427, N367);
nor NOR4 (N453, N446, N174, N386, N346);
and AND3 (N454, N449, N434, N348);
xor XOR2 (N455, N310, N42);
not NOT1 (N456, N435);
not NOT1 (N457, N448);
nor NOR3 (N458, N453, N112, N237);
not NOT1 (N459, N452);
buf BUF1 (N460, N436);
and AND4 (N461, N459, N439, N353, N371);
nor NOR4 (N462, N457, N371, N446, N182);
and AND3 (N463, N415, N233, N260);
not NOT1 (N464, N455);
nor NOR4 (N465, N447, N56, N335, N209);
nor NOR4 (N466, N456, N233, N421, N95);
not NOT1 (N467, N466);
buf BUF1 (N468, N458);
nand NAND2 (N469, N468, N240);
or OR3 (N470, N467, N351, N243);
buf BUF1 (N471, N464);
buf BUF1 (N472, N460);
nand NAND4 (N473, N472, N255, N42, N298);
or OR2 (N474, N454, N57);
and AND2 (N475, N462, N302);
or OR3 (N476, N465, N3, N338);
xor XOR2 (N477, N469, N349);
nand NAND3 (N478, N451, N196, N432);
not NOT1 (N479, N471);
and AND2 (N480, N463, N230);
buf BUF1 (N481, N480);
nor NOR4 (N482, N474, N345, N197, N380);
not NOT1 (N483, N481);
nand NAND2 (N484, N482, N327);
xor XOR2 (N485, N461, N98);
xor XOR2 (N486, N476, N420);
nand NAND3 (N487, N479, N229, N277);
buf BUF1 (N488, N477);
xor XOR2 (N489, N478, N371);
nand NAND2 (N490, N486, N331);
nor NOR2 (N491, N488, N401);
nand NAND4 (N492, N485, N38, N333, N311);
not NOT1 (N493, N489);
xor XOR2 (N494, N483, N63);
not NOT1 (N495, N492);
or OR3 (N496, N494, N400, N405);
and AND4 (N497, N491, N297, N434, N115);
or OR4 (N498, N484, N19, N463, N204);
buf BUF1 (N499, N496);
nor NOR3 (N500, N487, N170, N31);
nor NOR4 (N501, N490, N450, N12, N84);
nor NOR2 (N502, N475, N275);
nand NAND4 (N503, N502, N17, N386, N122);
and AND2 (N504, N499, N29);
nand NAND2 (N505, N497, N28);
or OR2 (N506, N503, N99);
nor NOR4 (N507, N495, N227, N227, N355);
or OR3 (N508, N470, N185, N260);
nand NAND4 (N509, N493, N494, N507, N215);
xor XOR2 (N510, N111, N402);
buf BUF1 (N511, N473);
buf BUF1 (N512, N500);
and AND3 (N513, N511, N134, N288);
and AND3 (N514, N512, N238, N204);
buf BUF1 (N515, N514);
nand NAND4 (N516, N508, N244, N195, N393);
or OR2 (N517, N515, N394);
or OR3 (N518, N498, N179, N500);
or OR3 (N519, N506, N276, N90);
not NOT1 (N520, N516);
or OR4 (N521, N518, N98, N63, N226);
not NOT1 (N522, N509);
and AND2 (N523, N517, N274);
nand NAND4 (N524, N522, N281, N140, N195);
buf BUF1 (N525, N524);
or OR2 (N526, N513, N168);
nand NAND3 (N527, N520, N13, N85);
and AND4 (N528, N505, N292, N215, N116);
nand NAND4 (N529, N510, N314, N46, N390);
or OR3 (N530, N528, N250, N412);
xor XOR2 (N531, N526, N379);
and AND4 (N532, N523, N465, N340, N123);
buf BUF1 (N533, N501);
or OR3 (N534, N521, N116, N74);
or OR3 (N535, N534, N178, N5);
nor NOR2 (N536, N519, N139);
and AND2 (N537, N531, N220);
or OR4 (N538, N537, N532, N472, N40);
buf BUF1 (N539, N178);
and AND2 (N540, N504, N36);
and AND2 (N541, N525, N505);
or OR4 (N542, N539, N88, N141, N476);
nor NOR4 (N543, N540, N267, N487, N343);
or OR4 (N544, N536, N376, N256, N324);
nand NAND4 (N545, N533, N233, N417, N41);
buf BUF1 (N546, N538);
and AND4 (N547, N544, N243, N537, N526);
xor XOR2 (N548, N527, N494);
and AND4 (N549, N541, N145, N299, N245);
or OR2 (N550, N542, N235);
nand NAND3 (N551, N529, N539, N316);
or OR4 (N552, N530, N328, N455, N157);
nor NOR4 (N553, N548, N220, N520, N166);
buf BUF1 (N554, N535);
buf BUF1 (N555, N547);
nand NAND4 (N556, N549, N132, N389, N331);
or OR3 (N557, N546, N379, N422);
xor XOR2 (N558, N551, N418);
buf BUF1 (N559, N553);
buf BUF1 (N560, N545);
xor XOR2 (N561, N559, N448);
and AND2 (N562, N558, N225);
nand NAND2 (N563, N557, N551);
or OR2 (N564, N561, N292);
nor NOR4 (N565, N555, N318, N13, N532);
not NOT1 (N566, N543);
not NOT1 (N567, N560);
xor XOR2 (N568, N556, N54);
or OR2 (N569, N552, N212);
xor XOR2 (N570, N563, N554);
and AND4 (N571, N372, N184, N378, N17);
xor XOR2 (N572, N562, N23);
and AND2 (N573, N568, N70);
nand NAND3 (N574, N567, N221, N548);
or OR4 (N575, N550, N433, N115, N449);
buf BUF1 (N576, N571);
and AND4 (N577, N564, N354, N135, N408);
buf BUF1 (N578, N577);
buf BUF1 (N579, N575);
nor NOR3 (N580, N576, N87, N321);
and AND2 (N581, N580, N354);
nand NAND3 (N582, N578, N64, N194);
and AND3 (N583, N566, N336, N499);
or OR2 (N584, N569, N72);
and AND4 (N585, N584, N265, N339, N133);
and AND2 (N586, N573, N147);
xor XOR2 (N587, N586, N316);
or OR3 (N588, N570, N48, N586);
xor XOR2 (N589, N587, N170);
xor XOR2 (N590, N565, N206);
or OR3 (N591, N588, N251, N570);
nand NAND2 (N592, N590, N120);
not NOT1 (N593, N582);
nand NAND2 (N594, N593, N84);
nand NAND3 (N595, N574, N507, N209);
nand NAND3 (N596, N595, N316, N194);
not NOT1 (N597, N579);
nand NAND2 (N598, N585, N424);
and AND4 (N599, N591, N228, N135, N340);
xor XOR2 (N600, N599, N367);
nand NAND2 (N601, N594, N67);
nand NAND2 (N602, N598, N466);
xor XOR2 (N603, N589, N137);
buf BUF1 (N604, N596);
xor XOR2 (N605, N603, N346);
not NOT1 (N606, N572);
not NOT1 (N607, N581);
buf BUF1 (N608, N605);
or OR3 (N609, N601, N599, N271);
or OR4 (N610, N602, N598, N362, N402);
buf BUF1 (N611, N597);
xor XOR2 (N612, N610, N241);
buf BUF1 (N613, N604);
or OR3 (N614, N583, N447, N389);
nor NOR4 (N615, N592, N176, N192, N282);
xor XOR2 (N616, N612, N197);
nor NOR4 (N617, N614, N509, N84, N601);
buf BUF1 (N618, N615);
and AND2 (N619, N609, N512);
xor XOR2 (N620, N619, N384);
nor NOR4 (N621, N606, N590, N129, N47);
xor XOR2 (N622, N611, N516);
or OR2 (N623, N621, N381);
and AND2 (N624, N613, N272);
xor XOR2 (N625, N616, N358);
nor NOR2 (N626, N622, N177);
not NOT1 (N627, N626);
and AND2 (N628, N617, N22);
nor NOR2 (N629, N627, N232);
nor NOR2 (N630, N618, N467);
not NOT1 (N631, N607);
or OR3 (N632, N624, N625, N617);
not NOT1 (N633, N413);
nand NAND3 (N634, N631, N146, N94);
xor XOR2 (N635, N630, N172);
xor XOR2 (N636, N620, N356);
not NOT1 (N637, N629);
and AND4 (N638, N636, N549, N608, N503);
and AND2 (N639, N201, N56);
xor XOR2 (N640, N634, N457);
and AND4 (N641, N632, N558, N239, N515);
buf BUF1 (N642, N638);
or OR4 (N643, N639, N73, N289, N74);
buf BUF1 (N644, N643);
nor NOR4 (N645, N600, N240, N260, N318);
buf BUF1 (N646, N645);
buf BUF1 (N647, N642);
buf BUF1 (N648, N635);
xor XOR2 (N649, N646, N127);
buf BUF1 (N650, N640);
not NOT1 (N651, N633);
nand NAND4 (N652, N650, N470, N565, N50);
not NOT1 (N653, N649);
or OR2 (N654, N652, N220);
buf BUF1 (N655, N647);
and AND2 (N656, N655, N67);
nand NAND3 (N657, N641, N359, N48);
and AND4 (N658, N648, N617, N612, N161);
nand NAND3 (N659, N656, N421, N241);
nor NOR2 (N660, N653, N2);
xor XOR2 (N661, N659, N334);
not NOT1 (N662, N628);
nor NOR3 (N663, N657, N418, N517);
or OR3 (N664, N637, N616, N216);
and AND4 (N665, N654, N261, N587, N39);
nand NAND2 (N666, N623, N554);
buf BUF1 (N667, N651);
nand NAND2 (N668, N667, N500);
or OR3 (N669, N666, N303, N336);
not NOT1 (N670, N663);
not NOT1 (N671, N665);
nand NAND4 (N672, N669, N50, N317, N367);
xor XOR2 (N673, N660, N332);
nand NAND2 (N674, N673, N281);
and AND3 (N675, N658, N296, N473);
not NOT1 (N676, N661);
or OR3 (N677, N664, N640, N8);
not NOT1 (N678, N644);
buf BUF1 (N679, N674);
buf BUF1 (N680, N670);
not NOT1 (N681, N668);
and AND2 (N682, N679, N651);
not NOT1 (N683, N682);
or OR4 (N684, N675, N502, N349, N143);
not NOT1 (N685, N676);
nand NAND2 (N686, N681, N396);
not NOT1 (N687, N683);
not NOT1 (N688, N672);
nor NOR3 (N689, N684, N333, N25);
not NOT1 (N690, N687);
or OR2 (N691, N680, N119);
nand NAND2 (N692, N688, N365);
or OR3 (N693, N692, N377, N346);
or OR4 (N694, N689, N523, N528, N292);
xor XOR2 (N695, N677, N684);
not NOT1 (N696, N678);
or OR3 (N697, N694, N212, N360);
or OR2 (N698, N691, N338);
nor NOR3 (N699, N671, N677, N405);
not NOT1 (N700, N686);
or OR2 (N701, N698, N13);
not NOT1 (N702, N695);
buf BUF1 (N703, N662);
nand NAND2 (N704, N685, N314);
and AND4 (N705, N697, N532, N249, N546);
and AND4 (N706, N703, N223, N490, N696);
nand NAND2 (N707, N157, N210);
not NOT1 (N708, N705);
or OR3 (N709, N707, N377, N580);
and AND4 (N710, N702, N352, N81, N662);
or OR2 (N711, N701, N51);
or OR2 (N712, N711, N205);
or OR2 (N713, N710, N581);
not NOT1 (N714, N713);
buf BUF1 (N715, N690);
or OR3 (N716, N714, N583, N604);
not NOT1 (N717, N708);
or OR2 (N718, N700, N697);
buf BUF1 (N719, N709);
nand NAND3 (N720, N704, N5, N661);
not NOT1 (N721, N706);
buf BUF1 (N722, N716);
not NOT1 (N723, N721);
or OR3 (N724, N718, N178, N497);
buf BUF1 (N725, N712);
or OR2 (N726, N723, N206);
nor NOR4 (N727, N717, N350, N697, N434);
not NOT1 (N728, N724);
buf BUF1 (N729, N725);
or OR4 (N730, N726, N546, N126, N406);
buf BUF1 (N731, N727);
xor XOR2 (N732, N728, N618);
or OR3 (N733, N729, N415, N574);
or OR3 (N734, N715, N173, N577);
buf BUF1 (N735, N720);
buf BUF1 (N736, N731);
or OR2 (N737, N734, N111);
nor NOR4 (N738, N737, N152, N492, N551);
buf BUF1 (N739, N693);
xor XOR2 (N740, N730, N30);
xor XOR2 (N741, N740, N256);
not NOT1 (N742, N699);
buf BUF1 (N743, N732);
and AND3 (N744, N736, N589, N136);
nand NAND2 (N745, N735, N558);
nor NOR4 (N746, N741, N74, N513, N739);
buf BUF1 (N747, N505);
nand NAND3 (N748, N742, N479, N520);
not NOT1 (N749, N748);
nand NAND3 (N750, N719, N468, N325);
not NOT1 (N751, N749);
and AND2 (N752, N746, N488);
or OR3 (N753, N750, N537, N267);
nor NOR3 (N754, N753, N592, N27);
and AND4 (N755, N754, N275, N497, N428);
nand NAND4 (N756, N738, N117, N83, N727);
nor NOR2 (N757, N722, N506);
not NOT1 (N758, N752);
xor XOR2 (N759, N747, N108);
not NOT1 (N760, N751);
xor XOR2 (N761, N745, N398);
buf BUF1 (N762, N744);
xor XOR2 (N763, N762, N745);
and AND4 (N764, N757, N614, N496, N310);
xor XOR2 (N765, N743, N719);
and AND2 (N766, N733, N221);
buf BUF1 (N767, N758);
and AND4 (N768, N759, N132, N270, N618);
not NOT1 (N769, N755);
nand NAND3 (N770, N764, N423, N276);
not NOT1 (N771, N756);
buf BUF1 (N772, N769);
and AND2 (N773, N772, N588);
buf BUF1 (N774, N773);
not NOT1 (N775, N766);
nand NAND2 (N776, N771, N643);
not NOT1 (N777, N767);
buf BUF1 (N778, N777);
not NOT1 (N779, N774);
buf BUF1 (N780, N779);
and AND4 (N781, N778, N99, N307, N111);
nor NOR4 (N782, N760, N587, N730, N28);
and AND2 (N783, N765, N654);
not NOT1 (N784, N776);
not NOT1 (N785, N781);
xor XOR2 (N786, N784, N163);
nand NAND2 (N787, N768, N7);
nand NAND2 (N788, N780, N150);
not NOT1 (N789, N763);
and AND2 (N790, N789, N12);
xor XOR2 (N791, N782, N280);
or OR4 (N792, N787, N638, N224, N785);
xor XOR2 (N793, N75, N413);
nor NOR3 (N794, N791, N467, N401);
nand NAND4 (N795, N786, N777, N419, N279);
xor XOR2 (N796, N792, N229);
xor XOR2 (N797, N761, N622);
nand NAND4 (N798, N790, N361, N75, N221);
xor XOR2 (N799, N788, N786);
not NOT1 (N800, N770);
xor XOR2 (N801, N796, N597);
xor XOR2 (N802, N775, N630);
not NOT1 (N803, N802);
not NOT1 (N804, N799);
buf BUF1 (N805, N783);
buf BUF1 (N806, N797);
buf BUF1 (N807, N798);
or OR2 (N808, N801, N764);
and AND4 (N809, N803, N806, N774, N314);
buf BUF1 (N810, N89);
xor XOR2 (N811, N810, N590);
nor NOR4 (N812, N807, N218, N803, N551);
not NOT1 (N813, N808);
nor NOR2 (N814, N813, N677);
buf BUF1 (N815, N800);
not NOT1 (N816, N814);
nand NAND2 (N817, N804, N253);
xor XOR2 (N818, N817, N4);
not NOT1 (N819, N795);
and AND3 (N820, N793, N727, N552);
nand NAND2 (N821, N815, N638);
nand NAND3 (N822, N811, N498, N583);
or OR3 (N823, N818, N788, N481);
or OR2 (N824, N823, N804);
nand NAND4 (N825, N824, N629, N53, N200);
nor NOR4 (N826, N820, N489, N764, N427);
buf BUF1 (N827, N794);
not NOT1 (N828, N826);
or OR2 (N829, N828, N737);
not NOT1 (N830, N827);
and AND4 (N831, N822, N28, N521, N74);
not NOT1 (N832, N812);
nor NOR3 (N833, N825, N295, N524);
or OR4 (N834, N832, N370, N236, N825);
xor XOR2 (N835, N834, N500);
nor NOR4 (N836, N821, N739, N133, N586);
and AND4 (N837, N809, N232, N508, N545);
nand NAND3 (N838, N837, N267, N796);
nand NAND2 (N839, N819, N644);
and AND4 (N840, N805, N289, N670, N203);
buf BUF1 (N841, N830);
xor XOR2 (N842, N838, N431);
xor XOR2 (N843, N842, N802);
or OR3 (N844, N843, N548, N773);
xor XOR2 (N845, N833, N258);
or OR2 (N846, N841, N354);
nand NAND3 (N847, N831, N457, N836);
buf BUF1 (N848, N614);
xor XOR2 (N849, N846, N492);
or OR2 (N850, N847, N37);
and AND3 (N851, N848, N603, N358);
buf BUF1 (N852, N835);
and AND3 (N853, N839, N107, N113);
or OR3 (N854, N844, N71, N228);
or OR2 (N855, N854, N454);
xor XOR2 (N856, N855, N312);
and AND3 (N857, N829, N348, N753);
not NOT1 (N858, N852);
xor XOR2 (N859, N851, N550);
and AND4 (N860, N856, N435, N55, N683);
xor XOR2 (N861, N859, N788);
buf BUF1 (N862, N860);
xor XOR2 (N863, N858, N117);
xor XOR2 (N864, N853, N640);
nor NOR3 (N865, N849, N814, N656);
xor XOR2 (N866, N864, N814);
not NOT1 (N867, N865);
nor NOR3 (N868, N862, N823, N113);
not NOT1 (N869, N863);
nand NAND4 (N870, N840, N824, N106, N739);
and AND3 (N871, N868, N376, N319);
not NOT1 (N872, N850);
nand NAND3 (N873, N857, N598, N285);
xor XOR2 (N874, N869, N855);
and AND4 (N875, N874, N700, N479, N304);
not NOT1 (N876, N866);
or OR3 (N877, N867, N316, N429);
nand NAND3 (N878, N870, N535, N704);
buf BUF1 (N879, N878);
and AND3 (N880, N845, N355, N414);
nor NOR2 (N881, N880, N332);
xor XOR2 (N882, N877, N481);
and AND4 (N883, N879, N10, N626, N578);
nand NAND2 (N884, N881, N392);
nor NOR2 (N885, N884, N414);
nand NAND3 (N886, N883, N763, N136);
or OR2 (N887, N871, N101);
buf BUF1 (N888, N885);
not NOT1 (N889, N816);
and AND3 (N890, N875, N586, N355);
nand NAND4 (N891, N890, N337, N361, N289);
or OR2 (N892, N886, N186);
and AND2 (N893, N889, N247);
xor XOR2 (N894, N872, N734);
not NOT1 (N895, N892);
and AND2 (N896, N876, N530);
not NOT1 (N897, N873);
not NOT1 (N898, N896);
and AND3 (N899, N894, N893, N143);
and AND3 (N900, N591, N503, N844);
nand NAND3 (N901, N887, N774, N61);
or OR4 (N902, N901, N40, N766, N351);
nor NOR3 (N903, N891, N658, N83);
nor NOR3 (N904, N882, N333, N678);
xor XOR2 (N905, N900, N467);
not NOT1 (N906, N888);
buf BUF1 (N907, N895);
or OR4 (N908, N905, N154, N56, N600);
or OR4 (N909, N898, N455, N592, N592);
xor XOR2 (N910, N909, N218);
xor XOR2 (N911, N903, N447);
xor XOR2 (N912, N904, N759);
or OR4 (N913, N911, N407, N874, N274);
xor XOR2 (N914, N912, N689);
and AND2 (N915, N913, N435);
nand NAND3 (N916, N902, N128, N741);
buf BUF1 (N917, N897);
nor NOR2 (N918, N915, N624);
nor NOR2 (N919, N861, N50);
not NOT1 (N920, N917);
buf BUF1 (N921, N910);
buf BUF1 (N922, N920);
buf BUF1 (N923, N914);
nand NAND4 (N924, N907, N27, N790, N788);
nor NOR2 (N925, N899, N240);
and AND2 (N926, N919, N373);
or OR2 (N927, N918, N390);
xor XOR2 (N928, N916, N592);
or OR2 (N929, N926, N841);
nor NOR3 (N930, N924, N767, N365);
buf BUF1 (N931, N930);
xor XOR2 (N932, N929, N417);
xor XOR2 (N933, N923, N314);
nand NAND3 (N934, N922, N462, N752);
nor NOR4 (N935, N928, N124, N257, N736);
xor XOR2 (N936, N927, N897);
nor NOR4 (N937, N925, N191, N436, N667);
or OR3 (N938, N934, N424, N404);
xor XOR2 (N939, N938, N272);
not NOT1 (N940, N932);
nand NAND3 (N941, N940, N849, N392);
not NOT1 (N942, N921);
buf BUF1 (N943, N931);
xor XOR2 (N944, N936, N250);
buf BUF1 (N945, N935);
not NOT1 (N946, N941);
or OR2 (N947, N937, N770);
nor NOR3 (N948, N933, N743, N857);
and AND4 (N949, N946, N698, N767, N232);
xor XOR2 (N950, N939, N576);
or OR2 (N951, N947, N53);
buf BUF1 (N952, N945);
nor NOR4 (N953, N944, N795, N61, N606);
nand NAND3 (N954, N948, N852, N949);
or OR3 (N955, N904, N806, N581);
nand NAND3 (N956, N943, N246, N183);
not NOT1 (N957, N908);
xor XOR2 (N958, N957, N30);
xor XOR2 (N959, N906, N461);
nor NOR3 (N960, N959, N38, N208);
nor NOR4 (N961, N950, N333, N555, N222);
nor NOR4 (N962, N942, N300, N682, N264);
xor XOR2 (N963, N954, N54);
nand NAND2 (N964, N962, N837);
nand NAND4 (N965, N952, N463, N113, N705);
and AND2 (N966, N965, N154);
not NOT1 (N967, N961);
nand NAND4 (N968, N956, N296, N842, N860);
or OR3 (N969, N953, N843, N555);
xor XOR2 (N970, N963, N31);
xor XOR2 (N971, N967, N858);
buf BUF1 (N972, N960);
buf BUF1 (N973, N951);
and AND4 (N974, N971, N432, N737, N75);
and AND4 (N975, N973, N110, N283, N819);
nor NOR3 (N976, N955, N91, N619);
buf BUF1 (N977, N974);
nor NOR2 (N978, N975, N533);
not NOT1 (N979, N968);
nand NAND4 (N980, N979, N448, N849, N847);
xor XOR2 (N981, N977, N160);
xor XOR2 (N982, N980, N544);
buf BUF1 (N983, N969);
buf BUF1 (N984, N983);
and AND4 (N985, N982, N329, N185, N749);
not NOT1 (N986, N966);
xor XOR2 (N987, N986, N919);
or OR4 (N988, N976, N369, N688, N453);
not NOT1 (N989, N964);
nand NAND3 (N990, N978, N344, N63);
xor XOR2 (N991, N985, N790);
and AND2 (N992, N984, N594);
nand NAND4 (N993, N970, N100, N709, N786);
nand NAND3 (N994, N972, N108, N720);
and AND4 (N995, N994, N395, N626, N585);
nor NOR4 (N996, N992, N444, N494, N926);
or OR4 (N997, N989, N751, N386, N654);
nand NAND4 (N998, N997, N455, N946, N925);
not NOT1 (N999, N988);
xor XOR2 (N1000, N987, N32);
nor NOR4 (N1001, N999, N1000, N965, N5);
nand NAND4 (N1002, N148, N301, N255, N595);
not NOT1 (N1003, N958);
nand NAND3 (N1004, N990, N540, N8);
buf BUF1 (N1005, N1004);
and AND4 (N1006, N1005, N713, N425, N334);
xor XOR2 (N1007, N995, N934);
buf BUF1 (N1008, N1002);
nand NAND3 (N1009, N1008, N1, N930);
buf BUF1 (N1010, N1001);
buf BUF1 (N1011, N1007);
xor XOR2 (N1012, N1006, N460);
nor NOR2 (N1013, N1009, N9);
nand NAND3 (N1014, N981, N579, N385);
or OR2 (N1015, N1003, N700);
nand NAND2 (N1016, N1015, N307);
not NOT1 (N1017, N996);
and AND4 (N1018, N1017, N908, N711, N722);
not NOT1 (N1019, N1018);
buf BUF1 (N1020, N1011);
nand NAND3 (N1021, N1012, N567, N485);
nand NAND4 (N1022, N1010, N585, N984, N678);
nand NAND4 (N1023, N1021, N159, N363, N783);
not NOT1 (N1024, N998);
not NOT1 (N1025, N1023);
not NOT1 (N1026, N1016);
xor XOR2 (N1027, N991, N133);
nand NAND2 (N1028, N1027, N964);
nor NOR2 (N1029, N1024, N502);
and AND2 (N1030, N1019, N94);
or OR2 (N1031, N1025, N975);
buf BUF1 (N1032, N1028);
nand NAND4 (N1033, N1029, N413, N220, N514);
or OR2 (N1034, N993, N645);
nand NAND2 (N1035, N1026, N751);
or OR2 (N1036, N1020, N748);
not NOT1 (N1037, N1032);
and AND3 (N1038, N1033, N980, N146);
xor XOR2 (N1039, N1037, N578);
or OR4 (N1040, N1031, N131, N917, N98);
not NOT1 (N1041, N1014);
not NOT1 (N1042, N1013);
not NOT1 (N1043, N1036);
not NOT1 (N1044, N1034);
nand NAND4 (N1045, N1043, N461, N900, N586);
and AND4 (N1046, N1044, N102, N564, N164);
nand NAND2 (N1047, N1042, N47);
nand NAND3 (N1048, N1039, N606, N183);
xor XOR2 (N1049, N1022, N984);
nand NAND4 (N1050, N1045, N781, N278, N1036);
buf BUF1 (N1051, N1048);
or OR4 (N1052, N1051, N202, N876, N954);
xor XOR2 (N1053, N1052, N989);
buf BUF1 (N1054, N1035);
and AND4 (N1055, N1053, N336, N909, N751);
or OR3 (N1056, N1040, N634, N630);
not NOT1 (N1057, N1041);
not NOT1 (N1058, N1056);
xor XOR2 (N1059, N1049, N797);
nor NOR3 (N1060, N1057, N111, N991);
nand NAND2 (N1061, N1050, N781);
nor NOR4 (N1062, N1058, N552, N471, N451);
or OR4 (N1063, N1062, N908, N856, N661);
and AND2 (N1064, N1046, N779);
xor XOR2 (N1065, N1063, N637);
xor XOR2 (N1066, N1030, N682);
or OR2 (N1067, N1064, N893);
nand NAND2 (N1068, N1055, N161);
buf BUF1 (N1069, N1060);
or OR2 (N1070, N1038, N764);
nor NOR3 (N1071, N1068, N456, N255);
and AND2 (N1072, N1047, N956);
nor NOR3 (N1073, N1054, N276, N698);
or OR4 (N1074, N1069, N285, N956, N321);
nor NOR2 (N1075, N1073, N461);
or OR2 (N1076, N1065, N394);
buf BUF1 (N1077, N1076);
buf BUF1 (N1078, N1066);
nand NAND2 (N1079, N1059, N954);
nor NOR3 (N1080, N1078, N1049, N236);
or OR2 (N1081, N1061, N107);
not NOT1 (N1082, N1081);
nand NAND4 (N1083, N1067, N197, N528, N767);
nor NOR3 (N1084, N1079, N810, N48);
and AND3 (N1085, N1072, N799, N294);
nor NOR2 (N1086, N1071, N501);
not NOT1 (N1087, N1082);
nor NOR4 (N1088, N1086, N617, N844, N488);
nor NOR4 (N1089, N1088, N944, N909, N305);
nand NAND4 (N1090, N1070, N942, N129, N576);
and AND2 (N1091, N1077, N356);
buf BUF1 (N1092, N1087);
nor NOR3 (N1093, N1083, N889, N764);
buf BUF1 (N1094, N1089);
not NOT1 (N1095, N1084);
or OR2 (N1096, N1075, N743);
and AND4 (N1097, N1090, N347, N311, N779);
and AND2 (N1098, N1096, N87);
and AND4 (N1099, N1094, N328, N924, N374);
or OR3 (N1100, N1085, N1057, N525);
not NOT1 (N1101, N1074);
or OR2 (N1102, N1080, N7);
and AND2 (N1103, N1092, N270);
and AND3 (N1104, N1091, N3, N864);
or OR4 (N1105, N1099, N415, N285, N689);
not NOT1 (N1106, N1095);
buf BUF1 (N1107, N1100);
or OR2 (N1108, N1101, N91);
buf BUF1 (N1109, N1098);
or OR2 (N1110, N1097, N629);
or OR2 (N1111, N1108, N246);
xor XOR2 (N1112, N1107, N264);
and AND3 (N1113, N1111, N787, N492);
buf BUF1 (N1114, N1109);
nor NOR4 (N1115, N1106, N533, N454, N540);
nor NOR2 (N1116, N1102, N612);
nor NOR2 (N1117, N1103, N936);
not NOT1 (N1118, N1114);
and AND4 (N1119, N1115, N117, N957, N997);
nor NOR2 (N1120, N1112, N994);
nand NAND3 (N1121, N1118, N15, N906);
and AND4 (N1122, N1104, N905, N641, N1079);
xor XOR2 (N1123, N1093, N832);
or OR2 (N1124, N1116, N287);
and AND4 (N1125, N1105, N816, N286, N1063);
nand NAND2 (N1126, N1110, N611);
nor NOR2 (N1127, N1124, N483);
nand NAND3 (N1128, N1122, N1076, N115);
nor NOR3 (N1129, N1121, N226, N478);
not NOT1 (N1130, N1117);
buf BUF1 (N1131, N1128);
or OR4 (N1132, N1123, N868, N516, N253);
and AND3 (N1133, N1119, N96, N167);
and AND3 (N1134, N1131, N879, N992);
and AND4 (N1135, N1113, N831, N916, N596);
buf BUF1 (N1136, N1129);
and AND3 (N1137, N1134, N565, N614);
buf BUF1 (N1138, N1135);
or OR2 (N1139, N1132, N118);
nor NOR4 (N1140, N1133, N93, N957, N793);
not NOT1 (N1141, N1127);
buf BUF1 (N1142, N1141);
buf BUF1 (N1143, N1126);
and AND4 (N1144, N1137, N61, N637, N762);
nand NAND4 (N1145, N1143, N568, N929, N359);
nor NOR3 (N1146, N1142, N156, N853);
buf BUF1 (N1147, N1130);
xor XOR2 (N1148, N1140, N1079);
xor XOR2 (N1149, N1138, N744);
not NOT1 (N1150, N1147);
and AND2 (N1151, N1120, N215);
and AND3 (N1152, N1139, N521, N365);
nor NOR2 (N1153, N1146, N652);
and AND2 (N1154, N1144, N167);
nand NAND2 (N1155, N1136, N996);
not NOT1 (N1156, N1152);
buf BUF1 (N1157, N1151);
xor XOR2 (N1158, N1145, N440);
and AND2 (N1159, N1157, N1154);
buf BUF1 (N1160, N467);
buf BUF1 (N1161, N1148);
buf BUF1 (N1162, N1149);
nor NOR4 (N1163, N1161, N1142, N499, N373);
xor XOR2 (N1164, N1159, N818);
or OR2 (N1165, N1158, N584);
not NOT1 (N1166, N1163);
xor XOR2 (N1167, N1150, N72);
and AND4 (N1168, N1166, N340, N156, N1005);
nor NOR2 (N1169, N1155, N1132);
buf BUF1 (N1170, N1164);
or OR3 (N1171, N1165, N162, N104);
or OR3 (N1172, N1153, N552, N379);
xor XOR2 (N1173, N1171, N266);
nand NAND3 (N1174, N1172, N121, N460);
and AND2 (N1175, N1168, N507);
not NOT1 (N1176, N1175);
or OR2 (N1177, N1174, N867);
or OR2 (N1178, N1177, N1100);
nor NOR2 (N1179, N1169, N201);
xor XOR2 (N1180, N1170, N481);
buf BUF1 (N1181, N1173);
nor NOR2 (N1182, N1162, N841);
nand NAND3 (N1183, N1160, N1172, N1011);
xor XOR2 (N1184, N1182, N702);
nand NAND2 (N1185, N1167, N824);
nand NAND3 (N1186, N1179, N884, N598);
not NOT1 (N1187, N1184);
and AND3 (N1188, N1187, N660, N722);
nor NOR4 (N1189, N1185, N30, N395, N830);
not NOT1 (N1190, N1125);
nand NAND2 (N1191, N1188, N563);
or OR2 (N1192, N1189, N958);
not NOT1 (N1193, N1180);
or OR2 (N1194, N1192, N375);
nor NOR4 (N1195, N1178, N1168, N177, N3);
and AND4 (N1196, N1193, N1141, N410, N910);
xor XOR2 (N1197, N1191, N943);
not NOT1 (N1198, N1195);
and AND4 (N1199, N1197, N967, N472, N1155);
and AND2 (N1200, N1198, N604);
xor XOR2 (N1201, N1199, N945);
or OR2 (N1202, N1194, N322);
nand NAND2 (N1203, N1186, N1143);
nor NOR4 (N1204, N1203, N625, N713, N1076);
and AND2 (N1205, N1201, N91);
and AND4 (N1206, N1156, N966, N740, N566);
or OR4 (N1207, N1181, N363, N121, N800);
and AND2 (N1208, N1200, N274);
nor NOR4 (N1209, N1208, N1149, N864, N592);
buf BUF1 (N1210, N1196);
nand NAND2 (N1211, N1210, N886);
not NOT1 (N1212, N1183);
xor XOR2 (N1213, N1202, N252);
nor NOR3 (N1214, N1206, N28, N981);
buf BUF1 (N1215, N1176);
not NOT1 (N1216, N1215);
buf BUF1 (N1217, N1216);
and AND4 (N1218, N1213, N572, N117, N828);
nand NAND2 (N1219, N1212, N1);
not NOT1 (N1220, N1205);
and AND3 (N1221, N1190, N49, N324);
buf BUF1 (N1222, N1204);
and AND3 (N1223, N1222, N1174, N187);
not NOT1 (N1224, N1218);
xor XOR2 (N1225, N1214, N324);
xor XOR2 (N1226, N1223, N2);
nand NAND2 (N1227, N1226, N899);
nand NAND2 (N1228, N1225, N231);
not NOT1 (N1229, N1227);
not NOT1 (N1230, N1220);
or OR3 (N1231, N1228, N886, N878);
nor NOR3 (N1232, N1221, N913, N720);
or OR2 (N1233, N1219, N200);
buf BUF1 (N1234, N1231);
buf BUF1 (N1235, N1233);
nor NOR3 (N1236, N1209, N32, N119);
nand NAND2 (N1237, N1207, N93);
buf BUF1 (N1238, N1235);
nand NAND4 (N1239, N1230, N463, N168, N964);
nor NOR2 (N1240, N1211, N104);
or OR4 (N1241, N1240, N505, N1040, N861);
or OR4 (N1242, N1234, N609, N946, N108);
nand NAND4 (N1243, N1232, N1220, N675, N1073);
nor NOR4 (N1244, N1242, N102, N1063, N532);
or OR2 (N1245, N1229, N1208);
and AND2 (N1246, N1243, N880);
nor NOR2 (N1247, N1246, N247);
nor NOR4 (N1248, N1244, N1230, N1145, N1015);
nand NAND2 (N1249, N1245, N456);
buf BUF1 (N1250, N1241);
or OR2 (N1251, N1248, N847);
nand NAND2 (N1252, N1217, N412);
or OR2 (N1253, N1249, N1203);
or OR4 (N1254, N1247, N750, N893, N647);
nand NAND3 (N1255, N1238, N124, N416);
buf BUF1 (N1256, N1224);
not NOT1 (N1257, N1256);
xor XOR2 (N1258, N1237, N859);
or OR3 (N1259, N1236, N348, N688);
buf BUF1 (N1260, N1251);
not NOT1 (N1261, N1239);
nand NAND4 (N1262, N1260, N517, N1224, N525);
nand NAND3 (N1263, N1258, N858, N525);
or OR4 (N1264, N1257, N79, N813, N38);
buf BUF1 (N1265, N1259);
not NOT1 (N1266, N1255);
not NOT1 (N1267, N1252);
xor XOR2 (N1268, N1254, N683);
not NOT1 (N1269, N1261);
and AND3 (N1270, N1263, N785, N1015);
or OR3 (N1271, N1268, N886, N1117);
or OR3 (N1272, N1266, N1259, N115);
or OR4 (N1273, N1267, N339, N89, N549);
or OR2 (N1274, N1269, N950);
xor XOR2 (N1275, N1274, N1174);
and AND3 (N1276, N1273, N275, N989);
buf BUF1 (N1277, N1253);
and AND3 (N1278, N1275, N152, N244);
nor NOR2 (N1279, N1262, N109);
buf BUF1 (N1280, N1277);
nand NAND2 (N1281, N1276, N675);
xor XOR2 (N1282, N1280, N503);
and AND4 (N1283, N1272, N70, N1187, N301);
nand NAND3 (N1284, N1271, N1218, N1280);
or OR2 (N1285, N1281, N703);
or OR4 (N1286, N1284, N1167, N841, N725);
nand NAND2 (N1287, N1282, N809);
buf BUF1 (N1288, N1250);
not NOT1 (N1289, N1285);
nor NOR4 (N1290, N1278, N1026, N1194, N335);
or OR4 (N1291, N1287, N1083, N58, N314);
or OR2 (N1292, N1291, N583);
xor XOR2 (N1293, N1288, N337);
not NOT1 (N1294, N1270);
nand NAND4 (N1295, N1264, N41, N576, N208);
nand NAND4 (N1296, N1283, N1067, N399, N446);
nand NAND2 (N1297, N1293, N465);
and AND4 (N1298, N1286, N116, N644, N1200);
not NOT1 (N1299, N1265);
xor XOR2 (N1300, N1279, N1150);
nand NAND4 (N1301, N1292, N908, N199, N487);
nand NAND2 (N1302, N1300, N758);
nand NAND4 (N1303, N1295, N210, N374, N994);
buf BUF1 (N1304, N1299);
buf BUF1 (N1305, N1303);
and AND4 (N1306, N1304, N464, N840, N835);
nand NAND3 (N1307, N1289, N1169, N247);
and AND2 (N1308, N1301, N284);
buf BUF1 (N1309, N1306);
nor NOR2 (N1310, N1307, N728);
nor NOR3 (N1311, N1296, N909, N276);
and AND4 (N1312, N1302, N878, N1190, N894);
nand NAND4 (N1313, N1309, N225, N166, N551);
and AND2 (N1314, N1305, N445);
nor NOR3 (N1315, N1313, N1050, N26);
buf BUF1 (N1316, N1290);
nor NOR3 (N1317, N1314, N152, N353);
not NOT1 (N1318, N1297);
nand NAND3 (N1319, N1312, N6, N888);
not NOT1 (N1320, N1315);
and AND3 (N1321, N1311, N69, N178);
xor XOR2 (N1322, N1310, N378);
nand NAND3 (N1323, N1298, N952, N806);
not NOT1 (N1324, N1308);
not NOT1 (N1325, N1317);
buf BUF1 (N1326, N1321);
buf BUF1 (N1327, N1320);
nor NOR2 (N1328, N1325, N466);
nor NOR2 (N1329, N1324, N308);
nor NOR4 (N1330, N1323, N306, N749, N1029);
or OR4 (N1331, N1318, N1205, N218, N238);
xor XOR2 (N1332, N1319, N752);
not NOT1 (N1333, N1328);
buf BUF1 (N1334, N1322);
and AND4 (N1335, N1294, N192, N578, N421);
or OR2 (N1336, N1332, N1248);
not NOT1 (N1337, N1327);
or OR4 (N1338, N1335, N1122, N1168, N1094);
buf BUF1 (N1339, N1337);
and AND4 (N1340, N1330, N161, N898, N451);
buf BUF1 (N1341, N1334);
or OR3 (N1342, N1338, N383, N862);
nand NAND2 (N1343, N1329, N436);
nor NOR2 (N1344, N1342, N583);
or OR4 (N1345, N1333, N662, N1268, N765);
or OR2 (N1346, N1340, N171);
nand NAND3 (N1347, N1344, N347, N877);
nand NAND2 (N1348, N1341, N696);
or OR4 (N1349, N1331, N409, N317, N885);
xor XOR2 (N1350, N1316, N460);
buf BUF1 (N1351, N1336);
xor XOR2 (N1352, N1348, N628);
nand NAND4 (N1353, N1350, N404, N626, N1264);
nor NOR3 (N1354, N1346, N1124, N1045);
and AND3 (N1355, N1353, N446, N55);
xor XOR2 (N1356, N1339, N926);
buf BUF1 (N1357, N1343);
and AND2 (N1358, N1326, N612);
nand NAND2 (N1359, N1352, N758);
nand NAND4 (N1360, N1351, N957, N496, N1231);
nand NAND4 (N1361, N1356, N262, N661, N998);
nand NAND3 (N1362, N1354, N927, N381);
not NOT1 (N1363, N1358);
or OR4 (N1364, N1355, N1047, N293, N88);
nor NOR3 (N1365, N1345, N992, N715);
nand NAND4 (N1366, N1359, N1195, N143, N613);
or OR2 (N1367, N1347, N720);
and AND3 (N1368, N1365, N676, N414);
or OR3 (N1369, N1360, N1354, N512);
or OR4 (N1370, N1366, N477, N1117, N887);
buf BUF1 (N1371, N1361);
xor XOR2 (N1372, N1362, N800);
xor XOR2 (N1373, N1369, N710);
nand NAND3 (N1374, N1363, N1202, N908);
nor NOR2 (N1375, N1371, N26);
nor NOR4 (N1376, N1367, N775, N1008, N104);
nor NOR4 (N1377, N1374, N1282, N614, N801);
nand NAND3 (N1378, N1364, N78, N187);
or OR4 (N1379, N1370, N193, N814, N428);
and AND3 (N1380, N1375, N817, N136);
and AND2 (N1381, N1377, N787);
nor NOR4 (N1382, N1380, N500, N15, N866);
buf BUF1 (N1383, N1378);
or OR3 (N1384, N1379, N423, N1077);
buf BUF1 (N1385, N1384);
buf BUF1 (N1386, N1357);
and AND3 (N1387, N1373, N587, N472);
not NOT1 (N1388, N1381);
or OR3 (N1389, N1382, N744, N78);
or OR3 (N1390, N1385, N683, N588);
not NOT1 (N1391, N1368);
buf BUF1 (N1392, N1372);
nor NOR2 (N1393, N1388, N354);
buf BUF1 (N1394, N1376);
or OR4 (N1395, N1386, N868, N622, N269);
nand NAND2 (N1396, N1392, N791);
or OR4 (N1397, N1391, N166, N598, N975);
or OR3 (N1398, N1394, N1143, N548);
or OR3 (N1399, N1393, N1006, N1001);
xor XOR2 (N1400, N1349, N357);
xor XOR2 (N1401, N1383, N872);
nor NOR3 (N1402, N1390, N1071, N612);
nor NOR3 (N1403, N1396, N631, N1204);
nor NOR3 (N1404, N1395, N901, N768);
xor XOR2 (N1405, N1401, N694);
xor XOR2 (N1406, N1400, N360);
buf BUF1 (N1407, N1399);
xor XOR2 (N1408, N1405, N1238);
or OR4 (N1409, N1406, N529, N1220, N858);
or OR4 (N1410, N1397, N340, N725, N413);
or OR2 (N1411, N1403, N784);
not NOT1 (N1412, N1410);
nand NAND2 (N1413, N1412, N539);
xor XOR2 (N1414, N1407, N1202);
buf BUF1 (N1415, N1414);
xor XOR2 (N1416, N1389, N493);
and AND4 (N1417, N1408, N1195, N11, N769);
nand NAND3 (N1418, N1398, N173, N551);
nand NAND2 (N1419, N1404, N610);
buf BUF1 (N1420, N1411);
and AND2 (N1421, N1416, N1227);
and AND3 (N1422, N1418, N588, N276);
not NOT1 (N1423, N1415);
not NOT1 (N1424, N1413);
or OR3 (N1425, N1417, N861, N784);
or OR4 (N1426, N1402, N664, N1183, N1023);
xor XOR2 (N1427, N1424, N958);
nand NAND3 (N1428, N1421, N80, N130);
and AND3 (N1429, N1426, N213, N326);
nand NAND3 (N1430, N1422, N1420, N49);
not NOT1 (N1431, N1339);
not NOT1 (N1432, N1423);
nand NAND3 (N1433, N1431, N878, N1073);
nand NAND2 (N1434, N1433, N1134);
xor XOR2 (N1435, N1425, N164);
nand NAND4 (N1436, N1430, N450, N655, N461);
not NOT1 (N1437, N1419);
nor NOR3 (N1438, N1409, N1292, N225);
nand NAND3 (N1439, N1434, N913, N127);
buf BUF1 (N1440, N1432);
not NOT1 (N1441, N1438);
nor NOR3 (N1442, N1440, N1200, N1015);
xor XOR2 (N1443, N1427, N438);
nand NAND4 (N1444, N1439, N1121, N1336, N307);
nor NOR4 (N1445, N1436, N510, N41, N731);
and AND4 (N1446, N1429, N1140, N1046, N852);
or OR3 (N1447, N1445, N874, N567);
not NOT1 (N1448, N1446);
not NOT1 (N1449, N1443);
nand NAND3 (N1450, N1444, N970, N543);
nand NAND3 (N1451, N1449, N1141, N23);
nand NAND3 (N1452, N1448, N101, N416);
xor XOR2 (N1453, N1387, N1181);
buf BUF1 (N1454, N1441);
nor NOR4 (N1455, N1450, N265, N895, N1078);
or OR3 (N1456, N1447, N757, N668);
and AND2 (N1457, N1437, N15);
or OR3 (N1458, N1435, N738, N330);
buf BUF1 (N1459, N1455);
or OR2 (N1460, N1452, N542);
nor NOR2 (N1461, N1459, N1089);
or OR2 (N1462, N1453, N119);
or OR4 (N1463, N1461, N924, N424, N686);
not NOT1 (N1464, N1458);
nand NAND3 (N1465, N1454, N1075, N836);
and AND4 (N1466, N1463, N480, N137, N488);
and AND2 (N1467, N1442, N1065);
buf BUF1 (N1468, N1456);
nor NOR3 (N1469, N1428, N600, N1299);
xor XOR2 (N1470, N1460, N1045);
not NOT1 (N1471, N1468);
xor XOR2 (N1472, N1457, N722);
nor NOR3 (N1473, N1467, N627, N1116);
or OR3 (N1474, N1462, N797, N291);
or OR4 (N1475, N1474, N153, N540, N1302);
buf BUF1 (N1476, N1471);
nand NAND4 (N1477, N1472, N526, N1176, N1267);
or OR3 (N1478, N1477, N1274, N771);
buf BUF1 (N1479, N1465);
buf BUF1 (N1480, N1469);
not NOT1 (N1481, N1479);
not NOT1 (N1482, N1475);
not NOT1 (N1483, N1473);
nand NAND4 (N1484, N1464, N487, N677, N575);
xor XOR2 (N1485, N1483, N829);
xor XOR2 (N1486, N1466, N244);
xor XOR2 (N1487, N1476, N1062);
xor XOR2 (N1488, N1470, N768);
buf BUF1 (N1489, N1487);
xor XOR2 (N1490, N1451, N828);
not NOT1 (N1491, N1482);
nor NOR2 (N1492, N1478, N1126);
xor XOR2 (N1493, N1485, N824);
buf BUF1 (N1494, N1484);
xor XOR2 (N1495, N1492, N199);
not NOT1 (N1496, N1493);
or OR4 (N1497, N1494, N687, N797, N301);
xor XOR2 (N1498, N1491, N1003);
xor XOR2 (N1499, N1488, N151);
buf BUF1 (N1500, N1481);
and AND4 (N1501, N1486, N699, N247, N602);
buf BUF1 (N1502, N1498);
nand NAND3 (N1503, N1480, N91, N1474);
and AND4 (N1504, N1489, N425, N1112, N507);
and AND4 (N1505, N1500, N585, N1051, N905);
and AND3 (N1506, N1505, N339, N1156);
nand NAND2 (N1507, N1490, N771);
nor NOR4 (N1508, N1503, N323, N1492, N689);
not NOT1 (N1509, N1508);
xor XOR2 (N1510, N1501, N529);
xor XOR2 (N1511, N1506, N349);
buf BUF1 (N1512, N1496);
and AND2 (N1513, N1510, N252);
not NOT1 (N1514, N1497);
xor XOR2 (N1515, N1509, N85);
xor XOR2 (N1516, N1504, N933);
buf BUF1 (N1517, N1516);
nand NAND3 (N1518, N1511, N287, N574);
buf BUF1 (N1519, N1499);
nand NAND2 (N1520, N1502, N973);
or OR2 (N1521, N1495, N716);
and AND4 (N1522, N1513, N400, N975, N672);
xor XOR2 (N1523, N1519, N73);
or OR2 (N1524, N1523, N341);
or OR3 (N1525, N1512, N1476, N1448);
buf BUF1 (N1526, N1521);
and AND2 (N1527, N1522, N413);
xor XOR2 (N1528, N1518, N960);
not NOT1 (N1529, N1514);
nor NOR4 (N1530, N1524, N231, N1445, N1188);
not NOT1 (N1531, N1525);
or OR4 (N1532, N1526, N702, N1318, N1171);
or OR3 (N1533, N1528, N345, N1257);
buf BUF1 (N1534, N1529);
nand NAND2 (N1535, N1507, N49);
and AND3 (N1536, N1527, N1140, N1260);
nor NOR2 (N1537, N1533, N76);
and AND2 (N1538, N1531, N486);
xor XOR2 (N1539, N1517, N811);
xor XOR2 (N1540, N1530, N1284);
or OR2 (N1541, N1534, N584);
or OR2 (N1542, N1515, N1232);
buf BUF1 (N1543, N1536);
and AND2 (N1544, N1535, N585);
or OR2 (N1545, N1538, N1004);
xor XOR2 (N1546, N1541, N1241);
not NOT1 (N1547, N1540);
buf BUF1 (N1548, N1532);
nor NOR3 (N1549, N1543, N889, N1270);
not NOT1 (N1550, N1545);
or OR2 (N1551, N1520, N300);
nor NOR3 (N1552, N1537, N717, N132);
nand NAND3 (N1553, N1542, N592, N1214);
and AND3 (N1554, N1550, N41, N290);
not NOT1 (N1555, N1552);
buf BUF1 (N1556, N1554);
and AND4 (N1557, N1546, N363, N963, N1135);
buf BUF1 (N1558, N1549);
not NOT1 (N1559, N1557);
buf BUF1 (N1560, N1558);
or OR4 (N1561, N1560, N733, N583, N315);
nor NOR2 (N1562, N1556, N1033);
not NOT1 (N1563, N1562);
buf BUF1 (N1564, N1563);
or OR4 (N1565, N1539, N1275, N795, N1560);
buf BUF1 (N1566, N1544);
xor XOR2 (N1567, N1547, N1518);
xor XOR2 (N1568, N1567, N226);
buf BUF1 (N1569, N1568);
and AND4 (N1570, N1559, N633, N343, N1071);
or OR4 (N1571, N1555, N767, N139, N283);
not NOT1 (N1572, N1565);
xor XOR2 (N1573, N1564, N192);
not NOT1 (N1574, N1572);
or OR4 (N1575, N1553, N601, N912, N348);
xor XOR2 (N1576, N1569, N1573);
nor NOR2 (N1577, N1243, N1296);
nand NAND3 (N1578, N1561, N101, N338);
xor XOR2 (N1579, N1574, N1111);
or OR3 (N1580, N1575, N1215, N1432);
not NOT1 (N1581, N1579);
xor XOR2 (N1582, N1571, N45);
nor NOR3 (N1583, N1548, N299, N329);
xor XOR2 (N1584, N1566, N1563);
not NOT1 (N1585, N1578);
nand NAND2 (N1586, N1570, N287);
nor NOR4 (N1587, N1576, N241, N372, N230);
not NOT1 (N1588, N1581);
not NOT1 (N1589, N1580);
xor XOR2 (N1590, N1588, N968);
or OR3 (N1591, N1587, N1226, N996);
buf BUF1 (N1592, N1551);
not NOT1 (N1593, N1584);
nor NOR3 (N1594, N1589, N199, N1318);
and AND3 (N1595, N1583, N714, N1017);
xor XOR2 (N1596, N1592, N256);
buf BUF1 (N1597, N1591);
and AND4 (N1598, N1597, N1539, N1072, N90);
buf BUF1 (N1599, N1582);
and AND3 (N1600, N1593, N55, N447);
buf BUF1 (N1601, N1598);
and AND3 (N1602, N1577, N767, N1500);
xor XOR2 (N1603, N1600, N669);
buf BUF1 (N1604, N1603);
xor XOR2 (N1605, N1596, N1040);
or OR2 (N1606, N1601, N1314);
nand NAND2 (N1607, N1595, N1424);
xor XOR2 (N1608, N1605, N537);
or OR3 (N1609, N1607, N1177, N1234);
xor XOR2 (N1610, N1609, N1047);
xor XOR2 (N1611, N1594, N1088);
or OR2 (N1612, N1606, N358);
and AND4 (N1613, N1585, N82, N1299, N28);
nand NAND4 (N1614, N1613, N348, N792, N1062);
or OR3 (N1615, N1611, N1402, N341);
and AND4 (N1616, N1602, N226, N1095, N1340);
not NOT1 (N1617, N1615);
nor NOR2 (N1618, N1590, N562);
and AND2 (N1619, N1604, N1150);
not NOT1 (N1620, N1610);
buf BUF1 (N1621, N1599);
nor NOR3 (N1622, N1612, N24, N454);
and AND4 (N1623, N1617, N735, N131, N942);
buf BUF1 (N1624, N1621);
or OR4 (N1625, N1614, N293, N339, N742);
xor XOR2 (N1626, N1625, N410);
nand NAND3 (N1627, N1624, N355, N640);
nand NAND3 (N1628, N1618, N1181, N62);
and AND4 (N1629, N1626, N54, N552, N834);
or OR4 (N1630, N1629, N500, N1424, N903);
nand NAND3 (N1631, N1616, N405, N274);
and AND3 (N1632, N1619, N1212, N907);
not NOT1 (N1633, N1628);
nor NOR3 (N1634, N1586, N1160, N1590);
nand NAND4 (N1635, N1620, N950, N416, N264);
buf BUF1 (N1636, N1631);
buf BUF1 (N1637, N1623);
and AND2 (N1638, N1637, N1469);
or OR2 (N1639, N1633, N28);
buf BUF1 (N1640, N1630);
buf BUF1 (N1641, N1638);
not NOT1 (N1642, N1641);
not NOT1 (N1643, N1622);
buf BUF1 (N1644, N1627);
and AND4 (N1645, N1642, N1464, N1110, N157);
nor NOR3 (N1646, N1644, N393, N934);
nand NAND2 (N1647, N1645, N303);
not NOT1 (N1648, N1634);
and AND2 (N1649, N1636, N372);
xor XOR2 (N1650, N1649, N127);
not NOT1 (N1651, N1647);
xor XOR2 (N1652, N1643, N247);
buf BUF1 (N1653, N1652);
nor NOR3 (N1654, N1650, N1143, N109);
nand NAND4 (N1655, N1654, N786, N1425, N404);
nor NOR2 (N1656, N1640, N30);
buf BUF1 (N1657, N1651);
nand NAND4 (N1658, N1648, N410, N1547, N33);
not NOT1 (N1659, N1655);
or OR3 (N1660, N1608, N1287, N1158);
and AND2 (N1661, N1635, N576);
not NOT1 (N1662, N1660);
buf BUF1 (N1663, N1658);
not NOT1 (N1664, N1661);
nor NOR2 (N1665, N1659, N1656);
or OR3 (N1666, N1524, N370, N1332);
and AND2 (N1667, N1663, N990);
buf BUF1 (N1668, N1667);
nand NAND3 (N1669, N1657, N1466, N461);
nand NAND3 (N1670, N1664, N404, N543);
nor NOR3 (N1671, N1632, N406, N458);
nand NAND4 (N1672, N1669, N1189, N627, N625);
xor XOR2 (N1673, N1639, N367);
nor NOR4 (N1674, N1670, N43, N1015, N63);
nor NOR3 (N1675, N1672, N1412, N1007);
not NOT1 (N1676, N1671);
nor NOR4 (N1677, N1675, N577, N177, N13);
not NOT1 (N1678, N1662);
or OR3 (N1679, N1665, N207, N599);
nand NAND3 (N1680, N1677, N597, N1006);
xor XOR2 (N1681, N1666, N134);
nor NOR3 (N1682, N1653, N291, N808);
xor XOR2 (N1683, N1674, N1113);
xor XOR2 (N1684, N1683, N1119);
xor XOR2 (N1685, N1681, N1107);
buf BUF1 (N1686, N1646);
nor NOR2 (N1687, N1678, N409);
not NOT1 (N1688, N1685);
nand NAND4 (N1689, N1673, N1439, N774, N1538);
nand NAND2 (N1690, N1688, N826);
nor NOR2 (N1691, N1682, N1045);
buf BUF1 (N1692, N1679);
nand NAND4 (N1693, N1676, N776, N62, N528);
nor NOR4 (N1694, N1687, N1192, N972, N663);
or OR3 (N1695, N1691, N610, N149);
xor XOR2 (N1696, N1693, N582);
buf BUF1 (N1697, N1694);
not NOT1 (N1698, N1684);
buf BUF1 (N1699, N1696);
nand NAND4 (N1700, N1690, N644, N433, N396);
xor XOR2 (N1701, N1680, N254);
not NOT1 (N1702, N1668);
xor XOR2 (N1703, N1689, N619);
xor XOR2 (N1704, N1692, N1228);
not NOT1 (N1705, N1698);
and AND2 (N1706, N1703, N697);
buf BUF1 (N1707, N1701);
xor XOR2 (N1708, N1700, N786);
not NOT1 (N1709, N1706);
not NOT1 (N1710, N1709);
nand NAND3 (N1711, N1705, N112, N13);
nor NOR4 (N1712, N1697, N674, N762, N782);
nand NAND2 (N1713, N1702, N1369);
and AND2 (N1714, N1699, N1027);
and AND2 (N1715, N1714, N1488);
nor NOR2 (N1716, N1713, N451);
and AND2 (N1717, N1708, N1245);
nand NAND2 (N1718, N1711, N381);
and AND2 (N1719, N1686, N256);
xor XOR2 (N1720, N1716, N412);
nand NAND4 (N1721, N1707, N58, N991, N129);
nand NAND3 (N1722, N1715, N776, N10);
xor XOR2 (N1723, N1717, N213);
or OR4 (N1724, N1718, N1400, N1631, N399);
xor XOR2 (N1725, N1719, N1252);
xor XOR2 (N1726, N1695, N343);
xor XOR2 (N1727, N1710, N1341);
xor XOR2 (N1728, N1725, N340);
or OR2 (N1729, N1712, N1006);
nand NAND4 (N1730, N1704, N1208, N765, N1638);
xor XOR2 (N1731, N1730, N807);
nand NAND3 (N1732, N1731, N652, N1515);
nand NAND2 (N1733, N1721, N776);
nand NAND3 (N1734, N1720, N1555, N289);
xor XOR2 (N1735, N1722, N655);
nor NOR2 (N1736, N1734, N684);
and AND3 (N1737, N1727, N1318, N55);
nand NAND2 (N1738, N1736, N629);
buf BUF1 (N1739, N1729);
nand NAND4 (N1740, N1728, N211, N790, N446);
nand NAND4 (N1741, N1733, N1681, N1254, N1315);
nand NAND2 (N1742, N1740, N824);
nand NAND3 (N1743, N1735, N1085, N488);
not NOT1 (N1744, N1738);
and AND2 (N1745, N1741, N1625);
and AND2 (N1746, N1744, N427);
and AND2 (N1747, N1732, N1405);
and AND4 (N1748, N1745, N1, N1524, N138);
nor NOR3 (N1749, N1743, N151, N760);
not NOT1 (N1750, N1746);
not NOT1 (N1751, N1739);
or OR3 (N1752, N1723, N221, N863);
nand NAND4 (N1753, N1750, N528, N1268, N882);
and AND3 (N1754, N1753, N511, N870);
nand NAND3 (N1755, N1742, N385, N1400);
not NOT1 (N1756, N1749);
or OR3 (N1757, N1726, N1343, N742);
buf BUF1 (N1758, N1724);
nor NOR3 (N1759, N1748, N1534, N1083);
or OR4 (N1760, N1759, N538, N454, N673);
nand NAND2 (N1761, N1751, N1180);
nand NAND3 (N1762, N1758, N12, N1096);
nand NAND2 (N1763, N1755, N664);
nor NOR4 (N1764, N1747, N86, N978, N865);
and AND3 (N1765, N1754, N1411, N1206);
and AND4 (N1766, N1765, N217, N446, N1704);
and AND3 (N1767, N1737, N1589, N726);
nand NAND4 (N1768, N1767, N1036, N575, N1303);
not NOT1 (N1769, N1752);
or OR3 (N1770, N1766, N220, N389);
nand NAND4 (N1771, N1770, N136, N1464, N777);
nor NOR2 (N1772, N1768, N1123);
buf BUF1 (N1773, N1756);
and AND2 (N1774, N1771, N725);
nand NAND2 (N1775, N1760, N1244);
not NOT1 (N1776, N1773);
buf BUF1 (N1777, N1776);
xor XOR2 (N1778, N1762, N83);
and AND3 (N1779, N1774, N76, N502);
not NOT1 (N1780, N1761);
buf BUF1 (N1781, N1763);
not NOT1 (N1782, N1780);
not NOT1 (N1783, N1764);
xor XOR2 (N1784, N1779, N502);
buf BUF1 (N1785, N1782);
buf BUF1 (N1786, N1781);
nor NOR2 (N1787, N1777, N1414);
nor NOR4 (N1788, N1757, N659, N1707, N394);
and AND2 (N1789, N1785, N726);
and AND4 (N1790, N1769, N1259, N208, N1204);
not NOT1 (N1791, N1775);
nand NAND4 (N1792, N1778, N107, N1122, N1595);
xor XOR2 (N1793, N1790, N653);
nand NAND2 (N1794, N1772, N268);
or OR4 (N1795, N1794, N1730, N965, N728);
buf BUF1 (N1796, N1786);
and AND3 (N1797, N1792, N508, N90);
not NOT1 (N1798, N1784);
and AND2 (N1799, N1793, N1540);
not NOT1 (N1800, N1788);
and AND4 (N1801, N1800, N624, N1311, N91);
not NOT1 (N1802, N1791);
nor NOR3 (N1803, N1801, N944, N427);
xor XOR2 (N1804, N1789, N784);
and AND3 (N1805, N1798, N420, N916);
not NOT1 (N1806, N1795);
or OR4 (N1807, N1803, N1007, N1771, N806);
xor XOR2 (N1808, N1805, N1464);
and AND3 (N1809, N1796, N1153, N1240);
nor NOR2 (N1810, N1808, N1306);
buf BUF1 (N1811, N1799);
and AND2 (N1812, N1807, N1151);
nor NOR2 (N1813, N1812, N1285);
or OR4 (N1814, N1809, N836, N1214, N432);
nor NOR3 (N1815, N1783, N314, N253);
nand NAND2 (N1816, N1802, N900);
or OR2 (N1817, N1806, N1188);
not NOT1 (N1818, N1813);
nor NOR2 (N1819, N1797, N1503);
nor NOR2 (N1820, N1816, N117);
or OR3 (N1821, N1817, N1219, N501);
nand NAND4 (N1822, N1804, N1749, N327, N1234);
or OR3 (N1823, N1822, N800, N324);
not NOT1 (N1824, N1820);
buf BUF1 (N1825, N1810);
and AND4 (N1826, N1787, N1140, N1650, N1452);
xor XOR2 (N1827, N1819, N93);
nand NAND2 (N1828, N1815, N724);
xor XOR2 (N1829, N1821, N1416);
not NOT1 (N1830, N1827);
or OR4 (N1831, N1830, N677, N1610, N175);
not NOT1 (N1832, N1828);
nand NAND3 (N1833, N1825, N1495, N955);
nand NAND4 (N1834, N1826, N1621, N955, N396);
nand NAND4 (N1835, N1811, N1415, N121, N358);
buf BUF1 (N1836, N1824);
not NOT1 (N1837, N1833);
nor NOR3 (N1838, N1835, N77, N1834);
not NOT1 (N1839, N1467);
nor NOR3 (N1840, N1837, N282, N451);
buf BUF1 (N1841, N1814);
and AND3 (N1842, N1836, N604, N851);
nand NAND3 (N1843, N1840, N182, N574);
or OR4 (N1844, N1831, N1399, N1328, N1282);
and AND4 (N1845, N1832, N563, N1534, N554);
buf BUF1 (N1846, N1823);
xor XOR2 (N1847, N1842, N220);
and AND2 (N1848, N1845, N1133);
not NOT1 (N1849, N1843);
buf BUF1 (N1850, N1847);
or OR4 (N1851, N1846, N1217, N271, N662);
or OR3 (N1852, N1838, N594, N210);
nor NOR2 (N1853, N1850, N530);
or OR2 (N1854, N1829, N786);
not NOT1 (N1855, N1852);
not NOT1 (N1856, N1855);
nor NOR2 (N1857, N1841, N24);
not NOT1 (N1858, N1844);
or OR2 (N1859, N1857, N351);
not NOT1 (N1860, N1859);
xor XOR2 (N1861, N1839, N1561);
nor NOR3 (N1862, N1860, N500, N1545);
and AND4 (N1863, N1851, N1806, N296, N1123);
buf BUF1 (N1864, N1848);
nor NOR4 (N1865, N1864, N1797, N735, N1712);
xor XOR2 (N1866, N1863, N707);
nand NAND2 (N1867, N1853, N1158);
nand NAND4 (N1868, N1865, N1066, N1460, N1165);
nand NAND4 (N1869, N1856, N1147, N416, N1137);
nand NAND3 (N1870, N1869, N308, N1516);
nor NOR2 (N1871, N1854, N1091);
not NOT1 (N1872, N1818);
not NOT1 (N1873, N1868);
or OR2 (N1874, N1873, N1107);
nor NOR3 (N1875, N1861, N1418, N760);
nand NAND3 (N1876, N1866, N1080, N1582);
xor XOR2 (N1877, N1875, N1536);
and AND2 (N1878, N1871, N406);
nor NOR3 (N1879, N1874, N305, N1007);
nand NAND4 (N1880, N1867, N879, N56, N1805);
or OR4 (N1881, N1878, N1460, N936, N1079);
or OR4 (N1882, N1870, N522, N876, N1788);
and AND4 (N1883, N1879, N1636, N1052, N447);
buf BUF1 (N1884, N1881);
or OR4 (N1885, N1849, N349, N1576, N1706);
nand NAND2 (N1886, N1862, N262);
or OR3 (N1887, N1880, N192, N1066);
not NOT1 (N1888, N1886);
xor XOR2 (N1889, N1882, N124);
not NOT1 (N1890, N1877);
nand NAND3 (N1891, N1889, N1648, N317);
xor XOR2 (N1892, N1891, N1875);
nor NOR2 (N1893, N1858, N1604);
not NOT1 (N1894, N1876);
nand NAND2 (N1895, N1872, N856);
and AND3 (N1896, N1895, N812, N1546);
buf BUF1 (N1897, N1894);
or OR3 (N1898, N1885, N169, N1106);
not NOT1 (N1899, N1892);
buf BUF1 (N1900, N1888);
nand NAND3 (N1901, N1898, N1515, N48);
xor XOR2 (N1902, N1900, N352);
xor XOR2 (N1903, N1893, N1710);
nand NAND4 (N1904, N1890, N578, N1647, N1010);
xor XOR2 (N1905, N1901, N1425);
nand NAND4 (N1906, N1897, N505, N1273, N128);
or OR2 (N1907, N1884, N748);
xor XOR2 (N1908, N1904, N719);
not NOT1 (N1909, N1905);
xor XOR2 (N1910, N1896, N553);
or OR4 (N1911, N1903, N692, N960, N229);
and AND2 (N1912, N1887, N859);
not NOT1 (N1913, N1911);
xor XOR2 (N1914, N1910, N1085);
or OR4 (N1915, N1907, N1783, N300, N800);
or OR2 (N1916, N1899, N793);
xor XOR2 (N1917, N1906, N675);
buf BUF1 (N1918, N1916);
buf BUF1 (N1919, N1914);
buf BUF1 (N1920, N1913);
or OR3 (N1921, N1902, N1529, N1791);
or OR4 (N1922, N1919, N945, N1800, N844);
or OR3 (N1923, N1909, N694, N574);
or OR4 (N1924, N1918, N1141, N699, N361);
nand NAND2 (N1925, N1922, N1016);
nor NOR4 (N1926, N1912, N827, N1675, N1907);
or OR2 (N1927, N1917, N1396);
buf BUF1 (N1928, N1925);
buf BUF1 (N1929, N1924);
nor NOR3 (N1930, N1923, N688, N866);
nand NAND4 (N1931, N1929, N1587, N558, N271);
buf BUF1 (N1932, N1908);
xor XOR2 (N1933, N1930, N1220);
xor XOR2 (N1934, N1932, N499);
buf BUF1 (N1935, N1915);
or OR2 (N1936, N1931, N182);
xor XOR2 (N1937, N1935, N216);
xor XOR2 (N1938, N1934, N822);
or OR3 (N1939, N1928, N1506, N1293);
nor NOR4 (N1940, N1938, N264, N1555, N1853);
nand NAND3 (N1941, N1940, N1688, N1559);
xor XOR2 (N1942, N1926, N358);
or OR2 (N1943, N1936, N1428);
nand NAND3 (N1944, N1942, N924, N1582);
xor XOR2 (N1945, N1944, N101);
xor XOR2 (N1946, N1921, N1860);
xor XOR2 (N1947, N1927, N568);
xor XOR2 (N1948, N1939, N261);
nor NOR3 (N1949, N1883, N860, N800);
xor XOR2 (N1950, N1920, N1394);
and AND4 (N1951, N1950, N793, N774, N737);
or OR3 (N1952, N1937, N1914, N556);
buf BUF1 (N1953, N1947);
xor XOR2 (N1954, N1952, N568);
nand NAND4 (N1955, N1941, N320, N1280, N412);
buf BUF1 (N1956, N1949);
xor XOR2 (N1957, N1946, N1340);
buf BUF1 (N1958, N1955);
xor XOR2 (N1959, N1943, N695);
nor NOR4 (N1960, N1945, N716, N698, N1828);
not NOT1 (N1961, N1951);
buf BUF1 (N1962, N1960);
nor NOR3 (N1963, N1954, N735, N1893);
nor NOR3 (N1964, N1956, N1483, N14);
xor XOR2 (N1965, N1959, N688);
nor NOR4 (N1966, N1965, N1896, N817, N708);
and AND4 (N1967, N1953, N1327, N365, N1858);
and AND4 (N1968, N1963, N747, N1531, N539);
and AND2 (N1969, N1958, N1364);
xor XOR2 (N1970, N1964, N1786);
nand NAND4 (N1971, N1970, N862, N1156, N127);
nand NAND4 (N1972, N1961, N1830, N442, N1554);
or OR2 (N1973, N1933, N1688);
nor NOR3 (N1974, N1968, N957, N1720);
buf BUF1 (N1975, N1948);
nand NAND3 (N1976, N1962, N965, N65);
and AND4 (N1977, N1966, N1462, N894, N1498);
nor NOR4 (N1978, N1976, N141, N582, N1339);
nand NAND4 (N1979, N1971, N1389, N110, N1600);
buf BUF1 (N1980, N1957);
or OR3 (N1981, N1969, N1850, N1419);
nor NOR2 (N1982, N1972, N645);
nor NOR4 (N1983, N1981, N1338, N1140, N387);
nor NOR3 (N1984, N1979, N958, N633);
nor NOR4 (N1985, N1980, N868, N149, N418);
xor XOR2 (N1986, N1967, N268);
and AND3 (N1987, N1978, N1458, N1512);
and AND2 (N1988, N1973, N692);
nor NOR3 (N1989, N1974, N1193, N648);
or OR2 (N1990, N1987, N1203);
xor XOR2 (N1991, N1985, N1535);
nand NAND3 (N1992, N1982, N361, N436);
or OR3 (N1993, N1977, N1862, N123);
nand NAND2 (N1994, N1983, N1004);
xor XOR2 (N1995, N1975, N573);
buf BUF1 (N1996, N1995);
or OR4 (N1997, N1996, N1860, N1081, N1750);
xor XOR2 (N1998, N1990, N1983);
or OR2 (N1999, N1991, N1117);
not NOT1 (N2000, N1992);
nor NOR2 (N2001, N1984, N21);
xor XOR2 (N2002, N2001, N1017);
not NOT1 (N2003, N1994);
nor NOR2 (N2004, N1993, N1863);
buf BUF1 (N2005, N2004);
xor XOR2 (N2006, N1997, N518);
or OR2 (N2007, N2003, N1083);
buf BUF1 (N2008, N1999);
or OR2 (N2009, N2002, N1025);
nand NAND2 (N2010, N2000, N411);
and AND3 (N2011, N2007, N788, N561);
xor XOR2 (N2012, N2009, N874);
nand NAND2 (N2013, N1988, N1264);
not NOT1 (N2014, N2010);
nor NOR2 (N2015, N1989, N477);
nand NAND2 (N2016, N1986, N1926);
or OR3 (N2017, N2008, N659, N498);
nand NAND3 (N2018, N2006, N1985, N1190);
buf BUF1 (N2019, N2011);
nor NOR2 (N2020, N2005, N1355);
buf BUF1 (N2021, N2014);
buf BUF1 (N2022, N2018);
buf BUF1 (N2023, N2022);
or OR4 (N2024, N2017, N858, N314, N1065);
nand NAND2 (N2025, N2013, N85);
not NOT1 (N2026, N2023);
not NOT1 (N2027, N2015);
xor XOR2 (N2028, N2021, N303);
nor NOR3 (N2029, N2027, N807, N1449);
buf BUF1 (N2030, N2016);
nor NOR4 (N2031, N2030, N24, N1598, N1506);
not NOT1 (N2032, N2026);
and AND2 (N2033, N2031, N448);
not NOT1 (N2034, N2020);
or OR2 (N2035, N2033, N579);
not NOT1 (N2036, N1998);
not NOT1 (N2037, N2032);
xor XOR2 (N2038, N2012, N698);
xor XOR2 (N2039, N2035, N645);
xor XOR2 (N2040, N2028, N453);
nor NOR2 (N2041, N2024, N18);
and AND4 (N2042, N2034, N1518, N43, N1133);
xor XOR2 (N2043, N2041, N220);
xor XOR2 (N2044, N2042, N903);
and AND2 (N2045, N2037, N1882);
and AND2 (N2046, N2043, N53);
or OR4 (N2047, N2039, N2043, N382, N891);
nor NOR2 (N2048, N2036, N1304);
buf BUF1 (N2049, N2047);
not NOT1 (N2050, N2048);
buf BUF1 (N2051, N2046);
xor XOR2 (N2052, N2040, N379);
not NOT1 (N2053, N2029);
nor NOR4 (N2054, N2045, N1128, N1733, N1304);
and AND3 (N2055, N2025, N886, N1724);
xor XOR2 (N2056, N2053, N1558);
nand NAND2 (N2057, N2054, N779);
xor XOR2 (N2058, N2019, N608);
or OR2 (N2059, N2056, N1314);
nor NOR4 (N2060, N2059, N1740, N671, N1995);
nand NAND4 (N2061, N2060, N1388, N480, N1070);
nand NAND4 (N2062, N2051, N1580, N1246, N988);
not NOT1 (N2063, N2052);
xor XOR2 (N2064, N2062, N315);
nor NOR4 (N2065, N2044, N867, N561, N1826);
nor NOR2 (N2066, N2050, N1470);
xor XOR2 (N2067, N2066, N771);
and AND4 (N2068, N2063, N2019, N1582, N733);
not NOT1 (N2069, N2067);
nand NAND3 (N2070, N2069, N800, N1534);
not NOT1 (N2071, N2065);
xor XOR2 (N2072, N2057, N996);
nand NAND4 (N2073, N2058, N1912, N1999, N533);
not NOT1 (N2074, N2071);
xor XOR2 (N2075, N2055, N2024);
xor XOR2 (N2076, N2061, N76);
buf BUF1 (N2077, N2072);
or OR4 (N2078, N2064, N446, N840, N1022);
and AND2 (N2079, N2068, N1416);
xor XOR2 (N2080, N2079, N825);
and AND4 (N2081, N2075, N274, N1258, N397);
and AND2 (N2082, N2078, N270);
xor XOR2 (N2083, N2070, N918);
and AND4 (N2084, N2049, N837, N813, N545);
nand NAND2 (N2085, N2082, N336);
or OR4 (N2086, N2080, N1662, N1915, N591);
buf BUF1 (N2087, N2076);
nand NAND2 (N2088, N2038, N1238);
buf BUF1 (N2089, N2084);
not NOT1 (N2090, N2086);
nand NAND3 (N2091, N2088, N298, N1172);
and AND2 (N2092, N2085, N244);
or OR2 (N2093, N2091, N575);
buf BUF1 (N2094, N2074);
or OR4 (N2095, N2077, N224, N758, N1628);
nor NOR4 (N2096, N2090, N1431, N132, N1373);
not NOT1 (N2097, N2081);
buf BUF1 (N2098, N2083);
xor XOR2 (N2099, N2096, N1440);
or OR4 (N2100, N2092, N1631, N498, N2060);
not NOT1 (N2101, N2100);
and AND2 (N2102, N2094, N294);
not NOT1 (N2103, N2101);
and AND4 (N2104, N2093, N1314, N1907, N1703);
nand NAND2 (N2105, N2097, N37);
nand NAND4 (N2106, N2095, N383, N1298, N1973);
xor XOR2 (N2107, N2089, N955);
nand NAND2 (N2108, N2102, N664);
xor XOR2 (N2109, N2104, N214);
or OR4 (N2110, N2087, N394, N567, N869);
buf BUF1 (N2111, N2098);
nor NOR2 (N2112, N2099, N1793);
and AND4 (N2113, N2109, N1726, N1568, N129);
or OR3 (N2114, N2108, N662, N1996);
buf BUF1 (N2115, N2103);
not NOT1 (N2116, N2112);
and AND4 (N2117, N2115, N220, N1087, N162);
and AND3 (N2118, N2117, N1805, N1053);
buf BUF1 (N2119, N2110);
and AND2 (N2120, N2116, N1899);
nand NAND2 (N2121, N2073, N415);
not NOT1 (N2122, N2105);
nor NOR2 (N2123, N2120, N320);
buf BUF1 (N2124, N2119);
nor NOR4 (N2125, N2114, N495, N1915, N894);
xor XOR2 (N2126, N2125, N1807);
not NOT1 (N2127, N2124);
nand NAND4 (N2128, N2107, N1505, N214, N439);
xor XOR2 (N2129, N2106, N22);
xor XOR2 (N2130, N2128, N1973);
buf BUF1 (N2131, N2126);
nand NAND2 (N2132, N2122, N1430);
buf BUF1 (N2133, N2111);
and AND3 (N2134, N2130, N534, N1581);
nand NAND2 (N2135, N2132, N1767);
buf BUF1 (N2136, N2123);
xor XOR2 (N2137, N2127, N1997);
nand NAND2 (N2138, N2133, N1165);
or OR4 (N2139, N2113, N1199, N872, N1431);
buf BUF1 (N2140, N2129);
nand NAND2 (N2141, N2140, N61);
not NOT1 (N2142, N2136);
or OR3 (N2143, N2131, N108, N1872);
buf BUF1 (N2144, N2118);
and AND3 (N2145, N2137, N48, N248);
nand NAND3 (N2146, N2141, N854, N636);
and AND3 (N2147, N2134, N1957, N48);
buf BUF1 (N2148, N2138);
and AND3 (N2149, N2144, N1126, N1911);
not NOT1 (N2150, N2135);
not NOT1 (N2151, N2143);
or OR4 (N2152, N2139, N851, N1117, N206);
and AND4 (N2153, N2148, N1720, N345, N66);
not NOT1 (N2154, N2153);
or OR2 (N2155, N2145, N1690);
nor NOR2 (N2156, N2154, N1681);
xor XOR2 (N2157, N2146, N1938);
xor XOR2 (N2158, N2155, N1954);
xor XOR2 (N2159, N2121, N780);
not NOT1 (N2160, N2151);
xor XOR2 (N2161, N2159, N38);
xor XOR2 (N2162, N2156, N1379);
and AND4 (N2163, N2161, N438, N1966, N1442);
and AND3 (N2164, N2163, N317, N172);
xor XOR2 (N2165, N2164, N733);
not NOT1 (N2166, N2160);
and AND4 (N2167, N2142, N1616, N1468, N268);
or OR4 (N2168, N2167, N1440, N1571, N1677);
or OR2 (N2169, N2165, N1547);
and AND2 (N2170, N2158, N1642);
xor XOR2 (N2171, N2169, N1608);
nand NAND4 (N2172, N2168, N903, N1027, N881);
nor NOR2 (N2173, N2171, N421);
or OR4 (N2174, N2147, N1441, N377, N1014);
not NOT1 (N2175, N2173);
or OR2 (N2176, N2166, N2081);
or OR3 (N2177, N2152, N1396, N137);
nor NOR4 (N2178, N2174, N622, N138, N1740);
or OR2 (N2179, N2177, N1732);
nor NOR2 (N2180, N2170, N1527);
and AND2 (N2181, N2178, N2041);
or OR2 (N2182, N2149, N1175);
and AND2 (N2183, N2181, N1966);
buf BUF1 (N2184, N2172);
nor NOR4 (N2185, N2175, N39, N1792, N1929);
xor XOR2 (N2186, N2157, N1017);
buf BUF1 (N2187, N2183);
and AND3 (N2188, N2150, N929, N339);
not NOT1 (N2189, N2184);
nand NAND4 (N2190, N2188, N994, N1425, N7);
xor XOR2 (N2191, N2182, N1608);
nand NAND4 (N2192, N2176, N953, N168, N1807);
not NOT1 (N2193, N2187);
xor XOR2 (N2194, N2162, N1040);
or OR2 (N2195, N2186, N321);
buf BUF1 (N2196, N2190);
nand NAND3 (N2197, N2180, N1679, N1304);
and AND2 (N2198, N2189, N366);
xor XOR2 (N2199, N2191, N757);
nor NOR3 (N2200, N2197, N368, N1746);
or OR4 (N2201, N2193, N1789, N2077, N589);
nand NAND4 (N2202, N2198, N1375, N1410, N1583);
xor XOR2 (N2203, N2201, N468);
buf BUF1 (N2204, N2192);
xor XOR2 (N2205, N2203, N312);
or OR2 (N2206, N2179, N956);
and AND2 (N2207, N2194, N1774);
nand NAND4 (N2208, N2196, N1512, N1122, N1422);
and AND2 (N2209, N2205, N523);
and AND4 (N2210, N2195, N178, N362, N911);
and AND2 (N2211, N2202, N2152);
and AND2 (N2212, N2210, N919);
nor NOR4 (N2213, N2204, N1643, N2115, N2064);
nand NAND2 (N2214, N2211, N1093);
nand NAND3 (N2215, N2207, N1402, N708);
and AND4 (N2216, N2208, N1970, N1108, N548);
or OR2 (N2217, N2199, N1316);
nand NAND2 (N2218, N2216, N983);
and AND2 (N2219, N2218, N1415);
buf BUF1 (N2220, N2215);
nor NOR2 (N2221, N2217, N2044);
and AND3 (N2222, N2221, N1629, N645);
or OR3 (N2223, N2213, N1174, N1944);
xor XOR2 (N2224, N2206, N1517);
or OR3 (N2225, N2200, N1388, N1864);
and AND4 (N2226, N2220, N703, N20, N432);
buf BUF1 (N2227, N2222);
buf BUF1 (N2228, N2185);
not NOT1 (N2229, N2225);
not NOT1 (N2230, N2209);
or OR2 (N2231, N2228, N1371);
xor XOR2 (N2232, N2230, N1800);
xor XOR2 (N2233, N2219, N309);
or OR3 (N2234, N2227, N297, N320);
not NOT1 (N2235, N2232);
nor NOR3 (N2236, N2223, N329, N1320);
and AND4 (N2237, N2229, N1040, N545, N128);
nor NOR2 (N2238, N2234, N337);
buf BUF1 (N2239, N2212);
or OR4 (N2240, N2239, N700, N1008, N1837);
or OR2 (N2241, N2235, N2014);
nor NOR3 (N2242, N2236, N2055, N1514);
nand NAND2 (N2243, N2226, N797);
nand NAND2 (N2244, N2238, N372);
xor XOR2 (N2245, N2214, N107);
xor XOR2 (N2246, N2242, N487);
or OR2 (N2247, N2241, N2186);
and AND3 (N2248, N2244, N1455, N1461);
buf BUF1 (N2249, N2233);
buf BUF1 (N2250, N2248);
and AND4 (N2251, N2240, N385, N1213, N1445);
or OR4 (N2252, N2231, N1150, N19, N580);
xor XOR2 (N2253, N2249, N611);
or OR4 (N2254, N2247, N1894, N1214, N582);
and AND4 (N2255, N2253, N1024, N76, N601);
nor NOR2 (N2256, N2237, N2061);
or OR3 (N2257, N2256, N2097, N1422);
nor NOR3 (N2258, N2224, N721, N1019);
and AND4 (N2259, N2243, N28, N2121, N2157);
or OR2 (N2260, N2259, N495);
nor NOR2 (N2261, N2245, N1765);
xor XOR2 (N2262, N2255, N1728);
and AND4 (N2263, N2254, N1505, N1620, N1977);
nand NAND2 (N2264, N2252, N675);
or OR3 (N2265, N2251, N383, N841);
buf BUF1 (N2266, N2265);
xor XOR2 (N2267, N2264, N101);
and AND2 (N2268, N2250, N1476);
buf BUF1 (N2269, N2267);
not NOT1 (N2270, N2260);
buf BUF1 (N2271, N2246);
buf BUF1 (N2272, N2258);
buf BUF1 (N2273, N2263);
buf BUF1 (N2274, N2268);
nor NOR2 (N2275, N2269, N1781);
not NOT1 (N2276, N2261);
and AND3 (N2277, N2274, N1056, N2032);
nand NAND2 (N2278, N2262, N2141);
not NOT1 (N2279, N2271);
xor XOR2 (N2280, N2279, N953);
nand NAND2 (N2281, N2280, N36);
not NOT1 (N2282, N2275);
or OR3 (N2283, N2281, N2015, N57);
nand NAND3 (N2284, N2257, N768, N1451);
nand NAND3 (N2285, N2276, N175, N1758);
buf BUF1 (N2286, N2277);
nand NAND4 (N2287, N2286, N1085, N2000, N942);
not NOT1 (N2288, N2282);
or OR3 (N2289, N2278, N1367, N2243);
xor XOR2 (N2290, N2289, N561);
nand NAND2 (N2291, N2272, N656);
buf BUF1 (N2292, N2273);
nor NOR4 (N2293, N2285, N939, N1774, N1935);
buf BUF1 (N2294, N2290);
or OR3 (N2295, N2292, N665, N1590);
not NOT1 (N2296, N2287);
xor XOR2 (N2297, N2284, N307);
not NOT1 (N2298, N2295);
nor NOR2 (N2299, N2294, N1124);
xor XOR2 (N2300, N2291, N67);
nand NAND2 (N2301, N2283, N1874);
nor NOR3 (N2302, N2270, N385, N1535);
not NOT1 (N2303, N2296);
nor NOR2 (N2304, N2298, N368);
buf BUF1 (N2305, N2302);
xor XOR2 (N2306, N2303, N1986);
nor NOR3 (N2307, N2293, N498, N1345);
nand NAND4 (N2308, N2299, N2, N1103, N1172);
nand NAND4 (N2309, N2305, N1799, N1941, N1273);
or OR3 (N2310, N2300, N829, N1515);
not NOT1 (N2311, N2307);
xor XOR2 (N2312, N2308, N1576);
buf BUF1 (N2313, N2311);
or OR2 (N2314, N2309, N1663);
nor NOR2 (N2315, N2304, N2140);
buf BUF1 (N2316, N2288);
nor NOR3 (N2317, N2313, N1526, N1219);
and AND3 (N2318, N2314, N1384, N2178);
and AND4 (N2319, N2266, N285, N1159, N783);
or OR2 (N2320, N2306, N184);
and AND2 (N2321, N2315, N166);
buf BUF1 (N2322, N2301);
and AND2 (N2323, N2317, N603);
not NOT1 (N2324, N2310);
buf BUF1 (N2325, N2324);
and AND2 (N2326, N2325, N1169);
buf BUF1 (N2327, N2318);
and AND2 (N2328, N2327, N2003);
nor NOR3 (N2329, N2320, N1899, N1655);
or OR3 (N2330, N2319, N1760, N1094);
nand NAND3 (N2331, N2330, N2118, N2175);
nand NAND2 (N2332, N2326, N2213);
nand NAND4 (N2333, N2323, N1942, N1533, N2272);
nor NOR2 (N2334, N2312, N1834);
nand NAND4 (N2335, N2322, N242, N1569, N11);
or OR4 (N2336, N2331, N1378, N2128, N1455);
not NOT1 (N2337, N2336);
xor XOR2 (N2338, N2337, N1513);
xor XOR2 (N2339, N2329, N301);
or OR4 (N2340, N2328, N1099, N687, N1299);
buf BUF1 (N2341, N2332);
buf BUF1 (N2342, N2339);
xor XOR2 (N2343, N2334, N1688);
or OR2 (N2344, N2297, N2052);
xor XOR2 (N2345, N2344, N1220);
or OR4 (N2346, N2333, N1778, N1399, N2174);
nand NAND4 (N2347, N2345, N1019, N1209, N658);
not NOT1 (N2348, N2342);
buf BUF1 (N2349, N2338);
not NOT1 (N2350, N2340);
or OR4 (N2351, N2349, N1359, N1351, N1171);
and AND2 (N2352, N2341, N1995);
not NOT1 (N2353, N2335);
nor NOR2 (N2354, N2316, N1264);
nand NAND4 (N2355, N2348, N962, N598, N1259);
or OR4 (N2356, N2353, N1702, N1408, N720);
or OR3 (N2357, N2356, N1942, N1789);
not NOT1 (N2358, N2346);
and AND3 (N2359, N2347, N223, N1359);
buf BUF1 (N2360, N2355);
and AND2 (N2361, N2321, N1520);
or OR2 (N2362, N2357, N1046);
nand NAND2 (N2363, N2358, N76);
xor XOR2 (N2364, N2361, N503);
not NOT1 (N2365, N2362);
or OR2 (N2366, N2351, N692);
nor NOR3 (N2367, N2360, N1971, N200);
xor XOR2 (N2368, N2365, N1761);
nand NAND3 (N2369, N2350, N965, N909);
nor NOR4 (N2370, N2368, N173, N174, N2225);
xor XOR2 (N2371, N2370, N1600);
and AND3 (N2372, N2359, N692, N553);
nand NAND4 (N2373, N2369, N179, N807, N1878);
or OR4 (N2374, N2343, N86, N1167, N1870);
and AND4 (N2375, N2363, N1588, N698, N863);
xor XOR2 (N2376, N2374, N943);
xor XOR2 (N2377, N2375, N1551);
nand NAND3 (N2378, N2376, N2322, N591);
xor XOR2 (N2379, N2378, N1815);
and AND4 (N2380, N2379, N1759, N1568, N1328);
nand NAND2 (N2381, N2373, N850);
and AND3 (N2382, N2364, N516, N1131);
buf BUF1 (N2383, N2382);
not NOT1 (N2384, N2380);
buf BUF1 (N2385, N2372);
not NOT1 (N2386, N2383);
or OR2 (N2387, N2352, N1796);
xor XOR2 (N2388, N2366, N238);
buf BUF1 (N2389, N2387);
buf BUF1 (N2390, N2371);
nand NAND3 (N2391, N2389, N1810, N1064);
buf BUF1 (N2392, N2367);
xor XOR2 (N2393, N2381, N1214);
and AND2 (N2394, N2386, N135);
nand NAND4 (N2395, N2391, N1122, N1867, N1130);
not NOT1 (N2396, N2388);
buf BUF1 (N2397, N2395);
not NOT1 (N2398, N2377);
or OR3 (N2399, N2390, N1790, N1443);
xor XOR2 (N2400, N2399, N1887);
buf BUF1 (N2401, N2392);
and AND4 (N2402, N2385, N669, N750, N815);
not NOT1 (N2403, N2402);
not NOT1 (N2404, N2393);
xor XOR2 (N2405, N2401, N2090);
or OR4 (N2406, N2396, N1880, N1770, N2266);
buf BUF1 (N2407, N2384);
buf BUF1 (N2408, N2394);
not NOT1 (N2409, N2407);
nand NAND4 (N2410, N2400, N1030, N1082, N729);
or OR4 (N2411, N2398, N1665, N1240, N1266);
nor NOR3 (N2412, N2397, N1647, N942);
xor XOR2 (N2413, N2411, N1043);
buf BUF1 (N2414, N2403);
buf BUF1 (N2415, N2414);
xor XOR2 (N2416, N2413, N278);
nand NAND3 (N2417, N2409, N2414, N610);
nor NOR4 (N2418, N2410, N2355, N827, N1782);
xor XOR2 (N2419, N2404, N1675);
buf BUF1 (N2420, N2417);
nand NAND3 (N2421, N2418, N1536, N850);
xor XOR2 (N2422, N2420, N811);
not NOT1 (N2423, N2415);
or OR2 (N2424, N2412, N2190);
xor XOR2 (N2425, N2421, N1612);
and AND2 (N2426, N2405, N1018);
nand NAND3 (N2427, N2406, N421, N497);
and AND2 (N2428, N2426, N19);
nor NOR3 (N2429, N2408, N1121, N1798);
nand NAND2 (N2430, N2428, N667);
nand NAND3 (N2431, N2416, N449, N2068);
xor XOR2 (N2432, N2419, N2081);
nand NAND2 (N2433, N2432, N797);
and AND2 (N2434, N2431, N2197);
nor NOR2 (N2435, N2423, N1833);
and AND3 (N2436, N2435, N694, N1679);
xor XOR2 (N2437, N2424, N2331);
nor NOR4 (N2438, N2433, N2263, N963, N1057);
not NOT1 (N2439, N2437);
nand NAND2 (N2440, N2438, N935);
or OR3 (N2441, N2429, N2386, N1077);
and AND2 (N2442, N2427, N2293);
or OR2 (N2443, N2425, N895);
xor XOR2 (N2444, N2436, N1594);
nor NOR2 (N2445, N2422, N798);
buf BUF1 (N2446, N2440);
not NOT1 (N2447, N2444);
nand NAND2 (N2448, N2434, N1487);
nor NOR3 (N2449, N2354, N808, N1422);
xor XOR2 (N2450, N2430, N923);
or OR4 (N2451, N2447, N952, N1006, N1964);
nor NOR4 (N2452, N2445, N698, N2444, N1606);
xor XOR2 (N2453, N2449, N1188);
or OR4 (N2454, N2446, N1645, N1534, N632);
or OR2 (N2455, N2450, N1989);
not NOT1 (N2456, N2442);
nor NOR2 (N2457, N2441, N1661);
nor NOR4 (N2458, N2457, N1354, N2341, N2435);
nor NOR3 (N2459, N2456, N1649, N1893);
nor NOR3 (N2460, N2448, N705, N999);
nor NOR2 (N2461, N2455, N1524);
nor NOR4 (N2462, N2459, N745, N1161, N780);
nor NOR4 (N2463, N2460, N1418, N1431, N812);
not NOT1 (N2464, N2463);
or OR4 (N2465, N2458, N227, N471, N1829);
nand NAND4 (N2466, N2461, N1371, N1861, N588);
and AND3 (N2467, N2466, N24, N1562);
and AND3 (N2468, N2443, N1545, N793);
or OR2 (N2469, N2454, N1307);
buf BUF1 (N2470, N2452);
nor NOR3 (N2471, N2439, N541, N1258);
nand NAND2 (N2472, N2464, N1101);
and AND3 (N2473, N2472, N725, N872);
nand NAND2 (N2474, N2473, N1216);
xor XOR2 (N2475, N2467, N663);
not NOT1 (N2476, N2471);
nand NAND4 (N2477, N2475, N2365, N1401, N1166);
nand NAND4 (N2478, N2451, N2306, N1277, N1985);
and AND2 (N2479, N2469, N1081);
not NOT1 (N2480, N2479);
nor NOR2 (N2481, N2468, N883);
or OR3 (N2482, N2453, N99, N833);
and AND3 (N2483, N2481, N762, N2233);
nor NOR4 (N2484, N2478, N1303, N881, N1766);
or OR4 (N2485, N2465, N2453, N1413, N2298);
xor XOR2 (N2486, N2485, N409);
nand NAND4 (N2487, N2480, N1829, N1960, N1929);
nor NOR2 (N2488, N2486, N746);
nor NOR2 (N2489, N2487, N2436);
xor XOR2 (N2490, N2482, N2473);
not NOT1 (N2491, N2483);
nand NAND4 (N2492, N2474, N2286, N2340, N173);
not NOT1 (N2493, N2491);
not NOT1 (N2494, N2477);
nand NAND4 (N2495, N2476, N205, N999, N739);
and AND4 (N2496, N2493, N1890, N747, N2209);
not NOT1 (N2497, N2490);
buf BUF1 (N2498, N2496);
xor XOR2 (N2499, N2488, N1679);
or OR4 (N2500, N2470, N1556, N1137, N985);
xor XOR2 (N2501, N2494, N1288);
xor XOR2 (N2502, N2492, N132);
and AND3 (N2503, N2497, N1884, N1850);
nand NAND2 (N2504, N2498, N2308);
buf BUF1 (N2505, N2499);
or OR2 (N2506, N2484, N2397);
nand NAND3 (N2507, N2495, N1255, N1828);
xor XOR2 (N2508, N2501, N1392);
or OR2 (N2509, N2503, N2161);
and AND2 (N2510, N2500, N1250);
not NOT1 (N2511, N2506);
and AND3 (N2512, N2502, N2021, N2287);
xor XOR2 (N2513, N2512, N1669);
and AND2 (N2514, N2508, N664);
nand NAND3 (N2515, N2507, N1024, N1082);
nor NOR4 (N2516, N2489, N1026, N2306, N1155);
nor NOR2 (N2517, N2510, N544);
and AND3 (N2518, N2511, N370, N985);
or OR3 (N2519, N2505, N875, N2502);
and AND2 (N2520, N2509, N232);
not NOT1 (N2521, N2514);
not NOT1 (N2522, N2513);
buf BUF1 (N2523, N2462);
and AND4 (N2524, N2520, N417, N560, N1107);
xor XOR2 (N2525, N2523, N1937);
buf BUF1 (N2526, N2524);
not NOT1 (N2527, N2504);
and AND4 (N2528, N2515, N1125, N917, N675);
or OR4 (N2529, N2525, N2351, N574, N1533);
nor NOR4 (N2530, N2516, N1736, N2268, N2436);
and AND2 (N2531, N2517, N2006);
buf BUF1 (N2532, N2526);
buf BUF1 (N2533, N2531);
nand NAND4 (N2534, N2530, N729, N837, N1461);
buf BUF1 (N2535, N2518);
nor NOR3 (N2536, N2522, N228, N320);
not NOT1 (N2537, N2527);
nor NOR4 (N2538, N2528, N1914, N1430, N1395);
or OR4 (N2539, N2529, N947, N262, N949);
nor NOR2 (N2540, N2532, N431);
buf BUF1 (N2541, N2537);
nand NAND3 (N2542, N2535, N2373, N1608);
and AND4 (N2543, N2542, N1923, N778, N1129);
not NOT1 (N2544, N2521);
buf BUF1 (N2545, N2533);
xor XOR2 (N2546, N2536, N909);
and AND4 (N2547, N2543, N1756, N377, N1815);
or OR3 (N2548, N2538, N1818, N873);
buf BUF1 (N2549, N2541);
xor XOR2 (N2550, N2548, N34);
and AND4 (N2551, N2546, N789, N2289, N365);
xor XOR2 (N2552, N2519, N294);
not NOT1 (N2553, N2550);
nand NAND2 (N2554, N2534, N1670);
nor NOR2 (N2555, N2540, N1420);
nor NOR3 (N2556, N2549, N51, N2527);
nor NOR4 (N2557, N2553, N17, N2177, N1259);
or OR4 (N2558, N2555, N1949, N566, N217);
or OR4 (N2559, N2557, N1277, N1138, N2353);
or OR4 (N2560, N2539, N140, N1971, N2137);
buf BUF1 (N2561, N2558);
nand NAND3 (N2562, N2545, N2113, N915);
xor XOR2 (N2563, N2560, N1051);
not NOT1 (N2564, N2554);
or OR4 (N2565, N2552, N533, N1400, N1618);
buf BUF1 (N2566, N2562);
and AND4 (N2567, N2559, N1897, N1571, N1496);
nand NAND4 (N2568, N2563, N650, N1890, N630);
buf BUF1 (N2569, N2561);
not NOT1 (N2570, N2569);
nor NOR3 (N2571, N2566, N2081, N1839);
and AND2 (N2572, N2544, N2011);
nor NOR4 (N2573, N2570, N660, N1862, N434);
and AND2 (N2574, N2565, N2146);
nor NOR3 (N2575, N2574, N2273, N2430);
nor NOR3 (N2576, N2572, N1403, N1554);
or OR4 (N2577, N2556, N1883, N1713, N1647);
and AND2 (N2578, N2567, N2049);
and AND4 (N2579, N2575, N154, N2299, N1816);
xor XOR2 (N2580, N2547, N299);
or OR3 (N2581, N2551, N1626, N1978);
not NOT1 (N2582, N2571);
and AND3 (N2583, N2582, N647, N2535);
buf BUF1 (N2584, N2564);
or OR3 (N2585, N2577, N1340, N740);
buf BUF1 (N2586, N2579);
nand NAND3 (N2587, N2568, N2343, N1025);
not NOT1 (N2588, N2586);
or OR4 (N2589, N2581, N1604, N679, N105);
nand NAND4 (N2590, N2580, N7, N1345, N243);
nor NOR3 (N2591, N2576, N1989, N308);
nor NOR3 (N2592, N2578, N79, N1650);
buf BUF1 (N2593, N2589);
and AND4 (N2594, N2593, N322, N1783, N2149);
nor NOR2 (N2595, N2592, N311);
xor XOR2 (N2596, N2584, N299);
and AND4 (N2597, N2587, N2022, N1342, N70);
not NOT1 (N2598, N2597);
xor XOR2 (N2599, N2585, N557);
xor XOR2 (N2600, N2599, N1641);
not NOT1 (N2601, N2595);
not NOT1 (N2602, N2596);
not NOT1 (N2603, N2594);
not NOT1 (N2604, N2598);
and AND4 (N2605, N2602, N460, N972, N1345);
nand NAND3 (N2606, N2604, N1568, N195);
or OR3 (N2607, N2588, N1364, N1580);
not NOT1 (N2608, N2590);
xor XOR2 (N2609, N2608, N246);
xor XOR2 (N2610, N2609, N70);
nand NAND2 (N2611, N2601, N1306);
not NOT1 (N2612, N2606);
or OR2 (N2613, N2600, N2344);
and AND3 (N2614, N2613, N1044, N1331);
xor XOR2 (N2615, N2611, N2118);
buf BUF1 (N2616, N2583);
or OR4 (N2617, N2605, N1609, N853, N2520);
not NOT1 (N2618, N2615);
xor XOR2 (N2619, N2607, N1067);
xor XOR2 (N2620, N2612, N2242);
buf BUF1 (N2621, N2618);
not NOT1 (N2622, N2614);
nor NOR4 (N2623, N2619, N116, N920, N592);
buf BUF1 (N2624, N2591);
xor XOR2 (N2625, N2617, N835);
and AND3 (N2626, N2610, N1822, N1325);
nor NOR2 (N2627, N2620, N643);
not NOT1 (N2628, N2627);
or OR4 (N2629, N2625, N1333, N1830, N555);
xor XOR2 (N2630, N2626, N1744);
xor XOR2 (N2631, N2622, N2192);
or OR2 (N2632, N2573, N965);
nand NAND3 (N2633, N2616, N2325, N1805);
buf BUF1 (N2634, N2624);
or OR2 (N2635, N2633, N2094);
not NOT1 (N2636, N2634);
xor XOR2 (N2637, N2621, N1146);
not NOT1 (N2638, N2632);
not NOT1 (N2639, N2638);
and AND3 (N2640, N2639, N1414, N1880);
or OR3 (N2641, N2637, N199, N2112);
nor NOR4 (N2642, N2623, N213, N2569, N446);
or OR2 (N2643, N2629, N663);
xor XOR2 (N2644, N2636, N1842);
buf BUF1 (N2645, N2628);
and AND3 (N2646, N2631, N2450, N2560);
xor XOR2 (N2647, N2640, N1792);
xor XOR2 (N2648, N2647, N2430);
not NOT1 (N2649, N2643);
and AND3 (N2650, N2644, N2171, N2240);
xor XOR2 (N2651, N2641, N1947);
nand NAND3 (N2652, N2603, N287, N829);
or OR4 (N2653, N2642, N2333, N2321, N370);
xor XOR2 (N2654, N2649, N1709);
buf BUF1 (N2655, N2654);
not NOT1 (N2656, N2650);
buf BUF1 (N2657, N2645);
nor NOR2 (N2658, N2652, N44);
nand NAND4 (N2659, N2655, N174, N1824, N1581);
nand NAND3 (N2660, N2659, N1564, N280);
and AND3 (N2661, N2653, N2292, N215);
buf BUF1 (N2662, N2648);
and AND4 (N2663, N2662, N998, N426, N839);
not NOT1 (N2664, N2658);
and AND2 (N2665, N2656, N1422);
not NOT1 (N2666, N2664);
or OR2 (N2667, N2666, N687);
xor XOR2 (N2668, N2651, N2264);
xor XOR2 (N2669, N2646, N267);
buf BUF1 (N2670, N2669);
and AND3 (N2671, N2635, N219, N2482);
not NOT1 (N2672, N2663);
nand NAND2 (N2673, N2661, N1258);
buf BUF1 (N2674, N2670);
buf BUF1 (N2675, N2665);
buf BUF1 (N2676, N2675);
nand NAND4 (N2677, N2660, N2537, N1860, N1371);
nor NOR4 (N2678, N2674, N1927, N2430, N1983);
and AND2 (N2679, N2672, N1265);
and AND3 (N2680, N2678, N740, N2571);
not NOT1 (N2681, N2667);
or OR3 (N2682, N2673, N431, N744);
nor NOR3 (N2683, N2680, N1048, N87);
xor XOR2 (N2684, N2679, N1543);
not NOT1 (N2685, N2683);
not NOT1 (N2686, N2677);
nor NOR4 (N2687, N2671, N577, N698, N2386);
xor XOR2 (N2688, N2687, N2469);
buf BUF1 (N2689, N2630);
or OR2 (N2690, N2668, N2637);
nor NOR4 (N2691, N2682, N201, N1916, N652);
nand NAND3 (N2692, N2681, N1467, N171);
nor NOR4 (N2693, N2686, N1243, N204, N2203);
or OR4 (N2694, N2688, N1861, N1486, N2547);
nor NOR3 (N2695, N2692, N16, N1383);
and AND4 (N2696, N2695, N2570, N131, N203);
not NOT1 (N2697, N2691);
nor NOR4 (N2698, N2684, N1389, N912, N1880);
nand NAND3 (N2699, N2696, N1872, N991);
nand NAND4 (N2700, N2676, N2593, N1234, N1381);
nand NAND4 (N2701, N2700, N2005, N2457, N64);
not NOT1 (N2702, N2699);
xor XOR2 (N2703, N2694, N878);
nor NOR3 (N2704, N2657, N2321, N2270);
not NOT1 (N2705, N2701);
buf BUF1 (N2706, N2705);
and AND3 (N2707, N2704, N2492, N426);
nor NOR4 (N2708, N2690, N1975, N1437, N1948);
nand NAND4 (N2709, N2689, N69, N1897, N2513);
xor XOR2 (N2710, N2697, N304);
nor NOR4 (N2711, N2693, N2229, N2086, N2466);
nor NOR3 (N2712, N2685, N436, N638);
or OR3 (N2713, N2706, N2356, N2284);
buf BUF1 (N2714, N2710);
nand NAND3 (N2715, N2709, N631, N608);
or OR2 (N2716, N2707, N2603);
nand NAND4 (N2717, N2715, N1029, N1296, N941);
nand NAND4 (N2718, N2708, N836, N1330, N352);
and AND2 (N2719, N2711, N2569);
not NOT1 (N2720, N2714);
and AND2 (N2721, N2718, N2201);
buf BUF1 (N2722, N2702);
not NOT1 (N2723, N2720);
buf BUF1 (N2724, N2716);
not NOT1 (N2725, N2713);
not NOT1 (N2726, N2725);
nor NOR3 (N2727, N2717, N301, N1511);
xor XOR2 (N2728, N2721, N984);
buf BUF1 (N2729, N2719);
xor XOR2 (N2730, N2729, N1978);
xor XOR2 (N2731, N2728, N293);
xor XOR2 (N2732, N2698, N1532);
and AND4 (N2733, N2703, N203, N1262, N2370);
and AND3 (N2734, N2724, N1459, N359);
xor XOR2 (N2735, N2722, N2220);
nand NAND4 (N2736, N2731, N1464, N418, N1831);
and AND4 (N2737, N2733, N578, N597, N1385);
buf BUF1 (N2738, N2734);
not NOT1 (N2739, N2730);
nor NOR2 (N2740, N2723, N854);
buf BUF1 (N2741, N2740);
or OR3 (N2742, N2738, N1740, N1454);
nand NAND4 (N2743, N2736, N661, N819, N562);
or OR2 (N2744, N2737, N724);
nand NAND3 (N2745, N2726, N1185, N1814);
or OR3 (N2746, N2735, N1030, N2629);
nor NOR4 (N2747, N2745, N914, N1086, N1517);
buf BUF1 (N2748, N2747);
nand NAND2 (N2749, N2743, N337);
nor NOR2 (N2750, N2742, N1451);
not NOT1 (N2751, N2746);
or OR4 (N2752, N2727, N178, N1639, N1266);
and AND2 (N2753, N2750, N1620);
xor XOR2 (N2754, N2732, N532);
buf BUF1 (N2755, N2752);
and AND3 (N2756, N2748, N1789, N89);
nor NOR3 (N2757, N2751, N1363, N2535);
not NOT1 (N2758, N2741);
or OR4 (N2759, N2749, N185, N2231, N1291);
and AND3 (N2760, N2754, N2173, N2338);
nand NAND2 (N2761, N2759, N1916);
xor XOR2 (N2762, N2712, N272);
not NOT1 (N2763, N2762);
or OR4 (N2764, N2739, N643, N2413, N1629);
or OR3 (N2765, N2744, N568, N165);
buf BUF1 (N2766, N2753);
or OR3 (N2767, N2758, N1022, N1802);
and AND2 (N2768, N2763, N510);
and AND4 (N2769, N2760, N1286, N2571, N2195);
xor XOR2 (N2770, N2756, N1891);
not NOT1 (N2771, N2768);
nand NAND4 (N2772, N2769, N2089, N2702, N1437);
and AND4 (N2773, N2765, N2471, N2439, N1480);
and AND3 (N2774, N2766, N1354, N2539);
and AND2 (N2775, N2774, N770);
xor XOR2 (N2776, N2755, N2598);
and AND3 (N2777, N2776, N2219, N964);
xor XOR2 (N2778, N2761, N2670);
nand NAND2 (N2779, N2773, N2302);
and AND4 (N2780, N2778, N2709, N2610, N1068);
not NOT1 (N2781, N2770);
buf BUF1 (N2782, N2772);
nand NAND2 (N2783, N2757, N1499);
or OR3 (N2784, N2781, N1235, N1597);
or OR2 (N2785, N2771, N2521);
or OR4 (N2786, N2777, N1069, N2677, N263);
and AND3 (N2787, N2782, N1152, N180);
nor NOR2 (N2788, N2780, N2371);
nand NAND3 (N2789, N2783, N1003, N1560);
not NOT1 (N2790, N2788);
or OR2 (N2791, N2764, N2292);
nor NOR3 (N2792, N2767, N2333, N2691);
xor XOR2 (N2793, N2791, N862);
nor NOR2 (N2794, N2775, N658);
nand NAND2 (N2795, N2784, N1325);
xor XOR2 (N2796, N2789, N1622);
nand NAND3 (N2797, N2779, N2100, N946);
xor XOR2 (N2798, N2796, N1895);
or OR4 (N2799, N2787, N1815, N765, N224);
nor NOR2 (N2800, N2785, N1089);
or OR2 (N2801, N2798, N2096);
not NOT1 (N2802, N2801);
not NOT1 (N2803, N2795);
or OR4 (N2804, N2802, N1519, N1960, N581);
buf BUF1 (N2805, N2794);
nor NOR3 (N2806, N2804, N2507, N1628);
nand NAND4 (N2807, N2786, N1300, N770, N1112);
not NOT1 (N2808, N2793);
xor XOR2 (N2809, N2797, N1176);
xor XOR2 (N2810, N2803, N1682);
buf BUF1 (N2811, N2790);
buf BUF1 (N2812, N2799);
and AND3 (N2813, N2800, N1613, N113);
xor XOR2 (N2814, N2805, N260);
not NOT1 (N2815, N2806);
nor NOR4 (N2816, N2807, N2753, N2600, N374);
buf BUF1 (N2817, N2813);
nand NAND3 (N2818, N2815, N2761, N240);
nor NOR3 (N2819, N2816, N2353, N121);
nand NAND3 (N2820, N2819, N2005, N169);
xor XOR2 (N2821, N2814, N1440);
nand NAND4 (N2822, N2808, N2519, N1293, N336);
nand NAND3 (N2823, N2822, N648, N388);
nor NOR2 (N2824, N2792, N2377);
and AND4 (N2825, N2811, N139, N1155, N927);
buf BUF1 (N2826, N2821);
xor XOR2 (N2827, N2820, N1675);
or OR4 (N2828, N2823, N1373, N1166, N1015);
nand NAND4 (N2829, N2825, N665, N2177, N2069);
and AND2 (N2830, N2810, N393);
or OR3 (N2831, N2827, N2126, N1551);
xor XOR2 (N2832, N2812, N2570);
or OR4 (N2833, N2831, N1592, N1942, N2579);
and AND2 (N2834, N2809, N965);
or OR4 (N2835, N2818, N1086, N2085, N678);
nand NAND2 (N2836, N2817, N2502);
nor NOR4 (N2837, N2836, N83, N175, N61);
xor XOR2 (N2838, N2830, N939);
xor XOR2 (N2839, N2838, N2528);
not NOT1 (N2840, N2824);
not NOT1 (N2841, N2832);
nand NAND3 (N2842, N2828, N31, N1652);
buf BUF1 (N2843, N2834);
buf BUF1 (N2844, N2833);
nor NOR2 (N2845, N2835, N1658);
buf BUF1 (N2846, N2826);
and AND3 (N2847, N2844, N2579, N689);
not NOT1 (N2848, N2829);
or OR3 (N2849, N2840, N754, N892);
not NOT1 (N2850, N2849);
nand NAND4 (N2851, N2846, N1836, N591, N1346);
or OR4 (N2852, N2842, N2016, N2349, N789);
buf BUF1 (N2853, N2851);
not NOT1 (N2854, N2839);
nand NAND2 (N2855, N2847, N1803);
and AND3 (N2856, N2852, N2538, N2840);
nand NAND4 (N2857, N2856, N2188, N2499, N1012);
and AND4 (N2858, N2845, N1711, N852, N1924);
buf BUF1 (N2859, N2837);
buf BUF1 (N2860, N2855);
buf BUF1 (N2861, N2860);
or OR3 (N2862, N2854, N2209, N2367);
and AND3 (N2863, N2862, N1674, N2657);
nor NOR2 (N2864, N2853, N2357);
or OR3 (N2865, N2857, N1991, N2371);
and AND3 (N2866, N2848, N2696, N2171);
nand NAND4 (N2867, N2866, N838, N267, N1766);
and AND3 (N2868, N2861, N1498, N605);
not NOT1 (N2869, N2864);
not NOT1 (N2870, N2843);
and AND2 (N2871, N2869, N2437);
not NOT1 (N2872, N2865);
nand NAND4 (N2873, N2872, N2685, N2662, N2417);
buf BUF1 (N2874, N2873);
nand NAND4 (N2875, N2874, N2653, N469, N2436);
not NOT1 (N2876, N2870);
not NOT1 (N2877, N2859);
not NOT1 (N2878, N2867);
and AND4 (N2879, N2878, N1293, N911, N931);
buf BUF1 (N2880, N2876);
xor XOR2 (N2881, N2879, N571);
buf BUF1 (N2882, N2881);
not NOT1 (N2883, N2882);
buf BUF1 (N2884, N2841);
nand NAND4 (N2885, N2871, N105, N2308, N753);
or OR2 (N2886, N2868, N881);
nor NOR3 (N2887, N2877, N517, N2355);
and AND3 (N2888, N2886, N309, N382);
not NOT1 (N2889, N2884);
and AND3 (N2890, N2880, N2877, N1513);
nor NOR2 (N2891, N2887, N491);
or OR4 (N2892, N2885, N795, N84, N2792);
xor XOR2 (N2893, N2889, N171);
buf BUF1 (N2894, N2888);
nor NOR3 (N2895, N2892, N1866, N346);
nand NAND4 (N2896, N2895, N549, N2210, N2575);
xor XOR2 (N2897, N2893, N2247);
buf BUF1 (N2898, N2858);
not NOT1 (N2899, N2850);
nor NOR4 (N2900, N2894, N522, N1083, N2156);
nor NOR2 (N2901, N2897, N1376);
not NOT1 (N2902, N2890);
and AND4 (N2903, N2901, N2767, N1456, N393);
nand NAND4 (N2904, N2902, N1205, N1581, N1986);
nand NAND3 (N2905, N2903, N2610, N1410);
and AND3 (N2906, N2883, N2425, N483);
xor XOR2 (N2907, N2896, N1855);
buf BUF1 (N2908, N2898);
or OR4 (N2909, N2875, N614, N1598, N2619);
or OR2 (N2910, N2900, N1790);
buf BUF1 (N2911, N2907);
or OR2 (N2912, N2863, N1170);
not NOT1 (N2913, N2909);
or OR3 (N2914, N2904, N1712, N1753);
not NOT1 (N2915, N2891);
buf BUF1 (N2916, N2914);
xor XOR2 (N2917, N2911, N1508);
buf BUF1 (N2918, N2912);
nor NOR4 (N2919, N2913, N1983, N886, N1060);
nor NOR2 (N2920, N2917, N1620);
buf BUF1 (N2921, N2919);
nor NOR3 (N2922, N2920, N2106, N2624);
not NOT1 (N2923, N2908);
xor XOR2 (N2924, N2918, N1223);
and AND2 (N2925, N2923, N349);
xor XOR2 (N2926, N2924, N990);
nand NAND3 (N2927, N2921, N738, N2682);
not NOT1 (N2928, N2927);
buf BUF1 (N2929, N2905);
not NOT1 (N2930, N2899);
xor XOR2 (N2931, N2906, N108);
nor NOR4 (N2932, N2915, N1578, N42, N787);
not NOT1 (N2933, N2928);
buf BUF1 (N2934, N2926);
nor NOR4 (N2935, N2922, N1792, N2761, N1141);
and AND2 (N2936, N2930, N513);
or OR4 (N2937, N2925, N2487, N916, N1050);
nor NOR3 (N2938, N2935, N747, N1890);
or OR3 (N2939, N2936, N2403, N105);
not NOT1 (N2940, N2934);
and AND2 (N2941, N2938, N571);
buf BUF1 (N2942, N2933);
or OR2 (N2943, N2910, N1381);
and AND4 (N2944, N2943, N1193, N2888, N1);
not NOT1 (N2945, N2942);
buf BUF1 (N2946, N2940);
not NOT1 (N2947, N2944);
nand NAND4 (N2948, N2939, N859, N690, N2223);
xor XOR2 (N2949, N2932, N2400);
xor XOR2 (N2950, N2931, N28);
and AND3 (N2951, N2947, N942, N2122);
and AND4 (N2952, N2950, N1442, N1191, N481);
nand NAND4 (N2953, N2945, N977, N1189, N2220);
not NOT1 (N2954, N2949);
xor XOR2 (N2955, N2941, N1983);
not NOT1 (N2956, N2937);
or OR2 (N2957, N2956, N783);
xor XOR2 (N2958, N2951, N842);
not NOT1 (N2959, N2952);
nor NOR4 (N2960, N2955, N2598, N881, N1728);
xor XOR2 (N2961, N2957, N2434);
buf BUF1 (N2962, N2958);
or OR4 (N2963, N2962, N593, N1232, N2413);
buf BUF1 (N2964, N2954);
or OR4 (N2965, N2953, N2324, N756, N2067);
nand NAND2 (N2966, N2929, N1263);
nor NOR3 (N2967, N2959, N1802, N2537);
nand NAND4 (N2968, N2964, N695, N1197, N1380);
nand NAND4 (N2969, N2967, N198, N234, N27);
xor XOR2 (N2970, N2946, N1574);
nor NOR4 (N2971, N2966, N2091, N451, N239);
buf BUF1 (N2972, N2971);
and AND4 (N2973, N2960, N2406, N313, N2964);
or OR2 (N2974, N2963, N2548);
nand NAND3 (N2975, N2916, N1149, N2202);
nor NOR4 (N2976, N2973, N2204, N1476, N215);
nand NAND4 (N2977, N2968, N2812, N1377, N1497);
and AND4 (N2978, N2948, N998, N973, N645);
not NOT1 (N2979, N2970);
xor XOR2 (N2980, N2961, N2914);
or OR3 (N2981, N2965, N1482, N393);
xor XOR2 (N2982, N2972, N1142);
xor XOR2 (N2983, N2974, N402);
xor XOR2 (N2984, N2979, N1178);
and AND4 (N2985, N2978, N440, N121, N2276);
xor XOR2 (N2986, N2976, N2533);
buf BUF1 (N2987, N2982);
or OR2 (N2988, N2987, N995);
xor XOR2 (N2989, N2986, N387);
nand NAND4 (N2990, N2977, N1277, N1084, N1844);
not NOT1 (N2991, N2984);
nand NAND2 (N2992, N2975, N257);
buf BUF1 (N2993, N2981);
nor NOR2 (N2994, N2993, N599);
and AND3 (N2995, N2983, N689, N1883);
nor NOR2 (N2996, N2990, N2263);
and AND4 (N2997, N2988, N313, N568, N2961);
nor NOR2 (N2998, N2980, N496);
buf BUF1 (N2999, N2969);
nand NAND3 (N3000, N2989, N1716, N1300);
nor NOR4 (N3001, N2997, N1516, N1241, N545);
not NOT1 (N3002, N2991);
nand NAND4 (N3003, N2998, N1598, N879, N2483);
and AND2 (N3004, N2994, N2289);
nand NAND2 (N3005, N3002, N1374);
nor NOR3 (N3006, N2996, N2721, N2933);
nor NOR3 (N3007, N3004, N1940, N1437);
nand NAND4 (N3008, N3000, N396, N368, N1671);
buf BUF1 (N3009, N2995);
and AND2 (N3010, N3001, N1414);
nor NOR4 (N3011, N3008, N2231, N765, N1548);
or OR3 (N3012, N3010, N2580, N135);
buf BUF1 (N3013, N3003);
or OR3 (N3014, N3013, N2693, N1902);
xor XOR2 (N3015, N2999, N356);
nand NAND4 (N3016, N3014, N2385, N2727, N1453);
nor NOR4 (N3017, N3006, N2453, N492, N2157);
not NOT1 (N3018, N2992);
nor NOR4 (N3019, N3005, N8, N1560, N2847);
or OR2 (N3020, N3019, N1560);
nand NAND4 (N3021, N3016, N185, N1757, N2858);
xor XOR2 (N3022, N3012, N1671);
nand NAND2 (N3023, N3007, N2920);
nor NOR2 (N3024, N3021, N1642);
not NOT1 (N3025, N3017);
not NOT1 (N3026, N3011);
and AND3 (N3027, N3015, N1810, N519);
not NOT1 (N3028, N3025);
buf BUF1 (N3029, N3009);
not NOT1 (N3030, N3027);
not NOT1 (N3031, N3029);
buf BUF1 (N3032, N3030);
nor NOR2 (N3033, N3032, N2976);
and AND4 (N3034, N3031, N1298, N2984, N553);
or OR2 (N3035, N2985, N1782);
or OR4 (N3036, N3024, N2056, N639, N246);
or OR3 (N3037, N3023, N1966, N1274);
or OR2 (N3038, N3035, N2116);
buf BUF1 (N3039, N3026);
buf BUF1 (N3040, N3037);
not NOT1 (N3041, N3022);
or OR3 (N3042, N3040, N2919, N376);
xor XOR2 (N3043, N3018, N1607);
and AND4 (N3044, N3034, N440, N1320, N2234);
nand NAND4 (N3045, N3043, N2339, N915, N1927);
nand NAND2 (N3046, N3038, N2007);
buf BUF1 (N3047, N3039);
nand NAND2 (N3048, N3042, N2868);
or OR4 (N3049, N3044, N2661, N981, N542);
nor NOR4 (N3050, N3020, N1867, N1642, N502);
and AND4 (N3051, N3049, N1694, N2524, N67);
nor NOR4 (N3052, N3048, N32, N2453, N1355);
and AND3 (N3053, N3033, N1006, N831);
xor XOR2 (N3054, N3050, N124);
buf BUF1 (N3055, N3046);
or OR4 (N3056, N3052, N725, N166, N1368);
or OR2 (N3057, N3041, N2931);
not NOT1 (N3058, N3057);
not NOT1 (N3059, N3051);
nand NAND3 (N3060, N3045, N615, N1214);
nor NOR3 (N3061, N3058, N845, N1320);
xor XOR2 (N3062, N3056, N1817);
not NOT1 (N3063, N3054);
nand NAND3 (N3064, N3060, N1817, N2372);
and AND4 (N3065, N3055, N1345, N2342, N1757);
buf BUF1 (N3066, N3062);
buf BUF1 (N3067, N3063);
nand NAND2 (N3068, N3047, N2278);
not NOT1 (N3069, N3059);
buf BUF1 (N3070, N3064);
buf BUF1 (N3071, N3070);
buf BUF1 (N3072, N3066);
xor XOR2 (N3073, N3071, N1570);
nor NOR3 (N3074, N3065, N2038, N1018);
and AND3 (N3075, N3036, N1345, N1872);
xor XOR2 (N3076, N3068, N2410);
and AND2 (N3077, N3069, N2633);
nand NAND2 (N3078, N3073, N2367);
nor NOR3 (N3079, N3075, N2889, N787);
nand NAND4 (N3080, N3074, N1796, N2850, N1815);
not NOT1 (N3081, N3078);
buf BUF1 (N3082, N3067);
buf BUF1 (N3083, N3082);
or OR3 (N3084, N3053, N705, N2848);
and AND3 (N3085, N3080, N1696, N227);
nor NOR4 (N3086, N3072, N3057, N1698, N2907);
or OR2 (N3087, N3028, N2196);
and AND4 (N3088, N3076, N635, N202, N1191);
buf BUF1 (N3089, N3088);
not NOT1 (N3090, N3079);
nor NOR3 (N3091, N3084, N1362, N991);
nand NAND4 (N3092, N3086, N156, N1055, N1053);
nand NAND3 (N3093, N3077, N1403, N935);
xor XOR2 (N3094, N3083, N406);
and AND2 (N3095, N3092, N2897);
nand NAND2 (N3096, N3094, N2932);
nor NOR4 (N3097, N3081, N2797, N2322, N1770);
or OR4 (N3098, N3061, N2527, N2465, N1922);
nor NOR3 (N3099, N3090, N1879, N942);
xor XOR2 (N3100, N3093, N2582);
nor NOR2 (N3101, N3087, N2052);
buf BUF1 (N3102, N3095);
or OR3 (N3103, N3102, N2666, N2681);
nor NOR4 (N3104, N3100, N907, N2188, N1761);
and AND3 (N3105, N3096, N1019, N721);
not NOT1 (N3106, N3099);
nand NAND4 (N3107, N3103, N200, N1158, N351);
and AND2 (N3108, N3101, N2029);
not NOT1 (N3109, N3106);
nand NAND4 (N3110, N3098, N951, N39, N2794);
nor NOR2 (N3111, N3091, N719);
nor NOR4 (N3112, N3104, N1341, N1929, N2268);
buf BUF1 (N3113, N3107);
not NOT1 (N3114, N3111);
xor XOR2 (N3115, N3089, N2001);
xor XOR2 (N3116, N3113, N1967);
buf BUF1 (N3117, N3108);
nor NOR2 (N3118, N3085, N539);
not NOT1 (N3119, N3118);
xor XOR2 (N3120, N3112, N1368);
not NOT1 (N3121, N3110);
nor NOR3 (N3122, N3105, N724, N271);
nand NAND4 (N3123, N3115, N2402, N661, N835);
nand NAND2 (N3124, N3120, N1230);
nand NAND2 (N3125, N3109, N21);
buf BUF1 (N3126, N3097);
or OR4 (N3127, N3117, N662, N2773, N232);
xor XOR2 (N3128, N3127, N2667);
buf BUF1 (N3129, N3119);
not NOT1 (N3130, N3125);
nor NOR3 (N3131, N3130, N2305, N980);
nand NAND4 (N3132, N3131, N1960, N2760, N212);
buf BUF1 (N3133, N3123);
and AND3 (N3134, N3129, N304, N574);
or OR4 (N3135, N3124, N2454, N967, N2804);
or OR4 (N3136, N3134, N2160, N2357, N1729);
buf BUF1 (N3137, N3126);
nand NAND4 (N3138, N3136, N2562, N708, N531);
not NOT1 (N3139, N3135);
nand NAND3 (N3140, N3138, N1877, N1145);
buf BUF1 (N3141, N3122);
not NOT1 (N3142, N3139);
nand NAND3 (N3143, N3121, N1055, N2391);
buf BUF1 (N3144, N3132);
buf BUF1 (N3145, N3137);
not NOT1 (N3146, N3143);
nand NAND2 (N3147, N3128, N2653);
not NOT1 (N3148, N3147);
buf BUF1 (N3149, N3144);
xor XOR2 (N3150, N3148, N1104);
nand NAND4 (N3151, N3141, N2525, N2618, N503);
not NOT1 (N3152, N3150);
or OR2 (N3153, N3133, N2643);
nand NAND2 (N3154, N3145, N1899);
and AND2 (N3155, N3152, N1930);
and AND2 (N3156, N3114, N1601);
nand NAND3 (N3157, N3155, N753, N1682);
not NOT1 (N3158, N3116);
nand NAND2 (N3159, N3151, N547);
nor NOR4 (N3160, N3157, N682, N2341, N218);
or OR3 (N3161, N3158, N958, N1885);
nor NOR4 (N3162, N3154, N38, N2961, N3030);
or OR2 (N3163, N3140, N1444);
not NOT1 (N3164, N3149);
nor NOR3 (N3165, N3142, N2622, N2402);
buf BUF1 (N3166, N3160);
not NOT1 (N3167, N3159);
or OR4 (N3168, N3165, N2291, N2255, N2680);
buf BUF1 (N3169, N3168);
or OR2 (N3170, N3163, N1450);
not NOT1 (N3171, N3161);
and AND2 (N3172, N3171, N1440);
nand NAND3 (N3173, N3153, N2575, N1226);
nand NAND3 (N3174, N3146, N2918, N2217);
xor XOR2 (N3175, N3173, N726);
nand NAND2 (N3176, N3174, N2110);
and AND2 (N3177, N3169, N2434);
xor XOR2 (N3178, N3166, N237);
buf BUF1 (N3179, N3170);
and AND2 (N3180, N3175, N672);
buf BUF1 (N3181, N3167);
or OR2 (N3182, N3156, N3013);
xor XOR2 (N3183, N3172, N510);
not NOT1 (N3184, N3183);
nand NAND3 (N3185, N3181, N1441, N1583);
buf BUF1 (N3186, N3178);
nand NAND4 (N3187, N3182, N2050, N185, N311);
and AND3 (N3188, N3187, N3132, N723);
buf BUF1 (N3189, N3186);
buf BUF1 (N3190, N3184);
and AND4 (N3191, N3162, N2472, N2292, N2090);
or OR2 (N3192, N3188, N970);
nand NAND4 (N3193, N3164, N35, N1467, N1466);
buf BUF1 (N3194, N3189);
xor XOR2 (N3195, N3191, N1102);
buf BUF1 (N3196, N3177);
not NOT1 (N3197, N3196);
nor NOR4 (N3198, N3192, N2975, N167, N2326);
not NOT1 (N3199, N3179);
buf BUF1 (N3200, N3198);
nor NOR4 (N3201, N3190, N2297, N646, N2563);
buf BUF1 (N3202, N3180);
nand NAND2 (N3203, N3176, N360);
nor NOR4 (N3204, N3201, N1887, N1205, N1483);
and AND2 (N3205, N3185, N3016);
and AND3 (N3206, N3195, N2562, N574);
or OR4 (N3207, N3203, N1215, N2357, N2915);
or OR2 (N3208, N3202, N445);
not NOT1 (N3209, N3208);
not NOT1 (N3210, N3209);
not NOT1 (N3211, N3193);
and AND4 (N3212, N3194, N2697, N2654, N1523);
not NOT1 (N3213, N3211);
nand NAND2 (N3214, N3200, N1640);
and AND2 (N3215, N3214, N2650);
nand NAND3 (N3216, N3210, N435, N63);
or OR3 (N3217, N3197, N3046, N3065);
nand NAND4 (N3218, N3217, N1505, N972, N1187);
or OR2 (N3219, N3213, N2672);
not NOT1 (N3220, N3204);
buf BUF1 (N3221, N3218);
nor NOR2 (N3222, N3207, N86);
xor XOR2 (N3223, N3215, N1856);
xor XOR2 (N3224, N3221, N603);
and AND4 (N3225, N3223, N2532, N2775, N2537);
nand NAND2 (N3226, N3199, N582);
or OR4 (N3227, N3212, N1810, N1377, N2657);
not NOT1 (N3228, N3205);
nor NOR3 (N3229, N3219, N3026, N2714);
and AND3 (N3230, N3222, N2654, N1093);
buf BUF1 (N3231, N3216);
or OR4 (N3232, N3226, N1609, N308, N2563);
not NOT1 (N3233, N3232);
nor NOR4 (N3234, N3229, N1461, N1221, N2335);
nor NOR3 (N3235, N3231, N735, N1951);
nand NAND3 (N3236, N3234, N939, N1750);
and AND4 (N3237, N3225, N961, N1482, N1833);
or OR3 (N3238, N3206, N2219, N2243);
xor XOR2 (N3239, N3228, N1447);
not NOT1 (N3240, N3224);
or OR4 (N3241, N3227, N2524, N1619, N2571);
xor XOR2 (N3242, N3240, N1541);
or OR2 (N3243, N3236, N1983);
nor NOR3 (N3244, N3241, N10, N1988);
and AND4 (N3245, N3238, N560, N1285, N749);
or OR3 (N3246, N3242, N732, N2231);
xor XOR2 (N3247, N3239, N1379);
buf BUF1 (N3248, N3237);
not NOT1 (N3249, N3248);
nand NAND2 (N3250, N3230, N1734);
nand NAND2 (N3251, N3233, N1679);
or OR3 (N3252, N3243, N2659, N1192);
not NOT1 (N3253, N3235);
buf BUF1 (N3254, N3250);
nand NAND3 (N3255, N3220, N2806, N805);
nor NOR4 (N3256, N3252, N1311, N2246, N602);
buf BUF1 (N3257, N3253);
nor NOR2 (N3258, N3247, N3199);
or OR4 (N3259, N3246, N2816, N1038, N2052);
nor NOR2 (N3260, N3254, N2872);
buf BUF1 (N3261, N3260);
nand NAND2 (N3262, N3244, N2881);
not NOT1 (N3263, N3261);
not NOT1 (N3264, N3258);
xor XOR2 (N3265, N3255, N1450);
nand NAND3 (N3266, N3264, N3013, N1845);
nor NOR4 (N3267, N3262, N1835, N986, N449);
nand NAND3 (N3268, N3265, N675, N1566);
buf BUF1 (N3269, N3251);
nand NAND3 (N3270, N3268, N2456, N503);
buf BUF1 (N3271, N3266);
nand NAND4 (N3272, N3263, N3100, N2327, N442);
buf BUF1 (N3273, N3256);
and AND4 (N3274, N3271, N701, N400, N960);
nor NOR3 (N3275, N3273, N523, N1944);
nand NAND2 (N3276, N3274, N2331);
xor XOR2 (N3277, N3269, N2996);
or OR2 (N3278, N3257, N2901);
buf BUF1 (N3279, N3272);
nand NAND3 (N3280, N3245, N257, N1545);
xor XOR2 (N3281, N3270, N676);
xor XOR2 (N3282, N3280, N2553);
xor XOR2 (N3283, N3282, N3241);
buf BUF1 (N3284, N3277);
or OR4 (N3285, N3283, N3121, N547, N2528);
nand NAND2 (N3286, N3276, N1164);
nand NAND2 (N3287, N3279, N1790);
and AND4 (N3288, N3286, N2103, N1312, N1904);
buf BUF1 (N3289, N3288);
nand NAND2 (N3290, N3267, N1849);
not NOT1 (N3291, N3284);
xor XOR2 (N3292, N3289, N279);
buf BUF1 (N3293, N3278);
nor NOR3 (N3294, N3259, N2388, N3151);
or OR3 (N3295, N3292, N2821, N728);
not NOT1 (N3296, N3281);
not NOT1 (N3297, N3296);
nor NOR4 (N3298, N3295, N2729, N1842, N2982);
nand NAND3 (N3299, N3297, N1230, N1330);
or OR4 (N3300, N3299, N243, N2637, N405);
and AND2 (N3301, N3293, N1750);
nand NAND4 (N3302, N3294, N2241, N292, N2591);
nor NOR3 (N3303, N3301, N2768, N936);
or OR2 (N3304, N3287, N3115);
xor XOR2 (N3305, N3249, N1370);
and AND4 (N3306, N3304, N622, N2509, N1590);
or OR4 (N3307, N3302, N1587, N1387, N1453);
and AND3 (N3308, N3291, N565, N259);
xor XOR2 (N3309, N3275, N360);
buf BUF1 (N3310, N3306);
not NOT1 (N3311, N3310);
nor NOR2 (N3312, N3285, N2186);
and AND3 (N3313, N3308, N1251, N2677);
nand NAND4 (N3314, N3305, N2087, N2134, N2916);
buf BUF1 (N3315, N3309);
nor NOR3 (N3316, N3307, N1200, N1726);
and AND2 (N3317, N3303, N2232);
and AND2 (N3318, N3314, N1250);
buf BUF1 (N3319, N3312);
nand NAND3 (N3320, N3315, N3260, N1738);
or OR2 (N3321, N3319, N2112);
buf BUF1 (N3322, N3298);
and AND4 (N3323, N3321, N42, N2353, N630);
buf BUF1 (N3324, N3313);
xor XOR2 (N3325, N3322, N2567);
nor NOR3 (N3326, N3311, N2458, N335);
not NOT1 (N3327, N3324);
xor XOR2 (N3328, N3325, N973);
nand NAND2 (N3329, N3318, N2995);
and AND4 (N3330, N3327, N2906, N966, N2979);
buf BUF1 (N3331, N3317);
nand NAND2 (N3332, N3290, N2262);
not NOT1 (N3333, N3332);
or OR4 (N3334, N3329, N3140, N149, N1541);
nor NOR2 (N3335, N3323, N2839);
and AND2 (N3336, N3335, N309);
buf BUF1 (N3337, N3333);
nand NAND2 (N3338, N3331, N1598);
buf BUF1 (N3339, N3336);
buf BUF1 (N3340, N3339);
buf BUF1 (N3341, N3340);
buf BUF1 (N3342, N3330);
xor XOR2 (N3343, N3337, N1335);
nand NAND4 (N3344, N3300, N1975, N256, N1208);
or OR4 (N3345, N3344, N361, N746, N373);
nand NAND3 (N3346, N3320, N2749, N997);
and AND2 (N3347, N3334, N2812);
not NOT1 (N3348, N3338);
buf BUF1 (N3349, N3345);
nor NOR2 (N3350, N3346, N3133);
and AND4 (N3351, N3348, N649, N1942, N145);
nor NOR3 (N3352, N3350, N172, N736);
not NOT1 (N3353, N3316);
or OR3 (N3354, N3328, N1109, N2311);
not NOT1 (N3355, N3347);
buf BUF1 (N3356, N3351);
not NOT1 (N3357, N3342);
nand NAND2 (N3358, N3353, N2404);
nand NAND3 (N3359, N3358, N382, N1069);
and AND4 (N3360, N3341, N3352, N1260, N3107);
nor NOR4 (N3361, N1211, N3330, N3216, N2990);
not NOT1 (N3362, N3355);
buf BUF1 (N3363, N3354);
buf BUF1 (N3364, N3360);
or OR4 (N3365, N3364, N2085, N2921, N2297);
nand NAND4 (N3366, N3362, N1944, N545, N2912);
not NOT1 (N3367, N3366);
nor NOR4 (N3368, N3343, N2983, N2845, N3331);
buf BUF1 (N3369, N3357);
and AND4 (N3370, N3326, N831, N2431, N574);
buf BUF1 (N3371, N3349);
nand NAND3 (N3372, N3368, N784, N3290);
buf BUF1 (N3373, N3372);
nand NAND2 (N3374, N3363, N2230);
xor XOR2 (N3375, N3369, N79);
or OR3 (N3376, N3374, N1733, N3299);
xor XOR2 (N3377, N3370, N1283);
not NOT1 (N3378, N3367);
not NOT1 (N3379, N3371);
nor NOR2 (N3380, N3373, N872);
and AND2 (N3381, N3376, N2975);
buf BUF1 (N3382, N3375);
or OR4 (N3383, N3377, N2280, N2937, N1935);
buf BUF1 (N3384, N3378);
xor XOR2 (N3385, N3379, N1197);
or OR3 (N3386, N3384, N2188, N1501);
xor XOR2 (N3387, N3381, N1653);
buf BUF1 (N3388, N3386);
or OR4 (N3389, N3387, N945, N288, N1649);
buf BUF1 (N3390, N3388);
buf BUF1 (N3391, N3385);
nand NAND3 (N3392, N3365, N1981, N2669);
xor XOR2 (N3393, N3380, N1428);
buf BUF1 (N3394, N3356);
nor NOR3 (N3395, N3361, N1933, N2880);
xor XOR2 (N3396, N3389, N1640);
not NOT1 (N3397, N3390);
xor XOR2 (N3398, N3397, N3096);
nor NOR4 (N3399, N3392, N11, N1540, N3214);
or OR2 (N3400, N3399, N2418);
nor NOR2 (N3401, N3398, N3123);
buf BUF1 (N3402, N3359);
or OR2 (N3403, N3396, N1610);
not NOT1 (N3404, N3393);
nor NOR3 (N3405, N3402, N1942, N3067);
buf BUF1 (N3406, N3394);
nand NAND4 (N3407, N3404, N3053, N1563, N866);
not NOT1 (N3408, N3400);
and AND3 (N3409, N3407, N3161, N1968);
nor NOR3 (N3410, N3408, N51, N1099);
buf BUF1 (N3411, N3410);
nand NAND4 (N3412, N3391, N1784, N2504, N2426);
buf BUF1 (N3413, N3406);
nor NOR3 (N3414, N3409, N1017, N2254);
xor XOR2 (N3415, N3382, N710);
or OR2 (N3416, N3413, N2896);
and AND3 (N3417, N3411, N1324, N1681);
nand NAND4 (N3418, N3405, N3219, N440, N239);
xor XOR2 (N3419, N3414, N1732);
and AND3 (N3420, N3418, N2962, N3132);
and AND4 (N3421, N3416, N1594, N1094, N798);
buf BUF1 (N3422, N3415);
nor NOR2 (N3423, N3420, N2651);
and AND2 (N3424, N3422, N1675);
or OR3 (N3425, N3401, N3133, N3277);
or OR2 (N3426, N3383, N1226);
buf BUF1 (N3427, N3419);
not NOT1 (N3428, N3395);
or OR2 (N3429, N3426, N516);
buf BUF1 (N3430, N3424);
not NOT1 (N3431, N3430);
xor XOR2 (N3432, N3428, N1769);
xor XOR2 (N3433, N3423, N595);
buf BUF1 (N3434, N3425);
xor XOR2 (N3435, N3431, N1481);
nand NAND2 (N3436, N3435, N2333);
and AND2 (N3437, N3436, N671);
nor NOR2 (N3438, N3417, N2130);
xor XOR2 (N3439, N3434, N1379);
nand NAND3 (N3440, N3421, N2622, N91);
or OR2 (N3441, N3440, N2333);
nor NOR2 (N3442, N3439, N2666);
not NOT1 (N3443, N3441);
or OR4 (N3444, N3403, N92, N792, N2883);
nor NOR2 (N3445, N3444, N1822);
buf BUF1 (N3446, N3432);
or OR3 (N3447, N3429, N3254, N2851);
buf BUF1 (N3448, N3442);
not NOT1 (N3449, N3412);
nand NAND3 (N3450, N3448, N3077, N3088);
and AND2 (N3451, N3446, N2222);
buf BUF1 (N3452, N3449);
nor NOR2 (N3453, N3450, N4);
not NOT1 (N3454, N3453);
and AND3 (N3455, N3447, N2021, N3337);
xor XOR2 (N3456, N3443, N453);
nand NAND3 (N3457, N3433, N2252, N1721);
not NOT1 (N3458, N3452);
xor XOR2 (N3459, N3437, N67);
or OR3 (N3460, N3459, N675, N731);
xor XOR2 (N3461, N3445, N2054);
or OR4 (N3462, N3456, N2889, N3456, N2404);
or OR3 (N3463, N3451, N1965, N1149);
nor NOR4 (N3464, N3458, N3296, N871, N1661);
xor XOR2 (N3465, N3462, N3025);
or OR3 (N3466, N3454, N367, N1732);
xor XOR2 (N3467, N3466, N1125);
nand NAND3 (N3468, N3457, N3055, N3311);
xor XOR2 (N3469, N3465, N2069);
xor XOR2 (N3470, N3460, N1614);
xor XOR2 (N3471, N3470, N300);
nand NAND3 (N3472, N3461, N1571, N80);
nand NAND4 (N3473, N3468, N1747, N3365, N1615);
not NOT1 (N3474, N3467);
nor NOR3 (N3475, N3427, N1818, N1914);
nor NOR2 (N3476, N3475, N2605);
not NOT1 (N3477, N3463);
not NOT1 (N3478, N3474);
buf BUF1 (N3479, N3472);
nor NOR4 (N3480, N3477, N2328, N1288, N70);
nand NAND4 (N3481, N3473, N352, N220, N2817);
or OR4 (N3482, N3464, N141, N2071, N207);
nand NAND4 (N3483, N3480, N1074, N1334, N2803);
buf BUF1 (N3484, N3455);
not NOT1 (N3485, N3476);
or OR4 (N3486, N3484, N2938, N2461, N2982);
nor NOR2 (N3487, N3469, N872);
xor XOR2 (N3488, N3487, N181);
and AND3 (N3489, N3483, N1874, N873);
buf BUF1 (N3490, N3486);
nor NOR4 (N3491, N3482, N2096, N3140, N2341);
buf BUF1 (N3492, N3489);
and AND2 (N3493, N3471, N923);
buf BUF1 (N3494, N3488);
xor XOR2 (N3495, N3491, N1186);
not NOT1 (N3496, N3481);
nand NAND2 (N3497, N3490, N2595);
nand NAND3 (N3498, N3438, N847, N866);
not NOT1 (N3499, N3496);
buf BUF1 (N3500, N3495);
xor XOR2 (N3501, N3485, N220);
xor XOR2 (N3502, N3492, N1076);
or OR4 (N3503, N3479, N231, N2263, N1356);
buf BUF1 (N3504, N3478);
nand NAND4 (N3505, N3493, N1735, N1886, N496);
xor XOR2 (N3506, N3505, N342);
and AND2 (N3507, N3494, N2961);
xor XOR2 (N3508, N3507, N2475);
xor XOR2 (N3509, N3498, N1012);
nand NAND4 (N3510, N3508, N2786, N793, N2235);
xor XOR2 (N3511, N3506, N962);
nand NAND4 (N3512, N3510, N1924, N2868, N1177);
and AND2 (N3513, N3504, N1361);
nor NOR4 (N3514, N3512, N210, N2461, N3029);
and AND2 (N3515, N3502, N1364);
xor XOR2 (N3516, N3501, N1160);
and AND3 (N3517, N3509, N2179, N554);
nor NOR3 (N3518, N3503, N1265, N1724);
nand NAND4 (N3519, N3500, N3104, N1814, N2905);
or OR4 (N3520, N3499, N1824, N2526, N1681);
nand NAND2 (N3521, N3519, N1085);
nand NAND3 (N3522, N3520, N2980, N1339);
or OR3 (N3523, N3513, N64, N2092);
and AND2 (N3524, N3522, N578);
xor XOR2 (N3525, N3524, N1243);
nor NOR4 (N3526, N3523, N2282, N3455, N1783);
xor XOR2 (N3527, N3518, N2138);
not NOT1 (N3528, N3525);
or OR4 (N3529, N3527, N1885, N2033, N240);
and AND2 (N3530, N3528, N1234);
nand NAND2 (N3531, N3529, N2540);
xor XOR2 (N3532, N3514, N347);
not NOT1 (N3533, N3526);
not NOT1 (N3534, N3517);
and AND3 (N3535, N3497, N153, N1749);
nand NAND2 (N3536, N3532, N4);
or OR3 (N3537, N3521, N128, N1288);
xor XOR2 (N3538, N3535, N764);
buf BUF1 (N3539, N3538);
not NOT1 (N3540, N3536);
nand NAND3 (N3541, N3511, N2058, N1006);
or OR3 (N3542, N3516, N1269, N3114);
and AND3 (N3543, N3539, N253, N1437);
buf BUF1 (N3544, N3515);
xor XOR2 (N3545, N3531, N2505);
nor NOR3 (N3546, N3545, N2705, N1399);
xor XOR2 (N3547, N3543, N898);
nand NAND4 (N3548, N3547, N96, N1477, N1107);
or OR3 (N3549, N3540, N2528, N347);
xor XOR2 (N3550, N3544, N1857);
not NOT1 (N3551, N3549);
xor XOR2 (N3552, N3550, N1522);
nand NAND3 (N3553, N3530, N510, N2472);
xor XOR2 (N3554, N3553, N2437);
buf BUF1 (N3555, N3551);
not NOT1 (N3556, N3537);
xor XOR2 (N3557, N3555, N114);
xor XOR2 (N3558, N3557, N1338);
and AND3 (N3559, N3541, N1689, N324);
nand NAND4 (N3560, N3558, N113, N843, N897);
nand NAND2 (N3561, N3554, N2753);
or OR2 (N3562, N3534, N3357);
or OR4 (N3563, N3548, N2795, N2714, N1868);
not NOT1 (N3564, N3563);
and AND4 (N3565, N3542, N183, N1032, N820);
or OR4 (N3566, N3533, N1726, N2745, N3332);
not NOT1 (N3567, N3564);
nor NOR3 (N3568, N3560, N766, N2661);
or OR2 (N3569, N3561, N2638);
nor NOR3 (N3570, N3565, N1336, N1976);
nor NOR2 (N3571, N3570, N720);
and AND4 (N3572, N3552, N2743, N1437, N470);
or OR4 (N3573, N3571, N1291, N2439, N2613);
buf BUF1 (N3574, N3567);
nand NAND4 (N3575, N3574, N1167, N1441, N3341);
buf BUF1 (N3576, N3556);
xor XOR2 (N3577, N3566, N1140);
nand NAND4 (N3578, N3575, N1187, N1928, N138);
not NOT1 (N3579, N3569);
nor NOR2 (N3580, N3577, N1712);
and AND4 (N3581, N3576, N2748, N2149, N2768);
buf BUF1 (N3582, N3580);
or OR3 (N3583, N3559, N2863, N2135);
nand NAND3 (N3584, N3562, N632, N3364);
and AND2 (N3585, N3573, N2945);
and AND3 (N3586, N3583, N630, N2558);
nor NOR2 (N3587, N3586, N2147);
buf BUF1 (N3588, N3578);
not NOT1 (N3589, N3584);
or OR3 (N3590, N3572, N757, N3560);
nand NAND3 (N3591, N3590, N1628, N2835);
xor XOR2 (N3592, N3591, N892);
or OR2 (N3593, N3589, N1309);
buf BUF1 (N3594, N3582);
nor NOR3 (N3595, N3587, N3064, N2396);
xor XOR2 (N3596, N3592, N660);
and AND3 (N3597, N3596, N698, N2385);
nor NOR3 (N3598, N3585, N3004, N2435);
xor XOR2 (N3599, N3593, N538);
and AND3 (N3600, N3595, N539, N1649);
xor XOR2 (N3601, N3546, N1283);
xor XOR2 (N3602, N3581, N2950);
and AND2 (N3603, N3579, N2874);
buf BUF1 (N3604, N3602);
xor XOR2 (N3605, N3599, N2158);
not NOT1 (N3606, N3588);
buf BUF1 (N3607, N3568);
nor NOR3 (N3608, N3594, N2181, N3288);
nand NAND4 (N3609, N3608, N410, N2742, N1259);
not NOT1 (N3610, N3597);
nand NAND2 (N3611, N3609, N3133);
not NOT1 (N3612, N3607);
nor NOR4 (N3613, N3603, N2631, N341, N1962);
nand NAND2 (N3614, N3605, N195);
not NOT1 (N3615, N3611);
nand NAND4 (N3616, N3598, N193, N267, N3105);
nor NOR2 (N3617, N3601, N2966);
nand NAND4 (N3618, N3614, N3119, N2074, N389);
buf BUF1 (N3619, N3613);
buf BUF1 (N3620, N3616);
buf BUF1 (N3621, N3600);
buf BUF1 (N3622, N3604);
and AND3 (N3623, N3619, N1405, N1620);
or OR2 (N3624, N3620, N1904);
xor XOR2 (N3625, N3621, N3529);
nor NOR4 (N3626, N3618, N2138, N2884, N1534);
not NOT1 (N3627, N3617);
xor XOR2 (N3628, N3623, N761);
or OR4 (N3629, N3615, N1932, N1179, N3153);
and AND3 (N3630, N3629, N391, N3627);
or OR2 (N3631, N2954, N2243);
nand NAND4 (N3632, N3612, N189, N453, N1532);
buf BUF1 (N3633, N3626);
xor XOR2 (N3634, N3625, N2340);
not NOT1 (N3635, N3633);
nand NAND3 (N3636, N3634, N3321, N2935);
xor XOR2 (N3637, N3610, N800);
nand NAND4 (N3638, N3636, N1048, N2169, N326);
or OR3 (N3639, N3631, N158, N1565);
buf BUF1 (N3640, N3638);
xor XOR2 (N3641, N3640, N264);
and AND3 (N3642, N3632, N3121, N1130);
and AND2 (N3643, N3628, N38);
nor NOR2 (N3644, N3624, N1654);
buf BUF1 (N3645, N3606);
xor XOR2 (N3646, N3635, N171);
or OR2 (N3647, N3622, N3147);
xor XOR2 (N3648, N3637, N2481);
not NOT1 (N3649, N3630);
buf BUF1 (N3650, N3642);
or OR3 (N3651, N3645, N640, N278);
and AND4 (N3652, N3643, N137, N2155, N1102);
or OR2 (N3653, N3641, N882);
nand NAND2 (N3654, N3650, N1951);
or OR3 (N3655, N3653, N1763, N526);
nor NOR2 (N3656, N3649, N1011);
nor NOR2 (N3657, N3656, N1171);
buf BUF1 (N3658, N3651);
nand NAND2 (N3659, N3657, N289);
not NOT1 (N3660, N3647);
or OR2 (N3661, N3655, N1492);
nand NAND4 (N3662, N3646, N2364, N2089, N1801);
buf BUF1 (N3663, N3662);
and AND2 (N3664, N3639, N123);
or OR2 (N3665, N3654, N3182);
xor XOR2 (N3666, N3664, N2544);
xor XOR2 (N3667, N3661, N2135);
nand NAND3 (N3668, N3658, N3405, N313);
not NOT1 (N3669, N3648);
nor NOR3 (N3670, N3663, N3418, N3504);
xor XOR2 (N3671, N3670, N2996);
not NOT1 (N3672, N3666);
and AND3 (N3673, N3665, N1533, N849);
and AND4 (N3674, N3667, N634, N444, N3277);
or OR4 (N3675, N3652, N1446, N540, N624);
nor NOR3 (N3676, N3675, N575, N2977);
buf BUF1 (N3677, N3668);
and AND2 (N3678, N3676, N2624);
not NOT1 (N3679, N3660);
or OR3 (N3680, N3659, N3611, N2577);
or OR2 (N3681, N3672, N1069);
and AND3 (N3682, N3678, N3049, N143);
and AND4 (N3683, N3669, N590, N2664, N1916);
or OR2 (N3684, N3671, N2533);
xor XOR2 (N3685, N3644, N1703);
nor NOR2 (N3686, N3677, N2359);
nand NAND3 (N3687, N3674, N1327, N322);
or OR4 (N3688, N3687, N3663, N3000, N3229);
nor NOR3 (N3689, N3688, N497, N1721);
buf BUF1 (N3690, N3682);
xor XOR2 (N3691, N3679, N1678);
nand NAND2 (N3692, N3685, N2588);
not NOT1 (N3693, N3690);
or OR3 (N3694, N3673, N3247, N3013);
buf BUF1 (N3695, N3686);
xor XOR2 (N3696, N3692, N2827);
buf BUF1 (N3697, N3681);
xor XOR2 (N3698, N3697, N742);
buf BUF1 (N3699, N3695);
nand NAND3 (N3700, N3694, N292, N3594);
nor NOR2 (N3701, N3691, N2962);
and AND2 (N3702, N3699, N1079);
nor NOR2 (N3703, N3698, N996);
xor XOR2 (N3704, N3702, N475);
buf BUF1 (N3705, N3680);
xor XOR2 (N3706, N3684, N20);
xor XOR2 (N3707, N3700, N1384);
xor XOR2 (N3708, N3703, N2972);
nor NOR4 (N3709, N3693, N232, N1737, N2741);
and AND3 (N3710, N3701, N3483, N1973);
or OR2 (N3711, N3710, N1689);
nor NOR4 (N3712, N3708, N2090, N3082, N2390);
not NOT1 (N3713, N3712);
and AND2 (N3714, N3696, N2938);
not NOT1 (N3715, N3706);
xor XOR2 (N3716, N3683, N2234);
and AND2 (N3717, N3705, N985);
buf BUF1 (N3718, N3717);
or OR4 (N3719, N3689, N1904, N1134, N2319);
nand NAND2 (N3720, N3713, N681);
and AND3 (N3721, N3718, N2283, N3068);
and AND4 (N3722, N3711, N2260, N1774, N3582);
and AND4 (N3723, N3722, N1476, N2297, N3436);
xor XOR2 (N3724, N3709, N1754);
xor XOR2 (N3725, N3719, N1496);
xor XOR2 (N3726, N3707, N880);
and AND2 (N3727, N3725, N2963);
xor XOR2 (N3728, N3715, N2652);
or OR3 (N3729, N3723, N762, N1907);
and AND4 (N3730, N3714, N2493, N3257, N3203);
not NOT1 (N3731, N3730);
xor XOR2 (N3732, N3720, N3236);
buf BUF1 (N3733, N3728);
not NOT1 (N3734, N3733);
buf BUF1 (N3735, N3724);
and AND3 (N3736, N3732, N325, N798);
not NOT1 (N3737, N3735);
not NOT1 (N3738, N3721);
nand NAND4 (N3739, N3704, N2094, N1727, N2299);
not NOT1 (N3740, N3727);
not NOT1 (N3741, N3740);
nand NAND4 (N3742, N3741, N2686, N2699, N2377);
or OR4 (N3743, N3742, N924, N3042, N2317);
nor NOR3 (N3744, N3729, N1366, N3717);
nand NAND4 (N3745, N3738, N1969, N644, N3476);
and AND3 (N3746, N3731, N1724, N2881);
nand NAND3 (N3747, N3744, N2079, N2120);
or OR3 (N3748, N3739, N199, N2923);
nor NOR4 (N3749, N3737, N2520, N1919, N2162);
or OR2 (N3750, N3743, N2948);
nand NAND3 (N3751, N3734, N2487, N343);
nand NAND2 (N3752, N3736, N2582);
and AND3 (N3753, N3716, N364, N1455);
or OR4 (N3754, N3750, N1213, N541, N3440);
xor XOR2 (N3755, N3752, N3080);
and AND2 (N3756, N3726, N1397);
not NOT1 (N3757, N3748);
not NOT1 (N3758, N3754);
nand NAND2 (N3759, N3755, N630);
xor XOR2 (N3760, N3749, N1139);
nand NAND2 (N3761, N3759, N2176);
and AND4 (N3762, N3757, N1438, N3113, N1142);
xor XOR2 (N3763, N3753, N2743);
nor NOR4 (N3764, N3763, N2382, N3606, N2467);
xor XOR2 (N3765, N3747, N436);
nor NOR2 (N3766, N3745, N210);
nand NAND2 (N3767, N3751, N3289);
and AND2 (N3768, N3765, N1516);
nand NAND4 (N3769, N3761, N2676, N1181, N3175);
nand NAND4 (N3770, N3769, N1550, N2571, N3184);
nor NOR2 (N3771, N3758, N3398);
buf BUF1 (N3772, N3756);
nor NOR2 (N3773, N3770, N3712);
xor XOR2 (N3774, N3767, N335);
and AND4 (N3775, N3772, N1309, N844, N3058);
and AND3 (N3776, N3768, N1524, N1215);
buf BUF1 (N3777, N3760);
buf BUF1 (N3778, N3764);
or OR2 (N3779, N3762, N2460);
buf BUF1 (N3780, N3774);
not NOT1 (N3781, N3775);
nor NOR2 (N3782, N3773, N1653);
or OR3 (N3783, N3780, N1633, N689);
and AND2 (N3784, N3777, N324);
and AND2 (N3785, N3776, N3646);
buf BUF1 (N3786, N3784);
buf BUF1 (N3787, N3786);
nor NOR3 (N3788, N3782, N2404, N3692);
buf BUF1 (N3789, N3788);
or OR2 (N3790, N3766, N161);
or OR4 (N3791, N3779, N2760, N1332, N907);
xor XOR2 (N3792, N3781, N228);
nand NAND3 (N3793, N3787, N973, N880);
nor NOR3 (N3794, N3789, N1392, N1135);
or OR2 (N3795, N3794, N1881);
and AND4 (N3796, N3746, N191, N1369, N3733);
nor NOR3 (N3797, N3771, N2068, N1878);
and AND2 (N3798, N3793, N1443);
buf BUF1 (N3799, N3785);
not NOT1 (N3800, N3783);
not NOT1 (N3801, N3792);
xor XOR2 (N3802, N3797, N2061);
not NOT1 (N3803, N3801);
buf BUF1 (N3804, N3790);
buf BUF1 (N3805, N3791);
buf BUF1 (N3806, N3803);
nand NAND3 (N3807, N3800, N3084, N1438);
and AND2 (N3808, N3778, N875);
buf BUF1 (N3809, N3807);
not NOT1 (N3810, N3802);
and AND4 (N3811, N3796, N909, N2014, N781);
and AND4 (N3812, N3795, N3633, N2449, N3654);
and AND2 (N3813, N3804, N2885);
buf BUF1 (N3814, N3798);
nand NAND2 (N3815, N3814, N372);
nand NAND3 (N3816, N3805, N1334, N80);
buf BUF1 (N3817, N3810);
and AND3 (N3818, N3811, N112, N3324);
buf BUF1 (N3819, N3812);
xor XOR2 (N3820, N3815, N1349);
or OR2 (N3821, N3816, N2224);
and AND3 (N3822, N3818, N3044, N2784);
and AND3 (N3823, N3819, N1764, N162);
or OR2 (N3824, N3821, N1708);
buf BUF1 (N3825, N3799);
xor XOR2 (N3826, N3817, N2252);
and AND2 (N3827, N3820, N1749);
not NOT1 (N3828, N3825);
nand NAND2 (N3829, N3809, N3744);
buf BUF1 (N3830, N3829);
buf BUF1 (N3831, N3808);
nand NAND2 (N3832, N3813, N2075);
nand NAND3 (N3833, N3828, N3252, N3547);
nand NAND3 (N3834, N3831, N403, N2356);
buf BUF1 (N3835, N3826);
nand NAND3 (N3836, N3822, N497, N2877);
nand NAND4 (N3837, N3806, N2575, N3597, N3833);
nor NOR2 (N3838, N2090, N1638);
or OR2 (N3839, N3837, N2941);
xor XOR2 (N3840, N3835, N1862);
not NOT1 (N3841, N3823);
not NOT1 (N3842, N3827);
nand NAND2 (N3843, N3830, N3099);
nor NOR4 (N3844, N3839, N3843, N1851, N1137);
xor XOR2 (N3845, N1038, N251);
nor NOR4 (N3846, N3841, N3404, N3609, N1773);
xor XOR2 (N3847, N3824, N2081);
xor XOR2 (N3848, N3838, N1557);
buf BUF1 (N3849, N3836);
buf BUF1 (N3850, N3845);
or OR4 (N3851, N3844, N2541, N1864, N43);
not NOT1 (N3852, N3840);
or OR3 (N3853, N3846, N2542, N2587);
not NOT1 (N3854, N3852);
not NOT1 (N3855, N3854);
xor XOR2 (N3856, N3834, N3033);
buf BUF1 (N3857, N3847);
buf BUF1 (N3858, N3855);
nor NOR4 (N3859, N3851, N1086, N3073, N3764);
nand NAND2 (N3860, N3857, N2076);
and AND3 (N3861, N3856, N3278, N3588);
nand NAND3 (N3862, N3842, N2062, N2082);
not NOT1 (N3863, N3860);
or OR3 (N3864, N3832, N539, N3493);
nand NAND2 (N3865, N3853, N2651);
buf BUF1 (N3866, N3858);
nand NAND3 (N3867, N3865, N3813, N1324);
nand NAND2 (N3868, N3859, N1584);
or OR4 (N3869, N3850, N192, N3642, N1000);
not NOT1 (N3870, N3868);
nor NOR4 (N3871, N3866, N2705, N1135, N1076);
nor NOR3 (N3872, N3871, N2919, N2104);
or OR4 (N3873, N3849, N386, N1740, N360);
xor XOR2 (N3874, N3864, N2792);
nor NOR4 (N3875, N3863, N1434, N916, N1137);
not NOT1 (N3876, N3874);
xor XOR2 (N3877, N3861, N802);
xor XOR2 (N3878, N3862, N3762);
xor XOR2 (N3879, N3873, N425);
xor XOR2 (N3880, N3870, N2097);
nand NAND4 (N3881, N3879, N1747, N2515, N999);
xor XOR2 (N3882, N3869, N610);
buf BUF1 (N3883, N3877);
or OR2 (N3884, N3867, N3344);
and AND2 (N3885, N3880, N2502);
or OR2 (N3886, N3878, N3341);
xor XOR2 (N3887, N3876, N2497);
or OR2 (N3888, N3883, N3516);
nor NOR2 (N3889, N3887, N1190);
buf BUF1 (N3890, N3875);
and AND2 (N3891, N3881, N638);
not NOT1 (N3892, N3890);
or OR2 (N3893, N3891, N2649);
and AND2 (N3894, N3886, N1417);
not NOT1 (N3895, N3892);
or OR4 (N3896, N3872, N1934, N1371, N2462);
or OR3 (N3897, N3882, N387, N2335);
not NOT1 (N3898, N3848);
not NOT1 (N3899, N3894);
and AND4 (N3900, N3888, N1500, N12, N2400);
or OR2 (N3901, N3896, N2392);
buf BUF1 (N3902, N3901);
or OR3 (N3903, N3897, N733, N2673);
not NOT1 (N3904, N3903);
nor NOR2 (N3905, N3900, N1596);
not NOT1 (N3906, N3899);
nor NOR2 (N3907, N3906, N1528);
not NOT1 (N3908, N3895);
and AND4 (N3909, N3904, N3712, N3123, N2658);
or OR4 (N3910, N3898, N1380, N1557, N1995);
not NOT1 (N3911, N3908);
xor XOR2 (N3912, N3911, N2251);
and AND2 (N3913, N3912, N3696);
buf BUF1 (N3914, N3889);
nand NAND3 (N3915, N3902, N1042, N3177);
and AND3 (N3916, N3913, N2248, N3284);
nand NAND4 (N3917, N3907, N822, N3808, N3618);
nand NAND4 (N3918, N3916, N1224, N1940, N2704);
or OR3 (N3919, N3917, N2383, N1284);
xor XOR2 (N3920, N3884, N1366);
buf BUF1 (N3921, N3885);
or OR4 (N3922, N3921, N953, N2355, N262);
buf BUF1 (N3923, N3922);
not NOT1 (N3924, N3905);
nor NOR3 (N3925, N3923, N2348, N1626);
nand NAND2 (N3926, N3909, N3445);
not NOT1 (N3927, N3910);
xor XOR2 (N3928, N3924, N2102);
not NOT1 (N3929, N3914);
or OR4 (N3930, N3915, N3863, N3461, N3287);
nand NAND3 (N3931, N3919, N944, N209);
nor NOR2 (N3932, N3925, N2870);
xor XOR2 (N3933, N3918, N3121);
and AND2 (N3934, N3933, N320);
not NOT1 (N3935, N3920);
xor XOR2 (N3936, N3934, N910);
not NOT1 (N3937, N3931);
nand NAND3 (N3938, N3928, N1046, N1018);
or OR3 (N3939, N3893, N1089, N3660);
xor XOR2 (N3940, N3937, N2132);
and AND2 (N3941, N3939, N3595);
or OR3 (N3942, N3936, N1708, N3593);
not NOT1 (N3943, N3938);
nor NOR2 (N3944, N3927, N1366);
buf BUF1 (N3945, N3942);
buf BUF1 (N3946, N3944);
or OR3 (N3947, N3926, N1293, N1337);
nand NAND4 (N3948, N3935, N1663, N1439, N732);
not NOT1 (N3949, N3948);
not NOT1 (N3950, N3949);
or OR3 (N3951, N3940, N1622, N164);
not NOT1 (N3952, N3951);
or OR4 (N3953, N3945, N3836, N3116, N3710);
and AND4 (N3954, N3947, N793, N227, N592);
xor XOR2 (N3955, N3953, N3722);
and AND3 (N3956, N3943, N1126, N1651);
not NOT1 (N3957, N3932);
buf BUF1 (N3958, N3952);
and AND2 (N3959, N3957, N1422);
buf BUF1 (N3960, N3930);
xor XOR2 (N3961, N3946, N3478);
or OR3 (N3962, N3960, N1656, N338);
or OR4 (N3963, N3954, N58, N2152, N3070);
not NOT1 (N3964, N3941);
buf BUF1 (N3965, N3964);
xor XOR2 (N3966, N3959, N1764);
and AND4 (N3967, N3929, N147, N3209, N3374);
xor XOR2 (N3968, N3962, N3743);
buf BUF1 (N3969, N3956);
or OR4 (N3970, N3950, N3681, N3920, N2875);
and AND3 (N3971, N3967, N923, N3368);
nand NAND3 (N3972, N3969, N3857, N2080);
nand NAND2 (N3973, N3966, N3820);
nand NAND3 (N3974, N3968, N2443, N2729);
nor NOR3 (N3975, N3961, N2800, N2939);
xor XOR2 (N3976, N3973, N3232);
or OR2 (N3977, N3971, N3209);
nor NOR3 (N3978, N3977, N3753, N313);
not NOT1 (N3979, N3978);
or OR3 (N3980, N3974, N1817, N1280);
and AND4 (N3981, N3963, N1411, N973, N2915);
not NOT1 (N3982, N3972);
nand NAND2 (N3983, N3980, N3866);
xor XOR2 (N3984, N3976, N3808);
xor XOR2 (N3985, N3981, N35);
and AND2 (N3986, N3965, N275);
buf BUF1 (N3987, N3985);
xor XOR2 (N3988, N3987, N3378);
or OR2 (N3989, N3958, N2137);
and AND4 (N3990, N3989, N1888, N536, N3134);
nand NAND3 (N3991, N3979, N2096, N1048);
nor NOR4 (N3992, N3970, N1752, N2975, N1096);
and AND2 (N3993, N3991, N76);
xor XOR2 (N3994, N3975, N331);
and AND3 (N3995, N3986, N3111, N2512);
buf BUF1 (N3996, N3982);
buf BUF1 (N3997, N3988);
nand NAND2 (N3998, N3992, N2461);
buf BUF1 (N3999, N3983);
and AND4 (N4000, N3990, N176, N2597, N1196);
nand NAND4 (N4001, N3998, N917, N3614, N3662);
xor XOR2 (N4002, N3995, N1817);
nor NOR4 (N4003, N4002, N2595, N1063, N122);
not NOT1 (N4004, N4001);
nand NAND3 (N4005, N3993, N1450, N2724);
nand NAND3 (N4006, N4005, N831, N1229);
xor XOR2 (N4007, N3996, N1393);
and AND3 (N4008, N4004, N3128, N2989);
buf BUF1 (N4009, N4003);
and AND4 (N4010, N4007, N2095, N3193, N2954);
and AND2 (N4011, N4009, N3320);
buf BUF1 (N4012, N3999);
buf BUF1 (N4013, N4000);
xor XOR2 (N4014, N3984, N1370);
xor XOR2 (N4015, N4012, N191);
and AND3 (N4016, N3997, N3277, N3392);
nand NAND3 (N4017, N4015, N1074, N3194);
or OR3 (N4018, N4008, N3750, N1030);
buf BUF1 (N4019, N4011);
nor NOR2 (N4020, N4013, N3381);
nor NOR2 (N4021, N4014, N3748);
buf BUF1 (N4022, N4010);
and AND3 (N4023, N4022, N1944, N1728);
and AND2 (N4024, N4006, N2510);
or OR2 (N4025, N4021, N396);
buf BUF1 (N4026, N4018);
not NOT1 (N4027, N4019);
nand NAND3 (N4028, N4025, N1840, N2326);
and AND4 (N4029, N4027, N2874, N979, N1470);
buf BUF1 (N4030, N4026);
nor NOR3 (N4031, N3994, N3919, N2037);
buf BUF1 (N4032, N4020);
buf BUF1 (N4033, N4028);
buf BUF1 (N4034, N4023);
and AND4 (N4035, N4033, N1483, N1294, N25);
xor XOR2 (N4036, N4024, N3424);
not NOT1 (N4037, N3955);
or OR2 (N4038, N4031, N1118);
buf BUF1 (N4039, N4032);
xor XOR2 (N4040, N4039, N3453);
nand NAND2 (N4041, N4016, N3039);
buf BUF1 (N4042, N4041);
not NOT1 (N4043, N4038);
nor NOR4 (N4044, N4034, N3646, N3329, N2947);
or OR4 (N4045, N4037, N279, N3168, N1873);
buf BUF1 (N4046, N4042);
or OR2 (N4047, N4040, N580);
or OR4 (N4048, N4035, N523, N2079, N3258);
xor XOR2 (N4049, N4045, N960);
nor NOR4 (N4050, N4030, N3413, N1890, N718);
xor XOR2 (N4051, N4044, N2096);
or OR4 (N4052, N4046, N3499, N2060, N549);
or OR3 (N4053, N4029, N1167, N2256);
nand NAND4 (N4054, N4047, N3911, N962, N593);
xor XOR2 (N4055, N4053, N61);
xor XOR2 (N4056, N4017, N1187);
and AND2 (N4057, N4052, N1642);
nand NAND4 (N4058, N4054, N414, N2848, N301);
nand NAND3 (N4059, N4058, N3970, N35);
or OR2 (N4060, N4036, N1544);
xor XOR2 (N4061, N4050, N3134);
or OR4 (N4062, N4055, N396, N345, N100);
xor XOR2 (N4063, N4043, N328);
nor NOR3 (N4064, N4048, N3332, N3165);
nor NOR2 (N4065, N4060, N1307);
buf BUF1 (N4066, N4056);
nand NAND4 (N4067, N4061, N2889, N3873, N2653);
nand NAND4 (N4068, N4059, N567, N1091, N642);
nor NOR4 (N4069, N4065, N1934, N1231, N2909);
or OR4 (N4070, N4051, N169, N458, N2861);
xor XOR2 (N4071, N4057, N2280);
or OR3 (N4072, N4049, N1736, N2009);
not NOT1 (N4073, N4069);
and AND3 (N4074, N4063, N35, N1041);
nor NOR3 (N4075, N4071, N3091, N3418);
buf BUF1 (N4076, N4067);
nand NAND3 (N4077, N4062, N2836, N2539);
or OR4 (N4078, N4064, N878, N766, N1742);
nand NAND2 (N4079, N4066, N216);
nand NAND2 (N4080, N4075, N2117);
and AND3 (N4081, N4073, N3924, N1676);
not NOT1 (N4082, N4076);
nor NOR4 (N4083, N4074, N1424, N3840, N2973);
nand NAND3 (N4084, N4078, N843, N3302);
or OR4 (N4085, N4072, N2057, N1612, N3229);
not NOT1 (N4086, N4080);
nor NOR4 (N4087, N4079, N534, N257, N3934);
buf BUF1 (N4088, N4082);
not NOT1 (N4089, N4086);
nand NAND3 (N4090, N4083, N296, N265);
buf BUF1 (N4091, N4084);
not NOT1 (N4092, N4070);
and AND3 (N4093, N4081, N484, N3840);
and AND4 (N4094, N4090, N3233, N445, N2693);
nand NAND3 (N4095, N4089, N1334, N1064);
buf BUF1 (N4096, N4093);
nor NOR2 (N4097, N4091, N1502);
xor XOR2 (N4098, N4097, N414);
not NOT1 (N4099, N4068);
not NOT1 (N4100, N4094);
not NOT1 (N4101, N4099);
nand NAND4 (N4102, N4087, N3136, N3122, N2699);
xor XOR2 (N4103, N4088, N2870);
nor NOR3 (N4104, N4096, N3225, N369);
buf BUF1 (N4105, N4100);
nand NAND2 (N4106, N4085, N2263);
and AND3 (N4107, N4095, N3682, N2040);
nand NAND4 (N4108, N4107, N622, N1102, N3265);
nor NOR2 (N4109, N4106, N364);
buf BUF1 (N4110, N4104);
xor XOR2 (N4111, N4105, N3559);
or OR3 (N4112, N4103, N726, N1038);
xor XOR2 (N4113, N4110, N42);
nand NAND3 (N4114, N4102, N1303, N2693);
not NOT1 (N4115, N4092);
not NOT1 (N4116, N4109);
nor NOR4 (N4117, N4114, N3122, N376, N1586);
buf BUF1 (N4118, N4111);
nand NAND2 (N4119, N4116, N1711);
xor XOR2 (N4120, N4118, N505);
nand NAND3 (N4121, N4098, N3965, N1392);
nor NOR4 (N4122, N4108, N1920, N1737, N267);
not NOT1 (N4123, N4077);
nand NAND2 (N4124, N4121, N1701);
not NOT1 (N4125, N4124);
not NOT1 (N4126, N4119);
and AND2 (N4127, N4101, N586);
not NOT1 (N4128, N4117);
buf BUF1 (N4129, N4127);
buf BUF1 (N4130, N4128);
xor XOR2 (N4131, N4126, N1798);
not NOT1 (N4132, N4113);
nand NAND4 (N4133, N4132, N3866, N2508, N186);
not NOT1 (N4134, N4115);
buf BUF1 (N4135, N4123);
or OR3 (N4136, N4130, N3069, N3122);
nand NAND3 (N4137, N4120, N1, N723);
xor XOR2 (N4138, N4131, N3283);
nor NOR3 (N4139, N4125, N1945, N1559);
buf BUF1 (N4140, N4135);
nor NOR4 (N4141, N4112, N279, N3629, N1318);
or OR4 (N4142, N4134, N1025, N1343, N3137);
nor NOR4 (N4143, N4136, N4020, N1189, N725);
buf BUF1 (N4144, N4141);
xor XOR2 (N4145, N4144, N3695);
nor NOR3 (N4146, N4137, N1942, N3131);
buf BUF1 (N4147, N4122);
xor XOR2 (N4148, N4138, N3475);
and AND3 (N4149, N4147, N3641, N2768);
and AND2 (N4150, N4140, N3253);
xor XOR2 (N4151, N4129, N13);
not NOT1 (N4152, N4151);
buf BUF1 (N4153, N4145);
buf BUF1 (N4154, N4152);
xor XOR2 (N4155, N4146, N1898);
or OR3 (N4156, N4148, N3638, N754);
not NOT1 (N4157, N4154);
or OR3 (N4158, N4155, N933, N342);
xor XOR2 (N4159, N4158, N495);
or OR2 (N4160, N4157, N1626);
not NOT1 (N4161, N4139);
nand NAND4 (N4162, N4160, N1324, N3986, N1994);
nor NOR3 (N4163, N4156, N2612, N3888);
and AND4 (N4164, N4161, N3018, N673, N2181);
buf BUF1 (N4165, N4133);
or OR2 (N4166, N4165, N3320);
and AND2 (N4167, N4164, N956);
not NOT1 (N4168, N4159);
buf BUF1 (N4169, N4149);
not NOT1 (N4170, N4142);
buf BUF1 (N4171, N4170);
buf BUF1 (N4172, N4163);
and AND4 (N4173, N4143, N1740, N1959, N3550);
nor NOR4 (N4174, N4171, N2467, N3750, N907);
nand NAND4 (N4175, N4166, N48, N3580, N1631);
nand NAND4 (N4176, N4169, N1241, N1303, N1166);
buf BUF1 (N4177, N4176);
nand NAND3 (N4178, N4174, N3099, N2175);
or OR4 (N4179, N4178, N3048, N3484, N1644);
nor NOR2 (N4180, N4162, N2973);
not NOT1 (N4181, N4167);
not NOT1 (N4182, N4177);
or OR4 (N4183, N4175, N1799, N1681, N3267);
nand NAND4 (N4184, N4173, N2957, N1365, N1226);
nand NAND2 (N4185, N4181, N2256);
nand NAND4 (N4186, N4168, N628, N849, N2664);
not NOT1 (N4187, N4172);
xor XOR2 (N4188, N4184, N3661);
xor XOR2 (N4189, N4150, N1525);
nand NAND2 (N4190, N4188, N3083);
or OR2 (N4191, N4187, N3094);
nand NAND4 (N4192, N4180, N3311, N2893, N2605);
nand NAND3 (N4193, N4191, N1576, N2893);
buf BUF1 (N4194, N4186);
not NOT1 (N4195, N4183);
and AND3 (N4196, N4190, N1064, N1360);
nor NOR3 (N4197, N4195, N3996, N2794);
nand NAND3 (N4198, N4189, N1248, N1456);
or OR2 (N4199, N4193, N359);
nor NOR3 (N4200, N4194, N3895, N3307);
xor XOR2 (N4201, N4199, N1318);
buf BUF1 (N4202, N4200);
not NOT1 (N4203, N4196);
or OR3 (N4204, N4198, N2823, N54);
nand NAND4 (N4205, N4185, N2719, N3782, N1957);
or OR3 (N4206, N4202, N1417, N1658);
not NOT1 (N4207, N4206);
xor XOR2 (N4208, N4201, N1545);
nand NAND4 (N4209, N4205, N1110, N3408, N1798);
or OR2 (N4210, N4197, N1273);
and AND4 (N4211, N4210, N2822, N3748, N3832);
buf BUF1 (N4212, N4209);
not NOT1 (N4213, N4192);
not NOT1 (N4214, N4203);
nor NOR4 (N4215, N4212, N3963, N182, N493);
xor XOR2 (N4216, N4207, N3774);
xor XOR2 (N4217, N4179, N3818);
and AND3 (N4218, N4211, N1212, N2810);
buf BUF1 (N4219, N4208);
buf BUF1 (N4220, N4218);
xor XOR2 (N4221, N4219, N2015);
or OR2 (N4222, N4204, N2272);
not NOT1 (N4223, N4213);
nor NOR4 (N4224, N4153, N3316, N2258, N3932);
nor NOR4 (N4225, N4215, N2307, N3607, N1878);
or OR4 (N4226, N4217, N1907, N3981, N2195);
nor NOR4 (N4227, N4222, N2221, N1973, N1220);
nand NAND2 (N4228, N4214, N2981);
xor XOR2 (N4229, N4216, N2289);
xor XOR2 (N4230, N4228, N2911);
not NOT1 (N4231, N4229);
xor XOR2 (N4232, N4230, N1478);
or OR4 (N4233, N4227, N1028, N1860, N1349);
and AND3 (N4234, N4221, N2627, N1952);
nand NAND2 (N4235, N4234, N1658);
or OR3 (N4236, N4223, N914, N3558);
and AND2 (N4237, N4182, N2899);
nand NAND4 (N4238, N4236, N1014, N4222, N2766);
xor XOR2 (N4239, N4233, N3586);
or OR2 (N4240, N4226, N336);
not NOT1 (N4241, N4220);
or OR4 (N4242, N4224, N1591, N2889, N1828);
or OR3 (N4243, N4232, N4075, N3714);
nor NOR2 (N4244, N4231, N1671);
buf BUF1 (N4245, N4240);
not NOT1 (N4246, N4239);
nor NOR2 (N4247, N4246, N2279);
buf BUF1 (N4248, N4245);
buf BUF1 (N4249, N4242);
not NOT1 (N4250, N4237);
nand NAND2 (N4251, N4238, N643);
nor NOR4 (N4252, N4249, N241, N1324, N2637);
xor XOR2 (N4253, N4248, N3215);
and AND2 (N4254, N4253, N169);
buf BUF1 (N4255, N4247);
or OR4 (N4256, N4252, N4171, N1947, N2160);
not NOT1 (N4257, N4244);
nand NAND3 (N4258, N4257, N872, N578);
nor NOR3 (N4259, N4251, N2832, N2109);
or OR2 (N4260, N4250, N4258);
not NOT1 (N4261, N3923);
buf BUF1 (N4262, N4260);
buf BUF1 (N4263, N4255);
nand NAND3 (N4264, N4225, N1653, N3338);
xor XOR2 (N4265, N4262, N341);
xor XOR2 (N4266, N4263, N4062);
not NOT1 (N4267, N4256);
not NOT1 (N4268, N4265);
buf BUF1 (N4269, N4235);
or OR2 (N4270, N4267, N402);
xor XOR2 (N4271, N4243, N574);
nand NAND3 (N4272, N4254, N4037, N2980);
xor XOR2 (N4273, N4259, N319);
nand NAND4 (N4274, N4270, N3674, N3016, N2750);
not NOT1 (N4275, N4266);
nor NOR2 (N4276, N4272, N345);
not NOT1 (N4277, N4264);
buf BUF1 (N4278, N4241);
nand NAND4 (N4279, N4275, N2534, N2599, N697);
or OR3 (N4280, N4276, N1522, N2625);
xor XOR2 (N4281, N4279, N3974);
nor NOR2 (N4282, N4273, N1744);
nand NAND3 (N4283, N4274, N4177, N52);
xor XOR2 (N4284, N4271, N342);
not NOT1 (N4285, N4269);
xor XOR2 (N4286, N4282, N949);
not NOT1 (N4287, N4285);
nand NAND2 (N4288, N4281, N3488);
buf BUF1 (N4289, N4268);
xor XOR2 (N4290, N4278, N1988);
not NOT1 (N4291, N4286);
xor XOR2 (N4292, N4280, N2409);
and AND3 (N4293, N4284, N310, N3688);
nand NAND2 (N4294, N4287, N2504);
buf BUF1 (N4295, N4288);
xor XOR2 (N4296, N4277, N3550);
nor NOR3 (N4297, N4283, N2933, N216);
buf BUF1 (N4298, N4289);
buf BUF1 (N4299, N4291);
or OR4 (N4300, N4299, N3864, N2190, N550);
not NOT1 (N4301, N4261);
nand NAND2 (N4302, N4298, N3218);
or OR4 (N4303, N4290, N870, N2345, N878);
nand NAND3 (N4304, N4296, N4130, N2881);
buf BUF1 (N4305, N4297);
nor NOR4 (N4306, N4305, N1448, N2055, N1138);
and AND4 (N4307, N4303, N2767, N582, N278);
nor NOR2 (N4308, N4304, N4268);
or OR4 (N4309, N4293, N2425, N3854, N1286);
and AND3 (N4310, N4302, N1764, N1868);
not NOT1 (N4311, N4310);
nand NAND4 (N4312, N4307, N2878, N1059, N1728);
nand NAND2 (N4313, N4312, N3887);
buf BUF1 (N4314, N4306);
or OR2 (N4315, N4308, N3839);
or OR3 (N4316, N4314, N1493, N2747);
nand NAND3 (N4317, N4313, N294, N3768);
and AND2 (N4318, N4301, N4045);
nand NAND4 (N4319, N4292, N379, N3898, N3510);
not NOT1 (N4320, N4316);
nand NAND2 (N4321, N4319, N998);
nor NOR4 (N4322, N4309, N3984, N3394, N2287);
xor XOR2 (N4323, N4311, N356);
or OR4 (N4324, N4317, N91, N3209, N1667);
buf BUF1 (N4325, N4323);
buf BUF1 (N4326, N4295);
nor NOR2 (N4327, N4325, N1826);
not NOT1 (N4328, N4327);
and AND4 (N4329, N4315, N716, N1762, N1417);
or OR4 (N4330, N4324, N416, N274, N637);
not NOT1 (N4331, N4320);
buf BUF1 (N4332, N4329);
xor XOR2 (N4333, N4300, N1654);
or OR2 (N4334, N4322, N632);
not NOT1 (N4335, N4331);
or OR3 (N4336, N4328, N2369, N3880);
xor XOR2 (N4337, N4332, N1222);
or OR4 (N4338, N4326, N3212, N288, N1729);
or OR4 (N4339, N4335, N1304, N3161, N4258);
xor XOR2 (N4340, N4337, N3200);
nand NAND2 (N4341, N4294, N40);
and AND2 (N4342, N4338, N3803);
xor XOR2 (N4343, N4333, N3237);
or OR4 (N4344, N4339, N163, N3857, N1840);
and AND4 (N4345, N4341, N253, N871, N100);
xor XOR2 (N4346, N4345, N1900);
xor XOR2 (N4347, N4342, N208);
buf BUF1 (N4348, N4321);
nand NAND4 (N4349, N4334, N275, N262, N3318);
nand NAND2 (N4350, N4330, N1153);
nand NAND3 (N4351, N4346, N4240, N729);
buf BUF1 (N4352, N4318);
or OR2 (N4353, N4347, N609);
xor XOR2 (N4354, N4340, N511);
xor XOR2 (N4355, N4344, N1561);
and AND3 (N4356, N4343, N3445, N4345);
xor XOR2 (N4357, N4356, N436);
nand NAND4 (N4358, N4357, N100, N1502, N1935);
not NOT1 (N4359, N4354);
nor NOR2 (N4360, N4352, N4016);
and AND3 (N4361, N4355, N1776, N195);
nor NOR4 (N4362, N4361, N2439, N1438, N1863);
nor NOR3 (N4363, N4351, N1093, N4164);
xor XOR2 (N4364, N4353, N3313);
not NOT1 (N4365, N4348);
nand NAND4 (N4366, N4363, N1889, N176, N882);
or OR2 (N4367, N4362, N2313);
buf BUF1 (N4368, N4365);
xor XOR2 (N4369, N4364, N1103);
nand NAND3 (N4370, N4366, N1807, N3119);
xor XOR2 (N4371, N4350, N4124);
nor NOR4 (N4372, N4367, N3044, N2607, N464);
not NOT1 (N4373, N4371);
not NOT1 (N4374, N4373);
nor NOR3 (N4375, N4360, N1482, N2648);
and AND2 (N4376, N4358, N1263);
or OR2 (N4377, N4359, N4339);
nand NAND3 (N4378, N4370, N2592, N1069);
xor XOR2 (N4379, N4376, N2202);
and AND2 (N4380, N4378, N692);
or OR2 (N4381, N4377, N111);
xor XOR2 (N4382, N4368, N1934);
xor XOR2 (N4383, N4336, N602);
or OR2 (N4384, N4381, N3974);
nand NAND2 (N4385, N4384, N1982);
nor NOR4 (N4386, N4369, N2808, N3668, N688);
xor XOR2 (N4387, N4372, N470);
and AND3 (N4388, N4375, N350, N4030);
nand NAND2 (N4389, N4382, N4086);
or OR4 (N4390, N4387, N4155, N1593, N113);
nor NOR4 (N4391, N4388, N3862, N2324, N1072);
and AND3 (N4392, N4380, N4248, N1172);
xor XOR2 (N4393, N4379, N3634);
nand NAND2 (N4394, N4390, N3026);
buf BUF1 (N4395, N4393);
nor NOR2 (N4396, N4389, N1124);
buf BUF1 (N4397, N4383);
nand NAND2 (N4398, N4395, N572);
buf BUF1 (N4399, N4392);
nor NOR4 (N4400, N4386, N886, N3890, N276);
not NOT1 (N4401, N4400);
or OR3 (N4402, N4398, N1080, N835);
xor XOR2 (N4403, N4397, N3648);
nand NAND2 (N4404, N4391, N2290);
buf BUF1 (N4405, N4385);
buf BUF1 (N4406, N4349);
nand NAND2 (N4407, N4403, N494);
and AND2 (N4408, N4399, N345);
nand NAND4 (N4409, N4402, N373, N381, N3719);
not NOT1 (N4410, N4406);
and AND2 (N4411, N4409, N2246);
and AND2 (N4412, N4374, N3400);
nor NOR4 (N4413, N4394, N4178, N1454, N550);
not NOT1 (N4414, N4408);
and AND2 (N4415, N4413, N2794);
nor NOR4 (N4416, N4411, N437, N2538, N3638);
not NOT1 (N4417, N4410);
buf BUF1 (N4418, N4404);
buf BUF1 (N4419, N4416);
xor XOR2 (N4420, N4405, N1188);
xor XOR2 (N4421, N4396, N3715);
buf BUF1 (N4422, N4418);
or OR2 (N4423, N4422, N4205);
xor XOR2 (N4424, N4412, N1486);
or OR2 (N4425, N4423, N663);
buf BUF1 (N4426, N4415);
and AND2 (N4427, N4401, N4138);
xor XOR2 (N4428, N4407, N2751);
and AND4 (N4429, N4417, N1370, N2991, N1558);
buf BUF1 (N4430, N4421);
nor NOR4 (N4431, N4426, N1390, N1853, N2973);
buf BUF1 (N4432, N4430);
xor XOR2 (N4433, N4424, N4047);
or OR4 (N4434, N4429, N857, N3697, N2630);
buf BUF1 (N4435, N4419);
buf BUF1 (N4436, N4425);
and AND4 (N4437, N4414, N1646, N814, N2861);
buf BUF1 (N4438, N4433);
xor XOR2 (N4439, N4420, N3463);
xor XOR2 (N4440, N4437, N3637);
or OR3 (N4441, N4440, N568, N1832);
and AND3 (N4442, N4432, N2445, N1497);
xor XOR2 (N4443, N4431, N579);
xor XOR2 (N4444, N4436, N3319);
and AND2 (N4445, N4434, N2923);
nor NOR2 (N4446, N4442, N2461);
xor XOR2 (N4447, N4444, N3498);
not NOT1 (N4448, N4447);
buf BUF1 (N4449, N4445);
buf BUF1 (N4450, N4438);
or OR2 (N4451, N4441, N2654);
and AND2 (N4452, N4443, N2018);
nor NOR2 (N4453, N4451, N3372);
nand NAND2 (N4454, N4450, N3261);
nor NOR3 (N4455, N4439, N1858, N1079);
and AND2 (N4456, N4452, N2199);
nand NAND4 (N4457, N4446, N2542, N3904, N1725);
and AND2 (N4458, N4457, N3137);
buf BUF1 (N4459, N4454);
or OR2 (N4460, N4435, N49);
buf BUF1 (N4461, N4460);
nand NAND3 (N4462, N4453, N2295, N1725);
nand NAND3 (N4463, N4461, N405, N2757);
or OR2 (N4464, N4459, N3964);
or OR3 (N4465, N4427, N68, N2411);
and AND4 (N4466, N4428, N2618, N2203, N4272);
nor NOR3 (N4467, N4448, N817, N4394);
or OR4 (N4468, N4458, N947, N1290, N2272);
nor NOR4 (N4469, N4463, N648, N2587, N3401);
and AND3 (N4470, N4465, N1307, N2703);
nand NAND3 (N4471, N4455, N2351, N2895);
buf BUF1 (N4472, N4471);
nor NOR3 (N4473, N4464, N3110, N1243);
and AND3 (N4474, N4456, N4372, N3877);
nand NAND2 (N4475, N4466, N1174);
or OR4 (N4476, N4469, N3596, N2596, N2276);
nand NAND2 (N4477, N4473, N4438);
buf BUF1 (N4478, N4470);
xor XOR2 (N4479, N4477, N2057);
not NOT1 (N4480, N4474);
nand NAND2 (N4481, N4472, N2599);
xor XOR2 (N4482, N4480, N1770);
nor NOR2 (N4483, N4468, N1157);
buf BUF1 (N4484, N4481);
and AND2 (N4485, N4478, N2515);
buf BUF1 (N4486, N4482);
and AND3 (N4487, N4467, N1321, N462);
not NOT1 (N4488, N4485);
or OR4 (N4489, N4484, N2665, N2650, N4399);
xor XOR2 (N4490, N4483, N162);
nand NAND2 (N4491, N4488, N4339);
nor NOR3 (N4492, N4489, N4331, N998);
xor XOR2 (N4493, N4476, N1773);
not NOT1 (N4494, N4492);
nand NAND2 (N4495, N4494, N558);
not NOT1 (N4496, N4490);
nand NAND4 (N4497, N4491, N4311, N2765, N1892);
buf BUF1 (N4498, N4493);
not NOT1 (N4499, N4498);
xor XOR2 (N4500, N4495, N1041);
and AND3 (N4501, N4496, N39, N2558);
or OR3 (N4502, N4479, N3392, N1825);
nor NOR3 (N4503, N4475, N2100, N1170);
or OR3 (N4504, N4487, N1765, N4294);
not NOT1 (N4505, N4499);
or OR4 (N4506, N4462, N2453, N4351, N3295);
nor NOR4 (N4507, N4504, N2463, N2145, N3231);
and AND2 (N4508, N4501, N4137);
not NOT1 (N4509, N4497);
not NOT1 (N4510, N4449);
nand NAND4 (N4511, N4507, N1677, N1597, N345);
or OR2 (N4512, N4500, N4472);
and AND3 (N4513, N4502, N421, N3075);
xor XOR2 (N4514, N4512, N1122);
or OR2 (N4515, N4508, N4057);
xor XOR2 (N4516, N4510, N1665);
nand NAND4 (N4517, N4509, N567, N1386, N3094);
xor XOR2 (N4518, N4517, N2872);
and AND3 (N4519, N4516, N1813, N2790);
nor NOR4 (N4520, N4486, N2139, N3397, N4303);
buf BUF1 (N4521, N4503);
and AND2 (N4522, N4514, N687);
and AND4 (N4523, N4522, N252, N999, N3875);
xor XOR2 (N4524, N4518, N972);
xor XOR2 (N4525, N4520, N2324);
xor XOR2 (N4526, N4506, N1949);
xor XOR2 (N4527, N4524, N642);
or OR4 (N4528, N4523, N4506, N1980, N4413);
and AND4 (N4529, N4519, N1730, N3798, N1031);
or OR2 (N4530, N4515, N2447);
nand NAND2 (N4531, N4505, N3200);
xor XOR2 (N4532, N4527, N1737);
or OR2 (N4533, N4525, N4099);
and AND4 (N4534, N4533, N4423, N3830, N3394);
buf BUF1 (N4535, N4534);
nand NAND3 (N4536, N4526, N1673, N3904);
not NOT1 (N4537, N4535);
xor XOR2 (N4538, N4513, N395);
nor NOR4 (N4539, N4531, N2398, N292, N3914);
xor XOR2 (N4540, N4538, N1237);
or OR2 (N4541, N4532, N3053);
nand NAND4 (N4542, N4528, N1877, N3762, N3361);
not NOT1 (N4543, N4530);
buf BUF1 (N4544, N4540);
not NOT1 (N4545, N4537);
nor NOR4 (N4546, N4521, N1407, N2989, N1270);
or OR2 (N4547, N4511, N2071);
xor XOR2 (N4548, N4546, N3462);
or OR4 (N4549, N4543, N3756, N3716, N732);
and AND4 (N4550, N4545, N1720, N4303, N177);
buf BUF1 (N4551, N4547);
xor XOR2 (N4552, N4529, N1724);
nand NAND2 (N4553, N4551, N4040);
or OR2 (N4554, N4544, N475);
and AND4 (N4555, N4553, N4514, N4398, N4367);
or OR4 (N4556, N4555, N3508, N117, N1205);
buf BUF1 (N4557, N4541);
nand NAND4 (N4558, N4542, N2561, N73, N486);
or OR4 (N4559, N4552, N2563, N723, N712);
nand NAND3 (N4560, N4558, N331, N3520);
buf BUF1 (N4561, N4560);
xor XOR2 (N4562, N4556, N1895);
or OR4 (N4563, N4557, N4086, N3863, N2450);
and AND3 (N4564, N4548, N186, N3227);
buf BUF1 (N4565, N4536);
xor XOR2 (N4566, N4559, N2893);
nand NAND4 (N4567, N4565, N1083, N1471, N3315);
nand NAND4 (N4568, N4554, N4042, N2675, N2927);
or OR3 (N4569, N4562, N868, N2893);
nand NAND4 (N4570, N4566, N1941, N2928, N3451);
nand NAND4 (N4571, N4569, N4175, N2403, N451);
or OR4 (N4572, N4549, N428, N4462, N2208);
and AND3 (N4573, N4567, N763, N1926);
not NOT1 (N4574, N4539);
nor NOR4 (N4575, N4568, N3747, N749, N476);
buf BUF1 (N4576, N4573);
or OR4 (N4577, N4571, N3491, N237, N2161);
nor NOR2 (N4578, N4574, N1134);
not NOT1 (N4579, N4561);
and AND2 (N4580, N4550, N2311);
nor NOR3 (N4581, N4579, N2356, N3549);
not NOT1 (N4582, N4578);
nand NAND3 (N4583, N4563, N3863, N3564);
xor XOR2 (N4584, N4583, N1953);
buf BUF1 (N4585, N4576);
and AND2 (N4586, N4564, N3018);
nand NAND3 (N4587, N4570, N2462, N1069);
and AND4 (N4588, N4580, N4226, N570, N1572);
not NOT1 (N4589, N4585);
nor NOR2 (N4590, N4575, N237);
buf BUF1 (N4591, N4581);
or OR2 (N4592, N4588, N2076);
not NOT1 (N4593, N4589);
buf BUF1 (N4594, N4590);
xor XOR2 (N4595, N4594, N3793);
buf BUF1 (N4596, N4593);
xor XOR2 (N4597, N4584, N3086);
nand NAND3 (N4598, N4595, N1097, N1604);
not NOT1 (N4599, N4591);
nor NOR2 (N4600, N4577, N1222);
xor XOR2 (N4601, N4598, N3034);
xor XOR2 (N4602, N4596, N3762);
nand NAND4 (N4603, N4600, N2007, N3690, N985);
and AND4 (N4604, N4603, N505, N3933, N2480);
buf BUF1 (N4605, N4601);
nor NOR3 (N4606, N4605, N1266, N1037);
xor XOR2 (N4607, N4606, N3627);
buf BUF1 (N4608, N4586);
buf BUF1 (N4609, N4607);
buf BUF1 (N4610, N4599);
nor NOR3 (N4611, N4592, N1741, N2822);
nand NAND3 (N4612, N4611, N4238, N2802);
nor NOR2 (N4613, N4612, N406);
buf BUF1 (N4614, N4608);
not NOT1 (N4615, N4597);
not NOT1 (N4616, N4587);
buf BUF1 (N4617, N4610);
xor XOR2 (N4618, N4572, N2214);
nand NAND4 (N4619, N4618, N1249, N2329, N2416);
nand NAND4 (N4620, N4619, N2650, N4525, N1986);
nand NAND2 (N4621, N4609, N4094);
buf BUF1 (N4622, N4616);
or OR4 (N4623, N4602, N8, N2091, N69);
buf BUF1 (N4624, N4613);
and AND3 (N4625, N4621, N3062, N1063);
buf BUF1 (N4626, N4624);
xor XOR2 (N4627, N4615, N1533);
and AND3 (N4628, N4622, N1685, N1532);
xor XOR2 (N4629, N4627, N3509);
and AND3 (N4630, N4614, N3273, N1295);
nor NOR3 (N4631, N4625, N943, N2722);
buf BUF1 (N4632, N4630);
buf BUF1 (N4633, N4632);
nand NAND4 (N4634, N4626, N4274, N2379, N3875);
xor XOR2 (N4635, N4617, N4379);
buf BUF1 (N4636, N4628);
or OR2 (N4637, N4623, N653);
xor XOR2 (N4638, N4620, N9);
buf BUF1 (N4639, N4582);
nor NOR3 (N4640, N4634, N4005, N2142);
and AND4 (N4641, N4638, N4472, N3143, N3240);
and AND3 (N4642, N4635, N1334, N1604);
nand NAND2 (N4643, N4642, N2503);
not NOT1 (N4644, N4633);
buf BUF1 (N4645, N4644);
not NOT1 (N4646, N4641);
not NOT1 (N4647, N4645);
not NOT1 (N4648, N4629);
or OR4 (N4649, N4647, N2926, N4462, N2753);
xor XOR2 (N4650, N4640, N3288);
or OR2 (N4651, N4631, N3587);
not NOT1 (N4652, N4651);
xor XOR2 (N4653, N4636, N893);
buf BUF1 (N4654, N4639);
and AND3 (N4655, N4649, N2988, N4523);
nand NAND2 (N4656, N4604, N3451);
xor XOR2 (N4657, N4637, N3878);
or OR2 (N4658, N4650, N2769);
nor NOR2 (N4659, N4643, N2411);
buf BUF1 (N4660, N4654);
not NOT1 (N4661, N4648);
nand NAND2 (N4662, N4655, N1291);
or OR4 (N4663, N4656, N1902, N441, N2969);
xor XOR2 (N4664, N4653, N1246);
xor XOR2 (N4665, N4661, N4569);
and AND2 (N4666, N4646, N349);
not NOT1 (N4667, N4658);
or OR4 (N4668, N4659, N4184, N1069, N262);
buf BUF1 (N4669, N4665);
xor XOR2 (N4670, N4657, N217);
and AND3 (N4671, N4652, N457, N3521);
or OR4 (N4672, N4671, N2518, N2801, N1874);
nor NOR3 (N4673, N4664, N3313, N4342);
xor XOR2 (N4674, N4667, N3062);
nand NAND2 (N4675, N4660, N1084);
or OR4 (N4676, N4669, N1715, N3004, N3392);
xor XOR2 (N4677, N4662, N2283);
and AND3 (N4678, N4673, N3820, N2584);
xor XOR2 (N4679, N4663, N3075);
nor NOR4 (N4680, N4679, N2848, N173, N3435);
not NOT1 (N4681, N4666);
not NOT1 (N4682, N4670);
nand NAND4 (N4683, N4680, N2191, N2312, N1267);
buf BUF1 (N4684, N4672);
nand NAND2 (N4685, N4682, N2272);
buf BUF1 (N4686, N4668);
not NOT1 (N4687, N4678);
not NOT1 (N4688, N4674);
or OR3 (N4689, N4685, N3159, N739);
buf BUF1 (N4690, N4686);
and AND2 (N4691, N4681, N2954);
and AND4 (N4692, N4677, N2763, N1011, N4190);
or OR2 (N4693, N4689, N411);
not NOT1 (N4694, N4683);
and AND2 (N4695, N4690, N419);
xor XOR2 (N4696, N4693, N3872);
not NOT1 (N4697, N4676);
nand NAND2 (N4698, N4694, N1334);
not NOT1 (N4699, N4695);
and AND2 (N4700, N4698, N2612);
nor NOR3 (N4701, N4691, N740, N1965);
nand NAND2 (N4702, N4675, N1127);
nand NAND4 (N4703, N4687, N97, N1059, N3168);
and AND4 (N4704, N4692, N1190, N4552, N2402);
nor NOR2 (N4705, N4684, N3968);
nor NOR3 (N4706, N4697, N4200, N4177);
xor XOR2 (N4707, N4699, N2107);
or OR4 (N4708, N4696, N1861, N1119, N147);
and AND4 (N4709, N4708, N2491, N3350, N741);
buf BUF1 (N4710, N4707);
nand NAND4 (N4711, N4701, N2072, N4545, N2673);
and AND2 (N4712, N4703, N4244);
buf BUF1 (N4713, N4706);
and AND2 (N4714, N4711, N1196);
or OR3 (N4715, N4700, N395, N4025);
buf BUF1 (N4716, N4714);
xor XOR2 (N4717, N4716, N2836);
nand NAND3 (N4718, N4702, N1459, N3919);
buf BUF1 (N4719, N4688);
nor NOR2 (N4720, N4719, N3421);
and AND3 (N4721, N4713, N3055, N1822);
buf BUF1 (N4722, N4721);
not NOT1 (N4723, N4718);
xor XOR2 (N4724, N4715, N3716);
buf BUF1 (N4725, N4704);
buf BUF1 (N4726, N4723);
xor XOR2 (N4727, N4722, N4265);
nand NAND2 (N4728, N4710, N380);
nand NAND2 (N4729, N4720, N2707);
nor NOR3 (N4730, N4717, N4440, N3834);
nor NOR2 (N4731, N4712, N4719);
and AND3 (N4732, N4730, N1598, N4196);
nand NAND2 (N4733, N4725, N1406);
or OR3 (N4734, N4732, N2992, N541);
nand NAND2 (N4735, N4734, N2474);
xor XOR2 (N4736, N4733, N353);
and AND3 (N4737, N4726, N4469, N437);
xor XOR2 (N4738, N4705, N605);
not NOT1 (N4739, N4731);
or OR2 (N4740, N4737, N3137);
and AND3 (N4741, N4724, N3784, N3286);
not NOT1 (N4742, N4735);
not NOT1 (N4743, N4728);
and AND2 (N4744, N4739, N2144);
not NOT1 (N4745, N4727);
nand NAND4 (N4746, N4729, N3610, N3908, N4202);
or OR2 (N4747, N4744, N3573);
xor XOR2 (N4748, N4736, N3477);
nor NOR2 (N4749, N4745, N3834);
nand NAND2 (N4750, N4743, N951);
and AND2 (N4751, N4748, N2049);
and AND3 (N4752, N4751, N312, N3467);
and AND4 (N4753, N4746, N2334, N4550, N838);
nand NAND4 (N4754, N4741, N1593, N4219, N3856);
or OR2 (N4755, N4752, N1472);
nand NAND3 (N4756, N4738, N918, N1911);
not NOT1 (N4757, N4754);
buf BUF1 (N4758, N4747);
not NOT1 (N4759, N4757);
xor XOR2 (N4760, N4740, N4568);
or OR3 (N4761, N4756, N4045, N3806);
and AND4 (N4762, N4742, N1123, N4745, N3838);
nor NOR2 (N4763, N4753, N4303);
buf BUF1 (N4764, N4758);
not NOT1 (N4765, N4764);
nand NAND3 (N4766, N4762, N3126, N4726);
or OR2 (N4767, N4765, N2486);
or OR4 (N4768, N4761, N1220, N2299, N3776);
or OR3 (N4769, N4759, N1244, N2646);
xor XOR2 (N4770, N4750, N4283);
buf BUF1 (N4771, N4709);
nand NAND3 (N4772, N4749, N4109, N2088);
or OR3 (N4773, N4772, N4144, N3774);
xor XOR2 (N4774, N4773, N2363);
buf BUF1 (N4775, N4763);
xor XOR2 (N4776, N4755, N1932);
or OR3 (N4777, N4767, N2751, N4614);
nor NOR4 (N4778, N4760, N2981, N1726, N1718);
nand NAND4 (N4779, N4776, N249, N1754, N3680);
and AND2 (N4780, N4769, N1033);
not NOT1 (N4781, N4774);
or OR3 (N4782, N4766, N1328, N1603);
nand NAND3 (N4783, N4775, N1638, N2284);
nor NOR3 (N4784, N4780, N994, N949);
not NOT1 (N4785, N4782);
xor XOR2 (N4786, N4784, N3896);
and AND4 (N4787, N4778, N2506, N4172, N3468);
buf BUF1 (N4788, N4771);
xor XOR2 (N4789, N4770, N3294);
buf BUF1 (N4790, N4786);
and AND3 (N4791, N4781, N184, N1080);
nor NOR4 (N4792, N4783, N527, N3212, N1974);
buf BUF1 (N4793, N4787);
buf BUF1 (N4794, N4768);
nor NOR4 (N4795, N4794, N3026, N4582, N4539);
nand NAND3 (N4796, N4789, N1676, N823);
nor NOR2 (N4797, N4793, N2965);
nand NAND3 (N4798, N4796, N4151, N326);
nand NAND4 (N4799, N4779, N2497, N4349, N207);
xor XOR2 (N4800, N4788, N1348);
and AND2 (N4801, N4785, N601);
buf BUF1 (N4802, N4790);
not NOT1 (N4803, N4791);
xor XOR2 (N4804, N4798, N251);
and AND3 (N4805, N4797, N1902, N494);
or OR3 (N4806, N4792, N2410, N1287);
xor XOR2 (N4807, N4802, N4597);
xor XOR2 (N4808, N4777, N2525);
or OR3 (N4809, N4805, N1384, N3539);
xor XOR2 (N4810, N4807, N105);
or OR2 (N4811, N4795, N803);
or OR3 (N4812, N4808, N284, N3600);
not NOT1 (N4813, N4810);
xor XOR2 (N4814, N4812, N1506);
not NOT1 (N4815, N4806);
nand NAND2 (N4816, N4811, N1331);
buf BUF1 (N4817, N4809);
and AND2 (N4818, N4804, N2800);
and AND3 (N4819, N4800, N1915, N449);
and AND3 (N4820, N4818, N1463, N3255);
buf BUF1 (N4821, N4803);
nand NAND2 (N4822, N4815, N3254);
and AND2 (N4823, N4820, N3037);
nor NOR2 (N4824, N4819, N748);
nand NAND2 (N4825, N4823, N3413);
buf BUF1 (N4826, N4813);
nand NAND4 (N4827, N4826, N406, N3644, N1053);
buf BUF1 (N4828, N4824);
or OR3 (N4829, N4821, N2468, N4066);
nor NOR3 (N4830, N4828, N530, N4375);
or OR4 (N4831, N4827, N3052, N2880, N1614);
nor NOR2 (N4832, N4814, N4042);
buf BUF1 (N4833, N4817);
xor XOR2 (N4834, N4816, N489);
xor XOR2 (N4835, N4833, N878);
or OR4 (N4836, N4799, N754, N1197, N4728);
not NOT1 (N4837, N4829);
or OR3 (N4838, N4830, N4650, N1342);
and AND4 (N4839, N4822, N1750, N4613, N3122);
nor NOR2 (N4840, N4832, N1099);
nor NOR2 (N4841, N4834, N3651);
and AND3 (N4842, N4836, N3173, N3219);
xor XOR2 (N4843, N4831, N3274);
nand NAND2 (N4844, N4835, N3850);
nor NOR2 (N4845, N4801, N3253);
nand NAND2 (N4846, N4825, N410);
nand NAND3 (N4847, N4838, N4172, N942);
not NOT1 (N4848, N4846);
nor NOR4 (N4849, N4847, N3458, N4565, N2965);
or OR4 (N4850, N4841, N2369, N4468, N1395);
buf BUF1 (N4851, N4849);
nor NOR3 (N4852, N4837, N2961, N2419);
and AND3 (N4853, N4851, N4517, N325);
xor XOR2 (N4854, N4844, N2542);
nand NAND2 (N4855, N4848, N4205);
or OR3 (N4856, N4839, N2240, N575);
not NOT1 (N4857, N4842);
nor NOR3 (N4858, N4856, N3342, N2078);
xor XOR2 (N4859, N4857, N4856);
nand NAND4 (N4860, N4850, N2050, N136, N3546);
not NOT1 (N4861, N4853);
buf BUF1 (N4862, N4858);
not NOT1 (N4863, N4855);
not NOT1 (N4864, N4854);
not NOT1 (N4865, N4860);
not NOT1 (N4866, N4861);
nand NAND4 (N4867, N4864, N4702, N3958, N876);
nor NOR3 (N4868, N4862, N1137, N3331);
or OR2 (N4869, N4840, N2662);
not NOT1 (N4870, N4867);
nand NAND2 (N4871, N4869, N2769);
nand NAND4 (N4872, N4868, N4854, N2436, N2515);
xor XOR2 (N4873, N4872, N2968);
xor XOR2 (N4874, N4871, N3392);
xor XOR2 (N4875, N4859, N4750);
nor NOR3 (N4876, N4866, N1221, N2199);
xor XOR2 (N4877, N4865, N1705);
not NOT1 (N4878, N4873);
not NOT1 (N4879, N4878);
nor NOR2 (N4880, N4875, N1751);
xor XOR2 (N4881, N4880, N1284);
and AND4 (N4882, N4843, N3487, N3839, N1756);
buf BUF1 (N4883, N4852);
and AND4 (N4884, N4881, N2751, N4239, N3985);
not NOT1 (N4885, N4877);
buf BUF1 (N4886, N4874);
nand NAND4 (N4887, N4845, N3732, N3731, N3652);
and AND3 (N4888, N4885, N1144, N1727);
not NOT1 (N4889, N4886);
nor NOR3 (N4890, N4876, N3801, N2989);
nor NOR4 (N4891, N4889, N4000, N1326, N1974);
xor XOR2 (N4892, N4888, N2567);
xor XOR2 (N4893, N4884, N174);
not NOT1 (N4894, N4883);
nand NAND3 (N4895, N4882, N15, N2898);
xor XOR2 (N4896, N4887, N382);
nand NAND2 (N4897, N4894, N4232);
buf BUF1 (N4898, N4893);
and AND3 (N4899, N4892, N3073, N1777);
buf BUF1 (N4900, N4899);
and AND4 (N4901, N4895, N2632, N4475, N117);
and AND4 (N4902, N4901, N2691, N2861, N1855);
buf BUF1 (N4903, N4870);
nand NAND4 (N4904, N4890, N4634, N761, N3155);
xor XOR2 (N4905, N4904, N3365);
buf BUF1 (N4906, N4897);
or OR4 (N4907, N4879, N4243, N432, N4593);
nor NOR3 (N4908, N4906, N3906, N2175);
or OR3 (N4909, N4905, N1595, N3400);
nor NOR3 (N4910, N4903, N4186, N1695);
xor XOR2 (N4911, N4907, N2531);
nand NAND2 (N4912, N4910, N4372);
not NOT1 (N4913, N4909);
not NOT1 (N4914, N4891);
and AND3 (N4915, N4914, N4793, N1518);
nand NAND4 (N4916, N4898, N1096, N1868, N4264);
not NOT1 (N4917, N4908);
nor NOR2 (N4918, N4917, N219);
or OR2 (N4919, N4918, N2491);
xor XOR2 (N4920, N4900, N1316);
nand NAND4 (N4921, N4912, N1500, N2179, N1403);
xor XOR2 (N4922, N4913, N755);
not NOT1 (N4923, N4863);
not NOT1 (N4924, N4916);
buf BUF1 (N4925, N4922);
nor NOR2 (N4926, N4924, N888);
or OR4 (N4927, N4923, N4580, N2879, N963);
or OR4 (N4928, N4920, N3278, N3074, N2878);
not NOT1 (N4929, N4896);
xor XOR2 (N4930, N4919, N39);
not NOT1 (N4931, N4929);
or OR4 (N4932, N4928, N2052, N2527, N1260);
buf BUF1 (N4933, N4931);
xor XOR2 (N4934, N4921, N3123);
nand NAND4 (N4935, N4932, N2508, N2266, N3255);
xor XOR2 (N4936, N4935, N3918);
not NOT1 (N4937, N4934);
not NOT1 (N4938, N4925);
nand NAND4 (N4939, N4936, N274, N4145, N3201);
or OR3 (N4940, N4937, N457, N3376);
not NOT1 (N4941, N4911);
xor XOR2 (N4942, N4939, N1871);
nand NAND2 (N4943, N4930, N4872);
not NOT1 (N4944, N4940);
and AND4 (N4945, N4944, N1506, N1391, N2382);
xor XOR2 (N4946, N4945, N385);
xor XOR2 (N4947, N4938, N1091);
and AND3 (N4948, N4933, N34, N2505);
not NOT1 (N4949, N4902);
buf BUF1 (N4950, N4946);
buf BUF1 (N4951, N4949);
xor XOR2 (N4952, N4941, N4618);
or OR2 (N4953, N4952, N1449);
or OR2 (N4954, N4950, N3905);
not NOT1 (N4955, N4926);
or OR3 (N4956, N4943, N4099, N4819);
or OR3 (N4957, N4915, N4035, N4114);
and AND2 (N4958, N4957, N1237);
nor NOR3 (N4959, N4942, N1923, N2733);
buf BUF1 (N4960, N4947);
not NOT1 (N4961, N4948);
and AND3 (N4962, N4955, N3112, N2713);
nor NOR2 (N4963, N4954, N3654);
xor XOR2 (N4964, N4953, N2304);
xor XOR2 (N4965, N4927, N2152);
or OR2 (N4966, N4959, N3284);
nand NAND4 (N4967, N4964, N2261, N3585, N4687);
and AND2 (N4968, N4951, N2675);
nor NOR4 (N4969, N4968, N3157, N4193, N4363);
nand NAND3 (N4970, N4963, N3407, N3633);
not NOT1 (N4971, N4961);
xor XOR2 (N4972, N4969, N379);
nor NOR3 (N4973, N4960, N4561, N2901);
or OR4 (N4974, N4956, N4621, N2234, N3639);
nor NOR3 (N4975, N4962, N943, N1405);
not NOT1 (N4976, N4972);
nor NOR3 (N4977, N4965, N946, N2843);
xor XOR2 (N4978, N4977, N1149);
nor NOR3 (N4979, N4966, N3275, N1795);
and AND3 (N4980, N4967, N3534, N4624);
nor NOR2 (N4981, N4973, N4704);
and AND4 (N4982, N4970, N3820, N2837, N953);
xor XOR2 (N4983, N4976, N2008);
xor XOR2 (N4984, N4974, N2705);
and AND2 (N4985, N4978, N1723);
buf BUF1 (N4986, N4984);
not NOT1 (N4987, N4975);
not NOT1 (N4988, N4980);
nor NOR4 (N4989, N4985, N2976, N2661, N1837);
and AND2 (N4990, N4958, N3339);
not NOT1 (N4991, N4989);
xor XOR2 (N4992, N4983, N1259);
not NOT1 (N4993, N4981);
nor NOR3 (N4994, N4992, N3570, N632);
not NOT1 (N4995, N4987);
xor XOR2 (N4996, N4979, N214);
and AND2 (N4997, N4982, N3300);
and AND3 (N4998, N4994, N4001, N2823);
or OR3 (N4999, N4998, N4019, N2195);
and AND2 (N5000, N4986, N4573);
or OR4 (N5001, N5000, N570, N2165, N3012);
buf BUF1 (N5002, N4993);
nand NAND3 (N5003, N4991, N2627, N4694);
and AND3 (N5004, N5001, N2002, N4339);
xor XOR2 (N5005, N4988, N739);
and AND2 (N5006, N4997, N4749);
not NOT1 (N5007, N5003);
buf BUF1 (N5008, N4990);
xor XOR2 (N5009, N4995, N2354);
buf BUF1 (N5010, N5005);
not NOT1 (N5011, N4996);
xor XOR2 (N5012, N5007, N365);
buf BUF1 (N5013, N4999);
not NOT1 (N5014, N5008);
and AND4 (N5015, N5004, N2056, N4372, N4308);
nor NOR2 (N5016, N5014, N4012);
or OR3 (N5017, N5009, N2159, N717);
and AND4 (N5018, N5006, N348, N1103, N2199);
nor NOR3 (N5019, N5018, N1723, N4060);
or OR2 (N5020, N5012, N4720);
not NOT1 (N5021, N5011);
or OR4 (N5022, N5010, N196, N487, N3881);
nand NAND2 (N5023, N5015, N4318);
nor NOR4 (N5024, N5002, N1629, N2286, N216);
nand NAND2 (N5025, N4971, N3747);
not NOT1 (N5026, N5019);
xor XOR2 (N5027, N5017, N1829);
or OR3 (N5028, N5025, N3843, N4983);
and AND3 (N5029, N5022, N4495, N301);
buf BUF1 (N5030, N5021);
nor NOR3 (N5031, N5028, N736, N2470);
nor NOR2 (N5032, N5023, N1049);
or OR3 (N5033, N5026, N1105, N4268);
and AND3 (N5034, N5016, N3569, N3337);
buf BUF1 (N5035, N5020);
and AND3 (N5036, N5031, N101, N2665);
not NOT1 (N5037, N5034);
xor XOR2 (N5038, N5032, N2757);
not NOT1 (N5039, N5033);
nor NOR3 (N5040, N5037, N3400, N2677);
nor NOR4 (N5041, N5029, N1948, N1940, N775);
nor NOR3 (N5042, N5024, N2701, N1224);
and AND2 (N5043, N5035, N1959);
xor XOR2 (N5044, N5036, N4856);
not NOT1 (N5045, N5040);
or OR4 (N5046, N5027, N2623, N261, N4806);
buf BUF1 (N5047, N5046);
or OR3 (N5048, N5039, N1951, N4996);
nand NAND2 (N5049, N5045, N2926);
nand NAND2 (N5050, N5043, N1676);
or OR4 (N5051, N5038, N3263, N4596, N664);
xor XOR2 (N5052, N5051, N3712);
or OR2 (N5053, N5050, N598);
nand NAND3 (N5054, N5041, N1340, N3092);
and AND4 (N5055, N5044, N2096, N1923, N992);
nor NOR2 (N5056, N5047, N2249);
nand NAND3 (N5057, N5053, N3334, N778);
not NOT1 (N5058, N5048);
and AND3 (N5059, N5013, N4913, N1947);
buf BUF1 (N5060, N5056);
nor NOR4 (N5061, N5055, N5060, N2566, N656);
nor NOR3 (N5062, N3251, N3433, N1898);
buf BUF1 (N5063, N5054);
xor XOR2 (N5064, N5057, N2947);
not NOT1 (N5065, N5059);
nand NAND3 (N5066, N5058, N383, N2245);
buf BUF1 (N5067, N5030);
nor NOR3 (N5068, N5063, N1342, N1139);
nand NAND4 (N5069, N5068, N2005, N3391, N1829);
and AND2 (N5070, N5052, N3222);
xor XOR2 (N5071, N5065, N3582);
not NOT1 (N5072, N5061);
buf BUF1 (N5073, N5072);
buf BUF1 (N5074, N5062);
and AND2 (N5075, N5049, N1311);
buf BUF1 (N5076, N5073);
or OR2 (N5077, N5069, N1906);
xor XOR2 (N5078, N5075, N174);
xor XOR2 (N5079, N5070, N2026);
buf BUF1 (N5080, N5064);
and AND4 (N5081, N5076, N3911, N534, N1683);
nand NAND2 (N5082, N5077, N824);
nand NAND4 (N5083, N5042, N950, N1011, N4900);
not NOT1 (N5084, N5071);
xor XOR2 (N5085, N5084, N2823);
xor XOR2 (N5086, N5066, N2791);
xor XOR2 (N5087, N5085, N3880);
nor NOR4 (N5088, N5079, N3626, N1046, N2324);
and AND2 (N5089, N5080, N1661);
not NOT1 (N5090, N5083);
nand NAND4 (N5091, N5078, N2501, N3662, N2663);
xor XOR2 (N5092, N5088, N901);
nor NOR4 (N5093, N5089, N1079, N4123, N2569);
nor NOR4 (N5094, N5087, N2203, N3400, N4679);
and AND3 (N5095, N5086, N4792, N3097);
nor NOR2 (N5096, N5082, N4229);
and AND4 (N5097, N5093, N4771, N1777, N4021);
or OR3 (N5098, N5097, N4917, N4326);
and AND2 (N5099, N5095, N3058);
nor NOR2 (N5100, N5090, N3636);
or OR2 (N5101, N5094, N3224);
nand NAND4 (N5102, N5092, N3115, N4898, N2519);
buf BUF1 (N5103, N5074);
not NOT1 (N5104, N5102);
nand NAND2 (N5105, N5081, N4283);
not NOT1 (N5106, N5099);
buf BUF1 (N5107, N5098);
and AND3 (N5108, N5103, N2631, N3083);
buf BUF1 (N5109, N5105);
or OR3 (N5110, N5101, N3620, N2962);
nand NAND4 (N5111, N5109, N333, N4850, N1339);
nor NOR2 (N5112, N5100, N2949);
nor NOR2 (N5113, N5067, N753);
buf BUF1 (N5114, N5107);
nor NOR3 (N5115, N5114, N1512, N3785);
buf BUF1 (N5116, N5112);
xor XOR2 (N5117, N5096, N3348);
xor XOR2 (N5118, N5108, N3286);
not NOT1 (N5119, N5111);
nand NAND3 (N5120, N5106, N487, N2240);
nand NAND3 (N5121, N5116, N1896, N2249);
and AND2 (N5122, N5104, N1386);
buf BUF1 (N5123, N5091);
or OR4 (N5124, N5117, N2141, N2656, N1853);
buf BUF1 (N5125, N5118);
buf BUF1 (N5126, N5125);
or OR3 (N5127, N5115, N1016, N3877);
and AND4 (N5128, N5113, N2499, N3421, N2507);
xor XOR2 (N5129, N5126, N2687);
buf BUF1 (N5130, N5110);
or OR4 (N5131, N5121, N2899, N4149, N1050);
nand NAND3 (N5132, N5123, N4399, N3038);
xor XOR2 (N5133, N5120, N3975);
or OR4 (N5134, N5119, N142, N1295, N2456);
buf BUF1 (N5135, N5128);
nor NOR4 (N5136, N5133, N279, N4329, N1500);
nor NOR3 (N5137, N5127, N2428, N4274);
or OR3 (N5138, N5131, N130, N144);
xor XOR2 (N5139, N5138, N2717);
xor XOR2 (N5140, N5132, N273);
buf BUF1 (N5141, N5122);
or OR3 (N5142, N5141, N137, N1572);
and AND4 (N5143, N5129, N286, N2659, N4913);
or OR3 (N5144, N5137, N2612, N2604);
nor NOR2 (N5145, N5143, N68);
or OR2 (N5146, N5144, N2227);
xor XOR2 (N5147, N5134, N2532);
nor NOR3 (N5148, N5146, N5042, N2850);
nor NOR4 (N5149, N5140, N2777, N1784, N4935);
xor XOR2 (N5150, N5147, N4688);
nor NOR3 (N5151, N5142, N2312, N4118);
xor XOR2 (N5152, N5149, N465);
and AND2 (N5153, N5151, N4321);
nor NOR2 (N5154, N5148, N2521);
buf BUF1 (N5155, N5150);
buf BUF1 (N5156, N5145);
not NOT1 (N5157, N5136);
or OR2 (N5158, N5153, N588);
buf BUF1 (N5159, N5157);
xor XOR2 (N5160, N5155, N847);
nor NOR2 (N5161, N5152, N2202);
not NOT1 (N5162, N5130);
and AND4 (N5163, N5159, N1128, N750, N3902);
nand NAND3 (N5164, N5135, N1000, N3309);
or OR4 (N5165, N5139, N2294, N1435, N4600);
xor XOR2 (N5166, N5156, N4208);
nand NAND2 (N5167, N5164, N297);
nor NOR2 (N5168, N5165, N4382);
or OR3 (N5169, N5166, N4684, N751);
buf BUF1 (N5170, N5162);
or OR2 (N5171, N5161, N2477);
xor XOR2 (N5172, N5169, N2714);
buf BUF1 (N5173, N5171);
not NOT1 (N5174, N5168);
and AND4 (N5175, N5167, N4164, N2491, N3851);
xor XOR2 (N5176, N5124, N2843);
and AND2 (N5177, N5176, N3547);
or OR2 (N5178, N5177, N3059);
nor NOR3 (N5179, N5158, N4496, N3239);
nand NAND2 (N5180, N5172, N418);
nor NOR4 (N5181, N5174, N3720, N4174, N5125);
nor NOR2 (N5182, N5163, N2532);
xor XOR2 (N5183, N5181, N1920);
xor XOR2 (N5184, N5179, N271);
or OR3 (N5185, N5180, N3073, N3166);
and AND2 (N5186, N5182, N672);
nand NAND2 (N5187, N5186, N4267);
nand NAND3 (N5188, N5173, N4817, N967);
nand NAND3 (N5189, N5178, N4197, N715);
nor NOR4 (N5190, N5188, N4202, N3471, N1244);
not NOT1 (N5191, N5184);
nand NAND2 (N5192, N5183, N4567);
nor NOR4 (N5193, N5192, N2838, N3031, N4862);
nand NAND4 (N5194, N5185, N4051, N3396, N3061);
buf BUF1 (N5195, N5190);
nand NAND4 (N5196, N5154, N3928, N284, N487);
nor NOR4 (N5197, N5160, N4374, N3241, N1682);
nor NOR3 (N5198, N5175, N961, N3198);
not NOT1 (N5199, N5193);
buf BUF1 (N5200, N5198);
buf BUF1 (N5201, N5189);
and AND4 (N5202, N5191, N4904, N4499, N3281);
xor XOR2 (N5203, N5170, N5056);
nor NOR4 (N5204, N5195, N2542, N2145, N3254);
buf BUF1 (N5205, N5187);
or OR3 (N5206, N5203, N3084, N2062);
xor XOR2 (N5207, N5202, N4412);
nor NOR3 (N5208, N5206, N3722, N3727);
or OR4 (N5209, N5197, N1939, N953, N2837);
buf BUF1 (N5210, N5200);
not NOT1 (N5211, N5207);
nand NAND2 (N5212, N5194, N679);
or OR2 (N5213, N5211, N4783);
not NOT1 (N5214, N5204);
xor XOR2 (N5215, N5208, N2326);
not NOT1 (N5216, N5214);
xor XOR2 (N5217, N5210, N4828);
nor NOR3 (N5218, N5196, N4396, N3267);
nand NAND4 (N5219, N5213, N3715, N2948, N2037);
and AND3 (N5220, N5199, N2930, N3647);
buf BUF1 (N5221, N5220);
and AND3 (N5222, N5219, N4608, N4402);
not NOT1 (N5223, N5218);
and AND2 (N5224, N5221, N4076);
not NOT1 (N5225, N5205);
and AND4 (N5226, N5216, N2622, N3174, N1361);
xor XOR2 (N5227, N5222, N4258);
xor XOR2 (N5228, N5209, N4817);
nand NAND4 (N5229, N5227, N1643, N2125, N1603);
and AND2 (N5230, N5212, N4234);
buf BUF1 (N5231, N5229);
nor NOR3 (N5232, N5201, N2854, N2181);
nand NAND4 (N5233, N5215, N14, N577, N1796);
buf BUF1 (N5234, N5233);
nand NAND2 (N5235, N5217, N1697);
nand NAND4 (N5236, N5231, N1956, N3202, N1521);
nand NAND2 (N5237, N5228, N2779);
xor XOR2 (N5238, N5224, N3904);
or OR2 (N5239, N5226, N4439);
nor NOR3 (N5240, N5234, N3104, N900);
nand NAND3 (N5241, N5232, N2280, N3516);
or OR4 (N5242, N5236, N5183, N656, N887);
and AND4 (N5243, N5241, N3788, N3461, N1628);
and AND2 (N5244, N5230, N1461);
buf BUF1 (N5245, N5237);
not NOT1 (N5246, N5243);
nand NAND2 (N5247, N5239, N800);
nor NOR3 (N5248, N5223, N2840, N1194);
or OR4 (N5249, N5238, N3537, N5162, N3569);
and AND2 (N5250, N5247, N4244);
not NOT1 (N5251, N5250);
nor NOR4 (N5252, N5242, N4926, N1507, N4195);
xor XOR2 (N5253, N5244, N3331);
xor XOR2 (N5254, N5248, N1684);
not NOT1 (N5255, N5235);
nor NOR2 (N5256, N5225, N3830);
or OR4 (N5257, N5253, N3439, N4279, N4102);
nand NAND2 (N5258, N5252, N4777);
nand NAND2 (N5259, N5255, N253);
not NOT1 (N5260, N5240);
nand NAND4 (N5261, N5246, N2475, N1934, N4914);
nor NOR3 (N5262, N5256, N3952, N2286);
nand NAND3 (N5263, N5260, N3936, N4776);
nand NAND2 (N5264, N5251, N1474);
nor NOR2 (N5265, N5254, N4617);
nand NAND2 (N5266, N5262, N800);
not NOT1 (N5267, N5261);
not NOT1 (N5268, N5249);
xor XOR2 (N5269, N5264, N361);
nand NAND2 (N5270, N5263, N2050);
buf BUF1 (N5271, N5258);
buf BUF1 (N5272, N5269);
not NOT1 (N5273, N5265);
not NOT1 (N5274, N5266);
or OR3 (N5275, N5267, N537, N310);
nand NAND3 (N5276, N5257, N1619, N3102);
or OR3 (N5277, N5272, N483, N4895);
nor NOR4 (N5278, N5245, N1568, N657, N1138);
buf BUF1 (N5279, N5277);
xor XOR2 (N5280, N5271, N2760);
or OR2 (N5281, N5276, N497);
or OR3 (N5282, N5259, N1294, N3288);
and AND2 (N5283, N5279, N4043);
or OR3 (N5284, N5282, N614, N5015);
xor XOR2 (N5285, N5284, N1278);
nand NAND4 (N5286, N5274, N3108, N2401, N2906);
nor NOR4 (N5287, N5278, N1378, N2825, N830);
nand NAND3 (N5288, N5273, N918, N2812);
not NOT1 (N5289, N5280);
buf BUF1 (N5290, N5283);
buf BUF1 (N5291, N5288);
xor XOR2 (N5292, N5275, N1970);
not NOT1 (N5293, N5289);
nand NAND4 (N5294, N5285, N1500, N2405, N3109);
nor NOR3 (N5295, N5286, N2540, N1285);
nor NOR4 (N5296, N5281, N4928, N399, N5214);
and AND3 (N5297, N5294, N2784, N3803);
or OR3 (N5298, N5290, N2442, N877);
buf BUF1 (N5299, N5296);
and AND3 (N5300, N5270, N3355, N5204);
nor NOR2 (N5301, N5297, N294);
and AND2 (N5302, N5301, N2920);
xor XOR2 (N5303, N5302, N3119);
not NOT1 (N5304, N5300);
nand NAND4 (N5305, N5291, N1364, N3133, N3957);
nand NAND4 (N5306, N5299, N3595, N898, N1224);
nand NAND4 (N5307, N5295, N1302, N946, N3766);
nor NOR3 (N5308, N5287, N1781, N1451);
xor XOR2 (N5309, N5298, N2722);
xor XOR2 (N5310, N5304, N380);
not NOT1 (N5311, N5309);
nand NAND3 (N5312, N5310, N5236, N868);
xor XOR2 (N5313, N5303, N1773);
nand NAND4 (N5314, N5311, N3259, N1261, N5302);
and AND3 (N5315, N5307, N3545, N2991);
xor XOR2 (N5316, N5293, N775);
nor NOR3 (N5317, N5292, N289, N2967);
xor XOR2 (N5318, N5315, N1015);
and AND2 (N5319, N5268, N4684);
nor NOR4 (N5320, N5318, N4766, N2504, N3128);
or OR3 (N5321, N5313, N1032, N931);
or OR4 (N5322, N5308, N2379, N3081, N4235);
buf BUF1 (N5323, N5317);
not NOT1 (N5324, N5323);
nor NOR4 (N5325, N5324, N1010, N4071, N3775);
nor NOR3 (N5326, N5316, N1836, N3593);
buf BUF1 (N5327, N5319);
not NOT1 (N5328, N5314);
xor XOR2 (N5329, N5305, N5212);
buf BUF1 (N5330, N5320);
xor XOR2 (N5331, N5312, N4778);
nor NOR2 (N5332, N5326, N1737);
not NOT1 (N5333, N5325);
or OR4 (N5334, N5322, N1127, N1233, N202);
not NOT1 (N5335, N5333);
nor NOR2 (N5336, N5329, N4398);
nor NOR4 (N5337, N5306, N3144, N1251, N3709);
xor XOR2 (N5338, N5331, N1000);
xor XOR2 (N5339, N5335, N4177);
nand NAND2 (N5340, N5338, N5064);
or OR2 (N5341, N5327, N4942);
or OR2 (N5342, N5336, N2136);
or OR4 (N5343, N5321, N3947, N3806, N4481);
and AND3 (N5344, N5341, N3303, N1805);
nand NAND4 (N5345, N5334, N559, N106, N3191);
nand NAND2 (N5346, N5332, N2990);
or OR4 (N5347, N5342, N5007, N14, N3067);
and AND4 (N5348, N5337, N94, N3090, N2633);
xor XOR2 (N5349, N5345, N2677);
or OR3 (N5350, N5346, N526, N2061);
not NOT1 (N5351, N5344);
buf BUF1 (N5352, N5339);
and AND4 (N5353, N5330, N103, N820, N1988);
or OR4 (N5354, N5350, N3089, N3796, N4229);
or OR4 (N5355, N5352, N2834, N4228, N4347);
buf BUF1 (N5356, N5328);
not NOT1 (N5357, N5351);
nand NAND4 (N5358, N5343, N4610, N2081, N2440);
buf BUF1 (N5359, N5347);
nor NOR3 (N5360, N5358, N2734, N779);
nand NAND4 (N5361, N5357, N2347, N3549, N5133);
not NOT1 (N5362, N5340);
buf BUF1 (N5363, N5362);
nor NOR2 (N5364, N5353, N2333);
nor NOR3 (N5365, N5355, N4376, N191);
nand NAND4 (N5366, N5359, N2409, N4840, N4291);
nor NOR3 (N5367, N5349, N1863, N4919);
not NOT1 (N5368, N5361);
buf BUF1 (N5369, N5367);
not NOT1 (N5370, N5363);
nor NOR2 (N5371, N5348, N1910);
xor XOR2 (N5372, N5356, N5072);
and AND2 (N5373, N5364, N1791);
nor NOR2 (N5374, N5366, N384);
buf BUF1 (N5375, N5373);
xor XOR2 (N5376, N5369, N2267);
and AND4 (N5377, N5360, N4150, N5318, N3556);
nand NAND3 (N5378, N5377, N5057, N2155);
xor XOR2 (N5379, N5372, N4660);
xor XOR2 (N5380, N5368, N400);
not NOT1 (N5381, N5374);
buf BUF1 (N5382, N5379);
nand NAND3 (N5383, N5382, N1350, N1368);
not NOT1 (N5384, N5383);
buf BUF1 (N5385, N5371);
buf BUF1 (N5386, N5376);
or OR4 (N5387, N5365, N4866, N2137, N2173);
buf BUF1 (N5388, N5385);
nand NAND3 (N5389, N5370, N5333, N5320);
nand NAND2 (N5390, N5386, N270);
buf BUF1 (N5391, N5390);
and AND4 (N5392, N5375, N2608, N5026, N1389);
nand NAND2 (N5393, N5388, N5321);
xor XOR2 (N5394, N5392, N1702);
and AND4 (N5395, N5354, N278, N164, N5099);
and AND3 (N5396, N5387, N1657, N1977);
nor NOR4 (N5397, N5391, N352, N5127, N201);
buf BUF1 (N5398, N5394);
nand NAND3 (N5399, N5381, N1524, N3687);
and AND2 (N5400, N5378, N3992);
buf BUF1 (N5401, N5380);
nor NOR2 (N5402, N5401, N4302);
nand NAND3 (N5403, N5395, N3957, N2661);
and AND4 (N5404, N5384, N1627, N3014, N3848);
nor NOR3 (N5405, N5403, N2699, N203);
nor NOR4 (N5406, N5404, N2004, N2565, N574);
xor XOR2 (N5407, N5406, N1875);
nand NAND2 (N5408, N5397, N1968);
buf BUF1 (N5409, N5396);
nor NOR4 (N5410, N5400, N4643, N1306, N1671);
not NOT1 (N5411, N5399);
nor NOR4 (N5412, N5389, N186, N4639, N4113);
and AND4 (N5413, N5398, N4539, N1410, N3857);
xor XOR2 (N5414, N5411, N5072);
nand NAND3 (N5415, N5405, N4454, N196);
and AND4 (N5416, N5393, N5284, N1174, N4207);
buf BUF1 (N5417, N5407);
and AND3 (N5418, N5413, N4871, N2016);
xor XOR2 (N5419, N5417, N1895);
buf BUF1 (N5420, N5412);
nand NAND2 (N5421, N5416, N2610);
xor XOR2 (N5422, N5414, N3468);
not NOT1 (N5423, N5409);
or OR4 (N5424, N5421, N3252, N2368, N4837);
and AND2 (N5425, N5419, N2762);
not NOT1 (N5426, N5420);
or OR4 (N5427, N5418, N3787, N1237, N2199);
nor NOR2 (N5428, N5425, N389);
buf BUF1 (N5429, N5402);
or OR2 (N5430, N5428, N1646);
or OR3 (N5431, N5429, N4964, N4922);
nand NAND2 (N5432, N5427, N4256);
and AND3 (N5433, N5423, N3244, N2127);
or OR4 (N5434, N5433, N369, N522, N633);
nor NOR3 (N5435, N5426, N1393, N2234);
xor XOR2 (N5436, N5435, N1104);
buf BUF1 (N5437, N5434);
or OR4 (N5438, N5410, N2972, N2298, N416);
and AND3 (N5439, N5436, N3370, N4548);
nor NOR3 (N5440, N5432, N4535, N2970);
nand NAND2 (N5441, N5424, N4711);
nor NOR4 (N5442, N5415, N4376, N1620, N2150);
xor XOR2 (N5443, N5442, N2309);
not NOT1 (N5444, N5422);
or OR3 (N5445, N5430, N415, N682);
nor NOR3 (N5446, N5443, N1441, N4077);
nand NAND2 (N5447, N5441, N5071);
xor XOR2 (N5448, N5438, N2269);
nor NOR4 (N5449, N5445, N1727, N2009, N2082);
not NOT1 (N5450, N5446);
xor XOR2 (N5451, N5439, N4408);
not NOT1 (N5452, N5449);
nor NOR3 (N5453, N5440, N4634, N536);
and AND3 (N5454, N5437, N1807, N351);
nand NAND2 (N5455, N5452, N1057);
nand NAND3 (N5456, N5455, N3886, N5349);
xor XOR2 (N5457, N5456, N141);
nand NAND3 (N5458, N5408, N2788, N796);
or OR2 (N5459, N5448, N1239);
nor NOR2 (N5460, N5453, N1932);
not NOT1 (N5461, N5458);
buf BUF1 (N5462, N5454);
buf BUF1 (N5463, N5462);
nand NAND2 (N5464, N5450, N3452);
buf BUF1 (N5465, N5460);
xor XOR2 (N5466, N5465, N1074);
nand NAND2 (N5467, N5466, N4125);
not NOT1 (N5468, N5457);
not NOT1 (N5469, N5463);
nand NAND3 (N5470, N5451, N1621, N1901);
xor XOR2 (N5471, N5468, N4739);
xor XOR2 (N5472, N5464, N1247);
nor NOR2 (N5473, N5447, N1054);
or OR2 (N5474, N5459, N5435);
xor XOR2 (N5475, N5431, N4218);
not NOT1 (N5476, N5472);
and AND2 (N5477, N5474, N2999);
or OR2 (N5478, N5469, N2059);
or OR4 (N5479, N5475, N2663, N794, N2811);
xor XOR2 (N5480, N5473, N3984);
nor NOR3 (N5481, N5444, N3153, N2835);
and AND4 (N5482, N5470, N3745, N1811, N4804);
and AND2 (N5483, N5480, N627);
xor XOR2 (N5484, N5471, N2557);
nor NOR2 (N5485, N5461, N2231);
nor NOR2 (N5486, N5476, N4122);
or OR2 (N5487, N5483, N585);
buf BUF1 (N5488, N5479);
and AND4 (N5489, N5477, N3231, N1520, N752);
or OR3 (N5490, N5487, N4860, N187);
not NOT1 (N5491, N5481);
or OR2 (N5492, N5478, N1846);
or OR3 (N5493, N5486, N1536, N4575);
or OR2 (N5494, N5493, N4120);
nor NOR2 (N5495, N5491, N4012);
and AND3 (N5496, N5485, N2919, N4392);
and AND2 (N5497, N5494, N4758);
xor XOR2 (N5498, N5489, N3977);
buf BUF1 (N5499, N5484);
or OR4 (N5500, N5496, N1670, N2422, N1036);
xor XOR2 (N5501, N5467, N869);
xor XOR2 (N5502, N5495, N2150);
nand NAND4 (N5503, N5492, N5274, N517, N91);
nor NOR3 (N5504, N5501, N2787, N1528);
or OR2 (N5505, N5488, N1759);
xor XOR2 (N5506, N5505, N1277);
nor NOR4 (N5507, N5498, N4093, N5290, N799);
xor XOR2 (N5508, N5506, N4829);
not NOT1 (N5509, N5497);
or OR3 (N5510, N5504, N2316, N654);
or OR3 (N5511, N5499, N5482, N5264);
not NOT1 (N5512, N4508);
not NOT1 (N5513, N5511);
not NOT1 (N5514, N5512);
buf BUF1 (N5515, N5503);
not NOT1 (N5516, N5490);
not NOT1 (N5517, N5509);
nand NAND3 (N5518, N5513, N5074, N4963);
xor XOR2 (N5519, N5514, N169);
not NOT1 (N5520, N5516);
xor XOR2 (N5521, N5517, N500);
and AND4 (N5522, N5500, N232, N778, N4605);
not NOT1 (N5523, N5515);
xor XOR2 (N5524, N5508, N3533);
nand NAND2 (N5525, N5518, N1275);
and AND2 (N5526, N5510, N5183);
not NOT1 (N5527, N5526);
not NOT1 (N5528, N5525);
nand NAND4 (N5529, N5527, N3467, N981, N2087);
xor XOR2 (N5530, N5521, N662);
buf BUF1 (N5531, N5528);
not NOT1 (N5532, N5530);
not NOT1 (N5533, N5507);
xor XOR2 (N5534, N5524, N2515);
buf BUF1 (N5535, N5520);
and AND2 (N5536, N5522, N4066);
xor XOR2 (N5537, N5523, N4819);
xor XOR2 (N5538, N5536, N636);
nor NOR4 (N5539, N5519, N2094, N2649, N3903);
nor NOR3 (N5540, N5538, N3577, N824);
or OR4 (N5541, N5535, N4814, N1016, N2377);
nand NAND2 (N5542, N5534, N1558);
nor NOR4 (N5543, N5539, N2479, N3296, N3670);
nor NOR2 (N5544, N5541, N3633);
and AND2 (N5545, N5532, N3389);
xor XOR2 (N5546, N5529, N5495);
nand NAND4 (N5547, N5546, N5179, N3121, N107);
nand NAND4 (N5548, N5544, N184, N2725, N3990);
buf BUF1 (N5549, N5540);
not NOT1 (N5550, N5543);
xor XOR2 (N5551, N5502, N4865);
nand NAND3 (N5552, N5550, N4896, N432);
xor XOR2 (N5553, N5547, N1475);
nor NOR3 (N5554, N5545, N762, N4456);
or OR2 (N5555, N5549, N3964);
buf BUF1 (N5556, N5552);
xor XOR2 (N5557, N5533, N386);
xor XOR2 (N5558, N5555, N2856);
not NOT1 (N5559, N5557);
not NOT1 (N5560, N5551);
or OR2 (N5561, N5542, N3353);
nor NOR4 (N5562, N5548, N1502, N3905, N1797);
buf BUF1 (N5563, N5553);
nor NOR2 (N5564, N5563, N1204);
buf BUF1 (N5565, N5560);
nand NAND4 (N5566, N5537, N3738, N1190, N115);
nor NOR3 (N5567, N5561, N5262, N412);
nand NAND4 (N5568, N5559, N32, N1781, N1878);
nor NOR3 (N5569, N5566, N2147, N305);
not NOT1 (N5570, N5565);
and AND4 (N5571, N5569, N5136, N4612, N340);
or OR2 (N5572, N5558, N1588);
nand NAND2 (N5573, N5570, N2146);
and AND2 (N5574, N5572, N3447);
nor NOR3 (N5575, N5571, N210, N3132);
xor XOR2 (N5576, N5567, N3361);
not NOT1 (N5577, N5575);
xor XOR2 (N5578, N5554, N39);
buf BUF1 (N5579, N5573);
and AND3 (N5580, N5577, N1482, N2771);
buf BUF1 (N5581, N5578);
nor NOR2 (N5582, N5579, N2863);
or OR3 (N5583, N5562, N4703, N2853);
xor XOR2 (N5584, N5531, N4631);
and AND4 (N5585, N5581, N926, N3157, N741);
and AND3 (N5586, N5574, N3615, N1348);
not NOT1 (N5587, N5568);
not NOT1 (N5588, N5583);
and AND4 (N5589, N5585, N2968, N3150, N4649);
not NOT1 (N5590, N5582);
not NOT1 (N5591, N5588);
buf BUF1 (N5592, N5591);
and AND4 (N5593, N5564, N3086, N5424, N504);
or OR2 (N5594, N5580, N103);
and AND4 (N5595, N5593, N1949, N1381, N4784);
nor NOR4 (N5596, N5556, N2307, N951, N1636);
xor XOR2 (N5597, N5592, N4389);
buf BUF1 (N5598, N5596);
not NOT1 (N5599, N5595);
or OR4 (N5600, N5587, N5211, N4504, N3280);
buf BUF1 (N5601, N5590);
xor XOR2 (N5602, N5584, N2736);
xor XOR2 (N5603, N5602, N1580);
nand NAND4 (N5604, N5600, N1502, N4476, N1169);
buf BUF1 (N5605, N5603);
xor XOR2 (N5606, N5589, N4011);
or OR3 (N5607, N5601, N1391, N5028);
xor XOR2 (N5608, N5605, N3307);
nand NAND2 (N5609, N5598, N1004);
nor NOR3 (N5610, N5586, N5023, N4279);
xor XOR2 (N5611, N5607, N479);
nor NOR3 (N5612, N5604, N1025, N3342);
and AND4 (N5613, N5576, N1953, N3673, N4916);
and AND4 (N5614, N5599, N628, N4285, N398);
and AND3 (N5615, N5614, N2520, N915);
not NOT1 (N5616, N5611);
not NOT1 (N5617, N5616);
nor NOR2 (N5618, N5606, N145);
xor XOR2 (N5619, N5597, N4438);
nor NOR2 (N5620, N5609, N1711);
and AND4 (N5621, N5610, N3090, N2825, N1657);
and AND2 (N5622, N5612, N1568);
xor XOR2 (N5623, N5619, N5068);
nand NAND4 (N5624, N5622, N4129, N918, N3052);
not NOT1 (N5625, N5623);
xor XOR2 (N5626, N5624, N1379);
nand NAND3 (N5627, N5626, N1298, N1159);
nor NOR2 (N5628, N5627, N1660);
buf BUF1 (N5629, N5621);
buf BUF1 (N5630, N5628);
xor XOR2 (N5631, N5613, N2297);
xor XOR2 (N5632, N5594, N679);
nor NOR2 (N5633, N5631, N2076);
and AND3 (N5634, N5625, N1661, N345);
and AND2 (N5635, N5615, N5502);
and AND3 (N5636, N5618, N5555, N2935);
buf BUF1 (N5637, N5608);
and AND4 (N5638, N5635, N2119, N1808, N2217);
buf BUF1 (N5639, N5617);
and AND3 (N5640, N5630, N8, N3785);
and AND2 (N5641, N5632, N186);
nor NOR3 (N5642, N5634, N5536, N1862);
nor NOR2 (N5643, N5633, N1850);
or OR4 (N5644, N5639, N4014, N1109, N3627);
or OR4 (N5645, N5638, N4801, N4839, N670);
and AND4 (N5646, N5629, N3903, N2793, N4392);
xor XOR2 (N5647, N5644, N506);
xor XOR2 (N5648, N5637, N1651);
nand NAND2 (N5649, N5641, N645);
and AND4 (N5650, N5642, N3916, N4501, N5249);
not NOT1 (N5651, N5646);
xor XOR2 (N5652, N5647, N1875);
or OR4 (N5653, N5648, N2164, N2729, N5395);
xor XOR2 (N5654, N5649, N2114);
not NOT1 (N5655, N5654);
nor NOR4 (N5656, N5655, N1774, N1455, N3483);
nand NAND3 (N5657, N5650, N5023, N4757);
buf BUF1 (N5658, N5656);
nor NOR2 (N5659, N5652, N2382);
buf BUF1 (N5660, N5636);
and AND4 (N5661, N5657, N1693, N570, N4905);
and AND2 (N5662, N5643, N3611);
and AND4 (N5663, N5640, N5422, N2534, N1331);
and AND3 (N5664, N5658, N4213, N2252);
and AND3 (N5665, N5661, N4621, N3584);
and AND3 (N5666, N5662, N4267, N5415);
buf BUF1 (N5667, N5663);
nor NOR4 (N5668, N5651, N1898, N221, N4483);
xor XOR2 (N5669, N5666, N4074);
xor XOR2 (N5670, N5664, N4165);
xor XOR2 (N5671, N5670, N2047);
nor NOR2 (N5672, N5665, N3226);
or OR4 (N5673, N5671, N2647, N4942, N2633);
nor NOR3 (N5674, N5669, N5122, N1876);
not NOT1 (N5675, N5668);
xor XOR2 (N5676, N5667, N3262);
nand NAND2 (N5677, N5659, N1295);
and AND3 (N5678, N5673, N1266, N3707);
buf BUF1 (N5679, N5676);
not NOT1 (N5680, N5679);
nor NOR4 (N5681, N5675, N1543, N4588, N2942);
buf BUF1 (N5682, N5620);
buf BUF1 (N5683, N5674);
and AND2 (N5684, N5678, N3155);
not NOT1 (N5685, N5645);
nand NAND2 (N5686, N5672, N4526);
buf BUF1 (N5687, N5681);
or OR2 (N5688, N5682, N4831);
or OR4 (N5689, N5680, N3281, N3661, N1312);
nor NOR4 (N5690, N5653, N1528, N622, N1454);
and AND2 (N5691, N5683, N1134);
nor NOR3 (N5692, N5691, N2087, N3451);
nand NAND4 (N5693, N5688, N5330, N2166, N3202);
buf BUF1 (N5694, N5692);
or OR3 (N5695, N5694, N3517, N774);
buf BUF1 (N5696, N5660);
nor NOR4 (N5697, N5685, N135, N340, N4841);
nand NAND2 (N5698, N5686, N3895);
not NOT1 (N5699, N5687);
nor NOR4 (N5700, N5684, N4550, N3334, N2152);
and AND2 (N5701, N5693, N2828);
nor NOR4 (N5702, N5695, N2389, N1042, N5353);
not NOT1 (N5703, N5690);
and AND4 (N5704, N5696, N2080, N3197, N5619);
and AND2 (N5705, N5699, N2565);
nand NAND2 (N5706, N5677, N1700);
or OR2 (N5707, N5703, N1819);
buf BUF1 (N5708, N5706);
and AND2 (N5709, N5701, N1645);
or OR2 (N5710, N5705, N4668);
not NOT1 (N5711, N5702);
or OR2 (N5712, N5708, N321);
nand NAND3 (N5713, N5711, N1194, N4851);
or OR3 (N5714, N5700, N4421, N2690);
or OR4 (N5715, N5698, N4538, N2439, N5005);
xor XOR2 (N5716, N5709, N2854);
not NOT1 (N5717, N5714);
nor NOR4 (N5718, N5712, N650, N3050, N809);
or OR3 (N5719, N5717, N2023, N1612);
or OR4 (N5720, N5704, N2435, N4492, N3132);
not NOT1 (N5721, N5707);
nor NOR4 (N5722, N5718, N148, N5010, N5162);
xor XOR2 (N5723, N5710, N1688);
not NOT1 (N5724, N5716);
nor NOR2 (N5725, N5713, N4084);
or OR2 (N5726, N5724, N3591);
buf BUF1 (N5727, N5689);
xor XOR2 (N5728, N5721, N3009);
xor XOR2 (N5729, N5722, N3709);
not NOT1 (N5730, N5729);
and AND3 (N5731, N5697, N2726, N3869);
nand NAND2 (N5732, N5730, N5388);
buf BUF1 (N5733, N5725);
not NOT1 (N5734, N5723);
not NOT1 (N5735, N5733);
or OR3 (N5736, N5734, N4059, N2459);
buf BUF1 (N5737, N5735);
or OR3 (N5738, N5726, N3488, N3234);
xor XOR2 (N5739, N5731, N2336);
buf BUF1 (N5740, N5737);
or OR2 (N5741, N5715, N325);
or OR2 (N5742, N5736, N783);
and AND4 (N5743, N5719, N4583, N4078, N2284);
or OR4 (N5744, N5740, N5112, N5282, N596);
xor XOR2 (N5745, N5744, N691);
or OR3 (N5746, N5739, N2199, N5634);
or OR2 (N5747, N5728, N472);
nor NOR3 (N5748, N5741, N4465, N4305);
or OR3 (N5749, N5748, N3030, N3675);
nor NOR3 (N5750, N5720, N3928, N3100);
buf BUF1 (N5751, N5749);
xor XOR2 (N5752, N5743, N5241);
not NOT1 (N5753, N5738);
nor NOR4 (N5754, N5752, N4757, N3977, N3028);
not NOT1 (N5755, N5747);
nand NAND4 (N5756, N5755, N2162, N3532, N1087);
nand NAND3 (N5757, N5746, N3494, N60);
not NOT1 (N5758, N5742);
buf BUF1 (N5759, N5745);
nand NAND4 (N5760, N5756, N1632, N5543, N539);
xor XOR2 (N5761, N5732, N894);
buf BUF1 (N5762, N5757);
nand NAND2 (N5763, N5761, N1423);
nand NAND3 (N5764, N5762, N2825, N3161);
buf BUF1 (N5765, N5754);
buf BUF1 (N5766, N5727);
and AND4 (N5767, N5759, N1506, N2992, N3840);
and AND4 (N5768, N5767, N801, N864, N4773);
nand NAND4 (N5769, N5764, N910, N2592, N3003);
nor NOR4 (N5770, N5769, N299, N4848, N2212);
buf BUF1 (N5771, N5753);
or OR2 (N5772, N5750, N2990);
and AND4 (N5773, N5751, N858, N4902, N290);
xor XOR2 (N5774, N5765, N2823);
xor XOR2 (N5775, N5773, N2041);
and AND2 (N5776, N5771, N5565);
nor NOR4 (N5777, N5758, N3048, N2746, N5568);
not NOT1 (N5778, N5768);
nand NAND2 (N5779, N5777, N91);
buf BUF1 (N5780, N5778);
xor XOR2 (N5781, N5775, N2722);
buf BUF1 (N5782, N5770);
buf BUF1 (N5783, N5781);
buf BUF1 (N5784, N5782);
buf BUF1 (N5785, N5780);
xor XOR2 (N5786, N5774, N5440);
or OR3 (N5787, N5766, N4182, N2282);
and AND3 (N5788, N5776, N2912, N2300);
nand NAND4 (N5789, N5783, N2536, N34, N284);
nand NAND3 (N5790, N5787, N4718, N2571);
xor XOR2 (N5791, N5790, N3128);
xor XOR2 (N5792, N5772, N450);
or OR3 (N5793, N5784, N5568, N608);
buf BUF1 (N5794, N5785);
nand NAND3 (N5795, N5788, N3179, N4324);
xor XOR2 (N5796, N5779, N1541);
xor XOR2 (N5797, N5763, N5739);
and AND2 (N5798, N5797, N2264);
xor XOR2 (N5799, N5789, N4993);
and AND4 (N5800, N5798, N2789, N1999, N3457);
nand NAND3 (N5801, N5796, N2305, N3338);
nor NOR2 (N5802, N5786, N882);
nand NAND3 (N5803, N5791, N788, N2521);
and AND4 (N5804, N5792, N1976, N2357, N4833);
xor XOR2 (N5805, N5795, N2851);
buf BUF1 (N5806, N5804);
xor XOR2 (N5807, N5800, N547);
nand NAND2 (N5808, N5794, N2483);
or OR3 (N5809, N5801, N4963, N3566);
and AND4 (N5810, N5760, N3326, N4962, N242);
and AND4 (N5811, N5802, N3170, N2786, N5259);
or OR3 (N5812, N5808, N4882, N3958);
xor XOR2 (N5813, N5809, N1989);
nor NOR3 (N5814, N5806, N5694, N1054);
buf BUF1 (N5815, N5812);
not NOT1 (N5816, N5805);
or OR2 (N5817, N5813, N3215);
and AND4 (N5818, N5807, N4191, N1205, N4058);
xor XOR2 (N5819, N5817, N1986);
and AND3 (N5820, N5816, N2555, N5077);
or OR4 (N5821, N5810, N2610, N2833, N1365);
or OR3 (N5822, N5820, N4785, N2041);
nand NAND2 (N5823, N5793, N1151);
nand NAND2 (N5824, N5821, N588);
not NOT1 (N5825, N5818);
or OR4 (N5826, N5825, N4106, N4610, N621);
buf BUF1 (N5827, N5826);
buf BUF1 (N5828, N5811);
and AND3 (N5829, N5827, N3772, N4228);
not NOT1 (N5830, N5799);
or OR2 (N5831, N5823, N1141);
nor NOR3 (N5832, N5803, N5201, N3843);
nor NOR4 (N5833, N5832, N796, N2111, N3434);
or OR2 (N5834, N5814, N1431);
or OR2 (N5835, N5815, N5602);
or OR2 (N5836, N5830, N5183);
or OR4 (N5837, N5833, N2222, N4956, N2544);
or OR3 (N5838, N5836, N800, N2579);
and AND4 (N5839, N5838, N4964, N1228, N3268);
buf BUF1 (N5840, N5837);
nor NOR3 (N5841, N5831, N3406, N1083);
or OR2 (N5842, N5824, N3653);
nand NAND4 (N5843, N5840, N5107, N4088, N1557);
buf BUF1 (N5844, N5839);
nor NOR3 (N5845, N5828, N5403, N1157);
buf BUF1 (N5846, N5843);
nor NOR2 (N5847, N5846, N4212);
xor XOR2 (N5848, N5842, N3547);
nand NAND3 (N5849, N5829, N371, N3525);
buf BUF1 (N5850, N5848);
and AND2 (N5851, N5844, N4001);
nor NOR2 (N5852, N5841, N4147);
or OR3 (N5853, N5822, N5035, N3515);
nor NOR4 (N5854, N5819, N2839, N1595, N2538);
not NOT1 (N5855, N5850);
nand NAND2 (N5856, N5849, N1671);
buf BUF1 (N5857, N5834);
not NOT1 (N5858, N5847);
nor NOR2 (N5859, N5835, N989);
xor XOR2 (N5860, N5853, N3904);
buf BUF1 (N5861, N5845);
or OR3 (N5862, N5861, N3560, N5571);
or OR2 (N5863, N5856, N2059);
xor XOR2 (N5864, N5863, N1086);
nor NOR2 (N5865, N5864, N2544);
xor XOR2 (N5866, N5857, N4451);
buf BUF1 (N5867, N5852);
buf BUF1 (N5868, N5860);
not NOT1 (N5869, N5868);
buf BUF1 (N5870, N5855);
not NOT1 (N5871, N5867);
buf BUF1 (N5872, N5870);
not NOT1 (N5873, N5854);
nand NAND3 (N5874, N5872, N2432, N2575);
nor NOR2 (N5875, N5862, N1902);
xor XOR2 (N5876, N5873, N4362);
not NOT1 (N5877, N5851);
buf BUF1 (N5878, N5858);
nand NAND3 (N5879, N5866, N963, N5231);
nor NOR2 (N5880, N5879, N1718);
not NOT1 (N5881, N5877);
buf BUF1 (N5882, N5865);
not NOT1 (N5883, N5871);
or OR4 (N5884, N5882, N3534, N1154, N534);
xor XOR2 (N5885, N5859, N4554);
and AND3 (N5886, N5869, N1949, N4195);
xor XOR2 (N5887, N5874, N1480);
nand NAND2 (N5888, N5876, N3254);
not NOT1 (N5889, N5880);
xor XOR2 (N5890, N5886, N4199);
nor NOR3 (N5891, N5878, N4146, N2076);
not NOT1 (N5892, N5883);
not NOT1 (N5893, N5892);
nor NOR3 (N5894, N5889, N3287, N4722);
and AND2 (N5895, N5885, N5216);
buf BUF1 (N5896, N5881);
not NOT1 (N5897, N5893);
buf BUF1 (N5898, N5890);
xor XOR2 (N5899, N5891, N5828);
nand NAND2 (N5900, N5894, N5000);
nor NOR3 (N5901, N5888, N2811, N4);
or OR2 (N5902, N5900, N4741);
buf BUF1 (N5903, N5902);
not NOT1 (N5904, N5884);
or OR3 (N5905, N5903, N1866, N3501);
nand NAND4 (N5906, N5901, N5658, N2551, N3492);
nand NAND2 (N5907, N5875, N1555);
not NOT1 (N5908, N5895);
nand NAND3 (N5909, N5896, N1048, N5623);
nand NAND2 (N5910, N5905, N699);
nor NOR3 (N5911, N5908, N5040, N4167);
or OR3 (N5912, N5898, N5247, N1559);
nand NAND4 (N5913, N5909, N1780, N1174, N2976);
nand NAND4 (N5914, N5910, N2876, N33, N5174);
nor NOR2 (N5915, N5913, N670);
not NOT1 (N5916, N5887);
nor NOR4 (N5917, N5907, N3979, N5387, N4239);
not NOT1 (N5918, N5897);
and AND4 (N5919, N5904, N3415, N4294, N3668);
nor NOR3 (N5920, N5916, N4874, N2910);
not NOT1 (N5921, N5906);
not NOT1 (N5922, N5921);
xor XOR2 (N5923, N5920, N1990);
xor XOR2 (N5924, N5923, N151);
and AND2 (N5925, N5911, N4382);
xor XOR2 (N5926, N5922, N1891);
nand NAND4 (N5927, N5924, N1525, N1509, N1760);
xor XOR2 (N5928, N5912, N2433);
nor NOR4 (N5929, N5927, N4807, N3930, N5885);
or OR3 (N5930, N5914, N4586, N1977);
not NOT1 (N5931, N5919);
or OR2 (N5932, N5926, N3029);
buf BUF1 (N5933, N5929);
xor XOR2 (N5934, N5918, N811);
nor NOR3 (N5935, N5917, N3931, N1610);
not NOT1 (N5936, N5931);
nand NAND4 (N5937, N5928, N665, N432, N1099);
or OR3 (N5938, N5937, N616, N448);
nand NAND3 (N5939, N5938, N1670, N1456);
or OR3 (N5940, N5925, N3642, N2479);
not NOT1 (N5941, N5930);
nor NOR3 (N5942, N5932, N3862, N5220);
not NOT1 (N5943, N5934);
nand NAND3 (N5944, N5933, N3536, N1108);
and AND3 (N5945, N5936, N3128, N3136);
not NOT1 (N5946, N5935);
nand NAND3 (N5947, N5915, N3067, N4547);
nor NOR3 (N5948, N5945, N5583, N2356);
nand NAND3 (N5949, N5946, N542, N2100);
xor XOR2 (N5950, N5943, N2047);
xor XOR2 (N5951, N5899, N4835);
not NOT1 (N5952, N5949);
nand NAND3 (N5953, N5941, N1133, N5694);
and AND3 (N5954, N5940, N2446, N4761);
nand NAND3 (N5955, N5952, N1129, N4583);
nand NAND2 (N5956, N5939, N357);
not NOT1 (N5957, N5955);
nand NAND2 (N5958, N5950, N2904);
not NOT1 (N5959, N5944);
xor XOR2 (N5960, N5959, N193);
xor XOR2 (N5961, N5956, N4965);
buf BUF1 (N5962, N5942);
and AND2 (N5963, N5947, N3407);
not NOT1 (N5964, N5951);
xor XOR2 (N5965, N5963, N1896);
not NOT1 (N5966, N5954);
or OR3 (N5967, N5961, N553, N4239);
and AND2 (N5968, N5960, N5148);
or OR4 (N5969, N5953, N4339, N5245, N372);
and AND2 (N5970, N5957, N5288);
buf BUF1 (N5971, N5948);
nand NAND3 (N5972, N5969, N3705, N5453);
buf BUF1 (N5973, N5964);
not NOT1 (N5974, N5973);
and AND3 (N5975, N5971, N1108, N4427);
xor XOR2 (N5976, N5972, N4239);
nand NAND4 (N5977, N5958, N2422, N1533, N5677);
nand NAND2 (N5978, N5974, N2334);
nor NOR4 (N5979, N5976, N2172, N1423, N2645);
and AND3 (N5980, N5979, N2407, N3430);
not NOT1 (N5981, N5962);
or OR2 (N5982, N5977, N4748);
or OR3 (N5983, N5982, N5479, N1326);
or OR4 (N5984, N5983, N3305, N3260, N3809);
not NOT1 (N5985, N5970);
buf BUF1 (N5986, N5984);
xor XOR2 (N5987, N5968, N1291);
or OR4 (N5988, N5978, N3397, N5481, N3306);
buf BUF1 (N5989, N5988);
not NOT1 (N5990, N5987);
buf BUF1 (N5991, N5985);
and AND2 (N5992, N5991, N3229);
buf BUF1 (N5993, N5989);
nor NOR3 (N5994, N5986, N5129, N5005);
xor XOR2 (N5995, N5990, N651);
not NOT1 (N5996, N5967);
buf BUF1 (N5997, N5981);
or OR4 (N5998, N5975, N2070, N5995, N3935);
nor NOR4 (N5999, N29, N5662, N573, N3738);
not NOT1 (N6000, N5994);
not NOT1 (N6001, N5992);
and AND3 (N6002, N5993, N4728, N2496);
and AND2 (N6003, N5980, N1867);
nand NAND3 (N6004, N6000, N3774, N5086);
not NOT1 (N6005, N6004);
not NOT1 (N6006, N5965);
or OR4 (N6007, N5997, N632, N2422, N881);
not NOT1 (N6008, N6006);
not NOT1 (N6009, N6001);
and AND3 (N6010, N5966, N3096, N295);
and AND4 (N6011, N5998, N5082, N3266, N2372);
nor NOR3 (N6012, N6011, N4492, N3336);
not NOT1 (N6013, N6007);
buf BUF1 (N6014, N6008);
or OR2 (N6015, N6003, N2568);
or OR4 (N6016, N6013, N1361, N2715, N2191);
and AND4 (N6017, N6014, N5162, N4450, N2180);
xor XOR2 (N6018, N6002, N2458);
nor NOR3 (N6019, N6012, N733, N5690);
nand NAND4 (N6020, N6019, N1868, N565, N4926);
and AND3 (N6021, N6005, N5447, N2492);
not NOT1 (N6022, N6015);
not NOT1 (N6023, N6021);
nand NAND4 (N6024, N6020, N5608, N4643, N1713);
xor XOR2 (N6025, N6024, N5994);
nor NOR4 (N6026, N5996, N5912, N5735, N1183);
and AND2 (N6027, N6026, N3033);
buf BUF1 (N6028, N6017);
nor NOR4 (N6029, N6028, N4603, N4738, N4224);
xor XOR2 (N6030, N6029, N5122);
and AND4 (N6031, N6030, N825, N4921, N2308);
not NOT1 (N6032, N6031);
xor XOR2 (N6033, N6032, N5088);
nand NAND3 (N6034, N6025, N4051, N1908);
or OR3 (N6035, N6016, N1710, N1828);
nand NAND4 (N6036, N6009, N3416, N3712, N742);
or OR4 (N6037, N6035, N1822, N5117, N5872);
and AND4 (N6038, N6027, N2245, N1455, N5953);
and AND2 (N6039, N6034, N764);
or OR3 (N6040, N6036, N1248, N229);
and AND4 (N6041, N6010, N3173, N4308, N1);
nor NOR4 (N6042, N6033, N3447, N4346, N2573);
or OR3 (N6043, N6023, N2640, N2935);
nand NAND2 (N6044, N6041, N787);
nand NAND2 (N6045, N6040, N660);
and AND4 (N6046, N6044, N1650, N3019, N3063);
nor NOR3 (N6047, N6043, N1082, N5824);
buf BUF1 (N6048, N6047);
nor NOR3 (N6049, N5999, N1035, N2595);
or OR4 (N6050, N6022, N2917, N3092, N5240);
or OR4 (N6051, N6042, N1655, N971, N307);
and AND4 (N6052, N6046, N1170, N2915, N4826);
nand NAND3 (N6053, N6049, N399, N4194);
xor XOR2 (N6054, N6037, N5392);
xor XOR2 (N6055, N6039, N355);
buf BUF1 (N6056, N6055);
nand NAND3 (N6057, N6048, N5609, N5925);
buf BUF1 (N6058, N6018);
not NOT1 (N6059, N6056);
nor NOR3 (N6060, N6052, N3679, N2263);
not NOT1 (N6061, N6038);
nor NOR4 (N6062, N6054, N1439, N3602, N4916);
xor XOR2 (N6063, N6051, N171);
buf BUF1 (N6064, N6062);
and AND4 (N6065, N6057, N2591, N1929, N2187);
xor XOR2 (N6066, N6063, N4022);
or OR3 (N6067, N6065, N5710, N3054);
or OR4 (N6068, N6059, N217, N4973, N4260);
xor XOR2 (N6069, N6053, N1035);
nand NAND3 (N6070, N6058, N4379, N1851);
nand NAND2 (N6071, N6070, N890);
xor XOR2 (N6072, N6068, N1624);
buf BUF1 (N6073, N6069);
nand NAND2 (N6074, N6050, N5510);
or OR4 (N6075, N6061, N4854, N5938, N993);
buf BUF1 (N6076, N6072);
or OR2 (N6077, N6071, N5536);
and AND3 (N6078, N6066, N5840, N4343);
buf BUF1 (N6079, N6067);
nand NAND4 (N6080, N6078, N816, N6072, N161);
nand NAND3 (N6081, N6045, N3854, N1563);
xor XOR2 (N6082, N6060, N1988);
or OR2 (N6083, N6080, N617);
not NOT1 (N6084, N6073);
or OR4 (N6085, N6076, N5688, N5137, N443);
nand NAND2 (N6086, N6084, N3701);
buf BUF1 (N6087, N6077);
nor NOR3 (N6088, N6087, N2377, N2418);
buf BUF1 (N6089, N6079);
buf BUF1 (N6090, N6083);
or OR2 (N6091, N6064, N5932);
nand NAND3 (N6092, N6089, N2143, N5886);
and AND4 (N6093, N6092, N3389, N3689, N1965);
buf BUF1 (N6094, N6086);
nor NOR4 (N6095, N6074, N4900, N5205, N2709);
and AND4 (N6096, N6090, N5648, N4539, N835);
and AND3 (N6097, N6094, N3235, N3860);
nor NOR3 (N6098, N6088, N1682, N2199);
not NOT1 (N6099, N6098);
nor NOR3 (N6100, N6099, N5476, N4788);
xor XOR2 (N6101, N6093, N425);
or OR4 (N6102, N6101, N1026, N157, N4662);
xor XOR2 (N6103, N6075, N4133);
xor XOR2 (N6104, N6096, N2686);
xor XOR2 (N6105, N6082, N5079);
or OR2 (N6106, N6104, N841);
and AND4 (N6107, N6081, N166, N1379, N140);
nand NAND3 (N6108, N6105, N5763, N665);
nor NOR3 (N6109, N6100, N2275, N2762);
nor NOR2 (N6110, N6095, N1931);
nor NOR2 (N6111, N6108, N5595);
nand NAND3 (N6112, N6110, N1371, N476);
xor XOR2 (N6113, N6097, N1131);
xor XOR2 (N6114, N6113, N2962);
not NOT1 (N6115, N6102);
not NOT1 (N6116, N6106);
xor XOR2 (N6117, N6114, N3020);
not NOT1 (N6118, N6085);
xor XOR2 (N6119, N6103, N2619);
not NOT1 (N6120, N6118);
nor NOR2 (N6121, N6111, N3159);
xor XOR2 (N6122, N6117, N4500);
nand NAND4 (N6123, N6109, N2629, N5297, N5121);
and AND3 (N6124, N6122, N4085, N80);
nor NOR2 (N6125, N6091, N926);
nand NAND2 (N6126, N6123, N1550);
and AND4 (N6127, N6115, N3391, N944, N1384);
buf BUF1 (N6128, N6120);
nor NOR3 (N6129, N6128, N456, N4129);
nor NOR2 (N6130, N6107, N5060);
or OR4 (N6131, N6119, N5220, N769, N389);
buf BUF1 (N6132, N6127);
buf BUF1 (N6133, N6131);
or OR4 (N6134, N6112, N1201, N4622, N1962);
nor NOR4 (N6135, N6116, N582, N3, N315);
and AND3 (N6136, N6129, N478, N5645);
and AND2 (N6137, N6126, N94);
buf BUF1 (N6138, N6130);
and AND3 (N6139, N6134, N1928, N1383);
nand NAND3 (N6140, N6125, N819, N2796);
xor XOR2 (N6141, N6133, N4544);
nor NOR2 (N6142, N6121, N4895);
or OR4 (N6143, N6140, N5046, N2481, N3084);
and AND2 (N6144, N6142, N5587);
and AND4 (N6145, N6136, N3768, N2987, N2972);
xor XOR2 (N6146, N6138, N1489);
and AND4 (N6147, N6124, N5869, N343, N2560);
nand NAND2 (N6148, N6146, N627);
not NOT1 (N6149, N6132);
xor XOR2 (N6150, N6144, N2521);
xor XOR2 (N6151, N6145, N3705);
not NOT1 (N6152, N6139);
or OR2 (N6153, N6149, N4788);
buf BUF1 (N6154, N6141);
not NOT1 (N6155, N6143);
or OR2 (N6156, N6153, N2980);
nand NAND3 (N6157, N6150, N4320, N1479);
nand NAND3 (N6158, N6135, N3005, N3615);
and AND3 (N6159, N6137, N5620, N2698);
xor XOR2 (N6160, N6156, N3788);
or OR3 (N6161, N6155, N2563, N4076);
nor NOR2 (N6162, N6147, N2953);
buf BUF1 (N6163, N6159);
nand NAND3 (N6164, N6160, N2554, N2391);
not NOT1 (N6165, N6148);
xor XOR2 (N6166, N6163, N1136);
or OR2 (N6167, N6166, N693);
and AND3 (N6168, N6165, N809, N1255);
and AND3 (N6169, N6157, N2172, N1496);
and AND4 (N6170, N6168, N1349, N1486, N2654);
nor NOR3 (N6171, N6167, N2952, N5115);
nand NAND2 (N6172, N6171, N5120);
xor XOR2 (N6173, N6154, N1666);
buf BUF1 (N6174, N6170);
not NOT1 (N6175, N6152);
and AND2 (N6176, N6169, N3586);
nand NAND4 (N6177, N6151, N3122, N430, N2457);
or OR3 (N6178, N6158, N5198, N5686);
not NOT1 (N6179, N6161);
nand NAND2 (N6180, N6178, N3275);
nor NOR4 (N6181, N6175, N117, N3819, N4771);
and AND2 (N6182, N6173, N3842);
xor XOR2 (N6183, N6177, N1586);
xor XOR2 (N6184, N6172, N2281);
or OR4 (N6185, N6180, N3250, N4704, N3776);
and AND2 (N6186, N6181, N3514);
nand NAND4 (N6187, N6183, N3126, N1987, N5194);
or OR4 (N6188, N6186, N3340, N1347, N3580);
or OR2 (N6189, N6162, N3522);
and AND4 (N6190, N6182, N6168, N4406, N5392);
nand NAND4 (N6191, N6174, N618, N2582, N3925);
buf BUF1 (N6192, N6185);
and AND2 (N6193, N6179, N1041);
and AND2 (N6194, N6184, N3901);
buf BUF1 (N6195, N6188);
and AND4 (N6196, N6189, N2029, N5850, N3407);
nand NAND2 (N6197, N6164, N6009);
nor NOR4 (N6198, N6191, N5146, N4674, N4832);
nor NOR2 (N6199, N6195, N722);
not NOT1 (N6200, N6190);
and AND4 (N6201, N6198, N2529, N3878, N2416);
nor NOR3 (N6202, N6187, N1386, N5586);
nand NAND3 (N6203, N6193, N5838, N5927);
and AND3 (N6204, N6203, N4062, N1957);
not NOT1 (N6205, N6200);
xor XOR2 (N6206, N6192, N672);
and AND3 (N6207, N6206, N4729, N1745);
xor XOR2 (N6208, N6194, N3262);
and AND2 (N6209, N6197, N1200);
xor XOR2 (N6210, N6199, N5888);
not NOT1 (N6211, N6201);
nor NOR4 (N6212, N6204, N3841, N5599, N5849);
not NOT1 (N6213, N6209);
and AND3 (N6214, N6207, N1773, N4543);
xor XOR2 (N6215, N6214, N6132);
xor XOR2 (N6216, N6208, N5981);
nor NOR3 (N6217, N6213, N3001, N4395);
or OR2 (N6218, N6176, N2737);
buf BUF1 (N6219, N6205);
nand NAND3 (N6220, N6219, N5227, N588);
and AND2 (N6221, N6215, N3743);
xor XOR2 (N6222, N6212, N1092);
or OR4 (N6223, N6196, N3252, N5807, N5740);
and AND2 (N6224, N6211, N2331);
xor XOR2 (N6225, N6224, N195);
buf BUF1 (N6226, N6217);
and AND4 (N6227, N6226, N96, N5219, N3105);
or OR4 (N6228, N6227, N5570, N3632, N4272);
buf BUF1 (N6229, N6225);
or OR2 (N6230, N6210, N1854);
buf BUF1 (N6231, N6218);
nor NOR3 (N6232, N6223, N4333, N3729);
nand NAND2 (N6233, N6202, N4979);
and AND4 (N6234, N6228, N4158, N5987, N4577);
xor XOR2 (N6235, N6222, N4697);
xor XOR2 (N6236, N6235, N512);
xor XOR2 (N6237, N6230, N436);
nand NAND2 (N6238, N6231, N5127);
xor XOR2 (N6239, N6229, N1223);
xor XOR2 (N6240, N6239, N4388);
or OR2 (N6241, N6233, N6046);
buf BUF1 (N6242, N6216);
nand NAND2 (N6243, N6241, N2875);
xor XOR2 (N6244, N6220, N1470);
nand NAND2 (N6245, N6242, N1168);
and AND3 (N6246, N6245, N3931, N3259);
buf BUF1 (N6247, N6244);
buf BUF1 (N6248, N6238);
nand NAND3 (N6249, N6247, N2736, N2607);
not NOT1 (N6250, N6248);
and AND2 (N6251, N6234, N6061);
and AND4 (N6252, N6243, N43, N5988, N3273);
or OR2 (N6253, N6236, N5668);
not NOT1 (N6254, N6221);
nor NOR3 (N6255, N6254, N611, N3753);
xor XOR2 (N6256, N6237, N155);
or OR2 (N6257, N6252, N2127);
and AND3 (N6258, N6256, N588, N1387);
buf BUF1 (N6259, N6249);
and AND4 (N6260, N6255, N2253, N1776, N582);
nor NOR2 (N6261, N6232, N3952);
xor XOR2 (N6262, N6240, N6261);
nor NOR3 (N6263, N3124, N6240, N5786);
or OR3 (N6264, N6246, N3840, N1286);
nand NAND4 (N6265, N6251, N4197, N449, N3118);
buf BUF1 (N6266, N6262);
and AND2 (N6267, N6263, N3026);
buf BUF1 (N6268, N6265);
xor XOR2 (N6269, N6257, N6211);
nand NAND2 (N6270, N6269, N3784);
nor NOR4 (N6271, N6259, N4385, N4357, N40);
buf BUF1 (N6272, N6258);
nand NAND2 (N6273, N6266, N3324);
or OR3 (N6274, N6273, N5758, N5633);
and AND2 (N6275, N6250, N5936);
and AND2 (N6276, N6270, N5749);
xor XOR2 (N6277, N6275, N5092);
not NOT1 (N6278, N6271);
buf BUF1 (N6279, N6267);
nor NOR4 (N6280, N6268, N5387, N3333, N5205);
and AND4 (N6281, N6277, N4326, N6072, N2922);
and AND2 (N6282, N6274, N2038);
buf BUF1 (N6283, N6282);
buf BUF1 (N6284, N6283);
not NOT1 (N6285, N6281);
and AND3 (N6286, N6260, N618, N5962);
or OR2 (N6287, N6253, N1795);
buf BUF1 (N6288, N6287);
nor NOR3 (N6289, N6278, N2251, N2388);
nand NAND3 (N6290, N6284, N5676, N4889);
or OR3 (N6291, N6276, N2529, N1501);
and AND4 (N6292, N6279, N1404, N5159, N3742);
and AND3 (N6293, N6292, N3438, N6084);
xor XOR2 (N6294, N6291, N2538);
xor XOR2 (N6295, N6264, N773);
and AND2 (N6296, N6294, N5761);
nand NAND3 (N6297, N6293, N2973, N6069);
or OR3 (N6298, N6280, N4796, N335);
xor XOR2 (N6299, N6272, N2119);
and AND4 (N6300, N6286, N3169, N3602, N5655);
or OR4 (N6301, N6288, N4664, N3237, N2247);
nor NOR2 (N6302, N6300, N670);
or OR3 (N6303, N6296, N1347, N5544);
and AND3 (N6304, N6302, N414, N734);
buf BUF1 (N6305, N6290);
and AND2 (N6306, N6289, N5669);
xor XOR2 (N6307, N6304, N3207);
or OR4 (N6308, N6297, N3981, N2161, N6017);
xor XOR2 (N6309, N6308, N1481);
and AND3 (N6310, N6309, N5367, N3955);
xor XOR2 (N6311, N6298, N1391);
nor NOR4 (N6312, N6306, N613, N6020, N6148);
not NOT1 (N6313, N6307);
not NOT1 (N6314, N6305);
and AND3 (N6315, N6314, N1457, N2906);
not NOT1 (N6316, N6299);
nor NOR4 (N6317, N6315, N2720, N782, N3852);
buf BUF1 (N6318, N6285);
or OR2 (N6319, N6303, N1585);
and AND4 (N6320, N6313, N903, N5866, N5085);
xor XOR2 (N6321, N6301, N818);
xor XOR2 (N6322, N6295, N3596);
or OR4 (N6323, N6317, N125, N3542, N6200);
nor NOR2 (N6324, N6318, N316);
xor XOR2 (N6325, N6319, N3823);
xor XOR2 (N6326, N6323, N4961);
xor XOR2 (N6327, N6322, N6008);
not NOT1 (N6328, N6316);
buf BUF1 (N6329, N6327);
and AND3 (N6330, N6324, N1707, N2671);
nand NAND4 (N6331, N6311, N5073, N4432, N3060);
buf BUF1 (N6332, N6310);
nor NOR2 (N6333, N6331, N6283);
nand NAND4 (N6334, N6326, N2531, N5313, N144);
nor NOR2 (N6335, N6334, N4006);
and AND4 (N6336, N6312, N614, N4540, N3605);
not NOT1 (N6337, N6325);
buf BUF1 (N6338, N6336);
nand NAND4 (N6339, N6338, N3699, N912, N3231);
buf BUF1 (N6340, N6333);
or OR4 (N6341, N6339, N1996, N3295, N1870);
or OR3 (N6342, N6328, N3489, N2023);
and AND4 (N6343, N6340, N3112, N3343, N5371);
and AND4 (N6344, N6337, N4370, N29, N4961);
buf BUF1 (N6345, N6341);
and AND2 (N6346, N6332, N3500);
and AND2 (N6347, N6345, N6045);
not NOT1 (N6348, N6344);
nor NOR4 (N6349, N6330, N618, N5592, N837);
nor NOR2 (N6350, N6349, N4611);
buf BUF1 (N6351, N6346);
or OR4 (N6352, N6351, N5889, N3825, N721);
buf BUF1 (N6353, N6329);
or OR3 (N6354, N6347, N5171, N2257);
buf BUF1 (N6355, N6353);
nand NAND3 (N6356, N6335, N1377, N2528);
buf BUF1 (N6357, N6354);
not NOT1 (N6358, N6350);
and AND4 (N6359, N6357, N5575, N3369, N6052);
nor NOR4 (N6360, N6356, N1290, N4488, N2741);
and AND3 (N6361, N6348, N4407, N1184);
buf BUF1 (N6362, N6360);
xor XOR2 (N6363, N6343, N5613);
buf BUF1 (N6364, N6321);
xor XOR2 (N6365, N6359, N2413);
nand NAND2 (N6366, N6361, N3578);
xor XOR2 (N6367, N6362, N4234);
buf BUF1 (N6368, N6367);
not NOT1 (N6369, N6342);
nand NAND2 (N6370, N6366, N2694);
nor NOR4 (N6371, N6320, N1735, N5831, N6017);
nand NAND4 (N6372, N6368, N3989, N1253, N6151);
nand NAND3 (N6373, N6358, N2861, N514);
buf BUF1 (N6374, N6369);
xor XOR2 (N6375, N6374, N4233);
and AND2 (N6376, N6372, N2337);
nand NAND4 (N6377, N6365, N344, N4058, N719);
and AND2 (N6378, N6364, N1639);
nand NAND4 (N6379, N6363, N2535, N5670, N5274);
and AND4 (N6380, N6352, N6083, N2383, N6297);
nand NAND3 (N6381, N6378, N1096, N3626);
nor NOR4 (N6382, N6373, N2945, N4947, N3194);
xor XOR2 (N6383, N6371, N2980);
nor NOR3 (N6384, N6370, N3248, N2782);
not NOT1 (N6385, N6381);
nand NAND3 (N6386, N6383, N857, N96);
buf BUF1 (N6387, N6377);
and AND4 (N6388, N6379, N1530, N2619, N1548);
nand NAND4 (N6389, N6376, N3604, N4158, N2128);
buf BUF1 (N6390, N6385);
and AND3 (N6391, N6387, N6125, N1851);
nor NOR4 (N6392, N6390, N2971, N1606, N3973);
nor NOR4 (N6393, N6391, N1933, N3383, N5018);
or OR3 (N6394, N6375, N4097, N3655);
not NOT1 (N6395, N6392);
buf BUF1 (N6396, N6388);
nand NAND4 (N6397, N6380, N2565, N5864, N3025);
not NOT1 (N6398, N6393);
and AND4 (N6399, N6395, N1774, N2656, N6041);
or OR3 (N6400, N6394, N2045, N4708);
nand NAND3 (N6401, N6355, N2157, N1857);
and AND4 (N6402, N6384, N4502, N4164, N4090);
buf BUF1 (N6403, N6386);
nor NOR3 (N6404, N6403, N706, N5520);
buf BUF1 (N6405, N6397);
and AND2 (N6406, N6399, N1320);
nor NOR2 (N6407, N6400, N4011);
nor NOR3 (N6408, N6406, N2090, N1646);
nor NOR3 (N6409, N6404, N6019, N4372);
or OR2 (N6410, N6396, N4369);
buf BUF1 (N6411, N6382);
not NOT1 (N6412, N6408);
nand NAND2 (N6413, N6410, N802);
or OR3 (N6414, N6412, N3823, N3696);
and AND2 (N6415, N6411, N2404);
and AND2 (N6416, N6407, N5617);
and AND4 (N6417, N6402, N3948, N2060, N3433);
or OR4 (N6418, N6398, N1888, N5911, N4247);
or OR3 (N6419, N6401, N1849, N4663);
or OR3 (N6420, N6417, N1914, N1959);
nor NOR4 (N6421, N6413, N4172, N4233, N4522);
nand NAND3 (N6422, N6414, N2840, N4708);
nand NAND3 (N6423, N6389, N5402, N1907);
xor XOR2 (N6424, N6421, N3994);
or OR2 (N6425, N6419, N4091);
nor NOR2 (N6426, N6416, N330);
not NOT1 (N6427, N6425);
buf BUF1 (N6428, N6427);
xor XOR2 (N6429, N6424, N1216);
buf BUF1 (N6430, N6426);
buf BUF1 (N6431, N6409);
buf BUF1 (N6432, N6422);
not NOT1 (N6433, N6415);
buf BUF1 (N6434, N6423);
xor XOR2 (N6435, N6429, N804);
nor NOR2 (N6436, N6434, N4620);
nand NAND3 (N6437, N6418, N2616, N3348);
nor NOR4 (N6438, N6435, N5804, N4872, N5857);
buf BUF1 (N6439, N6433);
or OR4 (N6440, N6430, N6346, N3755, N1796);
not NOT1 (N6441, N6439);
and AND4 (N6442, N6437, N1629, N5366, N6119);
buf BUF1 (N6443, N6432);
not NOT1 (N6444, N6428);
nand NAND3 (N6445, N6436, N3249, N3656);
and AND4 (N6446, N6440, N3807, N793, N1573);
and AND2 (N6447, N6405, N4756);
xor XOR2 (N6448, N6438, N1924);
or OR2 (N6449, N6443, N1369);
buf BUF1 (N6450, N6420);
nand NAND2 (N6451, N6446, N4591);
or OR3 (N6452, N6445, N3114, N4536);
nand NAND2 (N6453, N6444, N1650);
nor NOR2 (N6454, N6447, N5397);
xor XOR2 (N6455, N6452, N4738);
or OR2 (N6456, N6449, N2346);
or OR4 (N6457, N6442, N2794, N3548, N2767);
nor NOR2 (N6458, N6455, N2742);
not NOT1 (N6459, N6448);
buf BUF1 (N6460, N6453);
nor NOR3 (N6461, N6457, N3224, N2527);
nand NAND3 (N6462, N6461, N2452, N3187);
nand NAND4 (N6463, N6460, N4630, N4297, N6281);
nand NAND2 (N6464, N6462, N2550);
buf BUF1 (N6465, N6451);
nor NOR3 (N6466, N6456, N206, N4076);
nand NAND4 (N6467, N6464, N5836, N2282, N1689);
not NOT1 (N6468, N6431);
or OR3 (N6469, N6463, N3438, N4884);
buf BUF1 (N6470, N6469);
and AND3 (N6471, N6454, N5680, N931);
not NOT1 (N6472, N6466);
nor NOR4 (N6473, N6441, N2048, N4, N2374);
not NOT1 (N6474, N6468);
xor XOR2 (N6475, N6450, N5857);
not NOT1 (N6476, N6471);
or OR2 (N6477, N6459, N2284);
buf BUF1 (N6478, N6474);
buf BUF1 (N6479, N6477);
nor NOR4 (N6480, N6473, N5482, N6263, N3092);
xor XOR2 (N6481, N6467, N6057);
nand NAND2 (N6482, N6481, N998);
not NOT1 (N6483, N6475);
and AND4 (N6484, N6476, N3181, N4234, N72);
and AND2 (N6485, N6480, N2265);
and AND4 (N6486, N6458, N2610, N190, N1059);
and AND4 (N6487, N6485, N1230, N4594, N3935);
nand NAND2 (N6488, N6486, N3588);
buf BUF1 (N6489, N6484);
or OR2 (N6490, N6472, N2950);
and AND2 (N6491, N6483, N934);
and AND3 (N6492, N6491, N5999, N4338);
not NOT1 (N6493, N6492);
not NOT1 (N6494, N6488);
not NOT1 (N6495, N6490);
nor NOR2 (N6496, N6478, N6447);
or OR2 (N6497, N6493, N5587);
not NOT1 (N6498, N6479);
buf BUF1 (N6499, N6465);
not NOT1 (N6500, N6482);
or OR3 (N6501, N6494, N3142, N18);
xor XOR2 (N6502, N6470, N5495);
nor NOR3 (N6503, N6495, N5730, N147);
xor XOR2 (N6504, N6503, N3034);
buf BUF1 (N6505, N6502);
xor XOR2 (N6506, N6501, N117);
buf BUF1 (N6507, N6489);
or OR3 (N6508, N6499, N569, N1389);
xor XOR2 (N6509, N6504, N4315);
nor NOR4 (N6510, N6487, N790, N117, N1730);
nand NAND3 (N6511, N6498, N4421, N3380);
nor NOR4 (N6512, N6497, N1961, N3422, N456);
and AND3 (N6513, N6512, N6239, N4226);
and AND2 (N6514, N6507, N4431);
not NOT1 (N6515, N6508);
or OR3 (N6516, N6496, N413, N3129);
and AND2 (N6517, N6511, N3614);
xor XOR2 (N6518, N6500, N1277);
and AND2 (N6519, N6510, N1421);
not NOT1 (N6520, N6505);
buf BUF1 (N6521, N6517);
buf BUF1 (N6522, N6509);
or OR2 (N6523, N6519, N6140);
or OR3 (N6524, N6514, N6512, N2879);
xor XOR2 (N6525, N6523, N1735);
nor NOR3 (N6526, N6524, N3998, N4098);
and AND2 (N6527, N6525, N5650);
or OR2 (N6528, N6521, N6143);
or OR4 (N6529, N6518, N4548, N5395, N4452);
and AND3 (N6530, N6527, N59, N2179);
not NOT1 (N6531, N6513);
buf BUF1 (N6532, N6529);
buf BUF1 (N6533, N6522);
not NOT1 (N6534, N6515);
nand NAND4 (N6535, N6516, N4852, N5217, N546);
nand NAND2 (N6536, N6531, N3023);
nand NAND3 (N6537, N6506, N1225, N4235);
nand NAND3 (N6538, N6536, N4783, N4701);
and AND4 (N6539, N6528, N3045, N5072, N4758);
and AND3 (N6540, N6520, N2890, N1930);
buf BUF1 (N6541, N6534);
or OR2 (N6542, N6540, N1657);
buf BUF1 (N6543, N6526);
or OR3 (N6544, N6543, N38, N2774);
and AND3 (N6545, N6538, N2256, N2275);
not NOT1 (N6546, N6541);
nand NAND3 (N6547, N6539, N2513, N4885);
xor XOR2 (N6548, N6532, N2388);
buf BUF1 (N6549, N6544);
not NOT1 (N6550, N6542);
buf BUF1 (N6551, N6545);
nor NOR3 (N6552, N6548, N1617, N3784);
nand NAND2 (N6553, N6533, N5193);
xor XOR2 (N6554, N6549, N5215);
and AND4 (N6555, N6537, N3819, N5513, N3899);
nand NAND3 (N6556, N6551, N5923, N2696);
xor XOR2 (N6557, N6546, N3356);
xor XOR2 (N6558, N6556, N2228);
xor XOR2 (N6559, N6554, N6217);
nand NAND2 (N6560, N6547, N1771);
and AND4 (N6561, N6530, N3252, N6115, N1965);
nand NAND4 (N6562, N6559, N6247, N1766, N934);
nand NAND4 (N6563, N6562, N1237, N4381, N1722);
nor NOR4 (N6564, N6561, N113, N2315, N4557);
xor XOR2 (N6565, N6552, N4478);
buf BUF1 (N6566, N6553);
nand NAND3 (N6567, N6560, N5162, N1070);
buf BUF1 (N6568, N6565);
xor XOR2 (N6569, N6564, N3868);
or OR4 (N6570, N6550, N4668, N1455, N353);
xor XOR2 (N6571, N6567, N5941);
buf BUF1 (N6572, N6571);
or OR4 (N6573, N6535, N3722, N1449, N5918);
nor NOR4 (N6574, N6569, N2027, N5921, N3923);
or OR3 (N6575, N6568, N2715, N4819);
nor NOR4 (N6576, N6566, N3027, N5292, N1647);
xor XOR2 (N6577, N6572, N4314);
nor NOR4 (N6578, N6555, N4034, N768, N741);
xor XOR2 (N6579, N6570, N4076);
nand NAND3 (N6580, N6577, N1135, N1770);
nand NAND3 (N6581, N6573, N6182, N392);
not NOT1 (N6582, N6558);
buf BUF1 (N6583, N6580);
or OR2 (N6584, N6557, N1319);
nand NAND4 (N6585, N6583, N6441, N1695, N2652);
not NOT1 (N6586, N6563);
or OR2 (N6587, N6576, N2716);
nand NAND2 (N6588, N6584, N6371);
not NOT1 (N6589, N6585);
and AND2 (N6590, N6575, N3919);
nor NOR2 (N6591, N6586, N2680);
not NOT1 (N6592, N6581);
nand NAND3 (N6593, N6590, N2322, N2757);
buf BUF1 (N6594, N6592);
nand NAND4 (N6595, N6578, N1228, N1413, N581);
nand NAND4 (N6596, N6587, N6172, N3004, N6302);
and AND2 (N6597, N6589, N930);
xor XOR2 (N6598, N6574, N425);
xor XOR2 (N6599, N6597, N5495);
buf BUF1 (N6600, N6591);
not NOT1 (N6601, N6593);
and AND3 (N6602, N6601, N3877, N2179);
and AND4 (N6603, N6595, N4642, N340, N964);
not NOT1 (N6604, N6588);
buf BUF1 (N6605, N6600);
xor XOR2 (N6606, N6596, N2383);
nand NAND2 (N6607, N6604, N4335);
nand NAND2 (N6608, N6582, N3646);
buf BUF1 (N6609, N6606);
nor NOR2 (N6610, N6579, N1541);
or OR2 (N6611, N6607, N4139);
xor XOR2 (N6612, N6598, N2548);
nand NAND2 (N6613, N6608, N3587);
nor NOR2 (N6614, N6594, N4514);
nand NAND3 (N6615, N6614, N228, N3699);
nor NOR4 (N6616, N6610, N6149, N5965, N5452);
xor XOR2 (N6617, N6605, N2172);
and AND3 (N6618, N6611, N4140, N4676);
nor NOR4 (N6619, N6616, N4049, N6417, N3031);
not NOT1 (N6620, N6615);
or OR3 (N6621, N6609, N2516, N4646);
nor NOR2 (N6622, N6618, N3541);
nand NAND2 (N6623, N6602, N1971);
not NOT1 (N6624, N6599);
not NOT1 (N6625, N6603);
nand NAND4 (N6626, N6623, N3900, N104, N1228);
nand NAND2 (N6627, N6626, N2470);
and AND2 (N6628, N6624, N4820);
xor XOR2 (N6629, N6627, N6609);
xor XOR2 (N6630, N6612, N2448);
nor NOR4 (N6631, N6621, N1296, N5033, N1859);
not NOT1 (N6632, N6628);
nand NAND3 (N6633, N6617, N99, N5095);
nor NOR2 (N6634, N6619, N673);
not NOT1 (N6635, N6631);
not NOT1 (N6636, N6632);
not NOT1 (N6637, N6634);
or OR4 (N6638, N6622, N5264, N3351, N3278);
xor XOR2 (N6639, N6620, N3454);
or OR4 (N6640, N6633, N761, N5658, N1109);
and AND2 (N6641, N6638, N1076);
nor NOR4 (N6642, N6637, N228, N4465, N951);
nor NOR4 (N6643, N6636, N5190, N3834, N5739);
nor NOR2 (N6644, N6643, N4252);
or OR2 (N6645, N6644, N5407);
nor NOR4 (N6646, N6639, N5658, N2547, N5778);
nand NAND3 (N6647, N6640, N2298, N942);
or OR2 (N6648, N6613, N3916);
not NOT1 (N6649, N6647);
not NOT1 (N6650, N6646);
xor XOR2 (N6651, N6629, N2427);
xor XOR2 (N6652, N6635, N5505);
xor XOR2 (N6653, N6630, N6438);
nand NAND3 (N6654, N6625, N5688, N2197);
or OR4 (N6655, N6653, N3093, N4592, N6109);
buf BUF1 (N6656, N6642);
xor XOR2 (N6657, N6648, N5885);
and AND2 (N6658, N6645, N3333);
nor NOR2 (N6659, N6656, N2400);
not NOT1 (N6660, N6657);
xor XOR2 (N6661, N6651, N2445);
xor XOR2 (N6662, N6659, N1891);
and AND2 (N6663, N6661, N4206);
and AND4 (N6664, N6654, N2482, N5045, N4724);
nand NAND3 (N6665, N6664, N4133, N179);
and AND2 (N6666, N6641, N3916);
xor XOR2 (N6667, N6652, N1967);
and AND3 (N6668, N6665, N2866, N224);
or OR4 (N6669, N6649, N4546, N1430, N679);
or OR4 (N6670, N6660, N843, N2846, N3638);
nor NOR4 (N6671, N6667, N2306, N4673, N457);
buf BUF1 (N6672, N6655);
or OR3 (N6673, N6671, N6363, N487);
nand NAND3 (N6674, N6668, N5876, N5477);
nand NAND4 (N6675, N6658, N2316, N4104, N6249);
buf BUF1 (N6676, N6650);
or OR2 (N6677, N6672, N3344);
not NOT1 (N6678, N6676);
nand NAND2 (N6679, N6674, N5960);
nand NAND4 (N6680, N6678, N4025, N2919, N838);
nor NOR3 (N6681, N6679, N1218, N2725);
and AND4 (N6682, N6666, N3107, N2496, N3026);
and AND3 (N6683, N6663, N887, N6039);
and AND3 (N6684, N6669, N523, N1062);
or OR3 (N6685, N6673, N926, N2323);
nand NAND3 (N6686, N6681, N5259, N3937);
nor NOR2 (N6687, N6684, N906);
nor NOR2 (N6688, N6662, N320);
xor XOR2 (N6689, N6688, N6479);
nand NAND4 (N6690, N6687, N2005, N3658, N1199);
xor XOR2 (N6691, N6689, N2394);
and AND4 (N6692, N6670, N3303, N6377, N2021);
not NOT1 (N6693, N6691);
and AND4 (N6694, N6683, N3230, N2510, N4396);
not NOT1 (N6695, N6680);
nor NOR4 (N6696, N6686, N1550, N6459, N1350);
or OR2 (N6697, N6696, N1819);
xor XOR2 (N6698, N6685, N6024);
xor XOR2 (N6699, N6692, N1917);
or OR2 (N6700, N6698, N2736);
not NOT1 (N6701, N6700);
and AND3 (N6702, N6699, N4660, N6468);
and AND2 (N6703, N6675, N6408);
and AND4 (N6704, N6682, N6174, N6161, N3425);
buf BUF1 (N6705, N6702);
or OR2 (N6706, N6677, N5761);
not NOT1 (N6707, N6706);
nand NAND3 (N6708, N6697, N4774, N5945);
not NOT1 (N6709, N6705);
and AND2 (N6710, N6695, N2838);
nand NAND2 (N6711, N6710, N3914);
xor XOR2 (N6712, N6704, N6140);
not NOT1 (N6713, N6703);
nand NAND2 (N6714, N6701, N3222);
nor NOR4 (N6715, N6694, N6648, N3719, N3145);
not NOT1 (N6716, N6713);
or OR4 (N6717, N6690, N5544, N3866, N6080);
buf BUF1 (N6718, N6716);
or OR4 (N6719, N6707, N6060, N2837, N2899);
not NOT1 (N6720, N6693);
nor NOR2 (N6721, N6717, N4796);
xor XOR2 (N6722, N6720, N5807);
xor XOR2 (N6723, N6722, N5426);
xor XOR2 (N6724, N6718, N4682);
not NOT1 (N6725, N6712);
or OR2 (N6726, N6708, N4287);
xor XOR2 (N6727, N6723, N3546);
or OR4 (N6728, N6711, N2525, N206, N1300);
and AND2 (N6729, N6727, N4410);
nor NOR4 (N6730, N6725, N6254, N6098, N698);
xor XOR2 (N6731, N6719, N2251);
not NOT1 (N6732, N6721);
xor XOR2 (N6733, N6731, N4590);
buf BUF1 (N6734, N6714);
nor NOR4 (N6735, N6733, N5538, N3169, N4096);
xor XOR2 (N6736, N6728, N1911);
and AND3 (N6737, N6734, N516, N1585);
not NOT1 (N6738, N6735);
or OR2 (N6739, N6737, N4508);
and AND4 (N6740, N6715, N2121, N4747, N485);
buf BUF1 (N6741, N6709);
not NOT1 (N6742, N6732);
and AND4 (N6743, N6730, N1928, N5507, N5326);
xor XOR2 (N6744, N6742, N2681);
or OR4 (N6745, N6724, N395, N3354, N157);
buf BUF1 (N6746, N6743);
and AND4 (N6747, N6729, N5355, N1766, N1017);
or OR4 (N6748, N6739, N5202, N431, N4844);
buf BUF1 (N6749, N6736);
and AND2 (N6750, N6747, N1821);
nand NAND4 (N6751, N6740, N1321, N2505, N3423);
buf BUF1 (N6752, N6745);
and AND4 (N6753, N6741, N1091, N2519, N5014);
or OR4 (N6754, N6749, N2577, N923, N5426);
nor NOR3 (N6755, N6752, N5532, N1324);
buf BUF1 (N6756, N6748);
not NOT1 (N6757, N6755);
not NOT1 (N6758, N6746);
xor XOR2 (N6759, N6756, N1441);
and AND4 (N6760, N6751, N4846, N6404, N5965);
not NOT1 (N6761, N6757);
buf BUF1 (N6762, N6761);
or OR2 (N6763, N6759, N6287);
nor NOR4 (N6764, N6744, N3559, N2299, N4505);
buf BUF1 (N6765, N6762);
nand NAND3 (N6766, N6754, N6545, N3641);
buf BUF1 (N6767, N6738);
nor NOR3 (N6768, N6767, N1480, N1548);
or OR4 (N6769, N6766, N2506, N838, N4152);
or OR2 (N6770, N6763, N6768);
xor XOR2 (N6771, N1346, N3349);
xor XOR2 (N6772, N6726, N2015);
nand NAND3 (N6773, N6753, N1621, N1422);
xor XOR2 (N6774, N6758, N3183);
nor NOR4 (N6775, N6770, N3970, N5134, N6144);
nand NAND3 (N6776, N6775, N2036, N78);
nand NAND4 (N6777, N6771, N73, N2643, N4616);
xor XOR2 (N6778, N6776, N3909);
buf BUF1 (N6779, N6778);
not NOT1 (N6780, N6772);
and AND2 (N6781, N6764, N5196);
and AND3 (N6782, N6760, N87, N4219);
or OR4 (N6783, N6773, N846, N3065, N1921);
or OR4 (N6784, N6781, N2701, N513, N6124);
or OR4 (N6785, N6765, N5963, N3101, N394);
or OR4 (N6786, N6782, N1535, N1262, N5135);
nand NAND3 (N6787, N6774, N3311, N5696);
not NOT1 (N6788, N6785);
nor NOR4 (N6789, N6783, N6064, N406, N16);
buf BUF1 (N6790, N6786);
nand NAND3 (N6791, N6784, N928, N883);
or OR2 (N6792, N6787, N3621);
not NOT1 (N6793, N6780);
xor XOR2 (N6794, N6790, N6721);
buf BUF1 (N6795, N6791);
or OR4 (N6796, N6779, N1353, N1378, N962);
nand NAND3 (N6797, N6769, N145, N1362);
nor NOR3 (N6798, N6788, N4178, N114);
and AND2 (N6799, N6792, N1982);
or OR3 (N6800, N6793, N4513, N622);
or OR4 (N6801, N6795, N2319, N642, N6384);
and AND4 (N6802, N6798, N2131, N4955, N3081);
not NOT1 (N6803, N6796);
nor NOR2 (N6804, N6794, N5584);
and AND4 (N6805, N6777, N3455, N5100, N763);
or OR4 (N6806, N6800, N5431, N1902, N3216);
buf BUF1 (N6807, N6803);
nor NOR4 (N6808, N6807, N5334, N1452, N6090);
and AND4 (N6809, N6789, N2047, N4237, N108);
and AND2 (N6810, N6797, N2069);
or OR3 (N6811, N6801, N2192, N639);
not NOT1 (N6812, N6804);
not NOT1 (N6813, N6811);
buf BUF1 (N6814, N6808);
not NOT1 (N6815, N6809);
and AND2 (N6816, N6805, N5198);
buf BUF1 (N6817, N6799);
and AND3 (N6818, N6750, N2473, N5022);
and AND2 (N6819, N6812, N5092);
xor XOR2 (N6820, N6817, N3551);
nand NAND2 (N6821, N6815, N6371);
not NOT1 (N6822, N6818);
not NOT1 (N6823, N6802);
xor XOR2 (N6824, N6821, N1184);
and AND2 (N6825, N6822, N234);
not NOT1 (N6826, N6825);
xor XOR2 (N6827, N6814, N996);
xor XOR2 (N6828, N6819, N1769);
xor XOR2 (N6829, N6828, N1501);
not NOT1 (N6830, N6810);
nor NOR4 (N6831, N6823, N1280, N2483, N1107);
and AND2 (N6832, N6816, N6485);
nand NAND2 (N6833, N6832, N6479);
and AND3 (N6834, N6826, N422, N2769);
xor XOR2 (N6835, N6820, N2043);
not NOT1 (N6836, N6806);
or OR4 (N6837, N6827, N2834, N3105, N3528);
nand NAND2 (N6838, N6835, N5878);
xor XOR2 (N6839, N6837, N6674);
buf BUF1 (N6840, N6824);
nor NOR3 (N6841, N6833, N5186, N3811);
xor XOR2 (N6842, N6830, N3931);
nand NAND4 (N6843, N6838, N6708, N875, N3307);
xor XOR2 (N6844, N6842, N3243);
or OR3 (N6845, N6840, N2368, N2748);
buf BUF1 (N6846, N6841);
buf BUF1 (N6847, N6834);
not NOT1 (N6848, N6836);
and AND3 (N6849, N6845, N6161, N4657);
or OR2 (N6850, N6839, N5978);
buf BUF1 (N6851, N6831);
or OR4 (N6852, N6846, N450, N6252, N809);
not NOT1 (N6853, N6813);
and AND2 (N6854, N6851, N2790);
and AND2 (N6855, N6853, N5724);
nand NAND4 (N6856, N6843, N5749, N5244, N4419);
xor XOR2 (N6857, N6852, N2563);
not NOT1 (N6858, N6829);
and AND2 (N6859, N6850, N4331);
xor XOR2 (N6860, N6857, N3924);
buf BUF1 (N6861, N6847);
nor NOR4 (N6862, N6854, N872, N4819, N1229);
buf BUF1 (N6863, N6855);
and AND4 (N6864, N6859, N3546, N5993, N2375);
or OR4 (N6865, N6861, N1559, N3136, N145);
nor NOR3 (N6866, N6858, N2129, N2929);
and AND2 (N6867, N6848, N3865);
buf BUF1 (N6868, N6864);
xor XOR2 (N6869, N6866, N4790);
or OR4 (N6870, N6844, N19, N5992, N147);
and AND3 (N6871, N6869, N3950, N2447);
or OR3 (N6872, N6856, N1803, N6862);
nand NAND2 (N6873, N3939, N4704);
buf BUF1 (N6874, N6849);
xor XOR2 (N6875, N6872, N2042);
nor NOR4 (N6876, N6867, N89, N237, N1003);
and AND2 (N6877, N6874, N1608);
or OR4 (N6878, N6871, N1665, N919, N5026);
nor NOR2 (N6879, N6877, N1432);
nor NOR3 (N6880, N6863, N1305, N3482);
nand NAND3 (N6881, N6870, N5392, N6229);
buf BUF1 (N6882, N6875);
nand NAND4 (N6883, N6880, N5622, N5990, N6598);
buf BUF1 (N6884, N6868);
not NOT1 (N6885, N6876);
xor XOR2 (N6886, N6878, N6533);
nor NOR4 (N6887, N6865, N489, N571, N2668);
nor NOR2 (N6888, N6884, N1819);
or OR4 (N6889, N6887, N43, N155, N248);
buf BUF1 (N6890, N6879);
buf BUF1 (N6891, N6886);
nor NOR3 (N6892, N6873, N771, N5118);
and AND2 (N6893, N6883, N1944);
buf BUF1 (N6894, N6893);
buf BUF1 (N6895, N6891);
nor NOR3 (N6896, N6888, N706, N6861);
nand NAND2 (N6897, N6889, N2151);
nand NAND4 (N6898, N6882, N3605, N803, N4519);
or OR3 (N6899, N6885, N4869, N1652);
or OR2 (N6900, N6881, N2060);
xor XOR2 (N6901, N6899, N1671);
or OR4 (N6902, N6896, N5105, N2515, N272);
xor XOR2 (N6903, N6900, N6846);
buf BUF1 (N6904, N6898);
xor XOR2 (N6905, N6903, N2972);
and AND3 (N6906, N6901, N6645, N6500);
nor NOR2 (N6907, N6890, N1771);
and AND4 (N6908, N6860, N4219, N1963, N2971);
not NOT1 (N6909, N6902);
buf BUF1 (N6910, N6894);
buf BUF1 (N6911, N6897);
buf BUF1 (N6912, N6911);
nand NAND2 (N6913, N6895, N5511);
not NOT1 (N6914, N6892);
and AND2 (N6915, N6905, N6440);
not NOT1 (N6916, N6912);
xor XOR2 (N6917, N6904, N2421);
and AND3 (N6918, N6906, N5040, N3108);
not NOT1 (N6919, N6907);
buf BUF1 (N6920, N6919);
xor XOR2 (N6921, N6908, N2376);
buf BUF1 (N6922, N6921);
buf BUF1 (N6923, N6913);
or OR2 (N6924, N6915, N1789);
not NOT1 (N6925, N6922);
buf BUF1 (N6926, N6925);
and AND4 (N6927, N6926, N3679, N4276, N5630);
buf BUF1 (N6928, N6914);
buf BUF1 (N6929, N6924);
not NOT1 (N6930, N6928);
not NOT1 (N6931, N6910);
nor NOR2 (N6932, N6909, N3277);
nand NAND2 (N6933, N6929, N3448);
buf BUF1 (N6934, N6920);
buf BUF1 (N6935, N6934);
nand NAND2 (N6936, N6917, N6147);
nor NOR3 (N6937, N6918, N3143, N3118);
buf BUF1 (N6938, N6916);
or OR3 (N6939, N6932, N3742, N4124);
nand NAND2 (N6940, N6935, N6784);
nand NAND3 (N6941, N6933, N40, N6608);
buf BUF1 (N6942, N6941);
not NOT1 (N6943, N6939);
or OR2 (N6944, N6938, N3371);
buf BUF1 (N6945, N6930);
nor NOR4 (N6946, N6944, N4606, N3293, N4676);
not NOT1 (N6947, N6936);
or OR4 (N6948, N6923, N4528, N4789, N2631);
nand NAND2 (N6949, N6946, N2859);
nor NOR2 (N6950, N6948, N3468);
or OR3 (N6951, N6942, N2884, N5000);
buf BUF1 (N6952, N6940);
buf BUF1 (N6953, N6952);
xor XOR2 (N6954, N6950, N4846);
nand NAND2 (N6955, N6943, N3068);
or OR2 (N6956, N6953, N638);
buf BUF1 (N6957, N6954);
or OR4 (N6958, N6945, N1233, N321, N6775);
nor NOR4 (N6959, N6957, N35, N541, N5526);
and AND2 (N6960, N6949, N1295);
xor XOR2 (N6961, N6937, N4260);
or OR2 (N6962, N6958, N2325);
buf BUF1 (N6963, N6961);
nor NOR2 (N6964, N6931, N3061);
nand NAND2 (N6965, N6927, N1091);
nand NAND3 (N6966, N6951, N5497, N3594);
xor XOR2 (N6967, N6963, N2645);
and AND4 (N6968, N6955, N5620, N2333, N297);
nand NAND4 (N6969, N6960, N4885, N5108, N6037);
or OR3 (N6970, N6967, N1924, N6108);
xor XOR2 (N6971, N6970, N402);
not NOT1 (N6972, N6956);
xor XOR2 (N6973, N6962, N2392);
nand NAND4 (N6974, N6966, N5113, N2501, N1415);
nand NAND2 (N6975, N6973, N4972);
nand NAND3 (N6976, N6947, N1865, N4872);
nand NAND2 (N6977, N6959, N4525);
xor XOR2 (N6978, N6974, N2684);
buf BUF1 (N6979, N6965);
or OR4 (N6980, N6971, N4010, N4698, N4302);
not NOT1 (N6981, N6977);
buf BUF1 (N6982, N6975);
nand NAND4 (N6983, N6981, N3924, N488, N3333);
nor NOR2 (N6984, N6976, N1656);
xor XOR2 (N6985, N6979, N1859);
not NOT1 (N6986, N6978);
not NOT1 (N6987, N6985);
and AND2 (N6988, N6982, N6589);
or OR3 (N6989, N6964, N6581, N6562);
xor XOR2 (N6990, N6980, N1403);
buf BUF1 (N6991, N6968);
xor XOR2 (N6992, N6984, N889);
nand NAND4 (N6993, N6972, N5555, N2630, N337);
nand NAND2 (N6994, N6992, N6148);
or OR4 (N6995, N6993, N105, N5715, N6085);
not NOT1 (N6996, N6969);
nor NOR2 (N6997, N6991, N445);
nor NOR2 (N6998, N6996, N991);
not NOT1 (N6999, N6987);
nand NAND3 (N7000, N6989, N3039, N6862);
or OR2 (N7001, N6998, N5415);
not NOT1 (N7002, N6990);
not NOT1 (N7003, N6994);
not NOT1 (N7004, N6983);
nor NOR4 (N7005, N7004, N6084, N4911, N1518);
xor XOR2 (N7006, N6999, N3415);
and AND4 (N7007, N7005, N1787, N5909, N5645);
or OR2 (N7008, N6986, N6140);
nand NAND2 (N7009, N7001, N5217);
xor XOR2 (N7010, N7006, N1596);
nand NAND2 (N7011, N6995, N6570);
and AND4 (N7012, N7008, N6021, N1582, N604);
or OR3 (N7013, N7007, N1852, N937);
or OR2 (N7014, N6988, N5810);
buf BUF1 (N7015, N7010);
and AND4 (N7016, N7011, N823, N4790, N3181);
or OR4 (N7017, N6997, N6370, N1682, N2107);
nor NOR3 (N7018, N7002, N2235, N1271);
buf BUF1 (N7019, N7003);
buf BUF1 (N7020, N7013);
not NOT1 (N7021, N7020);
and AND2 (N7022, N7016, N6114);
xor XOR2 (N7023, N7015, N294);
not NOT1 (N7024, N7018);
not NOT1 (N7025, N7014);
nand NAND4 (N7026, N7000, N313, N5361, N4881);
or OR2 (N7027, N7025, N3029);
and AND3 (N7028, N7021, N3907, N3653);
nor NOR2 (N7029, N7009, N5851);
buf BUF1 (N7030, N7024);
xor XOR2 (N7031, N7029, N3890);
or OR4 (N7032, N7023, N2309, N4654, N6110);
not NOT1 (N7033, N7032);
nand NAND4 (N7034, N7027, N5121, N6503, N5977);
or OR3 (N7035, N7012, N1610, N1585);
not NOT1 (N7036, N7035);
not NOT1 (N7037, N7028);
buf BUF1 (N7038, N7019);
xor XOR2 (N7039, N7038, N5922);
nand NAND3 (N7040, N7017, N3695, N1393);
nor NOR4 (N7041, N7037, N6100, N2025, N1572);
nor NOR3 (N7042, N7030, N414, N4804);
xor XOR2 (N7043, N7042, N4748);
or OR3 (N7044, N7031, N1218, N144);
buf BUF1 (N7045, N7044);
xor XOR2 (N7046, N7034, N2397);
buf BUF1 (N7047, N7043);
or OR4 (N7048, N7036, N3927, N4016, N446);
buf BUF1 (N7049, N7045);
nor NOR2 (N7050, N7026, N5211);
and AND3 (N7051, N7040, N6063, N178);
buf BUF1 (N7052, N7050);
nor NOR2 (N7053, N7052, N520);
xor XOR2 (N7054, N7046, N6772);
not NOT1 (N7055, N7051);
nand NAND3 (N7056, N7033, N1105, N6023);
xor XOR2 (N7057, N7041, N1183);
buf BUF1 (N7058, N7057);
or OR4 (N7059, N7049, N5909, N861, N5017);
not NOT1 (N7060, N7039);
or OR3 (N7061, N7056, N6297, N6106);
xor XOR2 (N7062, N7059, N922);
nand NAND3 (N7063, N7054, N2006, N6596);
not NOT1 (N7064, N7048);
not NOT1 (N7065, N7060);
nand NAND2 (N7066, N7053, N436);
nor NOR3 (N7067, N7061, N4675, N5776);
nand NAND2 (N7068, N7066, N510);
and AND4 (N7069, N7022, N4912, N5218, N1895);
nor NOR4 (N7070, N7068, N5847, N4623, N4462);
xor XOR2 (N7071, N7047, N1564);
or OR4 (N7072, N7065, N665, N1915, N4553);
not NOT1 (N7073, N7058);
not NOT1 (N7074, N7069);
or OR2 (N7075, N7071, N23);
and AND4 (N7076, N7062, N5131, N5303, N6949);
xor XOR2 (N7077, N7072, N892);
nor NOR4 (N7078, N7063, N2455, N3414, N2825);
not NOT1 (N7079, N7073);
nor NOR2 (N7080, N7067, N2336);
and AND4 (N7081, N7055, N4638, N632, N1704);
or OR3 (N7082, N7078, N6323, N2097);
nand NAND4 (N7083, N7070, N5831, N5359, N5493);
nor NOR2 (N7084, N7074, N1927);
buf BUF1 (N7085, N7075);
not NOT1 (N7086, N7079);
not NOT1 (N7087, N7064);
xor XOR2 (N7088, N7077, N6935);
nand NAND4 (N7089, N7087, N5787, N5702, N3988);
not NOT1 (N7090, N7082);
nand NAND3 (N7091, N7081, N6019, N1651);
or OR3 (N7092, N7089, N2980, N5680);
or OR3 (N7093, N7076, N4815, N3526);
not NOT1 (N7094, N7085);
xor XOR2 (N7095, N7092, N6051);
buf BUF1 (N7096, N7086);
or OR4 (N7097, N7096, N6811, N1856, N957);
xor XOR2 (N7098, N7097, N6931);
not NOT1 (N7099, N7083);
buf BUF1 (N7100, N7095);
nand NAND2 (N7101, N7098, N3542);
nor NOR4 (N7102, N7084, N839, N4989, N6511);
nand NAND3 (N7103, N7094, N6387, N2649);
and AND2 (N7104, N7100, N1783);
or OR3 (N7105, N7093, N3008, N706);
buf BUF1 (N7106, N7102);
or OR3 (N7107, N7099, N2677, N444);
and AND4 (N7108, N7103, N7104, N2420, N614);
and AND4 (N7109, N5427, N3749, N1114, N3794);
nor NOR3 (N7110, N7108, N367, N5394);
nand NAND3 (N7111, N7101, N492, N961);
buf BUF1 (N7112, N7080);
xor XOR2 (N7113, N7106, N1995);
not NOT1 (N7114, N7113);
buf BUF1 (N7115, N7110);
buf BUF1 (N7116, N7114);
or OR4 (N7117, N7115, N119, N4209, N3757);
nand NAND4 (N7118, N7112, N4297, N1924, N6849);
nor NOR4 (N7119, N7109, N670, N5764, N2453);
or OR4 (N7120, N7119, N6803, N4375, N4066);
and AND4 (N7121, N7105, N6819, N5485, N1588);
nor NOR3 (N7122, N7117, N3679, N3477);
and AND2 (N7123, N7088, N1914);
and AND2 (N7124, N7121, N2833);
and AND2 (N7125, N7091, N5881);
nand NAND4 (N7126, N7122, N3836, N3204, N4479);
and AND3 (N7127, N7090, N6993, N6668);
buf BUF1 (N7128, N7118);
or OR4 (N7129, N7125, N4198, N6227, N2931);
not NOT1 (N7130, N7129);
not NOT1 (N7131, N7111);
not NOT1 (N7132, N7107);
or OR2 (N7133, N7116, N1824);
buf BUF1 (N7134, N7126);
or OR2 (N7135, N7131, N3998);
or OR4 (N7136, N7120, N6511, N957, N6369);
xor XOR2 (N7137, N7132, N5298);
not NOT1 (N7138, N7130);
buf BUF1 (N7139, N7138);
not NOT1 (N7140, N7123);
xor XOR2 (N7141, N7124, N3996);
nand NAND2 (N7142, N7139, N2428);
nor NOR3 (N7143, N7133, N4375, N6194);
nand NAND3 (N7144, N7134, N472, N2463);
or OR4 (N7145, N7127, N2936, N1922, N6428);
not NOT1 (N7146, N7137);
not NOT1 (N7147, N7142);
xor XOR2 (N7148, N7136, N3698);
not NOT1 (N7149, N7147);
nand NAND2 (N7150, N7128, N2065);
buf BUF1 (N7151, N7143);
xor XOR2 (N7152, N7135, N6313);
xor XOR2 (N7153, N7150, N2713);
nand NAND3 (N7154, N7148, N6714, N3830);
nand NAND4 (N7155, N7144, N337, N3189, N1173);
xor XOR2 (N7156, N7153, N6498);
not NOT1 (N7157, N7151);
or OR4 (N7158, N7156, N2578, N4273, N5850);
nor NOR3 (N7159, N7157, N2500, N1673);
nor NOR2 (N7160, N7140, N4843);
nor NOR2 (N7161, N7145, N2103);
and AND4 (N7162, N7161, N1987, N3339, N1840);
buf BUF1 (N7163, N7141);
buf BUF1 (N7164, N7163);
buf BUF1 (N7165, N7164);
nor NOR3 (N7166, N7152, N1752, N4851);
xor XOR2 (N7167, N7166, N4308);
xor XOR2 (N7168, N7162, N2593);
xor XOR2 (N7169, N7167, N6791);
or OR3 (N7170, N7169, N4388, N5460);
not NOT1 (N7171, N7146);
not NOT1 (N7172, N7165);
and AND2 (N7173, N7168, N520);
nor NOR3 (N7174, N7173, N598, N6621);
buf BUF1 (N7175, N7172);
and AND4 (N7176, N7170, N4643, N30, N1378);
buf BUF1 (N7177, N7159);
and AND2 (N7178, N7174, N5411);
buf BUF1 (N7179, N7154);
and AND4 (N7180, N7171, N5097, N5159, N71);
nor NOR4 (N7181, N7178, N807, N3890, N5896);
nand NAND2 (N7182, N7160, N4778);
not NOT1 (N7183, N7179);
nand NAND4 (N7184, N7182, N933, N3762, N5125);
nand NAND3 (N7185, N7149, N6500, N4184);
nor NOR4 (N7186, N7177, N2955, N1549, N1948);
xor XOR2 (N7187, N7183, N3880);
and AND2 (N7188, N7180, N5825);
nor NOR3 (N7189, N7187, N3729, N5828);
and AND2 (N7190, N7155, N4164);
and AND3 (N7191, N7190, N2794, N112);
xor XOR2 (N7192, N7175, N6079);
not NOT1 (N7193, N7189);
nand NAND4 (N7194, N7181, N6929, N2643, N709);
not NOT1 (N7195, N7158);
or OR2 (N7196, N7191, N4772);
buf BUF1 (N7197, N7192);
buf BUF1 (N7198, N7184);
not NOT1 (N7199, N7193);
xor XOR2 (N7200, N7198, N3524);
not NOT1 (N7201, N7200);
buf BUF1 (N7202, N7197);
or OR4 (N7203, N7176, N906, N6616, N465);
xor XOR2 (N7204, N7203, N4233);
buf BUF1 (N7205, N7201);
buf BUF1 (N7206, N7185);
not NOT1 (N7207, N7196);
xor XOR2 (N7208, N7199, N5466);
and AND2 (N7209, N7194, N6742);
or OR2 (N7210, N7186, N4983);
buf BUF1 (N7211, N7188);
xor XOR2 (N7212, N7208, N1851);
nand NAND2 (N7213, N7206, N4456);
xor XOR2 (N7214, N7202, N1430);
and AND2 (N7215, N7209, N6416);
or OR2 (N7216, N7195, N3139);
nand NAND4 (N7217, N7210, N3533, N2509, N546);
or OR2 (N7218, N7216, N2094);
and AND4 (N7219, N7207, N4600, N3943, N2295);
not NOT1 (N7220, N7214);
xor XOR2 (N7221, N7215, N3114);
or OR4 (N7222, N7204, N2662, N6072, N2794);
nor NOR2 (N7223, N7220, N5962);
nor NOR2 (N7224, N7213, N849);
not NOT1 (N7225, N7218);
and AND4 (N7226, N7211, N213, N6341, N3752);
and AND4 (N7227, N7217, N3658, N6491, N1144);
not NOT1 (N7228, N7225);
xor XOR2 (N7229, N7227, N878);
xor XOR2 (N7230, N7205, N6130);
nor NOR4 (N7231, N7223, N2730, N5546, N5362);
xor XOR2 (N7232, N7226, N5550);
not NOT1 (N7233, N7232);
not NOT1 (N7234, N7221);
and AND4 (N7235, N7212, N586, N1531, N3671);
nor NOR2 (N7236, N7235, N1617);
and AND2 (N7237, N7236, N260);
nor NOR2 (N7238, N7222, N3492);
not NOT1 (N7239, N7228);
nand NAND4 (N7240, N7224, N1210, N6820, N535);
nand NAND3 (N7241, N7230, N5580, N3485);
xor XOR2 (N7242, N7241, N973);
not NOT1 (N7243, N7238);
buf BUF1 (N7244, N7219);
xor XOR2 (N7245, N7231, N4068);
or OR2 (N7246, N7244, N5069);
or OR3 (N7247, N7233, N3524, N2110);
nor NOR2 (N7248, N7247, N1571);
nand NAND3 (N7249, N7248, N6077, N2892);
and AND4 (N7250, N7229, N2073, N5363, N268);
xor XOR2 (N7251, N7243, N7196);
nor NOR3 (N7252, N7242, N2795, N2241);
nand NAND4 (N7253, N7245, N2626, N4481, N714);
and AND3 (N7254, N7251, N4374, N5559);
buf BUF1 (N7255, N7250);
nor NOR4 (N7256, N7249, N4314, N4697, N4882);
xor XOR2 (N7257, N7240, N633);
buf BUF1 (N7258, N7237);
buf BUF1 (N7259, N7255);
xor XOR2 (N7260, N7239, N71);
nand NAND2 (N7261, N7246, N1168);
nand NAND4 (N7262, N7261, N5501, N145, N6065);
xor XOR2 (N7263, N7256, N5414);
xor XOR2 (N7264, N7257, N2243);
nand NAND2 (N7265, N7260, N5150);
not NOT1 (N7266, N7265);
nand NAND3 (N7267, N7252, N4262, N5922);
nor NOR2 (N7268, N7267, N4728);
nand NAND3 (N7269, N7258, N1422, N2867);
xor XOR2 (N7270, N7268, N5306);
and AND3 (N7271, N7234, N2545, N2429);
buf BUF1 (N7272, N7266);
or OR4 (N7273, N7263, N4685, N6904, N5883);
nand NAND2 (N7274, N7269, N5177);
or OR3 (N7275, N7273, N216, N2264);
nor NOR3 (N7276, N7264, N5218, N6672);
not NOT1 (N7277, N7254);
xor XOR2 (N7278, N7272, N2136);
nand NAND3 (N7279, N7270, N619, N1511);
nand NAND3 (N7280, N7274, N6904, N6060);
or OR3 (N7281, N7279, N3288, N2465);
xor XOR2 (N7282, N7280, N2592);
and AND3 (N7283, N7253, N4634, N6698);
nor NOR2 (N7284, N7275, N1614);
and AND3 (N7285, N7271, N3916, N3319);
xor XOR2 (N7286, N7277, N2276);
not NOT1 (N7287, N7285);
nand NAND4 (N7288, N7287, N4350, N4924, N3749);
nand NAND2 (N7289, N7281, N3655);
and AND3 (N7290, N7259, N6815, N6325);
and AND2 (N7291, N7262, N4418);
xor XOR2 (N7292, N7276, N1464);
buf BUF1 (N7293, N7288);
not NOT1 (N7294, N7291);
nand NAND3 (N7295, N7292, N6921, N4371);
or OR3 (N7296, N7294, N5417, N7238);
xor XOR2 (N7297, N7290, N6194);
xor XOR2 (N7298, N7286, N3759);
buf BUF1 (N7299, N7296);
or OR4 (N7300, N7278, N5647, N708, N1906);
and AND4 (N7301, N7284, N4934, N4292, N3724);
xor XOR2 (N7302, N7301, N4370);
nand NAND4 (N7303, N7300, N2247, N948, N4713);
not NOT1 (N7304, N7303);
xor XOR2 (N7305, N7282, N2285);
nand NAND3 (N7306, N7297, N7185, N6562);
not NOT1 (N7307, N7293);
not NOT1 (N7308, N7305);
or OR3 (N7309, N7283, N6194, N3155);
or OR2 (N7310, N7299, N6523);
nor NOR4 (N7311, N7307, N3323, N84, N666);
xor XOR2 (N7312, N7308, N4512);
and AND2 (N7313, N7289, N7281);
and AND4 (N7314, N7306, N3187, N2838, N6031);
xor XOR2 (N7315, N7310, N203);
and AND3 (N7316, N7311, N3843, N587);
nor NOR3 (N7317, N7314, N1755, N4161);
buf BUF1 (N7318, N7302);
xor XOR2 (N7319, N7316, N4497);
nor NOR4 (N7320, N7298, N2148, N6582, N7294);
buf BUF1 (N7321, N7313);
or OR3 (N7322, N7321, N319, N4119);
buf BUF1 (N7323, N7322);
or OR2 (N7324, N7317, N5038);
nor NOR4 (N7325, N7320, N6941, N4936, N3014);
nand NAND4 (N7326, N7312, N5403, N6627, N7098);
buf BUF1 (N7327, N7309);
or OR4 (N7328, N7327, N1056, N2626, N1582);
nand NAND2 (N7329, N7295, N1573);
or OR2 (N7330, N7315, N6636);
nand NAND3 (N7331, N7328, N4607, N6940);
not NOT1 (N7332, N7325);
nand NAND3 (N7333, N7318, N1317, N1298);
and AND3 (N7334, N7319, N925, N773);
buf BUF1 (N7335, N7332);
and AND4 (N7336, N7304, N2341, N3944, N6084);
buf BUF1 (N7337, N7329);
and AND3 (N7338, N7333, N5866, N2244);
or OR4 (N7339, N7326, N1638, N141, N6769);
nor NOR3 (N7340, N7323, N4556, N4612);
nor NOR4 (N7341, N7338, N508, N5301, N6490);
and AND4 (N7342, N7337, N695, N6353, N2819);
and AND4 (N7343, N7341, N6419, N4282, N2991);
buf BUF1 (N7344, N7339);
and AND4 (N7345, N7331, N2955, N7110, N6364);
xor XOR2 (N7346, N7345, N5875);
buf BUF1 (N7347, N7342);
buf BUF1 (N7348, N7336);
buf BUF1 (N7349, N7348);
nand NAND3 (N7350, N7343, N4336, N3482);
or OR2 (N7351, N7344, N5971);
buf BUF1 (N7352, N7349);
buf BUF1 (N7353, N7346);
and AND2 (N7354, N7351, N7257);
not NOT1 (N7355, N7334);
nor NOR4 (N7356, N7350, N2356, N6944, N1530);
not NOT1 (N7357, N7354);
buf BUF1 (N7358, N7356);
nand NAND3 (N7359, N7335, N6154, N5830);
nand NAND2 (N7360, N7359, N3306);
not NOT1 (N7361, N7340);
or OR4 (N7362, N7324, N1916, N4540, N6854);
nor NOR3 (N7363, N7330, N3966, N2994);
or OR2 (N7364, N7355, N1622);
nor NOR4 (N7365, N7358, N6341, N1404, N7042);
and AND3 (N7366, N7357, N995, N5973);
nor NOR2 (N7367, N7347, N3858);
buf BUF1 (N7368, N7366);
nand NAND3 (N7369, N7362, N4142, N5682);
nand NAND2 (N7370, N7368, N2933);
not NOT1 (N7371, N7364);
nor NOR4 (N7372, N7353, N5398, N5803, N6091);
nand NAND3 (N7373, N7367, N3767, N7129);
xor XOR2 (N7374, N7370, N2746);
not NOT1 (N7375, N7365);
not NOT1 (N7376, N7369);
nand NAND4 (N7377, N7375, N2527, N2225, N3621);
xor XOR2 (N7378, N7360, N1894);
nand NAND3 (N7379, N7371, N6299, N5984);
not NOT1 (N7380, N7376);
nor NOR4 (N7381, N7380, N4300, N1757, N1073);
not NOT1 (N7382, N7363);
nand NAND2 (N7383, N7377, N4292);
xor XOR2 (N7384, N7374, N1640);
nand NAND3 (N7385, N7361, N3581, N4271);
xor XOR2 (N7386, N7382, N3867);
nor NOR4 (N7387, N7383, N832, N2205, N6032);
nand NAND2 (N7388, N7373, N3897);
not NOT1 (N7389, N7381);
nand NAND3 (N7390, N7352, N681, N264);
or OR2 (N7391, N7379, N1195);
xor XOR2 (N7392, N7384, N1670);
not NOT1 (N7393, N7372);
xor XOR2 (N7394, N7392, N4732);
nand NAND3 (N7395, N7385, N392, N569);
nand NAND3 (N7396, N7393, N1013, N7189);
xor XOR2 (N7397, N7378, N1249);
or OR4 (N7398, N7391, N1184, N4629, N6796);
xor XOR2 (N7399, N7386, N6721);
not NOT1 (N7400, N7397);
not NOT1 (N7401, N7394);
nand NAND3 (N7402, N7396, N2811, N3678);
buf BUF1 (N7403, N7387);
or OR4 (N7404, N7403, N7062, N1162, N2085);
nand NAND4 (N7405, N7401, N6265, N6743, N698);
buf BUF1 (N7406, N7389);
nand NAND4 (N7407, N7405, N5340, N4229, N2311);
not NOT1 (N7408, N7402);
buf BUF1 (N7409, N7407);
not NOT1 (N7410, N7395);
xor XOR2 (N7411, N7404, N5443);
xor XOR2 (N7412, N7409, N6993);
and AND3 (N7413, N7400, N6922, N3072);
nand NAND4 (N7414, N7406, N6795, N15, N2071);
xor XOR2 (N7415, N7388, N1317);
or OR3 (N7416, N7410, N931, N5003);
not NOT1 (N7417, N7398);
nand NAND3 (N7418, N7415, N6487, N489);
or OR3 (N7419, N7408, N1339, N4423);
nand NAND2 (N7420, N7419, N1650);
nand NAND4 (N7421, N7411, N468, N3226, N4183);
and AND2 (N7422, N7414, N5609);
nor NOR4 (N7423, N7418, N2663, N6528, N6454);
not NOT1 (N7424, N7413);
nand NAND3 (N7425, N7420, N1972, N3170);
or OR2 (N7426, N7425, N6161);
nand NAND4 (N7427, N7423, N5545, N4748, N5779);
not NOT1 (N7428, N7416);
and AND3 (N7429, N7399, N949, N3825);
buf BUF1 (N7430, N7421);
not NOT1 (N7431, N7390);
xor XOR2 (N7432, N7417, N1716);
buf BUF1 (N7433, N7422);
and AND2 (N7434, N7412, N6412);
not NOT1 (N7435, N7424);
xor XOR2 (N7436, N7429, N7184);
or OR4 (N7437, N7436, N3021, N38, N2969);
nand NAND2 (N7438, N7428, N3731);
xor XOR2 (N7439, N7435, N2580);
and AND3 (N7440, N7426, N4271, N7226);
and AND3 (N7441, N7433, N235, N2514);
buf BUF1 (N7442, N7430);
or OR4 (N7443, N7439, N5928, N3103, N974);
not NOT1 (N7444, N7431);
nand NAND3 (N7445, N7427, N6915, N1801);
or OR3 (N7446, N7441, N4260, N906);
buf BUF1 (N7447, N7443);
xor XOR2 (N7448, N7437, N4398);
and AND4 (N7449, N7444, N854, N3697, N1414);
xor XOR2 (N7450, N7432, N5491);
or OR2 (N7451, N7448, N4110);
buf BUF1 (N7452, N7445);
buf BUF1 (N7453, N7438);
or OR3 (N7454, N7440, N4418, N4316);
and AND4 (N7455, N7454, N3279, N1172, N2889);
and AND2 (N7456, N7442, N887);
and AND3 (N7457, N7453, N4190, N1842);
nand NAND4 (N7458, N7456, N2402, N3116, N393);
nand NAND3 (N7459, N7446, N2665, N1697);
nor NOR3 (N7460, N7447, N4004, N2676);
not NOT1 (N7461, N7449);
buf BUF1 (N7462, N7459);
xor XOR2 (N7463, N7450, N7366);
buf BUF1 (N7464, N7457);
not NOT1 (N7465, N7460);
nor NOR2 (N7466, N7434, N3009);
and AND2 (N7467, N7455, N4503);
nor NOR2 (N7468, N7466, N2686);
nand NAND4 (N7469, N7465, N2060, N1313, N1605);
nor NOR3 (N7470, N7462, N3327, N4895);
nand NAND2 (N7471, N7452, N4284);
nor NOR4 (N7472, N7461, N240, N1083, N2564);
and AND4 (N7473, N7469, N6247, N7412, N5322);
nand NAND3 (N7474, N7451, N5367, N2438);
nor NOR4 (N7475, N7473, N3142, N1220, N6251);
and AND3 (N7476, N7472, N6456, N5863);
or OR4 (N7477, N7475, N2543, N2368, N3539);
xor XOR2 (N7478, N7458, N2669);
buf BUF1 (N7479, N7478);
and AND2 (N7480, N7476, N659);
nand NAND3 (N7481, N7474, N1415, N6073);
and AND4 (N7482, N7471, N1099, N1450, N2605);
nand NAND3 (N7483, N7482, N6624, N2);
not NOT1 (N7484, N7481);
buf BUF1 (N7485, N7480);
xor XOR2 (N7486, N7477, N5088);
and AND3 (N7487, N7486, N1100, N6470);
buf BUF1 (N7488, N7468);
nor NOR4 (N7489, N7464, N827, N2052, N1323);
nand NAND4 (N7490, N7467, N3454, N1796, N5082);
nor NOR2 (N7491, N7484, N2376);
or OR2 (N7492, N7485, N1154);
or OR2 (N7493, N7490, N4190);
nand NAND2 (N7494, N7470, N33);
xor XOR2 (N7495, N7491, N5741);
xor XOR2 (N7496, N7488, N7023);
nand NAND2 (N7497, N7495, N1630);
nand NAND2 (N7498, N7494, N2463);
nand NAND4 (N7499, N7479, N7393, N1927, N570);
nor NOR2 (N7500, N7493, N2515);
and AND4 (N7501, N7498, N417, N5145, N5797);
nand NAND4 (N7502, N7492, N5161, N1948, N4836);
not NOT1 (N7503, N7501);
nand NAND4 (N7504, N7483, N3155, N3971, N7363);
not NOT1 (N7505, N7504);
not NOT1 (N7506, N7487);
or OR3 (N7507, N7496, N5885, N2835);
buf BUF1 (N7508, N7489);
not NOT1 (N7509, N7506);
not NOT1 (N7510, N7499);
nand NAND3 (N7511, N7502, N1687, N5453);
and AND3 (N7512, N7509, N6663, N4458);
or OR3 (N7513, N7497, N4333, N5018);
not NOT1 (N7514, N7513);
xor XOR2 (N7515, N7505, N1519);
and AND3 (N7516, N7500, N2148, N5582);
nor NOR2 (N7517, N7516, N3280);
xor XOR2 (N7518, N7511, N7257);
or OR4 (N7519, N7463, N5929, N1727, N5174);
nor NOR2 (N7520, N7510, N1484);
xor XOR2 (N7521, N7515, N6535);
nand NAND3 (N7522, N7512, N2341, N1518);
xor XOR2 (N7523, N7521, N7320);
nor NOR2 (N7524, N7508, N7195);
or OR2 (N7525, N7519, N1760);
xor XOR2 (N7526, N7523, N2826);
xor XOR2 (N7527, N7522, N6027);
xor XOR2 (N7528, N7503, N1502);
nor NOR4 (N7529, N7517, N3485, N4926, N629);
nand NAND4 (N7530, N7518, N6544, N7511, N3335);
and AND4 (N7531, N7529, N4857, N4738, N4203);
buf BUF1 (N7532, N7531);
and AND4 (N7533, N7527, N5269, N7063, N2440);
nand NAND2 (N7534, N7533, N991);
xor XOR2 (N7535, N7525, N5152);
or OR3 (N7536, N7530, N2991, N5642);
buf BUF1 (N7537, N7535);
and AND2 (N7538, N7514, N1668);
xor XOR2 (N7539, N7537, N7126);
xor XOR2 (N7540, N7526, N7464);
nand NAND2 (N7541, N7534, N703);
not NOT1 (N7542, N7520);
not NOT1 (N7543, N7539);
or OR3 (N7544, N7542, N6713, N254);
and AND2 (N7545, N7536, N4951);
xor XOR2 (N7546, N7524, N2120);
and AND3 (N7547, N7541, N3025, N2570);
or OR3 (N7548, N7538, N4145, N1552);
or OR4 (N7549, N7507, N4432, N5159, N2348);
not NOT1 (N7550, N7540);
not NOT1 (N7551, N7544);
and AND4 (N7552, N7546, N4757, N3243, N1933);
and AND3 (N7553, N7528, N5441, N5344);
nor NOR4 (N7554, N7551, N7487, N2755, N5943);
nor NOR4 (N7555, N7543, N1200, N5048, N938);
nand NAND3 (N7556, N7549, N5403, N116);
nand NAND3 (N7557, N7553, N6472, N6802);
xor XOR2 (N7558, N7547, N7530);
not NOT1 (N7559, N7554);
and AND4 (N7560, N7555, N5204, N4319, N3515);
nand NAND4 (N7561, N7532, N3786, N4102, N634);
or OR2 (N7562, N7557, N337);
and AND2 (N7563, N7548, N1532);
not NOT1 (N7564, N7563);
and AND3 (N7565, N7561, N7229, N5537);
nand NAND4 (N7566, N7564, N1583, N5673, N6572);
not NOT1 (N7567, N7566);
and AND4 (N7568, N7562, N3496, N4685, N6180);
buf BUF1 (N7569, N7560);
nor NOR2 (N7570, N7558, N749);
and AND2 (N7571, N7550, N6376);
and AND3 (N7572, N7570, N2010, N6254);
or OR3 (N7573, N7571, N4901, N6218);
xor XOR2 (N7574, N7552, N5518);
and AND3 (N7575, N7569, N13, N4763);
and AND3 (N7576, N7574, N2621, N2886);
or OR4 (N7577, N7567, N4654, N153, N222);
not NOT1 (N7578, N7559);
xor XOR2 (N7579, N7578, N400);
not NOT1 (N7580, N7577);
xor XOR2 (N7581, N7580, N2054);
not NOT1 (N7582, N7581);
or OR4 (N7583, N7579, N6373, N1760, N120);
nor NOR4 (N7584, N7573, N2618, N2674, N5564);
and AND3 (N7585, N7575, N6110, N4763);
and AND2 (N7586, N7584, N3565);
and AND3 (N7587, N7585, N5942, N2521);
and AND2 (N7588, N7545, N5296);
xor XOR2 (N7589, N7576, N978);
nor NOR4 (N7590, N7583, N1901, N5465, N6733);
nand NAND3 (N7591, N7589, N5382, N2110);
or OR3 (N7592, N7586, N3017, N668);
not NOT1 (N7593, N7592);
or OR4 (N7594, N7591, N3165, N2426, N3850);
nor NOR3 (N7595, N7593, N2525, N5360);
buf BUF1 (N7596, N7590);
not NOT1 (N7597, N7596);
nand NAND2 (N7598, N7572, N2762);
and AND2 (N7599, N7582, N3347);
xor XOR2 (N7600, N7594, N4109);
nand NAND4 (N7601, N7598, N670, N3976, N250);
not NOT1 (N7602, N7601);
buf BUF1 (N7603, N7599);
nor NOR4 (N7604, N7565, N7296, N2054, N5586);
buf BUF1 (N7605, N7588);
nor NOR3 (N7606, N7595, N5904, N5463);
nand NAND2 (N7607, N7587, N7330);
or OR2 (N7608, N7604, N2247);
xor XOR2 (N7609, N7600, N2550);
nand NAND2 (N7610, N7605, N6885);
or OR2 (N7611, N7609, N3315);
or OR3 (N7612, N7606, N4320, N5669);
not NOT1 (N7613, N7603);
and AND2 (N7614, N7613, N3123);
and AND4 (N7615, N7607, N6003, N7361, N1934);
or OR3 (N7616, N7611, N3740, N1819);
xor XOR2 (N7617, N7616, N710);
not NOT1 (N7618, N7597);
not NOT1 (N7619, N7618);
and AND3 (N7620, N7619, N670, N2712);
buf BUF1 (N7621, N7617);
or OR4 (N7622, N7621, N2567, N4295, N3486);
and AND3 (N7623, N7615, N5084, N2937);
nor NOR2 (N7624, N7622, N3103);
not NOT1 (N7625, N7624);
nor NOR2 (N7626, N7614, N6783);
or OR3 (N7627, N7625, N933, N3000);
xor XOR2 (N7628, N7626, N4460);
nand NAND3 (N7629, N7610, N2188, N7371);
xor XOR2 (N7630, N7629, N2449);
xor XOR2 (N7631, N7630, N3829);
or OR2 (N7632, N7631, N7558);
or OR4 (N7633, N7620, N4571, N622, N7555);
or OR2 (N7634, N7568, N2415);
and AND2 (N7635, N7633, N4071);
buf BUF1 (N7636, N7608);
and AND4 (N7637, N7635, N5170, N2050, N4551);
buf BUF1 (N7638, N7623);
or OR3 (N7639, N7627, N2116, N3512);
nor NOR3 (N7640, N7602, N677, N5988);
not NOT1 (N7641, N7612);
xor XOR2 (N7642, N7632, N1790);
and AND4 (N7643, N7639, N3449, N1939, N6063);
or OR3 (N7644, N7643, N5204, N3612);
nand NAND3 (N7645, N7644, N1814, N3503);
nor NOR2 (N7646, N7628, N5728);
xor XOR2 (N7647, N7556, N6095);
nor NOR2 (N7648, N7646, N6739);
nor NOR2 (N7649, N7648, N5208);
nand NAND4 (N7650, N7638, N4227, N5098, N4030);
not NOT1 (N7651, N7642);
buf BUF1 (N7652, N7637);
or OR2 (N7653, N7645, N34);
not NOT1 (N7654, N7653);
xor XOR2 (N7655, N7649, N1924);
nand NAND4 (N7656, N7655, N4854, N1086, N3738);
or OR3 (N7657, N7656, N782, N3458);
or OR3 (N7658, N7634, N2537, N2340);
not NOT1 (N7659, N7636);
nand NAND3 (N7660, N7647, N11, N4086);
buf BUF1 (N7661, N7654);
xor XOR2 (N7662, N7658, N5508);
nor NOR2 (N7663, N7651, N1075);
not NOT1 (N7664, N7640);
not NOT1 (N7665, N7661);
or OR4 (N7666, N7650, N1780, N595, N2900);
buf BUF1 (N7667, N7663);
xor XOR2 (N7668, N7666, N3851);
and AND3 (N7669, N7657, N3003, N267);
xor XOR2 (N7670, N7669, N3153);
buf BUF1 (N7671, N7652);
and AND3 (N7672, N7641, N2031, N667);
nand NAND4 (N7673, N7670, N6101, N7459, N6404);
nor NOR4 (N7674, N7662, N7356, N1344, N676);
xor XOR2 (N7675, N7674, N1016);
xor XOR2 (N7676, N7660, N2013);
buf BUF1 (N7677, N7675);
not NOT1 (N7678, N7672);
buf BUF1 (N7679, N7665);
nand NAND2 (N7680, N7668, N4998);
nand NAND4 (N7681, N7680, N1930, N3246, N2850);
or OR2 (N7682, N7664, N3296);
nor NOR2 (N7683, N7677, N2647);
nor NOR4 (N7684, N7676, N1395, N533, N5332);
not NOT1 (N7685, N7678);
not NOT1 (N7686, N7673);
not NOT1 (N7687, N7684);
not NOT1 (N7688, N7679);
xor XOR2 (N7689, N7687, N6962);
xor XOR2 (N7690, N7659, N2085);
or OR3 (N7691, N7671, N3074, N5074);
not NOT1 (N7692, N7685);
buf BUF1 (N7693, N7686);
nand NAND4 (N7694, N7688, N2675, N7222, N51);
nand NAND3 (N7695, N7689, N7005, N6571);
not NOT1 (N7696, N7692);
nand NAND4 (N7697, N7691, N5599, N3000, N1606);
not NOT1 (N7698, N7667);
and AND4 (N7699, N7695, N2405, N885, N7520);
buf BUF1 (N7700, N7696);
buf BUF1 (N7701, N7681);
nand NAND4 (N7702, N7699, N7092, N2889, N5787);
buf BUF1 (N7703, N7682);
xor XOR2 (N7704, N7694, N5001);
and AND3 (N7705, N7690, N207, N6011);
or OR2 (N7706, N7697, N2122);
nor NOR4 (N7707, N7700, N5864, N451, N519);
buf BUF1 (N7708, N7698);
or OR2 (N7709, N7705, N99);
buf BUF1 (N7710, N7709);
buf BUF1 (N7711, N7701);
xor XOR2 (N7712, N7706, N6264);
buf BUF1 (N7713, N7683);
and AND2 (N7714, N7713, N2640);
nand NAND4 (N7715, N7714, N2604, N4481, N6441);
buf BUF1 (N7716, N7711);
xor XOR2 (N7717, N7716, N7570);
nor NOR3 (N7718, N7715, N6383, N482);
nor NOR4 (N7719, N7710, N618, N810, N1911);
xor XOR2 (N7720, N7712, N6792);
buf BUF1 (N7721, N7707);
buf BUF1 (N7722, N7720);
buf BUF1 (N7723, N7718);
nor NOR2 (N7724, N7703, N6101);
not NOT1 (N7725, N7702);
and AND2 (N7726, N7704, N1699);
nor NOR4 (N7727, N7693, N515, N1859, N2166);
buf BUF1 (N7728, N7717);
and AND4 (N7729, N7726, N3171, N6128, N6381);
not NOT1 (N7730, N7727);
nand NAND4 (N7731, N7724, N5925, N3006, N2732);
not NOT1 (N7732, N7721);
xor XOR2 (N7733, N7728, N4733);
nand NAND2 (N7734, N7733, N7122);
xor XOR2 (N7735, N7722, N2553);
xor XOR2 (N7736, N7719, N797);
xor XOR2 (N7737, N7708, N6541);
not NOT1 (N7738, N7729);
nand NAND2 (N7739, N7738, N5500);
nor NOR2 (N7740, N7725, N802);
nor NOR4 (N7741, N7739, N3368, N2309, N4727);
nand NAND4 (N7742, N7736, N3768, N7090, N7011);
and AND2 (N7743, N7732, N5304);
and AND2 (N7744, N7730, N4965);
not NOT1 (N7745, N7731);
or OR2 (N7746, N7743, N5725);
and AND2 (N7747, N7742, N649);
and AND3 (N7748, N7737, N3370, N697);
nand NAND3 (N7749, N7745, N4294, N5442);
nor NOR4 (N7750, N7723, N39, N643, N2206);
nand NAND2 (N7751, N7747, N2331);
and AND2 (N7752, N7746, N2265);
or OR4 (N7753, N7752, N2367, N4935, N1309);
xor XOR2 (N7754, N7753, N1324);
xor XOR2 (N7755, N7744, N3752);
and AND2 (N7756, N7755, N2150);
xor XOR2 (N7757, N7756, N2432);
nor NOR3 (N7758, N7741, N5412, N4958);
or OR4 (N7759, N7750, N1591, N2033, N1230);
nor NOR4 (N7760, N7751, N4185, N2530, N2181);
buf BUF1 (N7761, N7748);
or OR2 (N7762, N7734, N333);
nor NOR3 (N7763, N7759, N993, N980);
not NOT1 (N7764, N7762);
nand NAND3 (N7765, N7764, N5741, N6977);
nor NOR2 (N7766, N7758, N2736);
xor XOR2 (N7767, N7763, N1581);
nor NOR4 (N7768, N7749, N5016, N4819, N3157);
nor NOR2 (N7769, N7754, N440);
buf BUF1 (N7770, N7735);
xor XOR2 (N7771, N7740, N5514);
or OR3 (N7772, N7766, N700, N3187);
or OR3 (N7773, N7767, N6094, N6411);
and AND3 (N7774, N7761, N3014, N5791);
and AND4 (N7775, N7771, N400, N1080, N7729);
not NOT1 (N7776, N7757);
or OR4 (N7777, N7769, N3187, N2712, N1101);
buf BUF1 (N7778, N7774);
buf BUF1 (N7779, N7765);
and AND4 (N7780, N7778, N4197, N4238, N277);
nand NAND4 (N7781, N7780, N2284, N4943, N3729);
xor XOR2 (N7782, N7775, N1246);
xor XOR2 (N7783, N7772, N4451);
nor NOR2 (N7784, N7781, N3995);
and AND2 (N7785, N7773, N2518);
and AND4 (N7786, N7760, N2343, N1591, N5622);
nand NAND3 (N7787, N7785, N6733, N806);
buf BUF1 (N7788, N7784);
nor NOR2 (N7789, N7788, N7335);
not NOT1 (N7790, N7777);
nor NOR3 (N7791, N7789, N566, N1536);
and AND2 (N7792, N7786, N3395);
and AND3 (N7793, N7779, N5881, N4071);
or OR4 (N7794, N7782, N6387, N3503, N3601);
and AND2 (N7795, N7794, N2457);
nor NOR4 (N7796, N7790, N531, N2597, N5858);
and AND4 (N7797, N7795, N5461, N2675, N6365);
or OR4 (N7798, N7768, N1362, N2690, N4951);
buf BUF1 (N7799, N7791);
nor NOR4 (N7800, N7796, N3571, N2563, N5118);
or OR2 (N7801, N7797, N5272);
or OR2 (N7802, N7770, N6028);
or OR3 (N7803, N7800, N7766, N579);
buf BUF1 (N7804, N7783);
buf BUF1 (N7805, N7792);
xor XOR2 (N7806, N7804, N1016);
or OR2 (N7807, N7806, N7266);
and AND4 (N7808, N7798, N946, N4051, N2170);
xor XOR2 (N7809, N7787, N4082);
nor NOR3 (N7810, N7808, N3064, N5829);
and AND4 (N7811, N7801, N4002, N7172, N2048);
nand NAND3 (N7812, N7802, N6911, N6081);
buf BUF1 (N7813, N7807);
nand NAND3 (N7814, N7811, N163, N5065);
nor NOR4 (N7815, N7793, N5710, N3625, N6552);
not NOT1 (N7816, N7814);
not NOT1 (N7817, N7813);
and AND4 (N7818, N7803, N5071, N6830, N4901);
nand NAND4 (N7819, N7816, N2058, N2156, N1745);
not NOT1 (N7820, N7810);
not NOT1 (N7821, N7812);
nand NAND3 (N7822, N7799, N6659, N6203);
nor NOR4 (N7823, N7805, N1064, N4829, N5285);
nor NOR4 (N7824, N7822, N1077, N2291, N805);
or OR3 (N7825, N7824, N265, N5885);
xor XOR2 (N7826, N7819, N7412);
nor NOR2 (N7827, N7817, N797);
xor XOR2 (N7828, N7818, N3245);
xor XOR2 (N7829, N7821, N2231);
nor NOR4 (N7830, N7820, N7100, N4930, N2307);
nand NAND4 (N7831, N7776, N1673, N5651, N6955);
and AND2 (N7832, N7809, N3456);
xor XOR2 (N7833, N7831, N896);
nor NOR3 (N7834, N7828, N2006, N6033);
xor XOR2 (N7835, N7826, N309);
not NOT1 (N7836, N7829);
not NOT1 (N7837, N7815);
xor XOR2 (N7838, N7837, N7243);
and AND4 (N7839, N7823, N2181, N4639, N2250);
nand NAND4 (N7840, N7833, N6649, N4304, N1061);
or OR2 (N7841, N7825, N1041);
not NOT1 (N7842, N7838);
or OR2 (N7843, N7835, N7525);
xor XOR2 (N7844, N7843, N1997);
xor XOR2 (N7845, N7844, N4456);
and AND4 (N7846, N7836, N3622, N6127, N6570);
nand NAND3 (N7847, N7830, N3715, N7400);
not NOT1 (N7848, N7839);
buf BUF1 (N7849, N7832);
and AND3 (N7850, N7840, N5257, N3178);
and AND2 (N7851, N7842, N1753);
not NOT1 (N7852, N7846);
nor NOR2 (N7853, N7845, N86);
not NOT1 (N7854, N7848);
xor XOR2 (N7855, N7851, N3085);
or OR2 (N7856, N7853, N1036);
xor XOR2 (N7857, N7841, N1570);
buf BUF1 (N7858, N7850);
not NOT1 (N7859, N7855);
nor NOR2 (N7860, N7859, N2653);
nand NAND3 (N7861, N7849, N7199, N5851);
buf BUF1 (N7862, N7857);
nand NAND3 (N7863, N7827, N2611, N3328);
buf BUF1 (N7864, N7863);
or OR4 (N7865, N7847, N330, N5385, N7816);
or OR4 (N7866, N7865, N1098, N3601, N6930);
nor NOR2 (N7867, N7856, N6077);
nand NAND4 (N7868, N7834, N6108, N6563, N5403);
nand NAND2 (N7869, N7866, N1043);
buf BUF1 (N7870, N7868);
or OR2 (N7871, N7858, N6380);
nor NOR3 (N7872, N7852, N6822, N3665);
not NOT1 (N7873, N7860);
xor XOR2 (N7874, N7861, N5812);
and AND2 (N7875, N7854, N1310);
xor XOR2 (N7876, N7869, N758);
xor XOR2 (N7877, N7867, N7629);
nor NOR4 (N7878, N7872, N3537, N3199, N7641);
nand NAND3 (N7879, N7874, N5351, N4762);
xor XOR2 (N7880, N7873, N7458);
nand NAND2 (N7881, N7864, N3306);
not NOT1 (N7882, N7862);
nor NOR3 (N7883, N7871, N3320, N6957);
xor XOR2 (N7884, N7875, N1870);
xor XOR2 (N7885, N7880, N1818);
nand NAND3 (N7886, N7877, N2226, N3443);
and AND4 (N7887, N7876, N1676, N1948, N7599);
buf BUF1 (N7888, N7887);
or OR4 (N7889, N7882, N4656, N4493, N1113);
nor NOR2 (N7890, N7885, N3483);
not NOT1 (N7891, N7884);
and AND4 (N7892, N7891, N2436, N7473, N7143);
buf BUF1 (N7893, N7892);
or OR4 (N7894, N7879, N1228, N4623, N6535);
and AND2 (N7895, N7878, N1258);
xor XOR2 (N7896, N7893, N3622);
and AND4 (N7897, N7886, N4010, N307, N1771);
and AND3 (N7898, N7888, N6507, N5289);
or OR3 (N7899, N7897, N4399, N658);
buf BUF1 (N7900, N7898);
xor XOR2 (N7901, N7870, N6912);
nand NAND2 (N7902, N7881, N1825);
xor XOR2 (N7903, N7900, N650);
and AND4 (N7904, N7899, N7858, N7249, N6662);
buf BUF1 (N7905, N7895);
nand NAND4 (N7906, N7902, N1420, N2854, N1208);
and AND4 (N7907, N7901, N852, N7189, N2211);
and AND2 (N7908, N7889, N2385);
xor XOR2 (N7909, N7904, N6736);
nand NAND3 (N7910, N7909, N5546, N4531);
buf BUF1 (N7911, N7910);
or OR2 (N7912, N7905, N1329);
nand NAND3 (N7913, N7896, N3087, N6348);
nand NAND2 (N7914, N7912, N5322);
or OR2 (N7915, N7908, N7111);
not NOT1 (N7916, N7915);
or OR3 (N7917, N7907, N3850, N1819);
not NOT1 (N7918, N7917);
buf BUF1 (N7919, N7913);
not NOT1 (N7920, N7911);
nor NOR3 (N7921, N7903, N3057, N3973);
not NOT1 (N7922, N7918);
and AND4 (N7923, N7920, N4698, N4600, N1636);
buf BUF1 (N7924, N7921);
nor NOR2 (N7925, N7914, N3664);
nand NAND3 (N7926, N7894, N1853, N5415);
nand NAND2 (N7927, N7906, N3275);
not NOT1 (N7928, N7926);
buf BUF1 (N7929, N7927);
nand NAND4 (N7930, N7923, N1879, N7348, N3134);
xor XOR2 (N7931, N7925, N1249);
nand NAND4 (N7932, N7924, N2297, N1565, N1677);
and AND2 (N7933, N7922, N5152);
buf BUF1 (N7934, N7919);
nor NOR4 (N7935, N7931, N3847, N4337, N2582);
buf BUF1 (N7936, N7929);
not NOT1 (N7937, N7928);
and AND2 (N7938, N7934, N7359);
and AND4 (N7939, N7932, N7212, N4354, N5642);
nor NOR3 (N7940, N7936, N3871, N6837);
nor NOR3 (N7941, N7916, N6761, N2383);
nor NOR4 (N7942, N7940, N3591, N2451, N7932);
nand NAND4 (N7943, N7937, N889, N7585, N329);
buf BUF1 (N7944, N7943);
not NOT1 (N7945, N7942);
or OR3 (N7946, N7939, N5964, N3833);
or OR3 (N7947, N7935, N4696, N6945);
not NOT1 (N7948, N7883);
not NOT1 (N7949, N7947);
xor XOR2 (N7950, N7941, N6788);
xor XOR2 (N7951, N7948, N356);
and AND3 (N7952, N7890, N7710, N3346);
nand NAND2 (N7953, N7951, N4159);
and AND2 (N7954, N7949, N6386);
buf BUF1 (N7955, N7930);
not NOT1 (N7956, N7944);
and AND2 (N7957, N7954, N5516);
xor XOR2 (N7958, N7952, N2232);
and AND4 (N7959, N7933, N599, N5778, N441);
buf BUF1 (N7960, N7953);
nor NOR3 (N7961, N7950, N2378, N727);
xor XOR2 (N7962, N7955, N3870);
and AND2 (N7963, N7945, N7146);
not NOT1 (N7964, N7956);
and AND2 (N7965, N7946, N4753);
and AND4 (N7966, N7960, N2666, N4100, N5501);
xor XOR2 (N7967, N7963, N3406);
nand NAND2 (N7968, N7959, N3110);
xor XOR2 (N7969, N7958, N2651);
nand NAND2 (N7970, N7969, N2921);
nor NOR4 (N7971, N7962, N6102, N134, N5288);
buf BUF1 (N7972, N7968);
or OR2 (N7973, N7972, N6088);
not NOT1 (N7974, N7961);
xor XOR2 (N7975, N7971, N7509);
nor NOR3 (N7976, N7957, N576, N6919);
not NOT1 (N7977, N7970);
buf BUF1 (N7978, N7967);
xor XOR2 (N7979, N7965, N7763);
and AND2 (N7980, N7974, N3415);
not NOT1 (N7981, N7978);
xor XOR2 (N7982, N7976, N547);
and AND2 (N7983, N7973, N6926);
not NOT1 (N7984, N7982);
buf BUF1 (N7985, N7980);
not NOT1 (N7986, N7979);
buf BUF1 (N7987, N7975);
xor XOR2 (N7988, N7983, N6632);
nor NOR2 (N7989, N7981, N3078);
nand NAND3 (N7990, N7985, N1948, N7655);
nand NAND3 (N7991, N7986, N490, N4501);
xor XOR2 (N7992, N7977, N1632);
not NOT1 (N7993, N7984);
nand NAND2 (N7994, N7987, N6276);
nand NAND4 (N7995, N7994, N3483, N4800, N759);
xor XOR2 (N7996, N7990, N1024);
and AND2 (N7997, N7988, N7377);
or OR2 (N7998, N7992, N5766);
nor NOR3 (N7999, N7998, N3731, N1992);
nor NOR2 (N8000, N7991, N4635);
or OR2 (N8001, N7993, N5027);
xor XOR2 (N8002, N8001, N26);
not NOT1 (N8003, N7997);
or OR2 (N8004, N7999, N893);
nand NAND4 (N8005, N8004, N1760, N956, N6601);
not NOT1 (N8006, N7966);
and AND4 (N8007, N7995, N1029, N6911, N4389);
buf BUF1 (N8008, N7964);
or OR3 (N8009, N7996, N6493, N3774);
xor XOR2 (N8010, N8000, N2177);
nor NOR4 (N8011, N7989, N6862, N75, N4132);
or OR3 (N8012, N8008, N2743, N2312);
not NOT1 (N8013, N8011);
and AND3 (N8014, N8002, N1753, N3841);
nor NOR3 (N8015, N8007, N3303, N3149);
buf BUF1 (N8016, N7938);
and AND3 (N8017, N8006, N5056, N5049);
nand NAND3 (N8018, N8009, N3753, N3287);
nor NOR4 (N8019, N8016, N418, N1440, N429);
nand NAND3 (N8020, N8015, N189, N7389);
nor NOR2 (N8021, N8003, N2409);
xor XOR2 (N8022, N8021, N5979);
xor XOR2 (N8023, N8020, N5711);
nand NAND3 (N8024, N8019, N704, N3012);
and AND4 (N8025, N8023, N3731, N6067, N6488);
and AND2 (N8026, N8022, N3525);
and AND3 (N8027, N8010, N2109, N1232);
nand NAND4 (N8028, N8025, N3706, N4506, N2239);
nor NOR3 (N8029, N8013, N5207, N4675);
not NOT1 (N8030, N8027);
xor XOR2 (N8031, N8005, N7017);
xor XOR2 (N8032, N8017, N5672);
nor NOR3 (N8033, N8028, N350, N4331);
buf BUF1 (N8034, N8018);
xor XOR2 (N8035, N8029, N5564);
xor XOR2 (N8036, N8034, N5370);
nand NAND4 (N8037, N8032, N745, N2535, N7821);
xor XOR2 (N8038, N8035, N7606);
or OR4 (N8039, N8036, N3962, N1664, N2492);
xor XOR2 (N8040, N8014, N3315);
or OR2 (N8041, N8038, N6307);
xor XOR2 (N8042, N8037, N652);
or OR4 (N8043, N8033, N679, N7005, N4371);
xor XOR2 (N8044, N8039, N4723);
nor NOR4 (N8045, N8041, N1052, N1563, N6383);
or OR2 (N8046, N8045, N291);
nor NOR4 (N8047, N8030, N3611, N4407, N3623);
nand NAND4 (N8048, N8012, N5460, N6476, N2890);
xor XOR2 (N8049, N8040, N3432);
or OR3 (N8050, N8026, N60, N7738);
nand NAND4 (N8051, N8042, N4167, N7957, N1015);
or OR3 (N8052, N8031, N4065, N4891);
nor NOR4 (N8053, N8044, N849, N6478, N1032);
and AND2 (N8054, N8046, N2318);
and AND4 (N8055, N8024, N5057, N2428, N760);
or OR4 (N8056, N8049, N3816, N7929, N330);
nand NAND2 (N8057, N8055, N1024);
not NOT1 (N8058, N8052);
or OR4 (N8059, N8048, N6775, N19, N3998);
and AND3 (N8060, N8059, N4547, N2027);
nand NAND3 (N8061, N8057, N2715, N5050);
xor XOR2 (N8062, N8058, N6321);
or OR2 (N8063, N8051, N2512);
buf BUF1 (N8064, N8047);
buf BUF1 (N8065, N8062);
nand NAND2 (N8066, N8056, N2931);
not NOT1 (N8067, N8060);
xor XOR2 (N8068, N8064, N3004);
xor XOR2 (N8069, N8050, N5065);
nand NAND4 (N8070, N8069, N4791, N278, N6215);
nand NAND3 (N8071, N8067, N3919, N2975);
or OR3 (N8072, N8068, N7935, N5147);
not NOT1 (N8073, N8061);
nor NOR4 (N8074, N8066, N4657, N1874, N1228);
not NOT1 (N8075, N8053);
xor XOR2 (N8076, N8072, N462);
xor XOR2 (N8077, N8075, N578);
nand NAND4 (N8078, N8077, N5311, N1493, N3590);
not NOT1 (N8079, N8071);
or OR4 (N8080, N8043, N6597, N6742, N6150);
xor XOR2 (N8081, N8063, N7069);
buf BUF1 (N8082, N8079);
or OR2 (N8083, N8073, N6655);
or OR4 (N8084, N8070, N553, N5841, N6431);
buf BUF1 (N8085, N8054);
xor XOR2 (N8086, N8076, N5276);
or OR2 (N8087, N8081, N7748);
xor XOR2 (N8088, N8074, N844);
and AND4 (N8089, N8088, N5234, N3852, N6522);
buf BUF1 (N8090, N8089);
nand NAND3 (N8091, N8086, N1813, N7133);
xor XOR2 (N8092, N8078, N177);
nand NAND2 (N8093, N8090, N4746);
and AND3 (N8094, N8091, N5334, N4182);
nand NAND4 (N8095, N8084, N225, N6807, N3504);
or OR2 (N8096, N8083, N6061);
or OR4 (N8097, N8065, N2015, N6760, N6437);
nor NOR4 (N8098, N8082, N5200, N3623, N1371);
not NOT1 (N8099, N8098);
xor XOR2 (N8100, N8096, N5661);
buf BUF1 (N8101, N8099);
nor NOR2 (N8102, N8097, N2867);
buf BUF1 (N8103, N8100);
nand NAND3 (N8104, N8103, N5542, N3109);
nand NAND2 (N8105, N8080, N4938);
nor NOR2 (N8106, N8104, N2194);
not NOT1 (N8107, N8085);
and AND2 (N8108, N8087, N7545);
nor NOR4 (N8109, N8092, N7333, N7277, N574);
and AND4 (N8110, N8094, N4902, N7685, N7784);
and AND4 (N8111, N8105, N5493, N7210, N5047);
xor XOR2 (N8112, N8109, N2479);
and AND3 (N8113, N8102, N529, N6935);
and AND4 (N8114, N8108, N5162, N7230, N998);
buf BUF1 (N8115, N8112);
buf BUF1 (N8116, N8115);
nand NAND2 (N8117, N8106, N5251);
not NOT1 (N8118, N8110);
buf BUF1 (N8119, N8114);
and AND3 (N8120, N8119, N5059, N1232);
nor NOR3 (N8121, N8111, N7891, N7444);
or OR4 (N8122, N8117, N2499, N1200, N1935);
not NOT1 (N8123, N8116);
and AND3 (N8124, N8113, N6928, N7898);
not NOT1 (N8125, N8118);
and AND3 (N8126, N8122, N4644, N7028);
xor XOR2 (N8127, N8093, N2398);
and AND2 (N8128, N8126, N2295);
xor XOR2 (N8129, N8128, N5184);
not NOT1 (N8130, N8095);
nand NAND3 (N8131, N8127, N5264, N2924);
and AND2 (N8132, N8124, N4167);
or OR2 (N8133, N8123, N521);
buf BUF1 (N8134, N8129);
nand NAND3 (N8135, N8101, N2666, N4808);
buf BUF1 (N8136, N8134);
xor XOR2 (N8137, N8125, N4550);
not NOT1 (N8138, N8132);
nor NOR2 (N8139, N8133, N1201);
nand NAND2 (N8140, N8137, N311);
nand NAND3 (N8141, N8107, N2239, N7597);
and AND4 (N8142, N8130, N2496, N3410, N4165);
nor NOR2 (N8143, N8120, N3829);
xor XOR2 (N8144, N8131, N1966);
or OR2 (N8145, N8136, N43);
buf BUF1 (N8146, N8139);
buf BUF1 (N8147, N8146);
nor NOR3 (N8148, N8135, N4766, N2644);
nand NAND2 (N8149, N8121, N7909);
xor XOR2 (N8150, N8148, N8075);
xor XOR2 (N8151, N8147, N4272);
nand NAND4 (N8152, N8144, N2049, N716, N2792);
nor NOR2 (N8153, N8142, N881);
or OR3 (N8154, N8152, N5447, N2789);
nand NAND3 (N8155, N8150, N6663, N5124);
xor XOR2 (N8156, N8153, N6827);
xor XOR2 (N8157, N8155, N1401);
or OR3 (N8158, N8143, N6463, N3994);
buf BUF1 (N8159, N8138);
nor NOR3 (N8160, N8140, N4267, N1678);
xor XOR2 (N8161, N8154, N6513);
buf BUF1 (N8162, N8141);
and AND4 (N8163, N8162, N6372, N6979, N1297);
nand NAND3 (N8164, N8151, N1726, N1747);
nand NAND3 (N8165, N8158, N4813, N7754);
and AND2 (N8166, N8149, N6057);
or OR2 (N8167, N8166, N1403);
and AND3 (N8168, N8159, N7221, N5716);
and AND2 (N8169, N8145, N2619);
not NOT1 (N8170, N8167);
not NOT1 (N8171, N8164);
or OR4 (N8172, N8165, N7009, N6259, N5097);
not NOT1 (N8173, N8163);
buf BUF1 (N8174, N8173);
xor XOR2 (N8175, N8172, N4927);
or OR3 (N8176, N8161, N7771, N4846);
xor XOR2 (N8177, N8168, N1895);
and AND4 (N8178, N8169, N6073, N1414, N1539);
nand NAND3 (N8179, N8157, N1888, N399);
nand NAND3 (N8180, N8175, N485, N1036);
not NOT1 (N8181, N8171);
xor XOR2 (N8182, N8179, N922);
nor NOR2 (N8183, N8156, N7548);
buf BUF1 (N8184, N8182);
nor NOR2 (N8185, N8184, N2014);
buf BUF1 (N8186, N8176);
and AND2 (N8187, N8180, N2287);
not NOT1 (N8188, N8174);
and AND3 (N8189, N8188, N1914, N2466);
and AND4 (N8190, N8186, N5458, N7739, N4165);
xor XOR2 (N8191, N8183, N5981);
nor NOR4 (N8192, N8170, N8071, N1295, N3879);
or OR4 (N8193, N8189, N6161, N125, N7073);
not NOT1 (N8194, N8187);
buf BUF1 (N8195, N8191);
and AND4 (N8196, N8178, N2295, N7058, N4567);
not NOT1 (N8197, N8195);
and AND3 (N8198, N8160, N86, N2770);
or OR3 (N8199, N8192, N1988, N4257);
nand NAND3 (N8200, N8198, N2387, N1257);
nor NOR2 (N8201, N8193, N112);
nor NOR4 (N8202, N8201, N5712, N931, N3127);
or OR2 (N8203, N8181, N1145);
nor NOR2 (N8204, N8194, N1961);
and AND4 (N8205, N8202, N2835, N2256, N4345);
buf BUF1 (N8206, N8199);
xor XOR2 (N8207, N8196, N3530);
or OR2 (N8208, N8206, N5454);
buf BUF1 (N8209, N8185);
buf BUF1 (N8210, N8207);
xor XOR2 (N8211, N8200, N1356);
not NOT1 (N8212, N8203);
buf BUF1 (N8213, N8205);
buf BUF1 (N8214, N8190);
or OR3 (N8215, N8211, N208, N3494);
nor NOR2 (N8216, N8215, N7895);
buf BUF1 (N8217, N8212);
and AND4 (N8218, N8216, N4011, N7196, N1460);
nor NOR4 (N8219, N8218, N1363, N7370, N4544);
or OR3 (N8220, N8208, N5733, N4462);
xor XOR2 (N8221, N8210, N2931);
and AND2 (N8222, N8220, N2737);
xor XOR2 (N8223, N8214, N1135);
and AND4 (N8224, N8219, N703, N1985, N2286);
nor NOR2 (N8225, N8224, N707);
nor NOR2 (N8226, N8197, N3567);
nand NAND4 (N8227, N8204, N2300, N6160, N19);
and AND4 (N8228, N8222, N2535, N5224, N7879);
nor NOR2 (N8229, N8226, N2717);
buf BUF1 (N8230, N8217);
nor NOR3 (N8231, N8177, N5100, N8097);
xor XOR2 (N8232, N8223, N5434);
not NOT1 (N8233, N8213);
nand NAND4 (N8234, N8228, N6810, N717, N3631);
and AND3 (N8235, N8231, N3394, N7107);
xor XOR2 (N8236, N8227, N2333);
or OR4 (N8237, N8229, N59, N7336, N2820);
nand NAND3 (N8238, N8237, N729, N6854);
and AND3 (N8239, N8221, N2317, N5360);
or OR4 (N8240, N8225, N1112, N3910, N6905);
or OR2 (N8241, N8230, N7131);
xor XOR2 (N8242, N8239, N5849);
xor XOR2 (N8243, N8209, N2181);
buf BUF1 (N8244, N8241);
xor XOR2 (N8245, N8243, N1364);
xor XOR2 (N8246, N8232, N8240);
or OR4 (N8247, N4287, N4897, N2345, N4638);
xor XOR2 (N8248, N8242, N3075);
nand NAND4 (N8249, N8235, N1260, N7168, N512);
nand NAND3 (N8250, N8246, N840, N358);
nand NAND4 (N8251, N8236, N6465, N5319, N3780);
xor XOR2 (N8252, N8238, N8237);
not NOT1 (N8253, N8233);
or OR3 (N8254, N8244, N3743, N6688);
or OR2 (N8255, N8248, N6914);
xor XOR2 (N8256, N8252, N5960);
nand NAND3 (N8257, N8247, N2639, N7904);
nand NAND2 (N8258, N8257, N2731);
nand NAND3 (N8259, N8250, N171, N4407);
not NOT1 (N8260, N8234);
xor XOR2 (N8261, N8253, N3702);
not NOT1 (N8262, N8251);
nand NAND2 (N8263, N8254, N7917);
and AND3 (N8264, N8258, N2142, N5562);
nand NAND3 (N8265, N8263, N4718, N3351);
nor NOR3 (N8266, N8255, N1053, N2133);
or OR4 (N8267, N8266, N7631, N1270, N4736);
xor XOR2 (N8268, N8256, N6316);
nor NOR2 (N8269, N8260, N412);
nand NAND4 (N8270, N8245, N4368, N1205, N3896);
buf BUF1 (N8271, N8270);
not NOT1 (N8272, N8249);
nor NOR3 (N8273, N8264, N6352, N6855);
nor NOR2 (N8274, N8273, N2615);
not NOT1 (N8275, N8267);
xor XOR2 (N8276, N8261, N3989);
buf BUF1 (N8277, N8262);
and AND4 (N8278, N8269, N8115, N1040, N413);
xor XOR2 (N8279, N8276, N6168);
and AND3 (N8280, N8277, N7212, N6840);
and AND4 (N8281, N8259, N7930, N7165, N7800);
or OR3 (N8282, N8278, N5916, N1276);
buf BUF1 (N8283, N8272);
and AND3 (N8284, N8281, N846, N1623);
xor XOR2 (N8285, N8282, N6303);
xor XOR2 (N8286, N8275, N883);
not NOT1 (N8287, N8268);
nor NOR2 (N8288, N8283, N2241);
not NOT1 (N8289, N8285);
xor XOR2 (N8290, N8280, N6773);
or OR3 (N8291, N8265, N191, N5961);
nand NAND4 (N8292, N8279, N1298, N8134, N1268);
xor XOR2 (N8293, N8274, N851);
buf BUF1 (N8294, N8289);
not NOT1 (N8295, N8291);
not NOT1 (N8296, N8292);
not NOT1 (N8297, N8296);
nor NOR2 (N8298, N8271, N7204);
not NOT1 (N8299, N8293);
nand NAND2 (N8300, N8284, N193);
and AND2 (N8301, N8287, N6847);
and AND2 (N8302, N8299, N3359);
nor NOR2 (N8303, N8300, N4397);
xor XOR2 (N8304, N8302, N5547);
not NOT1 (N8305, N8297);
xor XOR2 (N8306, N8295, N7840);
xor XOR2 (N8307, N8303, N4246);
xor XOR2 (N8308, N8298, N2497);
buf BUF1 (N8309, N8304);
not NOT1 (N8310, N8307);
buf BUF1 (N8311, N8310);
or OR2 (N8312, N8301, N7270);
not NOT1 (N8313, N8286);
nand NAND4 (N8314, N8305, N3464, N4069, N666);
nand NAND4 (N8315, N8290, N7144, N3304, N6784);
nor NOR2 (N8316, N8294, N7389);
or OR4 (N8317, N8315, N7206, N8229, N5806);
nand NAND3 (N8318, N8288, N5946, N4767);
or OR2 (N8319, N8311, N7149);
not NOT1 (N8320, N8314);
and AND4 (N8321, N8319, N1031, N5623, N835);
or OR4 (N8322, N8309, N6858, N692, N661);
xor XOR2 (N8323, N8322, N603);
nor NOR3 (N8324, N8306, N7783, N3408);
or OR4 (N8325, N8316, N2213, N5398, N8166);
xor XOR2 (N8326, N8308, N5233);
and AND2 (N8327, N8325, N2374);
or OR4 (N8328, N8317, N6527, N6904, N2139);
and AND3 (N8329, N8312, N6650, N4611);
nand NAND3 (N8330, N8313, N7834, N894);
xor XOR2 (N8331, N8320, N1466);
and AND2 (N8332, N8328, N159);
buf BUF1 (N8333, N8329);
not NOT1 (N8334, N8331);
buf BUF1 (N8335, N8334);
and AND2 (N8336, N8324, N1030);
nand NAND4 (N8337, N8330, N3642, N5045, N280);
buf BUF1 (N8338, N8337);
nor NOR3 (N8339, N8318, N6230, N6763);
and AND4 (N8340, N8326, N8242, N4273, N1702);
buf BUF1 (N8341, N8327);
nor NOR2 (N8342, N8338, N1587);
nand NAND4 (N8343, N8342, N2878, N737, N6093);
or OR2 (N8344, N8340, N7127);
xor XOR2 (N8345, N8339, N4171);
not NOT1 (N8346, N8343);
nand NAND3 (N8347, N8344, N4479, N7394);
not NOT1 (N8348, N8335);
buf BUF1 (N8349, N8341);
nand NAND2 (N8350, N8333, N8031);
or OR2 (N8351, N8347, N3619);
buf BUF1 (N8352, N8350);
nor NOR4 (N8353, N8336, N966, N3071, N3639);
nor NOR2 (N8354, N8349, N2276);
buf BUF1 (N8355, N8346);
buf BUF1 (N8356, N8345);
and AND3 (N8357, N8351, N1527, N4829);
not NOT1 (N8358, N8356);
buf BUF1 (N8359, N8323);
xor XOR2 (N8360, N8353, N3973);
and AND3 (N8361, N8352, N2427, N6375);
or OR3 (N8362, N8358, N6976, N5545);
or OR2 (N8363, N8332, N3666);
buf BUF1 (N8364, N8360);
and AND2 (N8365, N8362, N7388);
not NOT1 (N8366, N8364);
and AND3 (N8367, N8363, N4587, N1825);
buf BUF1 (N8368, N8367);
nand NAND3 (N8369, N8355, N3553, N1970);
buf BUF1 (N8370, N8348);
xor XOR2 (N8371, N8366, N6012);
nor NOR4 (N8372, N8357, N1996, N2363, N5736);
or OR2 (N8373, N8371, N2469);
not NOT1 (N8374, N8369);
not NOT1 (N8375, N8374);
and AND3 (N8376, N8372, N6974, N5927);
xor XOR2 (N8377, N8361, N7183);
not NOT1 (N8378, N8373);
or OR3 (N8379, N8368, N7938, N2960);
xor XOR2 (N8380, N8370, N864);
buf BUF1 (N8381, N8321);
or OR3 (N8382, N8359, N2110, N5287);
not NOT1 (N8383, N8378);
buf BUF1 (N8384, N8375);
xor XOR2 (N8385, N8382, N655);
not NOT1 (N8386, N8380);
and AND4 (N8387, N8379, N2750, N2848, N4382);
xor XOR2 (N8388, N8385, N7620);
and AND2 (N8389, N8388, N1262);
xor XOR2 (N8390, N8354, N1968);
not NOT1 (N8391, N8384);
or OR4 (N8392, N8377, N1993, N3240, N5232);
nor NOR2 (N8393, N8365, N8120);
not NOT1 (N8394, N8393);
xor XOR2 (N8395, N8383, N8062);
and AND3 (N8396, N8381, N800, N2601);
buf BUF1 (N8397, N8396);
xor XOR2 (N8398, N8392, N1441);
buf BUF1 (N8399, N8397);
not NOT1 (N8400, N8391);
or OR2 (N8401, N8399, N8372);
and AND3 (N8402, N8389, N2682, N5735);
nor NOR4 (N8403, N8390, N22, N2611, N5951);
nand NAND3 (N8404, N8402, N688, N6992);
not NOT1 (N8405, N8404);
xor XOR2 (N8406, N8401, N3789);
and AND4 (N8407, N8398, N3962, N955, N7273);
or OR2 (N8408, N8394, N7119);
nor NOR4 (N8409, N8400, N6084, N836, N4974);
nand NAND3 (N8410, N8409, N7796, N2449);
buf BUF1 (N8411, N8376);
nor NOR3 (N8412, N8386, N5122, N6582);
not NOT1 (N8413, N8411);
or OR4 (N8414, N8406, N3643, N4656, N2355);
buf BUF1 (N8415, N8408);
nor NOR4 (N8416, N8410, N323, N2053, N2237);
xor XOR2 (N8417, N8412, N1902);
buf BUF1 (N8418, N8405);
nand NAND4 (N8419, N8407, N6599, N8198, N5991);
xor XOR2 (N8420, N8416, N742);
buf BUF1 (N8421, N8420);
not NOT1 (N8422, N8403);
buf BUF1 (N8423, N8419);
nand NAND3 (N8424, N8423, N2605, N8038);
nor NOR2 (N8425, N8421, N2362);
nand NAND2 (N8426, N8395, N3275);
xor XOR2 (N8427, N8414, N3633);
nand NAND2 (N8428, N8413, N6599);
or OR4 (N8429, N8428, N4949, N546, N6756);
buf BUF1 (N8430, N8387);
xor XOR2 (N8431, N8417, N2740);
nand NAND2 (N8432, N8422, N506);
nor NOR4 (N8433, N8424, N4997, N240, N3196);
or OR2 (N8434, N8430, N5273);
buf BUF1 (N8435, N8426);
nand NAND3 (N8436, N8432, N6910, N734);
nand NAND2 (N8437, N8429, N1844);
buf BUF1 (N8438, N8437);
or OR4 (N8439, N8438, N4413, N5788, N5428);
nor NOR4 (N8440, N8415, N3781, N1434, N4019);
nor NOR3 (N8441, N8431, N1328, N3608);
buf BUF1 (N8442, N8418);
xor XOR2 (N8443, N8442, N7341);
or OR2 (N8444, N8427, N3830);
and AND2 (N8445, N8425, N5354);
buf BUF1 (N8446, N8436);
nand NAND2 (N8447, N8439, N3801);
and AND3 (N8448, N8444, N1745, N161);
not NOT1 (N8449, N8447);
xor XOR2 (N8450, N8446, N5352);
or OR4 (N8451, N8450, N4145, N943, N5745);
buf BUF1 (N8452, N8443);
or OR4 (N8453, N8445, N4888, N2741, N1540);
or OR4 (N8454, N8451, N4599, N8380, N2013);
buf BUF1 (N8455, N8433);
nor NOR4 (N8456, N8449, N6241, N1163, N5756);
and AND4 (N8457, N8448, N6809, N6938, N7291);
and AND2 (N8458, N8434, N4548);
not NOT1 (N8459, N8453);
and AND2 (N8460, N8440, N1038);
not NOT1 (N8461, N8441);
buf BUF1 (N8462, N8461);
buf BUF1 (N8463, N8457);
not NOT1 (N8464, N8462);
and AND2 (N8465, N8456, N7803);
nand NAND3 (N8466, N8458, N4573, N3559);
nor NOR3 (N8467, N8463, N5168, N4411);
buf BUF1 (N8468, N8452);
or OR3 (N8469, N8467, N1786, N202);
buf BUF1 (N8470, N8455);
nand NAND4 (N8471, N8469, N933, N3655, N8382);
xor XOR2 (N8472, N8466, N2570);
and AND2 (N8473, N8459, N7716);
nor NOR3 (N8474, N8471, N3886, N8391);
and AND2 (N8475, N8474, N1372);
not NOT1 (N8476, N8473);
nor NOR4 (N8477, N8468, N7547, N3036, N7804);
buf BUF1 (N8478, N8472);
not NOT1 (N8479, N8460);
nor NOR3 (N8480, N8435, N1820, N7267);
and AND4 (N8481, N8465, N1823, N5287, N6423);
buf BUF1 (N8482, N8480);
not NOT1 (N8483, N8478);
nor NOR3 (N8484, N8454, N6984, N5002);
xor XOR2 (N8485, N8475, N5848);
xor XOR2 (N8486, N8464, N1305);
or OR3 (N8487, N8470, N1666, N3145);
xor XOR2 (N8488, N8485, N6563);
or OR2 (N8489, N8479, N3901);
nor NOR3 (N8490, N8481, N6529, N52);
nor NOR2 (N8491, N8487, N7308);
nor NOR4 (N8492, N8489, N2009, N3491, N42);
nand NAND2 (N8493, N8488, N7481);
nand NAND3 (N8494, N8490, N7216, N3353);
or OR2 (N8495, N8486, N2188);
buf BUF1 (N8496, N8493);
and AND4 (N8497, N8496, N3231, N1794, N5270);
and AND3 (N8498, N8484, N3678, N6495);
and AND2 (N8499, N8483, N5534);
and AND4 (N8500, N8498, N4876, N3099, N7915);
nor NOR3 (N8501, N8482, N950, N1125);
nor NOR2 (N8502, N8497, N6635);
not NOT1 (N8503, N8495);
and AND3 (N8504, N8500, N5729, N6932);
and AND2 (N8505, N8502, N2095);
buf BUF1 (N8506, N8503);
buf BUF1 (N8507, N8492);
and AND2 (N8508, N8477, N3268);
buf BUF1 (N8509, N8494);
not NOT1 (N8510, N8504);
nand NAND3 (N8511, N8507, N3731, N7246);
nor NOR3 (N8512, N8511, N7397, N7507);
not NOT1 (N8513, N8491);
nand NAND2 (N8514, N8508, N8276);
buf BUF1 (N8515, N8509);
nor NOR4 (N8516, N8501, N3974, N3478, N6078);
buf BUF1 (N8517, N8514);
not NOT1 (N8518, N8517);
or OR3 (N8519, N8506, N1609, N4592);
xor XOR2 (N8520, N8513, N574);
nor NOR2 (N8521, N8499, N3802);
nor NOR2 (N8522, N8510, N7372);
or OR2 (N8523, N8512, N2257);
xor XOR2 (N8524, N8516, N5615);
or OR4 (N8525, N8522, N8276, N3394, N8204);
or OR4 (N8526, N8518, N793, N2328, N412);
buf BUF1 (N8527, N8476);
and AND2 (N8528, N8523, N6075);
buf BUF1 (N8529, N8519);
not NOT1 (N8530, N8525);
xor XOR2 (N8531, N8520, N2578);
or OR3 (N8532, N8526, N5714, N1161);
xor XOR2 (N8533, N8531, N3175);
not NOT1 (N8534, N8515);
nor NOR2 (N8535, N8528, N6403);
nor NOR2 (N8536, N8535, N146);
or OR3 (N8537, N8534, N3254, N4193);
nand NAND3 (N8538, N8532, N7952, N4771);
not NOT1 (N8539, N8536);
or OR2 (N8540, N8537, N7319);
buf BUF1 (N8541, N8538);
nor NOR3 (N8542, N8505, N7001, N1148);
nand NAND3 (N8543, N8539, N8042, N2919);
and AND2 (N8544, N8529, N6285);
nor NOR3 (N8545, N8524, N5287, N6237);
xor XOR2 (N8546, N8545, N6727);
not NOT1 (N8547, N8530);
xor XOR2 (N8548, N8533, N3093);
nand NAND3 (N8549, N8521, N3730, N4674);
nor NOR3 (N8550, N8546, N5996, N919);
buf BUF1 (N8551, N8547);
nand NAND2 (N8552, N8527, N7842);
nor NOR2 (N8553, N8540, N2933);
not NOT1 (N8554, N8551);
and AND4 (N8555, N8549, N8115, N1702, N4846);
nand NAND4 (N8556, N8543, N810, N2429, N472);
and AND3 (N8557, N8556, N377, N198);
and AND4 (N8558, N8541, N1087, N4526, N6934);
and AND4 (N8559, N8558, N4426, N5103, N8431);
and AND2 (N8560, N8542, N7159);
nor NOR3 (N8561, N8548, N6087, N6120);
and AND2 (N8562, N8550, N4287);
nor NOR2 (N8563, N8562, N1511);
and AND2 (N8564, N8554, N5680);
and AND2 (N8565, N8555, N8471);
or OR2 (N8566, N8559, N8083);
nand NAND4 (N8567, N8560, N736, N1075, N5838);
xor XOR2 (N8568, N8567, N8241);
or OR3 (N8569, N8553, N3717, N6266);
or OR2 (N8570, N8544, N2715);
and AND4 (N8571, N8564, N4420, N1787, N2260);
buf BUF1 (N8572, N8569);
not NOT1 (N8573, N8561);
xor XOR2 (N8574, N8563, N8392);
nor NOR4 (N8575, N8573, N8546, N7362, N2863);
and AND4 (N8576, N8572, N3360, N1529, N7136);
or OR3 (N8577, N8566, N3011, N5738);
nand NAND3 (N8578, N8557, N7119, N2673);
and AND3 (N8579, N8570, N2181, N2740);
buf BUF1 (N8580, N8571);
nor NOR3 (N8581, N8574, N8096, N5682);
nor NOR2 (N8582, N8578, N1195);
nand NAND3 (N8583, N8575, N5874, N4324);
nor NOR3 (N8584, N8552, N1763, N730);
or OR2 (N8585, N8583, N2285);
not NOT1 (N8586, N8585);
nor NOR4 (N8587, N8584, N1792, N8142, N4849);
not NOT1 (N8588, N8581);
buf BUF1 (N8589, N8579);
nor NOR4 (N8590, N8587, N7573, N8277, N4632);
buf BUF1 (N8591, N8577);
nand NAND4 (N8592, N8576, N1690, N5675, N4865);
or OR4 (N8593, N8590, N1612, N6949, N4106);
nor NOR2 (N8594, N8565, N6963);
not NOT1 (N8595, N8586);
nor NOR3 (N8596, N8588, N2530, N615);
not NOT1 (N8597, N8596);
nand NAND4 (N8598, N8580, N4710, N6093, N1174);
nor NOR2 (N8599, N8594, N3353);
and AND2 (N8600, N8568, N3036);
xor XOR2 (N8601, N8593, N3880);
and AND2 (N8602, N8600, N6604);
and AND2 (N8603, N8599, N2464);
buf BUF1 (N8604, N8589);
and AND4 (N8605, N8604, N2430, N4882, N567);
or OR3 (N8606, N8603, N3432, N7101);
or OR4 (N8607, N8591, N1171, N7730, N8303);
buf BUF1 (N8608, N8607);
xor XOR2 (N8609, N8608, N5620);
nor NOR2 (N8610, N8595, N8144);
buf BUF1 (N8611, N8592);
xor XOR2 (N8612, N8609, N2665);
xor XOR2 (N8613, N8612, N8181);
xor XOR2 (N8614, N8582, N1622);
xor XOR2 (N8615, N8610, N4163);
nand NAND3 (N8616, N8614, N1310, N3785);
buf BUF1 (N8617, N8601);
nand NAND4 (N8618, N8606, N3181, N470, N3600);
xor XOR2 (N8619, N8617, N2807);
xor XOR2 (N8620, N8615, N423);
xor XOR2 (N8621, N8598, N4542);
nor NOR3 (N8622, N8613, N1907, N8310);
or OR3 (N8623, N8605, N6688, N5569);
not NOT1 (N8624, N8621);
nand NAND3 (N8625, N8616, N6386, N3444);
buf BUF1 (N8626, N8623);
not NOT1 (N8627, N8626);
nor NOR4 (N8628, N8627, N2860, N3194, N6668);
nor NOR3 (N8629, N8611, N8207, N6950);
buf BUF1 (N8630, N8619);
nand NAND2 (N8631, N8618, N7375);
not NOT1 (N8632, N8622);
xor XOR2 (N8633, N8629, N2449);
buf BUF1 (N8634, N8620);
nor NOR3 (N8635, N8602, N1639, N3803);
nand NAND2 (N8636, N8597, N6386);
nor NOR3 (N8637, N8634, N975, N3107);
not NOT1 (N8638, N8633);
nand NAND4 (N8639, N8638, N4640, N3293, N8107);
and AND3 (N8640, N8624, N4235, N5129);
buf BUF1 (N8641, N8636);
nor NOR3 (N8642, N8641, N2717, N2475);
nor NOR3 (N8643, N8632, N310, N2815);
not NOT1 (N8644, N8630);
nor NOR3 (N8645, N8643, N4913, N6890);
buf BUF1 (N8646, N8645);
not NOT1 (N8647, N8637);
not NOT1 (N8648, N8644);
or OR3 (N8649, N8646, N7220, N6051);
buf BUF1 (N8650, N8628);
nor NOR4 (N8651, N8640, N6117, N7061, N8289);
or OR2 (N8652, N8642, N7750);
not NOT1 (N8653, N8647);
and AND2 (N8654, N8631, N2661);
and AND4 (N8655, N8648, N7104, N7685, N5448);
not NOT1 (N8656, N8653);
xor XOR2 (N8657, N8656, N1503);
not NOT1 (N8658, N8651);
not NOT1 (N8659, N8639);
not NOT1 (N8660, N8659);
nor NOR4 (N8661, N8635, N6524, N4436, N7733);
nand NAND3 (N8662, N8661, N5686, N6535);
nand NAND2 (N8663, N8655, N497);
xor XOR2 (N8664, N8658, N7492);
not NOT1 (N8665, N8625);
nand NAND2 (N8666, N8652, N3789);
or OR2 (N8667, N8657, N3420);
nand NAND3 (N8668, N8660, N4236, N4873);
buf BUF1 (N8669, N8665);
or OR4 (N8670, N8666, N6203, N5480, N4322);
not NOT1 (N8671, N8663);
and AND2 (N8672, N8654, N4576);
nor NOR4 (N8673, N8669, N1516, N2885, N6661);
buf BUF1 (N8674, N8664);
not NOT1 (N8675, N8662);
not NOT1 (N8676, N8673);
buf BUF1 (N8677, N8668);
not NOT1 (N8678, N8672);
and AND4 (N8679, N8677, N3883, N2507, N3937);
not NOT1 (N8680, N8675);
not NOT1 (N8681, N8670);
not NOT1 (N8682, N8676);
and AND2 (N8683, N8650, N1957);
or OR2 (N8684, N8671, N1651);
not NOT1 (N8685, N8683);
buf BUF1 (N8686, N8678);
not NOT1 (N8687, N8667);
buf BUF1 (N8688, N8681);
xor XOR2 (N8689, N8679, N7149);
buf BUF1 (N8690, N8685);
xor XOR2 (N8691, N8687, N5111);
nand NAND3 (N8692, N8649, N7175, N759);
buf BUF1 (N8693, N8680);
and AND3 (N8694, N8693, N4580, N3723);
or OR4 (N8695, N8688, N4548, N4618, N5770);
and AND3 (N8696, N8692, N1573, N8391);
not NOT1 (N8697, N8689);
xor XOR2 (N8698, N8694, N2523);
nor NOR3 (N8699, N8695, N3035, N2841);
buf BUF1 (N8700, N8691);
or OR3 (N8701, N8696, N5578, N7747);
or OR3 (N8702, N8698, N5193, N41);
or OR2 (N8703, N8702, N4958);
nor NOR3 (N8704, N8686, N2838, N5341);
not NOT1 (N8705, N8690);
nor NOR4 (N8706, N8699, N7056, N5944, N7236);
or OR3 (N8707, N8700, N2022, N6912);
nand NAND2 (N8708, N8707, N691);
xor XOR2 (N8709, N8706, N677);
not NOT1 (N8710, N8701);
nand NAND2 (N8711, N8704, N6944);
nor NOR3 (N8712, N8697, N8281, N6949);
buf BUF1 (N8713, N8684);
xor XOR2 (N8714, N8709, N2612);
buf BUF1 (N8715, N8705);
and AND4 (N8716, N8703, N5572, N317, N6349);
or OR2 (N8717, N8674, N7604);
xor XOR2 (N8718, N8714, N2953);
not NOT1 (N8719, N8713);
buf BUF1 (N8720, N8710);
and AND4 (N8721, N8712, N3509, N7015, N7958);
not NOT1 (N8722, N8711);
or OR2 (N8723, N8715, N2051);
xor XOR2 (N8724, N8721, N1916);
not NOT1 (N8725, N8720);
xor XOR2 (N8726, N8724, N698);
xor XOR2 (N8727, N8719, N1457);
nand NAND2 (N8728, N8717, N8631);
nor NOR2 (N8729, N8708, N8008);
or OR4 (N8730, N8729, N5588, N3555, N7667);
nand NAND4 (N8731, N8716, N7174, N6158, N5528);
buf BUF1 (N8732, N8718);
buf BUF1 (N8733, N8726);
xor XOR2 (N8734, N8728, N6439);
xor XOR2 (N8735, N8722, N5956);
nor NOR3 (N8736, N8733, N5857, N1850);
or OR2 (N8737, N8734, N7752);
or OR4 (N8738, N8732, N8142, N2663, N3714);
not NOT1 (N8739, N8731);
and AND2 (N8740, N8727, N1147);
not NOT1 (N8741, N8738);
buf BUF1 (N8742, N8740);
nand NAND3 (N8743, N8725, N3180, N5599);
and AND4 (N8744, N8735, N6905, N6813, N2661);
not NOT1 (N8745, N8743);
nand NAND4 (N8746, N8741, N784, N4476, N225);
buf BUF1 (N8747, N8730);
nand NAND4 (N8748, N8744, N1195, N5995, N2640);
nand NAND4 (N8749, N8682, N1460, N8524, N4407);
and AND3 (N8750, N8749, N3611, N8136);
and AND3 (N8751, N8748, N183, N1799);
nor NOR2 (N8752, N8739, N6818);
or OR2 (N8753, N8747, N641);
not NOT1 (N8754, N8750);
or OR2 (N8755, N8751, N1330);
not NOT1 (N8756, N8753);
and AND2 (N8757, N8755, N2645);
nand NAND4 (N8758, N8754, N772, N7749, N5570);
nor NOR4 (N8759, N8737, N8419, N5952, N899);
not NOT1 (N8760, N8742);
xor XOR2 (N8761, N8756, N411);
buf BUF1 (N8762, N8752);
nand NAND3 (N8763, N8762, N1375, N2270);
xor XOR2 (N8764, N8763, N2157);
nor NOR4 (N8765, N8760, N1916, N6725, N3262);
xor XOR2 (N8766, N8758, N7685);
not NOT1 (N8767, N8765);
nor NOR4 (N8768, N8723, N8598, N875, N6350);
and AND2 (N8769, N8767, N755);
buf BUF1 (N8770, N8736);
buf BUF1 (N8771, N8764);
xor XOR2 (N8772, N8771, N6320);
nand NAND3 (N8773, N8745, N5092, N5105);
xor XOR2 (N8774, N8766, N8540);
buf BUF1 (N8775, N8770);
nor NOR2 (N8776, N8775, N6747);
xor XOR2 (N8777, N8746, N1876);
nor NOR4 (N8778, N8772, N7952, N7055, N3929);
not NOT1 (N8779, N8776);
xor XOR2 (N8780, N8779, N4994);
not NOT1 (N8781, N8769);
buf BUF1 (N8782, N8781);
and AND4 (N8783, N8774, N7152, N1326, N1586);
nor NOR3 (N8784, N8759, N458, N1195);
not NOT1 (N8785, N8780);
nor NOR2 (N8786, N8768, N6880);
buf BUF1 (N8787, N8761);
nand NAND2 (N8788, N8787, N8778);
nor NOR4 (N8789, N4162, N3415, N585, N3177);
nand NAND4 (N8790, N8788, N102, N4568, N2201);
nor NOR3 (N8791, N8790, N3267, N6764);
nor NOR3 (N8792, N8783, N4003, N4631);
nand NAND3 (N8793, N8786, N4133, N1074);
or OR4 (N8794, N8777, N527, N4390, N5022);
nand NAND2 (N8795, N8785, N7200);
not NOT1 (N8796, N8784);
or OR4 (N8797, N8757, N6290, N6487, N3268);
not NOT1 (N8798, N8795);
nor NOR3 (N8799, N8798, N3973, N8783);
buf BUF1 (N8800, N8782);
not NOT1 (N8801, N8793);
buf BUF1 (N8802, N8797);
or OR3 (N8803, N8799, N4003, N3457);
xor XOR2 (N8804, N8800, N1697);
nand NAND3 (N8805, N8773, N8308, N5226);
and AND4 (N8806, N8803, N4471, N1914, N5037);
nor NOR2 (N8807, N8796, N2750);
xor XOR2 (N8808, N8801, N4550);
or OR2 (N8809, N8808, N5835);
xor XOR2 (N8810, N8806, N7828);
nor NOR3 (N8811, N8792, N1165, N6929);
xor XOR2 (N8812, N8807, N3353);
nor NOR4 (N8813, N8810, N1007, N5258, N68);
and AND2 (N8814, N8804, N6040);
nand NAND2 (N8815, N8812, N7863);
nand NAND4 (N8816, N8811, N775, N677, N3396);
buf BUF1 (N8817, N8815);
not NOT1 (N8818, N8809);
nor NOR2 (N8819, N8805, N1737);
nor NOR3 (N8820, N8814, N5298, N3714);
or OR3 (N8821, N8816, N1738, N3363);
and AND4 (N8822, N8789, N6918, N3601, N2211);
not NOT1 (N8823, N8821);
not NOT1 (N8824, N8802);
xor XOR2 (N8825, N8818, N6512);
not NOT1 (N8826, N8813);
or OR4 (N8827, N8820, N3154, N6984, N320);
or OR2 (N8828, N8794, N5830);
and AND3 (N8829, N8825, N7880, N3352);
buf BUF1 (N8830, N8822);
nand NAND4 (N8831, N8823, N8800, N2113, N3134);
xor XOR2 (N8832, N8826, N2055);
and AND4 (N8833, N8830, N964, N2920, N2856);
or OR3 (N8834, N8827, N5507, N7660);
nor NOR4 (N8835, N8791, N3810, N984, N374);
buf BUF1 (N8836, N8833);
nor NOR2 (N8837, N8817, N3622);
buf BUF1 (N8838, N8836);
buf BUF1 (N8839, N8819);
nor NOR4 (N8840, N8829, N3359, N2643, N1398);
and AND2 (N8841, N8831, N3921);
nor NOR4 (N8842, N8839, N2298, N7695, N6746);
nor NOR3 (N8843, N8837, N7413, N2477);
nor NOR4 (N8844, N8842, N4134, N4885, N2367);
nor NOR3 (N8845, N8834, N1360, N4494);
not NOT1 (N8846, N8843);
nor NOR3 (N8847, N8840, N5539, N2411);
xor XOR2 (N8848, N8832, N162);
xor XOR2 (N8849, N8845, N6517);
buf BUF1 (N8850, N8849);
nand NAND3 (N8851, N8848, N5523, N165);
and AND2 (N8852, N8844, N7334);
or OR4 (N8853, N8852, N400, N8793, N8664);
xor XOR2 (N8854, N8846, N3785);
xor XOR2 (N8855, N8824, N7654);
not NOT1 (N8856, N8835);
not NOT1 (N8857, N8851);
buf BUF1 (N8858, N8838);
buf BUF1 (N8859, N8855);
not NOT1 (N8860, N8856);
or OR4 (N8861, N8828, N5568, N8829, N8135);
and AND4 (N8862, N8850, N6925, N3246, N7536);
and AND4 (N8863, N8854, N2094, N3218, N8127);
nor NOR2 (N8864, N8858, N3265);
and AND4 (N8865, N8853, N5876, N190, N2854);
xor XOR2 (N8866, N8861, N3049);
nand NAND2 (N8867, N8866, N5735);
nand NAND3 (N8868, N8860, N3433, N7226);
and AND3 (N8869, N8868, N6722, N6060);
and AND2 (N8870, N8847, N1979);
nor NOR3 (N8871, N8869, N5222, N8803);
or OR3 (N8872, N8857, N5288, N2746);
buf BUF1 (N8873, N8863);
and AND2 (N8874, N8864, N4449);
buf BUF1 (N8875, N8870);
not NOT1 (N8876, N8873);
xor XOR2 (N8877, N8871, N2586);
xor XOR2 (N8878, N8859, N3032);
not NOT1 (N8879, N8841);
nor NOR3 (N8880, N8877, N1620, N1786);
buf BUF1 (N8881, N8865);
and AND4 (N8882, N8862, N7117, N1262, N3520);
or OR2 (N8883, N8879, N3032);
xor XOR2 (N8884, N8874, N2988);
xor XOR2 (N8885, N8881, N6279);
and AND2 (N8886, N8872, N6515);
and AND3 (N8887, N8884, N6184, N2891);
nor NOR4 (N8888, N8876, N4490, N1961, N5558);
nand NAND4 (N8889, N8878, N4238, N6675, N6276);
not NOT1 (N8890, N8880);
nor NOR4 (N8891, N8875, N4412, N5863, N3578);
or OR3 (N8892, N8887, N5458, N2119);
nor NOR2 (N8893, N8889, N1483);
nand NAND2 (N8894, N8892, N181);
buf BUF1 (N8895, N8885);
buf BUF1 (N8896, N8888);
xor XOR2 (N8897, N8867, N4905);
buf BUF1 (N8898, N8893);
or OR4 (N8899, N8891, N3669, N3236, N6012);
nand NAND4 (N8900, N8890, N6284, N5768, N7195);
nand NAND4 (N8901, N8886, N4467, N5713, N8058);
xor XOR2 (N8902, N8896, N2439);
nand NAND2 (N8903, N8901, N2098);
or OR2 (N8904, N8882, N5080);
buf BUF1 (N8905, N8903);
nand NAND2 (N8906, N8900, N6495);
and AND4 (N8907, N8898, N5391, N5854, N4032);
buf BUF1 (N8908, N8883);
nand NAND4 (N8909, N8902, N3579, N5797, N6372);
xor XOR2 (N8910, N8906, N7565);
and AND3 (N8911, N8895, N7679, N2290);
buf BUF1 (N8912, N8911);
and AND4 (N8913, N8904, N452, N7572, N2938);
nor NOR3 (N8914, N8894, N1449, N5975);
nor NOR2 (N8915, N8909, N2767);
nand NAND2 (N8916, N8905, N1558);
buf BUF1 (N8917, N8912);
not NOT1 (N8918, N8914);
not NOT1 (N8919, N8907);
xor XOR2 (N8920, N8919, N4835);
not NOT1 (N8921, N8899);
nand NAND3 (N8922, N8897, N7799, N708);
nand NAND4 (N8923, N8921, N6060, N6429, N4600);
not NOT1 (N8924, N8913);
buf BUF1 (N8925, N8917);
nand NAND2 (N8926, N8923, N8661);
xor XOR2 (N8927, N8916, N3500);
nor NOR4 (N8928, N8908, N1865, N6342, N7150);
or OR4 (N8929, N8925, N705, N7453, N8621);
buf BUF1 (N8930, N8927);
or OR2 (N8931, N8918, N7447);
buf BUF1 (N8932, N8922);
nand NAND2 (N8933, N8932, N7394);
or OR2 (N8934, N8926, N3930);
nand NAND2 (N8935, N8929, N246);
or OR3 (N8936, N8935, N1560, N3218);
xor XOR2 (N8937, N8915, N6218);
nor NOR3 (N8938, N8936, N2762, N3848);
xor XOR2 (N8939, N8938, N6810);
buf BUF1 (N8940, N8920);
xor XOR2 (N8941, N8939, N6219);
and AND2 (N8942, N8924, N4215);
xor XOR2 (N8943, N8931, N3161);
or OR4 (N8944, N8941, N2475, N5257, N3988);
nor NOR4 (N8945, N8942, N7356, N8016, N6687);
and AND2 (N8946, N8933, N8789);
and AND4 (N8947, N8910, N8761, N6268, N4522);
and AND3 (N8948, N8928, N7344, N2513);
nand NAND3 (N8949, N8946, N6294, N1387);
xor XOR2 (N8950, N8937, N1138);
xor XOR2 (N8951, N8947, N2083);
and AND4 (N8952, N8930, N2347, N4807, N1850);
nor NOR2 (N8953, N8949, N6381);
xor XOR2 (N8954, N8940, N5278);
buf BUF1 (N8955, N8950);
xor XOR2 (N8956, N8954, N5859);
not NOT1 (N8957, N8951);
xor XOR2 (N8958, N8956, N2579);
nor NOR2 (N8959, N8943, N6129);
nor NOR3 (N8960, N8959, N7647, N6831);
and AND2 (N8961, N8934, N2788);
xor XOR2 (N8962, N8953, N5662);
and AND2 (N8963, N8952, N6746);
and AND2 (N8964, N8944, N2048);
and AND3 (N8965, N8945, N6786, N4034);
buf BUF1 (N8966, N8963);
not NOT1 (N8967, N8957);
xor XOR2 (N8968, N8960, N2409);
nor NOR4 (N8969, N8968, N3792, N8962, N3268);
nor NOR4 (N8970, N4869, N8831, N4746, N4628);
xor XOR2 (N8971, N8961, N2489);
buf BUF1 (N8972, N8970);
xor XOR2 (N8973, N8965, N4103);
or OR4 (N8974, N8967, N7694, N1815, N2861);
nor NOR4 (N8975, N8969, N7897, N4324, N8156);
or OR3 (N8976, N8971, N6036, N6539);
buf BUF1 (N8977, N8964);
nand NAND2 (N8978, N8975, N8312);
nor NOR3 (N8979, N8976, N7530, N8371);
nand NAND2 (N8980, N8979, N3229);
and AND3 (N8981, N8974, N4604, N957);
xor XOR2 (N8982, N8972, N8212);
buf BUF1 (N8983, N8977);
nand NAND3 (N8984, N8966, N2972, N4206);
not NOT1 (N8985, N8982);
or OR2 (N8986, N8955, N8832);
buf BUF1 (N8987, N8981);
and AND4 (N8988, N8987, N1697, N1590, N1258);
or OR2 (N8989, N8984, N5905);
xor XOR2 (N8990, N8978, N6472);
nand NAND3 (N8991, N8990, N7288, N2062);
xor XOR2 (N8992, N8986, N2043);
nand NAND4 (N8993, N8992, N5519, N6677, N3127);
nand NAND4 (N8994, N8980, N7358, N7302, N7955);
or OR3 (N8995, N8988, N55, N7015);
nand NAND4 (N8996, N8989, N5865, N3146, N6652);
nand NAND4 (N8997, N8996, N7120, N6620, N8440);
xor XOR2 (N8998, N8985, N2204);
nand NAND2 (N8999, N8995, N4818);
nor NOR3 (N9000, N8948, N2341, N648);
nand NAND3 (N9001, N9000, N6027, N8685);
and AND4 (N9002, N8998, N7625, N8264, N5911);
buf BUF1 (N9003, N9002);
xor XOR2 (N9004, N8973, N1997);
nor NOR3 (N9005, N8994, N667, N5819);
buf BUF1 (N9006, N8993);
buf BUF1 (N9007, N8991);
not NOT1 (N9008, N8997);
nand NAND3 (N9009, N9006, N3123, N7647);
xor XOR2 (N9010, N9001, N3889);
not NOT1 (N9011, N8983);
nor NOR2 (N9012, N8958, N5364);
nand NAND3 (N9013, N9010, N498, N2366);
and AND4 (N9014, N9005, N1092, N7738, N3895);
and AND3 (N9015, N9007, N5320, N5207);
buf BUF1 (N9016, N9011);
or OR2 (N9017, N9016, N2724);
xor XOR2 (N9018, N9009, N5753);
not NOT1 (N9019, N9015);
nand NAND2 (N9020, N9008, N4086);
buf BUF1 (N9021, N9004);
nand NAND4 (N9022, N9021, N4428, N5046, N1986);
or OR2 (N9023, N9019, N4393);
xor XOR2 (N9024, N9003, N3548);
nor NOR3 (N9025, N9014, N1881, N3594);
and AND4 (N9026, N9018, N3440, N8107, N4416);
buf BUF1 (N9027, N9012);
not NOT1 (N9028, N9027);
nand NAND4 (N9029, N9023, N37, N6023, N8656);
buf BUF1 (N9030, N9029);
nor NOR3 (N9031, N9013, N3742, N303);
not NOT1 (N9032, N9024);
buf BUF1 (N9033, N9020);
nand NAND3 (N9034, N9032, N2219, N1760);
or OR3 (N9035, N9034, N6821, N101);
and AND2 (N9036, N9030, N4954);
or OR2 (N9037, N9022, N6369);
nor NOR4 (N9038, N9026, N1196, N4965, N4158);
buf BUF1 (N9039, N9033);
not NOT1 (N9040, N9037);
buf BUF1 (N9041, N9036);
or OR4 (N9042, N9039, N1483, N5362, N2149);
and AND2 (N9043, N9042, N6379);
not NOT1 (N9044, N9040);
and AND2 (N9045, N9038, N7195);
and AND2 (N9046, N9035, N4179);
nor NOR4 (N9047, N9046, N7288, N7171, N6580);
nor NOR3 (N9048, N8999, N8235, N2891);
xor XOR2 (N9049, N9044, N8861);
and AND4 (N9050, N9041, N1078, N3993, N8468);
nor NOR4 (N9051, N9043, N2966, N2932, N6725);
buf BUF1 (N9052, N9047);
or OR2 (N9053, N9017, N273);
xor XOR2 (N9054, N9045, N6646);
xor XOR2 (N9055, N9031, N5057);
nand NAND2 (N9056, N9025, N2369);
buf BUF1 (N9057, N9055);
not NOT1 (N9058, N9049);
and AND3 (N9059, N9053, N706, N230);
nor NOR4 (N9060, N9059, N1715, N3586, N4726);
buf BUF1 (N9061, N9060);
and AND2 (N9062, N9028, N7600);
nor NOR2 (N9063, N9054, N2468);
nand NAND2 (N9064, N9063, N4542);
xor XOR2 (N9065, N9050, N5334);
and AND2 (N9066, N9058, N5904);
not NOT1 (N9067, N9065);
not NOT1 (N9068, N9056);
or OR2 (N9069, N9067, N1359);
not NOT1 (N9070, N9061);
xor XOR2 (N9071, N9066, N1889);
nor NOR2 (N9072, N9057, N3819);
nand NAND2 (N9073, N9064, N3878);
buf BUF1 (N9074, N9048);
nand NAND3 (N9075, N9071, N2017, N5363);
or OR4 (N9076, N9073, N2745, N6752, N4671);
buf BUF1 (N9077, N9074);
buf BUF1 (N9078, N9051);
not NOT1 (N9079, N9052);
nand NAND4 (N9080, N9077, N5262, N3487, N4734);
nand NAND4 (N9081, N9068, N7334, N4505, N7336);
nor NOR2 (N9082, N9079, N3279);
nor NOR2 (N9083, N9082, N867);
xor XOR2 (N9084, N9081, N7723);
not NOT1 (N9085, N9080);
buf BUF1 (N9086, N9076);
or OR3 (N9087, N9078, N3524, N3936);
nand NAND3 (N9088, N9086, N8451, N2015);
xor XOR2 (N9089, N9084, N6332);
buf BUF1 (N9090, N9072);
nand NAND2 (N9091, N9083, N3382);
not NOT1 (N9092, N9070);
buf BUF1 (N9093, N9085);
nand NAND2 (N9094, N9089, N4524);
not NOT1 (N9095, N9092);
buf BUF1 (N9096, N9075);
or OR4 (N9097, N9069, N8612, N5010, N1577);
nand NAND4 (N9098, N9095, N2354, N7763, N3730);
not NOT1 (N9099, N9093);
xor XOR2 (N9100, N9097, N1973);
and AND3 (N9101, N9099, N1007, N5850);
or OR3 (N9102, N9101, N6506, N90);
or OR3 (N9103, N9100, N6585, N5582);
and AND3 (N9104, N9087, N1122, N8611);
buf BUF1 (N9105, N9090);
nor NOR4 (N9106, N9104, N8605, N6092, N1014);
not NOT1 (N9107, N9088);
and AND4 (N9108, N9103, N2549, N7750, N7456);
and AND4 (N9109, N9091, N999, N7637, N7061);
buf BUF1 (N9110, N9098);
not NOT1 (N9111, N9110);
and AND3 (N9112, N9111, N5546, N7058);
and AND4 (N9113, N9096, N8962, N4225, N5562);
nand NAND2 (N9114, N9112, N5947);
xor XOR2 (N9115, N9062, N6985);
and AND4 (N9116, N9106, N493, N6421, N1758);
or OR2 (N9117, N9116, N3798);
not NOT1 (N9118, N9117);
nor NOR3 (N9119, N9105, N2665, N2375);
nor NOR4 (N9120, N9115, N7485, N5641, N3136);
xor XOR2 (N9121, N9120, N6799);
buf BUF1 (N9122, N9107);
buf BUF1 (N9123, N9109);
buf BUF1 (N9124, N9108);
or OR2 (N9125, N9118, N2760);
buf BUF1 (N9126, N9094);
buf BUF1 (N9127, N9114);
and AND3 (N9128, N9124, N6804, N4339);
xor XOR2 (N9129, N9127, N6869);
nand NAND4 (N9130, N9121, N2115, N3805, N2789);
buf BUF1 (N9131, N9122);
nor NOR4 (N9132, N9125, N5614, N5159, N2291);
nor NOR3 (N9133, N9119, N1833, N7085);
buf BUF1 (N9134, N9133);
or OR4 (N9135, N9126, N7411, N718, N7460);
xor XOR2 (N9136, N9113, N772);
nor NOR2 (N9137, N9129, N6855);
nand NAND3 (N9138, N9136, N5789, N4420);
buf BUF1 (N9139, N9137);
nand NAND2 (N9140, N9138, N619);
and AND3 (N9141, N9132, N3138, N8556);
nand NAND3 (N9142, N9123, N2758, N7691);
nand NAND2 (N9143, N9102, N982);
not NOT1 (N9144, N9141);
buf BUF1 (N9145, N9142);
buf BUF1 (N9146, N9139);
xor XOR2 (N9147, N9130, N8143);
xor XOR2 (N9148, N9131, N8206);
buf BUF1 (N9149, N9146);
nor NOR3 (N9150, N9144, N591, N2758);
nor NOR4 (N9151, N9150, N3962, N319, N5809);
buf BUF1 (N9152, N9147);
and AND3 (N9153, N9143, N1297, N3273);
buf BUF1 (N9154, N9140);
buf BUF1 (N9155, N9148);
or OR3 (N9156, N9152, N8978, N2305);
nor NOR4 (N9157, N9149, N7538, N3172, N8756);
or OR2 (N9158, N9151, N6037);
not NOT1 (N9159, N9156);
and AND3 (N9160, N9158, N804, N737);
nand NAND3 (N9161, N9128, N4726, N6818);
and AND4 (N9162, N9145, N3614, N2957, N3864);
buf BUF1 (N9163, N9153);
not NOT1 (N9164, N9159);
nand NAND4 (N9165, N9161, N7114, N7782, N1419);
buf BUF1 (N9166, N9157);
and AND3 (N9167, N9134, N2651, N4730);
xor XOR2 (N9168, N9164, N201);
and AND2 (N9169, N9135, N2597);
nor NOR2 (N9170, N9167, N7822);
nand NAND3 (N9171, N9165, N2991, N6886);
nor NOR2 (N9172, N9170, N3393);
buf BUF1 (N9173, N9169);
nand NAND4 (N9174, N9171, N338, N2636, N921);
and AND2 (N9175, N9173, N8886);
not NOT1 (N9176, N9160);
or OR2 (N9177, N9176, N4358);
xor XOR2 (N9178, N9172, N948);
not NOT1 (N9179, N9163);
xor XOR2 (N9180, N9162, N7198);
nand NAND2 (N9181, N9155, N1351);
xor XOR2 (N9182, N9181, N7011);
or OR4 (N9183, N9182, N7045, N1073, N487);
buf BUF1 (N9184, N9179);
not NOT1 (N9185, N9175);
xor XOR2 (N9186, N9185, N3917);
nor NOR2 (N9187, N9186, N4602);
and AND4 (N9188, N9187, N4682, N2117, N7485);
buf BUF1 (N9189, N9168);
or OR2 (N9190, N9180, N8482);
nor NOR3 (N9191, N9178, N2420, N6254);
or OR2 (N9192, N9184, N767);
buf BUF1 (N9193, N9166);
or OR4 (N9194, N9188, N248, N1339, N2035);
nand NAND4 (N9195, N9154, N3260, N8188, N7657);
xor XOR2 (N9196, N9189, N7838);
nand NAND2 (N9197, N9191, N8205);
and AND3 (N9198, N9174, N4028, N6355);
buf BUF1 (N9199, N9177);
or OR3 (N9200, N9192, N8911, N7387);
nor NOR4 (N9201, N9190, N5182, N5070, N7868);
buf BUF1 (N9202, N9200);
not NOT1 (N9203, N9183);
not NOT1 (N9204, N9194);
buf BUF1 (N9205, N9197);
buf BUF1 (N9206, N9203);
or OR4 (N9207, N9201, N576, N6126, N6750);
xor XOR2 (N9208, N9205, N5448);
or OR2 (N9209, N9206, N5277);
and AND2 (N9210, N9198, N7385);
not NOT1 (N9211, N9193);
not NOT1 (N9212, N9207);
nand NAND2 (N9213, N9209, N1111);
xor XOR2 (N9214, N9210, N5422);
nor NOR4 (N9215, N9208, N3432, N226, N1222);
nand NAND4 (N9216, N9214, N3816, N2920, N8262);
and AND4 (N9217, N9202, N7668, N7263, N5141);
nor NOR4 (N9218, N9212, N484, N5443, N2722);
nand NAND4 (N9219, N9211, N5928, N4299, N354);
and AND4 (N9220, N9218, N998, N4046, N3798);
or OR3 (N9221, N9217, N5547, N8358);
xor XOR2 (N9222, N9213, N8138);
xor XOR2 (N9223, N9220, N5257);
xor XOR2 (N9224, N9219, N7035);
nor NOR3 (N9225, N9224, N2677, N5214);
xor XOR2 (N9226, N9199, N4133);
nor NOR2 (N9227, N9225, N8218);
and AND4 (N9228, N9227, N5654, N5987, N7789);
or OR4 (N9229, N9228, N1124, N6417, N5067);
nor NOR4 (N9230, N9223, N3369, N7709, N7415);
nand NAND3 (N9231, N9215, N3406, N2003);
nand NAND4 (N9232, N9222, N6513, N393, N4380);
or OR3 (N9233, N9226, N7963, N2239);
buf BUF1 (N9234, N9221);
nand NAND3 (N9235, N9229, N2004, N464);
nand NAND2 (N9236, N9234, N939);
nand NAND3 (N9237, N9231, N8262, N6251);
and AND4 (N9238, N9232, N2934, N7101, N2742);
buf BUF1 (N9239, N9196);
xor XOR2 (N9240, N9238, N6799);
buf BUF1 (N9241, N9204);
or OR2 (N9242, N9241, N1133);
xor XOR2 (N9243, N9195, N3891);
buf BUF1 (N9244, N9237);
not NOT1 (N9245, N9233);
buf BUF1 (N9246, N9243);
nand NAND4 (N9247, N9242, N8389, N1038, N3704);
and AND4 (N9248, N9245, N5114, N5890, N6283);
and AND3 (N9249, N9246, N9176, N5039);
and AND3 (N9250, N9244, N3883, N4747);
buf BUF1 (N9251, N9240);
buf BUF1 (N9252, N9239);
nor NOR2 (N9253, N9248, N6999);
buf BUF1 (N9254, N9235);
nor NOR3 (N9255, N9230, N9205, N5604);
xor XOR2 (N9256, N9216, N6548);
buf BUF1 (N9257, N9253);
nor NOR4 (N9258, N9255, N8399, N6066, N4674);
nor NOR3 (N9259, N9252, N4114, N3292);
and AND4 (N9260, N9250, N7466, N3474, N4887);
nand NAND4 (N9261, N9251, N6306, N6731, N5819);
buf BUF1 (N9262, N9256);
nor NOR3 (N9263, N9258, N126, N2962);
nor NOR4 (N9264, N9261, N2134, N3180, N8048);
nand NAND4 (N9265, N9257, N843, N7090, N565);
nand NAND3 (N9266, N9259, N232, N7454);
and AND4 (N9267, N9266, N8275, N5420, N3697);
and AND4 (N9268, N9236, N4423, N5500, N8892);
nor NOR3 (N9269, N9249, N2934, N6187);
buf BUF1 (N9270, N9260);
nand NAND2 (N9271, N9268, N7022);
and AND3 (N9272, N9267, N4248, N2347);
nand NAND2 (N9273, N9272, N8392);
nand NAND2 (N9274, N9264, N6550);
not NOT1 (N9275, N9274);
nor NOR4 (N9276, N9270, N7813, N4800, N7707);
buf BUF1 (N9277, N9254);
and AND2 (N9278, N9271, N8536);
not NOT1 (N9279, N9276);
or OR3 (N9280, N9277, N2113, N6484);
nor NOR3 (N9281, N9275, N4736, N5797);
or OR2 (N9282, N9281, N9162);
or OR3 (N9283, N9273, N5934, N2192);
not NOT1 (N9284, N9280);
or OR4 (N9285, N9282, N6482, N7650, N5055);
or OR3 (N9286, N9263, N1398, N262);
not NOT1 (N9287, N9286);
nor NOR3 (N9288, N9269, N3646, N5638);
or OR4 (N9289, N9284, N3920, N3996, N4973);
not NOT1 (N9290, N9285);
nand NAND3 (N9291, N9278, N7092, N2742);
not NOT1 (N9292, N9289);
xor XOR2 (N9293, N9265, N5977);
and AND3 (N9294, N9293, N164, N4993);
nor NOR3 (N9295, N9291, N9023, N3273);
buf BUF1 (N9296, N9295);
xor XOR2 (N9297, N9247, N8740);
and AND4 (N9298, N9297, N4109, N5055, N6539);
and AND3 (N9299, N9290, N2601, N594);
xor XOR2 (N9300, N9296, N7228);
and AND2 (N9301, N9298, N1346);
and AND4 (N9302, N9292, N8658, N2683, N6615);
xor XOR2 (N9303, N9287, N4512);
and AND4 (N9304, N9288, N7227, N6418, N85);
nor NOR3 (N9305, N9303, N6139, N5291);
buf BUF1 (N9306, N9283);
and AND3 (N9307, N9299, N4071, N3401);
or OR2 (N9308, N9305, N9232);
not NOT1 (N9309, N9307);
nand NAND4 (N9310, N9309, N5666, N8219, N3096);
not NOT1 (N9311, N9294);
or OR3 (N9312, N9302, N7636, N7316);
not NOT1 (N9313, N9306);
and AND2 (N9314, N9310, N919);
not NOT1 (N9315, N9312);
xor XOR2 (N9316, N9279, N5719);
nand NAND3 (N9317, N9314, N954, N8870);
buf BUF1 (N9318, N9300);
buf BUF1 (N9319, N9315);
not NOT1 (N9320, N9304);
not NOT1 (N9321, N9320);
and AND3 (N9322, N9317, N96, N62);
nand NAND2 (N9323, N9301, N2616);
not NOT1 (N9324, N9319);
nand NAND3 (N9325, N9322, N1618, N4266);
xor XOR2 (N9326, N9311, N8467);
or OR4 (N9327, N9313, N7408, N4989, N2101);
nand NAND3 (N9328, N9324, N3517, N5142);
or OR4 (N9329, N9328, N1933, N8423, N2625);
xor XOR2 (N9330, N9326, N6121);
nand NAND4 (N9331, N9327, N8139, N4833, N6040);
xor XOR2 (N9332, N9318, N7733);
xor XOR2 (N9333, N9331, N5352);
buf BUF1 (N9334, N9321);
and AND4 (N9335, N9308, N7570, N8612, N3811);
and AND2 (N9336, N9335, N5664);
buf BUF1 (N9337, N9333);
buf BUF1 (N9338, N9316);
nor NOR4 (N9339, N9332, N3078, N8956, N3807);
buf BUF1 (N9340, N9330);
not NOT1 (N9341, N9338);
nand NAND2 (N9342, N9323, N8024);
nand NAND4 (N9343, N9337, N9257, N613, N4528);
and AND4 (N9344, N9334, N3861, N240, N1662);
xor XOR2 (N9345, N9329, N2074);
or OR2 (N9346, N9340, N5375);
and AND4 (N9347, N9262, N8369, N360, N3699);
buf BUF1 (N9348, N9343);
xor XOR2 (N9349, N9344, N5713);
not NOT1 (N9350, N9341);
buf BUF1 (N9351, N9348);
xor XOR2 (N9352, N9339, N2676);
and AND4 (N9353, N9349, N6103, N8623, N3517);
xor XOR2 (N9354, N9352, N2314);
xor XOR2 (N9355, N9345, N2217);
not NOT1 (N9356, N9354);
buf BUF1 (N9357, N9347);
xor XOR2 (N9358, N9351, N1706);
and AND2 (N9359, N9346, N5633);
or OR4 (N9360, N9359, N3260, N8416, N1860);
nor NOR4 (N9361, N9357, N2745, N6947, N447);
and AND4 (N9362, N9361, N4958, N4596, N4977);
nand NAND2 (N9363, N9336, N5397);
buf BUF1 (N9364, N9360);
xor XOR2 (N9365, N9353, N1868);
nor NOR4 (N9366, N9325, N1395, N7273, N1232);
and AND2 (N9367, N9365, N9298);
nand NAND4 (N9368, N9364, N8446, N3513, N9345);
nand NAND4 (N9369, N9368, N1914, N4807, N2565);
and AND2 (N9370, N9363, N6152);
or OR3 (N9371, N9366, N151, N3151);
not NOT1 (N9372, N9350);
not NOT1 (N9373, N9371);
nand NAND2 (N9374, N9367, N2394);
buf BUF1 (N9375, N9369);
nand NAND2 (N9376, N9375, N8863);
or OR4 (N9377, N9373, N6729, N3481, N6348);
or OR4 (N9378, N9374, N1886, N8562, N2473);
or OR4 (N9379, N9376, N320, N1510, N6105);
nor NOR3 (N9380, N9370, N8452, N4276);
not NOT1 (N9381, N9356);
not NOT1 (N9382, N9378);
and AND4 (N9383, N9362, N6883, N7645, N1519);
or OR4 (N9384, N9379, N1290, N6582, N3536);
buf BUF1 (N9385, N9384);
nand NAND3 (N9386, N9380, N7396, N249);
xor XOR2 (N9387, N9385, N8553);
nand NAND4 (N9388, N9372, N2728, N5650, N593);
not NOT1 (N9389, N9387);
buf BUF1 (N9390, N9386);
xor XOR2 (N9391, N9358, N7994);
and AND3 (N9392, N9381, N7116, N6867);
nor NOR3 (N9393, N9382, N7286, N817);
or OR4 (N9394, N9355, N5701, N8689, N1334);
xor XOR2 (N9395, N9392, N6979);
nor NOR2 (N9396, N9393, N843);
not NOT1 (N9397, N9388);
nor NOR2 (N9398, N9396, N4485);
xor XOR2 (N9399, N9342, N3826);
nand NAND3 (N9400, N9398, N8198, N9208);
xor XOR2 (N9401, N9397, N4748);
nand NAND3 (N9402, N9377, N3985, N1936);
nand NAND2 (N9403, N9399, N153);
or OR4 (N9404, N9389, N5221, N1208, N1150);
nor NOR2 (N9405, N9401, N4984);
nand NAND3 (N9406, N9405, N1067, N8470);
not NOT1 (N9407, N9383);
xor XOR2 (N9408, N9400, N3484);
nand NAND3 (N9409, N9407, N9074, N2083);
and AND4 (N9410, N9404, N7420, N3747, N9063);
nor NOR4 (N9411, N9409, N6950, N4943, N1826);
nor NOR3 (N9412, N9406, N7795, N3960);
buf BUF1 (N9413, N9394);
nand NAND2 (N9414, N9402, N8312);
not NOT1 (N9415, N9412);
buf BUF1 (N9416, N9395);
nor NOR3 (N9417, N9416, N537, N3581);
and AND2 (N9418, N9403, N1485);
xor XOR2 (N9419, N9408, N7927);
and AND4 (N9420, N9418, N2769, N3209, N4567);
nor NOR4 (N9421, N9391, N8297, N4623, N5871);
and AND3 (N9422, N9419, N3497, N8478);
and AND3 (N9423, N9422, N4475, N1716);
xor XOR2 (N9424, N9410, N8139);
nand NAND4 (N9425, N9415, N3883, N8122, N9228);
buf BUF1 (N9426, N9423);
not NOT1 (N9427, N9420);
and AND2 (N9428, N9425, N9337);
xor XOR2 (N9429, N9421, N6720);
or OR4 (N9430, N9428, N7367, N5784, N4112);
xor XOR2 (N9431, N9426, N3218);
not NOT1 (N9432, N9413);
and AND3 (N9433, N9431, N4191, N6048);
not NOT1 (N9434, N9424);
and AND2 (N9435, N9414, N8504);
buf BUF1 (N9436, N9390);
not NOT1 (N9437, N9436);
xor XOR2 (N9438, N9417, N7434);
nor NOR4 (N9439, N9435, N2197, N727, N469);
buf BUF1 (N9440, N9429);
nand NAND3 (N9441, N9437, N7284, N1623);
buf BUF1 (N9442, N9411);
nand NAND2 (N9443, N9439, N6163);
nand NAND3 (N9444, N9443, N936, N3017);
nor NOR3 (N9445, N9432, N5150, N2229);
xor XOR2 (N9446, N9430, N8436);
nor NOR2 (N9447, N9440, N5226);
buf BUF1 (N9448, N9438);
xor XOR2 (N9449, N9434, N1581);
not NOT1 (N9450, N9442);
not NOT1 (N9451, N9433);
nor NOR3 (N9452, N9451, N4342, N7640);
nor NOR2 (N9453, N9448, N618);
xor XOR2 (N9454, N9452, N5639);
nand NAND3 (N9455, N9446, N7392, N5949);
or OR3 (N9456, N9441, N8950, N871);
nand NAND3 (N9457, N9449, N8201, N101);
or OR2 (N9458, N9427, N133);
and AND2 (N9459, N9458, N9033);
buf BUF1 (N9460, N9455);
xor XOR2 (N9461, N9456, N160);
or OR2 (N9462, N9447, N4143);
buf BUF1 (N9463, N9454);
buf BUF1 (N9464, N9453);
not NOT1 (N9465, N9450);
nand NAND4 (N9466, N9461, N5093, N7707, N5638);
or OR4 (N9467, N9457, N7909, N807, N6079);
xor XOR2 (N9468, N9462, N8636);
xor XOR2 (N9469, N9465, N3082);
or OR2 (N9470, N9467, N6781);
not NOT1 (N9471, N9459);
or OR4 (N9472, N9445, N266, N2023, N4082);
nand NAND2 (N9473, N9470, N4051);
and AND4 (N9474, N9473, N8728, N8289, N5730);
and AND3 (N9475, N9474, N3784, N672);
nand NAND4 (N9476, N9466, N4657, N2960, N3360);
nor NOR2 (N9477, N9444, N5828);
not NOT1 (N9478, N9471);
buf BUF1 (N9479, N9464);
nand NAND3 (N9480, N9477, N34, N3014);
or OR3 (N9481, N9472, N7528, N7325);
nor NOR3 (N9482, N9460, N7910, N1952);
xor XOR2 (N9483, N9463, N5034);
or OR4 (N9484, N9480, N5231, N7029, N5196);
and AND3 (N9485, N9478, N8983, N6300);
nand NAND2 (N9486, N9476, N7408);
or OR3 (N9487, N9482, N1176, N4599);
nand NAND3 (N9488, N9484, N4347, N5955);
nand NAND3 (N9489, N9488, N6079, N4474);
and AND4 (N9490, N9479, N2685, N220, N9146);
and AND2 (N9491, N9489, N761);
and AND4 (N9492, N9468, N8766, N5698, N5117);
nor NOR2 (N9493, N9481, N3610);
xor XOR2 (N9494, N9492, N834);
buf BUF1 (N9495, N9485);
buf BUF1 (N9496, N9483);
buf BUF1 (N9497, N9496);
not NOT1 (N9498, N9487);
buf BUF1 (N9499, N9495);
xor XOR2 (N9500, N9494, N7064);
xor XOR2 (N9501, N9498, N2115);
and AND4 (N9502, N9497, N3552, N8849, N8279);
and AND2 (N9503, N9499, N6545);
not NOT1 (N9504, N9475);
nand NAND2 (N9505, N9501, N2248);
xor XOR2 (N9506, N9469, N6250);
nor NOR3 (N9507, N9486, N8356, N5492);
xor XOR2 (N9508, N9503, N8890);
nor NOR4 (N9509, N9507, N4964, N2374, N8573);
nand NAND2 (N9510, N9500, N9347);
not NOT1 (N9511, N9505);
nor NOR2 (N9512, N9491, N5788);
not NOT1 (N9513, N9506);
nor NOR4 (N9514, N9504, N8386, N7035, N8190);
or OR4 (N9515, N9510, N9361, N8759, N1726);
nor NOR3 (N9516, N9493, N7492, N8084);
xor XOR2 (N9517, N9502, N6477);
nand NAND4 (N9518, N9516, N2869, N4408, N5575);
or OR2 (N9519, N9517, N6017);
buf BUF1 (N9520, N9490);
nand NAND2 (N9521, N9514, N8471);
and AND2 (N9522, N9518, N2289);
or OR3 (N9523, N9508, N5558, N2188);
or OR3 (N9524, N9520, N693, N6714);
not NOT1 (N9525, N9519);
or OR2 (N9526, N9509, N9297);
not NOT1 (N9527, N9513);
or OR4 (N9528, N9524, N5782, N7768, N2271);
not NOT1 (N9529, N9522);
not NOT1 (N9530, N9515);
nor NOR2 (N9531, N9528, N5037);
xor XOR2 (N9532, N9523, N6596);
and AND3 (N9533, N9529, N5772, N4023);
xor XOR2 (N9534, N9526, N79);
not NOT1 (N9535, N9530);
xor XOR2 (N9536, N9534, N4177);
nand NAND2 (N9537, N9511, N4412);
nand NAND2 (N9538, N9532, N4617);
buf BUF1 (N9539, N9536);
and AND4 (N9540, N9537, N2418, N107, N7103);
not NOT1 (N9541, N9531);
not NOT1 (N9542, N9525);
nor NOR3 (N9543, N9533, N2124, N4399);
nor NOR4 (N9544, N9538, N4194, N7766, N885);
and AND2 (N9545, N9543, N2120);
nor NOR3 (N9546, N9539, N5710, N659);
xor XOR2 (N9547, N9540, N4159);
xor XOR2 (N9548, N9544, N4782);
and AND2 (N9549, N9548, N3147);
buf BUF1 (N9550, N9527);
and AND2 (N9551, N9512, N9523);
buf BUF1 (N9552, N9549);
or OR4 (N9553, N9546, N5449, N8783, N1503);
nor NOR4 (N9554, N9545, N9249, N3111, N4600);
nor NOR2 (N9555, N9551, N5377);
nand NAND3 (N9556, N9550, N4204, N6452);
nand NAND3 (N9557, N9547, N6119, N6650);
or OR2 (N9558, N9521, N15);
nand NAND2 (N9559, N9557, N8592);
nor NOR4 (N9560, N9555, N1464, N7391, N3153);
nand NAND2 (N9561, N9560, N7596);
or OR2 (N9562, N9535, N8497);
buf BUF1 (N9563, N9541);
and AND2 (N9564, N9559, N873);
xor XOR2 (N9565, N9556, N448);
nor NOR3 (N9566, N9563, N8818, N8615);
nand NAND3 (N9567, N9554, N8981, N9317);
nor NOR2 (N9568, N9566, N536);
buf BUF1 (N9569, N9564);
nand NAND2 (N9570, N9552, N3049);
or OR4 (N9571, N9542, N1539, N6267, N969);
xor XOR2 (N9572, N9553, N4536);
not NOT1 (N9573, N9562);
and AND2 (N9574, N9567, N5258);
not NOT1 (N9575, N9571);
xor XOR2 (N9576, N9570, N7789);
or OR2 (N9577, N9569, N6301);
nand NAND2 (N9578, N9565, N239);
not NOT1 (N9579, N9578);
nand NAND2 (N9580, N9572, N4954);
nand NAND3 (N9581, N9576, N4801, N9207);
xor XOR2 (N9582, N9581, N9526);
not NOT1 (N9583, N9579);
buf BUF1 (N9584, N9580);
buf BUF1 (N9585, N9568);
nor NOR2 (N9586, N9577, N602);
buf BUF1 (N9587, N9561);
nand NAND2 (N9588, N9585, N3992);
nand NAND2 (N9589, N9584, N5906);
or OR4 (N9590, N9586, N5135, N4134, N1140);
not NOT1 (N9591, N9587);
not NOT1 (N9592, N9589);
buf BUF1 (N9593, N9583);
not NOT1 (N9594, N9582);
nand NAND3 (N9595, N9592, N4585, N5143);
buf BUF1 (N9596, N9595);
nand NAND2 (N9597, N9574, N1899);
and AND3 (N9598, N9558, N749, N5881);
nor NOR2 (N9599, N9597, N5135);
xor XOR2 (N9600, N9573, N6688);
buf BUF1 (N9601, N9593);
not NOT1 (N9602, N9596);
not NOT1 (N9603, N9602);
xor XOR2 (N9604, N9601, N8710);
or OR4 (N9605, N9603, N5911, N8445, N4034);
buf BUF1 (N9606, N9590);
buf BUF1 (N9607, N9604);
and AND4 (N9608, N9605, N7741, N4652, N6039);
nor NOR4 (N9609, N9598, N6880, N5433, N6170);
or OR4 (N9610, N9608, N4302, N6191, N7426);
nand NAND4 (N9611, N9609, N1751, N948, N2882);
xor XOR2 (N9612, N9600, N9452);
or OR2 (N9613, N9594, N4502);
buf BUF1 (N9614, N9613);
or OR3 (N9615, N9614, N2085, N3425);
xor XOR2 (N9616, N9588, N1482);
buf BUF1 (N9617, N9606);
not NOT1 (N9618, N9617);
and AND2 (N9619, N9607, N7173);
nor NOR2 (N9620, N9616, N3355);
buf BUF1 (N9621, N9618);
or OR3 (N9622, N9599, N293, N1821);
nor NOR3 (N9623, N9610, N5094, N7488);
nor NOR3 (N9624, N9612, N9407, N3807);
xor XOR2 (N9625, N9623, N4446);
not NOT1 (N9626, N9624);
and AND2 (N9627, N9611, N4344);
xor XOR2 (N9628, N9626, N1328);
not NOT1 (N9629, N9625);
and AND4 (N9630, N9628, N9426, N6098, N5277);
nand NAND2 (N9631, N9575, N6944);
and AND2 (N9632, N9615, N8731);
or OR3 (N9633, N9591, N6686, N6697);
and AND4 (N9634, N9620, N9512, N1131, N5316);
not NOT1 (N9635, N9633);
nand NAND2 (N9636, N9630, N9526);
nor NOR2 (N9637, N9636, N8520);
xor XOR2 (N9638, N9635, N3624);
or OR2 (N9639, N9634, N4215);
and AND4 (N9640, N9639, N5836, N6295, N1492);
buf BUF1 (N9641, N9622);
buf BUF1 (N9642, N9631);
not NOT1 (N9643, N9627);
nor NOR4 (N9644, N9638, N5655, N1521, N3817);
xor XOR2 (N9645, N9641, N4246);
not NOT1 (N9646, N9645);
nand NAND2 (N9647, N9632, N659);
not NOT1 (N9648, N9619);
not NOT1 (N9649, N9644);
or OR2 (N9650, N9647, N54);
not NOT1 (N9651, N9642);
buf BUF1 (N9652, N9649);
and AND4 (N9653, N9637, N2675, N8530, N4742);
buf BUF1 (N9654, N9621);
xor XOR2 (N9655, N9643, N3259);
and AND2 (N9656, N9654, N237);
buf BUF1 (N9657, N9653);
xor XOR2 (N9658, N9652, N2464);
xor XOR2 (N9659, N9656, N7854);
not NOT1 (N9660, N9651);
nor NOR3 (N9661, N9657, N5416, N1527);
buf BUF1 (N9662, N9655);
nand NAND2 (N9663, N9629, N212);
or OR4 (N9664, N9650, N453, N3761, N4384);
not NOT1 (N9665, N9663);
nor NOR4 (N9666, N9658, N5903, N720, N2762);
xor XOR2 (N9667, N9646, N8007);
nor NOR3 (N9668, N9664, N4363, N9336);
xor XOR2 (N9669, N9668, N4702);
nand NAND2 (N9670, N9667, N6189);
and AND3 (N9671, N9660, N4372, N7403);
xor XOR2 (N9672, N9670, N9595);
or OR3 (N9673, N9659, N952, N6610);
nand NAND4 (N9674, N9648, N24, N9510, N6971);
xor XOR2 (N9675, N9640, N5834);
and AND4 (N9676, N9665, N9066, N1525, N3293);
nand NAND3 (N9677, N9674, N3527, N60);
nor NOR4 (N9678, N9675, N4771, N3311, N7812);
nand NAND2 (N9679, N9671, N7304);
and AND3 (N9680, N9669, N5934, N6636);
and AND2 (N9681, N9672, N8117);
xor XOR2 (N9682, N9679, N8554);
nand NAND4 (N9683, N9682, N7034, N5060, N8680);
nor NOR2 (N9684, N9662, N1616);
nor NOR3 (N9685, N9677, N8261, N4778);
not NOT1 (N9686, N9661);
buf BUF1 (N9687, N9683);
not NOT1 (N9688, N9676);
or OR3 (N9689, N9684, N9552, N3462);
or OR4 (N9690, N9681, N5668, N7766, N7894);
nor NOR3 (N9691, N9678, N6722, N4469);
and AND3 (N9692, N9686, N6054, N767);
or OR4 (N9693, N9690, N1601, N5704, N866);
nand NAND3 (N9694, N9685, N164, N8797);
and AND4 (N9695, N9691, N3045, N8086, N8303);
not NOT1 (N9696, N9673);
nor NOR4 (N9697, N9688, N4822, N6878, N8480);
and AND2 (N9698, N9694, N5019);
nand NAND4 (N9699, N9698, N8555, N5214, N6884);
not NOT1 (N9700, N9692);
buf BUF1 (N9701, N9700);
nor NOR3 (N9702, N9696, N8854, N3397);
xor XOR2 (N9703, N9702, N1189);
or OR4 (N9704, N9695, N4601, N2878, N7876);
or OR4 (N9705, N9687, N8204, N7550, N8123);
and AND3 (N9706, N9680, N1026, N1187);
not NOT1 (N9707, N9666);
or OR4 (N9708, N9705, N66, N3664, N6764);
or OR2 (N9709, N9699, N3979);
xor XOR2 (N9710, N9689, N1049);
nor NOR4 (N9711, N9693, N5110, N840, N9388);
buf BUF1 (N9712, N9710);
or OR4 (N9713, N9708, N8650, N6090, N1867);
buf BUF1 (N9714, N9709);
xor XOR2 (N9715, N9706, N6432);
or OR3 (N9716, N9701, N9404, N5967);
xor XOR2 (N9717, N9715, N8842);
buf BUF1 (N9718, N9697);
nor NOR3 (N9719, N9711, N6922, N4167);
or OR4 (N9720, N9718, N1251, N5627, N4840);
xor XOR2 (N9721, N9716, N6329);
buf BUF1 (N9722, N9719);
nor NOR2 (N9723, N9704, N4317);
nand NAND2 (N9724, N9723, N5521);
or OR3 (N9725, N9721, N5312, N427);
and AND4 (N9726, N9720, N3458, N5065, N9546);
xor XOR2 (N9727, N9703, N4090);
not NOT1 (N9728, N9727);
not NOT1 (N9729, N9724);
not NOT1 (N9730, N9712);
nand NAND4 (N9731, N9730, N1266, N9356, N5054);
buf BUF1 (N9732, N9726);
and AND3 (N9733, N9707, N5620, N1676);
buf BUF1 (N9734, N9717);
buf BUF1 (N9735, N9728);
nor NOR2 (N9736, N9713, N9660);
nor NOR3 (N9737, N9729, N5223, N1964);
nor NOR4 (N9738, N9725, N4158, N4572, N1374);
xor XOR2 (N9739, N9738, N6248);
not NOT1 (N9740, N9734);
not NOT1 (N9741, N9737);
not NOT1 (N9742, N9735);
and AND3 (N9743, N9736, N2760, N2591);
buf BUF1 (N9744, N9743);
not NOT1 (N9745, N9739);
and AND3 (N9746, N9742, N9174, N5995);
not NOT1 (N9747, N9731);
nand NAND2 (N9748, N9714, N1821);
nand NAND3 (N9749, N9744, N2596, N7847);
nand NAND3 (N9750, N9740, N3576, N2402);
nand NAND2 (N9751, N9746, N8820);
or OR4 (N9752, N9732, N606, N4515, N9299);
or OR3 (N9753, N9750, N790, N897);
and AND4 (N9754, N9733, N7021, N3291, N566);
nand NAND3 (N9755, N9754, N6883, N9195);
not NOT1 (N9756, N9741);
not NOT1 (N9757, N9755);
and AND2 (N9758, N9722, N7316);
buf BUF1 (N9759, N9747);
or OR2 (N9760, N9759, N1158);
nand NAND2 (N9761, N9753, N1878);
or OR3 (N9762, N9758, N7548, N7708);
buf BUF1 (N9763, N9760);
not NOT1 (N9764, N9749);
nand NAND2 (N9765, N9745, N1174);
nor NOR2 (N9766, N9762, N8047);
nor NOR3 (N9767, N9751, N3849, N7502);
xor XOR2 (N9768, N9765, N2392);
nor NOR3 (N9769, N9761, N5601, N7847);
buf BUF1 (N9770, N9763);
buf BUF1 (N9771, N9766);
and AND3 (N9772, N9767, N7235, N8098);
nor NOR3 (N9773, N9757, N3977, N5612);
buf BUF1 (N9774, N9772);
or OR2 (N9775, N9771, N847);
or OR4 (N9776, N9752, N191, N7825, N7529);
buf BUF1 (N9777, N9774);
not NOT1 (N9778, N9756);
and AND4 (N9779, N9748, N7212, N1560, N1987);
buf BUF1 (N9780, N9778);
buf BUF1 (N9781, N9764);
not NOT1 (N9782, N9781);
or OR4 (N9783, N9773, N4266, N7883, N8883);
or OR2 (N9784, N9770, N7011);
or OR3 (N9785, N9782, N137, N7412);
or OR3 (N9786, N9779, N2144, N9242);
nor NOR3 (N9787, N9768, N7681, N7458);
nand NAND2 (N9788, N9780, N4214);
xor XOR2 (N9789, N9775, N3410);
or OR3 (N9790, N9776, N8042, N6777);
nand NAND2 (N9791, N9787, N3607);
nor NOR4 (N9792, N9785, N2747, N619, N4425);
and AND4 (N9793, N9791, N3624, N6997, N1865);
nor NOR4 (N9794, N9786, N4282, N4746, N8588);
nor NOR3 (N9795, N9794, N5861, N1839);
and AND3 (N9796, N9795, N5965, N2229);
nor NOR2 (N9797, N9769, N7377);
buf BUF1 (N9798, N9784);
not NOT1 (N9799, N9792);
or OR4 (N9800, N9793, N3670, N77, N8543);
nor NOR2 (N9801, N9798, N7685);
not NOT1 (N9802, N9783);
nand NAND4 (N9803, N9788, N5391, N2875, N3777);
nor NOR2 (N9804, N9797, N89);
buf BUF1 (N9805, N9777);
nand NAND4 (N9806, N9789, N9181, N8311, N337);
nor NOR2 (N9807, N9806, N7082);
xor XOR2 (N9808, N9801, N9456);
nor NOR4 (N9809, N9790, N5135, N4398, N4690);
and AND3 (N9810, N9807, N450, N237);
or OR4 (N9811, N9810, N6314, N9138, N7211);
or OR3 (N9812, N9802, N7577, N6721);
xor XOR2 (N9813, N9808, N7139);
nor NOR3 (N9814, N9800, N6289, N7968);
not NOT1 (N9815, N9813);
nand NAND3 (N9816, N9804, N2433, N9472);
or OR4 (N9817, N9809, N2135, N2792, N7807);
buf BUF1 (N9818, N9796);
and AND2 (N9819, N9803, N4572);
and AND2 (N9820, N9814, N1061);
xor XOR2 (N9821, N9799, N3434);
not NOT1 (N9822, N9812);
and AND2 (N9823, N9811, N6638);
or OR3 (N9824, N9819, N8413, N4183);
or OR4 (N9825, N9822, N2197, N8408, N9658);
nor NOR4 (N9826, N9824, N950, N7989, N287);
nor NOR4 (N9827, N9823, N7584, N7389, N821);
or OR4 (N9828, N9815, N2860, N5481, N1086);
or OR2 (N9829, N9805, N4531);
nor NOR2 (N9830, N9821, N4319);
not NOT1 (N9831, N9825);
nand NAND2 (N9832, N9818, N8849);
and AND2 (N9833, N9830, N8237);
not NOT1 (N9834, N9833);
xor XOR2 (N9835, N9829, N6063);
buf BUF1 (N9836, N9820);
nor NOR3 (N9837, N9828, N671, N1369);
buf BUF1 (N9838, N9832);
xor XOR2 (N9839, N9834, N3288);
not NOT1 (N9840, N9816);
and AND2 (N9841, N9826, N7730);
and AND3 (N9842, N9839, N7495, N4607);
nand NAND2 (N9843, N9841, N311);
buf BUF1 (N9844, N9840);
not NOT1 (N9845, N9843);
and AND2 (N9846, N9831, N8859);
nand NAND3 (N9847, N9838, N3331, N212);
and AND3 (N9848, N9846, N1226, N3875);
and AND4 (N9849, N9837, N3707, N1759, N7273);
or OR2 (N9850, N9848, N875);
buf BUF1 (N9851, N9842);
nor NOR2 (N9852, N9847, N7507);
or OR2 (N9853, N9850, N6642);
nand NAND2 (N9854, N9836, N8414);
or OR2 (N9855, N9854, N2933);
xor XOR2 (N9856, N9845, N3171);
xor XOR2 (N9857, N9852, N2802);
not NOT1 (N9858, N9835);
nor NOR3 (N9859, N9858, N3694, N2141);
and AND2 (N9860, N9849, N472);
xor XOR2 (N9861, N9827, N7759);
or OR2 (N9862, N9817, N4896);
xor XOR2 (N9863, N9860, N4728);
xor XOR2 (N9864, N9851, N6148);
nand NAND3 (N9865, N9859, N1417, N2195);
or OR3 (N9866, N9862, N9725, N9451);
not NOT1 (N9867, N9866);
buf BUF1 (N9868, N9855);
nor NOR3 (N9869, N9856, N9829, N947);
or OR3 (N9870, N9857, N5089, N6247);
or OR2 (N9871, N9865, N6745);
buf BUF1 (N9872, N9853);
not NOT1 (N9873, N9868);
nand NAND3 (N9874, N9864, N7880, N3194);
nor NOR4 (N9875, N9863, N7514, N4718, N5339);
nand NAND4 (N9876, N9869, N681, N1550, N8961);
and AND2 (N9877, N9874, N4568);
xor XOR2 (N9878, N9873, N5637);
or OR2 (N9879, N9872, N781);
nor NOR3 (N9880, N9844, N2754, N1897);
nor NOR3 (N9881, N9875, N9501, N1351);
not NOT1 (N9882, N9880);
not NOT1 (N9883, N9870);
or OR3 (N9884, N9883, N7609, N8575);
not NOT1 (N9885, N9878);
nor NOR2 (N9886, N9876, N1397);
not NOT1 (N9887, N9871);
xor XOR2 (N9888, N9886, N6055);
not NOT1 (N9889, N9877);
or OR2 (N9890, N9885, N9622);
buf BUF1 (N9891, N9882);
buf BUF1 (N9892, N9890);
xor XOR2 (N9893, N9887, N8077);
nand NAND3 (N9894, N9881, N8253, N3260);
or OR3 (N9895, N9888, N912, N7788);
buf BUF1 (N9896, N9879);
nand NAND3 (N9897, N9867, N8880, N4882);
and AND3 (N9898, N9861, N5947, N7755);
xor XOR2 (N9899, N9894, N6123);
buf BUF1 (N9900, N9895);
buf BUF1 (N9901, N9891);
not NOT1 (N9902, N9899);
and AND4 (N9903, N9897, N4266, N6387, N4722);
or OR3 (N9904, N9900, N6481, N9397);
nor NOR4 (N9905, N9892, N6755, N3619, N7016);
or OR2 (N9906, N9884, N326);
and AND4 (N9907, N9889, N5598, N1271, N9685);
xor XOR2 (N9908, N9901, N7416);
nand NAND2 (N9909, N9903, N2805);
and AND2 (N9910, N9907, N5021);
xor XOR2 (N9911, N9902, N1041);
or OR2 (N9912, N9906, N4856);
buf BUF1 (N9913, N9905);
xor XOR2 (N9914, N9904, N3126);
and AND3 (N9915, N9914, N9155, N335);
xor XOR2 (N9916, N9912, N5019);
xor XOR2 (N9917, N9913, N3470);
buf BUF1 (N9918, N9898);
not NOT1 (N9919, N9908);
nand NAND4 (N9920, N9896, N7933, N8540, N8281);
xor XOR2 (N9921, N9919, N430);
buf BUF1 (N9922, N9909);
not NOT1 (N9923, N9910);
nor NOR2 (N9924, N9916, N6575);
or OR3 (N9925, N9918, N4490, N6025);
nand NAND2 (N9926, N9924, N6320);
not NOT1 (N9927, N9922);
buf BUF1 (N9928, N9920);
buf BUF1 (N9929, N9917);
not NOT1 (N9930, N9921);
and AND4 (N9931, N9923, N8928, N5029, N4708);
buf BUF1 (N9932, N9925);
and AND4 (N9933, N9928, N4681, N1702, N2160);
and AND2 (N9934, N9929, N9592);
nor NOR4 (N9935, N9934, N7660, N8581, N6281);
nand NAND4 (N9936, N9932, N1696, N1683, N3197);
buf BUF1 (N9937, N9911);
nand NAND4 (N9938, N9893, N4841, N8501, N5075);
buf BUF1 (N9939, N9936);
xor XOR2 (N9940, N9930, N8400);
or OR3 (N9941, N9937, N4316, N3459);
buf BUF1 (N9942, N9939);
xor XOR2 (N9943, N9938, N1152);
buf BUF1 (N9944, N9935);
buf BUF1 (N9945, N9933);
not NOT1 (N9946, N9931);
xor XOR2 (N9947, N9941, N5240);
or OR3 (N9948, N9945, N2193, N5064);
not NOT1 (N9949, N9942);
and AND4 (N9950, N9943, N5882, N3571, N7613);
buf BUF1 (N9951, N9940);
and AND3 (N9952, N9927, N1656, N8943);
and AND4 (N9953, N9951, N2982, N2418, N9741);
nand NAND4 (N9954, N9952, N2313, N3269, N149);
nand NAND3 (N9955, N9926, N3195, N9879);
not NOT1 (N9956, N9953);
and AND3 (N9957, N9949, N8615, N8408);
xor XOR2 (N9958, N9955, N2772);
nor NOR4 (N9959, N9956, N8667, N5959, N8265);
xor XOR2 (N9960, N9958, N7709);
not NOT1 (N9961, N9950);
xor XOR2 (N9962, N9957, N3697);
nand NAND2 (N9963, N9954, N5039);
nor NOR3 (N9964, N9948, N2866, N5926);
or OR2 (N9965, N9962, N3183);
not NOT1 (N9966, N9961);
xor XOR2 (N9967, N9964, N9240);
or OR4 (N9968, N9959, N310, N8980, N7424);
buf BUF1 (N9969, N9915);
xor XOR2 (N9970, N9946, N7692);
and AND4 (N9971, N9944, N967, N203, N5132);
xor XOR2 (N9972, N9970, N8937);
not NOT1 (N9973, N9965);
nor NOR4 (N9974, N9966, N3294, N9110, N3411);
xor XOR2 (N9975, N9973, N9187);
not NOT1 (N9976, N9967);
xor XOR2 (N9977, N9974, N3055);
or OR4 (N9978, N9975, N7128, N7206, N3159);
not NOT1 (N9979, N9947);
not NOT1 (N9980, N9969);
nand NAND2 (N9981, N9960, N2714);
nand NAND2 (N9982, N9977, N2327);
and AND2 (N9983, N9971, N1124);
not NOT1 (N9984, N9981);
not NOT1 (N9985, N9982);
xor XOR2 (N9986, N9976, N6860);
xor XOR2 (N9987, N9968, N3603);
or OR3 (N9988, N9987, N3334, N6783);
nor NOR4 (N9989, N9978, N8515, N4388, N8513);
and AND2 (N9990, N9985, N7215);
nand NAND2 (N9991, N9963, N6674);
and AND3 (N9992, N9979, N2916, N1625);
nor NOR2 (N9993, N9988, N8210);
xor XOR2 (N9994, N9992, N4745);
not NOT1 (N9995, N9980);
or OR3 (N9996, N9983, N4802, N290);
buf BUF1 (N9997, N9986);
xor XOR2 (N9998, N9991, N7680);
xor XOR2 (N9999, N9996, N9798);
and AND3 (N10000, N9997, N1361, N3540);
nor NOR4 (N10001, N9993, N7010, N5437, N2570);
or OR2 (N10002, N9999, N208);
nand NAND2 (N10003, N9972, N4249);
or OR4 (N10004, N9994, N9363, N2740, N2794);
or OR2 (N10005, N10003, N2966);
buf BUF1 (N10006, N9984);
or OR2 (N10007, N10006, N3470);
nand NAND3 (N10008, N10001, N5301, N665);
xor XOR2 (N10009, N9990, N4427);
or OR3 (N10010, N10007, N1091, N3438);
xor XOR2 (N10011, N10005, N1146);
xor XOR2 (N10012, N10010, N2499);
nand NAND2 (N10013, N9998, N3732);
xor XOR2 (N10014, N9995, N3452);
nor NOR2 (N10015, N10012, N2588);
nor NOR4 (N10016, N10011, N100, N3608, N437);
or OR3 (N10017, N10002, N9272, N1137);
buf BUF1 (N10018, N10000);
or OR3 (N10019, N10004, N1005, N5115);
xor XOR2 (N10020, N10018, N6371);
nor NOR2 (N10021, N10014, N9729);
xor XOR2 (N10022, N10016, N9181);
xor XOR2 (N10023, N10013, N8987);
buf BUF1 (N10024, N10021);
or OR2 (N10025, N10020, N9279);
nor NOR4 (N10026, N10025, N2094, N6852, N7756);
not NOT1 (N10027, N10015);
not NOT1 (N10028, N10019);
nand NAND4 (N10029, N10024, N10008, N6318, N4071);
and AND2 (N10030, N5419, N8449);
nor NOR3 (N10031, N10022, N7135, N543);
not NOT1 (N10032, N9989);
nor NOR4 (N10033, N10026, N8213, N1939, N6843);
or OR4 (N10034, N10033, N1495, N4378, N3567);
and AND4 (N10035, N10030, N7902, N3877, N7921);
and AND4 (N10036, N10023, N2788, N1716, N7870);
nor NOR3 (N10037, N10031, N5769, N9060);
nand NAND4 (N10038, N10029, N273, N5313, N6281);
buf BUF1 (N10039, N10017);
nand NAND2 (N10040, N10034, N7105);
and AND2 (N10041, N10038, N2585);
and AND2 (N10042, N10036, N6067);
xor XOR2 (N10043, N10040, N4388);
buf BUF1 (N10044, N10032);
nand NAND2 (N10045, N10027, N8516);
and AND3 (N10046, N10044, N9409, N2146);
and AND3 (N10047, N10043, N6719, N9457);
not NOT1 (N10048, N10045);
not NOT1 (N10049, N10037);
xor XOR2 (N10050, N10048, N416);
buf BUF1 (N10051, N10046);
not NOT1 (N10052, N10051);
or OR3 (N10053, N10028, N2412, N18);
nor NOR3 (N10054, N10039, N1587, N7425);
not NOT1 (N10055, N10035);
nand NAND4 (N10056, N10041, N4500, N1392, N633);
not NOT1 (N10057, N10042);
not NOT1 (N10058, N10052);
xor XOR2 (N10059, N10050, N7655);
buf BUF1 (N10060, N10056);
nor NOR4 (N10061, N10009, N7595, N2342, N4959);
not NOT1 (N10062, N10061);
and AND2 (N10063, N10053, N9757);
and AND4 (N10064, N10063, N9078, N12, N9466);
nor NOR4 (N10065, N10055, N6300, N2836, N524);
nand NAND4 (N10066, N10059, N2575, N2413, N7399);
or OR3 (N10067, N10058, N626, N409);
xor XOR2 (N10068, N10049, N3338);
or OR4 (N10069, N10047, N5381, N7226, N1184);
not NOT1 (N10070, N10060);
buf BUF1 (N10071, N10067);
xor XOR2 (N10072, N10068, N982);
nor NOR4 (N10073, N10062, N5163, N9311, N1727);
or OR2 (N10074, N10069, N716);
not NOT1 (N10075, N10066);
buf BUF1 (N10076, N10073);
and AND3 (N10077, N10071, N8362, N2267);
not NOT1 (N10078, N10075);
xor XOR2 (N10079, N10074, N2124);
nor NOR3 (N10080, N10057, N7133, N3182);
nand NAND2 (N10081, N10078, N8308);
nand NAND2 (N10082, N10077, N9099);
not NOT1 (N10083, N10081);
buf BUF1 (N10084, N10076);
or OR2 (N10085, N10082, N214);
buf BUF1 (N10086, N10085);
or OR4 (N10087, N10065, N8261, N4417, N7223);
and AND2 (N10088, N10054, N5827);
not NOT1 (N10089, N10064);
or OR4 (N10090, N10089, N1026, N4881, N822);
nand NAND3 (N10091, N10090, N5329, N4972);
or OR2 (N10092, N10088, N718);
nor NOR4 (N10093, N10091, N3242, N371, N7232);
and AND2 (N10094, N10070, N7387);
nand NAND2 (N10095, N10086, N7940);
nor NOR4 (N10096, N10095, N6900, N6087, N2504);
buf BUF1 (N10097, N10072);
nand NAND3 (N10098, N10097, N8482, N3797);
and AND4 (N10099, N10098, N6999, N5875, N5435);
or OR2 (N10100, N10094, N9834);
or OR4 (N10101, N10092, N1823, N7638, N4246);
nor NOR2 (N10102, N10101, N9420);
or OR3 (N10103, N10093, N7885, N1478);
or OR3 (N10104, N10084, N4540, N3453);
nand NAND2 (N10105, N10079, N517);
buf BUF1 (N10106, N10080);
or OR3 (N10107, N10103, N2986, N3324);
not NOT1 (N10108, N10083);
not NOT1 (N10109, N10104);
buf BUF1 (N10110, N10107);
not NOT1 (N10111, N10106);
or OR2 (N10112, N10102, N9398);
and AND3 (N10113, N10108, N4323, N6585);
buf BUF1 (N10114, N10100);
xor XOR2 (N10115, N10112, N809);
buf BUF1 (N10116, N10114);
nor NOR4 (N10117, N10087, N9431, N5125, N3126);
buf BUF1 (N10118, N10113);
buf BUF1 (N10119, N10099);
nand NAND2 (N10120, N10111, N3309);
nand NAND4 (N10121, N10116, N9408, N2841, N9909);
nand NAND4 (N10122, N10120, N4484, N9616, N3102);
and AND4 (N10123, N10096, N9980, N8289, N8978);
buf BUF1 (N10124, N10122);
or OR2 (N10125, N10109, N1278);
or OR3 (N10126, N10125, N5368, N2396);
nand NAND3 (N10127, N10119, N2228, N5982);
not NOT1 (N10128, N10118);
buf BUF1 (N10129, N10127);
nor NOR3 (N10130, N10128, N7124, N5260);
not NOT1 (N10131, N10124);
nand NAND3 (N10132, N10126, N961, N3483);
or OR4 (N10133, N10105, N3189, N5481, N2581);
nand NAND2 (N10134, N10121, N4472);
buf BUF1 (N10135, N10123);
and AND2 (N10136, N10131, N7436);
not NOT1 (N10137, N10133);
or OR4 (N10138, N10115, N8247, N3389, N5370);
buf BUF1 (N10139, N10110);
nand NAND4 (N10140, N10139, N3081, N9564, N4679);
buf BUF1 (N10141, N10134);
buf BUF1 (N10142, N10130);
or OR3 (N10143, N10137, N4476, N7175);
or OR2 (N10144, N10136, N9322);
or OR4 (N10145, N10138, N3609, N6370, N6425);
not NOT1 (N10146, N10141);
xor XOR2 (N10147, N10132, N9486);
nor NOR2 (N10148, N10146, N331);
and AND2 (N10149, N10147, N689);
xor XOR2 (N10150, N10145, N3437);
buf BUF1 (N10151, N10149);
xor XOR2 (N10152, N10150, N778);
and AND2 (N10153, N10148, N3056);
nor NOR2 (N10154, N10140, N3369);
not NOT1 (N10155, N10129);
and AND2 (N10156, N10144, N6960);
or OR3 (N10157, N10154, N9841, N3209);
buf BUF1 (N10158, N10117);
nor NOR4 (N10159, N10153, N906, N9287, N7695);
nor NOR3 (N10160, N10143, N8108, N2089);
nand NAND4 (N10161, N10156, N5240, N2711, N9474);
and AND2 (N10162, N10155, N7389);
and AND4 (N10163, N10158, N4430, N2345, N5896);
nor NOR4 (N10164, N10151, N6639, N6937, N3991);
xor XOR2 (N10165, N10164, N5505);
and AND3 (N10166, N10159, N7662, N5978);
nand NAND2 (N10167, N10160, N7402);
nand NAND2 (N10168, N10142, N1603);
nor NOR4 (N10169, N10135, N7764, N5597, N2647);
nor NOR4 (N10170, N10163, N3815, N1765, N4944);
or OR4 (N10171, N10166, N5224, N4231, N5910);
nand NAND3 (N10172, N10170, N1610, N1765);
buf BUF1 (N10173, N10161);
not NOT1 (N10174, N10171);
and AND2 (N10175, N10165, N2697);
nand NAND4 (N10176, N10174, N5113, N8489, N10112);
buf BUF1 (N10177, N10157);
nand NAND2 (N10178, N10175, N3308);
and AND4 (N10179, N10169, N5096, N9379, N1583);
not NOT1 (N10180, N10178);
or OR4 (N10181, N10179, N5440, N9775, N3192);
nand NAND3 (N10182, N10152, N2284, N7940);
or OR4 (N10183, N10182, N2264, N5122, N4223);
nand NAND4 (N10184, N10162, N827, N653, N4978);
nand NAND4 (N10185, N10181, N215, N4476, N1102);
or OR4 (N10186, N10177, N4296, N4047, N584);
nand NAND2 (N10187, N10184, N4325);
buf BUF1 (N10188, N10167);
and AND2 (N10189, N10180, N3343);
nor NOR2 (N10190, N10188, N7768);
nand NAND4 (N10191, N10185, N7183, N9183, N7879);
or OR4 (N10192, N10190, N3036, N4597, N8656);
nor NOR3 (N10193, N10183, N7942, N5303);
and AND2 (N10194, N10189, N5968);
nor NOR4 (N10195, N10186, N557, N3791, N715);
nor NOR4 (N10196, N10194, N9013, N3889, N3905);
not NOT1 (N10197, N10195);
or OR3 (N10198, N10172, N6326, N3803);
xor XOR2 (N10199, N10196, N709);
and AND4 (N10200, N10187, N1289, N5862, N2830);
buf BUF1 (N10201, N10168);
buf BUF1 (N10202, N10198);
nand NAND3 (N10203, N10173, N2710, N7869);
nand NAND2 (N10204, N10193, N8904);
buf BUF1 (N10205, N10199);
or OR4 (N10206, N10176, N6103, N6548, N10030);
xor XOR2 (N10207, N10191, N1930);
and AND2 (N10208, N10200, N4294);
nor NOR3 (N10209, N10203, N5958, N4463);
xor XOR2 (N10210, N10201, N27);
nor NOR2 (N10211, N10208, N3705);
nor NOR4 (N10212, N10204, N6933, N9958, N6018);
not NOT1 (N10213, N10197);
buf BUF1 (N10214, N10206);
not NOT1 (N10215, N10213);
nand NAND4 (N10216, N10202, N633, N3852, N6964);
buf BUF1 (N10217, N10214);
buf BUF1 (N10218, N10212);
buf BUF1 (N10219, N10205);
and AND4 (N10220, N10210, N6005, N8029, N6675);
and AND2 (N10221, N10215, N1603);
buf BUF1 (N10222, N10220);
buf BUF1 (N10223, N10222);
buf BUF1 (N10224, N10192);
or OR4 (N10225, N10223, N1659, N8916, N2653);
or OR4 (N10226, N10207, N5616, N2261, N10088);
not NOT1 (N10227, N10219);
nand NAND4 (N10228, N10217, N8523, N723, N7137);
nand NAND3 (N10229, N10228, N4164, N2558);
not NOT1 (N10230, N10211);
buf BUF1 (N10231, N10218);
and AND3 (N10232, N10230, N1673, N6734);
xor XOR2 (N10233, N10224, N9370);
or OR4 (N10234, N10209, N7577, N745, N383);
or OR3 (N10235, N10227, N9361, N2765);
xor XOR2 (N10236, N10234, N937);
nor NOR2 (N10237, N10226, N3638);
xor XOR2 (N10238, N10221, N1853);
xor XOR2 (N10239, N10216, N3217);
not NOT1 (N10240, N10225);
buf BUF1 (N10241, N10236);
nor NOR2 (N10242, N10241, N2191);
buf BUF1 (N10243, N10229);
nand NAND4 (N10244, N10242, N8081, N7288, N2347);
not NOT1 (N10245, N10233);
nand NAND4 (N10246, N10231, N2859, N23, N5547);
and AND3 (N10247, N10240, N10190, N7141);
not NOT1 (N10248, N10244);
nand NAND4 (N10249, N10239, N166, N6788, N4727);
xor XOR2 (N10250, N10237, N10016);
nor NOR4 (N10251, N10238, N7672, N9998, N2836);
not NOT1 (N10252, N10245);
buf BUF1 (N10253, N10249);
and AND4 (N10254, N10251, N7345, N4359, N9910);
not NOT1 (N10255, N10232);
not NOT1 (N10256, N10247);
nor NOR3 (N10257, N10254, N5215, N4164);
buf BUF1 (N10258, N10235);
buf BUF1 (N10259, N10250);
not NOT1 (N10260, N10252);
and AND4 (N10261, N10248, N6925, N351, N479);
nor NOR3 (N10262, N10255, N5728, N1205);
buf BUF1 (N10263, N10261);
not NOT1 (N10264, N10243);
nand NAND2 (N10265, N10256, N1661);
not NOT1 (N10266, N10259);
not NOT1 (N10267, N10265);
nand NAND2 (N10268, N10267, N8238);
not NOT1 (N10269, N10246);
buf BUF1 (N10270, N10263);
or OR4 (N10271, N10253, N395, N9129, N6737);
xor XOR2 (N10272, N10266, N3413);
nor NOR3 (N10273, N10268, N2070, N8626);
nor NOR4 (N10274, N10264, N8150, N4799, N4443);
xor XOR2 (N10275, N10271, N1760);
nand NAND4 (N10276, N10272, N8816, N259, N7602);
or OR2 (N10277, N10260, N2488);
or OR4 (N10278, N10262, N4634, N6713, N7799);
nand NAND3 (N10279, N10277, N5231, N4139);
or OR4 (N10280, N10276, N7014, N7123, N98);
and AND3 (N10281, N10270, N8415, N2821);
not NOT1 (N10282, N10281);
xor XOR2 (N10283, N10274, N5360);
and AND4 (N10284, N10278, N992, N8967, N2443);
not NOT1 (N10285, N10269);
xor XOR2 (N10286, N10285, N1561);
xor XOR2 (N10287, N10280, N4716);
xor XOR2 (N10288, N10283, N3479);
not NOT1 (N10289, N10273);
not NOT1 (N10290, N10279);
nor NOR2 (N10291, N10282, N7419);
and AND4 (N10292, N10291, N1248, N5652, N953);
and AND4 (N10293, N10257, N853, N9313, N5831);
nor NOR4 (N10294, N10292, N7531, N6118, N3147);
not NOT1 (N10295, N10290);
and AND4 (N10296, N10295, N9768, N2007, N9218);
not NOT1 (N10297, N10293);
not NOT1 (N10298, N10286);
or OR2 (N10299, N10258, N9735);
nand NAND2 (N10300, N10294, N5775);
and AND3 (N10301, N10300, N3762, N1020);
or OR4 (N10302, N10288, N3024, N49, N3289);
and AND2 (N10303, N10284, N8292);
buf BUF1 (N10304, N10287);
or OR3 (N10305, N10275, N6009, N2859);
nand NAND2 (N10306, N10303, N4540);
or OR3 (N10307, N10305, N9973, N4793);
not NOT1 (N10308, N10296);
buf BUF1 (N10309, N10304);
not NOT1 (N10310, N10307);
or OR2 (N10311, N10306, N4819);
buf BUF1 (N10312, N10310);
nand NAND4 (N10313, N10309, N3069, N5329, N3209);
and AND4 (N10314, N10299, N7541, N3193, N3998);
and AND4 (N10315, N10298, N8251, N4673, N7978);
xor XOR2 (N10316, N10312, N1222);
and AND3 (N10317, N10289, N6038, N273);
nor NOR2 (N10318, N10313, N2810);
and AND3 (N10319, N10315, N2995, N4666);
buf BUF1 (N10320, N10301);
buf BUF1 (N10321, N10318);
xor XOR2 (N10322, N10314, N1391);
xor XOR2 (N10323, N10308, N1912);
nor NOR2 (N10324, N10297, N3133);
and AND2 (N10325, N10302, N563);
xor XOR2 (N10326, N10320, N234);
xor XOR2 (N10327, N10323, N1780);
not NOT1 (N10328, N10326);
nand NAND3 (N10329, N10319, N2066, N6039);
or OR4 (N10330, N10324, N29, N457, N6805);
buf BUF1 (N10331, N10330);
and AND2 (N10332, N10325, N8803);
and AND4 (N10333, N10327, N5922, N10094, N1450);
buf BUF1 (N10334, N10321);
xor XOR2 (N10335, N10316, N6026);
xor XOR2 (N10336, N10322, N9479);
and AND2 (N10337, N10336, N3881);
buf BUF1 (N10338, N10328);
and AND3 (N10339, N10311, N5189, N3685);
buf BUF1 (N10340, N10317);
nand NAND3 (N10341, N10331, N7800, N10102);
and AND3 (N10342, N10329, N8705, N441);
and AND3 (N10343, N10341, N4096, N7876);
nand NAND4 (N10344, N10334, N1415, N3147, N6677);
not NOT1 (N10345, N10338);
nor NOR2 (N10346, N10343, N8797);
or OR4 (N10347, N10332, N1202, N8956, N9333);
nand NAND4 (N10348, N10333, N2382, N9471, N10000);
not NOT1 (N10349, N10335);
xor XOR2 (N10350, N10346, N2629);
not NOT1 (N10351, N10339);
nand NAND4 (N10352, N10351, N2764, N5617, N749);
not NOT1 (N10353, N10349);
xor XOR2 (N10354, N10350, N9997);
xor XOR2 (N10355, N10347, N7911);
nand NAND3 (N10356, N10340, N5525, N10073);
or OR4 (N10357, N10353, N7662, N3119, N4560);
not NOT1 (N10358, N10344);
nor NOR3 (N10359, N10352, N7937, N9596);
not NOT1 (N10360, N10359);
xor XOR2 (N10361, N10358, N6256);
nor NOR4 (N10362, N10342, N5747, N8250, N493);
xor XOR2 (N10363, N10362, N3546);
nor NOR4 (N10364, N10356, N10117, N9420, N2331);
buf BUF1 (N10365, N10361);
not NOT1 (N10366, N10355);
xor XOR2 (N10367, N10364, N3623);
or OR4 (N10368, N10365, N4435, N3793, N6117);
or OR2 (N10369, N10366, N7204);
or OR3 (N10370, N10357, N8208, N118);
nand NAND2 (N10371, N10360, N5438);
or OR3 (N10372, N10368, N5004, N10188);
and AND4 (N10373, N10337, N2711, N6101, N611);
xor XOR2 (N10374, N10345, N2600);
nor NOR4 (N10375, N10371, N5908, N7543, N2190);
nor NOR2 (N10376, N10367, N9513);
xor XOR2 (N10377, N10370, N10068);
not NOT1 (N10378, N10373);
not NOT1 (N10379, N10348);
not NOT1 (N10380, N10379);
buf BUF1 (N10381, N10378);
nand NAND2 (N10382, N10372, N9333);
nor NOR4 (N10383, N10375, N2562, N3897, N836);
xor XOR2 (N10384, N10377, N2454);
nor NOR2 (N10385, N10369, N2734);
or OR3 (N10386, N10363, N2480, N10062);
nand NAND4 (N10387, N10374, N1392, N6605, N4257);
nand NAND2 (N10388, N10387, N2290);
not NOT1 (N10389, N10383);
buf BUF1 (N10390, N10388);
nor NOR4 (N10391, N10382, N6366, N3235, N7896);
xor XOR2 (N10392, N10381, N552);
buf BUF1 (N10393, N10389);
nor NOR2 (N10394, N10384, N9523);
nor NOR2 (N10395, N10380, N2945);
nand NAND2 (N10396, N10394, N7741);
xor XOR2 (N10397, N10386, N6880);
buf BUF1 (N10398, N10391);
nand NAND3 (N10399, N10398, N7804, N9021);
and AND4 (N10400, N10397, N3363, N2660, N3403);
nand NAND4 (N10401, N10393, N4207, N3669, N9516);
nand NAND2 (N10402, N10395, N9540);
buf BUF1 (N10403, N10354);
buf BUF1 (N10404, N10396);
nor NOR2 (N10405, N10402, N2995);
not NOT1 (N10406, N10399);
nand NAND2 (N10407, N10401, N7936);
nand NAND4 (N10408, N10376, N6844, N9938, N47);
xor XOR2 (N10409, N10390, N2609);
not NOT1 (N10410, N10404);
or OR2 (N10411, N10405, N9364);
not NOT1 (N10412, N10392);
nand NAND2 (N10413, N10409, N3539);
buf BUF1 (N10414, N10408);
or OR2 (N10415, N10403, N6933);
not NOT1 (N10416, N10407);
or OR2 (N10417, N10414, N3824);
buf BUF1 (N10418, N10417);
nand NAND3 (N10419, N10413, N8751, N9854);
or OR4 (N10420, N10418, N7440, N6776, N7502);
and AND3 (N10421, N10406, N2693, N6378);
buf BUF1 (N10422, N10419);
nand NAND4 (N10423, N10410, N4519, N3057, N6181);
xor XOR2 (N10424, N10411, N5897);
not NOT1 (N10425, N10420);
xor XOR2 (N10426, N10423, N8775);
buf BUF1 (N10427, N10426);
nand NAND2 (N10428, N10422, N7556);
nor NOR2 (N10429, N10385, N5102);
nand NAND2 (N10430, N10424, N6009);
nor NOR4 (N10431, N10430, N5363, N7282, N9395);
nor NOR2 (N10432, N10416, N5815);
or OR4 (N10433, N10415, N5111, N4568, N7811);
not NOT1 (N10434, N10431);
not NOT1 (N10435, N10433);
xor XOR2 (N10436, N10427, N4052);
and AND4 (N10437, N10421, N8369, N8744, N3815);
buf BUF1 (N10438, N10412);
nand NAND4 (N10439, N10432, N1077, N155, N9914);
and AND2 (N10440, N10436, N9640);
not NOT1 (N10441, N10439);
nand NAND2 (N10442, N10425, N4067);
or OR3 (N10443, N10442, N4460, N9547);
and AND3 (N10444, N10438, N8131, N7569);
xor XOR2 (N10445, N10441, N7716);
not NOT1 (N10446, N10440);
xor XOR2 (N10447, N10400, N5311);
nand NAND4 (N10448, N10447, N3460, N4163, N2647);
not NOT1 (N10449, N10444);
not NOT1 (N10450, N10449);
not NOT1 (N10451, N10434);
or OR4 (N10452, N10428, N9270, N5726, N10093);
nand NAND2 (N10453, N10429, N4265);
buf BUF1 (N10454, N10445);
or OR3 (N10455, N10435, N6828, N7283);
not NOT1 (N10456, N10437);
xor XOR2 (N10457, N10456, N10034);
not NOT1 (N10458, N10451);
and AND2 (N10459, N10458, N2273);
and AND2 (N10460, N10450, N4674);
nor NOR3 (N10461, N10443, N1009, N6935);
nor NOR4 (N10462, N10455, N1632, N10424, N7195);
and AND4 (N10463, N10460, N4551, N7755, N6439);
buf BUF1 (N10464, N10457);
not NOT1 (N10465, N10454);
nor NOR3 (N10466, N10459, N1035, N4234);
and AND2 (N10467, N10463, N6157);
and AND3 (N10468, N10464, N2935, N9599);
xor XOR2 (N10469, N10465, N772);
nand NAND2 (N10470, N10452, N3530);
buf BUF1 (N10471, N10461);
nor NOR4 (N10472, N10471, N10309, N88, N7323);
nand NAND4 (N10473, N10472, N1670, N7114, N2914);
not NOT1 (N10474, N10467);
not NOT1 (N10475, N10453);
and AND3 (N10476, N10446, N2379, N9422);
nor NOR2 (N10477, N10475, N10461);
not NOT1 (N10478, N10470);
nor NOR2 (N10479, N10477, N3026);
and AND3 (N10480, N10448, N865, N2509);
nand NAND4 (N10481, N10480, N7278, N8280, N7999);
not NOT1 (N10482, N10479);
not NOT1 (N10483, N10466);
not NOT1 (N10484, N10483);
nor NOR3 (N10485, N10482, N2199, N4969);
not NOT1 (N10486, N10481);
nand NAND3 (N10487, N10484, N6588, N2742);
or OR4 (N10488, N10462, N6773, N6749, N2502);
nand NAND4 (N10489, N10476, N8052, N974, N10301);
or OR4 (N10490, N10486, N8053, N46, N1148);
or OR2 (N10491, N10487, N4680);
buf BUF1 (N10492, N10491);
nand NAND4 (N10493, N10469, N4398, N1407, N6136);
nand NAND4 (N10494, N10485, N8571, N2113, N3790);
or OR3 (N10495, N10473, N3169, N9477);
or OR3 (N10496, N10494, N8209, N7722);
xor XOR2 (N10497, N10490, N7602);
buf BUF1 (N10498, N10474);
nand NAND4 (N10499, N10488, N575, N9693, N6153);
nand NAND3 (N10500, N10493, N10114, N9531);
xor XOR2 (N10501, N10489, N10472);
nor NOR2 (N10502, N10497, N6705);
not NOT1 (N10503, N10496);
or OR3 (N10504, N10502, N7564, N8475);
not NOT1 (N10505, N10503);
buf BUF1 (N10506, N10501);
buf BUF1 (N10507, N10498);
or OR3 (N10508, N10504, N1660, N379);
nor NOR2 (N10509, N10508, N10321);
and AND2 (N10510, N10505, N1545);
and AND2 (N10511, N10492, N9613);
and AND3 (N10512, N10499, N4674, N6088);
and AND3 (N10513, N10468, N2964, N4880);
nor NOR2 (N10514, N10500, N1018);
nand NAND2 (N10515, N10506, N8757);
xor XOR2 (N10516, N10514, N1019);
xor XOR2 (N10517, N10478, N8267);
nor NOR2 (N10518, N10515, N5581);
or OR2 (N10519, N10517, N5857);
and AND2 (N10520, N10513, N5977);
and AND2 (N10521, N10510, N9610);
xor XOR2 (N10522, N10511, N9886);
or OR3 (N10523, N10512, N1324, N6810);
or OR4 (N10524, N10507, N8773, N1745, N9085);
buf BUF1 (N10525, N10524);
or OR2 (N10526, N10522, N5150);
and AND3 (N10527, N10525, N2506, N4784);
buf BUF1 (N10528, N10526);
not NOT1 (N10529, N10521);
and AND2 (N10530, N10509, N9928);
not NOT1 (N10531, N10530);
buf BUF1 (N10532, N10531);
nor NOR3 (N10533, N10529, N1315, N1471);
or OR4 (N10534, N10528, N5716, N8068, N4773);
xor XOR2 (N10535, N10516, N5596);
xor XOR2 (N10536, N10527, N9158);
or OR3 (N10537, N10520, N4033, N3174);
nor NOR4 (N10538, N10518, N6603, N6305, N8198);
nand NAND2 (N10539, N10532, N8371);
or OR3 (N10540, N10539, N3043, N180);
nor NOR3 (N10541, N10535, N5234, N8703);
xor XOR2 (N10542, N10540, N7529);
buf BUF1 (N10543, N10534);
not NOT1 (N10544, N10523);
buf BUF1 (N10545, N10495);
nand NAND3 (N10546, N10537, N9808, N6505);
not NOT1 (N10547, N10538);
buf BUF1 (N10548, N10542);
not NOT1 (N10549, N10541);
not NOT1 (N10550, N10519);
buf BUF1 (N10551, N10546);
and AND4 (N10552, N10543, N2619, N2318, N879);
nand NAND3 (N10553, N10533, N1658, N7791);
not NOT1 (N10554, N10536);
xor XOR2 (N10555, N10544, N910);
buf BUF1 (N10556, N10547);
nand NAND2 (N10557, N10556, N9695);
buf BUF1 (N10558, N10550);
xor XOR2 (N10559, N10552, N5437);
buf BUF1 (N10560, N10554);
and AND3 (N10561, N10549, N5628, N1037);
nor NOR2 (N10562, N10548, N3115);
and AND4 (N10563, N10559, N8511, N177, N5801);
xor XOR2 (N10564, N10553, N9981);
nor NOR2 (N10565, N10562, N6161);
xor XOR2 (N10566, N10557, N2638);
nand NAND3 (N10567, N10563, N4838, N744);
not NOT1 (N10568, N10561);
buf BUF1 (N10569, N10567);
or OR3 (N10570, N10565, N632, N8081);
nor NOR2 (N10571, N10566, N8369);
nor NOR4 (N10572, N10551, N9909, N1124, N10153);
xor XOR2 (N10573, N10560, N3117);
nand NAND4 (N10574, N10568, N3426, N8346, N1221);
nand NAND4 (N10575, N10572, N2912, N10295, N4752);
xor XOR2 (N10576, N10555, N3163);
not NOT1 (N10577, N10558);
not NOT1 (N10578, N10564);
buf BUF1 (N10579, N10578);
xor XOR2 (N10580, N10569, N5966);
xor XOR2 (N10581, N10574, N3927);
buf BUF1 (N10582, N10575);
xor XOR2 (N10583, N10579, N7023);
not NOT1 (N10584, N10576);
xor XOR2 (N10585, N10545, N9098);
nor NOR4 (N10586, N10570, N5542, N1787, N10215);
buf BUF1 (N10587, N10580);
xor XOR2 (N10588, N10586, N1387);
nand NAND3 (N10589, N10582, N9071, N9413);
xor XOR2 (N10590, N10585, N4415);
and AND3 (N10591, N10590, N1513, N9744);
nor NOR4 (N10592, N10583, N8519, N5586, N2814);
and AND3 (N10593, N10587, N9394, N3952);
buf BUF1 (N10594, N10588);
buf BUF1 (N10595, N10591);
or OR3 (N10596, N10592, N4323, N10060);
and AND3 (N10597, N10571, N5487, N7287);
and AND4 (N10598, N10594, N6284, N7271, N243);
nor NOR2 (N10599, N10577, N5584);
nor NOR4 (N10600, N10595, N29, N856, N8707);
or OR4 (N10601, N10581, N7247, N3891, N4327);
xor XOR2 (N10602, N10599, N3070);
nor NOR3 (N10603, N10584, N8115, N8258);
nor NOR4 (N10604, N10601, N2630, N10491, N791);
xor XOR2 (N10605, N10600, N8867);
not NOT1 (N10606, N10602);
xor XOR2 (N10607, N10596, N3881);
not NOT1 (N10608, N10606);
and AND2 (N10609, N10573, N2494);
and AND3 (N10610, N10609, N5366, N9192);
nand NAND3 (N10611, N10603, N5138, N2709);
nand NAND2 (N10612, N10598, N6356);
or OR2 (N10613, N10597, N2071);
xor XOR2 (N10614, N10605, N2778);
and AND4 (N10615, N10610, N2034, N2192, N6410);
nor NOR3 (N10616, N10611, N9781, N9290);
or OR3 (N10617, N10614, N9653, N10604);
buf BUF1 (N10618, N4435);
nor NOR3 (N10619, N10617, N10237, N7257);
nand NAND3 (N10620, N10607, N4293, N6115);
xor XOR2 (N10621, N10615, N7685);
not NOT1 (N10622, N10621);
and AND3 (N10623, N10589, N1094, N6779);
or OR2 (N10624, N10620, N9946);
nor NOR3 (N10625, N10616, N8440, N10511);
and AND2 (N10626, N10622, N1416);
buf BUF1 (N10627, N10623);
nor NOR2 (N10628, N10593, N7887);
nor NOR2 (N10629, N10627, N7556);
nor NOR3 (N10630, N10619, N10178, N6976);
nor NOR3 (N10631, N10628, N10256, N3208);
nor NOR2 (N10632, N10626, N656);
nand NAND4 (N10633, N10630, N9744, N1356, N10536);
xor XOR2 (N10634, N10608, N4696);
nand NAND2 (N10635, N10633, N8653);
buf BUF1 (N10636, N10631);
buf BUF1 (N10637, N10634);
xor XOR2 (N10638, N10612, N230);
nand NAND4 (N10639, N10629, N2460, N8887, N1801);
or OR4 (N10640, N10632, N2651, N3329, N3537);
buf BUF1 (N10641, N10624);
and AND2 (N10642, N10639, N8764);
not NOT1 (N10643, N10638);
and AND2 (N10644, N10637, N9520);
and AND4 (N10645, N10613, N9294, N250, N9768);
nor NOR3 (N10646, N10642, N1694, N3020);
or OR3 (N10647, N10644, N7218, N1770);
buf BUF1 (N10648, N10643);
buf BUF1 (N10649, N10625);
nor NOR3 (N10650, N10649, N2691, N2922);
nor NOR2 (N10651, N10635, N6758);
and AND4 (N10652, N10646, N8071, N326, N8627);
or OR3 (N10653, N10636, N5883, N6017);
and AND4 (N10654, N10645, N5649, N1430, N3266);
buf BUF1 (N10655, N10641);
buf BUF1 (N10656, N10653);
not NOT1 (N10657, N10640);
and AND4 (N10658, N10647, N1152, N9987, N6122);
not NOT1 (N10659, N10655);
nor NOR2 (N10660, N10618, N4676);
buf BUF1 (N10661, N10660);
nor NOR4 (N10662, N10656, N1225, N6425, N5360);
buf BUF1 (N10663, N10657);
or OR2 (N10664, N10651, N3179);
nor NOR4 (N10665, N10662, N8752, N6753, N5965);
and AND3 (N10666, N10648, N5982, N3761);
and AND4 (N10667, N10650, N2052, N4398, N3607);
and AND2 (N10668, N10664, N458);
nand NAND3 (N10669, N10666, N4342, N8800);
xor XOR2 (N10670, N10663, N6627);
not NOT1 (N10671, N10668);
or OR2 (N10672, N10665, N9190);
nor NOR4 (N10673, N10661, N6644, N9078, N533);
not NOT1 (N10674, N10671);
nand NAND3 (N10675, N10654, N6134, N10459);
buf BUF1 (N10676, N10675);
buf BUF1 (N10677, N10673);
xor XOR2 (N10678, N10670, N2489);
or OR3 (N10679, N10658, N9481, N7335);
and AND3 (N10680, N10659, N8555, N3329);
buf BUF1 (N10681, N10667);
xor XOR2 (N10682, N10679, N7607);
and AND3 (N10683, N10677, N5122, N10028);
nand NAND4 (N10684, N10669, N7488, N10181, N3963);
or OR2 (N10685, N10680, N554);
or OR3 (N10686, N10678, N8915, N2361);
and AND2 (N10687, N10674, N5957);
not NOT1 (N10688, N10687);
or OR3 (N10689, N10688, N6128, N583);
nor NOR3 (N10690, N10681, N4183, N7301);
xor XOR2 (N10691, N10676, N5107);
xor XOR2 (N10692, N10689, N3561);
buf BUF1 (N10693, N10685);
xor XOR2 (N10694, N10692, N791);
buf BUF1 (N10695, N10683);
or OR3 (N10696, N10693, N2177, N3665);
nand NAND3 (N10697, N10686, N9523, N2044);
nor NOR2 (N10698, N10652, N3208);
buf BUF1 (N10699, N10682);
nor NOR2 (N10700, N10697, N9289);
nand NAND4 (N10701, N10684, N3922, N6736, N3781);
buf BUF1 (N10702, N10672);
not NOT1 (N10703, N10696);
or OR4 (N10704, N10691, N5784, N10298, N6240);
not NOT1 (N10705, N10699);
nand NAND4 (N10706, N10694, N7186, N4451, N8402);
or OR2 (N10707, N10705, N2465);
nor NOR2 (N10708, N10703, N8977);
buf BUF1 (N10709, N10701);
xor XOR2 (N10710, N10709, N6314);
buf BUF1 (N10711, N10708);
xor XOR2 (N10712, N10706, N2993);
nor NOR3 (N10713, N10711, N9118, N614);
xor XOR2 (N10714, N10690, N5377);
not NOT1 (N10715, N10700);
xor XOR2 (N10716, N10713, N3962);
or OR3 (N10717, N10714, N6312, N9269);
xor XOR2 (N10718, N10715, N9734);
not NOT1 (N10719, N10716);
buf BUF1 (N10720, N10707);
xor XOR2 (N10721, N10718, N8562);
buf BUF1 (N10722, N10698);
not NOT1 (N10723, N10719);
or OR2 (N10724, N10710, N10091);
nor NOR2 (N10725, N10712, N2234);
buf BUF1 (N10726, N10717);
and AND4 (N10727, N10720, N8099, N8770, N2402);
and AND4 (N10728, N10702, N8368, N3618, N6348);
or OR2 (N10729, N10722, N4234);
nor NOR4 (N10730, N10729, N5367, N10620, N5078);
not NOT1 (N10731, N10724);
nor NOR2 (N10732, N10721, N7124);
nor NOR4 (N10733, N10730, N9805, N7300, N5743);
nor NOR2 (N10734, N10695, N10560);
and AND2 (N10735, N10733, N2478);
nand NAND2 (N10736, N10704, N875);
not NOT1 (N10737, N10725);
or OR2 (N10738, N10723, N4606);
and AND2 (N10739, N10734, N4606);
or OR3 (N10740, N10731, N3535, N717);
xor XOR2 (N10741, N10739, N3730);
xor XOR2 (N10742, N10740, N5379);
or OR2 (N10743, N10736, N2201);
xor XOR2 (N10744, N10728, N5072);
or OR3 (N10745, N10738, N9572, N2393);
or OR4 (N10746, N10737, N1154, N1618, N3180);
nor NOR4 (N10747, N10745, N2992, N9165, N5272);
or OR2 (N10748, N10744, N6954);
and AND2 (N10749, N10746, N8940);
buf BUF1 (N10750, N10732);
nand NAND2 (N10751, N10727, N9572);
and AND4 (N10752, N10742, N1827, N4811, N664);
and AND2 (N10753, N10741, N8121);
xor XOR2 (N10754, N10726, N8228);
and AND3 (N10755, N10743, N2761, N6891);
buf BUF1 (N10756, N10747);
not NOT1 (N10757, N10754);
nor NOR4 (N10758, N10735, N5560, N2287, N6996);
or OR3 (N10759, N10752, N5224, N5674);
nor NOR3 (N10760, N10750, N2830, N9324);
xor XOR2 (N10761, N10758, N1294);
buf BUF1 (N10762, N10753);
nand NAND4 (N10763, N10761, N1123, N5902, N3802);
or OR3 (N10764, N10748, N1355, N9990);
or OR2 (N10765, N10755, N10280);
xor XOR2 (N10766, N10756, N7035);
nand NAND4 (N10767, N10765, N7249, N1506, N6031);
buf BUF1 (N10768, N10767);
nand NAND3 (N10769, N10751, N9843, N2224);
or OR4 (N10770, N10768, N3337, N7507, N3669);
nand NAND3 (N10771, N10757, N7431, N3674);
nand NAND4 (N10772, N10763, N1521, N8151, N3895);
and AND3 (N10773, N10771, N1030, N5146);
or OR2 (N10774, N10766, N4591);
or OR4 (N10775, N10759, N6298, N3117, N9014);
buf BUF1 (N10776, N10769);
or OR3 (N10777, N10762, N6238, N1736);
and AND4 (N10778, N10775, N5304, N9773, N7033);
not NOT1 (N10779, N10772);
nor NOR2 (N10780, N10770, N8363);
buf BUF1 (N10781, N10773);
nand NAND3 (N10782, N10774, N8850, N5183);
xor XOR2 (N10783, N10777, N4680);
xor XOR2 (N10784, N10781, N2613);
xor XOR2 (N10785, N10749, N2292);
buf BUF1 (N10786, N10785);
or OR2 (N10787, N10764, N7991);
xor XOR2 (N10788, N10782, N6338);
xor XOR2 (N10789, N10787, N9062);
or OR2 (N10790, N10784, N3241);
or OR4 (N10791, N10790, N8324, N4680, N8319);
not NOT1 (N10792, N10791);
nor NOR4 (N10793, N10760, N6073, N5347, N10521);
or OR2 (N10794, N10778, N8144);
not NOT1 (N10795, N10788);
and AND2 (N10796, N10783, N4815);
or OR2 (N10797, N10796, N7799);
xor XOR2 (N10798, N10779, N8489);
nor NOR2 (N10799, N10798, N2952);
xor XOR2 (N10800, N10780, N4288);
not NOT1 (N10801, N10789);
not NOT1 (N10802, N10792);
nand NAND4 (N10803, N10786, N6225, N4590, N4275);
xor XOR2 (N10804, N10795, N525);
nand NAND3 (N10805, N10776, N2694, N3307);
nor NOR4 (N10806, N10801, N8033, N2626, N6792);
or OR4 (N10807, N10803, N1104, N5933, N9704);
buf BUF1 (N10808, N10807);
or OR2 (N10809, N10806, N2440);
nand NAND4 (N10810, N10799, N5039, N7611, N4317);
not NOT1 (N10811, N10805);
not NOT1 (N10812, N10811);
nor NOR4 (N10813, N10808, N1091, N10233, N4669);
not NOT1 (N10814, N10793);
buf BUF1 (N10815, N10809);
and AND2 (N10816, N10814, N4999);
or OR2 (N10817, N10797, N174);
xor XOR2 (N10818, N10794, N6829);
not NOT1 (N10819, N10804);
or OR2 (N10820, N10818, N9239);
nor NOR4 (N10821, N10815, N10027, N10130, N8251);
or OR3 (N10822, N10813, N2050, N53);
nor NOR3 (N10823, N10822, N5209, N557);
buf BUF1 (N10824, N10802);
nor NOR4 (N10825, N10820, N8233, N3126, N4186);
not NOT1 (N10826, N10817);
or OR2 (N10827, N10812, N1483);
nand NAND2 (N10828, N10800, N938);
buf BUF1 (N10829, N10810);
xor XOR2 (N10830, N10816, N5680);
nor NOR4 (N10831, N10824, N5511, N689, N6727);
buf BUF1 (N10832, N10826);
nor NOR2 (N10833, N10830, N1668);
and AND2 (N10834, N10825, N5239);
not NOT1 (N10835, N10821);
xor XOR2 (N10836, N10823, N7479);
xor XOR2 (N10837, N10835, N9502);
nor NOR3 (N10838, N10837, N5621, N3717);
nor NOR3 (N10839, N10819, N611, N9810);
nand NAND4 (N10840, N10838, N725, N7919, N2697);
xor XOR2 (N10841, N10834, N2698);
or OR2 (N10842, N10840, N4680);
nor NOR3 (N10843, N10842, N4988, N5974);
xor XOR2 (N10844, N10836, N7719);
xor XOR2 (N10845, N10832, N3906);
xor XOR2 (N10846, N10845, N1520);
and AND4 (N10847, N10831, N2245, N995, N7815);
nor NOR3 (N10848, N10846, N8961, N4162);
xor XOR2 (N10849, N10827, N2428);
not NOT1 (N10850, N10829);
or OR2 (N10851, N10849, N1046);
or OR4 (N10852, N10847, N5203, N10421, N9827);
buf BUF1 (N10853, N10852);
buf BUF1 (N10854, N10848);
xor XOR2 (N10855, N10853, N10159);
xor XOR2 (N10856, N10854, N10397);
buf BUF1 (N10857, N10851);
nand NAND3 (N10858, N10828, N10570, N10071);
nand NAND3 (N10859, N10841, N2033, N1065);
nor NOR2 (N10860, N10833, N9021);
buf BUF1 (N10861, N10860);
or OR2 (N10862, N10857, N149);
or OR2 (N10863, N10856, N720);
not NOT1 (N10864, N10844);
nand NAND3 (N10865, N10864, N10123, N8521);
nor NOR2 (N10866, N10861, N2573);
xor XOR2 (N10867, N10859, N3225);
not NOT1 (N10868, N10855);
not NOT1 (N10869, N10866);
nor NOR4 (N10870, N10843, N4213, N5047, N9072);
nor NOR4 (N10871, N10870, N6594, N3813, N9297);
nor NOR2 (N10872, N10863, N10780);
nand NAND2 (N10873, N10839, N3892);
nand NAND2 (N10874, N10862, N4910);
and AND2 (N10875, N10872, N5570);
nor NOR4 (N10876, N10867, N4047, N632, N8887);
buf BUF1 (N10877, N10858);
or OR4 (N10878, N10877, N577, N5667, N1055);
xor XOR2 (N10879, N10850, N4881);
nand NAND3 (N10880, N10871, N5025, N1689);
or OR2 (N10881, N10865, N10217);
nor NOR4 (N10882, N10878, N10115, N7697, N7108);
or OR4 (N10883, N10873, N6352, N1892, N3389);
nand NAND3 (N10884, N10876, N2966, N2397);
or OR2 (N10885, N10881, N8010);
not NOT1 (N10886, N10875);
nor NOR3 (N10887, N10882, N6048, N2020);
xor XOR2 (N10888, N10885, N8035);
buf BUF1 (N10889, N10879);
nor NOR2 (N10890, N10888, N1533);
or OR4 (N10891, N10880, N622, N6994, N9714);
buf BUF1 (N10892, N10868);
buf BUF1 (N10893, N10883);
and AND2 (N10894, N10892, N7118);
nand NAND4 (N10895, N10890, N66, N10678, N8604);
not NOT1 (N10896, N10894);
and AND4 (N10897, N10869, N6162, N10256, N9846);
nor NOR4 (N10898, N10874, N9346, N2072, N3180);
and AND3 (N10899, N10884, N10624, N6063);
nor NOR3 (N10900, N10887, N10587, N6329);
nand NAND2 (N10901, N10895, N1582);
not NOT1 (N10902, N10889);
nor NOR3 (N10903, N10893, N9319, N647);
buf BUF1 (N10904, N10899);
or OR4 (N10905, N10891, N875, N1756, N9336);
not NOT1 (N10906, N10900);
xor XOR2 (N10907, N10898, N6251);
buf BUF1 (N10908, N10906);
not NOT1 (N10909, N10907);
buf BUF1 (N10910, N10904);
or OR2 (N10911, N10909, N3803);
nand NAND3 (N10912, N10897, N4774, N4644);
buf BUF1 (N10913, N10911);
xor XOR2 (N10914, N10913, N8892);
or OR3 (N10915, N10910, N2828, N8128);
or OR4 (N10916, N10903, N5357, N8390, N575);
buf BUF1 (N10917, N10901);
and AND2 (N10918, N10916, N8689);
xor XOR2 (N10919, N10912, N5186);
nor NOR3 (N10920, N10917, N9021, N606);
buf BUF1 (N10921, N10918);
or OR4 (N10922, N10902, N6816, N1439, N7398);
nand NAND4 (N10923, N10886, N6513, N620, N2812);
xor XOR2 (N10924, N10922, N884);
nor NOR2 (N10925, N10914, N3200);
not NOT1 (N10926, N10921);
not NOT1 (N10927, N10915);
not NOT1 (N10928, N10923);
and AND3 (N10929, N10920, N75, N6028);
not NOT1 (N10930, N10928);
or OR2 (N10931, N10905, N7074);
buf BUF1 (N10932, N10896);
xor XOR2 (N10933, N10927, N10120);
not NOT1 (N10934, N10919);
buf BUF1 (N10935, N10924);
or OR3 (N10936, N10932, N3409, N3574);
not NOT1 (N10937, N10908);
nor NOR3 (N10938, N10926, N1463, N1636);
xor XOR2 (N10939, N10936, N7123);
buf BUF1 (N10940, N10931);
not NOT1 (N10941, N10930);
nor NOR2 (N10942, N10925, N4412);
xor XOR2 (N10943, N10937, N8295);
buf BUF1 (N10944, N10934);
or OR3 (N10945, N10941, N9334, N7379);
and AND3 (N10946, N10939, N163, N4169);
and AND4 (N10947, N10938, N8013, N1000, N7575);
or OR3 (N10948, N10944, N3923, N4368);
not NOT1 (N10949, N10946);
or OR2 (N10950, N10929, N4780);
not NOT1 (N10951, N10943);
nand NAND4 (N10952, N10940, N6025, N8315, N8631);
or OR4 (N10953, N10950, N5812, N4352, N7311);
or OR4 (N10954, N10952, N4945, N10839, N5514);
or OR2 (N10955, N10942, N5734);
or OR3 (N10956, N10935, N6102, N4208);
not NOT1 (N10957, N10953);
nor NOR2 (N10958, N10957, N2185);
and AND2 (N10959, N10933, N9213);
xor XOR2 (N10960, N10956, N8449);
nor NOR3 (N10961, N10951, N4677, N5856);
and AND3 (N10962, N10961, N7965, N6761);
nor NOR2 (N10963, N10958, N4925);
or OR4 (N10964, N10945, N9477, N10464, N8210);
or OR2 (N10965, N10959, N6771);
or OR3 (N10966, N10949, N172, N2936);
or OR3 (N10967, N10960, N4372, N3573);
xor XOR2 (N10968, N10955, N3544);
or OR3 (N10969, N10954, N8963, N2304);
or OR2 (N10970, N10963, N455);
buf BUF1 (N10971, N10970);
and AND2 (N10972, N10969, N10101);
not NOT1 (N10973, N10966);
nor NOR4 (N10974, N10971, N3146, N8810, N3085);
buf BUF1 (N10975, N10972);
and AND4 (N10976, N10968, N6388, N10576, N4937);
nand NAND4 (N10977, N10967, N10088, N3989, N8163);
buf BUF1 (N10978, N10948);
nor NOR3 (N10979, N10976, N2028, N7681);
buf BUF1 (N10980, N10979);
and AND4 (N10981, N10964, N1288, N10057, N354);
and AND3 (N10982, N10980, N6728, N9837);
nand NAND4 (N10983, N10974, N5845, N6375, N710);
or OR2 (N10984, N10947, N7263);
buf BUF1 (N10985, N10977);
nand NAND2 (N10986, N10982, N2938);
buf BUF1 (N10987, N10965);
nand NAND4 (N10988, N10987, N852, N573, N5930);
not NOT1 (N10989, N10962);
buf BUF1 (N10990, N10973);
or OR4 (N10991, N10989, N4252, N3862, N2864);
or OR2 (N10992, N10988, N3917);
or OR2 (N10993, N10981, N3396);
buf BUF1 (N10994, N10978);
or OR2 (N10995, N10975, N10410);
nand NAND3 (N10996, N10995, N10042, N3058);
and AND2 (N10997, N10992, N3721);
nand NAND4 (N10998, N10996, N3091, N6839, N3382);
or OR2 (N10999, N10990, N878);
not NOT1 (N11000, N10986);
nand NAND4 (N11001, N10991, N2600, N1055, N8345);
buf BUF1 (N11002, N11000);
buf BUF1 (N11003, N10984);
and AND4 (N11004, N10994, N7327, N4105, N4398);
not NOT1 (N11005, N10985);
nand NAND4 (N11006, N11003, N2771, N10271, N9670);
nor NOR3 (N11007, N11004, N3516, N8608);
and AND4 (N11008, N10998, N8308, N7757, N9755);
xor XOR2 (N11009, N10999, N9574);
or OR2 (N11010, N11002, N3823);
buf BUF1 (N11011, N10993);
or OR3 (N11012, N11010, N2654, N5537);
and AND3 (N11013, N11012, N9746, N3542);
xor XOR2 (N11014, N10997, N1266);
nand NAND4 (N11015, N11006, N513, N685, N8771);
buf BUF1 (N11016, N11001);
buf BUF1 (N11017, N11005);
buf BUF1 (N11018, N11009);
buf BUF1 (N11019, N11013);
xor XOR2 (N11020, N11016, N7277);
nand NAND3 (N11021, N11008, N1730, N8172);
not NOT1 (N11022, N11015);
nand NAND3 (N11023, N11021, N3765, N10714);
buf BUF1 (N11024, N11020);
not NOT1 (N11025, N11022);
or OR3 (N11026, N11018, N967, N7682);
buf BUF1 (N11027, N11025);
buf BUF1 (N11028, N11014);
and AND4 (N11029, N11028, N5598, N2693, N1107);
nand NAND3 (N11030, N11029, N6515, N6544);
xor XOR2 (N11031, N11023, N9359);
or OR4 (N11032, N11007, N3566, N3705, N8336);
or OR2 (N11033, N11030, N5961);
xor XOR2 (N11034, N11017, N9962);
or OR2 (N11035, N11034, N10820);
nor NOR3 (N11036, N11035, N562, N3357);
buf BUF1 (N11037, N11011);
xor XOR2 (N11038, N11027, N8780);
not NOT1 (N11039, N11036);
xor XOR2 (N11040, N11033, N118);
not NOT1 (N11041, N11026);
buf BUF1 (N11042, N11019);
and AND3 (N11043, N11032, N4131, N9330);
xor XOR2 (N11044, N11031, N5866);
and AND2 (N11045, N11039, N6742);
nor NOR4 (N11046, N11038, N1107, N9052, N3342);
xor XOR2 (N11047, N11024, N10944);
or OR3 (N11048, N11046, N1189, N3773);
xor XOR2 (N11049, N11037, N2814);
nand NAND2 (N11050, N11040, N9459);
buf BUF1 (N11051, N11049);
buf BUF1 (N11052, N11050);
nand NAND2 (N11053, N11051, N5651);
nand NAND4 (N11054, N11043, N6603, N2092, N8896);
nor NOR4 (N11055, N11053, N10499, N1504, N5980);
xor XOR2 (N11056, N11052, N635);
or OR3 (N11057, N11047, N3209, N5971);
not NOT1 (N11058, N11044);
not NOT1 (N11059, N11056);
and AND3 (N11060, N11048, N9088, N842);
not NOT1 (N11061, N11060);
nand NAND3 (N11062, N11041, N297, N1644);
xor XOR2 (N11063, N11061, N2115);
and AND4 (N11064, N11055, N3247, N3077, N7493);
buf BUF1 (N11065, N11058);
or OR4 (N11066, N11065, N8939, N3998, N10966);
nor NOR2 (N11067, N11059, N3149);
or OR4 (N11068, N11054, N4691, N7864, N7975);
nand NAND2 (N11069, N11067, N10302);
or OR4 (N11070, N11063, N3842, N10459, N10540);
or OR3 (N11071, N10983, N567, N5511);
or OR2 (N11072, N11042, N9261);
buf BUF1 (N11073, N11069);
and AND3 (N11074, N11066, N139, N5655);
or OR4 (N11075, N11045, N8305, N8880, N994);
not NOT1 (N11076, N11062);
nand NAND3 (N11077, N11070, N8583, N1029);
not NOT1 (N11078, N11071);
or OR2 (N11079, N11073, N4531);
nand NAND4 (N11080, N11068, N1272, N6329, N2279);
nor NOR2 (N11081, N11077, N4809);
nand NAND2 (N11082, N11078, N8028);
not NOT1 (N11083, N11075);
nor NOR2 (N11084, N11080, N9651);
or OR2 (N11085, N11076, N5226);
xor XOR2 (N11086, N11072, N8945);
nand NAND4 (N11087, N11081, N1816, N1446, N6725);
buf BUF1 (N11088, N11074);
or OR2 (N11089, N11086, N5173);
or OR3 (N11090, N11082, N378, N5042);
buf BUF1 (N11091, N11087);
buf BUF1 (N11092, N11084);
and AND2 (N11093, N11088, N4528);
xor XOR2 (N11094, N11057, N885);
nor NOR2 (N11095, N11083, N6417);
and AND3 (N11096, N11064, N7864, N2449);
nand NAND2 (N11097, N11093, N6555);
not NOT1 (N11098, N11092);
nand NAND3 (N11099, N11097, N8431, N4024);
nor NOR4 (N11100, N11089, N9576, N553, N922);
xor XOR2 (N11101, N11090, N1237);
xor XOR2 (N11102, N11085, N9225);
buf BUF1 (N11103, N11096);
nand NAND4 (N11104, N11099, N10232, N901, N10123);
buf BUF1 (N11105, N11104);
nand NAND3 (N11106, N11094, N7510, N1060);
nand NAND2 (N11107, N11103, N2635);
xor XOR2 (N11108, N11105, N10669);
nor NOR2 (N11109, N11108, N400);
nand NAND2 (N11110, N11098, N6157);
nand NAND2 (N11111, N11100, N2315);
buf BUF1 (N11112, N11095);
nor NOR4 (N11113, N11110, N7355, N8224, N1286);
xor XOR2 (N11114, N11101, N6417);
not NOT1 (N11115, N11106);
buf BUF1 (N11116, N11114);
xor XOR2 (N11117, N11079, N4010);
xor XOR2 (N11118, N11115, N9208);
nor NOR4 (N11119, N11109, N1932, N287, N1130);
nor NOR3 (N11120, N11091, N956, N8901);
not NOT1 (N11121, N11102);
or OR2 (N11122, N11117, N574);
and AND3 (N11123, N11122, N1661, N6946);
nor NOR3 (N11124, N11121, N637, N5461);
buf BUF1 (N11125, N11118);
and AND2 (N11126, N11123, N9586);
and AND2 (N11127, N11107, N10586);
nand NAND4 (N11128, N11127, N2134, N3998, N4307);
and AND3 (N11129, N11112, N3815, N1523);
not NOT1 (N11130, N11119);
or OR3 (N11131, N11125, N7064, N9044);
xor XOR2 (N11132, N11124, N5935);
buf BUF1 (N11133, N11128);
nor NOR4 (N11134, N11130, N4836, N10104, N5368);
nor NOR4 (N11135, N11126, N6084, N5470, N2630);
buf BUF1 (N11136, N11134);
nand NAND2 (N11137, N11132, N7416);
buf BUF1 (N11138, N11129);
or OR3 (N11139, N11131, N10292, N10421);
or OR4 (N11140, N11116, N141, N2730, N3100);
nor NOR3 (N11141, N11136, N2351, N8117);
buf BUF1 (N11142, N11137);
buf BUF1 (N11143, N11139);
buf BUF1 (N11144, N11143);
nor NOR3 (N11145, N11120, N2462, N2363);
buf BUF1 (N11146, N11142);
xor XOR2 (N11147, N11138, N4624);
xor XOR2 (N11148, N11141, N4815);
nand NAND4 (N11149, N11144, N117, N3278, N3012);
xor XOR2 (N11150, N11148, N10114);
not NOT1 (N11151, N11133);
buf BUF1 (N11152, N11146);
nor NOR4 (N11153, N11152, N324, N2650, N752);
nand NAND4 (N11154, N11145, N5669, N1680, N4246);
buf BUF1 (N11155, N11154);
not NOT1 (N11156, N11150);
buf BUF1 (N11157, N11151);
xor XOR2 (N11158, N11140, N2059);
and AND4 (N11159, N11156, N2288, N6163, N4632);
nand NAND3 (N11160, N11113, N10379, N9785);
buf BUF1 (N11161, N11157);
nor NOR2 (N11162, N11149, N4970);
buf BUF1 (N11163, N11158);
nand NAND2 (N11164, N11111, N5146);
or OR3 (N11165, N11163, N10950, N6634);
xor XOR2 (N11166, N11159, N9530);
nor NOR4 (N11167, N11153, N10497, N327, N163);
nor NOR4 (N11168, N11135, N4567, N4183, N9806);
xor XOR2 (N11169, N11168, N4981);
and AND2 (N11170, N11160, N2288);
xor XOR2 (N11171, N11165, N2228);
nand NAND4 (N11172, N11170, N6457, N10152, N8710);
nand NAND2 (N11173, N11171, N8611);
and AND2 (N11174, N11164, N7147);
nand NAND3 (N11175, N11147, N5022, N3547);
buf BUF1 (N11176, N11169);
nand NAND3 (N11177, N11155, N2934, N7591);
nand NAND4 (N11178, N11167, N7117, N6130, N225);
or OR2 (N11179, N11161, N9979);
nand NAND4 (N11180, N11176, N1311, N821, N2079);
nand NAND2 (N11181, N11175, N458);
or OR4 (N11182, N11172, N687, N8199, N595);
nor NOR4 (N11183, N11179, N10564, N4339, N7931);
buf BUF1 (N11184, N11174);
or OR4 (N11185, N11182, N5540, N710, N5987);
xor XOR2 (N11186, N11173, N6903);
nor NOR4 (N11187, N11181, N4030, N2630, N727);
buf BUF1 (N11188, N11178);
or OR3 (N11189, N11177, N10743, N7559);
not NOT1 (N11190, N11187);
and AND3 (N11191, N11186, N7001, N10184);
nor NOR3 (N11192, N11190, N5479, N11065);
and AND3 (N11193, N11189, N5567, N6154);
not NOT1 (N11194, N11162);
or OR4 (N11195, N11180, N8750, N53, N3071);
buf BUF1 (N11196, N11188);
or OR4 (N11197, N11192, N8509, N2968, N4550);
and AND3 (N11198, N11196, N4614, N9013);
nor NOR3 (N11199, N11166, N5824, N1690);
nor NOR4 (N11200, N11194, N5239, N10128, N690);
nor NOR4 (N11201, N11199, N6183, N2050, N5955);
or OR4 (N11202, N11185, N1908, N6610, N4377);
nor NOR4 (N11203, N11201, N10579, N7329, N6105);
and AND4 (N11204, N11202, N9906, N865, N7297);
buf BUF1 (N11205, N11200);
nand NAND2 (N11206, N11197, N10938);
xor XOR2 (N11207, N11193, N5558);
nor NOR2 (N11208, N11184, N6508);
or OR2 (N11209, N11195, N9678);
and AND4 (N11210, N11183, N10077, N11106, N7535);
not NOT1 (N11211, N11203);
nand NAND4 (N11212, N11198, N1079, N2228, N930);
or OR4 (N11213, N11205, N1937, N2197, N510);
nand NAND2 (N11214, N11204, N10480);
or OR4 (N11215, N11208, N6331, N6989, N8683);
or OR2 (N11216, N11215, N8518);
nor NOR2 (N11217, N11210, N7656);
and AND3 (N11218, N11191, N6982, N9425);
nand NAND3 (N11219, N11206, N5951, N1367);
nor NOR2 (N11220, N11213, N1685);
not NOT1 (N11221, N11209);
or OR2 (N11222, N11219, N4615);
not NOT1 (N11223, N11211);
or OR2 (N11224, N11220, N3830);
buf BUF1 (N11225, N11214);
nand NAND2 (N11226, N11218, N2303);
or OR4 (N11227, N11222, N5894, N10795, N5862);
nor NOR2 (N11228, N11226, N2123);
buf BUF1 (N11229, N11228);
nor NOR2 (N11230, N11217, N8359);
or OR2 (N11231, N11225, N2692);
and AND2 (N11232, N11212, N713);
not NOT1 (N11233, N11227);
or OR4 (N11234, N11229, N6430, N10795, N5744);
nor NOR3 (N11235, N11233, N9543, N819);
or OR3 (N11236, N11232, N1432, N5564);
xor XOR2 (N11237, N11221, N8212);
and AND2 (N11238, N11224, N6398);
nor NOR2 (N11239, N11216, N946);
buf BUF1 (N11240, N11223);
xor XOR2 (N11241, N11236, N2538);
not NOT1 (N11242, N11231);
or OR4 (N11243, N11230, N7969, N10407, N8557);
buf BUF1 (N11244, N11241);
nor NOR4 (N11245, N11235, N1756, N6660, N937);
nor NOR3 (N11246, N11237, N7234, N10505);
nor NOR3 (N11247, N11207, N7974, N8503);
buf BUF1 (N11248, N11238);
not NOT1 (N11249, N11234);
xor XOR2 (N11250, N11244, N10808);
nand NAND3 (N11251, N11248, N5914, N6134);
xor XOR2 (N11252, N11249, N9623);
and AND4 (N11253, N11242, N6552, N996, N8912);
xor XOR2 (N11254, N11246, N11074);
buf BUF1 (N11255, N11247);
or OR2 (N11256, N11251, N4122);
nand NAND2 (N11257, N11240, N9243);
or OR3 (N11258, N11257, N8909, N8267);
nor NOR2 (N11259, N11253, N2574);
not NOT1 (N11260, N11245);
not NOT1 (N11261, N11260);
nor NOR4 (N11262, N11255, N11176, N5586, N4753);
nor NOR4 (N11263, N11258, N5256, N1736, N803);
nand NAND2 (N11264, N11243, N7401);
or OR2 (N11265, N11261, N5664);
xor XOR2 (N11266, N11250, N1925);
xor XOR2 (N11267, N11264, N4215);
nand NAND3 (N11268, N11254, N7635, N2168);
nand NAND2 (N11269, N11265, N10559);
or OR2 (N11270, N11259, N10271);
not NOT1 (N11271, N11252);
not NOT1 (N11272, N11239);
xor XOR2 (N11273, N11268, N9114);
nor NOR3 (N11274, N11271, N6681, N502);
nor NOR2 (N11275, N11273, N744);
buf BUF1 (N11276, N11272);
xor XOR2 (N11277, N11266, N3222);
or OR3 (N11278, N11277, N5014, N8747);
and AND2 (N11279, N11267, N8888);
not NOT1 (N11280, N11274);
xor XOR2 (N11281, N11269, N11038);
not NOT1 (N11282, N11262);
xor XOR2 (N11283, N11282, N4476);
and AND3 (N11284, N11278, N1770, N1361);
or OR2 (N11285, N11279, N3886);
or OR4 (N11286, N11281, N10890, N3784, N6150);
not NOT1 (N11287, N11284);
not NOT1 (N11288, N11263);
and AND4 (N11289, N11280, N5611, N229, N7307);
not NOT1 (N11290, N11275);
nand NAND4 (N11291, N11285, N10542, N4510, N1845);
xor XOR2 (N11292, N11291, N4920);
or OR3 (N11293, N11290, N9078, N2284);
xor XOR2 (N11294, N11289, N9827);
or OR2 (N11295, N11293, N9101);
and AND3 (N11296, N11283, N9973, N3038);
nor NOR4 (N11297, N11292, N5561, N8896, N1702);
or OR4 (N11298, N11286, N3330, N2874, N4954);
xor XOR2 (N11299, N11294, N3631);
nor NOR4 (N11300, N11297, N9929, N10997, N9801);
nor NOR2 (N11301, N11295, N5260);
not NOT1 (N11302, N11270);
nand NAND3 (N11303, N11302, N3942, N5006);
xor XOR2 (N11304, N11298, N5940);
nor NOR4 (N11305, N11299, N9277, N10899, N3683);
not NOT1 (N11306, N11276);
xor XOR2 (N11307, N11300, N7159);
not NOT1 (N11308, N11296);
nand NAND2 (N11309, N11301, N2895);
nor NOR4 (N11310, N11288, N322, N7560, N1484);
or OR4 (N11311, N11304, N2228, N5108, N5524);
and AND3 (N11312, N11303, N2668, N5988);
not NOT1 (N11313, N11287);
xor XOR2 (N11314, N11305, N5769);
nand NAND3 (N11315, N11309, N5596, N2054);
nand NAND2 (N11316, N11310, N6967);
and AND2 (N11317, N11314, N3066);
or OR4 (N11318, N11315, N8944, N2193, N1040);
buf BUF1 (N11319, N11317);
nor NOR4 (N11320, N11307, N9482, N4483, N3916);
xor XOR2 (N11321, N11318, N4858);
not NOT1 (N11322, N11311);
nor NOR4 (N11323, N11319, N8070, N1588, N1335);
and AND2 (N11324, N11323, N7183);
nand NAND2 (N11325, N11308, N2391);
and AND4 (N11326, N11322, N8686, N11239, N6544);
or OR3 (N11327, N11321, N2235, N11232);
xor XOR2 (N11328, N11256, N3701);
not NOT1 (N11329, N11326);
nand NAND3 (N11330, N11328, N9013, N6312);
buf BUF1 (N11331, N11313);
buf BUF1 (N11332, N11324);
buf BUF1 (N11333, N11330);
nand NAND3 (N11334, N11325, N5541, N9510);
nand NAND4 (N11335, N11306, N698, N252, N11221);
xor XOR2 (N11336, N11327, N1756);
nand NAND2 (N11337, N11332, N7412);
and AND3 (N11338, N11336, N7955, N10691);
buf BUF1 (N11339, N11312);
or OR4 (N11340, N11339, N4667, N3306, N4640);
or OR2 (N11341, N11333, N9990);
xor XOR2 (N11342, N11335, N10589);
xor XOR2 (N11343, N11331, N4735);
xor XOR2 (N11344, N11329, N2894);
nor NOR3 (N11345, N11343, N155, N2065);
not NOT1 (N11346, N11344);
nand NAND3 (N11347, N11345, N4827, N3190);
xor XOR2 (N11348, N11340, N613);
not NOT1 (N11349, N11341);
nor NOR4 (N11350, N11342, N9247, N6166, N10543);
or OR4 (N11351, N11337, N11204, N1545, N751);
nor NOR2 (N11352, N11334, N690);
nor NOR2 (N11353, N11338, N6352);
not NOT1 (N11354, N11320);
nor NOR4 (N11355, N11351, N1340, N3339, N3966);
and AND4 (N11356, N11349, N10186, N4658, N6612);
xor XOR2 (N11357, N11355, N8835);
nor NOR3 (N11358, N11356, N5523, N864);
not NOT1 (N11359, N11346);
buf BUF1 (N11360, N11348);
buf BUF1 (N11361, N11347);
xor XOR2 (N11362, N11354, N8432);
nand NAND2 (N11363, N11316, N2298);
not NOT1 (N11364, N11360);
buf BUF1 (N11365, N11361);
xor XOR2 (N11366, N11363, N5136);
and AND2 (N11367, N11365, N6208);
not NOT1 (N11368, N11366);
buf BUF1 (N11369, N11368);
not NOT1 (N11370, N11362);
buf BUF1 (N11371, N11350);
and AND2 (N11372, N11358, N10771);
xor XOR2 (N11373, N11359, N3914);
not NOT1 (N11374, N11373);
or OR4 (N11375, N11367, N9833, N5304, N2189);
buf BUF1 (N11376, N11370);
not NOT1 (N11377, N11372);
and AND3 (N11378, N11352, N10908, N4889);
buf BUF1 (N11379, N11374);
buf BUF1 (N11380, N11353);
nor NOR4 (N11381, N11376, N7366, N7930, N6616);
buf BUF1 (N11382, N11379);
nand NAND2 (N11383, N11378, N11008);
or OR3 (N11384, N11381, N4277, N3488);
nand NAND2 (N11385, N11357, N963);
or OR2 (N11386, N11384, N7962);
not NOT1 (N11387, N11369);
not NOT1 (N11388, N11383);
nand NAND4 (N11389, N11388, N3912, N11197, N2858);
not NOT1 (N11390, N11364);
xor XOR2 (N11391, N11387, N5876);
and AND2 (N11392, N11385, N8848);
not NOT1 (N11393, N11390);
xor XOR2 (N11394, N11393, N7684);
not NOT1 (N11395, N11389);
nor NOR4 (N11396, N11382, N711, N9627, N4660);
nand NAND3 (N11397, N11392, N10468, N1199);
xor XOR2 (N11398, N11377, N10038);
nor NOR2 (N11399, N11398, N5586);
not NOT1 (N11400, N11375);
or OR3 (N11401, N11397, N34, N2714);
nand NAND4 (N11402, N11399, N10503, N6653, N2886);
buf BUF1 (N11403, N11391);
or OR2 (N11404, N11395, N501);
or OR2 (N11405, N11404, N2598);
nand NAND3 (N11406, N11402, N1411, N6147);
nand NAND2 (N11407, N11380, N2073);
not NOT1 (N11408, N11371);
or OR2 (N11409, N11400, N6571);
and AND3 (N11410, N11394, N7950, N10154);
nor NOR3 (N11411, N11386, N8126, N9824);
nor NOR3 (N11412, N11396, N7905, N10836);
buf BUF1 (N11413, N11408);
nor NOR2 (N11414, N11401, N5852);
not NOT1 (N11415, N11406);
and AND2 (N11416, N11407, N2695);
and AND4 (N11417, N11414, N9138, N4201, N5905);
buf BUF1 (N11418, N11412);
not NOT1 (N11419, N11418);
nand NAND3 (N11420, N11415, N900, N7985);
nand NAND2 (N11421, N11409, N6731);
nand NAND3 (N11422, N11416, N10894, N6460);
nand NAND2 (N11423, N11420, N11353);
and AND2 (N11424, N11422, N133);
nand NAND4 (N11425, N11421, N4511, N8719, N4261);
xor XOR2 (N11426, N11417, N10779);
and AND3 (N11427, N11405, N9816, N5517);
and AND2 (N11428, N11425, N10581);
xor XOR2 (N11429, N11403, N11044);
and AND4 (N11430, N11424, N4751, N7320, N7822);
or OR3 (N11431, N11411, N1022, N8998);
nand NAND4 (N11432, N11419, N7741, N9908, N3404);
or OR4 (N11433, N11413, N847, N6607, N8810);
or OR2 (N11434, N11410, N9419);
buf BUF1 (N11435, N11431);
xor XOR2 (N11436, N11435, N9531);
xor XOR2 (N11437, N11433, N3237);
xor XOR2 (N11438, N11427, N10952);
or OR3 (N11439, N11436, N9154, N3192);
or OR4 (N11440, N11438, N852, N9615, N4581);
nand NAND2 (N11441, N11430, N5529);
buf BUF1 (N11442, N11437);
nor NOR4 (N11443, N11432, N10797, N3847, N2236);
and AND2 (N11444, N11434, N3868);
nor NOR4 (N11445, N11442, N3588, N3617, N534);
xor XOR2 (N11446, N11439, N6768);
nor NOR3 (N11447, N11446, N3883, N7471);
and AND4 (N11448, N11429, N6159, N1770, N8516);
nand NAND2 (N11449, N11441, N4301);
buf BUF1 (N11450, N11448);
xor XOR2 (N11451, N11444, N7438);
not NOT1 (N11452, N11445);
not NOT1 (N11453, N11423);
not NOT1 (N11454, N11443);
xor XOR2 (N11455, N11440, N4292);
xor XOR2 (N11456, N11452, N1554);
buf BUF1 (N11457, N11428);
nand NAND3 (N11458, N11456, N4087, N4640);
buf BUF1 (N11459, N11447);
xor XOR2 (N11460, N11459, N8314);
not NOT1 (N11461, N11451);
or OR2 (N11462, N11458, N3830);
buf BUF1 (N11463, N11450);
or OR2 (N11464, N11454, N6392);
buf BUF1 (N11465, N11453);
or OR3 (N11466, N11463, N6522, N7570);
or OR2 (N11467, N11466, N7584);
not NOT1 (N11468, N11426);
nor NOR4 (N11469, N11457, N1899, N5220, N1951);
nand NAND4 (N11470, N11462, N8404, N6792, N9153);
buf BUF1 (N11471, N11449);
nand NAND2 (N11472, N11468, N8985);
and AND4 (N11473, N11465, N7707, N8571, N6856);
nor NOR4 (N11474, N11472, N9406, N242, N3893);
nor NOR3 (N11475, N11473, N5938, N7081);
nor NOR2 (N11476, N11464, N6264);
nand NAND2 (N11477, N11474, N36);
xor XOR2 (N11478, N11475, N4695);
and AND4 (N11479, N11476, N8595, N3158, N3088);
and AND4 (N11480, N11461, N11223, N5384, N5503);
not NOT1 (N11481, N11480);
nor NOR3 (N11482, N11460, N9258, N7095);
or OR2 (N11483, N11477, N4628);
xor XOR2 (N11484, N11482, N4701);
not NOT1 (N11485, N11484);
nor NOR2 (N11486, N11469, N2627);
nor NOR4 (N11487, N11470, N8360, N8964, N10077);
buf BUF1 (N11488, N11487);
nor NOR3 (N11489, N11488, N8803, N5875);
not NOT1 (N11490, N11483);
buf BUF1 (N11491, N11467);
and AND4 (N11492, N11489, N4318, N5427, N3580);
buf BUF1 (N11493, N11481);
xor XOR2 (N11494, N11485, N2148);
and AND2 (N11495, N11455, N10420);
nand NAND3 (N11496, N11492, N5753, N2987);
buf BUF1 (N11497, N11496);
nor NOR3 (N11498, N11495, N3810, N10517);
not NOT1 (N11499, N11497);
nor NOR2 (N11500, N11478, N8995);
xor XOR2 (N11501, N11498, N9119);
buf BUF1 (N11502, N11479);
xor XOR2 (N11503, N11493, N8640);
nor NOR4 (N11504, N11502, N9503, N9071, N11134);
xor XOR2 (N11505, N11490, N136);
nand NAND4 (N11506, N11491, N4353, N10058, N10674);
and AND4 (N11507, N11471, N1754, N10961, N3049);
not NOT1 (N11508, N11505);
nand NAND2 (N11509, N11501, N5756);
buf BUF1 (N11510, N11503);
nand NAND3 (N11511, N11504, N4063, N3096);
xor XOR2 (N11512, N11510, N4399);
nand NAND3 (N11513, N11500, N4548, N2140);
not NOT1 (N11514, N11512);
or OR2 (N11515, N11509, N4580);
nor NOR2 (N11516, N11513, N11068);
not NOT1 (N11517, N11507);
xor XOR2 (N11518, N11506, N8316);
and AND3 (N11519, N11514, N10255, N759);
buf BUF1 (N11520, N11519);
nor NOR4 (N11521, N11511, N6491, N4488, N2772);
and AND4 (N11522, N11515, N10588, N5812, N734);
buf BUF1 (N11523, N11517);
and AND2 (N11524, N11523, N139);
not NOT1 (N11525, N11521);
and AND3 (N11526, N11486, N4894, N5118);
xor XOR2 (N11527, N11524, N691);
buf BUF1 (N11528, N11508);
or OR3 (N11529, N11518, N9682, N10897);
and AND3 (N11530, N11525, N4109, N420);
nand NAND4 (N11531, N11499, N2844, N10795, N11070);
nand NAND3 (N11532, N11522, N11243, N5732);
nor NOR3 (N11533, N11494, N10618, N9509);
xor XOR2 (N11534, N11532, N5573);
nand NAND3 (N11535, N11534, N2694, N960);
nor NOR4 (N11536, N11520, N3052, N5301, N11324);
or OR2 (N11537, N11535, N4763);
nor NOR4 (N11538, N11530, N10308, N7618, N2836);
xor XOR2 (N11539, N11536, N2182);
nand NAND2 (N11540, N11516, N9884);
and AND2 (N11541, N11531, N8873);
nor NOR2 (N11542, N11541, N10974);
not NOT1 (N11543, N11529);
nand NAND3 (N11544, N11542, N8383, N3697);
buf BUF1 (N11545, N11528);
xor XOR2 (N11546, N11533, N218);
nand NAND3 (N11547, N11546, N385, N10572);
buf BUF1 (N11548, N11539);
buf BUF1 (N11549, N11540);
xor XOR2 (N11550, N11526, N5779);
nor NOR2 (N11551, N11545, N3906);
nor NOR3 (N11552, N11537, N5000, N9079);
buf BUF1 (N11553, N11549);
nand NAND3 (N11554, N11548, N5716, N6655);
and AND2 (N11555, N11543, N6561);
not NOT1 (N11556, N11550);
and AND3 (N11557, N11538, N4185, N6830);
or OR4 (N11558, N11552, N10161, N2167, N47);
nand NAND2 (N11559, N11527, N4931);
nand NAND2 (N11560, N11559, N7742);
and AND3 (N11561, N11547, N10705, N2418);
or OR4 (N11562, N11555, N5783, N11398, N2610);
nand NAND4 (N11563, N11562, N7016, N3019, N3531);
buf BUF1 (N11564, N11557);
nand NAND3 (N11565, N11554, N1033, N3990);
nor NOR3 (N11566, N11563, N2943, N3799);
nor NOR3 (N11567, N11560, N4549, N2220);
nand NAND2 (N11568, N11544, N4271);
or OR4 (N11569, N11566, N6649, N10122, N3659);
and AND2 (N11570, N11564, N4821);
nand NAND2 (N11571, N11556, N6115);
xor XOR2 (N11572, N11567, N6528);
and AND3 (N11573, N11570, N10322, N6391);
nor NOR3 (N11574, N11553, N2962, N8200);
xor XOR2 (N11575, N11569, N7425);
nor NOR4 (N11576, N11571, N11504, N11391, N4565);
or OR2 (N11577, N11568, N4774);
nand NAND3 (N11578, N11573, N8184, N6725);
nor NOR4 (N11579, N11576, N11209, N4431, N11513);
xor XOR2 (N11580, N11575, N9128);
xor XOR2 (N11581, N11561, N7029);
buf BUF1 (N11582, N11579);
nand NAND4 (N11583, N11581, N1734, N2010, N1725);
buf BUF1 (N11584, N11580);
xor XOR2 (N11585, N11572, N3572);
xor XOR2 (N11586, N11558, N5068);
buf BUF1 (N11587, N11574);
or OR4 (N11588, N11584, N3107, N5722, N1185);
not NOT1 (N11589, N11582);
buf BUF1 (N11590, N11577);
xor XOR2 (N11591, N11551, N2190);
and AND4 (N11592, N11587, N8633, N456, N8984);
not NOT1 (N11593, N11590);
buf BUF1 (N11594, N11588);
not NOT1 (N11595, N11592);
and AND3 (N11596, N11578, N7085, N820);
nor NOR4 (N11597, N11586, N2490, N1419, N6076);
nor NOR4 (N11598, N11565, N3820, N1986, N6811);
xor XOR2 (N11599, N11595, N2081);
or OR3 (N11600, N11599, N2176, N587);
not NOT1 (N11601, N11589);
nor NOR2 (N11602, N11596, N9082);
nor NOR3 (N11603, N11601, N3618, N2419);
xor XOR2 (N11604, N11602, N813);
nor NOR4 (N11605, N11604, N4226, N1579, N10711);
buf BUF1 (N11606, N11597);
not NOT1 (N11607, N11594);
nor NOR3 (N11608, N11598, N8227, N2548);
xor XOR2 (N11609, N11608, N9853);
xor XOR2 (N11610, N11591, N10222);
buf BUF1 (N11611, N11603);
not NOT1 (N11612, N11600);
buf BUF1 (N11613, N11585);
nor NOR2 (N11614, N11606, N2509);
nor NOR4 (N11615, N11607, N4238, N4906, N10962);
buf BUF1 (N11616, N11583);
nand NAND4 (N11617, N11593, N10429, N3451, N6785);
nor NOR3 (N11618, N11613, N7160, N8542);
nor NOR3 (N11619, N11614, N6619, N10703);
not NOT1 (N11620, N11610);
nand NAND4 (N11621, N11605, N5162, N361, N1649);
not NOT1 (N11622, N11615);
xor XOR2 (N11623, N11609, N9133);
and AND2 (N11624, N11611, N9331);
xor XOR2 (N11625, N11612, N10976);
xor XOR2 (N11626, N11625, N7073);
buf BUF1 (N11627, N11621);
xor XOR2 (N11628, N11616, N7967);
not NOT1 (N11629, N11624);
and AND4 (N11630, N11629, N6060, N9670, N10429);
not NOT1 (N11631, N11618);
not NOT1 (N11632, N11630);
and AND4 (N11633, N11620, N7592, N2341, N6484);
and AND2 (N11634, N11619, N6214);
buf BUF1 (N11635, N11633);
xor XOR2 (N11636, N11623, N10986);
not NOT1 (N11637, N11622);
and AND4 (N11638, N11631, N8476, N1077, N4797);
nor NOR3 (N11639, N11628, N1183, N3552);
xor XOR2 (N11640, N11632, N4382);
buf BUF1 (N11641, N11639);
nand NAND2 (N11642, N11635, N896);
and AND2 (N11643, N11627, N2031);
or OR4 (N11644, N11638, N7455, N6864, N11484);
nor NOR3 (N11645, N11640, N10917, N4805);
and AND3 (N11646, N11626, N5625, N631);
nor NOR4 (N11647, N11642, N2486, N9836, N8973);
xor XOR2 (N11648, N11647, N2326);
or OR2 (N11649, N11648, N10282);
nor NOR2 (N11650, N11637, N2475);
nand NAND3 (N11651, N11617, N1755, N7987);
not NOT1 (N11652, N11644);
not NOT1 (N11653, N11646);
and AND2 (N11654, N11651, N1059);
and AND4 (N11655, N11641, N10458, N8054, N1897);
and AND4 (N11656, N11643, N9087, N3225, N6633);
nor NOR2 (N11657, N11652, N4741);
buf BUF1 (N11658, N11634);
buf BUF1 (N11659, N11658);
buf BUF1 (N11660, N11657);
xor XOR2 (N11661, N11659, N8870);
buf BUF1 (N11662, N11649);
and AND2 (N11663, N11660, N2275);
not NOT1 (N11664, N11653);
nor NOR2 (N11665, N11656, N3279);
nand NAND3 (N11666, N11663, N98, N66);
or OR3 (N11667, N11662, N2488, N9638);
or OR2 (N11668, N11665, N697);
nor NOR4 (N11669, N11666, N9176, N10818, N2888);
nor NOR4 (N11670, N11664, N2152, N10947, N2625);
xor XOR2 (N11671, N11636, N11414);
or OR2 (N11672, N11671, N3065);
nand NAND4 (N11673, N11650, N8429, N10314, N6942);
not NOT1 (N11674, N11654);
buf BUF1 (N11675, N11645);
nor NOR4 (N11676, N11672, N2111, N7559, N6156);
and AND4 (N11677, N11655, N5444, N9895, N1899);
or OR2 (N11678, N11673, N7785);
xor XOR2 (N11679, N11675, N4594);
nor NOR2 (N11680, N11678, N4743);
xor XOR2 (N11681, N11674, N8762);
nand NAND4 (N11682, N11670, N10427, N4170, N1520);
buf BUF1 (N11683, N11679);
nand NAND2 (N11684, N11667, N4660);
buf BUF1 (N11685, N11683);
nor NOR3 (N11686, N11685, N8790, N1239);
and AND2 (N11687, N11680, N9732);
and AND4 (N11688, N11661, N1539, N3641, N9818);
and AND2 (N11689, N11668, N6278);
buf BUF1 (N11690, N11686);
nand NAND3 (N11691, N11669, N2465, N2592);
nor NOR2 (N11692, N11690, N271);
and AND4 (N11693, N11687, N8612, N6926, N10031);
or OR2 (N11694, N11677, N2406);
xor XOR2 (N11695, N11689, N1516);
or OR3 (N11696, N11684, N5290, N7022);
nor NOR4 (N11697, N11694, N9524, N3614, N4795);
nor NOR2 (N11698, N11692, N10711);
nor NOR3 (N11699, N11697, N542, N4053);
nand NAND3 (N11700, N11691, N5333, N1537);
or OR4 (N11701, N11695, N4614, N10076, N9805);
and AND3 (N11702, N11700, N57, N3878);
or OR2 (N11703, N11681, N3989);
nand NAND3 (N11704, N11693, N11183, N559);
and AND3 (N11705, N11682, N5555, N10162);
not NOT1 (N11706, N11705);
buf BUF1 (N11707, N11706);
not NOT1 (N11708, N11704);
and AND4 (N11709, N11699, N4944, N6782, N7109);
nor NOR2 (N11710, N11676, N5918);
nor NOR2 (N11711, N11709, N4274);
or OR2 (N11712, N11696, N11248);
nor NOR4 (N11713, N11703, N4787, N8099, N9027);
xor XOR2 (N11714, N11710, N10132);
or OR2 (N11715, N11688, N8218);
nor NOR2 (N11716, N11711, N1214);
buf BUF1 (N11717, N11707);
nand NAND4 (N11718, N11715, N941, N318, N11324);
and AND4 (N11719, N11717, N719, N11218, N2437);
xor XOR2 (N11720, N11719, N7768);
not NOT1 (N11721, N11701);
nand NAND4 (N11722, N11714, N10089, N6413, N2534);
or OR4 (N11723, N11712, N5158, N8944, N11247);
or OR3 (N11724, N11716, N9644, N1169);
buf BUF1 (N11725, N11722);
xor XOR2 (N11726, N11708, N9443);
and AND3 (N11727, N11698, N2628, N8734);
xor XOR2 (N11728, N11702, N987);
or OR2 (N11729, N11713, N9495);
not NOT1 (N11730, N11724);
xor XOR2 (N11731, N11720, N7036);
or OR4 (N11732, N11729, N4887, N917, N8465);
nand NAND4 (N11733, N11731, N4542, N40, N8791);
buf BUF1 (N11734, N11718);
or OR2 (N11735, N11728, N986);
or OR3 (N11736, N11726, N9596, N11653);
not NOT1 (N11737, N11733);
buf BUF1 (N11738, N11727);
buf BUF1 (N11739, N11738);
nand NAND4 (N11740, N11739, N6117, N9915, N9174);
buf BUF1 (N11741, N11732);
nor NOR3 (N11742, N11741, N4931, N11353);
or OR2 (N11743, N11721, N8193);
not NOT1 (N11744, N11737);
xor XOR2 (N11745, N11736, N7249);
nand NAND2 (N11746, N11735, N2768);
not NOT1 (N11747, N11723);
or OR4 (N11748, N11734, N5387, N6408, N50);
xor XOR2 (N11749, N11744, N3125);
nand NAND2 (N11750, N11725, N3520);
and AND3 (N11751, N11748, N6408, N9787);
and AND4 (N11752, N11745, N9820, N2193, N8312);
not NOT1 (N11753, N11750);
xor XOR2 (N11754, N11749, N6866);
nand NAND3 (N11755, N11742, N5484, N5145);
nand NAND4 (N11756, N11751, N4900, N6817, N5330);
nand NAND3 (N11757, N11743, N3582, N6317);
xor XOR2 (N11758, N11752, N2749);
and AND2 (N11759, N11753, N2180);
or OR3 (N11760, N11754, N9033, N3774);
buf BUF1 (N11761, N11758);
nand NAND2 (N11762, N11759, N9776);
xor XOR2 (N11763, N11747, N10061);
and AND3 (N11764, N11762, N1237, N9653);
or OR2 (N11765, N11764, N5318);
or OR4 (N11766, N11761, N3244, N3403, N8949);
xor XOR2 (N11767, N11746, N11698);
or OR4 (N11768, N11730, N9612, N5835, N3646);
not NOT1 (N11769, N11768);
xor XOR2 (N11770, N11756, N6359);
or OR2 (N11771, N11755, N9858);
and AND3 (N11772, N11770, N8562, N4303);
or OR2 (N11773, N11772, N7244);
buf BUF1 (N11774, N11763);
not NOT1 (N11775, N11771);
nor NOR4 (N11776, N11769, N9579, N8227, N11228);
nand NAND3 (N11777, N11776, N4787, N6916);
buf BUF1 (N11778, N11775);
not NOT1 (N11779, N11767);
nand NAND4 (N11780, N11778, N1635, N3452, N458);
or OR2 (N11781, N11766, N11289);
xor XOR2 (N11782, N11780, N9108);
xor XOR2 (N11783, N11779, N1445);
nand NAND4 (N11784, N11774, N503, N6405, N7292);
buf BUF1 (N11785, N11757);
xor XOR2 (N11786, N11784, N6135);
or OR2 (N11787, N11783, N2903);
xor XOR2 (N11788, N11781, N5311);
nand NAND2 (N11789, N11777, N3472);
buf BUF1 (N11790, N11787);
nand NAND2 (N11791, N11786, N11572);
and AND3 (N11792, N11782, N365, N7756);
and AND3 (N11793, N11785, N430, N6072);
not NOT1 (N11794, N11773);
not NOT1 (N11795, N11793);
not NOT1 (N11796, N11792);
and AND3 (N11797, N11790, N6269, N4758);
not NOT1 (N11798, N11765);
not NOT1 (N11799, N11788);
or OR4 (N11800, N11791, N957, N9949, N4249);
nor NOR3 (N11801, N11800, N9519, N1495);
or OR2 (N11802, N11794, N892);
xor XOR2 (N11803, N11796, N2111);
nand NAND4 (N11804, N11740, N3570, N8362, N5466);
xor XOR2 (N11805, N11802, N4946);
xor XOR2 (N11806, N11804, N2822);
buf BUF1 (N11807, N11795);
or OR3 (N11808, N11789, N108, N9696);
not NOT1 (N11809, N11799);
nor NOR3 (N11810, N11807, N7079, N11031);
xor XOR2 (N11811, N11809, N5794);
or OR4 (N11812, N11801, N7826, N4556, N1860);
nand NAND4 (N11813, N11798, N1852, N389, N992);
nor NOR2 (N11814, N11760, N4014);
xor XOR2 (N11815, N11814, N7635);
xor XOR2 (N11816, N11812, N10010);
and AND4 (N11817, N11811, N10481, N2728, N5231);
xor XOR2 (N11818, N11815, N2704);
not NOT1 (N11819, N11806);
and AND4 (N11820, N11810, N6206, N10020, N4790);
nor NOR2 (N11821, N11816, N7204);
nand NAND2 (N11822, N11821, N586);
nor NOR2 (N11823, N11817, N500);
and AND4 (N11824, N11819, N10295, N8635, N4859);
xor XOR2 (N11825, N11818, N1930);
xor XOR2 (N11826, N11822, N8304);
xor XOR2 (N11827, N11820, N7417);
not NOT1 (N11828, N11803);
nand NAND4 (N11829, N11824, N6756, N1861, N10790);
not NOT1 (N11830, N11813);
buf BUF1 (N11831, N11823);
not NOT1 (N11832, N11829);
not NOT1 (N11833, N11825);
and AND3 (N11834, N11827, N2514, N6728);
nand NAND3 (N11835, N11830, N5451, N6437);
xor XOR2 (N11836, N11831, N11192);
nor NOR4 (N11837, N11808, N3339, N11020, N5100);
nand NAND2 (N11838, N11826, N4367);
or OR2 (N11839, N11838, N2595);
buf BUF1 (N11840, N11833);
nand NAND2 (N11841, N11834, N11152);
not NOT1 (N11842, N11828);
xor XOR2 (N11843, N11837, N6972);
not NOT1 (N11844, N11840);
nor NOR3 (N11845, N11839, N8578, N3027);
nand NAND2 (N11846, N11841, N5574);
nand NAND3 (N11847, N11844, N5706, N8111);
nand NAND4 (N11848, N11846, N3360, N3634, N1462);
and AND3 (N11849, N11797, N8717, N8936);
nand NAND4 (N11850, N11849, N8049, N11612, N708);
nor NOR4 (N11851, N11835, N9845, N6453, N6774);
and AND3 (N11852, N11836, N6280, N10822);
and AND3 (N11853, N11845, N8876, N11455);
nor NOR4 (N11854, N11850, N605, N13, N7156);
nand NAND3 (N11855, N11848, N1053, N8914);
or OR4 (N11856, N11854, N11158, N6213, N4081);
or OR2 (N11857, N11852, N1208);
buf BUF1 (N11858, N11805);
nand NAND4 (N11859, N11832, N3536, N7732, N2502);
nand NAND2 (N11860, N11847, N10399);
and AND3 (N11861, N11856, N147, N5297);
nand NAND4 (N11862, N11859, N8848, N555, N2581);
or OR2 (N11863, N11853, N10894);
nand NAND3 (N11864, N11862, N3175, N1926);
xor XOR2 (N11865, N11860, N3268);
buf BUF1 (N11866, N11861);
nor NOR3 (N11867, N11858, N1982, N6409);
nor NOR3 (N11868, N11863, N2506, N6745);
nand NAND3 (N11869, N11865, N10249, N10262);
not NOT1 (N11870, N11843);
and AND3 (N11871, N11870, N7072, N2491);
nand NAND2 (N11872, N11857, N4057);
nand NAND2 (N11873, N11867, N9005);
or OR2 (N11874, N11842, N4487);
xor XOR2 (N11875, N11851, N7773);
nor NOR2 (N11876, N11873, N11205);
or OR4 (N11877, N11875, N3179, N2508, N3512);
nand NAND4 (N11878, N11868, N1601, N10100, N7460);
nor NOR2 (N11879, N11877, N7562);
nand NAND3 (N11880, N11878, N4929, N6199);
xor XOR2 (N11881, N11871, N7138);
not NOT1 (N11882, N11864);
not NOT1 (N11883, N11880);
not NOT1 (N11884, N11881);
xor XOR2 (N11885, N11879, N2372);
xor XOR2 (N11886, N11876, N7102);
xor XOR2 (N11887, N11855, N24);
nor NOR4 (N11888, N11883, N2175, N8450, N10243);
and AND4 (N11889, N11888, N2515, N2707, N6605);
nand NAND2 (N11890, N11882, N8629);
nor NOR3 (N11891, N11884, N5394, N11356);
not NOT1 (N11892, N11885);
or OR2 (N11893, N11890, N2329);
nand NAND4 (N11894, N11866, N857, N10969, N430);
buf BUF1 (N11895, N11872);
nor NOR2 (N11896, N11891, N4935);
nand NAND2 (N11897, N11889, N5137);
or OR4 (N11898, N11893, N8283, N6557, N7091);
buf BUF1 (N11899, N11896);
and AND3 (N11900, N11892, N6642, N6446);
buf BUF1 (N11901, N11887);
nand NAND3 (N11902, N11894, N11632, N11336);
nor NOR2 (N11903, N11897, N7612);
or OR2 (N11904, N11886, N4190);
not NOT1 (N11905, N11900);
nor NOR4 (N11906, N11902, N4071, N7246, N1789);
nor NOR2 (N11907, N11874, N2263);
buf BUF1 (N11908, N11905);
nand NAND2 (N11909, N11907, N4415);
or OR3 (N11910, N11906, N11424, N418);
nor NOR3 (N11911, N11898, N530, N1471);
xor XOR2 (N11912, N11910, N2048);
not NOT1 (N11913, N11903);
nand NAND2 (N11914, N11908, N11077);
nor NOR4 (N11915, N11899, N11006, N11657, N7875);
buf BUF1 (N11916, N11911);
xor XOR2 (N11917, N11909, N6669);
and AND3 (N11918, N11913, N6226, N1187);
nor NOR3 (N11919, N11912, N664, N6736);
nor NOR2 (N11920, N11918, N885);
buf BUF1 (N11921, N11914);
nor NOR4 (N11922, N11869, N1090, N6054, N3696);
or OR3 (N11923, N11922, N11787, N6088);
not NOT1 (N11924, N11919);
or OR4 (N11925, N11917, N9750, N10477, N4153);
buf BUF1 (N11926, N11921);
or OR2 (N11927, N11915, N11682);
xor XOR2 (N11928, N11904, N2430);
not NOT1 (N11929, N11901);
not NOT1 (N11930, N11925);
nand NAND2 (N11931, N11926, N1211);
and AND3 (N11932, N11927, N7854, N1328);
not NOT1 (N11933, N11931);
xor XOR2 (N11934, N11928, N165);
and AND3 (N11935, N11932, N5264, N3665);
and AND4 (N11936, N11923, N4178, N11731, N10122);
nor NOR2 (N11937, N11936, N6558);
nor NOR3 (N11938, N11935, N11578, N7301);
and AND2 (N11939, N11929, N1300);
not NOT1 (N11940, N11934);
not NOT1 (N11941, N11937);
nor NOR2 (N11942, N11895, N9391);
or OR2 (N11943, N11942, N853);
buf BUF1 (N11944, N11916);
buf BUF1 (N11945, N11939);
nor NOR4 (N11946, N11945, N9157, N1837, N8727);
or OR4 (N11947, N11924, N11481, N1486, N10448);
nand NAND2 (N11948, N11938, N168);
not NOT1 (N11949, N11946);
nor NOR2 (N11950, N11944, N5168);
not NOT1 (N11951, N11930);
or OR4 (N11952, N11948, N1751, N3285, N6889);
not NOT1 (N11953, N11933);
nand NAND3 (N11954, N11947, N2976, N8881);
not NOT1 (N11955, N11940);
buf BUF1 (N11956, N11950);
xor XOR2 (N11957, N11955, N7916);
and AND2 (N11958, N11957, N7845);
or OR4 (N11959, N11952, N2653, N5096, N3286);
xor XOR2 (N11960, N11958, N1030);
buf BUF1 (N11961, N11949);
buf BUF1 (N11962, N11959);
nand NAND4 (N11963, N11961, N9125, N3245, N7673);
nor NOR3 (N11964, N11962, N7410, N1711);
buf BUF1 (N11965, N11953);
buf BUF1 (N11966, N11965);
nand NAND4 (N11967, N11943, N4281, N5512, N7407);
xor XOR2 (N11968, N11967, N6266);
buf BUF1 (N11969, N11954);
nor NOR4 (N11970, N11956, N462, N3494, N6467);
not NOT1 (N11971, N11969);
xor XOR2 (N11972, N11951, N6268);
xor XOR2 (N11973, N11920, N4896);
not NOT1 (N11974, N11972);
not NOT1 (N11975, N11964);
xor XOR2 (N11976, N11974, N2521);
and AND3 (N11977, N11970, N7839, N7568);
buf BUF1 (N11978, N11975);
nor NOR3 (N11979, N11973, N1985, N3388);
or OR2 (N11980, N11971, N3586);
not NOT1 (N11981, N11963);
nand NAND4 (N11982, N11980, N1017, N5408, N3308);
or OR2 (N11983, N11981, N7518);
or OR4 (N11984, N11977, N7005, N668, N5538);
xor XOR2 (N11985, N11983, N7933);
and AND2 (N11986, N11978, N1200);
or OR3 (N11987, N11941, N10407, N2852);
xor XOR2 (N11988, N11979, N7187);
not NOT1 (N11989, N11984);
or OR2 (N11990, N11960, N11154);
or OR2 (N11991, N11985, N4267);
nor NOR3 (N11992, N11988, N5962, N8094);
not NOT1 (N11993, N11991);
buf BUF1 (N11994, N11986);
nand NAND2 (N11995, N11968, N9472);
xor XOR2 (N11996, N11982, N5111);
nor NOR4 (N11997, N11987, N11341, N2262, N11533);
or OR3 (N11998, N11993, N1464, N1124);
nand NAND2 (N11999, N11989, N11959);
not NOT1 (N12000, N11997);
nand NAND2 (N12001, N11998, N2493);
and AND4 (N12002, N12001, N545, N1439, N4382);
or OR4 (N12003, N11966, N11148, N10436, N1000);
buf BUF1 (N12004, N12002);
nand NAND3 (N12005, N11996, N1143, N3770);
not NOT1 (N12006, N12003);
or OR3 (N12007, N12004, N11884, N1517);
or OR4 (N12008, N11994, N8655, N8677, N4977);
not NOT1 (N12009, N11992);
xor XOR2 (N12010, N11999, N6207);
buf BUF1 (N12011, N11976);
nor NOR3 (N12012, N12008, N6445, N4052);
and AND2 (N12013, N11995, N860);
xor XOR2 (N12014, N12006, N11167);
not NOT1 (N12015, N12007);
not NOT1 (N12016, N12010);
not NOT1 (N12017, N12016);
not NOT1 (N12018, N12015);
or OR2 (N12019, N12005, N8736);
nand NAND4 (N12020, N12012, N7003, N5829, N11171);
or OR2 (N12021, N12000, N8690);
nor NOR4 (N12022, N12018, N9231, N1294, N3963);
buf BUF1 (N12023, N12011);
buf BUF1 (N12024, N12013);
nor NOR4 (N12025, N12017, N6665, N9599, N10872);
or OR4 (N12026, N12019, N1620, N10480, N5565);
not NOT1 (N12027, N12021);
xor XOR2 (N12028, N12020, N2808);
buf BUF1 (N12029, N12028);
nor NOR3 (N12030, N12027, N8868, N5252);
not NOT1 (N12031, N12030);
xor XOR2 (N12032, N12022, N10033);
nand NAND3 (N12033, N12031, N165, N3963);
nor NOR3 (N12034, N12023, N3141, N4361);
xor XOR2 (N12035, N11990, N5201);
not NOT1 (N12036, N12032);
and AND3 (N12037, N12024, N11393, N6554);
and AND3 (N12038, N12037, N6131, N5733);
not NOT1 (N12039, N12009);
buf BUF1 (N12040, N12029);
nor NOR2 (N12041, N12034, N1859);
or OR3 (N12042, N12036, N5099, N3440);
or OR4 (N12043, N12040, N9420, N165, N10466);
or OR2 (N12044, N12042, N546);
buf BUF1 (N12045, N12038);
or OR3 (N12046, N12025, N2129, N4324);
buf BUF1 (N12047, N12046);
and AND3 (N12048, N12041, N5115, N4414);
and AND2 (N12049, N12035, N8172);
nand NAND4 (N12050, N12043, N7378, N9232, N1601);
nor NOR4 (N12051, N12045, N2848, N9508, N2006);
xor XOR2 (N12052, N12049, N52);
nand NAND2 (N12053, N12047, N4653);
not NOT1 (N12054, N12044);
nor NOR4 (N12055, N12039, N6349, N9017, N6329);
buf BUF1 (N12056, N12014);
buf BUF1 (N12057, N12026);
nor NOR4 (N12058, N12053, N5133, N8774, N5664);
and AND2 (N12059, N12054, N9589);
or OR3 (N12060, N12050, N10920, N3687);
not NOT1 (N12061, N12055);
not NOT1 (N12062, N12058);
nor NOR4 (N12063, N12060, N7134, N11627, N1311);
not NOT1 (N12064, N12061);
not NOT1 (N12065, N12063);
xor XOR2 (N12066, N12057, N398);
not NOT1 (N12067, N12051);
nand NAND4 (N12068, N12065, N9998, N10415, N3519);
nand NAND4 (N12069, N12033, N6828, N11593, N11385);
not NOT1 (N12070, N12059);
buf BUF1 (N12071, N12067);
and AND3 (N12072, N12048, N4397, N8794);
nor NOR2 (N12073, N12069, N4014);
nand NAND4 (N12074, N12066, N8520, N10384, N7574);
nor NOR3 (N12075, N12070, N2457, N2493);
not NOT1 (N12076, N12068);
or OR3 (N12077, N12056, N587, N2106);
or OR3 (N12078, N12073, N11942, N10626);
xor XOR2 (N12079, N12062, N2236);
xor XOR2 (N12080, N12075, N4808);
or OR3 (N12081, N12076, N2518, N9721);
and AND2 (N12082, N12081, N5838);
not NOT1 (N12083, N12080);
buf BUF1 (N12084, N12071);
not NOT1 (N12085, N12077);
xor XOR2 (N12086, N12074, N1638);
nor NOR3 (N12087, N12052, N4840, N5095);
buf BUF1 (N12088, N12072);
xor XOR2 (N12089, N12064, N8870);
nor NOR2 (N12090, N12088, N2399);
and AND4 (N12091, N12078, N8196, N9948, N705);
buf BUF1 (N12092, N12089);
buf BUF1 (N12093, N12083);
and AND2 (N12094, N12091, N6379);
xor XOR2 (N12095, N12094, N9260);
nand NAND2 (N12096, N12093, N11173);
nor NOR4 (N12097, N12095, N6858, N11342, N9512);
xor XOR2 (N12098, N12096, N3290);
xor XOR2 (N12099, N12098, N5892);
and AND4 (N12100, N12092, N1526, N1949, N4529);
and AND4 (N12101, N12082, N2759, N1967, N854);
nor NOR4 (N12102, N12097, N9961, N8841, N4626);
not NOT1 (N12103, N12100);
nor NOR4 (N12104, N12103, N944, N6162, N9424);
or OR2 (N12105, N12079, N4487);
not NOT1 (N12106, N12087);
buf BUF1 (N12107, N12085);
buf BUF1 (N12108, N12086);
not NOT1 (N12109, N12105);
buf BUF1 (N12110, N12099);
not NOT1 (N12111, N12104);
buf BUF1 (N12112, N12107);
not NOT1 (N12113, N12102);
not NOT1 (N12114, N12113);
xor XOR2 (N12115, N12111, N4960);
buf BUF1 (N12116, N12108);
and AND3 (N12117, N12090, N9040, N9062);
and AND4 (N12118, N12116, N8511, N6414, N8556);
nor NOR2 (N12119, N12109, N10250);
nor NOR4 (N12120, N12112, N6214, N4931, N11440);
and AND3 (N12121, N12118, N2572, N5855);
not NOT1 (N12122, N12084);
not NOT1 (N12123, N12121);
and AND3 (N12124, N12120, N10819, N637);
and AND3 (N12125, N12114, N9824, N9967);
not NOT1 (N12126, N12123);
not NOT1 (N12127, N12119);
or OR2 (N12128, N12127, N2540);
or OR4 (N12129, N12128, N1979, N111, N10641);
nor NOR2 (N12130, N12126, N5204);
buf BUF1 (N12131, N12124);
not NOT1 (N12132, N12131);
nand NAND4 (N12133, N12132, N7853, N2195, N9773);
and AND3 (N12134, N12129, N10509, N10848);
not NOT1 (N12135, N12130);
and AND2 (N12136, N12133, N6572);
and AND2 (N12137, N12117, N11659);
not NOT1 (N12138, N12110);
nor NOR3 (N12139, N12134, N12055, N1569);
nand NAND2 (N12140, N12139, N1242);
and AND2 (N12141, N12115, N6065);
nand NAND4 (N12142, N12101, N9360, N10354, N9560);
nand NAND3 (N12143, N12122, N4338, N4550);
not NOT1 (N12144, N12135);
and AND4 (N12145, N12143, N5947, N918, N11460);
and AND2 (N12146, N12144, N6588);
or OR2 (N12147, N12140, N6211);
nand NAND4 (N12148, N12125, N10852, N274, N3217);
xor XOR2 (N12149, N12141, N11582);
nor NOR2 (N12150, N12149, N2040);
nor NOR4 (N12151, N12146, N11054, N7058, N11135);
nand NAND3 (N12152, N12145, N5032, N5783);
or OR3 (N12153, N12150, N5193, N12064);
nand NAND2 (N12154, N12152, N3060);
nand NAND2 (N12155, N12106, N7477);
nand NAND2 (N12156, N12148, N2985);
buf BUF1 (N12157, N12137);
not NOT1 (N12158, N12157);
not NOT1 (N12159, N12156);
not NOT1 (N12160, N12151);
not NOT1 (N12161, N12138);
nand NAND4 (N12162, N12136, N8782, N8182, N541);
not NOT1 (N12163, N12154);
or OR2 (N12164, N12163, N2862);
or OR2 (N12165, N12142, N7541);
or OR3 (N12166, N12158, N8734, N3516);
nand NAND3 (N12167, N12165, N3140, N9794);
nor NOR2 (N12168, N12159, N7479);
or OR3 (N12169, N12164, N8017, N4316);
xor XOR2 (N12170, N12161, N279);
and AND3 (N12171, N12155, N6936, N4854);
nand NAND4 (N12172, N12162, N10374, N11594, N4549);
not NOT1 (N12173, N12168);
nor NOR4 (N12174, N12147, N3898, N8364, N1999);
buf BUF1 (N12175, N12160);
nor NOR2 (N12176, N12170, N11013);
nand NAND3 (N12177, N12174, N10152, N2224);
or OR2 (N12178, N12176, N12000);
not NOT1 (N12179, N12173);
or OR3 (N12180, N12169, N9527, N7992);
nand NAND3 (N12181, N12153, N2242, N4147);
and AND2 (N12182, N12166, N11809);
and AND3 (N12183, N12177, N7307, N9995);
buf BUF1 (N12184, N12182);
nor NOR3 (N12185, N12183, N7847, N2082);
not NOT1 (N12186, N12178);
nand NAND3 (N12187, N12172, N9933, N1408);
and AND2 (N12188, N12186, N12050);
not NOT1 (N12189, N12167);
buf BUF1 (N12190, N12175);
and AND2 (N12191, N12181, N4829);
or OR2 (N12192, N12185, N6197);
xor XOR2 (N12193, N12179, N4147);
buf BUF1 (N12194, N12184);
and AND2 (N12195, N12192, N6888);
nand NAND2 (N12196, N12188, N9354);
xor XOR2 (N12197, N12195, N612);
not NOT1 (N12198, N12197);
or OR4 (N12199, N12187, N2196, N3405, N2994);
xor XOR2 (N12200, N12193, N7149);
xor XOR2 (N12201, N12199, N9506);
nor NOR3 (N12202, N12198, N1362, N5696);
nor NOR4 (N12203, N12189, N4302, N8689, N921);
buf BUF1 (N12204, N12201);
nand NAND4 (N12205, N12203, N620, N8290, N8656);
xor XOR2 (N12206, N12204, N10291);
nor NOR3 (N12207, N12196, N3726, N2096);
nand NAND3 (N12208, N12190, N8063, N1697);
and AND4 (N12209, N12171, N9816, N132, N1506);
and AND4 (N12210, N12208, N1168, N6965, N2335);
not NOT1 (N12211, N12206);
and AND4 (N12212, N12210, N7874, N10022, N3839);
buf BUF1 (N12213, N12209);
or OR3 (N12214, N12191, N9081, N11928);
nand NAND3 (N12215, N12205, N5945, N170);
and AND4 (N12216, N12212, N879, N5819, N11837);
xor XOR2 (N12217, N12211, N5634);
and AND2 (N12218, N12217, N5584);
or OR4 (N12219, N12200, N408, N10123, N2495);
nand NAND3 (N12220, N12219, N6030, N2333);
xor XOR2 (N12221, N12202, N11575);
xor XOR2 (N12222, N12214, N1657);
and AND2 (N12223, N12222, N1381);
buf BUF1 (N12224, N12220);
or OR2 (N12225, N12224, N8775);
not NOT1 (N12226, N12225);
buf BUF1 (N12227, N12180);
not NOT1 (N12228, N12218);
or OR3 (N12229, N12194, N11771, N12020);
nor NOR3 (N12230, N12213, N10199, N6211);
nand NAND3 (N12231, N12227, N933, N4253);
xor XOR2 (N12232, N12215, N10627);
xor XOR2 (N12233, N12207, N9520);
and AND3 (N12234, N12229, N9148, N2156);
not NOT1 (N12235, N12221);
not NOT1 (N12236, N12226);
not NOT1 (N12237, N12234);
or OR4 (N12238, N12233, N2233, N2169, N7535);
nor NOR2 (N12239, N12236, N4772);
buf BUF1 (N12240, N12232);
xor XOR2 (N12241, N12216, N8854);
and AND2 (N12242, N12223, N3623);
and AND4 (N12243, N12230, N2910, N1460, N12028);
and AND4 (N12244, N12242, N134, N7211, N7021);
and AND4 (N12245, N12228, N1387, N828, N6394);
or OR4 (N12246, N12243, N6640, N3846, N2800);
and AND2 (N12247, N12231, N4527);
nor NOR2 (N12248, N12240, N7318);
nand NAND3 (N12249, N12238, N3565, N4243);
nor NOR2 (N12250, N12235, N10715);
nand NAND2 (N12251, N12247, N1494);
not NOT1 (N12252, N12244);
and AND4 (N12253, N12246, N7013, N9812, N11002);
and AND3 (N12254, N12250, N2728, N7168);
xor XOR2 (N12255, N12239, N9031);
not NOT1 (N12256, N12255);
nor NOR3 (N12257, N12254, N274, N11450);
nand NAND3 (N12258, N12237, N1680, N9362);
xor XOR2 (N12259, N12252, N832);
or OR2 (N12260, N12241, N139);
or OR4 (N12261, N12256, N5062, N371, N3586);
or OR4 (N12262, N12259, N1650, N9130, N3502);
or OR4 (N12263, N12253, N5108, N5942, N7037);
nand NAND4 (N12264, N12260, N1363, N1557, N1403);
xor XOR2 (N12265, N12262, N3537);
nand NAND3 (N12266, N12261, N669, N11);
not NOT1 (N12267, N12263);
xor XOR2 (N12268, N12264, N5331);
and AND3 (N12269, N12248, N685, N7100);
nand NAND4 (N12270, N12251, N1057, N7251, N1496);
or OR4 (N12271, N12267, N2558, N7945, N6422);
not NOT1 (N12272, N12249);
and AND2 (N12273, N12271, N8692);
nor NOR3 (N12274, N12265, N10943, N887);
buf BUF1 (N12275, N12258);
buf BUF1 (N12276, N12269);
not NOT1 (N12277, N12275);
and AND2 (N12278, N12274, N1582);
not NOT1 (N12279, N12268);
and AND2 (N12280, N12273, N11271);
not NOT1 (N12281, N12272);
nand NAND3 (N12282, N12281, N1677, N6565);
not NOT1 (N12283, N12257);
not NOT1 (N12284, N12279);
and AND3 (N12285, N12277, N8415, N3986);
buf BUF1 (N12286, N12276);
not NOT1 (N12287, N12285);
or OR3 (N12288, N12287, N1683, N5299);
not NOT1 (N12289, N12288);
not NOT1 (N12290, N12283);
xor XOR2 (N12291, N12290, N2924);
nand NAND4 (N12292, N12245, N7111, N3352, N538);
buf BUF1 (N12293, N12278);
nor NOR4 (N12294, N12270, N130, N2869, N271);
not NOT1 (N12295, N12293);
xor XOR2 (N12296, N12289, N10432);
buf BUF1 (N12297, N12286);
xor XOR2 (N12298, N12294, N1646);
not NOT1 (N12299, N12282);
xor XOR2 (N12300, N12298, N4421);
nand NAND3 (N12301, N12296, N10046, N1546);
nand NAND3 (N12302, N12280, N2788, N9669);
not NOT1 (N12303, N12302);
and AND2 (N12304, N12295, N9590);
xor XOR2 (N12305, N12303, N5171);
not NOT1 (N12306, N12284);
not NOT1 (N12307, N12301);
nor NOR2 (N12308, N12297, N742);
and AND2 (N12309, N12266, N6083);
xor XOR2 (N12310, N12309, N8454);
nand NAND2 (N12311, N12305, N4574);
not NOT1 (N12312, N12292);
or OR4 (N12313, N12312, N10032, N53, N4551);
not NOT1 (N12314, N12300);
nand NAND3 (N12315, N12311, N4567, N721);
nand NAND2 (N12316, N12308, N2190);
or OR3 (N12317, N12313, N3409, N8006);
nand NAND4 (N12318, N12306, N8998, N11085, N679);
and AND3 (N12319, N12315, N6363, N1151);
and AND2 (N12320, N12310, N5469);
and AND2 (N12321, N12317, N7893);
xor XOR2 (N12322, N12320, N2277);
xor XOR2 (N12323, N12304, N1940);
xor XOR2 (N12324, N12307, N4110);
not NOT1 (N12325, N12299);
and AND4 (N12326, N12321, N3943, N238, N4392);
not NOT1 (N12327, N12314);
and AND2 (N12328, N12324, N12314);
nand NAND3 (N12329, N12326, N2521, N6858);
xor XOR2 (N12330, N12291, N7269);
not NOT1 (N12331, N12318);
nand NAND4 (N12332, N12330, N10517, N1311, N1929);
xor XOR2 (N12333, N12332, N10312);
nor NOR4 (N12334, N12329, N10091, N8737, N7877);
nand NAND2 (N12335, N12327, N3085);
not NOT1 (N12336, N12319);
nand NAND4 (N12337, N12333, N8850, N1151, N10731);
and AND2 (N12338, N12316, N12154);
and AND2 (N12339, N12325, N5975);
not NOT1 (N12340, N12328);
xor XOR2 (N12341, N12337, N8470);
nor NOR3 (N12342, N12323, N9971, N11081);
buf BUF1 (N12343, N12336);
nand NAND3 (N12344, N12341, N4220, N57);
not NOT1 (N12345, N12344);
not NOT1 (N12346, N12334);
and AND4 (N12347, N12345, N5854, N7140, N4078);
not NOT1 (N12348, N12335);
or OR3 (N12349, N12347, N972, N3552);
nor NOR4 (N12350, N12339, N6671, N8830, N11740);
xor XOR2 (N12351, N12346, N3135);
nand NAND2 (N12352, N12348, N6283);
xor XOR2 (N12353, N12331, N8713);
not NOT1 (N12354, N12342);
nand NAND4 (N12355, N12338, N6012, N6956, N8751);
nand NAND3 (N12356, N12353, N4870, N287);
not NOT1 (N12357, N12343);
and AND4 (N12358, N12356, N1792, N12245, N6110);
or OR4 (N12359, N12354, N5290, N4234, N2121);
or OR2 (N12360, N12357, N7083);
not NOT1 (N12361, N12359);
buf BUF1 (N12362, N12361);
buf BUF1 (N12363, N12350);
nor NOR3 (N12364, N12349, N358, N3099);
not NOT1 (N12365, N12364);
nand NAND3 (N12366, N12365, N10260, N11004);
nor NOR3 (N12367, N12340, N4078, N1073);
buf BUF1 (N12368, N12322);
xor XOR2 (N12369, N12366, N5065);
and AND3 (N12370, N12367, N4595, N1146);
buf BUF1 (N12371, N12352);
buf BUF1 (N12372, N12355);
nand NAND4 (N12373, N12370, N1511, N11069, N8961);
and AND3 (N12374, N12351, N1280, N9163);
not NOT1 (N12375, N12369);
xor XOR2 (N12376, N12358, N8863);
buf BUF1 (N12377, N12360);
nor NOR2 (N12378, N12374, N7770);
nand NAND4 (N12379, N12368, N294, N6752, N7986);
nand NAND4 (N12380, N12372, N9277, N7820, N5012);
xor XOR2 (N12381, N12373, N4573);
nor NOR4 (N12382, N12377, N3853, N7804, N1151);
buf BUF1 (N12383, N12378);
not NOT1 (N12384, N12383);
nand NAND4 (N12385, N12376, N3477, N2237, N5620);
and AND2 (N12386, N12384, N5563);
and AND4 (N12387, N12380, N4742, N7485, N1462);
nor NOR2 (N12388, N12385, N6715);
or OR4 (N12389, N12375, N721, N7790, N11077);
buf BUF1 (N12390, N12363);
nand NAND4 (N12391, N12386, N8279, N6354, N7781);
and AND2 (N12392, N12379, N9037);
xor XOR2 (N12393, N12390, N4389);
xor XOR2 (N12394, N12362, N4210);
xor XOR2 (N12395, N12392, N4628);
or OR4 (N12396, N12382, N9123, N9551, N8498);
or OR4 (N12397, N12395, N5996, N11553, N9320);
and AND3 (N12398, N12393, N7042, N1483);
buf BUF1 (N12399, N12388);
not NOT1 (N12400, N12391);
nor NOR2 (N12401, N12399, N10792);
nor NOR4 (N12402, N12381, N5423, N310, N4928);
or OR2 (N12403, N12397, N12307);
and AND4 (N12404, N12401, N8400, N10095, N9852);
nand NAND4 (N12405, N12389, N4733, N6903, N1939);
buf BUF1 (N12406, N12403);
not NOT1 (N12407, N12394);
xor XOR2 (N12408, N12407, N8682);
not NOT1 (N12409, N12396);
nor NOR2 (N12410, N12387, N4145);
buf BUF1 (N12411, N12405);
nand NAND3 (N12412, N12406, N5001, N9408);
xor XOR2 (N12413, N12371, N10358);
and AND3 (N12414, N12398, N10284, N6559);
nor NOR2 (N12415, N12409, N1186);
or OR2 (N12416, N12415, N8116);
nand NAND3 (N12417, N12411, N1507, N8748);
or OR2 (N12418, N12400, N2592);
and AND4 (N12419, N12417, N10315, N7707, N7801);
and AND4 (N12420, N12408, N9906, N7659, N11644);
buf BUF1 (N12421, N12418);
xor XOR2 (N12422, N12419, N11011);
not NOT1 (N12423, N12404);
nand NAND4 (N12424, N12422, N8410, N4549, N3675);
and AND2 (N12425, N12424, N7082);
not NOT1 (N12426, N12413);
and AND4 (N12427, N12412, N10118, N10882, N2436);
buf BUF1 (N12428, N12427);
not NOT1 (N12429, N12425);
buf BUF1 (N12430, N12420);
xor XOR2 (N12431, N12428, N2233);
and AND3 (N12432, N12426, N11469, N4706);
not NOT1 (N12433, N12423);
nor NOR4 (N12434, N12432, N6131, N5236, N1463);
xor XOR2 (N12435, N12431, N11721);
not NOT1 (N12436, N12433);
nand NAND3 (N12437, N12421, N11867, N10743);
and AND3 (N12438, N12414, N10829, N9171);
and AND2 (N12439, N12434, N10324);
and AND2 (N12440, N12438, N9100);
and AND4 (N12441, N12416, N8582, N2909, N3932);
buf BUF1 (N12442, N12437);
and AND2 (N12443, N12442, N8443);
nor NOR2 (N12444, N12429, N9839);
and AND3 (N12445, N12402, N4336, N4164);
buf BUF1 (N12446, N12441);
and AND4 (N12447, N12439, N10548, N1033, N7895);
and AND2 (N12448, N12447, N10150);
buf BUF1 (N12449, N12410);
buf BUF1 (N12450, N12436);
or OR4 (N12451, N12443, N8343, N4157, N9233);
nand NAND4 (N12452, N12451, N2328, N2606, N3394);
or OR4 (N12453, N12430, N1851, N8222, N2040);
buf BUF1 (N12454, N12440);
and AND3 (N12455, N12444, N6826, N1677);
or OR3 (N12456, N12455, N5142, N11078);
and AND2 (N12457, N12452, N4378);
xor XOR2 (N12458, N12448, N11115);
or OR4 (N12459, N12457, N4006, N961, N9795);
not NOT1 (N12460, N12459);
nor NOR2 (N12461, N12460, N10836);
nor NOR2 (N12462, N12456, N11981);
nor NOR4 (N12463, N12435, N10720, N2142, N11641);
nand NAND4 (N12464, N12461, N4541, N11248, N4851);
xor XOR2 (N12465, N12464, N4009);
xor XOR2 (N12466, N12465, N10676);
xor XOR2 (N12467, N12454, N8091);
nand NAND2 (N12468, N12445, N9459);
buf BUF1 (N12469, N12463);
and AND2 (N12470, N12469, N3474);
xor XOR2 (N12471, N12468, N6386);
and AND2 (N12472, N12471, N418);
nand NAND2 (N12473, N12450, N11044);
nor NOR4 (N12474, N12473, N9941, N11894, N10493);
buf BUF1 (N12475, N12470);
xor XOR2 (N12476, N12474, N8157);
nand NAND2 (N12477, N12472, N7545);
and AND3 (N12478, N12466, N3983, N12121);
nor NOR4 (N12479, N12446, N7306, N11638, N11782);
buf BUF1 (N12480, N12462);
buf BUF1 (N12481, N12476);
nor NOR4 (N12482, N12453, N4147, N5140, N4737);
nor NOR3 (N12483, N12467, N4427, N2784);
or OR2 (N12484, N12449, N9408);
nor NOR2 (N12485, N12475, N11986);
xor XOR2 (N12486, N12477, N6583);
nor NOR4 (N12487, N12486, N7329, N158, N12077);
or OR3 (N12488, N12480, N2139, N10569);
nor NOR4 (N12489, N12487, N12098, N11559, N4565);
nand NAND3 (N12490, N12478, N7391, N11537);
xor XOR2 (N12491, N12484, N10626);
buf BUF1 (N12492, N12479);
buf BUF1 (N12493, N12482);
buf BUF1 (N12494, N12488);
not NOT1 (N12495, N12489);
and AND4 (N12496, N12494, N5665, N8834, N838);
xor XOR2 (N12497, N12485, N9370);
nand NAND2 (N12498, N12481, N3368);
not NOT1 (N12499, N12493);
or OR3 (N12500, N12492, N5538, N3826);
nand NAND2 (N12501, N12458, N4621);
and AND4 (N12502, N12499, N6366, N9843, N8089);
or OR2 (N12503, N12500, N2922);
and AND3 (N12504, N12502, N4945, N12333);
xor XOR2 (N12505, N12483, N4405);
buf BUF1 (N12506, N12501);
and AND3 (N12507, N12505, N4764, N3062);
xor XOR2 (N12508, N12495, N2836);
nor NOR2 (N12509, N12507, N1541);
and AND4 (N12510, N12498, N3926, N2860, N11503);
buf BUF1 (N12511, N12503);
or OR4 (N12512, N12509, N11964, N6532, N3173);
nand NAND4 (N12513, N12508, N7794, N11804, N5153);
xor XOR2 (N12514, N12490, N11772);
nor NOR4 (N12515, N12511, N11360, N732, N12451);
nor NOR4 (N12516, N12514, N11095, N961, N11215);
and AND4 (N12517, N12491, N1265, N8610, N1277);
nand NAND3 (N12518, N12506, N1749, N10715);
and AND2 (N12519, N12497, N9901);
nand NAND2 (N12520, N12515, N265);
buf BUF1 (N12521, N12496);
or OR2 (N12522, N12516, N3172);
or OR4 (N12523, N12517, N9961, N4053, N7531);
or OR4 (N12524, N12521, N801, N3994, N7804);
or OR4 (N12525, N12518, N12023, N9961, N5282);
buf BUF1 (N12526, N12524);
xor XOR2 (N12527, N12522, N2148);
or OR3 (N12528, N12504, N6983, N2488);
xor XOR2 (N12529, N12519, N526);
or OR2 (N12530, N12526, N6774);
buf BUF1 (N12531, N12512);
buf BUF1 (N12532, N12530);
buf BUF1 (N12533, N12513);
and AND3 (N12534, N12525, N6162, N6530);
and AND3 (N12535, N12534, N8043, N7267);
nor NOR4 (N12536, N12510, N3495, N8783, N5040);
nand NAND2 (N12537, N12535, N11392);
and AND3 (N12538, N12520, N4516, N6575);
and AND2 (N12539, N12531, N8354);
nor NOR3 (N12540, N12538, N6309, N466);
nand NAND3 (N12541, N12529, N7113, N7573);
not NOT1 (N12542, N12537);
nand NAND4 (N12543, N12542, N2272, N8135, N10468);
buf BUF1 (N12544, N12536);
not NOT1 (N12545, N12532);
buf BUF1 (N12546, N12544);
buf BUF1 (N12547, N12545);
not NOT1 (N12548, N12527);
or OR4 (N12549, N12541, N1480, N10203, N10663);
xor XOR2 (N12550, N12533, N4009);
xor XOR2 (N12551, N12549, N9697);
nand NAND2 (N12552, N12523, N3858);
or OR3 (N12553, N12546, N9981, N1737);
nand NAND4 (N12554, N12553, N232, N9156, N1852);
xor XOR2 (N12555, N12552, N3081);
nand NAND2 (N12556, N12543, N7771);
or OR4 (N12557, N12548, N2464, N5819, N5948);
and AND3 (N12558, N12557, N6437, N3407);
or OR4 (N12559, N12556, N2688, N12341, N4118);
nand NAND2 (N12560, N12551, N395);
and AND3 (N12561, N12540, N6664, N1723);
not NOT1 (N12562, N12550);
not NOT1 (N12563, N12562);
and AND2 (N12564, N12558, N10944);
nor NOR3 (N12565, N12560, N8746, N5169);
and AND4 (N12566, N12561, N10859, N10765, N9434);
not NOT1 (N12567, N12528);
and AND2 (N12568, N12565, N9713);
buf BUF1 (N12569, N12559);
xor XOR2 (N12570, N12569, N3244);
and AND2 (N12571, N12570, N6804);
nand NAND2 (N12572, N12571, N5853);
nand NAND2 (N12573, N12563, N9796);
and AND4 (N12574, N12554, N9535, N10949, N7837);
xor XOR2 (N12575, N12574, N2494);
nor NOR3 (N12576, N12567, N2486, N9185);
xor XOR2 (N12577, N12576, N5514);
and AND3 (N12578, N12547, N5420, N11370);
nor NOR2 (N12579, N12539, N2993);
nor NOR2 (N12580, N12579, N10351);
not NOT1 (N12581, N12564);
or OR2 (N12582, N12575, N7557);
nand NAND4 (N12583, N12568, N8973, N1501, N10693);
nor NOR3 (N12584, N12582, N4361, N747);
and AND2 (N12585, N12577, N7845);
nand NAND2 (N12586, N12580, N1367);
not NOT1 (N12587, N12566);
nor NOR2 (N12588, N12587, N6728);
not NOT1 (N12589, N12572);
and AND4 (N12590, N12578, N1037, N4702, N4968);
nand NAND3 (N12591, N12588, N5140, N1974);
buf BUF1 (N12592, N12590);
and AND2 (N12593, N12591, N11963);
not NOT1 (N12594, N12589);
nand NAND4 (N12595, N12555, N1981, N10580, N4778);
nor NOR3 (N12596, N12585, N734, N842);
buf BUF1 (N12597, N12581);
or OR2 (N12598, N12592, N2040);
or OR4 (N12599, N12598, N1267, N360, N11394);
xor XOR2 (N12600, N12586, N9908);
or OR4 (N12601, N12600, N7850, N7205, N9533);
and AND2 (N12602, N12597, N2468);
not NOT1 (N12603, N12599);
and AND4 (N12604, N12594, N306, N2838, N5274);
xor XOR2 (N12605, N12602, N9726);
nand NAND2 (N12606, N12595, N2213);
nor NOR4 (N12607, N12584, N8942, N254, N11314);
nor NOR4 (N12608, N12604, N5524, N12312, N616);
not NOT1 (N12609, N12607);
nor NOR4 (N12610, N12606, N614, N8294, N8319);
nand NAND2 (N12611, N12583, N7561);
xor XOR2 (N12612, N12603, N8669);
not NOT1 (N12613, N12610);
nand NAND3 (N12614, N12601, N635, N7170);
buf BUF1 (N12615, N12573);
or OR4 (N12616, N12609, N9483, N4267, N5412);
nand NAND3 (N12617, N12615, N5656, N4872);
or OR4 (N12618, N12613, N3256, N11233, N900);
xor XOR2 (N12619, N12617, N36);
nor NOR2 (N12620, N12614, N11042);
or OR3 (N12621, N12616, N1668, N1034);
xor XOR2 (N12622, N12620, N6534);
nor NOR3 (N12623, N12611, N1790, N6616);
and AND4 (N12624, N12593, N11474, N10779, N5857);
nand NAND4 (N12625, N12618, N2959, N6569, N6659);
and AND3 (N12626, N12622, N1707, N10001);
xor XOR2 (N12627, N12623, N6928);
buf BUF1 (N12628, N12605);
and AND4 (N12629, N12621, N10568, N10939, N9727);
or OR4 (N12630, N12629, N3041, N2548, N7042);
and AND3 (N12631, N12619, N8940, N46);
xor XOR2 (N12632, N12625, N6463);
and AND3 (N12633, N12596, N10268, N104);
and AND3 (N12634, N12608, N2167, N7310);
buf BUF1 (N12635, N12633);
and AND4 (N12636, N12627, N9159, N9867, N4814);
or OR2 (N12637, N12612, N1320);
or OR3 (N12638, N12626, N11216, N5952);
and AND4 (N12639, N12638, N11450, N10933, N2425);
nand NAND4 (N12640, N12624, N5278, N9125, N2752);
not NOT1 (N12641, N12635);
and AND3 (N12642, N12640, N7654, N11283);
or OR2 (N12643, N12630, N10961);
or OR4 (N12644, N12632, N649, N11882, N28);
nand NAND4 (N12645, N12642, N23, N8738, N7219);
buf BUF1 (N12646, N12637);
not NOT1 (N12647, N12644);
nand NAND2 (N12648, N12639, N4939);
xor XOR2 (N12649, N12634, N6133);
xor XOR2 (N12650, N12643, N9020);
nor NOR2 (N12651, N12646, N3580);
or OR2 (N12652, N12647, N6008);
not NOT1 (N12653, N12651);
or OR4 (N12654, N12636, N1536, N2041, N11502);
buf BUF1 (N12655, N12650);
and AND4 (N12656, N12654, N5136, N8692, N1905);
and AND4 (N12657, N12653, N2813, N5356, N8660);
or OR4 (N12658, N12641, N2298, N8963, N4577);
and AND4 (N12659, N12628, N3406, N67, N5215);
and AND3 (N12660, N12658, N10666, N152);
and AND2 (N12661, N12659, N8005);
nand NAND4 (N12662, N12648, N8061, N2543, N1025);
nand NAND2 (N12663, N12631, N11423);
xor XOR2 (N12664, N12656, N5543);
or OR2 (N12665, N12662, N4215);
and AND2 (N12666, N12645, N10240);
and AND3 (N12667, N12663, N6490, N8015);
and AND2 (N12668, N12660, N6573);
and AND2 (N12669, N12666, N12562);
buf BUF1 (N12670, N12661);
xor XOR2 (N12671, N12669, N6777);
xor XOR2 (N12672, N12657, N10818);
and AND2 (N12673, N12655, N10918);
xor XOR2 (N12674, N12672, N11132);
nand NAND3 (N12675, N12649, N1566, N12044);
not NOT1 (N12676, N12664);
nor NOR3 (N12677, N12667, N10049, N403);
buf BUF1 (N12678, N12670);
not NOT1 (N12679, N12665);
or OR3 (N12680, N12668, N5604, N11869);
nor NOR3 (N12681, N12680, N980, N2821);
xor XOR2 (N12682, N12652, N1531);
buf BUF1 (N12683, N12671);
xor XOR2 (N12684, N12682, N8589);
nor NOR4 (N12685, N12673, N8705, N2583, N8395);
nand NAND3 (N12686, N12685, N4724, N2636);
buf BUF1 (N12687, N12686);
not NOT1 (N12688, N12687);
or OR3 (N12689, N12683, N3188, N4390);
buf BUF1 (N12690, N12676);
buf BUF1 (N12691, N12674);
and AND4 (N12692, N12677, N8009, N3374, N7934);
or OR3 (N12693, N12690, N551, N7429);
buf BUF1 (N12694, N12692);
or OR2 (N12695, N12688, N7084);
xor XOR2 (N12696, N12691, N12341);
nand NAND3 (N12697, N12693, N11014, N11109);
nor NOR2 (N12698, N12697, N9311);
nand NAND4 (N12699, N12675, N9539, N5675, N7346);
or OR4 (N12700, N12695, N9833, N11721, N8117);
nor NOR2 (N12701, N12681, N5459);
xor XOR2 (N12702, N12684, N3287);
or OR2 (N12703, N12698, N10850);
nand NAND2 (N12704, N12702, N512);
nor NOR2 (N12705, N12678, N516);
nor NOR3 (N12706, N12701, N3452, N132);
and AND4 (N12707, N12703, N6525, N3622, N4912);
buf BUF1 (N12708, N12706);
xor XOR2 (N12709, N12705, N2260);
nor NOR2 (N12710, N12694, N8063);
xor XOR2 (N12711, N12689, N1071);
xor XOR2 (N12712, N12709, N9532);
buf BUF1 (N12713, N12704);
nor NOR2 (N12714, N12712, N9198);
xor XOR2 (N12715, N12711, N2470);
not NOT1 (N12716, N12679);
xor XOR2 (N12717, N12716, N9493);
buf BUF1 (N12718, N12715);
not NOT1 (N12719, N12707);
or OR3 (N12720, N12710, N10588, N1825);
nand NAND4 (N12721, N12699, N5860, N5607, N7341);
nand NAND3 (N12722, N12717, N2787, N7896);
xor XOR2 (N12723, N12696, N10359);
nor NOR4 (N12724, N12718, N6481, N12296, N8533);
buf BUF1 (N12725, N12719);
buf BUF1 (N12726, N12708);
xor XOR2 (N12727, N12726, N1798);
not NOT1 (N12728, N12723);
or OR3 (N12729, N12722, N5212, N681);
xor XOR2 (N12730, N12724, N4577);
nand NAND3 (N12731, N12727, N135, N8478);
nor NOR2 (N12732, N12730, N1076);
buf BUF1 (N12733, N12713);
and AND2 (N12734, N12720, N7759);
or OR4 (N12735, N12721, N1848, N88, N11530);
xor XOR2 (N12736, N12731, N4139);
or OR3 (N12737, N12728, N4965, N4228);
nand NAND3 (N12738, N12734, N7483, N2144);
nor NOR3 (N12739, N12725, N4025, N9828);
xor XOR2 (N12740, N12729, N10924);
not NOT1 (N12741, N12737);
nand NAND2 (N12742, N12700, N1696);
or OR3 (N12743, N12741, N3449, N12317);
or OR4 (N12744, N12736, N8721, N11748, N4377);
and AND3 (N12745, N12744, N8185, N4316);
and AND3 (N12746, N12733, N10955, N7802);
or OR3 (N12747, N12746, N11177, N8233);
xor XOR2 (N12748, N12742, N2726);
xor XOR2 (N12749, N12735, N29);
nor NOR4 (N12750, N12714, N7659, N974, N6222);
nand NAND3 (N12751, N12748, N10878, N12514);
xor XOR2 (N12752, N12743, N9859);
buf BUF1 (N12753, N12740);
or OR3 (N12754, N12745, N4720, N1245);
xor XOR2 (N12755, N12747, N9842);
nor NOR3 (N12756, N12750, N3935, N9653);
and AND3 (N12757, N12732, N5999, N11927);
not NOT1 (N12758, N12751);
xor XOR2 (N12759, N12739, N7801);
not NOT1 (N12760, N12757);
not NOT1 (N12761, N12755);
nor NOR2 (N12762, N12738, N9558);
nor NOR2 (N12763, N12760, N11857);
and AND4 (N12764, N12761, N2975, N11654, N8438);
nor NOR3 (N12765, N12764, N12705, N2061);
nor NOR3 (N12766, N12749, N3523, N11262);
nand NAND2 (N12767, N12765, N495);
buf BUF1 (N12768, N12766);
nand NAND2 (N12769, N12768, N4810);
xor XOR2 (N12770, N12759, N1491);
xor XOR2 (N12771, N12762, N1097);
nor NOR4 (N12772, N12756, N4254, N12375, N5808);
not NOT1 (N12773, N12763);
nor NOR4 (N12774, N12771, N9622, N11689, N12120);
and AND2 (N12775, N12752, N5225);
xor XOR2 (N12776, N12773, N2184);
or OR2 (N12777, N12770, N2196);
and AND4 (N12778, N12753, N6805, N20, N3835);
or OR4 (N12779, N12777, N3563, N11747, N3900);
not NOT1 (N12780, N12776);
buf BUF1 (N12781, N12758);
and AND4 (N12782, N12774, N12535, N9197, N2515);
not NOT1 (N12783, N12779);
not NOT1 (N12784, N12775);
nor NOR2 (N12785, N12767, N4990);
or OR4 (N12786, N12784, N10475, N4087, N7249);
and AND3 (N12787, N12769, N3413, N11394);
nand NAND4 (N12788, N12783, N6312, N2417, N4982);
xor XOR2 (N12789, N12786, N12188);
nand NAND4 (N12790, N12788, N8218, N9044, N10970);
or OR2 (N12791, N12781, N6480);
and AND3 (N12792, N12772, N11658, N5716);
xor XOR2 (N12793, N12778, N1004);
nor NOR2 (N12794, N12789, N2366);
and AND2 (N12795, N12787, N5920);
or OR4 (N12796, N12792, N9138, N10373, N4174);
or OR4 (N12797, N12754, N2939, N9819, N9182);
xor XOR2 (N12798, N12785, N12456);
not NOT1 (N12799, N12798);
xor XOR2 (N12800, N12796, N5684);
nand NAND4 (N12801, N12797, N1949, N1075, N11298);
nor NOR2 (N12802, N12801, N9614);
and AND3 (N12803, N12782, N8393, N5783);
nand NAND4 (N12804, N12793, N10901, N7018, N342);
xor XOR2 (N12805, N12804, N2345);
not NOT1 (N12806, N12780);
nand NAND3 (N12807, N12791, N3974, N1984);
buf BUF1 (N12808, N12790);
nand NAND4 (N12809, N12806, N652, N7339, N10199);
nor NOR4 (N12810, N12808, N12724, N3575, N629);
buf BUF1 (N12811, N12805);
buf BUF1 (N12812, N12809);
not NOT1 (N12813, N12812);
or OR4 (N12814, N12811, N10108, N12178, N8864);
buf BUF1 (N12815, N12800);
xor XOR2 (N12816, N12795, N7641);
or OR2 (N12817, N12807, N11896);
or OR3 (N12818, N12815, N4414, N12006);
nand NAND2 (N12819, N12814, N9093);
or OR3 (N12820, N12817, N8276, N11523);
xor XOR2 (N12821, N12803, N2367);
xor XOR2 (N12822, N12820, N5253);
buf BUF1 (N12823, N12816);
not NOT1 (N12824, N12802);
not NOT1 (N12825, N12799);
buf BUF1 (N12826, N12823);
buf BUF1 (N12827, N12821);
buf BUF1 (N12828, N12810);
buf BUF1 (N12829, N12813);
or OR4 (N12830, N12828, N2362, N7720, N1433);
or OR2 (N12831, N12829, N10650);
not NOT1 (N12832, N12827);
not NOT1 (N12833, N12794);
or OR2 (N12834, N12832, N5887);
nand NAND4 (N12835, N12824, N8868, N572, N10127);
or OR3 (N12836, N12826, N4443, N1035);
xor XOR2 (N12837, N12825, N7284);
buf BUF1 (N12838, N12834);
not NOT1 (N12839, N12835);
xor XOR2 (N12840, N12830, N4688);
buf BUF1 (N12841, N12838);
xor XOR2 (N12842, N12840, N8022);
nor NOR2 (N12843, N12819, N12550);
nand NAND4 (N12844, N12842, N5182, N1514, N7822);
not NOT1 (N12845, N12822);
buf BUF1 (N12846, N12844);
xor XOR2 (N12847, N12836, N8320);
not NOT1 (N12848, N12845);
nand NAND2 (N12849, N12837, N10063);
and AND2 (N12850, N12833, N1340);
xor XOR2 (N12851, N12839, N490);
xor XOR2 (N12852, N12851, N3257);
and AND2 (N12853, N12841, N4648);
or OR4 (N12854, N12843, N7942, N6347, N11953);
nor NOR3 (N12855, N12853, N3527, N3516);
and AND3 (N12856, N12848, N4219, N3253);
and AND2 (N12857, N12849, N3081);
and AND3 (N12858, N12854, N4848, N10720);
or OR2 (N12859, N12850, N12730);
not NOT1 (N12860, N12856);
nand NAND2 (N12861, N12831, N636);
not NOT1 (N12862, N12861);
xor XOR2 (N12863, N12847, N6036);
buf BUF1 (N12864, N12860);
or OR4 (N12865, N12846, N565, N8841, N4439);
nand NAND2 (N12866, N12857, N8254);
not NOT1 (N12867, N12863);
or OR4 (N12868, N12865, N11895, N6456, N4255);
not NOT1 (N12869, N12855);
and AND2 (N12870, N12866, N12435);
nor NOR2 (N12871, N12858, N10486);
xor XOR2 (N12872, N12852, N10550);
xor XOR2 (N12873, N12869, N9149);
or OR4 (N12874, N12872, N2122, N11432, N11093);
nand NAND4 (N12875, N12818, N3150, N9877, N2202);
xor XOR2 (N12876, N12875, N565);
buf BUF1 (N12877, N12862);
not NOT1 (N12878, N12859);
buf BUF1 (N12879, N12868);
not NOT1 (N12880, N12867);
nor NOR4 (N12881, N12874, N10212, N3494, N8989);
buf BUF1 (N12882, N12877);
or OR2 (N12883, N12871, N7498);
nand NAND4 (N12884, N12878, N3454, N7488, N1556);
and AND4 (N12885, N12873, N4455, N9620, N6940);
nor NOR2 (N12886, N12879, N550);
not NOT1 (N12887, N12883);
not NOT1 (N12888, N12885);
xor XOR2 (N12889, N12870, N1470);
or OR2 (N12890, N12881, N3275);
not NOT1 (N12891, N12890);
nand NAND2 (N12892, N12886, N1292);
nand NAND3 (N12893, N12892, N5373, N1249);
nand NAND2 (N12894, N12889, N9220);
buf BUF1 (N12895, N12893);
and AND4 (N12896, N12880, N3130, N12694, N1761);
xor XOR2 (N12897, N12891, N8058);
nor NOR4 (N12898, N12896, N7052, N2278, N4689);
buf BUF1 (N12899, N12888);
buf BUF1 (N12900, N12895);
nor NOR3 (N12901, N12887, N5903, N4771);
and AND3 (N12902, N12898, N9508, N4933);
and AND3 (N12903, N12884, N11597, N10922);
not NOT1 (N12904, N12876);
and AND2 (N12905, N12900, N643);
buf BUF1 (N12906, N12899);
buf BUF1 (N12907, N12905);
nor NOR4 (N12908, N12901, N1222, N2933, N9741);
and AND2 (N12909, N12894, N5195);
not NOT1 (N12910, N12864);
nor NOR3 (N12911, N12906, N226, N12864);
not NOT1 (N12912, N12903);
or OR2 (N12913, N12910, N8716);
and AND2 (N12914, N12909, N3170);
nand NAND2 (N12915, N12904, N3574);
xor XOR2 (N12916, N12897, N3966);
and AND3 (N12917, N12915, N6660, N11294);
or OR4 (N12918, N12908, N9945, N9796, N6986);
nand NAND3 (N12919, N12912, N2450, N9877);
buf BUF1 (N12920, N12911);
and AND4 (N12921, N12882, N5193, N5933, N12230);
or OR2 (N12922, N12907, N10664);
and AND3 (N12923, N12919, N5478, N8400);
or OR2 (N12924, N12921, N2265);
buf BUF1 (N12925, N12916);
nor NOR3 (N12926, N12917, N8479, N4927);
xor XOR2 (N12927, N12918, N11559);
buf BUF1 (N12928, N12913);
not NOT1 (N12929, N12924);
and AND3 (N12930, N12922, N5631, N5521);
or OR2 (N12931, N12923, N6995);
and AND3 (N12932, N12927, N476, N9834);
or OR2 (N12933, N12925, N1432);
nand NAND2 (N12934, N12932, N10446);
xor XOR2 (N12935, N12930, N959);
buf BUF1 (N12936, N12933);
nor NOR4 (N12937, N12902, N10219, N2950, N3541);
nand NAND4 (N12938, N12914, N5467, N6126, N9014);
xor XOR2 (N12939, N12936, N3808);
nand NAND3 (N12940, N12931, N12870, N12421);
nor NOR4 (N12941, N12939, N8554, N10225, N11392);
or OR2 (N12942, N12920, N8251);
or OR2 (N12943, N12929, N11072);
nand NAND2 (N12944, N12942, N8821);
or OR2 (N12945, N12940, N1923);
buf BUF1 (N12946, N12945);
xor XOR2 (N12947, N12944, N7153);
or OR3 (N12948, N12943, N9694, N10046);
and AND4 (N12949, N12941, N8561, N12056, N3173);
xor XOR2 (N12950, N12938, N9379);
nand NAND3 (N12951, N12934, N7419, N7750);
nor NOR4 (N12952, N12926, N9843, N5228, N3771);
nor NOR3 (N12953, N12937, N2282, N9535);
not NOT1 (N12954, N12935);
nand NAND4 (N12955, N12947, N9470, N1907, N2604);
buf BUF1 (N12956, N12949);
buf BUF1 (N12957, N12928);
nor NOR4 (N12958, N12957, N10562, N11598, N4751);
nor NOR3 (N12959, N12948, N10245, N8092);
not NOT1 (N12960, N12959);
and AND3 (N12961, N12958, N7580, N3482);
and AND4 (N12962, N12951, N1298, N12275, N8291);
not NOT1 (N12963, N12950);
buf BUF1 (N12964, N12953);
nor NOR4 (N12965, N12955, N11440, N4450, N10079);
not NOT1 (N12966, N12961);
nand NAND3 (N12967, N12965, N680, N1377);
and AND4 (N12968, N12967, N3335, N4580, N1314);
nor NOR2 (N12969, N12952, N12092);
nor NOR2 (N12970, N12956, N3493);
xor XOR2 (N12971, N12968, N9500);
and AND3 (N12972, N12971, N6857, N5183);
not NOT1 (N12973, N12972);
buf BUF1 (N12974, N12969);
not NOT1 (N12975, N12963);
or OR3 (N12976, N12964, N7977, N3355);
or OR2 (N12977, N12946, N3190);
or OR2 (N12978, N12973, N464);
nor NOR2 (N12979, N12970, N8365);
not NOT1 (N12980, N12979);
nor NOR2 (N12981, N12977, N7246);
and AND4 (N12982, N12966, N6650, N12749, N9494);
xor XOR2 (N12983, N12975, N1712);
or OR2 (N12984, N12974, N4448);
nand NAND4 (N12985, N12982, N2236, N6102, N9248);
xor XOR2 (N12986, N12984, N5673);
buf BUF1 (N12987, N12962);
or OR3 (N12988, N12960, N10401, N12796);
xor XOR2 (N12989, N12987, N4295);
xor XOR2 (N12990, N12954, N4746);
xor XOR2 (N12991, N12981, N7817);
not NOT1 (N12992, N12988);
not NOT1 (N12993, N12990);
not NOT1 (N12994, N12976);
or OR3 (N12995, N12986, N791, N12003);
not NOT1 (N12996, N12995);
nand NAND4 (N12997, N12993, N9851, N5179, N9717);
xor XOR2 (N12998, N12994, N11816);
nor NOR4 (N12999, N12991, N244, N12733, N10979);
nand NAND3 (N13000, N12996, N5790, N11996);
not NOT1 (N13001, N12983);
nor NOR2 (N13002, N12989, N9079);
nand NAND2 (N13003, N12978, N10250);
xor XOR2 (N13004, N12985, N12868);
nor NOR2 (N13005, N12992, N1711);
and AND4 (N13006, N12999, N12158, N3812, N11598);
xor XOR2 (N13007, N13003, N1439);
not NOT1 (N13008, N13007);
not NOT1 (N13009, N13005);
nand NAND2 (N13010, N13006, N1427);
xor XOR2 (N13011, N12980, N9703);
and AND2 (N13012, N13009, N4843);
nand NAND2 (N13013, N13012, N573);
and AND3 (N13014, N12997, N4858, N12633);
and AND3 (N13015, N13011, N7071, N1317);
xor XOR2 (N13016, N13004, N12952);
nand NAND4 (N13017, N13015, N2981, N6573, N10894);
and AND4 (N13018, N13002, N7942, N10498, N1259);
nor NOR2 (N13019, N13018, N10071);
xor XOR2 (N13020, N12998, N6725);
nand NAND3 (N13021, N13020, N11807, N2868);
nand NAND4 (N13022, N13008, N4267, N8148, N1404);
and AND4 (N13023, N13016, N10799, N10289, N105);
and AND3 (N13024, N13019, N2431, N9637);
nand NAND4 (N13025, N13024, N8682, N10606, N2090);
and AND4 (N13026, N13017, N10348, N6397, N10757);
not NOT1 (N13027, N13013);
nor NOR4 (N13028, N13022, N7209, N4098, N2326);
and AND3 (N13029, N13014, N8145, N2525);
buf BUF1 (N13030, N13028);
xor XOR2 (N13031, N13023, N1021);
and AND4 (N13032, N13027, N2520, N8619, N6128);
nand NAND4 (N13033, N13010, N10177, N2203, N7264);
or OR4 (N13034, N13001, N2413, N8741, N7867);
nor NOR2 (N13035, N13029, N3370);
not NOT1 (N13036, N13031);
or OR2 (N13037, N13036, N12249);
buf BUF1 (N13038, N13037);
or OR2 (N13039, N13025, N2792);
nor NOR2 (N13040, N13034, N8113);
and AND4 (N13041, N13026, N11424, N7853, N9992);
nor NOR3 (N13042, N13030, N828, N911);
buf BUF1 (N13043, N13041);
xor XOR2 (N13044, N13000, N3143);
and AND4 (N13045, N13040, N1175, N4821, N940);
nor NOR2 (N13046, N13045, N10196);
nor NOR3 (N13047, N13043, N1230, N7988);
xor XOR2 (N13048, N13021, N10503);
buf BUF1 (N13049, N13039);
and AND3 (N13050, N13046, N7312, N7650);
nand NAND3 (N13051, N13033, N11274, N12974);
or OR3 (N13052, N13035, N12065, N1765);
nand NAND3 (N13053, N13048, N6151, N3596);
xor XOR2 (N13054, N13047, N9186);
nand NAND4 (N13055, N13052, N9072, N11792, N4388);
nand NAND4 (N13056, N13051, N4760, N8686, N6010);
nor NOR3 (N13057, N13042, N8089, N4586);
nand NAND3 (N13058, N13056, N2912, N6029);
nor NOR2 (N13059, N13058, N2657);
and AND4 (N13060, N13044, N5256, N1411, N3792);
nor NOR2 (N13061, N13049, N3259);
buf BUF1 (N13062, N13038);
or OR2 (N13063, N13061, N7254);
and AND2 (N13064, N13062, N4718);
xor XOR2 (N13065, N13032, N11404);
xor XOR2 (N13066, N13065, N9638);
nor NOR3 (N13067, N13050, N5313, N931);
or OR2 (N13068, N13055, N4003);
buf BUF1 (N13069, N13067);
xor XOR2 (N13070, N13066, N3082);
or OR2 (N13071, N13070, N4876);
xor XOR2 (N13072, N13069, N9733);
nand NAND3 (N13073, N13068, N5634, N1273);
nor NOR2 (N13074, N13072, N935);
or OR3 (N13075, N13071, N10552, N9454);
and AND4 (N13076, N13074, N2649, N4397, N7452);
xor XOR2 (N13077, N13054, N11148);
buf BUF1 (N13078, N13060);
not NOT1 (N13079, N13064);
xor XOR2 (N13080, N13079, N6782);
and AND2 (N13081, N13077, N11857);
nor NOR4 (N13082, N13073, N280, N12580, N2754);
buf BUF1 (N13083, N13081);
or OR4 (N13084, N13053, N6343, N938, N9496);
not NOT1 (N13085, N13057);
and AND2 (N13086, N13080, N12838);
or OR3 (N13087, N13075, N4424, N9689);
nor NOR3 (N13088, N13063, N3577, N11509);
and AND2 (N13089, N13084, N11734);
or OR2 (N13090, N13082, N3541);
or OR4 (N13091, N13085, N10613, N6765, N2137);
xor XOR2 (N13092, N13059, N1931);
or OR4 (N13093, N13089, N12555, N5191, N4825);
xor XOR2 (N13094, N13083, N6168);
and AND3 (N13095, N13094, N11282, N4609);
or OR2 (N13096, N13087, N2420);
nand NAND4 (N13097, N13086, N374, N3523, N5553);
or OR2 (N13098, N13078, N7525);
not NOT1 (N13099, N13076);
and AND2 (N13100, N13090, N2745);
not NOT1 (N13101, N13091);
and AND2 (N13102, N13095, N9727);
buf BUF1 (N13103, N13099);
nor NOR2 (N13104, N13088, N3274);
or OR4 (N13105, N13093, N9543, N6552, N10734);
not NOT1 (N13106, N13105);
not NOT1 (N13107, N13092);
nor NOR2 (N13108, N13097, N10791);
or OR4 (N13109, N13103, N5511, N1802, N1068);
nor NOR3 (N13110, N13101, N12295, N9638);
nand NAND3 (N13111, N13100, N6291, N11327);
or OR2 (N13112, N13107, N3626);
or OR4 (N13113, N13096, N149, N1415, N9423);
nor NOR3 (N13114, N13108, N9807, N7855);
or OR4 (N13115, N13114, N1224, N5370, N9427);
buf BUF1 (N13116, N13113);
or OR2 (N13117, N13112, N10823);
buf BUF1 (N13118, N13098);
and AND3 (N13119, N13104, N110, N3423);
nor NOR2 (N13120, N13116, N10016);
not NOT1 (N13121, N13111);
nor NOR3 (N13122, N13117, N12528, N10500);
and AND4 (N13123, N13122, N1010, N7529, N992);
not NOT1 (N13124, N13120);
buf BUF1 (N13125, N13123);
or OR4 (N13126, N13109, N7638, N3612, N4611);
xor XOR2 (N13127, N13126, N5415);
buf BUF1 (N13128, N13124);
and AND2 (N13129, N13121, N3082);
or OR2 (N13130, N13129, N5873);
nor NOR4 (N13131, N13125, N10372, N10047, N10253);
not NOT1 (N13132, N13102);
nor NOR3 (N13133, N13115, N7957, N6637);
not NOT1 (N13134, N13119);
not NOT1 (N13135, N13127);
nor NOR3 (N13136, N13132, N11435, N8537);
or OR3 (N13137, N13110, N9259, N3490);
or OR4 (N13138, N13106, N10372, N10544, N5017);
and AND3 (N13139, N13135, N9595, N3138);
not NOT1 (N13140, N13138);
nor NOR4 (N13141, N13128, N10610, N5301, N3548);
and AND3 (N13142, N13141, N5, N5265);
xor XOR2 (N13143, N13136, N6871);
xor XOR2 (N13144, N13130, N12550);
and AND4 (N13145, N13144, N11011, N12831, N5046);
or OR4 (N13146, N13137, N6314, N11490, N10816);
nand NAND2 (N13147, N13139, N6445);
and AND4 (N13148, N13118, N10885, N9942, N2885);
and AND2 (N13149, N13140, N5049);
and AND2 (N13150, N13133, N9239);
nand NAND3 (N13151, N13134, N5599, N9477);
nor NOR2 (N13152, N13149, N2347);
buf BUF1 (N13153, N13152);
or OR3 (N13154, N13131, N1192, N403);
xor XOR2 (N13155, N13153, N4550);
and AND2 (N13156, N13146, N8097);
buf BUF1 (N13157, N13148);
nor NOR3 (N13158, N13147, N5860, N2233);
xor XOR2 (N13159, N13157, N5494);
nand NAND3 (N13160, N13155, N8385, N5586);
and AND2 (N13161, N13151, N7271);
or OR3 (N13162, N13142, N8678, N5925);
and AND2 (N13163, N13159, N10570);
xor XOR2 (N13164, N13150, N10608);
buf BUF1 (N13165, N13145);
nand NAND3 (N13166, N13160, N4671, N10001);
or OR4 (N13167, N13143, N5935, N9217, N7095);
nand NAND2 (N13168, N13164, N4776);
or OR2 (N13169, N13167, N8387);
and AND3 (N13170, N13161, N10387, N12313);
and AND3 (N13171, N13162, N5064, N9683);
nand NAND3 (N13172, N13158, N6266, N10180);
and AND2 (N13173, N13166, N4105);
and AND2 (N13174, N13154, N3333);
buf BUF1 (N13175, N13165);
and AND3 (N13176, N13168, N7204, N199);
buf BUF1 (N13177, N13174);
buf BUF1 (N13178, N13156);
or OR2 (N13179, N13176, N5043);
and AND2 (N13180, N13169, N5753);
nor NOR4 (N13181, N13179, N9843, N5913, N12751);
xor XOR2 (N13182, N13175, N4343);
and AND2 (N13183, N13170, N8266);
nor NOR2 (N13184, N13180, N12984);
nor NOR2 (N13185, N13172, N7589);
buf BUF1 (N13186, N13177);
not NOT1 (N13187, N13171);
or OR2 (N13188, N13181, N10209);
nand NAND2 (N13189, N13184, N648);
buf BUF1 (N13190, N13182);
nand NAND3 (N13191, N13183, N8263, N6291);
xor XOR2 (N13192, N13186, N2366);
nor NOR2 (N13193, N13185, N4355);
or OR2 (N13194, N13193, N2801);
nand NAND4 (N13195, N13163, N8559, N7076, N2765);
not NOT1 (N13196, N13194);
or OR2 (N13197, N13192, N11752);
not NOT1 (N13198, N13187);
xor XOR2 (N13199, N13191, N4343);
not NOT1 (N13200, N13199);
nand NAND3 (N13201, N13197, N7124, N284);
nand NAND2 (N13202, N13195, N9154);
nand NAND2 (N13203, N13198, N12970);
nand NAND4 (N13204, N13188, N8075, N4143, N8200);
nand NAND2 (N13205, N13200, N5280);
or OR4 (N13206, N13201, N5066, N9856, N6289);
nor NOR4 (N13207, N13196, N6630, N12208, N5441);
or OR3 (N13208, N13189, N7928, N8257);
buf BUF1 (N13209, N13205);
not NOT1 (N13210, N13190);
buf BUF1 (N13211, N13178);
xor XOR2 (N13212, N13202, N11366);
xor XOR2 (N13213, N13203, N4817);
nand NAND2 (N13214, N13207, N7687);
buf BUF1 (N13215, N13173);
nand NAND2 (N13216, N13208, N7789);
nor NOR4 (N13217, N13216, N4741, N6543, N10379);
and AND4 (N13218, N13214, N9935, N5764, N7695);
buf BUF1 (N13219, N13212);
buf BUF1 (N13220, N13206);
not NOT1 (N13221, N13211);
nor NOR3 (N13222, N13221, N6973, N8732);
nor NOR4 (N13223, N13222, N4360, N8678, N8707);
or OR2 (N13224, N13220, N8843);
xor XOR2 (N13225, N13209, N7014);
or OR2 (N13226, N13217, N10076);
nand NAND2 (N13227, N13215, N1009);
nand NAND2 (N13228, N13227, N4860);
nand NAND4 (N13229, N13204, N2330, N11018, N4617);
buf BUF1 (N13230, N13223);
nor NOR4 (N13231, N13224, N8542, N9418, N4002);
and AND4 (N13232, N13229, N8664, N3945, N983);
and AND3 (N13233, N13230, N781, N5604);
nand NAND4 (N13234, N13228, N4091, N521, N1931);
nand NAND3 (N13235, N13210, N201, N604);
buf BUF1 (N13236, N13226);
or OR4 (N13237, N13236, N3728, N7801, N786);
not NOT1 (N13238, N13234);
and AND3 (N13239, N13231, N5948, N936);
and AND2 (N13240, N13235, N12758);
xor XOR2 (N13241, N13219, N306);
xor XOR2 (N13242, N13225, N6062);
nand NAND4 (N13243, N13233, N2861, N11277, N4404);
buf BUF1 (N13244, N13218);
buf BUF1 (N13245, N13239);
and AND2 (N13246, N13245, N4057);
buf BUF1 (N13247, N13241);
and AND3 (N13248, N13242, N2794, N11079);
xor XOR2 (N13249, N13248, N2352);
not NOT1 (N13250, N13232);
nor NOR4 (N13251, N13243, N9603, N7106, N7379);
buf BUF1 (N13252, N13244);
nor NOR2 (N13253, N13237, N9180);
buf BUF1 (N13254, N13253);
or OR3 (N13255, N13240, N4337, N11626);
xor XOR2 (N13256, N13254, N8109);
and AND3 (N13257, N13249, N1442, N1876);
or OR2 (N13258, N13251, N6571);
nor NOR4 (N13259, N13213, N10196, N9134, N6404);
nor NOR3 (N13260, N13247, N6696, N7167);
nand NAND4 (N13261, N13246, N7620, N4341, N13012);
nor NOR4 (N13262, N13257, N12601, N8780, N786);
not NOT1 (N13263, N13262);
or OR4 (N13264, N13263, N10972, N1222, N5554);
and AND2 (N13265, N13258, N8441);
xor XOR2 (N13266, N13259, N627);
or OR3 (N13267, N13260, N2223, N9099);
or OR3 (N13268, N13252, N9504, N12812);
or OR4 (N13269, N13256, N1860, N5184, N2760);
buf BUF1 (N13270, N13238);
and AND4 (N13271, N13265, N135, N221, N6798);
xor XOR2 (N13272, N13271, N11111);
or OR3 (N13273, N13261, N8644, N608);
not NOT1 (N13274, N13255);
or OR4 (N13275, N13268, N1601, N13274, N4406);
not NOT1 (N13276, N8156);
not NOT1 (N13277, N13250);
nand NAND3 (N13278, N13267, N9826, N12624);
nand NAND3 (N13279, N13273, N7396, N4086);
nand NAND2 (N13280, N13264, N1520);
and AND3 (N13281, N13269, N10211, N9738);
xor XOR2 (N13282, N13278, N4452);
xor XOR2 (N13283, N13272, N9686);
nand NAND3 (N13284, N13277, N12224, N6365);
buf BUF1 (N13285, N13266);
nor NOR2 (N13286, N13276, N6131);
and AND2 (N13287, N13280, N1069);
buf BUF1 (N13288, N13286);
and AND2 (N13289, N13287, N7402);
nand NAND2 (N13290, N13285, N4084);
and AND4 (N13291, N13282, N11395, N8208, N1932);
nand NAND4 (N13292, N13284, N4073, N8274, N7015);
nor NOR2 (N13293, N13289, N12093);
xor XOR2 (N13294, N13291, N1011);
xor XOR2 (N13295, N13288, N1258);
nand NAND2 (N13296, N13290, N13054);
buf BUF1 (N13297, N13294);
or OR2 (N13298, N13283, N6077);
nand NAND3 (N13299, N13297, N2401, N5656);
not NOT1 (N13300, N13296);
nor NOR3 (N13301, N13295, N5467, N10206);
xor XOR2 (N13302, N13298, N3487);
nand NAND3 (N13303, N13300, N10987, N8454);
or OR3 (N13304, N13299, N5661, N9127);
and AND3 (N13305, N13301, N1006, N2717);
buf BUF1 (N13306, N13292);
nand NAND4 (N13307, N13279, N11440, N3329, N10887);
nand NAND2 (N13308, N13275, N476);
nor NOR2 (N13309, N13281, N5868);
nand NAND3 (N13310, N13309, N7273, N4676);
nor NOR2 (N13311, N13303, N4682);
nand NAND2 (N13312, N13293, N9702);
and AND2 (N13313, N13270, N3103);
xor XOR2 (N13314, N13306, N8213);
not NOT1 (N13315, N13314);
nor NOR2 (N13316, N13310, N11598);
xor XOR2 (N13317, N13315, N5606);
not NOT1 (N13318, N13316);
not NOT1 (N13319, N13308);
buf BUF1 (N13320, N13305);
xor XOR2 (N13321, N13320, N10974);
not NOT1 (N13322, N13302);
nand NAND2 (N13323, N13321, N8147);
or OR4 (N13324, N13318, N10884, N11831, N12248);
xor XOR2 (N13325, N13313, N11570);
nor NOR4 (N13326, N13324, N11193, N1057, N91);
nand NAND2 (N13327, N13311, N7359);
buf BUF1 (N13328, N13319);
buf BUF1 (N13329, N13317);
nor NOR2 (N13330, N13327, N10920);
nand NAND3 (N13331, N13307, N6489, N716);
or OR3 (N13332, N13323, N5004, N8941);
buf BUF1 (N13333, N13304);
xor XOR2 (N13334, N13312, N5876);
and AND4 (N13335, N13330, N6712, N5800, N10245);
xor XOR2 (N13336, N13331, N4940);
nor NOR4 (N13337, N13329, N9331, N6983, N95);
or OR3 (N13338, N13336, N2967, N9068);
not NOT1 (N13339, N13326);
nor NOR4 (N13340, N13337, N11625, N966, N2430);
nor NOR2 (N13341, N13328, N12414);
buf BUF1 (N13342, N13339);
xor XOR2 (N13343, N13342, N2510);
and AND3 (N13344, N13322, N12445, N1196);
nor NOR2 (N13345, N13338, N4794);
xor XOR2 (N13346, N13325, N2202);
buf BUF1 (N13347, N13343);
not NOT1 (N13348, N13340);
buf BUF1 (N13349, N13341);
xor XOR2 (N13350, N13348, N10375);
nand NAND3 (N13351, N13333, N104, N9159);
nor NOR2 (N13352, N13351, N12115);
xor XOR2 (N13353, N13344, N5899);
xor XOR2 (N13354, N13346, N9424);
nor NOR3 (N13355, N13345, N9593, N5234);
xor XOR2 (N13356, N13355, N960);
or OR2 (N13357, N13353, N10456);
nor NOR4 (N13358, N13347, N7542, N700, N12229);
and AND3 (N13359, N13358, N7717, N6103);
nand NAND3 (N13360, N13356, N7257, N8289);
not NOT1 (N13361, N13360);
nand NAND2 (N13362, N13354, N6651);
not NOT1 (N13363, N13350);
xor XOR2 (N13364, N13352, N978);
nor NOR4 (N13365, N13349, N2802, N7768, N11247);
xor XOR2 (N13366, N13361, N5319);
or OR3 (N13367, N13366, N6831, N680);
buf BUF1 (N13368, N13367);
and AND4 (N13369, N13362, N12553, N5233, N10408);
nor NOR2 (N13370, N13332, N7336);
nand NAND4 (N13371, N13363, N9710, N6312, N775);
and AND3 (N13372, N13371, N11255, N3140);
nor NOR3 (N13373, N13357, N7274, N1400);
not NOT1 (N13374, N13372);
xor XOR2 (N13375, N13335, N6593);
not NOT1 (N13376, N13370);
and AND2 (N13377, N13375, N8197);
nand NAND4 (N13378, N13373, N12272, N11655, N8646);
nor NOR3 (N13379, N13368, N1376, N1606);
and AND2 (N13380, N13374, N7269);
or OR2 (N13381, N13380, N802);
not NOT1 (N13382, N13359);
and AND3 (N13383, N13334, N7273, N6454);
buf BUF1 (N13384, N13364);
not NOT1 (N13385, N13381);
xor XOR2 (N13386, N13385, N1689);
buf BUF1 (N13387, N13376);
nor NOR3 (N13388, N13378, N13081, N9639);
nand NAND4 (N13389, N13382, N7685, N10289, N12099);
and AND3 (N13390, N13377, N13259, N9012);
or OR4 (N13391, N13389, N4992, N8427, N5769);
nor NOR3 (N13392, N13384, N12387, N1438);
not NOT1 (N13393, N13386);
or OR2 (N13394, N13391, N7304);
or OR2 (N13395, N13369, N6687);
or OR3 (N13396, N13395, N389, N6539);
buf BUF1 (N13397, N13365);
not NOT1 (N13398, N13388);
not NOT1 (N13399, N13393);
and AND4 (N13400, N13398, N10900, N1627, N10915);
xor XOR2 (N13401, N13397, N11464);
not NOT1 (N13402, N13401);
buf BUF1 (N13403, N13396);
not NOT1 (N13404, N13399);
nand NAND3 (N13405, N13404, N2185, N752);
and AND2 (N13406, N13403, N4762);
and AND3 (N13407, N13394, N11182, N12430);
nand NAND2 (N13408, N13379, N8849);
nand NAND2 (N13409, N13405, N5592);
buf BUF1 (N13410, N13402);
buf BUF1 (N13411, N13407);
nand NAND3 (N13412, N13408, N691, N5646);
nand NAND3 (N13413, N13411, N12016, N10931);
nor NOR3 (N13414, N13392, N1249, N7987);
not NOT1 (N13415, N13409);
nor NOR4 (N13416, N13390, N6469, N10890, N684);
or OR4 (N13417, N13413, N1277, N10460, N2322);
nor NOR2 (N13418, N13412, N11003);
xor XOR2 (N13419, N13406, N9122);
nor NOR2 (N13420, N13419, N5161);
and AND2 (N13421, N13415, N7989);
and AND3 (N13422, N13416, N7171, N11589);
nand NAND3 (N13423, N13420, N2230, N9912);
or OR4 (N13424, N13422, N12382, N5451, N4990);
buf BUF1 (N13425, N13418);
nand NAND4 (N13426, N13423, N11626, N11232, N9879);
not NOT1 (N13427, N13400);
xor XOR2 (N13428, N13414, N4920);
nand NAND3 (N13429, N13425, N928, N11831);
nand NAND4 (N13430, N13421, N10253, N1766, N2886);
or OR2 (N13431, N13383, N11106);
xor XOR2 (N13432, N13429, N276);
and AND3 (N13433, N13427, N4604, N4086);
xor XOR2 (N13434, N13433, N8191);
not NOT1 (N13435, N13387);
xor XOR2 (N13436, N13426, N2562);
and AND3 (N13437, N13410, N13016, N5888);
xor XOR2 (N13438, N13430, N9978);
or OR4 (N13439, N13434, N4623, N1114, N629);
nand NAND2 (N13440, N13432, N2719);
buf BUF1 (N13441, N13437);
xor XOR2 (N13442, N13428, N4107);
xor XOR2 (N13443, N13436, N2376);
nor NOR3 (N13444, N13417, N2066, N3413);
or OR4 (N13445, N13431, N874, N7060, N3442);
and AND3 (N13446, N13435, N1387, N9681);
not NOT1 (N13447, N13446);
xor XOR2 (N13448, N13441, N4867);
not NOT1 (N13449, N13442);
xor XOR2 (N13450, N13445, N5639);
or OR3 (N13451, N13449, N4892, N335);
and AND2 (N13452, N13443, N1396);
nand NAND4 (N13453, N13444, N9559, N9237, N8913);
and AND3 (N13454, N13448, N9760, N1428);
nor NOR2 (N13455, N13451, N6686);
buf BUF1 (N13456, N13440);
nand NAND2 (N13457, N13439, N4182);
nor NOR4 (N13458, N13453, N2560, N1323, N7647);
nor NOR2 (N13459, N13454, N235);
xor XOR2 (N13460, N13450, N12479);
not NOT1 (N13461, N13457);
and AND3 (N13462, N13456, N118, N1712);
and AND4 (N13463, N13452, N7441, N5071, N9148);
xor XOR2 (N13464, N13459, N11897);
xor XOR2 (N13465, N13424, N13403);
xor XOR2 (N13466, N13458, N11131);
xor XOR2 (N13467, N13462, N8019);
or OR2 (N13468, N13455, N1395);
or OR2 (N13469, N13461, N11520);
buf BUF1 (N13470, N13447);
or OR3 (N13471, N13465, N2376, N1877);
xor XOR2 (N13472, N13464, N4038);
xor XOR2 (N13473, N13460, N9335);
and AND4 (N13474, N13472, N8836, N9433, N10126);
or OR2 (N13475, N13438, N9840);
and AND4 (N13476, N13474, N12948, N787, N771);
nor NOR4 (N13477, N13468, N3072, N1791, N11226);
nand NAND3 (N13478, N13476, N9571, N11209);
not NOT1 (N13479, N13478);
or OR3 (N13480, N13466, N10232, N545);
and AND4 (N13481, N13480, N6968, N5594, N13070);
not NOT1 (N13482, N13479);
nor NOR2 (N13483, N13477, N6655);
buf BUF1 (N13484, N13482);
buf BUF1 (N13485, N13484);
buf BUF1 (N13486, N13483);
buf BUF1 (N13487, N13485);
not NOT1 (N13488, N13475);
and AND4 (N13489, N13473, N6439, N9933, N4455);
and AND4 (N13490, N13467, N1264, N1117, N9634);
and AND3 (N13491, N13489, N1162, N10450);
xor XOR2 (N13492, N13486, N11900);
buf BUF1 (N13493, N13490);
and AND3 (N13494, N13487, N10647, N2371);
nor NOR4 (N13495, N13492, N6272, N4422, N1623);
and AND3 (N13496, N13493, N2662, N4160);
buf BUF1 (N13497, N13463);
nand NAND4 (N13498, N13481, N8682, N4493, N12646);
and AND3 (N13499, N13495, N1168, N5995);
nor NOR4 (N13500, N13499, N5206, N5518, N6463);
and AND2 (N13501, N13471, N7673);
nand NAND3 (N13502, N13496, N8431, N13012);
xor XOR2 (N13503, N13500, N3008);
nor NOR2 (N13504, N13503, N9803);
not NOT1 (N13505, N13469);
or OR2 (N13506, N13470, N10596);
nor NOR3 (N13507, N13497, N4331, N747);
buf BUF1 (N13508, N13498);
nor NOR4 (N13509, N13501, N8572, N12906, N6698);
and AND4 (N13510, N13504, N5703, N3928, N9574);
nand NAND4 (N13511, N13508, N13407, N10575, N9690);
and AND2 (N13512, N13509, N5432);
nand NAND4 (N13513, N13491, N4766, N10878, N5221);
not NOT1 (N13514, N13511);
and AND3 (N13515, N13488, N4559, N8204);
nand NAND2 (N13516, N13513, N7468);
nor NOR2 (N13517, N13515, N2990);
buf BUF1 (N13518, N13494);
and AND3 (N13519, N13506, N4903, N839);
or OR3 (N13520, N13507, N12998, N6315);
nand NAND2 (N13521, N13514, N7010);
buf BUF1 (N13522, N13505);
xor XOR2 (N13523, N13510, N8862);
nand NAND4 (N13524, N13523, N788, N7895, N2719);
xor XOR2 (N13525, N13502, N4543);
or OR4 (N13526, N13512, N2007, N12488, N2065);
nand NAND2 (N13527, N13520, N9734);
nand NAND3 (N13528, N13526, N5555, N8617);
nand NAND2 (N13529, N13516, N6045);
and AND3 (N13530, N13521, N1466, N3199);
and AND2 (N13531, N13528, N9842);
buf BUF1 (N13532, N13524);
nor NOR2 (N13533, N13525, N13033);
and AND3 (N13534, N13530, N1146, N1627);
nand NAND3 (N13535, N13519, N12684, N9904);
or OR2 (N13536, N13532, N2833);
and AND3 (N13537, N13522, N3131, N5222);
and AND4 (N13538, N13531, N12151, N9084, N2946);
xor XOR2 (N13539, N13529, N8292);
not NOT1 (N13540, N13539);
or OR2 (N13541, N13518, N10175);
nand NAND2 (N13542, N13527, N1931);
buf BUF1 (N13543, N13534);
buf BUF1 (N13544, N13538);
xor XOR2 (N13545, N13537, N11276);
and AND3 (N13546, N13544, N3841, N9211);
xor XOR2 (N13547, N13533, N8017);
or OR4 (N13548, N13536, N12721, N2935, N5839);
not NOT1 (N13549, N13535);
not NOT1 (N13550, N13542);
nor NOR3 (N13551, N13517, N6986, N11521);
or OR4 (N13552, N13548, N3894, N10766, N9659);
xor XOR2 (N13553, N13547, N6839);
xor XOR2 (N13554, N13550, N10018);
or OR4 (N13555, N13540, N9060, N9686, N5404);
nor NOR2 (N13556, N13545, N5304);
nor NOR2 (N13557, N13541, N8928);
not NOT1 (N13558, N13556);
buf BUF1 (N13559, N13549);
not NOT1 (N13560, N13554);
xor XOR2 (N13561, N13560, N6622);
xor XOR2 (N13562, N13552, N10300);
and AND4 (N13563, N13562, N8758, N7067, N4771);
nand NAND3 (N13564, N13546, N10077, N11692);
nand NAND2 (N13565, N13561, N5995);
nand NAND2 (N13566, N13557, N602);
nor NOR2 (N13567, N13543, N12855);
buf BUF1 (N13568, N13553);
or OR3 (N13569, N13567, N24, N9955);
or OR4 (N13570, N13555, N13536, N12557, N10145);
nand NAND3 (N13571, N13568, N8624, N1701);
nand NAND4 (N13572, N13570, N1671, N4858, N10355);
not NOT1 (N13573, N13564);
not NOT1 (N13574, N13558);
or OR3 (N13575, N13565, N4310, N4309);
not NOT1 (N13576, N13575);
buf BUF1 (N13577, N13563);
nand NAND4 (N13578, N13576, N8819, N10796, N7225);
not NOT1 (N13579, N13577);
xor XOR2 (N13580, N13571, N6027);
and AND4 (N13581, N13566, N7739, N5625, N11885);
not NOT1 (N13582, N13559);
nor NOR2 (N13583, N13551, N12192);
nand NAND2 (N13584, N13578, N10307);
not NOT1 (N13585, N13569);
and AND2 (N13586, N13581, N1362);
not NOT1 (N13587, N13572);
xor XOR2 (N13588, N13579, N1871);
buf BUF1 (N13589, N13574);
nor NOR2 (N13590, N13585, N6554);
xor XOR2 (N13591, N13589, N2180);
and AND4 (N13592, N13586, N4961, N8416, N960);
and AND2 (N13593, N13590, N10859);
not NOT1 (N13594, N13584);
buf BUF1 (N13595, N13591);
not NOT1 (N13596, N13580);
buf BUF1 (N13597, N13596);
xor XOR2 (N13598, N13592, N173);
not NOT1 (N13599, N13594);
or OR3 (N13600, N13599, N4205, N7743);
xor XOR2 (N13601, N13587, N1730);
or OR2 (N13602, N13573, N10351);
not NOT1 (N13603, N13602);
and AND3 (N13604, N13595, N12882, N3423);
xor XOR2 (N13605, N13597, N4155);
or OR4 (N13606, N13588, N5752, N9589, N1164);
nor NOR4 (N13607, N13582, N6041, N12257, N2079);
and AND4 (N13608, N13603, N10389, N6456, N4597);
and AND3 (N13609, N13608, N7239, N3491);
nor NOR3 (N13610, N13593, N566, N10636);
or OR2 (N13611, N13610, N74);
nor NOR2 (N13612, N13611, N6516);
nand NAND2 (N13613, N13606, N9985);
not NOT1 (N13614, N13607);
xor XOR2 (N13615, N13583, N9628);
not NOT1 (N13616, N13614);
xor XOR2 (N13617, N13615, N12572);
nand NAND2 (N13618, N13604, N1843);
nand NAND4 (N13619, N13601, N5252, N12887, N380);
or OR2 (N13620, N13612, N10764);
nor NOR2 (N13621, N13609, N5660);
not NOT1 (N13622, N13605);
or OR4 (N13623, N13617, N2870, N12380, N7642);
nor NOR4 (N13624, N13620, N12599, N9347, N1718);
xor XOR2 (N13625, N13623, N5403);
and AND2 (N13626, N13622, N4987);
xor XOR2 (N13627, N13616, N3438);
nand NAND4 (N13628, N13619, N799, N79, N9319);
not NOT1 (N13629, N13613);
xor XOR2 (N13630, N13621, N12335);
not NOT1 (N13631, N13626);
xor XOR2 (N13632, N13630, N11885);
xor XOR2 (N13633, N13627, N1280);
and AND4 (N13634, N13631, N6044, N11745, N5476);
not NOT1 (N13635, N13600);
nand NAND2 (N13636, N13598, N6);
and AND4 (N13637, N13634, N11408, N11571, N12555);
and AND4 (N13638, N13629, N4219, N9746, N513);
or OR2 (N13639, N13633, N7322);
and AND2 (N13640, N13638, N3765);
or OR2 (N13641, N13636, N3812);
and AND2 (N13642, N13625, N4325);
nor NOR3 (N13643, N13639, N4919, N6889);
and AND3 (N13644, N13635, N5641, N8817);
nand NAND3 (N13645, N13628, N7534, N5228);
and AND2 (N13646, N13632, N7632);
xor XOR2 (N13647, N13642, N7523);
nand NAND3 (N13648, N13647, N1354, N10896);
and AND3 (N13649, N13643, N6014, N6707);
xor XOR2 (N13650, N13649, N2527);
nor NOR3 (N13651, N13650, N12720, N4412);
nand NAND3 (N13652, N13646, N12796, N2700);
nand NAND4 (N13653, N13644, N2831, N6383, N1045);
xor XOR2 (N13654, N13645, N1456);
and AND3 (N13655, N13651, N12408, N12508);
nor NOR4 (N13656, N13624, N5295, N6621, N1514);
xor XOR2 (N13657, N13637, N6331);
and AND2 (N13658, N13653, N10562);
not NOT1 (N13659, N13656);
nor NOR2 (N13660, N13648, N5669);
nand NAND3 (N13661, N13658, N7818, N2820);
xor XOR2 (N13662, N13618, N2318);
buf BUF1 (N13663, N13641);
buf BUF1 (N13664, N13652);
or OR2 (N13665, N13654, N1354);
and AND2 (N13666, N13660, N9083);
or OR4 (N13667, N13659, N7813, N11632, N12577);
nor NOR3 (N13668, N13657, N7302, N5300);
not NOT1 (N13669, N13661);
nand NAND2 (N13670, N13662, N471);
and AND2 (N13671, N13664, N4885);
nor NOR3 (N13672, N13668, N785, N7855);
nor NOR2 (N13673, N13665, N1243);
xor XOR2 (N13674, N13671, N12708);
buf BUF1 (N13675, N13640);
nor NOR4 (N13676, N13666, N7141, N1170, N10999);
nand NAND2 (N13677, N13663, N7290);
not NOT1 (N13678, N13674);
or OR2 (N13679, N13672, N11822);
nand NAND4 (N13680, N13677, N4327, N12798, N6614);
xor XOR2 (N13681, N13680, N10071);
or OR2 (N13682, N13679, N4182);
nor NOR3 (N13683, N13667, N4460, N4701);
nand NAND3 (N13684, N13678, N1743, N11852);
not NOT1 (N13685, N13655);
or OR3 (N13686, N13676, N8691, N6794);
nor NOR4 (N13687, N13673, N6158, N500, N1139);
xor XOR2 (N13688, N13687, N6746);
nor NOR2 (N13689, N13688, N99);
xor XOR2 (N13690, N13684, N7438);
nor NOR2 (N13691, N13690, N4300);
nand NAND2 (N13692, N13683, N8274);
not NOT1 (N13693, N13675);
nand NAND4 (N13694, N13691, N4613, N4834, N10176);
or OR2 (N13695, N13689, N96);
nor NOR3 (N13696, N13695, N13415, N5224);
buf BUF1 (N13697, N13670);
buf BUF1 (N13698, N13693);
and AND2 (N13699, N13692, N2833);
buf BUF1 (N13700, N13699);
xor XOR2 (N13701, N13700, N7231);
buf BUF1 (N13702, N13701);
nand NAND3 (N13703, N13685, N1071, N3170);
not NOT1 (N13704, N13686);
not NOT1 (N13705, N13704);
or OR4 (N13706, N13682, N6761, N9548, N1959);
xor XOR2 (N13707, N13698, N4311);
and AND3 (N13708, N13702, N5107, N11460);
not NOT1 (N13709, N13694);
nand NAND3 (N13710, N13708, N8164, N9446);
xor XOR2 (N13711, N13697, N8228);
nor NOR3 (N13712, N13711, N8394, N12393);
and AND3 (N13713, N13706, N12392, N11258);
or OR4 (N13714, N13703, N11540, N8633, N12648);
nor NOR3 (N13715, N13713, N11345, N9080);
or OR4 (N13716, N13710, N1760, N2535, N11296);
xor XOR2 (N13717, N13669, N3137);
nor NOR2 (N13718, N13712, N7489);
not NOT1 (N13719, N13707);
nor NOR2 (N13720, N13681, N4256);
buf BUF1 (N13721, N13705);
not NOT1 (N13722, N13716);
not NOT1 (N13723, N13717);
buf BUF1 (N13724, N13723);
nor NOR4 (N13725, N13709, N11436, N8120, N11458);
or OR4 (N13726, N13724, N4769, N3535, N13139);
nor NOR2 (N13727, N13719, N12933);
xor XOR2 (N13728, N13727, N1089);
or OR2 (N13729, N13714, N12309);
buf BUF1 (N13730, N13728);
nor NOR4 (N13731, N13720, N12441, N6052, N6180);
or OR2 (N13732, N13729, N749);
not NOT1 (N13733, N13732);
buf BUF1 (N13734, N13721);
nand NAND3 (N13735, N13726, N7302, N10908);
not NOT1 (N13736, N13735);
and AND4 (N13737, N13725, N7287, N9503, N13700);
xor XOR2 (N13738, N13718, N6997);
buf BUF1 (N13739, N13730);
nor NOR2 (N13740, N13736, N1706);
and AND3 (N13741, N13715, N13294, N13198);
or OR2 (N13742, N13739, N10181);
and AND3 (N13743, N13731, N611, N9567);
nand NAND4 (N13744, N13742, N3455, N13626, N290);
xor XOR2 (N13745, N13741, N1378);
xor XOR2 (N13746, N13740, N4660);
xor XOR2 (N13747, N13744, N5570);
not NOT1 (N13748, N13734);
not NOT1 (N13749, N13748);
buf BUF1 (N13750, N13743);
not NOT1 (N13751, N13750);
xor XOR2 (N13752, N13747, N6954);
nor NOR2 (N13753, N13746, N11140);
and AND2 (N13754, N13751, N2062);
nand NAND2 (N13755, N13737, N10428);
nand NAND3 (N13756, N13753, N13389, N492);
buf BUF1 (N13757, N13755);
not NOT1 (N13758, N13722);
nor NOR3 (N13759, N13738, N11815, N9594);
not NOT1 (N13760, N13752);
xor XOR2 (N13761, N13696, N10386);
buf BUF1 (N13762, N13754);
nor NOR4 (N13763, N13756, N5278, N6694, N12714);
nor NOR2 (N13764, N13733, N12075);
not NOT1 (N13765, N13761);
not NOT1 (N13766, N13764);
buf BUF1 (N13767, N13759);
buf BUF1 (N13768, N13766);
buf BUF1 (N13769, N13763);
nand NAND2 (N13770, N13757, N685);
buf BUF1 (N13771, N13769);
not NOT1 (N13772, N13768);
not NOT1 (N13773, N13770);
nor NOR2 (N13774, N13772, N13182);
not NOT1 (N13775, N13745);
xor XOR2 (N13776, N13760, N4831);
xor XOR2 (N13777, N13771, N535);
or OR2 (N13778, N13774, N6622);
xor XOR2 (N13779, N13776, N1046);
not NOT1 (N13780, N13767);
or OR2 (N13781, N13779, N7782);
buf BUF1 (N13782, N13758);
and AND2 (N13783, N13781, N13148);
nor NOR2 (N13784, N13773, N2014);
nand NAND2 (N13785, N13778, N3272);
buf BUF1 (N13786, N13782);
buf BUF1 (N13787, N13749);
and AND4 (N13788, N13762, N1341, N901, N11939);
or OR3 (N13789, N13775, N2612, N13304);
buf BUF1 (N13790, N13788);
or OR3 (N13791, N13790, N8162, N13758);
and AND2 (N13792, N13783, N1675);
nand NAND2 (N13793, N13784, N3227);
or OR2 (N13794, N13789, N9408);
not NOT1 (N13795, N13765);
and AND4 (N13796, N13785, N10804, N2153, N5643);
buf BUF1 (N13797, N13777);
nor NOR3 (N13798, N13787, N12121, N5035);
xor XOR2 (N13799, N13795, N5341);
buf BUF1 (N13800, N13793);
buf BUF1 (N13801, N13800);
buf BUF1 (N13802, N13791);
nand NAND4 (N13803, N13792, N6337, N166, N6354);
or OR4 (N13804, N13797, N441, N5261, N124);
xor XOR2 (N13805, N13803, N8159);
or OR2 (N13806, N13798, N4080);
and AND3 (N13807, N13786, N1206, N10034);
nor NOR3 (N13808, N13799, N10005, N5419);
not NOT1 (N13809, N13802);
nor NOR4 (N13810, N13801, N12869, N11396, N7074);
not NOT1 (N13811, N13807);
buf BUF1 (N13812, N13780);
nor NOR3 (N13813, N13794, N1605, N2712);
nand NAND4 (N13814, N13811, N7669, N12105, N9607);
or OR2 (N13815, N13813, N11841);
or OR4 (N13816, N13808, N9465, N6618, N101);
not NOT1 (N13817, N13796);
nand NAND3 (N13818, N13805, N3335, N10619);
xor XOR2 (N13819, N13814, N8799);
buf BUF1 (N13820, N13809);
or OR4 (N13821, N13819, N8142, N8648, N3369);
xor XOR2 (N13822, N13815, N3158);
xor XOR2 (N13823, N13821, N1459);
nand NAND3 (N13824, N13817, N7434, N11094);
nor NOR4 (N13825, N13810, N7551, N11317, N5452);
nand NAND3 (N13826, N13806, N9087, N3884);
nor NOR4 (N13827, N13804, N4853, N8711, N8113);
and AND4 (N13828, N13827, N3187, N9896, N10807);
not NOT1 (N13829, N13820);
and AND3 (N13830, N13826, N1237, N2688);
nand NAND3 (N13831, N13816, N13062, N8294);
nor NOR4 (N13832, N13829, N2883, N2748, N3762);
and AND2 (N13833, N13818, N5440);
and AND4 (N13834, N13828, N3561, N1343, N6984);
xor XOR2 (N13835, N13831, N9751);
or OR3 (N13836, N13830, N12669, N8369);
and AND4 (N13837, N13833, N5739, N6083, N12914);
buf BUF1 (N13838, N13832);
not NOT1 (N13839, N13825);
not NOT1 (N13840, N13812);
nand NAND4 (N13841, N13838, N10374, N3491, N11742);
and AND2 (N13842, N13822, N10599);
nand NAND2 (N13843, N13842, N1812);
or OR3 (N13844, N13839, N12521, N4109);
nand NAND2 (N13845, N13837, N11312);
buf BUF1 (N13846, N13836);
buf BUF1 (N13847, N13844);
nor NOR4 (N13848, N13835, N11979, N4626, N13797);
not NOT1 (N13849, N13847);
xor XOR2 (N13850, N13834, N25);
nand NAND4 (N13851, N13850, N662, N6831, N11698);
buf BUF1 (N13852, N13823);
nand NAND4 (N13853, N13845, N2931, N6942, N4330);
nor NOR3 (N13854, N13841, N9236, N11298);
or OR3 (N13855, N13846, N436, N3595);
and AND4 (N13856, N13843, N10516, N450, N2970);
buf BUF1 (N13857, N13824);
xor XOR2 (N13858, N13848, N9948);
and AND4 (N13859, N13840, N3824, N9447, N3964);
and AND3 (N13860, N13853, N8679, N2169);
or OR2 (N13861, N13856, N12783);
or OR3 (N13862, N13857, N12133, N4777);
and AND2 (N13863, N13861, N1421);
nand NAND2 (N13864, N13859, N1828);
and AND2 (N13865, N13855, N3963);
buf BUF1 (N13866, N13864);
and AND4 (N13867, N13862, N6497, N4962, N8350);
not NOT1 (N13868, N13860);
nand NAND4 (N13869, N13867, N12005, N1112, N3340);
not NOT1 (N13870, N13863);
xor XOR2 (N13871, N13849, N5756);
not NOT1 (N13872, N13851);
nor NOR2 (N13873, N13871, N7944);
buf BUF1 (N13874, N13854);
nor NOR3 (N13875, N13872, N89, N6878);
xor XOR2 (N13876, N13858, N13053);
and AND3 (N13877, N13874, N12565, N857);
nor NOR2 (N13878, N13877, N5454);
nand NAND2 (N13879, N13873, N7490);
not NOT1 (N13880, N13875);
or OR3 (N13881, N13866, N2941, N8555);
or OR2 (N13882, N13879, N9817);
xor XOR2 (N13883, N13869, N491);
xor XOR2 (N13884, N13882, N3926);
not NOT1 (N13885, N13868);
or OR2 (N13886, N13881, N9610);
nand NAND2 (N13887, N13885, N1232);
buf BUF1 (N13888, N13887);
xor XOR2 (N13889, N13865, N5848);
buf BUF1 (N13890, N13884);
or OR4 (N13891, N13883, N9848, N1648, N5695);
not NOT1 (N13892, N13878);
or OR4 (N13893, N13852, N9646, N7980, N11994);
buf BUF1 (N13894, N13890);
and AND3 (N13895, N13892, N6985, N11914);
or OR2 (N13896, N13889, N8505);
buf BUF1 (N13897, N13886);
or OR3 (N13898, N13876, N6405, N12460);
buf BUF1 (N13899, N13888);
or OR4 (N13900, N13896, N8752, N5176, N8631);
not NOT1 (N13901, N13900);
not NOT1 (N13902, N13880);
buf BUF1 (N13903, N13898);
buf BUF1 (N13904, N13895);
not NOT1 (N13905, N13897);
xor XOR2 (N13906, N13905, N5383);
nor NOR3 (N13907, N13903, N10107, N4314);
buf BUF1 (N13908, N13891);
or OR3 (N13909, N13906, N2095, N5542);
nand NAND3 (N13910, N13907, N635, N6667);
nand NAND2 (N13911, N13909, N5733);
xor XOR2 (N13912, N13904, N5194);
nor NOR4 (N13913, N13902, N5035, N4511, N949);
not NOT1 (N13914, N13910);
or OR4 (N13915, N13870, N13521, N6020, N1481);
buf BUF1 (N13916, N13893);
and AND3 (N13917, N13913, N9181, N9236);
not NOT1 (N13918, N13908);
xor XOR2 (N13919, N13916, N6654);
nand NAND2 (N13920, N13901, N7746);
nand NAND2 (N13921, N13894, N12451);
not NOT1 (N13922, N13912);
xor XOR2 (N13923, N13919, N11661);
and AND3 (N13924, N13921, N13624, N12908);
nand NAND4 (N13925, N13917, N599, N3177, N9963);
and AND2 (N13926, N13899, N8617);
not NOT1 (N13927, N13923);
xor XOR2 (N13928, N13914, N11822);
or OR2 (N13929, N13922, N1126);
or OR4 (N13930, N13911, N13596, N5804, N12258);
or OR3 (N13931, N13925, N13051, N822);
or OR3 (N13932, N13920, N10933, N4079);
or OR4 (N13933, N13918, N3891, N4877, N394);
and AND4 (N13934, N13929, N9065, N10663, N8887);
and AND3 (N13935, N13915, N1307, N9219);
not NOT1 (N13936, N13935);
xor XOR2 (N13937, N13928, N12695);
or OR2 (N13938, N13933, N1961);
and AND2 (N13939, N13930, N13534);
xor XOR2 (N13940, N13938, N752);
or OR4 (N13941, N13940, N10552, N5155, N2998);
nand NAND3 (N13942, N13934, N13865, N1986);
nand NAND2 (N13943, N13927, N3665);
and AND2 (N13944, N13942, N13124);
nor NOR4 (N13945, N13943, N10645, N5349, N12854);
not NOT1 (N13946, N13939);
xor XOR2 (N13947, N13926, N3391);
nor NOR3 (N13948, N13946, N11834, N6791);
xor XOR2 (N13949, N13947, N13553);
xor XOR2 (N13950, N13931, N3270);
xor XOR2 (N13951, N13945, N1808);
and AND4 (N13952, N13948, N5486, N736, N2212);
nand NAND4 (N13953, N13936, N10961, N9776, N4100);
or OR4 (N13954, N13953, N5342, N9844, N11072);
buf BUF1 (N13955, N13937);
not NOT1 (N13956, N13955);
buf BUF1 (N13957, N13949);
and AND2 (N13958, N13951, N6189);
or OR4 (N13959, N13950, N8048, N8405, N4863);
and AND2 (N13960, N13924, N4006);
not NOT1 (N13961, N13941);
and AND4 (N13962, N13932, N1052, N328, N2504);
nand NAND2 (N13963, N13957, N13111);
or OR4 (N13964, N13952, N12463, N3271, N3010);
not NOT1 (N13965, N13961);
or OR4 (N13966, N13965, N1886, N4574, N1612);
nor NOR4 (N13967, N13960, N4356, N4316, N3571);
nor NOR4 (N13968, N13967, N10357, N8272, N4418);
nor NOR4 (N13969, N13964, N6420, N1275, N9925);
nor NOR4 (N13970, N13944, N8724, N241, N6914);
or OR2 (N13971, N13963, N11336);
and AND4 (N13972, N13956, N13948, N6348, N4863);
buf BUF1 (N13973, N13966);
not NOT1 (N13974, N13954);
nand NAND4 (N13975, N13974, N2075, N1737, N6218);
nand NAND4 (N13976, N13975, N8846, N7604, N10902);
or OR2 (N13977, N13970, N2557);
nand NAND3 (N13978, N13976, N5529, N3213);
not NOT1 (N13979, N13968);
or OR2 (N13980, N13959, N7751);
not NOT1 (N13981, N13973);
buf BUF1 (N13982, N13958);
not NOT1 (N13983, N13981);
nand NAND4 (N13984, N13972, N3970, N6904, N1667);
buf BUF1 (N13985, N13969);
and AND4 (N13986, N13980, N9377, N8985, N6077);
not NOT1 (N13987, N13985);
buf BUF1 (N13988, N13978);
xor XOR2 (N13989, N13977, N3294);
not NOT1 (N13990, N13988);
xor XOR2 (N13991, N13990, N1689);
nor NOR4 (N13992, N13991, N2393, N9057, N9078);
or OR3 (N13993, N13989, N9507, N7837);
xor XOR2 (N13994, N13993, N11372);
not NOT1 (N13995, N13982);
or OR4 (N13996, N13994, N6162, N11168, N12916);
xor XOR2 (N13997, N13962, N558);
nand NAND3 (N13998, N13983, N1188, N6765);
and AND4 (N13999, N13971, N5264, N7544, N1066);
or OR4 (N14000, N13995, N429, N12792, N13418);
and AND3 (N14001, N13996, N7328, N11600);
or OR4 (N14002, N13986, N8518, N9347, N2322);
buf BUF1 (N14003, N13987);
nor NOR2 (N14004, N13992, N10959);
nor NOR4 (N14005, N13999, N2013, N7479, N6007);
not NOT1 (N14006, N13979);
not NOT1 (N14007, N14000);
or OR4 (N14008, N14006, N8254, N13717, N4893);
buf BUF1 (N14009, N13998);
buf BUF1 (N14010, N14008);
nor NOR3 (N14011, N13997, N5205, N4380);
or OR2 (N14012, N14005, N10717);
or OR2 (N14013, N14004, N2723);
buf BUF1 (N14014, N14012);
nor NOR4 (N14015, N13984, N1857, N443, N8219);
buf BUF1 (N14016, N14009);
nor NOR3 (N14017, N14007, N12525, N11600);
or OR3 (N14018, N14017, N2973, N7848);
nand NAND4 (N14019, N14014, N10495, N1510, N11319);
nand NAND3 (N14020, N14010, N10168, N3651);
and AND3 (N14021, N14019, N1531, N8487);
nor NOR4 (N14022, N14013, N1686, N5951, N1722);
xor XOR2 (N14023, N14021, N13114);
nand NAND3 (N14024, N14001, N11746, N5136);
or OR2 (N14025, N14023, N12813);
xor XOR2 (N14026, N14015, N992);
buf BUF1 (N14027, N14016);
nor NOR3 (N14028, N14011, N3167, N4235);
buf BUF1 (N14029, N14003);
xor XOR2 (N14030, N14026, N10965);
and AND4 (N14031, N14030, N8821, N4244, N12170);
buf BUF1 (N14032, N14020);
nand NAND3 (N14033, N14025, N7017, N5131);
not NOT1 (N14034, N14024);
xor XOR2 (N14035, N14027, N13981);
and AND3 (N14036, N14032, N13826, N5843);
or OR4 (N14037, N14034, N2579, N13126, N10264);
not NOT1 (N14038, N14028);
or OR4 (N14039, N14018, N13259, N12596, N3853);
or OR2 (N14040, N14037, N9541);
xor XOR2 (N14041, N14036, N10499);
nand NAND2 (N14042, N14041, N4464);
nand NAND3 (N14043, N14022, N9870, N2822);
nand NAND4 (N14044, N14040, N5527, N8582, N6254);
or OR3 (N14045, N14039, N3934, N6049);
nand NAND3 (N14046, N14038, N9396, N470);
nor NOR2 (N14047, N14002, N4685);
xor XOR2 (N14048, N14035, N5472);
or OR3 (N14049, N14045, N12161, N1442);
buf BUF1 (N14050, N14047);
nor NOR4 (N14051, N14044, N8023, N14007, N6065);
and AND2 (N14052, N14051, N3602);
or OR2 (N14053, N14052, N8159);
not NOT1 (N14054, N14033);
or OR2 (N14055, N14042, N11671);
not NOT1 (N14056, N14048);
and AND4 (N14057, N14029, N10363, N5676, N13574);
or OR3 (N14058, N14056, N12181, N12503);
or OR3 (N14059, N14058, N11210, N5274);
or OR3 (N14060, N14049, N13786, N9575);
buf BUF1 (N14061, N14050);
xor XOR2 (N14062, N14053, N7226);
and AND4 (N14063, N14062, N5805, N894, N12676);
nor NOR2 (N14064, N14057, N12617);
or OR2 (N14065, N14046, N13777);
and AND2 (N14066, N14064, N10190);
nand NAND3 (N14067, N14065, N11307, N11382);
not NOT1 (N14068, N14055);
not NOT1 (N14069, N14043);
buf BUF1 (N14070, N14063);
xor XOR2 (N14071, N14060, N2152);
nand NAND2 (N14072, N14054, N2560);
xor XOR2 (N14073, N14066, N9727);
or OR4 (N14074, N14071, N1626, N12183, N7284);
buf BUF1 (N14075, N14067);
nand NAND4 (N14076, N14031, N1553, N12812, N1185);
xor XOR2 (N14077, N14068, N737);
nand NAND3 (N14078, N14070, N6108, N3372);
or OR2 (N14079, N14072, N1110);
nor NOR2 (N14080, N14059, N4094);
nor NOR2 (N14081, N14079, N4969);
nand NAND2 (N14082, N14076, N1156);
buf BUF1 (N14083, N14080);
not NOT1 (N14084, N14061);
nand NAND3 (N14085, N14074, N2574, N6135);
not NOT1 (N14086, N14073);
or OR2 (N14087, N14081, N2403);
not NOT1 (N14088, N14069);
nor NOR2 (N14089, N14084, N5445);
nor NOR2 (N14090, N14078, N5265);
or OR4 (N14091, N14089, N4770, N8027, N13097);
buf BUF1 (N14092, N14085);
or OR3 (N14093, N14090, N3129, N5388);
nor NOR4 (N14094, N14077, N143, N4552, N4438);
or OR4 (N14095, N14082, N9597, N600, N1705);
or OR3 (N14096, N14083, N5501, N9900);
xor XOR2 (N14097, N14091, N1798);
not NOT1 (N14098, N14097);
buf BUF1 (N14099, N14088);
or OR4 (N14100, N14094, N3838, N6951, N1269);
or OR3 (N14101, N14096, N13319, N9952);
and AND2 (N14102, N14098, N1005);
nor NOR2 (N14103, N14093, N5296);
or OR2 (N14104, N14075, N4152);
buf BUF1 (N14105, N14104);
nor NOR4 (N14106, N14087, N10753, N1810, N741);
nor NOR2 (N14107, N14101, N13167);
not NOT1 (N14108, N14095);
nand NAND3 (N14109, N14092, N942, N13073);
buf BUF1 (N14110, N14108);
not NOT1 (N14111, N14099);
or OR4 (N14112, N14110, N3815, N2741, N8948);
and AND3 (N14113, N14102, N9242, N7171);
nor NOR3 (N14114, N14107, N1933, N12016);
nand NAND3 (N14115, N14109, N11642, N7330);
nand NAND4 (N14116, N14106, N6358, N12449, N4966);
nand NAND3 (N14117, N14113, N6818, N6252);
nor NOR3 (N14118, N14105, N2797, N4785);
not NOT1 (N14119, N14115);
not NOT1 (N14120, N14112);
nand NAND3 (N14121, N14114, N7278, N12898);
buf BUF1 (N14122, N14120);
nor NOR4 (N14123, N14118, N6831, N4028, N6486);
xor XOR2 (N14124, N14121, N3522);
nand NAND3 (N14125, N14103, N4175, N1252);
and AND4 (N14126, N14086, N9444, N8601, N9125);
xor XOR2 (N14127, N14111, N13252);
xor XOR2 (N14128, N14127, N4961);
buf BUF1 (N14129, N14123);
nor NOR2 (N14130, N14119, N9725);
nand NAND3 (N14131, N14124, N8252, N9328);
nor NOR3 (N14132, N14122, N10930, N12093);
nand NAND2 (N14133, N14128, N5019);
not NOT1 (N14134, N14126);
and AND2 (N14135, N14130, N10873);
or OR3 (N14136, N14133, N1717, N151);
buf BUF1 (N14137, N14131);
xor XOR2 (N14138, N14136, N6720);
buf BUF1 (N14139, N14134);
or OR3 (N14140, N14138, N11953, N13394);
xor XOR2 (N14141, N14116, N7650);
and AND4 (N14142, N14132, N5815, N6325, N1132);
not NOT1 (N14143, N14140);
or OR2 (N14144, N14125, N4708);
not NOT1 (N14145, N14129);
or OR2 (N14146, N14144, N10720);
buf BUF1 (N14147, N14137);
nor NOR2 (N14148, N14141, N13699);
nand NAND2 (N14149, N14100, N12053);
nor NOR3 (N14150, N14142, N3819, N8244);
buf BUF1 (N14151, N14150);
nand NAND4 (N14152, N14145, N7031, N11045, N3922);
nand NAND2 (N14153, N14139, N1112);
or OR4 (N14154, N14135, N7541, N1493, N7357);
and AND4 (N14155, N14154, N11463, N9844, N13236);
buf BUF1 (N14156, N14117);
xor XOR2 (N14157, N14152, N516);
nand NAND2 (N14158, N14147, N13144);
or OR3 (N14159, N14157, N12078, N9626);
or OR2 (N14160, N14159, N13850);
not NOT1 (N14161, N14143);
nor NOR4 (N14162, N14151, N4881, N6136, N8123);
or OR2 (N14163, N14161, N9351);
xor XOR2 (N14164, N14162, N10433);
nand NAND4 (N14165, N14163, N1938, N4834, N7130);
not NOT1 (N14166, N14158);
and AND2 (N14167, N14156, N11276);
xor XOR2 (N14168, N14146, N3793);
xor XOR2 (N14169, N14168, N13860);
not NOT1 (N14170, N14148);
buf BUF1 (N14171, N14170);
nand NAND2 (N14172, N14155, N3706);
nor NOR4 (N14173, N14171, N10856, N3328, N6572);
not NOT1 (N14174, N14165);
and AND3 (N14175, N14164, N5331, N5347);
buf BUF1 (N14176, N14172);
nor NOR2 (N14177, N14173, N802);
not NOT1 (N14178, N14177);
nand NAND4 (N14179, N14149, N10095, N7182, N7917);
and AND2 (N14180, N14179, N9211);
not NOT1 (N14181, N14153);
not NOT1 (N14182, N14160);
and AND3 (N14183, N14169, N12529, N11919);
nand NAND4 (N14184, N14180, N2856, N1068, N6103);
and AND3 (N14185, N14183, N8382, N8241);
nand NAND4 (N14186, N14166, N1109, N2018, N12237);
not NOT1 (N14187, N14174);
not NOT1 (N14188, N14186);
and AND2 (N14189, N14188, N2260);
nor NOR3 (N14190, N14167, N8225, N2287);
nand NAND3 (N14191, N14189, N4922, N1645);
and AND2 (N14192, N14175, N3186);
nand NAND3 (N14193, N14192, N14142, N4080);
nand NAND4 (N14194, N14185, N8045, N11009, N2934);
not NOT1 (N14195, N14182);
buf BUF1 (N14196, N14181);
nor NOR2 (N14197, N14193, N4280);
nand NAND4 (N14198, N14190, N4160, N1276, N8823);
nand NAND4 (N14199, N14196, N14024, N711, N12722);
or OR3 (N14200, N14197, N901, N10689);
buf BUF1 (N14201, N14195);
not NOT1 (N14202, N14187);
and AND2 (N14203, N14202, N3902);
xor XOR2 (N14204, N14200, N526);
buf BUF1 (N14205, N14203);
or OR4 (N14206, N14191, N13493, N2596, N6522);
and AND2 (N14207, N14204, N1764);
xor XOR2 (N14208, N14178, N8691);
nand NAND3 (N14209, N14206, N6575, N7381);
not NOT1 (N14210, N14208);
nor NOR3 (N14211, N14210, N4480, N1948);
nor NOR3 (N14212, N14199, N5908, N5034);
not NOT1 (N14213, N14212);
xor XOR2 (N14214, N14209, N1698);
xor XOR2 (N14215, N14198, N2412);
nand NAND2 (N14216, N14176, N2771);
xor XOR2 (N14217, N14194, N665);
and AND4 (N14218, N14215, N6784, N11736, N2759);
or OR3 (N14219, N14201, N13183, N13467);
nand NAND3 (N14220, N14211, N4218, N2863);
nand NAND2 (N14221, N14220, N8424);
and AND4 (N14222, N14205, N5506, N1122, N11642);
nor NOR3 (N14223, N14184, N521, N13249);
nand NAND2 (N14224, N14217, N3360);
not NOT1 (N14225, N14207);
not NOT1 (N14226, N14222);
and AND2 (N14227, N14224, N5870);
or OR3 (N14228, N14219, N6500, N4717);
and AND2 (N14229, N14216, N6529);
and AND2 (N14230, N14228, N13558);
xor XOR2 (N14231, N14230, N2464);
nand NAND3 (N14232, N14229, N13099, N5046);
xor XOR2 (N14233, N14223, N9656);
and AND2 (N14234, N14231, N5457);
not NOT1 (N14235, N14221);
and AND2 (N14236, N14233, N7072);
nand NAND4 (N14237, N14227, N6975, N9737, N3804);
and AND2 (N14238, N14214, N5738);
xor XOR2 (N14239, N14225, N8848);
xor XOR2 (N14240, N14213, N10757);
buf BUF1 (N14241, N14238);
nor NOR2 (N14242, N14226, N5574);
not NOT1 (N14243, N14232);
nor NOR4 (N14244, N14235, N13212, N7581, N8482);
nand NAND4 (N14245, N14243, N4902, N7730, N6534);
nand NAND3 (N14246, N14218, N624, N10036);
or OR2 (N14247, N14241, N8192);
or OR3 (N14248, N14240, N223, N11964);
not NOT1 (N14249, N14246);
xor XOR2 (N14250, N14239, N10740);
not NOT1 (N14251, N14236);
or OR3 (N14252, N14251, N4541, N1659);
not NOT1 (N14253, N14247);
buf BUF1 (N14254, N14250);
buf BUF1 (N14255, N14254);
xor XOR2 (N14256, N14242, N13972);
or OR2 (N14257, N14244, N11815);
nor NOR4 (N14258, N14256, N11607, N12426, N255);
nor NOR4 (N14259, N14258, N10899, N11447, N12649);
nor NOR3 (N14260, N14237, N1533, N8528);
not NOT1 (N14261, N14234);
nor NOR2 (N14262, N14245, N12703);
nand NAND4 (N14263, N14260, N5278, N9359, N10890);
nand NAND2 (N14264, N14255, N13626);
and AND3 (N14265, N14262, N4721, N13740);
nand NAND3 (N14266, N14252, N12835, N6135);
xor XOR2 (N14267, N14264, N5131);
buf BUF1 (N14268, N14266);
nand NAND3 (N14269, N14257, N12527, N10872);
nand NAND3 (N14270, N14267, N13729, N4177);
buf BUF1 (N14271, N14265);
not NOT1 (N14272, N14263);
or OR3 (N14273, N14249, N7062, N5758);
or OR4 (N14274, N14272, N1915, N13260, N10719);
nand NAND2 (N14275, N14274, N3081);
buf BUF1 (N14276, N14261);
nand NAND4 (N14277, N14270, N3374, N6714, N5087);
and AND4 (N14278, N14248, N1876, N10518, N6572);
nand NAND4 (N14279, N14268, N5078, N8282, N6660);
nor NOR4 (N14280, N14253, N4693, N5531, N1993);
buf BUF1 (N14281, N14271);
and AND3 (N14282, N14280, N7948, N11621);
buf BUF1 (N14283, N14273);
not NOT1 (N14284, N14276);
xor XOR2 (N14285, N14269, N4595);
and AND4 (N14286, N14281, N11536, N219, N12052);
and AND4 (N14287, N14259, N75, N4568, N8483);
buf BUF1 (N14288, N14282);
not NOT1 (N14289, N14275);
and AND2 (N14290, N14283, N6512);
buf BUF1 (N14291, N14290);
and AND3 (N14292, N14287, N4169, N5600);
xor XOR2 (N14293, N14289, N13666);
xor XOR2 (N14294, N14285, N14252);
nor NOR4 (N14295, N14277, N7110, N8819, N8795);
nor NOR4 (N14296, N14295, N5965, N10238, N3477);
and AND4 (N14297, N14279, N9202, N6773, N1706);
not NOT1 (N14298, N14286);
buf BUF1 (N14299, N14284);
and AND2 (N14300, N14297, N2826);
or OR3 (N14301, N14288, N9717, N1177);
nand NAND4 (N14302, N14301, N6561, N9625, N9917);
or OR4 (N14303, N14291, N10507, N508, N2838);
buf BUF1 (N14304, N14293);
not NOT1 (N14305, N14303);
nand NAND4 (N14306, N14299, N5218, N9924, N2439);
xor XOR2 (N14307, N14292, N12356);
or OR2 (N14308, N14305, N14273);
buf BUF1 (N14309, N14308);
not NOT1 (N14310, N14306);
nand NAND4 (N14311, N14309, N2850, N3827, N7440);
buf BUF1 (N14312, N14310);
not NOT1 (N14313, N14300);
buf BUF1 (N14314, N14294);
not NOT1 (N14315, N14296);
and AND4 (N14316, N14302, N10725, N10331, N4668);
not NOT1 (N14317, N14278);
not NOT1 (N14318, N14304);
not NOT1 (N14319, N14316);
nand NAND4 (N14320, N14315, N10588, N1301, N9763);
xor XOR2 (N14321, N14314, N13347);
nor NOR2 (N14322, N14312, N7614);
not NOT1 (N14323, N14321);
or OR4 (N14324, N14318, N8774, N2727, N2469);
nor NOR3 (N14325, N14313, N9219, N8927);
and AND2 (N14326, N14325, N13996);
xor XOR2 (N14327, N14307, N5842);
nor NOR2 (N14328, N14311, N1946);
xor XOR2 (N14329, N14317, N3074);
buf BUF1 (N14330, N14323);
not NOT1 (N14331, N14329);
not NOT1 (N14332, N14320);
xor XOR2 (N14333, N14330, N3385);
nand NAND2 (N14334, N14322, N5438);
xor XOR2 (N14335, N14324, N12538);
and AND2 (N14336, N14328, N13535);
buf BUF1 (N14337, N14334);
not NOT1 (N14338, N14336);
xor XOR2 (N14339, N14333, N8945);
xor XOR2 (N14340, N14332, N13895);
or OR2 (N14341, N14331, N14286);
buf BUF1 (N14342, N14341);
and AND4 (N14343, N14335, N6027, N6708, N7267);
buf BUF1 (N14344, N14340);
and AND3 (N14345, N14319, N6705, N6671);
not NOT1 (N14346, N14298);
xor XOR2 (N14347, N14327, N4371);
or OR2 (N14348, N14343, N4821);
nand NAND4 (N14349, N14339, N4407, N6890, N13243);
not NOT1 (N14350, N14326);
nor NOR4 (N14351, N14348, N13796, N6966, N9073);
not NOT1 (N14352, N14349);
and AND2 (N14353, N14338, N6680);
buf BUF1 (N14354, N14351);
xor XOR2 (N14355, N14350, N5989);
buf BUF1 (N14356, N14342);
buf BUF1 (N14357, N14346);
nand NAND3 (N14358, N14357, N1923, N503);
nand NAND3 (N14359, N14337, N10345, N2686);
or OR4 (N14360, N14345, N6641, N5414, N8346);
not NOT1 (N14361, N14358);
xor XOR2 (N14362, N14360, N12006);
nor NOR4 (N14363, N14354, N9912, N5928, N1558);
nor NOR3 (N14364, N14347, N8453, N1170);
and AND2 (N14365, N14352, N13994);
or OR2 (N14366, N14364, N2371);
and AND2 (N14367, N14355, N6206);
xor XOR2 (N14368, N14367, N3100);
or OR2 (N14369, N14362, N7989);
xor XOR2 (N14370, N14353, N8486);
not NOT1 (N14371, N14370);
nor NOR4 (N14372, N14366, N9199, N14158, N4369);
and AND4 (N14373, N14365, N11744, N1394, N2855);
nand NAND2 (N14374, N14372, N10777);
and AND4 (N14375, N14374, N8035, N10213, N8047);
nand NAND4 (N14376, N14363, N3859, N9763, N5500);
xor XOR2 (N14377, N14344, N6876);
nor NOR4 (N14378, N14371, N10069, N1514, N9618);
buf BUF1 (N14379, N14378);
xor XOR2 (N14380, N14369, N11525);
and AND4 (N14381, N14373, N6637, N3515, N7341);
not NOT1 (N14382, N14381);
not NOT1 (N14383, N14361);
xor XOR2 (N14384, N14377, N10785);
buf BUF1 (N14385, N14384);
not NOT1 (N14386, N14368);
xor XOR2 (N14387, N14356, N12435);
and AND2 (N14388, N14385, N9343);
and AND4 (N14389, N14386, N7857, N8458, N8415);
nor NOR4 (N14390, N14380, N10084, N8796, N3517);
buf BUF1 (N14391, N14389);
buf BUF1 (N14392, N14383);
nand NAND3 (N14393, N14391, N6403, N6116);
nor NOR2 (N14394, N14390, N6191);
nor NOR2 (N14395, N14387, N8491);
and AND3 (N14396, N14394, N10229, N3741);
buf BUF1 (N14397, N14388);
nand NAND2 (N14398, N14359, N12187);
buf BUF1 (N14399, N14396);
and AND2 (N14400, N14376, N6506);
buf BUF1 (N14401, N14398);
or OR3 (N14402, N14379, N4488, N8253);
and AND2 (N14403, N14395, N3432);
xor XOR2 (N14404, N14397, N5168);
not NOT1 (N14405, N14399);
and AND3 (N14406, N14393, N11673, N1637);
xor XOR2 (N14407, N14404, N10380);
and AND2 (N14408, N14400, N12306);
buf BUF1 (N14409, N14406);
nand NAND3 (N14410, N14409, N4349, N13200);
xor XOR2 (N14411, N14401, N11623);
not NOT1 (N14412, N14410);
nand NAND3 (N14413, N14405, N1683, N11212);
and AND2 (N14414, N14412, N10574);
or OR4 (N14415, N14382, N13962, N13918, N8128);
and AND4 (N14416, N14414, N241, N12211, N153);
buf BUF1 (N14417, N14402);
and AND2 (N14418, N14408, N10322);
or OR4 (N14419, N14413, N14280, N9310, N12245);
buf BUF1 (N14420, N14419);
xor XOR2 (N14421, N14375, N8695);
buf BUF1 (N14422, N14403);
buf BUF1 (N14423, N14417);
nand NAND2 (N14424, N14411, N7623);
or OR3 (N14425, N14418, N10726, N12939);
buf BUF1 (N14426, N14407);
not NOT1 (N14427, N14392);
not NOT1 (N14428, N14423);
or OR2 (N14429, N14427, N7966);
and AND2 (N14430, N14428, N313);
or OR3 (N14431, N14424, N13273, N4517);
not NOT1 (N14432, N14422);
or OR4 (N14433, N14426, N11917, N1028, N12669);
nor NOR3 (N14434, N14429, N6718, N282);
buf BUF1 (N14435, N14421);
xor XOR2 (N14436, N14420, N12515);
nor NOR2 (N14437, N14430, N167);
nand NAND2 (N14438, N14432, N9619);
nand NAND4 (N14439, N14425, N3578, N13944, N9566);
buf BUF1 (N14440, N14435);
nand NAND3 (N14441, N14436, N12351, N13812);
nor NOR4 (N14442, N14440, N11219, N8814, N5892);
buf BUF1 (N14443, N14416);
xor XOR2 (N14444, N14442, N2799);
nand NAND4 (N14445, N14439, N174, N1875, N10735);
buf BUF1 (N14446, N14434);
nand NAND3 (N14447, N14444, N5529, N6842);
or OR4 (N14448, N14445, N7094, N1431, N3766);
buf BUF1 (N14449, N14446);
not NOT1 (N14450, N14415);
nor NOR4 (N14451, N14447, N1223, N4734, N8068);
not NOT1 (N14452, N14438);
or OR4 (N14453, N14449, N5394, N10728, N2581);
xor XOR2 (N14454, N14433, N13652);
not NOT1 (N14455, N14453);
or OR2 (N14456, N14454, N10915);
or OR3 (N14457, N14443, N2747, N5076);
xor XOR2 (N14458, N14448, N2541);
and AND2 (N14459, N14452, N13205);
buf BUF1 (N14460, N14450);
xor XOR2 (N14461, N14455, N5995);
or OR3 (N14462, N14456, N11617, N7673);
and AND3 (N14463, N14459, N5817, N785);
or OR2 (N14464, N14441, N13272);
and AND4 (N14465, N14437, N6297, N576, N13779);
nand NAND2 (N14466, N14431, N224);
nand NAND2 (N14467, N14464, N12058);
nor NOR3 (N14468, N14461, N10694, N10052);
or OR2 (N14469, N14451, N14277);
buf BUF1 (N14470, N14458);
not NOT1 (N14471, N14465);
not NOT1 (N14472, N14470);
not NOT1 (N14473, N14472);
and AND2 (N14474, N14463, N3670);
and AND3 (N14475, N14469, N3991, N1480);
or OR3 (N14476, N14460, N8665, N12465);
nand NAND4 (N14477, N14473, N13841, N1860, N4948);
or OR2 (N14478, N14467, N7339);
xor XOR2 (N14479, N14466, N12518);
xor XOR2 (N14480, N14457, N11221);
nor NOR4 (N14481, N14471, N12726, N6704, N7558);
nor NOR3 (N14482, N14480, N1063, N7217);
and AND2 (N14483, N14476, N11629);
or OR3 (N14484, N14479, N11645, N4108);
or OR3 (N14485, N14462, N13165, N7452);
nand NAND2 (N14486, N14482, N14122);
and AND2 (N14487, N14484, N6375);
and AND3 (N14488, N14478, N5752, N5571);
xor XOR2 (N14489, N14488, N6577);
buf BUF1 (N14490, N14481);
buf BUF1 (N14491, N14477);
nor NOR2 (N14492, N14483, N11189);
not NOT1 (N14493, N14475);
and AND4 (N14494, N14485, N11346, N14120, N5093);
or OR3 (N14495, N14492, N5735, N12207);
or OR2 (N14496, N14495, N14246);
nor NOR4 (N14497, N14487, N9183, N6452, N614);
xor XOR2 (N14498, N14494, N407);
buf BUF1 (N14499, N14496);
and AND2 (N14500, N14489, N1427);
or OR4 (N14501, N14500, N12181, N8470, N13446);
nor NOR4 (N14502, N14474, N12656, N4055, N14231);
not NOT1 (N14503, N14501);
buf BUF1 (N14504, N14493);
or OR2 (N14505, N14504, N384);
not NOT1 (N14506, N14486);
or OR3 (N14507, N14505, N11344, N931);
buf BUF1 (N14508, N14503);
or OR4 (N14509, N14507, N9943, N11829, N14250);
and AND2 (N14510, N14491, N12323);
nor NOR2 (N14511, N14468, N10823);
and AND4 (N14512, N14497, N2251, N4531, N4773);
xor XOR2 (N14513, N14506, N5234);
or OR2 (N14514, N14508, N11544);
not NOT1 (N14515, N14513);
not NOT1 (N14516, N14515);
not NOT1 (N14517, N14512);
nor NOR4 (N14518, N14516, N12810, N5240, N9523);
nor NOR4 (N14519, N14517, N12538, N9062, N14033);
buf BUF1 (N14520, N14499);
buf BUF1 (N14521, N14514);
nand NAND3 (N14522, N14490, N4265, N12400);
nor NOR4 (N14523, N14511, N6788, N9687, N4658);
nand NAND4 (N14524, N14518, N11239, N822, N8847);
nor NOR2 (N14525, N14520, N12064);
nor NOR4 (N14526, N14502, N1560, N14108, N6526);
buf BUF1 (N14527, N14522);
buf BUF1 (N14528, N14509);
nor NOR3 (N14529, N14528, N1065, N12509);
nand NAND2 (N14530, N14510, N5089);
or OR3 (N14531, N14526, N4099, N14462);
nor NOR4 (N14532, N14498, N12073, N8095, N13999);
nor NOR4 (N14533, N14521, N5978, N9682, N799);
not NOT1 (N14534, N14519);
nand NAND2 (N14535, N14527, N2675);
xor XOR2 (N14536, N14525, N6578);
and AND2 (N14537, N14536, N3571);
and AND3 (N14538, N14531, N834, N5245);
buf BUF1 (N14539, N14534);
not NOT1 (N14540, N14523);
nor NOR3 (N14541, N14533, N1541, N5996);
not NOT1 (N14542, N14529);
and AND2 (N14543, N14532, N11640);
not NOT1 (N14544, N14543);
not NOT1 (N14545, N14542);
nand NAND2 (N14546, N14541, N9233);
and AND3 (N14547, N14538, N10765, N14023);
buf BUF1 (N14548, N14544);
xor XOR2 (N14549, N14537, N7667);
or OR2 (N14550, N14547, N3466);
not NOT1 (N14551, N14550);
buf BUF1 (N14552, N14524);
buf BUF1 (N14553, N14548);
xor XOR2 (N14554, N14535, N13920);
xor XOR2 (N14555, N14553, N7667);
buf BUF1 (N14556, N14554);
not NOT1 (N14557, N14539);
or OR2 (N14558, N14549, N13426);
nor NOR4 (N14559, N14530, N8265, N2670, N13326);
xor XOR2 (N14560, N14546, N7634);
not NOT1 (N14561, N14545);
nand NAND4 (N14562, N14560, N6515, N4035, N8202);
buf BUF1 (N14563, N14557);
not NOT1 (N14564, N14556);
and AND2 (N14565, N14540, N9545);
not NOT1 (N14566, N14562);
nand NAND2 (N14567, N14566, N395);
buf BUF1 (N14568, N14555);
nor NOR2 (N14569, N14567, N10122);
nor NOR3 (N14570, N14563, N9094, N13417);
xor XOR2 (N14571, N14559, N4670);
and AND3 (N14572, N14552, N2817, N184);
nor NOR4 (N14573, N14551, N12555, N11647, N4278);
or OR2 (N14574, N14558, N10386);
not NOT1 (N14575, N14573);
or OR4 (N14576, N14571, N12001, N1105, N216);
and AND2 (N14577, N14569, N11369);
buf BUF1 (N14578, N14577);
not NOT1 (N14579, N14574);
nor NOR4 (N14580, N14564, N10837, N2389, N3146);
nor NOR2 (N14581, N14579, N5076);
nand NAND2 (N14582, N14581, N2053);
and AND4 (N14583, N14565, N189, N10696, N9360);
not NOT1 (N14584, N14572);
not NOT1 (N14585, N14568);
nor NOR3 (N14586, N14578, N3921, N12578);
nand NAND3 (N14587, N14570, N1054, N14485);
and AND2 (N14588, N14561, N8395);
or OR4 (N14589, N14585, N1169, N11169, N1030);
not NOT1 (N14590, N14576);
xor XOR2 (N14591, N14589, N1078);
nor NOR3 (N14592, N14582, N1865, N4880);
and AND2 (N14593, N14586, N4742);
xor XOR2 (N14594, N14592, N5809);
and AND4 (N14595, N14588, N3680, N8937, N13196);
or OR4 (N14596, N14590, N6838, N2985, N4216);
not NOT1 (N14597, N14587);
nand NAND2 (N14598, N14591, N8709);
nor NOR3 (N14599, N14595, N6680, N13019);
not NOT1 (N14600, N14593);
xor XOR2 (N14601, N14596, N5689);
and AND2 (N14602, N14601, N741);
or OR3 (N14603, N14600, N14447, N4788);
buf BUF1 (N14604, N14603);
nor NOR2 (N14605, N14597, N14222);
xor XOR2 (N14606, N14584, N12471);
or OR4 (N14607, N14594, N228, N6122, N7336);
not NOT1 (N14608, N14583);
nor NOR3 (N14609, N14608, N8378, N8748);
buf BUF1 (N14610, N14598);
not NOT1 (N14611, N14605);
nor NOR2 (N14612, N14602, N1027);
not NOT1 (N14613, N14599);
xor XOR2 (N14614, N14607, N4109);
nand NAND3 (N14615, N14611, N10374, N8585);
buf BUF1 (N14616, N14615);
and AND3 (N14617, N14614, N6816, N13574);
not NOT1 (N14618, N14613);
and AND4 (N14619, N14609, N3962, N6291, N8705);
and AND2 (N14620, N14606, N20);
or OR3 (N14621, N14610, N6580, N6138);
nand NAND2 (N14622, N14619, N3053);
or OR3 (N14623, N14575, N3891, N629);
or OR2 (N14624, N14618, N9652);
nand NAND3 (N14625, N14623, N5748, N2531);
and AND4 (N14626, N14621, N10026, N5147, N9683);
and AND4 (N14627, N14626, N3617, N11603, N14178);
or OR2 (N14628, N14612, N8827);
and AND4 (N14629, N14604, N617, N6092, N4436);
buf BUF1 (N14630, N14620);
nand NAND2 (N14631, N14627, N9721);
nor NOR2 (N14632, N14629, N14463);
nand NAND3 (N14633, N14632, N11587, N5290);
buf BUF1 (N14634, N14624);
xor XOR2 (N14635, N14580, N457);
nand NAND2 (N14636, N14635, N11255);
buf BUF1 (N14637, N14628);
not NOT1 (N14638, N14630);
or OR3 (N14639, N14634, N2364, N3181);
and AND2 (N14640, N14625, N7714);
buf BUF1 (N14641, N14631);
xor XOR2 (N14642, N14639, N11270);
not NOT1 (N14643, N14642);
nand NAND4 (N14644, N14643, N5613, N11340, N311);
or OR4 (N14645, N14636, N12999, N11226, N361);
buf BUF1 (N14646, N14637);
not NOT1 (N14647, N14646);
not NOT1 (N14648, N14633);
or OR4 (N14649, N14644, N11650, N2867, N3391);
xor XOR2 (N14650, N14649, N6708);
buf BUF1 (N14651, N14622);
not NOT1 (N14652, N14645);
not NOT1 (N14653, N14616);
or OR3 (N14654, N14652, N10769, N6206);
nand NAND2 (N14655, N14641, N11641);
nor NOR3 (N14656, N14648, N13703, N12687);
or OR2 (N14657, N14650, N1935);
nand NAND4 (N14658, N14656, N1967, N5705, N2960);
xor XOR2 (N14659, N14651, N6378);
and AND4 (N14660, N14638, N595, N2971, N10852);
or OR4 (N14661, N14617, N1518, N4297, N12593);
xor XOR2 (N14662, N14654, N1379);
not NOT1 (N14663, N14662);
buf BUF1 (N14664, N14661);
or OR2 (N14665, N14658, N6783);
or OR3 (N14666, N14640, N7544, N550);
nand NAND3 (N14667, N14666, N8074, N5275);
xor XOR2 (N14668, N14664, N1294);
and AND2 (N14669, N14668, N3574);
nor NOR3 (N14670, N14667, N3617, N10914);
buf BUF1 (N14671, N14669);
buf BUF1 (N14672, N14659);
and AND3 (N14673, N14647, N10536, N1574);
or OR3 (N14674, N14655, N4097, N6897);
xor XOR2 (N14675, N14663, N5642);
or OR3 (N14676, N14672, N13606, N12203);
and AND4 (N14677, N14674, N10201, N9568, N7170);
and AND2 (N14678, N14665, N10862);
xor XOR2 (N14679, N14676, N5164);
and AND4 (N14680, N14673, N8360, N170, N836);
nand NAND3 (N14681, N14675, N2041, N9733);
nor NOR4 (N14682, N14670, N2646, N3077, N12763);
buf BUF1 (N14683, N14653);
nand NAND3 (N14684, N14678, N1313, N11387);
xor XOR2 (N14685, N14677, N2282);
and AND2 (N14686, N14682, N3883);
nand NAND4 (N14687, N14681, N179, N8026, N6570);
nand NAND2 (N14688, N14657, N10003);
not NOT1 (N14689, N14684);
xor XOR2 (N14690, N14686, N7345);
buf BUF1 (N14691, N14690);
nor NOR3 (N14692, N14688, N13326, N11341);
nand NAND2 (N14693, N14687, N11419);
not NOT1 (N14694, N14692);
nand NAND4 (N14695, N14671, N8075, N14376, N9101);
nand NAND3 (N14696, N14679, N13237, N3913);
and AND2 (N14697, N14691, N10333);
or OR4 (N14698, N14697, N6857, N3582, N9906);
and AND2 (N14699, N14689, N5819);
xor XOR2 (N14700, N14699, N1738);
and AND2 (N14701, N14680, N13221);
not NOT1 (N14702, N14660);
nor NOR3 (N14703, N14700, N2467, N10770);
not NOT1 (N14704, N14701);
or OR4 (N14705, N14683, N1173, N12284, N9108);
nor NOR4 (N14706, N14702, N9425, N9559, N2123);
not NOT1 (N14707, N14706);
or OR3 (N14708, N14693, N1024, N8099);
or OR4 (N14709, N14696, N14143, N11096, N14524);
nand NAND4 (N14710, N14705, N3917, N4259, N6276);
nand NAND2 (N14711, N14685, N2242);
or OR3 (N14712, N14695, N10407, N8319);
nor NOR4 (N14713, N14709, N12010, N6375, N3480);
xor XOR2 (N14714, N14704, N8160);
nor NOR3 (N14715, N14713, N7302, N11813);
nand NAND3 (N14716, N14714, N2990, N5954);
nand NAND3 (N14717, N14707, N9822, N7321);
or OR4 (N14718, N14694, N8289, N14237, N7819);
buf BUF1 (N14719, N14711);
not NOT1 (N14720, N14718);
and AND2 (N14721, N14708, N12731);
or OR3 (N14722, N14717, N488, N13416);
not NOT1 (N14723, N14720);
nand NAND2 (N14724, N14723, N3947);
or OR2 (N14725, N14721, N13233);
nand NAND3 (N14726, N14698, N2428, N4462);
xor XOR2 (N14727, N14716, N3841);
nor NOR3 (N14728, N14727, N2188, N5622);
or OR2 (N14729, N14722, N7807);
and AND3 (N14730, N14712, N7236, N10746);
or OR3 (N14731, N14710, N8762, N3922);
xor XOR2 (N14732, N14725, N2159);
and AND4 (N14733, N14726, N10124, N11235, N13928);
and AND3 (N14734, N14731, N1743, N4534);
nand NAND2 (N14735, N14730, N14096);
or OR4 (N14736, N14734, N58, N9714, N8494);
or OR2 (N14737, N14724, N7141);
and AND3 (N14738, N14715, N3739, N5790);
not NOT1 (N14739, N14719);
nor NOR3 (N14740, N14737, N7795, N2052);
not NOT1 (N14741, N14732);
not NOT1 (N14742, N14729);
and AND2 (N14743, N14740, N13679);
or OR2 (N14744, N14742, N14274);
buf BUF1 (N14745, N14743);
or OR3 (N14746, N14741, N4370, N1836);
xor XOR2 (N14747, N14744, N12864);
xor XOR2 (N14748, N14735, N13040);
nor NOR3 (N14749, N14739, N455, N8287);
or OR2 (N14750, N14738, N10471);
xor XOR2 (N14751, N14703, N1128);
and AND2 (N14752, N14733, N1349);
and AND3 (N14753, N14736, N10099, N12876);
nand NAND4 (N14754, N14750, N1111, N7734, N1164);
and AND2 (N14755, N14747, N12351);
or OR3 (N14756, N14749, N181, N14473);
nand NAND3 (N14757, N14753, N920, N6271);
xor XOR2 (N14758, N14757, N2320);
nand NAND2 (N14759, N14728, N12326);
nand NAND3 (N14760, N14752, N6174, N7530);
buf BUF1 (N14761, N14758);
buf BUF1 (N14762, N14751);
not NOT1 (N14763, N14755);
not NOT1 (N14764, N14745);
not NOT1 (N14765, N14748);
nand NAND3 (N14766, N14746, N9990, N11664);
nor NOR3 (N14767, N14754, N8117, N1747);
buf BUF1 (N14768, N14763);
nand NAND4 (N14769, N14762, N10136, N1056, N13893);
or OR2 (N14770, N14768, N8244);
and AND3 (N14771, N14769, N927, N13944);
and AND3 (N14772, N14767, N10217, N9995);
buf BUF1 (N14773, N14759);
xor XOR2 (N14774, N14764, N12080);
nor NOR2 (N14775, N14773, N3536);
nor NOR4 (N14776, N14766, N1819, N9645, N7680);
or OR2 (N14777, N14775, N913);
nor NOR2 (N14778, N14770, N1783);
xor XOR2 (N14779, N14765, N8244);
and AND4 (N14780, N14778, N7646, N10405, N10329);
not NOT1 (N14781, N14777);
not NOT1 (N14782, N14761);
not NOT1 (N14783, N14774);
buf BUF1 (N14784, N14780);
and AND2 (N14785, N14779, N6551);
or OR4 (N14786, N14756, N4984, N10697, N3864);
buf BUF1 (N14787, N14776);
buf BUF1 (N14788, N14786);
xor XOR2 (N14789, N14784, N8349);
buf BUF1 (N14790, N14760);
nor NOR2 (N14791, N14789, N10339);
buf BUF1 (N14792, N14790);
and AND4 (N14793, N14772, N4399, N13540, N5626);
xor XOR2 (N14794, N14791, N3873);
or OR4 (N14795, N14794, N1170, N1392, N9654);
not NOT1 (N14796, N14785);
or OR2 (N14797, N14782, N5522);
buf BUF1 (N14798, N14787);
not NOT1 (N14799, N14788);
not NOT1 (N14800, N14799);
and AND3 (N14801, N14781, N9005, N2356);
buf BUF1 (N14802, N14801);
not NOT1 (N14803, N14797);
not NOT1 (N14804, N14798);
xor XOR2 (N14805, N14803, N717);
nor NOR4 (N14806, N14792, N13732, N235, N3849);
buf BUF1 (N14807, N14783);
and AND3 (N14808, N14807, N14637, N1633);
nand NAND2 (N14809, N14800, N11273);
nor NOR3 (N14810, N14802, N3739, N3284);
not NOT1 (N14811, N14771);
not NOT1 (N14812, N14796);
buf BUF1 (N14813, N14806);
nand NAND4 (N14814, N14812, N6600, N7474, N1369);
buf BUF1 (N14815, N14793);
nor NOR4 (N14816, N14795, N7228, N1843, N8033);
or OR2 (N14817, N14809, N10215);
buf BUF1 (N14818, N14817);
and AND4 (N14819, N14813, N13412, N2730, N9608);
not NOT1 (N14820, N14811);
or OR3 (N14821, N14820, N1628, N4697);
xor XOR2 (N14822, N14821, N1976);
and AND3 (N14823, N14818, N4700, N5926);
not NOT1 (N14824, N14810);
or OR2 (N14825, N14804, N5092);
xor XOR2 (N14826, N14824, N2449);
or OR4 (N14827, N14808, N8515, N7714, N11747);
buf BUF1 (N14828, N14827);
xor XOR2 (N14829, N14825, N9647);
nand NAND4 (N14830, N14822, N1401, N12255, N10520);
and AND4 (N14831, N14816, N4512, N8536, N10880);
or OR3 (N14832, N14829, N4915, N4928);
not NOT1 (N14833, N14830);
nor NOR3 (N14834, N14826, N10321, N6177);
and AND2 (N14835, N14805, N12247);
not NOT1 (N14836, N14835);
nor NOR2 (N14837, N14828, N10236);
nand NAND4 (N14838, N14837, N6799, N13463, N4515);
or OR4 (N14839, N14833, N2896, N10451, N13754);
or OR4 (N14840, N14838, N8541, N9756, N13898);
nor NOR2 (N14841, N14840, N6698);
or OR2 (N14842, N14841, N3540);
nand NAND2 (N14843, N14815, N13330);
xor XOR2 (N14844, N14823, N2513);
nor NOR3 (N14845, N14819, N5758, N3645);
not NOT1 (N14846, N14839);
nand NAND3 (N14847, N14814, N11775, N7872);
not NOT1 (N14848, N14832);
or OR2 (N14849, N14834, N14226);
buf BUF1 (N14850, N14847);
and AND3 (N14851, N14844, N1976, N1770);
xor XOR2 (N14852, N14842, N2904);
nor NOR4 (N14853, N14852, N13938, N13416, N12469);
not NOT1 (N14854, N14836);
or OR4 (N14855, N14850, N1205, N8552, N5669);
not NOT1 (N14856, N14855);
not NOT1 (N14857, N14845);
nand NAND4 (N14858, N14849, N2283, N30, N7841);
xor XOR2 (N14859, N14857, N10311);
xor XOR2 (N14860, N14846, N8125);
nand NAND3 (N14861, N14831, N11303, N8001);
nand NAND4 (N14862, N14854, N14635, N7787, N13124);
nor NOR2 (N14863, N14851, N4437);
or OR4 (N14864, N14848, N11323, N14301, N4782);
nand NAND3 (N14865, N14861, N10611, N11358);
not NOT1 (N14866, N14865);
and AND2 (N14867, N14860, N200);
not NOT1 (N14868, N14853);
xor XOR2 (N14869, N14858, N17);
nor NOR2 (N14870, N14856, N13004);
and AND3 (N14871, N14862, N6831, N8549);
and AND4 (N14872, N14871, N3927, N14144, N9400);
and AND2 (N14873, N14872, N3858);
or OR3 (N14874, N14864, N9173, N2729);
or OR2 (N14875, N14870, N10898);
and AND4 (N14876, N14874, N591, N7178, N1670);
buf BUF1 (N14877, N14868);
or OR2 (N14878, N14869, N6652);
nor NOR3 (N14879, N14877, N5426, N7309);
nor NOR3 (N14880, N14843, N11401, N4778);
xor XOR2 (N14881, N14879, N14280);
buf BUF1 (N14882, N14881);
or OR2 (N14883, N14882, N10980);
not NOT1 (N14884, N14867);
buf BUF1 (N14885, N14883);
and AND3 (N14886, N14884, N450, N14065);
nand NAND2 (N14887, N14863, N10834);
not NOT1 (N14888, N14885);
not NOT1 (N14889, N14875);
buf BUF1 (N14890, N14876);
nor NOR3 (N14891, N14873, N10201, N127);
nor NOR4 (N14892, N14891, N9795, N7630, N7789);
xor XOR2 (N14893, N14886, N7694);
buf BUF1 (N14894, N14887);
or OR3 (N14895, N14893, N6387, N14813);
not NOT1 (N14896, N14880);
not NOT1 (N14897, N14896);
not NOT1 (N14898, N14890);
not NOT1 (N14899, N14894);
or OR3 (N14900, N14897, N9152, N14787);
nand NAND3 (N14901, N14900, N7782, N10913);
nor NOR4 (N14902, N14888, N10591, N3967, N4488);
and AND2 (N14903, N14878, N2747);
or OR4 (N14904, N14903, N11767, N11004, N6236);
nand NAND3 (N14905, N14899, N6649, N5385);
or OR4 (N14906, N14859, N8453, N8616, N1986);
nor NOR3 (N14907, N14902, N9713, N11323);
nor NOR4 (N14908, N14906, N9639, N1948, N5225);
buf BUF1 (N14909, N14889);
and AND2 (N14910, N14866, N9018);
and AND2 (N14911, N14908, N425);
or OR2 (N14912, N14901, N6792);
nand NAND2 (N14913, N14898, N3034);
buf BUF1 (N14914, N14907);
xor XOR2 (N14915, N14895, N4609);
nand NAND2 (N14916, N14909, N9876);
buf BUF1 (N14917, N14912);
not NOT1 (N14918, N14892);
xor XOR2 (N14919, N14905, N2813);
or OR3 (N14920, N14910, N9374, N5177);
and AND4 (N14921, N14911, N5895, N2907, N2927);
nand NAND4 (N14922, N14919, N12048, N1520, N5275);
xor XOR2 (N14923, N14921, N7504);
not NOT1 (N14924, N14918);
and AND3 (N14925, N14917, N14577, N14314);
xor XOR2 (N14926, N14916, N2741);
buf BUF1 (N14927, N14925);
xor XOR2 (N14928, N14922, N5619);
or OR2 (N14929, N14913, N275);
not NOT1 (N14930, N14926);
buf BUF1 (N14931, N14920);
and AND2 (N14932, N14930, N636);
or OR2 (N14933, N14914, N3103);
and AND3 (N14934, N14928, N7429, N12141);
nand NAND2 (N14935, N14929, N11574);
not NOT1 (N14936, N14923);
buf BUF1 (N14937, N14932);
or OR3 (N14938, N14931, N6551, N9879);
and AND3 (N14939, N14936, N564, N14134);
xor XOR2 (N14940, N14937, N11890);
nand NAND2 (N14941, N14924, N8482);
and AND2 (N14942, N14934, N6318);
nand NAND2 (N14943, N14938, N9587);
or OR2 (N14944, N14941, N13499);
buf BUF1 (N14945, N14942);
and AND2 (N14946, N14927, N7835);
nor NOR3 (N14947, N14946, N4365, N14249);
nand NAND3 (N14948, N14904, N8040, N1012);
buf BUF1 (N14949, N14933);
and AND3 (N14950, N14947, N12329, N558);
not NOT1 (N14951, N14948);
xor XOR2 (N14952, N14939, N12994);
or OR4 (N14953, N14945, N8567, N14473, N5432);
and AND3 (N14954, N14950, N14703, N8193);
buf BUF1 (N14955, N14954);
xor XOR2 (N14956, N14952, N11124);
nand NAND4 (N14957, N14943, N6188, N11931, N1601);
buf BUF1 (N14958, N14944);
xor XOR2 (N14959, N14953, N13776);
and AND4 (N14960, N14955, N9082, N10529, N13730);
xor XOR2 (N14961, N14951, N95);
or OR3 (N14962, N14940, N4557, N9884);
not NOT1 (N14963, N14935);
or OR3 (N14964, N14960, N2533, N8634);
not NOT1 (N14965, N14962);
nor NOR3 (N14966, N14949, N1436, N10611);
nand NAND3 (N14967, N14966, N3191, N4284);
buf BUF1 (N14968, N14957);
not NOT1 (N14969, N14958);
xor XOR2 (N14970, N14964, N14484);
xor XOR2 (N14971, N14956, N1063);
xor XOR2 (N14972, N14963, N10441);
and AND3 (N14973, N14968, N14061, N11665);
buf BUF1 (N14974, N14973);
or OR2 (N14975, N14974, N2167);
nor NOR4 (N14976, N14915, N7107, N2284, N9521);
nor NOR4 (N14977, N14975, N1542, N9945, N14645);
nor NOR3 (N14978, N14977, N11972, N2364);
buf BUF1 (N14979, N14965);
xor XOR2 (N14980, N14978, N10295);
nor NOR2 (N14981, N14976, N21);
or OR4 (N14982, N14970, N7044, N4607, N7635);
nand NAND4 (N14983, N14979, N10587, N14332, N4484);
nor NOR4 (N14984, N14959, N3505, N9387, N14203);
buf BUF1 (N14985, N14981);
not NOT1 (N14986, N14969);
nand NAND2 (N14987, N14982, N9071);
and AND4 (N14988, N14986, N8172, N1272, N161);
and AND4 (N14989, N14988, N13255, N2303, N12584);
or OR3 (N14990, N14985, N13046, N9608);
nand NAND2 (N14991, N14967, N9034);
nor NOR3 (N14992, N14987, N7095, N8711);
xor XOR2 (N14993, N14989, N6191);
and AND2 (N14994, N14980, N3000);
nor NOR2 (N14995, N14991, N13178);
nor NOR4 (N14996, N14984, N7379, N7979, N212);
and AND4 (N14997, N14993, N7366, N1996, N1988);
xor XOR2 (N14998, N14992, N10748);
or OR4 (N14999, N14995, N10610, N14907, N5947);
xor XOR2 (N15000, N14971, N3388);
nand NAND3 (N15001, N14972, N8927, N9392);
nor NOR4 (N15002, N15000, N188, N7402, N9418);
nor NOR3 (N15003, N14996, N391, N14987);
not NOT1 (N15004, N14998);
and AND2 (N15005, N15002, N6858);
or OR4 (N15006, N15001, N4433, N5702, N2427);
nand NAND3 (N15007, N14994, N12806, N5046);
nor NOR3 (N15008, N14999, N5879, N4430);
nor NOR2 (N15009, N14961, N602);
not NOT1 (N15010, N14990);
or OR2 (N15011, N14983, N1132);
xor XOR2 (N15012, N15004, N2615);
nor NOR3 (N15013, N15010, N7787, N10504);
nand NAND3 (N15014, N15011, N5356, N4206);
and AND2 (N15015, N15007, N13339);
buf BUF1 (N15016, N15009);
xor XOR2 (N15017, N15015, N1826);
buf BUF1 (N15018, N15006);
or OR3 (N15019, N15016, N2571, N4371);
buf BUF1 (N15020, N15017);
buf BUF1 (N15021, N15018);
nor NOR3 (N15022, N15005, N830, N12940);
buf BUF1 (N15023, N15008);
and AND2 (N15024, N15019, N1506);
and AND2 (N15025, N15022, N14923);
not NOT1 (N15026, N15020);
nand NAND3 (N15027, N14997, N8432, N14465);
and AND4 (N15028, N15021, N13152, N10367, N6947);
and AND4 (N15029, N15023, N10855, N13045, N3032);
not NOT1 (N15030, N15029);
or OR3 (N15031, N15030, N13844, N2513);
not NOT1 (N15032, N15027);
xor XOR2 (N15033, N15032, N6944);
nand NAND2 (N15034, N15033, N10218);
or OR3 (N15035, N15031, N10741, N8686);
nand NAND3 (N15036, N15024, N6220, N1231);
nor NOR3 (N15037, N15013, N4263, N1920);
not NOT1 (N15038, N15036);
buf BUF1 (N15039, N15014);
xor XOR2 (N15040, N15003, N1905);
nor NOR4 (N15041, N15025, N4490, N10936, N6603);
and AND3 (N15042, N15037, N1335, N9975);
nand NAND2 (N15043, N15038, N14340);
or OR3 (N15044, N15040, N99, N5366);
nand NAND4 (N15045, N15044, N2557, N3432, N6479);
or OR2 (N15046, N15045, N10575);
and AND3 (N15047, N15041, N7589, N2264);
and AND2 (N15048, N15028, N7410);
and AND3 (N15049, N15047, N7398, N6173);
xor XOR2 (N15050, N15046, N11399);
buf BUF1 (N15051, N15050);
nor NOR2 (N15052, N15049, N4317);
buf BUF1 (N15053, N15042);
nand NAND3 (N15054, N15051, N5658, N14434);
or OR4 (N15055, N15034, N14044, N12125, N14373);
xor XOR2 (N15056, N15043, N9736);
nand NAND2 (N15057, N15026, N1836);
xor XOR2 (N15058, N15039, N11823);
and AND3 (N15059, N15055, N9365, N4519);
buf BUF1 (N15060, N15012);
nor NOR4 (N15061, N15052, N11716, N8917, N1326);
and AND3 (N15062, N15054, N10442, N4177);
nor NOR4 (N15063, N15061, N3876, N14730, N9650);
xor XOR2 (N15064, N15058, N1440);
xor XOR2 (N15065, N15053, N10357);
not NOT1 (N15066, N15064);
or OR2 (N15067, N15035, N10180);
buf BUF1 (N15068, N15060);
and AND4 (N15069, N15059, N13802, N13661, N3807);
buf BUF1 (N15070, N15066);
buf BUF1 (N15071, N15067);
nand NAND3 (N15072, N15063, N4156, N476);
and AND2 (N15073, N15062, N5244);
nor NOR2 (N15074, N15069, N7695);
nor NOR4 (N15075, N15065, N11432, N11542, N4041);
not NOT1 (N15076, N15056);
xor XOR2 (N15077, N15068, N5412);
nor NOR3 (N15078, N15057, N4964, N8395);
nand NAND2 (N15079, N15076, N6274);
nor NOR3 (N15080, N15078, N157, N13636);
buf BUF1 (N15081, N15080);
nand NAND4 (N15082, N15074, N9192, N8875, N4321);
buf BUF1 (N15083, N15070);
nand NAND2 (N15084, N15083, N1387);
nand NAND4 (N15085, N15079, N1188, N10844, N3948);
or OR3 (N15086, N15085, N3111, N4731);
and AND2 (N15087, N15082, N15010);
nor NOR4 (N15088, N15073, N6167, N7500, N13196);
and AND4 (N15089, N15072, N1083, N10527, N9062);
xor XOR2 (N15090, N15077, N12683);
and AND3 (N15091, N15086, N9357, N200);
and AND2 (N15092, N15084, N11259);
nor NOR3 (N15093, N15089, N2193, N2663);
xor XOR2 (N15094, N15071, N4115);
nand NAND4 (N15095, N15091, N6778, N3811, N277);
and AND4 (N15096, N15094, N5177, N14846, N12368);
buf BUF1 (N15097, N15095);
and AND4 (N15098, N15088, N14046, N5862, N5292);
xor XOR2 (N15099, N15087, N7761);
buf BUF1 (N15100, N15075);
buf BUF1 (N15101, N15096);
or OR2 (N15102, N15097, N10492);
buf BUF1 (N15103, N15098);
nor NOR3 (N15104, N15093, N12718, N11965);
xor XOR2 (N15105, N15100, N7318);
and AND3 (N15106, N15102, N1642, N5994);
not NOT1 (N15107, N15090);
nand NAND3 (N15108, N15105, N14985, N9142);
buf BUF1 (N15109, N15101);
buf BUF1 (N15110, N15048);
and AND2 (N15111, N15103, N7566);
buf BUF1 (N15112, N15099);
not NOT1 (N15113, N15081);
xor XOR2 (N15114, N15109, N7247);
nor NOR4 (N15115, N15110, N7437, N14598, N9924);
buf BUF1 (N15116, N15108);
or OR2 (N15117, N15092, N6311);
not NOT1 (N15118, N15113);
not NOT1 (N15119, N15116);
not NOT1 (N15120, N15114);
or OR4 (N15121, N15107, N5573, N3181, N3380);
nand NAND3 (N15122, N15119, N1346, N10358);
nand NAND3 (N15123, N15104, N12155, N5021);
and AND2 (N15124, N15112, N6168);
buf BUF1 (N15125, N15115);
xor XOR2 (N15126, N15123, N7969);
nand NAND2 (N15127, N15111, N999);
and AND3 (N15128, N15127, N9002, N4163);
or OR2 (N15129, N15106, N9745);
nand NAND4 (N15130, N15121, N6749, N11801, N11950);
buf BUF1 (N15131, N15124);
and AND4 (N15132, N15126, N6515, N11199, N2761);
xor XOR2 (N15133, N15129, N2827);
buf BUF1 (N15134, N15117);
nor NOR4 (N15135, N15134, N13520, N9500, N14348);
not NOT1 (N15136, N15131);
and AND2 (N15137, N15135, N11112);
xor XOR2 (N15138, N15130, N10981);
or OR4 (N15139, N15137, N9451, N1119, N1188);
nand NAND2 (N15140, N15132, N3754);
nor NOR2 (N15141, N15118, N10248);
or OR3 (N15142, N15138, N6878, N14763);
not NOT1 (N15143, N15120);
nand NAND3 (N15144, N15122, N13915, N13682);
or OR2 (N15145, N15133, N4556);
xor XOR2 (N15146, N15144, N10480);
and AND4 (N15147, N15142, N14356, N13911, N14681);
buf BUF1 (N15148, N15141);
xor XOR2 (N15149, N15146, N7987);
nor NOR2 (N15150, N15149, N3660);
not NOT1 (N15151, N15140);
or OR2 (N15152, N15139, N8670);
not NOT1 (N15153, N15128);
nand NAND4 (N15154, N15147, N895, N857, N7330);
or OR2 (N15155, N15153, N4526);
xor XOR2 (N15156, N15150, N14106);
nor NOR4 (N15157, N15145, N7745, N11990, N3854);
nor NOR4 (N15158, N15157, N8367, N5783, N8374);
xor XOR2 (N15159, N15158, N11294);
buf BUF1 (N15160, N15151);
or OR3 (N15161, N15143, N5285, N8133);
and AND4 (N15162, N15154, N13245, N11384, N1710);
and AND3 (N15163, N15161, N4452, N13938);
nor NOR4 (N15164, N15156, N8311, N10007, N10885);
not NOT1 (N15165, N15159);
or OR2 (N15166, N15136, N13034);
buf BUF1 (N15167, N15164);
or OR3 (N15168, N15152, N5844, N9099);
or OR2 (N15169, N15166, N1993);
or OR3 (N15170, N15165, N5602, N14997);
and AND4 (N15171, N15155, N12581, N5577, N3070);
buf BUF1 (N15172, N15160);
or OR3 (N15173, N15168, N5439, N15165);
nor NOR4 (N15174, N15162, N2882, N9945, N11455);
buf BUF1 (N15175, N15163);
not NOT1 (N15176, N15172);
nand NAND2 (N15177, N15171, N14511);
and AND3 (N15178, N15175, N3391, N3308);
or OR4 (N15179, N15176, N1828, N12948, N2211);
nand NAND3 (N15180, N15179, N12419, N13851);
and AND4 (N15181, N15125, N5578, N12882, N12456);
buf BUF1 (N15182, N15181);
or OR4 (N15183, N15167, N3362, N14220, N5735);
xor XOR2 (N15184, N15173, N6851);
nor NOR2 (N15185, N15178, N11717);
nor NOR2 (N15186, N15174, N14293);
nor NOR4 (N15187, N15180, N3552, N7928, N13026);
nand NAND3 (N15188, N15185, N7561, N8726);
buf BUF1 (N15189, N15184);
xor XOR2 (N15190, N15188, N2077);
or OR2 (N15191, N15189, N3496);
buf BUF1 (N15192, N15177);
nor NOR2 (N15193, N15190, N10143);
nor NOR3 (N15194, N15183, N6565, N11655);
and AND2 (N15195, N15169, N10528);
xor XOR2 (N15196, N15182, N4931);
and AND4 (N15197, N15186, N3943, N13902, N6686);
nand NAND4 (N15198, N15170, N5699, N8142, N927);
and AND2 (N15199, N15196, N13876);
xor XOR2 (N15200, N15193, N14514);
nor NOR2 (N15201, N15148, N11129);
xor XOR2 (N15202, N15200, N3374);
or OR4 (N15203, N15195, N7763, N11269, N5754);
nor NOR3 (N15204, N15199, N6276, N6471);
buf BUF1 (N15205, N15187);
xor XOR2 (N15206, N15204, N5122);
xor XOR2 (N15207, N15197, N11310);
and AND2 (N15208, N15203, N9633);
and AND2 (N15209, N15208, N192);
xor XOR2 (N15210, N15191, N1862);
nand NAND2 (N15211, N15192, N575);
nor NOR3 (N15212, N15210, N2031, N1189);
buf BUF1 (N15213, N15201);
nor NOR3 (N15214, N15207, N9049, N4949);
and AND4 (N15215, N15214, N6906, N12138, N4425);
nor NOR3 (N15216, N15209, N2451, N12236);
and AND4 (N15217, N15211, N732, N6582, N9663);
or OR2 (N15218, N15216, N6358);
buf BUF1 (N15219, N15217);
not NOT1 (N15220, N15218);
nand NAND4 (N15221, N15194, N13261, N428, N2667);
nand NAND2 (N15222, N15206, N5785);
and AND4 (N15223, N15220, N469, N2533, N3999);
or OR4 (N15224, N15205, N1450, N10148, N9670);
not NOT1 (N15225, N15215);
or OR4 (N15226, N15213, N5228, N5277, N1618);
xor XOR2 (N15227, N15222, N7857);
nand NAND3 (N15228, N15202, N1827, N3584);
nand NAND4 (N15229, N15219, N6649, N2663, N11925);
buf BUF1 (N15230, N15229);
nand NAND4 (N15231, N15221, N9934, N6832, N1793);
xor XOR2 (N15232, N15223, N14558);
nor NOR3 (N15233, N15226, N12520, N3295);
xor XOR2 (N15234, N15227, N3976);
nand NAND2 (N15235, N15198, N9467);
nor NOR3 (N15236, N15232, N14195, N15096);
and AND2 (N15237, N15225, N4870);
xor XOR2 (N15238, N15212, N4549);
nand NAND3 (N15239, N15235, N8725, N1820);
nand NAND3 (N15240, N15231, N10296, N4788);
nor NOR4 (N15241, N15240, N11702, N1056, N3095);
nand NAND4 (N15242, N15239, N770, N6869, N11501);
not NOT1 (N15243, N15242);
nor NOR3 (N15244, N15230, N278, N7315);
and AND3 (N15245, N15237, N2487, N5027);
and AND2 (N15246, N15234, N6634);
buf BUF1 (N15247, N15244);
and AND3 (N15248, N15245, N6015, N4929);
xor XOR2 (N15249, N15247, N5031);
xor XOR2 (N15250, N15243, N9202);
nor NOR3 (N15251, N15250, N14119, N10148);
nand NAND3 (N15252, N15233, N3385, N13175);
nor NOR3 (N15253, N15228, N11326, N10552);
nand NAND2 (N15254, N15238, N11982);
or OR2 (N15255, N15251, N6741);
nor NOR3 (N15256, N15253, N1571, N5649);
xor XOR2 (N15257, N15256, N3516);
buf BUF1 (N15258, N15224);
not NOT1 (N15259, N15241);
or OR3 (N15260, N15254, N10425, N12611);
xor XOR2 (N15261, N15259, N2235);
nor NOR2 (N15262, N15260, N4509);
nand NAND3 (N15263, N15252, N14551, N5686);
nand NAND2 (N15264, N15257, N1930);
and AND3 (N15265, N15262, N15008, N9247);
or OR3 (N15266, N15264, N1958, N606);
nor NOR4 (N15267, N15246, N1368, N5758, N1381);
xor XOR2 (N15268, N15249, N7889);
and AND3 (N15269, N15248, N12241, N14338);
xor XOR2 (N15270, N15265, N1574);
nand NAND2 (N15271, N15270, N14423);
buf BUF1 (N15272, N15263);
or OR4 (N15273, N15267, N9126, N1235, N12832);
buf BUF1 (N15274, N15269);
buf BUF1 (N15275, N15255);
buf BUF1 (N15276, N15271);
and AND4 (N15277, N15268, N8123, N12959, N13532);
and AND2 (N15278, N15275, N5905);
and AND3 (N15279, N15274, N6218, N7401);
nand NAND4 (N15280, N15278, N9812, N2569, N1196);
buf BUF1 (N15281, N15261);
and AND3 (N15282, N15273, N8353, N13452);
nor NOR4 (N15283, N15266, N3347, N2959, N12461);
buf BUF1 (N15284, N15281);
buf BUF1 (N15285, N15282);
and AND3 (N15286, N15285, N13394, N4124);
nor NOR4 (N15287, N15279, N2761, N5992, N12047);
nor NOR4 (N15288, N15272, N13696, N11865, N12607);
or OR3 (N15289, N15287, N11759, N776);
nor NOR2 (N15290, N15236, N13616);
not NOT1 (N15291, N15280);
nor NOR4 (N15292, N15283, N6939, N57, N838);
xor XOR2 (N15293, N15277, N8792);
xor XOR2 (N15294, N15293, N725);
or OR2 (N15295, N15286, N1199);
nand NAND4 (N15296, N15290, N11048, N2771, N13877);
or OR3 (N15297, N15276, N12354, N6139);
and AND3 (N15298, N15294, N1088, N9626);
and AND4 (N15299, N15288, N1568, N5089, N10328);
buf BUF1 (N15300, N15291);
buf BUF1 (N15301, N15299);
and AND4 (N15302, N15300, N14999, N7244, N8178);
or OR3 (N15303, N15258, N10895, N1286);
not NOT1 (N15304, N15297);
or OR2 (N15305, N15289, N13276);
not NOT1 (N15306, N15295);
not NOT1 (N15307, N15306);
not NOT1 (N15308, N15284);
nor NOR4 (N15309, N15303, N12702, N7965, N4447);
or OR4 (N15310, N15305, N10450, N4782, N13427);
not NOT1 (N15311, N15298);
xor XOR2 (N15312, N15310, N14606);
nand NAND4 (N15313, N15308, N13446, N5700, N4890);
nand NAND2 (N15314, N15309, N4866);
nor NOR2 (N15315, N15301, N3833);
not NOT1 (N15316, N15313);
nor NOR3 (N15317, N15315, N7031, N5795);
not NOT1 (N15318, N15312);
nand NAND4 (N15319, N15302, N10604, N14111, N3288);
nor NOR2 (N15320, N15318, N5978);
xor XOR2 (N15321, N15307, N5694);
xor XOR2 (N15322, N15296, N15014);
not NOT1 (N15323, N15314);
nand NAND4 (N15324, N15316, N2591, N2666, N397);
xor XOR2 (N15325, N15322, N8310);
buf BUF1 (N15326, N15324);
not NOT1 (N15327, N15320);
and AND3 (N15328, N15321, N10287, N9102);
or OR4 (N15329, N15304, N14445, N5491, N6495);
nand NAND3 (N15330, N15328, N9, N15188);
xor XOR2 (N15331, N15329, N9735);
xor XOR2 (N15332, N15325, N13046);
not NOT1 (N15333, N15323);
not NOT1 (N15334, N15326);
and AND4 (N15335, N15330, N1108, N9211, N6134);
xor XOR2 (N15336, N15292, N9559);
not NOT1 (N15337, N15317);
nor NOR4 (N15338, N15336, N7804, N11109, N1401);
buf BUF1 (N15339, N15337);
buf BUF1 (N15340, N15339);
nand NAND2 (N15341, N15340, N2271);
nor NOR4 (N15342, N15319, N3903, N3333, N11117);
and AND2 (N15343, N15333, N7774);
or OR3 (N15344, N15327, N8206, N88);
or OR3 (N15345, N15341, N3665, N8131);
nand NAND4 (N15346, N15334, N13704, N2367, N15149);
and AND4 (N15347, N15331, N10365, N2355, N6491);
not NOT1 (N15348, N15346);
not NOT1 (N15349, N15345);
and AND3 (N15350, N15343, N12740, N278);
nand NAND2 (N15351, N15338, N663);
xor XOR2 (N15352, N15335, N9873);
and AND2 (N15353, N15348, N8625);
and AND2 (N15354, N15350, N13373);
nor NOR2 (N15355, N15347, N5158);
not NOT1 (N15356, N15353);
not NOT1 (N15357, N15351);
buf BUF1 (N15358, N15352);
or OR4 (N15359, N15342, N15042, N1928, N5790);
nor NOR3 (N15360, N15356, N10233, N458);
nor NOR4 (N15361, N15360, N8807, N8031, N12265);
nand NAND3 (N15362, N15354, N9109, N4695);
or OR3 (N15363, N15344, N6786, N3878);
nor NOR4 (N15364, N15358, N8415, N1286, N15178);
buf BUF1 (N15365, N15357);
or OR2 (N15366, N15364, N5468);
xor XOR2 (N15367, N15363, N13817);
or OR3 (N15368, N15362, N13683, N4750);
not NOT1 (N15369, N15355);
and AND3 (N15370, N15311, N11805, N10619);
not NOT1 (N15371, N15368);
buf BUF1 (N15372, N15332);
nor NOR4 (N15373, N15372, N9718, N8400, N6835);
and AND3 (N15374, N15349, N14943, N5707);
and AND2 (N15375, N15359, N4293);
or OR3 (N15376, N15365, N14507, N10430);
not NOT1 (N15377, N15376);
nor NOR4 (N15378, N15366, N3289, N1362, N9632);
not NOT1 (N15379, N15374);
nor NOR3 (N15380, N15369, N1296, N6451);
buf BUF1 (N15381, N15370);
or OR3 (N15382, N15375, N6741, N7719);
xor XOR2 (N15383, N15377, N3617);
buf BUF1 (N15384, N15361);
buf BUF1 (N15385, N15367);
xor XOR2 (N15386, N15373, N6794);
or OR4 (N15387, N15385, N9886, N9922, N2666);
buf BUF1 (N15388, N15378);
or OR4 (N15389, N15381, N1853, N1922, N6483);
or OR4 (N15390, N15384, N4180, N14737, N14842);
buf BUF1 (N15391, N15389);
not NOT1 (N15392, N15371);
xor XOR2 (N15393, N15387, N12962);
not NOT1 (N15394, N15388);
not NOT1 (N15395, N15379);
nor NOR2 (N15396, N15382, N6118);
nand NAND3 (N15397, N15395, N3101, N175);
not NOT1 (N15398, N15380);
nand NAND2 (N15399, N15394, N8077);
xor XOR2 (N15400, N15397, N7224);
and AND2 (N15401, N15383, N14184);
nor NOR3 (N15402, N15386, N766, N12269);
and AND2 (N15403, N15398, N9831);
or OR2 (N15404, N15402, N11081);
xor XOR2 (N15405, N15393, N3476);
xor XOR2 (N15406, N15401, N1114);
nand NAND4 (N15407, N15399, N44, N6578, N11472);
or OR3 (N15408, N15392, N6891, N12530);
nor NOR4 (N15409, N15407, N6173, N5245, N9746);
not NOT1 (N15410, N15406);
nand NAND2 (N15411, N15405, N3470);
xor XOR2 (N15412, N15403, N2425);
nand NAND4 (N15413, N15410, N6918, N3428, N98);
or OR2 (N15414, N15408, N1905);
buf BUF1 (N15415, N15391);
or OR4 (N15416, N15400, N11497, N7804, N4893);
xor XOR2 (N15417, N15414, N15074);
nand NAND4 (N15418, N15412, N6059, N3228, N6615);
and AND3 (N15419, N15390, N8166, N5931);
nand NAND2 (N15420, N15413, N9512);
and AND3 (N15421, N15396, N12509, N8720);
not NOT1 (N15422, N15420);
and AND4 (N15423, N15422, N1436, N608, N2794);
and AND4 (N15424, N15419, N418, N6663, N10911);
not NOT1 (N15425, N15418);
buf BUF1 (N15426, N15416);
and AND4 (N15427, N15415, N4318, N3022, N13712);
not NOT1 (N15428, N15424);
or OR2 (N15429, N15417, N9139);
nand NAND4 (N15430, N15428, N13829, N2959, N5252);
or OR2 (N15431, N15430, N8315);
nand NAND2 (N15432, N15421, N11741);
buf BUF1 (N15433, N15425);
nor NOR4 (N15434, N15427, N13084, N2291, N11771);
or OR3 (N15435, N15423, N5804, N12780);
buf BUF1 (N15436, N15432);
or OR2 (N15437, N15409, N12427);
not NOT1 (N15438, N15426);
or OR2 (N15439, N15411, N1543);
nor NOR4 (N15440, N15435, N7360, N7530, N10182);
or OR4 (N15441, N15440, N6640, N1944, N1206);
xor XOR2 (N15442, N15404, N157);
nor NOR2 (N15443, N15434, N12407);
or OR3 (N15444, N15439, N6749, N8046);
and AND3 (N15445, N15437, N3330, N12923);
nand NAND3 (N15446, N15444, N13605, N6377);
nor NOR3 (N15447, N15433, N11719, N2650);
xor XOR2 (N15448, N15429, N8176);
buf BUF1 (N15449, N15448);
buf BUF1 (N15450, N15438);
or OR4 (N15451, N15441, N9440, N15175, N3157);
and AND2 (N15452, N15436, N5019);
nand NAND2 (N15453, N15447, N15259);
not NOT1 (N15454, N15450);
xor XOR2 (N15455, N15452, N4494);
xor XOR2 (N15456, N15453, N10462);
or OR2 (N15457, N15449, N14278);
and AND2 (N15458, N15442, N2634);
nand NAND4 (N15459, N15445, N9738, N8620, N4889);
xor XOR2 (N15460, N15454, N5430);
xor XOR2 (N15461, N15455, N13204);
or OR2 (N15462, N15443, N10176);
buf BUF1 (N15463, N15451);
nor NOR4 (N15464, N15457, N2552, N11647, N2448);
xor XOR2 (N15465, N15459, N5137);
buf BUF1 (N15466, N15456);
nand NAND2 (N15467, N15461, N10929);
xor XOR2 (N15468, N15446, N6848);
or OR2 (N15469, N15458, N12078);
and AND4 (N15470, N15463, N7786, N1717, N2774);
xor XOR2 (N15471, N15467, N2100);
and AND2 (N15472, N15466, N564);
and AND3 (N15473, N15471, N8117, N9589);
or OR4 (N15474, N15470, N3869, N8515, N4175);
buf BUF1 (N15475, N15465);
or OR3 (N15476, N15431, N12017, N6479);
buf BUF1 (N15477, N15474);
buf BUF1 (N15478, N15469);
and AND3 (N15479, N15468, N5992, N3480);
nor NOR4 (N15480, N15460, N13682, N9063, N7);
nand NAND2 (N15481, N15473, N13822);
not NOT1 (N15482, N15472);
buf BUF1 (N15483, N15475);
xor XOR2 (N15484, N15479, N445);
not NOT1 (N15485, N15480);
not NOT1 (N15486, N15485);
buf BUF1 (N15487, N15478);
nor NOR4 (N15488, N15481, N11898, N13718, N6753);
and AND4 (N15489, N15484, N12060, N8040, N6598);
and AND2 (N15490, N15483, N3327);
not NOT1 (N15491, N15462);
or OR2 (N15492, N15482, N5917);
not NOT1 (N15493, N15476);
nand NAND3 (N15494, N15489, N6833, N281);
not NOT1 (N15495, N15487);
buf BUF1 (N15496, N15477);
not NOT1 (N15497, N15488);
xor XOR2 (N15498, N15486, N12699);
xor XOR2 (N15499, N15498, N8255);
or OR4 (N15500, N15494, N8414, N8139, N9895);
not NOT1 (N15501, N15497);
or OR3 (N15502, N15490, N314, N307);
or OR4 (N15503, N15501, N1576, N10193, N14600);
buf BUF1 (N15504, N15464);
or OR2 (N15505, N15495, N1839);
or OR4 (N15506, N15492, N5271, N8418, N9373);
not NOT1 (N15507, N15500);
and AND3 (N15508, N15499, N6963, N13351);
nand NAND4 (N15509, N15505, N3364, N1165, N262);
nand NAND4 (N15510, N15508, N10282, N7603, N5174);
not NOT1 (N15511, N15506);
buf BUF1 (N15512, N15511);
or OR2 (N15513, N15512, N10911);
or OR3 (N15514, N15493, N2237, N5297);
nor NOR2 (N15515, N15514, N796);
and AND3 (N15516, N15502, N2986, N1027);
not NOT1 (N15517, N15510);
nor NOR4 (N15518, N15516, N10057, N13016, N6502);
not NOT1 (N15519, N15517);
buf BUF1 (N15520, N15504);
buf BUF1 (N15521, N15491);
and AND2 (N15522, N15496, N12393);
not NOT1 (N15523, N15519);
nor NOR3 (N15524, N15503, N8681, N1647);
and AND4 (N15525, N15523, N15353, N2715, N1875);
nand NAND2 (N15526, N15515, N13631);
or OR4 (N15527, N15507, N15170, N13407, N14041);
xor XOR2 (N15528, N15524, N15177);
not NOT1 (N15529, N15509);
nand NAND3 (N15530, N15527, N3029, N9656);
nand NAND4 (N15531, N15513, N12094, N5280, N12139);
or OR2 (N15532, N15525, N2901);
nand NAND2 (N15533, N15521, N3969);
buf BUF1 (N15534, N15522);
buf BUF1 (N15535, N15529);
or OR2 (N15536, N15520, N9753);
nand NAND3 (N15537, N15534, N986, N14211);
buf BUF1 (N15538, N15537);
buf BUF1 (N15539, N15531);
xor XOR2 (N15540, N15518, N6283);
and AND3 (N15541, N15533, N7345, N1461);
or OR4 (N15542, N15539, N12929, N11909, N3446);
buf BUF1 (N15543, N15532);
nand NAND4 (N15544, N15526, N14022, N764, N11007);
nand NAND3 (N15545, N15528, N2895, N13170);
nand NAND4 (N15546, N15535, N1143, N4252, N12724);
xor XOR2 (N15547, N15538, N1779);
and AND3 (N15548, N15536, N5868, N7140);
xor XOR2 (N15549, N15541, N12317);
nor NOR3 (N15550, N15530, N957, N7665);
nor NOR2 (N15551, N15548, N10422);
nor NOR2 (N15552, N15551, N14980);
or OR4 (N15553, N15542, N5174, N13422, N7145);
not NOT1 (N15554, N15543);
buf BUF1 (N15555, N15553);
not NOT1 (N15556, N15550);
buf BUF1 (N15557, N15555);
nor NOR3 (N15558, N15552, N7148, N6273);
buf BUF1 (N15559, N15558);
not NOT1 (N15560, N15557);
xor XOR2 (N15561, N15540, N14213);
and AND2 (N15562, N15547, N8563);
or OR4 (N15563, N15545, N691, N13712, N11711);
not NOT1 (N15564, N15560);
nor NOR3 (N15565, N15561, N9390, N4685);
xor XOR2 (N15566, N15564, N2184);
buf BUF1 (N15567, N15562);
buf BUF1 (N15568, N15554);
buf BUF1 (N15569, N15568);
not NOT1 (N15570, N15563);
buf BUF1 (N15571, N15567);
not NOT1 (N15572, N15569);
nand NAND4 (N15573, N15544, N14575, N8049, N4209);
buf BUF1 (N15574, N15565);
and AND4 (N15575, N15572, N5601, N9896, N6805);
xor XOR2 (N15576, N15556, N12639);
nor NOR3 (N15577, N15573, N8279, N13662);
buf BUF1 (N15578, N15570);
or OR3 (N15579, N15575, N2143, N7845);
buf BUF1 (N15580, N15579);
or OR2 (N15581, N15580, N605);
buf BUF1 (N15582, N15559);
or OR3 (N15583, N15546, N14573, N13927);
not NOT1 (N15584, N15581);
not NOT1 (N15585, N15566);
or OR4 (N15586, N15574, N10369, N4740, N7448);
nor NOR3 (N15587, N15586, N2981, N11339);
nand NAND4 (N15588, N15571, N2169, N156, N8338);
not NOT1 (N15589, N15583);
nor NOR3 (N15590, N15589, N956, N15385);
nor NOR4 (N15591, N15587, N4464, N4069, N4487);
xor XOR2 (N15592, N15591, N13857);
xor XOR2 (N15593, N15576, N13602);
and AND2 (N15594, N15592, N6937);
nand NAND2 (N15595, N15584, N10799);
nor NOR2 (N15596, N15588, N7332);
or OR3 (N15597, N15593, N11319, N9128);
and AND3 (N15598, N15582, N14560, N7042);
and AND2 (N15599, N15590, N8212);
or OR3 (N15600, N15549, N8768, N10095);
nand NAND2 (N15601, N15599, N3268);
nand NAND4 (N15602, N15596, N4555, N7053, N6874);
buf BUF1 (N15603, N15598);
not NOT1 (N15604, N15602);
nand NAND3 (N15605, N15595, N8032, N1713);
and AND3 (N15606, N15600, N12699, N13518);
nor NOR4 (N15607, N15577, N6635, N12491, N7209);
buf BUF1 (N15608, N15607);
xor XOR2 (N15609, N15605, N8452);
not NOT1 (N15610, N15606);
nor NOR2 (N15611, N15597, N2943);
nor NOR4 (N15612, N15594, N10001, N7685, N1616);
buf BUF1 (N15613, N15585);
xor XOR2 (N15614, N15608, N4828);
nor NOR3 (N15615, N15611, N13845, N1834);
and AND3 (N15616, N15614, N4738, N4444);
or OR2 (N15617, N15604, N4956);
nand NAND3 (N15618, N15615, N8181, N4813);
nor NOR3 (N15619, N15617, N3650, N8476);
buf BUF1 (N15620, N15613);
xor XOR2 (N15621, N15578, N9899);
not NOT1 (N15622, N15619);
nor NOR3 (N15623, N15618, N12171, N422);
xor XOR2 (N15624, N15603, N12098);
not NOT1 (N15625, N15609);
nand NAND2 (N15626, N15621, N15233);
nor NOR2 (N15627, N15610, N8972);
buf BUF1 (N15628, N15612);
xor XOR2 (N15629, N15624, N12087);
or OR4 (N15630, N15623, N6949, N6088, N14410);
xor XOR2 (N15631, N15628, N6426);
xor XOR2 (N15632, N15627, N7675);
buf BUF1 (N15633, N15616);
or OR4 (N15634, N15631, N10346, N13160, N6546);
nor NOR4 (N15635, N15634, N10300, N6304, N7105);
or OR2 (N15636, N15626, N9923);
or OR4 (N15637, N15632, N9668, N12981, N7);
xor XOR2 (N15638, N15636, N6466);
nor NOR4 (N15639, N15601, N11845, N7453, N11951);
not NOT1 (N15640, N15633);
and AND3 (N15641, N15622, N2844, N9123);
nand NAND2 (N15642, N15630, N2255);
nor NOR3 (N15643, N15637, N1721, N1548);
nand NAND2 (N15644, N15639, N4220);
nor NOR3 (N15645, N15643, N9288, N7180);
or OR2 (N15646, N15638, N6888);
nor NOR2 (N15647, N15644, N15131);
or OR4 (N15648, N15620, N9918, N9663, N12858);
or OR4 (N15649, N15646, N13917, N14681, N2355);
not NOT1 (N15650, N15641);
xor XOR2 (N15651, N15648, N7313);
and AND3 (N15652, N15625, N15368, N3361);
nand NAND4 (N15653, N15645, N375, N8711, N12894);
nand NAND3 (N15654, N15647, N9632, N9817);
xor XOR2 (N15655, N15651, N11315);
xor XOR2 (N15656, N15654, N5765);
buf BUF1 (N15657, N15640);
nor NOR3 (N15658, N15656, N13142, N6916);
and AND3 (N15659, N15642, N10303, N8252);
xor XOR2 (N15660, N15649, N9690);
and AND3 (N15661, N15650, N5163, N7393);
and AND4 (N15662, N15657, N10269, N6300, N2945);
xor XOR2 (N15663, N15658, N10561);
not NOT1 (N15664, N15653);
or OR3 (N15665, N15664, N11383, N9265);
and AND4 (N15666, N15661, N10454, N15037, N5317);
buf BUF1 (N15667, N15659);
xor XOR2 (N15668, N15662, N2913);
buf BUF1 (N15669, N15666);
and AND2 (N15670, N15652, N2955);
or OR2 (N15671, N15655, N416);
nor NOR3 (N15672, N15629, N10545, N15582);
xor XOR2 (N15673, N15635, N6685);
nor NOR2 (N15674, N15665, N204);
buf BUF1 (N15675, N15668);
or OR2 (N15676, N15667, N9118);
nor NOR2 (N15677, N15671, N10655);
not NOT1 (N15678, N15660);
not NOT1 (N15679, N15678);
and AND4 (N15680, N15663, N8657, N1660, N9624);
not NOT1 (N15681, N15672);
and AND2 (N15682, N15675, N6400);
not NOT1 (N15683, N15680);
or OR4 (N15684, N15679, N7660, N13293, N1160);
buf BUF1 (N15685, N15676);
buf BUF1 (N15686, N15674);
buf BUF1 (N15687, N15685);
xor XOR2 (N15688, N15670, N9985);
nor NOR2 (N15689, N15686, N202);
and AND3 (N15690, N15677, N11396, N2758);
buf BUF1 (N15691, N15669);
or OR2 (N15692, N15689, N8677);
not NOT1 (N15693, N15682);
or OR3 (N15694, N15687, N8135, N10528);
and AND2 (N15695, N15688, N6474);
not NOT1 (N15696, N15690);
buf BUF1 (N15697, N15691);
or OR2 (N15698, N15683, N7740);
xor XOR2 (N15699, N15694, N410);
nand NAND3 (N15700, N15692, N13404, N14309);
and AND4 (N15701, N15699, N8449, N13107, N12434);
xor XOR2 (N15702, N15695, N254);
nor NOR2 (N15703, N15673, N8372);
buf BUF1 (N15704, N15698);
xor XOR2 (N15705, N15704, N4929);
xor XOR2 (N15706, N15705, N11738);
nor NOR4 (N15707, N15684, N9684, N13143, N15588);
buf BUF1 (N15708, N15701);
or OR4 (N15709, N15706, N7208, N14783, N4841);
not NOT1 (N15710, N15700);
buf BUF1 (N15711, N15703);
xor XOR2 (N15712, N15697, N11224);
nand NAND3 (N15713, N15702, N8537, N2464);
xor XOR2 (N15714, N15713, N10525);
nand NAND2 (N15715, N15709, N14353);
xor XOR2 (N15716, N15707, N6785);
and AND3 (N15717, N15710, N7990, N4491);
nand NAND2 (N15718, N15693, N8298);
and AND4 (N15719, N15716, N9406, N9417, N14759);
xor XOR2 (N15720, N15714, N3770);
nor NOR4 (N15721, N15712, N2390, N4832, N12938);
nor NOR4 (N15722, N15721, N8383, N12579, N15646);
buf BUF1 (N15723, N15717);
or OR2 (N15724, N15719, N15433);
xor XOR2 (N15725, N15696, N250);
buf BUF1 (N15726, N15681);
nand NAND4 (N15727, N15725, N3505, N5850, N5183);
buf BUF1 (N15728, N15724);
and AND2 (N15729, N15715, N5843);
buf BUF1 (N15730, N15727);
xor XOR2 (N15731, N15726, N10809);
or OR4 (N15732, N15711, N4867, N12855, N1116);
not NOT1 (N15733, N15731);
not NOT1 (N15734, N15723);
or OR4 (N15735, N15722, N4293, N4359, N11354);
not NOT1 (N15736, N15718);
xor XOR2 (N15737, N15732, N1007);
not NOT1 (N15738, N15720);
or OR2 (N15739, N15734, N166);
or OR3 (N15740, N15729, N2866, N10128);
not NOT1 (N15741, N15708);
not NOT1 (N15742, N15740);
and AND4 (N15743, N15736, N13693, N7813, N13823);
nand NAND3 (N15744, N15730, N2714, N58);
xor XOR2 (N15745, N15733, N1542);
not NOT1 (N15746, N15738);
nor NOR4 (N15747, N15739, N13903, N9123, N7808);
xor XOR2 (N15748, N15728, N12727);
xor XOR2 (N15749, N15741, N8884);
and AND2 (N15750, N15749, N10602);
xor XOR2 (N15751, N15737, N14728);
or OR2 (N15752, N15745, N310);
nand NAND4 (N15753, N15748, N10631, N2066, N5668);
not NOT1 (N15754, N15735);
xor XOR2 (N15755, N15750, N3567);
nand NAND3 (N15756, N15751, N6219, N238);
buf BUF1 (N15757, N15753);
nand NAND3 (N15758, N15743, N5321, N9111);
not NOT1 (N15759, N15746);
and AND3 (N15760, N15756, N5210, N11009);
nor NOR2 (N15761, N15755, N9683);
not NOT1 (N15762, N15760);
not NOT1 (N15763, N15762);
xor XOR2 (N15764, N15759, N1632);
and AND3 (N15765, N15752, N13469, N15139);
not NOT1 (N15766, N15754);
and AND3 (N15767, N15757, N2015, N4609);
nand NAND4 (N15768, N15767, N4995, N225, N12569);
nand NAND4 (N15769, N15744, N459, N7096, N3290);
buf BUF1 (N15770, N15761);
not NOT1 (N15771, N15742);
nand NAND4 (N15772, N15766, N8385, N7635, N39);
not NOT1 (N15773, N15768);
nor NOR2 (N15774, N15763, N6974);
buf BUF1 (N15775, N15747);
not NOT1 (N15776, N15764);
buf BUF1 (N15777, N15774);
nand NAND2 (N15778, N15769, N10988);
nand NAND3 (N15779, N15758, N4678, N4363);
buf BUF1 (N15780, N15772);
not NOT1 (N15781, N15780);
nand NAND3 (N15782, N15770, N3301, N9770);
xor XOR2 (N15783, N15777, N10962);
nor NOR2 (N15784, N15778, N14366);
nor NOR3 (N15785, N15773, N13149, N2230);
nand NAND3 (N15786, N15782, N13443, N13260);
not NOT1 (N15787, N15771);
buf BUF1 (N15788, N15779);
not NOT1 (N15789, N15787);
nand NAND2 (N15790, N15785, N15024);
or OR3 (N15791, N15790, N9144, N9045);
xor XOR2 (N15792, N15783, N10213);
buf BUF1 (N15793, N15786);
xor XOR2 (N15794, N15793, N7716);
buf BUF1 (N15795, N15794);
and AND4 (N15796, N15792, N8706, N5994, N14887);
or OR4 (N15797, N15788, N12458, N7973, N11360);
and AND2 (N15798, N15795, N14830);
or OR3 (N15799, N15798, N39, N8234);
nand NAND3 (N15800, N15784, N12880, N6273);
nor NOR3 (N15801, N15797, N7991, N6219);
and AND3 (N15802, N15776, N9463, N10167);
nand NAND4 (N15803, N15801, N1730, N4579, N10088);
buf BUF1 (N15804, N15800);
and AND3 (N15805, N15799, N2149, N11631);
not NOT1 (N15806, N15791);
not NOT1 (N15807, N15803);
and AND2 (N15808, N15781, N4846);
or OR2 (N15809, N15806, N884);
and AND3 (N15810, N15802, N13419, N1805);
or OR4 (N15811, N15765, N13899, N13619, N11101);
and AND3 (N15812, N15807, N11061, N417);
and AND4 (N15813, N15775, N8666, N10532, N77);
or OR4 (N15814, N15809, N1723, N8464, N7037);
buf BUF1 (N15815, N15814);
not NOT1 (N15816, N15813);
nor NOR2 (N15817, N15789, N7812);
and AND4 (N15818, N15811, N9250, N4951, N4640);
and AND4 (N15819, N15817, N4375, N3960, N13186);
not NOT1 (N15820, N15796);
nand NAND4 (N15821, N15804, N5116, N8044, N12706);
or OR3 (N15822, N15805, N7567, N2385);
nor NOR3 (N15823, N15822, N9094, N13868);
or OR3 (N15824, N15823, N13700, N9924);
not NOT1 (N15825, N15821);
not NOT1 (N15826, N15810);
not NOT1 (N15827, N15812);
not NOT1 (N15828, N15819);
buf BUF1 (N15829, N15818);
buf BUF1 (N15830, N15824);
and AND4 (N15831, N15827, N10941, N274, N4830);
nor NOR4 (N15832, N15828, N15284, N12951, N9582);
nand NAND4 (N15833, N15830, N6298, N1828, N2402);
nor NOR3 (N15834, N15829, N1955, N13104);
and AND3 (N15835, N15831, N10928, N15632);
nor NOR3 (N15836, N15816, N2772, N8583);
nand NAND4 (N15837, N15825, N13798, N5348, N8465);
and AND3 (N15838, N15835, N11841, N5230);
xor XOR2 (N15839, N15834, N14880);
or OR2 (N15840, N15839, N3141);
nand NAND3 (N15841, N15826, N8307, N9861);
not NOT1 (N15842, N15841);
nor NOR4 (N15843, N15838, N3958, N2239, N6526);
nand NAND2 (N15844, N15808, N12958);
or OR2 (N15845, N15836, N5765);
buf BUF1 (N15846, N15844);
nor NOR4 (N15847, N15815, N9576, N12178, N13324);
nand NAND2 (N15848, N15842, N14915);
nor NOR4 (N15849, N15848, N5696, N2147, N9228);
or OR4 (N15850, N15845, N8074, N7113, N3263);
and AND4 (N15851, N15843, N10077, N10885, N6223);
and AND2 (N15852, N15820, N14147);
not NOT1 (N15853, N15851);
xor XOR2 (N15854, N15850, N40);
and AND3 (N15855, N15853, N13135, N12605);
not NOT1 (N15856, N15854);
buf BUF1 (N15857, N15856);
nand NAND2 (N15858, N15857, N13316);
or OR3 (N15859, N15832, N13115, N10134);
nand NAND2 (N15860, N15846, N9154);
nand NAND4 (N15861, N15847, N8101, N4639, N8969);
or OR4 (N15862, N15855, N8152, N303, N11608);
xor XOR2 (N15863, N15860, N864);
xor XOR2 (N15864, N15852, N14353);
not NOT1 (N15865, N15840);
and AND3 (N15866, N15865, N5166, N5613);
nor NOR2 (N15867, N15858, N10976);
nand NAND3 (N15868, N15833, N3160, N15076);
buf BUF1 (N15869, N15867);
buf BUF1 (N15870, N15864);
and AND3 (N15871, N15868, N9047, N462);
or OR3 (N15872, N15837, N6205, N6940);
not NOT1 (N15873, N15863);
xor XOR2 (N15874, N15869, N7379);
or OR3 (N15875, N15874, N2598, N577);
and AND2 (N15876, N15873, N14460);
buf BUF1 (N15877, N15870);
nor NOR4 (N15878, N15876, N3243, N9774, N2539);
or OR4 (N15879, N15859, N4041, N7951, N8893);
nor NOR3 (N15880, N15866, N2475, N12740);
buf BUF1 (N15881, N15849);
nand NAND4 (N15882, N15877, N7201, N9029, N4293);
or OR2 (N15883, N15871, N3648);
nor NOR2 (N15884, N15879, N8766);
xor XOR2 (N15885, N15882, N7513);
buf BUF1 (N15886, N15878);
not NOT1 (N15887, N15880);
xor XOR2 (N15888, N15885, N9352);
or OR4 (N15889, N15862, N86, N8977, N11677);
xor XOR2 (N15890, N15883, N1991);
nand NAND2 (N15891, N15887, N13308);
nor NOR3 (N15892, N15891, N9717, N1644);
not NOT1 (N15893, N15861);
nor NOR2 (N15894, N15886, N1341);
or OR3 (N15895, N15889, N14998, N7382);
not NOT1 (N15896, N15892);
not NOT1 (N15897, N15893);
nand NAND3 (N15898, N15872, N4436, N11383);
xor XOR2 (N15899, N15898, N5517);
buf BUF1 (N15900, N15881);
and AND2 (N15901, N15896, N13733);
and AND2 (N15902, N15894, N13030);
buf BUF1 (N15903, N15899);
not NOT1 (N15904, N15902);
not NOT1 (N15905, N15888);
nand NAND3 (N15906, N15895, N6365, N7140);
or OR2 (N15907, N15904, N561);
or OR3 (N15908, N15903, N3683, N5645);
buf BUF1 (N15909, N15907);
nor NOR2 (N15910, N15900, N3883);
buf BUF1 (N15911, N15905);
and AND3 (N15912, N15901, N984, N7284);
nand NAND2 (N15913, N15906, N809);
xor XOR2 (N15914, N15884, N8538);
and AND2 (N15915, N15914, N1163);
buf BUF1 (N15916, N15915);
buf BUF1 (N15917, N15916);
not NOT1 (N15918, N15912);
xor XOR2 (N15919, N15909, N14210);
nor NOR4 (N15920, N15910, N11879, N7430, N6318);
buf BUF1 (N15921, N15919);
or OR2 (N15922, N15917, N1730);
xor XOR2 (N15923, N15911, N6263);
and AND2 (N15924, N15897, N4853);
and AND2 (N15925, N15913, N2386);
buf BUF1 (N15926, N15875);
buf BUF1 (N15927, N15921);
xor XOR2 (N15928, N15922, N347);
or OR3 (N15929, N15926, N13209, N10930);
xor XOR2 (N15930, N15927, N9990);
and AND3 (N15931, N15908, N13933, N853);
buf BUF1 (N15932, N15920);
and AND2 (N15933, N15932, N4223);
xor XOR2 (N15934, N15890, N120);
nand NAND4 (N15935, N15931, N907, N13889, N12871);
not NOT1 (N15936, N15929);
nor NOR2 (N15937, N15930, N6692);
and AND2 (N15938, N15934, N4679);
and AND2 (N15939, N15923, N6765);
xor XOR2 (N15940, N15937, N10838);
not NOT1 (N15941, N15938);
nor NOR4 (N15942, N15935, N13268, N1547, N10824);
buf BUF1 (N15943, N15936);
nand NAND2 (N15944, N15925, N11687);
nand NAND3 (N15945, N15943, N14389, N4155);
nand NAND3 (N15946, N15940, N14175, N9692);
and AND3 (N15947, N15946, N2434, N1232);
xor XOR2 (N15948, N15939, N3793);
and AND4 (N15949, N15942, N4393, N12804, N4715);
and AND3 (N15950, N15924, N14761, N5361);
not NOT1 (N15951, N15941);
and AND4 (N15952, N15949, N8788, N15123, N10123);
xor XOR2 (N15953, N15950, N14693);
and AND4 (N15954, N15933, N3582, N4748, N8876);
or OR2 (N15955, N15944, N6231);
buf BUF1 (N15956, N15945);
and AND4 (N15957, N15956, N14988, N10228, N14560);
not NOT1 (N15958, N15954);
nand NAND4 (N15959, N15951, N5606, N4988, N11496);
buf BUF1 (N15960, N15918);
buf BUF1 (N15961, N15947);
not NOT1 (N15962, N15928);
buf BUF1 (N15963, N15962);
nand NAND2 (N15964, N15963, N586);
nor NOR4 (N15965, N15964, N14469, N4784, N10608);
and AND4 (N15966, N15953, N5694, N14392, N1478);
and AND3 (N15967, N15948, N5110, N8632);
xor XOR2 (N15968, N15965, N3675);
not NOT1 (N15969, N15968);
or OR2 (N15970, N15960, N5740);
or OR2 (N15971, N15969, N3189);
or OR2 (N15972, N15957, N7975);
buf BUF1 (N15973, N15971);
or OR4 (N15974, N15972, N4998, N9529, N575);
and AND3 (N15975, N15967, N12583, N14007);
nor NOR3 (N15976, N15966, N10480, N6088);
buf BUF1 (N15977, N15959);
or OR4 (N15978, N15952, N15697, N12127, N297);
not NOT1 (N15979, N15973);
or OR4 (N15980, N15978, N13321, N3622, N761);
nand NAND4 (N15981, N15979, N8158, N9072, N6173);
or OR3 (N15982, N15955, N9434, N6340);
not NOT1 (N15983, N15976);
not NOT1 (N15984, N15975);
and AND4 (N15985, N15982, N11576, N10046, N10477);
buf BUF1 (N15986, N15974);
xor XOR2 (N15987, N15958, N30);
and AND2 (N15988, N15980, N12677);
buf BUF1 (N15989, N15984);
or OR3 (N15990, N15988, N13510, N7515);
buf BUF1 (N15991, N15961);
nand NAND3 (N15992, N15983, N12721, N2288);
not NOT1 (N15993, N15992);
buf BUF1 (N15994, N15970);
and AND4 (N15995, N15987, N11615, N951, N10257);
not NOT1 (N15996, N15986);
not NOT1 (N15997, N15991);
not NOT1 (N15998, N15996);
nand NAND3 (N15999, N15993, N13096, N12063);
and AND4 (N16000, N15989, N15116, N13972, N6371);
or OR3 (N16001, N15999, N8761, N4684);
and AND3 (N16002, N15998, N6365, N13454);
and AND4 (N16003, N15981, N3721, N6340, N11380);
not NOT1 (N16004, N16000);
nor NOR3 (N16005, N15990, N4724, N6110);
not NOT1 (N16006, N16002);
nor NOR3 (N16007, N16006, N2016, N6078);
buf BUF1 (N16008, N16005);
xor XOR2 (N16009, N16001, N11874);
xor XOR2 (N16010, N15994, N7741);
or OR3 (N16011, N15985, N13225, N15797);
or OR4 (N16012, N16007, N4686, N10755, N3977);
not NOT1 (N16013, N15997);
and AND3 (N16014, N16012, N3021, N4604);
not NOT1 (N16015, N16004);
and AND4 (N16016, N16010, N13314, N14568, N14488);
or OR4 (N16017, N16008, N13610, N15840, N13556);
or OR4 (N16018, N16016, N11473, N2100, N5257);
or OR2 (N16019, N16013, N7787);
xor XOR2 (N16020, N16017, N12520);
not NOT1 (N16021, N16019);
nand NAND3 (N16022, N16011, N8437, N14902);
xor XOR2 (N16023, N16021, N951);
or OR4 (N16024, N16023, N8343, N10366, N10960);
or OR4 (N16025, N16014, N10450, N11822, N9471);
xor XOR2 (N16026, N16024, N1948);
and AND4 (N16027, N15995, N12438, N718, N9413);
or OR2 (N16028, N16020, N11360);
not NOT1 (N16029, N16018);
nor NOR4 (N16030, N16022, N10872, N5908, N5126);
nor NOR4 (N16031, N16025, N13729, N13110, N7368);
or OR4 (N16032, N16009, N101, N6748, N691);
or OR2 (N16033, N16028, N12240);
nand NAND3 (N16034, N16031, N11089, N15918);
buf BUF1 (N16035, N16026);
not NOT1 (N16036, N16027);
and AND3 (N16037, N16034, N15503, N8022);
and AND2 (N16038, N16035, N2841);
buf BUF1 (N16039, N16032);
xor XOR2 (N16040, N15977, N11702);
xor XOR2 (N16041, N16029, N6448);
or OR4 (N16042, N16015, N2748, N10114, N5655);
xor XOR2 (N16043, N16039, N7000);
and AND4 (N16044, N16038, N6789, N9558, N3999);
not NOT1 (N16045, N16042);
xor XOR2 (N16046, N16043, N10928);
xor XOR2 (N16047, N16036, N2216);
not NOT1 (N16048, N16040);
buf BUF1 (N16049, N16044);
not NOT1 (N16050, N16047);
not NOT1 (N16051, N16037);
buf BUF1 (N16052, N16030);
buf BUF1 (N16053, N16041);
not NOT1 (N16054, N16050);
or OR3 (N16055, N16048, N8612, N12879);
nor NOR2 (N16056, N16052, N6079);
or OR4 (N16057, N16045, N2483, N12153, N5066);
not NOT1 (N16058, N16054);
xor XOR2 (N16059, N16051, N14209);
buf BUF1 (N16060, N16057);
or OR3 (N16061, N16056, N15883, N8944);
nor NOR3 (N16062, N16033, N5219, N1889);
xor XOR2 (N16063, N16046, N13795);
xor XOR2 (N16064, N16060, N12444);
or OR4 (N16065, N16003, N11082, N1282, N13760);
xor XOR2 (N16066, N16064, N3408);
buf BUF1 (N16067, N16053);
or OR2 (N16068, N16067, N589);
xor XOR2 (N16069, N16055, N8912);
nand NAND2 (N16070, N16059, N11731);
buf BUF1 (N16071, N16069);
and AND2 (N16072, N16066, N7138);
buf BUF1 (N16073, N16068);
buf BUF1 (N16074, N16072);
not NOT1 (N16075, N16070);
or OR4 (N16076, N16062, N12693, N10796, N8994);
nor NOR3 (N16077, N16076, N3179, N1206);
not NOT1 (N16078, N16071);
or OR2 (N16079, N16078, N824);
nand NAND3 (N16080, N16049, N2621, N13143);
and AND4 (N16081, N16061, N9508, N1288, N7029);
not NOT1 (N16082, N16081);
or OR2 (N16083, N16058, N15559);
or OR3 (N16084, N16080, N10610, N5715);
and AND2 (N16085, N16065, N14665);
nor NOR3 (N16086, N16073, N11972, N7882);
not NOT1 (N16087, N16082);
xor XOR2 (N16088, N16087, N2938);
not NOT1 (N16089, N16079);
buf BUF1 (N16090, N16088);
not NOT1 (N16091, N16063);
buf BUF1 (N16092, N16084);
buf BUF1 (N16093, N16089);
nand NAND2 (N16094, N16093, N4005);
nand NAND4 (N16095, N16086, N9609, N5918, N11620);
nand NAND3 (N16096, N16077, N15980, N11344);
nand NAND4 (N16097, N16075, N7357, N5367, N7496);
buf BUF1 (N16098, N16085);
not NOT1 (N16099, N16097);
not NOT1 (N16100, N16098);
not NOT1 (N16101, N16095);
or OR3 (N16102, N16094, N9002, N14849);
or OR4 (N16103, N16099, N8449, N16039, N3848);
and AND3 (N16104, N16083, N11370, N5751);
not NOT1 (N16105, N16090);
nor NOR2 (N16106, N16100, N13926);
buf BUF1 (N16107, N16101);
and AND4 (N16108, N16102, N11255, N6358, N14055);
or OR2 (N16109, N16107, N16059);
or OR3 (N16110, N16092, N3020, N999);
and AND2 (N16111, N16096, N5540);
not NOT1 (N16112, N16091);
buf BUF1 (N16113, N16106);
and AND3 (N16114, N16108, N10620, N5285);
not NOT1 (N16115, N16113);
xor XOR2 (N16116, N16111, N9518);
buf BUF1 (N16117, N16109);
buf BUF1 (N16118, N16115);
and AND3 (N16119, N16118, N7047, N12355);
xor XOR2 (N16120, N16116, N1937);
nand NAND3 (N16121, N16074, N14532, N5740);
buf BUF1 (N16122, N16117);
and AND3 (N16123, N16121, N1876, N15538);
xor XOR2 (N16124, N16105, N9801);
nor NOR4 (N16125, N16103, N3881, N6330, N11519);
and AND4 (N16126, N16125, N4783, N3511, N12261);
buf BUF1 (N16127, N16110);
and AND4 (N16128, N16104, N11776, N7473, N7421);
buf BUF1 (N16129, N16114);
nand NAND4 (N16130, N16129, N2967, N5427, N12985);
not NOT1 (N16131, N16128);
nor NOR4 (N16132, N16126, N4110, N6584, N3678);
buf BUF1 (N16133, N16127);
or OR4 (N16134, N16132, N14731, N4592, N15309);
and AND4 (N16135, N16130, N6078, N15911, N11852);
nor NOR4 (N16136, N16131, N5774, N1525, N387);
nand NAND3 (N16137, N16119, N8539, N4709);
buf BUF1 (N16138, N16136);
not NOT1 (N16139, N16133);
nor NOR3 (N16140, N16120, N805, N5465);
and AND3 (N16141, N16137, N2027, N13084);
xor XOR2 (N16142, N16123, N3822);
nand NAND4 (N16143, N16134, N6182, N12914, N9909);
nand NAND2 (N16144, N16122, N1921);
nand NAND2 (N16145, N16135, N11388);
nand NAND3 (N16146, N16124, N13822, N16117);
and AND3 (N16147, N16138, N8031, N4503);
or OR2 (N16148, N16146, N8255);
buf BUF1 (N16149, N16142);
and AND4 (N16150, N16140, N1015, N1409, N227);
nand NAND4 (N16151, N16150, N7305, N7363, N9085);
or OR3 (N16152, N16112, N4840, N12744);
and AND4 (N16153, N16145, N13406, N13747, N16066);
nor NOR2 (N16154, N16149, N3699);
not NOT1 (N16155, N16154);
and AND2 (N16156, N16139, N12347);
and AND2 (N16157, N16151, N12472);
nor NOR2 (N16158, N16153, N8001);
xor XOR2 (N16159, N16157, N7074);
not NOT1 (N16160, N16156);
and AND2 (N16161, N16148, N5274);
buf BUF1 (N16162, N16143);
or OR4 (N16163, N16141, N15320, N9799, N9357);
nor NOR2 (N16164, N16147, N14354);
xor XOR2 (N16165, N16162, N12868);
xor XOR2 (N16166, N16164, N2069);
or OR2 (N16167, N16161, N15341);
xor XOR2 (N16168, N16159, N727);
nand NAND2 (N16169, N16158, N10597);
buf BUF1 (N16170, N16163);
not NOT1 (N16171, N16169);
nor NOR2 (N16172, N16170, N13390);
or OR2 (N16173, N16160, N7411);
not NOT1 (N16174, N16168);
and AND2 (N16175, N16167, N10470);
not NOT1 (N16176, N16152);
and AND4 (N16177, N16171, N5604, N4003, N2906);
or OR4 (N16178, N16174, N12644, N16131, N2682);
or OR3 (N16179, N16144, N6717, N10730);
not NOT1 (N16180, N16179);
nand NAND2 (N16181, N16165, N586);
xor XOR2 (N16182, N16173, N14581);
xor XOR2 (N16183, N16181, N1136);
xor XOR2 (N16184, N16175, N12134);
not NOT1 (N16185, N16180);
nor NOR3 (N16186, N16155, N10012, N15987);
and AND2 (N16187, N16186, N7210);
nand NAND3 (N16188, N16183, N11523, N8837);
xor XOR2 (N16189, N16177, N13005);
nand NAND2 (N16190, N16172, N7730);
and AND4 (N16191, N16166, N12045, N10051, N11641);
buf BUF1 (N16192, N16190);
nand NAND2 (N16193, N16184, N15886);
nor NOR3 (N16194, N16185, N13128, N4742);
not NOT1 (N16195, N16188);
buf BUF1 (N16196, N16194);
xor XOR2 (N16197, N16189, N2195);
nand NAND3 (N16198, N16187, N7615, N3239);
xor XOR2 (N16199, N16195, N6411);
buf BUF1 (N16200, N16197);
or OR4 (N16201, N16196, N5478, N2024, N15458);
not NOT1 (N16202, N16191);
nand NAND3 (N16203, N16200, N6437, N6112);
not NOT1 (N16204, N16182);
and AND3 (N16205, N16193, N3576, N14003);
nand NAND3 (N16206, N16201, N5297, N2300);
buf BUF1 (N16207, N16206);
nand NAND3 (N16208, N16199, N14073, N5473);
xor XOR2 (N16209, N16203, N4176);
not NOT1 (N16210, N16205);
not NOT1 (N16211, N16209);
xor XOR2 (N16212, N16192, N13025);
nor NOR4 (N16213, N16212, N5156, N9421, N4313);
and AND2 (N16214, N16178, N12825);
xor XOR2 (N16215, N16176, N5503);
and AND4 (N16216, N16215, N13520, N8355, N2668);
not NOT1 (N16217, N16214);
buf BUF1 (N16218, N16204);
nand NAND4 (N16219, N16202, N14492, N9753, N7817);
buf BUF1 (N16220, N16198);
nor NOR3 (N16221, N16216, N6816, N12006);
and AND4 (N16222, N16220, N13286, N2009, N8762);
nand NAND4 (N16223, N16208, N802, N3888, N9429);
nand NAND2 (N16224, N16213, N13447);
or OR4 (N16225, N16211, N10866, N597, N15581);
or OR4 (N16226, N16223, N15680, N16190, N13196);
not NOT1 (N16227, N16207);
and AND4 (N16228, N16227, N3636, N6850, N12018);
xor XOR2 (N16229, N16228, N15587);
not NOT1 (N16230, N16225);
or OR2 (N16231, N16224, N3908);
not NOT1 (N16232, N16221);
not NOT1 (N16233, N16230);
nand NAND2 (N16234, N16232, N4594);
and AND2 (N16235, N16218, N5207);
and AND2 (N16236, N16231, N5514);
nor NOR4 (N16237, N16222, N5494, N12462, N12191);
nor NOR4 (N16238, N16219, N5307, N14586, N818);
buf BUF1 (N16239, N16236);
or OR4 (N16240, N16234, N7539, N3427, N13810);
not NOT1 (N16241, N16229);
not NOT1 (N16242, N16235);
xor XOR2 (N16243, N16240, N2024);
buf BUF1 (N16244, N16243);
nor NOR4 (N16245, N16244, N2105, N8676, N14017);
buf BUF1 (N16246, N16233);
nor NOR4 (N16247, N16241, N11480, N3806, N10202);
xor XOR2 (N16248, N16242, N6892);
nor NOR3 (N16249, N16247, N5967, N2045);
and AND3 (N16250, N16246, N6628, N1897);
buf BUF1 (N16251, N16210);
buf BUF1 (N16252, N16217);
nor NOR3 (N16253, N16249, N10303, N8198);
and AND2 (N16254, N16248, N6571);
and AND4 (N16255, N16253, N10562, N1330, N11568);
nor NOR2 (N16256, N16226, N11714);
buf BUF1 (N16257, N16250);
nor NOR3 (N16258, N16252, N9451, N9227);
not NOT1 (N16259, N16258);
and AND4 (N16260, N16239, N13029, N13825, N14932);
not NOT1 (N16261, N16237);
xor XOR2 (N16262, N16256, N1108);
xor XOR2 (N16263, N16254, N15161);
nand NAND3 (N16264, N16255, N3423, N966);
buf BUF1 (N16265, N16261);
xor XOR2 (N16266, N16257, N5242);
and AND4 (N16267, N16265, N8380, N5692, N13881);
nor NOR3 (N16268, N16259, N2763, N301);
xor XOR2 (N16269, N16264, N3382);
buf BUF1 (N16270, N16268);
or OR3 (N16271, N16269, N8697, N14843);
buf BUF1 (N16272, N16263);
nor NOR4 (N16273, N16238, N8786, N12006, N6999);
nor NOR3 (N16274, N16262, N7396, N7815);
nor NOR3 (N16275, N16251, N13918, N15632);
or OR3 (N16276, N16270, N1573, N9577);
and AND2 (N16277, N16266, N360);
nor NOR2 (N16278, N16274, N6951);
xor XOR2 (N16279, N16275, N15139);
nand NAND2 (N16280, N16272, N8892);
or OR2 (N16281, N16245, N14310);
xor XOR2 (N16282, N16276, N484);
buf BUF1 (N16283, N16267);
xor XOR2 (N16284, N16283, N8005);
xor XOR2 (N16285, N16273, N14599);
or OR3 (N16286, N16285, N1420, N14714);
or OR4 (N16287, N16281, N11778, N5738, N12636);
nor NOR3 (N16288, N16284, N9683, N9490);
nand NAND3 (N16289, N16282, N12413, N6397);
and AND3 (N16290, N16288, N11437, N13889);
and AND2 (N16291, N16277, N8205);
nor NOR4 (N16292, N16291, N4640, N13828, N13327);
buf BUF1 (N16293, N16279);
and AND2 (N16294, N16280, N7078);
nand NAND2 (N16295, N16293, N1165);
or OR3 (N16296, N16294, N14521, N16214);
xor XOR2 (N16297, N16286, N11407);
nor NOR2 (N16298, N16292, N6350);
nand NAND2 (N16299, N16278, N6078);
not NOT1 (N16300, N16287);
xor XOR2 (N16301, N16300, N3687);
buf BUF1 (N16302, N16296);
xor XOR2 (N16303, N16289, N14473);
or OR2 (N16304, N16298, N14803);
or OR2 (N16305, N16295, N5095);
buf BUF1 (N16306, N16297);
not NOT1 (N16307, N16271);
nor NOR2 (N16308, N16305, N15892);
buf BUF1 (N16309, N16290);
xor XOR2 (N16310, N16302, N12032);
buf BUF1 (N16311, N16260);
buf BUF1 (N16312, N16306);
xor XOR2 (N16313, N16309, N891);
not NOT1 (N16314, N16307);
buf BUF1 (N16315, N16301);
or OR4 (N16316, N16303, N7404, N1947, N10261);
and AND2 (N16317, N16304, N1762);
buf BUF1 (N16318, N16316);
or OR3 (N16319, N16313, N5500, N1669);
nor NOR3 (N16320, N16312, N8035, N11860);
nand NAND3 (N16321, N16308, N15953, N9123);
nand NAND3 (N16322, N16319, N7578, N13254);
not NOT1 (N16323, N16310);
or OR2 (N16324, N16311, N3696);
buf BUF1 (N16325, N16318);
nand NAND4 (N16326, N16314, N6634, N1332, N6806);
xor XOR2 (N16327, N16299, N8677);
nor NOR3 (N16328, N16326, N12935, N4985);
nand NAND4 (N16329, N16324, N7728, N4610, N1570);
nand NAND4 (N16330, N16323, N8954, N6885, N10097);
or OR3 (N16331, N16327, N140, N53);
buf BUF1 (N16332, N16320);
not NOT1 (N16333, N16329);
nor NOR4 (N16334, N16321, N3757, N9962, N12685);
nor NOR2 (N16335, N16332, N1155);
buf BUF1 (N16336, N16325);
xor XOR2 (N16337, N16335, N8522);
or OR2 (N16338, N16331, N2190);
xor XOR2 (N16339, N16317, N8665);
and AND3 (N16340, N16330, N3213, N9852);
buf BUF1 (N16341, N16340);
and AND3 (N16342, N16315, N8653, N11382);
buf BUF1 (N16343, N16342);
buf BUF1 (N16344, N16338);
xor XOR2 (N16345, N16333, N10050);
buf BUF1 (N16346, N16328);
nor NOR4 (N16347, N16322, N3025, N5945, N4900);
nor NOR3 (N16348, N16341, N8801, N7593);
and AND4 (N16349, N16337, N3653, N8570, N7841);
nand NAND4 (N16350, N16345, N6982, N1016, N14896);
nand NAND3 (N16351, N16346, N6416, N15547);
buf BUF1 (N16352, N16334);
not NOT1 (N16353, N16347);
nor NOR4 (N16354, N16348, N14106, N1656, N5037);
and AND4 (N16355, N16354, N13659, N12135, N13480);
and AND3 (N16356, N16349, N6306, N858);
not NOT1 (N16357, N16339);
or OR4 (N16358, N16355, N7185, N13129, N12915);
or OR3 (N16359, N16353, N12032, N3155);
nand NAND2 (N16360, N16344, N542);
xor XOR2 (N16361, N16358, N11426);
or OR3 (N16362, N16350, N15899, N338);
not NOT1 (N16363, N16362);
and AND2 (N16364, N16359, N15250);
buf BUF1 (N16365, N16364);
buf BUF1 (N16366, N16365);
nand NAND3 (N16367, N16366, N15107, N12297);
and AND4 (N16368, N16363, N15950, N12809, N4543);
not NOT1 (N16369, N16361);
and AND2 (N16370, N16357, N10491);
nand NAND3 (N16371, N16356, N16212, N10084);
nor NOR2 (N16372, N16368, N1794);
and AND2 (N16373, N16369, N9268);
or OR3 (N16374, N16367, N5635, N8786);
buf BUF1 (N16375, N16360);
buf BUF1 (N16376, N16336);
or OR3 (N16377, N16376, N12358, N3067);
buf BUF1 (N16378, N16373);
and AND2 (N16379, N16377, N5520);
buf BUF1 (N16380, N16351);
or OR4 (N16381, N16372, N5535, N8665, N4214);
nor NOR4 (N16382, N16370, N3821, N2365, N540);
and AND2 (N16383, N16378, N4286);
buf BUF1 (N16384, N16371);
and AND4 (N16385, N16374, N6549, N7688, N1556);
not NOT1 (N16386, N16382);
xor XOR2 (N16387, N16380, N7397);
xor XOR2 (N16388, N16343, N13734);
nor NOR4 (N16389, N16352, N15818, N508, N7930);
nand NAND4 (N16390, N16386, N15544, N260, N11835);
and AND4 (N16391, N16381, N10035, N9891, N13570);
xor XOR2 (N16392, N16383, N4954);
buf BUF1 (N16393, N16375);
nand NAND3 (N16394, N16391, N9090, N5057);
xor XOR2 (N16395, N16387, N16302);
xor XOR2 (N16396, N16385, N2740);
not NOT1 (N16397, N16389);
or OR4 (N16398, N16390, N8929, N1416, N10767);
buf BUF1 (N16399, N16392);
buf BUF1 (N16400, N16396);
nand NAND4 (N16401, N16394, N12133, N12311, N2923);
nand NAND2 (N16402, N16401, N10117);
or OR2 (N16403, N16402, N11042);
nor NOR3 (N16404, N16403, N35, N10593);
not NOT1 (N16405, N16379);
and AND4 (N16406, N16398, N12297, N8114, N9750);
nand NAND3 (N16407, N16393, N3682, N15691);
nor NOR4 (N16408, N16406, N2870, N6210, N5622);
or OR3 (N16409, N16397, N14174, N4742);
xor XOR2 (N16410, N16400, N389);
not NOT1 (N16411, N16384);
nor NOR3 (N16412, N16399, N658, N3302);
and AND4 (N16413, N16404, N3832, N10478, N12332);
xor XOR2 (N16414, N16409, N8653);
not NOT1 (N16415, N16395);
or OR4 (N16416, N16412, N5819, N13456, N4517);
nand NAND2 (N16417, N16416, N8915);
nand NAND2 (N16418, N16413, N7436);
nor NOR2 (N16419, N16414, N3547);
nand NAND2 (N16420, N16411, N8014);
not NOT1 (N16421, N16420);
nand NAND2 (N16422, N16415, N5600);
xor XOR2 (N16423, N16418, N13001);
or OR2 (N16424, N16405, N8468);
or OR3 (N16425, N16407, N10857, N5379);
and AND4 (N16426, N16425, N8425, N14529, N13209);
nor NOR2 (N16427, N16426, N3730);
xor XOR2 (N16428, N16419, N5103);
not NOT1 (N16429, N16423);
and AND3 (N16430, N16427, N16270, N14050);
xor XOR2 (N16431, N16430, N8214);
buf BUF1 (N16432, N16424);
nor NOR4 (N16433, N16410, N10687, N13132, N7038);
nand NAND4 (N16434, N16431, N4187, N3278, N12967);
xor XOR2 (N16435, N16433, N6491);
buf BUF1 (N16436, N16408);
and AND3 (N16437, N16417, N6988, N2276);
buf BUF1 (N16438, N16437);
xor XOR2 (N16439, N16429, N3163);
and AND2 (N16440, N16428, N9100);
not NOT1 (N16441, N16438);
nor NOR4 (N16442, N16422, N5635, N12214, N10701);
and AND2 (N16443, N16441, N15805);
or OR2 (N16444, N16443, N5742);
nand NAND4 (N16445, N16439, N14672, N5923, N13873);
nor NOR4 (N16446, N16440, N10370, N2144, N14934);
or OR3 (N16447, N16442, N1896, N2290);
buf BUF1 (N16448, N16444);
and AND3 (N16449, N16388, N13151, N9489);
nor NOR2 (N16450, N16435, N11787);
xor XOR2 (N16451, N16445, N12082);
nand NAND4 (N16452, N16432, N13343, N8324, N2335);
buf BUF1 (N16453, N16446);
or OR2 (N16454, N16448, N6415);
nand NAND4 (N16455, N16434, N16122, N6329, N10022);
buf BUF1 (N16456, N16454);
buf BUF1 (N16457, N16453);
nor NOR2 (N16458, N16456, N14587);
and AND2 (N16459, N16449, N14906);
or OR4 (N16460, N16459, N6492, N8704, N1159);
buf BUF1 (N16461, N16450);
or OR4 (N16462, N16447, N10265, N13602, N6642);
buf BUF1 (N16463, N16458);
or OR3 (N16464, N16455, N662, N15491);
nor NOR3 (N16465, N16464, N6506, N7843);
xor XOR2 (N16466, N16421, N9831);
nand NAND3 (N16467, N16463, N263, N386);
buf BUF1 (N16468, N16467);
xor XOR2 (N16469, N16436, N3254);
nor NOR3 (N16470, N16460, N11810, N13797);
nand NAND4 (N16471, N16461, N93, N6185, N11578);
xor XOR2 (N16472, N16466, N5060);
or OR2 (N16473, N16468, N7571);
xor XOR2 (N16474, N16452, N7919);
xor XOR2 (N16475, N16474, N9460);
buf BUF1 (N16476, N16457);
not NOT1 (N16477, N16471);
buf BUF1 (N16478, N16465);
not NOT1 (N16479, N16470);
xor XOR2 (N16480, N16475, N15234);
not NOT1 (N16481, N16477);
xor XOR2 (N16482, N16479, N11262);
nor NOR2 (N16483, N16482, N1115);
xor XOR2 (N16484, N16451, N6484);
xor XOR2 (N16485, N16478, N12543);
nand NAND3 (N16486, N16485, N7350, N6095);
and AND4 (N16487, N16484, N4673, N3742, N4165);
and AND2 (N16488, N16472, N2644);
nand NAND4 (N16489, N16469, N16362, N7992, N3263);
not NOT1 (N16490, N16486);
and AND2 (N16491, N16462, N11705);
or OR2 (N16492, N16480, N1672);
and AND2 (N16493, N16490, N11772);
not NOT1 (N16494, N16473);
and AND4 (N16495, N16492, N6878, N3557, N15716);
and AND2 (N16496, N16489, N4767);
and AND2 (N16497, N16476, N414);
nand NAND2 (N16498, N16491, N12401);
and AND2 (N16499, N16495, N14219);
nor NOR4 (N16500, N16493, N1864, N14940, N10301);
or OR3 (N16501, N16499, N2429, N4917);
not NOT1 (N16502, N16498);
nor NOR2 (N16503, N16494, N12144);
or OR2 (N16504, N16481, N4392);
not NOT1 (N16505, N16488);
xor XOR2 (N16506, N16496, N5184);
nand NAND4 (N16507, N16483, N10603, N197, N7151);
or OR4 (N16508, N16487, N12345, N16450, N15873);
nor NOR3 (N16509, N16502, N13194, N10884);
or OR4 (N16510, N16504, N12567, N14216, N3938);
or OR4 (N16511, N16500, N5071, N13734, N6070);
nor NOR4 (N16512, N16501, N837, N1637, N5413);
buf BUF1 (N16513, N16512);
xor XOR2 (N16514, N16508, N550);
nand NAND4 (N16515, N16507, N8916, N213, N10926);
or OR2 (N16516, N16511, N3168);
xor XOR2 (N16517, N16503, N7637);
buf BUF1 (N16518, N16505);
xor XOR2 (N16519, N16497, N6276);
buf BUF1 (N16520, N16515);
not NOT1 (N16521, N16516);
buf BUF1 (N16522, N16518);
or OR3 (N16523, N16522, N4395, N13721);
and AND3 (N16524, N16510, N6875, N15840);
xor XOR2 (N16525, N16519, N13422);
nor NOR2 (N16526, N16523, N90);
not NOT1 (N16527, N16509);
and AND3 (N16528, N16514, N1454, N10037);
buf BUF1 (N16529, N16521);
nand NAND4 (N16530, N16520, N5696, N5520, N12598);
not NOT1 (N16531, N16517);
and AND3 (N16532, N16531, N15068, N5111);
buf BUF1 (N16533, N16530);
nand NAND2 (N16534, N16532, N3637);
and AND4 (N16535, N16524, N10559, N1686, N6307);
not NOT1 (N16536, N16527);
or OR2 (N16537, N16534, N5399);
not NOT1 (N16538, N16535);
buf BUF1 (N16539, N16529);
xor XOR2 (N16540, N16506, N5764);
nand NAND4 (N16541, N16540, N4707, N10342, N5405);
not NOT1 (N16542, N16528);
not NOT1 (N16543, N16539);
and AND4 (N16544, N16513, N5994, N1272, N141);
nor NOR3 (N16545, N16542, N14597, N10896);
nand NAND2 (N16546, N16544, N3980);
and AND4 (N16547, N16543, N11125, N16048, N951);
buf BUF1 (N16548, N16537);
xor XOR2 (N16549, N16536, N2238);
xor XOR2 (N16550, N16545, N13421);
or OR4 (N16551, N16538, N14179, N10914, N11141);
and AND4 (N16552, N16550, N2990, N13724, N1882);
not NOT1 (N16553, N16541);
xor XOR2 (N16554, N16526, N12528);
buf BUF1 (N16555, N16551);
buf BUF1 (N16556, N16548);
and AND4 (N16557, N16546, N515, N16176, N15529);
and AND3 (N16558, N16549, N7954, N12961);
nor NOR4 (N16559, N16553, N4429, N15254, N615);
nor NOR4 (N16560, N16555, N7951, N696, N3892);
xor XOR2 (N16561, N16560, N11612);
not NOT1 (N16562, N16552);
buf BUF1 (N16563, N16557);
not NOT1 (N16564, N16563);
xor XOR2 (N16565, N16547, N12289);
nand NAND2 (N16566, N16554, N7177);
not NOT1 (N16567, N16561);
buf BUF1 (N16568, N16564);
buf BUF1 (N16569, N16533);
and AND4 (N16570, N16569, N9552, N15095, N15773);
or OR2 (N16571, N16525, N652);
nor NOR3 (N16572, N16571, N12468, N932);
or OR3 (N16573, N16566, N7444, N15999);
nand NAND3 (N16574, N16573, N1404, N11070);
nand NAND2 (N16575, N16558, N8996);
xor XOR2 (N16576, N16570, N13035);
nand NAND2 (N16577, N16565, N14397);
not NOT1 (N16578, N16562);
not NOT1 (N16579, N16574);
nor NOR3 (N16580, N16556, N14811, N8465);
or OR4 (N16581, N16575, N1791, N6457, N3178);
nor NOR3 (N16582, N16559, N14054, N16010);
nand NAND4 (N16583, N16578, N2141, N15202, N6462);
and AND4 (N16584, N16576, N7510, N7382, N11782);
xor XOR2 (N16585, N16580, N10212);
xor XOR2 (N16586, N16579, N15901);
buf BUF1 (N16587, N16585);
xor XOR2 (N16588, N16572, N7333);
and AND4 (N16589, N16584, N6563, N15658, N13517);
buf BUF1 (N16590, N16581);
nand NAND3 (N16591, N16587, N15964, N10480);
nor NOR3 (N16592, N16590, N11869, N12984);
nor NOR4 (N16593, N16577, N2318, N2233, N7083);
nor NOR4 (N16594, N16567, N6294, N1248, N6464);
xor XOR2 (N16595, N16586, N14320);
nor NOR3 (N16596, N16588, N11094, N6705);
or OR3 (N16597, N16591, N7283, N11573);
buf BUF1 (N16598, N16594);
nor NOR3 (N16599, N16595, N10070, N13810);
or OR3 (N16600, N16589, N14067, N5587);
xor XOR2 (N16601, N16597, N7748);
nand NAND4 (N16602, N16593, N2010, N12187, N15251);
or OR3 (N16603, N16600, N7642, N3399);
not NOT1 (N16604, N16598);
xor XOR2 (N16605, N16582, N11743);
xor XOR2 (N16606, N16603, N14743);
not NOT1 (N16607, N16596);
or OR3 (N16608, N16583, N5453, N9608);
nor NOR3 (N16609, N16604, N7563, N13301);
or OR4 (N16610, N16606, N9530, N718, N2610);
nand NAND2 (N16611, N16605, N13108);
not NOT1 (N16612, N16568);
nand NAND2 (N16613, N16592, N9061);
or OR2 (N16614, N16601, N15630);
xor XOR2 (N16615, N16609, N16392);
nor NOR2 (N16616, N16602, N9478);
nor NOR3 (N16617, N16610, N4606, N15677);
xor XOR2 (N16618, N16608, N9845);
nor NOR3 (N16619, N16615, N12987, N6249);
buf BUF1 (N16620, N16616);
and AND3 (N16621, N16617, N1660, N12183);
and AND3 (N16622, N16607, N14216, N1780);
nand NAND4 (N16623, N16622, N11059, N9015, N3886);
nand NAND2 (N16624, N16618, N13342);
nand NAND3 (N16625, N16599, N8951, N10207);
and AND3 (N16626, N16624, N10135, N2212);
buf BUF1 (N16627, N16621);
and AND4 (N16628, N16623, N14225, N12833, N4222);
not NOT1 (N16629, N16619);
and AND3 (N16630, N16613, N13587, N13721);
not NOT1 (N16631, N16611);
and AND2 (N16632, N16612, N6512);
nand NAND3 (N16633, N16632, N2627, N1187);
and AND4 (N16634, N16631, N14102, N14753, N5926);
not NOT1 (N16635, N16626);
or OR4 (N16636, N16633, N3015, N14046, N7919);
xor XOR2 (N16637, N16635, N15032);
or OR4 (N16638, N16620, N8889, N14725, N2222);
buf BUF1 (N16639, N16637);
nor NOR4 (N16640, N16628, N911, N15410, N7736);
nor NOR2 (N16641, N16614, N2436);
nand NAND3 (N16642, N16634, N5319, N5021);
and AND4 (N16643, N16640, N3393, N13127, N8776);
nand NAND3 (N16644, N16643, N6284, N43);
nor NOR4 (N16645, N16625, N16543, N4338, N3717);
not NOT1 (N16646, N16642);
buf BUF1 (N16647, N16641);
buf BUF1 (N16648, N16647);
xor XOR2 (N16649, N16644, N15598);
not NOT1 (N16650, N16630);
or OR4 (N16651, N16648, N12052, N8491, N4096);
and AND3 (N16652, N16646, N3439, N9895);
not NOT1 (N16653, N16639);
not NOT1 (N16654, N16636);
or OR3 (N16655, N16651, N11977, N2375);
not NOT1 (N16656, N16627);
and AND2 (N16657, N16629, N10717);
buf BUF1 (N16658, N16657);
or OR3 (N16659, N16652, N1754, N8419);
not NOT1 (N16660, N16645);
or OR4 (N16661, N16660, N11426, N9545, N10618);
buf BUF1 (N16662, N16655);
and AND3 (N16663, N16662, N11594, N289);
or OR2 (N16664, N16663, N14462);
nor NOR2 (N16665, N16654, N14940);
not NOT1 (N16666, N16649);
and AND2 (N16667, N16665, N2923);
nor NOR3 (N16668, N16656, N5285, N7305);
nand NAND4 (N16669, N16650, N3426, N8482, N8650);
not NOT1 (N16670, N16666);
not NOT1 (N16671, N16659);
or OR3 (N16672, N16638, N9122, N5449);
nor NOR4 (N16673, N16653, N15422, N6554, N9277);
xor XOR2 (N16674, N16667, N1032);
buf BUF1 (N16675, N16673);
nand NAND3 (N16676, N16675, N11497, N2249);
not NOT1 (N16677, N16676);
xor XOR2 (N16678, N16677, N11408);
or OR4 (N16679, N16669, N3496, N10278, N5567);
or OR3 (N16680, N16678, N7138, N6406);
or OR4 (N16681, N16668, N2686, N4775, N3612);
nand NAND4 (N16682, N16671, N15084, N6656, N14098);
and AND3 (N16683, N16681, N11445, N9379);
or OR2 (N16684, N16680, N1913);
and AND3 (N16685, N16684, N14277, N15681);
nor NOR4 (N16686, N16682, N7412, N10976, N16073);
or OR2 (N16687, N16674, N7432);
buf BUF1 (N16688, N16685);
or OR2 (N16689, N16679, N8831);
or OR4 (N16690, N16664, N15947, N1018, N10006);
not NOT1 (N16691, N16670);
and AND3 (N16692, N16661, N10043, N5140);
nand NAND4 (N16693, N16687, N9071, N2355, N4786);
not NOT1 (N16694, N16689);
or OR4 (N16695, N16692, N10606, N2469, N16613);
not NOT1 (N16696, N16695);
not NOT1 (N16697, N16683);
nand NAND4 (N16698, N16697, N15397, N16454, N10550);
and AND4 (N16699, N16672, N7618, N7225, N5395);
and AND3 (N16700, N16694, N8977, N13996);
and AND3 (N16701, N16693, N15340, N8504);
and AND3 (N16702, N16688, N10239, N14824);
or OR4 (N16703, N16698, N11902, N15814, N13505);
not NOT1 (N16704, N16701);
nor NOR3 (N16705, N16696, N215, N4115);
not NOT1 (N16706, N16705);
not NOT1 (N16707, N16686);
xor XOR2 (N16708, N16700, N4700);
or OR2 (N16709, N16706, N9164);
and AND4 (N16710, N16691, N11159, N6169, N7645);
buf BUF1 (N16711, N16702);
and AND2 (N16712, N16690, N13125);
buf BUF1 (N16713, N16704);
or OR2 (N16714, N16708, N7721);
nor NOR4 (N16715, N16713, N13272, N4706, N15957);
xor XOR2 (N16716, N16707, N10754);
nand NAND4 (N16717, N16699, N1688, N6085, N6773);
and AND3 (N16718, N16711, N16279, N5856);
not NOT1 (N16719, N16703);
xor XOR2 (N16720, N16719, N8829);
or OR4 (N16721, N16714, N12915, N6282, N2441);
buf BUF1 (N16722, N16715);
or OR4 (N16723, N16718, N2254, N13865, N5532);
xor XOR2 (N16724, N16721, N453);
or OR2 (N16725, N16712, N8549);
or OR3 (N16726, N16710, N5217, N3334);
and AND2 (N16727, N16726, N13610);
xor XOR2 (N16728, N16727, N14255);
nand NAND4 (N16729, N16724, N1775, N7049, N10395);
and AND2 (N16730, N16717, N1717);
nand NAND4 (N16731, N16723, N8870, N8314, N4428);
nand NAND4 (N16732, N16716, N955, N11106, N10787);
xor XOR2 (N16733, N16720, N5917);
or OR4 (N16734, N16728, N11626, N14528, N1483);
or OR2 (N16735, N16658, N2126);
nand NAND2 (N16736, N16733, N9921);
xor XOR2 (N16737, N16732, N13989);
or OR3 (N16738, N16731, N6668, N15135);
buf BUF1 (N16739, N16736);
or OR4 (N16740, N16739, N6390, N12561, N3187);
or OR4 (N16741, N16737, N420, N14809, N8593);
or OR4 (N16742, N16741, N9874, N14133, N12623);
xor XOR2 (N16743, N16709, N10723);
not NOT1 (N16744, N16740);
xor XOR2 (N16745, N16744, N9133);
and AND4 (N16746, N16725, N6717, N16528, N6022);
or OR4 (N16747, N16722, N12782, N11855, N16665);
buf BUF1 (N16748, N16735);
xor XOR2 (N16749, N16748, N14525);
buf BUF1 (N16750, N16730);
nand NAND4 (N16751, N16746, N10385, N5404, N10531);
not NOT1 (N16752, N16729);
xor XOR2 (N16753, N16743, N12008);
xor XOR2 (N16754, N16753, N11730);
not NOT1 (N16755, N16752);
nand NAND3 (N16756, N16750, N4418, N11027);
nand NAND3 (N16757, N16747, N6876, N9450);
buf BUF1 (N16758, N16734);
and AND3 (N16759, N16757, N4434, N6940);
buf BUF1 (N16760, N16754);
nand NAND4 (N16761, N16756, N7969, N8577, N8756);
and AND4 (N16762, N16759, N16291, N16527, N8);
nand NAND3 (N16763, N16762, N8762, N6056);
and AND4 (N16764, N16755, N2691, N417, N9374);
not NOT1 (N16765, N16760);
nand NAND2 (N16766, N16745, N9184);
not NOT1 (N16767, N16761);
or OR3 (N16768, N16758, N7424, N15185);
or OR3 (N16769, N16749, N655, N4015);
or OR4 (N16770, N16764, N2034, N6906, N1296);
not NOT1 (N16771, N16769);
and AND4 (N16772, N16738, N10677, N14661, N5679);
and AND4 (N16773, N16770, N1224, N355, N8932);
not NOT1 (N16774, N16768);
and AND4 (N16775, N16742, N8924, N4016, N1547);
not NOT1 (N16776, N16772);
not NOT1 (N16777, N16763);
and AND2 (N16778, N16766, N2951);
nor NOR3 (N16779, N16767, N7056, N4590);
and AND4 (N16780, N16776, N5771, N14221, N1507);
and AND4 (N16781, N16775, N14737, N8329, N5580);
nor NOR2 (N16782, N16751, N10282);
or OR2 (N16783, N16781, N14931);
buf BUF1 (N16784, N16771);
nor NOR4 (N16785, N16782, N7062, N12365, N9369);
nand NAND4 (N16786, N16765, N14637, N13593, N10179);
not NOT1 (N16787, N16786);
buf BUF1 (N16788, N16773);
not NOT1 (N16789, N16785);
nand NAND4 (N16790, N16777, N14083, N5046, N10936);
buf BUF1 (N16791, N16787);
not NOT1 (N16792, N16778);
or OR3 (N16793, N16791, N13659, N14440);
nor NOR4 (N16794, N16789, N13491, N10548, N8626);
or OR4 (N16795, N16790, N2180, N10230, N6076);
not NOT1 (N16796, N16792);
or OR4 (N16797, N16795, N2982, N1818, N7526);
nor NOR2 (N16798, N16779, N10462);
nand NAND2 (N16799, N16774, N13808);
buf BUF1 (N16800, N16798);
buf BUF1 (N16801, N16788);
buf BUF1 (N16802, N16797);
not NOT1 (N16803, N16783);
xor XOR2 (N16804, N16799, N578);
nor NOR4 (N16805, N16793, N3710, N8431, N16210);
not NOT1 (N16806, N16805);
buf BUF1 (N16807, N16804);
xor XOR2 (N16808, N16796, N1161);
not NOT1 (N16809, N16808);
nand NAND2 (N16810, N16800, N12461);
nor NOR2 (N16811, N16784, N13354);
nand NAND2 (N16812, N16806, N8213);
xor XOR2 (N16813, N16809, N7367);
and AND4 (N16814, N16812, N7677, N15872, N9684);
or OR4 (N16815, N16813, N11485, N15419, N590);
nand NAND4 (N16816, N16803, N10981, N7573, N5837);
and AND2 (N16817, N16807, N14202);
xor XOR2 (N16818, N16810, N11516);
buf BUF1 (N16819, N16817);
nor NOR4 (N16820, N16802, N15629, N801, N6476);
and AND3 (N16821, N16819, N2061, N2890);
nand NAND3 (N16822, N16815, N5694, N3726);
nor NOR3 (N16823, N16780, N9459, N10011);
not NOT1 (N16824, N16794);
or OR3 (N16825, N16823, N8742, N5899);
and AND4 (N16826, N16801, N16653, N5568, N11439);
and AND2 (N16827, N16826, N6489);
nor NOR3 (N16828, N16825, N8429, N7621);
nand NAND4 (N16829, N16820, N13399, N4022, N9293);
not NOT1 (N16830, N16828);
nor NOR4 (N16831, N16811, N6462, N3345, N7303);
or OR4 (N16832, N16816, N13049, N15254, N11418);
and AND2 (N16833, N16829, N12579);
xor XOR2 (N16834, N16821, N1312);
and AND3 (N16835, N16824, N844, N13875);
not NOT1 (N16836, N16833);
xor XOR2 (N16837, N16830, N12308);
buf BUF1 (N16838, N16832);
buf BUF1 (N16839, N16831);
and AND3 (N16840, N16839, N4549, N6277);
or OR4 (N16841, N16814, N11577, N12269, N14217);
not NOT1 (N16842, N16836);
nor NOR3 (N16843, N16835, N3051, N15926);
xor XOR2 (N16844, N16843, N4122);
nand NAND3 (N16845, N16834, N2556, N9165);
or OR3 (N16846, N16838, N11180, N7578);
and AND4 (N16847, N16844, N4202, N266, N15608);
buf BUF1 (N16848, N16822);
buf BUF1 (N16849, N16840);
xor XOR2 (N16850, N16827, N917);
buf BUF1 (N16851, N16848);
nand NAND4 (N16852, N16851, N7468, N1437, N13921);
not NOT1 (N16853, N16818);
not NOT1 (N16854, N16841);
not NOT1 (N16855, N16846);
xor XOR2 (N16856, N16850, N2697);
or OR2 (N16857, N16856, N14109);
or OR4 (N16858, N16847, N212, N2646, N10636);
buf BUF1 (N16859, N16849);
nand NAND4 (N16860, N16852, N9891, N14181, N5573);
or OR3 (N16861, N16858, N13406, N6194);
xor XOR2 (N16862, N16855, N5963);
not NOT1 (N16863, N16859);
nand NAND2 (N16864, N16863, N4373);
buf BUF1 (N16865, N16864);
buf BUF1 (N16866, N16865);
xor XOR2 (N16867, N16842, N6285);
and AND4 (N16868, N16866, N13217, N1203, N8616);
or OR2 (N16869, N16860, N4752);
not NOT1 (N16870, N16845);
nor NOR2 (N16871, N16868, N831);
xor XOR2 (N16872, N16837, N11350);
xor XOR2 (N16873, N16867, N3119);
xor XOR2 (N16874, N16861, N6769);
xor XOR2 (N16875, N16869, N9512);
xor XOR2 (N16876, N16873, N6790);
buf BUF1 (N16877, N16876);
buf BUF1 (N16878, N16874);
xor XOR2 (N16879, N16877, N9998);
not NOT1 (N16880, N16862);
buf BUF1 (N16881, N16880);
or OR3 (N16882, N16853, N7026, N9361);
nand NAND3 (N16883, N16875, N6379, N13068);
nand NAND4 (N16884, N16871, N2112, N9319, N7323);
nor NOR2 (N16885, N16879, N11343);
nor NOR2 (N16886, N16881, N3376);
and AND2 (N16887, N16857, N13865);
buf BUF1 (N16888, N16886);
xor XOR2 (N16889, N16870, N4193);
buf BUF1 (N16890, N16882);
and AND2 (N16891, N16890, N8654);
or OR2 (N16892, N16888, N15191);
or OR3 (N16893, N16887, N6235, N277);
or OR3 (N16894, N16854, N15327, N5399);
nor NOR2 (N16895, N16892, N4711);
nand NAND2 (N16896, N16891, N4086);
not NOT1 (N16897, N16885);
nor NOR2 (N16898, N16884, N6338);
not NOT1 (N16899, N16895);
or OR2 (N16900, N16899, N16474);
xor XOR2 (N16901, N16872, N15084);
and AND3 (N16902, N16878, N10968, N6965);
and AND3 (N16903, N16900, N2488, N16227);
xor XOR2 (N16904, N16883, N7087);
nor NOR4 (N16905, N16889, N12092, N14643, N11349);
or OR4 (N16906, N16894, N16558, N8514, N15378);
or OR3 (N16907, N16898, N7771, N11138);
and AND4 (N16908, N16907, N13133, N14676, N15087);
buf BUF1 (N16909, N16904);
nand NAND3 (N16910, N16905, N16629, N8822);
buf BUF1 (N16911, N16906);
and AND3 (N16912, N16903, N15321, N8294);
nor NOR2 (N16913, N16901, N4876);
xor XOR2 (N16914, N16910, N9347);
not NOT1 (N16915, N16909);
nand NAND4 (N16916, N16896, N2, N1670, N11234);
nand NAND3 (N16917, N16897, N6128, N5517);
not NOT1 (N16918, N16911);
xor XOR2 (N16919, N16916, N4853);
and AND2 (N16920, N16902, N4378);
and AND2 (N16921, N16912, N11550);
xor XOR2 (N16922, N16913, N8097);
nand NAND2 (N16923, N16893, N9072);
nand NAND3 (N16924, N16919, N15402, N11403);
or OR2 (N16925, N16918, N7238);
not NOT1 (N16926, N16924);
nor NOR3 (N16927, N16917, N12600, N820);
buf BUF1 (N16928, N16920);
or OR4 (N16929, N16926, N15859, N7309, N8422);
not NOT1 (N16930, N16921);
and AND3 (N16931, N16929, N6523, N8713);
buf BUF1 (N16932, N16928);
xor XOR2 (N16933, N16927, N6189);
xor XOR2 (N16934, N16922, N5473);
or OR3 (N16935, N16933, N3928, N6160);
not NOT1 (N16936, N16931);
not NOT1 (N16937, N16915);
nand NAND3 (N16938, N16935, N3379, N2501);
not NOT1 (N16939, N16938);
nand NAND4 (N16940, N16937, N1596, N13607, N2962);
buf BUF1 (N16941, N16934);
xor XOR2 (N16942, N16939, N7994);
not NOT1 (N16943, N16942);
nand NAND3 (N16944, N16930, N9094, N9868);
buf BUF1 (N16945, N16925);
nor NOR2 (N16946, N16941, N16024);
not NOT1 (N16947, N16932);
nor NOR2 (N16948, N16923, N10038);
and AND2 (N16949, N16947, N2794);
buf BUF1 (N16950, N16936);
or OR3 (N16951, N16948, N13330, N1334);
xor XOR2 (N16952, N16949, N4794);
nor NOR4 (N16953, N16943, N9883, N10873, N13896);
xor XOR2 (N16954, N16952, N13642);
not NOT1 (N16955, N16953);
xor XOR2 (N16956, N16954, N3254);
not NOT1 (N16957, N16955);
xor XOR2 (N16958, N16914, N1546);
nand NAND3 (N16959, N16908, N7149, N9957);
xor XOR2 (N16960, N16940, N4463);
xor XOR2 (N16961, N16944, N12389);
nand NAND3 (N16962, N16958, N14453, N2016);
buf BUF1 (N16963, N16960);
and AND4 (N16964, N16946, N15039, N13753, N963);
buf BUF1 (N16965, N16956);
nand NAND3 (N16966, N16962, N15226, N13632);
nor NOR3 (N16967, N16961, N9946, N14719);
not NOT1 (N16968, N16950);
not NOT1 (N16969, N16964);
and AND2 (N16970, N16945, N7098);
buf BUF1 (N16971, N16970);
nand NAND2 (N16972, N16966, N6686);
nor NOR3 (N16973, N16968, N7852, N1655);
buf BUF1 (N16974, N16959);
buf BUF1 (N16975, N16967);
not NOT1 (N16976, N16951);
nor NOR3 (N16977, N16969, N3494, N1010);
not NOT1 (N16978, N16975);
and AND3 (N16979, N16977, N15398, N279);
and AND4 (N16980, N16974, N13610, N12329, N3954);
xor XOR2 (N16981, N16976, N12084);
not NOT1 (N16982, N16979);
and AND2 (N16983, N16972, N1164);
and AND4 (N16984, N16965, N7082, N3624, N16661);
buf BUF1 (N16985, N16984);
buf BUF1 (N16986, N16982);
not NOT1 (N16987, N16978);
nand NAND3 (N16988, N16973, N6690, N10246);
and AND2 (N16989, N16987, N2721);
buf BUF1 (N16990, N16963);
and AND2 (N16991, N16971, N14670);
nand NAND3 (N16992, N16990, N13119, N3812);
buf BUF1 (N16993, N16981);
nor NOR3 (N16994, N16980, N13193, N3557);
nor NOR2 (N16995, N16985, N12417);
nor NOR3 (N16996, N16991, N1602, N7867);
buf BUF1 (N16997, N16992);
xor XOR2 (N16998, N16997, N9357);
nand NAND2 (N16999, N16986, N13489);
nor NOR3 (N17000, N16983, N4871, N956);
or OR2 (N17001, N16989, N9098);
and AND3 (N17002, N17001, N4198, N5350);
or OR4 (N17003, N16988, N13193, N11190, N4592);
xor XOR2 (N17004, N16996, N7908);
or OR4 (N17005, N16999, N8539, N8817, N13384);
buf BUF1 (N17006, N17002);
or OR4 (N17007, N16993, N4459, N5285, N6779);
nor NOR4 (N17008, N16994, N10903, N13751, N13482);
not NOT1 (N17009, N17004);
nor NOR2 (N17010, N16995, N1913);
nor NOR3 (N17011, N17010, N15111, N2877);
buf BUF1 (N17012, N16957);
xor XOR2 (N17013, N17000, N15961);
buf BUF1 (N17014, N17011);
not NOT1 (N17015, N16998);
xor XOR2 (N17016, N17005, N908);
and AND3 (N17017, N17007, N16591, N14464);
nand NAND3 (N17018, N17014, N5178, N13150);
or OR3 (N17019, N17006, N4215, N624);
xor XOR2 (N17020, N17012, N15969);
and AND2 (N17021, N17016, N12794);
not NOT1 (N17022, N17018);
nand NAND2 (N17023, N17008, N10777);
nor NOR2 (N17024, N17019, N2651);
xor XOR2 (N17025, N17021, N6031);
nand NAND3 (N17026, N17003, N9528, N4311);
xor XOR2 (N17027, N17025, N8395);
nand NAND3 (N17028, N17015, N15620, N12472);
buf BUF1 (N17029, N17028);
buf BUF1 (N17030, N17023);
nor NOR4 (N17031, N17017, N10284, N3118, N9903);
xor XOR2 (N17032, N17031, N16867);
not NOT1 (N17033, N17013);
xor XOR2 (N17034, N17026, N7307);
not NOT1 (N17035, N17032);
xor XOR2 (N17036, N17030, N14039);
nor NOR4 (N17037, N17027, N8099, N12333, N5413);
buf BUF1 (N17038, N17034);
not NOT1 (N17039, N17038);
and AND4 (N17040, N17009, N16769, N14130, N4502);
buf BUF1 (N17041, N17035);
nand NAND4 (N17042, N17033, N3833, N11332, N7730);
and AND3 (N17043, N17029, N12793, N6302);
nand NAND3 (N17044, N17036, N16948, N9957);
nand NAND4 (N17045, N17044, N9261, N9638, N14780);
or OR3 (N17046, N17045, N5087, N7561);
not NOT1 (N17047, N17037);
xor XOR2 (N17048, N17047, N3060);
and AND3 (N17049, N17022, N1817, N5744);
xor XOR2 (N17050, N17043, N3563);
buf BUF1 (N17051, N17040);
nor NOR2 (N17052, N17024, N14082);
and AND3 (N17053, N17042, N11203, N5810);
or OR3 (N17054, N17039, N11786, N16080);
or OR3 (N17055, N17054, N592, N11132);
xor XOR2 (N17056, N17052, N4606);
nand NAND3 (N17057, N17048, N13541, N2362);
xor XOR2 (N17058, N17056, N4379);
xor XOR2 (N17059, N17046, N7711);
and AND4 (N17060, N17058, N8202, N1647, N2470);
nor NOR4 (N17061, N17050, N5515, N999, N16694);
nand NAND2 (N17062, N17061, N15651);
xor XOR2 (N17063, N17055, N16080);
buf BUF1 (N17064, N17059);
buf BUF1 (N17065, N17049);
and AND4 (N17066, N17065, N12146, N1685, N2367);
not NOT1 (N17067, N17051);
or OR2 (N17068, N17020, N421);
and AND4 (N17069, N17064, N14468, N1723, N15756);
not NOT1 (N17070, N17062);
nor NOR4 (N17071, N17063, N15553, N8281, N7842);
and AND3 (N17072, N17066, N13599, N14399);
or OR4 (N17073, N17041, N1888, N1826, N15964);
nand NAND3 (N17074, N17053, N9323, N3602);
buf BUF1 (N17075, N17067);
xor XOR2 (N17076, N17072, N9328);
and AND3 (N17077, N17068, N14686, N15901);
not NOT1 (N17078, N17077);
or OR2 (N17079, N17073, N3254);
or OR3 (N17080, N17078, N4688, N1375);
not NOT1 (N17081, N17060);
nor NOR3 (N17082, N17076, N2539, N9684);
nand NAND2 (N17083, N17057, N10824);
buf BUF1 (N17084, N17071);
nand NAND4 (N17085, N17084, N12056, N7256, N784);
nand NAND4 (N17086, N17069, N15981, N61, N13854);
or OR2 (N17087, N17080, N11267);
or OR4 (N17088, N17086, N11837, N7781, N14534);
not NOT1 (N17089, N17081);
not NOT1 (N17090, N17089);
nor NOR3 (N17091, N17088, N13520, N4239);
or OR3 (N17092, N17075, N10184, N767);
or OR3 (N17093, N17070, N4917, N7434);
nand NAND3 (N17094, N17082, N10960, N10681);
nand NAND4 (N17095, N17079, N14554, N9280, N7276);
and AND2 (N17096, N17095, N12999);
nand NAND4 (N17097, N17090, N15353, N31, N4079);
nor NOR4 (N17098, N17085, N10448, N13351, N4356);
buf BUF1 (N17099, N17091);
xor XOR2 (N17100, N17096, N16352);
nand NAND4 (N17101, N17083, N2069, N10963, N13942);
nand NAND2 (N17102, N17087, N11716);
xor XOR2 (N17103, N17099, N9698);
not NOT1 (N17104, N17097);
xor XOR2 (N17105, N17102, N15262);
nand NAND2 (N17106, N17101, N4621);
not NOT1 (N17107, N17074);
buf BUF1 (N17108, N17106);
or OR2 (N17109, N17107, N4148);
and AND4 (N17110, N17093, N6735, N2616, N15943);
nand NAND2 (N17111, N17109, N15833);
not NOT1 (N17112, N17104);
and AND4 (N17113, N17112, N15448, N1732, N4436);
xor XOR2 (N17114, N17113, N8765);
nand NAND4 (N17115, N17092, N4744, N2581, N15782);
and AND3 (N17116, N17111, N9052, N1903);
and AND4 (N17117, N17100, N14320, N6243, N11130);
xor XOR2 (N17118, N17117, N9332);
nand NAND2 (N17119, N17118, N5247);
or OR2 (N17120, N17114, N14075);
and AND4 (N17121, N17115, N7654, N15018, N14697);
or OR4 (N17122, N17098, N15176, N12349, N11574);
buf BUF1 (N17123, N17108);
and AND2 (N17124, N17103, N3193);
nor NOR2 (N17125, N17094, N2260);
and AND2 (N17126, N17110, N10408);
xor XOR2 (N17127, N17125, N3470);
buf BUF1 (N17128, N17122);
and AND2 (N17129, N17105, N5575);
and AND2 (N17130, N17126, N2523);
nand NAND3 (N17131, N17124, N9376, N3767);
or OR3 (N17132, N17131, N13023, N9953);
nand NAND4 (N17133, N17119, N11815, N13713, N49);
or OR4 (N17134, N17132, N5956, N7812, N98);
or OR4 (N17135, N17133, N11118, N4232, N4063);
xor XOR2 (N17136, N17134, N9632);
nor NOR2 (N17137, N17123, N11339);
nor NOR4 (N17138, N17137, N13620, N5262, N12670);
and AND2 (N17139, N17129, N13080);
nand NAND2 (N17140, N17128, N8889);
not NOT1 (N17141, N17135);
xor XOR2 (N17142, N17140, N11919);
nand NAND4 (N17143, N17116, N7175, N11214, N9523);
and AND4 (N17144, N17142, N10763, N6762, N13598);
and AND2 (N17145, N17130, N12746);
buf BUF1 (N17146, N17144);
nand NAND4 (N17147, N17121, N4609, N3559, N14508);
nand NAND2 (N17148, N17136, N13949);
not NOT1 (N17149, N17138);
or OR4 (N17150, N17149, N4486, N14622, N2588);
nand NAND3 (N17151, N17150, N7630, N14771);
not NOT1 (N17152, N17139);
not NOT1 (N17153, N17147);
nand NAND3 (N17154, N17153, N7834, N2356);
nor NOR3 (N17155, N17154, N16687, N11488);
nand NAND2 (N17156, N17141, N8544);
not NOT1 (N17157, N17156);
or OR2 (N17158, N17120, N1302);
and AND3 (N17159, N17143, N50, N6926);
and AND3 (N17160, N17151, N3162, N1703);
xor XOR2 (N17161, N17148, N4946);
or OR4 (N17162, N17152, N15899, N5216, N14545);
nor NOR3 (N17163, N17155, N1883, N15444);
or OR3 (N17164, N17159, N13543, N11731);
nand NAND3 (N17165, N17145, N2746, N8699);
buf BUF1 (N17166, N17127);
buf BUF1 (N17167, N17158);
buf BUF1 (N17168, N17167);
not NOT1 (N17169, N17164);
xor XOR2 (N17170, N17168, N7686);
and AND3 (N17171, N17146, N4464, N7540);
and AND4 (N17172, N17162, N6730, N2386, N552);
and AND4 (N17173, N17157, N7915, N2529, N9464);
buf BUF1 (N17174, N17161);
buf BUF1 (N17175, N17172);
not NOT1 (N17176, N17171);
not NOT1 (N17177, N17174);
nand NAND4 (N17178, N17170, N9526, N16042, N964);
or OR2 (N17179, N17175, N16653);
nor NOR3 (N17180, N17166, N12833, N1346);
nor NOR3 (N17181, N17177, N14818, N5114);
not NOT1 (N17182, N17169);
nor NOR4 (N17183, N17182, N2469, N13044, N14380);
and AND2 (N17184, N17160, N9395);
and AND3 (N17185, N17163, N11120, N3255);
xor XOR2 (N17186, N17176, N9907);
or OR2 (N17187, N17165, N489);
not NOT1 (N17188, N17180);
and AND2 (N17189, N17173, N1121);
and AND3 (N17190, N17187, N1108, N10597);
xor XOR2 (N17191, N17183, N122);
buf BUF1 (N17192, N17191);
xor XOR2 (N17193, N17179, N13515);
xor XOR2 (N17194, N17185, N13735);
buf BUF1 (N17195, N17189);
nand NAND3 (N17196, N17178, N13780, N15488);
not NOT1 (N17197, N17193);
nand NAND2 (N17198, N17194, N12699);
and AND2 (N17199, N17197, N2466);
nor NOR4 (N17200, N17190, N15598, N4599, N15625);
buf BUF1 (N17201, N17199);
or OR3 (N17202, N17192, N11832, N13896);
and AND3 (N17203, N17201, N13184, N9773);
nand NAND3 (N17204, N17181, N8153, N13863);
xor XOR2 (N17205, N17196, N3916);
and AND3 (N17206, N17195, N11965, N6487);
or OR3 (N17207, N17188, N5800, N13389);
buf BUF1 (N17208, N17198);
xor XOR2 (N17209, N17208, N7352);
or OR3 (N17210, N17186, N13689, N16896);
nor NOR3 (N17211, N17205, N16622, N10684);
nand NAND3 (N17212, N17184, N7440, N5689);
buf BUF1 (N17213, N17200);
xor XOR2 (N17214, N17207, N14138);
and AND4 (N17215, N17203, N16447, N8756, N11730);
buf BUF1 (N17216, N17215);
nor NOR2 (N17217, N17209, N4615);
nand NAND2 (N17218, N17214, N7137);
not NOT1 (N17219, N17202);
nand NAND3 (N17220, N17219, N15703, N9832);
and AND3 (N17221, N17206, N2077, N11982);
xor XOR2 (N17222, N17217, N14740);
buf BUF1 (N17223, N17212);
not NOT1 (N17224, N17220);
xor XOR2 (N17225, N17211, N2522);
and AND3 (N17226, N17216, N8435, N12164);
not NOT1 (N17227, N17223);
buf BUF1 (N17228, N17221);
buf BUF1 (N17229, N17218);
or OR3 (N17230, N17225, N8155, N5427);
nor NOR4 (N17231, N17230, N6792, N2166, N4156);
and AND2 (N17232, N17226, N12212);
nand NAND3 (N17233, N17210, N9538, N10392);
buf BUF1 (N17234, N17228);
not NOT1 (N17235, N17232);
buf BUF1 (N17236, N17231);
buf BUF1 (N17237, N17234);
nand NAND3 (N17238, N17204, N2191, N2961);
not NOT1 (N17239, N17233);
buf BUF1 (N17240, N17229);
xor XOR2 (N17241, N17235, N12522);
not NOT1 (N17242, N17240);
or OR4 (N17243, N17241, N14043, N3423, N5527);
or OR4 (N17244, N17242, N10883, N174, N14388);
or OR2 (N17245, N17236, N5887);
not NOT1 (N17246, N17238);
nor NOR2 (N17247, N17244, N5851);
or OR3 (N17248, N17243, N5156, N9390);
xor XOR2 (N17249, N17224, N3903);
buf BUF1 (N17250, N17239);
nor NOR3 (N17251, N17213, N13018, N11972);
not NOT1 (N17252, N17247);
buf BUF1 (N17253, N17246);
or OR2 (N17254, N17249, N3889);
xor XOR2 (N17255, N17227, N10873);
nor NOR3 (N17256, N17251, N4964, N17059);
buf BUF1 (N17257, N17254);
xor XOR2 (N17258, N17256, N485);
xor XOR2 (N17259, N17255, N2728);
or OR2 (N17260, N17252, N15737);
and AND2 (N17261, N17253, N12633);
xor XOR2 (N17262, N17237, N535);
buf BUF1 (N17263, N17257);
xor XOR2 (N17264, N17245, N3078);
nor NOR2 (N17265, N17248, N1009);
and AND3 (N17266, N17258, N16111, N16438);
not NOT1 (N17267, N17265);
not NOT1 (N17268, N17250);
xor XOR2 (N17269, N17263, N11990);
xor XOR2 (N17270, N17262, N14216);
or OR2 (N17271, N17269, N2210);
nand NAND4 (N17272, N17264, N8869, N4527, N2010);
nand NAND4 (N17273, N17271, N11268, N13964, N12443);
nand NAND3 (N17274, N17273, N12361, N8036);
and AND4 (N17275, N17222, N9900, N13588, N2942);
xor XOR2 (N17276, N17268, N6983);
not NOT1 (N17277, N17259);
buf BUF1 (N17278, N17260);
not NOT1 (N17279, N17270);
nor NOR4 (N17280, N17261, N4820, N16890, N2108);
nor NOR2 (N17281, N17278, N10775);
or OR3 (N17282, N17267, N5918, N15489);
or OR4 (N17283, N17280, N7956, N10411, N4334);
nor NOR2 (N17284, N17272, N14428);
and AND4 (N17285, N17282, N2824, N9281, N9522);
not NOT1 (N17286, N17275);
xor XOR2 (N17287, N17266, N16861);
and AND2 (N17288, N17284, N3558);
nand NAND3 (N17289, N17285, N3160, N6050);
or OR3 (N17290, N17289, N5173, N14806);
and AND4 (N17291, N17287, N3084, N17110, N744);
nand NAND4 (N17292, N17291, N2239, N2944, N25);
nand NAND2 (N17293, N17290, N7415);
or OR3 (N17294, N17281, N7035, N16874);
or OR4 (N17295, N17276, N10926, N3934, N11838);
not NOT1 (N17296, N17286);
buf BUF1 (N17297, N17288);
xor XOR2 (N17298, N17292, N293);
or OR2 (N17299, N17277, N9372);
and AND4 (N17300, N17294, N14818, N2430, N12315);
and AND2 (N17301, N17283, N6834);
or OR2 (N17302, N17295, N14795);
buf BUF1 (N17303, N17274);
nand NAND3 (N17304, N17298, N12107, N11258);
nor NOR4 (N17305, N17302, N4191, N13431, N10697);
not NOT1 (N17306, N17301);
buf BUF1 (N17307, N17297);
xor XOR2 (N17308, N17303, N14848);
or OR4 (N17309, N17305, N579, N90, N2585);
or OR3 (N17310, N17307, N1916, N6566);
and AND2 (N17311, N17296, N7819);
and AND4 (N17312, N17308, N12603, N5690, N16249);
xor XOR2 (N17313, N17299, N12255);
not NOT1 (N17314, N17311);
not NOT1 (N17315, N17293);
and AND2 (N17316, N17279, N10240);
nor NOR4 (N17317, N17306, N4962, N1927, N5283);
xor XOR2 (N17318, N17317, N7178);
buf BUF1 (N17319, N17309);
xor XOR2 (N17320, N17319, N13961);
buf BUF1 (N17321, N17313);
buf BUF1 (N17322, N17318);
nand NAND3 (N17323, N17322, N6366, N8640);
or OR4 (N17324, N17320, N235, N15952, N13863);
or OR4 (N17325, N17310, N4533, N13408, N6291);
nor NOR3 (N17326, N17323, N6028, N9586);
nor NOR4 (N17327, N17316, N12049, N4848, N3144);
and AND2 (N17328, N17324, N13501);
xor XOR2 (N17329, N17326, N4077);
nor NOR4 (N17330, N17304, N9253, N15961, N1048);
buf BUF1 (N17331, N17315);
nand NAND3 (N17332, N17329, N16966, N8614);
buf BUF1 (N17333, N17300);
nor NOR3 (N17334, N17332, N4047, N10787);
xor XOR2 (N17335, N17327, N14620);
not NOT1 (N17336, N17331);
nor NOR2 (N17337, N17333, N8840);
xor XOR2 (N17338, N17335, N17181);
or OR4 (N17339, N17334, N12062, N1989, N686);
nor NOR3 (N17340, N17325, N4373, N3203);
not NOT1 (N17341, N17312);
nor NOR4 (N17342, N17336, N493, N10773, N9854);
buf BUF1 (N17343, N17337);
nand NAND2 (N17344, N17342, N8592);
and AND2 (N17345, N17321, N955);
or OR2 (N17346, N17314, N8798);
or OR2 (N17347, N17346, N15262);
and AND2 (N17348, N17328, N4516);
or OR4 (N17349, N17340, N10203, N12436, N6553);
nand NAND3 (N17350, N17343, N11911, N12811);
and AND4 (N17351, N17330, N13588, N4752, N15947);
buf BUF1 (N17352, N17349);
buf BUF1 (N17353, N17345);
not NOT1 (N17354, N17347);
buf BUF1 (N17355, N17339);
nor NOR2 (N17356, N17348, N4642);
buf BUF1 (N17357, N17352);
buf BUF1 (N17358, N17341);
and AND3 (N17359, N17350, N13002, N12995);
nand NAND4 (N17360, N17338, N7866, N2773, N6248);
or OR2 (N17361, N17356, N40);
or OR2 (N17362, N17355, N3761);
or OR3 (N17363, N17351, N8826, N1806);
or OR2 (N17364, N17357, N12018);
xor XOR2 (N17365, N17353, N2627);
buf BUF1 (N17366, N17360);
xor XOR2 (N17367, N17362, N5137);
and AND2 (N17368, N17364, N6858);
or OR2 (N17369, N17363, N4965);
or OR3 (N17370, N17369, N4311, N3344);
not NOT1 (N17371, N17365);
xor XOR2 (N17372, N17367, N5092);
and AND2 (N17373, N17359, N17086);
nand NAND3 (N17374, N17371, N12537, N4517);
or OR4 (N17375, N17368, N8596, N3180, N5342);
xor XOR2 (N17376, N17370, N14541);
or OR3 (N17377, N17354, N16195, N12134);
nand NAND3 (N17378, N17361, N2655, N4345);
buf BUF1 (N17379, N17372);
buf BUF1 (N17380, N17373);
not NOT1 (N17381, N17376);
and AND3 (N17382, N17381, N7417, N14830);
and AND2 (N17383, N17358, N12885);
not NOT1 (N17384, N17383);
xor XOR2 (N17385, N17380, N2490);
or OR4 (N17386, N17375, N7043, N16916, N7617);
or OR3 (N17387, N17378, N10537, N6955);
buf BUF1 (N17388, N17386);
xor XOR2 (N17389, N17374, N14519);
or OR2 (N17390, N17388, N2265);
buf BUF1 (N17391, N17344);
and AND3 (N17392, N17385, N1262, N10851);
nor NOR3 (N17393, N17392, N67, N15331);
xor XOR2 (N17394, N17387, N1602);
buf BUF1 (N17395, N17389);
or OR2 (N17396, N17379, N8764);
nor NOR4 (N17397, N17393, N14274, N15500, N5555);
nand NAND3 (N17398, N17396, N9102, N16943);
buf BUF1 (N17399, N17377);
or OR4 (N17400, N17391, N549, N7636, N15678);
not NOT1 (N17401, N17398);
buf BUF1 (N17402, N17384);
xor XOR2 (N17403, N17395, N12909);
nor NOR2 (N17404, N17366, N9812);
nor NOR3 (N17405, N17399, N13721, N920);
not NOT1 (N17406, N17402);
buf BUF1 (N17407, N17394);
not NOT1 (N17408, N17382);
nor NOR4 (N17409, N17405, N2733, N7287, N14884);
nor NOR2 (N17410, N17407, N11872);
not NOT1 (N17411, N17397);
and AND4 (N17412, N17409, N13659, N15834, N5575);
not NOT1 (N17413, N17401);
buf BUF1 (N17414, N17411);
xor XOR2 (N17415, N17400, N4354);
xor XOR2 (N17416, N17403, N508);
nand NAND2 (N17417, N17408, N15563);
xor XOR2 (N17418, N17412, N12224);
not NOT1 (N17419, N17417);
nand NAND2 (N17420, N17410, N1159);
nand NAND2 (N17421, N17390, N1914);
or OR4 (N17422, N17414, N12654, N13168, N15046);
nand NAND4 (N17423, N17418, N1395, N6722, N15804);
buf BUF1 (N17424, N17416);
xor XOR2 (N17425, N17406, N12715);
nor NOR4 (N17426, N17413, N4430, N4193, N11145);
not NOT1 (N17427, N17426);
or OR2 (N17428, N17415, N9039);
or OR4 (N17429, N17425, N17082, N15284, N8274);
nand NAND3 (N17430, N17429, N12018, N13883);
nor NOR2 (N17431, N17422, N11805);
not NOT1 (N17432, N17423);
nor NOR4 (N17433, N17420, N3802, N8809, N13825);
nor NOR2 (N17434, N17433, N5166);
nor NOR4 (N17435, N17427, N840, N2704, N2620);
not NOT1 (N17436, N17430);
buf BUF1 (N17437, N17419);
or OR3 (N17438, N17431, N15237, N16671);
buf BUF1 (N17439, N17435);
xor XOR2 (N17440, N17432, N12018);
nor NOR3 (N17441, N17404, N8437, N6511);
or OR3 (N17442, N17421, N6534, N1954);
nand NAND4 (N17443, N17437, N9701, N3447, N17428);
buf BUF1 (N17444, N10217);
or OR4 (N17445, N17441, N13193, N9039, N5299);
not NOT1 (N17446, N17439);
xor XOR2 (N17447, N17442, N12165);
nand NAND4 (N17448, N17446, N7884, N4613, N10550);
xor XOR2 (N17449, N17436, N16381);
buf BUF1 (N17450, N17444);
not NOT1 (N17451, N17440);
or OR2 (N17452, N17438, N16688);
xor XOR2 (N17453, N17434, N13360);
and AND4 (N17454, N17448, N1378, N14496, N3896);
nor NOR2 (N17455, N17454, N6447);
and AND2 (N17456, N17449, N6643);
nor NOR4 (N17457, N17453, N9606, N1727, N12477);
not NOT1 (N17458, N17443);
nor NOR2 (N17459, N17451, N2970);
or OR2 (N17460, N17458, N15665);
not NOT1 (N17461, N17459);
not NOT1 (N17462, N17452);
buf BUF1 (N17463, N17424);
not NOT1 (N17464, N17462);
buf BUF1 (N17465, N17450);
nor NOR4 (N17466, N17465, N13551, N3308, N2050);
and AND3 (N17467, N17466, N12725, N11359);
and AND3 (N17468, N17457, N6389, N3195);
nand NAND4 (N17469, N17460, N5820, N7695, N1000);
xor XOR2 (N17470, N17455, N6417);
not NOT1 (N17471, N17467);
nand NAND3 (N17472, N17468, N2252, N15257);
xor XOR2 (N17473, N17470, N7386);
xor XOR2 (N17474, N17463, N7042);
and AND2 (N17475, N17469, N7814);
nand NAND3 (N17476, N17456, N2806, N11868);
nor NOR3 (N17477, N17445, N9080, N15381);
or OR4 (N17478, N17474, N2200, N14997, N12802);
and AND3 (N17479, N17472, N7865, N3014);
xor XOR2 (N17480, N17478, N14275);
buf BUF1 (N17481, N17447);
xor XOR2 (N17482, N17477, N2910);
and AND2 (N17483, N17464, N9102);
and AND3 (N17484, N17483, N4322, N14284);
and AND4 (N17485, N17475, N4983, N8629, N2522);
or OR4 (N17486, N17476, N2964, N6767, N3072);
not NOT1 (N17487, N17473);
xor XOR2 (N17488, N17471, N2898);
or OR2 (N17489, N17486, N168);
not NOT1 (N17490, N17485);
or OR2 (N17491, N17480, N15932);
nor NOR4 (N17492, N17461, N3979, N16270, N15473);
nand NAND4 (N17493, N17479, N726, N10920, N3332);
nor NOR4 (N17494, N17481, N5877, N6206, N7183);
nor NOR4 (N17495, N17482, N1199, N12605, N5808);
nor NOR2 (N17496, N17490, N7675);
buf BUF1 (N17497, N17495);
or OR4 (N17498, N17496, N3017, N15465, N7240);
and AND4 (N17499, N17492, N9918, N895, N4764);
and AND3 (N17500, N17487, N1739, N10125);
not NOT1 (N17501, N17488);
or OR3 (N17502, N17500, N14507, N12739);
nand NAND4 (N17503, N17494, N8494, N12770, N12890);
or OR2 (N17504, N17498, N12590);
nor NOR2 (N17505, N17491, N10021);
or OR3 (N17506, N17497, N6979, N10350);
xor XOR2 (N17507, N17506, N10347);
nor NOR3 (N17508, N17484, N12643, N12630);
buf BUF1 (N17509, N17493);
nor NOR3 (N17510, N17504, N14558, N3122);
or OR2 (N17511, N17508, N1890);
or OR3 (N17512, N17507, N14125, N6739);
or OR3 (N17513, N17502, N1422, N452);
nor NOR3 (N17514, N17509, N6154, N535);
and AND4 (N17515, N17503, N17467, N16926, N17210);
xor XOR2 (N17516, N17501, N5418);
nand NAND2 (N17517, N17499, N14580);
xor XOR2 (N17518, N17505, N14818);
or OR4 (N17519, N17516, N8999, N3839, N10021);
nand NAND3 (N17520, N17510, N6788, N6852);
nand NAND3 (N17521, N17519, N16836, N2843);
not NOT1 (N17522, N17515);
nor NOR3 (N17523, N17512, N11844, N8000);
nand NAND2 (N17524, N17521, N7097);
and AND4 (N17525, N17518, N13837, N2797, N2851);
buf BUF1 (N17526, N17514);
nor NOR2 (N17527, N17517, N7149);
not NOT1 (N17528, N17520);
buf BUF1 (N17529, N17525);
buf BUF1 (N17530, N17511);
and AND3 (N17531, N17527, N8109, N2891);
buf BUF1 (N17532, N17523);
and AND2 (N17533, N17524, N14152);
or OR4 (N17534, N17533, N7090, N9113, N17114);
nor NOR3 (N17535, N17489, N3147, N4379);
and AND3 (N17536, N17534, N4524, N8448);
nand NAND3 (N17537, N17531, N1412, N432);
and AND2 (N17538, N17536, N4157);
buf BUF1 (N17539, N17513);
nand NAND3 (N17540, N17528, N12259, N5085);
buf BUF1 (N17541, N17532);
and AND3 (N17542, N17539, N3460, N474);
xor XOR2 (N17543, N17542, N10538);
nand NAND2 (N17544, N17522, N1319);
nor NOR4 (N17545, N17529, N15807, N13057, N9293);
nor NOR3 (N17546, N17530, N7450, N13001);
nor NOR2 (N17547, N17545, N15564);
and AND2 (N17548, N17546, N8144);
nand NAND2 (N17549, N17538, N10420);
not NOT1 (N17550, N17544);
buf BUF1 (N17551, N17547);
or OR4 (N17552, N17540, N16681, N295, N11303);
nand NAND3 (N17553, N17551, N8970, N1877);
xor XOR2 (N17554, N17549, N13179);
xor XOR2 (N17555, N17553, N13511);
not NOT1 (N17556, N17537);
xor XOR2 (N17557, N17555, N13341);
or OR3 (N17558, N17557, N14420, N15565);
or OR2 (N17559, N17556, N3146);
nand NAND2 (N17560, N17526, N14944);
not NOT1 (N17561, N17560);
buf BUF1 (N17562, N17548);
or OR2 (N17563, N17543, N3898);
buf BUF1 (N17564, N17558);
not NOT1 (N17565, N17552);
buf BUF1 (N17566, N17561);
or OR3 (N17567, N17554, N5672, N9422);
nand NAND4 (N17568, N17567, N12767, N16098, N14309);
nor NOR4 (N17569, N17550, N898, N12716, N13927);
not NOT1 (N17570, N17564);
not NOT1 (N17571, N17541);
not NOT1 (N17572, N17569);
xor XOR2 (N17573, N17571, N2559);
nand NAND4 (N17574, N17563, N10328, N9639, N2734);
nor NOR2 (N17575, N17559, N8384);
or OR3 (N17576, N17562, N5690, N6705);
nand NAND3 (N17577, N17570, N3200, N4690);
or OR2 (N17578, N17573, N13973);
not NOT1 (N17579, N17577);
and AND4 (N17580, N17575, N3655, N15819, N8798);
and AND4 (N17581, N17565, N15278, N16809, N11015);
nand NAND4 (N17582, N17576, N12543, N2746, N4286);
nand NAND4 (N17583, N17574, N1745, N17017, N15267);
not NOT1 (N17584, N17582);
and AND4 (N17585, N17579, N6436, N3672, N7179);
xor XOR2 (N17586, N17572, N6603);
nor NOR2 (N17587, N17566, N3187);
buf BUF1 (N17588, N17585);
xor XOR2 (N17589, N17586, N4890);
nand NAND2 (N17590, N17583, N12681);
nand NAND2 (N17591, N17588, N1842);
xor XOR2 (N17592, N17535, N11310);
nor NOR2 (N17593, N17581, N17494);
nand NAND4 (N17594, N17580, N3455, N1674, N9694);
nor NOR3 (N17595, N17578, N11490, N10327);
xor XOR2 (N17596, N17595, N10548);
or OR2 (N17597, N17591, N9189);
and AND2 (N17598, N17590, N9819);
buf BUF1 (N17599, N17594);
nand NAND3 (N17600, N17597, N3132, N3598);
nor NOR2 (N17601, N17568, N10284);
and AND3 (N17602, N17598, N14295, N3355);
not NOT1 (N17603, N17593);
nand NAND4 (N17604, N17584, N4078, N6513, N15415);
and AND4 (N17605, N17599, N6332, N5982, N4364);
and AND3 (N17606, N17603, N390, N3745);
nand NAND4 (N17607, N17601, N7921, N4568, N7702);
and AND4 (N17608, N17596, N7069, N15069, N11234);
nand NAND4 (N17609, N17587, N8713, N13720, N1894);
xor XOR2 (N17610, N17592, N10770);
and AND2 (N17611, N17608, N1378);
buf BUF1 (N17612, N17611);
and AND2 (N17613, N17612, N14830);
or OR2 (N17614, N17602, N9138);
and AND3 (N17615, N17607, N13842, N14393);
buf BUF1 (N17616, N17600);
and AND4 (N17617, N17604, N12079, N7573, N140);
xor XOR2 (N17618, N17616, N7615);
xor XOR2 (N17619, N17589, N8792);
buf BUF1 (N17620, N17617);
nor NOR4 (N17621, N17619, N3633, N12606, N5372);
buf BUF1 (N17622, N17609);
not NOT1 (N17623, N17621);
xor XOR2 (N17624, N17606, N17515);
nor NOR2 (N17625, N17610, N15911);
not NOT1 (N17626, N17614);
not NOT1 (N17627, N17622);
xor XOR2 (N17628, N17605, N10531);
buf BUF1 (N17629, N17627);
and AND4 (N17630, N17623, N5140, N6387, N4072);
nand NAND4 (N17631, N17629, N7900, N11999, N6299);
and AND3 (N17632, N17615, N16807, N1853);
not NOT1 (N17633, N17628);
nor NOR3 (N17634, N17633, N15774, N6971);
and AND4 (N17635, N17620, N4649, N10146, N11046);
xor XOR2 (N17636, N17626, N16562);
or OR4 (N17637, N17624, N677, N7930, N14647);
and AND3 (N17638, N17634, N7015, N12634);
or OR3 (N17639, N17635, N6596, N1133);
nor NOR4 (N17640, N17630, N15437, N6151, N9347);
nor NOR4 (N17641, N17636, N13549, N5666, N11493);
nor NOR2 (N17642, N17618, N16244);
buf BUF1 (N17643, N17642);
nor NOR2 (N17644, N17643, N4056);
buf BUF1 (N17645, N17613);
nor NOR2 (N17646, N17641, N16728);
xor XOR2 (N17647, N17646, N13325);
buf BUF1 (N17648, N17637);
nor NOR4 (N17649, N17625, N11854, N11067, N2000);
not NOT1 (N17650, N17640);
nand NAND4 (N17651, N17644, N7986, N15527, N796);
nand NAND4 (N17652, N17650, N6711, N12217, N10959);
nor NOR3 (N17653, N17631, N3972, N5397);
not NOT1 (N17654, N17651);
and AND3 (N17655, N17653, N5640, N8105);
nand NAND3 (N17656, N17639, N4174, N3097);
and AND2 (N17657, N17632, N1471);
not NOT1 (N17658, N17649);
xor XOR2 (N17659, N17638, N16289);
not NOT1 (N17660, N17657);
nand NAND2 (N17661, N17652, N697);
buf BUF1 (N17662, N17647);
nor NOR2 (N17663, N17654, N12920);
xor XOR2 (N17664, N17645, N7835);
nand NAND4 (N17665, N17663, N3770, N10493, N16465);
not NOT1 (N17666, N17661);
nand NAND3 (N17667, N17660, N13622, N956);
not NOT1 (N17668, N17664);
nand NAND3 (N17669, N17662, N10270, N13666);
nor NOR4 (N17670, N17665, N14657, N9770, N2076);
nor NOR2 (N17671, N17667, N9322);
nor NOR4 (N17672, N17669, N15978, N4981, N11833);
nor NOR3 (N17673, N17648, N14830, N8815);
buf BUF1 (N17674, N17671);
not NOT1 (N17675, N17668);
nor NOR2 (N17676, N17655, N2664);
buf BUF1 (N17677, N17675);
xor XOR2 (N17678, N17673, N12838);
and AND4 (N17679, N17672, N11944, N10831, N16917);
not NOT1 (N17680, N17676);
nand NAND3 (N17681, N17679, N4992, N1425);
xor XOR2 (N17682, N17677, N1536);
or OR3 (N17683, N17678, N17238, N10145);
xor XOR2 (N17684, N17659, N8369);
not NOT1 (N17685, N17674);
buf BUF1 (N17686, N17670);
and AND3 (N17687, N17682, N13709, N9637);
nand NAND3 (N17688, N17683, N5275, N8722);
not NOT1 (N17689, N17684);
nor NOR4 (N17690, N17688, N15938, N15226, N6133);
nand NAND3 (N17691, N17681, N10338, N16953);
nor NOR2 (N17692, N17690, N14965);
nand NAND4 (N17693, N17691, N2346, N8575, N11428);
not NOT1 (N17694, N17692);
not NOT1 (N17695, N17687);
and AND3 (N17696, N17656, N16518, N7593);
nand NAND2 (N17697, N17695, N6064);
or OR3 (N17698, N17686, N2215, N17590);
or OR3 (N17699, N17693, N9987, N4672);
or OR2 (N17700, N17685, N15915);
buf BUF1 (N17701, N17696);
nor NOR3 (N17702, N17694, N7798, N17334);
or OR3 (N17703, N17680, N538, N15255);
nand NAND4 (N17704, N17658, N6163, N10681, N5383);
and AND2 (N17705, N17666, N7857);
nor NOR4 (N17706, N17705, N11259, N341, N11363);
nor NOR4 (N17707, N17703, N15446, N6588, N12573);
nand NAND3 (N17708, N17706, N6532, N4812);
xor XOR2 (N17709, N17698, N12491);
and AND4 (N17710, N17701, N11915, N3077, N7362);
xor XOR2 (N17711, N17707, N10149);
nor NOR3 (N17712, N17702, N15893, N7565);
not NOT1 (N17713, N17697);
xor XOR2 (N17714, N17711, N4380);
xor XOR2 (N17715, N17709, N5874);
nor NOR4 (N17716, N17712, N6052, N693, N8014);
xor XOR2 (N17717, N17699, N2931);
nand NAND3 (N17718, N17689, N7659, N2658);
buf BUF1 (N17719, N17718);
xor XOR2 (N17720, N17704, N13467);
and AND2 (N17721, N17717, N554);
xor XOR2 (N17722, N17715, N1172);
and AND3 (N17723, N17700, N4479, N15938);
xor XOR2 (N17724, N17721, N10114);
nor NOR3 (N17725, N17716, N11478, N10978);
xor XOR2 (N17726, N17724, N16165);
buf BUF1 (N17727, N17714);
or OR2 (N17728, N17722, N3073);
buf BUF1 (N17729, N17726);
buf BUF1 (N17730, N17708);
or OR2 (N17731, N17727, N7839);
buf BUF1 (N17732, N17713);
nand NAND4 (N17733, N17719, N59, N16469, N7825);
and AND2 (N17734, N17729, N1889);
nand NAND4 (N17735, N17728, N3291, N16665, N9338);
xor XOR2 (N17736, N17730, N4133);
not NOT1 (N17737, N17710);
not NOT1 (N17738, N17734);
or OR2 (N17739, N17733, N15459);
not NOT1 (N17740, N17732);
and AND4 (N17741, N17723, N10739, N107, N4178);
nor NOR4 (N17742, N17735, N844, N6297, N13587);
and AND2 (N17743, N17725, N7242);
nand NAND3 (N17744, N17737, N13558, N14083);
nor NOR2 (N17745, N17736, N2779);
xor XOR2 (N17746, N17742, N11021);
nand NAND4 (N17747, N17744, N4950, N9347, N11748);
xor XOR2 (N17748, N17740, N13459);
buf BUF1 (N17749, N17741);
and AND4 (N17750, N17739, N10150, N16899, N11554);
nand NAND4 (N17751, N17738, N9867, N2640, N7094);
or OR3 (N17752, N17731, N1037, N10136);
not NOT1 (N17753, N17720);
not NOT1 (N17754, N17747);
nand NAND2 (N17755, N17748, N2379);
xor XOR2 (N17756, N17755, N13342);
xor XOR2 (N17757, N17745, N13343);
nand NAND2 (N17758, N17746, N13481);
nand NAND3 (N17759, N17753, N17565, N4951);
buf BUF1 (N17760, N17754);
or OR4 (N17761, N17750, N5474, N3989, N17683);
or OR2 (N17762, N17758, N1900);
or OR2 (N17763, N17760, N11541);
nand NAND3 (N17764, N17749, N7501, N5969);
and AND4 (N17765, N17743, N11889, N12958, N12758);
not NOT1 (N17766, N17757);
xor XOR2 (N17767, N17756, N17542);
buf BUF1 (N17768, N17752);
or OR3 (N17769, N17766, N10319, N15310);
not NOT1 (N17770, N17768);
and AND3 (N17771, N17764, N3521, N7822);
nor NOR3 (N17772, N17765, N7267, N15839);
not NOT1 (N17773, N17772);
nor NOR2 (N17774, N17761, N5835);
and AND3 (N17775, N17769, N8644, N16947);
buf BUF1 (N17776, N17775);
xor XOR2 (N17777, N17771, N4741);
not NOT1 (N17778, N17773);
nand NAND4 (N17779, N17759, N6484, N16446, N15966);
nor NOR4 (N17780, N17779, N11108, N11755, N4423);
or OR3 (N17781, N17762, N7138, N7797);
and AND2 (N17782, N17780, N47);
xor XOR2 (N17783, N17782, N13054);
nand NAND4 (N17784, N17783, N16820, N4896, N5420);
xor XOR2 (N17785, N17781, N10160);
or OR4 (N17786, N17763, N13696, N5535, N2374);
nor NOR4 (N17787, N17770, N10095, N10696, N6428);
xor XOR2 (N17788, N17777, N8757);
nand NAND2 (N17789, N17787, N13605);
buf BUF1 (N17790, N17778);
not NOT1 (N17791, N17788);
nor NOR2 (N17792, N17784, N4041);
and AND2 (N17793, N17767, N1207);
or OR4 (N17794, N17793, N6813, N8780, N6896);
xor XOR2 (N17795, N17776, N13911);
or OR3 (N17796, N17795, N9260, N4309);
xor XOR2 (N17797, N17751, N13879);
nand NAND4 (N17798, N17792, N13453, N3488, N11870);
nor NOR3 (N17799, N17791, N4497, N12748);
or OR2 (N17800, N17774, N9044);
nor NOR3 (N17801, N17797, N382, N1882);
xor XOR2 (N17802, N17794, N9066);
xor XOR2 (N17803, N17790, N7703);
not NOT1 (N17804, N17798);
nor NOR4 (N17805, N17799, N10275, N9478, N12926);
xor XOR2 (N17806, N17802, N12576);
buf BUF1 (N17807, N17803);
or OR3 (N17808, N17796, N4275, N3773);
buf BUF1 (N17809, N17807);
buf BUF1 (N17810, N17800);
nor NOR3 (N17811, N17789, N5658, N9539);
nor NOR4 (N17812, N17809, N10866, N2496, N14569);
and AND2 (N17813, N17808, N11158);
or OR3 (N17814, N17806, N16411, N11605);
nor NOR2 (N17815, N17810, N8848);
nor NOR2 (N17816, N17804, N13729);
and AND2 (N17817, N17786, N13204);
xor XOR2 (N17818, N17812, N1377);
nand NAND3 (N17819, N17811, N7137, N8742);
and AND2 (N17820, N17805, N3461);
buf BUF1 (N17821, N17813);
xor XOR2 (N17822, N17785, N9875);
nor NOR3 (N17823, N17814, N6287, N1265);
nand NAND2 (N17824, N17801, N9655);
nand NAND4 (N17825, N17819, N17549, N8869, N13632);
xor XOR2 (N17826, N17818, N17602);
nand NAND3 (N17827, N17821, N14140, N7038);
not NOT1 (N17828, N17823);
and AND4 (N17829, N17828, N422, N8045, N11826);
nand NAND2 (N17830, N17829, N7540);
nor NOR2 (N17831, N17815, N5122);
or OR4 (N17832, N17826, N2619, N14208, N14653);
nor NOR3 (N17833, N17816, N5170, N11284);
buf BUF1 (N17834, N17817);
and AND3 (N17835, N17833, N9623, N1699);
or OR4 (N17836, N17825, N15253, N12336, N15281);
or OR4 (N17837, N17836, N15698, N1434, N15640);
xor XOR2 (N17838, N17837, N8601);
buf BUF1 (N17839, N17820);
nor NOR3 (N17840, N17835, N13391, N4872);
nor NOR2 (N17841, N17830, N2429);
and AND3 (N17842, N17824, N4670, N17323);
nor NOR3 (N17843, N17834, N4775, N1432);
and AND2 (N17844, N17832, N4966);
buf BUF1 (N17845, N17844);
nand NAND4 (N17846, N17841, N13795, N1511, N5511);
and AND4 (N17847, N17822, N16197, N16642, N5240);
nor NOR4 (N17848, N17842, N4707, N17561, N4272);
buf BUF1 (N17849, N17848);
nand NAND3 (N17850, N17831, N4965, N5112);
nand NAND3 (N17851, N17850, N13434, N10091);
and AND4 (N17852, N17843, N8072, N14863, N9142);
nand NAND4 (N17853, N17846, N12082, N916, N14657);
or OR4 (N17854, N17840, N14443, N7774, N14049);
not NOT1 (N17855, N17852);
and AND2 (N17856, N17851, N7361);
not NOT1 (N17857, N17854);
nor NOR4 (N17858, N17838, N5404, N2974, N7976);
nor NOR2 (N17859, N17827, N11204);
xor XOR2 (N17860, N17859, N9230);
nor NOR2 (N17861, N17845, N5351);
xor XOR2 (N17862, N17857, N10130);
nand NAND3 (N17863, N17856, N10697, N9010);
not NOT1 (N17864, N17847);
or OR4 (N17865, N17861, N6354, N14474, N10365);
or OR2 (N17866, N17863, N13515);
xor XOR2 (N17867, N17855, N7465);
not NOT1 (N17868, N17865);
nand NAND3 (N17869, N17866, N5576, N4992);
xor XOR2 (N17870, N17849, N14530);
or OR2 (N17871, N17860, N13696);
or OR3 (N17872, N17870, N12030, N14856);
or OR3 (N17873, N17872, N9132, N192);
or OR2 (N17874, N17868, N3225);
buf BUF1 (N17875, N17853);
nor NOR3 (N17876, N17873, N1538, N3235);
not NOT1 (N17877, N17869);
not NOT1 (N17878, N17876);
xor XOR2 (N17879, N17875, N16723);
nor NOR4 (N17880, N17862, N17223, N6523, N16288);
and AND4 (N17881, N17878, N7065, N16848, N6563);
not NOT1 (N17882, N17877);
or OR2 (N17883, N17867, N5242);
nand NAND4 (N17884, N17858, N11880, N5232, N2162);
not NOT1 (N17885, N17839);
buf BUF1 (N17886, N17871);
xor XOR2 (N17887, N17879, N10686);
nor NOR2 (N17888, N17885, N5798);
buf BUF1 (N17889, N17864);
and AND2 (N17890, N17888, N14780);
not NOT1 (N17891, N17890);
buf BUF1 (N17892, N17882);
nand NAND2 (N17893, N17880, N5992);
xor XOR2 (N17894, N17893, N420);
and AND4 (N17895, N17881, N1563, N4702, N7077);
nand NAND2 (N17896, N17892, N13169);
and AND4 (N17897, N17891, N16849, N10916, N7311);
xor XOR2 (N17898, N17897, N9995);
buf BUF1 (N17899, N17884);
and AND4 (N17900, N17889, N9936, N17466, N3240);
or OR2 (N17901, N17874, N16641);
or OR2 (N17902, N17883, N16621);
not NOT1 (N17903, N17894);
nor NOR3 (N17904, N17896, N14483, N4278);
nand NAND4 (N17905, N17904, N8980, N4849, N14233);
and AND4 (N17906, N17887, N14848, N7382, N6281);
and AND4 (N17907, N17901, N5836, N17791, N13192);
nand NAND4 (N17908, N17907, N1262, N13449, N2399);
nand NAND4 (N17909, N17900, N5038, N3470, N7388);
nand NAND4 (N17910, N17908, N14888, N2570, N3423);
nand NAND2 (N17911, N17905, N3309);
and AND3 (N17912, N17910, N12415, N13193);
or OR2 (N17913, N17902, N17134);
or OR2 (N17914, N17913, N6352);
or OR3 (N17915, N17898, N1180, N5407);
xor XOR2 (N17916, N17899, N4331);
buf BUF1 (N17917, N17912);
nand NAND4 (N17918, N17895, N10433, N6610, N6661);
nor NOR2 (N17919, N17886, N13458);
nor NOR4 (N17920, N17911, N12856, N3206, N261);
or OR3 (N17921, N17919, N13240, N311);
and AND2 (N17922, N17918, N10632);
and AND2 (N17923, N17921, N10947);
nor NOR4 (N17924, N17922, N7778, N7183, N13449);
not NOT1 (N17925, N17916);
or OR3 (N17926, N17923, N2869, N1392);
not NOT1 (N17927, N17926);
xor XOR2 (N17928, N17909, N15490);
or OR2 (N17929, N17903, N852);
nand NAND4 (N17930, N17924, N7124, N9374, N12018);
and AND2 (N17931, N17920, N17228);
buf BUF1 (N17932, N17931);
not NOT1 (N17933, N17917);
buf BUF1 (N17934, N17914);
nor NOR4 (N17935, N17915, N6036, N5718, N9346);
xor XOR2 (N17936, N17927, N7352);
or OR3 (N17937, N17932, N3732, N2885);
xor XOR2 (N17938, N17925, N911);
or OR4 (N17939, N17929, N8671, N3225, N11455);
not NOT1 (N17940, N17939);
buf BUF1 (N17941, N17906);
and AND2 (N17942, N17936, N9811);
nor NOR4 (N17943, N17941, N9958, N16850, N8104);
or OR3 (N17944, N17940, N6711, N12277);
and AND4 (N17945, N17928, N6428, N9594, N10109);
and AND4 (N17946, N17945, N17866, N11832, N13464);
not NOT1 (N17947, N17937);
nand NAND2 (N17948, N17938, N4160);
or OR4 (N17949, N17935, N6350, N6146, N6612);
or OR3 (N17950, N17948, N14, N4357);
xor XOR2 (N17951, N17933, N2096);
and AND3 (N17952, N17934, N4547, N2556);
nor NOR2 (N17953, N17930, N16703);
not NOT1 (N17954, N17947);
xor XOR2 (N17955, N17946, N9602);
or OR4 (N17956, N17952, N16379, N11372, N2824);
or OR2 (N17957, N17942, N11443);
buf BUF1 (N17958, N17957);
and AND3 (N17959, N17956, N810, N9794);
nand NAND2 (N17960, N17955, N511);
and AND2 (N17961, N17944, N16458);
not NOT1 (N17962, N17943);
nor NOR4 (N17963, N17949, N1513, N10463, N7699);
nor NOR2 (N17964, N17961, N16740);
not NOT1 (N17965, N17963);
nor NOR2 (N17966, N17959, N15067);
and AND2 (N17967, N17964, N8486);
and AND3 (N17968, N17954, N3154, N12437);
or OR4 (N17969, N17960, N1855, N11785, N5237);
and AND3 (N17970, N17950, N16451, N10939);
xor XOR2 (N17971, N17970, N13018);
or OR3 (N17972, N17971, N5363, N13315);
not NOT1 (N17973, N17953);
nor NOR2 (N17974, N17968, N13459);
or OR4 (N17975, N17969, N2202, N11835, N5064);
and AND2 (N17976, N17962, N11726);
or OR4 (N17977, N17951, N5154, N840, N1813);
not NOT1 (N17978, N17973);
buf BUF1 (N17979, N17972);
buf BUF1 (N17980, N17965);
not NOT1 (N17981, N17975);
buf BUF1 (N17982, N17958);
nor NOR4 (N17983, N17981, N4772, N15211, N4836);
nor NOR3 (N17984, N17980, N15841, N13452);
and AND2 (N17985, N17974, N13206);
nor NOR2 (N17986, N17967, N4376);
nor NOR3 (N17987, N17982, N917, N12217);
nor NOR3 (N17988, N17983, N8825, N6056);
nand NAND2 (N17989, N17976, N7445);
not NOT1 (N17990, N17988);
nor NOR2 (N17991, N17989, N5170);
nand NAND2 (N17992, N17991, N9346);
or OR2 (N17993, N17979, N119);
xor XOR2 (N17994, N17990, N13366);
nand NAND4 (N17995, N17977, N12203, N2142, N4657);
nand NAND2 (N17996, N17995, N10474);
buf BUF1 (N17997, N17984);
nor NOR2 (N17998, N17992, N17273);
buf BUF1 (N17999, N17978);
or OR3 (N18000, N17966, N9666, N17230);
or OR2 (N18001, N17987, N13866);
or OR4 (N18002, N17985, N17265, N2377, N1998);
not NOT1 (N18003, N17993);
and AND2 (N18004, N18002, N11202);
not NOT1 (N18005, N17997);
and AND2 (N18006, N18005, N11140);
not NOT1 (N18007, N17996);
nor NOR3 (N18008, N17994, N1159, N2269);
not NOT1 (N18009, N18008);
and AND3 (N18010, N18009, N17104, N15581);
or OR2 (N18011, N18010, N7741);
xor XOR2 (N18012, N17999, N6140);
not NOT1 (N18013, N17998);
buf BUF1 (N18014, N18003);
nand NAND4 (N18015, N18006, N11658, N1578, N8549);
or OR3 (N18016, N18011, N7030, N10270);
buf BUF1 (N18017, N18004);
or OR4 (N18018, N18001, N10695, N14821, N11130);
xor XOR2 (N18019, N18014, N14329);
nand NAND4 (N18020, N17986, N13081, N3938, N17931);
buf BUF1 (N18021, N18018);
xor XOR2 (N18022, N18021, N385);
xor XOR2 (N18023, N18012, N8985);
nand NAND4 (N18024, N18023, N15893, N11551, N1947);
nor NOR4 (N18025, N18019, N8310, N13461, N4983);
buf BUF1 (N18026, N18017);
or OR2 (N18027, N18016, N781);
or OR3 (N18028, N18000, N11856, N14578);
nand NAND2 (N18029, N18022, N4694);
xor XOR2 (N18030, N18029, N7386);
or OR3 (N18031, N18027, N16374, N1119);
buf BUF1 (N18032, N18013);
xor XOR2 (N18033, N18024, N16606);
not NOT1 (N18034, N18026);
and AND4 (N18035, N18025, N14120, N186, N17256);
nand NAND4 (N18036, N18035, N14901, N436, N3825);
xor XOR2 (N18037, N18032, N3626);
buf BUF1 (N18038, N18015);
not NOT1 (N18039, N18034);
not NOT1 (N18040, N18038);
xor XOR2 (N18041, N18007, N15761);
xor XOR2 (N18042, N18039, N5800);
nand NAND2 (N18043, N18036, N2925);
buf BUF1 (N18044, N18037);
buf BUF1 (N18045, N18042);
and AND2 (N18046, N18028, N6547);
or OR4 (N18047, N18020, N10527, N4667, N2634);
and AND4 (N18048, N18044, N528, N7280, N11687);
nand NAND4 (N18049, N18045, N9508, N3485, N6182);
nand NAND3 (N18050, N18046, N10348, N18021);
and AND2 (N18051, N18049, N12871);
or OR3 (N18052, N18048, N9990, N8574);
xor XOR2 (N18053, N18052, N11117);
not NOT1 (N18054, N18053);
or OR2 (N18055, N18051, N2151);
buf BUF1 (N18056, N18040);
buf BUF1 (N18057, N18054);
xor XOR2 (N18058, N18031, N1877);
or OR3 (N18059, N18041, N15766, N17782);
or OR4 (N18060, N18055, N652, N11910, N4597);
nor NOR2 (N18061, N18033, N9950);
buf BUF1 (N18062, N18061);
and AND4 (N18063, N18059, N10737, N12982, N8537);
or OR4 (N18064, N18058, N727, N3343, N16168);
nor NOR3 (N18065, N18057, N4655, N12273);
or OR2 (N18066, N18050, N3042);
or OR4 (N18067, N18056, N12760, N2379, N10538);
or OR4 (N18068, N18043, N10628, N10200, N12559);
not NOT1 (N18069, N18067);
buf BUF1 (N18070, N18062);
xor XOR2 (N18071, N18063, N7031);
buf BUF1 (N18072, N18065);
xor XOR2 (N18073, N18070, N6879);
xor XOR2 (N18074, N18030, N994);
not NOT1 (N18075, N18047);
not NOT1 (N18076, N18075);
or OR2 (N18077, N18069, N9224);
not NOT1 (N18078, N18064);
or OR3 (N18079, N18073, N9689, N13232);
nor NOR4 (N18080, N18078, N8829, N11382, N4480);
not NOT1 (N18081, N18060);
nor NOR2 (N18082, N18068, N16625);
not NOT1 (N18083, N18074);
buf BUF1 (N18084, N18066);
xor XOR2 (N18085, N18084, N8116);
or OR3 (N18086, N18079, N11909, N551);
xor XOR2 (N18087, N18083, N3753);
nand NAND4 (N18088, N18076, N6498, N4823, N15853);
xor XOR2 (N18089, N18085, N5134);
not NOT1 (N18090, N18086);
buf BUF1 (N18091, N18080);
buf BUF1 (N18092, N18087);
nor NOR4 (N18093, N18081, N5336, N17644, N4991);
not NOT1 (N18094, N18092);
nand NAND4 (N18095, N18071, N5490, N9892, N11477);
and AND4 (N18096, N18095, N6473, N3018, N10650);
not NOT1 (N18097, N18096);
or OR2 (N18098, N18088, N7118);
not NOT1 (N18099, N18094);
or OR3 (N18100, N18099, N5653, N3399);
nand NAND4 (N18101, N18089, N14069, N18057, N4412);
not NOT1 (N18102, N18072);
not NOT1 (N18103, N18101);
or OR4 (N18104, N18097, N11761, N6361, N3805);
nor NOR4 (N18105, N18091, N6935, N8823, N3966);
nand NAND4 (N18106, N18090, N5710, N938, N4835);
not NOT1 (N18107, N18100);
not NOT1 (N18108, N18102);
nor NOR3 (N18109, N18106, N16541, N7559);
or OR4 (N18110, N18109, N4424, N2612, N16470);
nor NOR4 (N18111, N18104, N18025, N5853, N16172);
nor NOR4 (N18112, N18103, N13484, N16069, N9967);
nand NAND4 (N18113, N18105, N4404, N6709, N7462);
xor XOR2 (N18114, N18098, N13192);
nand NAND3 (N18115, N18093, N2681, N13240);
buf BUF1 (N18116, N18113);
xor XOR2 (N18117, N18114, N1805);
not NOT1 (N18118, N18082);
nor NOR3 (N18119, N18077, N16994, N17541);
and AND2 (N18120, N18108, N1764);
and AND2 (N18121, N18120, N12047);
not NOT1 (N18122, N18119);
nor NOR3 (N18123, N18122, N11036, N11824);
nand NAND4 (N18124, N18117, N15927, N277, N17783);
and AND2 (N18125, N18115, N6948);
xor XOR2 (N18126, N18118, N2018);
and AND2 (N18127, N18110, N8812);
buf BUF1 (N18128, N18127);
nand NAND4 (N18129, N18112, N752, N16204, N1569);
nand NAND2 (N18130, N18107, N18035);
nor NOR2 (N18131, N18129, N14599);
nand NAND3 (N18132, N18128, N3901, N3216);
or OR2 (N18133, N18123, N11776);
not NOT1 (N18134, N18131);
nand NAND2 (N18135, N18130, N4759);
and AND4 (N18136, N18135, N284, N1858, N9423);
nand NAND2 (N18137, N18136, N18084);
or OR3 (N18138, N18137, N11678, N9980);
nand NAND2 (N18139, N18134, N10568);
not NOT1 (N18140, N18132);
buf BUF1 (N18141, N18111);
or OR4 (N18142, N18121, N3788, N7726, N17727);
nand NAND2 (N18143, N18142, N8530);
buf BUF1 (N18144, N18116);
nor NOR3 (N18145, N18140, N13653, N12552);
nand NAND2 (N18146, N18126, N16690);
not NOT1 (N18147, N18141);
buf BUF1 (N18148, N18144);
not NOT1 (N18149, N18146);
nor NOR4 (N18150, N18133, N2070, N8988, N766);
not NOT1 (N18151, N18150);
nand NAND2 (N18152, N18125, N644);
xor XOR2 (N18153, N18139, N31);
xor XOR2 (N18154, N18145, N14984);
and AND4 (N18155, N18147, N8451, N15312, N11793);
nor NOR3 (N18156, N18138, N123, N882);
and AND4 (N18157, N18153, N2791, N15388, N3378);
and AND3 (N18158, N18154, N8623, N2813);
xor XOR2 (N18159, N18151, N3642);
not NOT1 (N18160, N18155);
buf BUF1 (N18161, N18158);
nor NOR2 (N18162, N18152, N5758);
not NOT1 (N18163, N18156);
not NOT1 (N18164, N18143);
nand NAND3 (N18165, N18148, N2576, N1489);
and AND3 (N18166, N18149, N9126, N10840);
or OR3 (N18167, N18164, N14304, N1316);
nor NOR4 (N18168, N18160, N9012, N9038, N13590);
or OR4 (N18169, N18159, N14944, N12125, N11306);
and AND3 (N18170, N18124, N14926, N5215);
or OR3 (N18171, N18162, N7166, N9001);
xor XOR2 (N18172, N18167, N13791);
not NOT1 (N18173, N18172);
and AND2 (N18174, N18173, N6407);
buf BUF1 (N18175, N18165);
nand NAND4 (N18176, N18168, N3470, N2437, N12506);
nor NOR3 (N18177, N18174, N17730, N10110);
not NOT1 (N18178, N18157);
nor NOR4 (N18179, N18175, N12737, N2468, N9371);
xor XOR2 (N18180, N18176, N17530);
nor NOR3 (N18181, N18177, N2719, N3131);
nor NOR2 (N18182, N18169, N6602);
nand NAND3 (N18183, N18163, N5863, N9130);
xor XOR2 (N18184, N18183, N3965);
nand NAND2 (N18185, N18180, N2965);
nor NOR2 (N18186, N18178, N1071);
nand NAND3 (N18187, N18185, N7998, N16794);
not NOT1 (N18188, N18186);
not NOT1 (N18189, N18171);
and AND3 (N18190, N18161, N11701, N1221);
nor NOR2 (N18191, N18182, N17206);
buf BUF1 (N18192, N18187);
buf BUF1 (N18193, N18191);
nor NOR2 (N18194, N18192, N1358);
nor NOR2 (N18195, N18179, N3111);
xor XOR2 (N18196, N18181, N1809);
xor XOR2 (N18197, N18193, N6350);
nor NOR3 (N18198, N18184, N9299, N8922);
not NOT1 (N18199, N18196);
and AND2 (N18200, N18199, N14857);
nand NAND3 (N18201, N18189, N14589, N1005);
and AND4 (N18202, N18190, N16944, N12174, N16364);
buf BUF1 (N18203, N18188);
buf BUF1 (N18204, N18202);
and AND4 (N18205, N18194, N14514, N6227, N16877);
and AND3 (N18206, N18198, N9736, N3463);
or OR4 (N18207, N18204, N7636, N17052, N4015);
and AND3 (N18208, N18170, N2450, N8121);
or OR3 (N18209, N18166, N10362, N3515);
xor XOR2 (N18210, N18207, N11873);
not NOT1 (N18211, N18205);
xor XOR2 (N18212, N18195, N7850);
nor NOR4 (N18213, N18212, N2476, N5725, N574);
or OR4 (N18214, N18203, N10288, N15701, N9938);
xor XOR2 (N18215, N18211, N13166);
not NOT1 (N18216, N18206);
nor NOR4 (N18217, N18208, N8902, N2741, N5521);
and AND3 (N18218, N18216, N16939, N862);
or OR2 (N18219, N18213, N1460);
nor NOR4 (N18220, N18209, N5588, N11639, N15361);
and AND3 (N18221, N18200, N10324, N535);
or OR3 (N18222, N18217, N7594, N12059);
nor NOR3 (N18223, N18214, N3743, N6835);
nand NAND2 (N18224, N18215, N4674);
not NOT1 (N18225, N18220);
xor XOR2 (N18226, N18224, N4679);
and AND2 (N18227, N18201, N11526);
xor XOR2 (N18228, N18221, N6981);
not NOT1 (N18229, N18222);
buf BUF1 (N18230, N18225);
and AND3 (N18231, N18227, N3169, N4736);
xor XOR2 (N18232, N18219, N8992);
buf BUF1 (N18233, N18229);
not NOT1 (N18234, N18231);
and AND3 (N18235, N18233, N11742, N10418);
and AND3 (N18236, N18228, N11510, N8351);
buf BUF1 (N18237, N18236);
nor NOR2 (N18238, N18230, N8673);
buf BUF1 (N18239, N18238);
not NOT1 (N18240, N18234);
buf BUF1 (N18241, N18237);
and AND4 (N18242, N18240, N16412, N5792, N11417);
not NOT1 (N18243, N18210);
nor NOR3 (N18244, N18232, N14342, N8037);
buf BUF1 (N18245, N18197);
not NOT1 (N18246, N18242);
nand NAND2 (N18247, N18246, N3581);
xor XOR2 (N18248, N18241, N4180);
buf BUF1 (N18249, N18218);
buf BUF1 (N18250, N18239);
and AND2 (N18251, N18249, N11221);
not NOT1 (N18252, N18235);
nor NOR4 (N18253, N18251, N2545, N4715, N2365);
buf BUF1 (N18254, N18253);
xor XOR2 (N18255, N18243, N2682);
not NOT1 (N18256, N18245);
or OR4 (N18257, N18256, N14139, N15739, N4249);
not NOT1 (N18258, N18244);
buf BUF1 (N18259, N18252);
nand NAND3 (N18260, N18254, N16861, N7321);
and AND4 (N18261, N18248, N2, N15066, N16143);
or OR3 (N18262, N18223, N17551, N4367);
nor NOR4 (N18263, N18261, N527, N16344, N5138);
xor XOR2 (N18264, N18259, N14445);
xor XOR2 (N18265, N18264, N4385);
or OR3 (N18266, N18263, N10559, N15276);
buf BUF1 (N18267, N18258);
or OR4 (N18268, N18262, N8408, N4212, N6064);
not NOT1 (N18269, N18268);
buf BUF1 (N18270, N18257);
and AND2 (N18271, N18260, N12);
and AND4 (N18272, N18271, N6367, N5316, N11595);
or OR2 (N18273, N18226, N12359);
nor NOR2 (N18274, N18272, N8963);
xor XOR2 (N18275, N18273, N9990);
xor XOR2 (N18276, N18247, N2615);
nand NAND4 (N18277, N18267, N12565, N11104, N16238);
and AND3 (N18278, N18269, N9512, N13551);
or OR2 (N18279, N18276, N1268);
buf BUF1 (N18280, N18274);
and AND3 (N18281, N18266, N790, N11124);
nand NAND2 (N18282, N18278, N5655);
nor NOR2 (N18283, N18275, N6105);
and AND2 (N18284, N18255, N18051);
nor NOR2 (N18285, N18277, N9668);
or OR4 (N18286, N18250, N13620, N3835, N6343);
nand NAND4 (N18287, N18270, N13478, N15267, N14688);
buf BUF1 (N18288, N18285);
not NOT1 (N18289, N18282);
xor XOR2 (N18290, N18265, N15476);
nand NAND2 (N18291, N18289, N10802);
or OR2 (N18292, N18287, N17588);
and AND3 (N18293, N18281, N11055, N8806);
and AND3 (N18294, N18279, N3989, N6515);
nor NOR4 (N18295, N18293, N9478, N16794, N5310);
xor XOR2 (N18296, N18286, N7974);
buf BUF1 (N18297, N18283);
or OR2 (N18298, N18290, N3589);
nand NAND4 (N18299, N18297, N17528, N3080, N663);
nand NAND2 (N18300, N18298, N2875);
nor NOR2 (N18301, N18280, N1452);
nand NAND3 (N18302, N18284, N13548, N7346);
xor XOR2 (N18303, N18302, N586);
xor XOR2 (N18304, N18300, N7931);
not NOT1 (N18305, N18291);
xor XOR2 (N18306, N18292, N8198);
nand NAND4 (N18307, N18295, N6164, N9684, N3602);
nand NAND2 (N18308, N18294, N7846);
nor NOR2 (N18309, N18296, N9932);
nand NAND4 (N18310, N18303, N4154, N2669, N6180);
nor NOR2 (N18311, N18306, N12298);
and AND2 (N18312, N18305, N6094);
buf BUF1 (N18313, N18288);
xor XOR2 (N18314, N18312, N13520);
not NOT1 (N18315, N18310);
and AND3 (N18316, N18308, N15307, N13006);
buf BUF1 (N18317, N18309);
buf BUF1 (N18318, N18311);
buf BUF1 (N18319, N18314);
not NOT1 (N18320, N18304);
and AND3 (N18321, N18301, N15364, N11516);
nand NAND3 (N18322, N18320, N3454, N4321);
or OR3 (N18323, N18316, N11184, N16946);
buf BUF1 (N18324, N18323);
and AND4 (N18325, N18315, N3739, N15214, N5330);
not NOT1 (N18326, N18325);
not NOT1 (N18327, N18319);
xor XOR2 (N18328, N18321, N3239);
and AND2 (N18329, N18299, N14498);
or OR4 (N18330, N18326, N7905, N6118, N5630);
nand NAND2 (N18331, N18313, N13365);
nor NOR4 (N18332, N18329, N15529, N1283, N13524);
nand NAND3 (N18333, N18331, N3259, N15866);
xor XOR2 (N18334, N18318, N4811);
xor XOR2 (N18335, N18334, N13350);
buf BUF1 (N18336, N18332);
not NOT1 (N18337, N18322);
and AND4 (N18338, N18327, N562, N16828, N4118);
buf BUF1 (N18339, N18333);
buf BUF1 (N18340, N18330);
and AND4 (N18341, N18339, N15080, N5476, N15776);
or OR3 (N18342, N18338, N5134, N12212);
xor XOR2 (N18343, N18337, N11683);
and AND3 (N18344, N18335, N10940, N1497);
xor XOR2 (N18345, N18307, N13086);
and AND4 (N18346, N18336, N13969, N11035, N7771);
buf BUF1 (N18347, N18328);
xor XOR2 (N18348, N18324, N13432);
not NOT1 (N18349, N18348);
or OR2 (N18350, N18349, N32);
buf BUF1 (N18351, N18340);
buf BUF1 (N18352, N18317);
nand NAND2 (N18353, N18350, N12475);
nor NOR2 (N18354, N18353, N3877);
or OR4 (N18355, N18344, N12898, N11205, N7587);
nor NOR2 (N18356, N18343, N310);
and AND2 (N18357, N18341, N5817);
nand NAND4 (N18358, N18354, N17807, N12981, N6931);
nand NAND2 (N18359, N18357, N1608);
nor NOR2 (N18360, N18345, N2520);
not NOT1 (N18361, N18355);
nor NOR2 (N18362, N18358, N14694);
nor NOR2 (N18363, N18352, N8332);
xor XOR2 (N18364, N18360, N11741);
nand NAND2 (N18365, N18351, N4309);
xor XOR2 (N18366, N18346, N17059);
nand NAND2 (N18367, N18365, N8968);
or OR4 (N18368, N18364, N7593, N18340, N13914);
nor NOR3 (N18369, N18366, N7533, N2835);
nand NAND3 (N18370, N18342, N6084, N6604);
and AND4 (N18371, N18347, N1848, N3689, N5471);
nor NOR2 (N18372, N18359, N12671);
xor XOR2 (N18373, N18362, N1581);
nor NOR2 (N18374, N18373, N12606);
and AND4 (N18375, N18356, N9137, N11594, N10498);
nand NAND3 (N18376, N18369, N807, N11859);
nor NOR2 (N18377, N18374, N10824);
and AND2 (N18378, N18363, N4093);
nor NOR4 (N18379, N18372, N2302, N3697, N8693);
buf BUF1 (N18380, N18378);
nand NAND2 (N18381, N18368, N15511);
buf BUF1 (N18382, N18370);
buf BUF1 (N18383, N18380);
not NOT1 (N18384, N18377);
xor XOR2 (N18385, N18379, N2945);
buf BUF1 (N18386, N18376);
and AND3 (N18387, N18381, N7847, N14175);
nor NOR2 (N18388, N18387, N2142);
buf BUF1 (N18389, N18383);
not NOT1 (N18390, N18385);
nor NOR3 (N18391, N18390, N6775, N15729);
nor NOR3 (N18392, N18384, N14821, N9486);
xor XOR2 (N18393, N18392, N16130);
nor NOR2 (N18394, N18386, N3884);
or OR3 (N18395, N18367, N11637, N1341);
or OR3 (N18396, N18388, N2263, N11106);
or OR4 (N18397, N18361, N12568, N15427, N1640);
nand NAND4 (N18398, N18371, N6871, N6229, N4);
buf BUF1 (N18399, N18398);
nand NAND4 (N18400, N18391, N10430, N4197, N14835);
xor XOR2 (N18401, N18389, N427);
nor NOR3 (N18402, N18401, N17689, N920);
not NOT1 (N18403, N18396);
and AND2 (N18404, N18395, N10782);
or OR2 (N18405, N18393, N5430);
xor XOR2 (N18406, N18394, N3460);
not NOT1 (N18407, N18382);
nor NOR2 (N18408, N18404, N16779);
nand NAND2 (N18409, N18397, N558);
or OR2 (N18410, N18408, N985);
buf BUF1 (N18411, N18406);
nor NOR3 (N18412, N18409, N11838, N14747);
nand NAND3 (N18413, N18410, N15984, N10824);
nand NAND4 (N18414, N18407, N14588, N2601, N2547);
nor NOR2 (N18415, N18400, N5812);
or OR4 (N18416, N18412, N5425, N2190, N16765);
or OR4 (N18417, N18375, N17034, N6719, N10739);
not NOT1 (N18418, N18413);
nand NAND4 (N18419, N18415, N11676, N913, N2782);
or OR2 (N18420, N18414, N15213);
or OR4 (N18421, N18402, N3881, N18329, N13188);
xor XOR2 (N18422, N18419, N16796);
or OR4 (N18423, N18405, N9423, N1375, N13043);
or OR2 (N18424, N18422, N10788);
xor XOR2 (N18425, N18418, N12015);
buf BUF1 (N18426, N18416);
not NOT1 (N18427, N18424);
not NOT1 (N18428, N18399);
or OR4 (N18429, N18403, N5823, N11679, N16451);
not NOT1 (N18430, N18425);
buf BUF1 (N18431, N18426);
xor XOR2 (N18432, N18411, N12708);
xor XOR2 (N18433, N18430, N12795);
xor XOR2 (N18434, N18429, N7267);
or OR4 (N18435, N18423, N15993, N16810, N10300);
xor XOR2 (N18436, N18432, N7460);
not NOT1 (N18437, N18417);
nor NOR2 (N18438, N18428, N15708);
and AND2 (N18439, N18421, N15702);
and AND3 (N18440, N18434, N7248, N7888);
buf BUF1 (N18441, N18427);
not NOT1 (N18442, N18441);
buf BUF1 (N18443, N18433);
or OR2 (N18444, N18438, N14149);
buf BUF1 (N18445, N18443);
not NOT1 (N18446, N18445);
nor NOR4 (N18447, N18436, N13511, N2747, N11227);
nor NOR4 (N18448, N18440, N6138, N8928, N17179);
nor NOR3 (N18449, N18448, N9073, N12875);
xor XOR2 (N18450, N18420, N7324);
and AND2 (N18451, N18437, N933);
xor XOR2 (N18452, N18450, N16893);
not NOT1 (N18453, N18449);
nor NOR4 (N18454, N18452, N8716, N6209, N7347);
xor XOR2 (N18455, N18447, N10296);
or OR3 (N18456, N18439, N15801, N2413);
nand NAND3 (N18457, N18444, N759, N4534);
or OR4 (N18458, N18454, N17038, N6991, N9474);
not NOT1 (N18459, N18442);
nand NAND2 (N18460, N18431, N4046);
and AND2 (N18461, N18460, N6214);
buf BUF1 (N18462, N18451);
not NOT1 (N18463, N18456);
or OR2 (N18464, N18457, N2964);
nor NOR4 (N18465, N18435, N12358, N12084, N9190);
xor XOR2 (N18466, N18459, N4639);
nand NAND2 (N18467, N18462, N1998);
and AND3 (N18468, N18461, N1347, N7343);
and AND2 (N18469, N18468, N7579);
xor XOR2 (N18470, N18467, N8519);
nor NOR4 (N18471, N18455, N1932, N6688, N910);
not NOT1 (N18472, N18470);
buf BUF1 (N18473, N18463);
or OR3 (N18474, N18453, N2323, N2190);
or OR2 (N18475, N18469, N11330);
buf BUF1 (N18476, N18473);
not NOT1 (N18477, N18474);
and AND2 (N18478, N18458, N5908);
nand NAND3 (N18479, N18464, N841, N6669);
and AND3 (N18480, N18479, N1950, N16343);
and AND2 (N18481, N18472, N17974);
or OR3 (N18482, N18466, N13525, N10000);
nor NOR2 (N18483, N18478, N13911);
buf BUF1 (N18484, N18476);
buf BUF1 (N18485, N18480);
xor XOR2 (N18486, N18483, N5179);
nand NAND3 (N18487, N18484, N7972, N10522);
nor NOR4 (N18488, N18471, N15330, N13352, N8506);
buf BUF1 (N18489, N18486);
and AND4 (N18490, N18485, N8347, N18341, N1304);
nand NAND3 (N18491, N18490, N3985, N6822);
or OR3 (N18492, N18482, N17497, N6529);
not NOT1 (N18493, N18488);
and AND3 (N18494, N18487, N1512, N3780);
buf BUF1 (N18495, N18493);
nor NOR4 (N18496, N18475, N16513, N14261, N17502);
buf BUF1 (N18497, N18446);
nor NOR4 (N18498, N18489, N1379, N14514, N1306);
and AND3 (N18499, N18477, N11910, N159);
xor XOR2 (N18500, N18492, N9740);
and AND4 (N18501, N18465, N1292, N6100, N8646);
not NOT1 (N18502, N18494);
and AND3 (N18503, N18481, N6139, N9445);
buf BUF1 (N18504, N18498);
buf BUF1 (N18505, N18496);
and AND3 (N18506, N18503, N14477, N5183);
not NOT1 (N18507, N18500);
and AND4 (N18508, N18495, N17414, N5375, N761);
nand NAND3 (N18509, N18501, N3074, N6966);
and AND4 (N18510, N18507, N4494, N1955, N7103);
buf BUF1 (N18511, N18506);
or OR3 (N18512, N18497, N7637, N17439);
nand NAND4 (N18513, N18511, N5416, N11251, N2532);
or OR2 (N18514, N18510, N8259);
nor NOR3 (N18515, N18491, N2157, N15136);
and AND2 (N18516, N18505, N9925);
xor XOR2 (N18517, N18515, N2118);
buf BUF1 (N18518, N18499);
xor XOR2 (N18519, N18508, N10026);
nand NAND2 (N18520, N18502, N3264);
or OR4 (N18521, N18512, N15162, N2816, N9409);
not NOT1 (N18522, N18513);
or OR3 (N18523, N18514, N4607, N3392);
nor NOR2 (N18524, N18521, N9145);
xor XOR2 (N18525, N18523, N1133);
buf BUF1 (N18526, N18524);
nand NAND4 (N18527, N18518, N17945, N7409, N12353);
buf BUF1 (N18528, N18517);
buf BUF1 (N18529, N18522);
or OR2 (N18530, N18516, N9546);
xor XOR2 (N18531, N18527, N10451);
or OR3 (N18532, N18526, N5573, N926);
or OR3 (N18533, N18525, N13911, N9730);
nand NAND3 (N18534, N18520, N8353, N11320);
xor XOR2 (N18535, N18528, N9137);
nand NAND3 (N18536, N18529, N16190, N14317);
nor NOR4 (N18537, N18531, N10479, N3164, N10479);
not NOT1 (N18538, N18535);
nand NAND4 (N18539, N18534, N11190, N16188, N13897);
or OR2 (N18540, N18536, N10697);
nand NAND2 (N18541, N18504, N7413);
nand NAND3 (N18542, N18533, N11347, N1276);
or OR4 (N18543, N18530, N6225, N4144, N9608);
and AND3 (N18544, N18519, N3969, N10561);
or OR2 (N18545, N18537, N9012);
xor XOR2 (N18546, N18541, N11842);
nand NAND3 (N18547, N18532, N9232, N3650);
and AND3 (N18548, N18543, N14161, N7364);
and AND4 (N18549, N18540, N5300, N13407, N14882);
not NOT1 (N18550, N18549);
not NOT1 (N18551, N18548);
and AND2 (N18552, N18544, N13164);
nand NAND2 (N18553, N18551, N1299);
and AND3 (N18554, N18550, N13194, N3443);
xor XOR2 (N18555, N18542, N12996);
and AND4 (N18556, N18553, N10945, N12885, N4187);
nand NAND3 (N18557, N18547, N2522, N207);
and AND2 (N18558, N18545, N14577);
and AND3 (N18559, N18554, N4182, N11019);
not NOT1 (N18560, N18559);
buf BUF1 (N18561, N18560);
nand NAND4 (N18562, N18546, N15631, N2002, N3695);
or OR2 (N18563, N18562, N18267);
buf BUF1 (N18564, N18538);
and AND2 (N18565, N18555, N14038);
or OR4 (N18566, N18539, N14884, N2524, N17066);
or OR4 (N18567, N18563, N3006, N5127, N10235);
xor XOR2 (N18568, N18567, N6907);
xor XOR2 (N18569, N18558, N4609);
nor NOR3 (N18570, N18568, N12960, N1141);
buf BUF1 (N18571, N18561);
nand NAND4 (N18572, N18571, N4407, N12111, N4405);
xor XOR2 (N18573, N18565, N13749);
not NOT1 (N18574, N18564);
and AND3 (N18575, N18552, N16911, N18335);
nor NOR3 (N18576, N18574, N15289, N12214);
not NOT1 (N18577, N18569);
and AND4 (N18578, N18566, N3038, N13404, N18174);
buf BUF1 (N18579, N18570);
or OR2 (N18580, N18572, N16546);
nand NAND3 (N18581, N18579, N2649, N2447);
buf BUF1 (N18582, N18573);
and AND3 (N18583, N18577, N4446, N9045);
and AND4 (N18584, N18582, N14548, N3747, N6239);
buf BUF1 (N18585, N18509);
nor NOR3 (N18586, N18585, N7723, N12667);
nand NAND3 (N18587, N18583, N4966, N15621);
or OR3 (N18588, N18556, N8092, N7183);
xor XOR2 (N18589, N18557, N18046);
xor XOR2 (N18590, N18584, N319);
buf BUF1 (N18591, N18580);
not NOT1 (N18592, N18581);
not NOT1 (N18593, N18586);
xor XOR2 (N18594, N18593, N8285);
nand NAND2 (N18595, N18590, N18238);
nor NOR2 (N18596, N18595, N1590);
and AND2 (N18597, N18592, N3298);
xor XOR2 (N18598, N18576, N2746);
not NOT1 (N18599, N18587);
and AND3 (N18600, N18598, N5595, N4657);
buf BUF1 (N18601, N18600);
xor XOR2 (N18602, N18597, N26);
and AND3 (N18603, N18602, N17718, N3510);
xor XOR2 (N18604, N18575, N9179);
xor XOR2 (N18605, N18603, N17555);
buf BUF1 (N18606, N18591);
and AND4 (N18607, N18604, N14196, N10137, N4312);
nand NAND4 (N18608, N18596, N2786, N7301, N14816);
or OR2 (N18609, N18607, N2184);
not NOT1 (N18610, N18606);
or OR2 (N18611, N18601, N11538);
or OR2 (N18612, N18578, N16631);
nand NAND2 (N18613, N18599, N15711);
buf BUF1 (N18614, N18594);
or OR2 (N18615, N18613, N8759);
or OR2 (N18616, N18612, N10507);
xor XOR2 (N18617, N18609, N7962);
buf BUF1 (N18618, N18605);
and AND2 (N18619, N18589, N932);
buf BUF1 (N18620, N18617);
nand NAND4 (N18621, N18608, N18127, N13794, N258);
xor XOR2 (N18622, N18616, N5992);
and AND2 (N18623, N18618, N12760);
not NOT1 (N18624, N18615);
buf BUF1 (N18625, N18588);
not NOT1 (N18626, N18623);
nand NAND2 (N18627, N18626, N4011);
xor XOR2 (N18628, N18610, N11398);
nor NOR4 (N18629, N18621, N12090, N5921, N12793);
buf BUF1 (N18630, N18628);
and AND3 (N18631, N18611, N3741, N18489);
nor NOR4 (N18632, N18631, N16656, N6382, N2964);
nor NOR2 (N18633, N18630, N3161);
nor NOR2 (N18634, N18632, N3928);
not NOT1 (N18635, N18619);
xor XOR2 (N18636, N18622, N4993);
buf BUF1 (N18637, N18624);
nand NAND3 (N18638, N18625, N16440, N140);
and AND4 (N18639, N18636, N13970, N13054, N1508);
not NOT1 (N18640, N18634);
nor NOR3 (N18641, N18639, N18409, N12295);
buf BUF1 (N18642, N18637);
nand NAND3 (N18643, N18640, N16817, N4530);
xor XOR2 (N18644, N18620, N12882);
not NOT1 (N18645, N18644);
not NOT1 (N18646, N18635);
xor XOR2 (N18647, N18642, N9414);
xor XOR2 (N18648, N18643, N8284);
nand NAND3 (N18649, N18633, N10505, N8688);
or OR2 (N18650, N18649, N4456);
not NOT1 (N18651, N18648);
not NOT1 (N18652, N18645);
buf BUF1 (N18653, N18638);
xor XOR2 (N18654, N18646, N3541);
and AND2 (N18655, N18647, N17043);
xor XOR2 (N18656, N18629, N4721);
and AND4 (N18657, N18627, N16302, N6684, N4379);
and AND2 (N18658, N18655, N8705);
or OR4 (N18659, N18641, N16652, N4308, N3589);
and AND4 (N18660, N18651, N11897, N7233, N16317);
and AND2 (N18661, N18659, N13223);
buf BUF1 (N18662, N18654);
buf BUF1 (N18663, N18650);
or OR2 (N18664, N18661, N8064);
nor NOR4 (N18665, N18662, N8121, N16409, N14772);
or OR2 (N18666, N18614, N12605);
or OR4 (N18667, N18653, N1160, N5839, N5076);
not NOT1 (N18668, N18656);
nand NAND2 (N18669, N18658, N12297);
not NOT1 (N18670, N18652);
not NOT1 (N18671, N18657);
nand NAND2 (N18672, N18668, N18220);
buf BUF1 (N18673, N18670);
not NOT1 (N18674, N18665);
not NOT1 (N18675, N18660);
and AND2 (N18676, N18671, N8868);
nor NOR2 (N18677, N18663, N4042);
and AND3 (N18678, N18675, N10938, N17761);
not NOT1 (N18679, N18667);
buf BUF1 (N18680, N18664);
and AND3 (N18681, N18669, N3893, N16151);
nor NOR3 (N18682, N18680, N14940, N3931);
not NOT1 (N18683, N18673);
and AND3 (N18684, N18679, N12019, N7491);
nor NOR4 (N18685, N18678, N2915, N12357, N5799);
not NOT1 (N18686, N18685);
xor XOR2 (N18687, N18681, N1567);
and AND3 (N18688, N18683, N220, N11375);
buf BUF1 (N18689, N18686);
and AND3 (N18690, N18687, N9210, N9005);
or OR3 (N18691, N18684, N15417, N4081);
not NOT1 (N18692, N18677);
and AND4 (N18693, N18691, N17619, N130, N14463);
nand NAND4 (N18694, N18672, N1604, N17131, N5656);
and AND4 (N18695, N18693, N11, N3563, N16889);
or OR4 (N18696, N18674, N3950, N17844, N8991);
nor NOR3 (N18697, N18688, N15841, N9450);
and AND4 (N18698, N18695, N14640, N10251, N10933);
nor NOR3 (N18699, N18696, N9971, N1266);
not NOT1 (N18700, N18666);
not NOT1 (N18701, N18697);
xor XOR2 (N18702, N18699, N9099);
or OR2 (N18703, N18700, N18582);
xor XOR2 (N18704, N18703, N12970);
or OR3 (N18705, N18701, N17187, N15079);
nand NAND4 (N18706, N18690, N12752, N14479, N17963);
or OR4 (N18707, N18706, N17125, N12137, N15344);
nand NAND2 (N18708, N18705, N3050);
nand NAND2 (N18709, N18682, N15362);
and AND2 (N18710, N18689, N1474);
and AND3 (N18711, N18704, N13347, N8479);
not NOT1 (N18712, N18708);
xor XOR2 (N18713, N18676, N12817);
or OR2 (N18714, N18712, N8824);
and AND3 (N18715, N18709, N17221, N16213);
buf BUF1 (N18716, N18694);
nand NAND3 (N18717, N18702, N610, N15478);
not NOT1 (N18718, N18713);
buf BUF1 (N18719, N18714);
nand NAND4 (N18720, N18707, N17447, N2432, N17530);
and AND3 (N18721, N18711, N16066, N498);
or OR3 (N18722, N18710, N5774, N2387);
buf BUF1 (N18723, N18721);
xor XOR2 (N18724, N18719, N11151);
nand NAND2 (N18725, N18720, N9626);
xor XOR2 (N18726, N18725, N2166);
buf BUF1 (N18727, N18698);
and AND4 (N18728, N18724, N9700, N11672, N10289);
or OR3 (N18729, N18718, N15487, N14984);
nor NOR2 (N18730, N18715, N6510);
buf BUF1 (N18731, N18722);
xor XOR2 (N18732, N18692, N7911);
nand NAND2 (N18733, N18723, N2678);
not NOT1 (N18734, N18733);
buf BUF1 (N18735, N18727);
not NOT1 (N18736, N18729);
buf BUF1 (N18737, N18735);
xor XOR2 (N18738, N18716, N11761);
nand NAND2 (N18739, N18717, N17127);
nand NAND2 (N18740, N18731, N12266);
xor XOR2 (N18741, N18739, N15856);
not NOT1 (N18742, N18732);
not NOT1 (N18743, N18736);
or OR4 (N18744, N18738, N13962, N13232, N14791);
nand NAND3 (N18745, N18726, N17309, N11882);
nand NAND2 (N18746, N18730, N8508);
xor XOR2 (N18747, N18737, N13970);
and AND4 (N18748, N18744, N15347, N698, N9710);
xor XOR2 (N18749, N18728, N13865);
not NOT1 (N18750, N18743);
xor XOR2 (N18751, N18746, N6235);
buf BUF1 (N18752, N18747);
not NOT1 (N18753, N18734);
nor NOR4 (N18754, N18750, N16626, N4484, N10570);
and AND3 (N18755, N18753, N4004, N9655);
xor XOR2 (N18756, N18741, N343);
or OR2 (N18757, N18740, N5578);
nand NAND3 (N18758, N18757, N1368, N12231);
not NOT1 (N18759, N18755);
not NOT1 (N18760, N18758);
nor NOR3 (N18761, N18760, N2255, N2613);
or OR2 (N18762, N18761, N11288);
nor NOR2 (N18763, N18742, N12248);
and AND2 (N18764, N18749, N6551);
and AND2 (N18765, N18762, N8393);
nand NAND4 (N18766, N18752, N12155, N12364, N8337);
or OR3 (N18767, N18751, N4474, N15066);
nand NAND2 (N18768, N18765, N13494);
nor NOR2 (N18769, N18754, N12844);
xor XOR2 (N18770, N18756, N17277);
buf BUF1 (N18771, N18768);
or OR3 (N18772, N18748, N12900, N15546);
nor NOR2 (N18773, N18770, N5864);
buf BUF1 (N18774, N18771);
and AND2 (N18775, N18774, N15088);
nor NOR4 (N18776, N18766, N6948, N7920, N14967);
and AND2 (N18777, N18759, N16737);
nor NOR3 (N18778, N18767, N10370, N14917);
nand NAND4 (N18779, N18778, N13121, N15734, N15015);
nand NAND4 (N18780, N18769, N4791, N11290, N7363);
and AND4 (N18781, N18779, N13446, N14131, N3697);
buf BUF1 (N18782, N18764);
not NOT1 (N18783, N18763);
buf BUF1 (N18784, N18772);
or OR3 (N18785, N18777, N8876, N10862);
buf BUF1 (N18786, N18785);
or OR2 (N18787, N18784, N5457);
not NOT1 (N18788, N18781);
nor NOR2 (N18789, N18773, N15664);
not NOT1 (N18790, N18776);
nand NAND4 (N18791, N18787, N18653, N10421, N16842);
nor NOR2 (N18792, N18775, N7018);
or OR4 (N18793, N18786, N14145, N1290, N7418);
xor XOR2 (N18794, N18780, N17805);
nor NOR4 (N18795, N18782, N3622, N10078, N811);
or OR3 (N18796, N18793, N10227, N6687);
and AND4 (N18797, N18795, N14841, N4084, N8083);
nand NAND3 (N18798, N18797, N10126, N9246);
buf BUF1 (N18799, N18798);
nand NAND3 (N18800, N18788, N734, N17695);
nor NOR2 (N18801, N18783, N10095);
buf BUF1 (N18802, N18790);
xor XOR2 (N18803, N18800, N3053);
and AND3 (N18804, N18803, N14541, N8669);
not NOT1 (N18805, N18802);
xor XOR2 (N18806, N18804, N2996);
nand NAND2 (N18807, N18796, N8987);
nor NOR4 (N18808, N18789, N2669, N9239, N15681);
not NOT1 (N18809, N18801);
nor NOR3 (N18810, N18808, N9249, N12854);
nand NAND3 (N18811, N18745, N18784, N2949);
or OR3 (N18812, N18807, N8531, N14126);
xor XOR2 (N18813, N18791, N16206);
xor XOR2 (N18814, N18811, N391);
nor NOR4 (N18815, N18806, N140, N1423, N13383);
or OR3 (N18816, N18799, N3673, N5269);
and AND2 (N18817, N18812, N3895);
nand NAND3 (N18818, N18816, N2519, N17124);
nor NOR4 (N18819, N18805, N16876, N14031, N13016);
and AND4 (N18820, N18794, N6519, N14713, N12455);
nand NAND2 (N18821, N18792, N3807);
or OR4 (N18822, N18815, N2877, N14468, N10762);
not NOT1 (N18823, N18818);
and AND2 (N18824, N18813, N12717);
xor XOR2 (N18825, N18810, N10383);
xor XOR2 (N18826, N18821, N14476);
buf BUF1 (N18827, N18817);
and AND4 (N18828, N18823, N13726, N14286, N7940);
nor NOR4 (N18829, N18819, N13119, N11833, N10067);
xor XOR2 (N18830, N18824, N654);
or OR3 (N18831, N18820, N5211, N1812);
and AND4 (N18832, N18830, N11913, N6162, N3219);
not NOT1 (N18833, N18831);
xor XOR2 (N18834, N18833, N9761);
nand NAND3 (N18835, N18822, N9187, N6656);
xor XOR2 (N18836, N18809, N18468);
nor NOR4 (N18837, N18832, N15115, N13752, N11513);
nor NOR2 (N18838, N18836, N7674);
not NOT1 (N18839, N18837);
nor NOR4 (N18840, N18814, N3929, N13445, N15432);
and AND2 (N18841, N18825, N948);
nand NAND3 (N18842, N18841, N5206, N6363);
buf BUF1 (N18843, N18839);
xor XOR2 (N18844, N18843, N7764);
xor XOR2 (N18845, N18829, N8079);
xor XOR2 (N18846, N18827, N6010);
xor XOR2 (N18847, N18842, N5618);
or OR4 (N18848, N18845, N15243, N18513, N7881);
and AND2 (N18849, N18840, N6439);
and AND4 (N18850, N18847, N13263, N3692, N7277);
nand NAND4 (N18851, N18848, N7515, N16021, N10397);
not NOT1 (N18852, N18835);
nor NOR4 (N18853, N18826, N2212, N1970, N2955);
xor XOR2 (N18854, N18834, N8417);
nor NOR2 (N18855, N18853, N7972);
xor XOR2 (N18856, N18846, N12036);
buf BUF1 (N18857, N18855);
and AND4 (N18858, N18844, N12191, N1026, N13457);
not NOT1 (N18859, N18857);
buf BUF1 (N18860, N18828);
and AND2 (N18861, N18852, N3607);
and AND2 (N18862, N18860, N16958);
nand NAND3 (N18863, N18859, N12523, N8751);
nor NOR4 (N18864, N18856, N15934, N14174, N11033);
buf BUF1 (N18865, N18850);
nor NOR3 (N18866, N18849, N15195, N6082);
nor NOR4 (N18867, N18861, N2340, N4749, N13746);
and AND3 (N18868, N18864, N16322, N4308);
not NOT1 (N18869, N18863);
xor XOR2 (N18870, N18868, N6251);
or OR4 (N18871, N18870, N11538, N15524, N15308);
and AND2 (N18872, N18854, N7943);
not NOT1 (N18873, N18851);
xor XOR2 (N18874, N18869, N11066);
not NOT1 (N18875, N18858);
and AND3 (N18876, N18871, N9354, N8218);
buf BUF1 (N18877, N18874);
and AND4 (N18878, N18867, N16544, N11307, N14224);
nor NOR2 (N18879, N18873, N14869);
or OR3 (N18880, N18875, N1253, N17281);
not NOT1 (N18881, N18880);
nor NOR4 (N18882, N18877, N1242, N4300, N14487);
xor XOR2 (N18883, N18838, N14491);
and AND2 (N18884, N18865, N8163);
nor NOR4 (N18885, N18876, N11221, N3792, N18718);
buf BUF1 (N18886, N18878);
buf BUF1 (N18887, N18872);
not NOT1 (N18888, N18862);
nand NAND2 (N18889, N18883, N405);
buf BUF1 (N18890, N18888);
nand NAND2 (N18891, N18884, N4764);
nand NAND2 (N18892, N18866, N1310);
nor NOR4 (N18893, N18881, N9618, N17385, N8412);
or OR4 (N18894, N18885, N17724, N2948, N9862);
nor NOR4 (N18895, N18894, N14066, N3743, N6333);
not NOT1 (N18896, N18887);
or OR2 (N18897, N18891, N18890);
nand NAND2 (N18898, N12540, N3909);
xor XOR2 (N18899, N18886, N16162);
and AND2 (N18900, N18892, N9476);
and AND2 (N18901, N18897, N17616);
nor NOR3 (N18902, N18889, N2433, N1577);
xor XOR2 (N18903, N18901, N15258);
buf BUF1 (N18904, N18898);
not NOT1 (N18905, N18882);
xor XOR2 (N18906, N18903, N1739);
nand NAND2 (N18907, N18902, N1953);
xor XOR2 (N18908, N18893, N18183);
or OR3 (N18909, N18908, N15311, N4845);
and AND2 (N18910, N18905, N7301);
and AND4 (N18911, N18904, N4547, N12848, N5230);
nand NAND3 (N18912, N18899, N1183, N8002);
or OR2 (N18913, N18911, N273);
nand NAND2 (N18914, N18912, N438);
not NOT1 (N18915, N18913);
and AND4 (N18916, N18909, N18011, N16662, N4230);
or OR4 (N18917, N18907, N5215, N15753, N15405);
buf BUF1 (N18918, N18917);
buf BUF1 (N18919, N18896);
nor NOR4 (N18920, N18916, N8696, N9124, N92);
or OR4 (N18921, N18914, N4433, N6652, N11674);
nor NOR2 (N18922, N18900, N1502);
xor XOR2 (N18923, N18919, N11470);
and AND2 (N18924, N18915, N12099);
not NOT1 (N18925, N18924);
buf BUF1 (N18926, N18895);
nand NAND2 (N18927, N18925, N11470);
xor XOR2 (N18928, N18920, N2154);
nand NAND3 (N18929, N18926, N1200, N8087);
or OR3 (N18930, N18918, N6266, N7982);
xor XOR2 (N18931, N18927, N17540);
nor NOR4 (N18932, N18923, N2831, N6787, N15581);
and AND3 (N18933, N18921, N12996, N18822);
not NOT1 (N18934, N18929);
nor NOR3 (N18935, N18910, N10790, N10967);
buf BUF1 (N18936, N18932);
buf BUF1 (N18937, N18928);
and AND3 (N18938, N18933, N7496, N13801);
nand NAND2 (N18939, N18906, N3131);
or OR2 (N18940, N18922, N1671);
nand NAND3 (N18941, N18936, N10819, N5851);
nand NAND4 (N18942, N18938, N5361, N1819, N3577);
nor NOR4 (N18943, N18937, N689, N2327, N9632);
or OR4 (N18944, N18939, N12710, N18655, N15678);
buf BUF1 (N18945, N18940);
nand NAND2 (N18946, N18941, N9789);
xor XOR2 (N18947, N18942, N4880);
buf BUF1 (N18948, N18931);
buf BUF1 (N18949, N18943);
xor XOR2 (N18950, N18935, N456);
not NOT1 (N18951, N18879);
and AND2 (N18952, N18945, N1096);
nand NAND2 (N18953, N18944, N10184);
buf BUF1 (N18954, N18953);
buf BUF1 (N18955, N18950);
nor NOR2 (N18956, N18947, N11609);
nor NOR4 (N18957, N18956, N9084, N6941, N18690);
and AND3 (N18958, N18951, N4677, N3059);
not NOT1 (N18959, N18957);
and AND3 (N18960, N18934, N2465, N2962);
or OR4 (N18961, N18960, N902, N1173, N6440);
and AND3 (N18962, N18948, N5548, N16042);
or OR4 (N18963, N18949, N16759, N11347, N13516);
or OR3 (N18964, N18958, N8733, N8104);
buf BUF1 (N18965, N18946);
or OR2 (N18966, N18952, N12106);
xor XOR2 (N18967, N18959, N17659);
buf BUF1 (N18968, N18961);
not NOT1 (N18969, N18968);
nor NOR3 (N18970, N18930, N9795, N15117);
and AND2 (N18971, N18970, N10888);
or OR2 (N18972, N18962, N15580);
xor XOR2 (N18973, N18955, N16035);
not NOT1 (N18974, N18967);
buf BUF1 (N18975, N18973);
not NOT1 (N18976, N18964);
or OR3 (N18977, N18971, N18600, N8948);
buf BUF1 (N18978, N18963);
nor NOR3 (N18979, N18972, N5742, N10214);
buf BUF1 (N18980, N18977);
not NOT1 (N18981, N18965);
or OR2 (N18982, N18980, N6032);
nand NAND4 (N18983, N18978, N15648, N3762, N13830);
and AND2 (N18984, N18974, N10592);
or OR3 (N18985, N18982, N6833, N6577);
not NOT1 (N18986, N18976);
nor NOR4 (N18987, N18985, N13126, N13836, N2293);
xor XOR2 (N18988, N18969, N85);
xor XOR2 (N18989, N18954, N8852);
or OR3 (N18990, N18984, N515, N17363);
or OR4 (N18991, N18989, N4620, N14744, N15382);
buf BUF1 (N18992, N18990);
xor XOR2 (N18993, N18987, N9153);
not NOT1 (N18994, N18988);
and AND2 (N18995, N18979, N7481);
xor XOR2 (N18996, N18992, N352);
or OR2 (N18997, N18966, N18097);
nand NAND4 (N18998, N18994, N15557, N3636, N11325);
xor XOR2 (N18999, N18991, N8270);
not NOT1 (N19000, N18998);
xor XOR2 (N19001, N18986, N6208);
buf BUF1 (N19002, N18996);
xor XOR2 (N19003, N18997, N7489);
xor XOR2 (N19004, N18983, N4368);
or OR4 (N19005, N19000, N7779, N5317, N16943);
nand NAND2 (N19006, N18981, N11265);
nand NAND3 (N19007, N18993, N3783, N13575);
not NOT1 (N19008, N18995);
and AND3 (N19009, N19002, N3525, N3104);
xor XOR2 (N19010, N19004, N14962);
xor XOR2 (N19011, N19003, N14014);
not NOT1 (N19012, N19001);
or OR3 (N19013, N18975, N10578, N12001);
or OR3 (N19014, N19013, N11452, N9275);
nor NOR2 (N19015, N19011, N15185);
nor NOR4 (N19016, N19009, N1878, N13337, N2100);
or OR4 (N19017, N19006, N12165, N11952, N6500);
buf BUF1 (N19018, N19010);
and AND3 (N19019, N19008, N2221, N5739);
or OR3 (N19020, N19019, N4543, N17752);
buf BUF1 (N19021, N19017);
nor NOR4 (N19022, N19018, N14433, N7679, N18955);
xor XOR2 (N19023, N19012, N11440);
nand NAND4 (N19024, N19014, N7848, N14072, N16470);
and AND3 (N19025, N19007, N11546, N1953);
nand NAND4 (N19026, N19025, N9605, N6503, N5262);
or OR3 (N19027, N19005, N2533, N17877);
nand NAND3 (N19028, N19027, N11564, N108);
buf BUF1 (N19029, N19015);
xor XOR2 (N19030, N19016, N683);
and AND3 (N19031, N19021, N12613, N18534);
and AND4 (N19032, N19020, N13046, N15472, N13460);
buf BUF1 (N19033, N19022);
or OR4 (N19034, N19024, N16273, N12236, N11888);
nand NAND2 (N19035, N19033, N96);
or OR2 (N19036, N19034, N15447);
nor NOR4 (N19037, N19023, N3015, N4246, N10248);
and AND4 (N19038, N19032, N18059, N3929, N8044);
xor XOR2 (N19039, N19037, N7412);
not NOT1 (N19040, N19031);
nand NAND4 (N19041, N19036, N18871, N7009, N13218);
nor NOR3 (N19042, N19041, N11580, N15307);
not NOT1 (N19043, N19028);
and AND4 (N19044, N19026, N7794, N5906, N2343);
not NOT1 (N19045, N18999);
buf BUF1 (N19046, N19038);
xor XOR2 (N19047, N19043, N16324);
not NOT1 (N19048, N19030);
buf BUF1 (N19049, N19045);
and AND4 (N19050, N19049, N1320, N3036, N8178);
or OR2 (N19051, N19029, N15035);
and AND2 (N19052, N19050, N13757);
nor NOR2 (N19053, N19051, N9247);
nor NOR2 (N19054, N19044, N14141);
buf BUF1 (N19055, N19035);
nand NAND4 (N19056, N19055, N11715, N530, N10081);
or OR2 (N19057, N19046, N12068);
and AND2 (N19058, N19040, N8740);
or OR3 (N19059, N19058, N2390, N1911);
and AND2 (N19060, N19042, N6685);
nor NOR2 (N19061, N19057, N18874);
nor NOR4 (N19062, N19052, N2756, N6348, N17631);
buf BUF1 (N19063, N19059);
or OR4 (N19064, N19060, N18194, N10390, N6836);
buf BUF1 (N19065, N19054);
xor XOR2 (N19066, N19039, N6192);
xor XOR2 (N19067, N19063, N3777);
and AND4 (N19068, N19056, N11327, N12246, N6500);
buf BUF1 (N19069, N19068);
and AND3 (N19070, N19048, N5030, N11284);
and AND2 (N19071, N19047, N10868);
nor NOR3 (N19072, N19070, N11361, N9287);
and AND4 (N19073, N19071, N3308, N6949, N6571);
not NOT1 (N19074, N19064);
or OR3 (N19075, N19065, N10174, N11906);
not NOT1 (N19076, N19053);
not NOT1 (N19077, N19076);
and AND4 (N19078, N19062, N16926, N6933, N15632);
not NOT1 (N19079, N19072);
not NOT1 (N19080, N19067);
nor NOR3 (N19081, N19069, N14338, N2745);
buf BUF1 (N19082, N19073);
and AND3 (N19083, N19080, N18807, N16332);
and AND4 (N19084, N19066, N10412, N2437, N2458);
xor XOR2 (N19085, N19074, N7977);
nor NOR2 (N19086, N19082, N17913);
nor NOR2 (N19087, N19085, N7033);
and AND4 (N19088, N19075, N9009, N18197, N18042);
buf BUF1 (N19089, N19077);
xor XOR2 (N19090, N19084, N14854);
nand NAND3 (N19091, N19081, N12493, N6531);
and AND3 (N19092, N19079, N462, N16307);
not NOT1 (N19093, N19086);
nand NAND2 (N19094, N19091, N16300);
or OR2 (N19095, N19061, N3999);
xor XOR2 (N19096, N19083, N10161);
buf BUF1 (N19097, N19089);
or OR4 (N19098, N19088, N10528, N16960, N18983);
not NOT1 (N19099, N19096);
not NOT1 (N19100, N19087);
xor XOR2 (N19101, N19090, N15315);
not NOT1 (N19102, N19101);
or OR3 (N19103, N19093, N14755, N17086);
or OR4 (N19104, N19094, N10316, N13147, N14902);
or OR3 (N19105, N19102, N16638, N15817);
and AND4 (N19106, N19095, N12764, N9367, N13551);
or OR2 (N19107, N19078, N786);
buf BUF1 (N19108, N19104);
nor NOR3 (N19109, N19092, N16666, N9194);
not NOT1 (N19110, N19107);
nand NAND3 (N19111, N19103, N2898, N18138);
buf BUF1 (N19112, N19099);
not NOT1 (N19113, N19112);
or OR4 (N19114, N19105, N17837, N12425, N1853);
nor NOR3 (N19115, N19100, N12356, N5913);
or OR3 (N19116, N19111, N6210, N17068);
and AND3 (N19117, N19116, N4017, N78);
xor XOR2 (N19118, N19106, N4252);
not NOT1 (N19119, N19109);
buf BUF1 (N19120, N19118);
not NOT1 (N19121, N19110);
nand NAND2 (N19122, N19119, N6380);
nand NAND4 (N19123, N19121, N9611, N2794, N16141);
or OR4 (N19124, N19120, N7947, N3261, N15352);
and AND2 (N19125, N19114, N13687);
or OR3 (N19126, N19124, N11415, N1415);
nor NOR2 (N19127, N19126, N13320);
buf BUF1 (N19128, N19115);
nor NOR2 (N19129, N19127, N63);
nand NAND2 (N19130, N19113, N11389);
nand NAND2 (N19131, N19129, N12781);
and AND2 (N19132, N19128, N9772);
nor NOR4 (N19133, N19132, N14018, N17060, N10602);
or OR4 (N19134, N19117, N4013, N17613, N3302);
and AND3 (N19135, N19131, N11788, N8148);
not NOT1 (N19136, N19098);
and AND4 (N19137, N19135, N10660, N2539, N2461);
xor XOR2 (N19138, N19137, N11802);
and AND2 (N19139, N19138, N18209);
nand NAND2 (N19140, N19139, N13820);
not NOT1 (N19141, N19122);
buf BUF1 (N19142, N19108);
not NOT1 (N19143, N19133);
nor NOR4 (N19144, N19142, N15242, N19124, N8372);
nor NOR3 (N19145, N19140, N11825, N14434);
or OR2 (N19146, N19123, N4889);
nor NOR4 (N19147, N19145, N14319, N3570, N2228);
or OR2 (N19148, N19147, N11934);
xor XOR2 (N19149, N19148, N13332);
and AND3 (N19150, N19130, N11025, N15678);
buf BUF1 (N19151, N19149);
buf BUF1 (N19152, N19151);
and AND2 (N19153, N19144, N1806);
and AND3 (N19154, N19146, N9439, N6953);
and AND2 (N19155, N19125, N7635);
or OR3 (N19156, N19152, N6259, N56);
and AND2 (N19157, N19097, N12755);
nand NAND3 (N19158, N19153, N17293, N14775);
or OR4 (N19159, N19158, N14749, N8229, N7408);
buf BUF1 (N19160, N19143);
nand NAND4 (N19161, N19136, N1199, N7258, N7503);
not NOT1 (N19162, N19134);
buf BUF1 (N19163, N19161);
or OR2 (N19164, N19154, N1516);
nand NAND3 (N19165, N19157, N14470, N875);
nor NOR4 (N19166, N19160, N19109, N9071, N8055);
buf BUF1 (N19167, N19163);
nand NAND4 (N19168, N19165, N15121, N2337, N16277);
not NOT1 (N19169, N19167);
buf BUF1 (N19170, N19164);
and AND4 (N19171, N19162, N12318, N3255, N2352);
nand NAND4 (N19172, N19169, N3150, N875, N3561);
xor XOR2 (N19173, N19156, N9076);
nor NOR3 (N19174, N19173, N16373, N17281);
and AND3 (N19175, N19171, N502, N13960);
and AND4 (N19176, N19159, N3114, N16695, N9023);
and AND2 (N19177, N19176, N1831);
buf BUF1 (N19178, N19141);
nor NOR4 (N19179, N19170, N19, N17303, N7046);
xor XOR2 (N19180, N19150, N2379);
buf BUF1 (N19181, N19174);
nor NOR2 (N19182, N19179, N8952);
and AND2 (N19183, N19182, N6392);
not NOT1 (N19184, N19178);
nor NOR2 (N19185, N19177, N5120);
not NOT1 (N19186, N19166);
or OR2 (N19187, N19181, N4695);
not NOT1 (N19188, N19175);
buf BUF1 (N19189, N19168);
not NOT1 (N19190, N19186);
nor NOR3 (N19191, N19190, N18559, N15065);
xor XOR2 (N19192, N19184, N12501);
xor XOR2 (N19193, N19155, N4351);
xor XOR2 (N19194, N19191, N14059);
and AND3 (N19195, N19183, N15365, N6837);
not NOT1 (N19196, N19194);
or OR4 (N19197, N19188, N3461, N17825, N3613);
or OR3 (N19198, N19195, N11576, N7408);
or OR2 (N19199, N19185, N2834);
or OR3 (N19200, N19192, N786, N6294);
not NOT1 (N19201, N19196);
not NOT1 (N19202, N19200);
nand NAND3 (N19203, N19198, N1580, N6649);
buf BUF1 (N19204, N19202);
nand NAND4 (N19205, N19203, N14853, N7657, N12175);
and AND3 (N19206, N19205, N11081, N11238);
buf BUF1 (N19207, N19180);
buf BUF1 (N19208, N19189);
nor NOR3 (N19209, N19201, N1379, N4005);
nand NAND4 (N19210, N19172, N1335, N16773, N7115);
buf BUF1 (N19211, N19199);
xor XOR2 (N19212, N19193, N8823);
not NOT1 (N19213, N19209);
nor NOR4 (N19214, N19212, N18161, N11227, N16008);
buf BUF1 (N19215, N19207);
or OR4 (N19216, N19204, N10512, N13147, N984);
or OR2 (N19217, N19213, N1314);
and AND4 (N19218, N19206, N17940, N276, N9552);
not NOT1 (N19219, N19210);
not NOT1 (N19220, N19215);
buf BUF1 (N19221, N19216);
nand NAND4 (N19222, N19214, N8047, N8032, N9095);
or OR3 (N19223, N19197, N11121, N12387);
and AND2 (N19224, N19222, N10766);
nand NAND4 (N19225, N19187, N5469, N10334, N13592);
not NOT1 (N19226, N19211);
nor NOR4 (N19227, N19226, N3474, N11658, N15072);
not NOT1 (N19228, N19218);
and AND2 (N19229, N19208, N14865);
xor XOR2 (N19230, N19221, N18874);
buf BUF1 (N19231, N19220);
nor NOR3 (N19232, N19228, N1228, N19035);
buf BUF1 (N19233, N19227);
nand NAND3 (N19234, N19233, N185, N9677);
xor XOR2 (N19235, N19223, N2314);
xor XOR2 (N19236, N19231, N9058);
xor XOR2 (N19237, N19236, N18703);
nor NOR3 (N19238, N19219, N19230, N15779);
nand NAND3 (N19239, N11266, N13127, N2679);
buf BUF1 (N19240, N19234);
nand NAND2 (N19241, N19238, N12245);
xor XOR2 (N19242, N19237, N10918);
and AND3 (N19243, N19239, N19095, N3664);
nor NOR3 (N19244, N19229, N13725, N2059);
nand NAND3 (N19245, N19232, N15806, N6233);
buf BUF1 (N19246, N19244);
nor NOR2 (N19247, N19224, N13495);
or OR2 (N19248, N19246, N16127);
nor NOR2 (N19249, N19217, N8880);
buf BUF1 (N19250, N19242);
buf BUF1 (N19251, N19241);
nand NAND3 (N19252, N19245, N17398, N3052);
or OR4 (N19253, N19251, N2407, N14063, N7118);
buf BUF1 (N19254, N19249);
nor NOR3 (N19255, N19248, N8672, N7599);
buf BUF1 (N19256, N19254);
buf BUF1 (N19257, N19255);
not NOT1 (N19258, N19225);
xor XOR2 (N19259, N19256, N5087);
nand NAND4 (N19260, N19247, N8075, N1603, N13517);
nor NOR4 (N19261, N19240, N15922, N18083, N4756);
and AND2 (N19262, N19250, N12140);
buf BUF1 (N19263, N19243);
nand NAND3 (N19264, N19260, N2667, N4957);
nand NAND3 (N19265, N19235, N10264, N1797);
buf BUF1 (N19266, N19258);
and AND3 (N19267, N19265, N17144, N6276);
xor XOR2 (N19268, N19253, N1812);
xor XOR2 (N19269, N19252, N12792);
not NOT1 (N19270, N19268);
nand NAND2 (N19271, N19270, N4713);
or OR2 (N19272, N19262, N17470);
buf BUF1 (N19273, N19267);
nand NAND4 (N19274, N19271, N14647, N13240, N197);
xor XOR2 (N19275, N19261, N11767);
nor NOR3 (N19276, N19273, N15717, N5057);
not NOT1 (N19277, N19263);
nor NOR4 (N19278, N19272, N17478, N9467, N18865);
and AND4 (N19279, N19278, N10749, N14623, N13888);
not NOT1 (N19280, N19264);
nand NAND2 (N19281, N19257, N15645);
and AND2 (N19282, N19274, N11279);
buf BUF1 (N19283, N19281);
or OR3 (N19284, N19276, N813, N9281);
xor XOR2 (N19285, N19282, N8067);
or OR4 (N19286, N19266, N10936, N16476, N15051);
and AND3 (N19287, N19280, N15099, N5832);
nor NOR4 (N19288, N19259, N15979, N8728, N9470);
and AND4 (N19289, N19288, N12659, N7888, N5399);
or OR3 (N19290, N19275, N5488, N4976);
xor XOR2 (N19291, N19286, N1348);
xor XOR2 (N19292, N19291, N4752);
buf BUF1 (N19293, N19285);
or OR3 (N19294, N19293, N16068, N9885);
nor NOR4 (N19295, N19294, N13404, N1427, N13194);
nand NAND2 (N19296, N19295, N14141);
or OR2 (N19297, N19287, N2701);
nand NAND3 (N19298, N19283, N10314, N13497);
xor XOR2 (N19299, N19284, N18939);
xor XOR2 (N19300, N19292, N16033);
or OR3 (N19301, N19289, N13560, N16276);
nand NAND4 (N19302, N19301, N16882, N560, N10592);
nand NAND3 (N19303, N19269, N4410, N15743);
or OR2 (N19304, N19300, N16318);
nor NOR3 (N19305, N19297, N14422, N4708);
or OR3 (N19306, N19304, N18675, N11450);
nor NOR4 (N19307, N19306, N18327, N4877, N6374);
nor NOR4 (N19308, N19305, N11587, N3291, N9825);
xor XOR2 (N19309, N19308, N1776);
not NOT1 (N19310, N19298);
nor NOR3 (N19311, N19277, N11131, N6371);
not NOT1 (N19312, N19309);
not NOT1 (N19313, N19312);
xor XOR2 (N19314, N19279, N7598);
nor NOR2 (N19315, N19314, N14152);
xor XOR2 (N19316, N19290, N5432);
nor NOR3 (N19317, N19316, N3081, N615);
and AND3 (N19318, N19310, N18941, N228);
or OR4 (N19319, N19313, N17125, N13518, N5173);
buf BUF1 (N19320, N19318);
nor NOR3 (N19321, N19320, N19272, N515);
xor XOR2 (N19322, N19317, N18798);
xor XOR2 (N19323, N19311, N18986);
nor NOR3 (N19324, N19303, N10783, N16493);
nand NAND4 (N19325, N19302, N7266, N10779, N16689);
not NOT1 (N19326, N19307);
nand NAND3 (N19327, N19322, N11638, N16894);
or OR3 (N19328, N19319, N16502, N8341);
buf BUF1 (N19329, N19324);
nor NOR4 (N19330, N19327, N19046, N10053, N16917);
buf BUF1 (N19331, N19330);
buf BUF1 (N19332, N19323);
xor XOR2 (N19333, N19326, N14807);
nor NOR2 (N19334, N19299, N7571);
nand NAND2 (N19335, N19296, N1426);
xor XOR2 (N19336, N19329, N2712);
nor NOR2 (N19337, N19325, N1222);
not NOT1 (N19338, N19335);
nor NOR4 (N19339, N19333, N5257, N12340, N11415);
nand NAND4 (N19340, N19337, N3945, N11603, N8668);
nor NOR2 (N19341, N19332, N6372);
xor XOR2 (N19342, N19315, N16288);
buf BUF1 (N19343, N19331);
xor XOR2 (N19344, N19343, N13403);
xor XOR2 (N19345, N19339, N16341);
nor NOR2 (N19346, N19336, N11221);
nand NAND4 (N19347, N19342, N7680, N15, N12212);
nand NAND2 (N19348, N19346, N13562);
nor NOR3 (N19349, N19340, N15879, N4019);
or OR3 (N19350, N19345, N19313, N3743);
or OR4 (N19351, N19347, N14378, N18289, N16191);
not NOT1 (N19352, N19341);
or OR3 (N19353, N19334, N14436, N17317);
xor XOR2 (N19354, N19328, N14928);
and AND3 (N19355, N19344, N672, N14122);
not NOT1 (N19356, N19355);
nor NOR4 (N19357, N19356, N10136, N12076, N18795);
and AND3 (N19358, N19348, N13448, N9812);
buf BUF1 (N19359, N19358);
buf BUF1 (N19360, N19359);
buf BUF1 (N19361, N19338);
and AND3 (N19362, N19357, N19146, N18419);
and AND4 (N19363, N19321, N18130, N8881, N1902);
and AND2 (N19364, N19352, N12535);
xor XOR2 (N19365, N19349, N2814);
or OR2 (N19366, N19351, N18252);
and AND4 (N19367, N19361, N7201, N2066, N4034);
nand NAND2 (N19368, N19367, N11707);
or OR4 (N19369, N19368, N6150, N344, N6003);
xor XOR2 (N19370, N19350, N18016);
not NOT1 (N19371, N19360);
xor XOR2 (N19372, N19369, N2325);
nand NAND3 (N19373, N19362, N12941, N12630);
nor NOR4 (N19374, N19365, N14042, N17527, N13960);
nor NOR2 (N19375, N19354, N3562);
not NOT1 (N19376, N19353);
xor XOR2 (N19377, N19364, N1777);
and AND2 (N19378, N19366, N17726);
or OR3 (N19379, N19373, N14185, N5695);
and AND3 (N19380, N19378, N17236, N2079);
or OR4 (N19381, N19371, N15794, N5306, N6496);
or OR3 (N19382, N19376, N16808, N8326);
and AND3 (N19383, N19374, N18642, N9469);
and AND3 (N19384, N19363, N16623, N12177);
and AND4 (N19385, N19375, N7470, N13239, N6872);
buf BUF1 (N19386, N19384);
not NOT1 (N19387, N19385);
buf BUF1 (N19388, N19372);
and AND3 (N19389, N19370, N6734, N8732);
or OR3 (N19390, N19377, N18958, N19195);
not NOT1 (N19391, N19386);
or OR3 (N19392, N19381, N16389, N483);
xor XOR2 (N19393, N19392, N3746);
buf BUF1 (N19394, N19383);
nor NOR3 (N19395, N19382, N9326, N15868);
not NOT1 (N19396, N19389);
buf BUF1 (N19397, N19393);
xor XOR2 (N19398, N19391, N10114);
or OR3 (N19399, N19380, N16214, N17071);
xor XOR2 (N19400, N19398, N6326);
nor NOR3 (N19401, N19396, N13826, N17133);
not NOT1 (N19402, N19397);
nand NAND2 (N19403, N19387, N8651);
nand NAND2 (N19404, N19394, N8249);
buf BUF1 (N19405, N19399);
nand NAND2 (N19406, N19401, N9435);
xor XOR2 (N19407, N19388, N1737);
nor NOR4 (N19408, N19404, N5159, N11164, N15623);
xor XOR2 (N19409, N19405, N4744);
buf BUF1 (N19410, N19395);
buf BUF1 (N19411, N19406);
not NOT1 (N19412, N19379);
not NOT1 (N19413, N19403);
nand NAND2 (N19414, N19411, N16377);
xor XOR2 (N19415, N19414, N15367);
xor XOR2 (N19416, N19410, N13549);
buf BUF1 (N19417, N19415);
xor XOR2 (N19418, N19408, N14585);
not NOT1 (N19419, N19413);
and AND4 (N19420, N19402, N11990, N5984, N1132);
xor XOR2 (N19421, N19419, N16411);
or OR2 (N19422, N19407, N15989);
xor XOR2 (N19423, N19417, N9493);
buf BUF1 (N19424, N19416);
xor XOR2 (N19425, N19423, N15493);
and AND2 (N19426, N19400, N8423);
nor NOR2 (N19427, N19426, N6940);
not NOT1 (N19428, N19418);
nand NAND4 (N19429, N19409, N6515, N15585, N8434);
and AND2 (N19430, N19427, N11652);
buf BUF1 (N19431, N19421);
not NOT1 (N19432, N19390);
buf BUF1 (N19433, N19429);
or OR4 (N19434, N19431, N253, N7591, N4629);
and AND3 (N19435, N19425, N17401, N5127);
xor XOR2 (N19436, N19420, N19263);
not NOT1 (N19437, N19432);
buf BUF1 (N19438, N19435);
and AND3 (N19439, N19422, N18021, N17428);
not NOT1 (N19440, N19433);
and AND2 (N19441, N19436, N3520);
not NOT1 (N19442, N19440);
nand NAND2 (N19443, N19434, N15297);
not NOT1 (N19444, N19424);
and AND3 (N19445, N19442, N15268, N13163);
or OR4 (N19446, N19437, N18493, N18962, N10629);
buf BUF1 (N19447, N19438);
xor XOR2 (N19448, N19447, N15440);
nor NOR2 (N19449, N19441, N650);
nor NOR3 (N19450, N19412, N18801, N7021);
and AND3 (N19451, N19428, N17107, N6236);
not NOT1 (N19452, N19451);
xor XOR2 (N19453, N19448, N2568);
not NOT1 (N19454, N19453);
nand NAND3 (N19455, N19443, N7795, N17464);
xor XOR2 (N19456, N19446, N17384);
nand NAND3 (N19457, N19454, N16212, N12687);
and AND4 (N19458, N19449, N16771, N11753, N17472);
xor XOR2 (N19459, N19457, N2123);
or OR3 (N19460, N19455, N15384, N9971);
nor NOR3 (N19461, N19458, N9476, N531);
nor NOR4 (N19462, N19444, N5764, N2878, N2412);
nor NOR3 (N19463, N19452, N3789, N8845);
buf BUF1 (N19464, N19461);
not NOT1 (N19465, N19460);
and AND2 (N19466, N19439, N7801);
nand NAND2 (N19467, N19466, N13377);
not NOT1 (N19468, N19445);
not NOT1 (N19469, N19456);
nand NAND3 (N19470, N19430, N8512, N17029);
or OR3 (N19471, N19467, N10288, N15121);
buf BUF1 (N19472, N19469);
buf BUF1 (N19473, N19450);
or OR2 (N19474, N19462, N17379);
xor XOR2 (N19475, N19459, N5235);
and AND3 (N19476, N19468, N18983, N15135);
nor NOR4 (N19477, N19475, N3556, N1851, N5133);
not NOT1 (N19478, N19463);
xor XOR2 (N19479, N19473, N14327);
or OR2 (N19480, N19478, N150);
not NOT1 (N19481, N19472);
not NOT1 (N19482, N19481);
or OR3 (N19483, N19482, N19436, N5185);
nand NAND4 (N19484, N19474, N8414, N7790, N6133);
buf BUF1 (N19485, N19483);
or OR2 (N19486, N19471, N592);
buf BUF1 (N19487, N19477);
not NOT1 (N19488, N19465);
not NOT1 (N19489, N19464);
and AND4 (N19490, N19487, N8024, N1555, N15682);
or OR3 (N19491, N19486, N16160, N9785);
and AND4 (N19492, N19489, N14810, N12377, N6458);
nand NAND2 (N19493, N19485, N19333);
not NOT1 (N19494, N19492);
buf BUF1 (N19495, N19479);
not NOT1 (N19496, N19488);
nor NOR4 (N19497, N19494, N12146, N18711, N2017);
nor NOR3 (N19498, N19470, N14058, N13013);
or OR4 (N19499, N19476, N3396, N6138, N10448);
nor NOR3 (N19500, N19480, N15449, N11907);
or OR4 (N19501, N19491, N8572, N4202, N7414);
and AND3 (N19502, N19493, N876, N4897);
not NOT1 (N19503, N19490);
nand NAND4 (N19504, N19503, N10845, N3109, N2562);
nor NOR4 (N19505, N19500, N12087, N14072, N4732);
and AND2 (N19506, N19484, N17982);
and AND2 (N19507, N19505, N15146);
buf BUF1 (N19508, N19499);
not NOT1 (N19509, N19495);
nor NOR3 (N19510, N19508, N17318, N8428);
not NOT1 (N19511, N19509);
nand NAND3 (N19512, N19496, N10982, N11063);
and AND4 (N19513, N19507, N4546, N6669, N14019);
buf BUF1 (N19514, N19506);
or OR4 (N19515, N19510, N11358, N17196, N14988);
and AND3 (N19516, N19504, N12031, N4587);
buf BUF1 (N19517, N19502);
nor NOR4 (N19518, N19514, N8012, N2010, N10091);
nand NAND3 (N19519, N19511, N16803, N10817);
xor XOR2 (N19520, N19501, N9748);
and AND2 (N19521, N19519, N3826);
and AND2 (N19522, N19521, N11461);
xor XOR2 (N19523, N19522, N13989);
buf BUF1 (N19524, N19498);
xor XOR2 (N19525, N19518, N2517);
not NOT1 (N19526, N19524);
nand NAND3 (N19527, N19516, N8635, N12216);
nor NOR3 (N19528, N19497, N16637, N13222);
or OR2 (N19529, N19517, N666);
buf BUF1 (N19530, N19527);
nand NAND2 (N19531, N19513, N8736);
nand NAND3 (N19532, N19528, N10516, N2333);
nor NOR3 (N19533, N19526, N10219, N17693);
or OR4 (N19534, N19515, N8297, N4884, N14128);
buf BUF1 (N19535, N19523);
or OR4 (N19536, N19512, N11013, N10551, N7889);
not NOT1 (N19537, N19536);
and AND2 (N19538, N19533, N1644);
xor XOR2 (N19539, N19537, N15671);
and AND2 (N19540, N19539, N9719);
not NOT1 (N19541, N19534);
xor XOR2 (N19542, N19538, N10806);
and AND4 (N19543, N19531, N3288, N18687, N9973);
buf BUF1 (N19544, N19525);
and AND4 (N19545, N19540, N17737, N14882, N8937);
nand NAND4 (N19546, N19541, N5358, N15150, N9276);
or OR4 (N19547, N19530, N12823, N956, N233);
nand NAND4 (N19548, N19535, N1131, N5605, N683);
xor XOR2 (N19549, N19520, N6858);
nor NOR3 (N19550, N19548, N9457, N1350);
nand NAND4 (N19551, N19546, N12075, N675, N3765);
nor NOR4 (N19552, N19549, N10293, N8391, N5454);
buf BUF1 (N19553, N19552);
xor XOR2 (N19554, N19547, N3346);
nor NOR2 (N19555, N19551, N14234);
nor NOR3 (N19556, N19553, N1623, N7914);
xor XOR2 (N19557, N19556, N5206);
not NOT1 (N19558, N19554);
buf BUF1 (N19559, N19542);
or OR3 (N19560, N19545, N7615, N8707);
not NOT1 (N19561, N19544);
or OR2 (N19562, N19555, N15718);
nand NAND4 (N19563, N19557, N19100, N4596, N16677);
or OR3 (N19564, N19543, N412, N14092);
and AND3 (N19565, N19550, N7326, N16305);
buf BUF1 (N19566, N19532);
buf BUF1 (N19567, N19561);
or OR2 (N19568, N19562, N11948);
and AND4 (N19569, N19560, N5594, N2484, N7876);
xor XOR2 (N19570, N19559, N2252);
or OR2 (N19571, N19564, N4224);
nor NOR4 (N19572, N19565, N7009, N19244, N4350);
or OR3 (N19573, N19572, N11280, N2399);
nand NAND2 (N19574, N19569, N10801);
nor NOR3 (N19575, N19574, N10511, N19312);
and AND4 (N19576, N19568, N16470, N10296, N5210);
nand NAND2 (N19577, N19563, N19159);
nor NOR3 (N19578, N19566, N5558, N1813);
nor NOR3 (N19579, N19573, N18333, N12428);
not NOT1 (N19580, N19577);
nand NAND2 (N19581, N19578, N8000);
not NOT1 (N19582, N19529);
not NOT1 (N19583, N19571);
or OR2 (N19584, N19558, N4282);
xor XOR2 (N19585, N19576, N9738);
or OR3 (N19586, N19585, N16650, N9302);
nand NAND3 (N19587, N19582, N12718, N15777);
or OR4 (N19588, N19575, N4820, N19375, N12873);
not NOT1 (N19589, N19581);
nor NOR3 (N19590, N19589, N8138, N7080);
buf BUF1 (N19591, N19580);
xor XOR2 (N19592, N19583, N12121);
buf BUF1 (N19593, N19587);
nor NOR2 (N19594, N19591, N8827);
buf BUF1 (N19595, N19579);
xor XOR2 (N19596, N19593, N16530);
buf BUF1 (N19597, N19594);
not NOT1 (N19598, N19570);
nor NOR3 (N19599, N19590, N9136, N16189);
buf BUF1 (N19600, N19592);
xor XOR2 (N19601, N19584, N10996);
nand NAND4 (N19602, N19595, N5055, N747, N19073);
or OR4 (N19603, N19586, N13455, N6993, N14000);
buf BUF1 (N19604, N19588);
buf BUF1 (N19605, N19602);
xor XOR2 (N19606, N19567, N18625);
and AND3 (N19607, N19605, N12052, N2316);
nor NOR2 (N19608, N19598, N16147);
nand NAND2 (N19609, N19604, N7640);
nor NOR3 (N19610, N19608, N17367, N2073);
and AND2 (N19611, N19610, N13476);
nand NAND4 (N19612, N19609, N6915, N17988, N6970);
or OR2 (N19613, N19601, N7880);
nor NOR2 (N19614, N19599, N15227);
and AND4 (N19615, N19611, N11095, N17658, N3842);
buf BUF1 (N19616, N19600);
and AND2 (N19617, N19613, N6636);
buf BUF1 (N19618, N19596);
or OR2 (N19619, N19615, N9448);
and AND3 (N19620, N19616, N6544, N6654);
nand NAND2 (N19621, N19619, N5937);
buf BUF1 (N19622, N19620);
and AND3 (N19623, N19606, N10152, N19058);
and AND4 (N19624, N19607, N4968, N17966, N15765);
nand NAND4 (N19625, N19618, N914, N11916, N11176);
not NOT1 (N19626, N19625);
or OR3 (N19627, N19624, N9498, N4450);
or OR4 (N19628, N19626, N4272, N9417, N13111);
xor XOR2 (N19629, N19628, N2321);
nor NOR4 (N19630, N19617, N6434, N9733, N19272);
nor NOR3 (N19631, N19627, N16751, N4130);
nor NOR4 (N19632, N19597, N2072, N11324, N6203);
buf BUF1 (N19633, N19621);
xor XOR2 (N19634, N19623, N4911);
buf BUF1 (N19635, N19622);
nor NOR2 (N19636, N19635, N9644);
or OR2 (N19637, N19603, N14992);
buf BUF1 (N19638, N19612);
not NOT1 (N19639, N19636);
or OR2 (N19640, N19614, N17447);
and AND2 (N19641, N19638, N12644);
not NOT1 (N19642, N19630);
buf BUF1 (N19643, N19629);
and AND4 (N19644, N19631, N2149, N9176, N329);
and AND4 (N19645, N19644, N11237, N13375, N2710);
buf BUF1 (N19646, N19641);
xor XOR2 (N19647, N19634, N1415);
xor XOR2 (N19648, N19647, N3356);
not NOT1 (N19649, N19643);
not NOT1 (N19650, N19648);
or OR4 (N19651, N19642, N8937, N6062, N5334);
not NOT1 (N19652, N19632);
buf BUF1 (N19653, N19646);
not NOT1 (N19654, N19645);
not NOT1 (N19655, N19637);
buf BUF1 (N19656, N19640);
xor XOR2 (N19657, N19633, N17702);
nand NAND2 (N19658, N19639, N4993);
not NOT1 (N19659, N19658);
buf BUF1 (N19660, N19650);
not NOT1 (N19661, N19653);
nand NAND3 (N19662, N19661, N10320, N18295);
nor NOR2 (N19663, N19651, N12031);
nor NOR4 (N19664, N19662, N12069, N4083, N15685);
and AND3 (N19665, N19657, N9375, N4129);
buf BUF1 (N19666, N19660);
not NOT1 (N19667, N19659);
not NOT1 (N19668, N19665);
and AND4 (N19669, N19668, N48, N18154, N2911);
nand NAND4 (N19670, N19667, N488, N17037, N15206);
nor NOR2 (N19671, N19666, N16147);
xor XOR2 (N19672, N19656, N1542);
and AND2 (N19673, N19670, N16979);
xor XOR2 (N19674, N19649, N6402);
and AND4 (N19675, N19673, N1459, N19581, N13073);
xor XOR2 (N19676, N19671, N889);
nand NAND2 (N19677, N19672, N16401);
and AND2 (N19678, N19675, N17849);
buf BUF1 (N19679, N19664);
and AND4 (N19680, N19678, N8365, N10774, N5733);
not NOT1 (N19681, N19674);
nand NAND2 (N19682, N19676, N17893);
xor XOR2 (N19683, N19663, N3527);
or OR3 (N19684, N19683, N17512, N18201);
or OR4 (N19685, N19682, N16048, N9224, N17119);
and AND2 (N19686, N19654, N4221);
nor NOR4 (N19687, N19684, N10737, N19458, N2045);
not NOT1 (N19688, N19680);
nor NOR3 (N19689, N19681, N5752, N12060);
buf BUF1 (N19690, N19679);
nor NOR2 (N19691, N19655, N3352);
nand NAND4 (N19692, N19688, N9524, N19262, N17858);
buf BUF1 (N19693, N19686);
nor NOR4 (N19694, N19687, N14074, N1613, N4212);
and AND2 (N19695, N19694, N9202);
or OR3 (N19696, N19690, N13851, N17816);
or OR4 (N19697, N19652, N11805, N16703, N7527);
xor XOR2 (N19698, N19669, N17932);
not NOT1 (N19699, N19697);
and AND4 (N19700, N19696, N12483, N17053, N10965);
not NOT1 (N19701, N19693);
nand NAND3 (N19702, N19685, N4995, N9292);
nand NAND3 (N19703, N19700, N2252, N12931);
nor NOR2 (N19704, N19698, N5960);
nor NOR2 (N19705, N19699, N6445);
xor XOR2 (N19706, N19701, N12022);
not NOT1 (N19707, N19689);
xor XOR2 (N19708, N19704, N11051);
nand NAND2 (N19709, N19702, N16302);
nor NOR3 (N19710, N19677, N17021, N13974);
and AND2 (N19711, N19703, N8961);
or OR4 (N19712, N19692, N4385, N11521, N9414);
xor XOR2 (N19713, N19707, N19596);
xor XOR2 (N19714, N19695, N8844);
nor NOR2 (N19715, N19711, N16591);
buf BUF1 (N19716, N19714);
nor NOR2 (N19717, N19716, N17447);
and AND2 (N19718, N19710, N12686);
buf BUF1 (N19719, N19691);
or OR4 (N19720, N19708, N375, N1504, N11888);
or OR4 (N19721, N19709, N14986, N1288, N14793);
or OR4 (N19722, N19712, N16507, N11283, N17658);
nor NOR2 (N19723, N19713, N11225);
not NOT1 (N19724, N19723);
nand NAND2 (N19725, N19715, N19592);
nor NOR2 (N19726, N19706, N5927);
or OR2 (N19727, N19718, N14351);
buf BUF1 (N19728, N19719);
and AND3 (N19729, N19722, N2006, N14520);
and AND2 (N19730, N19729, N9346);
or OR3 (N19731, N19721, N16309, N2036);
nand NAND4 (N19732, N19727, N8777, N12135, N18327);
buf BUF1 (N19733, N19728);
xor XOR2 (N19734, N19720, N17856);
and AND2 (N19735, N19731, N6626);
and AND4 (N19736, N19733, N1924, N11373, N9244);
not NOT1 (N19737, N19724);
nor NOR4 (N19738, N19717, N16174, N223, N5626);
xor XOR2 (N19739, N19732, N10027);
not NOT1 (N19740, N19734);
xor XOR2 (N19741, N19735, N2042);
buf BUF1 (N19742, N19705);
and AND4 (N19743, N19740, N11549, N14696, N5408);
buf BUF1 (N19744, N19741);
nor NOR2 (N19745, N19737, N16562);
or OR2 (N19746, N19742, N19642);
buf BUF1 (N19747, N19736);
buf BUF1 (N19748, N19744);
not NOT1 (N19749, N19747);
buf BUF1 (N19750, N19746);
nand NAND3 (N19751, N19725, N8814, N7086);
buf BUF1 (N19752, N19751);
xor XOR2 (N19753, N19739, N17660);
nand NAND3 (N19754, N19726, N18276, N15935);
and AND3 (N19755, N19749, N1483, N142);
buf BUF1 (N19756, N19753);
nand NAND2 (N19757, N19752, N15182);
or OR3 (N19758, N19756, N17394, N3468);
and AND2 (N19759, N19745, N6921);
not NOT1 (N19760, N19738);
xor XOR2 (N19761, N19730, N5525);
and AND2 (N19762, N19750, N13232);
not NOT1 (N19763, N19760);
not NOT1 (N19764, N19763);
nand NAND4 (N19765, N19755, N19709, N8334, N15239);
not NOT1 (N19766, N19761);
buf BUF1 (N19767, N19757);
buf BUF1 (N19768, N19766);
xor XOR2 (N19769, N19743, N10293);
nand NAND4 (N19770, N19769, N484, N18513, N7966);
xor XOR2 (N19771, N19754, N9520);
and AND4 (N19772, N19771, N10476, N14994, N10337);
xor XOR2 (N19773, N19759, N407);
nand NAND4 (N19774, N19764, N14333, N15143, N12649);
buf BUF1 (N19775, N19758);
nand NAND4 (N19776, N19767, N3830, N18597, N6401);
nand NAND3 (N19777, N19775, N10830, N3361);
buf BUF1 (N19778, N19762);
xor XOR2 (N19779, N19748, N13007);
nor NOR2 (N19780, N19765, N12253);
and AND2 (N19781, N19774, N5375);
nand NAND4 (N19782, N19773, N15662, N3089, N18013);
buf BUF1 (N19783, N19772);
and AND3 (N19784, N19783, N2861, N11241);
not NOT1 (N19785, N19782);
not NOT1 (N19786, N19778);
or OR3 (N19787, N19770, N12657, N10060);
nor NOR3 (N19788, N19780, N1198, N11577);
nor NOR4 (N19789, N19788, N18662, N105, N19319);
and AND3 (N19790, N19768, N9679, N18713);
or OR3 (N19791, N19787, N6614, N14402);
nand NAND4 (N19792, N19790, N14515, N8070, N3147);
or OR2 (N19793, N19785, N16463);
or OR4 (N19794, N19791, N12030, N17129, N10185);
buf BUF1 (N19795, N19779);
nand NAND3 (N19796, N19784, N5842, N15530);
and AND4 (N19797, N19796, N3884, N17176, N9544);
or OR2 (N19798, N19786, N10429);
nand NAND2 (N19799, N19793, N17933);
buf BUF1 (N19800, N19781);
nand NAND3 (N19801, N19797, N3485, N14824);
xor XOR2 (N19802, N19800, N9494);
nor NOR4 (N19803, N19777, N7664, N6622, N10640);
nor NOR2 (N19804, N19776, N3227);
nand NAND2 (N19805, N19792, N16002);
not NOT1 (N19806, N19798);
or OR2 (N19807, N19789, N6872);
xor XOR2 (N19808, N19805, N5564);
nand NAND4 (N19809, N19803, N18606, N2297, N3650);
or OR2 (N19810, N19794, N19436);
nand NAND3 (N19811, N19807, N16291, N12325);
and AND3 (N19812, N19809, N7075, N13433);
and AND3 (N19813, N19801, N16234, N13763);
nand NAND2 (N19814, N19812, N637);
or OR3 (N19815, N19806, N2235, N7880);
or OR2 (N19816, N19802, N4266);
nand NAND3 (N19817, N19811, N5348, N19276);
nor NOR4 (N19818, N19799, N12078, N9898, N14618);
not NOT1 (N19819, N19810);
xor XOR2 (N19820, N19818, N10570);
buf BUF1 (N19821, N19795);
or OR2 (N19822, N19820, N9858);
not NOT1 (N19823, N19816);
buf BUF1 (N19824, N19808);
nor NOR3 (N19825, N19821, N5333, N661);
and AND2 (N19826, N19819, N4736);
not NOT1 (N19827, N19824);
not NOT1 (N19828, N19804);
buf BUF1 (N19829, N19828);
nor NOR4 (N19830, N19813, N12762, N19087, N4788);
nor NOR3 (N19831, N19827, N2804, N4798);
and AND4 (N19832, N19822, N5878, N1605, N11015);
nor NOR4 (N19833, N19832, N17286, N10799, N7093);
nor NOR3 (N19834, N19825, N4205, N10381);
nand NAND4 (N19835, N19817, N6655, N2422, N14814);
xor XOR2 (N19836, N19834, N4681);
buf BUF1 (N19837, N19829);
or OR2 (N19838, N19826, N10512);
and AND2 (N19839, N19814, N9019);
xor XOR2 (N19840, N19839, N3668);
nor NOR4 (N19841, N19815, N5783, N11237, N17255);
or OR2 (N19842, N19836, N6853);
and AND2 (N19843, N19831, N18563);
or OR2 (N19844, N19840, N71);
or OR2 (N19845, N19842, N1396);
xor XOR2 (N19846, N19844, N11428);
nor NOR3 (N19847, N19835, N9946, N5990);
and AND3 (N19848, N19845, N662, N8609);
and AND3 (N19849, N19823, N57, N15438);
nand NAND4 (N19850, N19837, N14830, N5129, N7267);
buf BUF1 (N19851, N19849);
and AND3 (N19852, N19846, N19465, N17767);
xor XOR2 (N19853, N19833, N13273);
xor XOR2 (N19854, N19841, N14272);
and AND2 (N19855, N19848, N16650);
or OR4 (N19856, N19838, N1628, N8992, N3003);
nand NAND3 (N19857, N19847, N5247, N19573);
nand NAND4 (N19858, N19850, N13796, N19059, N11947);
buf BUF1 (N19859, N19843);
nand NAND4 (N19860, N19856, N6162, N7091, N2604);
xor XOR2 (N19861, N19830, N14576);
and AND4 (N19862, N19854, N6516, N4236, N11677);
or OR2 (N19863, N19855, N12684);
buf BUF1 (N19864, N19860);
not NOT1 (N19865, N19862);
buf BUF1 (N19866, N19853);
xor XOR2 (N19867, N19864, N17318);
buf BUF1 (N19868, N19859);
not NOT1 (N19869, N19865);
buf BUF1 (N19870, N19851);
xor XOR2 (N19871, N19867, N4159);
and AND4 (N19872, N19869, N3444, N1653, N9139);
buf BUF1 (N19873, N19861);
nand NAND2 (N19874, N19852, N14876);
nor NOR2 (N19875, N19872, N1647);
not NOT1 (N19876, N19863);
not NOT1 (N19877, N19875);
nand NAND3 (N19878, N19870, N17632, N6114);
or OR4 (N19879, N19857, N13913, N12238, N11230);
buf BUF1 (N19880, N19879);
or OR2 (N19881, N19866, N7613);
nor NOR4 (N19882, N19858, N13065, N7340, N3142);
or OR4 (N19883, N19882, N3294, N14342, N15963);
xor XOR2 (N19884, N19873, N5760);
not NOT1 (N19885, N19874);
or OR3 (N19886, N19876, N19671, N13283);
xor XOR2 (N19887, N19883, N18709);
buf BUF1 (N19888, N19886);
nor NOR3 (N19889, N19885, N2117, N8587);
nand NAND4 (N19890, N19868, N2602, N8527, N2630);
and AND4 (N19891, N19877, N19769, N14550, N8073);
or OR4 (N19892, N19871, N10026, N11723, N7267);
nand NAND3 (N19893, N19890, N16956, N1661);
xor XOR2 (N19894, N19881, N19281);
and AND4 (N19895, N19880, N3320, N1269, N11463);
or OR4 (N19896, N19878, N2762, N14765, N9438);
xor XOR2 (N19897, N19889, N12961);
or OR4 (N19898, N19884, N14745, N6802, N14191);
nand NAND3 (N19899, N19898, N1645, N1132);
xor XOR2 (N19900, N19888, N8637);
nor NOR2 (N19901, N19887, N2466);
nor NOR3 (N19902, N19896, N10419, N3707);
not NOT1 (N19903, N19894);
and AND3 (N19904, N19899, N7175, N4575);
or OR2 (N19905, N19901, N10146);
xor XOR2 (N19906, N19905, N12058);
nand NAND2 (N19907, N19903, N2738);
nand NAND2 (N19908, N19900, N18099);
xor XOR2 (N19909, N19893, N15260);
or OR2 (N19910, N19909, N14317);
xor XOR2 (N19911, N19910, N18580);
xor XOR2 (N19912, N19892, N14358);
or OR3 (N19913, N19897, N18421, N9447);
nand NAND3 (N19914, N19913, N17504, N4889);
not NOT1 (N19915, N19908);
nor NOR3 (N19916, N19912, N5208, N5512);
and AND4 (N19917, N19916, N9345, N6442, N16800);
and AND2 (N19918, N19917, N14435);
not NOT1 (N19919, N19914);
nor NOR4 (N19920, N19911, N9067, N6823, N18609);
or OR3 (N19921, N19906, N15303, N18770);
or OR2 (N19922, N19918, N15502);
nand NAND4 (N19923, N19904, N2940, N18608, N9240);
nand NAND3 (N19924, N19895, N13253, N8375);
not NOT1 (N19925, N19920);
nor NOR2 (N19926, N19925, N18705);
and AND2 (N19927, N19919, N134);
nor NOR2 (N19928, N19891, N18346);
nor NOR3 (N19929, N19921, N7413, N17525);
nand NAND4 (N19930, N19928, N19834, N5263, N19748);
buf BUF1 (N19931, N19907);
nor NOR3 (N19932, N19922, N14189, N3705);
nor NOR4 (N19933, N19923, N7392, N18508, N18929);
nand NAND2 (N19934, N19902, N13993);
and AND2 (N19935, N19933, N10333);
nor NOR2 (N19936, N19935, N10384);
nor NOR4 (N19937, N19915, N18932, N15496, N1121);
or OR3 (N19938, N19929, N11455, N1892);
xor XOR2 (N19939, N19930, N15338);
or OR3 (N19940, N19936, N15254, N15955);
buf BUF1 (N19941, N19939);
nor NOR4 (N19942, N19931, N8879, N9091, N17016);
and AND3 (N19943, N19926, N12951, N10065);
nor NOR4 (N19944, N19932, N9220, N8869, N17490);
xor XOR2 (N19945, N19927, N14339);
xor XOR2 (N19946, N19941, N19287);
or OR3 (N19947, N19940, N3940, N9923);
nand NAND4 (N19948, N19947, N6187, N9370, N15689);
xor XOR2 (N19949, N19945, N4668);
buf BUF1 (N19950, N19946);
or OR4 (N19951, N19943, N4643, N11745, N14852);
and AND2 (N19952, N19937, N16678);
and AND4 (N19953, N19942, N12881, N16748, N11607);
and AND2 (N19954, N19944, N373);
nor NOR3 (N19955, N19948, N2802, N17283);
xor XOR2 (N19956, N19938, N10120);
or OR4 (N19957, N19924, N19784, N16846, N582);
nor NOR3 (N19958, N19956, N14859, N9298);
and AND4 (N19959, N19958, N5984, N19374, N9457);
nor NOR3 (N19960, N19952, N1050, N5913);
and AND2 (N19961, N19959, N1843);
and AND3 (N19962, N19960, N2408, N2773);
buf BUF1 (N19963, N19934);
not NOT1 (N19964, N19951);
xor XOR2 (N19965, N19955, N17454);
nand NAND3 (N19966, N19961, N5426, N8994);
and AND4 (N19967, N19964, N1109, N5891, N9924);
buf BUF1 (N19968, N19965);
not NOT1 (N19969, N19966);
not NOT1 (N19970, N19967);
nor NOR3 (N19971, N19950, N19074, N14551);
xor XOR2 (N19972, N19954, N5982);
or OR3 (N19973, N19969, N15675, N18890);
or OR2 (N19974, N19972, N847);
buf BUF1 (N19975, N19962);
and AND2 (N19976, N19971, N787);
buf BUF1 (N19977, N19953);
nor NOR3 (N19978, N19970, N9868, N9921);
and AND4 (N19979, N19976, N10591, N10236, N14806);
xor XOR2 (N19980, N19974, N7559);
xor XOR2 (N19981, N19968, N19422);
or OR4 (N19982, N19980, N7708, N6151, N7201);
buf BUF1 (N19983, N19957);
or OR3 (N19984, N19963, N14942, N3267);
buf BUF1 (N19985, N19973);
nor NOR2 (N19986, N19981, N1427);
and AND4 (N19987, N19979, N8588, N17712, N4393);
or OR2 (N19988, N19985, N6113);
nor NOR3 (N19989, N19975, N12408, N7556);
or OR3 (N19990, N19977, N19167, N2424);
buf BUF1 (N19991, N19987);
not NOT1 (N19992, N19988);
xor XOR2 (N19993, N19986, N779);
and AND4 (N19994, N19990, N16505, N11093, N10445);
xor XOR2 (N19995, N19993, N14143);
nand NAND4 (N19996, N19982, N16488, N12882, N1073);
not NOT1 (N19997, N19996);
nor NOR2 (N19998, N19949, N15080);
or OR3 (N19999, N19991, N7442, N10806);
nor NOR4 (N20000, N19989, N12076, N253, N12155);
not NOT1 (N20001, N19992);
buf BUF1 (N20002, N19998);
nand NAND3 (N20003, N19999, N9466, N14820);
and AND4 (N20004, N19984, N19147, N4994, N1355);
not NOT1 (N20005, N19978);
not NOT1 (N20006, N19983);
xor XOR2 (N20007, N20003, N1872);
nand NAND2 (N20008, N20001, N9154);
xor XOR2 (N20009, N20007, N10918);
nor NOR4 (N20010, N19997, N4935, N17418, N7034);
and AND2 (N20011, N20009, N16646);
nor NOR4 (N20012, N20011, N16787, N2895, N1907);
nor NOR2 (N20013, N19995, N18440);
not NOT1 (N20014, N20012);
nand NAND3 (N20015, N20008, N5324, N5041);
nor NOR3 (N20016, N20014, N13425, N15848);
nand NAND2 (N20017, N20015, N6337);
nand NAND2 (N20018, N20016, N4068);
and AND4 (N20019, N19994, N15164, N17205, N13682);
nor NOR3 (N20020, N20018, N3778, N17949);
and AND4 (N20021, N20020, N12053, N16172, N10803);
or OR4 (N20022, N20006, N7830, N17386, N8940);
or OR4 (N20023, N20004, N13918, N7446, N12021);
or OR3 (N20024, N20000, N6469, N1407);
not NOT1 (N20025, N20019);
nor NOR4 (N20026, N20024, N4019, N6474, N8786);
nor NOR4 (N20027, N20023, N8606, N8422, N6367);
and AND2 (N20028, N20026, N19885);
and AND4 (N20029, N20013, N15214, N17327, N18280);
not NOT1 (N20030, N20027);
or OR3 (N20031, N20005, N1427, N3112);
not NOT1 (N20032, N20028);
and AND2 (N20033, N20031, N13720);
and AND3 (N20034, N20030, N7509, N19519);
and AND4 (N20035, N20002, N17770, N490, N7589);
buf BUF1 (N20036, N20010);
and AND3 (N20037, N20032, N8253, N4662);
nand NAND4 (N20038, N20022, N2299, N19923, N12490);
nand NAND2 (N20039, N20036, N18513);
not NOT1 (N20040, N20029);
xor XOR2 (N20041, N20025, N19646);
nor NOR4 (N20042, N20039, N19165, N16064, N14582);
and AND4 (N20043, N20021, N13751, N13249, N17649);
and AND3 (N20044, N20043, N10715, N4795);
nand NAND3 (N20045, N20040, N2168, N18500);
xor XOR2 (N20046, N20034, N7161);
not NOT1 (N20047, N20038);
nand NAND4 (N20048, N20044, N16048, N16162, N7518);
buf BUF1 (N20049, N20033);
buf BUF1 (N20050, N20035);
xor XOR2 (N20051, N20047, N17795);
nor NOR4 (N20052, N20017, N18992, N14678, N11987);
nand NAND3 (N20053, N20052, N15919, N18712);
nor NOR3 (N20054, N20046, N11346, N13234);
xor XOR2 (N20055, N20050, N4443);
nor NOR4 (N20056, N20037, N6701, N3903, N3924);
and AND2 (N20057, N20041, N8305);
buf BUF1 (N20058, N20051);
nor NOR4 (N20059, N20057, N14088, N10317, N9555);
buf BUF1 (N20060, N20054);
nand NAND4 (N20061, N20059, N14943, N7106, N9628);
nand NAND4 (N20062, N20056, N2353, N14566, N14083);
not NOT1 (N20063, N20062);
and AND2 (N20064, N20049, N5016);
nor NOR4 (N20065, N20045, N8934, N4283, N8150);
nand NAND2 (N20066, N20053, N16380);
nor NOR3 (N20067, N20065, N1929, N3493);
not NOT1 (N20068, N20042);
nand NAND2 (N20069, N20060, N8807);
or OR3 (N20070, N20066, N16305, N16327);
nand NAND3 (N20071, N20055, N18345, N19166);
buf BUF1 (N20072, N20067);
and AND2 (N20073, N20072, N25);
not NOT1 (N20074, N20070);
nand NAND4 (N20075, N20048, N7648, N4433, N17788);
nor NOR4 (N20076, N20071, N6294, N736, N8400);
or OR4 (N20077, N20073, N6340, N13291, N4873);
nor NOR3 (N20078, N20064, N927, N15101);
nand NAND4 (N20079, N20069, N14954, N1870, N15051);
nand NAND2 (N20080, N20061, N16194);
nor NOR2 (N20081, N20077, N18104);
xor XOR2 (N20082, N20075, N17471);
and AND2 (N20083, N20068, N2322);
or OR4 (N20084, N20080, N9355, N6558, N2903);
and AND4 (N20085, N20084, N12847, N14166, N15516);
not NOT1 (N20086, N20085);
buf BUF1 (N20087, N20063);
and AND4 (N20088, N20087, N14597, N1909, N14586);
not NOT1 (N20089, N20076);
nor NOR2 (N20090, N20088, N1525);
not NOT1 (N20091, N20083);
xor XOR2 (N20092, N20091, N11249);
or OR2 (N20093, N20079, N8095);
and AND2 (N20094, N20058, N14477);
nor NOR4 (N20095, N20074, N444, N8223, N4477);
or OR2 (N20096, N20092, N5853);
or OR4 (N20097, N20090, N6596, N894, N2902);
nor NOR3 (N20098, N20096, N15266, N12214);
nand NAND4 (N20099, N20089, N1959, N16297, N7638);
buf BUF1 (N20100, N20098);
buf BUF1 (N20101, N20082);
buf BUF1 (N20102, N20100);
buf BUF1 (N20103, N20097);
and AND4 (N20104, N20101, N3247, N15744, N7771);
buf BUF1 (N20105, N20081);
or OR3 (N20106, N20094, N5987, N13796);
buf BUF1 (N20107, N20099);
nor NOR3 (N20108, N20107, N12870, N17693);
xor XOR2 (N20109, N20102, N2880);
and AND2 (N20110, N20086, N13941);
nand NAND3 (N20111, N20110, N2018, N18435);
nand NAND4 (N20112, N20095, N10024, N7785, N1435);
or OR2 (N20113, N20108, N19933);
nor NOR2 (N20114, N20113, N14897);
nand NAND2 (N20115, N20103, N7274);
or OR4 (N20116, N20109, N4571, N17611, N1619);
nor NOR2 (N20117, N20104, N1387);
and AND3 (N20118, N20116, N3906, N17199);
xor XOR2 (N20119, N20093, N8121);
nor NOR2 (N20120, N20078, N1607);
nand NAND3 (N20121, N20118, N1051, N1074);
or OR4 (N20122, N20105, N2779, N7387, N15112);
buf BUF1 (N20123, N20121);
nor NOR2 (N20124, N20119, N5670);
nor NOR3 (N20125, N20122, N1857, N19368);
not NOT1 (N20126, N20125);
nor NOR2 (N20127, N20114, N5421);
nand NAND4 (N20128, N20117, N4199, N8014, N19594);
nor NOR2 (N20129, N20127, N11414);
not NOT1 (N20130, N20120);
not NOT1 (N20131, N20123);
or OR2 (N20132, N20126, N8170);
xor XOR2 (N20133, N20111, N7528);
or OR3 (N20134, N20128, N13361, N14269);
or OR3 (N20135, N20115, N16083, N7436);
not NOT1 (N20136, N20131);
xor XOR2 (N20137, N20132, N19740);
or OR2 (N20138, N20134, N17363);
nand NAND4 (N20139, N20136, N6182, N4746, N3180);
not NOT1 (N20140, N20129);
or OR2 (N20141, N20139, N18269);
and AND2 (N20142, N20133, N14676);
xor XOR2 (N20143, N20130, N19131);
buf BUF1 (N20144, N20112);
not NOT1 (N20145, N20142);
xor XOR2 (N20146, N20140, N1128);
nor NOR2 (N20147, N20146, N14330);
nand NAND2 (N20148, N20137, N9530);
and AND3 (N20149, N20147, N9659, N4254);
or OR2 (N20150, N20145, N2253);
xor XOR2 (N20151, N20148, N17785);
or OR4 (N20152, N20138, N15416, N1524, N8644);
or OR2 (N20153, N20141, N5239);
xor XOR2 (N20154, N20150, N16626);
nor NOR2 (N20155, N20124, N3634);
nor NOR3 (N20156, N20151, N18576, N6112);
not NOT1 (N20157, N20135);
not NOT1 (N20158, N20152);
buf BUF1 (N20159, N20158);
buf BUF1 (N20160, N20154);
xor XOR2 (N20161, N20155, N10043);
buf BUF1 (N20162, N20157);
xor XOR2 (N20163, N20156, N7206);
nor NOR2 (N20164, N20161, N16356);
or OR3 (N20165, N20149, N9756, N9476);
buf BUF1 (N20166, N20106);
xor XOR2 (N20167, N20164, N15823);
not NOT1 (N20168, N20162);
buf BUF1 (N20169, N20166);
nor NOR2 (N20170, N20163, N4460);
nor NOR4 (N20171, N20143, N1870, N3773, N3472);
nor NOR3 (N20172, N20144, N11694, N10547);
or OR4 (N20173, N20168, N6454, N343, N17018);
xor XOR2 (N20174, N20165, N12527);
xor XOR2 (N20175, N20174, N6357);
xor XOR2 (N20176, N20171, N17869);
and AND3 (N20177, N20153, N12740, N653);
not NOT1 (N20178, N20170);
not NOT1 (N20179, N20175);
and AND2 (N20180, N20176, N1330);
not NOT1 (N20181, N20167);
nand NAND4 (N20182, N20178, N13093, N10903, N7213);
nand NAND4 (N20183, N20179, N61, N15159, N3124);
nor NOR4 (N20184, N20172, N14297, N18486, N7881);
not NOT1 (N20185, N20169);
nand NAND3 (N20186, N20180, N891, N13311);
buf BUF1 (N20187, N20181);
not NOT1 (N20188, N20173);
and AND3 (N20189, N20184, N15907, N2005);
buf BUF1 (N20190, N20189);
buf BUF1 (N20191, N20185);
xor XOR2 (N20192, N20177, N13746);
not NOT1 (N20193, N20190);
buf BUF1 (N20194, N20182);
or OR3 (N20195, N20194, N9125, N9689);
nand NAND2 (N20196, N20188, N18314);
xor XOR2 (N20197, N20186, N16816);
buf BUF1 (N20198, N20192);
or OR2 (N20199, N20198, N4443);
and AND4 (N20200, N20187, N6595, N256, N14472);
and AND2 (N20201, N20197, N20161);
or OR2 (N20202, N20159, N4571);
nor NOR4 (N20203, N20199, N19859, N8358, N10235);
xor XOR2 (N20204, N20196, N15505);
or OR4 (N20205, N20160, N9524, N8000, N14346);
xor XOR2 (N20206, N20191, N7306);
nand NAND3 (N20207, N20205, N2371, N17977);
nor NOR3 (N20208, N20203, N18736, N5553);
nand NAND3 (N20209, N20200, N12624, N13486);
xor XOR2 (N20210, N20204, N8966);
buf BUF1 (N20211, N20183);
buf BUF1 (N20212, N20195);
not NOT1 (N20213, N20201);
not NOT1 (N20214, N20212);
or OR4 (N20215, N20193, N12488, N8946, N5966);
and AND4 (N20216, N20206, N16777, N4113, N5000);
not NOT1 (N20217, N20214);
and AND2 (N20218, N20211, N2865);
nand NAND4 (N20219, N20209, N13599, N11953, N2215);
nand NAND3 (N20220, N20215, N14608, N10774);
buf BUF1 (N20221, N20210);
not NOT1 (N20222, N20219);
buf BUF1 (N20223, N20218);
nand NAND4 (N20224, N20220, N2042, N16291, N19774);
xor XOR2 (N20225, N20222, N16842);
xor XOR2 (N20226, N20225, N5421);
xor XOR2 (N20227, N20217, N9111);
xor XOR2 (N20228, N20223, N17034);
not NOT1 (N20229, N20224);
nand NAND3 (N20230, N20202, N1626, N11704);
and AND4 (N20231, N20226, N452, N7447, N15418);
nor NOR3 (N20232, N20221, N10309, N13382);
not NOT1 (N20233, N20232);
nand NAND4 (N20234, N20228, N3337, N6530, N9396);
and AND4 (N20235, N20227, N7477, N7825, N10844);
buf BUF1 (N20236, N20235);
buf BUF1 (N20237, N20236);
nor NOR4 (N20238, N20230, N7757, N14873, N2684);
nor NOR3 (N20239, N20237, N9286, N1133);
and AND4 (N20240, N20239, N20044, N11822, N1569);
nor NOR2 (N20241, N20216, N10771);
not NOT1 (N20242, N20234);
not NOT1 (N20243, N20241);
nand NAND4 (N20244, N20243, N506, N6989, N9061);
xor XOR2 (N20245, N20238, N5296);
or OR2 (N20246, N20208, N6560);
and AND3 (N20247, N20207, N18021, N14974);
not NOT1 (N20248, N20246);
buf BUF1 (N20249, N20247);
nor NOR4 (N20250, N20240, N5485, N4304, N6500);
nand NAND4 (N20251, N20248, N8649, N6302, N16471);
nand NAND2 (N20252, N20245, N7317);
buf BUF1 (N20253, N20252);
buf BUF1 (N20254, N20231);
and AND4 (N20255, N20244, N11139, N3869, N3987);
not NOT1 (N20256, N20249);
not NOT1 (N20257, N20213);
buf BUF1 (N20258, N20250);
or OR2 (N20259, N20257, N18428);
buf BUF1 (N20260, N20251);
nor NOR4 (N20261, N20256, N16570, N17611, N13414);
buf BUF1 (N20262, N20260);
and AND3 (N20263, N20255, N9341, N19693);
buf BUF1 (N20264, N20233);
nor NOR3 (N20265, N20253, N4005, N6325);
xor XOR2 (N20266, N20261, N10061);
and AND3 (N20267, N20258, N18579, N14359);
buf BUF1 (N20268, N20263);
buf BUF1 (N20269, N20264);
not NOT1 (N20270, N20242);
not NOT1 (N20271, N20268);
buf BUF1 (N20272, N20266);
nand NAND4 (N20273, N20262, N13393, N11747, N8480);
or OR3 (N20274, N20267, N12433, N13536);
or OR2 (N20275, N20269, N10029);
and AND2 (N20276, N20259, N7901);
not NOT1 (N20277, N20265);
or OR2 (N20278, N20254, N17369);
buf BUF1 (N20279, N20275);
not NOT1 (N20280, N20271);
nand NAND4 (N20281, N20277, N12359, N8731, N9515);
xor XOR2 (N20282, N20229, N360);
buf BUF1 (N20283, N20270);
not NOT1 (N20284, N20278);
and AND2 (N20285, N20274, N9360);
or OR2 (N20286, N20285, N711);
nand NAND3 (N20287, N20272, N18966, N5971);
nor NOR3 (N20288, N20281, N15870, N4282);
xor XOR2 (N20289, N20286, N15609);
nand NAND3 (N20290, N20280, N18844, N12278);
not NOT1 (N20291, N20283);
buf BUF1 (N20292, N20279);
xor XOR2 (N20293, N20290, N8538);
nand NAND2 (N20294, N20282, N16327);
nor NOR2 (N20295, N20288, N11675);
xor XOR2 (N20296, N20293, N12616);
or OR4 (N20297, N20287, N19869, N19562, N3116);
buf BUF1 (N20298, N20292);
and AND2 (N20299, N20295, N14263);
nand NAND2 (N20300, N20276, N17852);
xor XOR2 (N20301, N20296, N1441);
nand NAND3 (N20302, N20301, N8832, N7182);
and AND4 (N20303, N20297, N8984, N20130, N12611);
or OR2 (N20304, N20298, N1257);
nand NAND4 (N20305, N20289, N13104, N19943, N15398);
or OR4 (N20306, N20284, N14816, N8139, N9541);
and AND2 (N20307, N20304, N17628);
or OR2 (N20308, N20300, N14150);
nor NOR2 (N20309, N20302, N15780);
and AND3 (N20310, N20306, N2731, N16820);
buf BUF1 (N20311, N20307);
not NOT1 (N20312, N20308);
nand NAND3 (N20313, N20294, N3107, N6371);
or OR2 (N20314, N20313, N14396);
or OR2 (N20315, N20273, N5020);
not NOT1 (N20316, N20314);
nand NAND3 (N20317, N20311, N16798, N18398);
buf BUF1 (N20318, N20303);
buf BUF1 (N20319, N20309);
nor NOR2 (N20320, N20305, N13543);
not NOT1 (N20321, N20299);
xor XOR2 (N20322, N20310, N1556);
or OR2 (N20323, N20312, N12444);
or OR2 (N20324, N20319, N8323);
nor NOR3 (N20325, N20321, N2893, N2721);
nor NOR4 (N20326, N20316, N17501, N6185, N6837);
xor XOR2 (N20327, N20320, N12731);
not NOT1 (N20328, N20291);
buf BUF1 (N20329, N20325);
buf BUF1 (N20330, N20317);
and AND4 (N20331, N20329, N2310, N8864, N17398);
xor XOR2 (N20332, N20323, N2153);
buf BUF1 (N20333, N20331);
nand NAND4 (N20334, N20327, N2311, N17636, N1639);
buf BUF1 (N20335, N20330);
buf BUF1 (N20336, N20326);
and AND2 (N20337, N20318, N3385);
xor XOR2 (N20338, N20335, N6565);
nand NAND2 (N20339, N20315, N16352);
nand NAND3 (N20340, N20336, N7828, N5029);
or OR4 (N20341, N20337, N12736, N7965, N3328);
and AND2 (N20342, N20334, N11815);
xor XOR2 (N20343, N20342, N5696);
nor NOR3 (N20344, N20341, N13314, N15474);
nand NAND3 (N20345, N20332, N16109, N17384);
xor XOR2 (N20346, N20339, N19421);
not NOT1 (N20347, N20343);
xor XOR2 (N20348, N20347, N7817);
xor XOR2 (N20349, N20346, N17242);
xor XOR2 (N20350, N20333, N2526);
and AND3 (N20351, N20348, N2707, N19508);
not NOT1 (N20352, N20328);
buf BUF1 (N20353, N20345);
not NOT1 (N20354, N20338);
and AND2 (N20355, N20350, N12203);
and AND3 (N20356, N20355, N5457, N6246);
not NOT1 (N20357, N20322);
buf BUF1 (N20358, N20344);
nand NAND4 (N20359, N20352, N1343, N13161, N18081);
nor NOR3 (N20360, N20357, N10594, N18342);
buf BUF1 (N20361, N20349);
nor NOR2 (N20362, N20356, N7017);
and AND3 (N20363, N20359, N15689, N6908);
not NOT1 (N20364, N20362);
not NOT1 (N20365, N20361);
nor NOR4 (N20366, N20358, N16246, N17590, N10518);
xor XOR2 (N20367, N20366, N351);
and AND4 (N20368, N20340, N14377, N9308, N13555);
not NOT1 (N20369, N20363);
buf BUF1 (N20370, N20367);
nor NOR3 (N20371, N20324, N8442, N18069);
xor XOR2 (N20372, N20353, N6434);
and AND3 (N20373, N20354, N17222, N1791);
or OR3 (N20374, N20370, N16372, N6901);
not NOT1 (N20375, N20365);
nand NAND4 (N20376, N20372, N4722, N16274, N17290);
nand NAND2 (N20377, N20374, N9066);
xor XOR2 (N20378, N20360, N13600);
buf BUF1 (N20379, N20351);
and AND2 (N20380, N20378, N13810);
buf BUF1 (N20381, N20376);
xor XOR2 (N20382, N20375, N5399);
not NOT1 (N20383, N20369);
nand NAND4 (N20384, N20377, N14554, N8707, N811);
nand NAND4 (N20385, N20368, N9159, N17897, N9723);
not NOT1 (N20386, N20381);
nand NAND3 (N20387, N20382, N909, N11946);
not NOT1 (N20388, N20386);
not NOT1 (N20389, N20379);
nand NAND2 (N20390, N20387, N10784);
not NOT1 (N20391, N20373);
buf BUF1 (N20392, N20383);
and AND4 (N20393, N20380, N18, N17944, N3248);
or OR4 (N20394, N20393, N15708, N11627, N17935);
buf BUF1 (N20395, N20385);
buf BUF1 (N20396, N20391);
or OR4 (N20397, N20392, N4459, N7142, N11312);
and AND2 (N20398, N20395, N8079);
buf BUF1 (N20399, N20396);
xor XOR2 (N20400, N20390, N12156);
and AND4 (N20401, N20397, N4054, N20175, N11316);
and AND3 (N20402, N20398, N18294, N5702);
xor XOR2 (N20403, N20364, N2054);
nor NOR4 (N20404, N20389, N5966, N3129, N9262);
and AND2 (N20405, N20388, N12884);
or OR3 (N20406, N20402, N916, N10245);
not NOT1 (N20407, N20384);
nor NOR4 (N20408, N20401, N1689, N7838, N19560);
buf BUF1 (N20409, N20408);
xor XOR2 (N20410, N20404, N9842);
buf BUF1 (N20411, N20400);
not NOT1 (N20412, N20410);
and AND4 (N20413, N20409, N19304, N16314, N10173);
xor XOR2 (N20414, N20371, N18439);
or OR4 (N20415, N20411, N16801, N2042, N14286);
nand NAND3 (N20416, N20415, N2351, N1427);
nor NOR4 (N20417, N20414, N11885, N2097, N19286);
xor XOR2 (N20418, N20406, N858);
nand NAND3 (N20419, N20403, N13281, N12046);
not NOT1 (N20420, N20412);
or OR2 (N20421, N20419, N4641);
not NOT1 (N20422, N20417);
not NOT1 (N20423, N20399);
nand NAND4 (N20424, N20416, N4684, N9428, N12591);
buf BUF1 (N20425, N20405);
xor XOR2 (N20426, N20421, N17934);
nand NAND2 (N20427, N20418, N18086);
nand NAND4 (N20428, N20420, N7388, N44, N12837);
and AND2 (N20429, N20394, N2375);
buf BUF1 (N20430, N20424);
not NOT1 (N20431, N20427);
buf BUF1 (N20432, N20429);
not NOT1 (N20433, N20423);
nand NAND3 (N20434, N20430, N16842, N10476);
nand NAND2 (N20435, N20428, N13197);
nand NAND3 (N20436, N20435, N8158, N5314);
xor XOR2 (N20437, N20422, N11927);
nand NAND3 (N20438, N20437, N14504, N6471);
and AND4 (N20439, N20432, N8378, N1526, N8536);
not NOT1 (N20440, N20425);
not NOT1 (N20441, N20439);
and AND2 (N20442, N20407, N16281);
not NOT1 (N20443, N20413);
not NOT1 (N20444, N20440);
nor NOR2 (N20445, N20443, N14448);
xor XOR2 (N20446, N20434, N16109);
buf BUF1 (N20447, N20426);
xor XOR2 (N20448, N20442, N18489);
or OR3 (N20449, N20447, N13836, N463);
buf BUF1 (N20450, N20448);
nand NAND3 (N20451, N20449, N8809, N15338);
xor XOR2 (N20452, N20433, N5258);
or OR4 (N20453, N20450, N1294, N16630, N3984);
xor XOR2 (N20454, N20452, N11220);
xor XOR2 (N20455, N20441, N19038);
and AND3 (N20456, N20446, N14885, N4016);
nor NOR3 (N20457, N20451, N16110, N16089);
nor NOR3 (N20458, N20457, N3962, N16229);
not NOT1 (N20459, N20455);
and AND2 (N20460, N20458, N18746);
xor XOR2 (N20461, N20444, N18649);
nor NOR2 (N20462, N20461, N18423);
or OR4 (N20463, N20436, N7351, N6344, N18571);
buf BUF1 (N20464, N20459);
not NOT1 (N20465, N20454);
not NOT1 (N20466, N20431);
or OR4 (N20467, N20464, N20263, N20289, N8826);
nor NOR3 (N20468, N20466, N9086, N12085);
nor NOR3 (N20469, N20467, N4130, N10837);
or OR2 (N20470, N20465, N15098);
not NOT1 (N20471, N20460);
nor NOR4 (N20472, N20438, N18471, N4727, N13631);
nor NOR4 (N20473, N20469, N2932, N4966, N12849);
and AND3 (N20474, N20462, N15987, N13411);
buf BUF1 (N20475, N20472);
xor XOR2 (N20476, N20473, N18977);
or OR2 (N20477, N20453, N7142);
nor NOR2 (N20478, N20463, N13618);
xor XOR2 (N20479, N20478, N273);
and AND4 (N20480, N20476, N8487, N7994, N10131);
nor NOR4 (N20481, N20477, N14451, N327, N18701);
nor NOR4 (N20482, N20475, N11521, N2421, N1533);
xor XOR2 (N20483, N20481, N11166);
or OR2 (N20484, N20445, N11654);
buf BUF1 (N20485, N20479);
buf BUF1 (N20486, N20480);
nand NAND4 (N20487, N20484, N19454, N19116, N3649);
nor NOR2 (N20488, N20483, N18440);
and AND4 (N20489, N20468, N17591, N2122, N14719);
or OR4 (N20490, N20470, N12835, N11925, N17972);
and AND4 (N20491, N20482, N10377, N7623, N2547);
nand NAND2 (N20492, N20456, N5640);
xor XOR2 (N20493, N20488, N2802);
xor XOR2 (N20494, N20471, N14232);
nor NOR4 (N20495, N20490, N12001, N12080, N12096);
or OR2 (N20496, N20491, N19451);
buf BUF1 (N20497, N20487);
or OR3 (N20498, N20497, N11417, N9323);
xor XOR2 (N20499, N20496, N13260);
nand NAND3 (N20500, N20498, N15230, N5433);
nor NOR4 (N20501, N20474, N8033, N8637, N8187);
nor NOR4 (N20502, N20492, N3078, N12475, N9293);
and AND4 (N20503, N20500, N1356, N15280, N4772);
nor NOR4 (N20504, N20493, N14112, N9243, N15322);
nor NOR4 (N20505, N20495, N3426, N9904, N14567);
nor NOR3 (N20506, N20494, N10238, N5911);
not NOT1 (N20507, N20501);
nor NOR4 (N20508, N20486, N12426, N20166, N18972);
nor NOR3 (N20509, N20508, N9381, N5276);
not NOT1 (N20510, N20502);
nor NOR4 (N20511, N20503, N17327, N16658, N16970);
and AND4 (N20512, N20505, N11531, N13645, N337);
nor NOR4 (N20513, N20511, N4550, N6774, N345);
xor XOR2 (N20514, N20499, N4012);
nor NOR3 (N20515, N20485, N14698, N18168);
not NOT1 (N20516, N20515);
xor XOR2 (N20517, N20512, N15931);
buf BUF1 (N20518, N20514);
and AND4 (N20519, N20507, N8663, N6377, N9971);
xor XOR2 (N20520, N20517, N6145);
buf BUF1 (N20521, N20519);
buf BUF1 (N20522, N20506);
xor XOR2 (N20523, N20504, N5788);
or OR3 (N20524, N20521, N15962, N12259);
xor XOR2 (N20525, N20510, N17502);
or OR2 (N20526, N20489, N9868);
not NOT1 (N20527, N20523);
or OR3 (N20528, N20527, N643, N1580);
xor XOR2 (N20529, N20522, N10694);
or OR3 (N20530, N20526, N19184, N19637);
nor NOR4 (N20531, N20518, N4621, N4590, N17038);
nor NOR3 (N20532, N20528, N2820, N23);
nor NOR4 (N20533, N20524, N19829, N695, N5024);
not NOT1 (N20534, N20509);
or OR3 (N20535, N20532, N11595, N1157);
nor NOR4 (N20536, N20534, N2261, N8169, N8602);
xor XOR2 (N20537, N20530, N12055);
and AND4 (N20538, N20529, N8003, N15104, N4137);
xor XOR2 (N20539, N20535, N16476);
or OR2 (N20540, N20520, N4595);
not NOT1 (N20541, N20540);
nor NOR4 (N20542, N20541, N16267, N1068, N17817);
nand NAND3 (N20543, N20542, N19947, N6407);
or OR3 (N20544, N20516, N18044, N9268);
nand NAND2 (N20545, N20513, N10431);
and AND3 (N20546, N20536, N17096, N8388);
and AND2 (N20547, N20539, N16766);
not NOT1 (N20548, N20543);
xor XOR2 (N20549, N20525, N3081);
not NOT1 (N20550, N20546);
not NOT1 (N20551, N20547);
xor XOR2 (N20552, N20537, N4622);
not NOT1 (N20553, N20550);
or OR4 (N20554, N20548, N9186, N2234, N13984);
not NOT1 (N20555, N20544);
or OR3 (N20556, N20538, N4125, N15401);
nand NAND3 (N20557, N20531, N3550, N5614);
nor NOR3 (N20558, N20555, N6363, N870);
buf BUF1 (N20559, N20556);
and AND2 (N20560, N20551, N14707);
nand NAND4 (N20561, N20552, N15594, N11347, N7921);
nand NAND2 (N20562, N20561, N3148);
nor NOR2 (N20563, N20559, N334);
or OR2 (N20564, N20562, N6699);
not NOT1 (N20565, N20564);
nand NAND4 (N20566, N20549, N17996, N8700, N12287);
xor XOR2 (N20567, N20557, N8187);
nor NOR2 (N20568, N20565, N574);
not NOT1 (N20569, N20568);
buf BUF1 (N20570, N20554);
xor XOR2 (N20571, N20553, N5381);
or OR3 (N20572, N20567, N16759, N869);
not NOT1 (N20573, N20563);
nand NAND2 (N20574, N20571, N3165);
or OR4 (N20575, N20533, N11920, N2153, N6390);
buf BUF1 (N20576, N20545);
not NOT1 (N20577, N20575);
nand NAND3 (N20578, N20558, N425, N174);
or OR2 (N20579, N20573, N14202);
nor NOR2 (N20580, N20579, N18952);
buf BUF1 (N20581, N20560);
nor NOR3 (N20582, N20577, N14369, N7098);
xor XOR2 (N20583, N20569, N11265);
not NOT1 (N20584, N20570);
nor NOR4 (N20585, N20574, N176, N9239, N10799);
nor NOR2 (N20586, N20576, N10831);
or OR2 (N20587, N20585, N7198);
nor NOR2 (N20588, N20566, N20268);
buf BUF1 (N20589, N20583);
or OR4 (N20590, N20572, N12121, N20082, N9794);
or OR2 (N20591, N20584, N20362);
buf BUF1 (N20592, N20580);
nor NOR3 (N20593, N20578, N20147, N3502);
or OR3 (N20594, N20589, N4404, N5144);
buf BUF1 (N20595, N20592);
nor NOR4 (N20596, N20581, N12268, N16147, N4726);
xor XOR2 (N20597, N20593, N4032);
xor XOR2 (N20598, N20591, N11255);
nand NAND4 (N20599, N20597, N6065, N10829, N4673);
and AND4 (N20600, N20588, N5337, N11624, N11186);
nand NAND2 (N20601, N20598, N19820);
and AND2 (N20602, N20587, N6098);
and AND4 (N20603, N20600, N18250, N7118, N7917);
nand NAND3 (N20604, N20602, N935, N17696);
nor NOR3 (N20605, N20603, N19091, N16380);
xor XOR2 (N20606, N20594, N10052);
not NOT1 (N20607, N20599);
and AND4 (N20608, N20586, N18504, N7241, N16105);
and AND4 (N20609, N20608, N9367, N16357, N4310);
nor NOR4 (N20610, N20605, N20129, N2632, N1393);
buf BUF1 (N20611, N20604);
and AND2 (N20612, N20582, N16420);
buf BUF1 (N20613, N20612);
and AND3 (N20614, N20613, N11178, N3262);
xor XOR2 (N20615, N20614, N3799);
nor NOR3 (N20616, N20609, N3209, N5173);
not NOT1 (N20617, N20607);
nand NAND3 (N20618, N20616, N11996, N5567);
nand NAND4 (N20619, N20595, N4626, N4253, N3335);
xor XOR2 (N20620, N20618, N19263);
nor NOR4 (N20621, N20601, N12982, N20085, N7540);
nand NAND2 (N20622, N20610, N8383);
buf BUF1 (N20623, N20606);
and AND2 (N20624, N20590, N2488);
not NOT1 (N20625, N20617);
nor NOR2 (N20626, N20625, N96);
or OR3 (N20627, N20611, N20520, N11338);
and AND3 (N20628, N20622, N18485, N685);
buf BUF1 (N20629, N20624);
xor XOR2 (N20630, N20621, N745);
xor XOR2 (N20631, N20615, N12008);
and AND3 (N20632, N20627, N16861, N15189);
and AND4 (N20633, N20630, N17998, N3241, N10157);
xor XOR2 (N20634, N20619, N12905);
and AND3 (N20635, N20628, N15747, N11213);
nor NOR2 (N20636, N20633, N20314);
or OR4 (N20637, N20626, N6106, N7624, N4002);
nor NOR4 (N20638, N20623, N13885, N6334, N15362);
nor NOR2 (N20639, N20632, N18604);
nand NAND3 (N20640, N20636, N1056, N13329);
nor NOR2 (N20641, N20639, N12951);
or OR4 (N20642, N20635, N6824, N12790, N16233);
or OR3 (N20643, N20640, N14252, N14780);
not NOT1 (N20644, N20631);
nand NAND3 (N20645, N20642, N19574, N6952);
nor NOR4 (N20646, N20645, N3772, N7500, N12198);
or OR4 (N20647, N20620, N16720, N13079, N20440);
nor NOR4 (N20648, N20643, N10184, N6753, N3588);
xor XOR2 (N20649, N20644, N19322);
not NOT1 (N20650, N20647);
not NOT1 (N20651, N20648);
xor XOR2 (N20652, N20629, N9060);
nor NOR2 (N20653, N20638, N1346);
not NOT1 (N20654, N20651);
xor XOR2 (N20655, N20596, N5727);
nand NAND4 (N20656, N20637, N9856, N13774, N20355);
nand NAND3 (N20657, N20655, N19919, N1695);
not NOT1 (N20658, N20641);
or OR3 (N20659, N20652, N8222, N17440);
not NOT1 (N20660, N20650);
nand NAND3 (N20661, N20659, N19509, N9400);
nor NOR3 (N20662, N20653, N2361, N934);
not NOT1 (N20663, N20657);
xor XOR2 (N20664, N20634, N15482);
xor XOR2 (N20665, N20664, N9633);
or OR2 (N20666, N20649, N8834);
nor NOR2 (N20667, N20656, N7346);
or OR2 (N20668, N20662, N16657);
and AND3 (N20669, N20665, N8771, N8373);
or OR2 (N20670, N20658, N10078);
nor NOR2 (N20671, N20646, N9846);
nor NOR2 (N20672, N20661, N6797);
not NOT1 (N20673, N20654);
not NOT1 (N20674, N20667);
or OR2 (N20675, N20670, N20386);
buf BUF1 (N20676, N20674);
buf BUF1 (N20677, N20672);
or OR3 (N20678, N20660, N19968, N12202);
or OR2 (N20679, N20666, N5155);
and AND2 (N20680, N20663, N8496);
buf BUF1 (N20681, N20673);
buf BUF1 (N20682, N20675);
or OR4 (N20683, N20680, N13009, N16974, N3504);
not NOT1 (N20684, N20681);
and AND4 (N20685, N20676, N7240, N10373, N9626);
nor NOR3 (N20686, N20685, N12028, N18320);
xor XOR2 (N20687, N20671, N10145);
or OR4 (N20688, N20677, N17857, N6367, N16660);
and AND3 (N20689, N20678, N1352, N7502);
and AND3 (N20690, N20687, N500, N15242);
xor XOR2 (N20691, N20690, N6873);
or OR3 (N20692, N20684, N17674, N3989);
not NOT1 (N20693, N20668);
not NOT1 (N20694, N20689);
nor NOR3 (N20695, N20669, N234, N13125);
buf BUF1 (N20696, N20695);
nand NAND2 (N20697, N20693, N12224);
buf BUF1 (N20698, N20683);
nor NOR2 (N20699, N20694, N17719);
xor XOR2 (N20700, N20699, N659);
not NOT1 (N20701, N20700);
xor XOR2 (N20702, N20696, N10466);
not NOT1 (N20703, N20701);
or OR2 (N20704, N20703, N18759);
and AND4 (N20705, N20686, N17810, N15228, N19918);
xor XOR2 (N20706, N20698, N14394);
nor NOR4 (N20707, N20688, N1268, N14478, N7494);
nand NAND4 (N20708, N20691, N18670, N2501, N10813);
and AND4 (N20709, N20682, N14643, N15841, N9822);
xor XOR2 (N20710, N20705, N4374);
buf BUF1 (N20711, N20706);
buf BUF1 (N20712, N20702);
and AND2 (N20713, N20708, N6344);
xor XOR2 (N20714, N20710, N14666);
xor XOR2 (N20715, N20713, N17084);
nor NOR2 (N20716, N20697, N769);
nor NOR4 (N20717, N20715, N4588, N731, N19421);
xor XOR2 (N20718, N20679, N9075);
nor NOR3 (N20719, N20704, N11367, N2396);
nand NAND4 (N20720, N20711, N5720, N4931, N8891);
buf BUF1 (N20721, N20714);
nor NOR3 (N20722, N20720, N1608, N4482);
and AND2 (N20723, N20712, N17517);
nand NAND2 (N20724, N20721, N16873);
not NOT1 (N20725, N20707);
nand NAND3 (N20726, N20725, N16231, N13974);
nand NAND4 (N20727, N20716, N2120, N13083, N18919);
xor XOR2 (N20728, N20727, N13618);
buf BUF1 (N20729, N20718);
nand NAND4 (N20730, N20692, N15485, N16630, N18060);
not NOT1 (N20731, N20709);
buf BUF1 (N20732, N20726);
nand NAND4 (N20733, N20728, N4418, N18212, N39);
xor XOR2 (N20734, N20717, N6809);
not NOT1 (N20735, N20731);
nor NOR2 (N20736, N20722, N11826);
not NOT1 (N20737, N20724);
nand NAND3 (N20738, N20736, N13117, N10809);
not NOT1 (N20739, N20719);
or OR2 (N20740, N20738, N8748);
nand NAND2 (N20741, N20739, N18142);
xor XOR2 (N20742, N20729, N4525);
or OR3 (N20743, N20730, N6095, N11417);
buf BUF1 (N20744, N20741);
not NOT1 (N20745, N20733);
and AND2 (N20746, N20743, N7763);
not NOT1 (N20747, N20744);
not NOT1 (N20748, N20746);
nand NAND4 (N20749, N20732, N4032, N15161, N7476);
buf BUF1 (N20750, N20742);
nand NAND2 (N20751, N20749, N9385);
buf BUF1 (N20752, N20723);
xor XOR2 (N20753, N20740, N10481);
nor NOR2 (N20754, N20750, N13946);
and AND3 (N20755, N20753, N6434, N8393);
nand NAND2 (N20756, N20755, N5134);
xor XOR2 (N20757, N20754, N15920);
nor NOR4 (N20758, N20735, N9181, N5013, N12325);
xor XOR2 (N20759, N20758, N12938);
nand NAND3 (N20760, N20757, N13539, N14822);
and AND4 (N20761, N20751, N19804, N9679, N8565);
buf BUF1 (N20762, N20734);
not NOT1 (N20763, N20760);
nor NOR4 (N20764, N20761, N4962, N409, N1222);
buf BUF1 (N20765, N20748);
or OR2 (N20766, N20759, N9742);
buf BUF1 (N20767, N20765);
buf BUF1 (N20768, N20767);
nand NAND3 (N20769, N20768, N14159, N4102);
xor XOR2 (N20770, N20766, N9151);
nand NAND4 (N20771, N20752, N8658, N9383, N1450);
and AND3 (N20772, N20763, N1151, N14922);
or OR2 (N20773, N20747, N20194);
xor XOR2 (N20774, N20764, N9950);
or OR2 (N20775, N20774, N633);
and AND4 (N20776, N20769, N8060, N11636, N17889);
buf BUF1 (N20777, N20745);
xor XOR2 (N20778, N20772, N2897);
nand NAND4 (N20779, N20771, N14991, N3306, N13615);
nor NOR2 (N20780, N20775, N1044);
nor NOR3 (N20781, N20779, N12205, N13535);
nor NOR4 (N20782, N20777, N13725, N11872, N3869);
nand NAND2 (N20783, N20781, N13382);
xor XOR2 (N20784, N20782, N6052);
not NOT1 (N20785, N20737);
buf BUF1 (N20786, N20783);
not NOT1 (N20787, N20762);
or OR3 (N20788, N20776, N8367, N9615);
nor NOR2 (N20789, N20756, N5092);
nor NOR3 (N20790, N20785, N6893, N11733);
nor NOR4 (N20791, N20789, N14710, N6830, N8658);
not NOT1 (N20792, N20787);
or OR4 (N20793, N20792, N8423, N7083, N14662);
nand NAND2 (N20794, N20780, N3868);
or OR4 (N20795, N20770, N3681, N2767, N5683);
nor NOR2 (N20796, N20795, N394);
nor NOR3 (N20797, N20778, N17885, N4269);
nand NAND3 (N20798, N20791, N10109, N18898);
buf BUF1 (N20799, N20797);
and AND3 (N20800, N20796, N2143, N2727);
buf BUF1 (N20801, N20773);
nand NAND2 (N20802, N20794, N16498);
nand NAND2 (N20803, N20798, N11909);
xor XOR2 (N20804, N20800, N17260);
nand NAND3 (N20805, N20788, N10706, N10821);
xor XOR2 (N20806, N20784, N8618);
buf BUF1 (N20807, N20804);
or OR3 (N20808, N20786, N18201, N1633);
nand NAND4 (N20809, N20801, N12279, N8129, N12554);
xor XOR2 (N20810, N20809, N6665);
nor NOR3 (N20811, N20808, N19656, N18438);
and AND4 (N20812, N20807, N10830, N15589, N6513);
nor NOR2 (N20813, N20810, N4875);
xor XOR2 (N20814, N20811, N12660);
and AND4 (N20815, N20802, N5152, N13113, N20529);
and AND3 (N20816, N20806, N4093, N10903);
xor XOR2 (N20817, N20812, N50);
xor XOR2 (N20818, N20815, N8562);
not NOT1 (N20819, N20799);
not NOT1 (N20820, N20803);
not NOT1 (N20821, N20793);
nand NAND3 (N20822, N20805, N5656, N10270);
or OR3 (N20823, N20817, N15217, N9044);
nor NOR3 (N20824, N20819, N1862, N20436);
xor XOR2 (N20825, N20820, N17260);
nand NAND2 (N20826, N20818, N12399);
xor XOR2 (N20827, N20822, N8927);
and AND3 (N20828, N20814, N2961, N262);
nor NOR4 (N20829, N20816, N7632, N6366, N20706);
and AND3 (N20830, N20827, N14796, N9133);
and AND2 (N20831, N20821, N4228);
and AND4 (N20832, N20831, N17669, N5968, N4873);
xor XOR2 (N20833, N20832, N13209);
xor XOR2 (N20834, N20813, N11744);
not NOT1 (N20835, N20790);
nand NAND2 (N20836, N20829, N11188);
or OR2 (N20837, N20836, N11366);
not NOT1 (N20838, N20834);
not NOT1 (N20839, N20838);
xor XOR2 (N20840, N20830, N15554);
or OR4 (N20841, N20824, N301, N2811, N8542);
not NOT1 (N20842, N20840);
and AND2 (N20843, N20823, N9577);
and AND2 (N20844, N20841, N15836);
not NOT1 (N20845, N20833);
and AND2 (N20846, N20843, N17994);
xor XOR2 (N20847, N20842, N16110);
xor XOR2 (N20848, N20839, N7515);
or OR3 (N20849, N20846, N15164, N11786);
and AND3 (N20850, N20835, N17544, N19837);
or OR4 (N20851, N20826, N2861, N9260, N10451);
or OR4 (N20852, N20848, N4321, N639, N5129);
not NOT1 (N20853, N20851);
buf BUF1 (N20854, N20853);
xor XOR2 (N20855, N20837, N18158);
not NOT1 (N20856, N20828);
and AND3 (N20857, N20852, N5620, N17745);
xor XOR2 (N20858, N20857, N16743);
nand NAND2 (N20859, N20854, N6578);
xor XOR2 (N20860, N20844, N5837);
nand NAND2 (N20861, N20856, N20583);
or OR3 (N20862, N20825, N9012, N10273);
or OR4 (N20863, N20862, N8529, N19226, N17073);
nor NOR2 (N20864, N20850, N9380);
nand NAND2 (N20865, N20845, N11189);
nand NAND2 (N20866, N20865, N19001);
nor NOR3 (N20867, N20847, N20358, N16128);
nor NOR2 (N20868, N20864, N18260);
and AND3 (N20869, N20849, N7736, N5392);
xor XOR2 (N20870, N20861, N6482);
nand NAND4 (N20871, N20867, N10645, N15498, N3863);
not NOT1 (N20872, N20866);
buf BUF1 (N20873, N20870);
nor NOR3 (N20874, N20869, N9509, N12580);
and AND2 (N20875, N20872, N3999);
and AND2 (N20876, N20871, N11703);
buf BUF1 (N20877, N20860);
buf BUF1 (N20878, N20855);
or OR3 (N20879, N20875, N12445, N5099);
nand NAND3 (N20880, N20878, N2442, N18307);
nor NOR2 (N20881, N20858, N14098);
not NOT1 (N20882, N20879);
not NOT1 (N20883, N20876);
xor XOR2 (N20884, N20877, N1119);
nand NAND2 (N20885, N20868, N17671);
xor XOR2 (N20886, N20883, N11173);
or OR3 (N20887, N20873, N14490, N17732);
nand NAND2 (N20888, N20882, N1077);
and AND4 (N20889, N20886, N18559, N9753, N4504);
not NOT1 (N20890, N20874);
xor XOR2 (N20891, N20888, N19263);
nand NAND2 (N20892, N20889, N15438);
nor NOR4 (N20893, N20859, N6589, N12797, N5186);
or OR4 (N20894, N20863, N1642, N7515, N11672);
and AND3 (N20895, N20893, N15066, N17276);
not NOT1 (N20896, N20887);
xor XOR2 (N20897, N20892, N10881);
nor NOR3 (N20898, N20895, N18032, N11059);
buf BUF1 (N20899, N20881);
nand NAND2 (N20900, N20898, N11501);
or OR4 (N20901, N20885, N8490, N16201, N19686);
buf BUF1 (N20902, N20901);
and AND2 (N20903, N20897, N8068);
xor XOR2 (N20904, N20891, N19246);
and AND2 (N20905, N20896, N2860);
not NOT1 (N20906, N20890);
or OR4 (N20907, N20894, N15139, N9226, N18423);
xor XOR2 (N20908, N20902, N20405);
or OR2 (N20909, N20884, N12410);
buf BUF1 (N20910, N20900);
xor XOR2 (N20911, N20908, N16279);
buf BUF1 (N20912, N20907);
or OR4 (N20913, N20880, N1584, N15818, N10882);
and AND4 (N20914, N20910, N4184, N2758, N14413);
or OR4 (N20915, N20906, N10092, N14530, N14332);
buf BUF1 (N20916, N20909);
buf BUF1 (N20917, N20914);
buf BUF1 (N20918, N20903);
not NOT1 (N20919, N20915);
and AND4 (N20920, N20911, N3196, N13526, N6401);
or OR3 (N20921, N20920, N18844, N6341);
and AND3 (N20922, N20899, N13905, N2563);
xor XOR2 (N20923, N20921, N15640);
buf BUF1 (N20924, N20919);
or OR2 (N20925, N20917, N20376);
not NOT1 (N20926, N20922);
xor XOR2 (N20927, N20905, N6302);
nor NOR3 (N20928, N20926, N13450, N5566);
not NOT1 (N20929, N20913);
nor NOR4 (N20930, N20924, N17693, N6044, N12115);
xor XOR2 (N20931, N20918, N3418);
xor XOR2 (N20932, N20931, N1755);
nand NAND2 (N20933, N20904, N14241);
nor NOR2 (N20934, N20912, N18205);
xor XOR2 (N20935, N20933, N9970);
nand NAND3 (N20936, N20934, N13352, N7566);
buf BUF1 (N20937, N20916);
nand NAND3 (N20938, N20936, N19100, N4419);
or OR2 (N20939, N20923, N5889);
nand NAND2 (N20940, N20925, N4061);
and AND3 (N20941, N20940, N11627, N12157);
xor XOR2 (N20942, N20937, N8529);
nand NAND2 (N20943, N20927, N6395);
or OR3 (N20944, N20941, N18465, N8806);
buf BUF1 (N20945, N20930);
not NOT1 (N20946, N20938);
not NOT1 (N20947, N20946);
nand NAND3 (N20948, N20928, N2324, N2730);
nor NOR2 (N20949, N20942, N4093);
not NOT1 (N20950, N20949);
not NOT1 (N20951, N20939);
buf BUF1 (N20952, N20935);
or OR2 (N20953, N20945, N9361);
and AND4 (N20954, N20953, N19589, N16113, N8552);
and AND4 (N20955, N20944, N15118, N15278, N17986);
nand NAND2 (N20956, N20950, N14517);
not NOT1 (N20957, N20932);
not NOT1 (N20958, N20948);
nand NAND4 (N20959, N20929, N14305, N12855, N4400);
nor NOR3 (N20960, N20943, N15019, N14801);
buf BUF1 (N20961, N20952);
not NOT1 (N20962, N20958);
nor NOR2 (N20963, N20960, N7124);
and AND4 (N20964, N20957, N13091, N19787, N10485);
not NOT1 (N20965, N20961);
or OR2 (N20966, N20956, N10440);
and AND2 (N20967, N20964, N13652);
nand NAND4 (N20968, N20951, N19602, N861, N3761);
or OR2 (N20969, N20962, N6635);
buf BUF1 (N20970, N20967);
xor XOR2 (N20971, N20954, N11158);
nor NOR3 (N20972, N20969, N5073, N16254);
xor XOR2 (N20973, N20971, N11266);
or OR2 (N20974, N20973, N3808);
or OR4 (N20975, N20970, N10661, N13814, N6948);
buf BUF1 (N20976, N20947);
not NOT1 (N20977, N20966);
buf BUF1 (N20978, N20972);
buf BUF1 (N20979, N20955);
or OR4 (N20980, N20978, N20378, N1600, N18724);
nand NAND2 (N20981, N20968, N15535);
nand NAND2 (N20982, N20959, N4058);
buf BUF1 (N20983, N20979);
nor NOR3 (N20984, N20974, N5856, N10766);
and AND2 (N20985, N20983, N3159);
xor XOR2 (N20986, N20982, N19360);
and AND4 (N20987, N20975, N11353, N5181, N3179);
not NOT1 (N20988, N20981);
xor XOR2 (N20989, N20965, N14753);
buf BUF1 (N20990, N20980);
and AND3 (N20991, N20985, N5193, N3419);
and AND2 (N20992, N20984, N3346);
xor XOR2 (N20993, N20977, N17969);
or OR3 (N20994, N20963, N9634, N14725);
and AND4 (N20995, N20987, N16145, N13174, N8220);
nand NAND4 (N20996, N20976, N5098, N13192, N18300);
xor XOR2 (N20997, N20993, N6441);
or OR2 (N20998, N20992, N568);
and AND3 (N20999, N20994, N2879, N9487);
nand NAND3 (N21000, N20997, N4172, N3371);
buf BUF1 (N21001, N21000);
not NOT1 (N21002, N20998);
nor NOR4 (N21003, N20989, N13767, N6973, N165);
or OR4 (N21004, N20995, N14374, N13081, N19846);
not NOT1 (N21005, N20991);
nor NOR2 (N21006, N21001, N13063);
or OR4 (N21007, N21004, N3144, N6916, N20647);
buf BUF1 (N21008, N20999);
buf BUF1 (N21009, N21007);
not NOT1 (N21010, N21006);
buf BUF1 (N21011, N21005);
buf BUF1 (N21012, N20996);
or OR3 (N21013, N21010, N18060, N19018);
and AND3 (N21014, N20990, N4789, N20642);
not NOT1 (N21015, N21011);
or OR4 (N21016, N21014, N10176, N19877, N18463);
and AND4 (N21017, N21013, N20077, N20842, N2738);
or OR2 (N21018, N21008, N9033);
xor XOR2 (N21019, N21002, N12254);
nor NOR3 (N21020, N21016, N4320, N14820);
nor NOR4 (N21021, N21012, N11651, N2075, N1266);
buf BUF1 (N21022, N21003);
nand NAND2 (N21023, N21015, N12524);
and AND4 (N21024, N21017, N17855, N6818, N15464);
not NOT1 (N21025, N20988);
and AND4 (N21026, N21021, N20412, N13855, N6626);
nor NOR2 (N21027, N21023, N11230);
and AND3 (N21028, N21027, N12007, N15938);
xor XOR2 (N21029, N21018, N13620);
and AND4 (N21030, N21022, N2741, N2987, N13051);
buf BUF1 (N21031, N21028);
and AND2 (N21032, N21026, N3669);
not NOT1 (N21033, N21009);
nor NOR3 (N21034, N21030, N13598, N732);
or OR2 (N21035, N21029, N981);
or OR3 (N21036, N21031, N3898, N5766);
nand NAND3 (N21037, N21035, N3476, N20705);
buf BUF1 (N21038, N21020);
buf BUF1 (N21039, N21033);
not NOT1 (N21040, N21032);
xor XOR2 (N21041, N21040, N8810);
and AND3 (N21042, N21025, N290, N14324);
nand NAND3 (N21043, N21036, N10954, N2790);
or OR2 (N21044, N21024, N18473);
xor XOR2 (N21045, N21041, N16406);
nor NOR3 (N21046, N21039, N13384, N7008);
buf BUF1 (N21047, N21045);
xor XOR2 (N21048, N20986, N16774);
or OR4 (N21049, N21042, N19708, N8779, N10969);
buf BUF1 (N21050, N21048);
nor NOR2 (N21051, N21019, N2749);
and AND4 (N21052, N21050, N11982, N4997, N1536);
buf BUF1 (N21053, N21037);
nor NOR2 (N21054, N21051, N13306);
buf BUF1 (N21055, N21047);
and AND2 (N21056, N21055, N5980);
buf BUF1 (N21057, N21056);
and AND4 (N21058, N21053, N1540, N5453, N18978);
buf BUF1 (N21059, N21049);
nor NOR3 (N21060, N21058, N8666, N5699);
xor XOR2 (N21061, N21057, N7120);
and AND3 (N21062, N21059, N16074, N16850);
nor NOR2 (N21063, N21038, N19598);
not NOT1 (N21064, N21052);
buf BUF1 (N21065, N21062);
xor XOR2 (N21066, N21060, N7941);
or OR2 (N21067, N21061, N17534);
and AND4 (N21068, N21067, N13272, N10591, N20897);
and AND2 (N21069, N21065, N9117);
buf BUF1 (N21070, N21054);
not NOT1 (N21071, N21043);
xor XOR2 (N21072, N21069, N19974);
xor XOR2 (N21073, N21068, N19197);
buf BUF1 (N21074, N21063);
buf BUF1 (N21075, N21034);
buf BUF1 (N21076, N21074);
xor XOR2 (N21077, N21044, N316);
not NOT1 (N21078, N21064);
nand NAND2 (N21079, N21072, N10559);
nor NOR4 (N21080, N21046, N4767, N6658, N8981);
and AND2 (N21081, N21077, N17340);
or OR3 (N21082, N21071, N11189, N11168);
nand NAND3 (N21083, N21076, N2448, N2884);
nand NAND2 (N21084, N21073, N4943);
or OR4 (N21085, N21082, N10606, N8260, N2236);
nor NOR2 (N21086, N21080, N10507);
not NOT1 (N21087, N21070);
or OR4 (N21088, N21083, N5024, N11598, N11107);
or OR4 (N21089, N21086, N14449, N5360, N7840);
not NOT1 (N21090, N21079);
buf BUF1 (N21091, N21088);
xor XOR2 (N21092, N21066, N20218);
buf BUF1 (N21093, N21085);
and AND2 (N21094, N21093, N20840);
xor XOR2 (N21095, N21094, N19414);
not NOT1 (N21096, N21092);
buf BUF1 (N21097, N21090);
nand NAND2 (N21098, N21075, N9418);
nor NOR2 (N21099, N21087, N6548);
or OR2 (N21100, N21078, N834);
or OR2 (N21101, N21095, N19010);
and AND2 (N21102, N21091, N9341);
buf BUF1 (N21103, N21101);
xor XOR2 (N21104, N21097, N13302);
nand NAND2 (N21105, N21084, N11675);
not NOT1 (N21106, N21089);
not NOT1 (N21107, N21100);
nor NOR3 (N21108, N21104, N9588, N13873);
xor XOR2 (N21109, N21106, N16474);
nor NOR2 (N21110, N21103, N15640);
xor XOR2 (N21111, N21105, N1295);
and AND2 (N21112, N21109, N3641);
and AND4 (N21113, N21107, N11327, N106, N19438);
not NOT1 (N21114, N21096);
and AND3 (N21115, N21108, N16854, N2694);
nand NAND2 (N21116, N21112, N2484);
nor NOR2 (N21117, N21116, N9166);
or OR3 (N21118, N21099, N8394, N20022);
and AND2 (N21119, N21117, N13426);
not NOT1 (N21120, N21110);
xor XOR2 (N21121, N21115, N11346);
xor XOR2 (N21122, N21102, N11698);
nand NAND3 (N21123, N21121, N20456, N17388);
and AND2 (N21124, N21081, N13778);
or OR3 (N21125, N21120, N6275, N8788);
not NOT1 (N21126, N21122);
and AND2 (N21127, N21125, N18164);
and AND4 (N21128, N21126, N19982, N17958, N4102);
not NOT1 (N21129, N21111);
not NOT1 (N21130, N21118);
buf BUF1 (N21131, N21123);
nand NAND2 (N21132, N21128, N14972);
buf BUF1 (N21133, N21129);
not NOT1 (N21134, N21132);
and AND2 (N21135, N21133, N2351);
or OR2 (N21136, N21134, N260);
nand NAND2 (N21137, N21136, N7274);
nor NOR3 (N21138, N21113, N8016, N16343);
nand NAND4 (N21139, N21135, N18675, N17614, N3613);
nor NOR4 (N21140, N21119, N14113, N2503, N7891);
xor XOR2 (N21141, N21137, N16263);
and AND4 (N21142, N21140, N10402, N15197, N10472);
or OR2 (N21143, N21139, N14595);
nand NAND2 (N21144, N21127, N6539);
buf BUF1 (N21145, N21141);
or OR3 (N21146, N21143, N14139, N9225);
or OR2 (N21147, N21138, N5158);
xor XOR2 (N21148, N21098, N9986);
not NOT1 (N21149, N21142);
xor XOR2 (N21150, N21148, N8996);
not NOT1 (N21151, N21146);
xor XOR2 (N21152, N21145, N4590);
buf BUF1 (N21153, N21149);
or OR2 (N21154, N21150, N19183);
or OR3 (N21155, N21131, N15804, N17292);
nor NOR3 (N21156, N21147, N8777, N20801);
nand NAND3 (N21157, N21156, N9608, N11178);
or OR3 (N21158, N21124, N487, N1808);
xor XOR2 (N21159, N21151, N3612);
or OR4 (N21160, N21155, N13666, N12111, N4300);
buf BUF1 (N21161, N21152);
nand NAND2 (N21162, N21160, N14031);
nand NAND4 (N21163, N21161, N9318, N9922, N16824);
xor XOR2 (N21164, N21157, N10090);
nor NOR3 (N21165, N21114, N15780, N800);
and AND4 (N21166, N21163, N19026, N18137, N12787);
xor XOR2 (N21167, N21166, N16191);
nor NOR4 (N21168, N21162, N6600, N10046, N14786);
or OR2 (N21169, N21164, N16997);
and AND4 (N21170, N21154, N19062, N13861, N16565);
or OR2 (N21171, N21144, N9604);
xor XOR2 (N21172, N21158, N16740);
buf BUF1 (N21173, N21169);
not NOT1 (N21174, N21172);
and AND4 (N21175, N21167, N9183, N6517, N17416);
nor NOR3 (N21176, N21173, N16132, N2679);
and AND2 (N21177, N21153, N3572);
xor XOR2 (N21178, N21159, N16769);
xor XOR2 (N21179, N21170, N12094);
or OR2 (N21180, N21178, N14492);
xor XOR2 (N21181, N21175, N8916);
xor XOR2 (N21182, N21176, N12552);
nand NAND2 (N21183, N21168, N12846);
xor XOR2 (N21184, N21130, N21056);
xor XOR2 (N21185, N21180, N3897);
not NOT1 (N21186, N21171);
nand NAND4 (N21187, N21182, N14467, N7353, N2109);
or OR4 (N21188, N21179, N18579, N19378, N14670);
nor NOR3 (N21189, N21183, N14374, N7517);
or OR2 (N21190, N21189, N16616);
not NOT1 (N21191, N21177);
buf BUF1 (N21192, N21185);
buf BUF1 (N21193, N21192);
nand NAND3 (N21194, N21187, N18012, N383);
not NOT1 (N21195, N21190);
xor XOR2 (N21196, N21184, N18267);
and AND2 (N21197, N21165, N323);
and AND4 (N21198, N21197, N6837, N282, N13757);
or OR3 (N21199, N21198, N9320, N239);
xor XOR2 (N21200, N21186, N13254);
and AND4 (N21201, N21195, N5556, N3881, N12472);
and AND3 (N21202, N21188, N4667, N17832);
and AND4 (N21203, N21191, N17844, N2080, N13787);
nand NAND3 (N21204, N21202, N14389, N389);
or OR2 (N21205, N21196, N18347);
buf BUF1 (N21206, N21201);
nand NAND4 (N21207, N21174, N5524, N20970, N10702);
or OR2 (N21208, N21199, N1298);
xor XOR2 (N21209, N21206, N17254);
not NOT1 (N21210, N21205);
nand NAND3 (N21211, N21181, N3442, N17555);
or OR4 (N21212, N21211, N10436, N11291, N8867);
not NOT1 (N21213, N21210);
nor NOR3 (N21214, N21213, N12270, N17813);
buf BUF1 (N21215, N21204);
nor NOR2 (N21216, N21208, N16371);
not NOT1 (N21217, N21193);
and AND4 (N21218, N21215, N1931, N12415, N11840);
xor XOR2 (N21219, N21212, N21003);
buf BUF1 (N21220, N21200);
or OR4 (N21221, N21218, N8010, N15014, N16111);
or OR4 (N21222, N21220, N4860, N4758, N17692);
and AND2 (N21223, N21203, N14000);
or OR2 (N21224, N21221, N3479);
not NOT1 (N21225, N21214);
and AND3 (N21226, N21224, N6128, N17129);
buf BUF1 (N21227, N21209);
nand NAND3 (N21228, N21222, N7255, N9280);
or OR2 (N21229, N21194, N20649);
buf BUF1 (N21230, N21227);
xor XOR2 (N21231, N21229, N19107);
nor NOR3 (N21232, N21219, N11396, N18832);
and AND2 (N21233, N21225, N17570);
xor XOR2 (N21234, N21223, N869);
and AND2 (N21235, N21216, N9157);
buf BUF1 (N21236, N21232);
and AND3 (N21237, N21231, N8540, N6567);
or OR3 (N21238, N21233, N5360, N16994);
nand NAND4 (N21239, N21234, N6675, N1421, N19802);
and AND2 (N21240, N21226, N1832);
xor XOR2 (N21241, N21235, N12357);
buf BUF1 (N21242, N21241);
or OR3 (N21243, N21237, N18577, N9437);
xor XOR2 (N21244, N21243, N19679);
or OR3 (N21245, N21240, N21209, N3584);
not NOT1 (N21246, N21236);
or OR4 (N21247, N21228, N12474, N15987, N19238);
and AND2 (N21248, N21217, N13713);
not NOT1 (N21249, N21245);
not NOT1 (N21250, N21207);
or OR2 (N21251, N21239, N10028);
buf BUF1 (N21252, N21238);
not NOT1 (N21253, N21247);
buf BUF1 (N21254, N21246);
nor NOR2 (N21255, N21253, N6140);
or OR3 (N21256, N21251, N16354, N8749);
xor XOR2 (N21257, N21230, N19270);
nand NAND2 (N21258, N21250, N9182);
and AND4 (N21259, N21242, N20610, N19751, N18682);
nand NAND4 (N21260, N21259, N5368, N14356, N10916);
nand NAND2 (N21261, N21244, N9807);
buf BUF1 (N21262, N21261);
xor XOR2 (N21263, N21254, N13414);
xor XOR2 (N21264, N21249, N19698);
buf BUF1 (N21265, N21260);
nor NOR4 (N21266, N21255, N19736, N20094, N8941);
not NOT1 (N21267, N21263);
nand NAND2 (N21268, N21262, N7353);
xor XOR2 (N21269, N21248, N14424);
nand NAND2 (N21270, N21267, N14218);
nand NAND2 (N21271, N21265, N8471);
xor XOR2 (N21272, N21270, N20033);
nand NAND3 (N21273, N21264, N16249, N4309);
or OR3 (N21274, N21271, N7884, N652);
buf BUF1 (N21275, N21252);
nand NAND3 (N21276, N21274, N7991, N19969);
buf BUF1 (N21277, N21256);
or OR3 (N21278, N21258, N17337, N19223);
not NOT1 (N21279, N21278);
not NOT1 (N21280, N21272);
and AND4 (N21281, N21273, N13272, N4600, N7244);
nor NOR2 (N21282, N21268, N3746);
nor NOR4 (N21283, N21266, N4477, N5476, N11778);
not NOT1 (N21284, N21257);
or OR2 (N21285, N21277, N1038);
and AND3 (N21286, N21279, N11638, N11756);
not NOT1 (N21287, N21281);
buf BUF1 (N21288, N21286);
buf BUF1 (N21289, N21284);
nand NAND3 (N21290, N21275, N14547, N19547);
not NOT1 (N21291, N21288);
xor XOR2 (N21292, N21282, N783);
or OR4 (N21293, N21290, N7565, N4770, N1498);
buf BUF1 (N21294, N21287);
nor NOR4 (N21295, N21285, N795, N5514, N15345);
buf BUF1 (N21296, N21292);
nand NAND3 (N21297, N21289, N12046, N4439);
and AND2 (N21298, N21291, N4758);
xor XOR2 (N21299, N21298, N5804);
and AND4 (N21300, N21276, N14588, N5201, N11398);
not NOT1 (N21301, N21293);
xor XOR2 (N21302, N21301, N8537);
and AND3 (N21303, N21295, N1159, N1474);
not NOT1 (N21304, N21302);
and AND4 (N21305, N21304, N15639, N13972, N13701);
nor NOR2 (N21306, N21297, N7486);
nand NAND2 (N21307, N21280, N2297);
buf BUF1 (N21308, N21305);
buf BUF1 (N21309, N21269);
nor NOR4 (N21310, N21308, N11264, N10502, N15852);
nand NAND4 (N21311, N21307, N19796, N21042, N7853);
xor XOR2 (N21312, N21309, N12813);
buf BUF1 (N21313, N21283);
xor XOR2 (N21314, N21311, N382);
buf BUF1 (N21315, N21306);
nor NOR2 (N21316, N21314, N4042);
buf BUF1 (N21317, N21296);
xor XOR2 (N21318, N21299, N14933);
nor NOR3 (N21319, N21300, N15323, N640);
xor XOR2 (N21320, N21312, N10112);
not NOT1 (N21321, N21319);
or OR3 (N21322, N21294, N4818, N4258);
not NOT1 (N21323, N21321);
nor NOR3 (N21324, N21303, N17724, N16455);
nor NOR3 (N21325, N21322, N13173, N894);
buf BUF1 (N21326, N21324);
nor NOR4 (N21327, N21318, N10890, N16355, N16351);
and AND2 (N21328, N21310, N18526);
or OR3 (N21329, N21313, N1152, N565);
nor NOR4 (N21330, N21317, N20262, N20172, N12103);
buf BUF1 (N21331, N21316);
and AND3 (N21332, N21315, N2661, N6381);
nand NAND3 (N21333, N21329, N21303, N20884);
or OR2 (N21334, N21325, N20232);
or OR3 (N21335, N21320, N8887, N14141);
nand NAND4 (N21336, N21331, N17527, N18285, N18471);
nor NOR4 (N21337, N21336, N15171, N7909, N3081);
nor NOR4 (N21338, N21335, N5832, N5240, N17919);
nor NOR2 (N21339, N21328, N15714);
xor XOR2 (N21340, N21327, N20444);
xor XOR2 (N21341, N21340, N11981);
not NOT1 (N21342, N21334);
nand NAND3 (N21343, N21323, N13487, N1876);
xor XOR2 (N21344, N21332, N8481);
or OR3 (N21345, N21341, N1958, N6465);
xor XOR2 (N21346, N21326, N15924);
not NOT1 (N21347, N21345);
nor NOR4 (N21348, N21338, N10290, N13414, N14823);
buf BUF1 (N21349, N21339);
buf BUF1 (N21350, N21349);
xor XOR2 (N21351, N21344, N17816);
xor XOR2 (N21352, N21351, N12709);
nor NOR2 (N21353, N21337, N4400);
nor NOR2 (N21354, N21343, N15642);
nor NOR2 (N21355, N21333, N11469);
buf BUF1 (N21356, N21352);
or OR3 (N21357, N21355, N710, N9557);
or OR2 (N21358, N21354, N21207);
or OR4 (N21359, N21350, N6476, N17562, N15494);
and AND2 (N21360, N21347, N1800);
buf BUF1 (N21361, N21348);
nand NAND3 (N21362, N21358, N12060, N13351);
xor XOR2 (N21363, N21342, N7565);
xor XOR2 (N21364, N21353, N18571);
nor NOR3 (N21365, N21363, N2570, N19474);
nor NOR3 (N21366, N21362, N17359, N1338);
and AND3 (N21367, N21360, N17201, N4749);
or OR2 (N21368, N21366, N5698);
xor XOR2 (N21369, N21365, N9831);
not NOT1 (N21370, N21369);
buf BUF1 (N21371, N21367);
nor NOR2 (N21372, N21357, N14327);
and AND4 (N21373, N21368, N1636, N5288, N2723);
xor XOR2 (N21374, N21361, N4932);
not NOT1 (N21375, N21364);
or OR3 (N21376, N21346, N4392, N2674);
and AND4 (N21377, N21330, N13246, N14539, N18353);
and AND4 (N21378, N21373, N293, N3053, N17938);
and AND3 (N21379, N21372, N15201, N3763);
xor XOR2 (N21380, N21375, N13736);
nor NOR3 (N21381, N21377, N1771, N18156);
and AND3 (N21382, N21370, N13922, N807);
xor XOR2 (N21383, N21371, N13662);
not NOT1 (N21384, N21359);
nand NAND3 (N21385, N21356, N15057, N18881);
nand NAND4 (N21386, N21384, N17592, N12081, N18394);
or OR2 (N21387, N21378, N11077);
nor NOR4 (N21388, N21382, N11387, N3180, N16959);
not NOT1 (N21389, N21380);
nand NAND4 (N21390, N21387, N3814, N3476, N16588);
xor XOR2 (N21391, N21381, N20892);
nor NOR3 (N21392, N21379, N12216, N13482);
not NOT1 (N21393, N21386);
buf BUF1 (N21394, N21385);
nand NAND2 (N21395, N21389, N8125);
and AND3 (N21396, N21388, N10962, N7149);
or OR4 (N21397, N21396, N14131, N7670, N1631);
buf BUF1 (N21398, N21392);
nand NAND2 (N21399, N21394, N15301);
xor XOR2 (N21400, N21390, N19711);
not NOT1 (N21401, N21399);
nand NAND4 (N21402, N21398, N1757, N11791, N9007);
nor NOR4 (N21403, N21374, N15577, N3909, N9625);
xor XOR2 (N21404, N21383, N15903);
xor XOR2 (N21405, N21376, N6624);
nor NOR2 (N21406, N21391, N1769);
xor XOR2 (N21407, N21397, N13490);
nor NOR3 (N21408, N21407, N12406, N910);
or OR4 (N21409, N21405, N10708, N17019, N8566);
and AND3 (N21410, N21393, N18144, N6980);
buf BUF1 (N21411, N21409);
or OR4 (N21412, N21406, N2816, N18927, N12702);
nor NOR4 (N21413, N21401, N7167, N241, N18679);
xor XOR2 (N21414, N21402, N20816);
xor XOR2 (N21415, N21404, N18699);
nor NOR3 (N21416, N21414, N4384, N14450);
buf BUF1 (N21417, N21408);
nor NOR2 (N21418, N21403, N5305);
nor NOR4 (N21419, N21418, N21151, N18710, N4162);
nand NAND3 (N21420, N21417, N20610, N15810);
xor XOR2 (N21421, N21411, N11713);
nand NAND4 (N21422, N21412, N13380, N19921, N3823);
buf BUF1 (N21423, N21419);
nand NAND2 (N21424, N21400, N5843);
nor NOR4 (N21425, N21422, N19172, N3273, N11159);
buf BUF1 (N21426, N21413);
nor NOR4 (N21427, N21395, N3503, N13541, N18383);
xor XOR2 (N21428, N21426, N40);
buf BUF1 (N21429, N21427);
buf BUF1 (N21430, N21428);
buf BUF1 (N21431, N21416);
xor XOR2 (N21432, N21421, N14989);
and AND3 (N21433, N21423, N2358, N12680);
not NOT1 (N21434, N21429);
buf BUF1 (N21435, N21424);
not NOT1 (N21436, N21432);
and AND4 (N21437, N21430, N12195, N18840, N15437);
xor XOR2 (N21438, N21437, N13320);
nand NAND4 (N21439, N21420, N19480, N11694, N13358);
or OR4 (N21440, N21435, N3083, N14345, N5070);
nand NAND4 (N21441, N21415, N17271, N20890, N14013);
buf BUF1 (N21442, N21439);
nor NOR3 (N21443, N21436, N6104, N19354);
or OR3 (N21444, N21442, N4950, N10163);
buf BUF1 (N21445, N21438);
and AND4 (N21446, N21444, N9722, N719, N1378);
xor XOR2 (N21447, N21433, N4645);
nor NOR4 (N21448, N21441, N1108, N21157, N3703);
or OR4 (N21449, N21440, N19860, N9456, N2482);
nor NOR2 (N21450, N21410, N7630);
nand NAND3 (N21451, N21434, N20777, N16764);
or OR2 (N21452, N21449, N15161);
buf BUF1 (N21453, N21448);
buf BUF1 (N21454, N21452);
or OR2 (N21455, N21443, N3478);
not NOT1 (N21456, N21425);
buf BUF1 (N21457, N21446);
not NOT1 (N21458, N21456);
nor NOR2 (N21459, N21455, N19196);
nand NAND3 (N21460, N21458, N14047, N8444);
xor XOR2 (N21461, N21454, N2181);
nand NAND3 (N21462, N21450, N9203, N260);
and AND2 (N21463, N21431, N10324);
nand NAND3 (N21464, N21459, N9360, N2395);
not NOT1 (N21465, N21453);
or OR2 (N21466, N21465, N7479);
xor XOR2 (N21467, N21462, N9025);
nand NAND3 (N21468, N21463, N17558, N20025);
buf BUF1 (N21469, N21460);
xor XOR2 (N21470, N21469, N3486);
buf BUF1 (N21471, N21468);
or OR4 (N21472, N21470, N16340, N20570, N8323);
or OR3 (N21473, N21472, N14238, N14747);
and AND4 (N21474, N21447, N9784, N9929, N8633);
nor NOR3 (N21475, N21457, N21116, N20688);
nor NOR2 (N21476, N21473, N2212);
not NOT1 (N21477, N21467);
or OR2 (N21478, N21477, N2201);
nor NOR3 (N21479, N21466, N13441, N2302);
not NOT1 (N21480, N21461);
and AND2 (N21481, N21451, N8406);
nor NOR3 (N21482, N21476, N13728, N9752);
nor NOR2 (N21483, N21479, N8854);
nand NAND2 (N21484, N21475, N18837);
and AND3 (N21485, N21481, N3881, N734);
buf BUF1 (N21486, N21484);
nor NOR3 (N21487, N21480, N17507, N2299);
or OR4 (N21488, N21482, N1824, N17792, N7311);
xor XOR2 (N21489, N21464, N1466);
nor NOR4 (N21490, N21474, N16261, N16036, N20007);
nand NAND4 (N21491, N21471, N15316, N2652, N20083);
and AND3 (N21492, N21478, N9839, N3502);
and AND2 (N21493, N21490, N5423);
and AND3 (N21494, N21492, N6593, N16823);
nand NAND3 (N21495, N21488, N5042, N12686);
xor XOR2 (N21496, N21493, N1122);
xor XOR2 (N21497, N21496, N4435);
nand NAND3 (N21498, N21494, N7922, N20096);
nand NAND3 (N21499, N21445, N6002, N14093);
buf BUF1 (N21500, N21498);
nor NOR3 (N21501, N21483, N9163, N11461);
xor XOR2 (N21502, N21501, N6123);
and AND3 (N21503, N21486, N6526, N10506);
not NOT1 (N21504, N21485);
or OR3 (N21505, N21499, N11195, N2817);
nand NAND2 (N21506, N21497, N11288);
xor XOR2 (N21507, N21487, N15711);
buf BUF1 (N21508, N21503);
xor XOR2 (N21509, N21489, N17193);
and AND3 (N21510, N21495, N13134, N3874);
xor XOR2 (N21511, N21502, N6832);
nor NOR4 (N21512, N21508, N20205, N12664, N9924);
not NOT1 (N21513, N21505);
not NOT1 (N21514, N21504);
nor NOR2 (N21515, N21491, N7503);
xor XOR2 (N21516, N21515, N3442);
or OR3 (N21517, N21513, N10976, N16597);
and AND3 (N21518, N21507, N8184, N5372);
xor XOR2 (N21519, N21516, N13409);
buf BUF1 (N21520, N21510);
and AND3 (N21521, N21519, N19828, N4848);
nand NAND3 (N21522, N21500, N18398, N14241);
nand NAND3 (N21523, N21514, N9469, N16017);
not NOT1 (N21524, N21512);
and AND4 (N21525, N21522, N13430, N9479, N12511);
and AND3 (N21526, N21518, N6865, N13318);
nand NAND4 (N21527, N21521, N9090, N8716, N6602);
xor XOR2 (N21528, N21517, N7865);
or OR3 (N21529, N21511, N9611, N2298);
buf BUF1 (N21530, N21509);
buf BUF1 (N21531, N21506);
buf BUF1 (N21532, N21529);
xor XOR2 (N21533, N21525, N2359);
not NOT1 (N21534, N21527);
and AND4 (N21535, N21520, N1231, N14890, N14639);
buf BUF1 (N21536, N21532);
or OR3 (N21537, N21524, N16523, N15508);
or OR2 (N21538, N21533, N16000);
nand NAND4 (N21539, N21523, N11308, N13953, N6859);
buf BUF1 (N21540, N21528);
not NOT1 (N21541, N21537);
buf BUF1 (N21542, N21539);
xor XOR2 (N21543, N21530, N19440);
xor XOR2 (N21544, N21535, N17065);
or OR4 (N21545, N21534, N9806, N3122, N14724);
and AND3 (N21546, N21543, N17464, N1489);
nand NAND3 (N21547, N21542, N10134, N4448);
and AND3 (N21548, N21544, N6948, N13557);
and AND2 (N21549, N21545, N9902);
not NOT1 (N21550, N21536);
xor XOR2 (N21551, N21531, N17928);
nand NAND4 (N21552, N21547, N12936, N4360, N5278);
buf BUF1 (N21553, N21526);
and AND2 (N21554, N21550, N8811);
xor XOR2 (N21555, N21554, N8493);
nor NOR3 (N21556, N21549, N20473, N20458);
buf BUF1 (N21557, N21541);
and AND4 (N21558, N21546, N19218, N15094, N10962);
not NOT1 (N21559, N21552);
buf BUF1 (N21560, N21557);
nand NAND3 (N21561, N21538, N9707, N15740);
not NOT1 (N21562, N21561);
xor XOR2 (N21563, N21558, N10836);
and AND3 (N21564, N21559, N15333, N6386);
or OR3 (N21565, N21564, N13796, N9249);
and AND2 (N21566, N21560, N1656);
nand NAND3 (N21567, N21562, N4229, N15242);
buf BUF1 (N21568, N21566);
and AND4 (N21569, N21555, N18572, N3378, N13449);
nand NAND3 (N21570, N21540, N13095, N14289);
nor NOR2 (N21571, N21548, N4107);
xor XOR2 (N21572, N21563, N6098);
not NOT1 (N21573, N21556);
buf BUF1 (N21574, N21573);
and AND4 (N21575, N21569, N17545, N9975, N16708);
buf BUF1 (N21576, N21572);
xor XOR2 (N21577, N21576, N11183);
buf BUF1 (N21578, N21553);
xor XOR2 (N21579, N21571, N19539);
nor NOR4 (N21580, N21568, N11605, N14353, N9835);
not NOT1 (N21581, N21570);
nor NOR4 (N21582, N21581, N2315, N2626, N4913);
or OR2 (N21583, N21575, N15939);
or OR2 (N21584, N21551, N2609);
and AND2 (N21585, N21565, N20654);
nand NAND3 (N21586, N21584, N4034, N4254);
nor NOR4 (N21587, N21578, N13740, N11503, N19778);
nor NOR2 (N21588, N21577, N17817);
nand NAND2 (N21589, N21574, N11704);
and AND2 (N21590, N21582, N9938);
nor NOR4 (N21591, N21579, N10829, N6270, N12570);
nor NOR3 (N21592, N21587, N10094, N5930);
nor NOR4 (N21593, N21583, N17276, N19358, N1378);
xor XOR2 (N21594, N21591, N19998);
or OR2 (N21595, N21585, N17329);
nand NAND2 (N21596, N21592, N3010);
xor XOR2 (N21597, N21589, N14955);
not NOT1 (N21598, N21586);
or OR3 (N21599, N21593, N8269, N18990);
not NOT1 (N21600, N21599);
buf BUF1 (N21601, N21588);
nand NAND3 (N21602, N21600, N16976, N6146);
buf BUF1 (N21603, N21594);
nor NOR3 (N21604, N21603, N2551, N8259);
not NOT1 (N21605, N21598);
buf BUF1 (N21606, N21605);
not NOT1 (N21607, N21604);
nand NAND3 (N21608, N21567, N15162, N2172);
buf BUF1 (N21609, N21595);
or OR2 (N21610, N21597, N13413);
nor NOR2 (N21611, N21590, N14020);
buf BUF1 (N21612, N21580);
xor XOR2 (N21613, N21609, N2034);
buf BUF1 (N21614, N21612);
not NOT1 (N21615, N21614);
and AND2 (N21616, N21601, N12723);
or OR2 (N21617, N21610, N14715);
nor NOR4 (N21618, N21615, N2985, N7235, N12912);
not NOT1 (N21619, N21617);
or OR3 (N21620, N21607, N13004, N9723);
nand NAND2 (N21621, N21616, N408);
not NOT1 (N21622, N21618);
nor NOR4 (N21623, N21608, N7217, N7288, N19327);
nor NOR3 (N21624, N21613, N20037, N11476);
nand NAND3 (N21625, N21596, N14175, N12472);
nor NOR2 (N21626, N21621, N11920);
or OR3 (N21627, N21623, N14675, N2748);
nor NOR3 (N21628, N21625, N19471, N13288);
xor XOR2 (N21629, N21622, N1303);
and AND3 (N21630, N21627, N12432, N3980);
or OR3 (N21631, N21628, N9460, N15550);
and AND3 (N21632, N21619, N7470, N1667);
buf BUF1 (N21633, N21629);
nor NOR4 (N21634, N21624, N1765, N8169, N16558);
nor NOR4 (N21635, N21620, N5188, N8152, N13835);
xor XOR2 (N21636, N21626, N2205);
nand NAND2 (N21637, N21602, N17150);
buf BUF1 (N21638, N21631);
xor XOR2 (N21639, N21637, N5119);
or OR2 (N21640, N21639, N4480);
buf BUF1 (N21641, N21640);
xor XOR2 (N21642, N21636, N17343);
and AND2 (N21643, N21611, N6157);
nor NOR3 (N21644, N21630, N7932, N21008);
buf BUF1 (N21645, N21641);
buf BUF1 (N21646, N21642);
nand NAND2 (N21647, N21646, N21321);
not NOT1 (N21648, N21633);
and AND2 (N21649, N21638, N10588);
buf BUF1 (N21650, N21643);
or OR4 (N21651, N21650, N18888, N21519, N6116);
not NOT1 (N21652, N21651);
and AND3 (N21653, N21647, N2006, N1157);
nor NOR2 (N21654, N21652, N630);
or OR4 (N21655, N21649, N1509, N13938, N16323);
buf BUF1 (N21656, N21632);
nor NOR2 (N21657, N21656, N11729);
xor XOR2 (N21658, N21654, N16456);
not NOT1 (N21659, N21606);
not NOT1 (N21660, N21634);
nand NAND4 (N21661, N21645, N2933, N9759, N12823);
or OR2 (N21662, N21644, N15931);
buf BUF1 (N21663, N21660);
or OR4 (N21664, N21655, N20510, N12374, N6653);
and AND2 (N21665, N21661, N13543);
nor NOR3 (N21666, N21635, N12666, N6685);
nand NAND3 (N21667, N21666, N880, N20461);
nor NOR4 (N21668, N21664, N16022, N4032, N17882);
buf BUF1 (N21669, N21667);
buf BUF1 (N21670, N21648);
or OR2 (N21671, N21669, N21542);
or OR2 (N21672, N21659, N16994);
nor NOR3 (N21673, N21672, N11719, N729);
xor XOR2 (N21674, N21658, N19638);
and AND3 (N21675, N21671, N677, N21450);
not NOT1 (N21676, N21668);
and AND3 (N21677, N21653, N17750, N5513);
xor XOR2 (N21678, N21657, N14132);
nor NOR3 (N21679, N21674, N4891, N5726);
not NOT1 (N21680, N21662);
nand NAND4 (N21681, N21676, N17011, N13837, N12633);
nand NAND4 (N21682, N21663, N16928, N21360, N20845);
buf BUF1 (N21683, N21678);
nor NOR4 (N21684, N21677, N7246, N9592, N7073);
or OR2 (N21685, N21665, N17893);
nand NAND2 (N21686, N21675, N10489);
xor XOR2 (N21687, N21680, N5424);
and AND4 (N21688, N21679, N13419, N16074, N2897);
and AND4 (N21689, N21670, N20017, N370, N15201);
nand NAND4 (N21690, N21687, N2139, N9775, N11334);
xor XOR2 (N21691, N21690, N16275);
and AND2 (N21692, N21673, N13898);
xor XOR2 (N21693, N21691, N2341);
nor NOR2 (N21694, N21682, N9075);
not NOT1 (N21695, N21694);
nor NOR3 (N21696, N21689, N18859, N9284);
nand NAND2 (N21697, N21688, N11337);
or OR2 (N21698, N21685, N536);
xor XOR2 (N21699, N21695, N5277);
not NOT1 (N21700, N21681);
or OR4 (N21701, N21693, N11580, N664, N7835);
not NOT1 (N21702, N21684);
or OR3 (N21703, N21702, N14268, N11078);
and AND2 (N21704, N21697, N13083);
nor NOR4 (N21705, N21701, N1578, N16455, N7387);
nor NOR3 (N21706, N21699, N16593, N15814);
not NOT1 (N21707, N21696);
not NOT1 (N21708, N21705);
xor XOR2 (N21709, N21698, N7437);
buf BUF1 (N21710, N21706);
or OR3 (N21711, N21703, N2141, N4528);
or OR3 (N21712, N21708, N7663, N18902);
or OR2 (N21713, N21686, N19095);
and AND4 (N21714, N21692, N6928, N15269, N4558);
and AND3 (N21715, N21700, N15343, N14849);
nor NOR4 (N21716, N21709, N7056, N10977, N4556);
and AND3 (N21717, N21683, N3976, N16469);
nand NAND4 (N21718, N21713, N19381, N12913, N18435);
buf BUF1 (N21719, N21707);
nand NAND4 (N21720, N21718, N18997, N1590, N2929);
nand NAND4 (N21721, N21719, N581, N17767, N8087);
and AND4 (N21722, N21717, N999, N16327, N20344);
or OR4 (N21723, N21722, N12680, N8563, N19092);
xor XOR2 (N21724, N21711, N17899);
xor XOR2 (N21725, N21704, N2560);
and AND2 (N21726, N21725, N18327);
and AND3 (N21727, N21710, N15196, N19781);
nor NOR3 (N21728, N21716, N15430, N6996);
buf BUF1 (N21729, N21727);
not NOT1 (N21730, N21714);
nand NAND4 (N21731, N21723, N18898, N19988, N3918);
xor XOR2 (N21732, N21724, N1378);
and AND3 (N21733, N21721, N19232, N3275);
nand NAND3 (N21734, N21733, N5628, N5594);
buf BUF1 (N21735, N21729);
not NOT1 (N21736, N21732);
not NOT1 (N21737, N21730);
buf BUF1 (N21738, N21728);
buf BUF1 (N21739, N21715);
not NOT1 (N21740, N21738);
not NOT1 (N21741, N21720);
nand NAND2 (N21742, N21726, N3880);
nor NOR2 (N21743, N21737, N12823);
xor XOR2 (N21744, N21735, N7327);
buf BUF1 (N21745, N21734);
nand NAND2 (N21746, N21745, N12010);
nand NAND2 (N21747, N21736, N9585);
not NOT1 (N21748, N21739);
or OR4 (N21749, N21743, N20892, N21527, N20305);
not NOT1 (N21750, N21742);
not NOT1 (N21751, N21741);
and AND3 (N21752, N21712, N8417, N10508);
buf BUF1 (N21753, N21731);
xor XOR2 (N21754, N21749, N20522);
nand NAND4 (N21755, N21751, N12519, N9546, N19754);
nand NAND3 (N21756, N21747, N10195, N15189);
and AND4 (N21757, N21754, N1385, N14743, N4699);
xor XOR2 (N21758, N21752, N14650);
nor NOR2 (N21759, N21755, N15996);
buf BUF1 (N21760, N21740);
buf BUF1 (N21761, N21759);
not NOT1 (N21762, N21753);
xor XOR2 (N21763, N21750, N11463);
or OR4 (N21764, N21757, N5551, N4672, N13623);
nor NOR3 (N21765, N21746, N8936, N15265);
nor NOR3 (N21766, N21760, N7050, N14066);
buf BUF1 (N21767, N21744);
or OR3 (N21768, N21767, N2867, N20544);
or OR4 (N21769, N21765, N5102, N581, N5232);
buf BUF1 (N21770, N21762);
or OR2 (N21771, N21766, N17758);
nand NAND3 (N21772, N21756, N15540, N18704);
or OR4 (N21773, N21748, N15347, N4593, N13184);
and AND2 (N21774, N21761, N14143);
nand NAND2 (N21775, N21774, N10250);
nand NAND3 (N21776, N21771, N12638, N11251);
and AND3 (N21777, N21758, N1244, N4037);
nor NOR2 (N21778, N21769, N9115);
or OR4 (N21779, N21770, N1117, N15447, N15259);
or OR2 (N21780, N21778, N20124);
xor XOR2 (N21781, N21779, N1538);
and AND2 (N21782, N21772, N10588);
or OR3 (N21783, N21780, N204, N1666);
not NOT1 (N21784, N21773);
nand NAND4 (N21785, N21775, N18128, N15477, N15622);
and AND2 (N21786, N21784, N17351);
buf BUF1 (N21787, N21783);
xor XOR2 (N21788, N21781, N14707);
and AND4 (N21789, N21776, N12052, N7034, N15395);
not NOT1 (N21790, N21787);
nand NAND2 (N21791, N21790, N4562);
xor XOR2 (N21792, N21785, N10909);
xor XOR2 (N21793, N21788, N21615);
xor XOR2 (N21794, N21789, N21603);
xor XOR2 (N21795, N21764, N5122);
buf BUF1 (N21796, N21794);
and AND3 (N21797, N21792, N1837, N17364);
nand NAND4 (N21798, N21782, N967, N20934, N18016);
or OR2 (N21799, N21798, N18351);
xor XOR2 (N21800, N21777, N18883);
nand NAND3 (N21801, N21786, N20597, N24);
not NOT1 (N21802, N21795);
and AND2 (N21803, N21799, N9843);
not NOT1 (N21804, N21768);
or OR4 (N21805, N21802, N888, N11413, N20317);
nand NAND3 (N21806, N21803, N10442, N1944);
or OR4 (N21807, N21804, N16716, N842, N4436);
not NOT1 (N21808, N21807);
xor XOR2 (N21809, N21801, N10100);
xor XOR2 (N21810, N21796, N21291);
xor XOR2 (N21811, N21800, N20723);
and AND3 (N21812, N21808, N2426, N15296);
or OR4 (N21813, N21791, N545, N170, N1989);
nand NAND4 (N21814, N21793, N19163, N15720, N19948);
nor NOR3 (N21815, N21797, N4126, N17833);
not NOT1 (N21816, N21814);
buf BUF1 (N21817, N21815);
nor NOR2 (N21818, N21806, N5374);
nand NAND3 (N21819, N21812, N2894, N17898);
nor NOR2 (N21820, N21817, N12190);
or OR3 (N21821, N21811, N19141, N6298);
buf BUF1 (N21822, N21821);
nor NOR3 (N21823, N21818, N15942, N13883);
nor NOR2 (N21824, N21820, N15733);
not NOT1 (N21825, N21822);
buf BUF1 (N21826, N21819);
and AND3 (N21827, N21824, N6804, N15086);
not NOT1 (N21828, N21823);
xor XOR2 (N21829, N21828, N10565);
not NOT1 (N21830, N21825);
nor NOR4 (N21831, N21813, N18809, N20173, N16536);
not NOT1 (N21832, N21805);
or OR3 (N21833, N21832, N18862, N4628);
nand NAND3 (N21834, N21816, N9852, N14122);
or OR4 (N21835, N21833, N10964, N64, N11936);
nand NAND4 (N21836, N21829, N2807, N13152, N17525);
xor XOR2 (N21837, N21830, N2488);
buf BUF1 (N21838, N21827);
not NOT1 (N21839, N21763);
nor NOR2 (N21840, N21826, N12121);
nor NOR3 (N21841, N21809, N8901, N10498);
xor XOR2 (N21842, N21834, N15952);
and AND3 (N21843, N21841, N4848, N16189);
not NOT1 (N21844, N21835);
not NOT1 (N21845, N21843);
xor XOR2 (N21846, N21837, N1113);
and AND2 (N21847, N21842, N16876);
nand NAND2 (N21848, N21810, N12503);
buf BUF1 (N21849, N21845);
not NOT1 (N21850, N21846);
xor XOR2 (N21851, N21840, N9341);
not NOT1 (N21852, N21851);
and AND4 (N21853, N21839, N19009, N5875, N460);
and AND3 (N21854, N21844, N1440, N7556);
xor XOR2 (N21855, N21831, N11387);
nor NOR4 (N21856, N21855, N13097, N10550, N6309);
nor NOR4 (N21857, N21850, N5268, N4073, N7336);
not NOT1 (N21858, N21854);
xor XOR2 (N21859, N21857, N17967);
not NOT1 (N21860, N21836);
nor NOR4 (N21861, N21860, N7385, N8795, N18816);
buf BUF1 (N21862, N21838);
and AND2 (N21863, N21853, N3291);
or OR2 (N21864, N21849, N18339);
nor NOR3 (N21865, N21858, N2107, N21340);
nor NOR2 (N21866, N21865, N10961);
buf BUF1 (N21867, N21856);
not NOT1 (N21868, N21862);
nor NOR3 (N21869, N21847, N640, N17128);
and AND3 (N21870, N21863, N3697, N14457);
nand NAND2 (N21871, N21861, N7970);
buf BUF1 (N21872, N21852);
and AND3 (N21873, N21871, N15385, N8626);
nor NOR2 (N21874, N21859, N16349);
buf BUF1 (N21875, N21864);
nor NOR2 (N21876, N21874, N896);
nand NAND2 (N21877, N21867, N20125);
buf BUF1 (N21878, N21848);
and AND3 (N21879, N21872, N10346, N14793);
nand NAND4 (N21880, N21873, N7341, N17222, N3106);
not NOT1 (N21881, N21878);
and AND4 (N21882, N21868, N6493, N9797, N17593);
and AND4 (N21883, N21876, N2250, N232, N11647);
buf BUF1 (N21884, N21866);
not NOT1 (N21885, N21879);
or OR2 (N21886, N21870, N17677);
buf BUF1 (N21887, N21881);
buf BUF1 (N21888, N21886);
nor NOR4 (N21889, N21869, N7235, N17380, N11247);
or OR3 (N21890, N21875, N4399, N14126);
or OR4 (N21891, N21887, N13704, N10477, N12686);
buf BUF1 (N21892, N21883);
or OR2 (N21893, N21885, N19784);
or OR2 (N21894, N21892, N19439);
and AND4 (N21895, N21877, N14813, N7873, N7888);
buf BUF1 (N21896, N21893);
and AND4 (N21897, N21884, N12470, N5400, N14796);
not NOT1 (N21898, N21889);
or OR4 (N21899, N21891, N18998, N5660, N20238);
xor XOR2 (N21900, N21888, N7929);
buf BUF1 (N21901, N21895);
buf BUF1 (N21902, N21894);
and AND4 (N21903, N21896, N16529, N7625, N13589);
or OR4 (N21904, N21903, N13693, N4923, N17885);
nand NAND4 (N21905, N21897, N2838, N12839, N11670);
xor XOR2 (N21906, N21904, N15008);
or OR3 (N21907, N21901, N8770, N9187);
xor XOR2 (N21908, N21906, N10073);
xor XOR2 (N21909, N21890, N180);
buf BUF1 (N21910, N21907);
and AND4 (N21911, N21899, N19628, N8001, N1611);
nor NOR3 (N21912, N21880, N12291, N6309);
not NOT1 (N21913, N21912);
buf BUF1 (N21914, N21908);
buf BUF1 (N21915, N21902);
not NOT1 (N21916, N21882);
buf BUF1 (N21917, N21911);
xor XOR2 (N21918, N21915, N13966);
nor NOR3 (N21919, N21913, N8896, N18467);
nor NOR4 (N21920, N21916, N14078, N768, N14443);
nor NOR4 (N21921, N21920, N14201, N9811, N5048);
nor NOR2 (N21922, N21909, N18508);
nand NAND4 (N21923, N21917, N18993, N15379, N27);
buf BUF1 (N21924, N21921);
not NOT1 (N21925, N21923);
nand NAND3 (N21926, N21919, N5841, N12450);
nand NAND2 (N21927, N21926, N19675);
not NOT1 (N21928, N21900);
or OR4 (N21929, N21927, N6908, N5097, N11444);
not NOT1 (N21930, N21918);
xor XOR2 (N21931, N21910, N2373);
not NOT1 (N21932, N21929);
xor XOR2 (N21933, N21922, N244);
nand NAND3 (N21934, N21924, N20065, N17848);
or OR3 (N21935, N21905, N5289, N20425);
or OR2 (N21936, N21898, N6894);
and AND2 (N21937, N21914, N3505);
nor NOR4 (N21938, N21934, N11451, N20791, N4392);
nand NAND3 (N21939, N21930, N16596, N11132);
and AND4 (N21940, N21931, N19329, N21563, N13589);
not NOT1 (N21941, N21940);
or OR3 (N21942, N21933, N16414, N13610);
not NOT1 (N21943, N21937);
nand NAND3 (N21944, N21938, N16099, N3698);
nand NAND4 (N21945, N21936, N3803, N11228, N8923);
or OR2 (N21946, N21932, N4163);
nand NAND2 (N21947, N21943, N9258);
not NOT1 (N21948, N21944);
nor NOR3 (N21949, N21948, N2873, N2190);
xor XOR2 (N21950, N21941, N12143);
buf BUF1 (N21951, N21925);
not NOT1 (N21952, N21951);
not NOT1 (N21953, N21946);
and AND4 (N21954, N21952, N4665, N11537, N18185);
nand NAND3 (N21955, N21945, N3067, N5831);
not NOT1 (N21956, N21953);
and AND2 (N21957, N21954, N18286);
buf BUF1 (N21958, N21949);
not NOT1 (N21959, N21935);
xor XOR2 (N21960, N21928, N5163);
not NOT1 (N21961, N21960);
buf BUF1 (N21962, N21957);
xor XOR2 (N21963, N21959, N9385);
buf BUF1 (N21964, N21939);
xor XOR2 (N21965, N21942, N3977);
xor XOR2 (N21966, N21958, N12449);
and AND3 (N21967, N21965, N5445, N19731);
buf BUF1 (N21968, N21955);
nand NAND4 (N21969, N21961, N6282, N9923, N6879);
and AND3 (N21970, N21968, N3644, N11079);
buf BUF1 (N21971, N21947);
or OR2 (N21972, N21967, N20609);
not NOT1 (N21973, N21963);
not NOT1 (N21974, N21966);
xor XOR2 (N21975, N21956, N15740);
or OR4 (N21976, N21975, N5583, N10149, N20949);
nand NAND3 (N21977, N21964, N11837, N16089);
nand NAND3 (N21978, N21974, N15029, N16693);
nand NAND3 (N21979, N21973, N7733, N3068);
buf BUF1 (N21980, N21976);
xor XOR2 (N21981, N21971, N10390);
nand NAND2 (N21982, N21978, N17405);
nand NAND3 (N21983, N21979, N14406, N8929);
or OR3 (N21984, N21977, N1756, N12855);
xor XOR2 (N21985, N21970, N15361);
or OR4 (N21986, N21983, N15857, N17454, N8428);
xor XOR2 (N21987, N21962, N19692);
xor XOR2 (N21988, N21982, N4575);
or OR4 (N21989, N21986, N14705, N14419, N13025);
or OR3 (N21990, N21988, N1807, N8365);
xor XOR2 (N21991, N21989, N8713);
nor NOR4 (N21992, N21980, N4366, N6000, N15714);
not NOT1 (N21993, N21987);
buf BUF1 (N21994, N21993);
and AND3 (N21995, N21984, N13913, N20473);
and AND4 (N21996, N21969, N6308, N12380, N12443);
nand NAND3 (N21997, N21950, N18110, N12265);
xor XOR2 (N21998, N21996, N8700);
nor NOR2 (N21999, N21995, N19909);
or OR4 (N22000, N21992, N7028, N18269, N16001);
nor NOR3 (N22001, N21990, N1102, N7508);
and AND3 (N22002, N21991, N2007, N13922);
not NOT1 (N22003, N22002);
not NOT1 (N22004, N22000);
xor XOR2 (N22005, N21994, N21818);
xor XOR2 (N22006, N22003, N2362);
xor XOR2 (N22007, N21981, N14532);
and AND3 (N22008, N21997, N21920, N9860);
not NOT1 (N22009, N22004);
nand NAND3 (N22010, N21999, N21022, N21671);
or OR3 (N22011, N22010, N10749, N21527);
not NOT1 (N22012, N22001);
not NOT1 (N22013, N21985);
nand NAND2 (N22014, N21972, N13634);
or OR2 (N22015, N21998, N254);
xor XOR2 (N22016, N22006, N7380);
xor XOR2 (N22017, N22005, N4481);
buf BUF1 (N22018, N22009);
nand NAND3 (N22019, N22015, N20985, N888);
not NOT1 (N22020, N22013);
or OR4 (N22021, N22020, N10199, N13963, N7767);
xor XOR2 (N22022, N22008, N12609);
nor NOR3 (N22023, N22016, N17363, N9559);
nand NAND2 (N22024, N22019, N20517);
nor NOR2 (N22025, N22022, N10660);
buf BUF1 (N22026, N22021);
or OR2 (N22027, N22024, N2153);
nor NOR3 (N22028, N22017, N1472, N9741);
buf BUF1 (N22029, N22011);
buf BUF1 (N22030, N22023);
or OR3 (N22031, N22018, N1751, N10448);
not NOT1 (N22032, N22029);
xor XOR2 (N22033, N22025, N8514);
nor NOR2 (N22034, N22014, N19898);
or OR3 (N22035, N22032, N5489, N17169);
or OR3 (N22036, N22026, N9571, N6300);
not NOT1 (N22037, N22012);
xor XOR2 (N22038, N22036, N8244);
nand NAND2 (N22039, N22038, N1671);
nand NAND3 (N22040, N22037, N19227, N19173);
not NOT1 (N22041, N22039);
nor NOR3 (N22042, N22007, N1179, N6299);
nor NOR4 (N22043, N22027, N2174, N9048, N6608);
nor NOR3 (N22044, N22033, N11413, N3129);
buf BUF1 (N22045, N22044);
xor XOR2 (N22046, N22031, N5731);
nand NAND2 (N22047, N22035, N442);
nand NAND4 (N22048, N22042, N1241, N7037, N16122);
xor XOR2 (N22049, N22030, N20588);
nor NOR3 (N22050, N22043, N20772, N8747);
nor NOR3 (N22051, N22048, N4963, N12410);
and AND3 (N22052, N22028, N19498, N13368);
nand NAND4 (N22053, N22052, N8750, N12301, N13882);
and AND4 (N22054, N22040, N17888, N7960, N16875);
and AND4 (N22055, N22047, N20716, N8575, N11843);
not NOT1 (N22056, N22054);
xor XOR2 (N22057, N22041, N19215);
buf BUF1 (N22058, N22053);
buf BUF1 (N22059, N22058);
nand NAND3 (N22060, N22057, N18963, N19822);
and AND2 (N22061, N22051, N13328);
nand NAND3 (N22062, N22056, N3369, N16337);
nand NAND2 (N22063, N22050, N10729);
nand NAND2 (N22064, N22045, N198);
and AND3 (N22065, N22055, N17736, N18350);
and AND3 (N22066, N22049, N5140, N19538);
buf BUF1 (N22067, N22066);
buf BUF1 (N22068, N22034);
xor XOR2 (N22069, N22046, N10350);
or OR2 (N22070, N22063, N17425);
nor NOR4 (N22071, N22062, N1070, N4986, N14611);
nand NAND4 (N22072, N22069, N14102, N12387, N7920);
and AND4 (N22073, N22060, N2822, N15994, N7430);
nand NAND3 (N22074, N22072, N2156, N2658);
not NOT1 (N22075, N22070);
xor XOR2 (N22076, N22064, N20000);
not NOT1 (N22077, N22065);
nand NAND4 (N22078, N22075, N337, N13127, N7928);
nand NAND4 (N22079, N22068, N2849, N20750, N17192);
buf BUF1 (N22080, N22079);
not NOT1 (N22081, N22078);
buf BUF1 (N22082, N22073);
not NOT1 (N22083, N22080);
not NOT1 (N22084, N22059);
nand NAND3 (N22085, N22081, N14933, N11105);
and AND2 (N22086, N22085, N13611);
or OR4 (N22087, N22084, N5407, N13203, N19428);
nor NOR2 (N22088, N22086, N20509);
nand NAND3 (N22089, N22071, N12054, N19007);
buf BUF1 (N22090, N22067);
or OR2 (N22091, N22089, N17070);
not NOT1 (N22092, N22083);
or OR2 (N22093, N22077, N5516);
and AND3 (N22094, N22093, N5961, N6872);
xor XOR2 (N22095, N22087, N13363);
not NOT1 (N22096, N22082);
and AND2 (N22097, N22061, N1662);
nor NOR3 (N22098, N22094, N6467, N12444);
xor XOR2 (N22099, N22074, N11894);
xor XOR2 (N22100, N22091, N10032);
buf BUF1 (N22101, N22100);
nor NOR3 (N22102, N22095, N6451, N9873);
xor XOR2 (N22103, N22088, N3610);
nand NAND4 (N22104, N22097, N17083, N6808, N11137);
nor NOR2 (N22105, N22092, N20842);
xor XOR2 (N22106, N22076, N4649);
not NOT1 (N22107, N22104);
nor NOR3 (N22108, N22098, N1870, N13627);
nand NAND3 (N22109, N22096, N11567, N11365);
and AND4 (N22110, N22101, N2048, N18781, N11602);
or OR4 (N22111, N22103, N6156, N11182, N1477);
nor NOR2 (N22112, N22105, N2388);
nand NAND3 (N22113, N22090, N5528, N6464);
nand NAND2 (N22114, N22108, N13279);
xor XOR2 (N22115, N22099, N9009);
xor XOR2 (N22116, N22107, N232);
buf BUF1 (N22117, N22115);
or OR2 (N22118, N22112, N21060);
nor NOR3 (N22119, N22116, N21701, N8825);
or OR4 (N22120, N22110, N5652, N1560, N1526);
nand NAND4 (N22121, N22120, N14708, N9754, N7411);
nor NOR4 (N22122, N22119, N10874, N12832, N9963);
nor NOR4 (N22123, N22118, N19248, N6185, N1000);
nor NOR2 (N22124, N22113, N1455);
and AND3 (N22125, N22123, N11633, N3687);
and AND3 (N22126, N22106, N8635, N4654);
or OR4 (N22127, N22125, N8496, N1086, N4217);
nor NOR4 (N22128, N22111, N3971, N1176, N14350);
nand NAND2 (N22129, N22117, N5571);
buf BUF1 (N22130, N22121);
nor NOR4 (N22131, N22122, N6359, N8865, N3876);
nor NOR2 (N22132, N22130, N6508);
and AND4 (N22133, N22126, N1412, N18694, N20974);
and AND4 (N22134, N22109, N6170, N8490, N15183);
not NOT1 (N22135, N22134);
or OR4 (N22136, N22124, N12108, N16809, N20563);
xor XOR2 (N22137, N22129, N16925);
buf BUF1 (N22138, N22102);
buf BUF1 (N22139, N22132);
buf BUF1 (N22140, N22127);
nand NAND4 (N22141, N22138, N8372, N1799, N11881);
buf BUF1 (N22142, N22135);
buf BUF1 (N22143, N22142);
or OR2 (N22144, N22128, N6998);
or OR3 (N22145, N22139, N5180, N15246);
not NOT1 (N22146, N22136);
not NOT1 (N22147, N22131);
nor NOR4 (N22148, N22141, N15381, N18706, N17769);
nand NAND4 (N22149, N22114, N17836, N1937, N17961);
buf BUF1 (N22150, N22145);
buf BUF1 (N22151, N22149);
xor XOR2 (N22152, N22137, N10612);
or OR2 (N22153, N22146, N3522);
xor XOR2 (N22154, N22148, N20465);
nor NOR4 (N22155, N22133, N2933, N2235, N7125);
not NOT1 (N22156, N22151);
or OR4 (N22157, N22147, N17876, N14365, N19620);
nand NAND4 (N22158, N22152, N13453, N8400, N1809);
nor NOR3 (N22159, N22154, N10778, N15416);
not NOT1 (N22160, N22156);
xor XOR2 (N22161, N22140, N20081);
and AND4 (N22162, N22160, N18376, N10823, N10250);
not NOT1 (N22163, N22158);
and AND2 (N22164, N22157, N21253);
xor XOR2 (N22165, N22144, N9122);
not NOT1 (N22166, N22163);
nand NAND4 (N22167, N22166, N3170, N13483, N6751);
and AND2 (N22168, N22161, N5006);
and AND2 (N22169, N22165, N7950);
nor NOR2 (N22170, N22143, N13722);
not NOT1 (N22171, N22170);
and AND4 (N22172, N22169, N18432, N18342, N10782);
and AND3 (N22173, N22150, N10731, N6631);
buf BUF1 (N22174, N22155);
nor NOR3 (N22175, N22172, N15761, N16973);
not NOT1 (N22176, N22175);
nor NOR3 (N22177, N22159, N9687, N15022);
nor NOR4 (N22178, N22153, N3475, N3169, N19264);
nand NAND3 (N22179, N22167, N15856, N2260);
not NOT1 (N22180, N22173);
xor XOR2 (N22181, N22164, N15475);
buf BUF1 (N22182, N22180);
buf BUF1 (N22183, N22176);
nor NOR4 (N22184, N22181, N18506, N8116, N20275);
nand NAND3 (N22185, N22184, N12521, N7389);
buf BUF1 (N22186, N22178);
buf BUF1 (N22187, N22182);
buf BUF1 (N22188, N22185);
xor XOR2 (N22189, N22186, N14305);
or OR3 (N22190, N22189, N12670, N15557);
xor XOR2 (N22191, N22177, N20855);
xor XOR2 (N22192, N22171, N17836);
nor NOR2 (N22193, N22168, N5343);
nand NAND4 (N22194, N22193, N14021, N7478, N19145);
and AND4 (N22195, N22162, N19329, N7954, N9945);
not NOT1 (N22196, N22179);
or OR2 (N22197, N22174, N10184);
or OR4 (N22198, N22183, N5899, N1425, N14722);
buf BUF1 (N22199, N22187);
nand NAND4 (N22200, N22198, N21351, N20577, N9530);
or OR2 (N22201, N22197, N10572);
nand NAND3 (N22202, N22199, N11839, N6241);
nor NOR4 (N22203, N22202, N797, N13575, N6643);
nor NOR2 (N22204, N22200, N8995);
nor NOR3 (N22205, N22203, N13847, N6003);
xor XOR2 (N22206, N22190, N7409);
nor NOR4 (N22207, N22192, N16751, N11077, N4020);
nor NOR3 (N22208, N22201, N5050, N1917);
xor XOR2 (N22209, N22205, N15617);
nand NAND3 (N22210, N22206, N18932, N13819);
or OR3 (N22211, N22210, N510, N3960);
not NOT1 (N22212, N22188);
buf BUF1 (N22213, N22208);
nand NAND3 (N22214, N22213, N1809, N11803);
or OR3 (N22215, N22204, N18608, N8397);
xor XOR2 (N22216, N22191, N18590);
nor NOR2 (N22217, N22194, N8205);
nor NOR2 (N22218, N22209, N8116);
xor XOR2 (N22219, N22214, N13031);
nor NOR2 (N22220, N22212, N18777);
or OR2 (N22221, N22216, N17461);
or OR2 (N22222, N22207, N6266);
xor XOR2 (N22223, N22195, N9304);
and AND2 (N22224, N22218, N3906);
not NOT1 (N22225, N22211);
or OR2 (N22226, N22221, N5889);
xor XOR2 (N22227, N22224, N4057);
nand NAND2 (N22228, N22219, N21762);
nand NAND4 (N22229, N22220, N4929, N7634, N2405);
not NOT1 (N22230, N22223);
xor XOR2 (N22231, N22215, N16103);
xor XOR2 (N22232, N22217, N15068);
nand NAND2 (N22233, N22227, N4042);
nor NOR4 (N22234, N22231, N16532, N12193, N14545);
or OR4 (N22235, N22233, N1538, N13961, N18516);
not NOT1 (N22236, N22196);
nand NAND4 (N22237, N22232, N7392, N10615, N1094);
nand NAND2 (N22238, N22236, N5800);
or OR4 (N22239, N22226, N18731, N13957, N15269);
xor XOR2 (N22240, N22230, N21979);
xor XOR2 (N22241, N22238, N18276);
or OR2 (N22242, N22234, N16105);
not NOT1 (N22243, N22241);
or OR2 (N22244, N22229, N21093);
and AND4 (N22245, N22222, N17676, N1070, N1355);
or OR3 (N22246, N22242, N11441, N8721);
not NOT1 (N22247, N22246);
xor XOR2 (N22248, N22240, N19820);
xor XOR2 (N22249, N22248, N3594);
xor XOR2 (N22250, N22247, N8028);
nand NAND2 (N22251, N22245, N682);
xor XOR2 (N22252, N22249, N64);
buf BUF1 (N22253, N22235);
xor XOR2 (N22254, N22253, N18017);
buf BUF1 (N22255, N22251);
buf BUF1 (N22256, N22243);
nand NAND2 (N22257, N22250, N13393);
nand NAND4 (N22258, N22252, N10534, N7520, N9390);
not NOT1 (N22259, N22255);
not NOT1 (N22260, N22239);
not NOT1 (N22261, N22259);
not NOT1 (N22262, N22258);
buf BUF1 (N22263, N22260);
nor NOR3 (N22264, N22262, N12303, N10588);
and AND4 (N22265, N22256, N15350, N10947, N20765);
or OR3 (N22266, N22244, N13062, N6151);
not NOT1 (N22267, N22261);
nor NOR2 (N22268, N22263, N14899);
nand NAND2 (N22269, N22254, N16314);
and AND3 (N22270, N22266, N6668, N13523);
not NOT1 (N22271, N22268);
and AND4 (N22272, N22267, N7049, N18490, N5031);
or OR2 (N22273, N22272, N5573);
buf BUF1 (N22274, N22270);
xor XOR2 (N22275, N22273, N13863);
xor XOR2 (N22276, N22271, N2293);
xor XOR2 (N22277, N22265, N266);
and AND3 (N22278, N22237, N20706, N2882);
and AND3 (N22279, N22275, N14940, N20616);
buf BUF1 (N22280, N22264);
nand NAND4 (N22281, N22277, N568, N4257, N3287);
nand NAND3 (N22282, N22281, N18002, N5448);
not NOT1 (N22283, N22282);
nor NOR2 (N22284, N22283, N21879);
or OR2 (N22285, N22274, N17054);
or OR4 (N22286, N22278, N632, N20415, N10118);
or OR3 (N22287, N22228, N19802, N521);
not NOT1 (N22288, N22287);
xor XOR2 (N22289, N22279, N13939);
xor XOR2 (N22290, N22225, N6277);
buf BUF1 (N22291, N22269);
or OR2 (N22292, N22286, N6444);
and AND4 (N22293, N22292, N18126, N16005, N11227);
nor NOR3 (N22294, N22289, N21431, N570);
or OR2 (N22295, N22294, N13146);
xor XOR2 (N22296, N22288, N9802);
xor XOR2 (N22297, N22284, N18115);
nand NAND4 (N22298, N22295, N4582, N4015, N14838);
and AND4 (N22299, N22298, N6356, N3243, N18373);
nor NOR4 (N22300, N22291, N6278, N21048, N3403);
and AND3 (N22301, N22293, N177, N7024);
nand NAND2 (N22302, N22296, N21388);
xor XOR2 (N22303, N22285, N20852);
not NOT1 (N22304, N22300);
nand NAND2 (N22305, N22257, N10399);
buf BUF1 (N22306, N22297);
xor XOR2 (N22307, N22276, N21197);
nor NOR3 (N22308, N22299, N4267, N2135);
nor NOR3 (N22309, N22307, N18002, N8634);
nand NAND3 (N22310, N22305, N9211, N7421);
xor XOR2 (N22311, N22304, N7446);
and AND4 (N22312, N22290, N9317, N20804, N19127);
nor NOR4 (N22313, N22310, N20485, N17782, N18592);
buf BUF1 (N22314, N22302);
or OR3 (N22315, N22303, N2724, N14801);
nor NOR2 (N22316, N22301, N1647);
not NOT1 (N22317, N22280);
xor XOR2 (N22318, N22313, N4095);
xor XOR2 (N22319, N22312, N9246);
nand NAND4 (N22320, N22316, N13219, N3367, N22242);
not NOT1 (N22321, N22320);
xor XOR2 (N22322, N22319, N6538);
not NOT1 (N22323, N22306);
and AND3 (N22324, N22315, N15684, N17778);
and AND4 (N22325, N22308, N17886, N12192, N5973);
and AND3 (N22326, N22314, N12999, N19553);
buf BUF1 (N22327, N22317);
not NOT1 (N22328, N22318);
or OR2 (N22329, N22311, N9676);
not NOT1 (N22330, N22329);
not NOT1 (N22331, N22309);
nand NAND4 (N22332, N22322, N17808, N4093, N5623);
not NOT1 (N22333, N22327);
or OR3 (N22334, N22328, N8716, N3104);
nor NOR2 (N22335, N22323, N20396);
buf BUF1 (N22336, N22334);
nor NOR2 (N22337, N22335, N943);
and AND4 (N22338, N22332, N22243, N8056, N12453);
or OR4 (N22339, N22336, N15785, N15016, N5664);
xor XOR2 (N22340, N22324, N10074);
xor XOR2 (N22341, N22339, N20189);
not NOT1 (N22342, N22331);
not NOT1 (N22343, N22337);
nor NOR4 (N22344, N22330, N4638, N5006, N9259);
xor XOR2 (N22345, N22333, N2702);
xor XOR2 (N22346, N22341, N16994);
or OR2 (N22347, N22321, N18436);
or OR2 (N22348, N22344, N754);
nor NOR2 (N22349, N22340, N7122);
buf BUF1 (N22350, N22346);
nor NOR2 (N22351, N22348, N10845);
xor XOR2 (N22352, N22343, N4894);
not NOT1 (N22353, N22352);
not NOT1 (N22354, N22342);
nor NOR3 (N22355, N22354, N11419, N2029);
not NOT1 (N22356, N22353);
not NOT1 (N22357, N22325);
or OR2 (N22358, N22326, N303);
not NOT1 (N22359, N22356);
not NOT1 (N22360, N22349);
buf BUF1 (N22361, N22351);
xor XOR2 (N22362, N22347, N19925);
nor NOR2 (N22363, N22345, N11950);
or OR4 (N22364, N22361, N14299, N16687, N12196);
nor NOR4 (N22365, N22350, N1426, N1350, N20384);
not NOT1 (N22366, N22355);
and AND3 (N22367, N22362, N16728, N115);
nor NOR3 (N22368, N22359, N3351, N6223);
or OR3 (N22369, N22368, N18102, N9802);
not NOT1 (N22370, N22366);
nand NAND2 (N22371, N22360, N12566);
xor XOR2 (N22372, N22365, N8609);
xor XOR2 (N22373, N22371, N21994);
nand NAND4 (N22374, N22372, N4516, N13872, N5801);
or OR4 (N22375, N22374, N20901, N3459, N21735);
not NOT1 (N22376, N22375);
not NOT1 (N22377, N22358);
buf BUF1 (N22378, N22338);
and AND3 (N22379, N22370, N18950, N6407);
buf BUF1 (N22380, N22357);
and AND2 (N22381, N22378, N21563);
nand NAND3 (N22382, N22369, N4571, N16617);
buf BUF1 (N22383, N22373);
not NOT1 (N22384, N22376);
nand NAND2 (N22385, N22379, N4900);
not NOT1 (N22386, N22383);
nand NAND3 (N22387, N22367, N15149, N9204);
xor XOR2 (N22388, N22380, N5461);
xor XOR2 (N22389, N22387, N11221);
not NOT1 (N22390, N22377);
or OR2 (N22391, N22381, N18972);
buf BUF1 (N22392, N22385);
and AND2 (N22393, N22382, N7115);
or OR4 (N22394, N22384, N20954, N21150, N21934);
or OR2 (N22395, N22390, N1970);
and AND4 (N22396, N22395, N8085, N17965, N7180);
or OR3 (N22397, N22386, N14992, N14894);
nor NOR2 (N22398, N22364, N15930);
nor NOR4 (N22399, N22388, N16894, N700, N16574);
xor XOR2 (N22400, N22399, N9875);
xor XOR2 (N22401, N22396, N19300);
buf BUF1 (N22402, N22398);
not NOT1 (N22403, N22402);
and AND4 (N22404, N22401, N20610, N12974, N19379);
nor NOR4 (N22405, N22393, N18040, N1335, N10465);
not NOT1 (N22406, N22400);
nor NOR4 (N22407, N22403, N4428, N1176, N11763);
nand NAND4 (N22408, N22397, N9271, N16945, N12219);
nand NAND2 (N22409, N22405, N8766);
not NOT1 (N22410, N22408);
or OR3 (N22411, N22363, N17803, N16782);
nand NAND2 (N22412, N22404, N21851);
buf BUF1 (N22413, N22407);
xor XOR2 (N22414, N22412, N8205);
nor NOR2 (N22415, N22394, N16762);
xor XOR2 (N22416, N22409, N9335);
nor NOR2 (N22417, N22413, N9074);
not NOT1 (N22418, N22389);
buf BUF1 (N22419, N22417);
xor XOR2 (N22420, N22410, N9976);
and AND2 (N22421, N22419, N5828);
or OR3 (N22422, N22418, N8354, N12549);
and AND3 (N22423, N22421, N11456, N21065);
and AND2 (N22424, N22422, N3951);
nor NOR3 (N22425, N22414, N5486, N8441);
or OR2 (N22426, N22416, N5138);
not NOT1 (N22427, N22420);
nor NOR4 (N22428, N22423, N14724, N12253, N19971);
and AND4 (N22429, N22427, N8520, N10682, N20724);
nor NOR2 (N22430, N22426, N14988);
not NOT1 (N22431, N22429);
and AND3 (N22432, N22430, N4094, N20600);
not NOT1 (N22433, N22406);
and AND3 (N22434, N22428, N3643, N5247);
buf BUF1 (N22435, N22433);
xor XOR2 (N22436, N22392, N9277);
xor XOR2 (N22437, N22432, N2264);
xor XOR2 (N22438, N22436, N13726);
nand NAND4 (N22439, N22431, N4427, N12390, N17329);
or OR2 (N22440, N22425, N10926);
or OR3 (N22441, N22434, N4917, N1218);
nand NAND4 (N22442, N22438, N9342, N564, N5951);
not NOT1 (N22443, N22411);
buf BUF1 (N22444, N22391);
or OR3 (N22445, N22440, N588, N561);
nand NAND4 (N22446, N22442, N2682, N904, N16007);
or OR2 (N22447, N22437, N4683);
buf BUF1 (N22448, N22446);
nand NAND3 (N22449, N22443, N9585, N15296);
not NOT1 (N22450, N22449);
buf BUF1 (N22451, N22441);
nor NOR3 (N22452, N22424, N4016, N20655);
nor NOR2 (N22453, N22452, N10197);
nor NOR2 (N22454, N22445, N18883);
not NOT1 (N22455, N22454);
not NOT1 (N22456, N22439);
xor XOR2 (N22457, N22444, N6613);
not NOT1 (N22458, N22448);
nand NAND3 (N22459, N22451, N19855, N19635);
nand NAND4 (N22460, N22435, N18260, N5076, N12037);
and AND4 (N22461, N22455, N14902, N19388, N11821);
nand NAND3 (N22462, N22460, N5408, N4115);
or OR2 (N22463, N22461, N11177);
buf BUF1 (N22464, N22415);
or OR4 (N22465, N22456, N3477, N7936, N20878);
nor NOR4 (N22466, N22463, N5246, N16948, N3309);
buf BUF1 (N22467, N22458);
not NOT1 (N22468, N22457);
buf BUF1 (N22469, N22467);
xor XOR2 (N22470, N22453, N8488);
buf BUF1 (N22471, N22447);
xor XOR2 (N22472, N22471, N15057);
and AND3 (N22473, N22469, N11685, N19014);
and AND3 (N22474, N22450, N15048, N17934);
and AND2 (N22475, N22466, N14272);
nor NOR4 (N22476, N22465, N5699, N16065, N7224);
buf BUF1 (N22477, N22475);
xor XOR2 (N22478, N22476, N3282);
buf BUF1 (N22479, N22468);
nor NOR3 (N22480, N22474, N3200, N106);
nand NAND3 (N22481, N22462, N12307, N4815);
and AND2 (N22482, N22479, N19285);
nand NAND3 (N22483, N22464, N9601, N3576);
buf BUF1 (N22484, N22470);
xor XOR2 (N22485, N22477, N384);
or OR3 (N22486, N22482, N12079, N98);
nand NAND3 (N22487, N22483, N5144, N18624);
or OR2 (N22488, N22486, N17192);
buf BUF1 (N22489, N22488);
or OR4 (N22490, N22487, N19811, N6499, N10683);
xor XOR2 (N22491, N22473, N4494);
nor NOR2 (N22492, N22481, N15663);
nand NAND2 (N22493, N22480, N10982);
or OR2 (N22494, N22493, N4127);
nor NOR3 (N22495, N22484, N2931, N10249);
and AND3 (N22496, N22495, N7019, N14278);
not NOT1 (N22497, N22485);
xor XOR2 (N22498, N22494, N9242);
nand NAND4 (N22499, N22492, N13989, N10994, N502);
nor NOR2 (N22500, N22459, N19511);
not NOT1 (N22501, N22489);
buf BUF1 (N22502, N22498);
nor NOR3 (N22503, N22496, N3905, N5155);
nand NAND2 (N22504, N22478, N4875);
nor NOR2 (N22505, N22499, N13877);
and AND3 (N22506, N22497, N15301, N14977);
and AND3 (N22507, N22490, N19320, N16744);
nor NOR4 (N22508, N22503, N20240, N11991, N21065);
buf BUF1 (N22509, N22505);
and AND3 (N22510, N22504, N22499, N11298);
nor NOR2 (N22511, N22510, N2527);
nor NOR4 (N22512, N22507, N1040, N4175, N17679);
and AND4 (N22513, N22502, N15804, N16354, N10619);
buf BUF1 (N22514, N22472);
or OR2 (N22515, N22513, N8123);
and AND4 (N22516, N22512, N15666, N6789, N8751);
xor XOR2 (N22517, N22501, N9236);
buf BUF1 (N22518, N22511);
xor XOR2 (N22519, N22514, N10329);
xor XOR2 (N22520, N22517, N20081);
xor XOR2 (N22521, N22509, N1600);
xor XOR2 (N22522, N22520, N11372);
not NOT1 (N22523, N22518);
nand NAND2 (N22524, N22522, N2342);
nor NOR3 (N22525, N22491, N7447, N12505);
xor XOR2 (N22526, N22508, N21604);
and AND3 (N22527, N22521, N8291, N19859);
and AND3 (N22528, N22527, N14376, N833);
nor NOR3 (N22529, N22524, N6409, N11439);
xor XOR2 (N22530, N22523, N9509);
not NOT1 (N22531, N22528);
or OR2 (N22532, N22519, N9016);
or OR2 (N22533, N22531, N17575);
nand NAND2 (N22534, N22533, N13494);
or OR3 (N22535, N22516, N17279, N11162);
buf BUF1 (N22536, N22500);
buf BUF1 (N22537, N22526);
and AND3 (N22538, N22535, N11318, N21188);
nor NOR3 (N22539, N22538, N7421, N11747);
nand NAND3 (N22540, N22534, N17499, N3891);
nand NAND3 (N22541, N22530, N5162, N10879);
nor NOR4 (N22542, N22539, N20256, N17973, N16252);
and AND4 (N22543, N22541, N14396, N2597, N3380);
xor XOR2 (N22544, N22540, N16607);
buf BUF1 (N22545, N22532);
or OR2 (N22546, N22544, N1674);
xor XOR2 (N22547, N22529, N15131);
or OR4 (N22548, N22506, N12230, N17261, N14528);
nor NOR2 (N22549, N22547, N428);
xor XOR2 (N22550, N22542, N10001);
and AND2 (N22551, N22545, N19162);
or OR4 (N22552, N22550, N6405, N19069, N1599);
or OR3 (N22553, N22549, N7414, N6666);
buf BUF1 (N22554, N22551);
nand NAND4 (N22555, N22554, N6725, N6353, N14837);
nand NAND3 (N22556, N22555, N13422, N12944);
xor XOR2 (N22557, N22536, N8136);
xor XOR2 (N22558, N22543, N11370);
xor XOR2 (N22559, N22525, N7332);
nand NAND3 (N22560, N22537, N3175, N11935);
buf BUF1 (N22561, N22558);
buf BUF1 (N22562, N22515);
or OR3 (N22563, N22562, N16995, N8557);
and AND3 (N22564, N22561, N14553, N16228);
and AND3 (N22565, N22553, N21199, N13135);
nand NAND3 (N22566, N22565, N18211, N16332);
or OR4 (N22567, N22563, N18784, N16757, N17412);
and AND2 (N22568, N22546, N12883);
and AND3 (N22569, N22567, N5640, N8238);
buf BUF1 (N22570, N22556);
buf BUF1 (N22571, N22568);
xor XOR2 (N22572, N22570, N463);
nand NAND2 (N22573, N22552, N16839);
nor NOR4 (N22574, N22572, N11443, N20554, N8485);
nor NOR3 (N22575, N22557, N18139, N16254);
xor XOR2 (N22576, N22574, N11989);
and AND3 (N22577, N22575, N8508, N18013);
nor NOR2 (N22578, N22560, N1508);
not NOT1 (N22579, N22548);
nand NAND4 (N22580, N22576, N14642, N14692, N18059);
buf BUF1 (N22581, N22566);
xor XOR2 (N22582, N22573, N3536);
buf BUF1 (N22583, N22577);
buf BUF1 (N22584, N22559);
and AND3 (N22585, N22564, N8270, N12623);
nand NAND3 (N22586, N22578, N20967, N15382);
xor XOR2 (N22587, N22571, N11568);
buf BUF1 (N22588, N22582);
and AND4 (N22589, N22588, N3098, N14924, N17290);
or OR4 (N22590, N22586, N2342, N15813, N15526);
nand NAND4 (N22591, N22569, N20432, N18429, N19015);
nand NAND3 (N22592, N22579, N7630, N12872);
or OR2 (N22593, N22591, N2693);
buf BUF1 (N22594, N22590);
nand NAND3 (N22595, N22587, N11806, N8648);
not NOT1 (N22596, N22585);
buf BUF1 (N22597, N22580);
buf BUF1 (N22598, N22583);
buf BUF1 (N22599, N22594);
or OR2 (N22600, N22599, N10789);
xor XOR2 (N22601, N22600, N8643);
nand NAND4 (N22602, N22598, N1684, N15866, N12475);
xor XOR2 (N22603, N22602, N10462);
and AND2 (N22604, N22592, N554);
or OR3 (N22605, N22595, N7761, N18534);
nor NOR4 (N22606, N22601, N3553, N12853, N18800);
not NOT1 (N22607, N22604);
xor XOR2 (N22608, N22605, N17187);
xor XOR2 (N22609, N22597, N10372);
or OR3 (N22610, N22608, N7104, N20543);
buf BUF1 (N22611, N22603);
nor NOR4 (N22612, N22611, N16916, N9566, N14213);
buf BUF1 (N22613, N22609);
not NOT1 (N22614, N22607);
or OR2 (N22615, N22606, N1518);
nor NOR4 (N22616, N22584, N5009, N13862, N12080);
nor NOR3 (N22617, N22589, N11563, N9992);
or OR4 (N22618, N22596, N7246, N6198, N20537);
nor NOR3 (N22619, N22612, N14815, N1382);
xor XOR2 (N22620, N22610, N15888);
xor XOR2 (N22621, N22619, N297);
nand NAND3 (N22622, N22620, N3714, N11760);
and AND3 (N22623, N22621, N10233, N22330);
or OR2 (N22624, N22617, N10743);
nand NAND3 (N22625, N22615, N20325, N11199);
xor XOR2 (N22626, N22581, N22606);
not NOT1 (N22627, N22618);
buf BUF1 (N22628, N22613);
nand NAND4 (N22629, N22614, N18506, N16838, N14647);
not NOT1 (N22630, N22616);
buf BUF1 (N22631, N22629);
xor XOR2 (N22632, N22628, N12971);
nand NAND4 (N22633, N22593, N12217, N1868, N22363);
and AND2 (N22634, N22625, N5481);
buf BUF1 (N22635, N22630);
buf BUF1 (N22636, N22634);
xor XOR2 (N22637, N22627, N21934);
xor XOR2 (N22638, N22623, N22627);
nand NAND2 (N22639, N22637, N4970);
buf BUF1 (N22640, N22624);
xor XOR2 (N22641, N22639, N22451);
nor NOR2 (N22642, N22632, N14066);
and AND4 (N22643, N22633, N18564, N4521, N12550);
and AND2 (N22644, N22636, N22074);
nor NOR3 (N22645, N22638, N16013, N18138);
not NOT1 (N22646, N22643);
not NOT1 (N22647, N22635);
buf BUF1 (N22648, N22626);
buf BUF1 (N22649, N22642);
not NOT1 (N22650, N22622);
nor NOR2 (N22651, N22641, N17283);
or OR4 (N22652, N22650, N16755, N21462, N11474);
or OR2 (N22653, N22644, N19890);
xor XOR2 (N22654, N22648, N2422);
nand NAND4 (N22655, N22652, N1617, N17329, N16016);
buf BUF1 (N22656, N22645);
nor NOR3 (N22657, N22631, N2973, N7215);
and AND2 (N22658, N22640, N6870);
xor XOR2 (N22659, N22649, N20920);
nor NOR3 (N22660, N22655, N6774, N11365);
not NOT1 (N22661, N22660);
and AND3 (N22662, N22653, N22190, N21477);
and AND4 (N22663, N22657, N10376, N13182, N18986);
buf BUF1 (N22664, N22662);
or OR4 (N22665, N22658, N17042, N20827, N15832);
or OR4 (N22666, N22647, N6648, N8718, N406);
nand NAND2 (N22667, N22654, N9345);
nand NAND3 (N22668, N22646, N16916, N3750);
and AND4 (N22669, N22651, N506, N244, N629);
nor NOR4 (N22670, N22667, N13573, N18385, N13947);
or OR2 (N22671, N22668, N21440);
buf BUF1 (N22672, N22665);
nor NOR4 (N22673, N22669, N20759, N4588, N4719);
nand NAND4 (N22674, N22659, N4260, N17074, N8554);
nand NAND2 (N22675, N22656, N5155);
buf BUF1 (N22676, N22673);
buf BUF1 (N22677, N22664);
not NOT1 (N22678, N22670);
or OR3 (N22679, N22675, N8225, N4631);
xor XOR2 (N22680, N22671, N12401);
or OR4 (N22681, N22663, N11894, N4779, N15090);
and AND3 (N22682, N22666, N15022, N12974);
nand NAND3 (N22683, N22672, N3323, N17611);
nand NAND2 (N22684, N22679, N4348);
buf BUF1 (N22685, N22661);
not NOT1 (N22686, N22680);
and AND4 (N22687, N22674, N2189, N20247, N7694);
not NOT1 (N22688, N22682);
not NOT1 (N22689, N22688);
xor XOR2 (N22690, N22687, N1632);
not NOT1 (N22691, N22677);
or OR4 (N22692, N22683, N16579, N8640, N11870);
buf BUF1 (N22693, N22681);
nand NAND4 (N22694, N22691, N3075, N8966, N15767);
buf BUF1 (N22695, N22694);
and AND4 (N22696, N22689, N7572, N1042, N2644);
xor XOR2 (N22697, N22684, N8206);
and AND4 (N22698, N22696, N8802, N7160, N14220);
and AND4 (N22699, N22676, N2364, N8161, N17673);
or OR4 (N22700, N22695, N496, N13284, N21064);
buf BUF1 (N22701, N22690);
not NOT1 (N22702, N22697);
buf BUF1 (N22703, N22686);
not NOT1 (N22704, N22678);
nand NAND3 (N22705, N22702, N14077, N15488);
buf BUF1 (N22706, N22701);
xor XOR2 (N22707, N22705, N9053);
buf BUF1 (N22708, N22685);
or OR4 (N22709, N22692, N19976, N21373, N9537);
not NOT1 (N22710, N22698);
or OR4 (N22711, N22707, N10417, N2775, N2994);
or OR3 (N22712, N22710, N7813, N14137);
and AND2 (N22713, N22708, N6157);
xor XOR2 (N22714, N22706, N144);
nand NAND2 (N22715, N22703, N8775);
nor NOR2 (N22716, N22693, N1350);
nand NAND4 (N22717, N22713, N21302, N2974, N18780);
nor NOR3 (N22718, N22699, N4900, N11045);
xor XOR2 (N22719, N22712, N6741);
nor NOR4 (N22720, N22715, N1708, N1750, N32);
buf BUF1 (N22721, N22714);
buf BUF1 (N22722, N22711);
or OR4 (N22723, N22704, N1520, N8558, N18692);
nand NAND4 (N22724, N22716, N14843, N21430, N3908);
nand NAND4 (N22725, N22724, N15746, N13171, N16924);
nand NAND4 (N22726, N22722, N15130, N17320, N15767);
nand NAND4 (N22727, N22718, N7247, N22537, N6373);
nand NAND4 (N22728, N22727, N20539, N9115, N2448);
xor XOR2 (N22729, N22719, N21258);
xor XOR2 (N22730, N22717, N10521);
nor NOR2 (N22731, N22730, N1195);
nand NAND4 (N22732, N22720, N13327, N22127, N14591);
not NOT1 (N22733, N22731);
buf BUF1 (N22734, N22725);
nand NAND2 (N22735, N22734, N105);
buf BUF1 (N22736, N22732);
and AND2 (N22737, N22733, N1079);
and AND4 (N22738, N22736, N5228, N14638, N13032);
nor NOR4 (N22739, N22726, N1969, N22056, N9500);
and AND2 (N22740, N22737, N13509);
nor NOR4 (N22741, N22740, N8119, N715, N13953);
or OR4 (N22742, N22729, N21415, N6175, N7977);
and AND2 (N22743, N22738, N14794);
not NOT1 (N22744, N22728);
xor XOR2 (N22745, N22709, N21282);
nand NAND4 (N22746, N22744, N12746, N9469, N19569);
or OR4 (N22747, N22739, N2983, N5432, N8543);
xor XOR2 (N22748, N22721, N9388);
or OR4 (N22749, N22723, N8976, N5615, N16393);
nor NOR4 (N22750, N22747, N9976, N19760, N7863);
nor NOR4 (N22751, N22745, N5850, N7479, N2228);
nor NOR4 (N22752, N22741, N12348, N8988, N16222);
and AND2 (N22753, N22750, N9513);
buf BUF1 (N22754, N22743);
nand NAND4 (N22755, N22751, N22676, N3355, N9833);
nor NOR4 (N22756, N22700, N444, N6473, N22128);
and AND3 (N22757, N22756, N8182, N21616);
not NOT1 (N22758, N22735);
buf BUF1 (N22759, N22746);
and AND4 (N22760, N22748, N8772, N11636, N4517);
nor NOR3 (N22761, N22749, N2304, N21960);
nor NOR2 (N22762, N22759, N6752);
not NOT1 (N22763, N22753);
xor XOR2 (N22764, N22761, N7115);
buf BUF1 (N22765, N22754);
or OR2 (N22766, N22758, N22056);
xor XOR2 (N22767, N22765, N7298);
and AND4 (N22768, N22742, N10883, N12985, N1014);
not NOT1 (N22769, N22768);
xor XOR2 (N22770, N22762, N8390);
buf BUF1 (N22771, N22769);
nand NAND4 (N22772, N22763, N20821, N9833, N14295);
or OR4 (N22773, N22760, N845, N11705, N15978);
and AND2 (N22774, N22757, N14488);
nand NAND4 (N22775, N22774, N18784, N2606, N22671);
and AND2 (N22776, N22773, N3647);
xor XOR2 (N22777, N22770, N20295);
nor NOR3 (N22778, N22775, N10591, N16443);
xor XOR2 (N22779, N22771, N13773);
xor XOR2 (N22780, N22755, N16444);
xor XOR2 (N22781, N22776, N2361);
xor XOR2 (N22782, N22781, N8993);
nor NOR4 (N22783, N22779, N20183, N10767, N2618);
nand NAND2 (N22784, N22780, N20569);
nand NAND4 (N22785, N22777, N19116, N7487, N769);
or OR3 (N22786, N22782, N12662, N19294);
nor NOR2 (N22787, N22784, N20586);
nor NOR2 (N22788, N22752, N13085);
or OR4 (N22789, N22764, N3618, N20981, N7578);
buf BUF1 (N22790, N22786);
or OR2 (N22791, N22785, N172);
not NOT1 (N22792, N22778);
nor NOR3 (N22793, N22787, N6883, N16863);
and AND2 (N22794, N22766, N10474);
xor XOR2 (N22795, N22789, N4621);
or OR3 (N22796, N22783, N8744, N19264);
and AND2 (N22797, N22772, N3497);
nand NAND4 (N22798, N22794, N17983, N8704, N10571);
not NOT1 (N22799, N22767);
not NOT1 (N22800, N22793);
xor XOR2 (N22801, N22788, N20377);
not NOT1 (N22802, N22798);
buf BUF1 (N22803, N22790);
nor NOR2 (N22804, N22803, N15243);
and AND4 (N22805, N22800, N12659, N8644, N16412);
nor NOR2 (N22806, N22796, N11265);
or OR4 (N22807, N22805, N10116, N20297, N12012);
buf BUF1 (N22808, N22807);
xor XOR2 (N22809, N22808, N10847);
xor XOR2 (N22810, N22795, N12182);
and AND4 (N22811, N22799, N18152, N22609, N16797);
or OR3 (N22812, N22797, N1534, N14317);
not NOT1 (N22813, N22792);
buf BUF1 (N22814, N22801);
xor XOR2 (N22815, N22806, N552);
not NOT1 (N22816, N22811);
xor XOR2 (N22817, N22809, N3320);
and AND3 (N22818, N22816, N2173, N1823);
nor NOR2 (N22819, N22815, N7707);
not NOT1 (N22820, N22817);
not NOT1 (N22821, N22814);
and AND2 (N22822, N22818, N16903);
nand NAND4 (N22823, N22819, N6672, N21188, N16631);
and AND2 (N22824, N22822, N6259);
xor XOR2 (N22825, N22813, N8481);
and AND3 (N22826, N22821, N1035, N3831);
nand NAND3 (N22827, N22802, N17393, N3319);
or OR4 (N22828, N22825, N14342, N18626, N5507);
buf BUF1 (N22829, N22824);
and AND4 (N22830, N22804, N18384, N6205, N8247);
xor XOR2 (N22831, N22810, N7803);
or OR2 (N22832, N22830, N16765);
and AND4 (N22833, N22823, N22155, N11528, N12468);
and AND2 (N22834, N22826, N17049);
nor NOR3 (N22835, N22820, N16792, N6319);
nand NAND2 (N22836, N22791, N13343);
and AND3 (N22837, N22836, N7103, N22199);
nand NAND3 (N22838, N22833, N3890, N9863);
buf BUF1 (N22839, N22829);
and AND2 (N22840, N22827, N8267);
or OR4 (N22841, N22828, N1878, N8551, N8074);
buf BUF1 (N22842, N22835);
and AND2 (N22843, N22812, N11177);
or OR3 (N22844, N22840, N9343, N19121);
xor XOR2 (N22845, N22834, N14423);
nand NAND4 (N22846, N22844, N11348, N14933, N9630);
nand NAND3 (N22847, N22845, N12470, N22550);
or OR3 (N22848, N22841, N19185, N18978);
and AND2 (N22849, N22837, N4656);
not NOT1 (N22850, N22847);
not NOT1 (N22851, N22849);
xor XOR2 (N22852, N22831, N1100);
not NOT1 (N22853, N22852);
and AND4 (N22854, N22838, N3582, N15503, N4868);
not NOT1 (N22855, N22854);
and AND2 (N22856, N22846, N19242);
not NOT1 (N22857, N22853);
or OR2 (N22858, N22848, N6390);
buf BUF1 (N22859, N22850);
nor NOR3 (N22860, N22855, N17270, N8156);
not NOT1 (N22861, N22851);
xor XOR2 (N22862, N22839, N6764);
or OR4 (N22863, N22858, N16354, N3697, N7217);
and AND3 (N22864, N22863, N17372, N14417);
buf BUF1 (N22865, N22856);
and AND4 (N22866, N22832, N12881, N9361, N8387);
and AND2 (N22867, N22866, N6209);
xor XOR2 (N22868, N22867, N8416);
xor XOR2 (N22869, N22857, N5449);
or OR3 (N22870, N22842, N4077, N15386);
nand NAND2 (N22871, N22865, N13107);
buf BUF1 (N22872, N22864);
nand NAND3 (N22873, N22860, N18627, N15968);
buf BUF1 (N22874, N22859);
not NOT1 (N22875, N22873);
xor XOR2 (N22876, N22875, N16634);
or OR4 (N22877, N22869, N7025, N14436, N23);
and AND3 (N22878, N22861, N22340, N19002);
nor NOR4 (N22879, N22862, N13033, N11133, N19872);
nor NOR4 (N22880, N22872, N3002, N1155, N1646);
buf BUF1 (N22881, N22876);
and AND3 (N22882, N22878, N3739, N17589);
not NOT1 (N22883, N22880);
buf BUF1 (N22884, N22871);
or OR4 (N22885, N22843, N9178, N18533, N9390);
nand NAND2 (N22886, N22884, N975);
nand NAND4 (N22887, N22883, N19543, N8501, N17988);
xor XOR2 (N22888, N22885, N9102);
nor NOR2 (N22889, N22877, N19364);
nor NOR2 (N22890, N22887, N8566);
nor NOR4 (N22891, N22881, N16470, N18772, N1105);
nand NAND3 (N22892, N22886, N11834, N22680);
nand NAND3 (N22893, N22882, N20677, N16243);
buf BUF1 (N22894, N22868);
nor NOR3 (N22895, N22889, N5468, N6129);
and AND4 (N22896, N22895, N10424, N16903, N2543);
nand NAND4 (N22897, N22879, N16470, N16573, N16847);
nor NOR2 (N22898, N22896, N9859);
buf BUF1 (N22899, N22888);
and AND4 (N22900, N22893, N4243, N16988, N16529);
buf BUF1 (N22901, N22894);
xor XOR2 (N22902, N22899, N18610);
or OR4 (N22903, N22898, N14912, N6572, N16630);
nand NAND4 (N22904, N22892, N20834, N9212, N10704);
nor NOR4 (N22905, N22902, N12977, N426, N10399);
or OR2 (N22906, N22901, N8674);
not NOT1 (N22907, N22905);
xor XOR2 (N22908, N22874, N15163);
nand NAND4 (N22909, N22900, N16383, N9979, N21842);
nand NAND4 (N22910, N22907, N6528, N9419, N15231);
xor XOR2 (N22911, N22910, N1963);
or OR2 (N22912, N22891, N10922);
and AND4 (N22913, N22903, N8459, N15425, N14108);
buf BUF1 (N22914, N22908);
or OR2 (N22915, N22912, N1708);
nand NAND4 (N22916, N22915, N16895, N9046, N4182);
nor NOR3 (N22917, N22909, N4005, N14904);
buf BUF1 (N22918, N22897);
not NOT1 (N22919, N22890);
nor NOR2 (N22920, N22904, N5723);
and AND2 (N22921, N22917, N8987);
not NOT1 (N22922, N22918);
and AND2 (N22923, N22906, N6712);
nor NOR3 (N22924, N22870, N15176, N7268);
nor NOR2 (N22925, N22913, N4070);
nand NAND4 (N22926, N22923, N8163, N6069, N21809);
or OR2 (N22927, N22914, N5946);
and AND3 (N22928, N22911, N2775, N22047);
nand NAND3 (N22929, N22926, N11957, N5041);
xor XOR2 (N22930, N22925, N7993);
buf BUF1 (N22931, N22916);
nor NOR3 (N22932, N22919, N19299, N9324);
xor XOR2 (N22933, N22921, N2846);
buf BUF1 (N22934, N22933);
and AND3 (N22935, N22922, N19404, N4043);
xor XOR2 (N22936, N22931, N16050);
and AND3 (N22937, N22936, N10832, N11516);
nand NAND4 (N22938, N22934, N5480, N12778, N1726);
nor NOR3 (N22939, N22935, N3874, N6492);
not NOT1 (N22940, N22929);
buf BUF1 (N22941, N22939);
or OR2 (N22942, N22924, N5483);
xor XOR2 (N22943, N22938, N22282);
buf BUF1 (N22944, N22942);
and AND4 (N22945, N22930, N20656, N14727, N14027);
xor XOR2 (N22946, N22920, N15003);
not NOT1 (N22947, N22940);
not NOT1 (N22948, N22928);
xor XOR2 (N22949, N22943, N4324);
nand NAND2 (N22950, N22946, N19176);
or OR4 (N22951, N22950, N22251, N18189, N16671);
nor NOR2 (N22952, N22932, N20495);
not NOT1 (N22953, N22948);
buf BUF1 (N22954, N22945);
or OR4 (N22955, N22944, N17493, N17543, N22897);
not NOT1 (N22956, N22951);
xor XOR2 (N22957, N22955, N13023);
xor XOR2 (N22958, N22956, N13469);
or OR2 (N22959, N22958, N17335);
not NOT1 (N22960, N22941);
nor NOR2 (N22961, N22954, N9613);
xor XOR2 (N22962, N22927, N21796);
or OR3 (N22963, N22962, N20740, N19453);
and AND2 (N22964, N22949, N3891);
not NOT1 (N22965, N22953);
buf BUF1 (N22966, N22961);
xor XOR2 (N22967, N22959, N16930);
xor XOR2 (N22968, N22963, N5672);
or OR4 (N22969, N22964, N6071, N8745, N10148);
and AND4 (N22970, N22969, N17935, N10560, N22007);
xor XOR2 (N22971, N22952, N18831);
nor NOR4 (N22972, N22968, N7324, N2795, N7338);
xor XOR2 (N22973, N22965, N18773);
xor XOR2 (N22974, N22947, N13605);
and AND4 (N22975, N22957, N15494, N20903, N12001);
buf BUF1 (N22976, N22974);
and AND3 (N22977, N22972, N2523, N21869);
xor XOR2 (N22978, N22971, N8482);
nor NOR3 (N22979, N22967, N19209, N22000);
nand NAND2 (N22980, N22970, N7114);
or OR4 (N22981, N22966, N5338, N17359, N19930);
nor NOR4 (N22982, N22973, N5769, N12427, N19106);
xor XOR2 (N22983, N22979, N19351);
nor NOR2 (N22984, N22960, N17846);
nor NOR4 (N22985, N22983, N2821, N11214, N15360);
and AND4 (N22986, N22980, N19279, N7674, N6468);
not NOT1 (N22987, N22937);
nand NAND2 (N22988, N22978, N1560);
and AND3 (N22989, N22985, N9917, N14365);
xor XOR2 (N22990, N22982, N6213);
and AND2 (N22991, N22986, N361);
xor XOR2 (N22992, N22975, N16133);
not NOT1 (N22993, N22984);
not NOT1 (N22994, N22977);
nor NOR2 (N22995, N22988, N18090);
nor NOR2 (N22996, N22990, N15633);
not NOT1 (N22997, N22996);
buf BUF1 (N22998, N22992);
nand NAND3 (N22999, N22991, N2019, N20331);
nor NOR4 (N23000, N22995, N22482, N1080, N3809);
or OR3 (N23001, N22989, N22330, N8825);
or OR3 (N23002, N23001, N1937, N15474);
nand NAND2 (N23003, N22987, N22681);
xor XOR2 (N23004, N22994, N19933);
or OR4 (N23005, N23004, N17912, N18797, N13220);
buf BUF1 (N23006, N22976);
and AND4 (N23007, N23005, N20428, N2023, N2717);
xor XOR2 (N23008, N22998, N16316);
xor XOR2 (N23009, N23003, N14412);
and AND4 (N23010, N23009, N7733, N3911, N13221);
xor XOR2 (N23011, N23002, N3705);
and AND4 (N23012, N22993, N16382, N6266, N2618);
nor NOR4 (N23013, N23012, N8490, N2209, N11772);
buf BUF1 (N23014, N23010);
buf BUF1 (N23015, N22997);
xor XOR2 (N23016, N23014, N9515);
buf BUF1 (N23017, N23007);
or OR3 (N23018, N23013, N5834, N21952);
nand NAND2 (N23019, N23016, N3075);
nand NAND3 (N23020, N23017, N6038, N8012);
not NOT1 (N23021, N22981);
xor XOR2 (N23022, N22999, N21304);
nand NAND2 (N23023, N23006, N16110);
and AND4 (N23024, N23008, N12483, N12329, N19527);
nor NOR2 (N23025, N23011, N20274);
xor XOR2 (N23026, N23022, N17135);
not NOT1 (N23027, N23000);
xor XOR2 (N23028, N23024, N2154);
nor NOR2 (N23029, N23027, N19667);
and AND4 (N23030, N23023, N22072, N13517, N5077);
nor NOR3 (N23031, N23029, N18369, N10785);
or OR3 (N23032, N23030, N11314, N13066);
and AND4 (N23033, N23020, N9987, N19294, N5905);
or OR4 (N23034, N23031, N2030, N9129, N6189);
not NOT1 (N23035, N23026);
xor XOR2 (N23036, N23021, N4774);
buf BUF1 (N23037, N23019);
xor XOR2 (N23038, N23034, N2194);
or OR3 (N23039, N23025, N18096, N13435);
buf BUF1 (N23040, N23036);
and AND2 (N23041, N23032, N15936);
nand NAND3 (N23042, N23040, N19405, N18613);
and AND3 (N23043, N23033, N18505, N1039);
xor XOR2 (N23044, N23035, N4578);
nor NOR2 (N23045, N23041, N19025);
nor NOR3 (N23046, N23039, N9660, N16950);
nand NAND3 (N23047, N23038, N6844, N2768);
nor NOR4 (N23048, N23044, N15837, N14200, N5036);
not NOT1 (N23049, N23015);
or OR2 (N23050, N23048, N17923);
nand NAND4 (N23051, N23028, N1688, N21486, N920);
and AND3 (N23052, N23050, N5336, N16850);
xor XOR2 (N23053, N23042, N916);
and AND2 (N23054, N23047, N21827);
and AND2 (N23055, N23049, N17851);
not NOT1 (N23056, N23051);
xor XOR2 (N23057, N23043, N13533);
buf BUF1 (N23058, N23053);
xor XOR2 (N23059, N23046, N6250);
xor XOR2 (N23060, N23057, N13538);
nor NOR4 (N23061, N23054, N4382, N10291, N10477);
nand NAND4 (N23062, N23055, N21357, N2790, N18580);
nand NAND2 (N23063, N23060, N6570);
xor XOR2 (N23064, N23018, N11745);
xor XOR2 (N23065, N23037, N18255);
not NOT1 (N23066, N23056);
and AND3 (N23067, N23052, N8931, N22439);
buf BUF1 (N23068, N23066);
buf BUF1 (N23069, N23059);
or OR4 (N23070, N23045, N7567, N19957, N18654);
or OR2 (N23071, N23065, N13258);
and AND4 (N23072, N23063, N9202, N9578, N3185);
or OR3 (N23073, N23062, N12808, N22444);
nand NAND3 (N23074, N23064, N5722, N18841);
buf BUF1 (N23075, N23068);
and AND2 (N23076, N23058, N13091);
xor XOR2 (N23077, N23070, N1326);
buf BUF1 (N23078, N23074);
and AND2 (N23079, N23077, N14197);
not NOT1 (N23080, N23075);
and AND3 (N23081, N23071, N13993, N13715);
nor NOR4 (N23082, N23079, N21187, N5738, N15972);
buf BUF1 (N23083, N23061);
xor XOR2 (N23084, N23067, N21578);
buf BUF1 (N23085, N23082);
nor NOR4 (N23086, N23083, N2802, N9101, N18414);
not NOT1 (N23087, N23073);
nor NOR4 (N23088, N23084, N6523, N880, N10435);
nand NAND2 (N23089, N23080, N7734);
or OR2 (N23090, N23078, N21319);
not NOT1 (N23091, N23076);
or OR3 (N23092, N23088, N6588, N8455);
and AND2 (N23093, N23087, N1211);
not NOT1 (N23094, N23089);
buf BUF1 (N23095, N23093);
buf BUF1 (N23096, N23090);
nand NAND2 (N23097, N23072, N397);
buf BUF1 (N23098, N23092);
not NOT1 (N23099, N23098);
nand NAND2 (N23100, N23096, N9980);
buf BUF1 (N23101, N23069);
buf BUF1 (N23102, N23091);
not NOT1 (N23103, N23095);
xor XOR2 (N23104, N23100, N14343);
nand NAND2 (N23105, N23094, N22171);
not NOT1 (N23106, N23105);
buf BUF1 (N23107, N23104);
nor NOR4 (N23108, N23101, N6069, N7949, N3347);
nand NAND2 (N23109, N23081, N21029);
nand NAND4 (N23110, N23102, N3141, N8953, N15567);
and AND3 (N23111, N23085, N5616, N14592);
and AND2 (N23112, N23108, N22820);
or OR4 (N23113, N23109, N1937, N7382, N13353);
buf BUF1 (N23114, N23113);
and AND2 (N23115, N23099, N5078);
or OR3 (N23116, N23114, N1508, N14358);
buf BUF1 (N23117, N23107);
not NOT1 (N23118, N23112);
or OR3 (N23119, N23097, N5703, N2709);
nand NAND4 (N23120, N23111, N7707, N8738, N9340);
not NOT1 (N23121, N23106);
or OR4 (N23122, N23103, N10228, N6754, N19915);
buf BUF1 (N23123, N23122);
nor NOR3 (N23124, N23123, N10643, N3923);
and AND3 (N23125, N23124, N2734, N2022);
or OR2 (N23126, N23125, N4270);
nor NOR4 (N23127, N23119, N22618, N6037, N2210);
or OR2 (N23128, N23127, N9524);
nor NOR3 (N23129, N23115, N2007, N2368);
or OR3 (N23130, N23117, N7680, N11242);
and AND4 (N23131, N23110, N35, N21367, N14833);
nor NOR3 (N23132, N23086, N22510, N6443);
not NOT1 (N23133, N23121);
buf BUF1 (N23134, N23126);
not NOT1 (N23135, N23128);
not NOT1 (N23136, N23135);
or OR3 (N23137, N23130, N9952, N9800);
or OR4 (N23138, N23133, N12935, N8372, N8349);
nor NOR3 (N23139, N23132, N6311, N20682);
nand NAND4 (N23140, N23120, N6108, N2673, N18186);
buf BUF1 (N23141, N23134);
and AND2 (N23142, N23118, N4198);
buf BUF1 (N23143, N23137);
xor XOR2 (N23144, N23129, N15140);
and AND3 (N23145, N23138, N21579, N4959);
and AND3 (N23146, N23140, N687, N4426);
buf BUF1 (N23147, N23139);
xor XOR2 (N23148, N23142, N295);
and AND3 (N23149, N23143, N17962, N13188);
or OR2 (N23150, N23147, N4381);
nor NOR4 (N23151, N23145, N1913, N11982, N10198);
nand NAND2 (N23152, N23144, N18549);
not NOT1 (N23153, N23149);
not NOT1 (N23154, N23131);
nand NAND3 (N23155, N23154, N20434, N4896);
buf BUF1 (N23156, N23141);
xor XOR2 (N23157, N23156, N10378);
buf BUF1 (N23158, N23150);
buf BUF1 (N23159, N23146);
nor NOR4 (N23160, N23116, N20612, N15012, N9203);
xor XOR2 (N23161, N23152, N14527);
buf BUF1 (N23162, N23151);
nor NOR4 (N23163, N23153, N3372, N2410, N21061);
nand NAND3 (N23164, N23157, N2470, N2149);
buf BUF1 (N23165, N23164);
buf BUF1 (N23166, N23165);
or OR4 (N23167, N23159, N18196, N1888, N18194);
and AND3 (N23168, N23162, N10366, N10383);
and AND2 (N23169, N23167, N13887);
buf BUF1 (N23170, N23163);
nand NAND3 (N23171, N23148, N15143, N10910);
not NOT1 (N23172, N23160);
or OR2 (N23173, N23169, N17338);
nand NAND2 (N23174, N23155, N509);
or OR3 (N23175, N23171, N4492, N134);
or OR2 (N23176, N23136, N4247);
nand NAND3 (N23177, N23176, N16066, N3774);
and AND3 (N23178, N23174, N5845, N17101);
nor NOR4 (N23179, N23177, N11350, N4783, N8837);
or OR4 (N23180, N23179, N3115, N17201, N13185);
buf BUF1 (N23181, N23172);
or OR3 (N23182, N23161, N1377, N13873);
and AND2 (N23183, N23173, N18161);
buf BUF1 (N23184, N23170);
or OR3 (N23185, N23184, N10855, N632);
buf BUF1 (N23186, N23166);
buf BUF1 (N23187, N23178);
and AND4 (N23188, N23168, N22948, N19735, N6761);
not NOT1 (N23189, N23185);
buf BUF1 (N23190, N23182);
or OR2 (N23191, N23180, N9901);
nand NAND3 (N23192, N23158, N2322, N11638);
buf BUF1 (N23193, N23189);
nor NOR3 (N23194, N23192, N20085, N19550);
nand NAND2 (N23195, N23194, N350);
or OR4 (N23196, N23190, N10471, N19956, N17158);
nand NAND2 (N23197, N23188, N2655);
xor XOR2 (N23198, N23183, N11243);
xor XOR2 (N23199, N23193, N17813);
nor NOR2 (N23200, N23198, N21410);
not NOT1 (N23201, N23197);
nand NAND4 (N23202, N23186, N16800, N12764, N8170);
or OR4 (N23203, N23181, N697, N19170, N14636);
nand NAND3 (N23204, N23195, N2562, N11975);
xor XOR2 (N23205, N23200, N21531);
or OR2 (N23206, N23191, N261);
not NOT1 (N23207, N23199);
and AND3 (N23208, N23206, N489, N20);
and AND3 (N23209, N23202, N3326, N16388);
xor XOR2 (N23210, N23205, N13371);
or OR4 (N23211, N23196, N19933, N8203, N17771);
not NOT1 (N23212, N23210);
buf BUF1 (N23213, N23187);
xor XOR2 (N23214, N23212, N23121);
and AND4 (N23215, N23175, N4926, N3173, N6226);
nand NAND4 (N23216, N23207, N5483, N1970, N9090);
and AND4 (N23217, N23208, N1201, N1106, N20007);
nand NAND2 (N23218, N23204, N16967);
xor XOR2 (N23219, N23214, N834);
not NOT1 (N23220, N23216);
or OR4 (N23221, N23209, N14942, N21679, N8648);
or OR4 (N23222, N23211, N11286, N22661, N13102);
nor NOR3 (N23223, N23218, N8109, N22847);
and AND3 (N23224, N23203, N17075, N7774);
nand NAND2 (N23225, N23201, N8913);
or OR3 (N23226, N23215, N13984, N6010);
nor NOR3 (N23227, N23222, N17746, N17337);
nand NAND4 (N23228, N23221, N23104, N17965, N21144);
buf BUF1 (N23229, N23224);
buf BUF1 (N23230, N23226);
buf BUF1 (N23231, N23227);
not NOT1 (N23232, N23217);
not NOT1 (N23233, N23230);
and AND4 (N23234, N23225, N17789, N11851, N15981);
and AND4 (N23235, N23228, N4362, N11444, N17064);
or OR3 (N23236, N23229, N20108, N10458);
xor XOR2 (N23237, N23235, N22095);
or OR2 (N23238, N23220, N14658);
not NOT1 (N23239, N23232);
not NOT1 (N23240, N23233);
or OR3 (N23241, N23239, N22908, N14588);
xor XOR2 (N23242, N23213, N5133);
or OR2 (N23243, N23223, N12795);
nand NAND2 (N23244, N23234, N11695);
or OR3 (N23245, N23240, N7149, N18376);
xor XOR2 (N23246, N23236, N3059);
nor NOR2 (N23247, N23243, N1669);
xor XOR2 (N23248, N23247, N21591);
not NOT1 (N23249, N23219);
nand NAND2 (N23250, N23246, N15790);
not NOT1 (N23251, N23248);
not NOT1 (N23252, N23250);
nor NOR2 (N23253, N23231, N5642);
buf BUF1 (N23254, N23249);
or OR2 (N23255, N23254, N18572);
nor NOR3 (N23256, N23242, N16287, N3673);
and AND2 (N23257, N23255, N16887);
and AND2 (N23258, N23245, N4323);
nor NOR2 (N23259, N23258, N4093);
xor XOR2 (N23260, N23259, N1046);
or OR2 (N23261, N23237, N17941);
xor XOR2 (N23262, N23257, N13004);
nor NOR4 (N23263, N23253, N13616, N17040, N878);
buf BUF1 (N23264, N23252);
or OR2 (N23265, N23261, N19750);
xor XOR2 (N23266, N23262, N3984);
xor XOR2 (N23267, N23260, N4525);
or OR3 (N23268, N23251, N16551, N172);
buf BUF1 (N23269, N23266);
nand NAND2 (N23270, N23241, N4290);
xor XOR2 (N23271, N23238, N1160);
nand NAND4 (N23272, N23244, N4825, N15037, N5198);
nor NOR4 (N23273, N23271, N19751, N751, N15034);
nor NOR3 (N23274, N23269, N14447, N19132);
buf BUF1 (N23275, N23274);
nor NOR3 (N23276, N23263, N1221, N7638);
nand NAND4 (N23277, N23264, N9184, N16798, N12211);
nand NAND2 (N23278, N23273, N5404);
or OR2 (N23279, N23275, N2040);
not NOT1 (N23280, N23267);
not NOT1 (N23281, N23278);
buf BUF1 (N23282, N23256);
nor NOR3 (N23283, N23265, N13579, N12122);
xor XOR2 (N23284, N23279, N14662);
and AND2 (N23285, N23282, N20124);
not NOT1 (N23286, N23283);
nand NAND3 (N23287, N23285, N15420, N19735);
nor NOR4 (N23288, N23281, N6895, N3048, N7208);
not NOT1 (N23289, N23280);
or OR4 (N23290, N23268, N12346, N16916, N6090);
nand NAND4 (N23291, N23287, N11521, N1637, N2160);
xor XOR2 (N23292, N23276, N20480);
xor XOR2 (N23293, N23284, N11498);
or OR3 (N23294, N23288, N22011, N13878);
and AND4 (N23295, N23277, N8911, N19953, N11026);
xor XOR2 (N23296, N23290, N15337);
buf BUF1 (N23297, N23295);
nor NOR2 (N23298, N23297, N3308);
nand NAND4 (N23299, N23296, N5341, N2964, N1103);
nand NAND2 (N23300, N23272, N17571);
buf BUF1 (N23301, N23298);
buf BUF1 (N23302, N23291);
not NOT1 (N23303, N23300);
xor XOR2 (N23304, N23289, N12993);
and AND3 (N23305, N23304, N18205, N14816);
xor XOR2 (N23306, N23292, N15101);
not NOT1 (N23307, N23270);
xor XOR2 (N23308, N23305, N22233);
buf BUF1 (N23309, N23306);
nor NOR3 (N23310, N23301, N3068, N11487);
nand NAND2 (N23311, N23299, N12107);
nor NOR2 (N23312, N23286, N9862);
xor XOR2 (N23313, N23303, N17356);
nor NOR2 (N23314, N23309, N9153);
not NOT1 (N23315, N23308);
nand NAND2 (N23316, N23310, N16317);
not NOT1 (N23317, N23293);
nor NOR4 (N23318, N23316, N16035, N3691, N5356);
not NOT1 (N23319, N23318);
nand NAND2 (N23320, N23315, N2019);
and AND3 (N23321, N23317, N3551, N12469);
xor XOR2 (N23322, N23313, N19283);
nor NOR4 (N23323, N23312, N2177, N4657, N17528);
buf BUF1 (N23324, N23320);
not NOT1 (N23325, N23314);
and AND2 (N23326, N23311, N22239);
and AND3 (N23327, N23294, N9161, N10914);
or OR2 (N23328, N23327, N10927);
not NOT1 (N23329, N23323);
nor NOR4 (N23330, N23322, N21896, N19157, N498);
and AND2 (N23331, N23302, N10502);
buf BUF1 (N23332, N23324);
nand NAND3 (N23333, N23330, N22875, N8851);
and AND2 (N23334, N23307, N18761);
xor XOR2 (N23335, N23331, N11358);
buf BUF1 (N23336, N23334);
nor NOR2 (N23337, N23321, N12498);
xor XOR2 (N23338, N23337, N18856);
not NOT1 (N23339, N23338);
not NOT1 (N23340, N23335);
nor NOR4 (N23341, N23336, N21586, N454, N11056);
and AND2 (N23342, N23326, N7170);
not NOT1 (N23343, N23340);
not NOT1 (N23344, N23319);
not NOT1 (N23345, N23344);
buf BUF1 (N23346, N23329);
or OR2 (N23347, N23339, N22838);
xor XOR2 (N23348, N23345, N12869);
and AND4 (N23349, N23346, N11045, N21225, N22384);
nand NAND4 (N23350, N23325, N19336, N1472, N12504);
buf BUF1 (N23351, N23350);
nand NAND4 (N23352, N23332, N2238, N12280, N21960);
not NOT1 (N23353, N23351);
not NOT1 (N23354, N23348);
or OR2 (N23355, N23342, N19297);
not NOT1 (N23356, N23341);
or OR2 (N23357, N23354, N3018);
buf BUF1 (N23358, N23352);
nand NAND4 (N23359, N23349, N12623, N8756, N12301);
and AND3 (N23360, N23359, N274, N15425);
nor NOR3 (N23361, N23355, N11816, N12401);
not NOT1 (N23362, N23357);
or OR4 (N23363, N23347, N1563, N20595, N14170);
buf BUF1 (N23364, N23328);
or OR3 (N23365, N23333, N16273, N3487);
and AND2 (N23366, N23364, N4082);
or OR2 (N23367, N23358, N13226);
xor XOR2 (N23368, N23365, N21343);
buf BUF1 (N23369, N23361);
nor NOR4 (N23370, N23367, N7031, N2982, N15502);
nor NOR4 (N23371, N23363, N13577, N9936, N6153);
or OR2 (N23372, N23343, N10823);
nor NOR3 (N23373, N23353, N13392, N12036);
xor XOR2 (N23374, N23371, N14316);
buf BUF1 (N23375, N23360);
or OR3 (N23376, N23366, N2280, N23119);
not NOT1 (N23377, N23356);
xor XOR2 (N23378, N23368, N17758);
not NOT1 (N23379, N23376);
or OR3 (N23380, N23374, N3055, N9916);
nor NOR3 (N23381, N23370, N4928, N2807);
buf BUF1 (N23382, N23377);
or OR4 (N23383, N23382, N22927, N17996, N19407);
and AND3 (N23384, N23362, N14962, N20305);
nor NOR3 (N23385, N23380, N10270, N15339);
buf BUF1 (N23386, N23381);
nor NOR4 (N23387, N23378, N14555, N21674, N9495);
xor XOR2 (N23388, N23372, N5241);
and AND4 (N23389, N23386, N4139, N5852, N8514);
nor NOR3 (N23390, N23389, N15349, N8641);
and AND2 (N23391, N23385, N17438);
buf BUF1 (N23392, N23388);
or OR3 (N23393, N23375, N9131, N108);
nand NAND4 (N23394, N23379, N4205, N6189, N18485);
xor XOR2 (N23395, N23373, N19299);
nand NAND4 (N23396, N23384, N5468, N13374, N14030);
nand NAND3 (N23397, N23395, N4817, N22557);
xor XOR2 (N23398, N23369, N1098);
nor NOR2 (N23399, N23396, N766);
not NOT1 (N23400, N23399);
xor XOR2 (N23401, N23393, N431);
nor NOR4 (N23402, N23397, N17711, N13962, N22165);
nor NOR2 (N23403, N23400, N15299);
xor XOR2 (N23404, N23391, N13848);
nand NAND3 (N23405, N23387, N20149, N2771);
not NOT1 (N23406, N23394);
or OR3 (N23407, N23401, N10156, N2251);
or OR2 (N23408, N23402, N21330);
and AND4 (N23409, N23392, N3562, N3264, N10446);
or OR3 (N23410, N23406, N22040, N11750);
xor XOR2 (N23411, N23383, N17197);
not NOT1 (N23412, N23403);
nand NAND2 (N23413, N23390, N15253);
nor NOR3 (N23414, N23412, N21224, N21743);
and AND2 (N23415, N23407, N10580);
xor XOR2 (N23416, N23413, N22079);
and AND2 (N23417, N23404, N1254);
nor NOR2 (N23418, N23416, N16181);
and AND3 (N23419, N23405, N17819, N20325);
xor XOR2 (N23420, N23414, N9978);
and AND2 (N23421, N23408, N16221);
or OR2 (N23422, N23417, N21557);
and AND4 (N23423, N23415, N6129, N13878, N5317);
not NOT1 (N23424, N23422);
buf BUF1 (N23425, N23419);
nand NAND2 (N23426, N23424, N12302);
not NOT1 (N23427, N23411);
not NOT1 (N23428, N23426);
and AND2 (N23429, N23420, N16076);
nor NOR4 (N23430, N23425, N2475, N13632, N19062);
and AND4 (N23431, N23421, N18058, N6836, N8805);
nand NAND3 (N23432, N23418, N3411, N301);
nor NOR3 (N23433, N23430, N884, N3528);
and AND4 (N23434, N23432, N11769, N7829, N10886);
and AND4 (N23435, N23409, N20095, N2015, N4641);
nand NAND3 (N23436, N23427, N19650, N5800);
not NOT1 (N23437, N23423);
nor NOR3 (N23438, N23435, N14308, N10619);
and AND3 (N23439, N23431, N17456, N7330);
not NOT1 (N23440, N23398);
nor NOR4 (N23441, N23434, N20039, N338, N2316);
or OR3 (N23442, N23428, N17261, N2882);
buf BUF1 (N23443, N23433);
or OR4 (N23444, N23437, N10367, N19606, N11596);
nand NAND2 (N23445, N23442, N18099);
not NOT1 (N23446, N23429);
xor XOR2 (N23447, N23438, N12006);
or OR4 (N23448, N23439, N1981, N1587, N19863);
nor NOR2 (N23449, N23446, N23404);
not NOT1 (N23450, N23449);
or OR2 (N23451, N23450, N5136);
nor NOR4 (N23452, N23441, N8320, N370, N15908);
not NOT1 (N23453, N23445);
not NOT1 (N23454, N23448);
xor XOR2 (N23455, N23451, N17483);
or OR3 (N23456, N23410, N1557, N12513);
not NOT1 (N23457, N23453);
not NOT1 (N23458, N23447);
xor XOR2 (N23459, N23458, N23199);
xor XOR2 (N23460, N23444, N5303);
xor XOR2 (N23461, N23457, N4760);
xor XOR2 (N23462, N23443, N15998);
not NOT1 (N23463, N23440);
and AND4 (N23464, N23454, N16369, N15592, N4581);
not NOT1 (N23465, N23463);
nand NAND4 (N23466, N23460, N4378, N14017, N6720);
or OR3 (N23467, N23456, N12303, N3878);
buf BUF1 (N23468, N23465);
buf BUF1 (N23469, N23452);
nor NOR3 (N23470, N23469, N5858, N7209);
xor XOR2 (N23471, N23461, N22975);
and AND3 (N23472, N23459, N29, N2716);
xor XOR2 (N23473, N23472, N13877);
or OR4 (N23474, N23455, N16890, N5268, N22904);
not NOT1 (N23475, N23470);
and AND3 (N23476, N23468, N8968, N5378);
or OR4 (N23477, N23471, N14382, N8358, N12891);
nor NOR2 (N23478, N23476, N5038);
xor XOR2 (N23479, N23478, N5923);
buf BUF1 (N23480, N23479);
xor XOR2 (N23481, N23436, N22414);
or OR3 (N23482, N23481, N11952, N6921);
nand NAND2 (N23483, N23474, N17677);
xor XOR2 (N23484, N23466, N11071);
and AND2 (N23485, N23482, N6148);
nand NAND4 (N23486, N23483, N9967, N1668, N14359);
buf BUF1 (N23487, N23484);
nand NAND4 (N23488, N23487, N10186, N7156, N17230);
buf BUF1 (N23489, N23467);
nand NAND3 (N23490, N23489, N17667, N15360);
nor NOR3 (N23491, N23488, N15598, N7344);
or OR3 (N23492, N23480, N22649, N15077);
nor NOR3 (N23493, N23485, N4618, N9931);
and AND4 (N23494, N23475, N11920, N4502, N388);
nor NOR2 (N23495, N23462, N10765);
nand NAND4 (N23496, N23464, N18263, N8857, N18117);
and AND4 (N23497, N23491, N6655, N10301, N10351);
xor XOR2 (N23498, N23473, N8784);
nor NOR2 (N23499, N23486, N3903);
nor NOR4 (N23500, N23477, N17994, N7716, N14634);
buf BUF1 (N23501, N23498);
not NOT1 (N23502, N23494);
nand NAND2 (N23503, N23501, N16588);
or OR2 (N23504, N23492, N8961);
nor NOR4 (N23505, N23504, N19412, N10640, N23235);
or OR4 (N23506, N23502, N20568, N10068, N15679);
or OR2 (N23507, N23505, N17467);
and AND4 (N23508, N23500, N22404, N16304, N15962);
nand NAND3 (N23509, N23507, N6504, N19282);
nand NAND4 (N23510, N23508, N2980, N7296, N11634);
and AND2 (N23511, N23499, N21380);
nor NOR2 (N23512, N23511, N21148);
buf BUF1 (N23513, N23509);
nor NOR2 (N23514, N23506, N6932);
and AND3 (N23515, N23514, N21805, N18126);
not NOT1 (N23516, N23493);
and AND4 (N23517, N23513, N13745, N13051, N1181);
and AND2 (N23518, N23495, N5039);
buf BUF1 (N23519, N23515);
buf BUF1 (N23520, N23517);
and AND2 (N23521, N23520, N15634);
or OR3 (N23522, N23521, N20739, N4840);
not NOT1 (N23523, N23512);
xor XOR2 (N23524, N23516, N11563);
not NOT1 (N23525, N23496);
buf BUF1 (N23526, N23503);
buf BUF1 (N23527, N23526);
xor XOR2 (N23528, N23527, N19765);
not NOT1 (N23529, N23518);
buf BUF1 (N23530, N23528);
not NOT1 (N23531, N23497);
not NOT1 (N23532, N23522);
nand NAND2 (N23533, N23530, N9331);
and AND3 (N23534, N23531, N10709, N22280);
and AND4 (N23535, N23525, N2866, N6813, N17492);
xor XOR2 (N23536, N23532, N23090);
nor NOR3 (N23537, N23536, N17201, N7080);
and AND3 (N23538, N23535, N11210, N11188);
and AND4 (N23539, N23537, N18167, N11598, N13669);
nand NAND3 (N23540, N23519, N16322, N14290);
or OR2 (N23541, N23524, N4779);
xor XOR2 (N23542, N23523, N18991);
xor XOR2 (N23543, N23540, N3551);
not NOT1 (N23544, N23541);
xor XOR2 (N23545, N23543, N8432);
and AND3 (N23546, N23534, N11210, N22728);
xor XOR2 (N23547, N23546, N6932);
nand NAND3 (N23548, N23533, N7556, N15202);
not NOT1 (N23549, N23548);
buf BUF1 (N23550, N23544);
not NOT1 (N23551, N23529);
nor NOR2 (N23552, N23550, N21057);
or OR4 (N23553, N23539, N5076, N14681, N5830);
or OR2 (N23554, N23538, N14093);
or OR3 (N23555, N23552, N12179, N5029);
nor NOR3 (N23556, N23545, N9039, N4097);
buf BUF1 (N23557, N23549);
or OR2 (N23558, N23553, N20319);
nor NOR2 (N23559, N23551, N14523);
buf BUF1 (N23560, N23557);
xor XOR2 (N23561, N23556, N7907);
or OR2 (N23562, N23510, N6355);
nand NAND4 (N23563, N23555, N1361, N10119, N22508);
and AND3 (N23564, N23563, N17804, N241);
nor NOR2 (N23565, N23561, N13921);
and AND4 (N23566, N23554, N6738, N1545, N22089);
or OR4 (N23567, N23558, N7607, N5115, N15960);
xor XOR2 (N23568, N23564, N3086);
or OR2 (N23569, N23567, N11228);
or OR4 (N23570, N23547, N7082, N2747, N23143);
buf BUF1 (N23571, N23559);
and AND3 (N23572, N23571, N23128, N14260);
not NOT1 (N23573, N23568);
buf BUF1 (N23574, N23566);
nor NOR4 (N23575, N23565, N10767, N2063, N11158);
not NOT1 (N23576, N23573);
xor XOR2 (N23577, N23574, N10576);
and AND3 (N23578, N23577, N9451, N17832);
nand NAND3 (N23579, N23575, N21265, N21839);
and AND2 (N23580, N23579, N5233);
and AND4 (N23581, N23580, N5144, N1845, N12994);
nor NOR2 (N23582, N23581, N3602);
nand NAND2 (N23583, N23569, N4736);
or OR3 (N23584, N23583, N22080, N10761);
nand NAND2 (N23585, N23490, N21369);
nor NOR3 (N23586, N23584, N19427, N7021);
not NOT1 (N23587, N23576);
and AND4 (N23588, N23582, N16832, N9585, N13990);
and AND4 (N23589, N23585, N23541, N14421, N8074);
and AND4 (N23590, N23562, N6354, N4866, N17927);
not NOT1 (N23591, N23589);
not NOT1 (N23592, N23587);
buf BUF1 (N23593, N23560);
buf BUF1 (N23594, N23578);
nor NOR2 (N23595, N23594, N17514);
xor XOR2 (N23596, N23592, N16764);
and AND4 (N23597, N23570, N3822, N9321, N18859);
not NOT1 (N23598, N23597);
nor NOR2 (N23599, N23591, N11294);
not NOT1 (N23600, N23542);
not NOT1 (N23601, N23586);
nor NOR3 (N23602, N23600, N4383, N8175);
nand NAND2 (N23603, N23602, N15992);
not NOT1 (N23604, N23598);
or OR3 (N23605, N23588, N4989, N13594);
nand NAND3 (N23606, N23605, N7977, N2905);
xor XOR2 (N23607, N23604, N9359);
not NOT1 (N23608, N23593);
nand NAND4 (N23609, N23607, N19900, N23174, N1320);
xor XOR2 (N23610, N23572, N10033);
buf BUF1 (N23611, N23590);
xor XOR2 (N23612, N23601, N13442);
nand NAND4 (N23613, N23608, N10059, N5654, N8318);
xor XOR2 (N23614, N23599, N11006);
and AND4 (N23615, N23596, N13042, N22445, N7708);
buf BUF1 (N23616, N23613);
nand NAND4 (N23617, N23595, N16184, N18294, N16916);
not NOT1 (N23618, N23603);
nand NAND4 (N23619, N23614, N20358, N4559, N7993);
or OR2 (N23620, N23616, N2139);
xor XOR2 (N23621, N23612, N18145);
xor XOR2 (N23622, N23617, N16578);
nor NOR3 (N23623, N23621, N12913, N22492);
xor XOR2 (N23624, N23609, N1668);
xor XOR2 (N23625, N23619, N16196);
or OR3 (N23626, N23623, N14533, N6493);
buf BUF1 (N23627, N23620);
not NOT1 (N23628, N23615);
nor NOR2 (N23629, N23624, N10123);
or OR3 (N23630, N23628, N21320, N6661);
nor NOR3 (N23631, N23629, N8329, N11885);
not NOT1 (N23632, N23622);
or OR3 (N23633, N23630, N7487, N116);
buf BUF1 (N23634, N23625);
buf BUF1 (N23635, N23631);
nand NAND4 (N23636, N23618, N17412, N20971, N18354);
xor XOR2 (N23637, N23632, N21782);
or OR4 (N23638, N23635, N7586, N9193, N103);
and AND4 (N23639, N23610, N18441, N22779, N11170);
and AND4 (N23640, N23606, N17180, N4785, N6811);
nand NAND3 (N23641, N23626, N3094, N12108);
nor NOR4 (N23642, N23636, N4351, N17160, N3954);
xor XOR2 (N23643, N23611, N17483);
xor XOR2 (N23644, N23637, N19373);
nand NAND2 (N23645, N23634, N17395);
nor NOR4 (N23646, N23627, N21640, N7446, N14950);
xor XOR2 (N23647, N23645, N11203);
buf BUF1 (N23648, N23639);
xor XOR2 (N23649, N23643, N9287);
nor NOR3 (N23650, N23638, N12035, N16098);
xor XOR2 (N23651, N23650, N11264);
and AND2 (N23652, N23641, N21958);
or OR4 (N23653, N23648, N19829, N13520, N7154);
xor XOR2 (N23654, N23646, N17574);
and AND4 (N23655, N23644, N11453, N16399, N17330);
nand NAND4 (N23656, N23649, N21776, N22666, N16191);
buf BUF1 (N23657, N23633);
or OR2 (N23658, N23657, N15235);
and AND4 (N23659, N23658, N16250, N4497, N16372);
nand NAND4 (N23660, N23654, N13953, N13187, N9512);
or OR3 (N23661, N23659, N7170, N19350);
buf BUF1 (N23662, N23655);
not NOT1 (N23663, N23640);
nand NAND2 (N23664, N23647, N13055);
nand NAND4 (N23665, N23651, N7927, N12407, N3616);
nor NOR4 (N23666, N23656, N19165, N19185, N23185);
and AND2 (N23667, N23665, N20434);
and AND4 (N23668, N23661, N13483, N4451, N14591);
nor NOR3 (N23669, N23652, N6532, N22359);
or OR3 (N23670, N23660, N19769, N3681);
and AND3 (N23671, N23669, N14657, N9983);
buf BUF1 (N23672, N23671);
nand NAND3 (N23673, N23666, N10615, N18081);
not NOT1 (N23674, N23653);
nor NOR3 (N23675, N23672, N5454, N11644);
and AND4 (N23676, N23673, N14598, N1644, N16893);
or OR2 (N23677, N23675, N18196);
nand NAND3 (N23678, N23663, N12769, N11717);
and AND2 (N23679, N23676, N5580);
or OR3 (N23680, N23662, N7486, N12575);
nand NAND3 (N23681, N23667, N6445, N14762);
buf BUF1 (N23682, N23674);
nand NAND2 (N23683, N23678, N1982);
nor NOR2 (N23684, N23683, N9653);
nor NOR4 (N23685, N23682, N8037, N3675, N9973);
nand NAND3 (N23686, N23679, N6770, N15482);
and AND4 (N23687, N23684, N11488, N21100, N21118);
buf BUF1 (N23688, N23680);
nor NOR3 (N23689, N23688, N12775, N13457);
not NOT1 (N23690, N23664);
nand NAND2 (N23691, N23690, N7144);
nor NOR3 (N23692, N23691, N8823, N14384);
nor NOR3 (N23693, N23687, N15607, N964);
xor XOR2 (N23694, N23677, N22040);
nand NAND4 (N23695, N23642, N11001, N14828, N5395);
nor NOR2 (N23696, N23692, N10694);
and AND2 (N23697, N23695, N20387);
nand NAND3 (N23698, N23685, N6529, N15380);
or OR3 (N23699, N23668, N4072, N5758);
nor NOR4 (N23700, N23681, N22053, N7367, N13751);
and AND3 (N23701, N23696, N13079, N15387);
nand NAND4 (N23702, N23694, N19918, N22306, N148);
nor NOR3 (N23703, N23698, N5711, N7385);
buf BUF1 (N23704, N23697);
not NOT1 (N23705, N23702);
not NOT1 (N23706, N23689);
nand NAND3 (N23707, N23670, N13358, N1082);
nor NOR3 (N23708, N23707, N22804, N6679);
not NOT1 (N23709, N23699);
not NOT1 (N23710, N23700);
not NOT1 (N23711, N23704);
buf BUF1 (N23712, N23709);
and AND4 (N23713, N23711, N6334, N23181, N10925);
nand NAND3 (N23714, N23686, N6377, N6864);
buf BUF1 (N23715, N23693);
xor XOR2 (N23716, N23703, N11480);
nor NOR3 (N23717, N23708, N383, N8589);
not NOT1 (N23718, N23713);
and AND2 (N23719, N23705, N15537);
nor NOR2 (N23720, N23719, N6590);
nand NAND4 (N23721, N23715, N15977, N20580, N1810);
not NOT1 (N23722, N23720);
or OR4 (N23723, N23717, N1080, N16795, N1920);
nand NAND4 (N23724, N23723, N9025, N10217, N22889);
not NOT1 (N23725, N23714);
nor NOR2 (N23726, N23721, N16514);
nand NAND2 (N23727, N23712, N2335);
nand NAND4 (N23728, N23718, N9746, N11771, N2691);
nor NOR2 (N23729, N23727, N23095);
nand NAND2 (N23730, N23728, N3681);
xor XOR2 (N23731, N23726, N6796);
and AND3 (N23732, N23725, N532, N19324);
nand NAND4 (N23733, N23729, N1566, N11507, N5047);
nand NAND4 (N23734, N23724, N918, N18948, N15978);
nor NOR4 (N23735, N23716, N18295, N8972, N4766);
and AND2 (N23736, N23735, N8337);
or OR2 (N23737, N23736, N6721);
nand NAND3 (N23738, N23737, N4412, N17791);
buf BUF1 (N23739, N23734);
or OR2 (N23740, N23733, N19719);
nor NOR4 (N23741, N23738, N8633, N4466, N1377);
or OR4 (N23742, N23701, N5007, N23028, N2718);
xor XOR2 (N23743, N23710, N19594);
buf BUF1 (N23744, N23732);
not NOT1 (N23745, N23743);
buf BUF1 (N23746, N23741);
or OR2 (N23747, N23745, N19950);
xor XOR2 (N23748, N23742, N18148);
nor NOR4 (N23749, N23739, N1926, N3150, N15406);
and AND2 (N23750, N23722, N9672);
not NOT1 (N23751, N23706);
buf BUF1 (N23752, N23751);
xor XOR2 (N23753, N23752, N12965);
and AND2 (N23754, N23748, N16709);
nor NOR4 (N23755, N23750, N14577, N11408, N20632);
nor NOR4 (N23756, N23744, N14799, N16215, N19932);
nand NAND3 (N23757, N23756, N8897, N19179);
or OR4 (N23758, N23755, N12186, N8494, N23693);
nor NOR3 (N23759, N23731, N6053, N1292);
xor XOR2 (N23760, N23753, N22160);
or OR3 (N23761, N23760, N11924, N1980);
not NOT1 (N23762, N23730);
and AND2 (N23763, N23754, N6138);
and AND4 (N23764, N23740, N16946, N235, N18491);
or OR3 (N23765, N23761, N17718, N1254);
not NOT1 (N23766, N23758);
buf BUF1 (N23767, N23746);
or OR2 (N23768, N23759, N21717);
or OR4 (N23769, N23768, N21918, N9839, N17523);
or OR2 (N23770, N23765, N10691);
buf BUF1 (N23771, N23757);
nand NAND3 (N23772, N23747, N16242, N11899);
buf BUF1 (N23773, N23764);
xor XOR2 (N23774, N23770, N23147);
xor XOR2 (N23775, N23772, N11109);
nand NAND4 (N23776, N23773, N10824, N4979, N21768);
not NOT1 (N23777, N23749);
nand NAND3 (N23778, N23766, N21967, N13315);
nand NAND3 (N23779, N23775, N2746, N8816);
nand NAND3 (N23780, N23769, N17032, N5580);
and AND2 (N23781, N23780, N20374);
buf BUF1 (N23782, N23778);
nand NAND3 (N23783, N23771, N3784, N21202);
or OR2 (N23784, N23779, N2261);
nor NOR2 (N23785, N23776, N3204);
nand NAND3 (N23786, N23777, N18947, N3910);
nand NAND3 (N23787, N23767, N7620, N23102);
or OR3 (N23788, N23763, N14727, N21509);
nor NOR2 (N23789, N23781, N2677);
xor XOR2 (N23790, N23788, N16780);
nor NOR2 (N23791, N23782, N1372);
xor XOR2 (N23792, N23784, N1015);
or OR4 (N23793, N23785, N7992, N2126, N10685);
xor XOR2 (N23794, N23783, N15554);
nand NAND2 (N23795, N23794, N9962);
nor NOR2 (N23796, N23787, N20102);
buf BUF1 (N23797, N23774);
or OR3 (N23798, N23762, N16833, N17957);
nand NAND2 (N23799, N23789, N16395);
xor XOR2 (N23800, N23793, N17342);
nor NOR2 (N23801, N23791, N12509);
and AND4 (N23802, N23798, N22067, N16835, N12493);
nor NOR4 (N23803, N23790, N20781, N23775, N5427);
or OR4 (N23804, N23803, N2303, N4447, N11902);
buf BUF1 (N23805, N23792);
buf BUF1 (N23806, N23796);
buf BUF1 (N23807, N23786);
and AND3 (N23808, N23806, N13553, N18378);
or OR2 (N23809, N23807, N9126);
nand NAND2 (N23810, N23808, N4121);
buf BUF1 (N23811, N23797);
nor NOR4 (N23812, N23800, N2991, N5952, N22203);
buf BUF1 (N23813, N23795);
or OR2 (N23814, N23804, N3905);
xor XOR2 (N23815, N23813, N12267);
not NOT1 (N23816, N23809);
xor XOR2 (N23817, N23802, N6670);
buf BUF1 (N23818, N23814);
nand NAND3 (N23819, N23810, N18270, N18644);
and AND3 (N23820, N23819, N10974, N22592);
xor XOR2 (N23821, N23820, N16613);
xor XOR2 (N23822, N23817, N16579);
not NOT1 (N23823, N23805);
buf BUF1 (N23824, N23801);
and AND4 (N23825, N23816, N17635, N15781, N3354);
xor XOR2 (N23826, N23818, N6865);
nand NAND2 (N23827, N23821, N18989);
buf BUF1 (N23828, N23825);
not NOT1 (N23829, N23824);
and AND2 (N23830, N23815, N7801);
or OR4 (N23831, N23826, N5447, N21214, N12732);
not NOT1 (N23832, N23831);
nand NAND4 (N23833, N23812, N11722, N4692, N12248);
nand NAND4 (N23834, N23799, N3084, N10177, N19296);
not NOT1 (N23835, N23833);
nor NOR3 (N23836, N23835, N9642, N7454);
not NOT1 (N23837, N23823);
xor XOR2 (N23838, N23822, N13995);
nand NAND2 (N23839, N23832, N23091);
or OR2 (N23840, N23829, N11841);
nand NAND3 (N23841, N23839, N5102, N22665);
nor NOR3 (N23842, N23840, N19054, N14487);
buf BUF1 (N23843, N23834);
nor NOR4 (N23844, N23828, N10297, N23100, N22720);
and AND2 (N23845, N23838, N3902);
not NOT1 (N23846, N23842);
or OR3 (N23847, N23836, N12328, N12292);
nor NOR3 (N23848, N23844, N13435, N4917);
nor NOR4 (N23849, N23843, N13726, N14787, N23621);
and AND3 (N23850, N23837, N20888, N19490);
nand NAND2 (N23851, N23847, N13213);
nand NAND4 (N23852, N23850, N19239, N23782, N11622);
buf BUF1 (N23853, N23830);
buf BUF1 (N23854, N23852);
nand NAND2 (N23855, N23849, N15369);
not NOT1 (N23856, N23855);
xor XOR2 (N23857, N23846, N13641);
and AND4 (N23858, N23857, N21651, N22779, N8216);
or OR3 (N23859, N23858, N10834, N8013);
buf BUF1 (N23860, N23848);
nand NAND4 (N23861, N23827, N13489, N11025, N12560);
nor NOR2 (N23862, N23854, N22636);
xor XOR2 (N23863, N23860, N4875);
and AND2 (N23864, N23859, N16762);
buf BUF1 (N23865, N23811);
nand NAND4 (N23866, N23851, N1095, N7612, N18089);
nand NAND4 (N23867, N23864, N9089, N20654, N22630);
nand NAND4 (N23868, N23867, N16879, N7739, N18158);
and AND4 (N23869, N23868, N12688, N1453, N6481);
xor XOR2 (N23870, N23869, N12403);
or OR3 (N23871, N23870, N2845, N14352);
nand NAND4 (N23872, N23862, N19508, N7742, N3313);
not NOT1 (N23873, N23861);
or OR4 (N23874, N23853, N18977, N3963, N15277);
nor NOR3 (N23875, N23863, N10226, N14537);
nand NAND4 (N23876, N23871, N8595, N10279, N7605);
or OR2 (N23877, N23873, N21555);
not NOT1 (N23878, N23877);
nor NOR2 (N23879, N23872, N14421);
not NOT1 (N23880, N23866);
or OR2 (N23881, N23878, N9770);
xor XOR2 (N23882, N23876, N8676);
xor XOR2 (N23883, N23845, N10603);
xor XOR2 (N23884, N23841, N3430);
not NOT1 (N23885, N23882);
not NOT1 (N23886, N23875);
not NOT1 (N23887, N23879);
nor NOR2 (N23888, N23884, N13340);
or OR3 (N23889, N23887, N2947, N7045);
nand NAND3 (N23890, N23886, N12965, N10045);
and AND3 (N23891, N23874, N12470, N5153);
or OR4 (N23892, N23856, N5100, N4045, N23675);
xor XOR2 (N23893, N23891, N7720);
not NOT1 (N23894, N23890);
not NOT1 (N23895, N23883);
nand NAND4 (N23896, N23880, N22259, N281, N8580);
or OR3 (N23897, N23888, N7323, N7609);
or OR4 (N23898, N23881, N3178, N11077, N12514);
xor XOR2 (N23899, N23885, N13608);
and AND4 (N23900, N23898, N17822, N13439, N8245);
nor NOR3 (N23901, N23892, N6026, N9944);
xor XOR2 (N23902, N23865, N20757);
not NOT1 (N23903, N23897);
nand NAND4 (N23904, N23900, N2163, N13699, N19396);
buf BUF1 (N23905, N23896);
or OR3 (N23906, N23895, N15710, N13188);
buf BUF1 (N23907, N23906);
and AND3 (N23908, N23903, N19396, N20615);
xor XOR2 (N23909, N23894, N15648);
xor XOR2 (N23910, N23889, N21846);
buf BUF1 (N23911, N23910);
and AND2 (N23912, N23904, N16197);
not NOT1 (N23913, N23905);
nor NOR3 (N23914, N23913, N5009, N23728);
not NOT1 (N23915, N23912);
and AND4 (N23916, N23915, N991, N21238, N12434);
buf BUF1 (N23917, N23916);
nor NOR3 (N23918, N23908, N10302, N7406);
nor NOR3 (N23919, N23907, N17423, N245);
nand NAND3 (N23920, N23919, N11046, N22902);
nand NAND4 (N23921, N23909, N852, N5032, N21261);
nand NAND4 (N23922, N23914, N18001, N6629, N9463);
buf BUF1 (N23923, N23902);
not NOT1 (N23924, N23911);
buf BUF1 (N23925, N23922);
not NOT1 (N23926, N23920);
not NOT1 (N23927, N23926);
or OR3 (N23928, N23924, N636, N3833);
or OR3 (N23929, N23901, N15950, N18144);
nand NAND4 (N23930, N23923, N15585, N3377, N23018);
xor XOR2 (N23931, N23929, N13931);
or OR2 (N23932, N23921, N11208);
xor XOR2 (N23933, N23918, N8673);
or OR3 (N23934, N23931, N5118, N14199);
not NOT1 (N23935, N23933);
and AND2 (N23936, N23934, N6337);
buf BUF1 (N23937, N23927);
buf BUF1 (N23938, N23935);
and AND2 (N23939, N23928, N5596);
nand NAND2 (N23940, N23937, N1064);
xor XOR2 (N23941, N23925, N20413);
or OR3 (N23942, N23941, N16402, N12396);
xor XOR2 (N23943, N23940, N19328);
nor NOR2 (N23944, N23936, N22964);
nor NOR2 (N23945, N23942, N21023);
xor XOR2 (N23946, N23943, N10107);
nand NAND2 (N23947, N23938, N18775);
nor NOR4 (N23948, N23944, N5900, N8197, N11479);
buf BUF1 (N23949, N23930);
xor XOR2 (N23950, N23945, N11086);
or OR2 (N23951, N23946, N8859);
buf BUF1 (N23952, N23951);
nand NAND2 (N23953, N23948, N21350);
buf BUF1 (N23954, N23939);
or OR4 (N23955, N23952, N6141, N4458, N737);
not NOT1 (N23956, N23955);
nor NOR2 (N23957, N23893, N18950);
or OR3 (N23958, N23947, N19272, N22773);
and AND2 (N23959, N23957, N16371);
not NOT1 (N23960, N23950);
nand NAND2 (N23961, N23960, N4678);
xor XOR2 (N23962, N23953, N22990);
buf BUF1 (N23963, N23917);
not NOT1 (N23964, N23958);
xor XOR2 (N23965, N23954, N5464);
buf BUF1 (N23966, N23949);
nand NAND4 (N23967, N23932, N22620, N8629, N3366);
and AND3 (N23968, N23962, N9896, N5492);
not NOT1 (N23969, N23968);
nand NAND3 (N23970, N23899, N16427, N10372);
nor NOR3 (N23971, N23970, N5110, N13951);
not NOT1 (N23972, N23956);
not NOT1 (N23973, N23964);
not NOT1 (N23974, N23973);
nand NAND3 (N23975, N23961, N11033, N21636);
xor XOR2 (N23976, N23966, N17055);
xor XOR2 (N23977, N23959, N3081);
and AND4 (N23978, N23965, N6580, N17297, N19526);
or OR4 (N23979, N23972, N572, N22689, N14520);
not NOT1 (N23980, N23967);
xor XOR2 (N23981, N23976, N1117);
or OR4 (N23982, N23979, N20687, N10048, N5265);
not NOT1 (N23983, N23982);
or OR2 (N23984, N23978, N7677);
and AND3 (N23985, N23969, N21269, N10983);
xor XOR2 (N23986, N23971, N14356);
xor XOR2 (N23987, N23974, N8767);
nand NAND3 (N23988, N23985, N11456, N8875);
not NOT1 (N23989, N23983);
xor XOR2 (N23990, N23989, N13047);
nand NAND4 (N23991, N23984, N6110, N19465, N5311);
buf BUF1 (N23992, N23986);
or OR4 (N23993, N23990, N8217, N20630, N6797);
xor XOR2 (N23994, N23980, N12802);
nor NOR4 (N23995, N23977, N23837, N22901, N6205);
nor NOR4 (N23996, N23994, N1812, N1877, N22192);
buf BUF1 (N23997, N23963);
nand NAND3 (N23998, N23992, N4505, N16461);
or OR2 (N23999, N23987, N8908);
and AND2 (N24000, N23995, N8078);
and AND2 (N24001, N23998, N13419);
not NOT1 (N24002, N23997);
or OR3 (N24003, N23996, N15626, N15941);
buf BUF1 (N24004, N23975);
nor NOR2 (N24005, N23993, N3724);
nor NOR3 (N24006, N23999, N9931, N13102);
nand NAND4 (N24007, N23988, N1006, N22758, N1446);
and AND3 (N24008, N24002, N13720, N4446);
nand NAND4 (N24009, N24007, N252, N23175, N2075);
or OR3 (N24010, N24001, N2594, N16587);
or OR3 (N24011, N24009, N12992, N4075);
buf BUF1 (N24012, N23991);
and AND4 (N24013, N24003, N6072, N11196, N3095);
not NOT1 (N24014, N24013);
or OR4 (N24015, N24008, N14287, N2806, N12980);
and AND4 (N24016, N24015, N18159, N21444, N21411);
nor NOR3 (N24017, N24004, N23865, N7741);
nor NOR2 (N24018, N24010, N15627);
or OR3 (N24019, N24018, N20193, N11573);
or OR4 (N24020, N24005, N12361, N5282, N7956);
nand NAND4 (N24021, N23981, N15578, N1261, N21674);
and AND2 (N24022, N24014, N1516);
xor XOR2 (N24023, N24020, N16153);
buf BUF1 (N24024, N24006);
nand NAND3 (N24025, N24017, N1660, N20125);
buf BUF1 (N24026, N24025);
not NOT1 (N24027, N24024);
xor XOR2 (N24028, N24000, N21447);
and AND2 (N24029, N24023, N14110);
or OR3 (N24030, N24016, N15344, N6597);
and AND2 (N24031, N24012, N20752);
not NOT1 (N24032, N24021);
and AND4 (N24033, N24022, N6231, N9760, N8286);
xor XOR2 (N24034, N24033, N1871);
buf BUF1 (N24035, N24011);
and AND2 (N24036, N24035, N14085);
xor XOR2 (N24037, N24036, N2913);
not NOT1 (N24038, N24026);
nor NOR2 (N24039, N24034, N19282);
buf BUF1 (N24040, N24032);
buf BUF1 (N24041, N24037);
or OR2 (N24042, N24029, N3122);
xor XOR2 (N24043, N24028, N12515);
nor NOR4 (N24044, N24042, N10754, N2548, N18159);
or OR2 (N24045, N24031, N18810);
nor NOR4 (N24046, N24044, N21560, N834, N45);
nor NOR2 (N24047, N24027, N4734);
buf BUF1 (N24048, N24045);
not NOT1 (N24049, N24030);
or OR2 (N24050, N24039, N13585);
buf BUF1 (N24051, N24043);
or OR2 (N24052, N24041, N9865);
xor XOR2 (N24053, N24019, N16124);
buf BUF1 (N24054, N24050);
not NOT1 (N24055, N24051);
buf BUF1 (N24056, N24052);
nand NAND2 (N24057, N24046, N10828);
not NOT1 (N24058, N24047);
xor XOR2 (N24059, N24038, N5548);
or OR3 (N24060, N24054, N15683, N9506);
buf BUF1 (N24061, N24053);
xor XOR2 (N24062, N24048, N24027);
nand NAND2 (N24063, N24055, N6421);
or OR4 (N24064, N24056, N15492, N5334, N10013);
nor NOR4 (N24065, N24063, N7773, N22951, N8997);
not NOT1 (N24066, N24064);
xor XOR2 (N24067, N24060, N783);
nand NAND4 (N24068, N24059, N9386, N17351, N5984);
or OR4 (N24069, N24062, N3141, N19041, N13449);
buf BUF1 (N24070, N24065);
nand NAND2 (N24071, N24058, N8653);
nor NOR4 (N24072, N24071, N18430, N1893, N5247);
or OR2 (N24073, N24069, N6835);
or OR4 (N24074, N24073, N5093, N3230, N17490);
not NOT1 (N24075, N24049);
buf BUF1 (N24076, N24072);
buf BUF1 (N24077, N24040);
nand NAND3 (N24078, N24067, N14958, N7536);
buf BUF1 (N24079, N24066);
nand NAND4 (N24080, N24079, N4883, N22448, N22660);
nand NAND2 (N24081, N24077, N5510);
xor XOR2 (N24082, N24070, N8522);
not NOT1 (N24083, N24057);
or OR4 (N24084, N24081, N11687, N1734, N9772);
nor NOR4 (N24085, N24074, N5880, N17030, N18007);
nand NAND2 (N24086, N24084, N18116);
not NOT1 (N24087, N24086);
xor XOR2 (N24088, N24078, N21805);
not NOT1 (N24089, N24088);
and AND4 (N24090, N24061, N23633, N22032, N3759);
and AND4 (N24091, N24085, N12897, N23729, N13416);
or OR4 (N24092, N24076, N10014, N14003, N10805);
or OR2 (N24093, N24089, N8742);
and AND4 (N24094, N24091, N142, N10079, N1934);
nor NOR3 (N24095, N24080, N7432, N12861);
or OR4 (N24096, N24095, N20836, N10933, N21321);
and AND3 (N24097, N24090, N357, N20744);
not NOT1 (N24098, N24094);
or OR2 (N24099, N24075, N22354);
and AND4 (N24100, N24083, N4054, N19205, N6816);
and AND3 (N24101, N24087, N21002, N14950);
xor XOR2 (N24102, N24082, N6211);
nand NAND4 (N24103, N24093, N19085, N6025, N3071);
nand NAND4 (N24104, N24100, N15932, N16494, N2008);
or OR2 (N24105, N24103, N9328);
xor XOR2 (N24106, N24092, N20742);
buf BUF1 (N24107, N24068);
and AND3 (N24108, N24105, N1690, N1805);
and AND2 (N24109, N24099, N8103);
or OR3 (N24110, N24106, N2587, N20870);
or OR4 (N24111, N24108, N20775, N8247, N11273);
xor XOR2 (N24112, N24097, N8780);
and AND2 (N24113, N24104, N3550);
nand NAND2 (N24114, N24096, N23607);
nand NAND2 (N24115, N24111, N16011);
nor NOR4 (N24116, N24112, N13878, N17258, N10951);
nand NAND2 (N24117, N24114, N14259);
or OR2 (N24118, N24109, N20815);
xor XOR2 (N24119, N24110, N12571);
and AND2 (N24120, N24113, N15626);
buf BUF1 (N24121, N24118);
nor NOR2 (N24122, N24119, N15756);
and AND2 (N24123, N24122, N22410);
and AND2 (N24124, N24117, N17513);
buf BUF1 (N24125, N24102);
nand NAND4 (N24126, N24101, N22145, N15393, N22901);
xor XOR2 (N24127, N24125, N19975);
xor XOR2 (N24128, N24120, N12651);
buf BUF1 (N24129, N24123);
nand NAND2 (N24130, N24107, N17460);
nor NOR2 (N24131, N24121, N17415);
nor NOR4 (N24132, N24115, N3034, N21632, N10892);
and AND3 (N24133, N24131, N15741, N3478);
nor NOR3 (N24134, N24116, N3160, N3259);
and AND4 (N24135, N24132, N10080, N6136, N20966);
buf BUF1 (N24136, N24126);
buf BUF1 (N24137, N24130);
or OR4 (N24138, N24124, N23545, N263, N18659);
xor XOR2 (N24139, N24129, N9253);
or OR3 (N24140, N24128, N17373, N16778);
and AND3 (N24141, N24133, N1634, N7676);
nand NAND3 (N24142, N24137, N13839, N21444);
xor XOR2 (N24143, N24140, N1411);
not NOT1 (N24144, N24134);
buf BUF1 (N24145, N24098);
not NOT1 (N24146, N24127);
not NOT1 (N24147, N24143);
buf BUF1 (N24148, N24139);
buf BUF1 (N24149, N24145);
buf BUF1 (N24150, N24149);
or OR2 (N24151, N24141, N6664);
not NOT1 (N24152, N24147);
or OR3 (N24153, N24150, N8725, N5409);
and AND4 (N24154, N24144, N20559, N18224, N9114);
nor NOR4 (N24155, N24138, N15160, N21676, N2322);
not NOT1 (N24156, N24142);
xor XOR2 (N24157, N24136, N15894);
not NOT1 (N24158, N24156);
not NOT1 (N24159, N24154);
nand NAND2 (N24160, N24148, N7448);
not NOT1 (N24161, N24135);
not NOT1 (N24162, N24158);
nand NAND4 (N24163, N24161, N16772, N5201, N2972);
or OR2 (N24164, N24155, N12046);
and AND3 (N24165, N24151, N5543, N13586);
or OR3 (N24166, N24153, N6736, N3080);
and AND4 (N24167, N24152, N9635, N14894, N18250);
not NOT1 (N24168, N24160);
or OR2 (N24169, N24164, N8699);
buf BUF1 (N24170, N24157);
buf BUF1 (N24171, N24159);
and AND4 (N24172, N24165, N2539, N7983, N8995);
or OR3 (N24173, N24163, N16145, N6985);
nand NAND2 (N24174, N24171, N21726);
nor NOR4 (N24175, N24146, N6714, N1287, N21691);
buf BUF1 (N24176, N24166);
xor XOR2 (N24177, N24167, N6308);
xor XOR2 (N24178, N24175, N22561);
xor XOR2 (N24179, N24162, N14966);
xor XOR2 (N24180, N24172, N21808);
or OR3 (N24181, N24168, N10709, N14220);
nor NOR2 (N24182, N24170, N15730);
nor NOR4 (N24183, N24173, N16776, N6163, N7060);
or OR4 (N24184, N24179, N10610, N9700, N7672);
nor NOR2 (N24185, N24180, N20134);
nand NAND2 (N24186, N24177, N10934);
buf BUF1 (N24187, N24182);
xor XOR2 (N24188, N24176, N7420);
nand NAND3 (N24189, N24185, N2374, N20141);
and AND3 (N24190, N24169, N7680, N7899);
nand NAND3 (N24191, N24174, N1252, N14589);
nor NOR4 (N24192, N24183, N11117, N8821, N4718);
or OR2 (N24193, N24184, N2906);
xor XOR2 (N24194, N24191, N7260);
buf BUF1 (N24195, N24187);
and AND3 (N24196, N24195, N20000, N199);
or OR4 (N24197, N24181, N18424, N21010, N21408);
xor XOR2 (N24198, N24188, N1420);
nor NOR2 (N24199, N24198, N7760);
xor XOR2 (N24200, N24194, N3138);
nor NOR4 (N24201, N24193, N21006, N3927, N13995);
nand NAND3 (N24202, N24186, N10440, N4220);
nand NAND4 (N24203, N24202, N16205, N10713, N14674);
not NOT1 (N24204, N24178);
buf BUF1 (N24205, N24204);
or OR4 (N24206, N24199, N18852, N12189, N756);
nand NAND3 (N24207, N24203, N1938, N20298);
or OR4 (N24208, N24200, N18059, N11225, N3678);
nor NOR2 (N24209, N24197, N17515);
buf BUF1 (N24210, N24201);
nand NAND3 (N24211, N24189, N19298, N13683);
or OR3 (N24212, N24206, N3866, N14745);
nor NOR4 (N24213, N24210, N21478, N10597, N15218);
and AND2 (N24214, N24208, N691);
or OR3 (N24215, N24211, N14845, N1939);
buf BUF1 (N24216, N24214);
buf BUF1 (N24217, N24215);
and AND3 (N24218, N24192, N18125, N22665);
buf BUF1 (N24219, N24212);
nor NOR2 (N24220, N24205, N12747);
and AND4 (N24221, N24219, N8012, N23734, N21073);
and AND3 (N24222, N24190, N17760, N13076);
xor XOR2 (N24223, N24207, N464);
or OR3 (N24224, N24218, N4026, N10432);
and AND4 (N24225, N24216, N18002, N376, N20398);
or OR4 (N24226, N24209, N9954, N8013, N24190);
not NOT1 (N24227, N24225);
not NOT1 (N24228, N24220);
nand NAND3 (N24229, N24228, N18447, N9768);
buf BUF1 (N24230, N24221);
or OR4 (N24231, N24222, N1862, N19527, N10502);
and AND3 (N24232, N24213, N19107, N12136);
not NOT1 (N24233, N24224);
not NOT1 (N24234, N24227);
and AND4 (N24235, N24196, N6519, N15462, N19709);
and AND4 (N24236, N24217, N18032, N2546, N1418);
or OR2 (N24237, N24226, N10970);
xor XOR2 (N24238, N24231, N20898);
nand NAND2 (N24239, N24233, N22838);
not NOT1 (N24240, N24236);
xor XOR2 (N24241, N24235, N16778);
nor NOR3 (N24242, N24239, N1320, N5898);
and AND2 (N24243, N24223, N11317);
or OR3 (N24244, N24234, N14552, N6373);
nand NAND2 (N24245, N24242, N18989);
or OR3 (N24246, N24229, N6709, N1679);
buf BUF1 (N24247, N24245);
or OR4 (N24248, N24243, N4247, N905, N5633);
xor XOR2 (N24249, N24230, N11345);
not NOT1 (N24250, N24232);
nor NOR3 (N24251, N24240, N11933, N10645);
and AND4 (N24252, N24251, N5721, N4827, N4915);
nand NAND4 (N24253, N24237, N20829, N6027, N17975);
not NOT1 (N24254, N24246);
nor NOR3 (N24255, N24249, N3205, N13846);
nor NOR4 (N24256, N24253, N20377, N3872, N2978);
and AND3 (N24257, N24241, N21043, N6087);
and AND4 (N24258, N24254, N3622, N23632, N20442);
buf BUF1 (N24259, N24255);
xor XOR2 (N24260, N24259, N4098);
nor NOR4 (N24261, N24257, N21931, N18706, N2923);
not NOT1 (N24262, N24238);
nand NAND4 (N24263, N24262, N7128, N13183, N12901);
nor NOR4 (N24264, N24263, N9590, N897, N2793);
nand NAND3 (N24265, N24248, N12188, N21218);
or OR2 (N24266, N24256, N20691);
nand NAND3 (N24267, N24260, N14519, N16159);
nor NOR3 (N24268, N24261, N17207, N18578);
not NOT1 (N24269, N24266);
buf BUF1 (N24270, N24258);
not NOT1 (N24271, N24247);
buf BUF1 (N24272, N24264);
or OR3 (N24273, N24265, N18260, N19);
nand NAND4 (N24274, N24268, N2718, N5425, N8308);
and AND4 (N24275, N24273, N20709, N20191, N797);
not NOT1 (N24276, N24272);
not NOT1 (N24277, N24252);
buf BUF1 (N24278, N24271);
nor NOR2 (N24279, N24275, N20642);
buf BUF1 (N24280, N24276);
buf BUF1 (N24281, N24278);
and AND2 (N24282, N24269, N6344);
xor XOR2 (N24283, N24250, N12979);
buf BUF1 (N24284, N24274);
nor NOR2 (N24285, N24244, N6896);
nand NAND3 (N24286, N24280, N23583, N22654);
buf BUF1 (N24287, N24283);
xor XOR2 (N24288, N24279, N13583);
nor NOR2 (N24289, N24288, N22283);
nor NOR3 (N24290, N24281, N22348, N10822);
or OR3 (N24291, N24289, N15670, N21772);
nand NAND4 (N24292, N24287, N17906, N15992, N5979);
or OR4 (N24293, N24267, N7310, N8065, N4455);
nand NAND3 (N24294, N24290, N387, N18102);
and AND4 (N24295, N24294, N7228, N13123, N18919);
or OR4 (N24296, N24277, N23167, N7353, N7483);
not NOT1 (N24297, N24270);
not NOT1 (N24298, N24293);
buf BUF1 (N24299, N24296);
xor XOR2 (N24300, N24295, N5067);
and AND3 (N24301, N24282, N9803, N10091);
xor XOR2 (N24302, N24300, N10960);
xor XOR2 (N24303, N24301, N11106);
or OR3 (N24304, N24286, N7425, N24253);
and AND4 (N24305, N24304, N15586, N24055, N12822);
not NOT1 (N24306, N24305);
xor XOR2 (N24307, N24302, N15477);
not NOT1 (N24308, N24298);
nor NOR3 (N24309, N24299, N6022, N22180);
nand NAND3 (N24310, N24306, N11251, N3417);
nand NAND3 (N24311, N24307, N22852, N24209);
nand NAND2 (N24312, N24303, N780);
nand NAND2 (N24313, N24284, N18685);
nor NOR2 (N24314, N24309, N9120);
and AND4 (N24315, N24314, N23163, N1173, N16604);
or OR2 (N24316, N24310, N11121);
nand NAND2 (N24317, N24308, N13259);
or OR2 (N24318, N24311, N16364);
nor NOR3 (N24319, N24317, N1396, N19345);
xor XOR2 (N24320, N24291, N3823);
nor NOR4 (N24321, N24285, N23762, N2974, N14031);
buf BUF1 (N24322, N24316);
nor NOR3 (N24323, N24312, N21013, N11159);
buf BUF1 (N24324, N24318);
nand NAND2 (N24325, N24292, N516);
nand NAND3 (N24326, N24322, N4912, N10988);
or OR3 (N24327, N24315, N13073, N10967);
nand NAND4 (N24328, N24325, N19195, N21156, N4085);
buf BUF1 (N24329, N24323);
nor NOR2 (N24330, N24313, N17941);
nand NAND2 (N24331, N24319, N13614);
nor NOR4 (N24332, N24321, N8589, N19069, N18702);
buf BUF1 (N24333, N24297);
nor NOR2 (N24334, N24333, N8214);
nor NOR4 (N24335, N24328, N19887, N1966, N6522);
and AND2 (N24336, N24332, N576);
nor NOR4 (N24337, N24327, N10193, N18935, N20936);
not NOT1 (N24338, N24335);
nor NOR2 (N24339, N24337, N22598);
nand NAND3 (N24340, N24320, N5879, N536);
nor NOR3 (N24341, N24336, N12134, N16221);
not NOT1 (N24342, N24339);
nor NOR4 (N24343, N24330, N5377, N11670, N12770);
or OR3 (N24344, N24343, N2622, N11149);
or OR3 (N24345, N24342, N3717, N14029);
xor XOR2 (N24346, N24341, N1885);
and AND4 (N24347, N24338, N3382, N4046, N10409);
or OR3 (N24348, N24346, N15552, N13381);
or OR2 (N24349, N24345, N5607);
or OR3 (N24350, N24334, N24132, N3677);
nand NAND2 (N24351, N24347, N10473);
nand NAND2 (N24352, N24329, N5601);
xor XOR2 (N24353, N24326, N23077);
buf BUF1 (N24354, N24350);
or OR2 (N24355, N24351, N9522);
buf BUF1 (N24356, N24348);
buf BUF1 (N24357, N24356);
buf BUF1 (N24358, N24324);
buf BUF1 (N24359, N24344);
nand NAND2 (N24360, N24359, N22992);
nand NAND2 (N24361, N24340, N13977);
nand NAND4 (N24362, N24354, N8578, N21667, N17171);
not NOT1 (N24363, N24358);
not NOT1 (N24364, N24349);
nor NOR2 (N24365, N24363, N3553);
nor NOR2 (N24366, N24353, N21779);
and AND2 (N24367, N24352, N6733);
nor NOR2 (N24368, N24364, N16947);
nor NOR3 (N24369, N24357, N1295, N19251);
and AND4 (N24370, N24361, N10781, N10135, N8646);
nand NAND2 (N24371, N24355, N16220);
buf BUF1 (N24372, N24360);
xor XOR2 (N24373, N24368, N5190);
and AND4 (N24374, N24365, N15199, N12111, N18761);
nand NAND2 (N24375, N24331, N3744);
nor NOR2 (N24376, N24372, N2582);
not NOT1 (N24377, N24375);
nor NOR3 (N24378, N24366, N7735, N24357);
not NOT1 (N24379, N24369);
not NOT1 (N24380, N24373);
nand NAND3 (N24381, N24370, N484, N13723);
not NOT1 (N24382, N24378);
nand NAND2 (N24383, N24367, N12617);
nand NAND4 (N24384, N24382, N10270, N2883, N6968);
buf BUF1 (N24385, N24383);
and AND3 (N24386, N24380, N8207, N21616);
xor XOR2 (N24387, N24371, N9251);
nand NAND2 (N24388, N24387, N1071);
nand NAND2 (N24389, N24384, N19876);
buf BUF1 (N24390, N24377);
or OR2 (N24391, N24390, N8431);
not NOT1 (N24392, N24385);
xor XOR2 (N24393, N24388, N6604);
and AND2 (N24394, N24379, N185);
xor XOR2 (N24395, N24374, N18546);
buf BUF1 (N24396, N24381);
nand NAND3 (N24397, N24395, N4242, N17133);
xor XOR2 (N24398, N24396, N4786);
or OR3 (N24399, N24386, N10664, N7976);
not NOT1 (N24400, N24394);
nand NAND3 (N24401, N24391, N10486, N1537);
not NOT1 (N24402, N24398);
nor NOR2 (N24403, N24401, N14377);
nand NAND2 (N24404, N24399, N22296);
xor XOR2 (N24405, N24404, N23902);
nor NOR4 (N24406, N24403, N992, N16199, N3693);
nor NOR3 (N24407, N24389, N10961, N6223);
buf BUF1 (N24408, N24397);
xor XOR2 (N24409, N24406, N14061);
not NOT1 (N24410, N24393);
xor XOR2 (N24411, N24392, N14582);
nor NOR3 (N24412, N24410, N15188, N9419);
or OR3 (N24413, N24405, N590, N21954);
or OR4 (N24414, N24413, N13933, N5289, N21247);
buf BUF1 (N24415, N24402);
and AND3 (N24416, N24409, N9717, N6967);
nor NOR3 (N24417, N24415, N773, N18738);
nand NAND4 (N24418, N24417, N18202, N20820, N23119);
nand NAND4 (N24419, N24416, N10232, N12144, N3286);
xor XOR2 (N24420, N24414, N22067);
or OR2 (N24421, N24376, N7516);
and AND3 (N24422, N24411, N21590, N6601);
and AND2 (N24423, N24362, N23824);
buf BUF1 (N24424, N24408);
not NOT1 (N24425, N24423);
not NOT1 (N24426, N24400);
or OR3 (N24427, N24420, N4720, N17956);
or OR4 (N24428, N24407, N23072, N21338, N7475);
nand NAND4 (N24429, N24422, N22231, N19936, N24093);
and AND4 (N24430, N24424, N18399, N15440, N3521);
and AND4 (N24431, N24427, N9783, N17577, N346);
buf BUF1 (N24432, N24431);
nor NOR4 (N24433, N24426, N16463, N11458, N18495);
and AND3 (N24434, N24429, N20069, N6819);
and AND2 (N24435, N24432, N16630);
nor NOR3 (N24436, N24419, N6699, N17964);
xor XOR2 (N24437, N24421, N19783);
xor XOR2 (N24438, N24418, N360);
nand NAND4 (N24439, N24437, N15969, N18790, N3870);
xor XOR2 (N24440, N24438, N17813);
or OR4 (N24441, N24428, N3438, N9808, N21090);
buf BUF1 (N24442, N24425);
and AND2 (N24443, N24435, N2243);
or OR2 (N24444, N24440, N10334);
nand NAND2 (N24445, N24436, N493);
and AND2 (N24446, N24442, N16879);
not NOT1 (N24447, N24439);
nand NAND2 (N24448, N24447, N13273);
nand NAND4 (N24449, N24446, N6971, N15885, N16322);
nor NOR2 (N24450, N24433, N6300);
not NOT1 (N24451, N24450);
or OR3 (N24452, N24448, N18257, N14272);
nor NOR4 (N24453, N24452, N17040, N15888, N22165);
nor NOR3 (N24454, N24441, N11542, N10270);
buf BUF1 (N24455, N24443);
nand NAND4 (N24456, N24451, N19259, N14209, N23054);
not NOT1 (N24457, N24430);
nor NOR2 (N24458, N24445, N7432);
buf BUF1 (N24459, N24458);
nand NAND2 (N24460, N24412, N15777);
not NOT1 (N24461, N24457);
xor XOR2 (N24462, N24454, N8305);
buf BUF1 (N24463, N24449);
xor XOR2 (N24464, N24455, N24274);
xor XOR2 (N24465, N24460, N404);
not NOT1 (N24466, N24463);
or OR4 (N24467, N24456, N10556, N6460, N20363);
not NOT1 (N24468, N24465);
xor XOR2 (N24469, N24459, N10566);
and AND2 (N24470, N24467, N8568);
and AND2 (N24471, N24466, N18649);
not NOT1 (N24472, N24444);
buf BUF1 (N24473, N24434);
or OR4 (N24474, N24469, N12400, N21134, N4004);
and AND2 (N24475, N24464, N3623);
and AND3 (N24476, N24474, N17256, N24058);
xor XOR2 (N24477, N24475, N9488);
or OR3 (N24478, N24473, N22660, N14656);
not NOT1 (N24479, N24462);
nor NOR4 (N24480, N24476, N11456, N347, N2450);
buf BUF1 (N24481, N24472);
buf BUF1 (N24482, N24481);
nand NAND4 (N24483, N24470, N23568, N19867, N18902);
not NOT1 (N24484, N24479);
xor XOR2 (N24485, N24480, N20633);
not NOT1 (N24486, N24471);
xor XOR2 (N24487, N24484, N5043);
nand NAND4 (N24488, N24477, N20979, N12687, N4275);
xor XOR2 (N24489, N24487, N6955);
and AND3 (N24490, N24488, N23426, N16121);
xor XOR2 (N24491, N24461, N3605);
xor XOR2 (N24492, N24483, N9879);
or OR3 (N24493, N24478, N4722, N23651);
nor NOR3 (N24494, N24489, N22584, N9637);
or OR4 (N24495, N24493, N16669, N6280, N2397);
nand NAND3 (N24496, N24494, N524, N21848);
nor NOR3 (N24497, N24468, N11910, N5892);
nor NOR3 (N24498, N24496, N11966, N6929);
xor XOR2 (N24499, N24495, N4465);
or OR2 (N24500, N24492, N17978);
nand NAND4 (N24501, N24453, N24067, N3317, N24344);
xor XOR2 (N24502, N24482, N190);
xor XOR2 (N24503, N24485, N12457);
buf BUF1 (N24504, N24501);
buf BUF1 (N24505, N24497);
nand NAND4 (N24506, N24498, N19468, N12268, N4582);
or OR4 (N24507, N24503, N4109, N1822, N4743);
not NOT1 (N24508, N24491);
nand NAND3 (N24509, N24499, N15077, N2345);
xor XOR2 (N24510, N24508, N17323);
and AND4 (N24511, N24486, N2131, N7026, N15942);
nor NOR4 (N24512, N24500, N22528, N24417, N13712);
and AND4 (N24513, N24510, N12685, N6160, N11801);
nor NOR2 (N24514, N24511, N9893);
not NOT1 (N24515, N24514);
buf BUF1 (N24516, N24505);
nor NOR2 (N24517, N24515, N15164);
nand NAND4 (N24518, N24504, N10032, N17953, N18741);
or OR2 (N24519, N24506, N17784);
not NOT1 (N24520, N24516);
nor NOR3 (N24521, N24513, N8309, N17465);
or OR2 (N24522, N24507, N15371);
buf BUF1 (N24523, N24509);
nor NOR2 (N24524, N24512, N3220);
and AND4 (N24525, N24522, N10964, N14333, N17323);
not NOT1 (N24526, N24518);
nand NAND4 (N24527, N24525, N17308, N9478, N17244);
nand NAND3 (N24528, N24526, N11348, N22658);
buf BUF1 (N24529, N24527);
and AND4 (N24530, N24519, N17862, N20660, N2399);
and AND2 (N24531, N24521, N23274);
xor XOR2 (N24532, N24523, N529);
not NOT1 (N24533, N24502);
nor NOR3 (N24534, N24490, N20789, N816);
and AND3 (N24535, N24529, N18807, N14835);
and AND4 (N24536, N24532, N248, N23049, N20478);
nor NOR4 (N24537, N24534, N10942, N11086, N7962);
buf BUF1 (N24538, N24537);
or OR3 (N24539, N24524, N2492, N3650);
xor XOR2 (N24540, N24533, N23818);
nand NAND4 (N24541, N24531, N13562, N8159, N23784);
or OR2 (N24542, N24517, N1309);
and AND4 (N24543, N24536, N17789, N24489, N5879);
nor NOR4 (N24544, N24538, N17390, N15469, N23567);
nand NAND4 (N24545, N24543, N4060, N12241, N20958);
nor NOR2 (N24546, N24541, N13287);
buf BUF1 (N24547, N24540);
or OR3 (N24548, N24544, N3556, N11636);
nor NOR3 (N24549, N24520, N15929, N20835);
xor XOR2 (N24550, N24546, N13599);
xor XOR2 (N24551, N24547, N4827);
nor NOR4 (N24552, N24528, N23720, N10470, N15065);
nand NAND3 (N24553, N24550, N18136, N5525);
or OR4 (N24554, N24552, N1350, N9437, N23830);
nand NAND4 (N24555, N24551, N1690, N6608, N16896);
xor XOR2 (N24556, N24539, N1777);
nand NAND3 (N24557, N24548, N16621, N4946);
and AND4 (N24558, N24554, N11299, N19979, N7918);
xor XOR2 (N24559, N24558, N14768);
nand NAND4 (N24560, N24555, N8409, N13418, N77);
not NOT1 (N24561, N24559);
buf BUF1 (N24562, N24553);
buf BUF1 (N24563, N24545);
nor NOR4 (N24564, N24549, N1397, N12558, N12754);
or OR3 (N24565, N24556, N23915, N11188);
xor XOR2 (N24566, N24535, N11349);
xor XOR2 (N24567, N24565, N20568);
and AND4 (N24568, N24562, N1034, N18154, N19900);
buf BUF1 (N24569, N24560);
and AND4 (N24570, N24542, N6550, N20008, N16137);
nand NAND4 (N24571, N24570, N2346, N6375, N17479);
or OR3 (N24572, N24569, N14330, N392);
xor XOR2 (N24573, N24564, N4886);
buf BUF1 (N24574, N24568);
buf BUF1 (N24575, N24566);
xor XOR2 (N24576, N24561, N23634);
xor XOR2 (N24577, N24576, N12966);
or OR2 (N24578, N24563, N21360);
buf BUF1 (N24579, N24575);
nand NAND3 (N24580, N24578, N7690, N22351);
or OR2 (N24581, N24530, N1694);
buf BUF1 (N24582, N24580);
and AND2 (N24583, N24582, N5491);
not NOT1 (N24584, N24574);
or OR2 (N24585, N24557, N21371);
nor NOR3 (N24586, N24579, N13792, N11190);
xor XOR2 (N24587, N24584, N18429);
and AND4 (N24588, N24587, N8167, N15768, N24006);
xor XOR2 (N24589, N24588, N14323);
not NOT1 (N24590, N24573);
and AND3 (N24591, N24586, N17028, N956);
and AND3 (N24592, N24581, N10170, N10834);
not NOT1 (N24593, N24567);
not NOT1 (N24594, N24590);
nand NAND2 (N24595, N24585, N4954);
or OR4 (N24596, N24595, N1305, N5716, N21916);
not NOT1 (N24597, N24594);
nor NOR4 (N24598, N24571, N4054, N3641, N19056);
nor NOR4 (N24599, N24589, N12778, N14520, N8651);
nand NAND3 (N24600, N24591, N6353, N2778);
or OR3 (N24601, N24598, N16435, N6003);
nand NAND4 (N24602, N24600, N9554, N21748, N12121);
xor XOR2 (N24603, N24597, N5299);
and AND3 (N24604, N24596, N3644, N7445);
buf BUF1 (N24605, N24603);
nor NOR3 (N24606, N24572, N11525, N13124);
nand NAND2 (N24607, N24583, N1132);
or OR2 (N24608, N24606, N19543);
not NOT1 (N24609, N24599);
buf BUF1 (N24610, N24577);
or OR2 (N24611, N24602, N20408);
and AND2 (N24612, N24593, N21401);
and AND2 (N24613, N24604, N8797);
nand NAND4 (N24614, N24610, N9964, N15315, N5185);
buf BUF1 (N24615, N24612);
buf BUF1 (N24616, N24613);
or OR2 (N24617, N24592, N7296);
and AND3 (N24618, N24601, N3233, N16270);
xor XOR2 (N24619, N24608, N19160);
nor NOR4 (N24620, N24605, N18832, N3038, N15808);
not NOT1 (N24621, N24607);
nand NAND2 (N24622, N24618, N14597);
or OR2 (N24623, N24614, N13689);
buf BUF1 (N24624, N24617);
xor XOR2 (N24625, N24624, N9313);
and AND2 (N24626, N24616, N21779);
xor XOR2 (N24627, N24609, N1450);
nor NOR3 (N24628, N24622, N12801, N2148);
and AND2 (N24629, N24611, N5882);
or OR3 (N24630, N24615, N6249, N11538);
xor XOR2 (N24631, N24627, N19315);
not NOT1 (N24632, N24625);
nor NOR3 (N24633, N24631, N16990, N3112);
nor NOR4 (N24634, N24621, N12734, N18153, N20102);
nor NOR2 (N24635, N24628, N18140);
not NOT1 (N24636, N24620);
xor XOR2 (N24637, N24635, N9039);
nand NAND4 (N24638, N24637, N11906, N22765, N6825);
buf BUF1 (N24639, N24636);
buf BUF1 (N24640, N24630);
xor XOR2 (N24641, N24629, N11772);
and AND3 (N24642, N24632, N1694, N18055);
not NOT1 (N24643, N24641);
xor XOR2 (N24644, N24643, N17482);
nor NOR4 (N24645, N24640, N10176, N23226, N13236);
nand NAND4 (N24646, N24639, N8295, N1138, N1381);
nand NAND2 (N24647, N24645, N544);
and AND4 (N24648, N24646, N4294, N10961, N22154);
nand NAND4 (N24649, N24648, N21429, N22485, N10464);
buf BUF1 (N24650, N24626);
xor XOR2 (N24651, N24649, N9507);
or OR3 (N24652, N24619, N3405, N6677);
nand NAND2 (N24653, N24644, N16577);
nor NOR4 (N24654, N24642, N23348, N17352, N17106);
not NOT1 (N24655, N24652);
buf BUF1 (N24656, N24654);
nand NAND4 (N24657, N24651, N17845, N593, N16662);
nand NAND3 (N24658, N24647, N6539, N9066);
buf BUF1 (N24659, N24633);
nor NOR4 (N24660, N24634, N11974, N16727, N22067);
nor NOR4 (N24661, N24653, N703, N24524, N17763);
not NOT1 (N24662, N24659);
nand NAND3 (N24663, N24662, N2697, N16009);
nor NOR4 (N24664, N24656, N15627, N18527, N10798);
or OR3 (N24665, N24660, N3564, N21405);
or OR3 (N24666, N24623, N22192, N4095);
nand NAND2 (N24667, N24650, N18416);
buf BUF1 (N24668, N24667);
or OR2 (N24669, N24661, N21153);
buf BUF1 (N24670, N24638);
nor NOR4 (N24671, N24657, N14920, N23492, N8727);
nor NOR2 (N24672, N24666, N3787);
nand NAND4 (N24673, N24668, N21994, N3234, N21648);
nor NOR4 (N24674, N24665, N6508, N5041, N23937);
nand NAND4 (N24675, N24674, N14437, N5595, N8693);
nor NOR3 (N24676, N24655, N17635, N8431);
nand NAND3 (N24677, N24675, N2812, N21506);
buf BUF1 (N24678, N24658);
nor NOR4 (N24679, N24672, N6994, N23729, N8979);
not NOT1 (N24680, N24678);
or OR4 (N24681, N24680, N5060, N19740, N22748);
not NOT1 (N24682, N24677);
nand NAND4 (N24683, N24669, N18748, N16, N11730);
and AND4 (N24684, N24679, N4721, N799, N14892);
not NOT1 (N24685, N24671);
nor NOR4 (N24686, N24682, N22230, N16178, N21255);
nand NAND3 (N24687, N24663, N8840, N14342);
nand NAND3 (N24688, N24683, N7199, N23564);
and AND4 (N24689, N24687, N23445, N5918, N17498);
buf BUF1 (N24690, N24673);
nand NAND3 (N24691, N24685, N7719, N3670);
not NOT1 (N24692, N24676);
nor NOR2 (N24693, N24684, N532);
not NOT1 (N24694, N24690);
nand NAND3 (N24695, N24692, N5283, N10644);
xor XOR2 (N24696, N24694, N13458);
and AND3 (N24697, N24693, N20826, N491);
buf BUF1 (N24698, N24696);
or OR3 (N24699, N24689, N12601, N14931);
or OR4 (N24700, N24691, N19819, N16836, N9978);
nand NAND3 (N24701, N24697, N5940, N6035);
and AND2 (N24702, N24670, N3099);
xor XOR2 (N24703, N24698, N14816);
not NOT1 (N24704, N24681);
xor XOR2 (N24705, N24700, N662);
nor NOR2 (N24706, N24705, N1380);
or OR3 (N24707, N24704, N16317, N23190);
xor XOR2 (N24708, N24699, N138);
and AND4 (N24709, N24701, N21189, N14646, N14727);
not NOT1 (N24710, N24688);
not NOT1 (N24711, N24708);
xor XOR2 (N24712, N24703, N20647);
not NOT1 (N24713, N24707);
not NOT1 (N24714, N24702);
buf BUF1 (N24715, N24686);
buf BUF1 (N24716, N24706);
nor NOR2 (N24717, N24710, N22898);
not NOT1 (N24718, N24716);
or OR2 (N24719, N24711, N23851);
buf BUF1 (N24720, N24664);
and AND2 (N24721, N24720, N23528);
xor XOR2 (N24722, N24714, N11348);
nand NAND2 (N24723, N24719, N2121);
or OR3 (N24724, N24718, N11082, N11032);
nor NOR2 (N24725, N24709, N14245);
or OR3 (N24726, N24725, N16326, N7112);
not NOT1 (N24727, N24723);
nand NAND4 (N24728, N24726, N19552, N8785, N22956);
not NOT1 (N24729, N24724);
nor NOR2 (N24730, N24717, N15802);
nor NOR2 (N24731, N24727, N20229);
not NOT1 (N24732, N24722);
and AND3 (N24733, N24713, N555, N20712);
nand NAND3 (N24734, N24729, N17149, N11908);
not NOT1 (N24735, N24728);
or OR4 (N24736, N24732, N16963, N17897, N7651);
not NOT1 (N24737, N24731);
not NOT1 (N24738, N24735);
nor NOR2 (N24739, N24736, N11676);
not NOT1 (N24740, N24712);
xor XOR2 (N24741, N24733, N22509);
not NOT1 (N24742, N24740);
not NOT1 (N24743, N24738);
and AND3 (N24744, N24743, N13542, N19220);
nand NAND4 (N24745, N24741, N12254, N3771, N10608);
and AND4 (N24746, N24730, N9525, N18601, N15454);
nor NOR3 (N24747, N24745, N4081, N13402);
nor NOR3 (N24748, N24739, N13565, N8417);
not NOT1 (N24749, N24734);
xor XOR2 (N24750, N24695, N4038);
buf BUF1 (N24751, N24747);
buf BUF1 (N24752, N24737);
or OR4 (N24753, N24749, N3136, N6466, N19423);
nand NAND4 (N24754, N24746, N18636, N17675, N7606);
not NOT1 (N24755, N24754);
buf BUF1 (N24756, N24750);
xor XOR2 (N24757, N24755, N11026);
and AND4 (N24758, N24721, N23047, N4899, N8965);
nand NAND3 (N24759, N24744, N22626, N9802);
nor NOR2 (N24760, N24758, N7310);
buf BUF1 (N24761, N24753);
and AND3 (N24762, N24760, N18416, N17937);
buf BUF1 (N24763, N24761);
or OR2 (N24764, N24752, N19291);
not NOT1 (N24765, N24759);
xor XOR2 (N24766, N24742, N12940);
xor XOR2 (N24767, N24757, N3958);
not NOT1 (N24768, N24715);
and AND3 (N24769, N24766, N9978, N17936);
or OR4 (N24770, N24748, N21135, N21457, N24495);
or OR4 (N24771, N24763, N18890, N20846, N9436);
xor XOR2 (N24772, N24770, N1465);
nand NAND2 (N24773, N24756, N19517);
not NOT1 (N24774, N24772);
buf BUF1 (N24775, N24767);
xor XOR2 (N24776, N24768, N14230);
or OR3 (N24777, N24776, N3676, N21816);
and AND3 (N24778, N24771, N17079, N15511);
not NOT1 (N24779, N24765);
xor XOR2 (N24780, N24764, N23234);
buf BUF1 (N24781, N24773);
not NOT1 (N24782, N24774);
nand NAND3 (N24783, N24779, N17349, N1366);
nand NAND3 (N24784, N24769, N4901, N14260);
or OR4 (N24785, N24784, N12461, N11639, N2399);
xor XOR2 (N24786, N24783, N4893);
nor NOR3 (N24787, N24751, N12164, N16982);
nand NAND2 (N24788, N24775, N16771);
nand NAND2 (N24789, N24762, N19919);
and AND3 (N24790, N24786, N12262, N3518);
and AND2 (N24791, N24788, N4631);
and AND2 (N24792, N24787, N17107);
buf BUF1 (N24793, N24789);
xor XOR2 (N24794, N24782, N19836);
nand NAND4 (N24795, N24785, N14382, N220, N3866);
not NOT1 (N24796, N24791);
or OR4 (N24797, N24790, N473, N15415, N24488);
or OR4 (N24798, N24796, N2379, N20438, N18273);
buf BUF1 (N24799, N24781);
nor NOR3 (N24800, N24778, N1353, N9811);
nor NOR4 (N24801, N24793, N14111, N6395, N22307);
nand NAND2 (N24802, N24799, N2234);
nor NOR3 (N24803, N24795, N13096, N16903);
buf BUF1 (N24804, N24797);
or OR4 (N24805, N24794, N22972, N22972, N19998);
or OR4 (N24806, N24800, N3999, N20329, N6630);
and AND4 (N24807, N24777, N19023, N8423, N15079);
xor XOR2 (N24808, N24803, N999);
or OR3 (N24809, N24792, N8023, N23763);
nor NOR3 (N24810, N24780, N12891, N15959);
and AND2 (N24811, N24804, N3165);
buf BUF1 (N24812, N24802);
and AND3 (N24813, N24809, N10030, N544);
nor NOR4 (N24814, N24801, N6973, N8691, N4327);
nand NAND2 (N24815, N24806, N16254);
and AND4 (N24816, N24813, N13021, N21480, N21018);
nor NOR2 (N24817, N24812, N1803);
and AND3 (N24818, N24808, N1048, N12815);
nor NOR2 (N24819, N24807, N5990);
buf BUF1 (N24820, N24811);
buf BUF1 (N24821, N24817);
buf BUF1 (N24822, N24820);
not NOT1 (N24823, N24821);
xor XOR2 (N24824, N24805, N10039);
or OR4 (N24825, N24815, N17435, N6607, N18017);
not NOT1 (N24826, N24816);
nor NOR3 (N24827, N24798, N17831, N8639);
not NOT1 (N24828, N24823);
xor XOR2 (N24829, N24814, N7784);
nand NAND3 (N24830, N24819, N23785, N9129);
buf BUF1 (N24831, N24827);
or OR3 (N24832, N24831, N23144, N267);
not NOT1 (N24833, N24825);
or OR4 (N24834, N24832, N20363, N14848, N21921);
not NOT1 (N24835, N24810);
nor NOR3 (N24836, N24829, N14312, N3022);
nor NOR4 (N24837, N24834, N1394, N7990, N8949);
not NOT1 (N24838, N24830);
nor NOR2 (N24839, N24822, N1649);
or OR2 (N24840, N24828, N15789);
xor XOR2 (N24841, N24838, N24294);
or OR4 (N24842, N24818, N8959, N11309, N15497);
buf BUF1 (N24843, N24824);
or OR4 (N24844, N24835, N10194, N10039, N6761);
and AND4 (N24845, N24842, N21038, N4979, N24661);
nand NAND3 (N24846, N24837, N20094, N24536);
or OR4 (N24847, N24846, N4854, N13677, N565);
and AND3 (N24848, N24836, N3261, N17588);
not NOT1 (N24849, N24840);
nor NOR4 (N24850, N24843, N333, N10456, N4876);
or OR3 (N24851, N24844, N7202, N22905);
nand NAND4 (N24852, N24826, N5232, N12354, N2741);
or OR3 (N24853, N24851, N24113, N12564);
xor XOR2 (N24854, N24850, N15281);
not NOT1 (N24855, N24854);
xor XOR2 (N24856, N24849, N1946);
xor XOR2 (N24857, N24839, N3338);
xor XOR2 (N24858, N24841, N7192);
nor NOR3 (N24859, N24857, N21166, N14073);
and AND3 (N24860, N24855, N7011, N10277);
not NOT1 (N24861, N24858);
buf BUF1 (N24862, N24845);
buf BUF1 (N24863, N24861);
nor NOR2 (N24864, N24860, N20447);
nand NAND2 (N24865, N24859, N9223);
nand NAND4 (N24866, N24856, N8214, N10875, N21201);
nor NOR4 (N24867, N24862, N3102, N15020, N1751);
and AND2 (N24868, N24866, N4837);
buf BUF1 (N24869, N24868);
xor XOR2 (N24870, N24833, N19508);
xor XOR2 (N24871, N24852, N220);
nor NOR2 (N24872, N24848, N9786);
nand NAND4 (N24873, N24853, N11979, N4548, N13025);
nor NOR3 (N24874, N24870, N4458, N19471);
xor XOR2 (N24875, N24847, N22339);
buf BUF1 (N24876, N24863);
and AND4 (N24877, N24867, N20133, N11147, N24219);
nor NOR3 (N24878, N24864, N17789, N17634);
buf BUF1 (N24879, N24873);
nor NOR3 (N24880, N24876, N4, N21915);
xor XOR2 (N24881, N24871, N24161);
nor NOR3 (N24882, N24874, N6242, N14769);
nand NAND3 (N24883, N24877, N215, N9139);
and AND4 (N24884, N24883, N14067, N18905, N24781);
buf BUF1 (N24885, N24881);
not NOT1 (N24886, N24869);
nand NAND2 (N24887, N24885, N17962);
buf BUF1 (N24888, N24887);
nor NOR4 (N24889, N24878, N22927, N13465, N13609);
nand NAND2 (N24890, N24879, N11985);
nand NAND4 (N24891, N24886, N17132, N2407, N5838);
not NOT1 (N24892, N24891);
buf BUF1 (N24893, N24882);
not NOT1 (N24894, N24865);
or OR4 (N24895, N24894, N10545, N701, N426);
xor XOR2 (N24896, N24884, N3572);
buf BUF1 (N24897, N24889);
nor NOR2 (N24898, N24872, N12304);
or OR3 (N24899, N24890, N18785, N23399);
buf BUF1 (N24900, N24899);
nor NOR2 (N24901, N24893, N10563);
buf BUF1 (N24902, N24897);
not NOT1 (N24903, N24900);
nand NAND4 (N24904, N24901, N3595, N17927, N5785);
buf BUF1 (N24905, N24904);
nand NAND4 (N24906, N24888, N5134, N15638, N11951);
nor NOR2 (N24907, N24875, N18015);
nand NAND3 (N24908, N24892, N16806, N7412);
or OR2 (N24909, N24895, N7137);
not NOT1 (N24910, N24905);
and AND2 (N24911, N24909, N7520);
nand NAND3 (N24912, N24903, N13446, N8732);
nor NOR2 (N24913, N24910, N14168);
nor NOR4 (N24914, N24898, N4774, N11433, N9329);
nand NAND4 (N24915, N24896, N21573, N12932, N23665);
buf BUF1 (N24916, N24880);
not NOT1 (N24917, N24914);
or OR3 (N24918, N24913, N8383, N5614);
nor NOR4 (N24919, N24908, N13345, N4350, N24854);
not NOT1 (N24920, N24912);
and AND4 (N24921, N24902, N11883, N16814, N20879);
xor XOR2 (N24922, N24917, N7174);
or OR4 (N24923, N24922, N24196, N23545, N3840);
xor XOR2 (N24924, N24921, N21403);
xor XOR2 (N24925, N24915, N12713);
nand NAND4 (N24926, N24906, N7618, N21282, N7332);
nand NAND3 (N24927, N24920, N9541, N24740);
nand NAND4 (N24928, N24916, N23199, N3912, N18312);
or OR4 (N24929, N24911, N7523, N11463, N3088);
or OR2 (N24930, N24923, N24567);
or OR4 (N24931, N24907, N21366, N6686, N11412);
buf BUF1 (N24932, N24931);
and AND3 (N24933, N24928, N23012, N93);
buf BUF1 (N24934, N24919);
nand NAND4 (N24935, N24924, N181, N4587, N7956);
xor XOR2 (N24936, N24935, N11615);
buf BUF1 (N24937, N24933);
not NOT1 (N24938, N24936);
xor XOR2 (N24939, N24937, N9672);
or OR4 (N24940, N24932, N3391, N24766, N24588);
or OR3 (N24941, N24927, N14109, N14060);
nor NOR2 (N24942, N24926, N1937);
nand NAND4 (N24943, N24925, N20494, N9279, N5751);
buf BUF1 (N24944, N24939);
and AND2 (N24945, N24930, N23025);
xor XOR2 (N24946, N24945, N20879);
nand NAND2 (N24947, N24918, N16216);
nor NOR4 (N24948, N24946, N1024, N3030, N7800);
nor NOR3 (N24949, N24929, N12465, N15176);
not NOT1 (N24950, N24940);
buf BUF1 (N24951, N24949);
and AND2 (N24952, N24943, N1746);
nor NOR3 (N24953, N24942, N15917, N13269);
nand NAND2 (N24954, N24944, N443);
nor NOR4 (N24955, N24953, N4622, N4033, N7257);
and AND2 (N24956, N24950, N12411);
nand NAND4 (N24957, N24934, N1457, N15253, N11615);
nor NOR3 (N24958, N24954, N19546, N8067);
or OR4 (N24959, N24958, N12049, N15942, N21093);
xor XOR2 (N24960, N24955, N17475);
buf BUF1 (N24961, N24941);
buf BUF1 (N24962, N24957);
buf BUF1 (N24963, N24959);
buf BUF1 (N24964, N24960);
nand NAND4 (N24965, N24961, N14991, N23056, N13207);
xor XOR2 (N24966, N24938, N7335);
not NOT1 (N24967, N24947);
buf BUF1 (N24968, N24956);
nand NAND2 (N24969, N24963, N15457);
nand NAND3 (N24970, N24952, N15984, N379);
nor NOR4 (N24971, N24968, N4181, N16108, N15390);
xor XOR2 (N24972, N24966, N20989);
buf BUF1 (N24973, N24972);
not NOT1 (N24974, N24973);
nand NAND4 (N24975, N24971, N13712, N14144, N24434);
nand NAND4 (N24976, N24964, N9024, N11584, N3841);
xor XOR2 (N24977, N24975, N10977);
and AND2 (N24978, N24962, N361);
nand NAND3 (N24979, N24965, N6414, N10515);
nand NAND4 (N24980, N24951, N15303, N8054, N4634);
nand NAND2 (N24981, N24978, N17085);
nand NAND2 (N24982, N24980, N19326);
or OR3 (N24983, N24981, N23943, N23460);
and AND3 (N24984, N24974, N8523, N11073);
nor NOR4 (N24985, N24982, N22737, N21861, N2933);
buf BUF1 (N24986, N24976);
nor NOR2 (N24987, N24948, N3608);
or OR3 (N24988, N24985, N18682, N3940);
xor XOR2 (N24989, N24987, N16699);
buf BUF1 (N24990, N24983);
or OR4 (N24991, N24988, N21844, N22025, N4056);
and AND2 (N24992, N24990, N21677);
buf BUF1 (N24993, N24970);
xor XOR2 (N24994, N24989, N7933);
buf BUF1 (N24995, N24993);
buf BUF1 (N24996, N24969);
not NOT1 (N24997, N24992);
nor NOR3 (N24998, N24984, N18322, N2740);
or OR4 (N24999, N24986, N16700, N1254, N15981);
and AND4 (N25000, N24995, N3834, N19782, N124);
nand NAND4 (N25001, N24979, N12042, N23698, N21031);
or OR3 (N25002, N24996, N9258, N15097);
nor NOR2 (N25003, N24997, N16847);
nand NAND3 (N25004, N25000, N16903, N5923);
xor XOR2 (N25005, N25004, N24199);
and AND3 (N25006, N25005, N7224, N19267);
not NOT1 (N25007, N24991);
not NOT1 (N25008, N25001);
or OR3 (N25009, N25006, N21148, N18604);
nor NOR4 (N25010, N24998, N7396, N2580, N6715);
nand NAND4 (N25011, N25003, N13139, N6951, N6951);
xor XOR2 (N25012, N24999, N15911);
buf BUF1 (N25013, N25012);
buf BUF1 (N25014, N24977);
or OR2 (N25015, N25014, N13176);
buf BUF1 (N25016, N25009);
nor NOR2 (N25017, N25015, N8986);
not NOT1 (N25018, N25013);
nand NAND2 (N25019, N25002, N2700);
or OR2 (N25020, N25019, N5611);
xor XOR2 (N25021, N25018, N16196);
buf BUF1 (N25022, N25021);
nor NOR4 (N25023, N25022, N3208, N10693, N10485);
not NOT1 (N25024, N25007);
or OR4 (N25025, N25020, N11316, N12119, N23955);
buf BUF1 (N25026, N25017);
buf BUF1 (N25027, N25026);
or OR4 (N25028, N25011, N3646, N8836, N2116);
or OR3 (N25029, N25024, N14042, N17429);
or OR3 (N25030, N25028, N19280, N9069);
and AND3 (N25031, N25023, N1516, N2538);
or OR4 (N25032, N25030, N888, N11408, N11709);
nor NOR4 (N25033, N24994, N7115, N9131, N4610);
not NOT1 (N25034, N25032);
not NOT1 (N25035, N25033);
not NOT1 (N25036, N25016);
nand NAND4 (N25037, N25035, N20590, N7378, N1469);
nand NAND3 (N25038, N25036, N5921, N11632);
or OR3 (N25039, N25037, N20590, N14229);
or OR2 (N25040, N24967, N13633);
nand NAND3 (N25041, N25040, N12192, N9630);
and AND2 (N25042, N25029, N12496);
and AND4 (N25043, N25008, N2713, N16799, N12613);
nor NOR3 (N25044, N25038, N16513, N1283);
or OR3 (N25045, N25010, N22407, N18620);
and AND3 (N25046, N25044, N9631, N18299);
and AND3 (N25047, N25042, N3389, N10106);
nand NAND3 (N25048, N25027, N16929, N8118);
nand NAND2 (N25049, N25046, N19366);
xor XOR2 (N25050, N25045, N18651);
nand NAND3 (N25051, N25025, N18449, N12847);
nand NAND2 (N25052, N25039, N13);
not NOT1 (N25053, N25034);
xor XOR2 (N25054, N25041, N18260);
and AND4 (N25055, N25048, N18532, N24455, N14529);
nand NAND3 (N25056, N25047, N9149, N3967);
nand NAND3 (N25057, N25049, N13572, N14261);
or OR3 (N25058, N25055, N13084, N5484);
not NOT1 (N25059, N25053);
not NOT1 (N25060, N25043);
and AND2 (N25061, N25050, N19565);
xor XOR2 (N25062, N25059, N620);
nand NAND3 (N25063, N25061, N22280, N780);
and AND3 (N25064, N25052, N9526, N15290);
nand NAND3 (N25065, N25062, N18692, N13525);
nand NAND2 (N25066, N25060, N19577);
xor XOR2 (N25067, N25031, N2800);
nor NOR3 (N25068, N25065, N271, N3173);
nand NAND2 (N25069, N25058, N10260);
buf BUF1 (N25070, N25069);
not NOT1 (N25071, N25056);
xor XOR2 (N25072, N25071, N8720);
nand NAND2 (N25073, N25067, N10862);
nand NAND3 (N25074, N25072, N17982, N5592);
nand NAND4 (N25075, N25051, N11650, N22221, N9556);
nand NAND4 (N25076, N25075, N12047, N8943, N12767);
not NOT1 (N25077, N25054);
nor NOR2 (N25078, N25068, N2395);
nand NAND2 (N25079, N25077, N19236);
and AND4 (N25080, N25073, N7077, N3835, N22448);
or OR4 (N25081, N25078, N19923, N7542, N8259);
or OR3 (N25082, N25063, N5537, N10132);
nor NOR3 (N25083, N25070, N20402, N18547);
not NOT1 (N25084, N25080);
nor NOR3 (N25085, N25076, N8880, N11071);
nor NOR3 (N25086, N25081, N21740, N513);
not NOT1 (N25087, N25084);
and AND4 (N25088, N25082, N3674, N17294, N9734);
and AND3 (N25089, N25057, N24580, N15278);
and AND4 (N25090, N25064, N913, N15509, N7872);
nor NOR4 (N25091, N25086, N4200, N8306, N18428);
not NOT1 (N25092, N25090);
buf BUF1 (N25093, N25085);
nor NOR4 (N25094, N25089, N10234, N12076, N15119);
nor NOR3 (N25095, N25094, N24114, N19762);
xor XOR2 (N25096, N25095, N19876);
or OR3 (N25097, N25092, N24971, N16725);
and AND3 (N25098, N25097, N21309, N2306);
nand NAND2 (N25099, N25083, N5843);
nor NOR2 (N25100, N25066, N4052);
buf BUF1 (N25101, N25079);
buf BUF1 (N25102, N25100);
not NOT1 (N25103, N25102);
xor XOR2 (N25104, N25074, N13048);
xor XOR2 (N25105, N25099, N812);
or OR4 (N25106, N25093, N1485, N17198, N270);
or OR2 (N25107, N25087, N20577);
and AND4 (N25108, N25104, N3137, N1509, N14016);
not NOT1 (N25109, N25103);
nor NOR3 (N25110, N25088, N10235, N21967);
buf BUF1 (N25111, N25109);
nor NOR2 (N25112, N25096, N6208);
nand NAND2 (N25113, N25110, N22831);
nor NOR3 (N25114, N25105, N8364, N10912);
nand NAND2 (N25115, N25108, N19951);
or OR2 (N25116, N25101, N22421);
not NOT1 (N25117, N25098);
xor XOR2 (N25118, N25107, N21405);
nand NAND3 (N25119, N25115, N7560, N15850);
buf BUF1 (N25120, N25116);
and AND3 (N25121, N25113, N1614, N9608);
or OR4 (N25122, N25118, N8379, N7999, N1046);
or OR2 (N25123, N25122, N20621);
buf BUF1 (N25124, N25120);
or OR3 (N25125, N25091, N17533, N18630);
or OR2 (N25126, N25124, N9358);
and AND4 (N25127, N25125, N16785, N17885, N14939);
and AND2 (N25128, N25126, N16598);
or OR4 (N25129, N25119, N4256, N18304, N6741);
and AND3 (N25130, N25123, N7215, N5933);
or OR3 (N25131, N25121, N21011, N286);
xor XOR2 (N25132, N25129, N22297);
xor XOR2 (N25133, N25132, N24220);
or OR2 (N25134, N25112, N10920);
and AND4 (N25135, N25106, N12567, N7936, N6486);
or OR2 (N25136, N25114, N20031);
buf BUF1 (N25137, N25136);
nor NOR2 (N25138, N25131, N6917);
and AND3 (N25139, N25117, N11535, N20035);
not NOT1 (N25140, N25139);
not NOT1 (N25141, N25134);
nand NAND2 (N25142, N25137, N5394);
not NOT1 (N25143, N25142);
xor XOR2 (N25144, N25138, N12223);
or OR2 (N25145, N25127, N23580);
nand NAND3 (N25146, N25130, N23551, N12563);
nor NOR3 (N25147, N25128, N7082, N377);
not NOT1 (N25148, N25141);
nor NOR3 (N25149, N25146, N8606, N8415);
and AND4 (N25150, N25148, N17992, N6025, N13613);
not NOT1 (N25151, N25149);
nand NAND2 (N25152, N25111, N3702);
and AND2 (N25153, N25143, N18017);
xor XOR2 (N25154, N25151, N8969);
not NOT1 (N25155, N25140);
not NOT1 (N25156, N25135);
or OR3 (N25157, N25152, N1045, N10605);
and AND4 (N25158, N25155, N12855, N5802, N2658);
and AND2 (N25159, N25154, N6289);
or OR4 (N25160, N25158, N10564, N21269, N15210);
buf BUF1 (N25161, N25144);
buf BUF1 (N25162, N25147);
and AND4 (N25163, N25153, N24321, N13235, N20809);
xor XOR2 (N25164, N25145, N21911);
or OR2 (N25165, N25162, N20228);
nand NAND4 (N25166, N25164, N7984, N2683, N24312);
not NOT1 (N25167, N25160);
xor XOR2 (N25168, N25161, N17990);
and AND4 (N25169, N25159, N20761, N14582, N19505);
xor XOR2 (N25170, N25166, N23607);
xor XOR2 (N25171, N25169, N7781);
and AND3 (N25172, N25150, N20649, N22683);
nor NOR3 (N25173, N25172, N17263, N19847);
nor NOR3 (N25174, N25156, N17154, N12832);
or OR3 (N25175, N25165, N11901, N14071);
buf BUF1 (N25176, N25171);
nor NOR2 (N25177, N25170, N24193);
nor NOR3 (N25178, N25167, N14762, N4080);
nor NOR2 (N25179, N25133, N23437);
not NOT1 (N25180, N25173);
or OR3 (N25181, N25176, N9956, N15471);
or OR3 (N25182, N25157, N22740, N11247);
xor XOR2 (N25183, N25181, N19729);
not NOT1 (N25184, N25174);
or OR4 (N25185, N25179, N7663, N10277, N23439);
not NOT1 (N25186, N25175);
and AND2 (N25187, N25183, N10101);
or OR4 (N25188, N25178, N4144, N18844, N22962);
nor NOR4 (N25189, N25182, N8899, N2772, N14863);
buf BUF1 (N25190, N25177);
buf BUF1 (N25191, N25180);
not NOT1 (N25192, N25189);
nor NOR3 (N25193, N25186, N7010, N3506);
nor NOR4 (N25194, N25191, N10688, N24888, N17946);
or OR4 (N25195, N25188, N18689, N16832, N2138);
nor NOR3 (N25196, N25194, N5666, N10212);
buf BUF1 (N25197, N25187);
nand NAND4 (N25198, N25185, N7545, N5783, N14286);
buf BUF1 (N25199, N25197);
buf BUF1 (N25200, N25184);
not NOT1 (N25201, N25196);
nand NAND3 (N25202, N25195, N18862, N13036);
and AND3 (N25203, N25193, N16807, N7403);
nor NOR3 (N25204, N25200, N2979, N24738);
or OR4 (N25205, N25198, N22887, N7776, N13191);
and AND3 (N25206, N25168, N2263, N5511);
xor XOR2 (N25207, N25204, N4552);
buf BUF1 (N25208, N25202);
nand NAND4 (N25209, N25201, N12241, N11008, N2830);
nor NOR2 (N25210, N25163, N23462);
not NOT1 (N25211, N25190);
nand NAND3 (N25212, N25206, N2914, N5273);
nand NAND2 (N25213, N25209, N13899);
xor XOR2 (N25214, N25210, N14517);
and AND3 (N25215, N25208, N22327, N8246);
and AND2 (N25216, N25192, N19202);
xor XOR2 (N25217, N25211, N8435);
xor XOR2 (N25218, N25199, N5310);
buf BUF1 (N25219, N25205);
not NOT1 (N25220, N25216);
buf BUF1 (N25221, N25214);
xor XOR2 (N25222, N25217, N18305);
nor NOR2 (N25223, N25215, N9354);
xor XOR2 (N25224, N25203, N3024);
nor NOR4 (N25225, N25212, N5726, N6210, N20334);
buf BUF1 (N25226, N25223);
nor NOR3 (N25227, N25221, N24720, N4753);
xor XOR2 (N25228, N25220, N2447);
and AND2 (N25229, N25225, N4897);
and AND4 (N25230, N25226, N18410, N23632, N16875);
not NOT1 (N25231, N25207);
xor XOR2 (N25232, N25228, N5086);
not NOT1 (N25233, N25218);
and AND4 (N25234, N25231, N17337, N20644, N1145);
buf BUF1 (N25235, N25229);
nor NOR2 (N25236, N25230, N23307);
nor NOR3 (N25237, N25213, N17345, N1610);
or OR4 (N25238, N25227, N8855, N21871, N13859);
nand NAND4 (N25239, N25219, N14638, N7425, N24996);
nand NAND4 (N25240, N25238, N19283, N21862, N2483);
nand NAND4 (N25241, N25233, N23901, N10527, N76);
not NOT1 (N25242, N25234);
buf BUF1 (N25243, N25242);
nand NAND3 (N25244, N25239, N16752, N7679);
xor XOR2 (N25245, N25244, N6825);
or OR4 (N25246, N25232, N21901, N7123, N18603);
and AND4 (N25247, N25246, N23069, N6902, N11086);
not NOT1 (N25248, N25222);
or OR4 (N25249, N25241, N4910, N14693, N21506);
or OR3 (N25250, N25237, N15422, N2906);
buf BUF1 (N25251, N25224);
nor NOR2 (N25252, N25249, N3109);
nand NAND2 (N25253, N25240, N7482);
not NOT1 (N25254, N25250);
or OR4 (N25255, N25253, N24996, N15011, N519);
not NOT1 (N25256, N25248);
buf BUF1 (N25257, N25247);
or OR2 (N25258, N25254, N22260);
and AND2 (N25259, N25255, N24343);
buf BUF1 (N25260, N25257);
nor NOR2 (N25261, N25251, N3960);
or OR4 (N25262, N25258, N13060, N3352, N17266);
xor XOR2 (N25263, N25256, N7165);
buf BUF1 (N25264, N25252);
and AND3 (N25265, N25236, N21800, N6258);
or OR2 (N25266, N25262, N9724);
buf BUF1 (N25267, N25243);
and AND2 (N25268, N25266, N8340);
nand NAND2 (N25269, N25265, N5875);
buf BUF1 (N25270, N25269);
and AND3 (N25271, N25260, N336, N7921);
buf BUF1 (N25272, N25267);
xor XOR2 (N25273, N25263, N11817);
or OR2 (N25274, N25273, N9852);
nand NAND4 (N25275, N25272, N641, N1398, N18980);
or OR2 (N25276, N25268, N2045);
nor NOR4 (N25277, N25276, N5053, N19764, N21324);
not NOT1 (N25278, N25245);
buf BUF1 (N25279, N25275);
or OR2 (N25280, N25278, N8979);
not NOT1 (N25281, N25261);
xor XOR2 (N25282, N25280, N11584);
or OR3 (N25283, N25279, N18058, N14839);
and AND2 (N25284, N25282, N13240);
or OR4 (N25285, N25264, N6114, N24049, N15984);
xor XOR2 (N25286, N25283, N16292);
or OR4 (N25287, N25235, N3493, N20264, N19495);
or OR3 (N25288, N25287, N14409, N16858);
and AND2 (N25289, N25288, N4642);
xor XOR2 (N25290, N25271, N22357);
xor XOR2 (N25291, N25286, N11446);
nor NOR3 (N25292, N25281, N21565, N23230);
buf BUF1 (N25293, N25259);
nor NOR2 (N25294, N25285, N13359);
or OR4 (N25295, N25274, N24281, N3212, N19530);
or OR3 (N25296, N25277, N17975, N7560);
and AND2 (N25297, N25290, N3671);
not NOT1 (N25298, N25270);
nand NAND2 (N25299, N25284, N3710);
and AND4 (N25300, N25297, N22183, N17320, N2680);
xor XOR2 (N25301, N25295, N23577);
nor NOR2 (N25302, N25299, N13548);
buf BUF1 (N25303, N25300);
buf BUF1 (N25304, N25303);
buf BUF1 (N25305, N25296);
not NOT1 (N25306, N25301);
not NOT1 (N25307, N25289);
buf BUF1 (N25308, N25293);
xor XOR2 (N25309, N25307, N600);
xor XOR2 (N25310, N25292, N10985);
buf BUF1 (N25311, N25305);
nand NAND3 (N25312, N25308, N3969, N7257);
not NOT1 (N25313, N25294);
buf BUF1 (N25314, N25312);
not NOT1 (N25315, N25304);
nor NOR4 (N25316, N25311, N15081, N24318, N20026);
buf BUF1 (N25317, N25314);
or OR4 (N25318, N25302, N22469, N1629, N8320);
nand NAND3 (N25319, N25315, N17021, N11298);
nand NAND4 (N25320, N25319, N9085, N16854, N9917);
or OR4 (N25321, N25291, N3080, N24934, N17288);
nor NOR3 (N25322, N25317, N19709, N18771);
nor NOR2 (N25323, N25322, N4317);
nor NOR2 (N25324, N25309, N16284);
or OR4 (N25325, N25318, N1073, N2481, N15420);
and AND2 (N25326, N25320, N19327);
xor XOR2 (N25327, N25298, N3286);
buf BUF1 (N25328, N25310);
buf BUF1 (N25329, N25328);
nor NOR4 (N25330, N25313, N20248, N9759, N8036);
or OR2 (N25331, N25326, N15569);
not NOT1 (N25332, N25306);
not NOT1 (N25333, N25321);
buf BUF1 (N25334, N25329);
buf BUF1 (N25335, N25316);
not NOT1 (N25336, N25335);
or OR2 (N25337, N25332, N1046);
or OR4 (N25338, N25336, N6365, N19868, N3033);
xor XOR2 (N25339, N25331, N18342);
buf BUF1 (N25340, N25339);
nor NOR2 (N25341, N25327, N23887);
xor XOR2 (N25342, N25337, N12380);
buf BUF1 (N25343, N25325);
and AND2 (N25344, N25323, N23631);
not NOT1 (N25345, N25344);
buf BUF1 (N25346, N25340);
and AND4 (N25347, N25330, N23707, N7778, N5577);
nor NOR3 (N25348, N25324, N17142, N404);
nand NAND2 (N25349, N25334, N7207);
nand NAND2 (N25350, N25341, N22575);
not NOT1 (N25351, N25348);
nand NAND4 (N25352, N25338, N12233, N11635, N3456);
buf BUF1 (N25353, N25347);
not NOT1 (N25354, N25342);
not NOT1 (N25355, N25353);
buf BUF1 (N25356, N25345);
not NOT1 (N25357, N25346);
not NOT1 (N25358, N25352);
nor NOR3 (N25359, N25357, N1194, N3250);
or OR3 (N25360, N25355, N3567, N19727);
nand NAND3 (N25361, N25358, N20438, N8878);
buf BUF1 (N25362, N25354);
or OR4 (N25363, N25359, N1514, N6300, N12342);
xor XOR2 (N25364, N25349, N3543);
nand NAND4 (N25365, N25356, N11099, N10690, N19449);
nand NAND4 (N25366, N25365, N14945, N20997, N24443);
nand NAND2 (N25367, N25363, N13027);
buf BUF1 (N25368, N25350);
xor XOR2 (N25369, N25366, N9486);
nor NOR2 (N25370, N25343, N5114);
xor XOR2 (N25371, N25367, N23746);
or OR3 (N25372, N25370, N8141, N12663);
nand NAND2 (N25373, N25360, N3620);
nor NOR4 (N25374, N25362, N16837, N9577, N15534);
not NOT1 (N25375, N25364);
or OR2 (N25376, N25371, N10485);
nor NOR3 (N25377, N25333, N6086, N5345);
buf BUF1 (N25378, N25368);
nand NAND2 (N25379, N25373, N13261);
nor NOR4 (N25380, N25377, N13380, N4952, N8522);
buf BUF1 (N25381, N25379);
not NOT1 (N25382, N25376);
buf BUF1 (N25383, N25351);
xor XOR2 (N25384, N25375, N16284);
xor XOR2 (N25385, N25369, N20265);
xor XOR2 (N25386, N25372, N10801);
nand NAND4 (N25387, N25383, N20491, N8132, N17279);
nand NAND3 (N25388, N25374, N23453, N21047);
nand NAND3 (N25389, N25381, N4648, N20136);
buf BUF1 (N25390, N25388);
xor XOR2 (N25391, N25386, N25294);
not NOT1 (N25392, N25382);
not NOT1 (N25393, N25384);
xor XOR2 (N25394, N25385, N13895);
buf BUF1 (N25395, N25391);
not NOT1 (N25396, N25390);
nor NOR3 (N25397, N25395, N10598, N22235);
buf BUF1 (N25398, N25378);
and AND4 (N25399, N25389, N2095, N7289, N11115);
xor XOR2 (N25400, N25393, N17533);
and AND2 (N25401, N25400, N2389);
not NOT1 (N25402, N25387);
not NOT1 (N25403, N25401);
nand NAND4 (N25404, N25380, N3847, N13160, N3092);
nand NAND4 (N25405, N25392, N12661, N10550, N18116);
or OR3 (N25406, N25402, N219, N3677);
or OR3 (N25407, N25397, N18205, N3296);
not NOT1 (N25408, N25394);
buf BUF1 (N25409, N25407);
buf BUF1 (N25410, N25406);
nand NAND3 (N25411, N25405, N6236, N7622);
nor NOR2 (N25412, N25398, N23035);
not NOT1 (N25413, N25410);
buf BUF1 (N25414, N25412);
and AND3 (N25415, N25414, N18394, N23758);
not NOT1 (N25416, N25403);
not NOT1 (N25417, N25416);
or OR2 (N25418, N25408, N1858);
nor NOR3 (N25419, N25411, N13932, N13505);
nor NOR3 (N25420, N25419, N1231, N8797);
or OR4 (N25421, N25415, N12272, N20595, N13233);
and AND3 (N25422, N25417, N18118, N4894);
nand NAND4 (N25423, N25396, N8615, N23483, N11218);
and AND3 (N25424, N25404, N19312, N575);
buf BUF1 (N25425, N25399);
buf BUF1 (N25426, N25421);
nor NOR3 (N25427, N25423, N23423, N23201);
nor NOR4 (N25428, N25361, N15215, N13995, N13246);
xor XOR2 (N25429, N25424, N12339);
and AND4 (N25430, N25429, N22544, N12388, N4782);
xor XOR2 (N25431, N25409, N17714);
xor XOR2 (N25432, N25426, N19592);
nor NOR2 (N25433, N25413, N17231);
and AND2 (N25434, N25425, N12570);
and AND3 (N25435, N25434, N22730, N5849);
nor NOR2 (N25436, N25433, N22684);
xor XOR2 (N25437, N25422, N24686);
not NOT1 (N25438, N25432);
xor XOR2 (N25439, N25418, N10818);
xor XOR2 (N25440, N25420, N21095);
or OR3 (N25441, N25431, N503, N13520);
xor XOR2 (N25442, N25441, N24243);
nand NAND2 (N25443, N25435, N22926);
or OR2 (N25444, N25442, N1246);
or OR4 (N25445, N25440, N16506, N23602, N1027);
not NOT1 (N25446, N25443);
nor NOR4 (N25447, N25445, N4619, N12285, N7561);
xor XOR2 (N25448, N25428, N10892);
not NOT1 (N25449, N25439);
nand NAND2 (N25450, N25448, N14752);
xor XOR2 (N25451, N25450, N24374);
xor XOR2 (N25452, N25430, N3637);
not NOT1 (N25453, N25444);
or OR4 (N25454, N25438, N3197, N10492, N23050);
buf BUF1 (N25455, N25447);
xor XOR2 (N25456, N25446, N22573);
not NOT1 (N25457, N25451);
buf BUF1 (N25458, N25427);
or OR2 (N25459, N25454, N25335);
buf BUF1 (N25460, N25452);
buf BUF1 (N25461, N25460);
xor XOR2 (N25462, N25437, N230);
xor XOR2 (N25463, N25436, N18364);
nand NAND2 (N25464, N25461, N18401);
nor NOR4 (N25465, N25462, N538, N9663, N12989);
nand NAND2 (N25466, N25458, N3442);
nor NOR2 (N25467, N25463, N8049);
nand NAND2 (N25468, N25449, N5145);
nor NOR4 (N25469, N25456, N12930, N6372, N2474);
nand NAND4 (N25470, N25464, N2943, N15814, N20140);
buf BUF1 (N25471, N25465);
and AND4 (N25472, N25466, N24802, N13575, N3355);
nand NAND4 (N25473, N25470, N3755, N14851, N2299);
or OR2 (N25474, N25473, N13853);
nand NAND3 (N25475, N25472, N7604, N9002);
or OR3 (N25476, N25453, N17042, N23720);
and AND4 (N25477, N25468, N22402, N19505, N14226);
not NOT1 (N25478, N25471);
and AND2 (N25479, N25475, N23603);
xor XOR2 (N25480, N25469, N21988);
nand NAND4 (N25481, N25467, N18072, N22974, N12361);
and AND2 (N25482, N25477, N13190);
nand NAND2 (N25483, N25479, N24116);
and AND3 (N25484, N25478, N18001, N21879);
nand NAND3 (N25485, N25459, N16487, N24924);
xor XOR2 (N25486, N25476, N7368);
buf BUF1 (N25487, N25483);
xor XOR2 (N25488, N25486, N10289);
nor NOR2 (N25489, N25488, N20433);
or OR2 (N25490, N25484, N23739);
nor NOR2 (N25491, N25487, N12742);
not NOT1 (N25492, N25482);
not NOT1 (N25493, N25489);
nand NAND4 (N25494, N25455, N21664, N3621, N1871);
xor XOR2 (N25495, N25491, N17504);
and AND4 (N25496, N25495, N3404, N551, N11092);
nor NOR2 (N25497, N25480, N6032);
and AND3 (N25498, N25474, N6352, N14527);
nand NAND3 (N25499, N25485, N6035, N336);
nor NOR2 (N25500, N25496, N3269);
buf BUF1 (N25501, N25490);
not NOT1 (N25502, N25497);
buf BUF1 (N25503, N25492);
buf BUF1 (N25504, N25498);
or OR2 (N25505, N25500, N8883);
not NOT1 (N25506, N25457);
nand NAND3 (N25507, N25502, N7300, N2307);
nand NAND3 (N25508, N25504, N6383, N6348);
xor XOR2 (N25509, N25499, N568);
and AND4 (N25510, N25505, N5212, N1263, N20079);
xor XOR2 (N25511, N25494, N22280);
xor XOR2 (N25512, N25508, N4053);
xor XOR2 (N25513, N25510, N9901);
nor NOR2 (N25514, N25509, N13582);
buf BUF1 (N25515, N25514);
nand NAND3 (N25516, N25481, N12368, N6328);
or OR4 (N25517, N25512, N23069, N23924, N10200);
nand NAND2 (N25518, N25503, N25034);
buf BUF1 (N25519, N25507);
not NOT1 (N25520, N25516);
or OR3 (N25521, N25519, N8803, N12883);
buf BUF1 (N25522, N25515);
or OR4 (N25523, N25511, N19572, N24502, N15575);
nor NOR3 (N25524, N25520, N22156, N15166);
nor NOR3 (N25525, N25524, N25397, N8212);
or OR4 (N25526, N25513, N11217, N14173, N15407);
not NOT1 (N25527, N25493);
nand NAND3 (N25528, N25501, N7334, N10246);
nor NOR4 (N25529, N25506, N3058, N13962, N18786);
not NOT1 (N25530, N25525);
buf BUF1 (N25531, N25517);
nand NAND4 (N25532, N25518, N5602, N16032, N5650);
xor XOR2 (N25533, N25531, N5085);
nor NOR3 (N25534, N25533, N6174, N20728);
nor NOR2 (N25535, N25523, N18935);
not NOT1 (N25536, N25527);
and AND3 (N25537, N25529, N93, N16186);
and AND4 (N25538, N25526, N4108, N22344, N12406);
and AND3 (N25539, N25530, N20588, N12324);
nor NOR2 (N25540, N25537, N3538);
or OR3 (N25541, N25521, N2012, N1498);
nor NOR3 (N25542, N25539, N17818, N6753);
not NOT1 (N25543, N25534);
nor NOR2 (N25544, N25540, N15908);
nor NOR3 (N25545, N25544, N3669, N14090);
not NOT1 (N25546, N25528);
not NOT1 (N25547, N25536);
not NOT1 (N25548, N25545);
or OR3 (N25549, N25542, N22166, N17685);
buf BUF1 (N25550, N25535);
nor NOR2 (N25551, N25547, N5550);
nor NOR2 (N25552, N25550, N1281);
or OR4 (N25553, N25522, N10950, N6345, N20202);
not NOT1 (N25554, N25538);
nand NAND3 (N25555, N25554, N7276, N13992);
buf BUF1 (N25556, N25549);
not NOT1 (N25557, N25548);
and AND2 (N25558, N25543, N13671);
buf BUF1 (N25559, N25553);
nand NAND4 (N25560, N25556, N16205, N23002, N1680);
and AND2 (N25561, N25555, N4739);
buf BUF1 (N25562, N25561);
nand NAND4 (N25563, N25552, N18046, N8059, N19145);
xor XOR2 (N25564, N25551, N611);
not NOT1 (N25565, N25563);
not NOT1 (N25566, N25546);
and AND4 (N25567, N25560, N15417, N10309, N21641);
buf BUF1 (N25568, N25564);
not NOT1 (N25569, N25566);
not NOT1 (N25570, N25532);
xor XOR2 (N25571, N25558, N24773);
nand NAND4 (N25572, N25571, N1688, N22405, N18705);
not NOT1 (N25573, N25567);
nand NAND2 (N25574, N25573, N15701);
and AND3 (N25575, N25568, N7006, N19022);
nand NAND3 (N25576, N25541, N3142, N25430);
not NOT1 (N25577, N25569);
not NOT1 (N25578, N25574);
nor NOR3 (N25579, N25559, N7806, N6991);
not NOT1 (N25580, N25565);
and AND4 (N25581, N25580, N8176, N21442, N12166);
buf BUF1 (N25582, N25575);
nor NOR3 (N25583, N25572, N4130, N7645);
nand NAND3 (N25584, N25581, N17997, N17816);
nand NAND2 (N25585, N25576, N20651);
nand NAND2 (N25586, N25557, N17313);
nor NOR2 (N25587, N25577, N13061);
xor XOR2 (N25588, N25586, N18470);
nand NAND3 (N25589, N25579, N21894, N24402);
or OR3 (N25590, N25587, N20310, N1152);
xor XOR2 (N25591, N25589, N2416);
not NOT1 (N25592, N25584);
not NOT1 (N25593, N25590);
nand NAND3 (N25594, N25588, N7756, N4250);
and AND4 (N25595, N25593, N17851, N18257, N12219);
nand NAND2 (N25596, N25562, N20511);
xor XOR2 (N25597, N25570, N17939);
and AND4 (N25598, N25596, N9311, N2049, N18120);
buf BUF1 (N25599, N25578);
not NOT1 (N25600, N25582);
and AND3 (N25601, N25599, N21030, N2252);
xor XOR2 (N25602, N25594, N17043);
nand NAND4 (N25603, N25602, N19021, N14819, N20914);
nand NAND3 (N25604, N25597, N4717, N2129);
nand NAND3 (N25605, N25603, N19589, N19362);
not NOT1 (N25606, N25598);
or OR4 (N25607, N25600, N10285, N3519, N589);
and AND2 (N25608, N25601, N15261);
not NOT1 (N25609, N25591);
or OR3 (N25610, N25606, N18915, N10013);
buf BUF1 (N25611, N25583);
not NOT1 (N25612, N25592);
and AND4 (N25613, N25585, N18351, N16966, N23991);
buf BUF1 (N25614, N25608);
or OR4 (N25615, N25609, N18085, N19841, N21805);
buf BUF1 (N25616, N25595);
nand NAND4 (N25617, N25611, N21598, N7907, N16492);
buf BUF1 (N25618, N25612);
xor XOR2 (N25619, N25605, N18632);
and AND2 (N25620, N25604, N14889);
and AND2 (N25621, N25610, N5702);
endmodule