// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21;

output N16006,N16018,N16005,N16019,N16012,N16015,N16020,N16003,N16008,N16021;

and AND3 (N22, N3, N6, N6);
nand NAND3 (N23, N2, N19, N10);
nand NAND3 (N24, N2, N22, N5);
xor XOR2 (N25, N15, N4);
nand NAND4 (N26, N7, N1, N4, N15);
buf BUF1 (N27, N22);
and AND3 (N28, N24, N21, N7);
and AND4 (N29, N9, N21, N7, N23);
buf BUF1 (N30, N26);
xor XOR2 (N31, N23, N26);
nor NOR4 (N32, N10, N20, N7, N8);
buf BUF1 (N33, N23);
and AND4 (N34, N16, N19, N32, N7);
xor XOR2 (N35, N10, N11);
or OR4 (N36, N27, N19, N20, N35);
nor NOR4 (N37, N6, N28, N9, N4);
xor XOR2 (N38, N24, N4);
xor XOR2 (N39, N14, N28);
not NOT1 (N40, N29);
and AND4 (N41, N38, N1, N4, N25);
and AND4 (N42, N23, N32, N37, N24);
and AND2 (N43, N14, N17);
nor NOR4 (N44, N33, N6, N10, N39);
nand NAND4 (N45, N7, N20, N12, N1);
xor XOR2 (N46, N36, N5);
and AND2 (N47, N40, N6);
or OR2 (N48, N31, N3);
not NOT1 (N49, N43);
not NOT1 (N50, N30);
not NOT1 (N51, N50);
nor NOR3 (N52, N51, N43, N38);
buf BUF1 (N53, N48);
or OR4 (N54, N47, N52, N19, N52);
not NOT1 (N55, N27);
nand NAND2 (N56, N54, N16);
not NOT1 (N57, N44);
not NOT1 (N58, N34);
xor XOR2 (N59, N49, N50);
xor XOR2 (N60, N41, N4);
nor NOR3 (N61, N46, N21, N2);
nand NAND3 (N62, N55, N33, N30);
nor NOR4 (N63, N45, N46, N11, N4);
nand NAND4 (N64, N58, N42, N52, N7);
nor NOR4 (N65, N36, N26, N49, N16);
xor XOR2 (N66, N65, N44);
not NOT1 (N67, N66);
xor XOR2 (N68, N62, N39);
nor NOR4 (N69, N57, N51, N4, N10);
buf BUF1 (N70, N59);
not NOT1 (N71, N67);
or OR2 (N72, N61, N27);
xor XOR2 (N73, N56, N12);
not NOT1 (N74, N63);
nor NOR4 (N75, N68, N7, N56, N18);
not NOT1 (N76, N70);
xor XOR2 (N77, N64, N48);
nor NOR3 (N78, N69, N64, N4);
nor NOR4 (N79, N75, N2, N44, N15);
buf BUF1 (N80, N77);
xor XOR2 (N81, N76, N7);
not NOT1 (N82, N53);
xor XOR2 (N83, N72, N60);
and AND4 (N84, N59, N66, N47, N52);
or OR2 (N85, N80, N57);
xor XOR2 (N86, N85, N82);
and AND3 (N87, N7, N83, N24);
nand NAND4 (N88, N4, N7, N31, N84);
buf BUF1 (N89, N28);
nand NAND3 (N90, N79, N4, N42);
xor XOR2 (N91, N74, N44);
or OR2 (N92, N91, N42);
xor XOR2 (N93, N87, N24);
not NOT1 (N94, N86);
xor XOR2 (N95, N93, N26);
and AND4 (N96, N71, N44, N6, N66);
nor NOR4 (N97, N94, N10, N90, N3);
nor NOR4 (N98, N56, N53, N42, N48);
or OR2 (N99, N92, N54);
xor XOR2 (N100, N99, N91);
nor NOR3 (N101, N100, N79, N88);
nand NAND2 (N102, N13, N34);
nor NOR2 (N103, N73, N7);
nand NAND2 (N104, N81, N74);
nand NAND3 (N105, N104, N58, N6);
not NOT1 (N106, N96);
or OR2 (N107, N106, N77);
xor XOR2 (N108, N103, N42);
nor NOR3 (N109, N101, N54, N33);
buf BUF1 (N110, N107);
xor XOR2 (N111, N102, N33);
or OR2 (N112, N111, N3);
nand NAND3 (N113, N98, N93, N23);
or OR4 (N114, N108, N104, N99, N107);
buf BUF1 (N115, N105);
nor NOR2 (N116, N89, N24);
buf BUF1 (N117, N116);
not NOT1 (N118, N110);
or OR2 (N119, N78, N20);
and AND4 (N120, N113, N103, N105, N74);
nand NAND3 (N121, N118, N113, N61);
buf BUF1 (N122, N97);
nand NAND4 (N123, N109, N83, N30, N77);
buf BUF1 (N124, N115);
xor XOR2 (N125, N112, N114);
buf BUF1 (N126, N80);
xor XOR2 (N127, N117, N72);
nand NAND4 (N128, N127, N85, N78, N83);
and AND2 (N129, N120, N88);
not NOT1 (N130, N129);
nand NAND3 (N131, N123, N11, N32);
nand NAND4 (N132, N128, N42, N8, N95);
buf BUF1 (N133, N94);
not NOT1 (N134, N132);
not NOT1 (N135, N126);
and AND4 (N136, N134, N53, N64, N17);
xor XOR2 (N137, N133, N15);
nor NOR2 (N138, N122, N14);
nand NAND4 (N139, N135, N138, N35, N14);
buf BUF1 (N140, N112);
nand NAND2 (N141, N124, N51);
nand NAND2 (N142, N119, N44);
nand NAND2 (N143, N131, N51);
or OR2 (N144, N125, N26);
or OR2 (N145, N141, N131);
xor XOR2 (N146, N140, N67);
or OR3 (N147, N143, N50, N143);
xor XOR2 (N148, N142, N102);
buf BUF1 (N149, N136);
or OR2 (N150, N149, N90);
not NOT1 (N151, N139);
xor XOR2 (N152, N151, N60);
nand NAND3 (N153, N152, N66, N88);
nand NAND4 (N154, N145, N52, N93, N121);
nor NOR2 (N155, N36, N28);
not NOT1 (N156, N155);
xor XOR2 (N157, N146, N29);
xor XOR2 (N158, N148, N131);
and AND4 (N159, N157, N7, N54, N24);
and AND2 (N160, N159, N143);
and AND3 (N161, N160, N106, N80);
nor NOR3 (N162, N158, N79, N86);
not NOT1 (N163, N153);
not NOT1 (N164, N163);
nor NOR3 (N165, N164, N93, N120);
nor NOR3 (N166, N162, N5, N107);
not NOT1 (N167, N165);
nor NOR4 (N168, N144, N117, N153, N58);
buf BUF1 (N169, N168);
not NOT1 (N170, N130);
nor NOR2 (N171, N154, N62);
and AND4 (N172, N166, N74, N69, N157);
or OR4 (N173, N137, N62, N39, N140);
and AND2 (N174, N167, N18);
and AND3 (N175, N150, N82, N122);
nand NAND3 (N176, N161, N149, N14);
buf BUF1 (N177, N173);
or OR4 (N178, N170, N1, N90, N98);
not NOT1 (N179, N169);
nor NOR3 (N180, N175, N103, N134);
nand NAND4 (N181, N177, N111, N18, N51);
xor XOR2 (N182, N147, N94);
or OR4 (N183, N178, N160, N78, N6);
or OR3 (N184, N181, N106, N143);
nor NOR3 (N185, N176, N55, N163);
buf BUF1 (N186, N182);
and AND4 (N187, N179, N10, N137, N38);
nor NOR3 (N188, N183, N78, N179);
nor NOR3 (N189, N184, N159, N37);
not NOT1 (N190, N186);
nand NAND4 (N191, N174, N97, N190, N6);
xor XOR2 (N192, N121, N190);
buf BUF1 (N193, N172);
not NOT1 (N194, N180);
nand NAND4 (N195, N185, N46, N179, N115);
xor XOR2 (N196, N171, N2);
or OR3 (N197, N191, N80, N23);
nor NOR3 (N198, N156, N4, N106);
or OR3 (N199, N197, N10, N7);
or OR4 (N200, N195, N97, N91, N70);
nor NOR4 (N201, N196, N143, N102, N189);
nand NAND2 (N202, N178, N155);
xor XOR2 (N203, N200, N195);
nand NAND2 (N204, N193, N112);
and AND4 (N205, N202, N125, N155, N155);
or OR2 (N206, N199, N173);
nand NAND4 (N207, N188, N105, N74, N193);
xor XOR2 (N208, N205, N145);
nand NAND3 (N209, N208, N66, N115);
nand NAND3 (N210, N198, N200, N123);
not NOT1 (N211, N203);
or OR3 (N212, N209, N77, N82);
or OR4 (N213, N194, N74, N46, N109);
xor XOR2 (N214, N192, N45);
nor NOR2 (N215, N210, N78);
nand NAND4 (N216, N212, N19, N65, N164);
buf BUF1 (N217, N213);
nor NOR4 (N218, N214, N31, N121, N192);
nand NAND2 (N219, N216, N109);
and AND2 (N220, N201, N153);
or OR2 (N221, N215, N179);
and AND2 (N222, N221, N187);
not NOT1 (N223, N156);
xor XOR2 (N224, N207, N101);
nor NOR2 (N225, N211, N118);
xor XOR2 (N226, N204, N112);
not NOT1 (N227, N217);
nand NAND3 (N228, N218, N146, N23);
xor XOR2 (N229, N220, N106);
nor NOR3 (N230, N206, N104, N136);
buf BUF1 (N231, N222);
buf BUF1 (N232, N219);
nor NOR4 (N233, N228, N209, N147, N180);
or OR2 (N234, N224, N74);
buf BUF1 (N235, N223);
buf BUF1 (N236, N235);
or OR2 (N237, N227, N161);
nor NOR3 (N238, N229, N222, N7);
nor NOR2 (N239, N225, N105);
not NOT1 (N240, N232);
buf BUF1 (N241, N237);
nor NOR2 (N242, N240, N7);
not NOT1 (N243, N242);
not NOT1 (N244, N239);
and AND4 (N245, N236, N45, N90, N71);
nand NAND2 (N246, N230, N65);
xor XOR2 (N247, N234, N24);
and AND4 (N248, N246, N54, N183, N84);
or OR4 (N249, N233, N72, N181, N216);
nor NOR4 (N250, N226, N180, N96, N138);
buf BUF1 (N251, N231);
or OR4 (N252, N251, N37, N72, N213);
nand NAND3 (N253, N244, N171, N119);
nor NOR3 (N254, N249, N177, N64);
nand NAND4 (N255, N252, N72, N218, N140);
buf BUF1 (N256, N250);
xor XOR2 (N257, N255, N58);
not NOT1 (N258, N247);
nor NOR2 (N259, N248, N201);
xor XOR2 (N260, N243, N136);
xor XOR2 (N261, N253, N128);
nor NOR4 (N262, N254, N97, N89, N48);
nand NAND2 (N263, N256, N190);
nand NAND4 (N264, N245, N186, N211, N183);
nand NAND4 (N265, N238, N52, N119, N27);
xor XOR2 (N266, N265, N196);
nand NAND2 (N267, N241, N70);
nand NAND4 (N268, N258, N85, N37, N4);
nor NOR2 (N269, N260, N247);
xor XOR2 (N270, N269, N217);
xor XOR2 (N271, N266, N80);
not NOT1 (N272, N263);
or OR4 (N273, N262, N51, N224, N188);
buf BUF1 (N274, N273);
nand NAND3 (N275, N272, N198, N47);
nand NAND4 (N276, N270, N198, N40, N27);
and AND2 (N277, N268, N8);
not NOT1 (N278, N267);
or OR4 (N279, N257, N239, N110, N43);
nand NAND4 (N280, N275, N66, N5, N117);
or OR2 (N281, N279, N72);
or OR3 (N282, N276, N136, N194);
buf BUF1 (N283, N271);
nor NOR4 (N284, N261, N16, N67, N99);
nor NOR2 (N285, N283, N13);
and AND4 (N286, N277, N9, N60, N191);
nand NAND2 (N287, N282, N207);
xor XOR2 (N288, N280, N257);
not NOT1 (N289, N285);
nor NOR3 (N290, N286, N98, N162);
or OR4 (N291, N259, N229, N250, N50);
not NOT1 (N292, N264);
or OR2 (N293, N290, N162);
nand NAND2 (N294, N281, N104);
buf BUF1 (N295, N288);
buf BUF1 (N296, N293);
nor NOR3 (N297, N284, N130, N81);
and AND3 (N298, N297, N102, N235);
nand NAND4 (N299, N278, N7, N251, N199);
not NOT1 (N300, N298);
buf BUF1 (N301, N296);
buf BUF1 (N302, N292);
xor XOR2 (N303, N302, N250);
or OR2 (N304, N299, N228);
nand NAND2 (N305, N300, N149);
nand NAND3 (N306, N287, N95, N157);
nand NAND2 (N307, N274, N95);
nand NAND4 (N308, N306, N299, N30, N22);
and AND4 (N309, N291, N50, N214, N84);
nor NOR2 (N310, N301, N10);
and AND3 (N311, N303, N141, N149);
not NOT1 (N312, N310);
or OR2 (N313, N311, N211);
buf BUF1 (N314, N305);
buf BUF1 (N315, N313);
not NOT1 (N316, N309);
buf BUF1 (N317, N315);
buf BUF1 (N318, N312);
or OR4 (N319, N294, N241, N312, N71);
nor NOR4 (N320, N304, N126, N60, N38);
or OR3 (N321, N314, N237, N178);
and AND3 (N322, N318, N296, N69);
nand NAND3 (N323, N307, N65, N175);
not NOT1 (N324, N316);
and AND2 (N325, N324, N24);
nor NOR4 (N326, N325, N285, N196, N94);
buf BUF1 (N327, N295);
nor NOR3 (N328, N321, N289, N78);
or OR2 (N329, N259, N274);
or OR3 (N330, N308, N130, N238);
buf BUF1 (N331, N329);
xor XOR2 (N332, N320, N58);
buf BUF1 (N333, N331);
xor XOR2 (N334, N332, N320);
nor NOR2 (N335, N323, N82);
or OR4 (N336, N326, N112, N64, N198);
buf BUF1 (N337, N328);
nor NOR3 (N338, N336, N200, N91);
buf BUF1 (N339, N338);
buf BUF1 (N340, N330);
xor XOR2 (N341, N317, N81);
xor XOR2 (N342, N340, N101);
nor NOR3 (N343, N337, N88, N88);
nand NAND4 (N344, N327, N188, N80, N124);
nor NOR4 (N345, N322, N221, N178, N48);
or OR4 (N346, N345, N212, N210, N305);
not NOT1 (N347, N335);
and AND4 (N348, N343, N235, N97, N200);
nand NAND2 (N349, N346, N334);
not NOT1 (N350, N169);
nor NOR2 (N351, N344, N328);
or OR2 (N352, N348, N224);
nand NAND3 (N353, N350, N73, N314);
or OR4 (N354, N352, N116, N155, N258);
xor XOR2 (N355, N342, N215);
nand NAND4 (N356, N349, N341, N261, N188);
or OR3 (N357, N63, N10, N330);
nand NAND2 (N358, N354, N166);
buf BUF1 (N359, N357);
and AND3 (N360, N358, N71, N358);
not NOT1 (N361, N360);
and AND2 (N362, N359, N254);
xor XOR2 (N363, N355, N305);
and AND2 (N364, N356, N99);
and AND3 (N365, N333, N83, N181);
or OR2 (N366, N362, N207);
and AND3 (N367, N364, N43, N353);
xor XOR2 (N368, N363, N70);
and AND4 (N369, N296, N13, N194, N292);
and AND3 (N370, N347, N367, N37);
not NOT1 (N371, N101);
buf BUF1 (N372, N370);
xor XOR2 (N373, N361, N211);
or OR3 (N374, N366, N341, N311);
and AND3 (N375, N365, N39, N141);
or OR4 (N376, N368, N220, N283, N77);
nor NOR3 (N377, N373, N157, N368);
nand NAND3 (N378, N377, N14, N90);
not NOT1 (N379, N372);
xor XOR2 (N380, N379, N178);
nor NOR3 (N381, N380, N355, N284);
not NOT1 (N382, N339);
or OR4 (N383, N382, N103, N245, N176);
nand NAND2 (N384, N351, N49);
buf BUF1 (N385, N319);
xor XOR2 (N386, N384, N267);
buf BUF1 (N387, N374);
and AND3 (N388, N387, N304, N177);
xor XOR2 (N389, N388, N355);
not NOT1 (N390, N371);
and AND4 (N391, N378, N242, N64, N43);
xor XOR2 (N392, N383, N178);
xor XOR2 (N393, N392, N275);
or OR2 (N394, N390, N2);
nand NAND2 (N395, N375, N124);
buf BUF1 (N396, N391);
nand NAND3 (N397, N369, N262, N229);
nand NAND4 (N398, N385, N348, N79, N256);
or OR2 (N399, N393, N114);
buf BUF1 (N400, N397);
not NOT1 (N401, N395);
buf BUF1 (N402, N376);
and AND4 (N403, N399, N133, N393, N271);
nand NAND3 (N404, N400, N168, N64);
xor XOR2 (N405, N402, N235);
or OR2 (N406, N404, N228);
nand NAND4 (N407, N401, N185, N6, N406);
buf BUF1 (N408, N59);
nand NAND4 (N409, N394, N372, N108, N328);
and AND2 (N410, N409, N309);
xor XOR2 (N411, N381, N396);
buf BUF1 (N412, N32);
nor NOR2 (N413, N405, N359);
xor XOR2 (N414, N386, N184);
nor NOR2 (N415, N408, N279);
buf BUF1 (N416, N415);
nand NAND2 (N417, N410, N323);
nor NOR4 (N418, N414, N22, N9, N409);
nor NOR4 (N419, N412, N196, N258, N241);
nor NOR2 (N420, N403, N203);
or OR3 (N421, N407, N287, N37);
or OR3 (N422, N389, N294, N292);
not NOT1 (N423, N417);
nand NAND2 (N424, N413, N307);
and AND4 (N425, N411, N361, N394, N145);
nor NOR3 (N426, N418, N77, N141);
and AND3 (N427, N425, N290, N204);
nand NAND3 (N428, N423, N234, N328);
nor NOR3 (N429, N427, N295, N42);
xor XOR2 (N430, N416, N117);
xor XOR2 (N431, N421, N426);
buf BUF1 (N432, N153);
xor XOR2 (N433, N428, N29);
or OR2 (N434, N424, N102);
buf BUF1 (N435, N420);
or OR4 (N436, N431, N238, N204, N251);
nor NOR3 (N437, N432, N99, N341);
or OR4 (N438, N434, N417, N230, N310);
nor NOR4 (N439, N433, N268, N397, N173);
buf BUF1 (N440, N437);
buf BUF1 (N441, N436);
and AND2 (N442, N422, N246);
and AND3 (N443, N419, N374, N392);
buf BUF1 (N444, N441);
or OR4 (N445, N444, N23, N78, N360);
and AND3 (N446, N438, N416, N4);
not NOT1 (N447, N442);
xor XOR2 (N448, N446, N109);
xor XOR2 (N449, N445, N215);
nor NOR3 (N450, N439, N403, N92);
not NOT1 (N451, N448);
xor XOR2 (N452, N440, N435);
xor XOR2 (N453, N335, N17);
buf BUF1 (N454, N429);
nor NOR4 (N455, N449, N389, N91, N343);
nand NAND4 (N456, N430, N267, N144, N129);
nand NAND4 (N457, N447, N366, N77, N122);
not NOT1 (N458, N452);
xor XOR2 (N459, N455, N27);
xor XOR2 (N460, N456, N392);
not NOT1 (N461, N450);
buf BUF1 (N462, N461);
and AND4 (N463, N398, N128, N375, N124);
not NOT1 (N464, N460);
and AND2 (N465, N451, N114);
buf BUF1 (N466, N464);
and AND3 (N467, N465, N408, N164);
nor NOR2 (N468, N457, N401);
buf BUF1 (N469, N463);
not NOT1 (N470, N467);
buf BUF1 (N471, N458);
nand NAND2 (N472, N443, N164);
and AND4 (N473, N453, N431, N422, N355);
buf BUF1 (N474, N459);
nor NOR4 (N475, N471, N89, N33, N301);
or OR3 (N476, N475, N245, N381);
xor XOR2 (N477, N466, N370);
and AND2 (N478, N473, N105);
xor XOR2 (N479, N462, N304);
not NOT1 (N480, N454);
xor XOR2 (N481, N480, N295);
nor NOR2 (N482, N479, N50);
and AND3 (N483, N472, N265, N4);
nand NAND4 (N484, N474, N330, N41, N12);
nand NAND2 (N485, N481, N314);
nor NOR4 (N486, N485, N186, N150, N419);
nand NAND3 (N487, N469, N311, N468);
not NOT1 (N488, N121);
buf BUF1 (N489, N476);
buf BUF1 (N490, N482);
and AND4 (N491, N488, N326, N246, N326);
nand NAND2 (N492, N490, N442);
or OR2 (N493, N470, N250);
and AND2 (N494, N478, N181);
buf BUF1 (N495, N494);
and AND2 (N496, N489, N429);
and AND4 (N497, N492, N256, N65, N149);
not NOT1 (N498, N487);
buf BUF1 (N499, N477);
xor XOR2 (N500, N483, N441);
and AND2 (N501, N493, N374);
buf BUF1 (N502, N499);
xor XOR2 (N503, N498, N315);
or OR3 (N504, N486, N158, N72);
nor NOR2 (N505, N496, N396);
not NOT1 (N506, N497);
and AND4 (N507, N506, N289, N466, N476);
xor XOR2 (N508, N503, N366);
not NOT1 (N509, N484);
xor XOR2 (N510, N504, N39);
nor NOR3 (N511, N507, N378, N297);
and AND2 (N512, N495, N57);
buf BUF1 (N513, N509);
or OR2 (N514, N510, N225);
nor NOR2 (N515, N508, N7);
xor XOR2 (N516, N514, N287);
or OR2 (N517, N491, N121);
nand NAND4 (N518, N501, N79, N388, N294);
buf BUF1 (N519, N500);
or OR3 (N520, N516, N392, N192);
xor XOR2 (N521, N513, N402);
nand NAND3 (N522, N520, N195, N58);
and AND2 (N523, N511, N517);
or OR4 (N524, N346, N313, N16, N20);
not NOT1 (N525, N522);
buf BUF1 (N526, N523);
and AND4 (N527, N524, N408, N39, N427);
buf BUF1 (N528, N502);
not NOT1 (N529, N526);
or OR4 (N530, N527, N295, N1, N400);
buf BUF1 (N531, N518);
xor XOR2 (N532, N531, N406);
xor XOR2 (N533, N515, N122);
or OR4 (N534, N533, N429, N171, N449);
xor XOR2 (N535, N505, N57);
and AND4 (N536, N530, N265, N59, N65);
and AND2 (N537, N525, N376);
buf BUF1 (N538, N529);
nand NAND3 (N539, N535, N494, N257);
nand NAND2 (N540, N536, N293);
buf BUF1 (N541, N540);
nor NOR4 (N542, N519, N96, N530, N404);
and AND4 (N543, N541, N237, N105, N132);
xor XOR2 (N544, N512, N526);
and AND4 (N545, N542, N418, N424, N136);
nand NAND2 (N546, N534, N377);
not NOT1 (N547, N543);
not NOT1 (N548, N538);
or OR2 (N549, N548, N305);
or OR2 (N550, N546, N494);
nand NAND2 (N551, N521, N321);
or OR4 (N552, N550, N196, N139, N147);
xor XOR2 (N553, N552, N190);
not NOT1 (N554, N547);
nand NAND2 (N555, N551, N215);
and AND4 (N556, N537, N252, N411, N329);
or OR4 (N557, N544, N51, N99, N124);
buf BUF1 (N558, N557);
or OR2 (N559, N528, N545);
or OR3 (N560, N126, N111, N351);
nor NOR4 (N561, N555, N384, N245, N399);
not NOT1 (N562, N539);
nor NOR3 (N563, N556, N234, N404);
not NOT1 (N564, N553);
nand NAND4 (N565, N532, N9, N61, N320);
or OR3 (N566, N558, N44, N144);
or OR2 (N567, N562, N168);
or OR4 (N568, N567, N499, N263, N411);
and AND4 (N569, N568, N198, N203, N299);
xor XOR2 (N570, N549, N191);
nand NAND3 (N571, N565, N38, N434);
nand NAND4 (N572, N571, N65, N393, N276);
not NOT1 (N573, N566);
buf BUF1 (N574, N563);
xor XOR2 (N575, N573, N409);
xor XOR2 (N576, N575, N34);
nand NAND2 (N577, N576, N329);
nand NAND2 (N578, N560, N159);
nand NAND2 (N579, N564, N507);
nand NAND2 (N580, N561, N420);
not NOT1 (N581, N570);
nand NAND3 (N582, N569, N361, N38);
not NOT1 (N583, N574);
xor XOR2 (N584, N572, N127);
not NOT1 (N585, N584);
nand NAND3 (N586, N579, N19, N159);
buf BUF1 (N587, N586);
xor XOR2 (N588, N585, N217);
nand NAND4 (N589, N577, N17, N70, N251);
nand NAND2 (N590, N587, N81);
and AND3 (N591, N580, N235, N332);
buf BUF1 (N592, N554);
nor NOR2 (N593, N583, N576);
buf BUF1 (N594, N559);
buf BUF1 (N595, N589);
nor NOR2 (N596, N594, N97);
nand NAND3 (N597, N582, N533, N559);
not NOT1 (N598, N578);
or OR2 (N599, N581, N334);
not NOT1 (N600, N597);
not NOT1 (N601, N592);
xor XOR2 (N602, N591, N455);
or OR2 (N603, N590, N252);
and AND3 (N604, N595, N365, N438);
xor XOR2 (N605, N588, N34);
not NOT1 (N606, N604);
xor XOR2 (N607, N605, N523);
nand NAND4 (N608, N598, N169, N128, N173);
nand NAND2 (N609, N596, N148);
nand NAND2 (N610, N601, N50);
buf BUF1 (N611, N600);
not NOT1 (N612, N611);
not NOT1 (N613, N610);
or OR3 (N614, N606, N386, N535);
buf BUF1 (N615, N607);
or OR3 (N616, N613, N204, N582);
not NOT1 (N617, N609);
not NOT1 (N618, N599);
and AND4 (N619, N618, N254, N82, N518);
xor XOR2 (N620, N593, N123);
not NOT1 (N621, N615);
xor XOR2 (N622, N621, N202);
nand NAND3 (N623, N612, N602, N93);
and AND4 (N624, N474, N88, N296, N235);
not NOT1 (N625, N603);
not NOT1 (N626, N622);
or OR4 (N627, N617, N341, N198, N575);
nor NOR4 (N628, N614, N591, N423, N476);
xor XOR2 (N629, N620, N345);
buf BUF1 (N630, N625);
nand NAND2 (N631, N616, N523);
nor NOR3 (N632, N630, N85, N499);
nor NOR3 (N633, N624, N525, N455);
buf BUF1 (N634, N608);
nand NAND3 (N635, N626, N97, N197);
nand NAND3 (N636, N619, N631, N18);
not NOT1 (N637, N341);
and AND2 (N638, N632, N135);
and AND2 (N639, N629, N514);
and AND2 (N640, N633, N159);
nand NAND2 (N641, N637, N12);
buf BUF1 (N642, N641);
nand NAND4 (N643, N623, N226, N277, N426);
not NOT1 (N644, N638);
nand NAND4 (N645, N628, N388, N478, N166);
not NOT1 (N646, N635);
or OR4 (N647, N627, N74, N56, N525);
nor NOR4 (N648, N639, N91, N474, N524);
and AND2 (N649, N644, N373);
or OR4 (N650, N636, N504, N641, N266);
not NOT1 (N651, N649);
nand NAND3 (N652, N634, N91, N315);
nand NAND2 (N653, N650, N485);
buf BUF1 (N654, N646);
xor XOR2 (N655, N643, N384);
buf BUF1 (N656, N654);
buf BUF1 (N657, N645);
xor XOR2 (N658, N653, N489);
not NOT1 (N659, N647);
and AND3 (N660, N655, N215, N255);
and AND3 (N661, N640, N112, N48);
xor XOR2 (N662, N658, N9);
not NOT1 (N663, N661);
not NOT1 (N664, N656);
and AND2 (N665, N657, N70);
buf BUF1 (N666, N651);
nand NAND3 (N667, N648, N155, N151);
nand NAND2 (N668, N666, N635);
or OR4 (N669, N664, N189, N429, N239);
and AND3 (N670, N659, N72, N623);
buf BUF1 (N671, N652);
buf BUF1 (N672, N668);
nand NAND3 (N673, N672, N535, N368);
nand NAND4 (N674, N660, N151, N359, N32);
xor XOR2 (N675, N663, N231);
or OR2 (N676, N674, N481);
buf BUF1 (N677, N673);
or OR2 (N678, N675, N155);
not NOT1 (N679, N670);
nand NAND4 (N680, N662, N50, N402, N292);
buf BUF1 (N681, N671);
nand NAND3 (N682, N665, N147, N281);
nand NAND2 (N683, N642, N668);
nand NAND4 (N684, N678, N344, N412, N95);
not NOT1 (N685, N679);
not NOT1 (N686, N682);
buf BUF1 (N687, N681);
nand NAND4 (N688, N669, N382, N89, N545);
not NOT1 (N689, N683);
xor XOR2 (N690, N687, N559);
and AND3 (N691, N686, N53, N344);
or OR2 (N692, N690, N416);
buf BUF1 (N693, N691);
and AND4 (N694, N677, N292, N27, N218);
not NOT1 (N695, N694);
nand NAND4 (N696, N693, N397, N162, N308);
or OR3 (N697, N688, N689, N633);
nand NAND3 (N698, N302, N132, N396);
nand NAND2 (N699, N676, N320);
xor XOR2 (N700, N695, N429);
and AND4 (N701, N667, N42, N452, N46);
nor NOR2 (N702, N698, N659);
nor NOR2 (N703, N680, N147);
buf BUF1 (N704, N684);
and AND4 (N705, N704, N677, N699, N8);
nand NAND2 (N706, N400, N494);
and AND2 (N707, N700, N555);
or OR3 (N708, N696, N83, N368);
and AND3 (N709, N697, N301, N448);
not NOT1 (N710, N709);
nand NAND4 (N711, N703, N585, N337, N200);
not NOT1 (N712, N708);
nor NOR3 (N713, N711, N145, N633);
nor NOR4 (N714, N692, N202, N199, N279);
nand NAND4 (N715, N705, N35, N175, N165);
nor NOR3 (N716, N706, N331, N549);
buf BUF1 (N717, N702);
buf BUF1 (N718, N717);
xor XOR2 (N719, N715, N39);
xor XOR2 (N720, N713, N483);
xor XOR2 (N721, N712, N575);
and AND3 (N722, N714, N409, N280);
xor XOR2 (N723, N707, N667);
and AND2 (N724, N710, N647);
nand NAND2 (N725, N701, N390);
nand NAND2 (N726, N725, N292);
and AND2 (N727, N719, N571);
and AND2 (N728, N721, N48);
or OR4 (N729, N727, N538, N234, N391);
nand NAND4 (N730, N726, N167, N81, N516);
or OR4 (N731, N685, N237, N512, N214);
nor NOR3 (N732, N720, N638, N132);
nor NOR4 (N733, N723, N611, N43, N273);
or OR4 (N734, N716, N492, N630, N199);
not NOT1 (N735, N724);
or OR3 (N736, N734, N72, N584);
buf BUF1 (N737, N735);
and AND4 (N738, N729, N176, N230, N74);
buf BUF1 (N739, N737);
or OR3 (N740, N739, N340, N405);
buf BUF1 (N741, N731);
or OR2 (N742, N741, N131);
or OR4 (N743, N738, N475, N725, N29);
buf BUF1 (N744, N736);
or OR2 (N745, N730, N53);
or OR2 (N746, N733, N211);
or OR4 (N747, N743, N580, N532, N617);
xor XOR2 (N748, N718, N746);
buf BUF1 (N749, N118);
or OR4 (N750, N728, N528, N693, N380);
nor NOR3 (N751, N722, N191, N719);
or OR2 (N752, N747, N551);
xor XOR2 (N753, N751, N432);
and AND2 (N754, N742, N329);
nor NOR4 (N755, N750, N734, N161, N260);
xor XOR2 (N756, N749, N163);
nand NAND4 (N757, N732, N246, N9, N215);
or OR4 (N758, N744, N461, N703, N291);
or OR4 (N759, N753, N25, N497, N495);
not NOT1 (N760, N740);
nand NAND2 (N761, N754, N649);
or OR3 (N762, N752, N185, N106);
not NOT1 (N763, N760);
or OR3 (N764, N763, N376, N205);
nand NAND3 (N765, N758, N740, N360);
nand NAND3 (N766, N761, N296, N445);
xor XOR2 (N767, N762, N491);
or OR2 (N768, N755, N261);
or OR4 (N769, N764, N434, N9, N706);
xor XOR2 (N770, N768, N650);
and AND3 (N771, N766, N258, N54);
nor NOR4 (N772, N765, N596, N72, N616);
buf BUF1 (N773, N756);
and AND2 (N774, N748, N36);
and AND4 (N775, N767, N303, N90, N444);
and AND3 (N776, N774, N472, N289);
nor NOR2 (N777, N757, N280);
not NOT1 (N778, N773);
nand NAND3 (N779, N777, N310, N149);
xor XOR2 (N780, N771, N719);
nor NOR4 (N781, N780, N674, N757, N298);
nand NAND4 (N782, N769, N720, N138, N754);
or OR3 (N783, N778, N239, N745);
nand NAND3 (N784, N36, N290, N780);
nor NOR3 (N785, N781, N736, N321);
and AND3 (N786, N775, N228, N362);
and AND4 (N787, N770, N735, N760, N635);
or OR4 (N788, N786, N332, N173, N217);
nor NOR2 (N789, N785, N720);
and AND3 (N790, N779, N624, N241);
or OR3 (N791, N783, N91, N766);
not NOT1 (N792, N791);
not NOT1 (N793, N784);
nand NAND2 (N794, N792, N596);
nor NOR4 (N795, N793, N417, N447, N294);
nor NOR3 (N796, N759, N479, N584);
nand NAND3 (N797, N790, N435, N312);
nor NOR4 (N798, N772, N67, N187, N4);
not NOT1 (N799, N794);
or OR4 (N800, N776, N650, N607, N116);
xor XOR2 (N801, N797, N554);
or OR4 (N802, N787, N440, N295, N739);
not NOT1 (N803, N802);
nor NOR2 (N804, N800, N799);
nand NAND4 (N805, N546, N237, N482, N412);
buf BUF1 (N806, N796);
nand NAND4 (N807, N788, N9, N509, N126);
not NOT1 (N808, N806);
nand NAND2 (N809, N798, N351);
nand NAND4 (N810, N795, N607, N647, N409);
nand NAND4 (N811, N803, N795, N575, N16);
xor XOR2 (N812, N810, N22);
or OR2 (N813, N801, N415);
or OR4 (N814, N805, N81, N607, N577);
buf BUF1 (N815, N807);
or OR3 (N816, N782, N315, N438);
nand NAND2 (N817, N789, N267);
buf BUF1 (N818, N813);
nand NAND2 (N819, N814, N721);
nand NAND2 (N820, N804, N553);
or OR4 (N821, N808, N709, N602, N505);
nor NOR4 (N822, N815, N50, N452, N399);
not NOT1 (N823, N816);
not NOT1 (N824, N823);
or OR4 (N825, N821, N519, N536, N371);
nand NAND3 (N826, N812, N419, N113);
nand NAND4 (N827, N811, N336, N19, N311);
and AND2 (N828, N820, N109);
nor NOR4 (N829, N809, N60, N602, N523);
nand NAND4 (N830, N826, N220, N321, N103);
not NOT1 (N831, N827);
nand NAND4 (N832, N819, N670, N246, N405);
nor NOR2 (N833, N831, N325);
buf BUF1 (N834, N829);
buf BUF1 (N835, N833);
and AND2 (N836, N832, N48);
nor NOR4 (N837, N822, N827, N625, N109);
or OR2 (N838, N835, N18);
not NOT1 (N839, N828);
xor XOR2 (N840, N834, N255);
buf BUF1 (N841, N825);
nor NOR3 (N842, N836, N738, N501);
nand NAND4 (N843, N830, N651, N452, N820);
buf BUF1 (N844, N818);
xor XOR2 (N845, N843, N393);
and AND3 (N846, N837, N138, N832);
nor NOR4 (N847, N824, N520, N806, N30);
nor NOR3 (N848, N847, N192, N67);
xor XOR2 (N849, N844, N564);
nor NOR4 (N850, N845, N230, N590, N288);
nor NOR4 (N851, N840, N376, N355, N72);
nor NOR2 (N852, N841, N616);
and AND2 (N853, N817, N135);
and AND2 (N854, N838, N461);
xor XOR2 (N855, N848, N220);
and AND3 (N856, N851, N448, N472);
nand NAND2 (N857, N849, N117);
not NOT1 (N858, N852);
nand NAND2 (N859, N854, N383);
nor NOR2 (N860, N855, N810);
nor NOR4 (N861, N857, N236, N473, N371);
buf BUF1 (N862, N846);
or OR4 (N863, N862, N639, N592, N754);
nor NOR4 (N864, N863, N84, N769, N121);
or OR3 (N865, N860, N279, N597);
or OR2 (N866, N859, N854);
or OR3 (N867, N864, N61, N823);
nand NAND3 (N868, N856, N524, N691);
nor NOR2 (N869, N850, N333);
not NOT1 (N870, N869);
nand NAND2 (N871, N870, N800);
or OR2 (N872, N871, N725);
nand NAND3 (N873, N867, N410, N782);
xor XOR2 (N874, N861, N557);
or OR3 (N875, N858, N479, N82);
nand NAND4 (N876, N868, N62, N717, N586);
nor NOR2 (N877, N839, N646);
nand NAND3 (N878, N877, N32, N741);
xor XOR2 (N879, N853, N278);
buf BUF1 (N880, N873);
xor XOR2 (N881, N879, N557);
not NOT1 (N882, N875);
buf BUF1 (N883, N842);
or OR3 (N884, N865, N835, N757);
not NOT1 (N885, N872);
nor NOR2 (N886, N882, N746);
nand NAND2 (N887, N874, N262);
nand NAND2 (N888, N876, N120);
or OR3 (N889, N888, N30, N532);
nand NAND2 (N890, N889, N528);
buf BUF1 (N891, N885);
buf BUF1 (N892, N890);
nand NAND3 (N893, N892, N229, N672);
xor XOR2 (N894, N884, N229);
nor NOR3 (N895, N886, N557, N859);
nor NOR4 (N896, N880, N50, N760, N655);
and AND4 (N897, N893, N869, N506, N895);
not NOT1 (N898, N679);
buf BUF1 (N899, N887);
not NOT1 (N900, N866);
buf BUF1 (N901, N891);
xor XOR2 (N902, N898, N509);
not NOT1 (N903, N900);
xor XOR2 (N904, N896, N688);
and AND2 (N905, N897, N126);
nand NAND3 (N906, N894, N392, N862);
xor XOR2 (N907, N903, N346);
and AND2 (N908, N906, N769);
nand NAND3 (N909, N883, N79, N858);
nand NAND2 (N910, N904, N439);
xor XOR2 (N911, N901, N1);
xor XOR2 (N912, N905, N348);
buf BUF1 (N913, N909);
not NOT1 (N914, N913);
xor XOR2 (N915, N910, N311);
not NOT1 (N916, N908);
xor XOR2 (N917, N916, N730);
buf BUF1 (N918, N902);
buf BUF1 (N919, N911);
xor XOR2 (N920, N881, N121);
buf BUF1 (N921, N918);
not NOT1 (N922, N920);
nor NOR3 (N923, N878, N820, N144);
xor XOR2 (N924, N899, N548);
nor NOR4 (N925, N914, N626, N852, N325);
buf BUF1 (N926, N924);
nor NOR3 (N927, N922, N208, N99);
or OR3 (N928, N921, N892, N631);
nor NOR4 (N929, N928, N39, N326, N492);
buf BUF1 (N930, N917);
nor NOR2 (N931, N912, N141);
not NOT1 (N932, N926);
xor XOR2 (N933, N929, N213);
or OR2 (N934, N933, N717);
or OR2 (N935, N927, N598);
xor XOR2 (N936, N931, N832);
and AND3 (N937, N936, N922, N455);
nor NOR2 (N938, N923, N90);
not NOT1 (N939, N938);
not NOT1 (N940, N907);
nor NOR4 (N941, N915, N288, N154, N390);
buf BUF1 (N942, N935);
not NOT1 (N943, N925);
buf BUF1 (N944, N941);
or OR2 (N945, N937, N265);
nor NOR3 (N946, N940, N25, N818);
not NOT1 (N947, N939);
nand NAND3 (N948, N942, N174, N14);
not NOT1 (N949, N934);
buf BUF1 (N950, N943);
nor NOR4 (N951, N946, N281, N807, N64);
nor NOR3 (N952, N947, N883, N554);
nand NAND4 (N953, N944, N357, N948, N125);
nand NAND3 (N954, N220, N5, N512);
buf BUF1 (N955, N952);
buf BUF1 (N956, N953);
not NOT1 (N957, N954);
xor XOR2 (N958, N957, N775);
not NOT1 (N959, N950);
nor NOR3 (N960, N956, N562, N448);
buf BUF1 (N961, N958);
and AND4 (N962, N960, N824, N790, N654);
nor NOR4 (N963, N945, N493, N64, N21);
not NOT1 (N964, N930);
xor XOR2 (N965, N955, N577);
and AND3 (N966, N951, N279, N74);
xor XOR2 (N967, N961, N272);
buf BUF1 (N968, N964);
nand NAND4 (N969, N968, N395, N219, N706);
not NOT1 (N970, N966);
and AND4 (N971, N967, N230, N388, N40);
not NOT1 (N972, N959);
and AND4 (N973, N949, N345, N511, N73);
buf BUF1 (N974, N969);
and AND2 (N975, N965, N47);
xor XOR2 (N976, N975, N778);
or OR3 (N977, N974, N637, N803);
not NOT1 (N978, N976);
xor XOR2 (N979, N970, N467);
or OR2 (N980, N963, N230);
buf BUF1 (N981, N962);
not NOT1 (N982, N919);
xor XOR2 (N983, N981, N126);
nand NAND2 (N984, N972, N237);
nor NOR4 (N985, N973, N704, N207, N819);
nor NOR3 (N986, N980, N156, N579);
or OR4 (N987, N932, N711, N400, N693);
buf BUF1 (N988, N985);
nor NOR2 (N989, N983, N410);
xor XOR2 (N990, N979, N415);
nor NOR2 (N991, N988, N113);
or OR4 (N992, N987, N786, N470, N363);
and AND4 (N993, N990, N482, N560, N635);
xor XOR2 (N994, N986, N540);
or OR2 (N995, N978, N581);
xor XOR2 (N996, N971, N117);
and AND4 (N997, N995, N509, N996, N782);
nand NAND4 (N998, N807, N775, N464, N232);
and AND2 (N999, N993, N306);
and AND4 (N1000, N999, N5, N659, N820);
or OR2 (N1001, N992, N100);
or OR2 (N1002, N989, N751);
xor XOR2 (N1003, N982, N290);
not NOT1 (N1004, N977);
or OR2 (N1005, N991, N560);
buf BUF1 (N1006, N1000);
and AND4 (N1007, N1003, N849, N150, N344);
and AND2 (N1008, N1006, N669);
or OR2 (N1009, N994, N9);
nand NAND3 (N1010, N1008, N968, N279);
buf BUF1 (N1011, N984);
buf BUF1 (N1012, N1011);
xor XOR2 (N1013, N1001, N889);
and AND4 (N1014, N997, N153, N589, N579);
nor NOR2 (N1015, N1005, N952);
and AND3 (N1016, N1004, N587, N680);
nor NOR2 (N1017, N1016, N890);
xor XOR2 (N1018, N1012, N473);
buf BUF1 (N1019, N1002);
xor XOR2 (N1020, N1014, N667);
and AND4 (N1021, N1013, N795, N55, N853);
nor NOR2 (N1022, N1017, N69);
or OR2 (N1023, N1022, N749);
not NOT1 (N1024, N1023);
buf BUF1 (N1025, N1010);
nand NAND2 (N1026, N1020, N670);
xor XOR2 (N1027, N1015, N8);
nand NAND4 (N1028, N1025, N806, N1027, N1004);
buf BUF1 (N1029, N568);
not NOT1 (N1030, N1029);
nand NAND2 (N1031, N1030, N967);
nand NAND3 (N1032, N1031, N1021, N418);
nand NAND3 (N1033, N301, N749, N251);
and AND4 (N1034, N1024, N326, N5, N404);
buf BUF1 (N1035, N1009);
buf BUF1 (N1036, N998);
buf BUF1 (N1037, N1028);
not NOT1 (N1038, N1033);
and AND2 (N1039, N1007, N793);
nor NOR3 (N1040, N1032, N462, N393);
and AND4 (N1041, N1039, N988, N545, N636);
nor NOR3 (N1042, N1019, N203, N300);
not NOT1 (N1043, N1035);
xor XOR2 (N1044, N1042, N893);
buf BUF1 (N1045, N1034);
not NOT1 (N1046, N1018);
or OR3 (N1047, N1045, N209, N990);
buf BUF1 (N1048, N1043);
and AND4 (N1049, N1026, N259, N456, N898);
buf BUF1 (N1050, N1046);
and AND2 (N1051, N1041, N717);
xor XOR2 (N1052, N1044, N67);
nor NOR2 (N1053, N1038, N315);
nand NAND2 (N1054, N1050, N708);
nor NOR3 (N1055, N1049, N942, N268);
xor XOR2 (N1056, N1054, N884);
or OR4 (N1057, N1051, N1056, N818, N63);
nand NAND4 (N1058, N240, N802, N995, N642);
or OR3 (N1059, N1036, N1026, N50);
or OR2 (N1060, N1052, N810);
and AND2 (N1061, N1037, N268);
and AND4 (N1062, N1047, N804, N962, N834);
and AND2 (N1063, N1048, N997);
or OR4 (N1064, N1063, N966, N91, N106);
or OR3 (N1065, N1064, N868, N290);
or OR2 (N1066, N1061, N287);
buf BUF1 (N1067, N1057);
nor NOR2 (N1068, N1053, N753);
or OR2 (N1069, N1055, N285);
buf BUF1 (N1070, N1062);
or OR4 (N1071, N1060, N270, N1000, N404);
xor XOR2 (N1072, N1059, N837);
buf BUF1 (N1073, N1066);
nand NAND2 (N1074, N1067, N699);
not NOT1 (N1075, N1072);
or OR3 (N1076, N1070, N1068, N260);
buf BUF1 (N1077, N1034);
xor XOR2 (N1078, N1069, N1014);
xor XOR2 (N1079, N1071, N194);
nor NOR3 (N1080, N1077, N7, N77);
and AND2 (N1081, N1074, N157);
not NOT1 (N1082, N1079);
nor NOR4 (N1083, N1081, N329, N720, N656);
and AND4 (N1084, N1040, N996, N1044, N771);
buf BUF1 (N1085, N1073);
nand NAND2 (N1086, N1083, N726);
nor NOR2 (N1087, N1065, N147);
or OR4 (N1088, N1086, N138, N886, N706);
buf BUF1 (N1089, N1087);
or OR4 (N1090, N1085, N542, N809, N1058);
not NOT1 (N1091, N17);
or OR4 (N1092, N1089, N677, N119, N277);
nor NOR4 (N1093, N1091, N147, N784, N242);
and AND2 (N1094, N1092, N249);
nor NOR2 (N1095, N1076, N282);
xor XOR2 (N1096, N1093, N854);
or OR2 (N1097, N1080, N348);
and AND4 (N1098, N1084, N596, N106, N1097);
nor NOR3 (N1099, N610, N416, N299);
not NOT1 (N1100, N1094);
nand NAND2 (N1101, N1082, N763);
nand NAND3 (N1102, N1100, N406, N510);
nand NAND2 (N1103, N1075, N486);
and AND3 (N1104, N1101, N1021, N545);
buf BUF1 (N1105, N1104);
nor NOR2 (N1106, N1096, N67);
and AND4 (N1107, N1102, N742, N404, N1085);
not NOT1 (N1108, N1105);
nor NOR2 (N1109, N1106, N325);
nand NAND4 (N1110, N1090, N781, N446, N679);
or OR3 (N1111, N1095, N278, N915);
buf BUF1 (N1112, N1098);
xor XOR2 (N1113, N1078, N402);
xor XOR2 (N1114, N1109, N1093);
or OR4 (N1115, N1111, N722, N747, N328);
nand NAND3 (N1116, N1115, N80, N545);
or OR3 (N1117, N1114, N100, N961);
not NOT1 (N1118, N1108);
or OR4 (N1119, N1107, N770, N475, N547);
buf BUF1 (N1120, N1112);
buf BUF1 (N1121, N1117);
and AND2 (N1122, N1121, N952);
nand NAND2 (N1123, N1113, N133);
xor XOR2 (N1124, N1088, N311);
and AND2 (N1125, N1110, N150);
xor XOR2 (N1126, N1103, N996);
nor NOR2 (N1127, N1120, N618);
xor XOR2 (N1128, N1122, N136);
or OR2 (N1129, N1119, N1112);
not NOT1 (N1130, N1126);
not NOT1 (N1131, N1127);
and AND3 (N1132, N1118, N614, N61);
not NOT1 (N1133, N1124);
not NOT1 (N1134, N1116);
or OR4 (N1135, N1132, N750, N732, N542);
or OR3 (N1136, N1125, N938, N871);
not NOT1 (N1137, N1134);
or OR3 (N1138, N1130, N742, N1068);
nand NAND4 (N1139, N1137, N552, N255, N904);
xor XOR2 (N1140, N1133, N205);
buf BUF1 (N1141, N1138);
not NOT1 (N1142, N1123);
xor XOR2 (N1143, N1139, N305);
not NOT1 (N1144, N1136);
and AND4 (N1145, N1143, N72, N1002, N1000);
nor NOR4 (N1146, N1141, N287, N187, N862);
and AND3 (N1147, N1142, N389, N289);
nand NAND4 (N1148, N1131, N1023, N414, N268);
not NOT1 (N1149, N1099);
nand NAND2 (N1150, N1144, N184);
not NOT1 (N1151, N1146);
not NOT1 (N1152, N1135);
buf BUF1 (N1153, N1147);
nor NOR2 (N1154, N1149, N542);
or OR2 (N1155, N1145, N410);
nor NOR4 (N1156, N1128, N402, N767, N690);
not NOT1 (N1157, N1129);
xor XOR2 (N1158, N1153, N130);
not NOT1 (N1159, N1154);
not NOT1 (N1160, N1150);
or OR2 (N1161, N1158, N48);
xor XOR2 (N1162, N1151, N59);
buf BUF1 (N1163, N1157);
nor NOR3 (N1164, N1159, N896, N816);
not NOT1 (N1165, N1156);
xor XOR2 (N1166, N1161, N519);
buf BUF1 (N1167, N1166);
nor NOR2 (N1168, N1167, N937);
or OR3 (N1169, N1164, N94, N898);
or OR3 (N1170, N1163, N583, N138);
not NOT1 (N1171, N1170);
nand NAND2 (N1172, N1152, N785);
nor NOR3 (N1173, N1168, N1142, N774);
or OR4 (N1174, N1173, N539, N1155, N563);
nor NOR3 (N1175, N587, N849, N405);
nand NAND3 (N1176, N1169, N726, N1048);
or OR3 (N1177, N1176, N883, N499);
nand NAND3 (N1178, N1160, N532, N526);
buf BUF1 (N1179, N1140);
or OR4 (N1180, N1174, N1168, N272, N1034);
and AND4 (N1181, N1148, N1006, N612, N748);
and AND2 (N1182, N1180, N193);
xor XOR2 (N1183, N1178, N394);
buf BUF1 (N1184, N1171);
xor XOR2 (N1185, N1165, N45);
nor NOR2 (N1186, N1181, N768);
or OR4 (N1187, N1177, N245, N646, N561);
buf BUF1 (N1188, N1185);
nand NAND4 (N1189, N1186, N188, N1054, N511);
nor NOR4 (N1190, N1187, N179, N388, N448);
nand NAND3 (N1191, N1188, N1169, N415);
buf BUF1 (N1192, N1191);
or OR2 (N1193, N1175, N265);
nor NOR3 (N1194, N1172, N302, N361);
and AND4 (N1195, N1184, N728, N1088, N471);
buf BUF1 (N1196, N1162);
not NOT1 (N1197, N1189);
and AND2 (N1198, N1195, N1168);
nand NAND2 (N1199, N1190, N900);
and AND2 (N1200, N1197, N919);
xor XOR2 (N1201, N1182, N421);
or OR4 (N1202, N1196, N321, N569, N270);
and AND4 (N1203, N1201, N570, N513, N1033);
and AND2 (N1204, N1203, N1044);
xor XOR2 (N1205, N1194, N80);
not NOT1 (N1206, N1183);
buf BUF1 (N1207, N1204);
buf BUF1 (N1208, N1202);
nor NOR3 (N1209, N1205, N1068, N1153);
or OR4 (N1210, N1193, N389, N1206, N1112);
and AND4 (N1211, N998, N665, N816, N1146);
nor NOR3 (N1212, N1210, N700, N286);
nand NAND4 (N1213, N1200, N392, N677, N134);
xor XOR2 (N1214, N1213, N192);
or OR4 (N1215, N1198, N585, N1214, N953);
nor NOR4 (N1216, N494, N56, N28, N844);
and AND4 (N1217, N1199, N644, N201, N264);
nor NOR4 (N1218, N1211, N355, N678, N604);
nand NAND4 (N1219, N1216, N372, N328, N943);
buf BUF1 (N1220, N1179);
buf BUF1 (N1221, N1217);
and AND2 (N1222, N1215, N936);
not NOT1 (N1223, N1220);
nor NOR2 (N1224, N1218, N918);
or OR4 (N1225, N1209, N1052, N190, N172);
and AND2 (N1226, N1208, N1055);
buf BUF1 (N1227, N1224);
nand NAND4 (N1228, N1212, N518, N332, N187);
xor XOR2 (N1229, N1219, N39);
nand NAND4 (N1230, N1207, N1189, N409, N425);
xor XOR2 (N1231, N1229, N515);
buf BUF1 (N1232, N1192);
not NOT1 (N1233, N1226);
not NOT1 (N1234, N1230);
nor NOR4 (N1235, N1227, N40, N124, N409);
buf BUF1 (N1236, N1233);
nor NOR4 (N1237, N1225, N6, N232, N972);
buf BUF1 (N1238, N1223);
or OR3 (N1239, N1238, N1222, N1164);
not NOT1 (N1240, N698);
not NOT1 (N1241, N1236);
not NOT1 (N1242, N1235);
not NOT1 (N1243, N1231);
buf BUF1 (N1244, N1234);
nand NAND4 (N1245, N1221, N1231, N1076, N783);
nand NAND3 (N1246, N1245, N173, N331);
or OR3 (N1247, N1246, N909, N1234);
nor NOR3 (N1248, N1242, N583, N1001);
nand NAND4 (N1249, N1243, N794, N186, N462);
nand NAND2 (N1250, N1237, N877);
nand NAND3 (N1251, N1228, N139, N1165);
or OR2 (N1252, N1248, N649);
nor NOR2 (N1253, N1239, N1030);
nor NOR2 (N1254, N1247, N999);
and AND2 (N1255, N1241, N38);
nor NOR2 (N1256, N1252, N178);
or OR2 (N1257, N1253, N542);
nand NAND4 (N1258, N1232, N137, N1252, N162);
or OR2 (N1259, N1250, N1005);
xor XOR2 (N1260, N1254, N505);
buf BUF1 (N1261, N1257);
and AND3 (N1262, N1261, N271, N247);
nor NOR3 (N1263, N1259, N1041, N379);
xor XOR2 (N1264, N1255, N630);
nand NAND2 (N1265, N1263, N221);
not NOT1 (N1266, N1244);
nor NOR3 (N1267, N1240, N822, N82);
and AND2 (N1268, N1265, N488);
not NOT1 (N1269, N1249);
xor XOR2 (N1270, N1264, N305);
and AND4 (N1271, N1269, N73, N505, N543);
nand NAND2 (N1272, N1262, N1033);
buf BUF1 (N1273, N1266);
nor NOR4 (N1274, N1260, N636, N42, N556);
or OR3 (N1275, N1258, N693, N1174);
nand NAND2 (N1276, N1251, N1174);
nand NAND2 (N1277, N1270, N961);
buf BUF1 (N1278, N1256);
not NOT1 (N1279, N1273);
and AND3 (N1280, N1279, N908, N372);
or OR2 (N1281, N1277, N506);
xor XOR2 (N1282, N1280, N957);
nand NAND4 (N1283, N1276, N269, N279, N1161);
xor XOR2 (N1284, N1275, N845);
or OR3 (N1285, N1278, N260, N1081);
and AND4 (N1286, N1272, N792, N425, N83);
xor XOR2 (N1287, N1285, N748);
nand NAND2 (N1288, N1274, N336);
or OR2 (N1289, N1288, N47);
or OR4 (N1290, N1271, N930, N424, N496);
buf BUF1 (N1291, N1281);
nor NOR2 (N1292, N1268, N439);
buf BUF1 (N1293, N1289);
nand NAND2 (N1294, N1290, N1220);
not NOT1 (N1295, N1294);
nand NAND2 (N1296, N1287, N1098);
or OR3 (N1297, N1291, N546, N766);
buf BUF1 (N1298, N1296);
not NOT1 (N1299, N1297);
xor XOR2 (N1300, N1283, N838);
nor NOR3 (N1301, N1295, N961, N404);
not NOT1 (N1302, N1284);
nor NOR3 (N1303, N1267, N205, N350);
xor XOR2 (N1304, N1300, N683);
not NOT1 (N1305, N1292);
xor XOR2 (N1306, N1282, N457);
buf BUF1 (N1307, N1301);
and AND3 (N1308, N1305, N330, N1166);
nor NOR2 (N1309, N1304, N321);
not NOT1 (N1310, N1298);
nand NAND3 (N1311, N1293, N1, N951);
nand NAND4 (N1312, N1299, N247, N27, N64);
nor NOR2 (N1313, N1306, N1250);
xor XOR2 (N1314, N1308, N1299);
buf BUF1 (N1315, N1311);
nand NAND4 (N1316, N1313, N768, N966, N143);
nand NAND3 (N1317, N1307, N1171, N468);
buf BUF1 (N1318, N1314);
not NOT1 (N1319, N1318);
xor XOR2 (N1320, N1315, N820);
nor NOR2 (N1321, N1303, N44);
and AND3 (N1322, N1320, N35, N950);
xor XOR2 (N1323, N1319, N232);
nand NAND3 (N1324, N1316, N510, N476);
and AND2 (N1325, N1321, N1150);
nand NAND4 (N1326, N1322, N9, N924, N1266);
xor XOR2 (N1327, N1317, N685);
buf BUF1 (N1328, N1325);
buf BUF1 (N1329, N1327);
xor XOR2 (N1330, N1329, N932);
nand NAND2 (N1331, N1323, N948);
nor NOR2 (N1332, N1302, N607);
and AND4 (N1333, N1310, N690, N844, N1331);
nand NAND4 (N1334, N762, N1211, N473, N823);
nor NOR3 (N1335, N1333, N1164, N459);
or OR4 (N1336, N1335, N222, N635, N476);
xor XOR2 (N1337, N1336, N454);
not NOT1 (N1338, N1328);
or OR4 (N1339, N1286, N1302, N219, N504);
buf BUF1 (N1340, N1337);
buf BUF1 (N1341, N1309);
nor NOR3 (N1342, N1334, N952, N589);
not NOT1 (N1343, N1332);
nor NOR4 (N1344, N1312, N948, N183, N1039);
nor NOR4 (N1345, N1326, N826, N1268, N276);
or OR3 (N1346, N1340, N488, N1039);
nand NAND2 (N1347, N1330, N790);
xor XOR2 (N1348, N1338, N748);
not NOT1 (N1349, N1341);
xor XOR2 (N1350, N1339, N169);
xor XOR2 (N1351, N1324, N1259);
nor NOR4 (N1352, N1350, N795, N1271, N672);
not NOT1 (N1353, N1344);
nor NOR4 (N1354, N1351, N1261, N848, N831);
not NOT1 (N1355, N1352);
not NOT1 (N1356, N1342);
nor NOR4 (N1357, N1349, N321, N1325, N22);
and AND3 (N1358, N1357, N798, N543);
nor NOR4 (N1359, N1356, N343, N26, N703);
buf BUF1 (N1360, N1359);
or OR2 (N1361, N1346, N1202);
not NOT1 (N1362, N1348);
or OR2 (N1363, N1361, N548);
or OR2 (N1364, N1343, N345);
and AND2 (N1365, N1347, N376);
buf BUF1 (N1366, N1363);
not NOT1 (N1367, N1358);
nand NAND3 (N1368, N1353, N530, N800);
or OR2 (N1369, N1354, N1);
not NOT1 (N1370, N1355);
nor NOR2 (N1371, N1369, N267);
or OR2 (N1372, N1368, N589);
nor NOR3 (N1373, N1372, N20, N775);
or OR4 (N1374, N1345, N1188, N1289, N540);
nor NOR4 (N1375, N1362, N885, N1088, N1129);
not NOT1 (N1376, N1371);
or OR4 (N1377, N1370, N74, N138, N567);
or OR3 (N1378, N1366, N908, N571);
and AND4 (N1379, N1376, N970, N255, N1308);
nand NAND4 (N1380, N1379, N151, N1275, N824);
or OR3 (N1381, N1364, N99, N1291);
buf BUF1 (N1382, N1365);
buf BUF1 (N1383, N1373);
nor NOR4 (N1384, N1375, N1327, N1207, N603);
not NOT1 (N1385, N1381);
or OR2 (N1386, N1382, N963);
not NOT1 (N1387, N1374);
nand NAND4 (N1388, N1385, N149, N792, N1174);
buf BUF1 (N1389, N1360);
or OR4 (N1390, N1386, N471, N1310, N557);
buf BUF1 (N1391, N1377);
or OR4 (N1392, N1387, N487, N642, N188);
buf BUF1 (N1393, N1384);
and AND2 (N1394, N1378, N1323);
xor XOR2 (N1395, N1390, N194);
nor NOR4 (N1396, N1367, N602, N451, N585);
xor XOR2 (N1397, N1383, N468);
nor NOR3 (N1398, N1392, N299, N551);
nand NAND3 (N1399, N1398, N1258, N56);
not NOT1 (N1400, N1394);
xor XOR2 (N1401, N1397, N1030);
nor NOR3 (N1402, N1389, N1368, N674);
or OR4 (N1403, N1393, N777, N697, N953);
buf BUF1 (N1404, N1400);
nand NAND2 (N1405, N1399, N333);
xor XOR2 (N1406, N1402, N979);
or OR2 (N1407, N1405, N632);
nor NOR4 (N1408, N1404, N928, N1317, N1058);
xor XOR2 (N1409, N1391, N13);
and AND2 (N1410, N1408, N819);
xor XOR2 (N1411, N1407, N158);
not NOT1 (N1412, N1396);
not NOT1 (N1413, N1411);
or OR2 (N1414, N1403, N711);
nor NOR2 (N1415, N1410, N1041);
nor NOR4 (N1416, N1415, N811, N538, N621);
and AND4 (N1417, N1413, N316, N859, N575);
nor NOR4 (N1418, N1416, N679, N1360, N1231);
xor XOR2 (N1419, N1417, N562);
or OR4 (N1420, N1419, N462, N1351, N1344);
nor NOR2 (N1421, N1414, N1048);
not NOT1 (N1422, N1421);
not NOT1 (N1423, N1380);
nor NOR4 (N1424, N1420, N85, N85, N43);
nor NOR3 (N1425, N1395, N1246, N591);
and AND2 (N1426, N1401, N483);
buf BUF1 (N1427, N1388);
not NOT1 (N1428, N1426);
xor XOR2 (N1429, N1418, N325);
and AND2 (N1430, N1429, N1290);
xor XOR2 (N1431, N1412, N920);
or OR4 (N1432, N1430, N735, N1134, N609);
xor XOR2 (N1433, N1406, N301);
and AND3 (N1434, N1422, N91, N582);
not NOT1 (N1435, N1425);
xor XOR2 (N1436, N1434, N973);
and AND2 (N1437, N1431, N232);
nor NOR4 (N1438, N1437, N454, N473, N183);
or OR4 (N1439, N1435, N300, N249, N1339);
or OR3 (N1440, N1423, N412, N1355);
not NOT1 (N1441, N1433);
or OR3 (N1442, N1428, N1300, N631);
or OR3 (N1443, N1432, N511, N1075);
nand NAND3 (N1444, N1439, N210, N11);
buf BUF1 (N1445, N1444);
or OR2 (N1446, N1436, N217);
nand NAND2 (N1447, N1438, N314);
xor XOR2 (N1448, N1440, N315);
nor NOR2 (N1449, N1448, N1135);
and AND4 (N1450, N1445, N265, N564, N107);
buf BUF1 (N1451, N1424);
and AND4 (N1452, N1446, N228, N1262, N915);
nor NOR4 (N1453, N1409, N655, N386, N655);
nor NOR4 (N1454, N1449, N368, N1290, N411);
and AND3 (N1455, N1427, N1091, N371);
nor NOR2 (N1456, N1455, N851);
buf BUF1 (N1457, N1452);
nand NAND3 (N1458, N1442, N484, N1101);
and AND4 (N1459, N1450, N247, N358, N1449);
xor XOR2 (N1460, N1457, N1132);
not NOT1 (N1461, N1459);
nor NOR4 (N1462, N1461, N501, N124, N986);
not NOT1 (N1463, N1462);
not NOT1 (N1464, N1463);
nor NOR3 (N1465, N1458, N388, N632);
or OR3 (N1466, N1464, N1282, N1255);
nand NAND3 (N1467, N1454, N785, N420);
nand NAND2 (N1468, N1451, N1274);
nand NAND2 (N1469, N1466, N182);
xor XOR2 (N1470, N1441, N209);
or OR2 (N1471, N1467, N611);
xor XOR2 (N1472, N1471, N257);
nor NOR4 (N1473, N1453, N1393, N98, N1423);
nor NOR2 (N1474, N1456, N917);
nor NOR3 (N1475, N1447, N420, N1184);
nor NOR3 (N1476, N1470, N1336, N928);
xor XOR2 (N1477, N1460, N636);
nand NAND2 (N1478, N1465, N1279);
nor NOR2 (N1479, N1478, N800);
and AND3 (N1480, N1469, N774, N1413);
buf BUF1 (N1481, N1477);
nand NAND2 (N1482, N1443, N1228);
or OR3 (N1483, N1481, N1468, N302);
xor XOR2 (N1484, N1299, N932);
or OR2 (N1485, N1480, N1172);
or OR3 (N1486, N1474, N1345, N388);
nor NOR2 (N1487, N1485, N400);
or OR3 (N1488, N1487, N1295, N1148);
and AND3 (N1489, N1483, N559, N372);
nand NAND3 (N1490, N1482, N180, N219);
nor NOR2 (N1491, N1479, N1171);
xor XOR2 (N1492, N1491, N563);
buf BUF1 (N1493, N1472);
and AND4 (N1494, N1476, N1217, N125, N1380);
buf BUF1 (N1495, N1492);
and AND2 (N1496, N1489, N804);
nor NOR2 (N1497, N1494, N588);
xor XOR2 (N1498, N1486, N152);
xor XOR2 (N1499, N1475, N908);
or OR3 (N1500, N1484, N1, N1255);
and AND3 (N1501, N1499, N1421, N751);
and AND4 (N1502, N1493, N263, N33, N1279);
xor XOR2 (N1503, N1501, N1024);
not NOT1 (N1504, N1490);
or OR3 (N1505, N1496, N1036, N1411);
xor XOR2 (N1506, N1495, N721);
xor XOR2 (N1507, N1473, N1050);
not NOT1 (N1508, N1502);
buf BUF1 (N1509, N1503);
xor XOR2 (N1510, N1509, N266);
buf BUF1 (N1511, N1488);
xor XOR2 (N1512, N1505, N1435);
and AND2 (N1513, N1512, N1371);
not NOT1 (N1514, N1507);
or OR4 (N1515, N1497, N522, N872, N1242);
not NOT1 (N1516, N1511);
or OR4 (N1517, N1510, N1047, N386, N148);
nor NOR2 (N1518, N1504, N311);
or OR3 (N1519, N1506, N1295, N365);
or OR3 (N1520, N1516, N442, N1439);
and AND3 (N1521, N1519, N623, N471);
and AND3 (N1522, N1521, N1001, N656);
nor NOR2 (N1523, N1508, N1300);
and AND4 (N1524, N1518, N1328, N823, N268);
and AND3 (N1525, N1500, N378, N1156);
and AND3 (N1526, N1514, N1000, N1344);
not NOT1 (N1527, N1498);
or OR3 (N1528, N1525, N1130, N674);
not NOT1 (N1529, N1520);
buf BUF1 (N1530, N1526);
and AND3 (N1531, N1528, N563, N817);
not NOT1 (N1532, N1517);
buf BUF1 (N1533, N1531);
nand NAND2 (N1534, N1524, N356);
and AND3 (N1535, N1529, N455, N513);
and AND2 (N1536, N1533, N1500);
buf BUF1 (N1537, N1522);
or OR2 (N1538, N1534, N974);
not NOT1 (N1539, N1513);
not NOT1 (N1540, N1537);
buf BUF1 (N1541, N1538);
nand NAND4 (N1542, N1515, N1309, N723, N365);
not NOT1 (N1543, N1539);
buf BUF1 (N1544, N1535);
xor XOR2 (N1545, N1536, N1078);
nand NAND2 (N1546, N1523, N1078);
nor NOR3 (N1547, N1530, N319, N869);
and AND4 (N1548, N1540, N351, N600, N1466);
and AND2 (N1549, N1542, N1293);
xor XOR2 (N1550, N1546, N922);
and AND4 (N1551, N1549, N473, N159, N1189);
buf BUF1 (N1552, N1550);
buf BUF1 (N1553, N1532);
nand NAND2 (N1554, N1551, N660);
nor NOR3 (N1555, N1547, N677, N1502);
not NOT1 (N1556, N1541);
not NOT1 (N1557, N1527);
buf BUF1 (N1558, N1557);
buf BUF1 (N1559, N1543);
xor XOR2 (N1560, N1554, N1279);
nand NAND2 (N1561, N1544, N1291);
buf BUF1 (N1562, N1553);
or OR4 (N1563, N1558, N1315, N660, N325);
nand NAND3 (N1564, N1545, N231, N1435);
xor XOR2 (N1565, N1548, N1342);
not NOT1 (N1566, N1563);
and AND2 (N1567, N1564, N283);
nand NAND3 (N1568, N1555, N1420, N899);
nor NOR2 (N1569, N1559, N407);
xor XOR2 (N1570, N1566, N1114);
nand NAND4 (N1571, N1565, N1082, N821, N184);
nor NOR2 (N1572, N1568, N1427);
and AND3 (N1573, N1562, N945, N326);
buf BUF1 (N1574, N1567);
and AND4 (N1575, N1561, N469, N579, N379);
and AND4 (N1576, N1575, N969, N146, N144);
and AND4 (N1577, N1560, N802, N1235, N985);
or OR3 (N1578, N1574, N375, N1458);
not NOT1 (N1579, N1573);
or OR4 (N1580, N1552, N1500, N237, N697);
not NOT1 (N1581, N1571);
nor NOR2 (N1582, N1577, N1418);
or OR4 (N1583, N1581, N1480, N250, N1444);
buf BUF1 (N1584, N1578);
nor NOR3 (N1585, N1584, N455, N788);
and AND2 (N1586, N1579, N723);
not NOT1 (N1587, N1585);
nand NAND4 (N1588, N1572, N1531, N1114, N1211);
nor NOR4 (N1589, N1556, N225, N1072, N299);
nand NAND3 (N1590, N1583, N616, N846);
not NOT1 (N1591, N1589);
or OR3 (N1592, N1580, N1582, N905);
and AND4 (N1593, N13, N640, N157, N336);
nand NAND3 (N1594, N1576, N459, N515);
nand NAND4 (N1595, N1569, N1329, N1374, N783);
buf BUF1 (N1596, N1592);
not NOT1 (N1597, N1590);
or OR3 (N1598, N1587, N945, N313);
nor NOR4 (N1599, N1594, N902, N483, N90);
and AND3 (N1600, N1570, N1089, N543);
not NOT1 (N1601, N1596);
nor NOR4 (N1602, N1597, N401, N1163, N1389);
or OR2 (N1603, N1588, N1485);
xor XOR2 (N1604, N1600, N294);
and AND4 (N1605, N1593, N1432, N336, N291);
nor NOR4 (N1606, N1603, N1361, N692, N1097);
or OR2 (N1607, N1604, N553);
not NOT1 (N1608, N1591);
not NOT1 (N1609, N1605);
nor NOR4 (N1610, N1606, N913, N296, N1400);
and AND2 (N1611, N1595, N1201);
nand NAND4 (N1612, N1602, N58, N1186, N511);
nand NAND3 (N1613, N1599, N1084, N914);
buf BUF1 (N1614, N1609);
nor NOR2 (N1615, N1601, N1394);
buf BUF1 (N1616, N1607);
buf BUF1 (N1617, N1608);
xor XOR2 (N1618, N1614, N438);
not NOT1 (N1619, N1610);
nor NOR4 (N1620, N1612, N903, N167, N887);
or OR4 (N1621, N1611, N1172, N41, N288);
buf BUF1 (N1622, N1616);
buf BUF1 (N1623, N1615);
buf BUF1 (N1624, N1619);
and AND2 (N1625, N1617, N886);
xor XOR2 (N1626, N1618, N1105);
xor XOR2 (N1627, N1623, N196);
nor NOR4 (N1628, N1586, N997, N1205, N434);
and AND3 (N1629, N1625, N675, N1331);
nand NAND3 (N1630, N1628, N1241, N647);
buf BUF1 (N1631, N1630);
and AND3 (N1632, N1613, N1343, N1373);
nand NAND4 (N1633, N1631, N1196, N338, N739);
not NOT1 (N1634, N1622);
not NOT1 (N1635, N1633);
nand NAND3 (N1636, N1598, N1353, N1336);
nand NAND4 (N1637, N1627, N34, N495, N1015);
buf BUF1 (N1638, N1634);
or OR4 (N1639, N1638, N1507, N1043, N366);
nand NAND4 (N1640, N1636, N1578, N585, N84);
or OR2 (N1641, N1629, N499);
buf BUF1 (N1642, N1639);
buf BUF1 (N1643, N1642);
buf BUF1 (N1644, N1640);
not NOT1 (N1645, N1644);
nor NOR2 (N1646, N1641, N372);
buf BUF1 (N1647, N1621);
xor XOR2 (N1648, N1646, N590);
nor NOR2 (N1649, N1645, N904);
and AND4 (N1650, N1649, N667, N1277, N1485);
nor NOR2 (N1651, N1648, N459);
or OR3 (N1652, N1626, N515, N88);
not NOT1 (N1653, N1624);
and AND2 (N1654, N1632, N229);
or OR3 (N1655, N1643, N1178, N1417);
nor NOR2 (N1656, N1637, N1427);
nor NOR2 (N1657, N1655, N1363);
and AND4 (N1658, N1620, N1351, N884, N1615);
buf BUF1 (N1659, N1658);
or OR2 (N1660, N1647, N849);
nor NOR3 (N1661, N1654, N1352, N115);
buf BUF1 (N1662, N1653);
not NOT1 (N1663, N1659);
buf BUF1 (N1664, N1661);
xor XOR2 (N1665, N1663, N733);
not NOT1 (N1666, N1635);
or OR2 (N1667, N1666, N797);
not NOT1 (N1668, N1652);
nand NAND4 (N1669, N1664, N818, N624, N1649);
and AND4 (N1670, N1656, N1090, N1070, N237);
nand NAND2 (N1671, N1650, N93);
and AND3 (N1672, N1651, N402, N490);
and AND3 (N1673, N1669, N505, N1313);
xor XOR2 (N1674, N1671, N1322);
buf BUF1 (N1675, N1660);
xor XOR2 (N1676, N1667, N104);
xor XOR2 (N1677, N1670, N796);
or OR2 (N1678, N1673, N1026);
nand NAND4 (N1679, N1657, N1523, N630, N1357);
nor NOR2 (N1680, N1679, N1360);
or OR4 (N1681, N1675, N590, N913, N1496);
nor NOR3 (N1682, N1680, N1050, N1093);
buf BUF1 (N1683, N1678);
nand NAND3 (N1684, N1682, N1400, N65);
xor XOR2 (N1685, N1668, N439);
and AND3 (N1686, N1665, N322, N577);
nor NOR4 (N1687, N1683, N539, N1417, N106);
buf BUF1 (N1688, N1687);
buf BUF1 (N1689, N1674);
nand NAND2 (N1690, N1685, N590);
or OR3 (N1691, N1677, N500, N265);
not NOT1 (N1692, N1662);
buf BUF1 (N1693, N1684);
and AND3 (N1694, N1672, N113, N642);
xor XOR2 (N1695, N1690, N1052);
buf BUF1 (N1696, N1686);
or OR2 (N1697, N1681, N1002);
buf BUF1 (N1698, N1695);
xor XOR2 (N1699, N1697, N1398);
and AND2 (N1700, N1694, N1699);
nor NOR2 (N1701, N1544, N1393);
nor NOR4 (N1702, N1689, N37, N1340, N1524);
xor XOR2 (N1703, N1691, N573);
not NOT1 (N1704, N1701);
not NOT1 (N1705, N1688);
nor NOR2 (N1706, N1676, N136);
not NOT1 (N1707, N1700);
nand NAND2 (N1708, N1702, N424);
nand NAND3 (N1709, N1693, N1100, N1229);
and AND4 (N1710, N1696, N660, N940, N113);
buf BUF1 (N1711, N1708);
and AND2 (N1712, N1707, N154);
not NOT1 (N1713, N1704);
nor NOR3 (N1714, N1713, N711, N1082);
and AND4 (N1715, N1705, N1003, N1074, N482);
or OR3 (N1716, N1706, N872, N1219);
or OR4 (N1717, N1711, N44, N1494, N1409);
xor XOR2 (N1718, N1714, N1715);
nand NAND2 (N1719, N873, N1538);
nand NAND2 (N1720, N1698, N357);
or OR3 (N1721, N1720, N356, N955);
buf BUF1 (N1722, N1716);
not NOT1 (N1723, N1703);
or OR2 (N1724, N1717, N55);
nor NOR3 (N1725, N1724, N887, N123);
and AND2 (N1726, N1725, N105);
buf BUF1 (N1727, N1719);
xor XOR2 (N1728, N1726, N499);
and AND2 (N1729, N1692, N954);
xor XOR2 (N1730, N1722, N1110);
or OR3 (N1731, N1727, N1636, N904);
buf BUF1 (N1732, N1718);
and AND4 (N1733, N1728, N202, N1142, N572);
xor XOR2 (N1734, N1709, N1398);
and AND3 (N1735, N1729, N779, N1511);
or OR3 (N1736, N1734, N534, N1631);
not NOT1 (N1737, N1712);
nor NOR2 (N1738, N1737, N1209);
xor XOR2 (N1739, N1733, N635);
or OR2 (N1740, N1710, N1726);
nand NAND4 (N1741, N1738, N308, N801, N1167);
and AND4 (N1742, N1721, N602, N415, N394);
or OR2 (N1743, N1740, N830);
nand NAND2 (N1744, N1741, N195);
and AND3 (N1745, N1739, N1204, N276);
buf BUF1 (N1746, N1736);
nand NAND2 (N1747, N1742, N1521);
nand NAND2 (N1748, N1743, N932);
and AND2 (N1749, N1746, N1628);
or OR4 (N1750, N1744, N1164, N663, N653);
xor XOR2 (N1751, N1749, N1108);
or OR4 (N1752, N1731, N1176, N689, N121);
xor XOR2 (N1753, N1747, N411);
and AND4 (N1754, N1753, N1055, N1591, N754);
not NOT1 (N1755, N1730);
or OR4 (N1756, N1745, N415, N622, N926);
nand NAND4 (N1757, N1750, N1617, N407, N1016);
buf BUF1 (N1758, N1755);
xor XOR2 (N1759, N1756, N251);
nand NAND4 (N1760, N1732, N1200, N696, N1699);
buf BUF1 (N1761, N1723);
buf BUF1 (N1762, N1759);
xor XOR2 (N1763, N1751, N1567);
buf BUF1 (N1764, N1760);
buf BUF1 (N1765, N1757);
or OR3 (N1766, N1752, N568, N776);
or OR4 (N1767, N1735, N1304, N1660, N251);
not NOT1 (N1768, N1748);
buf BUF1 (N1769, N1761);
or OR2 (N1770, N1766, N628);
and AND2 (N1771, N1769, N372);
or OR3 (N1772, N1758, N1261, N858);
xor XOR2 (N1773, N1762, N1030);
xor XOR2 (N1774, N1770, N372);
buf BUF1 (N1775, N1763);
nand NAND4 (N1776, N1772, N1621, N1722, N619);
xor XOR2 (N1777, N1771, N35);
and AND3 (N1778, N1775, N947, N639);
and AND4 (N1779, N1773, N190, N13, N1147);
or OR4 (N1780, N1776, N927, N561, N665);
and AND3 (N1781, N1780, N1378, N782);
buf BUF1 (N1782, N1767);
and AND2 (N1783, N1778, N1313);
and AND4 (N1784, N1754, N643, N910, N20);
xor XOR2 (N1785, N1781, N750);
nor NOR4 (N1786, N1783, N1302, N1456, N568);
buf BUF1 (N1787, N1765);
nor NOR4 (N1788, N1768, N66, N556, N881);
nand NAND2 (N1789, N1785, N1274);
not NOT1 (N1790, N1786);
buf BUF1 (N1791, N1788);
nand NAND4 (N1792, N1791, N663, N1736, N509);
nor NOR2 (N1793, N1764, N118);
xor XOR2 (N1794, N1790, N930);
nor NOR2 (N1795, N1774, N838);
and AND3 (N1796, N1792, N140, N743);
nand NAND3 (N1797, N1796, N166, N831);
nor NOR3 (N1798, N1789, N859, N1185);
xor XOR2 (N1799, N1784, N1196);
buf BUF1 (N1800, N1797);
or OR2 (N1801, N1799, N398);
nor NOR3 (N1802, N1795, N1158, N318);
not NOT1 (N1803, N1777);
and AND2 (N1804, N1779, N536);
xor XOR2 (N1805, N1803, N1434);
xor XOR2 (N1806, N1801, N1271);
and AND4 (N1807, N1802, N93, N352, N1599);
buf BUF1 (N1808, N1800);
nand NAND2 (N1809, N1787, N675);
or OR2 (N1810, N1806, N929);
and AND4 (N1811, N1794, N214, N343, N734);
nor NOR4 (N1812, N1804, N987, N1528, N324);
not NOT1 (N1813, N1812);
not NOT1 (N1814, N1808);
and AND3 (N1815, N1782, N1575, N436);
xor XOR2 (N1816, N1811, N451);
and AND2 (N1817, N1809, N635);
xor XOR2 (N1818, N1814, N1711);
nor NOR2 (N1819, N1813, N1429);
or OR4 (N1820, N1816, N965, N1173, N528);
nand NAND3 (N1821, N1805, N96, N511);
and AND4 (N1822, N1817, N682, N81, N1233);
nand NAND2 (N1823, N1793, N890);
buf BUF1 (N1824, N1820);
xor XOR2 (N1825, N1798, N1480);
or OR2 (N1826, N1822, N1539);
not NOT1 (N1827, N1819);
xor XOR2 (N1828, N1807, N1117);
or OR2 (N1829, N1826, N559);
buf BUF1 (N1830, N1829);
not NOT1 (N1831, N1815);
nor NOR4 (N1832, N1810, N206, N86, N188);
xor XOR2 (N1833, N1824, N974);
not NOT1 (N1834, N1823);
buf BUF1 (N1835, N1830);
nor NOR2 (N1836, N1825, N816);
or OR3 (N1837, N1827, N183, N75);
and AND2 (N1838, N1831, N1779);
not NOT1 (N1839, N1834);
xor XOR2 (N1840, N1821, N766);
and AND2 (N1841, N1833, N1621);
nor NOR2 (N1842, N1828, N1331);
buf BUF1 (N1843, N1842);
nand NAND4 (N1844, N1835, N29, N113, N1185);
xor XOR2 (N1845, N1818, N598);
xor XOR2 (N1846, N1838, N252);
nor NOR2 (N1847, N1843, N964);
xor XOR2 (N1848, N1832, N363);
and AND4 (N1849, N1836, N726, N1149, N1275);
xor XOR2 (N1850, N1848, N21);
not NOT1 (N1851, N1840);
buf BUF1 (N1852, N1845);
xor XOR2 (N1853, N1850, N369);
nor NOR4 (N1854, N1853, N1243, N961, N696);
nand NAND3 (N1855, N1846, N1085, N888);
xor XOR2 (N1856, N1855, N1645);
nand NAND4 (N1857, N1837, N203, N1169, N822);
and AND3 (N1858, N1847, N298, N1603);
nand NAND2 (N1859, N1841, N521);
and AND3 (N1860, N1849, N661, N1344);
buf BUF1 (N1861, N1852);
xor XOR2 (N1862, N1854, N252);
buf BUF1 (N1863, N1859);
not NOT1 (N1864, N1858);
xor XOR2 (N1865, N1861, N1534);
xor XOR2 (N1866, N1862, N1516);
and AND3 (N1867, N1865, N1801, N1819);
xor XOR2 (N1868, N1866, N1363);
nor NOR3 (N1869, N1839, N475, N125);
and AND4 (N1870, N1851, N365, N23, N1771);
not NOT1 (N1871, N1868);
not NOT1 (N1872, N1856);
buf BUF1 (N1873, N1857);
nand NAND3 (N1874, N1844, N878, N425);
nor NOR3 (N1875, N1860, N303, N1693);
not NOT1 (N1876, N1875);
not NOT1 (N1877, N1872);
nand NAND3 (N1878, N1874, N1794, N1348);
nor NOR2 (N1879, N1864, N1818);
buf BUF1 (N1880, N1878);
not NOT1 (N1881, N1880);
buf BUF1 (N1882, N1876);
and AND3 (N1883, N1870, N934, N1356);
nand NAND3 (N1884, N1863, N1471, N552);
xor XOR2 (N1885, N1873, N1744);
not NOT1 (N1886, N1882);
and AND4 (N1887, N1886, N929, N1668, N603);
nand NAND4 (N1888, N1867, N1841, N315, N498);
xor XOR2 (N1889, N1883, N1369);
or OR3 (N1890, N1885, N695, N17);
not NOT1 (N1891, N1879);
or OR3 (N1892, N1884, N562, N371);
or OR4 (N1893, N1891, N712, N1238, N801);
nand NAND2 (N1894, N1892, N1564);
nor NOR4 (N1895, N1889, N700, N1415, N693);
not NOT1 (N1896, N1888);
nand NAND4 (N1897, N1871, N1703, N1643, N585);
xor XOR2 (N1898, N1894, N812);
and AND4 (N1899, N1895, N1409, N897, N699);
buf BUF1 (N1900, N1897);
and AND2 (N1901, N1887, N20);
not NOT1 (N1902, N1893);
buf BUF1 (N1903, N1881);
not NOT1 (N1904, N1877);
xor XOR2 (N1905, N1896, N1014);
buf BUF1 (N1906, N1869);
nor NOR3 (N1907, N1906, N1308, N535);
nand NAND4 (N1908, N1898, N1382, N1778, N1712);
not NOT1 (N1909, N1905);
nand NAND4 (N1910, N1899, N1350, N1830, N1846);
not NOT1 (N1911, N1902);
nand NAND4 (N1912, N1911, N197, N1666, N1655);
xor XOR2 (N1913, N1900, N1446);
not NOT1 (N1914, N1909);
not NOT1 (N1915, N1912);
buf BUF1 (N1916, N1914);
xor XOR2 (N1917, N1910, N792);
buf BUF1 (N1918, N1908);
buf BUF1 (N1919, N1903);
and AND3 (N1920, N1913, N210, N909);
or OR2 (N1921, N1916, N10);
and AND4 (N1922, N1921, N254, N341, N484);
nand NAND4 (N1923, N1907, N1297, N851, N1616);
nand NAND4 (N1924, N1890, N949, N1874, N515);
nand NAND3 (N1925, N1919, N404, N314);
not NOT1 (N1926, N1923);
xor XOR2 (N1927, N1924, N941);
not NOT1 (N1928, N1920);
not NOT1 (N1929, N1915);
or OR4 (N1930, N1904, N1740, N1148, N465);
buf BUF1 (N1931, N1928);
nor NOR4 (N1932, N1922, N779, N1700, N1654);
xor XOR2 (N1933, N1925, N503);
nand NAND3 (N1934, N1901, N710, N398);
xor XOR2 (N1935, N1927, N336);
and AND2 (N1936, N1932, N1618);
buf BUF1 (N1937, N1926);
nor NOR3 (N1938, N1930, N1716, N164);
nor NOR4 (N1939, N1931, N1150, N442, N15);
buf BUF1 (N1940, N1929);
xor XOR2 (N1941, N1938, N321);
xor XOR2 (N1942, N1940, N925);
not NOT1 (N1943, N1939);
or OR4 (N1944, N1917, N443, N991, N1297);
not NOT1 (N1945, N1936);
not NOT1 (N1946, N1934);
nand NAND3 (N1947, N1944, N197, N523);
nand NAND3 (N1948, N1946, N1619, N1121);
not NOT1 (N1949, N1943);
not NOT1 (N1950, N1935);
xor XOR2 (N1951, N1918, N380);
nor NOR2 (N1952, N1950, N410);
xor XOR2 (N1953, N1948, N926);
nor NOR3 (N1954, N1941, N533, N174);
nor NOR3 (N1955, N1933, N160, N1695);
nand NAND4 (N1956, N1945, N456, N1141, N842);
nor NOR2 (N1957, N1955, N1880);
nand NAND4 (N1958, N1942, N1417, N1605, N1636);
or OR3 (N1959, N1956, N1586, N449);
not NOT1 (N1960, N1953);
or OR2 (N1961, N1951, N948);
xor XOR2 (N1962, N1952, N754);
nor NOR2 (N1963, N1959, N1914);
nand NAND2 (N1964, N1937, N301);
and AND2 (N1965, N1957, N1350);
buf BUF1 (N1966, N1963);
nand NAND3 (N1967, N1954, N1043, N932);
or OR4 (N1968, N1967, N502, N429, N1872);
nor NOR3 (N1969, N1968, N1809, N157);
xor XOR2 (N1970, N1969, N825);
not NOT1 (N1971, N1949);
not NOT1 (N1972, N1960);
or OR3 (N1973, N1971, N1752, N575);
and AND3 (N1974, N1972, N669, N1685);
or OR2 (N1975, N1958, N1206);
and AND3 (N1976, N1973, N533, N1012);
xor XOR2 (N1977, N1966, N727);
or OR2 (N1978, N1975, N8);
nor NOR4 (N1979, N1976, N963, N916, N22);
nand NAND3 (N1980, N1977, N1240, N1127);
or OR4 (N1981, N1962, N730, N1465, N1715);
buf BUF1 (N1982, N1970);
nor NOR3 (N1983, N1980, N1219, N1243);
or OR4 (N1984, N1961, N981, N1003, N287);
nand NAND2 (N1985, N1983, N1741);
not NOT1 (N1986, N1978);
and AND2 (N1987, N1986, N1855);
not NOT1 (N1988, N1979);
or OR3 (N1989, N1964, N19, N1593);
and AND4 (N1990, N1985, N974, N1336, N856);
nor NOR2 (N1991, N1974, N1714);
nand NAND3 (N1992, N1982, N1538, N635);
not NOT1 (N1993, N1989);
nor NOR4 (N1994, N1993, N1868, N997, N133);
or OR2 (N1995, N1965, N1021);
nor NOR2 (N1996, N1994, N197);
or OR2 (N1997, N1947, N249);
and AND2 (N1998, N1997, N717);
nor NOR3 (N1999, N1981, N1640, N211);
or OR3 (N2000, N1998, N1420, N1473);
nand NAND2 (N2001, N1996, N899);
xor XOR2 (N2002, N1990, N1957);
or OR3 (N2003, N1992, N1660, N720);
xor XOR2 (N2004, N1991, N379);
or OR2 (N2005, N2001, N1891);
buf BUF1 (N2006, N2003);
or OR4 (N2007, N1995, N100, N1876, N1122);
not NOT1 (N2008, N2004);
xor XOR2 (N2009, N2005, N1917);
and AND3 (N2010, N2007, N1513, N669);
not NOT1 (N2011, N2010);
nor NOR4 (N2012, N2002, N1267, N1368, N244);
xor XOR2 (N2013, N2012, N1280);
buf BUF1 (N2014, N1999);
not NOT1 (N2015, N2008);
buf BUF1 (N2016, N1988);
buf BUF1 (N2017, N2013);
or OR4 (N2018, N2011, N643, N141, N1254);
buf BUF1 (N2019, N1984);
xor XOR2 (N2020, N1987, N1316);
nand NAND2 (N2021, N2016, N1322);
or OR4 (N2022, N2019, N1112, N1504, N298);
xor XOR2 (N2023, N2009, N967);
nand NAND3 (N2024, N2014, N1530, N1286);
not NOT1 (N2025, N2021);
or OR2 (N2026, N2018, N558);
nor NOR4 (N2027, N2022, N1289, N2025, N255);
or OR3 (N2028, N1198, N1473, N1532);
not NOT1 (N2029, N2026);
and AND4 (N2030, N2015, N1313, N145, N614);
buf BUF1 (N2031, N2017);
xor XOR2 (N2032, N2031, N1372);
or OR4 (N2033, N2027, N1491, N1010, N525);
nor NOR4 (N2034, N2033, N619, N1396, N6);
xor XOR2 (N2035, N2006, N911);
xor XOR2 (N2036, N2035, N1956);
xor XOR2 (N2037, N2029, N1027);
nor NOR3 (N2038, N2032, N1236, N1516);
nor NOR2 (N2039, N2000, N1544);
or OR2 (N2040, N2037, N1608);
xor XOR2 (N2041, N2034, N607);
or OR3 (N2042, N2020, N1010, N1145);
xor XOR2 (N2043, N2039, N397);
or OR4 (N2044, N2030, N1830, N407, N1257);
nor NOR3 (N2045, N2036, N891, N1248);
nand NAND4 (N2046, N2040, N1981, N1384, N215);
and AND2 (N2047, N2038, N934);
or OR3 (N2048, N2043, N165, N1842);
xor XOR2 (N2049, N2042, N531);
nor NOR3 (N2050, N2047, N1246, N321);
and AND3 (N2051, N2045, N52, N1200);
xor XOR2 (N2052, N2049, N1460);
buf BUF1 (N2053, N2046);
xor XOR2 (N2054, N2053, N208);
xor XOR2 (N2055, N2041, N1303);
and AND3 (N2056, N2051, N237, N601);
nor NOR4 (N2057, N2028, N413, N136, N1377);
and AND4 (N2058, N2050, N689, N59, N330);
xor XOR2 (N2059, N2055, N513);
and AND4 (N2060, N2056, N1883, N1475, N2037);
and AND2 (N2061, N2044, N1182);
and AND2 (N2062, N2060, N2007);
xor XOR2 (N2063, N2061, N1418);
nor NOR2 (N2064, N2023, N1053);
xor XOR2 (N2065, N2054, N1222);
and AND4 (N2066, N2024, N1351, N69, N1816);
nor NOR2 (N2067, N2057, N466);
xor XOR2 (N2068, N2052, N225);
or OR4 (N2069, N2063, N655, N1002, N1582);
nand NAND2 (N2070, N2048, N1571);
not NOT1 (N2071, N2070);
buf BUF1 (N2072, N2069);
not NOT1 (N2073, N2072);
and AND3 (N2074, N2058, N1696, N760);
and AND2 (N2075, N2066, N362);
and AND4 (N2076, N2074, N512, N38, N562);
xor XOR2 (N2077, N2076, N224);
not NOT1 (N2078, N2065);
buf BUF1 (N2079, N2071);
nor NOR4 (N2080, N2077, N1359, N1332, N809);
xor XOR2 (N2081, N2075, N422);
xor XOR2 (N2082, N2064, N1110);
or OR3 (N2083, N2079, N120, N923);
buf BUF1 (N2084, N2083);
not NOT1 (N2085, N2062);
buf BUF1 (N2086, N2078);
and AND3 (N2087, N2068, N2069, N553);
or OR4 (N2088, N2067, N149, N516, N277);
not NOT1 (N2089, N2081);
xor XOR2 (N2090, N2087, N1420);
buf BUF1 (N2091, N2082);
nor NOR2 (N2092, N2059, N285);
and AND4 (N2093, N2088, N907, N1134, N1859);
nand NAND3 (N2094, N2090, N1339, N593);
not NOT1 (N2095, N2091);
and AND4 (N2096, N2089, N1557, N1019, N784);
nor NOR4 (N2097, N2092, N247, N980, N758);
buf BUF1 (N2098, N2084);
and AND3 (N2099, N2098, N416, N1561);
not NOT1 (N2100, N2073);
and AND4 (N2101, N2096, N851, N1780, N263);
or OR3 (N2102, N2093, N830, N1475);
not NOT1 (N2103, N2097);
not NOT1 (N2104, N2095);
nor NOR2 (N2105, N2080, N1327);
and AND2 (N2106, N2094, N158);
buf BUF1 (N2107, N2101);
or OR4 (N2108, N2086, N2000, N329, N1055);
nand NAND4 (N2109, N2105, N1285, N1900, N1540);
nor NOR2 (N2110, N2085, N1440);
and AND4 (N2111, N2110, N1378, N1410, N2010);
buf BUF1 (N2112, N2099);
nor NOR3 (N2113, N2102, N432, N603);
buf BUF1 (N2114, N2103);
not NOT1 (N2115, N2114);
xor XOR2 (N2116, N2111, N1062);
xor XOR2 (N2117, N2115, N1293);
buf BUF1 (N2118, N2112);
buf BUF1 (N2119, N2118);
xor XOR2 (N2120, N2108, N206);
and AND3 (N2121, N2113, N908, N1494);
xor XOR2 (N2122, N2109, N1371);
and AND4 (N2123, N2100, N2028, N484, N983);
and AND3 (N2124, N2121, N661, N488);
and AND3 (N2125, N2122, N21, N1904);
nor NOR4 (N2126, N2104, N1809, N974, N427);
and AND3 (N2127, N2107, N916, N1754);
nand NAND4 (N2128, N2123, N389, N1020, N1972);
nand NAND4 (N2129, N2127, N1994, N832, N542);
nand NAND3 (N2130, N2119, N579, N2090);
or OR4 (N2131, N2124, N991, N1922, N107);
xor XOR2 (N2132, N2125, N237);
nand NAND2 (N2133, N2120, N137);
and AND2 (N2134, N2106, N1491);
not NOT1 (N2135, N2131);
and AND2 (N2136, N2132, N688);
nand NAND4 (N2137, N2133, N1573, N91, N421);
xor XOR2 (N2138, N2126, N158);
xor XOR2 (N2139, N2136, N250);
or OR2 (N2140, N2134, N1019);
not NOT1 (N2141, N2129);
nand NAND4 (N2142, N2137, N2023, N1231, N197);
or OR4 (N2143, N2117, N1064, N163, N333);
and AND4 (N2144, N2143, N292, N898, N613);
or OR4 (N2145, N2135, N1366, N1005, N177);
not NOT1 (N2146, N2138);
xor XOR2 (N2147, N2139, N484);
xor XOR2 (N2148, N2130, N1675);
buf BUF1 (N2149, N2148);
nand NAND4 (N2150, N2140, N615, N1905, N865);
xor XOR2 (N2151, N2116, N1650);
or OR3 (N2152, N2151, N1137, N2087);
and AND4 (N2153, N2147, N509, N954, N425);
xor XOR2 (N2154, N2149, N1213);
and AND3 (N2155, N2144, N550, N942);
or OR4 (N2156, N2153, N1981, N630, N40);
and AND2 (N2157, N2146, N1231);
and AND3 (N2158, N2128, N2020, N1518);
buf BUF1 (N2159, N2157);
or OR4 (N2160, N2159, N1361, N735, N2112);
not NOT1 (N2161, N2154);
nand NAND4 (N2162, N2156, N1718, N1460, N1856);
nor NOR3 (N2163, N2152, N359, N1236);
xor XOR2 (N2164, N2161, N857);
nand NAND4 (N2165, N2164, N105, N891, N528);
not NOT1 (N2166, N2165);
nor NOR3 (N2167, N2158, N1481, N505);
xor XOR2 (N2168, N2145, N1157);
nand NAND4 (N2169, N2155, N1880, N275, N984);
nand NAND4 (N2170, N2150, N811, N2031, N588);
not NOT1 (N2171, N2167);
not NOT1 (N2172, N2142);
not NOT1 (N2173, N2172);
not NOT1 (N2174, N2173);
nor NOR2 (N2175, N2166, N2147);
xor XOR2 (N2176, N2162, N1238);
nor NOR2 (N2177, N2175, N1005);
xor XOR2 (N2178, N2171, N2002);
xor XOR2 (N2179, N2174, N849);
and AND3 (N2180, N2170, N401, N983);
and AND3 (N2181, N2177, N484, N700);
nor NOR3 (N2182, N2176, N839, N1183);
or OR4 (N2183, N2181, N1023, N572, N1861);
xor XOR2 (N2184, N2179, N1694);
and AND2 (N2185, N2180, N1465);
and AND2 (N2186, N2184, N482);
or OR4 (N2187, N2186, N2158, N1924, N1218);
or OR2 (N2188, N2160, N2181);
or OR3 (N2189, N2185, N1642, N2049);
and AND3 (N2190, N2163, N1199, N49);
not NOT1 (N2191, N2169);
or OR4 (N2192, N2141, N190, N1026, N1688);
buf BUF1 (N2193, N2192);
nand NAND3 (N2194, N2191, N235, N859);
buf BUF1 (N2195, N2189);
or OR2 (N2196, N2178, N419);
nand NAND4 (N2197, N2168, N307, N1404, N580);
not NOT1 (N2198, N2187);
nand NAND3 (N2199, N2194, N1469, N986);
and AND2 (N2200, N2190, N749);
nand NAND3 (N2201, N2199, N670, N851);
not NOT1 (N2202, N2193);
xor XOR2 (N2203, N2201, N984);
or OR3 (N2204, N2183, N2118, N217);
xor XOR2 (N2205, N2196, N1743);
not NOT1 (N2206, N2205);
not NOT1 (N2207, N2188);
or OR3 (N2208, N2200, N689, N2191);
buf BUF1 (N2209, N2182);
xor XOR2 (N2210, N2195, N879);
nor NOR4 (N2211, N2210, N463, N624, N586);
nor NOR2 (N2212, N2197, N1027);
nand NAND4 (N2213, N2202, N1949, N662, N1570);
nand NAND2 (N2214, N2198, N1653);
and AND3 (N2215, N2213, N1430, N48);
buf BUF1 (N2216, N2204);
and AND3 (N2217, N2209, N1222, N356);
buf BUF1 (N2218, N2215);
nor NOR3 (N2219, N2211, N439, N63);
and AND3 (N2220, N2216, N739, N1023);
nand NAND2 (N2221, N2217, N97);
and AND3 (N2222, N2208, N820, N2039);
nor NOR3 (N2223, N2212, N1023, N990);
not NOT1 (N2224, N2207);
nand NAND3 (N2225, N2224, N1485, N396);
buf BUF1 (N2226, N2206);
xor XOR2 (N2227, N2220, N687);
and AND2 (N2228, N2219, N857);
buf BUF1 (N2229, N2222);
not NOT1 (N2230, N2228);
nor NOR2 (N2231, N2221, N638);
or OR2 (N2232, N2230, N2099);
nor NOR4 (N2233, N2225, N1913, N1848, N1811);
and AND3 (N2234, N2218, N2107, N613);
buf BUF1 (N2235, N2223);
xor XOR2 (N2236, N2227, N606);
xor XOR2 (N2237, N2236, N2123);
or OR4 (N2238, N2231, N1523, N1849, N1126);
not NOT1 (N2239, N2226);
or OR4 (N2240, N2214, N1683, N1785, N632);
xor XOR2 (N2241, N2233, N1787);
nor NOR2 (N2242, N2238, N410);
xor XOR2 (N2243, N2237, N1031);
not NOT1 (N2244, N2232);
and AND4 (N2245, N2240, N471, N1856, N1141);
buf BUF1 (N2246, N2234);
nor NOR4 (N2247, N2243, N1132, N2035, N1093);
nand NAND4 (N2248, N2229, N1262, N1894, N646);
nand NAND4 (N2249, N2239, N1262, N1354, N253);
buf BUF1 (N2250, N2241);
or OR2 (N2251, N2247, N1957);
nand NAND3 (N2252, N2249, N1079, N1622);
and AND4 (N2253, N2244, N718, N756, N475);
xor XOR2 (N2254, N2242, N1100);
xor XOR2 (N2255, N2251, N67);
nand NAND2 (N2256, N2254, N1403);
or OR4 (N2257, N2250, N1797, N471, N1830);
or OR3 (N2258, N2203, N1321, N211);
buf BUF1 (N2259, N2257);
nand NAND4 (N2260, N2245, N1034, N744, N1929);
not NOT1 (N2261, N2246);
nor NOR4 (N2262, N2235, N1205, N118, N1019);
or OR4 (N2263, N2256, N1433, N2042, N2061);
or OR3 (N2264, N2263, N639, N525);
not NOT1 (N2265, N2261);
nor NOR3 (N2266, N2255, N1476, N1388);
nor NOR3 (N2267, N2264, N875, N521);
xor XOR2 (N2268, N2253, N1433);
nor NOR2 (N2269, N2267, N1685);
not NOT1 (N2270, N2260);
and AND3 (N2271, N2259, N233, N1856);
buf BUF1 (N2272, N2265);
and AND4 (N2273, N2268, N1050, N339, N1951);
nand NAND3 (N2274, N2272, N1722, N996);
buf BUF1 (N2275, N2262);
not NOT1 (N2276, N2271);
or OR4 (N2277, N2274, N1571, N1136, N1997);
xor XOR2 (N2278, N2248, N1789);
xor XOR2 (N2279, N2273, N3);
nand NAND4 (N2280, N2270, N1173, N528, N2148);
and AND2 (N2281, N2277, N1984);
buf BUF1 (N2282, N2275);
and AND3 (N2283, N2269, N1090, N2191);
and AND3 (N2284, N2278, N1382, N2117);
and AND2 (N2285, N2279, N1907);
xor XOR2 (N2286, N2258, N503);
nand NAND4 (N2287, N2285, N1323, N1662, N719);
buf BUF1 (N2288, N2266);
nand NAND3 (N2289, N2288, N1794, N301);
not NOT1 (N2290, N2281);
not NOT1 (N2291, N2286);
nor NOR2 (N2292, N2252, N2146);
and AND3 (N2293, N2282, N445, N1113);
nand NAND2 (N2294, N2283, N1211);
buf BUF1 (N2295, N2291);
not NOT1 (N2296, N2294);
xor XOR2 (N2297, N2287, N1300);
nand NAND2 (N2298, N2296, N1845);
nand NAND4 (N2299, N2289, N632, N1368, N1478);
buf BUF1 (N2300, N2295);
buf BUF1 (N2301, N2298);
not NOT1 (N2302, N2293);
buf BUF1 (N2303, N2300);
xor XOR2 (N2304, N2280, N1598);
or OR4 (N2305, N2292, N1357, N119, N211);
buf BUF1 (N2306, N2302);
or OR4 (N2307, N2290, N1789, N1505, N70);
xor XOR2 (N2308, N2306, N1482);
nor NOR2 (N2309, N2303, N1954);
and AND4 (N2310, N2304, N1153, N1458, N1123);
buf BUF1 (N2311, N2310);
buf BUF1 (N2312, N2299);
and AND4 (N2313, N2308, N1555, N487, N1888);
and AND3 (N2314, N2305, N1812, N1666);
and AND2 (N2315, N2313, N1926);
nand NAND3 (N2316, N2297, N299, N1285);
not NOT1 (N2317, N2315);
nand NAND4 (N2318, N2314, N690, N1957, N1807);
xor XOR2 (N2319, N2284, N566);
and AND4 (N2320, N2316, N1886, N1906, N206);
nor NOR2 (N2321, N2312, N531);
xor XOR2 (N2322, N2311, N941);
or OR2 (N2323, N2318, N48);
buf BUF1 (N2324, N2321);
xor XOR2 (N2325, N2309, N57);
nand NAND4 (N2326, N2323, N374, N1178, N695);
not NOT1 (N2327, N2320);
nor NOR4 (N2328, N2327, N1947, N1669, N867);
xor XOR2 (N2329, N2328, N2025);
not NOT1 (N2330, N2325);
not NOT1 (N2331, N2324);
nand NAND3 (N2332, N2330, N2030, N1864);
or OR3 (N2333, N2319, N437, N316);
or OR4 (N2334, N2326, N2258, N871, N870);
and AND2 (N2335, N2332, N782);
nor NOR2 (N2336, N2331, N1523);
buf BUF1 (N2337, N2307);
buf BUF1 (N2338, N2337);
buf BUF1 (N2339, N2333);
or OR3 (N2340, N2322, N1932, N559);
nor NOR4 (N2341, N2301, N59, N1920, N110);
nand NAND4 (N2342, N2334, N536, N264, N1988);
not NOT1 (N2343, N2317);
xor XOR2 (N2344, N2329, N1323);
nor NOR4 (N2345, N2343, N1132, N386, N1717);
buf BUF1 (N2346, N2345);
xor XOR2 (N2347, N2339, N2132);
xor XOR2 (N2348, N2336, N4);
nor NOR3 (N2349, N2342, N2192, N1791);
xor XOR2 (N2350, N2347, N1500);
not NOT1 (N2351, N2349);
nor NOR2 (N2352, N2348, N2117);
not NOT1 (N2353, N2340);
nand NAND4 (N2354, N2353, N316, N521, N1475);
xor XOR2 (N2355, N2354, N484);
nor NOR2 (N2356, N2351, N774);
nand NAND4 (N2357, N2346, N683, N1127, N1630);
nand NAND4 (N2358, N2357, N1843, N980, N2209);
and AND4 (N2359, N2356, N1101, N1098, N1779);
not NOT1 (N2360, N2344);
nand NAND3 (N2361, N2338, N1144, N329);
and AND3 (N2362, N2358, N2074, N420);
not NOT1 (N2363, N2352);
nand NAND4 (N2364, N2350, N1507, N1511, N2090);
and AND2 (N2365, N2359, N1376);
xor XOR2 (N2366, N2355, N2242);
and AND4 (N2367, N2335, N601, N1319, N1762);
not NOT1 (N2368, N2360);
not NOT1 (N2369, N2365);
nor NOR3 (N2370, N2363, N642, N1669);
not NOT1 (N2371, N2368);
buf BUF1 (N2372, N2364);
and AND3 (N2373, N2369, N1784, N769);
and AND3 (N2374, N2371, N1720, N166);
and AND4 (N2375, N2341, N218, N1318, N661);
or OR3 (N2376, N2375, N1107, N1607);
or OR3 (N2377, N2370, N624, N1809);
xor XOR2 (N2378, N2372, N2205);
or OR4 (N2379, N2374, N1416, N404, N188);
xor XOR2 (N2380, N2379, N1193);
nand NAND3 (N2381, N2361, N1823, N441);
nand NAND2 (N2382, N2367, N2003);
nor NOR4 (N2383, N2377, N1677, N786, N1544);
buf BUF1 (N2384, N2362);
nor NOR3 (N2385, N2381, N351, N557);
buf BUF1 (N2386, N2382);
nor NOR4 (N2387, N2383, N1899, N1759, N519);
xor XOR2 (N2388, N2378, N1477);
xor XOR2 (N2389, N2366, N1175);
or OR3 (N2390, N2387, N689, N1004);
nor NOR3 (N2391, N2386, N37, N2345);
xor XOR2 (N2392, N2391, N11);
nor NOR2 (N2393, N2376, N190);
nand NAND4 (N2394, N2390, N622, N327, N1255);
buf BUF1 (N2395, N2394);
buf BUF1 (N2396, N2393);
and AND2 (N2397, N2392, N342);
or OR3 (N2398, N2397, N596, N1124);
buf BUF1 (N2399, N2276);
nor NOR3 (N2400, N2389, N1758, N256);
and AND4 (N2401, N2399, N651, N1286, N480);
buf BUF1 (N2402, N2380);
buf BUF1 (N2403, N2373);
buf BUF1 (N2404, N2396);
nand NAND2 (N2405, N2402, N76);
xor XOR2 (N2406, N2395, N998);
and AND4 (N2407, N2388, N2328, N1297, N1392);
xor XOR2 (N2408, N2404, N2394);
buf BUF1 (N2409, N2398);
or OR3 (N2410, N2403, N546, N2013);
nor NOR2 (N2411, N2384, N1929);
xor XOR2 (N2412, N2406, N1915);
buf BUF1 (N2413, N2385);
buf BUF1 (N2414, N2409);
buf BUF1 (N2415, N2413);
buf BUF1 (N2416, N2411);
or OR3 (N2417, N2405, N255, N2366);
and AND4 (N2418, N2415, N1611, N570, N507);
not NOT1 (N2419, N2412);
buf BUF1 (N2420, N2414);
xor XOR2 (N2421, N2416, N1167);
and AND4 (N2422, N2420, N944, N648, N2285);
nor NOR2 (N2423, N2407, N1492);
nand NAND4 (N2424, N2417, N154, N2158, N1471);
nor NOR4 (N2425, N2410, N1674, N2384, N294);
xor XOR2 (N2426, N2424, N1016);
or OR4 (N2427, N2421, N1316, N98, N2061);
nand NAND3 (N2428, N2408, N2279, N2110);
buf BUF1 (N2429, N2401);
or OR2 (N2430, N2426, N1221);
nand NAND4 (N2431, N2427, N2180, N1036, N1811);
or OR3 (N2432, N2428, N1760, N360);
buf BUF1 (N2433, N2429);
buf BUF1 (N2434, N2423);
nor NOR4 (N2435, N2431, N1176, N1532, N1);
buf BUF1 (N2436, N2422);
nand NAND2 (N2437, N2434, N2375);
xor XOR2 (N2438, N2435, N1312);
nor NOR2 (N2439, N2436, N1717);
nand NAND2 (N2440, N2425, N635);
xor XOR2 (N2441, N2430, N173);
nor NOR3 (N2442, N2438, N2430, N661);
not NOT1 (N2443, N2441);
or OR3 (N2444, N2432, N2124, N38);
nor NOR4 (N2445, N2418, N679, N1369, N1899);
nand NAND2 (N2446, N2439, N56);
xor XOR2 (N2447, N2443, N2145);
xor XOR2 (N2448, N2400, N36);
and AND3 (N2449, N2447, N1149, N1593);
not NOT1 (N2450, N2449);
buf BUF1 (N2451, N2442);
and AND2 (N2452, N2419, N2014);
buf BUF1 (N2453, N2446);
nand NAND4 (N2454, N2437, N139, N2264, N496);
nand NAND3 (N2455, N2448, N2373, N1473);
and AND2 (N2456, N2433, N2350);
not NOT1 (N2457, N2455);
nor NOR3 (N2458, N2453, N1589, N1660);
not NOT1 (N2459, N2451);
nor NOR4 (N2460, N2454, N668, N1592, N332);
and AND4 (N2461, N2440, N220, N1946, N2250);
xor XOR2 (N2462, N2452, N2078);
not NOT1 (N2463, N2450);
nand NAND3 (N2464, N2463, N1601, N1866);
nand NAND4 (N2465, N2459, N2084, N2329, N1830);
not NOT1 (N2466, N2462);
nand NAND3 (N2467, N2461, N1616, N2286);
nand NAND4 (N2468, N2467, N2116, N1212, N329);
buf BUF1 (N2469, N2445);
and AND2 (N2470, N2468, N195);
nand NAND2 (N2471, N2465, N1284);
or OR2 (N2472, N2471, N37);
xor XOR2 (N2473, N2457, N2466);
xor XOR2 (N2474, N2459, N854);
nand NAND3 (N2475, N2444, N1852, N59);
not NOT1 (N2476, N2458);
nand NAND3 (N2477, N2470, N918, N631);
nand NAND4 (N2478, N2476, N1149, N2133, N2241);
and AND2 (N2479, N2478, N2211);
not NOT1 (N2480, N2464);
or OR4 (N2481, N2456, N559, N2398, N512);
or OR4 (N2482, N2480, N1505, N1475, N1966);
and AND3 (N2483, N2460, N1959, N539);
and AND4 (N2484, N2474, N1474, N1121, N126);
buf BUF1 (N2485, N2484);
nor NOR3 (N2486, N2481, N1906, N2099);
nand NAND4 (N2487, N2482, N835, N2111, N1499);
or OR3 (N2488, N2487, N523, N613);
nand NAND2 (N2489, N2477, N307);
nor NOR2 (N2490, N2469, N321);
xor XOR2 (N2491, N2475, N2141);
nor NOR2 (N2492, N2490, N1026);
nand NAND4 (N2493, N2485, N500, N8, N756);
or OR2 (N2494, N2483, N2240);
nor NOR2 (N2495, N2473, N988);
nor NOR4 (N2496, N2472, N1373, N2456, N1798);
nand NAND2 (N2497, N2491, N1042);
nor NOR2 (N2498, N2489, N1990);
not NOT1 (N2499, N2492);
nor NOR3 (N2500, N2498, N50, N2298);
not NOT1 (N2501, N2494);
not NOT1 (N2502, N2488);
and AND3 (N2503, N2499, N980, N2412);
not NOT1 (N2504, N2486);
nand NAND3 (N2505, N2479, N198, N1462);
nand NAND4 (N2506, N2495, N2058, N2409, N1588);
buf BUF1 (N2507, N2496);
or OR4 (N2508, N2503, N2341, N1159, N1375);
and AND2 (N2509, N2507, N552);
or OR2 (N2510, N2502, N535);
or OR4 (N2511, N2501, N1509, N43, N1007);
xor XOR2 (N2512, N2505, N2437);
xor XOR2 (N2513, N2508, N880);
or OR4 (N2514, N2510, N654, N298, N1017);
xor XOR2 (N2515, N2509, N1294);
not NOT1 (N2516, N2497);
xor XOR2 (N2517, N2516, N2429);
nor NOR3 (N2518, N2511, N229, N1537);
not NOT1 (N2519, N2504);
nor NOR3 (N2520, N2518, N308, N1805);
buf BUF1 (N2521, N2520);
or OR2 (N2522, N2519, N1945);
or OR2 (N2523, N2515, N271);
nand NAND2 (N2524, N2506, N900);
not NOT1 (N2525, N2513);
or OR3 (N2526, N2525, N931, N1130);
nor NOR2 (N2527, N2493, N1075);
xor XOR2 (N2528, N2527, N1729);
or OR3 (N2529, N2526, N1859, N583);
xor XOR2 (N2530, N2524, N2328);
not NOT1 (N2531, N2512);
not NOT1 (N2532, N2530);
nand NAND2 (N2533, N2517, N534);
and AND2 (N2534, N2500, N1276);
and AND4 (N2535, N2532, N2221, N1644, N942);
xor XOR2 (N2536, N2531, N2005);
nor NOR4 (N2537, N2521, N1425, N216, N175);
and AND2 (N2538, N2536, N1190);
xor XOR2 (N2539, N2514, N1950);
not NOT1 (N2540, N2534);
nand NAND3 (N2541, N2538, N1411, N637);
and AND2 (N2542, N2528, N1390);
xor XOR2 (N2543, N2535, N1147);
not NOT1 (N2544, N2529);
not NOT1 (N2545, N2533);
and AND2 (N2546, N2523, N916);
buf BUF1 (N2547, N2546);
nor NOR2 (N2548, N2541, N877);
nand NAND2 (N2549, N2539, N1937);
buf BUF1 (N2550, N2522);
and AND3 (N2551, N2543, N1969, N1883);
nand NAND4 (N2552, N2548, N724, N1106, N952);
and AND3 (N2553, N2544, N299, N1287);
and AND4 (N2554, N2540, N2469, N274, N797);
xor XOR2 (N2555, N2545, N529);
not NOT1 (N2556, N2547);
not NOT1 (N2557, N2550);
nand NAND4 (N2558, N2551, N527, N2266, N1472);
and AND2 (N2559, N2542, N1281);
buf BUF1 (N2560, N2556);
not NOT1 (N2561, N2560);
not NOT1 (N2562, N2553);
not NOT1 (N2563, N2558);
nand NAND4 (N2564, N2563, N1888, N1332, N2356);
buf BUF1 (N2565, N2537);
nor NOR2 (N2566, N2559, N2297);
nand NAND2 (N2567, N2561, N2412);
and AND3 (N2568, N2565, N1938, N1066);
and AND4 (N2569, N2554, N2008, N937, N1352);
buf BUF1 (N2570, N2549);
buf BUF1 (N2571, N2569);
or OR4 (N2572, N2564, N1277, N1327, N851);
nand NAND4 (N2573, N2571, N380, N2121, N1448);
not NOT1 (N2574, N2567);
xor XOR2 (N2575, N2555, N373);
not NOT1 (N2576, N2574);
nor NOR4 (N2577, N2566, N1264, N1702, N1839);
nand NAND3 (N2578, N2562, N523, N582);
xor XOR2 (N2579, N2552, N1270);
xor XOR2 (N2580, N2578, N923);
buf BUF1 (N2581, N2570);
nor NOR3 (N2582, N2557, N2321, N2341);
nand NAND2 (N2583, N2573, N2246);
buf BUF1 (N2584, N2575);
xor XOR2 (N2585, N2581, N1018);
and AND4 (N2586, N2577, N419, N1629, N2121);
nor NOR3 (N2587, N2582, N951, N1615);
nor NOR2 (N2588, N2583, N649);
buf BUF1 (N2589, N2587);
nand NAND3 (N2590, N2586, N1710, N1652);
xor XOR2 (N2591, N2585, N394);
nor NOR2 (N2592, N2591, N2387);
nor NOR3 (N2593, N2589, N1078, N1385);
and AND4 (N2594, N2590, N168, N406, N1660);
nand NAND2 (N2595, N2568, N2577);
or OR3 (N2596, N2576, N1042, N651);
nand NAND2 (N2597, N2579, N234);
xor XOR2 (N2598, N2595, N1717);
buf BUF1 (N2599, N2572);
xor XOR2 (N2600, N2599, N1473);
xor XOR2 (N2601, N2584, N1148);
xor XOR2 (N2602, N2580, N2279);
and AND2 (N2603, N2600, N2024);
nor NOR3 (N2604, N2597, N15, N909);
not NOT1 (N2605, N2593);
buf BUF1 (N2606, N2604);
nand NAND3 (N2607, N2602, N2112, N881);
nand NAND4 (N2608, N2605, N1700, N50, N533);
nand NAND3 (N2609, N2608, N2453, N1480);
nand NAND2 (N2610, N2588, N1784);
nor NOR4 (N2611, N2592, N1311, N890, N1991);
xor XOR2 (N2612, N2607, N184);
nand NAND4 (N2613, N2612, N1534, N186, N1330);
or OR2 (N2614, N2598, N331);
nor NOR2 (N2615, N2596, N2285);
xor XOR2 (N2616, N2603, N1436);
buf BUF1 (N2617, N2615);
nor NOR2 (N2618, N2611, N1082);
and AND3 (N2619, N2594, N742, N1147);
nand NAND2 (N2620, N2619, N1379);
nor NOR2 (N2621, N2617, N1400);
or OR2 (N2622, N2620, N13);
nand NAND4 (N2623, N2609, N2478, N366, N2519);
or OR3 (N2624, N2623, N1938, N996);
nand NAND2 (N2625, N2624, N863);
buf BUF1 (N2626, N2613);
nand NAND2 (N2627, N2621, N955);
and AND3 (N2628, N2616, N1747, N688);
nor NOR2 (N2629, N2618, N1075);
buf BUF1 (N2630, N2628);
nor NOR3 (N2631, N2627, N938, N1275);
buf BUF1 (N2632, N2629);
buf BUF1 (N2633, N2625);
not NOT1 (N2634, N2626);
xor XOR2 (N2635, N2601, N1197);
xor XOR2 (N2636, N2633, N428);
xor XOR2 (N2637, N2635, N1526);
nor NOR4 (N2638, N2637, N2229, N2257, N381);
xor XOR2 (N2639, N2614, N38);
not NOT1 (N2640, N2631);
nand NAND3 (N2641, N2639, N1308, N1787);
xor XOR2 (N2642, N2641, N2563);
and AND4 (N2643, N2634, N925, N302, N1636);
nor NOR4 (N2644, N2632, N493, N693, N2191);
not NOT1 (N2645, N2644);
nand NAND2 (N2646, N2630, N983);
xor XOR2 (N2647, N2622, N301);
not NOT1 (N2648, N2636);
or OR2 (N2649, N2642, N456);
nand NAND3 (N2650, N2645, N582, N172);
xor XOR2 (N2651, N2646, N2159);
nor NOR2 (N2652, N2606, N1974);
xor XOR2 (N2653, N2649, N1147);
not NOT1 (N2654, N2643);
nor NOR3 (N2655, N2640, N1984, N2584);
nand NAND4 (N2656, N2651, N2557, N1015, N1277);
nand NAND4 (N2657, N2647, N244, N2626, N822);
nand NAND4 (N2658, N2653, N2233, N2593, N262);
xor XOR2 (N2659, N2658, N1005);
or OR3 (N2660, N2656, N2466, N1671);
buf BUF1 (N2661, N2659);
not NOT1 (N2662, N2655);
buf BUF1 (N2663, N2657);
or OR4 (N2664, N2661, N2351, N1833, N2523);
xor XOR2 (N2665, N2652, N2513);
and AND3 (N2666, N2654, N955, N2130);
and AND2 (N2667, N2663, N558);
xor XOR2 (N2668, N2650, N920);
or OR2 (N2669, N2665, N880);
or OR3 (N2670, N2669, N769, N7);
nor NOR2 (N2671, N2666, N639);
or OR4 (N2672, N2662, N448, N224, N1294);
nor NOR2 (N2673, N2668, N1665);
or OR3 (N2674, N2671, N1120, N148);
or OR2 (N2675, N2610, N1460);
not NOT1 (N2676, N2660);
not NOT1 (N2677, N2664);
nand NAND4 (N2678, N2648, N1108, N772, N2543);
and AND4 (N2679, N2678, N1107, N1206, N1644);
xor XOR2 (N2680, N2674, N1155);
or OR3 (N2681, N2667, N1099, N145);
xor XOR2 (N2682, N2672, N1542);
and AND3 (N2683, N2675, N2650, N305);
or OR4 (N2684, N2673, N2490, N1670, N1341);
nor NOR4 (N2685, N2676, N721, N370, N886);
or OR3 (N2686, N2684, N1232, N1048);
not NOT1 (N2687, N2683);
and AND3 (N2688, N2680, N599, N6);
not NOT1 (N2689, N2682);
or OR2 (N2690, N2689, N1257);
nand NAND2 (N2691, N2687, N865);
and AND3 (N2692, N2690, N2583, N1083);
or OR3 (N2693, N2670, N2316, N1072);
xor XOR2 (N2694, N2692, N1216);
nor NOR3 (N2695, N2693, N626, N1191);
or OR2 (N2696, N2688, N2071);
nand NAND4 (N2697, N2694, N138, N417, N2001);
nand NAND3 (N2698, N2685, N508, N2487);
nand NAND3 (N2699, N2695, N66, N345);
nor NOR3 (N2700, N2696, N1945, N1302);
and AND3 (N2701, N2681, N884, N1352);
or OR4 (N2702, N2677, N1117, N1954, N2493);
buf BUF1 (N2703, N2691);
xor XOR2 (N2704, N2638, N1191);
nand NAND2 (N2705, N2699, N1033);
buf BUF1 (N2706, N2704);
xor XOR2 (N2707, N2705, N2501);
and AND2 (N2708, N2700, N1856);
and AND3 (N2709, N2679, N617, N197);
and AND4 (N2710, N2697, N704, N2195, N399);
xor XOR2 (N2711, N2703, N790);
or OR3 (N2712, N2686, N2574, N1945);
and AND2 (N2713, N2711, N2529);
or OR4 (N2714, N2708, N857, N1117, N283);
nand NAND2 (N2715, N2712, N2200);
nor NOR4 (N2716, N2707, N1799, N1187, N1255);
nor NOR4 (N2717, N2698, N75, N2466, N1230);
and AND4 (N2718, N2715, N565, N336, N1653);
not NOT1 (N2719, N2710);
or OR2 (N2720, N2713, N1358);
and AND4 (N2721, N2709, N1488, N46, N1265);
nor NOR3 (N2722, N2706, N762, N1034);
nand NAND3 (N2723, N2719, N2425, N2048);
and AND2 (N2724, N2714, N2000);
nand NAND2 (N2725, N2720, N861);
buf BUF1 (N2726, N2701);
nand NAND3 (N2727, N2725, N347, N1313);
nor NOR4 (N2728, N2717, N2348, N1092, N385);
nor NOR3 (N2729, N2721, N1074, N2409);
nand NAND3 (N2730, N2722, N2064, N2394);
and AND3 (N2731, N2716, N680, N2403);
xor XOR2 (N2732, N2724, N1551);
not NOT1 (N2733, N2732);
xor XOR2 (N2734, N2726, N2722);
nor NOR3 (N2735, N2727, N674, N526);
nor NOR4 (N2736, N2718, N880, N959, N583);
buf BUF1 (N2737, N2702);
nor NOR3 (N2738, N2733, N2736, N104);
not NOT1 (N2739, N71);
or OR2 (N2740, N2728, N494);
or OR3 (N2741, N2737, N2145, N1231);
buf BUF1 (N2742, N2740);
buf BUF1 (N2743, N2729);
or OR4 (N2744, N2741, N2648, N695, N465);
nand NAND2 (N2745, N2738, N2321);
nor NOR2 (N2746, N2735, N49);
not NOT1 (N2747, N2723);
not NOT1 (N2748, N2745);
xor XOR2 (N2749, N2744, N940);
or OR4 (N2750, N2742, N1143, N2374, N32);
xor XOR2 (N2751, N2748, N1467);
or OR4 (N2752, N2743, N1460, N208, N225);
not NOT1 (N2753, N2734);
and AND3 (N2754, N2752, N1089, N1808);
not NOT1 (N2755, N2747);
xor XOR2 (N2756, N2746, N1656);
or OR3 (N2757, N2756, N837, N221);
nand NAND3 (N2758, N2731, N950, N70);
nor NOR4 (N2759, N2753, N2436, N1617, N2415);
nor NOR3 (N2760, N2751, N2460, N1769);
nand NAND2 (N2761, N2759, N1503);
or OR3 (N2762, N2755, N2233, N1799);
buf BUF1 (N2763, N2749);
nor NOR2 (N2764, N2763, N2211);
buf BUF1 (N2765, N2762);
nand NAND4 (N2766, N2739, N113, N1840, N573);
nor NOR2 (N2767, N2730, N197);
or OR2 (N2768, N2767, N1330);
nor NOR4 (N2769, N2765, N1060, N496, N1494);
xor XOR2 (N2770, N2754, N2571);
not NOT1 (N2771, N2769);
or OR3 (N2772, N2771, N533, N229);
xor XOR2 (N2773, N2761, N1168);
and AND4 (N2774, N2770, N1638, N1040, N1434);
nand NAND2 (N2775, N2760, N487);
and AND4 (N2776, N2764, N884, N1916, N1402);
not NOT1 (N2777, N2766);
nor NOR4 (N2778, N2777, N2659, N2288, N2252);
or OR3 (N2779, N2775, N2749, N182);
xor XOR2 (N2780, N2750, N976);
and AND3 (N2781, N2758, N1804, N52);
nand NAND2 (N2782, N2779, N930);
or OR2 (N2783, N2773, N135);
nor NOR2 (N2784, N2783, N533);
nand NAND3 (N2785, N2781, N1933, N1336);
nand NAND2 (N2786, N2772, N1045);
and AND4 (N2787, N2774, N1222, N1411, N706);
not NOT1 (N2788, N2780);
and AND2 (N2789, N2776, N1693);
nor NOR4 (N2790, N2757, N253, N477, N13);
xor XOR2 (N2791, N2768, N1218);
xor XOR2 (N2792, N2785, N1060);
nor NOR3 (N2793, N2790, N2742, N1792);
and AND4 (N2794, N2784, N1280, N1841, N1080);
or OR2 (N2795, N2794, N1866);
xor XOR2 (N2796, N2795, N1035);
not NOT1 (N2797, N2782);
or OR3 (N2798, N2797, N1817, N986);
nor NOR3 (N2799, N2778, N639, N1607);
or OR3 (N2800, N2791, N1686, N2133);
xor XOR2 (N2801, N2789, N1718);
not NOT1 (N2802, N2788);
buf BUF1 (N2803, N2798);
nand NAND4 (N2804, N2786, N1240, N381, N1847);
not NOT1 (N2805, N2804);
and AND4 (N2806, N2802, N1628, N2245, N2441);
or OR2 (N2807, N2792, N2554);
buf BUF1 (N2808, N2805);
or OR2 (N2809, N2787, N1435);
and AND3 (N2810, N2806, N1473, N497);
not NOT1 (N2811, N2810);
xor XOR2 (N2812, N2800, N339);
or OR2 (N2813, N2808, N344);
xor XOR2 (N2814, N2813, N2140);
nand NAND2 (N2815, N2812, N2144);
or OR3 (N2816, N2796, N1801, N2067);
and AND2 (N2817, N2803, N1782);
nor NOR3 (N2818, N2799, N1103, N2076);
and AND4 (N2819, N2807, N603, N2593, N1055);
not NOT1 (N2820, N2809);
and AND2 (N2821, N2814, N96);
not NOT1 (N2822, N2821);
xor XOR2 (N2823, N2819, N1147);
nand NAND3 (N2824, N2801, N2008, N1392);
not NOT1 (N2825, N2815);
buf BUF1 (N2826, N2820);
buf BUF1 (N2827, N2818);
nand NAND3 (N2828, N2825, N2392, N1087);
buf BUF1 (N2829, N2823);
buf BUF1 (N2830, N2816);
or OR3 (N2831, N2828, N1221, N92);
not NOT1 (N2832, N2824);
not NOT1 (N2833, N2817);
not NOT1 (N2834, N2811);
or OR2 (N2835, N2822, N2064);
nand NAND4 (N2836, N2832, N2620, N1585, N196);
nor NOR3 (N2837, N2831, N322, N2220);
buf BUF1 (N2838, N2830);
xor XOR2 (N2839, N2837, N1551);
nor NOR4 (N2840, N2835, N1100, N770, N2044);
buf BUF1 (N2841, N2839);
or OR2 (N2842, N2829, N738);
or OR4 (N2843, N2838, N2375, N1622, N2407);
and AND2 (N2844, N2836, N476);
or OR4 (N2845, N2834, N1038, N741, N59);
nand NAND3 (N2846, N2833, N1656, N2530);
not NOT1 (N2847, N2793);
nor NOR3 (N2848, N2827, N2227, N774);
nor NOR4 (N2849, N2845, N149, N1872, N1900);
nand NAND4 (N2850, N2844, N2641, N1405, N2150);
and AND4 (N2851, N2842, N2022, N117, N852);
nor NOR2 (N2852, N2849, N2330);
not NOT1 (N2853, N2850);
nor NOR4 (N2854, N2847, N1584, N1703, N177);
or OR3 (N2855, N2848, N2674, N107);
nand NAND2 (N2856, N2851, N989);
and AND4 (N2857, N2841, N824, N907, N1010);
and AND4 (N2858, N2846, N2397, N2269, N1750);
or OR3 (N2859, N2856, N1923, N1044);
not NOT1 (N2860, N2859);
buf BUF1 (N2861, N2854);
nor NOR2 (N2862, N2861, N206);
nor NOR3 (N2863, N2857, N170, N1972);
buf BUF1 (N2864, N2860);
or OR3 (N2865, N2862, N637, N2064);
and AND3 (N2866, N2863, N73, N261);
nor NOR2 (N2867, N2865, N576);
and AND3 (N2868, N2826, N310, N1691);
and AND4 (N2869, N2867, N1269, N1439, N1455);
xor XOR2 (N2870, N2864, N515);
and AND4 (N2871, N2840, N909, N2712, N666);
and AND3 (N2872, N2870, N353, N2035);
buf BUF1 (N2873, N2855);
not NOT1 (N2874, N2871);
nor NOR2 (N2875, N2873, N2505);
xor XOR2 (N2876, N2866, N2070);
buf BUF1 (N2877, N2874);
and AND4 (N2878, N2872, N2760, N2423, N2358);
xor XOR2 (N2879, N2853, N1548);
and AND3 (N2880, N2843, N1300, N1426);
or OR4 (N2881, N2875, N2098, N1021, N1920);
buf BUF1 (N2882, N2858);
or OR4 (N2883, N2878, N107, N519, N1098);
or OR3 (N2884, N2852, N1941, N2416);
and AND4 (N2885, N2876, N2647, N693, N2273);
and AND2 (N2886, N2868, N2610);
nor NOR4 (N2887, N2885, N2325, N186, N1190);
nor NOR2 (N2888, N2869, N2769);
and AND2 (N2889, N2877, N494);
nor NOR3 (N2890, N2883, N1637, N1783);
and AND2 (N2891, N2889, N65);
and AND2 (N2892, N2882, N2606);
xor XOR2 (N2893, N2881, N1495);
not NOT1 (N2894, N2884);
not NOT1 (N2895, N2886);
nand NAND2 (N2896, N2879, N2554);
buf BUF1 (N2897, N2895);
or OR4 (N2898, N2896, N2342, N1238, N704);
xor XOR2 (N2899, N2898, N1894);
nand NAND3 (N2900, N2893, N2274, N1955);
nor NOR3 (N2901, N2900, N503, N1967);
nor NOR2 (N2902, N2891, N44);
nor NOR2 (N2903, N2894, N1221);
nor NOR4 (N2904, N2887, N238, N1063, N1121);
and AND2 (N2905, N2880, N2071);
nor NOR4 (N2906, N2904, N1345, N356, N1929);
nand NAND3 (N2907, N2888, N48, N936);
buf BUF1 (N2908, N2899);
buf BUF1 (N2909, N2903);
or OR4 (N2910, N2907, N2234, N30, N1561);
and AND4 (N2911, N2892, N1142, N1753, N1698);
xor XOR2 (N2912, N2909, N1858);
or OR4 (N2913, N2905, N459, N1429, N2813);
and AND4 (N2914, N2911, N1003, N1, N2100);
nand NAND3 (N2915, N2890, N690, N367);
xor XOR2 (N2916, N2897, N642);
nand NAND2 (N2917, N2901, N1884);
buf BUF1 (N2918, N2910);
or OR3 (N2919, N2912, N97, N2613);
nand NAND2 (N2920, N2906, N2562);
not NOT1 (N2921, N2918);
or OR3 (N2922, N2920, N992, N934);
and AND2 (N2923, N2915, N2366);
buf BUF1 (N2924, N2908);
not NOT1 (N2925, N2917);
buf BUF1 (N2926, N2916);
xor XOR2 (N2927, N2926, N1811);
and AND3 (N2928, N2923, N2766, N167);
not NOT1 (N2929, N2921);
nor NOR4 (N2930, N2927, N283, N306, N1937);
not NOT1 (N2931, N2928);
nor NOR3 (N2932, N2931, N2179, N146);
xor XOR2 (N2933, N2924, N2930);
nor NOR2 (N2934, N2874, N293);
nand NAND2 (N2935, N2929, N1140);
or OR4 (N2936, N2935, N2389, N437, N1498);
nand NAND4 (N2937, N2936, N121, N32, N1386);
buf BUF1 (N2938, N2919);
buf BUF1 (N2939, N2934);
and AND2 (N2940, N2922, N2601);
not NOT1 (N2941, N2925);
buf BUF1 (N2942, N2932);
buf BUF1 (N2943, N2939);
nor NOR2 (N2944, N2933, N2278);
not NOT1 (N2945, N2913);
or OR3 (N2946, N2902, N2259, N1119);
nor NOR2 (N2947, N2943, N470);
xor XOR2 (N2948, N2937, N1141);
nor NOR2 (N2949, N2938, N43);
not NOT1 (N2950, N2948);
xor XOR2 (N2951, N2942, N2650);
or OR2 (N2952, N2950, N1466);
buf BUF1 (N2953, N2951);
and AND2 (N2954, N2944, N537);
or OR2 (N2955, N2946, N404);
nand NAND3 (N2956, N2947, N1628, N1110);
or OR4 (N2957, N2941, N2170, N2025, N2541);
or OR4 (N2958, N2945, N1963, N2298, N2484);
xor XOR2 (N2959, N2914, N2017);
xor XOR2 (N2960, N2953, N2897);
buf BUF1 (N2961, N2955);
not NOT1 (N2962, N2952);
xor XOR2 (N2963, N2954, N1192);
xor XOR2 (N2964, N2962, N532);
xor XOR2 (N2965, N2958, N1448);
nand NAND2 (N2966, N2965, N798);
nand NAND3 (N2967, N2949, N290, N1051);
nand NAND2 (N2968, N2960, N2940);
nand NAND2 (N2969, N1691, N2091);
and AND2 (N2970, N2969, N2331);
nor NOR3 (N2971, N2961, N2593, N1084);
nand NAND2 (N2972, N2971, N2937);
not NOT1 (N2973, N2957);
and AND4 (N2974, N2972, N1813, N550, N2140);
not NOT1 (N2975, N2973);
buf BUF1 (N2976, N2966);
or OR2 (N2977, N2968, N2149);
or OR3 (N2978, N2970, N864, N2732);
or OR2 (N2979, N2977, N1182);
xor XOR2 (N2980, N2975, N257);
nor NOR4 (N2981, N2978, N1862, N11, N1613);
not NOT1 (N2982, N2967);
buf BUF1 (N2983, N2979);
xor XOR2 (N2984, N2963, N1411);
not NOT1 (N2985, N2983);
xor XOR2 (N2986, N2959, N412);
or OR3 (N2987, N2964, N2482, N1942);
nor NOR2 (N2988, N2956, N1814);
xor XOR2 (N2989, N2980, N1325);
buf BUF1 (N2990, N2982);
xor XOR2 (N2991, N2987, N2833);
and AND2 (N2992, N2981, N173);
nor NOR2 (N2993, N2990, N1384);
nor NOR3 (N2994, N2989, N1346, N929);
or OR3 (N2995, N2992, N900, N101);
nand NAND3 (N2996, N2991, N1555, N235);
and AND4 (N2997, N2993, N1117, N898, N777);
xor XOR2 (N2998, N2974, N1900);
nand NAND4 (N2999, N2995, N722, N447, N1367);
nand NAND4 (N3000, N2998, N1943, N2768, N1016);
nor NOR4 (N3001, N2988, N2934, N1009, N2092);
buf BUF1 (N3002, N3001);
and AND2 (N3003, N3000, N1641);
and AND2 (N3004, N2999, N2329);
not NOT1 (N3005, N3002);
buf BUF1 (N3006, N2986);
nor NOR2 (N3007, N2976, N197);
nand NAND4 (N3008, N3005, N999, N633, N2249);
buf BUF1 (N3009, N3003);
xor XOR2 (N3010, N3006, N2731);
or OR4 (N3011, N2984, N2155, N236, N155);
and AND3 (N3012, N3011, N905, N1763);
buf BUF1 (N3013, N3004);
xor XOR2 (N3014, N3008, N1412);
or OR2 (N3015, N3007, N355);
xor XOR2 (N3016, N2996, N2037);
or OR2 (N3017, N3009, N1769);
buf BUF1 (N3018, N3010);
buf BUF1 (N3019, N3017);
and AND2 (N3020, N3014, N922);
xor XOR2 (N3021, N3016, N1263);
nor NOR2 (N3022, N2985, N409);
or OR3 (N3023, N3022, N1018, N788);
nand NAND2 (N3024, N2997, N2573);
and AND4 (N3025, N3013, N786, N21, N48);
buf BUF1 (N3026, N3015);
or OR3 (N3027, N3023, N982, N280);
or OR4 (N3028, N3018, N382, N600, N51);
not NOT1 (N3029, N2994);
xor XOR2 (N3030, N3012, N2142);
nor NOR3 (N3031, N3019, N468, N2463);
nor NOR4 (N3032, N3024, N2577, N2330, N191);
not NOT1 (N3033, N3020);
and AND2 (N3034, N3027, N2379);
or OR2 (N3035, N3029, N1988);
and AND4 (N3036, N3035, N2693, N1023, N2463);
nand NAND2 (N3037, N3030, N583);
not NOT1 (N3038, N3032);
xor XOR2 (N3039, N3026, N2160);
nor NOR2 (N3040, N3033, N1539);
xor XOR2 (N3041, N3040, N1497);
not NOT1 (N3042, N3034);
and AND3 (N3043, N3039, N2787, N2962);
and AND4 (N3044, N3031, N1971, N2107, N2018);
not NOT1 (N3045, N3041);
xor XOR2 (N3046, N3038, N2010);
and AND2 (N3047, N3042, N2347);
or OR3 (N3048, N3028, N110, N955);
buf BUF1 (N3049, N3044);
xor XOR2 (N3050, N3046, N192);
or OR2 (N3051, N3036, N3003);
nand NAND4 (N3052, N3043, N2195, N720, N1607);
not NOT1 (N3053, N3052);
and AND4 (N3054, N3048, N220, N2670, N2447);
or OR3 (N3055, N3049, N3048, N2959);
or OR3 (N3056, N3054, N806, N2816);
nor NOR4 (N3057, N3051, N442, N2550, N367);
and AND4 (N3058, N3045, N1437, N467, N219);
and AND2 (N3059, N3025, N162);
nand NAND4 (N3060, N3057, N2575, N1176, N1492);
not NOT1 (N3061, N3037);
buf BUF1 (N3062, N3021);
nand NAND2 (N3063, N3056, N732);
and AND3 (N3064, N3060, N996, N2463);
buf BUF1 (N3065, N3058);
buf BUF1 (N3066, N3059);
nor NOR2 (N3067, N3062, N291);
not NOT1 (N3068, N3066);
xor XOR2 (N3069, N3063, N672);
nand NAND2 (N3070, N3065, N3057);
not NOT1 (N3071, N3061);
nand NAND4 (N3072, N3050, N2453, N3012, N1073);
and AND4 (N3073, N3072, N2403, N2548, N516);
nand NAND4 (N3074, N3067, N1748, N2716, N2784);
nor NOR2 (N3075, N3070, N694);
nor NOR4 (N3076, N3064, N2243, N349, N927);
and AND2 (N3077, N3075, N2794);
buf BUF1 (N3078, N3074);
or OR4 (N3079, N3053, N2445, N2107, N2019);
xor XOR2 (N3080, N3076, N2910);
nand NAND2 (N3081, N3080, N1904);
xor XOR2 (N3082, N3071, N1883);
buf BUF1 (N3083, N3079);
nor NOR2 (N3084, N3069, N862);
or OR3 (N3085, N3077, N1284, N2418);
buf BUF1 (N3086, N3068);
not NOT1 (N3087, N3055);
or OR2 (N3088, N3082, N2776);
buf BUF1 (N3089, N3087);
xor XOR2 (N3090, N3083, N2493);
or OR4 (N3091, N3085, N2771, N649, N2366);
not NOT1 (N3092, N3091);
nand NAND4 (N3093, N3047, N590, N2960, N2116);
and AND2 (N3094, N3092, N1678);
and AND4 (N3095, N3073, N618, N351, N1518);
not NOT1 (N3096, N3078);
xor XOR2 (N3097, N3090, N1598);
xor XOR2 (N3098, N3093, N2584);
not NOT1 (N3099, N3098);
nand NAND2 (N3100, N3088, N290);
nand NAND4 (N3101, N3099, N2643, N2268, N740);
nand NAND2 (N3102, N3095, N916);
xor XOR2 (N3103, N3100, N346);
xor XOR2 (N3104, N3101, N164);
buf BUF1 (N3105, N3104);
and AND4 (N3106, N3102, N2003, N655, N1353);
not NOT1 (N3107, N3081);
or OR2 (N3108, N3107, N2364);
or OR2 (N3109, N3108, N1077);
xor XOR2 (N3110, N3096, N1613);
buf BUF1 (N3111, N3094);
nand NAND4 (N3112, N3084, N156, N1781, N3049);
nand NAND4 (N3113, N3106, N203, N1694, N2226);
or OR2 (N3114, N3112, N2537);
xor XOR2 (N3115, N3110, N1659);
and AND4 (N3116, N3103, N409, N1840, N1772);
nor NOR3 (N3117, N3114, N2785, N2878);
and AND3 (N3118, N3116, N3046, N2422);
or OR4 (N3119, N3113, N1582, N1162, N1347);
not NOT1 (N3120, N3097);
nand NAND2 (N3121, N3086, N1255);
nand NAND4 (N3122, N3118, N22, N1968, N892);
xor XOR2 (N3123, N3111, N2749);
nor NOR2 (N3124, N3120, N3039);
and AND4 (N3125, N3124, N2816, N215, N66);
nand NAND3 (N3126, N3125, N1654, N60);
xor XOR2 (N3127, N3105, N2811);
nor NOR2 (N3128, N3119, N1104);
not NOT1 (N3129, N3109);
xor XOR2 (N3130, N3089, N2268);
not NOT1 (N3131, N3123);
buf BUF1 (N3132, N3130);
and AND2 (N3133, N3132, N1794);
or OR3 (N3134, N3133, N1924, N2918);
or OR4 (N3135, N3131, N2526, N2003, N1395);
and AND2 (N3136, N3122, N430);
nand NAND2 (N3137, N3127, N1264);
buf BUF1 (N3138, N3117);
buf BUF1 (N3139, N3126);
nor NOR4 (N3140, N3121, N1065, N2998, N2791);
buf BUF1 (N3141, N3115);
nor NOR4 (N3142, N3138, N2368, N2560, N666);
or OR3 (N3143, N3136, N906, N1436);
nand NAND3 (N3144, N3139, N1639, N2409);
nand NAND3 (N3145, N3135, N656, N2751);
buf BUF1 (N3146, N3142);
nor NOR2 (N3147, N3141, N161);
not NOT1 (N3148, N3140);
buf BUF1 (N3149, N3137);
xor XOR2 (N3150, N3128, N1145);
or OR2 (N3151, N3149, N2399);
xor XOR2 (N3152, N3151, N2307);
xor XOR2 (N3153, N3145, N641);
nor NOR2 (N3154, N3129, N1609);
and AND3 (N3155, N3144, N3147, N1758);
not NOT1 (N3156, N226);
buf BUF1 (N3157, N3146);
nor NOR3 (N3158, N3153, N881, N1123);
xor XOR2 (N3159, N3158, N1175);
and AND2 (N3160, N3152, N44);
or OR4 (N3161, N3148, N2832, N182, N1621);
not NOT1 (N3162, N3156);
buf BUF1 (N3163, N3154);
not NOT1 (N3164, N3155);
not NOT1 (N3165, N3160);
nor NOR2 (N3166, N3163, N7);
xor XOR2 (N3167, N3134, N216);
xor XOR2 (N3168, N3165, N1668);
nor NOR2 (N3169, N3157, N1401);
nor NOR4 (N3170, N3162, N407, N1569, N2218);
nor NOR4 (N3171, N3159, N2615, N1262, N2570);
and AND4 (N3172, N3168, N29, N1169, N2344);
not NOT1 (N3173, N3172);
or OR3 (N3174, N3143, N1410, N2447);
or OR4 (N3175, N3170, N1720, N695, N963);
or OR3 (N3176, N3169, N957, N1587);
nand NAND4 (N3177, N3161, N916, N2932, N1343);
and AND4 (N3178, N3164, N2834, N2141, N2719);
nor NOR2 (N3179, N3166, N2378);
nand NAND2 (N3180, N3177, N3099);
xor XOR2 (N3181, N3176, N1214);
or OR4 (N3182, N3178, N162, N3080, N2191);
nor NOR3 (N3183, N3167, N2888, N3067);
buf BUF1 (N3184, N3175);
and AND4 (N3185, N3171, N1554, N600, N1121);
nor NOR4 (N3186, N3180, N2714, N1799, N386);
xor XOR2 (N3187, N3181, N1089);
nand NAND3 (N3188, N3184, N2961, N204);
and AND4 (N3189, N3185, N1261, N181, N1583);
nand NAND2 (N3190, N3183, N160);
not NOT1 (N3191, N3189);
xor XOR2 (N3192, N3150, N290);
not NOT1 (N3193, N3174);
nor NOR2 (N3194, N3173, N2472);
or OR4 (N3195, N3194, N1607, N1513, N653);
and AND4 (N3196, N3179, N901, N2314, N2662);
or OR2 (N3197, N3187, N587);
buf BUF1 (N3198, N3197);
and AND4 (N3199, N3190, N1986, N101, N1775);
and AND4 (N3200, N3195, N1209, N494, N2708);
nor NOR4 (N3201, N3182, N1626, N884, N1107);
nor NOR3 (N3202, N3186, N2663, N1683);
buf BUF1 (N3203, N3200);
not NOT1 (N3204, N3192);
not NOT1 (N3205, N3199);
buf BUF1 (N3206, N3204);
not NOT1 (N3207, N3191);
not NOT1 (N3208, N3196);
and AND2 (N3209, N3201, N2325);
nand NAND3 (N3210, N3207, N2711, N1514);
nor NOR4 (N3211, N3188, N995, N783, N3056);
nand NAND4 (N3212, N3193, N242, N194, N2459);
not NOT1 (N3213, N3203);
buf BUF1 (N3214, N3208);
and AND3 (N3215, N3210, N2381, N55);
and AND3 (N3216, N3205, N1009, N2936);
buf BUF1 (N3217, N3211);
not NOT1 (N3218, N3206);
and AND4 (N3219, N3214, N3048, N2447, N1604);
nor NOR4 (N3220, N3215, N2536, N1132, N2745);
nor NOR4 (N3221, N3220, N3125, N799, N2606);
not NOT1 (N3222, N3217);
or OR4 (N3223, N3216, N198, N1211, N1549);
and AND3 (N3224, N3218, N172, N1865);
not NOT1 (N3225, N3224);
not NOT1 (N3226, N3212);
buf BUF1 (N3227, N3223);
nor NOR4 (N3228, N3226, N2411, N1289, N1733);
and AND2 (N3229, N3198, N207);
not NOT1 (N3230, N3202);
buf BUF1 (N3231, N3230);
and AND3 (N3232, N3222, N1859, N1210);
not NOT1 (N3233, N3231);
xor XOR2 (N3234, N3213, N630);
or OR2 (N3235, N3229, N3129);
nand NAND4 (N3236, N3228, N3086, N2978, N1862);
and AND4 (N3237, N3233, N2502, N456, N2137);
xor XOR2 (N3238, N3234, N3195);
nand NAND2 (N3239, N3225, N1101);
not NOT1 (N3240, N3239);
and AND3 (N3241, N3232, N3127, N1986);
not NOT1 (N3242, N3241);
and AND3 (N3243, N3236, N1024, N1058);
buf BUF1 (N3244, N3240);
nand NAND3 (N3245, N3227, N956, N1257);
nand NAND2 (N3246, N3245, N1756);
buf BUF1 (N3247, N3237);
and AND3 (N3248, N3238, N2888, N540);
and AND3 (N3249, N3248, N174, N2580);
not NOT1 (N3250, N3235);
and AND4 (N3251, N3219, N1042, N115, N1555);
not NOT1 (N3252, N3242);
not NOT1 (N3253, N3250);
not NOT1 (N3254, N3243);
xor XOR2 (N3255, N3221, N1860);
nor NOR4 (N3256, N3246, N2814, N364, N2201);
or OR3 (N3257, N3209, N1388, N3174);
and AND2 (N3258, N3254, N2969);
and AND3 (N3259, N3247, N2419, N347);
nor NOR4 (N3260, N3259, N3157, N2062, N2656);
nand NAND3 (N3261, N3260, N2707, N2591);
or OR3 (N3262, N3256, N63, N1939);
and AND2 (N3263, N3255, N3249);
nand NAND3 (N3264, N2137, N98, N1356);
and AND3 (N3265, N3252, N2283, N2305);
and AND3 (N3266, N3244, N145, N2634);
buf BUF1 (N3267, N3263);
nor NOR4 (N3268, N3265, N1468, N2524, N1981);
or OR4 (N3269, N3258, N2735, N1680, N2913);
or OR2 (N3270, N3264, N1257);
or OR4 (N3271, N3269, N2810, N748, N2932);
not NOT1 (N3272, N3270);
buf BUF1 (N3273, N3261);
and AND2 (N3274, N3268, N3133);
not NOT1 (N3275, N3251);
xor XOR2 (N3276, N3271, N1305);
nor NOR2 (N3277, N3275, N1849);
and AND4 (N3278, N3276, N1913, N3233, N694);
nor NOR4 (N3279, N3277, N2909, N1374, N46);
buf BUF1 (N3280, N3279);
and AND3 (N3281, N3272, N2917, N1437);
not NOT1 (N3282, N3257);
xor XOR2 (N3283, N3253, N2109);
buf BUF1 (N3284, N3266);
and AND4 (N3285, N3273, N941, N1444, N614);
and AND3 (N3286, N3274, N2690, N828);
or OR4 (N3287, N3280, N461, N1604, N1806);
nor NOR3 (N3288, N3285, N324, N535);
and AND4 (N3289, N3288, N594, N1837, N2595);
or OR4 (N3290, N3278, N1456, N2019, N2736);
nor NOR4 (N3291, N3284, N2351, N1625, N1229);
nor NOR3 (N3292, N3289, N421, N2193);
or OR2 (N3293, N3287, N2986);
nand NAND3 (N3294, N3292, N115, N1467);
nor NOR2 (N3295, N3267, N2206);
not NOT1 (N3296, N3286);
xor XOR2 (N3297, N3282, N1782);
and AND2 (N3298, N3291, N1148);
and AND4 (N3299, N3293, N1121, N3084, N2809);
not NOT1 (N3300, N3298);
xor XOR2 (N3301, N3296, N502);
nor NOR2 (N3302, N3283, N2542);
or OR3 (N3303, N3301, N1748, N1949);
and AND3 (N3304, N3300, N944, N2526);
and AND2 (N3305, N3295, N930);
buf BUF1 (N3306, N3290);
nand NAND3 (N3307, N3306, N1645, N1252);
not NOT1 (N3308, N3303);
and AND4 (N3309, N3305, N624, N1160, N951);
nor NOR4 (N3310, N3299, N2172, N3020, N758);
and AND2 (N3311, N3308, N1939);
not NOT1 (N3312, N3311);
or OR3 (N3313, N3281, N947, N2258);
xor XOR2 (N3314, N3302, N1733);
not NOT1 (N3315, N3314);
xor XOR2 (N3316, N3262, N2689);
buf BUF1 (N3317, N3297);
nand NAND4 (N3318, N3307, N579, N1907, N3044);
nand NAND4 (N3319, N3309, N3091, N2238, N1213);
not NOT1 (N3320, N3304);
or OR4 (N3321, N3312, N1525, N2086, N2923);
buf BUF1 (N3322, N3315);
buf BUF1 (N3323, N3321);
or OR4 (N3324, N3318, N1682, N256, N611);
nand NAND2 (N3325, N3317, N1328);
and AND4 (N3326, N3319, N436, N2523, N1048);
xor XOR2 (N3327, N3322, N2357);
and AND4 (N3328, N3313, N748, N1815, N3159);
nand NAND2 (N3329, N3326, N2752);
buf BUF1 (N3330, N3327);
nor NOR2 (N3331, N3324, N1628);
nand NAND2 (N3332, N3328, N876);
nor NOR3 (N3333, N3331, N1564, N955);
nor NOR3 (N3334, N3294, N2487, N3164);
or OR3 (N3335, N3323, N2248, N90);
buf BUF1 (N3336, N3329);
nor NOR3 (N3337, N3333, N2216, N855);
and AND4 (N3338, N3320, N2829, N2489, N1744);
nand NAND2 (N3339, N3338, N2236);
and AND2 (N3340, N3325, N2170);
xor XOR2 (N3341, N3332, N3075);
buf BUF1 (N3342, N3316);
not NOT1 (N3343, N3310);
or OR2 (N3344, N3342, N1485);
nor NOR4 (N3345, N3340, N286, N2002, N1784);
not NOT1 (N3346, N3345);
or OR2 (N3347, N3336, N1318);
nor NOR4 (N3348, N3343, N414, N2927, N1913);
and AND4 (N3349, N3339, N2100, N2305, N305);
xor XOR2 (N3350, N3348, N1109);
xor XOR2 (N3351, N3347, N2776);
not NOT1 (N3352, N3341);
not NOT1 (N3353, N3334);
xor XOR2 (N3354, N3330, N487);
buf BUF1 (N3355, N3352);
buf BUF1 (N3356, N3351);
not NOT1 (N3357, N3346);
not NOT1 (N3358, N3354);
not NOT1 (N3359, N3356);
nor NOR4 (N3360, N3344, N1832, N1613, N2270);
or OR2 (N3361, N3359, N2998);
or OR4 (N3362, N3335, N3278, N209, N2757);
nor NOR3 (N3363, N3337, N3216, N1317);
buf BUF1 (N3364, N3362);
xor XOR2 (N3365, N3353, N3217);
nand NAND2 (N3366, N3364, N3168);
not NOT1 (N3367, N3350);
nand NAND4 (N3368, N3367, N864, N1099, N3260);
not NOT1 (N3369, N3357);
nand NAND4 (N3370, N3355, N1925, N601, N1822);
and AND4 (N3371, N3366, N2988, N1977, N684);
nand NAND4 (N3372, N3358, N3184, N590, N1560);
and AND3 (N3373, N3371, N3129, N2574);
nor NOR3 (N3374, N3368, N398, N1844);
xor XOR2 (N3375, N3363, N1094);
not NOT1 (N3376, N3372);
nand NAND3 (N3377, N3365, N3146, N1648);
nor NOR3 (N3378, N3374, N1098, N2732);
xor XOR2 (N3379, N3370, N1749);
not NOT1 (N3380, N3349);
xor XOR2 (N3381, N3361, N3284);
nand NAND2 (N3382, N3376, N1359);
nor NOR2 (N3383, N3379, N198);
nand NAND4 (N3384, N3373, N2101, N2949, N156);
nor NOR2 (N3385, N3381, N1957);
or OR2 (N3386, N3375, N580);
xor XOR2 (N3387, N3382, N1991);
xor XOR2 (N3388, N3385, N2237);
buf BUF1 (N3389, N3377);
not NOT1 (N3390, N3378);
nand NAND2 (N3391, N3369, N1745);
nor NOR4 (N3392, N3386, N1835, N2122, N340);
nor NOR4 (N3393, N3389, N2080, N1961, N2954);
nand NAND2 (N3394, N3384, N2754);
nand NAND4 (N3395, N3360, N2719, N1110, N2766);
nand NAND2 (N3396, N3390, N3118);
xor XOR2 (N3397, N3387, N2489);
nor NOR4 (N3398, N3388, N1113, N309, N2627);
buf BUF1 (N3399, N3395);
not NOT1 (N3400, N3391);
and AND2 (N3401, N3393, N2572);
buf BUF1 (N3402, N3394);
buf BUF1 (N3403, N3396);
nor NOR2 (N3404, N3392, N1819);
not NOT1 (N3405, N3401);
not NOT1 (N3406, N3400);
nor NOR2 (N3407, N3402, N1013);
nand NAND4 (N3408, N3397, N1231, N2966, N739);
buf BUF1 (N3409, N3380);
nand NAND2 (N3410, N3383, N3125);
xor XOR2 (N3411, N3408, N1318);
not NOT1 (N3412, N3403);
nand NAND4 (N3413, N3404, N1719, N1344, N414);
nand NAND4 (N3414, N3405, N2527, N377, N1887);
buf BUF1 (N3415, N3399);
and AND3 (N3416, N3407, N2687, N1215);
not NOT1 (N3417, N3409);
or OR2 (N3418, N3412, N2756);
xor XOR2 (N3419, N3406, N911);
and AND3 (N3420, N3417, N742, N804);
not NOT1 (N3421, N3414);
nand NAND4 (N3422, N3419, N671, N688, N1868);
buf BUF1 (N3423, N3398);
buf BUF1 (N3424, N3413);
or OR2 (N3425, N3416, N624);
buf BUF1 (N3426, N3420);
or OR2 (N3427, N3411, N2959);
buf BUF1 (N3428, N3424);
not NOT1 (N3429, N3425);
nor NOR3 (N3430, N3415, N440, N69);
or OR2 (N3431, N3421, N43);
or OR4 (N3432, N3418, N2197, N3051, N3272);
buf BUF1 (N3433, N3427);
or OR3 (N3434, N3431, N3112, N1545);
buf BUF1 (N3435, N3422);
nor NOR3 (N3436, N3434, N1105, N642);
buf BUF1 (N3437, N3430);
and AND4 (N3438, N3432, N10, N2195, N1386);
not NOT1 (N3439, N3410);
nand NAND3 (N3440, N3436, N1297, N2523);
nor NOR3 (N3441, N3440, N1403, N159);
nand NAND4 (N3442, N3437, N3419, N1915, N1059);
or OR3 (N3443, N3426, N765, N378);
and AND4 (N3444, N3429, N573, N295, N799);
xor XOR2 (N3445, N3439, N3280);
nand NAND3 (N3446, N3423, N461, N1480);
not NOT1 (N3447, N3435);
and AND4 (N3448, N3443, N2485, N1930, N1808);
not NOT1 (N3449, N3433);
nand NAND4 (N3450, N3441, N231, N1256, N763);
nand NAND3 (N3451, N3450, N2704, N359);
buf BUF1 (N3452, N3451);
buf BUF1 (N3453, N3445);
nand NAND3 (N3454, N3444, N2953, N3107);
xor XOR2 (N3455, N3446, N253);
xor XOR2 (N3456, N3438, N529);
and AND3 (N3457, N3455, N1197, N1668);
buf BUF1 (N3458, N3452);
xor XOR2 (N3459, N3449, N1317);
buf BUF1 (N3460, N3448);
and AND4 (N3461, N3459, N62, N2666, N1532);
and AND4 (N3462, N3458, N2445, N1157, N1690);
nor NOR2 (N3463, N3457, N844);
not NOT1 (N3464, N3456);
nand NAND3 (N3465, N3447, N1817, N637);
buf BUF1 (N3466, N3463);
nand NAND4 (N3467, N3442, N585, N2452, N2671);
nand NAND4 (N3468, N3465, N245, N3270, N951);
nor NOR4 (N3469, N3453, N817, N3112, N1220);
nor NOR3 (N3470, N3460, N2706, N837);
or OR2 (N3471, N3466, N2735);
or OR4 (N3472, N3428, N2173, N616, N228);
or OR4 (N3473, N3461, N1113, N415, N1614);
xor XOR2 (N3474, N3471, N514);
nor NOR3 (N3475, N3468, N2710, N192);
nand NAND3 (N3476, N3472, N380, N2870);
buf BUF1 (N3477, N3474);
xor XOR2 (N3478, N3475, N1703);
not NOT1 (N3479, N3470);
or OR4 (N3480, N3473, N1317, N2661, N1315);
nor NOR4 (N3481, N3478, N1671, N2610, N2955);
xor XOR2 (N3482, N3469, N41);
not NOT1 (N3483, N3462);
xor XOR2 (N3484, N3481, N3198);
not NOT1 (N3485, N3464);
or OR4 (N3486, N3477, N1647, N1461, N2036);
buf BUF1 (N3487, N3454);
buf BUF1 (N3488, N3486);
buf BUF1 (N3489, N3488);
nor NOR4 (N3490, N3476, N3292, N2915, N1613);
not NOT1 (N3491, N3490);
not NOT1 (N3492, N3480);
nor NOR3 (N3493, N3485, N335, N2718);
not NOT1 (N3494, N3479);
not NOT1 (N3495, N3467);
and AND2 (N3496, N3484, N2199);
nor NOR2 (N3497, N3496, N1130);
xor XOR2 (N3498, N3489, N1103);
or OR2 (N3499, N3498, N427);
nand NAND3 (N3500, N3495, N2496, N3394);
xor XOR2 (N3501, N3499, N1892);
and AND2 (N3502, N3501, N2498);
nand NAND4 (N3503, N3502, N3491, N1144, N3476);
buf BUF1 (N3504, N2625);
nor NOR3 (N3505, N3493, N2984, N792);
and AND3 (N3506, N3504, N2933, N711);
or OR4 (N3507, N3500, N728, N2404, N1263);
and AND3 (N3508, N3483, N3093, N2114);
buf BUF1 (N3509, N3505);
buf BUF1 (N3510, N3487);
and AND3 (N3511, N3503, N1993, N3409);
buf BUF1 (N3512, N3511);
not NOT1 (N3513, N3506);
nand NAND4 (N3514, N3509, N2540, N1634, N1723);
xor XOR2 (N3515, N3492, N324);
or OR3 (N3516, N3513, N1251, N420);
nor NOR3 (N3517, N3494, N560, N138);
or OR4 (N3518, N3516, N2437, N2060, N90);
or OR2 (N3519, N3497, N315);
xor XOR2 (N3520, N3519, N1085);
or OR3 (N3521, N3515, N725, N2080);
buf BUF1 (N3522, N3512);
nand NAND2 (N3523, N3521, N3321);
and AND2 (N3524, N3518, N1060);
buf BUF1 (N3525, N3482);
buf BUF1 (N3526, N3517);
not NOT1 (N3527, N3514);
xor XOR2 (N3528, N3522, N11);
or OR4 (N3529, N3523, N676, N3236, N1677);
nand NAND3 (N3530, N3529, N521, N124);
nand NAND3 (N3531, N3507, N2205, N226);
nand NAND4 (N3532, N3527, N2607, N2947, N893);
nand NAND4 (N3533, N3530, N1581, N2294, N3086);
and AND3 (N3534, N3533, N3226, N169);
and AND2 (N3535, N3520, N677);
buf BUF1 (N3536, N3528);
buf BUF1 (N3537, N3510);
or OR3 (N3538, N3532, N633, N755);
nor NOR2 (N3539, N3531, N2670);
and AND2 (N3540, N3537, N1443);
or OR4 (N3541, N3508, N2448, N1528, N2136);
xor XOR2 (N3542, N3541, N2484);
nand NAND4 (N3543, N3534, N530, N902, N3374);
or OR2 (N3544, N3542, N1481);
not NOT1 (N3545, N3526);
nand NAND2 (N3546, N3544, N2659);
and AND4 (N3547, N3540, N831, N1195, N1619);
xor XOR2 (N3548, N3536, N1805);
nand NAND2 (N3549, N3535, N2723);
xor XOR2 (N3550, N3525, N2037);
nor NOR4 (N3551, N3524, N3369, N457, N152);
nor NOR4 (N3552, N3543, N1801, N2523, N2792);
or OR3 (N3553, N3538, N3546, N1251);
nor NOR2 (N3554, N316, N1334);
xor XOR2 (N3555, N3550, N2173);
and AND3 (N3556, N3554, N590, N888);
nand NAND4 (N3557, N3555, N2423, N264, N1101);
nor NOR4 (N3558, N3548, N3112, N3382, N2933);
not NOT1 (N3559, N3545);
buf BUF1 (N3560, N3547);
buf BUF1 (N3561, N3539);
xor XOR2 (N3562, N3552, N261);
not NOT1 (N3563, N3560);
nand NAND4 (N3564, N3553, N2298, N1457, N3149);
xor XOR2 (N3565, N3558, N2559);
nor NOR4 (N3566, N3561, N1665, N1321, N2259);
not NOT1 (N3567, N3559);
and AND4 (N3568, N3565, N1439, N2765, N723);
nand NAND3 (N3569, N3551, N142, N1465);
nand NAND2 (N3570, N3569, N2914);
and AND3 (N3571, N3570, N1218, N803);
nor NOR4 (N3572, N3549, N812, N2426, N1213);
nor NOR2 (N3573, N3571, N2012);
nor NOR3 (N3574, N3563, N1952, N2932);
nand NAND4 (N3575, N3573, N3528, N1343, N3517);
and AND2 (N3576, N3564, N2563);
and AND3 (N3577, N3562, N3476, N2054);
not NOT1 (N3578, N3567);
nor NOR3 (N3579, N3566, N1605, N2669);
nor NOR3 (N3580, N3556, N178, N469);
and AND3 (N3581, N3579, N335, N2003);
xor XOR2 (N3582, N3557, N319);
not NOT1 (N3583, N3582);
or OR4 (N3584, N3581, N596, N2101, N2236);
nor NOR2 (N3585, N3572, N2508);
buf BUF1 (N3586, N3583);
nor NOR2 (N3587, N3574, N3317);
nor NOR3 (N3588, N3577, N582, N1395);
and AND3 (N3589, N3568, N518, N1775);
xor XOR2 (N3590, N3589, N819);
and AND2 (N3591, N3578, N266);
xor XOR2 (N3592, N3580, N2060);
buf BUF1 (N3593, N3586);
not NOT1 (N3594, N3585);
not NOT1 (N3595, N3593);
or OR4 (N3596, N3575, N1427, N1167, N1262);
xor XOR2 (N3597, N3590, N1737);
not NOT1 (N3598, N3594);
not NOT1 (N3599, N3584);
not NOT1 (N3600, N3587);
or OR2 (N3601, N3576, N1703);
nor NOR4 (N3602, N3597, N2579, N1399, N1748);
and AND4 (N3603, N3595, N168, N1446, N2135);
not NOT1 (N3604, N3592);
or OR4 (N3605, N3591, N2314, N2643, N529);
not NOT1 (N3606, N3604);
nor NOR4 (N3607, N3599, N3417, N1034, N469);
or OR2 (N3608, N3596, N528);
nand NAND3 (N3609, N3600, N2429, N3069);
nor NOR3 (N3610, N3608, N28, N1892);
not NOT1 (N3611, N3609);
nor NOR2 (N3612, N3611, N78);
and AND3 (N3613, N3606, N1914, N250);
or OR3 (N3614, N3602, N2640, N722);
and AND3 (N3615, N3613, N3443, N185);
nor NOR4 (N3616, N3610, N177, N2691, N1962);
nor NOR2 (N3617, N3615, N1905);
buf BUF1 (N3618, N3588);
xor XOR2 (N3619, N3598, N2677);
not NOT1 (N3620, N3619);
nor NOR3 (N3621, N3607, N329, N1551);
xor XOR2 (N3622, N3601, N2523);
not NOT1 (N3623, N3616);
nor NOR2 (N3624, N3614, N3374);
buf BUF1 (N3625, N3605);
or OR3 (N3626, N3622, N1164, N436);
xor XOR2 (N3627, N3603, N3132);
xor XOR2 (N3628, N3626, N3481);
buf BUF1 (N3629, N3612);
buf BUF1 (N3630, N3618);
xor XOR2 (N3631, N3625, N2167);
buf BUF1 (N3632, N3624);
nand NAND3 (N3633, N3629, N3194, N2042);
buf BUF1 (N3634, N3632);
buf BUF1 (N3635, N3621);
not NOT1 (N3636, N3633);
buf BUF1 (N3637, N3631);
buf BUF1 (N3638, N3635);
buf BUF1 (N3639, N3638);
nor NOR4 (N3640, N3639, N2586, N943, N2972);
and AND4 (N3641, N3636, N832, N2835, N1782);
or OR2 (N3642, N3630, N3317);
xor XOR2 (N3643, N3623, N1452);
and AND2 (N3644, N3640, N3298);
nand NAND4 (N3645, N3628, N2220, N2066, N3477);
nor NOR2 (N3646, N3643, N1408);
nand NAND4 (N3647, N3620, N2813, N1143, N1171);
nand NAND4 (N3648, N3641, N3135, N3467, N858);
xor XOR2 (N3649, N3637, N2404);
nand NAND2 (N3650, N3649, N2855);
or OR3 (N3651, N3627, N279, N2882);
and AND3 (N3652, N3651, N2175, N105);
xor XOR2 (N3653, N3645, N2050);
not NOT1 (N3654, N3617);
xor XOR2 (N3655, N3648, N1217);
or OR3 (N3656, N3644, N3338, N2067);
nand NAND2 (N3657, N3650, N2118);
nand NAND4 (N3658, N3657, N3331, N108, N405);
buf BUF1 (N3659, N3655);
xor XOR2 (N3660, N3653, N1062);
not NOT1 (N3661, N3658);
xor XOR2 (N3662, N3656, N3040);
buf BUF1 (N3663, N3647);
buf BUF1 (N3664, N3663);
xor XOR2 (N3665, N3654, N1116);
xor XOR2 (N3666, N3646, N2508);
and AND2 (N3667, N3662, N2013);
not NOT1 (N3668, N3659);
or OR4 (N3669, N3665, N3224, N3630, N2837);
xor XOR2 (N3670, N3634, N1134);
nor NOR2 (N3671, N3660, N119);
not NOT1 (N3672, N3652);
not NOT1 (N3673, N3671);
or OR2 (N3674, N3666, N3419);
and AND4 (N3675, N3664, N1032, N2253, N789);
nand NAND3 (N3676, N3670, N83, N3525);
and AND4 (N3677, N3672, N1934, N2959, N2242);
not NOT1 (N3678, N3674);
not NOT1 (N3679, N3668);
nand NAND3 (N3680, N3679, N1542, N11);
nor NOR4 (N3681, N3677, N1949, N631, N1138);
buf BUF1 (N3682, N3673);
nand NAND2 (N3683, N3667, N2814);
or OR2 (N3684, N3680, N2814);
buf BUF1 (N3685, N3676);
or OR3 (N3686, N3675, N1767, N2061);
nand NAND4 (N3687, N3642, N2459, N760, N1903);
nor NOR2 (N3688, N3686, N3409);
nand NAND3 (N3689, N3681, N2891, N3544);
xor XOR2 (N3690, N3685, N164);
xor XOR2 (N3691, N3682, N2259);
nand NAND4 (N3692, N3688, N2846, N3285, N1327);
buf BUF1 (N3693, N3691);
nand NAND4 (N3694, N3684, N3353, N2446, N3100);
buf BUF1 (N3695, N3669);
and AND2 (N3696, N3683, N973);
nor NOR4 (N3697, N3695, N871, N427, N2609);
or OR4 (N3698, N3693, N2449, N1164, N466);
xor XOR2 (N3699, N3689, N1848);
nor NOR4 (N3700, N3696, N3550, N64, N219);
not NOT1 (N3701, N3700);
and AND2 (N3702, N3687, N3476);
nand NAND2 (N3703, N3690, N2800);
or OR4 (N3704, N3692, N1505, N2250, N2003);
xor XOR2 (N3705, N3697, N1207);
nor NOR4 (N3706, N3705, N3124, N2116, N3650);
nor NOR2 (N3707, N3702, N3653);
buf BUF1 (N3708, N3661);
and AND2 (N3709, N3707, N2554);
and AND2 (N3710, N3694, N3355);
not NOT1 (N3711, N3709);
not NOT1 (N3712, N3699);
nor NOR3 (N3713, N3706, N3041, N1855);
nand NAND4 (N3714, N3713, N437, N2095, N3405);
buf BUF1 (N3715, N3678);
buf BUF1 (N3716, N3703);
nand NAND3 (N3717, N3698, N1554, N2796);
or OR3 (N3718, N3708, N2220, N256);
not NOT1 (N3719, N3710);
nand NAND4 (N3720, N3712, N3558, N2701, N2031);
nand NAND4 (N3721, N3718, N1314, N3049, N524);
or OR3 (N3722, N3714, N980, N3500);
xor XOR2 (N3723, N3715, N943);
or OR2 (N3724, N3720, N485);
and AND3 (N3725, N3704, N62, N3436);
xor XOR2 (N3726, N3711, N187);
xor XOR2 (N3727, N3719, N2248);
buf BUF1 (N3728, N3727);
nand NAND2 (N3729, N3721, N784);
and AND2 (N3730, N3729, N2395);
nand NAND3 (N3731, N3728, N2136, N1779);
nor NOR3 (N3732, N3725, N3076, N590);
nor NOR3 (N3733, N3701, N2718, N1065);
or OR3 (N3734, N3730, N3002, N689);
buf BUF1 (N3735, N3724);
not NOT1 (N3736, N3716);
or OR4 (N3737, N3734, N2235, N1818, N1264);
or OR2 (N3738, N3735, N1980);
nand NAND3 (N3739, N3726, N1899, N3704);
xor XOR2 (N3740, N3739, N1773);
nor NOR3 (N3741, N3731, N1239, N681);
and AND3 (N3742, N3717, N2455, N653);
not NOT1 (N3743, N3723);
and AND4 (N3744, N3743, N232, N85, N2596);
nand NAND3 (N3745, N3722, N2718, N2415);
nor NOR2 (N3746, N3740, N3119);
not NOT1 (N3747, N3737);
or OR2 (N3748, N3745, N637);
xor XOR2 (N3749, N3744, N1454);
and AND4 (N3750, N3738, N1236, N495, N1862);
nor NOR2 (N3751, N3733, N2293);
or OR3 (N3752, N3732, N304, N467);
or OR3 (N3753, N3751, N2008, N2341);
or OR4 (N3754, N3742, N3338, N48, N3430);
nand NAND4 (N3755, N3749, N2845, N362, N567);
xor XOR2 (N3756, N3750, N1771);
or OR3 (N3757, N3753, N1737, N2683);
xor XOR2 (N3758, N3757, N3656);
and AND2 (N3759, N3747, N20);
buf BUF1 (N3760, N3748);
and AND2 (N3761, N3741, N1252);
xor XOR2 (N3762, N3761, N3647);
nor NOR3 (N3763, N3752, N2235, N1492);
xor XOR2 (N3764, N3763, N1217);
xor XOR2 (N3765, N3755, N1684);
and AND4 (N3766, N3762, N2710, N1869, N1706);
or OR3 (N3767, N3760, N3162, N2999);
buf BUF1 (N3768, N3756);
nor NOR2 (N3769, N3736, N2186);
xor XOR2 (N3770, N3754, N1263);
nand NAND3 (N3771, N3769, N1875, N1206);
nand NAND4 (N3772, N3766, N1602, N906, N1053);
and AND2 (N3773, N3771, N3329);
buf BUF1 (N3774, N3746);
not NOT1 (N3775, N3767);
and AND2 (N3776, N3765, N894);
nor NOR2 (N3777, N3768, N484);
not NOT1 (N3778, N3770);
nand NAND2 (N3779, N3764, N1504);
nor NOR3 (N3780, N3758, N1760, N1330);
buf BUF1 (N3781, N3777);
xor XOR2 (N3782, N3775, N2341);
nand NAND2 (N3783, N3773, N822);
or OR3 (N3784, N3778, N529, N3748);
not NOT1 (N3785, N3782);
and AND4 (N3786, N3776, N523, N1505, N3702);
nand NAND3 (N3787, N3784, N417, N2255);
buf BUF1 (N3788, N3780);
nand NAND2 (N3789, N3786, N751);
buf BUF1 (N3790, N3772);
buf BUF1 (N3791, N3779);
xor XOR2 (N3792, N3785, N2802);
xor XOR2 (N3793, N3790, N2807);
xor XOR2 (N3794, N3789, N384);
nand NAND3 (N3795, N3794, N2767, N1051);
xor XOR2 (N3796, N3795, N3346);
buf BUF1 (N3797, N3792);
or OR3 (N3798, N3781, N3502, N1211);
not NOT1 (N3799, N3793);
and AND2 (N3800, N3788, N2912);
or OR2 (N3801, N3783, N11);
nand NAND2 (N3802, N3791, N300);
xor XOR2 (N3803, N3787, N1147);
nand NAND2 (N3804, N3801, N262);
xor XOR2 (N3805, N3774, N530);
nor NOR2 (N3806, N3804, N1444);
buf BUF1 (N3807, N3799);
nand NAND2 (N3808, N3805, N1039);
nand NAND3 (N3809, N3796, N2312, N611);
and AND3 (N3810, N3759, N2560, N3367);
buf BUF1 (N3811, N3803);
nor NOR4 (N3812, N3808, N714, N2805, N1570);
buf BUF1 (N3813, N3809);
buf BUF1 (N3814, N3811);
buf BUF1 (N3815, N3798);
nand NAND4 (N3816, N3797, N2330, N580, N222);
nor NOR4 (N3817, N3806, N1109, N3072, N978);
nor NOR3 (N3818, N3807, N2959, N2566);
buf BUF1 (N3819, N3800);
or OR3 (N3820, N3815, N2214, N1650);
or OR3 (N3821, N3810, N2785, N2640);
nand NAND2 (N3822, N3814, N2616);
nand NAND4 (N3823, N3821, N3679, N327, N2072);
xor XOR2 (N3824, N3819, N2268);
xor XOR2 (N3825, N3818, N2345);
buf BUF1 (N3826, N3813);
not NOT1 (N3827, N3812);
xor XOR2 (N3828, N3822, N1158);
and AND4 (N3829, N3828, N2392, N585, N1805);
xor XOR2 (N3830, N3826, N564);
xor XOR2 (N3831, N3816, N1864);
xor XOR2 (N3832, N3829, N1988);
xor XOR2 (N3833, N3824, N587);
and AND3 (N3834, N3832, N709, N1665);
and AND3 (N3835, N3825, N521, N2397);
buf BUF1 (N3836, N3823);
nand NAND3 (N3837, N3836, N1151, N3075);
nand NAND3 (N3838, N3817, N3473, N2602);
or OR2 (N3839, N3837, N334);
and AND3 (N3840, N3820, N1771, N1607);
not NOT1 (N3841, N3839);
nor NOR4 (N3842, N3827, N259, N3663, N3094);
nor NOR4 (N3843, N3841, N528, N1909, N985);
not NOT1 (N3844, N3843);
buf BUF1 (N3845, N3842);
xor XOR2 (N3846, N3833, N319);
nor NOR4 (N3847, N3838, N3398, N1794, N65);
or OR3 (N3848, N3847, N3, N3572);
nor NOR2 (N3849, N3840, N3074);
and AND4 (N3850, N3846, N2541, N3031, N2074);
nand NAND2 (N3851, N3802, N1194);
xor XOR2 (N3852, N3830, N2896);
not NOT1 (N3853, N3834);
not NOT1 (N3854, N3845);
nor NOR2 (N3855, N3835, N2742);
not NOT1 (N3856, N3851);
and AND4 (N3857, N3831, N747, N3592, N2547);
buf BUF1 (N3858, N3849);
xor XOR2 (N3859, N3858, N3556);
nor NOR2 (N3860, N3850, N3630);
and AND4 (N3861, N3848, N3206, N360, N2113);
nor NOR3 (N3862, N3853, N3252, N1468);
buf BUF1 (N3863, N3861);
not NOT1 (N3864, N3859);
not NOT1 (N3865, N3854);
xor XOR2 (N3866, N3865, N85);
or OR4 (N3867, N3863, N2168, N3066, N1514);
nand NAND3 (N3868, N3866, N400, N512);
and AND2 (N3869, N3868, N1472);
nor NOR4 (N3870, N3864, N1345, N947, N3697);
not NOT1 (N3871, N3856);
xor XOR2 (N3872, N3852, N2813);
nand NAND3 (N3873, N3862, N1492, N3563);
nand NAND2 (N3874, N3857, N577);
nand NAND3 (N3875, N3873, N2078, N2417);
not NOT1 (N3876, N3870);
nor NOR2 (N3877, N3875, N78);
or OR4 (N3878, N3872, N2207, N1770, N1131);
nand NAND4 (N3879, N3878, N1694, N542, N2775);
xor XOR2 (N3880, N3844, N2743);
nor NOR3 (N3881, N3871, N527, N2273);
buf BUF1 (N3882, N3876);
not NOT1 (N3883, N3881);
xor XOR2 (N3884, N3874, N1869);
and AND3 (N3885, N3884, N3374, N229);
or OR3 (N3886, N3882, N1171, N731);
xor XOR2 (N3887, N3855, N3369);
or OR4 (N3888, N3860, N1326, N3325, N2941);
buf BUF1 (N3889, N3869);
nor NOR3 (N3890, N3877, N3256, N3688);
and AND3 (N3891, N3885, N1366, N1528);
nand NAND3 (N3892, N3890, N2968, N385);
nand NAND4 (N3893, N3867, N3651, N963, N3701);
nor NOR3 (N3894, N3880, N3298, N547);
or OR4 (N3895, N3891, N2271, N255, N1979);
xor XOR2 (N3896, N3894, N2513);
xor XOR2 (N3897, N3896, N3055);
nor NOR3 (N3898, N3879, N143, N2507);
xor XOR2 (N3899, N3897, N3816);
and AND2 (N3900, N3886, N2728);
xor XOR2 (N3901, N3893, N3251);
nand NAND3 (N3902, N3895, N1167, N1099);
nand NAND2 (N3903, N3888, N2954);
not NOT1 (N3904, N3892);
xor XOR2 (N3905, N3899, N2175);
or OR3 (N3906, N3898, N3503, N1934);
and AND3 (N3907, N3904, N1629, N805);
not NOT1 (N3908, N3901);
and AND4 (N3909, N3883, N698, N2165, N792);
and AND4 (N3910, N3909, N1642, N837, N3133);
nand NAND4 (N3911, N3906, N3867, N1397, N1333);
or OR2 (N3912, N3902, N2484);
and AND3 (N3913, N3907, N3287, N784);
nor NOR3 (N3914, N3887, N3109, N154);
or OR3 (N3915, N3903, N2033, N1012);
buf BUF1 (N3916, N3915);
nor NOR3 (N3917, N3913, N2567, N866);
or OR4 (N3918, N3889, N632, N2953, N562);
buf BUF1 (N3919, N3916);
or OR4 (N3920, N3900, N2864, N344, N256);
nor NOR4 (N3921, N3920, N1537, N441, N1665);
nand NAND3 (N3922, N3921, N3756, N2020);
nor NOR4 (N3923, N3911, N1378, N2682, N1508);
not NOT1 (N3924, N3918);
xor XOR2 (N3925, N3922, N1705);
and AND3 (N3926, N3914, N252, N887);
not NOT1 (N3927, N3910);
or OR2 (N3928, N3905, N3303);
and AND3 (N3929, N3924, N3601, N3853);
xor XOR2 (N3930, N3912, N2651);
buf BUF1 (N3931, N3908);
nand NAND3 (N3932, N3929, N2752, N1832);
xor XOR2 (N3933, N3926, N3490);
not NOT1 (N3934, N3925);
nand NAND2 (N3935, N3930, N3494);
nand NAND3 (N3936, N3932, N1572, N527);
nand NAND3 (N3937, N3933, N3419, N177);
xor XOR2 (N3938, N3934, N3595);
buf BUF1 (N3939, N3931);
or OR4 (N3940, N3923, N2370, N2040, N2629);
buf BUF1 (N3941, N3939);
buf BUF1 (N3942, N3938);
nor NOR3 (N3943, N3927, N159, N1137);
and AND2 (N3944, N3940, N1368);
nor NOR3 (N3945, N3941, N1183, N1635);
and AND2 (N3946, N3919, N1559);
nand NAND4 (N3947, N3943, N2298, N3390, N3018);
not NOT1 (N3948, N3935);
nor NOR3 (N3949, N3946, N2797, N1641);
not NOT1 (N3950, N3949);
or OR4 (N3951, N3944, N157, N1389, N1958);
xor XOR2 (N3952, N3936, N801);
or OR4 (N3953, N3917, N2548, N1493, N996);
not NOT1 (N3954, N3947);
not NOT1 (N3955, N3928);
buf BUF1 (N3956, N3952);
and AND4 (N3957, N3951, N1350, N2454, N3277);
and AND2 (N3958, N3945, N3162);
nand NAND4 (N3959, N3937, N1467, N1714, N3027);
and AND3 (N3960, N3957, N1869, N654);
not NOT1 (N3961, N3942);
buf BUF1 (N3962, N3950);
or OR4 (N3963, N3960, N783, N112, N1174);
and AND2 (N3964, N3963, N2506);
nor NOR2 (N3965, N3958, N2678);
nand NAND2 (N3966, N3962, N572);
or OR4 (N3967, N3964, N2713, N3066, N714);
xor XOR2 (N3968, N3953, N2527);
or OR4 (N3969, N3968, N1665, N3134, N2113);
or OR4 (N3970, N3959, N1033, N252, N1031);
nand NAND3 (N3971, N3966, N392, N1687);
xor XOR2 (N3972, N3955, N283);
nand NAND4 (N3973, N3961, N706, N1581, N1948);
nand NAND3 (N3974, N3971, N3600, N1573);
nand NAND3 (N3975, N3970, N1117, N2366);
nor NOR2 (N3976, N3975, N3763);
nand NAND2 (N3977, N3972, N1252);
buf BUF1 (N3978, N3956);
nand NAND2 (N3979, N3954, N870);
xor XOR2 (N3980, N3969, N1590);
and AND2 (N3981, N3948, N842);
nor NOR2 (N3982, N3978, N3485);
not NOT1 (N3983, N3979);
nor NOR4 (N3984, N3977, N3534, N1264, N118);
not NOT1 (N3985, N3982);
nand NAND4 (N3986, N3976, N3441, N2080, N2697);
nand NAND2 (N3987, N3983, N2998);
buf BUF1 (N3988, N3980);
nand NAND2 (N3989, N3987, N3416);
or OR2 (N3990, N3988, N637);
buf BUF1 (N3991, N3989);
not NOT1 (N3992, N3974);
not NOT1 (N3993, N3965);
not NOT1 (N3994, N3993);
xor XOR2 (N3995, N3985, N295);
nand NAND2 (N3996, N3986, N1250);
nor NOR4 (N3997, N3990, N3609, N3152, N683);
not NOT1 (N3998, N3991);
or OR3 (N3999, N3994, N2051, N3752);
buf BUF1 (N4000, N3981);
and AND4 (N4001, N3996, N2464, N2383, N1308);
not NOT1 (N4002, N3992);
not NOT1 (N4003, N4002);
nor NOR4 (N4004, N4003, N2477, N572, N3633);
and AND2 (N4005, N4004, N2430);
nor NOR2 (N4006, N4005, N1519);
xor XOR2 (N4007, N4001, N65);
xor XOR2 (N4008, N3995, N1545);
xor XOR2 (N4009, N3973, N657);
xor XOR2 (N4010, N4000, N3419);
or OR3 (N4011, N3967, N3753, N781);
not NOT1 (N4012, N3997);
or OR2 (N4013, N4009, N3489);
not NOT1 (N4014, N4011);
xor XOR2 (N4015, N3984, N3276);
not NOT1 (N4016, N4010);
nand NAND4 (N4017, N4006, N3952, N3431, N736);
buf BUF1 (N4018, N4016);
buf BUF1 (N4019, N3998);
nor NOR3 (N4020, N4014, N3293, N1244);
not NOT1 (N4021, N4007);
buf BUF1 (N4022, N4018);
and AND2 (N4023, N4012, N3438);
xor XOR2 (N4024, N4017, N3046);
xor XOR2 (N4025, N3999, N3050);
and AND2 (N4026, N4008, N2730);
and AND3 (N4027, N4021, N388, N1660);
nand NAND3 (N4028, N4023, N2241, N1531);
and AND4 (N4029, N4015, N108, N1813, N1759);
xor XOR2 (N4030, N4029, N3054);
nand NAND4 (N4031, N4020, N1880, N368, N2152);
or OR4 (N4032, N4031, N3939, N647, N2010);
xor XOR2 (N4033, N4028, N2011);
xor XOR2 (N4034, N4019, N3563);
buf BUF1 (N4035, N4030);
nand NAND3 (N4036, N4027, N3505, N3647);
or OR3 (N4037, N4026, N2546, N474);
buf BUF1 (N4038, N4022);
nand NAND4 (N4039, N4032, N2318, N394, N3499);
buf BUF1 (N4040, N4036);
xor XOR2 (N4041, N4035, N1692);
nor NOR3 (N4042, N4013, N1672, N1938);
nor NOR2 (N4043, N4040, N3189);
or OR4 (N4044, N4042, N3285, N2658, N1328);
and AND2 (N4045, N4043, N3924);
xor XOR2 (N4046, N4041, N1890);
and AND4 (N4047, N4025, N1084, N1877, N2655);
nand NAND3 (N4048, N4038, N1775, N430);
nor NOR4 (N4049, N4047, N2334, N2640, N3567);
xor XOR2 (N4050, N4044, N1850);
nor NOR3 (N4051, N4024, N273, N2435);
xor XOR2 (N4052, N4049, N383);
or OR2 (N4053, N4033, N2519);
xor XOR2 (N4054, N4034, N2849);
and AND4 (N4055, N4037, N2013, N3053, N2310);
or OR4 (N4056, N4039, N2981, N3955, N2236);
not NOT1 (N4057, N4051);
and AND2 (N4058, N4050, N1318);
xor XOR2 (N4059, N4054, N3523);
buf BUF1 (N4060, N4048);
not NOT1 (N4061, N4052);
nand NAND4 (N4062, N4055, N2817, N3762, N2651);
xor XOR2 (N4063, N4046, N1355);
nor NOR3 (N4064, N4060, N1386, N4022);
nor NOR2 (N4065, N4045, N2125);
xor XOR2 (N4066, N4057, N2311);
nand NAND4 (N4067, N4061, N546, N1930, N2716);
nand NAND4 (N4068, N4062, N3979, N442, N3787);
and AND3 (N4069, N4053, N2804, N2329);
not NOT1 (N4070, N4056);
buf BUF1 (N4071, N4064);
nand NAND4 (N4072, N4070, N2700, N811, N3870);
nor NOR2 (N4073, N4066, N1870);
not NOT1 (N4074, N4067);
nand NAND4 (N4075, N4063, N2709, N1646, N974);
not NOT1 (N4076, N4059);
or OR4 (N4077, N4071, N3733, N1699, N2478);
not NOT1 (N4078, N4077);
xor XOR2 (N4079, N4072, N2864);
nand NAND4 (N4080, N4074, N1735, N3216, N617);
not NOT1 (N4081, N4068);
and AND3 (N4082, N4078, N2190, N1739);
xor XOR2 (N4083, N4076, N828);
not NOT1 (N4084, N4083);
and AND2 (N4085, N4075, N3976);
not NOT1 (N4086, N4085);
xor XOR2 (N4087, N4081, N1706);
xor XOR2 (N4088, N4073, N3427);
nand NAND3 (N4089, N4080, N2202, N2251);
or OR3 (N4090, N4065, N1810, N903);
or OR4 (N4091, N4089, N3810, N711, N999);
nor NOR3 (N4092, N4088, N434, N1185);
nand NAND4 (N4093, N4082, N3631, N87, N2967);
not NOT1 (N4094, N4091);
buf BUF1 (N4095, N4093);
xor XOR2 (N4096, N4058, N3962);
buf BUF1 (N4097, N4086);
xor XOR2 (N4098, N4092, N3374);
nor NOR3 (N4099, N4079, N3965, N2877);
buf BUF1 (N4100, N4084);
or OR4 (N4101, N4096, N1368, N2628, N74);
nand NAND2 (N4102, N4098, N1172);
buf BUF1 (N4103, N4094);
buf BUF1 (N4104, N4090);
not NOT1 (N4105, N4087);
buf BUF1 (N4106, N4095);
and AND4 (N4107, N4103, N4000, N2757, N116);
or OR4 (N4108, N4105, N1290, N3329, N3897);
nor NOR2 (N4109, N4104, N244);
buf BUF1 (N4110, N4069);
xor XOR2 (N4111, N4100, N1832);
nor NOR3 (N4112, N4099, N1403, N2056);
and AND4 (N4113, N4108, N728, N3843, N12);
buf BUF1 (N4114, N4097);
buf BUF1 (N4115, N4107);
nand NAND2 (N4116, N4106, N1929);
nand NAND3 (N4117, N4116, N3518, N2374);
nor NOR2 (N4118, N4114, N139);
and AND2 (N4119, N4112, N2626);
and AND3 (N4120, N4115, N362, N3021);
and AND4 (N4121, N4109, N2868, N3130, N915);
nor NOR3 (N4122, N4110, N563, N150);
and AND3 (N4123, N4101, N3109, N624);
nand NAND4 (N4124, N4117, N2761, N2231, N1576);
nor NOR3 (N4125, N4113, N1378, N1049);
and AND2 (N4126, N4121, N3211);
not NOT1 (N4127, N4122);
buf BUF1 (N4128, N4118);
nor NOR2 (N4129, N4125, N3265);
buf BUF1 (N4130, N4123);
buf BUF1 (N4131, N4127);
buf BUF1 (N4132, N4120);
nor NOR3 (N4133, N4124, N1350, N1597);
or OR4 (N4134, N4119, N966, N3074, N1809);
or OR3 (N4135, N4130, N1419, N2814);
nor NOR3 (N4136, N4134, N2674, N1961);
or OR3 (N4137, N4128, N125, N156);
nor NOR4 (N4138, N4137, N2506, N1726, N2709);
xor XOR2 (N4139, N4138, N371);
and AND2 (N4140, N4126, N431);
xor XOR2 (N4141, N4129, N810);
and AND2 (N4142, N4135, N1329);
nor NOR3 (N4143, N4132, N1933, N2129);
not NOT1 (N4144, N4140);
buf BUF1 (N4145, N4102);
or OR3 (N4146, N4139, N411, N1822);
or OR3 (N4147, N4144, N2554, N3409);
nor NOR2 (N4148, N4141, N992);
buf BUF1 (N4149, N4136);
xor XOR2 (N4150, N4147, N2391);
nor NOR2 (N4151, N4150, N1877);
buf BUF1 (N4152, N4111);
and AND3 (N4153, N4146, N1778, N395);
xor XOR2 (N4154, N4151, N3484);
nand NAND3 (N4155, N4142, N1238, N2453);
not NOT1 (N4156, N4148);
not NOT1 (N4157, N4152);
nor NOR2 (N4158, N4153, N3346);
not NOT1 (N4159, N4131);
not NOT1 (N4160, N4157);
not NOT1 (N4161, N4158);
xor XOR2 (N4162, N4155, N1864);
buf BUF1 (N4163, N4156);
and AND3 (N4164, N4145, N1816, N3187);
xor XOR2 (N4165, N4159, N3585);
or OR4 (N4166, N4163, N2404, N710, N1280);
nor NOR3 (N4167, N4162, N971, N2204);
buf BUF1 (N4168, N4165);
nor NOR2 (N4169, N4166, N1379);
nor NOR3 (N4170, N4149, N3626, N3225);
nand NAND4 (N4171, N4160, N326, N1736, N3874);
and AND4 (N4172, N4171, N2802, N3897, N4089);
not NOT1 (N4173, N4172);
or OR2 (N4174, N4169, N1743);
and AND2 (N4175, N4143, N2820);
not NOT1 (N4176, N4168);
nor NOR4 (N4177, N4133, N2823, N981, N1275);
or OR2 (N4178, N4176, N430);
nand NAND2 (N4179, N4167, N2672);
not NOT1 (N4180, N4177);
nand NAND2 (N4181, N4161, N3203);
not NOT1 (N4182, N4175);
xor XOR2 (N4183, N4181, N1565);
nand NAND4 (N4184, N4182, N2249, N2567, N3382);
not NOT1 (N4185, N4178);
or OR3 (N4186, N4170, N1108, N3834);
or OR2 (N4187, N4174, N3008);
or OR3 (N4188, N4164, N1219, N4181);
or OR3 (N4189, N4154, N1648, N1448);
nand NAND3 (N4190, N4184, N4100, N3170);
nand NAND2 (N4191, N4188, N3075);
xor XOR2 (N4192, N4185, N512);
nor NOR4 (N4193, N4190, N2841, N2759, N2487);
not NOT1 (N4194, N4187);
nor NOR3 (N4195, N4173, N2633, N2859);
buf BUF1 (N4196, N4195);
nor NOR3 (N4197, N4189, N3402, N2397);
or OR4 (N4198, N4196, N2818, N416, N3771);
or OR4 (N4199, N4197, N1187, N1741, N930);
or OR2 (N4200, N4194, N2551);
and AND3 (N4201, N4186, N2211, N3605);
xor XOR2 (N4202, N4198, N3375);
buf BUF1 (N4203, N4180);
or OR2 (N4204, N4193, N2767);
nor NOR3 (N4205, N4201, N2945, N2413);
buf BUF1 (N4206, N4204);
and AND4 (N4207, N4192, N673, N1619, N3701);
not NOT1 (N4208, N4179);
nor NOR4 (N4209, N4207, N1762, N3452, N1221);
or OR3 (N4210, N4206, N950, N3980);
and AND4 (N4211, N4210, N4071, N2993, N4042);
xor XOR2 (N4212, N4203, N2639);
nand NAND4 (N4213, N4183, N679, N1327, N288);
nor NOR3 (N4214, N4200, N1586, N3438);
and AND3 (N4215, N4191, N112, N1719);
or OR2 (N4216, N4214, N277);
nor NOR3 (N4217, N4215, N407, N1415);
nand NAND4 (N4218, N4209, N4124, N1466, N4033);
not NOT1 (N4219, N4202);
nand NAND3 (N4220, N4213, N688, N3425);
or OR3 (N4221, N4219, N1042, N2641);
buf BUF1 (N4222, N4220);
xor XOR2 (N4223, N4199, N2672);
not NOT1 (N4224, N4216);
buf BUF1 (N4225, N4205);
buf BUF1 (N4226, N4222);
or OR2 (N4227, N4221, N285);
or OR4 (N4228, N4223, N1238, N1854, N1125);
buf BUF1 (N4229, N4225);
xor XOR2 (N4230, N4212, N2524);
nor NOR4 (N4231, N4211, N214, N3429, N853);
nand NAND4 (N4232, N4230, N3838, N96, N2050);
nor NOR2 (N4233, N4217, N969);
not NOT1 (N4234, N4228);
nor NOR4 (N4235, N4208, N3943, N889, N3887);
nand NAND4 (N4236, N4231, N85, N4048, N4098);
not NOT1 (N4237, N4227);
not NOT1 (N4238, N4226);
or OR3 (N4239, N4229, N3778, N351);
nor NOR3 (N4240, N4239, N116, N14);
and AND4 (N4241, N4232, N51, N4208, N1637);
nand NAND4 (N4242, N4237, N3907, N448, N231);
and AND3 (N4243, N4224, N711, N1059);
or OR4 (N4244, N4233, N990, N3270, N1532);
xor XOR2 (N4245, N4242, N1948);
not NOT1 (N4246, N4243);
nand NAND4 (N4247, N4240, N1186, N3181, N699);
not NOT1 (N4248, N4238);
nand NAND4 (N4249, N4236, N4178, N3587, N1843);
xor XOR2 (N4250, N4247, N1828);
xor XOR2 (N4251, N4234, N3096);
not NOT1 (N4252, N4235);
or OR2 (N4253, N4252, N755);
nand NAND2 (N4254, N4245, N3044);
xor XOR2 (N4255, N4246, N2787);
nand NAND2 (N4256, N4253, N2174);
and AND4 (N4257, N4254, N73, N2687, N4235);
or OR2 (N4258, N4248, N2257);
and AND4 (N4259, N4249, N3629, N759, N3382);
and AND3 (N4260, N4250, N1916, N612);
or OR3 (N4261, N4259, N1967, N283);
and AND4 (N4262, N4257, N622, N4193, N4132);
xor XOR2 (N4263, N4251, N2128);
xor XOR2 (N4264, N4218, N2599);
buf BUF1 (N4265, N4260);
xor XOR2 (N4266, N4265, N2793);
nor NOR2 (N4267, N4241, N457);
nor NOR2 (N4268, N4261, N580);
buf BUF1 (N4269, N4267);
buf BUF1 (N4270, N4268);
nor NOR2 (N4271, N4269, N3194);
xor XOR2 (N4272, N4258, N330);
not NOT1 (N4273, N4266);
buf BUF1 (N4274, N4270);
or OR2 (N4275, N4264, N2183);
not NOT1 (N4276, N4255);
nor NOR3 (N4277, N4275, N2996, N103);
not NOT1 (N4278, N4276);
nor NOR2 (N4279, N4274, N2511);
nand NAND3 (N4280, N4273, N2791, N1147);
nor NOR3 (N4281, N4280, N2823, N191);
or OR2 (N4282, N4281, N297);
not NOT1 (N4283, N4262);
or OR4 (N4284, N4282, N1718, N3791, N1239);
nand NAND2 (N4285, N4256, N366);
or OR4 (N4286, N4285, N2612, N1544, N18);
or OR3 (N4287, N4286, N2238, N2939);
xor XOR2 (N4288, N4272, N595);
nor NOR4 (N4289, N4271, N1522, N3244, N98);
nor NOR4 (N4290, N4244, N100, N3792, N840);
nand NAND2 (N4291, N4287, N3021);
or OR3 (N4292, N4288, N2523, N182);
and AND2 (N4293, N4291, N1321);
xor XOR2 (N4294, N4283, N2414);
nor NOR2 (N4295, N4293, N2124);
nor NOR3 (N4296, N4290, N735, N3838);
and AND4 (N4297, N4289, N87, N2540, N3332);
or OR4 (N4298, N4263, N3496, N1212, N2607);
or OR2 (N4299, N4295, N3587);
nand NAND3 (N4300, N4297, N3621, N507);
not NOT1 (N4301, N4300);
and AND2 (N4302, N4284, N25);
not NOT1 (N4303, N4292);
not NOT1 (N4304, N4302);
buf BUF1 (N4305, N4277);
buf BUF1 (N4306, N4294);
nand NAND2 (N4307, N4296, N2489);
and AND2 (N4308, N4278, N2847);
nand NAND2 (N4309, N4301, N1505);
or OR2 (N4310, N4298, N1871);
nand NAND2 (N4311, N4310, N1347);
buf BUF1 (N4312, N4304);
nor NOR2 (N4313, N4307, N2121);
nand NAND3 (N4314, N4305, N1731, N1206);
or OR3 (N4315, N4303, N1798, N3025);
or OR4 (N4316, N4314, N2978, N2169, N4276);
buf BUF1 (N4317, N4312);
nand NAND2 (N4318, N4313, N964);
and AND2 (N4319, N4308, N776);
not NOT1 (N4320, N4306);
and AND3 (N4321, N4318, N308, N3366);
buf BUF1 (N4322, N4311);
nand NAND4 (N4323, N4321, N4063, N3092, N2850);
xor XOR2 (N4324, N4316, N3501);
xor XOR2 (N4325, N4324, N202);
nand NAND4 (N4326, N4279, N2074, N3578, N1809);
xor XOR2 (N4327, N4325, N2853);
not NOT1 (N4328, N4323);
nor NOR4 (N4329, N4319, N3591, N2391, N1754);
not NOT1 (N4330, N4327);
buf BUF1 (N4331, N4315);
not NOT1 (N4332, N4328);
nand NAND3 (N4333, N4330, N1298, N1785);
nor NOR2 (N4334, N4332, N2236);
xor XOR2 (N4335, N4326, N516);
or OR3 (N4336, N4329, N1541, N576);
or OR3 (N4337, N4331, N1399, N450);
nor NOR3 (N4338, N4335, N722, N985);
nor NOR3 (N4339, N4336, N3238, N1735);
nand NAND4 (N4340, N4320, N2630, N4331, N1230);
nand NAND2 (N4341, N4338, N3219);
or OR3 (N4342, N4341, N895, N3349);
xor XOR2 (N4343, N4299, N1527);
not NOT1 (N4344, N4339);
xor XOR2 (N4345, N4340, N1035);
and AND4 (N4346, N4333, N2167, N3428, N4227);
nand NAND4 (N4347, N4334, N635, N3657, N2198);
nand NAND4 (N4348, N4344, N3867, N2867, N3075);
not NOT1 (N4349, N4343);
and AND3 (N4350, N4347, N4094, N2810);
and AND2 (N4351, N4346, N1914);
or OR4 (N4352, N4337, N386, N987, N1839);
nand NAND2 (N4353, N4350, N762);
not NOT1 (N4354, N4317);
xor XOR2 (N4355, N4349, N1671);
nand NAND2 (N4356, N4352, N439);
and AND3 (N4357, N4354, N3931, N3822);
nor NOR2 (N4358, N4342, N3116);
nand NAND3 (N4359, N4356, N49, N3546);
nor NOR2 (N4360, N4355, N3350);
and AND4 (N4361, N4345, N860, N2232, N2392);
and AND4 (N4362, N4359, N1273, N3904, N1438);
or OR4 (N4363, N4362, N3227, N707, N2098);
or OR2 (N4364, N4357, N1725);
or OR3 (N4365, N4360, N1071, N614);
and AND4 (N4366, N4351, N1942, N3902, N4019);
buf BUF1 (N4367, N4309);
buf BUF1 (N4368, N4364);
xor XOR2 (N4369, N4322, N1681);
buf BUF1 (N4370, N4365);
and AND4 (N4371, N4348, N493, N613, N2361);
xor XOR2 (N4372, N4358, N499);
and AND4 (N4373, N4353, N1243, N3229, N658);
or OR2 (N4374, N4367, N541);
and AND2 (N4375, N4374, N90);
or OR4 (N4376, N4375, N4094, N2590, N3170);
xor XOR2 (N4377, N4372, N1729);
not NOT1 (N4378, N4371);
nand NAND3 (N4379, N4369, N1014, N990);
buf BUF1 (N4380, N4378);
buf BUF1 (N4381, N4373);
nand NAND4 (N4382, N4368, N4246, N130, N4119);
xor XOR2 (N4383, N4382, N3343);
nor NOR3 (N4384, N4383, N948, N3759);
nand NAND3 (N4385, N4380, N1243, N3149);
or OR2 (N4386, N4377, N2762);
buf BUF1 (N4387, N4379);
nand NAND4 (N4388, N4363, N2098, N1765, N4088);
nand NAND3 (N4389, N4366, N2709, N3502);
and AND3 (N4390, N4387, N2306, N3410);
and AND2 (N4391, N4370, N645);
nand NAND3 (N4392, N4386, N2639, N992);
and AND2 (N4393, N4381, N1951);
buf BUF1 (N4394, N4393);
nor NOR3 (N4395, N4376, N779, N2292);
and AND3 (N4396, N4390, N425, N1378);
or OR4 (N4397, N4389, N3301, N1140, N1837);
not NOT1 (N4398, N4384);
and AND2 (N4399, N4361, N3822);
or OR2 (N4400, N4388, N726);
nand NAND4 (N4401, N4385, N2490, N696, N2463);
nand NAND3 (N4402, N4398, N778, N1100);
or OR4 (N4403, N4394, N247, N4159, N3198);
not NOT1 (N4404, N4396);
buf BUF1 (N4405, N4403);
xor XOR2 (N4406, N4391, N112);
and AND2 (N4407, N4395, N1182);
buf BUF1 (N4408, N4400);
buf BUF1 (N4409, N4399);
and AND4 (N4410, N4406, N4291, N975, N311);
nor NOR2 (N4411, N4410, N3907);
or OR4 (N4412, N4411, N1971, N644, N2926);
nand NAND3 (N4413, N4404, N1325, N2971);
buf BUF1 (N4414, N4392);
nand NAND2 (N4415, N4401, N2243);
buf BUF1 (N4416, N4402);
or OR3 (N4417, N4415, N2806, N4221);
not NOT1 (N4418, N4412);
not NOT1 (N4419, N4397);
or OR4 (N4420, N4409, N360, N2783, N2980);
not NOT1 (N4421, N4419);
xor XOR2 (N4422, N4417, N156);
xor XOR2 (N4423, N4420, N1594);
not NOT1 (N4424, N4407);
nor NOR2 (N4425, N4422, N3787);
nand NAND4 (N4426, N4413, N1544, N2408, N3323);
or OR2 (N4427, N4416, N3738);
and AND2 (N4428, N4423, N836);
not NOT1 (N4429, N4428);
nand NAND4 (N4430, N4405, N2736, N1543, N2684);
and AND2 (N4431, N4427, N2065);
nand NAND3 (N4432, N4429, N1274, N1594);
and AND4 (N4433, N4408, N1510, N2846, N2937);
not NOT1 (N4434, N4421);
buf BUF1 (N4435, N4418);
and AND3 (N4436, N4432, N201, N1376);
or OR3 (N4437, N4431, N1608, N1847);
or OR2 (N4438, N4424, N3955);
nand NAND2 (N4439, N4425, N211);
and AND4 (N4440, N4435, N1877, N1181, N1461);
or OR3 (N4441, N4438, N254, N2207);
nand NAND2 (N4442, N4440, N2591);
not NOT1 (N4443, N4433);
buf BUF1 (N4444, N4434);
buf BUF1 (N4445, N4414);
nor NOR3 (N4446, N4426, N3331, N2766);
not NOT1 (N4447, N4445);
not NOT1 (N4448, N4446);
not NOT1 (N4449, N4448);
or OR3 (N4450, N4443, N2618, N2762);
xor XOR2 (N4451, N4439, N2017);
not NOT1 (N4452, N4430);
nand NAND2 (N4453, N4437, N1705);
or OR3 (N4454, N4452, N2258, N496);
or OR4 (N4455, N4451, N2069, N1196, N1623);
or OR4 (N4456, N4453, N3141, N1222, N3904);
nor NOR2 (N4457, N4441, N2184);
or OR2 (N4458, N4447, N2427);
or OR2 (N4459, N4449, N2579);
nand NAND3 (N4460, N4444, N1152, N855);
not NOT1 (N4461, N4458);
and AND2 (N4462, N4456, N1155);
nor NOR3 (N4463, N4442, N3611, N1259);
or OR2 (N4464, N4454, N150);
and AND3 (N4465, N4459, N4220, N3404);
or OR4 (N4466, N4457, N1608, N212, N879);
or OR4 (N4467, N4464, N830, N2058, N2910);
xor XOR2 (N4468, N4467, N858);
and AND2 (N4469, N4436, N157);
or OR3 (N4470, N4461, N2506, N1883);
buf BUF1 (N4471, N4460);
or OR2 (N4472, N4462, N1516);
not NOT1 (N4473, N4468);
and AND2 (N4474, N4463, N183);
nand NAND4 (N4475, N4469, N389, N2201, N1737);
xor XOR2 (N4476, N4474, N499);
nor NOR2 (N4477, N4450, N1461);
buf BUF1 (N4478, N4475);
nor NOR3 (N4479, N4478, N2711, N513);
buf BUF1 (N4480, N4473);
nor NOR3 (N4481, N4465, N2113, N3656);
not NOT1 (N4482, N4481);
nor NOR4 (N4483, N4466, N1590, N4312, N2788);
not NOT1 (N4484, N4472);
nand NAND2 (N4485, N4471, N3895);
buf BUF1 (N4486, N4482);
nand NAND4 (N4487, N4479, N3935, N3275, N2878);
nor NOR2 (N4488, N4485, N3673);
not NOT1 (N4489, N4477);
buf BUF1 (N4490, N4483);
nand NAND4 (N4491, N4476, N1427, N945, N2039);
nor NOR2 (N4492, N4455, N121);
buf BUF1 (N4493, N4490);
not NOT1 (N4494, N4480);
not NOT1 (N4495, N4486);
buf BUF1 (N4496, N4470);
and AND3 (N4497, N4493, N1638, N541);
nand NAND4 (N4498, N4492, N1236, N3383, N3922);
nor NOR4 (N4499, N4496, N3402, N2056, N2586);
not NOT1 (N4500, N4499);
nand NAND3 (N4501, N4498, N733, N3232);
and AND2 (N4502, N4489, N278);
and AND4 (N4503, N4491, N2905, N2797, N3840);
or OR4 (N4504, N4487, N2374, N613, N514);
nor NOR4 (N4505, N4504, N834, N187, N3645);
xor XOR2 (N4506, N4500, N4229);
nor NOR3 (N4507, N4495, N2743, N2230);
buf BUF1 (N4508, N4501);
or OR2 (N4509, N4497, N67);
nor NOR2 (N4510, N4506, N769);
not NOT1 (N4511, N4507);
or OR3 (N4512, N4511, N825, N2920);
not NOT1 (N4513, N4503);
and AND3 (N4514, N4488, N2712, N856);
or OR3 (N4515, N4508, N3358, N4095);
buf BUF1 (N4516, N4509);
buf BUF1 (N4517, N4516);
nor NOR3 (N4518, N4502, N454, N718);
buf BUF1 (N4519, N4505);
xor XOR2 (N4520, N4518, N1743);
nor NOR4 (N4521, N4512, N1337, N4094, N3437);
nand NAND2 (N4522, N4510, N3671);
and AND4 (N4523, N4522, N1089, N2009, N448);
not NOT1 (N4524, N4523);
and AND3 (N4525, N4519, N3337, N4298);
or OR2 (N4526, N4521, N4020);
and AND3 (N4527, N4520, N265, N929);
not NOT1 (N4528, N4526);
buf BUF1 (N4529, N4484);
buf BUF1 (N4530, N4517);
nand NAND3 (N4531, N4528, N815, N1587);
nor NOR4 (N4532, N4530, N3906, N31, N4335);
nand NAND2 (N4533, N4529, N4475);
nand NAND4 (N4534, N4524, N872, N171, N1740);
or OR4 (N4535, N4515, N1292, N3737, N3366);
nor NOR2 (N4536, N4525, N2514);
buf BUF1 (N4537, N4536);
nand NAND3 (N4538, N4535, N1763, N2167);
not NOT1 (N4539, N4534);
buf BUF1 (N4540, N4513);
buf BUF1 (N4541, N4527);
nor NOR4 (N4542, N4494, N1296, N3557, N2342);
not NOT1 (N4543, N4537);
buf BUF1 (N4544, N4540);
nor NOR2 (N4545, N4543, N4440);
nand NAND3 (N4546, N4544, N758, N572);
nor NOR3 (N4547, N4538, N3368, N768);
nor NOR2 (N4548, N4533, N483);
or OR4 (N4549, N4531, N3145, N1341, N1677);
and AND4 (N4550, N4545, N3711, N4506, N2069);
and AND2 (N4551, N4539, N3218);
not NOT1 (N4552, N4541);
or OR2 (N4553, N4532, N1910);
or OR3 (N4554, N4550, N488, N3800);
or OR3 (N4555, N4546, N261, N3338);
or OR2 (N4556, N4555, N1606);
nand NAND3 (N4557, N4547, N2201, N428);
or OR2 (N4558, N4553, N409);
buf BUF1 (N4559, N4556);
nand NAND4 (N4560, N4559, N573, N416, N2592);
and AND3 (N4561, N4557, N3924, N420);
or OR4 (N4562, N4561, N446, N3828, N2237);
buf BUF1 (N4563, N4562);
or OR4 (N4564, N4563, N2244, N913, N663);
buf BUF1 (N4565, N4542);
nand NAND3 (N4566, N4548, N2447, N2936);
or OR4 (N4567, N4560, N1767, N344, N723);
nand NAND4 (N4568, N4567, N3138, N2697, N568);
or OR2 (N4569, N4514, N206);
or OR4 (N4570, N4568, N136, N1270, N337);
nand NAND4 (N4571, N4566, N2402, N4386, N2538);
xor XOR2 (N4572, N4569, N4215);
xor XOR2 (N4573, N4565, N633);
nor NOR4 (N4574, N4573, N3712, N4000, N2402);
nor NOR2 (N4575, N4571, N4564);
not NOT1 (N4576, N4479);
and AND2 (N4577, N4574, N3757);
nand NAND3 (N4578, N4576, N504, N765);
xor XOR2 (N4579, N4551, N3705);
nand NAND4 (N4580, N4575, N2507, N1195, N100);
and AND3 (N4581, N4549, N4161, N36);
nand NAND4 (N4582, N4572, N4398, N2954, N3725);
nor NOR4 (N4583, N4580, N4246, N3309, N461);
and AND3 (N4584, N4554, N2490, N1291);
and AND4 (N4585, N4581, N4336, N424, N2811);
nand NAND3 (N4586, N4577, N2265, N4023);
nor NOR3 (N4587, N4582, N2214, N1690);
nor NOR4 (N4588, N4552, N3709, N486, N1624);
nor NOR3 (N4589, N4587, N1879, N4144);
and AND3 (N4590, N4570, N3809, N4144);
not NOT1 (N4591, N4579);
nor NOR4 (N4592, N4578, N3761, N986, N2420);
xor XOR2 (N4593, N4588, N997);
not NOT1 (N4594, N4584);
not NOT1 (N4595, N4592);
nand NAND4 (N4596, N4591, N4426, N2430, N164);
nand NAND3 (N4597, N4595, N133, N2394);
not NOT1 (N4598, N4589);
nand NAND4 (N4599, N4586, N348, N2126, N4010);
and AND3 (N4600, N4599, N3481, N4148);
or OR3 (N4601, N4596, N1651, N2611);
nor NOR3 (N4602, N4590, N3931, N1973);
buf BUF1 (N4603, N4594);
or OR2 (N4604, N4583, N4147);
nand NAND3 (N4605, N4601, N388, N4299);
xor XOR2 (N4606, N4585, N2097);
and AND3 (N4607, N4602, N1009, N348);
and AND2 (N4608, N4600, N2193);
and AND2 (N4609, N4606, N268);
nor NOR3 (N4610, N4603, N3966, N1837);
or OR3 (N4611, N4604, N520, N3261);
buf BUF1 (N4612, N4609);
nand NAND4 (N4613, N4558, N4001, N776, N857);
not NOT1 (N4614, N4610);
nor NOR2 (N4615, N4597, N1152);
nand NAND2 (N4616, N4598, N3065);
nand NAND3 (N4617, N4614, N3269, N837);
xor XOR2 (N4618, N4607, N3936);
and AND3 (N4619, N4593, N1540, N1126);
nand NAND4 (N4620, N4612, N629, N3152, N1422);
nor NOR4 (N4621, N4605, N2426, N4132, N68);
buf BUF1 (N4622, N4613);
and AND2 (N4623, N4616, N148);
xor XOR2 (N4624, N4608, N1189);
or OR3 (N4625, N4617, N2338, N540);
not NOT1 (N4626, N4623);
not NOT1 (N4627, N4615);
not NOT1 (N4628, N4626);
or OR2 (N4629, N4618, N3977);
nor NOR2 (N4630, N4611, N2622);
buf BUF1 (N4631, N4628);
not NOT1 (N4632, N4624);
buf BUF1 (N4633, N4625);
nor NOR4 (N4634, N4627, N4559, N1901, N2505);
not NOT1 (N4635, N4630);
and AND4 (N4636, N4629, N3047, N2079, N4349);
not NOT1 (N4637, N4636);
xor XOR2 (N4638, N4637, N614);
not NOT1 (N4639, N4633);
or OR4 (N4640, N4620, N3426, N3420, N4386);
nand NAND2 (N4641, N4621, N3465);
xor XOR2 (N4642, N4640, N3905);
xor XOR2 (N4643, N4619, N1893);
nor NOR3 (N4644, N4639, N4552, N1675);
nor NOR3 (N4645, N4635, N599, N2457);
not NOT1 (N4646, N4634);
buf BUF1 (N4647, N4642);
and AND3 (N4648, N4647, N701, N2831);
not NOT1 (N4649, N4643);
or OR2 (N4650, N4638, N692);
nor NOR4 (N4651, N4646, N1675, N4642, N2796);
or OR2 (N4652, N4632, N3821);
nand NAND4 (N4653, N4652, N3815, N4248, N2995);
not NOT1 (N4654, N4644);
buf BUF1 (N4655, N4648);
nand NAND4 (N4656, N4655, N4234, N2258, N2921);
buf BUF1 (N4657, N4622);
not NOT1 (N4658, N4651);
nand NAND4 (N4659, N4654, N2588, N2472, N385);
nand NAND4 (N4660, N4641, N4608, N239, N1372);
buf BUF1 (N4661, N4631);
and AND3 (N4662, N4661, N2768, N1337);
xor XOR2 (N4663, N4645, N4324);
nor NOR4 (N4664, N4657, N2840, N54, N4143);
nand NAND2 (N4665, N4658, N1485);
xor XOR2 (N4666, N4665, N4031);
buf BUF1 (N4667, N4659);
or OR2 (N4668, N4664, N1787);
nand NAND3 (N4669, N4656, N752, N2019);
and AND4 (N4670, N4660, N2693, N2262, N3952);
buf BUF1 (N4671, N4649);
and AND4 (N4672, N4653, N4185, N1506, N4627);
not NOT1 (N4673, N4663);
buf BUF1 (N4674, N4671);
not NOT1 (N4675, N4669);
or OR4 (N4676, N4672, N770, N1630, N135);
buf BUF1 (N4677, N4667);
nor NOR4 (N4678, N4676, N3743, N937, N999);
nor NOR4 (N4679, N4666, N3466, N1502, N449);
and AND4 (N4680, N4668, N3852, N107, N647);
nor NOR3 (N4681, N4678, N3006, N693);
and AND2 (N4682, N4680, N4272);
nand NAND2 (N4683, N4674, N345);
not NOT1 (N4684, N4673);
not NOT1 (N4685, N4677);
nand NAND4 (N4686, N4684, N3579, N523, N4248);
or OR2 (N4687, N4686, N2416);
xor XOR2 (N4688, N4675, N2524);
or OR2 (N4689, N4682, N607);
nand NAND4 (N4690, N4662, N2953, N654, N1151);
nor NOR3 (N4691, N4679, N4541, N1094);
nand NAND2 (N4692, N4685, N947);
buf BUF1 (N4693, N4681);
nor NOR3 (N4694, N4690, N1767, N1859);
nand NAND2 (N4695, N4688, N2178);
xor XOR2 (N4696, N4687, N803);
buf BUF1 (N4697, N4694);
nor NOR4 (N4698, N4693, N395, N2488, N4338);
nor NOR3 (N4699, N4698, N2762, N1037);
not NOT1 (N4700, N4683);
nand NAND4 (N4701, N4696, N843, N3682, N514);
not NOT1 (N4702, N4691);
nand NAND4 (N4703, N4702, N2418, N1220, N2007);
nand NAND3 (N4704, N4697, N4249, N4662);
nor NOR3 (N4705, N4692, N2928, N624);
buf BUF1 (N4706, N4705);
nor NOR3 (N4707, N4695, N4134, N1201);
or OR2 (N4708, N4670, N897);
nor NOR2 (N4709, N4707, N1069);
nand NAND2 (N4710, N4703, N1514);
buf BUF1 (N4711, N4708);
not NOT1 (N4712, N4709);
or OR2 (N4713, N4710, N739);
nand NAND2 (N4714, N4704, N1560);
buf BUF1 (N4715, N4712);
or OR2 (N4716, N4714, N4284);
buf BUF1 (N4717, N4711);
nand NAND4 (N4718, N4713, N4533, N1196, N2940);
xor XOR2 (N4719, N4700, N1290);
nand NAND3 (N4720, N4717, N3071, N849);
buf BUF1 (N4721, N4706);
nand NAND4 (N4722, N4716, N3802, N1179, N632);
buf BUF1 (N4723, N4722);
xor XOR2 (N4724, N4718, N2139);
not NOT1 (N4725, N4721);
xor XOR2 (N4726, N4701, N3658);
buf BUF1 (N4727, N4726);
xor XOR2 (N4728, N4725, N639);
nand NAND2 (N4729, N4689, N2744);
and AND2 (N4730, N4727, N4123);
or OR2 (N4731, N4730, N276);
nor NOR3 (N4732, N4720, N4559, N2252);
xor XOR2 (N4733, N4650, N541);
buf BUF1 (N4734, N4724);
nand NAND2 (N4735, N4719, N4008);
and AND2 (N4736, N4715, N3843);
and AND4 (N4737, N4734, N4510, N3611, N1443);
nand NAND4 (N4738, N4699, N1740, N700, N2313);
not NOT1 (N4739, N4732);
xor XOR2 (N4740, N4737, N4309);
xor XOR2 (N4741, N4728, N4574);
xor XOR2 (N4742, N4723, N482);
nand NAND2 (N4743, N4741, N3425);
or OR3 (N4744, N4738, N2726, N3376);
buf BUF1 (N4745, N4739);
xor XOR2 (N4746, N4731, N1097);
xor XOR2 (N4747, N4735, N4395);
and AND3 (N4748, N4740, N4079, N2346);
nand NAND4 (N4749, N4748, N2027, N1098, N2386);
nor NOR2 (N4750, N4747, N391);
and AND4 (N4751, N4736, N380, N2289, N2484);
not NOT1 (N4752, N4733);
buf BUF1 (N4753, N4744);
and AND2 (N4754, N4750, N3055);
xor XOR2 (N4755, N4729, N1736);
xor XOR2 (N4756, N4745, N1374);
xor XOR2 (N4757, N4751, N4369);
xor XOR2 (N4758, N4754, N24);
xor XOR2 (N4759, N4742, N1815);
nor NOR3 (N4760, N4746, N1543, N2195);
not NOT1 (N4761, N4756);
or OR4 (N4762, N4761, N1531, N551, N3808);
not NOT1 (N4763, N4743);
nor NOR3 (N4764, N4758, N2113, N3051);
and AND2 (N4765, N4753, N1952);
nand NAND4 (N4766, N4764, N804, N4223, N3132);
nand NAND4 (N4767, N4749, N3853, N2339, N608);
nor NOR3 (N4768, N4752, N3858, N2972);
or OR4 (N4769, N4762, N1193, N982, N4731);
nor NOR2 (N4770, N4767, N1017);
xor XOR2 (N4771, N4769, N141);
buf BUF1 (N4772, N4770);
or OR4 (N4773, N4759, N29, N4681, N2650);
or OR2 (N4774, N4773, N4291);
buf BUF1 (N4775, N4757);
nand NAND4 (N4776, N4760, N2665, N4368, N4522);
and AND2 (N4777, N4775, N1802);
xor XOR2 (N4778, N4755, N2997);
not NOT1 (N4779, N4763);
and AND4 (N4780, N4765, N1795, N94, N4158);
xor XOR2 (N4781, N4779, N3483);
or OR2 (N4782, N4774, N4560);
or OR4 (N4783, N4782, N759, N4044, N3991);
not NOT1 (N4784, N4778);
xor XOR2 (N4785, N4784, N2795);
nor NOR3 (N4786, N4776, N2930, N4113);
and AND2 (N4787, N4777, N540);
xor XOR2 (N4788, N4785, N3997);
not NOT1 (N4789, N4787);
buf BUF1 (N4790, N4780);
or OR4 (N4791, N4781, N1135, N309, N4544);
not NOT1 (N4792, N4766);
nand NAND2 (N4793, N4783, N801);
nand NAND3 (N4794, N4772, N18, N4584);
buf BUF1 (N4795, N4789);
xor XOR2 (N4796, N4792, N4655);
and AND2 (N4797, N4793, N2128);
and AND2 (N4798, N4795, N567);
not NOT1 (N4799, N4786);
nor NOR3 (N4800, N4798, N4041, N1970);
and AND4 (N4801, N4797, N4199, N4514, N2877);
or OR4 (N4802, N4771, N208, N2522, N3399);
nor NOR2 (N4803, N4791, N3401);
buf BUF1 (N4804, N4790);
buf BUF1 (N4805, N4804);
nor NOR3 (N4806, N4805, N1867, N2055);
nand NAND4 (N4807, N4799, N3343, N3158, N3775);
and AND2 (N4808, N4807, N1260);
and AND4 (N4809, N4801, N3520, N40, N3810);
nor NOR2 (N4810, N4788, N2752);
buf BUF1 (N4811, N4803);
xor XOR2 (N4812, N4810, N2787);
buf BUF1 (N4813, N4800);
xor XOR2 (N4814, N4796, N4207);
and AND3 (N4815, N4811, N1116, N1033);
and AND2 (N4816, N4812, N3554);
nand NAND3 (N4817, N4814, N2633, N2169);
or OR2 (N4818, N4817, N2976);
nand NAND3 (N4819, N4816, N2, N1425);
nand NAND3 (N4820, N4794, N3881, N1735);
not NOT1 (N4821, N4809);
or OR3 (N4822, N4813, N2790, N4035);
not NOT1 (N4823, N4818);
not NOT1 (N4824, N4821);
or OR2 (N4825, N4806, N65);
or OR2 (N4826, N4802, N975);
buf BUF1 (N4827, N4808);
and AND4 (N4828, N4768, N4289, N3422, N2657);
not NOT1 (N4829, N4826);
nand NAND4 (N4830, N4823, N1786, N2702, N1999);
or OR3 (N4831, N4820, N1326, N1460);
buf BUF1 (N4832, N4824);
or OR4 (N4833, N4815, N3307, N361, N1620);
buf BUF1 (N4834, N4829);
and AND4 (N4835, N4819, N1699, N2673, N3826);
nand NAND3 (N4836, N4830, N2771, N4459);
nor NOR4 (N4837, N4827, N975, N2798, N1050);
and AND4 (N4838, N4837, N668, N2557, N1454);
not NOT1 (N4839, N4838);
nor NOR3 (N4840, N4825, N3213, N1705);
not NOT1 (N4841, N4831);
and AND3 (N4842, N4839, N382, N4783);
not NOT1 (N4843, N4822);
or OR4 (N4844, N4834, N1138, N948, N1380);
buf BUF1 (N4845, N4840);
xor XOR2 (N4846, N4843, N572);
not NOT1 (N4847, N4833);
buf BUF1 (N4848, N4836);
not NOT1 (N4849, N4847);
and AND4 (N4850, N4846, N2013, N1049, N3106);
nand NAND4 (N4851, N4849, N362, N443, N1332);
not NOT1 (N4852, N4845);
nand NAND2 (N4853, N4844, N2349);
or OR3 (N4854, N4853, N31, N4729);
or OR3 (N4855, N4852, N707, N89);
not NOT1 (N4856, N4842);
not NOT1 (N4857, N4850);
buf BUF1 (N4858, N4857);
nand NAND3 (N4859, N4856, N1105, N3613);
or OR3 (N4860, N4828, N2043, N2118);
buf BUF1 (N4861, N4860);
not NOT1 (N4862, N4854);
nand NAND2 (N4863, N4861, N2780);
xor XOR2 (N4864, N4841, N2076);
nand NAND3 (N4865, N4835, N4593, N964);
buf BUF1 (N4866, N4848);
xor XOR2 (N4867, N4858, N2517);
nor NOR3 (N4868, N4863, N2523, N1879);
xor XOR2 (N4869, N4851, N658);
nand NAND2 (N4870, N4865, N2183);
xor XOR2 (N4871, N4866, N4317);
xor XOR2 (N4872, N4869, N1754);
nand NAND3 (N4873, N4832, N2985, N1736);
or OR3 (N4874, N4872, N2381, N1739);
or OR4 (N4875, N4873, N665, N223, N1127);
not NOT1 (N4876, N4864);
nor NOR2 (N4877, N4871, N1612);
xor XOR2 (N4878, N4855, N2083);
and AND2 (N4879, N4870, N154);
xor XOR2 (N4880, N4876, N4863);
and AND4 (N4881, N4874, N4445, N2596, N2919);
nor NOR2 (N4882, N4867, N4340);
not NOT1 (N4883, N4882);
and AND4 (N4884, N4883, N1814, N107, N2242);
nor NOR2 (N4885, N4862, N1251);
nor NOR4 (N4886, N4880, N271, N3639, N1056);
not NOT1 (N4887, N4886);
nand NAND4 (N4888, N4881, N4036, N214, N755);
or OR2 (N4889, N4875, N903);
not NOT1 (N4890, N4887);
not NOT1 (N4891, N4877);
not NOT1 (N4892, N4884);
nor NOR4 (N4893, N4892, N1001, N953, N2258);
or OR2 (N4894, N4859, N4786);
xor XOR2 (N4895, N4891, N2243);
buf BUF1 (N4896, N4868);
nor NOR3 (N4897, N4889, N2391, N2109);
and AND3 (N4898, N4896, N3302, N1648);
xor XOR2 (N4899, N4893, N3724);
xor XOR2 (N4900, N4897, N493);
and AND2 (N4901, N4879, N3318);
nor NOR3 (N4902, N4898, N3416, N4107);
buf BUF1 (N4903, N4894);
buf BUF1 (N4904, N4885);
nor NOR2 (N4905, N4903, N2254);
or OR3 (N4906, N4878, N3897, N733);
xor XOR2 (N4907, N4888, N1976);
buf BUF1 (N4908, N4899);
buf BUF1 (N4909, N4905);
or OR3 (N4910, N4909, N1825, N1387);
or OR4 (N4911, N4910, N2247, N976, N3533);
buf BUF1 (N4912, N4900);
buf BUF1 (N4913, N4904);
nor NOR2 (N4914, N4912, N576);
xor XOR2 (N4915, N4911, N3181);
nand NAND3 (N4916, N4890, N3787, N3827);
not NOT1 (N4917, N4913);
nor NOR4 (N4918, N4907, N2741, N214, N2927);
nand NAND4 (N4919, N4915, N1445, N599, N2325);
not NOT1 (N4920, N4914);
and AND3 (N4921, N4895, N3423, N3875);
and AND3 (N4922, N4917, N2857, N1329);
not NOT1 (N4923, N4916);
nor NOR3 (N4924, N4908, N794, N4835);
nand NAND3 (N4925, N4921, N975, N3001);
and AND4 (N4926, N4920, N2225, N3850, N3266);
nand NAND2 (N4927, N4906, N293);
buf BUF1 (N4928, N4925);
and AND4 (N4929, N4902, N373, N144, N353);
nor NOR4 (N4930, N4927, N1168, N3882, N85);
nor NOR4 (N4931, N4901, N1964, N1736, N2525);
buf BUF1 (N4932, N4926);
and AND2 (N4933, N4929, N2967);
xor XOR2 (N4934, N4932, N2818);
and AND4 (N4935, N4934, N1855, N4855, N1228);
buf BUF1 (N4936, N4928);
buf BUF1 (N4937, N4923);
xor XOR2 (N4938, N4933, N276);
and AND2 (N4939, N4937, N3277);
and AND3 (N4940, N4919, N217, N2986);
nor NOR4 (N4941, N4918, N3838, N1981, N190);
buf BUF1 (N4942, N4924);
and AND2 (N4943, N4939, N617);
and AND2 (N4944, N4942, N3287);
nand NAND4 (N4945, N4943, N4426, N352, N1314);
or OR2 (N4946, N4935, N372);
xor XOR2 (N4947, N4944, N2916);
and AND3 (N4948, N4940, N348, N3969);
not NOT1 (N4949, N4938);
or OR2 (N4950, N4936, N93);
or OR2 (N4951, N4922, N2428);
nand NAND3 (N4952, N4931, N2675, N3300);
buf BUF1 (N4953, N4950);
nor NOR2 (N4954, N4946, N1753);
nand NAND3 (N4955, N4930, N373, N3580);
buf BUF1 (N4956, N4952);
xor XOR2 (N4957, N4947, N2553);
buf BUF1 (N4958, N4941);
nand NAND3 (N4959, N4956, N3646, N1569);
xor XOR2 (N4960, N4948, N185);
xor XOR2 (N4961, N4951, N2212);
or OR2 (N4962, N4958, N3821);
and AND3 (N4963, N4954, N484, N4611);
buf BUF1 (N4964, N4961);
nor NOR2 (N4965, N4964, N3029);
or OR3 (N4966, N4962, N4196, N3267);
xor XOR2 (N4967, N4945, N412);
nor NOR2 (N4968, N4949, N2244);
xor XOR2 (N4969, N4957, N2924);
buf BUF1 (N4970, N4968);
xor XOR2 (N4971, N4969, N4826);
nor NOR3 (N4972, N4963, N2674, N2737);
nand NAND4 (N4973, N4965, N4326, N1662, N1160);
buf BUF1 (N4974, N4970);
nand NAND3 (N4975, N4972, N430, N2391);
or OR2 (N4976, N4967, N147);
or OR3 (N4977, N4976, N2592, N2034);
xor XOR2 (N4978, N4966, N407);
xor XOR2 (N4979, N4959, N3340);
buf BUF1 (N4980, N4955);
and AND4 (N4981, N4977, N507, N3631, N316);
not NOT1 (N4982, N4981);
nand NAND2 (N4983, N4979, N2090);
nor NOR3 (N4984, N4971, N3598, N642);
xor XOR2 (N4985, N4983, N565);
nand NAND3 (N4986, N4984, N3095, N3286);
nor NOR2 (N4987, N4975, N2289);
xor XOR2 (N4988, N4986, N4240);
buf BUF1 (N4989, N4988);
xor XOR2 (N4990, N4974, N4269);
not NOT1 (N4991, N4980);
xor XOR2 (N4992, N4982, N4530);
buf BUF1 (N4993, N4992);
and AND3 (N4994, N4960, N1166, N1876);
not NOT1 (N4995, N4978);
or OR4 (N4996, N4994, N4547, N2733, N1213);
nor NOR4 (N4997, N4993, N3438, N1631, N3076);
buf BUF1 (N4998, N4995);
and AND3 (N4999, N4953, N2544, N1033);
nor NOR2 (N5000, N4987, N1938);
or OR3 (N5001, N4996, N3724, N1227);
xor XOR2 (N5002, N4999, N1632);
buf BUF1 (N5003, N5002);
nand NAND4 (N5004, N5001, N1415, N4017, N2870);
xor XOR2 (N5005, N4998, N358);
not NOT1 (N5006, N4991);
buf BUF1 (N5007, N4989);
not NOT1 (N5008, N5004);
and AND2 (N5009, N5003, N1068);
or OR2 (N5010, N5000, N3757);
nor NOR2 (N5011, N5006, N2053);
nor NOR4 (N5012, N4973, N1610, N3957, N979);
xor XOR2 (N5013, N5007, N1441);
xor XOR2 (N5014, N5009, N3074);
not NOT1 (N5015, N4990);
nor NOR4 (N5016, N5014, N2416, N2694, N4058);
buf BUF1 (N5017, N5015);
xor XOR2 (N5018, N5008, N545);
and AND4 (N5019, N5010, N2803, N4747, N4305);
xor XOR2 (N5020, N4985, N1990);
xor XOR2 (N5021, N5016, N1719);
nand NAND3 (N5022, N5012, N4293, N3615);
and AND4 (N5023, N5005, N3707, N3442, N4351);
nor NOR2 (N5024, N5019, N4130);
or OR3 (N5025, N5011, N3958, N944);
xor XOR2 (N5026, N5021, N596);
not NOT1 (N5027, N5024);
nor NOR4 (N5028, N4997, N4223, N253, N873);
xor XOR2 (N5029, N5025, N1617);
and AND3 (N5030, N5017, N3304, N3329);
xor XOR2 (N5031, N5013, N643);
xor XOR2 (N5032, N5029, N2677);
and AND4 (N5033, N5030, N1932, N2709, N3372);
nor NOR2 (N5034, N5032, N3778);
xor XOR2 (N5035, N5018, N4978);
xor XOR2 (N5036, N5034, N576);
and AND3 (N5037, N5035, N3860, N1237);
and AND2 (N5038, N5022, N2111);
nand NAND2 (N5039, N5033, N2429);
nand NAND2 (N5040, N5027, N1342);
xor XOR2 (N5041, N5038, N4024);
buf BUF1 (N5042, N5037);
nand NAND3 (N5043, N5040, N1761, N2816);
or OR3 (N5044, N5026, N2645, N1269);
and AND4 (N5045, N5044, N404, N3136, N2320);
buf BUF1 (N5046, N5020);
or OR3 (N5047, N5031, N4133, N857);
nor NOR2 (N5048, N5047, N130);
xor XOR2 (N5049, N5046, N1241);
buf BUF1 (N5050, N5023);
and AND2 (N5051, N5043, N702);
not NOT1 (N5052, N5036);
not NOT1 (N5053, N5049);
buf BUF1 (N5054, N5051);
buf BUF1 (N5055, N5053);
nand NAND4 (N5056, N5054, N1184, N1257, N2669);
and AND2 (N5057, N5052, N2766);
xor XOR2 (N5058, N5042, N3467);
not NOT1 (N5059, N5057);
not NOT1 (N5060, N5048);
nor NOR3 (N5061, N5055, N3935, N185);
not NOT1 (N5062, N5045);
not NOT1 (N5063, N5059);
or OR3 (N5064, N5061, N2002, N3058);
nand NAND3 (N5065, N5062, N1692, N541);
or OR2 (N5066, N5041, N3674);
buf BUF1 (N5067, N5028);
and AND3 (N5068, N5039, N1843, N608);
not NOT1 (N5069, N5068);
and AND4 (N5070, N5069, N2644, N3400, N3040);
nor NOR3 (N5071, N5070, N3345, N4317);
and AND4 (N5072, N5050, N2564, N2338, N828);
xor XOR2 (N5073, N5072, N246);
and AND3 (N5074, N5060, N2402, N4869);
xor XOR2 (N5075, N5066, N3723);
and AND3 (N5076, N5063, N1206, N1501);
not NOT1 (N5077, N5075);
nor NOR4 (N5078, N5064, N2117, N2313, N4110);
xor XOR2 (N5079, N5067, N2590);
or OR2 (N5080, N5056, N1799);
buf BUF1 (N5081, N5071);
and AND2 (N5082, N5065, N2898);
nor NOR2 (N5083, N5074, N3534);
or OR2 (N5084, N5082, N1079);
xor XOR2 (N5085, N5077, N4615);
buf BUF1 (N5086, N5083);
nand NAND4 (N5087, N5085, N792, N3674, N2789);
nand NAND2 (N5088, N5076, N3169);
nand NAND3 (N5089, N5078, N1784, N2853);
and AND3 (N5090, N5089, N1375, N1172);
nand NAND4 (N5091, N5084, N2367, N2261, N3434);
xor XOR2 (N5092, N5081, N3695);
nor NOR3 (N5093, N5073, N283, N2651);
xor XOR2 (N5094, N5093, N1807);
not NOT1 (N5095, N5094);
xor XOR2 (N5096, N5095, N4276);
nor NOR4 (N5097, N5058, N4886, N3304, N4835);
nor NOR4 (N5098, N5087, N5027, N4950, N3924);
not NOT1 (N5099, N5091);
xor XOR2 (N5100, N5098, N4955);
nor NOR3 (N5101, N5079, N1909, N1853);
and AND2 (N5102, N5080, N170);
nor NOR2 (N5103, N5086, N2160);
nor NOR3 (N5104, N5097, N737, N1982);
xor XOR2 (N5105, N5102, N2594);
not NOT1 (N5106, N5088);
not NOT1 (N5107, N5090);
or OR3 (N5108, N5101, N3393, N2977);
nor NOR3 (N5109, N5099, N982, N4991);
not NOT1 (N5110, N5103);
buf BUF1 (N5111, N5109);
and AND3 (N5112, N5092, N2669, N1207);
buf BUF1 (N5113, N5108);
not NOT1 (N5114, N5104);
or OR2 (N5115, N5096, N4303);
xor XOR2 (N5116, N5105, N1823);
xor XOR2 (N5117, N5115, N442);
xor XOR2 (N5118, N5100, N550);
buf BUF1 (N5119, N5110);
nand NAND4 (N5120, N5112, N2861, N1884, N1372);
or OR2 (N5121, N5120, N1452);
xor XOR2 (N5122, N5116, N2105);
nand NAND3 (N5123, N5119, N624, N1482);
xor XOR2 (N5124, N5106, N2143);
buf BUF1 (N5125, N5121);
or OR4 (N5126, N5124, N3345, N3494, N125);
xor XOR2 (N5127, N5117, N2659);
buf BUF1 (N5128, N5118);
nand NAND2 (N5129, N5127, N5001);
not NOT1 (N5130, N5111);
xor XOR2 (N5131, N5128, N3682);
not NOT1 (N5132, N5130);
or OR3 (N5133, N5122, N350, N3460);
buf BUF1 (N5134, N5114);
nor NOR2 (N5135, N5126, N2093);
nand NAND3 (N5136, N5113, N4911, N4100);
xor XOR2 (N5137, N5136, N847);
not NOT1 (N5138, N5123);
not NOT1 (N5139, N5129);
not NOT1 (N5140, N5137);
buf BUF1 (N5141, N5133);
or OR2 (N5142, N5107, N4424);
xor XOR2 (N5143, N5132, N1404);
nor NOR2 (N5144, N5143, N2616);
not NOT1 (N5145, N5141);
xor XOR2 (N5146, N5142, N4429);
and AND2 (N5147, N5146, N1720);
buf BUF1 (N5148, N5125);
or OR3 (N5149, N5148, N2300, N925);
nor NOR3 (N5150, N5149, N1583, N1218);
nand NAND4 (N5151, N5138, N183, N284, N307);
not NOT1 (N5152, N5140);
xor XOR2 (N5153, N5134, N631);
buf BUF1 (N5154, N5152);
nand NAND2 (N5155, N5153, N4575);
xor XOR2 (N5156, N5131, N5148);
buf BUF1 (N5157, N5139);
nand NAND3 (N5158, N5151, N490, N1023);
not NOT1 (N5159, N5158);
and AND3 (N5160, N5135, N4522, N125);
not NOT1 (N5161, N5150);
or OR2 (N5162, N5161, N2378);
or OR2 (N5163, N5156, N2784);
nand NAND4 (N5164, N5157, N5161, N1722, N2859);
and AND3 (N5165, N5155, N1497, N906);
nor NOR3 (N5166, N5154, N6, N533);
nand NAND2 (N5167, N5163, N2536);
or OR2 (N5168, N5167, N958);
not NOT1 (N5169, N5144);
buf BUF1 (N5170, N5168);
nand NAND2 (N5171, N5165, N4038);
or OR4 (N5172, N5169, N2603, N679, N3617);
or OR3 (N5173, N5147, N768, N4806);
xor XOR2 (N5174, N5166, N2698);
nor NOR4 (N5175, N5171, N873, N1703, N278);
buf BUF1 (N5176, N5160);
xor XOR2 (N5177, N5174, N1138);
nor NOR2 (N5178, N5173, N2262);
buf BUF1 (N5179, N5159);
buf BUF1 (N5180, N5145);
nor NOR3 (N5181, N5180, N4346, N2569);
nand NAND3 (N5182, N5170, N2206, N1714);
xor XOR2 (N5183, N5162, N5063);
xor XOR2 (N5184, N5182, N2934);
nor NOR4 (N5185, N5177, N3184, N4596, N894);
and AND2 (N5186, N5164, N2856);
buf BUF1 (N5187, N5181);
and AND2 (N5188, N5176, N3966);
nor NOR2 (N5189, N5183, N1121);
not NOT1 (N5190, N5175);
xor XOR2 (N5191, N5179, N3539);
nand NAND2 (N5192, N5185, N3347);
nand NAND2 (N5193, N5187, N2126);
xor XOR2 (N5194, N5188, N1004);
xor XOR2 (N5195, N5192, N4332);
and AND3 (N5196, N5191, N2957, N4457);
not NOT1 (N5197, N5195);
xor XOR2 (N5198, N5184, N4696);
nor NOR2 (N5199, N5196, N2957);
not NOT1 (N5200, N5186);
or OR3 (N5201, N5200, N643, N2868);
nand NAND4 (N5202, N5198, N1427, N3219, N1323);
and AND2 (N5203, N5193, N3976);
not NOT1 (N5204, N5203);
or OR4 (N5205, N5189, N4068, N1641, N926);
or OR2 (N5206, N5202, N578);
and AND3 (N5207, N5197, N610, N359);
or OR4 (N5208, N5204, N656, N4667, N2175);
or OR3 (N5209, N5206, N1856, N1804);
nor NOR2 (N5210, N5194, N562);
nor NOR2 (N5211, N5172, N764);
xor XOR2 (N5212, N5190, N733);
xor XOR2 (N5213, N5207, N314);
or OR3 (N5214, N5213, N3051, N236);
nor NOR2 (N5215, N5178, N3459);
and AND4 (N5216, N5215, N3253, N1829, N3870);
or OR4 (N5217, N5209, N3144, N2900, N2133);
or OR4 (N5218, N5216, N279, N2673, N1551);
or OR2 (N5219, N5218, N3744);
nand NAND4 (N5220, N5212, N4437, N2788, N3132);
and AND3 (N5221, N5211, N602, N2615);
and AND3 (N5222, N5220, N2845, N4752);
or OR2 (N5223, N5222, N2877);
buf BUF1 (N5224, N5201);
xor XOR2 (N5225, N5217, N3211);
nor NOR4 (N5226, N5205, N3694, N3440, N3152);
buf BUF1 (N5227, N5208);
and AND2 (N5228, N5227, N3057);
nand NAND4 (N5229, N5214, N4767, N3304, N960);
and AND4 (N5230, N5199, N4629, N3842, N4338);
or OR4 (N5231, N5224, N3815, N4571, N4098);
nor NOR4 (N5232, N5226, N3247, N773, N4435);
or OR2 (N5233, N5223, N2141);
buf BUF1 (N5234, N5225);
nand NAND3 (N5235, N5229, N3034, N5179);
not NOT1 (N5236, N5233);
or OR4 (N5237, N5234, N4977, N2912, N1372);
xor XOR2 (N5238, N5232, N3477);
nand NAND4 (N5239, N5236, N4564, N697, N1500);
nand NAND4 (N5240, N5228, N2526, N1833, N625);
nor NOR3 (N5241, N5235, N2756, N2183);
nand NAND2 (N5242, N5237, N638);
nand NAND4 (N5243, N5210, N2498, N3286, N2179);
nor NOR4 (N5244, N5239, N4379, N3037, N4646);
nor NOR4 (N5245, N5230, N1249, N480, N981);
xor XOR2 (N5246, N5231, N3759);
buf BUF1 (N5247, N5243);
nor NOR3 (N5248, N5238, N1349, N3956);
and AND3 (N5249, N5240, N3461, N4008);
not NOT1 (N5250, N5221);
and AND3 (N5251, N5246, N1595, N1008);
and AND2 (N5252, N5250, N948);
or OR2 (N5253, N5252, N2964);
or OR4 (N5254, N5245, N2073, N1932, N302);
not NOT1 (N5255, N5249);
and AND4 (N5256, N5253, N3486, N3372, N3863);
and AND3 (N5257, N5219, N1577, N3722);
nor NOR3 (N5258, N5251, N1100, N2722);
and AND4 (N5259, N5248, N528, N2989, N1263);
nor NOR2 (N5260, N5259, N3291);
and AND3 (N5261, N5255, N976, N2245);
xor XOR2 (N5262, N5254, N3269);
or OR3 (N5263, N5247, N794, N559);
or OR3 (N5264, N5242, N2423, N4871);
not NOT1 (N5265, N5244);
or OR4 (N5266, N5261, N4875, N4910, N874);
xor XOR2 (N5267, N5258, N961);
or OR3 (N5268, N5266, N2254, N754);
or OR3 (N5269, N5265, N1124, N2778);
nor NOR4 (N5270, N5260, N4954, N5233, N4866);
and AND3 (N5271, N5262, N2153, N632);
nand NAND4 (N5272, N5270, N3832, N3075, N4790);
and AND3 (N5273, N5241, N3899, N1430);
xor XOR2 (N5274, N5267, N3230);
xor XOR2 (N5275, N5271, N220);
and AND4 (N5276, N5263, N4415, N2955, N3212);
buf BUF1 (N5277, N5276);
xor XOR2 (N5278, N5275, N1258);
buf BUF1 (N5279, N5277);
xor XOR2 (N5280, N5268, N2353);
xor XOR2 (N5281, N5257, N4346);
or OR3 (N5282, N5279, N1089, N5280);
or OR2 (N5283, N3905, N2220);
xor XOR2 (N5284, N5274, N1826);
xor XOR2 (N5285, N5278, N5004);
nand NAND2 (N5286, N5273, N4876);
and AND2 (N5287, N5283, N1038);
nor NOR2 (N5288, N5256, N3635);
xor XOR2 (N5289, N5269, N1178);
nand NAND2 (N5290, N5272, N5140);
and AND4 (N5291, N5286, N77, N293, N5134);
nand NAND4 (N5292, N5287, N2768, N3222, N3827);
nand NAND3 (N5293, N5289, N4885, N2682);
xor XOR2 (N5294, N5264, N2471);
or OR3 (N5295, N5292, N2425, N3473);
nand NAND4 (N5296, N5284, N1079, N1068, N5013);
or OR4 (N5297, N5285, N5254, N2350, N1870);
and AND4 (N5298, N5290, N4360, N2171, N4086);
and AND4 (N5299, N5298, N4447, N1248, N1865);
nand NAND3 (N5300, N5293, N4393, N3726);
and AND3 (N5301, N5296, N1629, N2418);
and AND2 (N5302, N5291, N3572);
and AND2 (N5303, N5297, N5195);
buf BUF1 (N5304, N5301);
and AND2 (N5305, N5300, N2902);
or OR4 (N5306, N5295, N2544, N2565, N1168);
buf BUF1 (N5307, N5302);
xor XOR2 (N5308, N5294, N1983);
and AND3 (N5309, N5307, N4760, N1525);
and AND2 (N5310, N5281, N4356);
or OR2 (N5311, N5305, N4261);
or OR3 (N5312, N5288, N40, N2386);
nand NAND2 (N5313, N5308, N401);
nand NAND3 (N5314, N5282, N720, N4996);
xor XOR2 (N5315, N5304, N3850);
and AND4 (N5316, N5303, N2888, N5166, N1324);
xor XOR2 (N5317, N5309, N1534);
nor NOR2 (N5318, N5310, N2151);
and AND3 (N5319, N5312, N1825, N4681);
buf BUF1 (N5320, N5313);
and AND2 (N5321, N5299, N1833);
nor NOR4 (N5322, N5316, N1184, N561, N1994);
and AND4 (N5323, N5317, N4115, N1008, N2089);
and AND2 (N5324, N5320, N1420);
nand NAND2 (N5325, N5311, N4435);
xor XOR2 (N5326, N5322, N4401);
xor XOR2 (N5327, N5315, N3232);
buf BUF1 (N5328, N5306);
or OR4 (N5329, N5327, N667, N5320, N4406);
buf BUF1 (N5330, N5323);
buf BUF1 (N5331, N5329);
nand NAND2 (N5332, N5328, N3346);
not NOT1 (N5333, N5324);
or OR4 (N5334, N5325, N658, N5138, N1398);
nand NAND2 (N5335, N5332, N4604);
nor NOR3 (N5336, N5319, N4135, N3368);
and AND4 (N5337, N5334, N2353, N862, N2715);
or OR3 (N5338, N5333, N1894, N5024);
xor XOR2 (N5339, N5338, N201);
not NOT1 (N5340, N5337);
buf BUF1 (N5341, N5331);
and AND2 (N5342, N5314, N4677);
nand NAND3 (N5343, N5340, N1, N135);
nor NOR3 (N5344, N5321, N2594, N367);
nand NAND3 (N5345, N5335, N3322, N3620);
nand NAND4 (N5346, N5326, N5291, N4991, N2089);
and AND3 (N5347, N5341, N722, N4587);
not NOT1 (N5348, N5339);
or OR3 (N5349, N5348, N1398, N1680);
or OR4 (N5350, N5343, N3181, N5051, N1764);
not NOT1 (N5351, N5330);
nand NAND3 (N5352, N5350, N3100, N4440);
xor XOR2 (N5353, N5352, N1558);
xor XOR2 (N5354, N5344, N4660);
or OR3 (N5355, N5342, N2621, N4014);
nor NOR2 (N5356, N5354, N4804);
or OR3 (N5357, N5351, N940, N4911);
xor XOR2 (N5358, N5347, N491);
and AND3 (N5359, N5336, N4351, N652);
not NOT1 (N5360, N5353);
nand NAND4 (N5361, N5356, N1304, N1003, N5294);
xor XOR2 (N5362, N5359, N2225);
or OR2 (N5363, N5361, N5026);
xor XOR2 (N5364, N5357, N4911);
and AND3 (N5365, N5363, N3558, N847);
xor XOR2 (N5366, N5365, N4773);
nand NAND2 (N5367, N5364, N2584);
nand NAND3 (N5368, N5355, N1089, N383);
buf BUF1 (N5369, N5318);
xor XOR2 (N5370, N5358, N4122);
nand NAND4 (N5371, N5360, N3504, N3722, N2412);
not NOT1 (N5372, N5345);
or OR3 (N5373, N5349, N4872, N1707);
nand NAND4 (N5374, N5368, N1334, N729, N3876);
or OR2 (N5375, N5372, N2366);
or OR2 (N5376, N5367, N131);
not NOT1 (N5377, N5370);
nand NAND3 (N5378, N5377, N2073, N5216);
buf BUF1 (N5379, N5376);
nand NAND2 (N5380, N5374, N3794);
nor NOR3 (N5381, N5362, N1334, N822);
nor NOR4 (N5382, N5380, N2736, N4777, N3647);
buf BUF1 (N5383, N5379);
and AND2 (N5384, N5378, N4542);
nand NAND3 (N5385, N5383, N4438, N2817);
nand NAND4 (N5386, N5371, N734, N2180, N3725);
buf BUF1 (N5387, N5369);
not NOT1 (N5388, N5375);
and AND4 (N5389, N5387, N378, N914, N3689);
not NOT1 (N5390, N5381);
buf BUF1 (N5391, N5385);
nand NAND2 (N5392, N5390, N1477);
nand NAND2 (N5393, N5346, N4279);
and AND3 (N5394, N5382, N4430, N742);
nor NOR3 (N5395, N5392, N2472, N5306);
buf BUF1 (N5396, N5394);
or OR2 (N5397, N5391, N4327);
not NOT1 (N5398, N5393);
xor XOR2 (N5399, N5373, N2001);
and AND4 (N5400, N5366, N5081, N1260, N1659);
and AND2 (N5401, N5388, N4763);
buf BUF1 (N5402, N5399);
nor NOR3 (N5403, N5397, N1939, N699);
buf BUF1 (N5404, N5402);
xor XOR2 (N5405, N5398, N435);
nor NOR4 (N5406, N5395, N4165, N2665, N1786);
xor XOR2 (N5407, N5400, N3658);
nor NOR4 (N5408, N5406, N883, N3731, N3186);
xor XOR2 (N5409, N5384, N4949);
buf BUF1 (N5410, N5401);
xor XOR2 (N5411, N5396, N1803);
and AND4 (N5412, N5389, N4672, N1767, N2733);
buf BUF1 (N5413, N5408);
nor NOR3 (N5414, N5412, N1966, N4376);
and AND3 (N5415, N5411, N1752, N2663);
or OR4 (N5416, N5414, N4666, N1764, N590);
xor XOR2 (N5417, N5410, N3880);
buf BUF1 (N5418, N5415);
buf BUF1 (N5419, N5409);
nor NOR4 (N5420, N5405, N2140, N3779, N8);
nand NAND4 (N5421, N5419, N126, N2937, N1997);
and AND3 (N5422, N5413, N851, N2635);
not NOT1 (N5423, N5418);
nor NOR3 (N5424, N5403, N1168, N5251);
and AND3 (N5425, N5416, N81, N4489);
nand NAND2 (N5426, N5425, N3522);
nand NAND3 (N5427, N5420, N371, N5395);
nor NOR2 (N5428, N5423, N1920);
buf BUF1 (N5429, N5424);
nand NAND2 (N5430, N5421, N435);
and AND2 (N5431, N5422, N5184);
xor XOR2 (N5432, N5430, N5382);
nor NOR4 (N5433, N5429, N1519, N5170, N436);
and AND2 (N5434, N5432, N3929);
or OR2 (N5435, N5426, N4687);
xor XOR2 (N5436, N5428, N3819);
not NOT1 (N5437, N5435);
and AND3 (N5438, N5417, N119, N1070);
buf BUF1 (N5439, N5404);
buf BUF1 (N5440, N5436);
xor XOR2 (N5441, N5433, N4008);
xor XOR2 (N5442, N5427, N5352);
buf BUF1 (N5443, N5438);
or OR3 (N5444, N5443, N2685, N4214);
nor NOR2 (N5445, N5440, N4782);
nor NOR3 (N5446, N5434, N1664, N1144);
not NOT1 (N5447, N5439);
buf BUF1 (N5448, N5442);
nand NAND2 (N5449, N5448, N471);
buf BUF1 (N5450, N5446);
nor NOR4 (N5451, N5450, N4858, N4531, N1098);
or OR4 (N5452, N5386, N2057, N3459, N434);
and AND3 (N5453, N5441, N1299, N3572);
xor XOR2 (N5454, N5407, N3722);
and AND2 (N5455, N5447, N5234);
nor NOR3 (N5456, N5437, N3865, N3435);
or OR3 (N5457, N5449, N1003, N2358);
buf BUF1 (N5458, N5444);
not NOT1 (N5459, N5455);
nand NAND4 (N5460, N5457, N4569, N1879, N1125);
not NOT1 (N5461, N5460);
and AND2 (N5462, N5454, N2714);
nor NOR4 (N5463, N5453, N4617, N2352, N5011);
and AND2 (N5464, N5456, N577);
nor NOR3 (N5465, N5452, N4632, N3301);
or OR4 (N5466, N5459, N3831, N1958, N5364);
buf BUF1 (N5467, N5431);
xor XOR2 (N5468, N5465, N1894);
nor NOR2 (N5469, N5468, N2878);
nor NOR4 (N5470, N5467, N1662, N810, N4634);
nor NOR2 (N5471, N5466, N3621);
not NOT1 (N5472, N5469);
and AND2 (N5473, N5463, N180);
nor NOR4 (N5474, N5451, N3597, N4074, N2523);
nor NOR2 (N5475, N5445, N4967);
and AND2 (N5476, N5458, N2947);
xor XOR2 (N5477, N5473, N2114);
and AND2 (N5478, N5462, N4475);
xor XOR2 (N5479, N5476, N1181);
not NOT1 (N5480, N5479);
xor XOR2 (N5481, N5474, N1329);
buf BUF1 (N5482, N5477);
xor XOR2 (N5483, N5478, N3851);
nand NAND2 (N5484, N5471, N5209);
not NOT1 (N5485, N5475);
buf BUF1 (N5486, N5485);
buf BUF1 (N5487, N5470);
buf BUF1 (N5488, N5487);
or OR3 (N5489, N5484, N5052, N2626);
buf BUF1 (N5490, N5489);
xor XOR2 (N5491, N5472, N2509);
buf BUF1 (N5492, N5486);
nor NOR2 (N5493, N5480, N868);
xor XOR2 (N5494, N5483, N310);
not NOT1 (N5495, N5493);
and AND2 (N5496, N5488, N3226);
buf BUF1 (N5497, N5494);
nor NOR2 (N5498, N5491, N1802);
xor XOR2 (N5499, N5482, N5144);
nor NOR3 (N5500, N5497, N1245, N671);
xor XOR2 (N5501, N5499, N3300);
and AND2 (N5502, N5500, N910);
and AND4 (N5503, N5492, N200, N957, N4459);
and AND2 (N5504, N5496, N3282);
xor XOR2 (N5505, N5461, N979);
xor XOR2 (N5506, N5495, N4259);
xor XOR2 (N5507, N5504, N5216);
nor NOR4 (N5508, N5505, N1924, N1894, N5185);
and AND2 (N5509, N5506, N2713);
and AND4 (N5510, N5502, N87, N3539, N3690);
nand NAND2 (N5511, N5501, N2028);
not NOT1 (N5512, N5509);
xor XOR2 (N5513, N5503, N1581);
and AND4 (N5514, N5510, N2527, N1605, N2812);
xor XOR2 (N5515, N5507, N4615);
nand NAND4 (N5516, N5481, N1796, N2541, N3452);
xor XOR2 (N5517, N5513, N4258);
and AND2 (N5518, N5516, N5372);
not NOT1 (N5519, N5514);
buf BUF1 (N5520, N5519);
xor XOR2 (N5521, N5508, N3054);
xor XOR2 (N5522, N5498, N2243);
nor NOR4 (N5523, N5511, N2743, N4609, N3792);
xor XOR2 (N5524, N5517, N2877);
nor NOR3 (N5525, N5464, N5224, N5409);
or OR4 (N5526, N5523, N1502, N3080, N2506);
or OR3 (N5527, N5521, N1657, N3732);
nor NOR4 (N5528, N5525, N4656, N4545, N1351);
nand NAND4 (N5529, N5527, N491, N5011, N4575);
and AND2 (N5530, N5515, N5345);
nor NOR2 (N5531, N5526, N1322);
not NOT1 (N5532, N5512);
xor XOR2 (N5533, N5524, N2186);
buf BUF1 (N5534, N5532);
nor NOR3 (N5535, N5530, N3893, N1408);
buf BUF1 (N5536, N5533);
nand NAND3 (N5537, N5490, N4269, N618);
and AND4 (N5538, N5531, N4547, N5516, N940);
or OR2 (N5539, N5536, N385);
and AND4 (N5540, N5534, N2019, N3938, N4827);
not NOT1 (N5541, N5535);
nand NAND3 (N5542, N5539, N2201, N2956);
nor NOR2 (N5543, N5529, N291);
nor NOR4 (N5544, N5541, N4689, N1182, N1592);
xor XOR2 (N5545, N5537, N4748);
or OR3 (N5546, N5520, N282, N1403);
not NOT1 (N5547, N5518);
or OR2 (N5548, N5546, N5269);
or OR2 (N5549, N5542, N1482);
nand NAND3 (N5550, N5545, N1885, N2119);
nor NOR3 (N5551, N5540, N3963, N4907);
or OR3 (N5552, N5548, N4147, N4405);
or OR4 (N5553, N5550, N2825, N5315, N2643);
buf BUF1 (N5554, N5522);
or OR3 (N5555, N5553, N5295, N3671);
buf BUF1 (N5556, N5544);
and AND4 (N5557, N5543, N1883, N1347, N5291);
and AND3 (N5558, N5551, N1308, N2242);
and AND3 (N5559, N5554, N3985, N5419);
not NOT1 (N5560, N5549);
and AND4 (N5561, N5557, N4791, N4718, N1039);
not NOT1 (N5562, N5560);
xor XOR2 (N5563, N5559, N4681);
nor NOR2 (N5564, N5558, N2508);
buf BUF1 (N5565, N5563);
not NOT1 (N5566, N5555);
nor NOR2 (N5567, N5538, N4167);
nor NOR3 (N5568, N5561, N1603, N4491);
nor NOR3 (N5569, N5564, N3951, N2753);
and AND2 (N5570, N5562, N2068);
and AND2 (N5571, N5570, N1128);
buf BUF1 (N5572, N5571);
not NOT1 (N5573, N5568);
buf BUF1 (N5574, N5569);
xor XOR2 (N5575, N5572, N4611);
buf BUF1 (N5576, N5547);
xor XOR2 (N5577, N5565, N5261);
nor NOR3 (N5578, N5556, N869, N696);
and AND2 (N5579, N5574, N4444);
or OR2 (N5580, N5573, N252);
nand NAND4 (N5581, N5552, N4998, N522, N1802);
xor XOR2 (N5582, N5579, N5446);
buf BUF1 (N5583, N5576);
not NOT1 (N5584, N5580);
not NOT1 (N5585, N5577);
buf BUF1 (N5586, N5584);
not NOT1 (N5587, N5582);
or OR3 (N5588, N5587, N5286, N1435);
not NOT1 (N5589, N5588);
and AND2 (N5590, N5578, N5067);
buf BUF1 (N5591, N5581);
or OR4 (N5592, N5586, N336, N945, N886);
or OR4 (N5593, N5583, N2400, N2271, N962);
buf BUF1 (N5594, N5591);
and AND2 (N5595, N5567, N3685);
buf BUF1 (N5596, N5566);
not NOT1 (N5597, N5594);
nand NAND3 (N5598, N5596, N3131, N1002);
nand NAND2 (N5599, N5593, N3918);
nand NAND4 (N5600, N5592, N4988, N1711, N5175);
nor NOR2 (N5601, N5595, N4348);
or OR3 (N5602, N5585, N4395, N4496);
nor NOR3 (N5603, N5598, N4091, N5168);
xor XOR2 (N5604, N5597, N2930);
not NOT1 (N5605, N5528);
xor XOR2 (N5606, N5589, N1958);
buf BUF1 (N5607, N5605);
nor NOR4 (N5608, N5575, N1557, N3259, N2413);
nand NAND4 (N5609, N5603, N5207, N2530, N5372);
buf BUF1 (N5610, N5599);
nor NOR2 (N5611, N5610, N2956);
or OR2 (N5612, N5609, N2808);
nand NAND2 (N5613, N5604, N2073);
xor XOR2 (N5614, N5608, N794);
xor XOR2 (N5615, N5611, N3427);
not NOT1 (N5616, N5601);
nor NOR4 (N5617, N5615, N3392, N1869, N1542);
nor NOR3 (N5618, N5590, N2345, N1176);
xor XOR2 (N5619, N5618, N1829);
buf BUF1 (N5620, N5606);
and AND3 (N5621, N5614, N3524, N4955);
not NOT1 (N5622, N5607);
nand NAND2 (N5623, N5616, N1573);
nor NOR3 (N5624, N5622, N5041, N4831);
not NOT1 (N5625, N5600);
nor NOR2 (N5626, N5619, N2789);
not NOT1 (N5627, N5625);
not NOT1 (N5628, N5602);
xor XOR2 (N5629, N5617, N3586);
xor XOR2 (N5630, N5623, N4787);
not NOT1 (N5631, N5612);
nand NAND2 (N5632, N5627, N1960);
or OR2 (N5633, N5631, N1155);
nand NAND4 (N5634, N5613, N3636, N5509, N2200);
not NOT1 (N5635, N5634);
not NOT1 (N5636, N5621);
nand NAND2 (N5637, N5633, N2795);
or OR2 (N5638, N5632, N1627);
nand NAND2 (N5639, N5626, N4945);
not NOT1 (N5640, N5624);
xor XOR2 (N5641, N5636, N899);
not NOT1 (N5642, N5620);
and AND3 (N5643, N5639, N3620, N1657);
buf BUF1 (N5644, N5643);
nor NOR2 (N5645, N5630, N165);
or OR4 (N5646, N5642, N5021, N1987, N2989);
nand NAND4 (N5647, N5637, N3462, N3464, N3130);
xor XOR2 (N5648, N5644, N1013);
buf BUF1 (N5649, N5646);
nand NAND4 (N5650, N5635, N4484, N2945, N1044);
nand NAND3 (N5651, N5647, N2316, N3990);
and AND2 (N5652, N5628, N1848);
xor XOR2 (N5653, N5645, N275);
nor NOR2 (N5654, N5629, N5367);
not NOT1 (N5655, N5640);
buf BUF1 (N5656, N5650);
nand NAND2 (N5657, N5654, N6);
nand NAND4 (N5658, N5656, N2693, N3158, N999);
not NOT1 (N5659, N5649);
or OR2 (N5660, N5651, N3433);
and AND4 (N5661, N5641, N4014, N4833, N2204);
buf BUF1 (N5662, N5653);
nor NOR3 (N5663, N5659, N904, N1871);
nor NOR2 (N5664, N5661, N5597);
xor XOR2 (N5665, N5652, N5531);
not NOT1 (N5666, N5662);
buf BUF1 (N5667, N5658);
not NOT1 (N5668, N5655);
buf BUF1 (N5669, N5657);
nand NAND4 (N5670, N5638, N2464, N4948, N1920);
and AND3 (N5671, N5648, N3918, N5475);
or OR4 (N5672, N5671, N628, N2629, N4497);
or OR3 (N5673, N5670, N2096, N2745);
or OR4 (N5674, N5672, N5338, N3205, N646);
xor XOR2 (N5675, N5669, N2467);
xor XOR2 (N5676, N5660, N4766);
buf BUF1 (N5677, N5664);
xor XOR2 (N5678, N5668, N3110);
xor XOR2 (N5679, N5676, N2817);
or OR2 (N5680, N5666, N924);
nand NAND3 (N5681, N5677, N5049, N1039);
or OR2 (N5682, N5679, N2117);
not NOT1 (N5683, N5674);
nor NOR2 (N5684, N5680, N2425);
xor XOR2 (N5685, N5675, N4578);
and AND4 (N5686, N5665, N2802, N5273, N1781);
buf BUF1 (N5687, N5678);
nand NAND2 (N5688, N5663, N2920);
or OR4 (N5689, N5682, N1085, N3532, N1177);
nor NOR4 (N5690, N5684, N4358, N2573, N3468);
xor XOR2 (N5691, N5683, N2705);
xor XOR2 (N5692, N5667, N560);
nand NAND4 (N5693, N5686, N2723, N1802, N3651);
or OR3 (N5694, N5693, N167, N2019);
or OR2 (N5695, N5681, N3430);
nand NAND2 (N5696, N5692, N1779);
and AND2 (N5697, N5695, N5222);
xor XOR2 (N5698, N5697, N23);
nor NOR2 (N5699, N5687, N5205);
not NOT1 (N5700, N5696);
and AND3 (N5701, N5689, N3197, N4465);
nor NOR4 (N5702, N5673, N200, N681, N5514);
nand NAND2 (N5703, N5698, N2112);
nand NAND4 (N5704, N5685, N2311, N2437, N206);
xor XOR2 (N5705, N5699, N2911);
or OR2 (N5706, N5694, N5466);
and AND4 (N5707, N5700, N5277, N625, N636);
xor XOR2 (N5708, N5707, N4072);
nor NOR4 (N5709, N5701, N1885, N4036, N1621);
not NOT1 (N5710, N5708);
or OR3 (N5711, N5704, N4706, N488);
and AND3 (N5712, N5710, N2548, N4864);
buf BUF1 (N5713, N5709);
not NOT1 (N5714, N5702);
or OR4 (N5715, N5690, N879, N1998, N2626);
nor NOR2 (N5716, N5713, N3552);
xor XOR2 (N5717, N5716, N2219);
or OR2 (N5718, N5712, N5087);
buf BUF1 (N5719, N5714);
and AND4 (N5720, N5715, N344, N4493, N1388);
xor XOR2 (N5721, N5705, N4639);
or OR4 (N5722, N5719, N4746, N3073, N1073);
or OR2 (N5723, N5688, N2029);
xor XOR2 (N5724, N5691, N5595);
nor NOR2 (N5725, N5722, N1651);
xor XOR2 (N5726, N5718, N5588);
not NOT1 (N5727, N5721);
nor NOR4 (N5728, N5720, N3716, N3756, N1647);
and AND2 (N5729, N5711, N2780);
buf BUF1 (N5730, N5717);
xor XOR2 (N5731, N5703, N785);
not NOT1 (N5732, N5729);
and AND4 (N5733, N5723, N4191, N2792, N1868);
nand NAND3 (N5734, N5706, N5671, N5463);
not NOT1 (N5735, N5732);
nor NOR4 (N5736, N5725, N2827, N1147, N717);
and AND4 (N5737, N5730, N4593, N1485, N2116);
and AND2 (N5738, N5728, N930);
or OR3 (N5739, N5737, N238, N4971);
or OR4 (N5740, N5739, N3814, N2697, N5163);
nor NOR3 (N5741, N5740, N3996, N3822);
or OR3 (N5742, N5736, N1041, N5584);
and AND2 (N5743, N5727, N402);
and AND3 (N5744, N5726, N5511, N494);
and AND2 (N5745, N5743, N2241);
nor NOR4 (N5746, N5724, N1677, N1657, N5362);
and AND2 (N5747, N5733, N2756);
or OR3 (N5748, N5741, N2697, N1277);
buf BUF1 (N5749, N5742);
or OR2 (N5750, N5731, N4092);
and AND2 (N5751, N5738, N1802);
buf BUF1 (N5752, N5734);
or OR2 (N5753, N5751, N234);
nand NAND2 (N5754, N5735, N5699);
buf BUF1 (N5755, N5747);
not NOT1 (N5756, N5753);
and AND4 (N5757, N5744, N4253, N3475, N3196);
not NOT1 (N5758, N5748);
nand NAND3 (N5759, N5758, N559, N1420);
buf BUF1 (N5760, N5749);
and AND4 (N5761, N5752, N4518, N1060, N1140);
nand NAND2 (N5762, N5745, N295);
and AND2 (N5763, N5757, N5705);
xor XOR2 (N5764, N5763, N2571);
or OR3 (N5765, N5754, N772, N197);
xor XOR2 (N5766, N5756, N4699);
nor NOR2 (N5767, N5761, N130);
nor NOR4 (N5768, N5760, N4147, N4978, N1269);
buf BUF1 (N5769, N5755);
or OR3 (N5770, N5766, N5417, N5216);
nand NAND4 (N5771, N5750, N5314, N628, N3136);
nor NOR2 (N5772, N5768, N4098);
nand NAND4 (N5773, N5765, N1603, N788, N1043);
not NOT1 (N5774, N5764);
nor NOR2 (N5775, N5770, N4832);
and AND3 (N5776, N5775, N5353, N5388);
not NOT1 (N5777, N5772);
and AND4 (N5778, N5767, N4305, N5732, N3590);
not NOT1 (N5779, N5759);
not NOT1 (N5780, N5774);
or OR4 (N5781, N5769, N1174, N4667, N356);
xor XOR2 (N5782, N5780, N2924);
and AND2 (N5783, N5782, N2841);
not NOT1 (N5784, N5779);
not NOT1 (N5785, N5746);
nor NOR2 (N5786, N5783, N4863);
buf BUF1 (N5787, N5762);
nor NOR3 (N5788, N5786, N576, N3477);
and AND3 (N5789, N5773, N752, N5751);
or OR3 (N5790, N5785, N3547, N4276);
buf BUF1 (N5791, N5789);
nor NOR3 (N5792, N5784, N1177, N2594);
not NOT1 (N5793, N5778);
xor XOR2 (N5794, N5788, N4581);
nand NAND2 (N5795, N5776, N5089);
nand NAND2 (N5796, N5794, N3781);
and AND4 (N5797, N5792, N1366, N56, N3444);
nand NAND3 (N5798, N5777, N5304, N1542);
and AND3 (N5799, N5771, N409, N4695);
nor NOR3 (N5800, N5787, N1376, N3444);
xor XOR2 (N5801, N5791, N723);
nand NAND4 (N5802, N5799, N4118, N587, N856);
nand NAND2 (N5803, N5802, N3177);
or OR3 (N5804, N5801, N2157, N3746);
not NOT1 (N5805, N5800);
nand NAND3 (N5806, N5797, N4726, N5670);
xor XOR2 (N5807, N5793, N3611);
not NOT1 (N5808, N5796);
nand NAND2 (N5809, N5807, N1998);
not NOT1 (N5810, N5805);
xor XOR2 (N5811, N5781, N5488);
xor XOR2 (N5812, N5809, N4421);
or OR4 (N5813, N5808, N665, N2344, N855);
nor NOR3 (N5814, N5804, N4720, N861);
nor NOR4 (N5815, N5790, N4680, N705, N5058);
xor XOR2 (N5816, N5811, N1096);
buf BUF1 (N5817, N5803);
buf BUF1 (N5818, N5814);
not NOT1 (N5819, N5812);
not NOT1 (N5820, N5819);
xor XOR2 (N5821, N5818, N5309);
not NOT1 (N5822, N5795);
and AND3 (N5823, N5813, N26, N656);
nor NOR3 (N5824, N5798, N2664, N190);
and AND2 (N5825, N5817, N1677);
nor NOR2 (N5826, N5824, N5033);
or OR3 (N5827, N5825, N5189, N4355);
and AND4 (N5828, N5810, N610, N2088, N2445);
buf BUF1 (N5829, N5828);
or OR3 (N5830, N5829, N1768, N2992);
and AND4 (N5831, N5816, N3961, N298, N1324);
nor NOR2 (N5832, N5820, N2411);
buf BUF1 (N5833, N5826);
nand NAND2 (N5834, N5823, N1975);
or OR2 (N5835, N5833, N277);
and AND4 (N5836, N5822, N5542, N804, N4214);
xor XOR2 (N5837, N5834, N4145);
not NOT1 (N5838, N5831);
buf BUF1 (N5839, N5815);
nand NAND4 (N5840, N5827, N3268, N4517, N3456);
and AND4 (N5841, N5838, N5749, N4233, N334);
xor XOR2 (N5842, N5806, N908);
xor XOR2 (N5843, N5841, N3954);
and AND2 (N5844, N5830, N1851);
buf BUF1 (N5845, N5840);
not NOT1 (N5846, N5837);
buf BUF1 (N5847, N5821);
and AND3 (N5848, N5839, N4025, N5669);
or OR4 (N5849, N5846, N448, N1765, N4457);
or OR2 (N5850, N5832, N4322);
and AND3 (N5851, N5847, N2893, N1363);
and AND3 (N5852, N5844, N4013, N5803);
xor XOR2 (N5853, N5849, N4696);
not NOT1 (N5854, N5852);
or OR3 (N5855, N5850, N4299, N4649);
buf BUF1 (N5856, N5842);
xor XOR2 (N5857, N5851, N1435);
nand NAND3 (N5858, N5848, N470, N3560);
not NOT1 (N5859, N5845);
nand NAND2 (N5860, N5857, N4281);
xor XOR2 (N5861, N5835, N239);
xor XOR2 (N5862, N5860, N4664);
buf BUF1 (N5863, N5861);
and AND2 (N5864, N5853, N3278);
or OR3 (N5865, N5859, N4051, N92);
not NOT1 (N5866, N5865);
nor NOR2 (N5867, N5843, N1213);
xor XOR2 (N5868, N5867, N5862);
nand NAND2 (N5869, N5831, N2672);
nor NOR3 (N5870, N5868, N2895, N4497);
not NOT1 (N5871, N5870);
buf BUF1 (N5872, N5836);
nand NAND4 (N5873, N5855, N4066, N684, N4538);
or OR3 (N5874, N5872, N4786, N2368);
nor NOR3 (N5875, N5866, N38, N5391);
xor XOR2 (N5876, N5863, N2577);
nor NOR4 (N5877, N5871, N2806, N4045, N179);
nand NAND4 (N5878, N5876, N3190, N313, N5624);
or OR4 (N5879, N5854, N1360, N3884, N5577);
or OR3 (N5880, N5875, N1677, N1939);
buf BUF1 (N5881, N5878);
nor NOR2 (N5882, N5873, N256);
xor XOR2 (N5883, N5880, N4846);
or OR4 (N5884, N5877, N604, N2316, N431);
nor NOR2 (N5885, N5883, N5050);
buf BUF1 (N5886, N5869);
or OR4 (N5887, N5881, N106, N184, N5151);
xor XOR2 (N5888, N5874, N4045);
or OR4 (N5889, N5882, N4630, N5321, N1150);
nor NOR2 (N5890, N5858, N4911);
nor NOR2 (N5891, N5879, N18);
not NOT1 (N5892, N5884);
buf BUF1 (N5893, N5889);
and AND3 (N5894, N5887, N82, N822);
nand NAND2 (N5895, N5864, N4019);
nor NOR3 (N5896, N5856, N4988, N1843);
or OR3 (N5897, N5896, N5082, N5345);
buf BUF1 (N5898, N5894);
and AND4 (N5899, N5885, N420, N3605, N3282);
not NOT1 (N5900, N5897);
nor NOR3 (N5901, N5891, N2044, N2638);
nor NOR4 (N5902, N5900, N2387, N151, N4971);
not NOT1 (N5903, N5890);
xor XOR2 (N5904, N5888, N2886);
and AND4 (N5905, N5899, N564, N5142, N3436);
buf BUF1 (N5906, N5905);
buf BUF1 (N5907, N5892);
and AND4 (N5908, N5898, N2859, N1931, N4305);
not NOT1 (N5909, N5893);
nand NAND4 (N5910, N5902, N5839, N1552, N3002);
or OR2 (N5911, N5907, N1235);
not NOT1 (N5912, N5895);
nor NOR3 (N5913, N5901, N1110, N4890);
not NOT1 (N5914, N5886);
not NOT1 (N5915, N5906);
not NOT1 (N5916, N5911);
buf BUF1 (N5917, N5908);
nor NOR3 (N5918, N5915, N5318, N4065);
and AND2 (N5919, N5918, N4395);
or OR2 (N5920, N5904, N5150);
nor NOR2 (N5921, N5919, N693);
or OR2 (N5922, N5912, N2365);
nor NOR4 (N5923, N5917, N4278, N1185, N822);
and AND3 (N5924, N5909, N2845, N5783);
or OR4 (N5925, N5910, N2921, N3967, N2336);
nor NOR3 (N5926, N5922, N5345, N3931);
and AND4 (N5927, N5920, N2960, N5917, N4126);
or OR4 (N5928, N5921, N990, N2572, N5119);
or OR3 (N5929, N5903, N1406, N3615);
buf BUF1 (N5930, N5916);
nand NAND3 (N5931, N5913, N1888, N2126);
not NOT1 (N5932, N5924);
nand NAND4 (N5933, N5923, N1944, N5228, N183);
not NOT1 (N5934, N5932);
and AND4 (N5935, N5925, N2405, N5373, N1261);
nor NOR2 (N5936, N5926, N951);
or OR4 (N5937, N5928, N5237, N1582, N4593);
and AND3 (N5938, N5931, N2367, N350);
nand NAND3 (N5939, N5929, N886, N210);
nand NAND3 (N5940, N5938, N5712, N2053);
xor XOR2 (N5941, N5914, N5284);
buf BUF1 (N5942, N5941);
not NOT1 (N5943, N5934);
nor NOR4 (N5944, N5939, N4099, N2090, N5834);
nor NOR3 (N5945, N5933, N4195, N2737);
nor NOR2 (N5946, N5945, N125);
nand NAND2 (N5947, N5943, N3436);
and AND3 (N5948, N5947, N5552, N2088);
xor XOR2 (N5949, N5940, N5790);
not NOT1 (N5950, N5948);
not NOT1 (N5951, N5949);
xor XOR2 (N5952, N5950, N5171);
not NOT1 (N5953, N5946);
not NOT1 (N5954, N5936);
and AND2 (N5955, N5942, N4860);
nand NAND3 (N5956, N5935, N121, N2776);
not NOT1 (N5957, N5944);
buf BUF1 (N5958, N5927);
xor XOR2 (N5959, N5954, N5763);
xor XOR2 (N5960, N5953, N380);
nand NAND2 (N5961, N5937, N182);
and AND4 (N5962, N5952, N5311, N3921, N3572);
and AND4 (N5963, N5956, N1689, N5809, N4663);
or OR4 (N5964, N5930, N1291, N1073, N1340);
nor NOR3 (N5965, N5958, N2102, N4074);
buf BUF1 (N5966, N5963);
not NOT1 (N5967, N5957);
nor NOR3 (N5968, N5951, N5486, N4051);
nor NOR4 (N5969, N5965, N4792, N146, N3455);
nand NAND3 (N5970, N5960, N4895, N4122);
not NOT1 (N5971, N5955);
xor XOR2 (N5972, N5969, N794);
or OR2 (N5973, N5970, N1743);
or OR3 (N5974, N5966, N2301, N4037);
xor XOR2 (N5975, N5974, N5193);
or OR4 (N5976, N5975, N3815, N3208, N5498);
not NOT1 (N5977, N5968);
nand NAND4 (N5978, N5972, N5600, N3742, N1297);
not NOT1 (N5979, N5978);
and AND2 (N5980, N5979, N2531);
nand NAND3 (N5981, N5977, N3652, N597);
and AND4 (N5982, N5971, N1085, N4872, N5890);
buf BUF1 (N5983, N5962);
or OR4 (N5984, N5976, N5498, N4713, N3644);
buf BUF1 (N5985, N5983);
buf BUF1 (N5986, N5967);
and AND2 (N5987, N5973, N1928);
nor NOR3 (N5988, N5986, N119, N3408);
xor XOR2 (N5989, N5987, N4616);
buf BUF1 (N5990, N5982);
xor XOR2 (N5991, N5985, N5407);
and AND3 (N5992, N5988, N923, N4294);
and AND4 (N5993, N5984, N3707, N2682, N1287);
buf BUF1 (N5994, N5959);
nand NAND2 (N5995, N5980, N2258);
not NOT1 (N5996, N5991);
buf BUF1 (N5997, N5993);
xor XOR2 (N5998, N5989, N2768);
or OR3 (N5999, N5964, N5475, N1398);
xor XOR2 (N6000, N5997, N1361);
or OR3 (N6001, N5994, N4591, N367);
or OR2 (N6002, N6001, N4169);
nand NAND4 (N6003, N5981, N2048, N291, N5390);
nor NOR2 (N6004, N6002, N699);
nand NAND4 (N6005, N6004, N691, N5769, N580);
nor NOR2 (N6006, N5998, N3747);
or OR2 (N6007, N5995, N5562);
xor XOR2 (N6008, N6000, N1618);
or OR2 (N6009, N6007, N1723);
buf BUF1 (N6010, N5996);
and AND4 (N6011, N5992, N640, N4521, N803);
not NOT1 (N6012, N6006);
buf BUF1 (N6013, N6011);
buf BUF1 (N6014, N6005);
and AND3 (N6015, N6009, N2025, N5128);
not NOT1 (N6016, N5999);
or OR4 (N6017, N5961, N6009, N2282, N670);
nand NAND2 (N6018, N6008, N2825);
nor NOR4 (N6019, N6015, N3893, N3942, N2526);
nor NOR4 (N6020, N6016, N119, N4390, N4452);
not NOT1 (N6021, N5990);
nand NAND4 (N6022, N6019, N2055, N1666, N3714);
buf BUF1 (N6023, N6020);
or OR2 (N6024, N6022, N2721);
and AND3 (N6025, N6018, N3459, N416);
nand NAND4 (N6026, N6013, N2041, N3985, N3166);
or OR3 (N6027, N6023, N5216, N2667);
nor NOR2 (N6028, N6012, N5262);
not NOT1 (N6029, N6026);
buf BUF1 (N6030, N6014);
and AND2 (N6031, N6017, N4344);
xor XOR2 (N6032, N6025, N5592);
xor XOR2 (N6033, N6030, N1670);
nor NOR3 (N6034, N6027, N1696, N4);
not NOT1 (N6035, N6010);
and AND2 (N6036, N6031, N4497);
nand NAND4 (N6037, N6028, N3565, N885, N148);
not NOT1 (N6038, N6037);
buf BUF1 (N6039, N6038);
not NOT1 (N6040, N6024);
nand NAND2 (N6041, N6035, N4711);
buf BUF1 (N6042, N6036);
nor NOR2 (N6043, N6021, N5290);
xor XOR2 (N6044, N6033, N1194);
nand NAND3 (N6045, N6003, N1528, N12);
buf BUF1 (N6046, N6042);
or OR4 (N6047, N6032, N5983, N1004, N3167);
nor NOR3 (N6048, N6043, N3571, N5520);
nor NOR2 (N6049, N6040, N3520);
and AND3 (N6050, N6034, N2925, N4261);
nand NAND3 (N6051, N6049, N3335, N4929);
buf BUF1 (N6052, N6048);
buf BUF1 (N6053, N6044);
xor XOR2 (N6054, N6051, N3651);
or OR4 (N6055, N6052, N2017, N1147, N1122);
not NOT1 (N6056, N6047);
nor NOR4 (N6057, N6029, N227, N5065, N5097);
buf BUF1 (N6058, N6039);
or OR3 (N6059, N6045, N3523, N5910);
xor XOR2 (N6060, N6054, N3956);
nor NOR4 (N6061, N6055, N5167, N2845, N51);
or OR4 (N6062, N6057, N682, N3681, N3501);
nor NOR4 (N6063, N6053, N1041, N5161, N4666);
buf BUF1 (N6064, N6060);
xor XOR2 (N6065, N6063, N4975);
nor NOR3 (N6066, N6059, N1765, N2201);
or OR3 (N6067, N6041, N4676, N5514);
or OR4 (N6068, N6062, N2962, N816, N106);
and AND3 (N6069, N6058, N2692, N639);
nand NAND3 (N6070, N6069, N4016, N5600);
and AND2 (N6071, N6065, N2245);
and AND3 (N6072, N6050, N5533, N4850);
and AND2 (N6073, N6046, N5406);
and AND2 (N6074, N6067, N4768);
xor XOR2 (N6075, N6071, N515);
buf BUF1 (N6076, N6068);
nand NAND2 (N6077, N6070, N6058);
nor NOR3 (N6078, N6073, N1045, N5403);
not NOT1 (N6079, N6072);
nor NOR2 (N6080, N6061, N1646);
buf BUF1 (N6081, N6078);
or OR4 (N6082, N6066, N3232, N5163, N5290);
not NOT1 (N6083, N6079);
nand NAND4 (N6084, N6082, N5562, N5769, N1901);
not NOT1 (N6085, N6081);
not NOT1 (N6086, N6056);
buf BUF1 (N6087, N6086);
xor XOR2 (N6088, N6084, N5116);
xor XOR2 (N6089, N6080, N1232);
not NOT1 (N6090, N6085);
or OR2 (N6091, N6088, N1044);
xor XOR2 (N6092, N6076, N5125);
nor NOR3 (N6093, N6077, N4633, N5268);
buf BUF1 (N6094, N6090);
or OR3 (N6095, N6087, N1242, N1097);
and AND2 (N6096, N6092, N5670);
and AND2 (N6097, N6091, N5575);
buf BUF1 (N6098, N6095);
or OR3 (N6099, N6094, N3357, N655);
and AND3 (N6100, N6093, N54, N4203);
xor XOR2 (N6101, N6083, N1741);
nand NAND2 (N6102, N6099, N5436);
xor XOR2 (N6103, N6102, N486);
or OR2 (N6104, N6098, N247);
nor NOR4 (N6105, N6074, N3356, N92, N3552);
not NOT1 (N6106, N6075);
nor NOR4 (N6107, N6064, N1651, N1168, N1997);
nand NAND3 (N6108, N6097, N2278, N4779);
or OR2 (N6109, N6106, N3695);
xor XOR2 (N6110, N6109, N3421);
xor XOR2 (N6111, N6107, N3284);
or OR2 (N6112, N6110, N2312);
nor NOR4 (N6113, N6100, N2291, N118, N1136);
and AND3 (N6114, N6101, N2, N2986);
nor NOR3 (N6115, N6108, N4569, N2405);
nand NAND3 (N6116, N6113, N233, N2103);
and AND3 (N6117, N6114, N1671, N556);
not NOT1 (N6118, N6115);
buf BUF1 (N6119, N6111);
and AND3 (N6120, N6104, N1391, N2215);
or OR4 (N6121, N6117, N554, N2000, N578);
and AND3 (N6122, N6096, N1526, N5891);
nand NAND4 (N6123, N6116, N366, N3929, N4320);
nor NOR4 (N6124, N6121, N4991, N5705, N766);
nor NOR2 (N6125, N6103, N573);
nor NOR4 (N6126, N6125, N2189, N84, N1348);
buf BUF1 (N6127, N6118);
nand NAND4 (N6128, N6127, N2467, N2000, N249);
not NOT1 (N6129, N6089);
and AND4 (N6130, N6120, N4941, N1833, N957);
xor XOR2 (N6131, N6126, N550);
nand NAND2 (N6132, N6131, N5446);
nand NAND2 (N6133, N6132, N4830);
or OR2 (N6134, N6124, N5340);
and AND3 (N6135, N6129, N837, N1696);
nand NAND3 (N6136, N6134, N6047, N5181);
and AND2 (N6137, N6128, N3724);
and AND2 (N6138, N6105, N4257);
nor NOR4 (N6139, N6135, N2176, N3441, N5354);
buf BUF1 (N6140, N6137);
nor NOR3 (N6141, N6133, N1362, N103);
or OR3 (N6142, N6130, N495, N1224);
or OR2 (N6143, N6112, N3925);
nand NAND2 (N6144, N6136, N5276);
and AND3 (N6145, N6144, N2330, N2048);
or OR2 (N6146, N6138, N2317);
nand NAND2 (N6147, N6122, N2850);
nand NAND2 (N6148, N6139, N6112);
and AND3 (N6149, N6142, N317, N2744);
buf BUF1 (N6150, N6141);
or OR2 (N6151, N6147, N3892);
nand NAND2 (N6152, N6123, N3145);
nand NAND3 (N6153, N6143, N4208, N1310);
nor NOR4 (N6154, N6145, N2074, N3466, N1209);
nor NOR2 (N6155, N6148, N2666);
buf BUF1 (N6156, N6151);
nand NAND4 (N6157, N6150, N4354, N1763, N2941);
or OR3 (N6158, N6140, N5417, N4884);
and AND2 (N6159, N6155, N1101);
nand NAND2 (N6160, N6153, N396);
not NOT1 (N6161, N6119);
nor NOR2 (N6162, N6157, N314);
buf BUF1 (N6163, N6152);
not NOT1 (N6164, N6161);
and AND2 (N6165, N6154, N1852);
and AND2 (N6166, N6146, N951);
nor NOR4 (N6167, N6166, N5122, N2937, N3624);
nor NOR2 (N6168, N6163, N1379);
and AND4 (N6169, N6156, N2825, N1868, N4935);
or OR3 (N6170, N6162, N2494, N3299);
and AND3 (N6171, N6149, N964, N4541);
nor NOR4 (N6172, N6158, N931, N2089, N1974);
xor XOR2 (N6173, N6159, N536);
buf BUF1 (N6174, N6172);
nor NOR3 (N6175, N6165, N4835, N3957);
or OR2 (N6176, N6175, N4046);
or OR2 (N6177, N6164, N1590);
not NOT1 (N6178, N6176);
or OR3 (N6179, N6174, N2891, N6123);
nor NOR3 (N6180, N6169, N2093, N4843);
or OR4 (N6181, N6180, N394, N3977, N2725);
nand NAND3 (N6182, N6167, N6180, N4180);
and AND4 (N6183, N6178, N599, N4281, N513);
nand NAND2 (N6184, N6168, N3854);
or OR4 (N6185, N6182, N2622, N1688, N3360);
not NOT1 (N6186, N6170);
not NOT1 (N6187, N6179);
buf BUF1 (N6188, N6185);
and AND2 (N6189, N6183, N4006);
not NOT1 (N6190, N6188);
or OR2 (N6191, N6173, N4280);
and AND2 (N6192, N6190, N3874);
nor NOR4 (N6193, N6160, N2522, N2757, N2721);
or OR4 (N6194, N6186, N3303, N916, N5751);
not NOT1 (N6195, N6189);
not NOT1 (N6196, N6184);
buf BUF1 (N6197, N6195);
nand NAND4 (N6198, N6192, N2206, N653, N1627);
nand NAND3 (N6199, N6198, N1041, N3300);
and AND2 (N6200, N6199, N939);
buf BUF1 (N6201, N6187);
and AND2 (N6202, N6194, N1012);
nand NAND4 (N6203, N6177, N723, N4286, N524);
buf BUF1 (N6204, N6201);
buf BUF1 (N6205, N6204);
nand NAND2 (N6206, N6191, N509);
nor NOR3 (N6207, N6171, N4455, N2911);
not NOT1 (N6208, N6202);
buf BUF1 (N6209, N6203);
nand NAND3 (N6210, N6197, N3674, N2740);
nor NOR2 (N6211, N6207, N2956);
nor NOR3 (N6212, N6181, N3387, N529);
buf BUF1 (N6213, N6196);
nand NAND2 (N6214, N6206, N4402);
nor NOR4 (N6215, N6211, N3732, N294, N2276);
not NOT1 (N6216, N6214);
nand NAND2 (N6217, N6216, N3424);
buf BUF1 (N6218, N6212);
xor XOR2 (N6219, N6217, N3019);
xor XOR2 (N6220, N6208, N5452);
and AND2 (N6221, N6193, N4848);
xor XOR2 (N6222, N6215, N3549);
nor NOR3 (N6223, N6213, N2241, N4784);
xor XOR2 (N6224, N6200, N5660);
xor XOR2 (N6225, N6205, N3535);
and AND4 (N6226, N6224, N493, N584, N713);
not NOT1 (N6227, N6221);
nor NOR3 (N6228, N6209, N3089, N5967);
xor XOR2 (N6229, N6226, N5724);
xor XOR2 (N6230, N6222, N458);
buf BUF1 (N6231, N6210);
and AND4 (N6232, N6223, N4732, N1960, N3422);
or OR2 (N6233, N6231, N2491);
nor NOR3 (N6234, N6229, N3206, N3776);
or OR4 (N6235, N6233, N5482, N1691, N4045);
nand NAND3 (N6236, N6225, N1551, N4642);
nand NAND3 (N6237, N6235, N5672, N4716);
or OR2 (N6238, N6232, N1523);
buf BUF1 (N6239, N6230);
and AND3 (N6240, N6218, N4651, N5376);
not NOT1 (N6241, N6234);
xor XOR2 (N6242, N6236, N4390);
buf BUF1 (N6243, N6219);
and AND4 (N6244, N6238, N6046, N2610, N4957);
nand NAND4 (N6245, N6244, N5464, N6107, N1884);
or OR3 (N6246, N6241, N4390, N3229);
buf BUF1 (N6247, N6237);
buf BUF1 (N6248, N6246);
nor NOR3 (N6249, N6243, N4907, N1700);
nor NOR4 (N6250, N6248, N5688, N4870, N909);
not NOT1 (N6251, N6227);
not NOT1 (N6252, N6239);
xor XOR2 (N6253, N6251, N98);
nand NAND3 (N6254, N6228, N1537, N5660);
not NOT1 (N6255, N6245);
not NOT1 (N6256, N6254);
or OR4 (N6257, N6252, N2244, N5398, N3851);
nand NAND4 (N6258, N6242, N5558, N1656, N2649);
buf BUF1 (N6259, N6249);
not NOT1 (N6260, N6259);
not NOT1 (N6261, N6258);
nor NOR2 (N6262, N6240, N5241);
or OR2 (N6263, N6261, N1595);
nand NAND4 (N6264, N6262, N90, N5774, N4293);
nand NAND3 (N6265, N6256, N665, N813);
not NOT1 (N6266, N6247);
or OR4 (N6267, N6264, N5441, N5907, N1138);
not NOT1 (N6268, N6266);
not NOT1 (N6269, N6268);
buf BUF1 (N6270, N6267);
xor XOR2 (N6271, N6255, N2731);
nand NAND3 (N6272, N6265, N529, N3254);
and AND2 (N6273, N6257, N4484);
buf BUF1 (N6274, N6250);
nor NOR4 (N6275, N6263, N3287, N6149, N512);
or OR3 (N6276, N6275, N2443, N1677);
nor NOR4 (N6277, N6276, N2859, N845, N1600);
not NOT1 (N6278, N6277);
buf BUF1 (N6279, N6220);
nor NOR3 (N6280, N6271, N3119, N1785);
nand NAND3 (N6281, N6272, N2172, N5617);
and AND4 (N6282, N6274, N6175, N4731, N5409);
xor XOR2 (N6283, N6269, N2948);
and AND4 (N6284, N6273, N6264, N1606, N5613);
buf BUF1 (N6285, N6260);
not NOT1 (N6286, N6284);
and AND2 (N6287, N6283, N2425);
buf BUF1 (N6288, N6279);
xor XOR2 (N6289, N6278, N5288);
nor NOR4 (N6290, N6281, N432, N3606, N925);
or OR4 (N6291, N6288, N2757, N4925, N2841);
and AND3 (N6292, N6270, N3540, N5715);
nand NAND3 (N6293, N6285, N4616, N3725);
and AND4 (N6294, N6286, N6151, N767, N3855);
or OR3 (N6295, N6253, N3106, N3645);
or OR3 (N6296, N6290, N1636, N4564);
nor NOR3 (N6297, N6287, N1926, N3304);
not NOT1 (N6298, N6282);
and AND3 (N6299, N6289, N3814, N447);
not NOT1 (N6300, N6295);
or OR2 (N6301, N6298, N4008);
and AND4 (N6302, N6299, N4107, N2347, N5885);
buf BUF1 (N6303, N6291);
and AND2 (N6304, N6280, N3953);
buf BUF1 (N6305, N6292);
nor NOR4 (N6306, N6305, N4836, N5355, N1836);
or OR2 (N6307, N6304, N4889);
nor NOR4 (N6308, N6300, N2621, N2733, N5874);
not NOT1 (N6309, N6308);
nand NAND3 (N6310, N6306, N5477, N4541);
or OR2 (N6311, N6310, N1806);
xor XOR2 (N6312, N6294, N4979);
and AND2 (N6313, N6296, N801);
buf BUF1 (N6314, N6311);
xor XOR2 (N6315, N6297, N2355);
nor NOR2 (N6316, N6302, N550);
not NOT1 (N6317, N6314);
not NOT1 (N6318, N6309);
buf BUF1 (N6319, N6307);
buf BUF1 (N6320, N6293);
nor NOR2 (N6321, N6313, N5585);
nand NAND2 (N6322, N6318, N2463);
not NOT1 (N6323, N6301);
xor XOR2 (N6324, N6303, N1005);
nand NAND3 (N6325, N6320, N2003, N4864);
or OR2 (N6326, N6312, N6156);
or OR2 (N6327, N6319, N618);
and AND3 (N6328, N6317, N1932, N813);
nand NAND2 (N6329, N6322, N5891);
not NOT1 (N6330, N6315);
not NOT1 (N6331, N6323);
not NOT1 (N6332, N6316);
nor NOR4 (N6333, N6328, N3734, N4449, N2004);
not NOT1 (N6334, N6331);
not NOT1 (N6335, N6324);
nand NAND2 (N6336, N6330, N2159);
xor XOR2 (N6337, N6336, N3684);
not NOT1 (N6338, N6327);
not NOT1 (N6339, N6326);
and AND2 (N6340, N6332, N6163);
not NOT1 (N6341, N6338);
and AND3 (N6342, N6333, N2571, N168);
nand NAND2 (N6343, N6339, N1950);
buf BUF1 (N6344, N6329);
buf BUF1 (N6345, N6340);
xor XOR2 (N6346, N6321, N199);
xor XOR2 (N6347, N6345, N3270);
buf BUF1 (N6348, N6343);
nand NAND2 (N6349, N6341, N3503);
nand NAND4 (N6350, N6342, N4811, N2940, N4905);
nor NOR4 (N6351, N6349, N1619, N400, N2066);
not NOT1 (N6352, N6346);
nand NAND2 (N6353, N6351, N5946);
not NOT1 (N6354, N6344);
not NOT1 (N6355, N6334);
not NOT1 (N6356, N6325);
and AND4 (N6357, N6356, N632, N656, N568);
or OR2 (N6358, N6347, N1578);
nor NOR4 (N6359, N6350, N3697, N2248, N4070);
nand NAND2 (N6360, N6337, N5570);
and AND4 (N6361, N6357, N4037, N4918, N5854);
nand NAND3 (N6362, N6355, N5, N4552);
or OR4 (N6363, N6353, N2981, N1952, N2601);
not NOT1 (N6364, N6363);
nand NAND4 (N6365, N6348, N5446, N4805, N563);
buf BUF1 (N6366, N6360);
xor XOR2 (N6367, N6361, N6156);
not NOT1 (N6368, N6358);
nand NAND4 (N6369, N6366, N4801, N4652, N659);
and AND4 (N6370, N6335, N6024, N6200, N4168);
nor NOR3 (N6371, N6368, N3050, N4389);
not NOT1 (N6372, N6370);
xor XOR2 (N6373, N6365, N2996);
or OR3 (N6374, N6372, N1136, N5276);
nor NOR3 (N6375, N6374, N5296, N5964);
nor NOR2 (N6376, N6359, N120);
or OR4 (N6377, N6371, N5815, N2765, N762);
nor NOR3 (N6378, N6377, N635, N4701);
nand NAND4 (N6379, N6364, N3319, N4269, N1494);
and AND4 (N6380, N6354, N781, N3553, N36);
nand NAND3 (N6381, N6380, N4262, N4445);
buf BUF1 (N6382, N6352);
buf BUF1 (N6383, N6362);
nand NAND3 (N6384, N6376, N3086, N1318);
nor NOR3 (N6385, N6369, N6296, N5600);
nand NAND4 (N6386, N6375, N2365, N3268, N2311);
xor XOR2 (N6387, N6384, N802);
not NOT1 (N6388, N6378);
not NOT1 (N6389, N6382);
or OR3 (N6390, N6389, N2726, N5930);
xor XOR2 (N6391, N6381, N670);
or OR4 (N6392, N6388, N4564, N2783, N609);
and AND2 (N6393, N6379, N6253);
nor NOR3 (N6394, N6385, N328, N4768);
nand NAND2 (N6395, N6391, N2267);
buf BUF1 (N6396, N6393);
nor NOR3 (N6397, N6373, N3858, N2347);
not NOT1 (N6398, N6390);
and AND2 (N6399, N6397, N1530);
nand NAND4 (N6400, N6383, N1047, N5942, N5821);
nand NAND2 (N6401, N6400, N2824);
buf BUF1 (N6402, N6398);
nand NAND2 (N6403, N6387, N4971);
nand NAND3 (N6404, N6401, N6159, N3558);
nand NAND2 (N6405, N6392, N423);
buf BUF1 (N6406, N6402);
not NOT1 (N6407, N6405);
or OR2 (N6408, N6399, N742);
nand NAND3 (N6409, N6396, N6194, N5791);
or OR2 (N6410, N6404, N2778);
not NOT1 (N6411, N6407);
nor NOR2 (N6412, N6410, N2205);
or OR2 (N6413, N6386, N1787);
and AND2 (N6414, N6394, N2201);
nor NOR3 (N6415, N6409, N304, N6203);
not NOT1 (N6416, N6367);
nor NOR3 (N6417, N6406, N3425, N6012);
buf BUF1 (N6418, N6413);
and AND3 (N6419, N6414, N2491, N2332);
nand NAND4 (N6420, N6416, N3425, N5095, N4062);
buf BUF1 (N6421, N6420);
not NOT1 (N6422, N6395);
buf BUF1 (N6423, N6422);
not NOT1 (N6424, N6408);
not NOT1 (N6425, N6418);
buf BUF1 (N6426, N6423);
xor XOR2 (N6427, N6412, N3891);
or OR4 (N6428, N6411, N2263, N3901, N5553);
and AND2 (N6429, N6419, N4474);
nand NAND3 (N6430, N6417, N1922, N6334);
nand NAND3 (N6431, N6415, N294, N2450);
or OR3 (N6432, N6421, N1548, N4530);
buf BUF1 (N6433, N6432);
not NOT1 (N6434, N6429);
or OR4 (N6435, N6433, N1133, N1222, N6370);
nor NOR2 (N6436, N6424, N6204);
xor XOR2 (N6437, N6426, N5527);
and AND4 (N6438, N6430, N1540, N1404, N6166);
nor NOR2 (N6439, N6403, N2151);
not NOT1 (N6440, N6439);
and AND3 (N6441, N6431, N2893, N1027);
nor NOR4 (N6442, N6434, N5350, N1646, N4212);
nor NOR2 (N6443, N6425, N2161);
or OR3 (N6444, N6428, N1865, N1820);
nand NAND4 (N6445, N6436, N4381, N5231, N2888);
or OR2 (N6446, N6438, N978);
not NOT1 (N6447, N6435);
nand NAND4 (N6448, N6443, N4615, N5827, N1310);
buf BUF1 (N6449, N6427);
nand NAND4 (N6450, N6449, N883, N1542, N3228);
not NOT1 (N6451, N6442);
nand NAND2 (N6452, N6451, N3646);
and AND4 (N6453, N6444, N2619, N5077, N3513);
nor NOR4 (N6454, N6437, N3978, N3270, N2280);
nor NOR2 (N6455, N6453, N5837);
xor XOR2 (N6456, N6450, N5673);
buf BUF1 (N6457, N6454);
not NOT1 (N6458, N6457);
or OR4 (N6459, N6448, N2398, N4167, N5488);
nor NOR4 (N6460, N6458, N3794, N2144, N2552);
xor XOR2 (N6461, N6447, N3565);
not NOT1 (N6462, N6452);
nor NOR2 (N6463, N6459, N5000);
or OR2 (N6464, N6455, N4243);
xor XOR2 (N6465, N6441, N5159);
nor NOR3 (N6466, N6440, N1813, N5212);
or OR4 (N6467, N6446, N3137, N251, N3765);
or OR2 (N6468, N6464, N2808);
nand NAND2 (N6469, N6466, N976);
and AND3 (N6470, N6462, N1839, N4607);
and AND2 (N6471, N6467, N5045);
nand NAND3 (N6472, N6469, N1228, N1480);
not NOT1 (N6473, N6461);
or OR2 (N6474, N6445, N2160);
nor NOR4 (N6475, N6474, N1024, N6325, N1425);
xor XOR2 (N6476, N6465, N4310);
buf BUF1 (N6477, N6470);
nand NAND4 (N6478, N6475, N3094, N5976, N705);
or OR3 (N6479, N6456, N2933, N414);
xor XOR2 (N6480, N6463, N5857);
nor NOR4 (N6481, N6473, N4406, N5941, N4889);
or OR2 (N6482, N6472, N1586);
and AND4 (N6483, N6468, N5588, N943, N2846);
not NOT1 (N6484, N6478);
xor XOR2 (N6485, N6482, N6339);
nand NAND3 (N6486, N6477, N2002, N3468);
xor XOR2 (N6487, N6479, N2492);
nor NOR4 (N6488, N6471, N1938, N5245, N6139);
or OR3 (N6489, N6480, N1588, N1895);
or OR2 (N6490, N6481, N2605);
xor XOR2 (N6491, N6485, N843);
xor XOR2 (N6492, N6486, N4431);
or OR4 (N6493, N6483, N140, N4291, N1353);
nand NAND3 (N6494, N6490, N5531, N155);
nor NOR4 (N6495, N6460, N1606, N4807, N282);
nand NAND3 (N6496, N6492, N187, N4872);
buf BUF1 (N6497, N6488);
buf BUF1 (N6498, N6495);
buf BUF1 (N6499, N6496);
xor XOR2 (N6500, N6487, N1144);
nand NAND4 (N6501, N6489, N5552, N5734, N5977);
buf BUF1 (N6502, N6493);
buf BUF1 (N6503, N6484);
and AND2 (N6504, N6498, N1881);
and AND2 (N6505, N6494, N5575);
xor XOR2 (N6506, N6491, N730);
nor NOR4 (N6507, N6505, N6394, N1268, N302);
or OR4 (N6508, N6501, N2783, N2475, N3619);
nor NOR4 (N6509, N6503, N183, N424, N1259);
buf BUF1 (N6510, N6509);
not NOT1 (N6511, N6497);
nor NOR4 (N6512, N6507, N3212, N2447, N2032);
nand NAND3 (N6513, N6506, N2509, N4031);
nor NOR2 (N6514, N6500, N6143);
nor NOR3 (N6515, N6513, N130, N6431);
nor NOR4 (N6516, N6499, N3180, N4351, N1605);
or OR4 (N6517, N6514, N1852, N983, N6200);
nor NOR4 (N6518, N6511, N2553, N2317, N5931);
buf BUF1 (N6519, N6508);
nor NOR4 (N6520, N6504, N2656, N2472, N4738);
not NOT1 (N6521, N6518);
not NOT1 (N6522, N6502);
xor XOR2 (N6523, N6515, N1600);
not NOT1 (N6524, N6512);
nor NOR4 (N6525, N6510, N5143, N4848, N5012);
and AND2 (N6526, N6516, N4921);
and AND4 (N6527, N6523, N466, N6112, N323);
xor XOR2 (N6528, N6521, N4917);
nand NAND4 (N6529, N6525, N4180, N6434, N1335);
buf BUF1 (N6530, N6526);
nor NOR4 (N6531, N6517, N1502, N3569, N5107);
nand NAND4 (N6532, N6527, N6503, N2404, N4881);
buf BUF1 (N6533, N6524);
and AND2 (N6534, N6528, N911);
xor XOR2 (N6535, N6522, N6500);
and AND3 (N6536, N6534, N3161, N3265);
buf BUF1 (N6537, N6532);
not NOT1 (N6538, N6529);
nor NOR3 (N6539, N6536, N2732, N4282);
buf BUF1 (N6540, N6538);
or OR2 (N6541, N6531, N6348);
nor NOR2 (N6542, N6520, N1322);
or OR2 (N6543, N6539, N3320);
nand NAND2 (N6544, N6541, N3518);
nand NAND2 (N6545, N6542, N1545);
not NOT1 (N6546, N6540);
nand NAND2 (N6547, N6535, N2123);
or OR3 (N6548, N6537, N5877, N4865);
nor NOR2 (N6549, N6543, N3387);
or OR4 (N6550, N6547, N4712, N3636, N390);
not NOT1 (N6551, N6533);
xor XOR2 (N6552, N6551, N3457);
nor NOR2 (N6553, N6530, N2515);
and AND2 (N6554, N6545, N332);
nor NOR3 (N6555, N6519, N2814, N1457);
nor NOR4 (N6556, N6550, N5312, N1873, N4925);
nand NAND2 (N6557, N6553, N2749);
xor XOR2 (N6558, N6549, N3934);
buf BUF1 (N6559, N6552);
nand NAND4 (N6560, N6558, N6114, N1349, N5864);
and AND4 (N6561, N6544, N2095, N4908, N4373);
and AND4 (N6562, N6556, N4108, N1294, N3116);
xor XOR2 (N6563, N6555, N1301);
or OR4 (N6564, N6557, N1246, N4922, N2066);
xor XOR2 (N6565, N6561, N6365);
nor NOR2 (N6566, N6476, N3907);
not NOT1 (N6567, N6548);
or OR2 (N6568, N6563, N4622);
and AND3 (N6569, N6559, N257, N5729);
not NOT1 (N6570, N6560);
not NOT1 (N6571, N6565);
nand NAND3 (N6572, N6567, N5293, N583);
or OR3 (N6573, N6570, N2291, N5468);
not NOT1 (N6574, N6568);
or OR2 (N6575, N6574, N2708);
nand NAND2 (N6576, N6569, N5817);
nand NAND4 (N6577, N6546, N3457, N6123, N4798);
xor XOR2 (N6578, N6573, N4538);
buf BUF1 (N6579, N6562);
buf BUF1 (N6580, N6578);
nand NAND3 (N6581, N6571, N3090, N6472);
nand NAND2 (N6582, N6577, N3654);
buf BUF1 (N6583, N6579);
nor NOR3 (N6584, N6583, N2842, N1770);
or OR4 (N6585, N6581, N1567, N526, N4864);
buf BUF1 (N6586, N6554);
nand NAND2 (N6587, N6584, N3242);
or OR3 (N6588, N6585, N4268, N4625);
not NOT1 (N6589, N6572);
nand NAND4 (N6590, N6586, N5796, N4747, N5026);
nor NOR3 (N6591, N6564, N6013, N6346);
or OR4 (N6592, N6591, N1000, N1081, N112);
nor NOR3 (N6593, N6592, N5449, N2969);
nor NOR4 (N6594, N6576, N6333, N6589, N5554);
xor XOR2 (N6595, N6070, N1483);
xor XOR2 (N6596, N6587, N1931);
nor NOR3 (N6597, N6575, N1742, N3952);
nor NOR2 (N6598, N6596, N2263);
and AND2 (N6599, N6594, N843);
nor NOR3 (N6600, N6599, N3614, N4406);
nor NOR4 (N6601, N6597, N3911, N4809, N1076);
nor NOR2 (N6602, N6600, N6359);
nor NOR2 (N6603, N6598, N3689);
buf BUF1 (N6604, N6601);
xor XOR2 (N6605, N6603, N5703);
not NOT1 (N6606, N6605);
or OR2 (N6607, N6590, N4627);
nand NAND2 (N6608, N6593, N3003);
or OR2 (N6609, N6604, N1972);
nand NAND3 (N6610, N6602, N4537, N5863);
nand NAND4 (N6611, N6610, N3138, N1067, N444);
xor XOR2 (N6612, N6609, N5369);
and AND4 (N6613, N6566, N1067, N650, N3585);
nor NOR3 (N6614, N6613, N5193, N4765);
nor NOR4 (N6615, N6595, N3850, N489, N1);
xor XOR2 (N6616, N6580, N1147);
not NOT1 (N6617, N6582);
or OR3 (N6618, N6616, N6606, N1059);
not NOT1 (N6619, N4443);
buf BUF1 (N6620, N6619);
not NOT1 (N6621, N6612);
buf BUF1 (N6622, N6607);
and AND4 (N6623, N6615, N3874, N1922, N3614);
xor XOR2 (N6624, N6621, N67);
or OR3 (N6625, N6624, N285, N6388);
nor NOR3 (N6626, N6625, N6186, N91);
or OR2 (N6627, N6608, N3042);
xor XOR2 (N6628, N6614, N1223);
not NOT1 (N6629, N6611);
nand NAND2 (N6630, N6618, N5338);
and AND3 (N6631, N6588, N6365, N1944);
xor XOR2 (N6632, N6629, N3337);
not NOT1 (N6633, N6620);
or OR2 (N6634, N6632, N246);
nand NAND4 (N6635, N6628, N2823, N1443, N2961);
not NOT1 (N6636, N6622);
nor NOR2 (N6637, N6626, N894);
nand NAND4 (N6638, N6635, N6302, N2282, N2491);
and AND3 (N6639, N6617, N6266, N4412);
not NOT1 (N6640, N6627);
or OR2 (N6641, N6637, N6229);
and AND2 (N6642, N6623, N5598);
and AND4 (N6643, N6636, N2115, N6616, N2511);
xor XOR2 (N6644, N6640, N3903);
not NOT1 (N6645, N6638);
buf BUF1 (N6646, N6645);
or OR2 (N6647, N6643, N6414);
nor NOR2 (N6648, N6639, N2649);
buf BUF1 (N6649, N6642);
and AND4 (N6650, N6633, N2161, N5061, N5832);
xor XOR2 (N6651, N6647, N2777);
buf BUF1 (N6652, N6650);
xor XOR2 (N6653, N6641, N4519);
xor XOR2 (N6654, N6653, N335);
xor XOR2 (N6655, N6654, N5920);
not NOT1 (N6656, N6655);
buf BUF1 (N6657, N6646);
and AND2 (N6658, N6634, N3300);
not NOT1 (N6659, N6648);
xor XOR2 (N6660, N6652, N2958);
nand NAND4 (N6661, N6658, N4916, N1325, N2558);
xor XOR2 (N6662, N6659, N4837);
nand NAND2 (N6663, N6631, N672);
xor XOR2 (N6664, N6660, N6485);
and AND4 (N6665, N6662, N4258, N5204, N456);
and AND2 (N6666, N6665, N4044);
buf BUF1 (N6667, N6661);
buf BUF1 (N6668, N6657);
nand NAND4 (N6669, N6666, N827, N5257, N5059);
nand NAND3 (N6670, N6656, N6548, N6017);
nor NOR3 (N6671, N6649, N2392, N3154);
and AND3 (N6672, N6671, N988, N2486);
or OR2 (N6673, N6664, N3684);
and AND4 (N6674, N6673, N1028, N634, N1810);
or OR4 (N6675, N6674, N5364, N4285, N5077);
or OR4 (N6676, N6644, N2712, N674, N3924);
or OR2 (N6677, N6630, N1083);
buf BUF1 (N6678, N6663);
or OR4 (N6679, N6669, N4662, N4006, N491);
or OR2 (N6680, N6676, N5912);
nand NAND4 (N6681, N6672, N2829, N5159, N201);
or OR4 (N6682, N6681, N946, N2841, N983);
xor XOR2 (N6683, N6667, N2679);
or OR3 (N6684, N6670, N2575, N2784);
not NOT1 (N6685, N6677);
nand NAND4 (N6686, N6680, N277, N3117, N3061);
and AND3 (N6687, N6686, N2568, N5483);
or OR2 (N6688, N6675, N4493);
or OR3 (N6689, N6687, N255, N1981);
nand NAND3 (N6690, N6668, N4778, N5648);
and AND4 (N6691, N6685, N5253, N6310, N2042);
xor XOR2 (N6692, N6678, N430);
buf BUF1 (N6693, N6683);
or OR3 (N6694, N6690, N6680, N1966);
and AND3 (N6695, N6689, N5952, N4689);
and AND4 (N6696, N6688, N1454, N3048, N5061);
nand NAND2 (N6697, N6692, N4748);
xor XOR2 (N6698, N6679, N1645);
xor XOR2 (N6699, N6682, N6692);
nand NAND4 (N6700, N6696, N4451, N1124, N5840);
nor NOR4 (N6701, N6684, N3447, N636, N6459);
nor NOR4 (N6702, N6693, N692, N1149, N6274);
or OR3 (N6703, N6697, N6401, N2067);
nor NOR3 (N6704, N6694, N114, N289);
nand NAND2 (N6705, N6703, N3138);
nand NAND2 (N6706, N6704, N3343);
not NOT1 (N6707, N6695);
xor XOR2 (N6708, N6701, N5032);
buf BUF1 (N6709, N6705);
buf BUF1 (N6710, N6691);
and AND2 (N6711, N6651, N9);
and AND4 (N6712, N6698, N1498, N6521, N5241);
buf BUF1 (N6713, N6702);
not NOT1 (N6714, N6711);
xor XOR2 (N6715, N6699, N3578);
and AND2 (N6716, N6700, N4953);
nand NAND3 (N6717, N6707, N6360, N3936);
and AND3 (N6718, N6709, N2939, N5172);
nor NOR2 (N6719, N6714, N3166);
buf BUF1 (N6720, N6717);
or OR2 (N6721, N6718, N5866);
not NOT1 (N6722, N6721);
not NOT1 (N6723, N6710);
or OR4 (N6724, N6712, N6259, N5734, N1407);
or OR3 (N6725, N6722, N1867, N2691);
buf BUF1 (N6726, N6719);
xor XOR2 (N6727, N6726, N3199);
nor NOR2 (N6728, N6723, N2124);
and AND3 (N6729, N6708, N4888, N2122);
not NOT1 (N6730, N6715);
buf BUF1 (N6731, N6730);
buf BUF1 (N6732, N6729);
not NOT1 (N6733, N6716);
or OR2 (N6734, N6733, N2224);
or OR2 (N6735, N6727, N5738);
nor NOR3 (N6736, N6734, N6194, N6273);
not NOT1 (N6737, N6731);
and AND4 (N6738, N6732, N4784, N3016, N237);
and AND4 (N6739, N6720, N3704, N4557, N5841);
and AND2 (N6740, N6725, N4997);
buf BUF1 (N6741, N6740);
not NOT1 (N6742, N6724);
and AND2 (N6743, N6739, N3950);
xor XOR2 (N6744, N6728, N2949);
or OR4 (N6745, N6742, N1723, N3938, N1529);
or OR3 (N6746, N6744, N1620, N2555);
or OR3 (N6747, N6713, N2813, N6399);
nand NAND3 (N6748, N6745, N1649, N3853);
not NOT1 (N6749, N6737);
and AND4 (N6750, N6735, N4774, N3635, N4167);
and AND4 (N6751, N6750, N5699, N149, N2947);
nor NOR3 (N6752, N6746, N2895, N4893);
nand NAND2 (N6753, N6752, N3874);
nand NAND2 (N6754, N6751, N4939);
not NOT1 (N6755, N6741);
nor NOR2 (N6756, N6749, N5767);
and AND3 (N6757, N6755, N1833, N5132);
and AND4 (N6758, N6757, N5650, N5589, N6404);
xor XOR2 (N6759, N6756, N4448);
nand NAND3 (N6760, N6738, N2672, N4606);
xor XOR2 (N6761, N6753, N2355);
not NOT1 (N6762, N6747);
xor XOR2 (N6763, N6754, N3113);
and AND2 (N6764, N6706, N5571);
or OR4 (N6765, N6762, N6676, N1358, N3970);
or OR4 (N6766, N6748, N2398, N3647, N6701);
nand NAND3 (N6767, N6766, N632, N2462);
xor XOR2 (N6768, N6765, N2138);
and AND2 (N6769, N6759, N2529);
not NOT1 (N6770, N6769);
buf BUF1 (N6771, N6743);
not NOT1 (N6772, N6758);
or OR2 (N6773, N6760, N1892);
and AND2 (N6774, N6736, N4635);
not NOT1 (N6775, N6772);
xor XOR2 (N6776, N6763, N485);
or OR2 (N6777, N6773, N2744);
not NOT1 (N6778, N6776);
not NOT1 (N6779, N6767);
nor NOR3 (N6780, N6764, N1938, N4490);
or OR2 (N6781, N6779, N4221);
and AND4 (N6782, N6761, N6482, N5165, N5533);
nand NAND4 (N6783, N6782, N2450, N3304, N2767);
nand NAND4 (N6784, N6781, N4027, N425, N1239);
or OR2 (N6785, N6771, N812);
or OR2 (N6786, N6777, N5869);
or OR2 (N6787, N6785, N2657);
nor NOR2 (N6788, N6770, N6521);
or OR3 (N6789, N6788, N2021, N3895);
and AND2 (N6790, N6787, N3556);
and AND3 (N6791, N6780, N2423, N1306);
not NOT1 (N6792, N6783);
and AND3 (N6793, N6790, N1100, N6308);
xor XOR2 (N6794, N6791, N5187);
buf BUF1 (N6795, N6775);
not NOT1 (N6796, N6774);
not NOT1 (N6797, N6795);
nor NOR3 (N6798, N6797, N5832, N5454);
or OR4 (N6799, N6798, N4737, N2338, N1863);
or OR4 (N6800, N6792, N997, N1236, N358);
nor NOR3 (N6801, N6768, N5635, N1693);
or OR4 (N6802, N6796, N5842, N4296, N3567);
nor NOR4 (N6803, N6802, N664, N362, N891);
or OR3 (N6804, N6789, N4630, N2546);
and AND4 (N6805, N6800, N4465, N506, N1581);
not NOT1 (N6806, N6801);
nand NAND3 (N6807, N6799, N5342, N6614);
xor XOR2 (N6808, N6794, N436);
buf BUF1 (N6809, N6784);
not NOT1 (N6810, N6786);
not NOT1 (N6811, N6808);
nor NOR2 (N6812, N6805, N4383);
nand NAND4 (N6813, N6807, N4837, N366, N3725);
nand NAND3 (N6814, N6804, N1611, N4611);
buf BUF1 (N6815, N6811);
and AND4 (N6816, N6814, N3445, N684, N2499);
xor XOR2 (N6817, N6815, N2180);
or OR2 (N6818, N6810, N587);
not NOT1 (N6819, N6817);
and AND2 (N6820, N6819, N4369);
nand NAND2 (N6821, N6816, N1540);
not NOT1 (N6822, N6818);
buf BUF1 (N6823, N6820);
and AND2 (N6824, N6813, N2845);
xor XOR2 (N6825, N6778, N1441);
buf BUF1 (N6826, N6824);
xor XOR2 (N6827, N6821, N5268);
and AND3 (N6828, N6806, N4811, N4828);
buf BUF1 (N6829, N6809);
or OR4 (N6830, N6803, N3056, N6212, N378);
and AND4 (N6831, N6828, N5836, N3166, N2292);
or OR4 (N6832, N6812, N1387, N5165, N6202);
and AND3 (N6833, N6826, N5343, N3577);
xor XOR2 (N6834, N6829, N2023);
and AND3 (N6835, N6834, N2711, N817);
nor NOR2 (N6836, N6827, N2943);
or OR4 (N6837, N6823, N3566, N5949, N4540);
nor NOR2 (N6838, N6793, N6328);
and AND2 (N6839, N6831, N613);
nor NOR4 (N6840, N6836, N3573, N74, N1553);
or OR4 (N6841, N6837, N4580, N4327, N3022);
not NOT1 (N6842, N6839);
and AND4 (N6843, N6832, N3894, N904, N497);
or OR2 (N6844, N6830, N5129);
or OR2 (N6845, N6833, N35);
and AND2 (N6846, N6844, N1611);
nand NAND3 (N6847, N6822, N1626, N2984);
nor NOR3 (N6848, N6841, N410, N5196);
nor NOR3 (N6849, N6825, N2232, N5076);
and AND2 (N6850, N6846, N1521);
and AND3 (N6851, N6847, N3325, N5744);
xor XOR2 (N6852, N6849, N3460);
and AND2 (N6853, N6850, N727);
and AND2 (N6854, N6843, N2098);
or OR3 (N6855, N6852, N259, N3453);
or OR2 (N6856, N6842, N6535);
xor XOR2 (N6857, N6851, N2317);
nand NAND4 (N6858, N6857, N3572, N1727, N5690);
nor NOR3 (N6859, N6856, N6818, N995);
xor XOR2 (N6860, N6859, N3325);
and AND3 (N6861, N6854, N5146, N6551);
buf BUF1 (N6862, N6860);
buf BUF1 (N6863, N6838);
and AND4 (N6864, N6853, N2555, N2458, N3653);
xor XOR2 (N6865, N6864, N67);
buf BUF1 (N6866, N6845);
not NOT1 (N6867, N6855);
not NOT1 (N6868, N6862);
and AND3 (N6869, N6835, N4597, N33);
nor NOR4 (N6870, N6863, N5452, N4582, N3687);
not NOT1 (N6871, N6868);
nor NOR3 (N6872, N6861, N917, N193);
nor NOR4 (N6873, N6871, N3491, N2068, N1460);
nand NAND3 (N6874, N6869, N289, N2754);
buf BUF1 (N6875, N6873);
buf BUF1 (N6876, N6858);
and AND4 (N6877, N6875, N4373, N6079, N2347);
xor XOR2 (N6878, N6848, N2574);
buf BUF1 (N6879, N6872);
buf BUF1 (N6880, N6874);
nor NOR4 (N6881, N6878, N506, N5380, N1606);
or OR4 (N6882, N6840, N4881, N1463, N2817);
not NOT1 (N6883, N6865);
xor XOR2 (N6884, N6880, N4700);
nor NOR2 (N6885, N6879, N2876);
nor NOR4 (N6886, N6877, N4582, N5656, N5817);
nand NAND3 (N6887, N6886, N3667, N5944);
and AND3 (N6888, N6881, N6688, N6645);
or OR3 (N6889, N6867, N3619, N6269);
or OR4 (N6890, N6887, N1371, N2940, N1755);
and AND2 (N6891, N6884, N5710);
nor NOR4 (N6892, N6876, N3616, N2994, N4644);
xor XOR2 (N6893, N6866, N6530);
buf BUF1 (N6894, N6890);
not NOT1 (N6895, N6894);
and AND3 (N6896, N6883, N3233, N1833);
not NOT1 (N6897, N6888);
buf BUF1 (N6898, N6892);
and AND3 (N6899, N6893, N2865, N2289);
xor XOR2 (N6900, N6882, N477);
or OR4 (N6901, N6895, N62, N5818, N2174);
and AND2 (N6902, N6896, N5609);
not NOT1 (N6903, N6885);
or OR3 (N6904, N6902, N4570, N616);
nor NOR3 (N6905, N6899, N1142, N5585);
nand NAND2 (N6906, N6900, N4576);
not NOT1 (N6907, N6897);
not NOT1 (N6908, N6907);
not NOT1 (N6909, N6903);
not NOT1 (N6910, N6908);
nand NAND4 (N6911, N6906, N1963, N4254, N3192);
xor XOR2 (N6912, N6911, N1023);
xor XOR2 (N6913, N6910, N5893);
nand NAND3 (N6914, N6898, N5166, N4278);
buf BUF1 (N6915, N6904);
or OR4 (N6916, N6915, N6406, N5034, N866);
nand NAND2 (N6917, N6870, N2371);
xor XOR2 (N6918, N6914, N2618);
and AND3 (N6919, N6905, N1888, N3702);
buf BUF1 (N6920, N6909);
not NOT1 (N6921, N6891);
xor XOR2 (N6922, N6916, N2730);
nor NOR3 (N6923, N6889, N4447, N3075);
xor XOR2 (N6924, N6917, N522);
or OR4 (N6925, N6924, N6194, N181, N3625);
or OR2 (N6926, N6922, N2377);
not NOT1 (N6927, N6919);
nor NOR3 (N6928, N6901, N5616, N124);
xor XOR2 (N6929, N6913, N4402);
xor XOR2 (N6930, N6925, N1435);
buf BUF1 (N6931, N6918);
buf BUF1 (N6932, N6929);
xor XOR2 (N6933, N6927, N2764);
xor XOR2 (N6934, N6933, N4027);
xor XOR2 (N6935, N6932, N6011);
buf BUF1 (N6936, N6935);
nand NAND4 (N6937, N6921, N4481, N3005, N2558);
and AND3 (N6938, N6920, N6131, N5738);
xor XOR2 (N6939, N6936, N3567);
or OR4 (N6940, N6912, N4890, N5347, N6081);
buf BUF1 (N6941, N6931);
nor NOR2 (N6942, N6940, N2655);
not NOT1 (N6943, N6937);
xor XOR2 (N6944, N6923, N4680);
buf BUF1 (N6945, N6941);
or OR2 (N6946, N6928, N4359);
or OR4 (N6947, N6943, N5425, N872, N295);
not NOT1 (N6948, N6947);
nor NOR2 (N6949, N6942, N5459);
nand NAND3 (N6950, N6944, N3579, N4473);
xor XOR2 (N6951, N6945, N2180);
nor NOR3 (N6952, N6950, N3540, N2665);
or OR4 (N6953, N6939, N3772, N4870, N3542);
not NOT1 (N6954, N6953);
and AND4 (N6955, N6948, N2701, N541, N3417);
nor NOR2 (N6956, N6955, N1016);
and AND3 (N6957, N6949, N2558, N2577);
nor NOR4 (N6958, N6946, N3441, N3514, N6281);
nor NOR2 (N6959, N6958, N4932);
nor NOR4 (N6960, N6951, N174, N1051, N2322);
buf BUF1 (N6961, N6934);
buf BUF1 (N6962, N6959);
or OR4 (N6963, N6957, N2190, N6500, N279);
nor NOR2 (N6964, N6938, N6545);
and AND4 (N6965, N6952, N2154, N949, N4968);
nand NAND2 (N6966, N6956, N294);
nand NAND4 (N6967, N6966, N454, N3191, N2189);
nor NOR4 (N6968, N6926, N1752, N6045, N3115);
nor NOR3 (N6969, N6962, N3360, N1339);
buf BUF1 (N6970, N6969);
not NOT1 (N6971, N6967);
not NOT1 (N6972, N6960);
nor NOR2 (N6973, N6968, N107);
xor XOR2 (N6974, N6971, N2471);
or OR3 (N6975, N6964, N4251, N5933);
xor XOR2 (N6976, N6974, N1900);
buf BUF1 (N6977, N6972);
or OR2 (N6978, N6961, N4909);
not NOT1 (N6979, N6970);
nor NOR3 (N6980, N6963, N6803, N3991);
buf BUF1 (N6981, N6973);
or OR2 (N6982, N6930, N1120);
xor XOR2 (N6983, N6982, N2201);
buf BUF1 (N6984, N6981);
nor NOR4 (N6985, N6983, N5005, N3972, N6510);
or OR4 (N6986, N6965, N939, N2545, N1638);
buf BUF1 (N6987, N6985);
not NOT1 (N6988, N6984);
or OR3 (N6989, N6954, N4327, N855);
nor NOR4 (N6990, N6977, N6067, N4918, N6359);
not NOT1 (N6991, N6988);
nand NAND3 (N6992, N6980, N4, N1395);
nor NOR3 (N6993, N6975, N2742, N2184);
not NOT1 (N6994, N6976);
xor XOR2 (N6995, N6987, N3160);
nand NAND3 (N6996, N6995, N1592, N5833);
nand NAND3 (N6997, N6990, N3933, N6093);
not NOT1 (N6998, N6996);
nand NAND2 (N6999, N6992, N6488);
nand NAND4 (N7000, N6994, N6366, N1859, N137);
nand NAND4 (N7001, N7000, N2524, N1015, N4237);
or OR3 (N7002, N6997, N4431, N6181);
nand NAND3 (N7003, N7002, N3988, N5112);
buf BUF1 (N7004, N6986);
nand NAND3 (N7005, N6989, N5377, N3964);
nor NOR4 (N7006, N6998, N287, N867, N1909);
buf BUF1 (N7007, N6978);
not NOT1 (N7008, N6993);
buf BUF1 (N7009, N6999);
nor NOR3 (N7010, N7009, N1708, N297);
nor NOR4 (N7011, N7001, N1651, N6726, N2717);
buf BUF1 (N7012, N7005);
not NOT1 (N7013, N7012);
nor NOR4 (N7014, N7006, N4536, N2706, N1410);
nor NOR4 (N7015, N7014, N196, N5952, N2766);
nand NAND2 (N7016, N7011, N3964);
xor XOR2 (N7017, N7007, N3110);
nand NAND4 (N7018, N6991, N7002, N4040, N5894);
buf BUF1 (N7019, N6979);
xor XOR2 (N7020, N7010, N1796);
buf BUF1 (N7021, N7017);
buf BUF1 (N7022, N7016);
xor XOR2 (N7023, N7018, N5766);
buf BUF1 (N7024, N7023);
buf BUF1 (N7025, N7019);
not NOT1 (N7026, N7015);
or OR3 (N7027, N7013, N5579, N1718);
not NOT1 (N7028, N7008);
not NOT1 (N7029, N7021);
not NOT1 (N7030, N7003);
nand NAND4 (N7031, N7020, N1517, N4728, N4766);
xor XOR2 (N7032, N7022, N1417);
xor XOR2 (N7033, N7028, N5536);
nand NAND2 (N7034, N7032, N5380);
and AND3 (N7035, N7033, N3105, N6533);
nand NAND3 (N7036, N7027, N2300, N499);
buf BUF1 (N7037, N7031);
buf BUF1 (N7038, N7004);
xor XOR2 (N7039, N7029, N2909);
buf BUF1 (N7040, N7030);
nand NAND4 (N7041, N7035, N5339, N3586, N3113);
and AND4 (N7042, N7026, N6997, N2259, N6229);
xor XOR2 (N7043, N7024, N3649);
buf BUF1 (N7044, N7041);
not NOT1 (N7045, N7025);
or OR2 (N7046, N7043, N5153);
buf BUF1 (N7047, N7045);
xor XOR2 (N7048, N7047, N1922);
not NOT1 (N7049, N7038);
xor XOR2 (N7050, N7048, N6334);
not NOT1 (N7051, N7044);
nor NOR3 (N7052, N7036, N4130, N1216);
xor XOR2 (N7053, N7037, N1061);
xor XOR2 (N7054, N7053, N1116);
xor XOR2 (N7055, N7049, N1468);
not NOT1 (N7056, N7040);
buf BUF1 (N7057, N7055);
or OR3 (N7058, N7051, N6978, N6721);
or OR3 (N7059, N7057, N2849, N419);
not NOT1 (N7060, N7056);
or OR4 (N7061, N7046, N467, N1626, N2438);
nor NOR2 (N7062, N7059, N613);
and AND2 (N7063, N7061, N1524);
buf BUF1 (N7064, N7052);
xor XOR2 (N7065, N7034, N2052);
and AND3 (N7066, N7050, N1173, N308);
and AND2 (N7067, N7039, N1329);
or OR3 (N7068, N7064, N5682, N497);
xor XOR2 (N7069, N7062, N1249);
not NOT1 (N7070, N7068);
xor XOR2 (N7071, N7066, N1131);
nand NAND4 (N7072, N7054, N6538, N5352, N1585);
xor XOR2 (N7073, N7070, N5315);
or OR2 (N7074, N7042, N4852);
not NOT1 (N7075, N7063);
xor XOR2 (N7076, N7060, N89);
nand NAND2 (N7077, N7065, N1494);
nand NAND3 (N7078, N7071, N1340, N1516);
nand NAND3 (N7079, N7072, N5114, N6490);
and AND4 (N7080, N7074, N4626, N2602, N3503);
and AND2 (N7081, N7067, N17);
and AND3 (N7082, N7069, N2391, N1267);
not NOT1 (N7083, N7081);
buf BUF1 (N7084, N7077);
nor NOR4 (N7085, N7083, N5517, N4582, N2390);
buf BUF1 (N7086, N7084);
nor NOR2 (N7087, N7073, N4717);
nor NOR3 (N7088, N7058, N1712, N6316);
nor NOR2 (N7089, N7086, N1424);
or OR2 (N7090, N7080, N50);
not NOT1 (N7091, N7079);
not NOT1 (N7092, N7078);
and AND4 (N7093, N7075, N7072, N172, N1404);
not NOT1 (N7094, N7091);
and AND2 (N7095, N7093, N4959);
or OR4 (N7096, N7087, N4718, N1169, N2019);
not NOT1 (N7097, N7082);
buf BUF1 (N7098, N7097);
nand NAND2 (N7099, N7098, N1931);
and AND3 (N7100, N7090, N3995, N6857);
not NOT1 (N7101, N7096);
or OR2 (N7102, N7099, N2724);
nand NAND3 (N7103, N7102, N3951, N4051);
buf BUF1 (N7104, N7095);
not NOT1 (N7105, N7076);
and AND2 (N7106, N7088, N5334);
and AND4 (N7107, N7085, N3257, N2330, N1931);
buf BUF1 (N7108, N7105);
nor NOR2 (N7109, N7103, N6928);
nor NOR4 (N7110, N7108, N5714, N4695, N3232);
not NOT1 (N7111, N7092);
not NOT1 (N7112, N7110);
buf BUF1 (N7113, N7107);
and AND2 (N7114, N7112, N1136);
not NOT1 (N7115, N7100);
not NOT1 (N7116, N7106);
nor NOR2 (N7117, N7104, N3072);
not NOT1 (N7118, N7116);
buf BUF1 (N7119, N7109);
and AND2 (N7120, N7111, N1874);
and AND2 (N7121, N7115, N2031);
nor NOR2 (N7122, N7117, N5997);
not NOT1 (N7123, N7121);
or OR4 (N7124, N7119, N6814, N6772, N1725);
and AND3 (N7125, N7122, N4195, N6873);
and AND4 (N7126, N7120, N4944, N3164, N3942);
nor NOR2 (N7127, N7113, N1547);
not NOT1 (N7128, N7118);
and AND4 (N7129, N7128, N6217, N6201, N1571);
or OR3 (N7130, N7125, N1309, N5103);
and AND2 (N7131, N7126, N4645);
buf BUF1 (N7132, N7127);
xor XOR2 (N7133, N7131, N6186);
nor NOR4 (N7134, N7133, N2426, N1648, N6001);
buf BUF1 (N7135, N7130);
not NOT1 (N7136, N7132);
buf BUF1 (N7137, N7089);
and AND3 (N7138, N7137, N5007, N1398);
nor NOR4 (N7139, N7114, N1670, N6089, N4808);
nand NAND3 (N7140, N7129, N3315, N5514);
not NOT1 (N7141, N7140);
nand NAND4 (N7142, N7124, N5307, N4657, N3265);
nor NOR4 (N7143, N7134, N6361, N4223, N2139);
nand NAND4 (N7144, N7094, N3612, N2985, N7046);
nand NAND3 (N7145, N7142, N6359, N2803);
xor XOR2 (N7146, N7144, N2713);
nand NAND4 (N7147, N7143, N2629, N2762, N2103);
not NOT1 (N7148, N7146);
or OR3 (N7149, N7145, N476, N1841);
or OR4 (N7150, N7148, N2094, N6623, N402);
or OR2 (N7151, N7139, N1082);
nand NAND4 (N7152, N7135, N735, N1722, N2974);
buf BUF1 (N7153, N7123);
nor NOR2 (N7154, N7152, N86);
xor XOR2 (N7155, N7149, N4315);
and AND2 (N7156, N7101, N289);
nand NAND4 (N7157, N7147, N3373, N4379, N2807);
xor XOR2 (N7158, N7136, N6701);
buf BUF1 (N7159, N7151);
and AND4 (N7160, N7156, N3023, N6802, N3422);
nor NOR3 (N7161, N7154, N5352, N4638);
not NOT1 (N7162, N7160);
nand NAND3 (N7163, N7161, N2626, N6418);
and AND4 (N7164, N7153, N3493, N3731, N4569);
nand NAND2 (N7165, N7141, N3953);
or OR2 (N7166, N7165, N6703);
buf BUF1 (N7167, N7159);
nand NAND3 (N7168, N7158, N4012, N3643);
not NOT1 (N7169, N7168);
buf BUF1 (N7170, N7164);
and AND4 (N7171, N7167, N4083, N3700, N6506);
nand NAND4 (N7172, N7163, N6441, N4121, N747);
xor XOR2 (N7173, N7162, N4112);
nand NAND3 (N7174, N7170, N282, N5569);
nand NAND4 (N7175, N7171, N5965, N3605, N853);
nor NOR3 (N7176, N7175, N2497, N1993);
or OR3 (N7177, N7176, N5363, N3569);
buf BUF1 (N7178, N7174);
and AND3 (N7179, N7138, N2440, N482);
buf BUF1 (N7180, N7155);
or OR2 (N7181, N7178, N321);
buf BUF1 (N7182, N7166);
not NOT1 (N7183, N7179);
nor NOR4 (N7184, N7172, N4306, N4687, N4674);
nor NOR2 (N7185, N7183, N4577);
and AND4 (N7186, N7150, N602, N5495, N640);
nor NOR2 (N7187, N7180, N3733);
xor XOR2 (N7188, N7184, N1975);
nor NOR4 (N7189, N7169, N6115, N1239, N5396);
nand NAND4 (N7190, N7188, N3123, N3324, N4394);
not NOT1 (N7191, N7173);
xor XOR2 (N7192, N7190, N4258);
nand NAND2 (N7193, N7187, N3166);
buf BUF1 (N7194, N7177);
xor XOR2 (N7195, N7189, N445);
and AND4 (N7196, N7192, N4506, N6785, N6247);
nand NAND3 (N7197, N7182, N6021, N6677);
buf BUF1 (N7198, N7181);
not NOT1 (N7199, N7195);
not NOT1 (N7200, N7199);
buf BUF1 (N7201, N7191);
xor XOR2 (N7202, N7157, N2712);
nor NOR3 (N7203, N7196, N1801, N2975);
or OR2 (N7204, N7193, N6263);
and AND3 (N7205, N7204, N1460, N4899);
nor NOR2 (N7206, N7201, N2534);
nor NOR4 (N7207, N7203, N1050, N237, N3287);
nand NAND4 (N7208, N7194, N3132, N3756, N794);
and AND3 (N7209, N7185, N6892, N5088);
xor XOR2 (N7210, N7208, N2886);
and AND3 (N7211, N7186, N2268, N2317);
and AND2 (N7212, N7198, N2383);
nand NAND4 (N7213, N7212, N5482, N7162, N3615);
nand NAND4 (N7214, N7202, N4572, N2479, N6472);
xor XOR2 (N7215, N7213, N4417);
buf BUF1 (N7216, N7215);
nor NOR4 (N7217, N7214, N6118, N6281, N5653);
and AND4 (N7218, N7200, N3753, N4282, N4160);
buf BUF1 (N7219, N7207);
buf BUF1 (N7220, N7218);
or OR4 (N7221, N7197, N2645, N1759, N6437);
or OR3 (N7222, N7209, N152, N5071);
xor XOR2 (N7223, N7216, N1331);
xor XOR2 (N7224, N7220, N6543);
or OR4 (N7225, N7210, N3374, N3742, N423);
xor XOR2 (N7226, N7224, N4381);
or OR3 (N7227, N7211, N3295, N2640);
nand NAND3 (N7228, N7222, N6316, N1040);
and AND4 (N7229, N7223, N5989, N602, N5361);
and AND3 (N7230, N7227, N1449, N6428);
xor XOR2 (N7231, N7205, N4933);
buf BUF1 (N7232, N7228);
and AND3 (N7233, N7232, N2094, N3994);
not NOT1 (N7234, N7229);
or OR3 (N7235, N7230, N1823, N5862);
and AND2 (N7236, N7225, N4589);
buf BUF1 (N7237, N7217);
nand NAND4 (N7238, N7235, N4846, N2908, N2656);
nand NAND3 (N7239, N7236, N5759, N2654);
xor XOR2 (N7240, N7238, N6044);
buf BUF1 (N7241, N7240);
or OR2 (N7242, N7221, N6584);
not NOT1 (N7243, N7241);
or OR4 (N7244, N7239, N6539, N3372, N4267);
or OR2 (N7245, N7226, N4710);
and AND4 (N7246, N7243, N943, N2621, N1799);
nor NOR4 (N7247, N7237, N6965, N1443, N150);
and AND3 (N7248, N7233, N220, N6197);
nand NAND3 (N7249, N7245, N6056, N1873);
and AND4 (N7250, N7246, N2303, N4556, N2750);
or OR3 (N7251, N7219, N1976, N5803);
nor NOR4 (N7252, N7250, N4770, N1486, N423);
nor NOR4 (N7253, N7206, N3892, N2282, N4090);
nand NAND2 (N7254, N7252, N1809);
or OR2 (N7255, N7231, N3129);
and AND3 (N7256, N7254, N1962, N2563);
not NOT1 (N7257, N7234);
xor XOR2 (N7258, N7253, N2928);
nor NOR4 (N7259, N7257, N2066, N5767, N3090);
not NOT1 (N7260, N7242);
nor NOR3 (N7261, N7256, N4665, N3780);
or OR3 (N7262, N7259, N3073, N6261);
buf BUF1 (N7263, N7249);
or OR3 (N7264, N7251, N26, N2233);
xor XOR2 (N7265, N7248, N23);
buf BUF1 (N7266, N7264);
nand NAND3 (N7267, N7258, N1108, N2517);
xor XOR2 (N7268, N7265, N4452);
nor NOR3 (N7269, N7262, N2346, N5733);
buf BUF1 (N7270, N7244);
not NOT1 (N7271, N7255);
and AND3 (N7272, N7267, N5940, N3605);
not NOT1 (N7273, N7260);
nand NAND3 (N7274, N7261, N4863, N5033);
and AND2 (N7275, N7269, N831);
not NOT1 (N7276, N7273);
nor NOR3 (N7277, N7271, N2290, N6813);
nand NAND2 (N7278, N7277, N1744);
not NOT1 (N7279, N7275);
nor NOR2 (N7280, N7272, N310);
xor XOR2 (N7281, N7263, N6438);
and AND4 (N7282, N7278, N4793, N437, N1213);
not NOT1 (N7283, N7268);
buf BUF1 (N7284, N7282);
nor NOR2 (N7285, N7270, N3071);
and AND3 (N7286, N7279, N702, N435);
or OR3 (N7287, N7281, N6603, N1663);
nor NOR3 (N7288, N7283, N771, N4142);
not NOT1 (N7289, N7276);
not NOT1 (N7290, N7285);
or OR2 (N7291, N7280, N4965);
or OR2 (N7292, N7288, N4827);
and AND4 (N7293, N7247, N4827, N4062, N1947);
nor NOR2 (N7294, N7266, N5196);
and AND3 (N7295, N7289, N4056, N651);
not NOT1 (N7296, N7287);
or OR3 (N7297, N7286, N5054, N3592);
buf BUF1 (N7298, N7295);
not NOT1 (N7299, N7297);
and AND3 (N7300, N7284, N4955, N1177);
not NOT1 (N7301, N7291);
xor XOR2 (N7302, N7293, N5202);
nand NAND4 (N7303, N7300, N5709, N6588, N4089);
nand NAND4 (N7304, N7296, N3009, N7082, N1179);
xor XOR2 (N7305, N7299, N6160);
or OR3 (N7306, N7290, N3790, N1511);
or OR4 (N7307, N7303, N3732, N2093, N5099);
and AND4 (N7308, N7298, N7208, N4240, N1411);
or OR3 (N7309, N7305, N4263, N6725);
or OR4 (N7310, N7294, N6067, N3536, N3697);
or OR2 (N7311, N7301, N3451);
not NOT1 (N7312, N7310);
nor NOR3 (N7313, N7307, N2158, N7049);
and AND2 (N7314, N7308, N3356);
buf BUF1 (N7315, N7309);
nor NOR4 (N7316, N7306, N5598, N688, N4957);
nand NAND3 (N7317, N7304, N5601, N857);
not NOT1 (N7318, N7274);
xor XOR2 (N7319, N7313, N923);
or OR4 (N7320, N7318, N1192, N2622, N780);
buf BUF1 (N7321, N7319);
xor XOR2 (N7322, N7311, N4321);
nor NOR4 (N7323, N7320, N3356, N3949, N2237);
and AND3 (N7324, N7321, N27, N3027);
nor NOR2 (N7325, N7324, N4486);
nor NOR3 (N7326, N7312, N3447, N4382);
and AND3 (N7327, N7292, N295, N5824);
buf BUF1 (N7328, N7326);
xor XOR2 (N7329, N7328, N119);
nor NOR3 (N7330, N7322, N3320, N623);
nor NOR3 (N7331, N7316, N6364, N3792);
not NOT1 (N7332, N7329);
buf BUF1 (N7333, N7327);
or OR4 (N7334, N7325, N2431, N1126, N402);
buf BUF1 (N7335, N7314);
nand NAND4 (N7336, N7315, N253, N4004, N5158);
and AND4 (N7337, N7336, N3582, N1626, N6246);
or OR2 (N7338, N7334, N1269);
or OR3 (N7339, N7323, N1404, N296);
not NOT1 (N7340, N7339);
and AND2 (N7341, N7302, N4928);
nand NAND2 (N7342, N7330, N5115);
and AND4 (N7343, N7335, N1254, N2442, N5808);
and AND2 (N7344, N7343, N6292);
not NOT1 (N7345, N7338);
not NOT1 (N7346, N7317);
or OR4 (N7347, N7345, N2271, N437, N5165);
buf BUF1 (N7348, N7333);
nand NAND3 (N7349, N7347, N1579, N6280);
xor XOR2 (N7350, N7344, N1360);
xor XOR2 (N7351, N7342, N5956);
or OR2 (N7352, N7349, N4906);
nand NAND3 (N7353, N7348, N5732, N5374);
not NOT1 (N7354, N7340);
and AND4 (N7355, N7346, N4464, N2516, N1402);
buf BUF1 (N7356, N7354);
or OR4 (N7357, N7332, N2627, N140, N5681);
nor NOR2 (N7358, N7356, N132);
nand NAND4 (N7359, N7350, N4476, N539, N4882);
not NOT1 (N7360, N7341);
and AND4 (N7361, N7359, N1288, N6409, N1763);
nor NOR3 (N7362, N7337, N2235, N2421);
nand NAND2 (N7363, N7351, N854);
nand NAND2 (N7364, N7352, N7190);
not NOT1 (N7365, N7357);
buf BUF1 (N7366, N7364);
nor NOR4 (N7367, N7366, N3538, N5837, N4522);
or OR3 (N7368, N7360, N1818, N1803);
nor NOR2 (N7369, N7358, N772);
nor NOR3 (N7370, N7367, N3145, N155);
xor XOR2 (N7371, N7363, N4616);
not NOT1 (N7372, N7370);
not NOT1 (N7373, N7361);
nor NOR2 (N7374, N7355, N3488);
not NOT1 (N7375, N7331);
nand NAND4 (N7376, N7372, N3504, N1044, N7326);
not NOT1 (N7377, N7362);
xor XOR2 (N7378, N7368, N2026);
buf BUF1 (N7379, N7369);
xor XOR2 (N7380, N7376, N1654);
buf BUF1 (N7381, N7371);
or OR4 (N7382, N7381, N221, N231, N6346);
not NOT1 (N7383, N7374);
xor XOR2 (N7384, N7373, N5966);
xor XOR2 (N7385, N7353, N305);
buf BUF1 (N7386, N7379);
nor NOR2 (N7387, N7377, N4124);
or OR2 (N7388, N7387, N6545);
nor NOR4 (N7389, N7378, N3016, N2356, N6015);
nor NOR3 (N7390, N7383, N7094, N4600);
not NOT1 (N7391, N7375);
not NOT1 (N7392, N7384);
xor XOR2 (N7393, N7391, N6813);
not NOT1 (N7394, N7392);
and AND3 (N7395, N7394, N127, N962);
xor XOR2 (N7396, N7386, N181);
and AND2 (N7397, N7365, N4183);
xor XOR2 (N7398, N7393, N3618);
or OR3 (N7399, N7396, N3390, N2795);
not NOT1 (N7400, N7380);
nor NOR4 (N7401, N7388, N6928, N4589, N408);
nand NAND2 (N7402, N7400, N3311);
and AND2 (N7403, N7390, N113);
buf BUF1 (N7404, N7401);
buf BUF1 (N7405, N7382);
nand NAND3 (N7406, N7389, N6093, N2408);
or OR2 (N7407, N7403, N1843);
or OR2 (N7408, N7407, N6457);
not NOT1 (N7409, N7405);
or OR3 (N7410, N7406, N4195, N1110);
xor XOR2 (N7411, N7395, N684);
buf BUF1 (N7412, N7408);
buf BUF1 (N7413, N7412);
xor XOR2 (N7414, N7385, N517);
nand NAND3 (N7415, N7399, N6527, N2018);
or OR3 (N7416, N7413, N6570, N3852);
xor XOR2 (N7417, N7416, N6911);
and AND2 (N7418, N7410, N5171);
and AND4 (N7419, N7418, N826, N2599, N3105);
or OR4 (N7420, N7411, N411, N4234, N3818);
xor XOR2 (N7421, N7404, N1567);
nor NOR2 (N7422, N7420, N3237);
not NOT1 (N7423, N7419);
nand NAND4 (N7424, N7422, N2946, N2074, N3482);
nand NAND2 (N7425, N7414, N6130);
xor XOR2 (N7426, N7415, N5029);
nand NAND2 (N7427, N7421, N5141);
not NOT1 (N7428, N7424);
xor XOR2 (N7429, N7428, N7393);
xor XOR2 (N7430, N7425, N6393);
and AND2 (N7431, N7417, N5805);
nor NOR4 (N7432, N7427, N2903, N5692, N3065);
nor NOR2 (N7433, N7431, N2705);
and AND2 (N7434, N7409, N1261);
nand NAND3 (N7435, N7430, N3091, N1474);
nand NAND3 (N7436, N7434, N4764, N641);
nand NAND4 (N7437, N7432, N1922, N5217, N3054);
nor NOR2 (N7438, N7423, N5846);
and AND4 (N7439, N7398, N5839, N1520, N6835);
and AND4 (N7440, N7397, N7381, N2989, N337);
nand NAND2 (N7441, N7433, N2051);
not NOT1 (N7442, N7439);
nor NOR2 (N7443, N7402, N6651);
nand NAND3 (N7444, N7438, N4481, N3176);
or OR3 (N7445, N7429, N5778, N2049);
or OR4 (N7446, N7444, N13, N4443, N3578);
and AND4 (N7447, N7440, N7045, N5818, N571);
nor NOR4 (N7448, N7441, N5851, N690, N6271);
not NOT1 (N7449, N7443);
nor NOR4 (N7450, N7437, N318, N1522, N5163);
xor XOR2 (N7451, N7436, N2585);
buf BUF1 (N7452, N7435);
not NOT1 (N7453, N7426);
nor NOR4 (N7454, N7452, N3982, N4654, N6688);
xor XOR2 (N7455, N7447, N2895);
and AND3 (N7456, N7445, N6195, N2052);
xor XOR2 (N7457, N7449, N1536);
or OR3 (N7458, N7442, N489, N1935);
or OR3 (N7459, N7448, N762, N5647);
nand NAND2 (N7460, N7451, N2540);
not NOT1 (N7461, N7457);
or OR4 (N7462, N7455, N4139, N2136, N720);
or OR2 (N7463, N7450, N1281);
xor XOR2 (N7464, N7461, N4136);
or OR3 (N7465, N7453, N2319, N3580);
nor NOR3 (N7466, N7459, N4641, N6904);
nor NOR3 (N7467, N7462, N6404, N4948);
not NOT1 (N7468, N7467);
or OR2 (N7469, N7465, N7381);
buf BUF1 (N7470, N7458);
nand NAND2 (N7471, N7460, N2180);
or OR3 (N7472, N7466, N1387, N3056);
xor XOR2 (N7473, N7456, N4546);
xor XOR2 (N7474, N7468, N4567);
not NOT1 (N7475, N7454);
nor NOR4 (N7476, N7446, N3067, N4552, N7248);
not NOT1 (N7477, N7472);
xor XOR2 (N7478, N7473, N1713);
and AND4 (N7479, N7477, N6102, N6436, N6506);
nand NAND3 (N7480, N7470, N6073, N1998);
buf BUF1 (N7481, N7478);
nand NAND3 (N7482, N7471, N5540, N3029);
nand NAND2 (N7483, N7479, N3723);
or OR2 (N7484, N7482, N2376);
xor XOR2 (N7485, N7483, N7001);
nor NOR4 (N7486, N7485, N2167, N5021, N5680);
buf BUF1 (N7487, N7474);
and AND4 (N7488, N7475, N4741, N2484, N3364);
and AND3 (N7489, N7488, N3685, N1995);
nand NAND2 (N7490, N7469, N797);
nor NOR2 (N7491, N7480, N6838);
or OR2 (N7492, N7490, N1583);
nand NAND3 (N7493, N7489, N1249, N2388);
or OR4 (N7494, N7492, N5672, N216, N2563);
nand NAND4 (N7495, N7487, N2021, N2396, N1049);
xor XOR2 (N7496, N7495, N2923);
nor NOR2 (N7497, N7491, N3174);
buf BUF1 (N7498, N7464);
or OR4 (N7499, N7493, N5002, N5045, N3093);
not NOT1 (N7500, N7494);
or OR3 (N7501, N7498, N6613, N1309);
nor NOR4 (N7502, N7463, N4852, N1740, N7410);
not NOT1 (N7503, N7496);
buf BUF1 (N7504, N7481);
buf BUF1 (N7505, N7501);
and AND2 (N7506, N7500, N4054);
nand NAND4 (N7507, N7502, N1718, N5351, N6419);
buf BUF1 (N7508, N7507);
not NOT1 (N7509, N7506);
or OR3 (N7510, N7486, N6989, N7319);
buf BUF1 (N7511, N7497);
and AND2 (N7512, N7510, N2554);
not NOT1 (N7513, N7511);
buf BUF1 (N7514, N7513);
xor XOR2 (N7515, N7509, N4895);
not NOT1 (N7516, N7508);
or OR4 (N7517, N7484, N519, N1289, N3314);
nand NAND3 (N7518, N7516, N6376, N6081);
buf BUF1 (N7519, N7476);
xor XOR2 (N7520, N7504, N3565);
not NOT1 (N7521, N7512);
nand NAND2 (N7522, N7505, N6117);
and AND2 (N7523, N7520, N6070);
nand NAND2 (N7524, N7514, N163);
buf BUF1 (N7525, N7515);
buf BUF1 (N7526, N7499);
or OR2 (N7527, N7525, N787);
nor NOR4 (N7528, N7518, N6701, N5551, N204);
and AND3 (N7529, N7526, N4815, N4985);
nand NAND3 (N7530, N7527, N2155, N7183);
not NOT1 (N7531, N7503);
buf BUF1 (N7532, N7522);
and AND3 (N7533, N7532, N1534, N6476);
nand NAND4 (N7534, N7517, N5377, N7249, N3929);
not NOT1 (N7535, N7524);
nand NAND3 (N7536, N7529, N1840, N1875);
not NOT1 (N7537, N7536);
and AND4 (N7538, N7535, N2924, N3403, N1259);
buf BUF1 (N7539, N7534);
not NOT1 (N7540, N7521);
buf BUF1 (N7541, N7540);
xor XOR2 (N7542, N7538, N47);
and AND3 (N7543, N7519, N6586, N465);
not NOT1 (N7544, N7531);
and AND3 (N7545, N7542, N408, N3470);
xor XOR2 (N7546, N7545, N818);
nor NOR2 (N7547, N7537, N2918);
buf BUF1 (N7548, N7541);
buf BUF1 (N7549, N7528);
nand NAND4 (N7550, N7548, N567, N2852, N683);
nor NOR4 (N7551, N7550, N3766, N1015, N5019);
not NOT1 (N7552, N7546);
nand NAND2 (N7553, N7547, N2132);
or OR4 (N7554, N7543, N3327, N6518, N2468);
nor NOR4 (N7555, N7523, N5528, N4810, N2137);
buf BUF1 (N7556, N7554);
xor XOR2 (N7557, N7553, N5445);
or OR4 (N7558, N7549, N1834, N5136, N7205);
or OR4 (N7559, N7558, N5795, N1245, N6762);
buf BUF1 (N7560, N7555);
not NOT1 (N7561, N7551);
buf BUF1 (N7562, N7552);
nor NOR4 (N7563, N7562, N6343, N2240, N5093);
and AND4 (N7564, N7560, N6729, N2637, N701);
or OR4 (N7565, N7561, N1365, N3752, N1396);
nor NOR3 (N7566, N7565, N3192, N3158);
xor XOR2 (N7567, N7557, N48);
and AND2 (N7568, N7539, N3251);
and AND4 (N7569, N7559, N1383, N4957, N2394);
nand NAND2 (N7570, N7567, N1201);
or OR2 (N7571, N7530, N3285);
nand NAND2 (N7572, N7556, N6257);
nor NOR2 (N7573, N7533, N1135);
and AND3 (N7574, N7573, N558, N284);
not NOT1 (N7575, N7572);
xor XOR2 (N7576, N7569, N3164);
nand NAND4 (N7577, N7575, N620, N3302, N1294);
buf BUF1 (N7578, N7563);
nor NOR3 (N7579, N7577, N1327, N6951);
nand NAND3 (N7580, N7579, N680, N2302);
and AND3 (N7581, N7564, N1641, N7029);
not NOT1 (N7582, N7578);
xor XOR2 (N7583, N7582, N3424);
or OR4 (N7584, N7576, N3747, N4627, N4726);
not NOT1 (N7585, N7568);
nor NOR2 (N7586, N7581, N119);
or OR4 (N7587, N7544, N5818, N3535, N1247);
and AND2 (N7588, N7580, N3234);
not NOT1 (N7589, N7574);
or OR3 (N7590, N7584, N3188, N164);
nor NOR3 (N7591, N7570, N6777, N5739);
and AND4 (N7592, N7571, N1858, N4184, N5922);
nand NAND2 (N7593, N7591, N5582);
nand NAND4 (N7594, N7588, N731, N2977, N3320);
and AND2 (N7595, N7566, N4441);
buf BUF1 (N7596, N7589);
nor NOR4 (N7597, N7583, N3707, N3151, N4667);
and AND2 (N7598, N7587, N5107);
xor XOR2 (N7599, N7595, N237);
or OR4 (N7600, N7593, N4727, N3379, N1526);
buf BUF1 (N7601, N7592);
xor XOR2 (N7602, N7586, N6833);
nand NAND2 (N7603, N7594, N5087);
and AND2 (N7604, N7585, N2387);
buf BUF1 (N7605, N7598);
not NOT1 (N7606, N7600);
nor NOR2 (N7607, N7590, N3486);
buf BUF1 (N7608, N7604);
nand NAND4 (N7609, N7599, N5723, N1109, N5072);
not NOT1 (N7610, N7609);
buf BUF1 (N7611, N7601);
buf BUF1 (N7612, N7602);
nor NOR4 (N7613, N7608, N2088, N7204, N1910);
nor NOR4 (N7614, N7612, N4956, N3310, N5277);
not NOT1 (N7615, N7607);
nand NAND2 (N7616, N7610, N6358);
nor NOR4 (N7617, N7616, N2689, N3947, N3599);
or OR3 (N7618, N7605, N435, N6438);
xor XOR2 (N7619, N7618, N6946);
buf BUF1 (N7620, N7614);
and AND2 (N7621, N7603, N8);
not NOT1 (N7622, N7619);
nand NAND4 (N7623, N7597, N2712, N6079, N4779);
not NOT1 (N7624, N7615);
nand NAND3 (N7625, N7624, N3366, N2766);
or OR4 (N7626, N7622, N1566, N5793, N6113);
nand NAND4 (N7627, N7621, N1387, N707, N4282);
not NOT1 (N7628, N7625);
or OR3 (N7629, N7606, N7237, N1382);
nor NOR3 (N7630, N7617, N5909, N7234);
not NOT1 (N7631, N7623);
nand NAND4 (N7632, N7628, N1756, N7182, N1415);
buf BUF1 (N7633, N7611);
xor XOR2 (N7634, N7626, N5135);
nor NOR2 (N7635, N7634, N7413);
nand NAND4 (N7636, N7613, N1735, N3142, N1247);
or OR4 (N7637, N7630, N6096, N6680, N6648);
not NOT1 (N7638, N7620);
not NOT1 (N7639, N7633);
and AND4 (N7640, N7596, N1980, N5844, N4637);
or OR2 (N7641, N7635, N5713);
or OR3 (N7642, N7629, N1604, N7040);
and AND4 (N7643, N7627, N3721, N3077, N1169);
buf BUF1 (N7644, N7641);
xor XOR2 (N7645, N7638, N958);
nand NAND4 (N7646, N7643, N2479, N3905, N7557);
xor XOR2 (N7647, N7646, N3639);
nand NAND2 (N7648, N7636, N1459);
not NOT1 (N7649, N7632);
buf BUF1 (N7650, N7645);
not NOT1 (N7651, N7640);
nand NAND2 (N7652, N7639, N4410);
not NOT1 (N7653, N7650);
nand NAND2 (N7654, N7653, N3756);
nand NAND3 (N7655, N7651, N7120, N7042);
or OR2 (N7656, N7654, N1524);
xor XOR2 (N7657, N7631, N4094);
buf BUF1 (N7658, N7648);
or OR2 (N7659, N7652, N6500);
nor NOR4 (N7660, N7655, N4171, N2925, N212);
or OR2 (N7661, N7660, N4163);
nand NAND4 (N7662, N7644, N6071, N265, N4452);
nor NOR3 (N7663, N7642, N2036, N34);
nor NOR4 (N7664, N7659, N5328, N4775, N5045);
buf BUF1 (N7665, N7661);
or OR2 (N7666, N7664, N6318);
buf BUF1 (N7667, N7666);
nand NAND2 (N7668, N7647, N6443);
or OR2 (N7669, N7657, N2274);
not NOT1 (N7670, N7668);
or OR2 (N7671, N7669, N1068);
and AND3 (N7672, N7656, N7393, N5300);
nand NAND3 (N7673, N7667, N2167, N6945);
nand NAND3 (N7674, N7671, N6769, N3911);
buf BUF1 (N7675, N7665);
buf BUF1 (N7676, N7675);
and AND2 (N7677, N7637, N94);
not NOT1 (N7678, N7662);
nand NAND3 (N7679, N7676, N4836, N5791);
not NOT1 (N7680, N7673);
buf BUF1 (N7681, N7680);
or OR4 (N7682, N7674, N3551, N763, N7476);
buf BUF1 (N7683, N7677);
not NOT1 (N7684, N7678);
nor NOR2 (N7685, N7679, N6919);
nand NAND3 (N7686, N7658, N3522, N6207);
or OR2 (N7687, N7686, N2283);
buf BUF1 (N7688, N7663);
nor NOR2 (N7689, N7670, N1649);
buf BUF1 (N7690, N7687);
xor XOR2 (N7691, N7682, N667);
xor XOR2 (N7692, N7690, N6203);
or OR2 (N7693, N7692, N3293);
xor XOR2 (N7694, N7685, N3843);
not NOT1 (N7695, N7694);
or OR3 (N7696, N7688, N1606, N474);
and AND4 (N7697, N7696, N5240, N5349, N441);
nor NOR4 (N7698, N7672, N3578, N2320, N2826);
not NOT1 (N7699, N7684);
not NOT1 (N7700, N7691);
or OR3 (N7701, N7693, N1563, N4725);
or OR3 (N7702, N7681, N6350, N5245);
or OR2 (N7703, N7702, N7549);
xor XOR2 (N7704, N7689, N759);
xor XOR2 (N7705, N7703, N7170);
buf BUF1 (N7706, N7697);
nor NOR3 (N7707, N7649, N593, N44);
nand NAND4 (N7708, N7695, N5574, N1779, N5118);
buf BUF1 (N7709, N7708);
nand NAND4 (N7710, N7705, N538, N1952, N5213);
xor XOR2 (N7711, N7699, N1065);
or OR2 (N7712, N7701, N4914);
and AND4 (N7713, N7710, N4619, N3009, N1006);
or OR2 (N7714, N7698, N6057);
not NOT1 (N7715, N7700);
not NOT1 (N7716, N7707);
not NOT1 (N7717, N7712);
nand NAND4 (N7718, N7709, N1490, N7335, N2017);
not NOT1 (N7719, N7706);
or OR2 (N7720, N7717, N2008);
nor NOR3 (N7721, N7719, N4001, N5431);
and AND3 (N7722, N7711, N1157, N6574);
xor XOR2 (N7723, N7715, N5465);
or OR4 (N7724, N7716, N5959, N3691, N5728);
xor XOR2 (N7725, N7723, N4248);
not NOT1 (N7726, N7704);
or OR2 (N7727, N7720, N31);
buf BUF1 (N7728, N7713);
nor NOR3 (N7729, N7718, N2038, N2627);
xor XOR2 (N7730, N7729, N1687);
not NOT1 (N7731, N7730);
or OR2 (N7732, N7714, N21);
not NOT1 (N7733, N7721);
buf BUF1 (N7734, N7726);
xor XOR2 (N7735, N7728, N1610);
nor NOR3 (N7736, N7734, N7131, N1697);
not NOT1 (N7737, N7725);
nor NOR2 (N7738, N7727, N6524);
nand NAND3 (N7739, N7738, N2629, N1283);
or OR3 (N7740, N7722, N3865, N2132);
or OR3 (N7741, N7739, N4732, N6511);
xor XOR2 (N7742, N7740, N3771);
nor NOR4 (N7743, N7724, N6865, N1687, N4386);
not NOT1 (N7744, N7735);
buf BUF1 (N7745, N7683);
xor XOR2 (N7746, N7736, N5618);
or OR2 (N7747, N7737, N1708);
buf BUF1 (N7748, N7745);
buf BUF1 (N7749, N7733);
xor XOR2 (N7750, N7748, N5964);
nor NOR3 (N7751, N7742, N1252, N6307);
nor NOR2 (N7752, N7732, N4785);
not NOT1 (N7753, N7750);
buf BUF1 (N7754, N7751);
and AND2 (N7755, N7746, N6229);
xor XOR2 (N7756, N7731, N5674);
buf BUF1 (N7757, N7744);
buf BUF1 (N7758, N7753);
and AND3 (N7759, N7757, N4285, N1723);
or OR4 (N7760, N7741, N4121, N2389, N3088);
not NOT1 (N7761, N7755);
or OR4 (N7762, N7756, N1885, N7696, N1369);
xor XOR2 (N7763, N7747, N350);
xor XOR2 (N7764, N7758, N6744);
or OR2 (N7765, N7749, N5068);
and AND4 (N7766, N7760, N3561, N3203, N3951);
xor XOR2 (N7767, N7762, N6321);
nand NAND3 (N7768, N7767, N6609, N916);
buf BUF1 (N7769, N7759);
nor NOR3 (N7770, N7768, N5980, N1676);
buf BUF1 (N7771, N7754);
not NOT1 (N7772, N7764);
or OR4 (N7773, N7770, N3411, N416, N4033);
nand NAND4 (N7774, N7772, N101, N6119, N3526);
not NOT1 (N7775, N7763);
nand NAND4 (N7776, N7765, N6355, N4184, N5788);
xor XOR2 (N7777, N7769, N1322);
not NOT1 (N7778, N7775);
nor NOR4 (N7779, N7771, N5688, N1279, N1747);
and AND2 (N7780, N7774, N6175);
not NOT1 (N7781, N7777);
or OR2 (N7782, N7778, N656);
nand NAND4 (N7783, N7761, N5113, N715, N725);
nor NOR3 (N7784, N7776, N4311, N5193);
nand NAND3 (N7785, N7752, N2441, N2802);
not NOT1 (N7786, N7779);
not NOT1 (N7787, N7784);
xor XOR2 (N7788, N7786, N1632);
not NOT1 (N7789, N7743);
nand NAND2 (N7790, N7787, N6293);
xor XOR2 (N7791, N7781, N2525);
buf BUF1 (N7792, N7785);
nand NAND4 (N7793, N7792, N430, N4504, N6379);
buf BUF1 (N7794, N7793);
nor NOR3 (N7795, N7790, N5849, N6947);
nand NAND4 (N7796, N7788, N3440, N2570, N7487);
nor NOR3 (N7797, N7782, N69, N3699);
or OR2 (N7798, N7796, N4522);
nor NOR4 (N7799, N7789, N3869, N4276, N646);
xor XOR2 (N7800, N7794, N2749);
and AND4 (N7801, N7799, N4721, N4502, N3810);
buf BUF1 (N7802, N7797);
nand NAND2 (N7803, N7800, N1164);
xor XOR2 (N7804, N7783, N5999);
or OR4 (N7805, N7804, N2144, N57, N3820);
not NOT1 (N7806, N7798);
or OR4 (N7807, N7805, N353, N7654, N591);
and AND4 (N7808, N7780, N290, N6739, N7099);
not NOT1 (N7809, N7766);
and AND2 (N7810, N7795, N6968);
or OR3 (N7811, N7809, N5017, N6139);
buf BUF1 (N7812, N7810);
buf BUF1 (N7813, N7811);
buf BUF1 (N7814, N7813);
nand NAND3 (N7815, N7812, N5561, N3580);
buf BUF1 (N7816, N7814);
xor XOR2 (N7817, N7801, N4778);
nor NOR3 (N7818, N7808, N1620, N4231);
not NOT1 (N7819, N7817);
nor NOR4 (N7820, N7802, N5846, N633, N2448);
buf BUF1 (N7821, N7816);
and AND2 (N7822, N7803, N2134);
not NOT1 (N7823, N7791);
and AND3 (N7824, N7823, N6398, N4101);
and AND4 (N7825, N7820, N5096, N2040, N2052);
nor NOR4 (N7826, N7807, N5012, N1088, N6986);
nor NOR3 (N7827, N7821, N1268, N5996);
buf BUF1 (N7828, N7824);
or OR3 (N7829, N7822, N4078, N6174);
nand NAND2 (N7830, N7825, N109);
xor XOR2 (N7831, N7819, N5482);
and AND4 (N7832, N7828, N1305, N5924, N1800);
buf BUF1 (N7833, N7829);
nand NAND4 (N7834, N7831, N3909, N6480, N3400);
buf BUF1 (N7835, N7773);
nand NAND4 (N7836, N7826, N3885, N5370, N2668);
and AND4 (N7837, N7815, N7554, N2733, N491);
nand NAND3 (N7838, N7830, N4934, N7152);
not NOT1 (N7839, N7836);
nor NOR4 (N7840, N7832, N6060, N659, N1882);
not NOT1 (N7841, N7835);
not NOT1 (N7842, N7840);
nand NAND2 (N7843, N7834, N7013);
and AND4 (N7844, N7833, N3913, N7609, N334);
nor NOR4 (N7845, N7818, N3082, N2615, N1332);
not NOT1 (N7846, N7841);
nand NAND4 (N7847, N7806, N1546, N5883, N6228);
nor NOR4 (N7848, N7845, N7079, N687, N566);
and AND2 (N7849, N7848, N5907);
buf BUF1 (N7850, N7847);
buf BUF1 (N7851, N7827);
buf BUF1 (N7852, N7837);
xor XOR2 (N7853, N7850, N1104);
buf BUF1 (N7854, N7843);
and AND3 (N7855, N7842, N7036, N7448);
nor NOR3 (N7856, N7852, N6272, N5960);
or OR2 (N7857, N7849, N6482);
not NOT1 (N7858, N7856);
or OR4 (N7859, N7839, N490, N1105, N6985);
nand NAND3 (N7860, N7853, N755, N5176);
not NOT1 (N7861, N7855);
not NOT1 (N7862, N7851);
not NOT1 (N7863, N7846);
and AND4 (N7864, N7859, N4091, N3172, N5111);
xor XOR2 (N7865, N7862, N3171);
or OR4 (N7866, N7864, N7461, N2599, N6155);
or OR3 (N7867, N7838, N28, N5267);
or OR3 (N7868, N7858, N5933, N2256);
or OR3 (N7869, N7865, N6553, N685);
buf BUF1 (N7870, N7861);
xor XOR2 (N7871, N7867, N7722);
nor NOR4 (N7872, N7870, N7700, N5002, N7185);
and AND3 (N7873, N7860, N2224, N190);
xor XOR2 (N7874, N7873, N3445);
nand NAND3 (N7875, N7863, N5284, N5835);
or OR3 (N7876, N7868, N2249, N3015);
not NOT1 (N7877, N7869);
buf BUF1 (N7878, N7876);
buf BUF1 (N7879, N7872);
nor NOR2 (N7880, N7879, N577);
or OR2 (N7881, N7866, N2479);
not NOT1 (N7882, N7844);
and AND3 (N7883, N7877, N2723, N2090);
buf BUF1 (N7884, N7878);
and AND3 (N7885, N7874, N3830, N4339);
nor NOR3 (N7886, N7871, N7026, N2559);
nor NOR4 (N7887, N7854, N3285, N4667, N3433);
nor NOR4 (N7888, N7875, N5243, N358, N5528);
nor NOR2 (N7889, N7882, N4495);
and AND4 (N7890, N7888, N4113, N1532, N6101);
or OR4 (N7891, N7880, N6514, N7190, N5728);
xor XOR2 (N7892, N7885, N4133);
and AND4 (N7893, N7889, N4760, N568, N3435);
xor XOR2 (N7894, N7891, N7533);
xor XOR2 (N7895, N7883, N973);
not NOT1 (N7896, N7857);
nor NOR3 (N7897, N7886, N5360, N2211);
nor NOR2 (N7898, N7894, N4248);
or OR3 (N7899, N7881, N451, N480);
and AND2 (N7900, N7898, N2235);
buf BUF1 (N7901, N7895);
or OR3 (N7902, N7887, N7226, N3732);
buf BUF1 (N7903, N7902);
buf BUF1 (N7904, N7896);
and AND4 (N7905, N7884, N6779, N895, N4541);
nand NAND3 (N7906, N7892, N6931, N6533);
xor XOR2 (N7907, N7904, N6096);
and AND4 (N7908, N7893, N3739, N2984, N7128);
and AND2 (N7909, N7905, N2373);
not NOT1 (N7910, N7907);
nor NOR3 (N7911, N7909, N2584, N2268);
nor NOR4 (N7912, N7906, N7678, N2148, N456);
nand NAND2 (N7913, N7899, N278);
and AND2 (N7914, N7912, N6950);
and AND4 (N7915, N7897, N4722, N7629, N2141);
nor NOR2 (N7916, N7890, N6024);
nor NOR4 (N7917, N7916, N6210, N2059, N4735);
nor NOR3 (N7918, N7917, N1903, N806);
xor XOR2 (N7919, N7903, N2342);
not NOT1 (N7920, N7915);
xor XOR2 (N7921, N7900, N4111);
and AND3 (N7922, N7919, N7255, N3543);
nand NAND2 (N7923, N7913, N4483);
or OR4 (N7924, N7921, N7777, N7666, N6523);
not NOT1 (N7925, N7911);
or OR3 (N7926, N7920, N2094, N1927);
and AND4 (N7927, N7918, N5658, N1558, N343);
xor XOR2 (N7928, N7901, N4219);
not NOT1 (N7929, N7924);
nand NAND3 (N7930, N7908, N7583, N2977);
nand NAND3 (N7931, N7914, N7857, N6825);
or OR3 (N7932, N7910, N7307, N4224);
buf BUF1 (N7933, N7928);
nor NOR3 (N7934, N7931, N3907, N1184);
xor XOR2 (N7935, N7923, N7479);
xor XOR2 (N7936, N7934, N1522);
nor NOR2 (N7937, N7936, N3433);
not NOT1 (N7938, N7937);
nand NAND2 (N7939, N7926, N1497);
and AND4 (N7940, N7925, N4619, N6323, N5209);
not NOT1 (N7941, N7939);
and AND3 (N7942, N7933, N2472, N185);
or OR2 (N7943, N7935, N6046);
nand NAND2 (N7944, N7940, N6326);
nor NOR4 (N7945, N7922, N4545, N2129, N5735);
nand NAND4 (N7946, N7941, N728, N1759, N1449);
or OR2 (N7947, N7927, N6994);
or OR3 (N7948, N7947, N5785, N5868);
and AND3 (N7949, N7942, N5289, N31);
not NOT1 (N7950, N7949);
xor XOR2 (N7951, N7948, N5598);
not NOT1 (N7952, N7938);
nand NAND4 (N7953, N7952, N736, N4002, N5567);
xor XOR2 (N7954, N7945, N1298);
nor NOR4 (N7955, N7932, N2604, N1922, N6653);
nor NOR2 (N7956, N7955, N4240);
xor XOR2 (N7957, N7950, N1606);
buf BUF1 (N7958, N7954);
and AND2 (N7959, N7944, N1919);
not NOT1 (N7960, N7958);
buf BUF1 (N7961, N7943);
not NOT1 (N7962, N7960);
buf BUF1 (N7963, N7946);
nor NOR3 (N7964, N7930, N6119, N7712);
nand NAND4 (N7965, N7962, N6635, N7726, N3033);
or OR4 (N7966, N7956, N7871, N7313, N671);
buf BUF1 (N7967, N7963);
not NOT1 (N7968, N7957);
nand NAND3 (N7969, N7968, N1110, N2610);
not NOT1 (N7970, N7953);
nor NOR3 (N7971, N7965, N5255, N3101);
buf BUF1 (N7972, N7959);
nor NOR2 (N7973, N7964, N6415);
and AND3 (N7974, N7973, N5022, N6599);
xor XOR2 (N7975, N7974, N5745);
or OR3 (N7976, N7969, N642, N49);
not NOT1 (N7977, N7961);
or OR3 (N7978, N7970, N687, N3677);
nor NOR2 (N7979, N7978, N1041);
and AND3 (N7980, N7971, N935, N6137);
not NOT1 (N7981, N7980);
buf BUF1 (N7982, N7979);
or OR3 (N7983, N7981, N4276, N1975);
not NOT1 (N7984, N7951);
or OR2 (N7985, N7977, N6804);
nor NOR4 (N7986, N7966, N2949, N5875, N407);
and AND4 (N7987, N7975, N4510, N985, N7323);
and AND4 (N7988, N7982, N3274, N5653, N5708);
nand NAND2 (N7989, N7988, N6212);
nor NOR4 (N7990, N7987, N1378, N1808, N415);
nand NAND3 (N7991, N7976, N7415, N5279);
or OR2 (N7992, N7984, N6745);
and AND2 (N7993, N7989, N5110);
nor NOR4 (N7994, N7967, N2212, N3266, N2913);
nor NOR3 (N7995, N7993, N38, N4360);
not NOT1 (N7996, N7983);
nand NAND3 (N7997, N7994, N3197, N6110);
buf BUF1 (N7998, N7929);
not NOT1 (N7999, N7986);
not NOT1 (N8000, N7997);
nand NAND3 (N8001, N7972, N843, N6582);
not NOT1 (N8002, N8000);
buf BUF1 (N8003, N8002);
nand NAND3 (N8004, N7990, N7015, N53);
not NOT1 (N8005, N7995);
or OR2 (N8006, N7992, N5330);
not NOT1 (N8007, N7999);
buf BUF1 (N8008, N8007);
and AND2 (N8009, N7996, N5323);
xor XOR2 (N8010, N8004, N7334);
buf BUF1 (N8011, N8010);
xor XOR2 (N8012, N8011, N3270);
xor XOR2 (N8013, N8006, N4534);
nor NOR2 (N8014, N8003, N3575);
nand NAND4 (N8015, N7998, N3377, N1303, N5865);
or OR3 (N8016, N8012, N7487, N4383);
buf BUF1 (N8017, N8013);
or OR3 (N8018, N8009, N2347, N6138);
not NOT1 (N8019, N7991);
nor NOR4 (N8020, N7985, N5372, N6748, N3073);
buf BUF1 (N8021, N8019);
xor XOR2 (N8022, N8021, N1550);
or OR4 (N8023, N8008, N3920, N6531, N3225);
nand NAND2 (N8024, N8015, N5201);
buf BUF1 (N8025, N8014);
or OR3 (N8026, N8024, N2040, N5466);
xor XOR2 (N8027, N8018, N1983);
and AND4 (N8028, N8016, N4759, N2955, N3612);
not NOT1 (N8029, N8026);
not NOT1 (N8030, N8028);
nor NOR3 (N8031, N8022, N3498, N2352);
nand NAND4 (N8032, N8027, N6462, N2942, N5598);
not NOT1 (N8033, N8032);
nor NOR4 (N8034, N8017, N796, N3496, N453);
nor NOR2 (N8035, N8001, N1419);
and AND4 (N8036, N8034, N6124, N1592, N5351);
xor XOR2 (N8037, N8005, N6402);
not NOT1 (N8038, N8037);
xor XOR2 (N8039, N8033, N5924);
xor XOR2 (N8040, N8020, N6882);
and AND3 (N8041, N8031, N1373, N7303);
nand NAND2 (N8042, N8036, N5245);
or OR3 (N8043, N8035, N1695, N5262);
nand NAND4 (N8044, N8042, N3713, N7853, N1710);
not NOT1 (N8045, N8030);
nand NAND2 (N8046, N8043, N2953);
and AND4 (N8047, N8038, N6304, N5785, N7150);
xor XOR2 (N8048, N8047, N6640);
and AND2 (N8049, N8044, N2144);
buf BUF1 (N8050, N8041);
or OR3 (N8051, N8046, N5840, N3331);
nor NOR3 (N8052, N8049, N4374, N1714);
not NOT1 (N8053, N8029);
or OR2 (N8054, N8045, N3389);
and AND2 (N8055, N8040, N1144);
xor XOR2 (N8056, N8054, N5965);
or OR3 (N8057, N8053, N741, N2610);
not NOT1 (N8058, N8051);
nand NAND2 (N8059, N8052, N2460);
or OR4 (N8060, N8048, N2608, N1435, N7240);
nor NOR2 (N8061, N8056, N6447);
nor NOR2 (N8062, N8061, N3684);
and AND3 (N8063, N8059, N7540, N857);
not NOT1 (N8064, N8062);
nor NOR4 (N8065, N8063, N868, N6979, N6997);
nor NOR2 (N8066, N8057, N606);
not NOT1 (N8067, N8050);
not NOT1 (N8068, N8066);
not NOT1 (N8069, N8067);
and AND2 (N8070, N8025, N907);
buf BUF1 (N8071, N8070);
nand NAND2 (N8072, N8069, N5321);
buf BUF1 (N8073, N8058);
buf BUF1 (N8074, N8064);
nor NOR2 (N8075, N8055, N2286);
nor NOR3 (N8076, N8071, N5486, N4922);
or OR3 (N8077, N8074, N5306, N6273);
or OR4 (N8078, N8072, N6140, N7805, N2933);
not NOT1 (N8079, N8039);
nand NAND4 (N8080, N8060, N3711, N5512, N7060);
and AND2 (N8081, N8078, N1181);
or OR2 (N8082, N8076, N1529);
or OR4 (N8083, N8079, N3063, N5963, N6195);
buf BUF1 (N8084, N8023);
nor NOR2 (N8085, N8083, N7851);
nand NAND4 (N8086, N8084, N5515, N2529, N3687);
and AND4 (N8087, N8082, N7887, N4833, N3406);
or OR4 (N8088, N8081, N4362, N3694, N3538);
buf BUF1 (N8089, N8088);
and AND4 (N8090, N8065, N231, N7506, N1136);
buf BUF1 (N8091, N8073);
and AND4 (N8092, N8068, N1726, N7653, N5836);
buf BUF1 (N8093, N8075);
and AND2 (N8094, N8091, N1685);
xor XOR2 (N8095, N8086, N6112);
buf BUF1 (N8096, N8077);
and AND3 (N8097, N8085, N2107, N6273);
buf BUF1 (N8098, N8087);
nor NOR2 (N8099, N8080, N7278);
not NOT1 (N8100, N8098);
xor XOR2 (N8101, N8095, N6777);
nand NAND3 (N8102, N8090, N6909, N5573);
or OR2 (N8103, N8097, N3166);
nand NAND3 (N8104, N8094, N7586, N878);
xor XOR2 (N8105, N8089, N6254);
not NOT1 (N8106, N8092);
nand NAND3 (N8107, N8100, N5514, N714);
not NOT1 (N8108, N8102);
not NOT1 (N8109, N8104);
nand NAND2 (N8110, N8108, N1198);
not NOT1 (N8111, N8099);
xor XOR2 (N8112, N8096, N2093);
xor XOR2 (N8113, N8110, N1449);
nor NOR4 (N8114, N8101, N7737, N800, N5423);
nand NAND2 (N8115, N8112, N6949);
xor XOR2 (N8116, N8113, N66);
and AND4 (N8117, N8114, N5483, N4543, N5900);
not NOT1 (N8118, N8107);
nand NAND4 (N8119, N8106, N7177, N4160, N802);
or OR4 (N8120, N8115, N3680, N4347, N1546);
xor XOR2 (N8121, N8120, N2081);
not NOT1 (N8122, N8105);
buf BUF1 (N8123, N8121);
not NOT1 (N8124, N8093);
and AND3 (N8125, N8116, N7734, N5235);
or OR3 (N8126, N8119, N7916, N7356);
xor XOR2 (N8127, N8125, N2833);
not NOT1 (N8128, N8111);
nor NOR2 (N8129, N8123, N6851);
nor NOR2 (N8130, N8109, N2256);
or OR4 (N8131, N8124, N7278, N5715, N2430);
or OR2 (N8132, N8128, N5479);
xor XOR2 (N8133, N8103, N7629);
buf BUF1 (N8134, N8133);
or OR2 (N8135, N8130, N3782);
nand NAND3 (N8136, N8131, N6968, N3562);
and AND4 (N8137, N8136, N1944, N6737, N7016);
or OR4 (N8138, N8122, N3845, N5928, N3699);
not NOT1 (N8139, N8127);
not NOT1 (N8140, N8132);
nor NOR2 (N8141, N8139, N2467);
not NOT1 (N8142, N8140);
nand NAND2 (N8143, N8135, N3188);
and AND3 (N8144, N8118, N4638, N5883);
nand NAND3 (N8145, N8129, N3091, N1165);
and AND3 (N8146, N8141, N4953, N3708);
xor XOR2 (N8147, N8138, N5835);
xor XOR2 (N8148, N8142, N6572);
nor NOR2 (N8149, N8137, N6065);
or OR2 (N8150, N8117, N4435);
xor XOR2 (N8151, N8149, N5921);
and AND3 (N8152, N8146, N148, N1983);
xor XOR2 (N8153, N8151, N4865);
nor NOR2 (N8154, N8148, N6354);
and AND2 (N8155, N8143, N6766);
nor NOR3 (N8156, N8147, N5253, N3060);
not NOT1 (N8157, N8145);
nand NAND2 (N8158, N8126, N3815);
not NOT1 (N8159, N8157);
and AND4 (N8160, N8156, N79, N6344, N3444);
not NOT1 (N8161, N8160);
and AND2 (N8162, N8134, N153);
and AND2 (N8163, N8158, N4455);
and AND2 (N8164, N8144, N4748);
buf BUF1 (N8165, N8155);
nor NOR3 (N8166, N8150, N3783, N65);
and AND3 (N8167, N8153, N2802, N6398);
not NOT1 (N8168, N8162);
not NOT1 (N8169, N8167);
xor XOR2 (N8170, N8159, N3402);
or OR3 (N8171, N8166, N6090, N4092);
nand NAND2 (N8172, N8152, N944);
not NOT1 (N8173, N8172);
or OR3 (N8174, N8165, N5193, N453);
xor XOR2 (N8175, N8171, N2791);
nor NOR4 (N8176, N8154, N1429, N5437, N3043);
or OR2 (N8177, N8174, N2641);
and AND4 (N8178, N8164, N7927, N6240, N2699);
or OR2 (N8179, N8161, N5829);
buf BUF1 (N8180, N8176);
not NOT1 (N8181, N8180);
buf BUF1 (N8182, N8173);
and AND4 (N8183, N8163, N6838, N4874, N7028);
nand NAND2 (N8184, N8183, N565);
and AND2 (N8185, N8177, N2298);
not NOT1 (N8186, N8168);
or OR4 (N8187, N8178, N7439, N1568, N2698);
buf BUF1 (N8188, N8182);
nand NAND4 (N8189, N8181, N5161, N3178, N712);
not NOT1 (N8190, N8188);
nor NOR4 (N8191, N8169, N7302, N4093, N3260);
or OR3 (N8192, N8189, N2927, N7116);
or OR4 (N8193, N8187, N6148, N8094, N7345);
nand NAND2 (N8194, N8190, N6134);
xor XOR2 (N8195, N8184, N3801);
or OR2 (N8196, N8192, N5007);
and AND4 (N8197, N8194, N2264, N2680, N1651);
not NOT1 (N8198, N8191);
nand NAND2 (N8199, N8193, N2803);
nand NAND3 (N8200, N8170, N3354, N1262);
nor NOR4 (N8201, N8195, N6313, N6735, N7726);
or OR2 (N8202, N8201, N7458);
nor NOR4 (N8203, N8175, N5309, N1214, N8171);
nand NAND3 (N8204, N8186, N602, N8115);
xor XOR2 (N8205, N8198, N558);
nor NOR3 (N8206, N8196, N4260, N472);
not NOT1 (N8207, N8185);
and AND3 (N8208, N8206, N2377, N2066);
or OR3 (N8209, N8179, N6737, N4884);
not NOT1 (N8210, N8209);
or OR4 (N8211, N8197, N2717, N3058, N1152);
xor XOR2 (N8212, N8207, N4602);
and AND4 (N8213, N8212, N5225, N7283, N512);
and AND3 (N8214, N8213, N7335, N1408);
buf BUF1 (N8215, N8202);
buf BUF1 (N8216, N8199);
buf BUF1 (N8217, N8204);
or OR4 (N8218, N8203, N636, N5852, N4299);
nor NOR3 (N8219, N8210, N1592, N3893);
buf BUF1 (N8220, N8218);
or OR3 (N8221, N8219, N5135, N7367);
buf BUF1 (N8222, N8217);
or OR3 (N8223, N8214, N6308, N4162);
and AND3 (N8224, N8220, N1356, N7215);
nor NOR3 (N8225, N8215, N6267, N5152);
nand NAND3 (N8226, N8200, N6958, N648);
buf BUF1 (N8227, N8205);
buf BUF1 (N8228, N8227);
nor NOR2 (N8229, N8216, N5711);
nand NAND4 (N8230, N8224, N7957, N3966, N952);
buf BUF1 (N8231, N8223);
nor NOR3 (N8232, N8221, N7906, N3554);
nand NAND3 (N8233, N8222, N4563, N2388);
nand NAND4 (N8234, N8211, N2542, N169, N6887);
not NOT1 (N8235, N8233);
nand NAND3 (N8236, N8228, N841, N5906);
nor NOR2 (N8237, N8229, N5892);
xor XOR2 (N8238, N8234, N4681);
not NOT1 (N8239, N8237);
xor XOR2 (N8240, N8231, N935);
nor NOR3 (N8241, N8208, N6903, N3229);
nor NOR3 (N8242, N8236, N45, N4854);
or OR2 (N8243, N8242, N1790);
nor NOR4 (N8244, N8230, N1739, N4974, N1561);
nor NOR2 (N8245, N8235, N12);
nand NAND3 (N8246, N8243, N4538, N5765);
not NOT1 (N8247, N8226);
nand NAND3 (N8248, N8241, N1348, N5374);
or OR3 (N8249, N8232, N2730, N7593);
nand NAND3 (N8250, N8240, N2577, N7144);
buf BUF1 (N8251, N8246);
nor NOR4 (N8252, N8250, N2449, N3143, N5306);
or OR4 (N8253, N8251, N7369, N627, N618);
and AND4 (N8254, N8225, N4890, N4034, N2850);
or OR2 (N8255, N8238, N6125);
or OR2 (N8256, N8247, N3448);
xor XOR2 (N8257, N8249, N2877);
xor XOR2 (N8258, N8257, N5186);
and AND3 (N8259, N8252, N1612, N6057);
buf BUF1 (N8260, N8245);
xor XOR2 (N8261, N8259, N7517);
not NOT1 (N8262, N8239);
buf BUF1 (N8263, N8256);
nor NOR3 (N8264, N8253, N4582, N3325);
buf BUF1 (N8265, N8258);
or OR3 (N8266, N8263, N1917, N3860);
nand NAND3 (N8267, N8244, N4631, N2341);
not NOT1 (N8268, N8262);
and AND2 (N8269, N8248, N1083);
nor NOR3 (N8270, N8267, N7278, N4037);
and AND4 (N8271, N8261, N770, N1118, N3397);
nor NOR4 (N8272, N8270, N3620, N4646, N5164);
xor XOR2 (N8273, N8264, N1729);
nor NOR2 (N8274, N8265, N852);
or OR2 (N8275, N8271, N3201);
xor XOR2 (N8276, N8266, N2078);
nand NAND2 (N8277, N8269, N4075);
not NOT1 (N8278, N8277);
xor XOR2 (N8279, N8273, N5358);
or OR2 (N8280, N8268, N4415);
nor NOR3 (N8281, N8260, N7845, N2335);
buf BUF1 (N8282, N8276);
not NOT1 (N8283, N8281);
and AND4 (N8284, N8272, N1624, N1252, N605);
nor NOR4 (N8285, N8275, N7271, N2773, N7279);
buf BUF1 (N8286, N8254);
or OR3 (N8287, N8284, N1132, N4187);
or OR4 (N8288, N8286, N3183, N1489, N6992);
nor NOR3 (N8289, N8283, N556, N6010);
and AND3 (N8290, N8289, N4416, N660);
and AND4 (N8291, N8282, N4480, N3222, N601);
nor NOR2 (N8292, N8279, N3488);
nor NOR3 (N8293, N8278, N4175, N2909);
or OR4 (N8294, N8287, N3155, N1862, N4747);
nand NAND3 (N8295, N8255, N3008, N5251);
nand NAND4 (N8296, N8292, N4067, N5907, N5789);
and AND4 (N8297, N8294, N3481, N4767, N7294);
nor NOR4 (N8298, N8295, N7554, N2812, N3403);
nor NOR3 (N8299, N8280, N6407, N5071);
buf BUF1 (N8300, N8288);
buf BUF1 (N8301, N8285);
xor XOR2 (N8302, N8301, N5235);
nand NAND2 (N8303, N8293, N6709);
xor XOR2 (N8304, N8290, N1747);
and AND3 (N8305, N8296, N1579, N3187);
not NOT1 (N8306, N8304);
not NOT1 (N8307, N8305);
and AND3 (N8308, N8298, N513, N7186);
nand NAND4 (N8309, N8291, N844, N7507, N1699);
buf BUF1 (N8310, N8306);
buf BUF1 (N8311, N8303);
nor NOR4 (N8312, N8307, N7466, N7137, N6189);
and AND2 (N8313, N8312, N1882);
not NOT1 (N8314, N8310);
nand NAND4 (N8315, N8308, N4137, N5223, N1298);
xor XOR2 (N8316, N8309, N6251);
xor XOR2 (N8317, N8300, N440);
not NOT1 (N8318, N8311);
buf BUF1 (N8319, N8317);
and AND2 (N8320, N8297, N75);
nor NOR4 (N8321, N8314, N6511, N7027, N5182);
and AND2 (N8322, N8319, N2004);
not NOT1 (N8323, N8274);
not NOT1 (N8324, N8315);
buf BUF1 (N8325, N8299);
and AND4 (N8326, N8322, N683, N8246, N30);
not NOT1 (N8327, N8325);
and AND3 (N8328, N8327, N3098, N8159);
nor NOR4 (N8329, N8321, N490, N1572, N5269);
or OR2 (N8330, N8313, N7571);
nand NAND2 (N8331, N8329, N3320);
nor NOR2 (N8332, N8323, N7822);
and AND3 (N8333, N8332, N107, N2613);
or OR4 (N8334, N8324, N7764, N4113, N6791);
not NOT1 (N8335, N8334);
buf BUF1 (N8336, N8335);
and AND3 (N8337, N8331, N3692, N1191);
or OR3 (N8338, N8318, N5959, N5472);
nor NOR2 (N8339, N8330, N5281);
nand NAND4 (N8340, N8337, N7718, N1713, N8271);
not NOT1 (N8341, N8316);
buf BUF1 (N8342, N8302);
xor XOR2 (N8343, N8340, N4288);
and AND3 (N8344, N8328, N1743, N2366);
nand NAND2 (N8345, N8326, N2643);
and AND2 (N8346, N8339, N7757);
and AND4 (N8347, N8338, N1789, N2443, N6759);
nor NOR3 (N8348, N8336, N7762, N1873);
nor NOR2 (N8349, N8333, N6872);
and AND3 (N8350, N8320, N5725, N714);
not NOT1 (N8351, N8346);
xor XOR2 (N8352, N8350, N1026);
nand NAND2 (N8353, N8343, N8278);
or OR3 (N8354, N8353, N1222, N377);
buf BUF1 (N8355, N8354);
or OR2 (N8356, N8342, N6555);
or OR2 (N8357, N8351, N143);
and AND4 (N8358, N8356, N4576, N5350, N4650);
or OR3 (N8359, N8344, N4777, N737);
or OR2 (N8360, N8357, N4613);
nor NOR2 (N8361, N8359, N330);
and AND3 (N8362, N8347, N6871, N3255);
not NOT1 (N8363, N8341);
and AND2 (N8364, N8355, N3051);
nor NOR2 (N8365, N8363, N4725);
not NOT1 (N8366, N8358);
not NOT1 (N8367, N8352);
and AND2 (N8368, N8345, N5928);
buf BUF1 (N8369, N8367);
nand NAND2 (N8370, N8360, N5077);
nor NOR2 (N8371, N8364, N8135);
xor XOR2 (N8372, N8349, N1264);
nand NAND3 (N8373, N8371, N2510, N2403);
nand NAND3 (N8374, N8373, N8161, N4979);
not NOT1 (N8375, N8365);
xor XOR2 (N8376, N8372, N4501);
nand NAND3 (N8377, N8375, N6130, N821);
xor XOR2 (N8378, N8374, N3131);
or OR3 (N8379, N8348, N4335, N6213);
buf BUF1 (N8380, N8379);
and AND2 (N8381, N8366, N8026);
and AND4 (N8382, N8378, N5829, N5613, N3452);
nor NOR2 (N8383, N8377, N3334);
or OR3 (N8384, N8370, N6413, N3394);
not NOT1 (N8385, N8380);
nand NAND2 (N8386, N8384, N2374);
not NOT1 (N8387, N8369);
nand NAND4 (N8388, N8361, N1683, N8021, N6259);
nand NAND4 (N8389, N8381, N7756, N1474, N2791);
and AND4 (N8390, N8382, N3607, N7986, N480);
buf BUF1 (N8391, N8390);
or OR3 (N8392, N8389, N2238, N188);
nor NOR3 (N8393, N8392, N7917, N8288);
nor NOR3 (N8394, N8393, N7776, N1370);
nand NAND3 (N8395, N8376, N8312, N3844);
not NOT1 (N8396, N8391);
nand NAND2 (N8397, N8386, N3590);
nor NOR2 (N8398, N8383, N717);
xor XOR2 (N8399, N8387, N5263);
and AND2 (N8400, N8385, N5019);
and AND4 (N8401, N8362, N3678, N7063, N2917);
or OR2 (N8402, N8401, N943);
not NOT1 (N8403, N8398);
xor XOR2 (N8404, N8395, N4879);
nand NAND4 (N8405, N8399, N3123, N3592, N6474);
xor XOR2 (N8406, N8396, N5513);
nand NAND4 (N8407, N8406, N277, N5309, N5308);
buf BUF1 (N8408, N8397);
xor XOR2 (N8409, N8408, N5434);
nand NAND2 (N8410, N8405, N1313);
or OR3 (N8411, N8407, N33, N8288);
nor NOR2 (N8412, N8409, N2924);
not NOT1 (N8413, N8368);
nand NAND4 (N8414, N8411, N439, N3261, N7467);
and AND3 (N8415, N8388, N1792, N1072);
nand NAND2 (N8416, N8400, N7600);
buf BUF1 (N8417, N8410);
nor NOR4 (N8418, N8417, N4486, N7335, N4536);
buf BUF1 (N8419, N8414);
nor NOR4 (N8420, N8415, N4900, N6729, N2244);
xor XOR2 (N8421, N8404, N2604);
and AND4 (N8422, N8412, N1856, N7150, N8206);
and AND4 (N8423, N8416, N7970, N6651, N6535);
nor NOR4 (N8424, N8413, N6343, N378, N187);
xor XOR2 (N8425, N8402, N2647);
and AND4 (N8426, N8423, N6365, N2127, N7308);
xor XOR2 (N8427, N8426, N8361);
nand NAND3 (N8428, N8422, N3174, N3485);
buf BUF1 (N8429, N8418);
nor NOR3 (N8430, N8425, N2515, N6926);
buf BUF1 (N8431, N8429);
and AND3 (N8432, N8427, N7151, N3835);
and AND4 (N8433, N8419, N1276, N2242, N326);
buf BUF1 (N8434, N8428);
xor XOR2 (N8435, N8403, N7124);
xor XOR2 (N8436, N8430, N4502);
nor NOR3 (N8437, N8433, N4058, N6956);
and AND3 (N8438, N8434, N2197, N938);
not NOT1 (N8439, N8431);
and AND2 (N8440, N8437, N1665);
nor NOR2 (N8441, N8394, N5931);
buf BUF1 (N8442, N8436);
nand NAND4 (N8443, N8420, N5812, N2689, N4284);
nand NAND2 (N8444, N8440, N2994);
nand NAND4 (N8445, N8442, N3273, N7084, N8326);
and AND3 (N8446, N8443, N938, N4085);
buf BUF1 (N8447, N8446);
nand NAND2 (N8448, N8439, N3041);
and AND4 (N8449, N8444, N2045, N3856, N6770);
buf BUF1 (N8450, N8445);
or OR3 (N8451, N8448, N770, N3485);
nand NAND2 (N8452, N8438, N3022);
nor NOR2 (N8453, N8447, N7651);
not NOT1 (N8454, N8424);
not NOT1 (N8455, N8450);
and AND3 (N8456, N8455, N1490, N5329);
or OR4 (N8457, N8441, N6717, N5372, N6822);
or OR3 (N8458, N8453, N755, N5259);
xor XOR2 (N8459, N8458, N7534);
buf BUF1 (N8460, N8435);
xor XOR2 (N8461, N8432, N5747);
and AND4 (N8462, N8452, N8435, N562, N8013);
nor NOR3 (N8463, N8456, N7084, N2781);
buf BUF1 (N8464, N8457);
and AND2 (N8465, N8449, N3636);
nor NOR4 (N8466, N8421, N4110, N2704, N7890);
not NOT1 (N8467, N8464);
nand NAND3 (N8468, N8459, N509, N990);
nor NOR3 (N8469, N8463, N7620, N642);
nand NAND2 (N8470, N8451, N5429);
nor NOR2 (N8471, N8469, N209);
buf BUF1 (N8472, N8460);
nand NAND2 (N8473, N8454, N5246);
nor NOR2 (N8474, N8462, N76);
buf BUF1 (N8475, N8461);
buf BUF1 (N8476, N8468);
nor NOR4 (N8477, N8473, N6333, N5, N1420);
or OR2 (N8478, N8477, N3097);
and AND2 (N8479, N8478, N1291);
and AND4 (N8480, N8465, N4712, N8040, N7549);
xor XOR2 (N8481, N8471, N1792);
not NOT1 (N8482, N8467);
or OR4 (N8483, N8475, N3312, N144, N813);
nor NOR2 (N8484, N8466, N4786);
buf BUF1 (N8485, N8481);
or OR2 (N8486, N8480, N368);
nor NOR3 (N8487, N8485, N1605, N5128);
nor NOR2 (N8488, N8470, N4786);
buf BUF1 (N8489, N8484);
xor XOR2 (N8490, N8489, N938);
not NOT1 (N8491, N8474);
buf BUF1 (N8492, N8491);
nor NOR3 (N8493, N8492, N2718, N6427);
buf BUF1 (N8494, N8487);
and AND2 (N8495, N8472, N2870);
xor XOR2 (N8496, N8476, N1760);
nand NAND2 (N8497, N8495, N7330);
xor XOR2 (N8498, N8483, N8473);
nor NOR4 (N8499, N8490, N6084, N3186, N6776);
and AND2 (N8500, N8494, N5161);
not NOT1 (N8501, N8493);
nand NAND4 (N8502, N8496, N6308, N1162, N7884);
nor NOR2 (N8503, N8498, N5175);
nor NOR4 (N8504, N8482, N7188, N3715, N5089);
and AND3 (N8505, N8502, N5878, N8246);
nor NOR2 (N8506, N8503, N4305);
or OR4 (N8507, N8504, N7631, N4399, N8148);
or OR3 (N8508, N8506, N6944, N4539);
xor XOR2 (N8509, N8505, N7892);
nand NAND2 (N8510, N8479, N3939);
nand NAND3 (N8511, N8508, N6377, N4756);
nand NAND2 (N8512, N8511, N2244);
xor XOR2 (N8513, N8512, N3615);
nand NAND3 (N8514, N8509, N5921, N5061);
nand NAND2 (N8515, N8510, N5308);
nand NAND2 (N8516, N8499, N8378);
nor NOR2 (N8517, N8514, N7284);
buf BUF1 (N8518, N8500);
not NOT1 (N8519, N8497);
nor NOR2 (N8520, N8518, N1184);
or OR4 (N8521, N8517, N5173, N6400, N3746);
not NOT1 (N8522, N8501);
buf BUF1 (N8523, N8516);
nor NOR2 (N8524, N8519, N4321);
nand NAND4 (N8525, N8523, N1834, N5099, N4596);
and AND3 (N8526, N8515, N3204, N1577);
not NOT1 (N8527, N8488);
nor NOR2 (N8528, N8526, N2302);
xor XOR2 (N8529, N8525, N2144);
nor NOR4 (N8530, N8520, N4047, N2561, N4941);
or OR3 (N8531, N8530, N3364, N2982);
buf BUF1 (N8532, N8531);
not NOT1 (N8533, N8527);
or OR4 (N8534, N8521, N7826, N3412, N4950);
not NOT1 (N8535, N8534);
nand NAND4 (N8536, N8533, N5292, N1075, N6365);
not NOT1 (N8537, N8532);
nand NAND2 (N8538, N8524, N4471);
or OR4 (N8539, N8536, N6196, N7774, N1444);
nand NAND3 (N8540, N8528, N6227, N148);
xor XOR2 (N8541, N8529, N7045);
or OR4 (N8542, N8540, N2016, N7824, N6220);
not NOT1 (N8543, N8542);
nor NOR3 (N8544, N8538, N3155, N2057);
xor XOR2 (N8545, N8513, N7008);
not NOT1 (N8546, N8522);
not NOT1 (N8547, N8539);
xor XOR2 (N8548, N8543, N4926);
buf BUF1 (N8549, N8486);
buf BUF1 (N8550, N8541);
not NOT1 (N8551, N8544);
nor NOR2 (N8552, N8551, N2945);
and AND3 (N8553, N8550, N5199, N2775);
nand NAND2 (N8554, N8537, N1920);
not NOT1 (N8555, N8546);
xor XOR2 (N8556, N8545, N6190);
nand NAND2 (N8557, N8507, N4967);
or OR2 (N8558, N8555, N2297);
buf BUF1 (N8559, N8554);
xor XOR2 (N8560, N8558, N3584);
and AND3 (N8561, N8552, N4702, N61);
nand NAND4 (N8562, N8561, N1943, N7149, N5240);
nor NOR4 (N8563, N8549, N390, N1822, N6926);
nand NAND4 (N8564, N8563, N6843, N2859, N3275);
buf BUF1 (N8565, N8564);
or OR2 (N8566, N8557, N5432);
and AND2 (N8567, N8560, N1439);
buf BUF1 (N8568, N8559);
and AND4 (N8569, N8535, N2058, N4089, N2782);
nor NOR3 (N8570, N8565, N5036, N8444);
nand NAND4 (N8571, N8547, N1726, N1476, N4392);
not NOT1 (N8572, N8562);
nand NAND4 (N8573, N8556, N6720, N2920, N721);
buf BUF1 (N8574, N8571);
and AND3 (N8575, N8573, N4874, N4290);
buf BUF1 (N8576, N8569);
or OR4 (N8577, N8574, N2289, N4190, N2712);
nand NAND3 (N8578, N8548, N4465, N2198);
or OR3 (N8579, N8576, N5851, N3375);
buf BUF1 (N8580, N8570);
nor NOR3 (N8581, N8580, N2147, N5734);
xor XOR2 (N8582, N8579, N8034);
not NOT1 (N8583, N8582);
or OR3 (N8584, N8567, N4521, N2922);
buf BUF1 (N8585, N8581);
nand NAND2 (N8586, N8575, N4123);
and AND3 (N8587, N8577, N5786, N7445);
nor NOR3 (N8588, N8566, N2650, N4730);
and AND3 (N8589, N8586, N1195, N5100);
buf BUF1 (N8590, N8584);
nand NAND4 (N8591, N8590, N5086, N391, N6738);
nor NOR3 (N8592, N8585, N2674, N5302);
nor NOR2 (N8593, N8578, N2577);
buf BUF1 (N8594, N8588);
buf BUF1 (N8595, N8583);
or OR4 (N8596, N8589, N1399, N7072, N608);
not NOT1 (N8597, N8587);
not NOT1 (N8598, N8553);
buf BUF1 (N8599, N8572);
buf BUF1 (N8600, N8596);
buf BUF1 (N8601, N8597);
or OR2 (N8602, N8593, N6082);
or OR4 (N8603, N8592, N8237, N2014, N1155);
or OR2 (N8604, N8600, N3755);
and AND3 (N8605, N8595, N6345, N437);
not NOT1 (N8606, N8591);
xor XOR2 (N8607, N8568, N3349);
nand NAND3 (N8608, N8599, N8039, N3157);
or OR2 (N8609, N8603, N6932);
and AND2 (N8610, N8598, N624);
nor NOR2 (N8611, N8594, N4592);
nand NAND4 (N8612, N8605, N8514, N560, N320);
or OR3 (N8613, N8611, N2546, N1757);
not NOT1 (N8614, N8606);
or OR3 (N8615, N8614, N7169, N427);
nor NOR3 (N8616, N8602, N6683, N4748);
buf BUF1 (N8617, N8601);
or OR2 (N8618, N8604, N695);
xor XOR2 (N8619, N8618, N6233);
buf BUF1 (N8620, N8609);
xor XOR2 (N8621, N8613, N5903);
and AND4 (N8622, N8610, N6310, N1595, N8153);
nand NAND4 (N8623, N8619, N1934, N533, N2383);
xor XOR2 (N8624, N8617, N8524);
xor XOR2 (N8625, N8616, N583);
nand NAND4 (N8626, N8615, N2255, N2828, N3610);
not NOT1 (N8627, N8608);
and AND3 (N8628, N8624, N4932, N6206);
buf BUF1 (N8629, N8623);
and AND2 (N8630, N8621, N338);
not NOT1 (N8631, N8629);
xor XOR2 (N8632, N8612, N2752);
buf BUF1 (N8633, N8632);
not NOT1 (N8634, N8633);
nor NOR3 (N8635, N8627, N5245, N1505);
not NOT1 (N8636, N8620);
xor XOR2 (N8637, N8622, N4716);
and AND2 (N8638, N8636, N4304);
and AND4 (N8639, N8625, N2916, N3685, N6513);
and AND2 (N8640, N8631, N764);
nand NAND2 (N8641, N8630, N3978);
nand NAND4 (N8642, N8637, N3941, N7237, N3782);
or OR2 (N8643, N8626, N6595);
xor XOR2 (N8644, N8639, N8244);
or OR2 (N8645, N8638, N1862);
xor XOR2 (N8646, N8634, N5544);
nor NOR2 (N8647, N8642, N3633);
buf BUF1 (N8648, N8643);
nor NOR2 (N8649, N8645, N5465);
not NOT1 (N8650, N8644);
not NOT1 (N8651, N8650);
xor XOR2 (N8652, N8641, N7408);
nor NOR3 (N8653, N8651, N3521, N4576);
or OR3 (N8654, N8628, N4059, N8574);
nor NOR4 (N8655, N8607, N1380, N2554, N64);
buf BUF1 (N8656, N8635);
not NOT1 (N8657, N8648);
nor NOR4 (N8658, N8656, N5283, N6093, N220);
not NOT1 (N8659, N8655);
or OR2 (N8660, N8652, N2838);
xor XOR2 (N8661, N8660, N186);
nand NAND3 (N8662, N8658, N2964, N4715);
not NOT1 (N8663, N8640);
nand NAND2 (N8664, N8646, N2656);
and AND3 (N8665, N8653, N6720, N2858);
buf BUF1 (N8666, N8662);
or OR4 (N8667, N8666, N1117, N8417, N292);
and AND3 (N8668, N8659, N7908, N4243);
xor XOR2 (N8669, N8657, N8077);
not NOT1 (N8670, N8664);
buf BUF1 (N8671, N8667);
nor NOR2 (N8672, N8668, N2852);
nor NOR3 (N8673, N8663, N7625, N8033);
buf BUF1 (N8674, N8654);
or OR2 (N8675, N8661, N6691);
buf BUF1 (N8676, N8670);
nor NOR2 (N8677, N8665, N2584);
and AND3 (N8678, N8672, N1369, N7305);
nand NAND3 (N8679, N8649, N4415, N6910);
xor XOR2 (N8680, N8669, N3427);
not NOT1 (N8681, N8673);
xor XOR2 (N8682, N8671, N4144);
buf BUF1 (N8683, N8674);
nand NAND2 (N8684, N8679, N8266);
nor NOR2 (N8685, N8680, N4890);
not NOT1 (N8686, N8647);
or OR4 (N8687, N8685, N3108, N6262, N1729);
or OR3 (N8688, N8676, N393, N5759);
nand NAND4 (N8689, N8684, N3031, N4878, N6857);
nand NAND4 (N8690, N8681, N1874, N1710, N7056);
not NOT1 (N8691, N8687);
buf BUF1 (N8692, N8690);
not NOT1 (N8693, N8691);
nand NAND3 (N8694, N8692, N860, N3596);
nand NAND4 (N8695, N8688, N7547, N784, N6323);
nor NOR3 (N8696, N8689, N8396, N6812);
xor XOR2 (N8697, N8695, N2663);
nand NAND3 (N8698, N8697, N1253, N6925);
buf BUF1 (N8699, N8675);
buf BUF1 (N8700, N8696);
or OR3 (N8701, N8700, N1070, N1886);
nor NOR2 (N8702, N8694, N7333);
not NOT1 (N8703, N8701);
not NOT1 (N8704, N8686);
or OR2 (N8705, N8677, N5695);
not NOT1 (N8706, N8682);
nor NOR2 (N8707, N8705, N4433);
nor NOR2 (N8708, N8698, N1580);
nand NAND4 (N8709, N8706, N4595, N820, N7347);
and AND2 (N8710, N8678, N2075);
nand NAND3 (N8711, N8683, N6559, N2466);
nand NAND4 (N8712, N8709, N3213, N613, N1695);
nor NOR4 (N8713, N8693, N3870, N5595, N2944);
and AND3 (N8714, N8702, N3614, N3621);
not NOT1 (N8715, N8710);
buf BUF1 (N8716, N8714);
nand NAND4 (N8717, N8712, N489, N7455, N4775);
and AND4 (N8718, N8708, N5410, N2457, N2360);
buf BUF1 (N8719, N8699);
nor NOR2 (N8720, N8715, N1005);
not NOT1 (N8721, N8719);
nand NAND2 (N8722, N8711, N7790);
nor NOR2 (N8723, N8721, N4325);
buf BUF1 (N8724, N8713);
or OR3 (N8725, N8720, N1302, N4690);
or OR3 (N8726, N8704, N11, N3898);
or OR3 (N8727, N8726, N6276, N5578);
not NOT1 (N8728, N8703);
buf BUF1 (N8729, N8707);
or OR4 (N8730, N8722, N6688, N5993, N7111);
or OR2 (N8731, N8730, N4098);
nand NAND3 (N8732, N8723, N1748, N1648);
buf BUF1 (N8733, N8716);
xor XOR2 (N8734, N8733, N1194);
nor NOR4 (N8735, N8724, N739, N5793, N5619);
not NOT1 (N8736, N8735);
xor XOR2 (N8737, N8728, N566);
xor XOR2 (N8738, N8737, N4025);
nor NOR2 (N8739, N8738, N1825);
xor XOR2 (N8740, N8732, N4584);
not NOT1 (N8741, N8725);
buf BUF1 (N8742, N8740);
xor XOR2 (N8743, N8742, N8301);
buf BUF1 (N8744, N8718);
xor XOR2 (N8745, N8741, N3308);
nor NOR2 (N8746, N8731, N6267);
not NOT1 (N8747, N8744);
and AND3 (N8748, N8727, N4341, N4718);
nand NAND2 (N8749, N8729, N5805);
nor NOR3 (N8750, N8747, N3179, N638);
not NOT1 (N8751, N8750);
and AND2 (N8752, N8748, N2962);
and AND3 (N8753, N8743, N5043, N3257);
nor NOR4 (N8754, N8739, N2226, N2717, N3251);
not NOT1 (N8755, N8734);
and AND4 (N8756, N8745, N5936, N3639, N477);
nor NOR2 (N8757, N8755, N2186);
not NOT1 (N8758, N8753);
or OR3 (N8759, N8749, N6815, N2941);
nor NOR4 (N8760, N8751, N2370, N458, N7816);
or OR3 (N8761, N8752, N2548, N4349);
and AND3 (N8762, N8761, N1770, N2915);
xor XOR2 (N8763, N8736, N7062);
or OR3 (N8764, N8757, N8155, N8318);
buf BUF1 (N8765, N8764);
not NOT1 (N8766, N8754);
xor XOR2 (N8767, N8756, N4986);
buf BUF1 (N8768, N8766);
and AND2 (N8769, N8763, N7970);
nand NAND3 (N8770, N8762, N7444, N8178);
nor NOR3 (N8771, N8769, N5307, N4640);
or OR2 (N8772, N8770, N1689);
nand NAND2 (N8773, N8760, N3553);
or OR2 (N8774, N8758, N2040);
or OR3 (N8775, N8759, N794, N4103);
and AND4 (N8776, N8746, N8411, N5909, N99);
not NOT1 (N8777, N8773);
buf BUF1 (N8778, N8767);
and AND3 (N8779, N8778, N3968, N1356);
nand NAND4 (N8780, N8777, N8025, N4456, N3558);
nand NAND4 (N8781, N8765, N572, N7512, N1940);
xor XOR2 (N8782, N8776, N5119);
xor XOR2 (N8783, N8780, N3725);
nor NOR4 (N8784, N8782, N6114, N7496, N1823);
or OR2 (N8785, N8768, N7840);
xor XOR2 (N8786, N8771, N1954);
xor XOR2 (N8787, N8774, N7282);
not NOT1 (N8788, N8785);
and AND4 (N8789, N8787, N2959, N1005, N7418);
and AND4 (N8790, N8788, N4386, N5666, N327);
not NOT1 (N8791, N8790);
not NOT1 (N8792, N8779);
nor NOR4 (N8793, N8783, N8116, N2192, N2446);
xor XOR2 (N8794, N8784, N5084);
buf BUF1 (N8795, N8793);
xor XOR2 (N8796, N8795, N321);
and AND2 (N8797, N8789, N1645);
nor NOR2 (N8798, N8794, N2757);
or OR3 (N8799, N8798, N2138, N8420);
not NOT1 (N8800, N8796);
nor NOR4 (N8801, N8797, N5935, N5825, N5602);
and AND3 (N8802, N8791, N6786, N7905);
or OR2 (N8803, N8781, N1649);
nand NAND3 (N8804, N8717, N8070, N644);
buf BUF1 (N8805, N8792);
nor NOR3 (N8806, N8775, N2676, N6694);
buf BUF1 (N8807, N8772);
or OR4 (N8808, N8800, N67, N7038, N1084);
or OR4 (N8809, N8802, N8770, N3319, N6728);
xor XOR2 (N8810, N8803, N3294);
nor NOR4 (N8811, N8786, N8319, N3961, N3865);
nor NOR3 (N8812, N8806, N4205, N1040);
buf BUF1 (N8813, N8811);
and AND2 (N8814, N8805, N2030);
not NOT1 (N8815, N8814);
or OR3 (N8816, N8813, N5146, N5969);
xor XOR2 (N8817, N8810, N4596);
buf BUF1 (N8818, N8801);
or OR2 (N8819, N8807, N4197);
not NOT1 (N8820, N8808);
or OR4 (N8821, N8812, N1759, N7402, N8345);
not NOT1 (N8822, N8809);
buf BUF1 (N8823, N8819);
xor XOR2 (N8824, N8816, N238);
nand NAND3 (N8825, N8824, N3000, N5294);
or OR2 (N8826, N8818, N3464);
nand NAND2 (N8827, N8826, N2173);
or OR3 (N8828, N8822, N5231, N5026);
nor NOR4 (N8829, N8804, N6304, N4537, N4552);
and AND3 (N8830, N8820, N688, N4785);
buf BUF1 (N8831, N8825);
nand NAND2 (N8832, N8799, N3107);
and AND4 (N8833, N8815, N797, N4001, N814);
or OR4 (N8834, N8821, N1484, N7707, N1846);
xor XOR2 (N8835, N8828, N7120);
nand NAND2 (N8836, N8831, N3875);
buf BUF1 (N8837, N8835);
buf BUF1 (N8838, N8817);
buf BUF1 (N8839, N8823);
or OR3 (N8840, N8839, N7192, N665);
xor XOR2 (N8841, N8838, N992);
nor NOR2 (N8842, N8833, N8509);
not NOT1 (N8843, N8836);
xor XOR2 (N8844, N8832, N7508);
xor XOR2 (N8845, N8841, N2653);
nand NAND4 (N8846, N8834, N289, N620, N6405);
nand NAND2 (N8847, N8840, N7112);
and AND2 (N8848, N8844, N8525);
nor NOR2 (N8849, N8827, N5713);
nand NAND3 (N8850, N8842, N6571, N4224);
or OR2 (N8851, N8846, N7099);
and AND3 (N8852, N8849, N1330, N2791);
buf BUF1 (N8853, N8851);
not NOT1 (N8854, N8829);
xor XOR2 (N8855, N8852, N6749);
and AND4 (N8856, N8850, N7755, N7900, N616);
and AND2 (N8857, N8837, N6919);
and AND4 (N8858, N8845, N7710, N3924, N7793);
not NOT1 (N8859, N8853);
not NOT1 (N8860, N8855);
xor XOR2 (N8861, N8857, N4784);
nand NAND4 (N8862, N8848, N1469, N7670, N4478);
nor NOR3 (N8863, N8860, N7273, N8410);
nor NOR4 (N8864, N8830, N775, N6126, N2777);
nor NOR3 (N8865, N8859, N8611, N2566);
not NOT1 (N8866, N8843);
or OR2 (N8867, N8866, N441);
nor NOR2 (N8868, N8861, N5313);
buf BUF1 (N8869, N8863);
or OR4 (N8870, N8864, N5219, N6345, N7400);
or OR4 (N8871, N8868, N6324, N174, N5881);
buf BUF1 (N8872, N8854);
buf BUF1 (N8873, N8871);
nand NAND4 (N8874, N8858, N3757, N991, N1998);
buf BUF1 (N8875, N8872);
nand NAND3 (N8876, N8862, N8635, N2118);
and AND3 (N8877, N8873, N873, N2142);
xor XOR2 (N8878, N8867, N2230);
buf BUF1 (N8879, N8847);
and AND3 (N8880, N8879, N8661, N1131);
xor XOR2 (N8881, N8880, N4302);
xor XOR2 (N8882, N8877, N5096);
xor XOR2 (N8883, N8870, N359);
xor XOR2 (N8884, N8882, N4038);
nand NAND3 (N8885, N8881, N6076, N8125);
xor XOR2 (N8886, N8878, N443);
buf BUF1 (N8887, N8875);
xor XOR2 (N8888, N8869, N3493);
not NOT1 (N8889, N8865);
nand NAND3 (N8890, N8856, N3887, N7483);
nand NAND2 (N8891, N8874, N5472);
not NOT1 (N8892, N8884);
nor NOR3 (N8893, N8891, N6077, N2972);
xor XOR2 (N8894, N8892, N7449);
xor XOR2 (N8895, N8876, N237);
nor NOR4 (N8896, N8895, N5552, N5408, N7220);
and AND4 (N8897, N8893, N3486, N3243, N6401);
nor NOR3 (N8898, N8887, N117, N5985);
nand NAND4 (N8899, N8897, N3275, N4738, N491);
not NOT1 (N8900, N8896);
nor NOR3 (N8901, N8886, N4834, N3261);
and AND2 (N8902, N8883, N1642);
or OR4 (N8903, N8894, N6638, N2319, N2558);
or OR4 (N8904, N8889, N5720, N4406, N8492);
or OR3 (N8905, N8898, N2144, N819);
or OR3 (N8906, N8905, N3368, N2418);
and AND2 (N8907, N8890, N917);
xor XOR2 (N8908, N8885, N4915);
or OR2 (N8909, N8907, N492);
nor NOR3 (N8910, N8899, N1727, N1459);
nand NAND4 (N8911, N8910, N8285, N7238, N4886);
and AND3 (N8912, N8909, N7178, N8811);
buf BUF1 (N8913, N8901);
nand NAND4 (N8914, N8903, N4686, N2928, N2976);
and AND2 (N8915, N8913, N6407);
buf BUF1 (N8916, N8902);
nand NAND3 (N8917, N8914, N3957, N654);
nor NOR4 (N8918, N8915, N4198, N4335, N7671);
nand NAND3 (N8919, N8904, N4226, N7163);
not NOT1 (N8920, N8912);
nand NAND3 (N8921, N8900, N1316, N4385);
buf BUF1 (N8922, N8906);
or OR4 (N8923, N8922, N6001, N4767, N2907);
nor NOR3 (N8924, N8918, N8045, N6573);
nor NOR4 (N8925, N8911, N5949, N6834, N3197);
or OR3 (N8926, N8921, N2156, N7508);
nor NOR3 (N8927, N8924, N8221, N1254);
or OR3 (N8928, N8926, N4598, N3516);
xor XOR2 (N8929, N8919, N8780);
nor NOR2 (N8930, N8928, N266);
not NOT1 (N8931, N8929);
xor XOR2 (N8932, N8917, N3784);
or OR3 (N8933, N8920, N4999, N3094);
nand NAND2 (N8934, N8908, N1315);
and AND4 (N8935, N8930, N7558, N5370, N4742);
not NOT1 (N8936, N8932);
nand NAND4 (N8937, N8934, N8805, N7255, N1038);
or OR3 (N8938, N8933, N5089, N2431);
and AND2 (N8939, N8888, N6301);
and AND4 (N8940, N8937, N7185, N3478, N4973);
buf BUF1 (N8941, N8936);
buf BUF1 (N8942, N8923);
not NOT1 (N8943, N8942);
xor XOR2 (N8944, N8931, N7277);
xor XOR2 (N8945, N8935, N4720);
and AND3 (N8946, N8941, N3432, N3924);
nand NAND3 (N8947, N8916, N8344, N7129);
buf BUF1 (N8948, N8943);
nor NOR3 (N8949, N8945, N7650, N2070);
nor NOR4 (N8950, N8944, N5954, N2158, N1850);
not NOT1 (N8951, N8946);
and AND4 (N8952, N8940, N8586, N7085, N3320);
and AND2 (N8953, N8948, N8634);
or OR2 (N8954, N8947, N4790);
or OR2 (N8955, N8949, N5779);
buf BUF1 (N8956, N8952);
nor NOR3 (N8957, N8954, N7001, N4095);
not NOT1 (N8958, N8957);
nand NAND3 (N8959, N8925, N8452, N8790);
and AND4 (N8960, N8938, N2296, N1875, N6817);
nand NAND3 (N8961, N8955, N463, N3881);
buf BUF1 (N8962, N8956);
xor XOR2 (N8963, N8950, N2424);
and AND3 (N8964, N8953, N1866, N2630);
nand NAND3 (N8965, N8951, N5808, N7480);
nand NAND3 (N8966, N8961, N4444, N5312);
buf BUF1 (N8967, N8927);
nand NAND3 (N8968, N8963, N1766, N4632);
nand NAND2 (N8969, N8939, N5396);
nor NOR4 (N8970, N8967, N25, N5547, N6764);
and AND3 (N8971, N8965, N675, N803);
and AND2 (N8972, N8966, N2626);
nor NOR3 (N8973, N8969, N5059, N1042);
nor NOR2 (N8974, N8972, N1992);
and AND2 (N8975, N8968, N6206);
not NOT1 (N8976, N8974);
buf BUF1 (N8977, N8962);
and AND4 (N8978, N8959, N4239, N4851, N4381);
nor NOR3 (N8979, N8975, N8507, N6210);
buf BUF1 (N8980, N8976);
and AND3 (N8981, N8958, N5475, N4748);
xor XOR2 (N8982, N8970, N7931);
or OR4 (N8983, N8978, N775, N5278, N6586);
or OR3 (N8984, N8960, N8408, N5781);
nand NAND2 (N8985, N8981, N1952);
xor XOR2 (N8986, N8973, N4206);
nor NOR3 (N8987, N8971, N7337, N1958);
or OR3 (N8988, N8987, N7728, N2894);
or OR2 (N8989, N8985, N4099);
xor XOR2 (N8990, N8984, N1367);
and AND4 (N8991, N8986, N8077, N765, N6975);
xor XOR2 (N8992, N8964, N6454);
or OR4 (N8993, N8977, N6507, N4874, N2104);
not NOT1 (N8994, N8993);
not NOT1 (N8995, N8983);
not NOT1 (N8996, N8979);
or OR3 (N8997, N8995, N4738, N4135);
or OR3 (N8998, N8992, N8346, N3482);
xor XOR2 (N8999, N8994, N5035);
not NOT1 (N9000, N8980);
xor XOR2 (N9001, N8998, N4957);
not NOT1 (N9002, N8991);
buf BUF1 (N9003, N8982);
not NOT1 (N9004, N8988);
nand NAND4 (N9005, N9002, N8253, N4677, N5258);
and AND3 (N9006, N8990, N2892, N2358);
and AND2 (N9007, N9005, N4414);
nand NAND4 (N9008, N9000, N1967, N5684, N5884);
or OR4 (N9009, N9001, N4210, N4283, N4862);
buf BUF1 (N9010, N9006);
not NOT1 (N9011, N9010);
xor XOR2 (N9012, N8996, N3962);
or OR3 (N9013, N9003, N8342, N8739);
nand NAND4 (N9014, N9008, N3334, N1707, N2017);
not NOT1 (N9015, N9011);
or OR4 (N9016, N9013, N4489, N5025, N5735);
or OR4 (N9017, N8989, N8276, N1148, N1853);
and AND2 (N9018, N9016, N4960);
or OR2 (N9019, N9009, N1655);
xor XOR2 (N9020, N9004, N6011);
buf BUF1 (N9021, N9012);
nand NAND3 (N9022, N8997, N6784, N2061);
nor NOR3 (N9023, N9022, N315, N7828);
and AND3 (N9024, N9020, N290, N4511);
and AND3 (N9025, N9021, N7341, N7050);
nor NOR2 (N9026, N9007, N7528);
or OR2 (N9027, N8999, N528);
or OR3 (N9028, N9015, N1903, N6185);
and AND3 (N9029, N9018, N2873, N8861);
buf BUF1 (N9030, N9019);
nor NOR3 (N9031, N9027, N6325, N7684);
buf BUF1 (N9032, N9029);
nand NAND2 (N9033, N9014, N1843);
xor XOR2 (N9034, N9025, N3956);
buf BUF1 (N9035, N9030);
nand NAND2 (N9036, N9023, N8048);
not NOT1 (N9037, N9024);
not NOT1 (N9038, N9034);
nand NAND2 (N9039, N9036, N2131);
or OR3 (N9040, N9038, N2187, N2297);
and AND2 (N9041, N9033, N486);
xor XOR2 (N9042, N9037, N8445);
xor XOR2 (N9043, N9039, N6782);
nand NAND2 (N9044, N9041, N6394);
nor NOR4 (N9045, N9043, N6826, N1916, N5050);
buf BUF1 (N9046, N9040);
buf BUF1 (N9047, N9032);
not NOT1 (N9048, N9031);
or OR4 (N9049, N9047, N1564, N1624, N727);
and AND2 (N9050, N9042, N2628);
and AND3 (N9051, N9017, N4696, N1823);
nand NAND4 (N9052, N9028, N4591, N3468, N8899);
nand NAND3 (N9053, N9035, N8745, N9022);
not NOT1 (N9054, N9026);
xor XOR2 (N9055, N9045, N8149);
or OR4 (N9056, N9053, N3212, N6098, N4109);
nand NAND4 (N9057, N9056, N3168, N2560, N7241);
buf BUF1 (N9058, N9054);
or OR4 (N9059, N9046, N3419, N7376, N4445);
not NOT1 (N9060, N9059);
and AND2 (N9061, N9049, N2186);
nand NAND3 (N9062, N9057, N3725, N3578);
nor NOR4 (N9063, N9062, N551, N3750, N1969);
xor XOR2 (N9064, N9063, N5269);
not NOT1 (N9065, N9060);
nand NAND3 (N9066, N9061, N8867, N3092);
or OR2 (N9067, N9051, N4553);
nand NAND2 (N9068, N9066, N7801);
nand NAND2 (N9069, N9068, N6989);
xor XOR2 (N9070, N9052, N421);
not NOT1 (N9071, N9067);
not NOT1 (N9072, N9048);
or OR3 (N9073, N9071, N6179, N1081);
nor NOR4 (N9074, N9073, N2874, N2951, N6418);
not NOT1 (N9075, N9044);
nand NAND4 (N9076, N9055, N8001, N2831, N1914);
nor NOR4 (N9077, N9065, N6046, N548, N6055);
or OR3 (N9078, N9064, N3325, N6533);
buf BUF1 (N9079, N9072);
and AND2 (N9080, N9070, N5763);
nand NAND3 (N9081, N9079, N2362, N5148);
buf BUF1 (N9082, N9069);
xor XOR2 (N9083, N9050, N1572);
nand NAND2 (N9084, N9074, N4972);
xor XOR2 (N9085, N9083, N7627);
xor XOR2 (N9086, N9075, N3614);
nand NAND2 (N9087, N9084, N6665);
nand NAND2 (N9088, N9085, N2180);
buf BUF1 (N9089, N9077);
buf BUF1 (N9090, N9088);
not NOT1 (N9091, N9082);
buf BUF1 (N9092, N9090);
and AND2 (N9093, N9086, N8177);
nor NOR2 (N9094, N9087, N1359);
nor NOR4 (N9095, N9080, N59, N4235, N2576);
not NOT1 (N9096, N9094);
nand NAND3 (N9097, N9095, N4755, N5246);
not NOT1 (N9098, N9089);
xor XOR2 (N9099, N9097, N6729);
not NOT1 (N9100, N9078);
not NOT1 (N9101, N9099);
xor XOR2 (N9102, N9100, N6023);
xor XOR2 (N9103, N9091, N818);
nor NOR2 (N9104, N9081, N1811);
or OR4 (N9105, N9093, N7778, N7560, N7415);
or OR3 (N9106, N9103, N8064, N189);
nor NOR2 (N9107, N9105, N52);
xor XOR2 (N9108, N9092, N4035);
and AND3 (N9109, N9058, N7369, N8271);
not NOT1 (N9110, N9076);
not NOT1 (N9111, N9098);
buf BUF1 (N9112, N9108);
nand NAND4 (N9113, N9106, N4203, N6562, N851);
not NOT1 (N9114, N9096);
nand NAND4 (N9115, N9109, N1429, N8307, N2769);
nand NAND4 (N9116, N9114, N4293, N227, N182);
and AND2 (N9117, N9112, N1134);
buf BUF1 (N9118, N9101);
or OR2 (N9119, N9116, N1517);
nand NAND2 (N9120, N9118, N3377);
or OR2 (N9121, N9102, N7949);
xor XOR2 (N9122, N9107, N4010);
and AND2 (N9123, N9120, N7180);
and AND2 (N9124, N9119, N7243);
nand NAND2 (N9125, N9122, N2098);
or OR4 (N9126, N9115, N4803, N3807, N2700);
and AND4 (N9127, N9126, N8446, N6936, N2143);
nand NAND2 (N9128, N9110, N8182);
xor XOR2 (N9129, N9117, N103);
or OR3 (N9130, N9111, N7585, N1939);
xor XOR2 (N9131, N9113, N5237);
buf BUF1 (N9132, N9121);
nand NAND3 (N9133, N9128, N3046, N7872);
and AND2 (N9134, N9104, N929);
not NOT1 (N9135, N9123);
or OR3 (N9136, N9133, N5209, N5935);
nand NAND4 (N9137, N9131, N5840, N3315, N8569);
and AND3 (N9138, N9137, N2077, N7551);
buf BUF1 (N9139, N9129);
buf BUF1 (N9140, N9134);
or OR4 (N9141, N9135, N2053, N7914, N1244);
nand NAND4 (N9142, N9140, N2644, N3562, N189);
nand NAND4 (N9143, N9139, N6782, N6989, N7090);
xor XOR2 (N9144, N9141, N895);
and AND3 (N9145, N9125, N5226, N7517);
xor XOR2 (N9146, N9138, N6750);
nand NAND2 (N9147, N9132, N5634);
and AND2 (N9148, N9147, N7580);
nand NAND3 (N9149, N9144, N1352, N3082);
nor NOR4 (N9150, N9145, N6147, N6320, N7971);
or OR4 (N9151, N9142, N1458, N7824, N8169);
xor XOR2 (N9152, N9127, N4201);
buf BUF1 (N9153, N9146);
or OR3 (N9154, N9130, N5987, N4403);
and AND4 (N9155, N9151, N1901, N6300, N6020);
nor NOR3 (N9156, N9149, N9109, N4636);
or OR2 (N9157, N9150, N3452);
and AND4 (N9158, N9154, N1983, N4602, N8051);
or OR4 (N9159, N9158, N7573, N7994, N7824);
nor NOR4 (N9160, N9136, N3980, N6022, N7141);
nor NOR3 (N9161, N9159, N2604, N8776);
and AND2 (N9162, N9148, N4570);
xor XOR2 (N9163, N9155, N9136);
nand NAND2 (N9164, N9160, N4139);
not NOT1 (N9165, N9153);
nor NOR2 (N9166, N9164, N6210);
xor XOR2 (N9167, N9165, N8896);
buf BUF1 (N9168, N9163);
nor NOR4 (N9169, N9143, N7007, N1756, N6989);
or OR2 (N9170, N9169, N2921);
not NOT1 (N9171, N9166);
or OR4 (N9172, N9161, N5252, N459, N6984);
or OR3 (N9173, N9152, N8378, N9064);
not NOT1 (N9174, N9173);
or OR3 (N9175, N9168, N6371, N3757);
or OR3 (N9176, N9156, N7403, N7494);
nand NAND2 (N9177, N9175, N3757);
buf BUF1 (N9178, N9172);
and AND4 (N9179, N9167, N1543, N8636, N2670);
not NOT1 (N9180, N9171);
nand NAND4 (N9181, N9174, N2965, N3753, N6986);
and AND4 (N9182, N9157, N7828, N5300, N6433);
or OR3 (N9183, N9176, N2392, N8305);
not NOT1 (N9184, N9181);
buf BUF1 (N9185, N9170);
or OR2 (N9186, N9179, N8674);
not NOT1 (N9187, N9186);
nand NAND4 (N9188, N9124, N6639, N6165, N719);
or OR3 (N9189, N9182, N8258, N8236);
nand NAND2 (N9190, N9177, N7903);
nor NOR4 (N9191, N9184, N8603, N3066, N4564);
buf BUF1 (N9192, N9189);
xor XOR2 (N9193, N9178, N6383);
nor NOR2 (N9194, N9180, N3809);
and AND4 (N9195, N9190, N7550, N7179, N5862);
nand NAND3 (N9196, N9185, N3145, N1500);
and AND4 (N9197, N9162, N4504, N42, N8965);
xor XOR2 (N9198, N9193, N5803);
xor XOR2 (N9199, N9197, N8207);
buf BUF1 (N9200, N9187);
nor NOR3 (N9201, N9195, N7813, N2046);
nand NAND2 (N9202, N9192, N7274);
xor XOR2 (N9203, N9188, N1739);
nor NOR2 (N9204, N9191, N3102);
and AND4 (N9205, N9202, N2654, N9147, N1874);
xor XOR2 (N9206, N9194, N3845);
buf BUF1 (N9207, N9183);
buf BUF1 (N9208, N9201);
or OR3 (N9209, N9203, N2538, N2377);
nor NOR4 (N9210, N9199, N8921, N6809, N4316);
not NOT1 (N9211, N9198);
and AND3 (N9212, N9209, N1253, N7925);
nor NOR4 (N9213, N9196, N1904, N3867, N8541);
not NOT1 (N9214, N9212);
and AND4 (N9215, N9204, N2036, N2281, N8970);
nand NAND4 (N9216, N9207, N5948, N7448, N1582);
and AND3 (N9217, N9213, N4425, N4865);
or OR3 (N9218, N9200, N4745, N3829);
buf BUF1 (N9219, N9217);
or OR4 (N9220, N9218, N1807, N7887, N6967);
buf BUF1 (N9221, N9211);
nand NAND2 (N9222, N9215, N8835);
nor NOR2 (N9223, N9221, N6235);
nand NAND2 (N9224, N9205, N2429);
nand NAND2 (N9225, N9210, N3494);
xor XOR2 (N9226, N9223, N2805);
nand NAND4 (N9227, N9225, N6921, N7689, N2579);
buf BUF1 (N9228, N9214);
nor NOR2 (N9229, N9224, N5704);
buf BUF1 (N9230, N9219);
not NOT1 (N9231, N9222);
buf BUF1 (N9232, N9206);
and AND4 (N9233, N9208, N5275, N3025, N4017);
or OR3 (N9234, N9220, N5356, N6007);
or OR2 (N9235, N9229, N5965);
nor NOR3 (N9236, N9235, N5955, N8175);
and AND4 (N9237, N9232, N3478, N4949, N52);
xor XOR2 (N9238, N9226, N1184);
or OR2 (N9239, N9236, N2920);
not NOT1 (N9240, N9238);
nor NOR3 (N9241, N9234, N1842, N1723);
nor NOR2 (N9242, N9227, N6248);
nor NOR3 (N9243, N9228, N2740, N8903);
not NOT1 (N9244, N9216);
nor NOR4 (N9245, N9230, N7217, N44, N3116);
nor NOR2 (N9246, N9239, N8945);
nor NOR4 (N9247, N9240, N295, N7749, N6232);
not NOT1 (N9248, N9237);
or OR2 (N9249, N9233, N4271);
nand NAND2 (N9250, N9241, N2260);
nor NOR4 (N9251, N9248, N6104, N963, N1041);
and AND3 (N9252, N9242, N2360, N7753);
nor NOR3 (N9253, N9251, N3458, N7388);
nand NAND3 (N9254, N9245, N9233, N1751);
and AND3 (N9255, N9249, N1883, N6687);
buf BUF1 (N9256, N9250);
not NOT1 (N9257, N9252);
nand NAND2 (N9258, N9231, N6576);
or OR2 (N9259, N9246, N3863);
nand NAND2 (N9260, N9243, N8940);
or OR4 (N9261, N9256, N535, N2544, N2511);
buf BUF1 (N9262, N9253);
buf BUF1 (N9263, N9259);
and AND4 (N9264, N9255, N4426, N8574, N8363);
or OR4 (N9265, N9254, N7047, N8374, N5951);
buf BUF1 (N9266, N9262);
xor XOR2 (N9267, N9266, N2305);
and AND4 (N9268, N9244, N4108, N9176, N7655);
or OR3 (N9269, N9260, N7712, N8862);
xor XOR2 (N9270, N9264, N5723);
buf BUF1 (N9271, N9257);
or OR3 (N9272, N9270, N7335, N846);
nand NAND3 (N9273, N9247, N5466, N4520);
buf BUF1 (N9274, N9269);
or OR3 (N9275, N9261, N8425, N3569);
nand NAND2 (N9276, N9268, N7836);
or OR3 (N9277, N9273, N7589, N2610);
not NOT1 (N9278, N9265);
buf BUF1 (N9279, N9275);
and AND4 (N9280, N9271, N8534, N3930, N5976);
nand NAND2 (N9281, N9267, N1406);
or OR2 (N9282, N9280, N9240);
not NOT1 (N9283, N9276);
not NOT1 (N9284, N9272);
and AND2 (N9285, N9263, N8593);
not NOT1 (N9286, N9283);
xor XOR2 (N9287, N9284, N364);
and AND2 (N9288, N9258, N5254);
not NOT1 (N9289, N9288);
buf BUF1 (N9290, N9289);
or OR2 (N9291, N9279, N4547);
and AND4 (N9292, N9290, N571, N3777, N1453);
buf BUF1 (N9293, N9291);
and AND2 (N9294, N9274, N4743);
not NOT1 (N9295, N9278);
nor NOR4 (N9296, N9282, N2050, N4859, N5789);
not NOT1 (N9297, N9294);
nand NAND3 (N9298, N9286, N7069, N7182);
xor XOR2 (N9299, N9285, N1459);
not NOT1 (N9300, N9298);
or OR4 (N9301, N9293, N864, N20, N4876);
nor NOR3 (N9302, N9295, N5360, N2351);
nor NOR4 (N9303, N9292, N3908, N549, N3266);
xor XOR2 (N9304, N9300, N5467);
buf BUF1 (N9305, N9287);
buf BUF1 (N9306, N9304);
nand NAND4 (N9307, N9281, N368, N7179, N5440);
not NOT1 (N9308, N9303);
buf BUF1 (N9309, N9297);
nand NAND4 (N9310, N9277, N3209, N6266, N4756);
and AND3 (N9311, N9308, N7653, N1322);
nand NAND3 (N9312, N9306, N774, N3257);
xor XOR2 (N9313, N9310, N609);
and AND2 (N9314, N9301, N357);
buf BUF1 (N9315, N9299);
buf BUF1 (N9316, N9312);
buf BUF1 (N9317, N9311);
buf BUF1 (N9318, N9315);
and AND2 (N9319, N9305, N6289);
nand NAND4 (N9320, N9296, N4059, N3408, N4554);
xor XOR2 (N9321, N9313, N1157);
xor XOR2 (N9322, N9302, N7477);
nor NOR2 (N9323, N9314, N4842);
or OR3 (N9324, N9317, N1091, N5885);
or OR4 (N9325, N9323, N8818, N3398, N8551);
and AND2 (N9326, N9316, N7317);
or OR2 (N9327, N9325, N3103);
and AND3 (N9328, N9321, N8093, N7923);
or OR4 (N9329, N9322, N9264, N7031, N3227);
not NOT1 (N9330, N9320);
buf BUF1 (N9331, N9319);
not NOT1 (N9332, N9326);
xor XOR2 (N9333, N9329, N1453);
or OR2 (N9334, N9307, N3197);
buf BUF1 (N9335, N9318);
nand NAND4 (N9336, N9330, N7808, N470, N70);
xor XOR2 (N9337, N9335, N4940);
nor NOR3 (N9338, N9334, N7866, N2915);
or OR2 (N9339, N9324, N4270);
or OR3 (N9340, N9332, N4188, N5687);
buf BUF1 (N9341, N9338);
not NOT1 (N9342, N9337);
not NOT1 (N9343, N9339);
xor XOR2 (N9344, N9340, N4432);
and AND4 (N9345, N9327, N2827, N5028, N6996);
nor NOR2 (N9346, N9342, N1129);
nor NOR4 (N9347, N9328, N1573, N7256, N2651);
and AND2 (N9348, N9331, N1400);
nand NAND2 (N9349, N9347, N5591);
nor NOR3 (N9350, N9333, N1444, N7506);
and AND4 (N9351, N9309, N4734, N7563, N2778);
not NOT1 (N9352, N9351);
xor XOR2 (N9353, N9349, N4406);
not NOT1 (N9354, N9344);
not NOT1 (N9355, N9343);
nor NOR3 (N9356, N9354, N819, N3622);
buf BUF1 (N9357, N9345);
not NOT1 (N9358, N9336);
or OR4 (N9359, N9348, N646, N6550, N7632);
or OR4 (N9360, N9359, N3759, N7899, N2483);
not NOT1 (N9361, N9346);
xor XOR2 (N9362, N9356, N1902);
nor NOR2 (N9363, N9358, N2860);
not NOT1 (N9364, N9350);
xor XOR2 (N9365, N9364, N8248);
nor NOR2 (N9366, N9365, N6202);
nor NOR2 (N9367, N9352, N204);
buf BUF1 (N9368, N9361);
buf BUF1 (N9369, N9357);
not NOT1 (N9370, N9355);
nor NOR3 (N9371, N9353, N7729, N2768);
not NOT1 (N9372, N9366);
or OR3 (N9373, N9372, N8407, N1878);
or OR2 (N9374, N9368, N5980);
and AND2 (N9375, N9341, N5633);
nor NOR3 (N9376, N9360, N6704, N2880);
or OR4 (N9377, N9367, N5119, N552, N5512);
nor NOR2 (N9378, N9374, N3199);
or OR3 (N9379, N9376, N6487, N8028);
nor NOR2 (N9380, N9362, N8265);
not NOT1 (N9381, N9375);
not NOT1 (N9382, N9381);
buf BUF1 (N9383, N9371);
xor XOR2 (N9384, N9383, N3333);
not NOT1 (N9385, N9377);
not NOT1 (N9386, N9385);
nor NOR2 (N9387, N9386, N306);
or OR4 (N9388, N9379, N3385, N2387, N7342);
nand NAND4 (N9389, N9388, N2566, N8183, N3950);
xor XOR2 (N9390, N9387, N1928);
and AND4 (N9391, N9378, N5139, N3675, N9376);
or OR3 (N9392, N9389, N2589, N5843);
not NOT1 (N9393, N9369);
and AND3 (N9394, N9392, N96, N1380);
buf BUF1 (N9395, N9393);
nor NOR3 (N9396, N9394, N7540, N4536);
buf BUF1 (N9397, N9395);
and AND4 (N9398, N9370, N6328, N5098, N8435);
and AND2 (N9399, N9396, N1243);
buf BUF1 (N9400, N9382);
nor NOR4 (N9401, N9391, N3471, N4447, N5181);
or OR4 (N9402, N9363, N1057, N5437, N3930);
nor NOR3 (N9403, N9398, N5894, N3412);
or OR4 (N9404, N9390, N9350, N2986, N7638);
or OR2 (N9405, N9404, N1178);
nor NOR2 (N9406, N9397, N413);
nand NAND3 (N9407, N9405, N1691, N5311);
or OR4 (N9408, N9399, N7496, N9265, N6550);
buf BUF1 (N9409, N9400);
xor XOR2 (N9410, N9408, N2952);
or OR2 (N9411, N9384, N5011);
nor NOR2 (N9412, N9411, N3210);
buf BUF1 (N9413, N9409);
or OR3 (N9414, N9410, N228, N1190);
not NOT1 (N9415, N9406);
nor NOR4 (N9416, N9373, N4319, N1906, N1008);
xor XOR2 (N9417, N9415, N28);
nand NAND4 (N9418, N9403, N4005, N1829, N8408);
and AND4 (N9419, N9418, N78, N6307, N6758);
nand NAND2 (N9420, N9401, N859);
buf BUF1 (N9421, N9407);
or OR4 (N9422, N9402, N265, N4689, N7765);
nor NOR2 (N9423, N9414, N2677);
xor XOR2 (N9424, N9413, N1851);
nor NOR3 (N9425, N9419, N2466, N5961);
nand NAND4 (N9426, N9422, N1119, N60, N6135);
xor XOR2 (N9427, N9412, N5498);
nor NOR2 (N9428, N9421, N3028);
xor XOR2 (N9429, N9426, N802);
nor NOR4 (N9430, N9416, N6307, N79, N8145);
nand NAND4 (N9431, N9424, N3994, N3773, N8374);
nand NAND2 (N9432, N9428, N805);
xor XOR2 (N9433, N9429, N6207);
nor NOR3 (N9434, N9417, N1709, N7797);
or OR3 (N9435, N9434, N2505, N8610);
buf BUF1 (N9436, N9423);
and AND2 (N9437, N9430, N971);
not NOT1 (N9438, N9437);
nand NAND3 (N9439, N9435, N2058, N7235);
nor NOR3 (N9440, N9433, N1840, N6974);
or OR3 (N9441, N9439, N4374, N4371);
buf BUF1 (N9442, N9425);
nor NOR3 (N9443, N9427, N6566, N3060);
buf BUF1 (N9444, N9436);
or OR3 (N9445, N9444, N1832, N6507);
and AND2 (N9446, N9420, N3132);
or OR4 (N9447, N9442, N247, N2419, N9312);
xor XOR2 (N9448, N9443, N8353);
xor XOR2 (N9449, N9448, N5680);
or OR4 (N9450, N9449, N9280, N5994, N2130);
xor XOR2 (N9451, N9431, N8825);
not NOT1 (N9452, N9380);
xor XOR2 (N9453, N9441, N4677);
or OR3 (N9454, N9453, N5609, N3684);
buf BUF1 (N9455, N9452);
xor XOR2 (N9456, N9450, N7184);
not NOT1 (N9457, N9456);
buf BUF1 (N9458, N9451);
not NOT1 (N9459, N9445);
buf BUF1 (N9460, N9459);
not NOT1 (N9461, N9455);
nor NOR4 (N9462, N9446, N3084, N857, N76);
buf BUF1 (N9463, N9458);
or OR4 (N9464, N9454, N7742, N2911, N1009);
not NOT1 (N9465, N9460);
buf BUF1 (N9466, N9463);
or OR3 (N9467, N9432, N4345, N3557);
and AND4 (N9468, N9465, N8270, N8945, N5504);
nor NOR2 (N9469, N9447, N4963);
not NOT1 (N9470, N9464);
and AND3 (N9471, N9467, N8577, N8542);
and AND2 (N9472, N9457, N5926);
nand NAND4 (N9473, N9471, N753, N4113, N370);
xor XOR2 (N9474, N9473, N3680);
xor XOR2 (N9475, N9438, N7363);
not NOT1 (N9476, N9469);
not NOT1 (N9477, N9462);
xor XOR2 (N9478, N9461, N2404);
not NOT1 (N9479, N9477);
buf BUF1 (N9480, N9474);
and AND3 (N9481, N9480, N1166, N5921);
and AND4 (N9482, N9475, N2967, N2135, N4539);
or OR4 (N9483, N9470, N8217, N8365, N676);
not NOT1 (N9484, N9440);
xor XOR2 (N9485, N9476, N6353);
or OR3 (N9486, N9485, N854, N1151);
nor NOR4 (N9487, N9486, N6975, N2479, N4366);
nand NAND2 (N9488, N9468, N2987);
nor NOR4 (N9489, N9487, N1058, N6841, N4354);
and AND2 (N9490, N9482, N8084);
or OR3 (N9491, N9466, N4068, N7248);
not NOT1 (N9492, N9489);
buf BUF1 (N9493, N9479);
and AND3 (N9494, N9492, N9103, N2395);
and AND3 (N9495, N9491, N2708, N8693);
not NOT1 (N9496, N9481);
nor NOR3 (N9497, N9493, N9420, N1610);
nor NOR2 (N9498, N9496, N5468);
nand NAND4 (N9499, N9488, N2283, N2476, N6451);
not NOT1 (N9500, N9495);
and AND3 (N9501, N9499, N2638, N3190);
buf BUF1 (N9502, N9484);
or OR2 (N9503, N9498, N3917);
buf BUF1 (N9504, N9503);
not NOT1 (N9505, N9494);
nand NAND3 (N9506, N9483, N4707, N7984);
nor NOR4 (N9507, N9497, N8568, N5696, N3741);
and AND4 (N9508, N9504, N6727, N4027, N3272);
and AND2 (N9509, N9472, N3095);
not NOT1 (N9510, N9505);
nand NAND3 (N9511, N9506, N2847, N1057);
not NOT1 (N9512, N9511);
nor NOR3 (N9513, N9500, N2041, N6182);
and AND2 (N9514, N9478, N8585);
not NOT1 (N9515, N9490);
or OR4 (N9516, N9512, N3981, N9477, N4497);
and AND3 (N9517, N9515, N2337, N3324);
nor NOR3 (N9518, N9509, N619, N4754);
nor NOR3 (N9519, N9516, N783, N7381);
buf BUF1 (N9520, N9514);
not NOT1 (N9521, N9513);
not NOT1 (N9522, N9517);
xor XOR2 (N9523, N9501, N4378);
buf BUF1 (N9524, N9521);
not NOT1 (N9525, N9522);
buf BUF1 (N9526, N9525);
nor NOR4 (N9527, N9518, N9107, N8083, N7939);
or OR3 (N9528, N9519, N3332, N947);
or OR2 (N9529, N9510, N310);
nand NAND4 (N9530, N9520, N7341, N7201, N8270);
or OR2 (N9531, N9527, N5489);
or OR3 (N9532, N9526, N5633, N7503);
buf BUF1 (N9533, N9508);
nand NAND4 (N9534, N9523, N3989, N8767, N8433);
not NOT1 (N9535, N9502);
xor XOR2 (N9536, N9524, N6337);
or OR3 (N9537, N9530, N4534, N6952);
buf BUF1 (N9538, N9537);
not NOT1 (N9539, N9532);
and AND4 (N9540, N9529, N5079, N7287, N8573);
not NOT1 (N9541, N9535);
buf BUF1 (N9542, N9507);
nand NAND3 (N9543, N9528, N7066, N3147);
and AND3 (N9544, N9534, N7847, N3733);
not NOT1 (N9545, N9538);
not NOT1 (N9546, N9540);
nor NOR3 (N9547, N9539, N255, N9020);
and AND4 (N9548, N9546, N4440, N3056, N7541);
buf BUF1 (N9549, N9533);
or OR3 (N9550, N9544, N5559, N3496);
nand NAND4 (N9551, N9549, N8552, N994, N2831);
nand NAND2 (N9552, N9551, N5303);
nor NOR2 (N9553, N9552, N1624);
nor NOR3 (N9554, N9545, N4022, N6892);
nand NAND4 (N9555, N9543, N7650, N2993, N6364);
buf BUF1 (N9556, N9550);
nor NOR2 (N9557, N9547, N9364);
and AND2 (N9558, N9554, N6892);
or OR4 (N9559, N9542, N7506, N8388, N9263);
buf BUF1 (N9560, N9558);
xor XOR2 (N9561, N9531, N7927);
buf BUF1 (N9562, N9553);
or OR2 (N9563, N9562, N1769);
and AND3 (N9564, N9563, N504, N571);
xor XOR2 (N9565, N9548, N7940);
nor NOR2 (N9566, N9555, N1893);
xor XOR2 (N9567, N9564, N6403);
buf BUF1 (N9568, N9556);
or OR3 (N9569, N9560, N1897, N604);
buf BUF1 (N9570, N9557);
buf BUF1 (N9571, N9565);
or OR3 (N9572, N9569, N7831, N8761);
nor NOR3 (N9573, N9566, N6260, N6121);
buf BUF1 (N9574, N9570);
nor NOR3 (N9575, N9574, N8531, N7205);
not NOT1 (N9576, N9573);
and AND3 (N9577, N9536, N4895, N2558);
xor XOR2 (N9578, N9568, N7751);
and AND3 (N9579, N9571, N3898, N2927);
xor XOR2 (N9580, N9575, N9302);
buf BUF1 (N9581, N9578);
or OR3 (N9582, N9581, N7370, N4669);
not NOT1 (N9583, N9559);
nor NOR3 (N9584, N9561, N8955, N150);
not NOT1 (N9585, N9579);
buf BUF1 (N9586, N9572);
and AND3 (N9587, N9577, N8613, N1235);
nor NOR2 (N9588, N9583, N4111);
and AND4 (N9589, N9580, N2081, N8047, N2026);
and AND2 (N9590, N9567, N8576);
and AND4 (N9591, N9587, N8851, N3477, N9180);
xor XOR2 (N9592, N9584, N4317);
not NOT1 (N9593, N9586);
or OR2 (N9594, N9541, N2972);
and AND2 (N9595, N9588, N6918);
and AND4 (N9596, N9590, N6220, N7741, N6421);
or OR3 (N9597, N9591, N5857, N9121);
nand NAND2 (N9598, N9593, N5873);
and AND3 (N9599, N9594, N6172, N3605);
and AND4 (N9600, N9595, N7212, N3938, N4408);
nand NAND3 (N9601, N9599, N7941, N8016);
not NOT1 (N9602, N9582);
and AND2 (N9603, N9596, N4565);
xor XOR2 (N9604, N9592, N16);
buf BUF1 (N9605, N9585);
not NOT1 (N9606, N9597);
buf BUF1 (N9607, N9598);
nand NAND2 (N9608, N9602, N8856);
buf BUF1 (N9609, N9606);
and AND4 (N9610, N9607, N3075, N922, N5302);
not NOT1 (N9611, N9610);
buf BUF1 (N9612, N9611);
not NOT1 (N9613, N9601);
and AND3 (N9614, N9605, N7108, N4147);
not NOT1 (N9615, N9612);
buf BUF1 (N9616, N9613);
and AND2 (N9617, N9614, N3708);
buf BUF1 (N9618, N9576);
xor XOR2 (N9619, N9615, N1322);
or OR3 (N9620, N9619, N5207, N6669);
xor XOR2 (N9621, N9589, N80);
and AND2 (N9622, N9620, N8898);
or OR3 (N9623, N9603, N102, N1357);
nand NAND4 (N9624, N9600, N254, N9483, N446);
buf BUF1 (N9625, N9618);
xor XOR2 (N9626, N9624, N8195);
not NOT1 (N9627, N9625);
nand NAND2 (N9628, N9627, N3637);
and AND2 (N9629, N9623, N7924);
not NOT1 (N9630, N9622);
buf BUF1 (N9631, N9628);
and AND4 (N9632, N9616, N3738, N8516, N6855);
or OR4 (N9633, N9632, N1508, N6403, N6174);
or OR3 (N9634, N9617, N4345, N7273);
xor XOR2 (N9635, N9608, N1433);
nand NAND2 (N9636, N9634, N9150);
buf BUF1 (N9637, N9609);
not NOT1 (N9638, N9633);
xor XOR2 (N9639, N9630, N7709);
buf BUF1 (N9640, N9636);
or OR3 (N9641, N9638, N2431, N3815);
and AND2 (N9642, N9604, N1242);
and AND4 (N9643, N9639, N7070, N5199, N7197);
not NOT1 (N9644, N9637);
nand NAND3 (N9645, N9629, N4574, N915);
buf BUF1 (N9646, N9621);
nand NAND4 (N9647, N9626, N9466, N3528, N8733);
nor NOR2 (N9648, N9644, N6577);
or OR2 (N9649, N9645, N3219);
nor NOR3 (N9650, N9642, N520, N5178);
nor NOR2 (N9651, N9650, N8238);
nand NAND4 (N9652, N9641, N9590, N2398, N9586);
and AND2 (N9653, N9652, N9414);
or OR2 (N9654, N9648, N281);
or OR2 (N9655, N9651, N5535);
nor NOR4 (N9656, N9631, N3192, N4595, N2432);
nand NAND2 (N9657, N9646, N5484);
nand NAND4 (N9658, N9655, N5714, N305, N4287);
or OR2 (N9659, N9635, N9643);
buf BUF1 (N9660, N3851);
buf BUF1 (N9661, N9656);
and AND3 (N9662, N9640, N4905, N5690);
buf BUF1 (N9663, N9647);
and AND2 (N9664, N9653, N3856);
or OR4 (N9665, N9662, N8614, N4445, N4524);
nand NAND3 (N9666, N9654, N8554, N2561);
and AND3 (N9667, N9664, N239, N2977);
xor XOR2 (N9668, N9665, N7581);
buf BUF1 (N9669, N9667);
not NOT1 (N9670, N9657);
not NOT1 (N9671, N9660);
or OR2 (N9672, N9666, N1609);
nand NAND4 (N9673, N9670, N6612, N8992, N9456);
not NOT1 (N9674, N9661);
and AND2 (N9675, N9674, N1624);
not NOT1 (N9676, N9659);
buf BUF1 (N9677, N9673);
nor NOR4 (N9678, N9672, N7297, N7682, N9362);
not NOT1 (N9679, N9658);
nand NAND3 (N9680, N9669, N5802, N2076);
or OR2 (N9681, N9677, N1745);
xor XOR2 (N9682, N9679, N903);
xor XOR2 (N9683, N9671, N9194);
nand NAND3 (N9684, N9668, N383, N793);
xor XOR2 (N9685, N9678, N9584);
and AND2 (N9686, N9675, N7516);
nand NAND2 (N9687, N9681, N8137);
buf BUF1 (N9688, N9649);
or OR4 (N9689, N9680, N8347, N3509, N4057);
xor XOR2 (N9690, N9686, N1466);
nor NOR3 (N9691, N9689, N4333, N3168);
nand NAND4 (N9692, N9684, N3797, N778, N6991);
and AND4 (N9693, N9691, N3582, N9546, N6288);
nand NAND2 (N9694, N9688, N6058);
and AND3 (N9695, N9685, N4404, N3614);
and AND2 (N9696, N9676, N7451);
buf BUF1 (N9697, N9683);
nor NOR2 (N9698, N9697, N8863);
buf BUF1 (N9699, N9696);
buf BUF1 (N9700, N9682);
not NOT1 (N9701, N9695);
xor XOR2 (N9702, N9694, N6120);
buf BUF1 (N9703, N9690);
nor NOR4 (N9704, N9693, N1037, N84, N9110);
and AND2 (N9705, N9699, N7258);
and AND3 (N9706, N9702, N6759, N2080);
nand NAND4 (N9707, N9704, N2637, N6268, N5709);
not NOT1 (N9708, N9706);
nand NAND4 (N9709, N9698, N7141, N1704, N1350);
xor XOR2 (N9710, N9701, N5751);
nand NAND3 (N9711, N9709, N9529, N1213);
or OR4 (N9712, N9687, N5178, N5693, N581);
not NOT1 (N9713, N9708);
xor XOR2 (N9714, N9713, N4024);
nand NAND2 (N9715, N9714, N952);
nand NAND2 (N9716, N9692, N2445);
not NOT1 (N9717, N9711);
xor XOR2 (N9718, N9700, N3998);
nand NAND2 (N9719, N9716, N2434);
and AND3 (N9720, N9718, N6971, N2162);
nor NOR4 (N9721, N9720, N6124, N3428, N2189);
xor XOR2 (N9722, N9721, N5788);
nor NOR4 (N9723, N9722, N1959, N1781, N7302);
nand NAND4 (N9724, N9703, N6691, N9709, N3114);
not NOT1 (N9725, N9723);
nand NAND3 (N9726, N9715, N6919, N5763);
or OR3 (N9727, N9726, N3777, N1525);
or OR2 (N9728, N9724, N9432);
and AND3 (N9729, N9707, N4173, N4688);
and AND3 (N9730, N9717, N9410, N6975);
xor XOR2 (N9731, N9705, N7474);
nor NOR2 (N9732, N9663, N5027);
nor NOR4 (N9733, N9731, N9666, N1533, N8819);
nand NAND2 (N9734, N9712, N5501);
xor XOR2 (N9735, N9732, N6089);
and AND2 (N9736, N9733, N1810);
nand NAND3 (N9737, N9728, N6891, N5885);
and AND2 (N9738, N9725, N2917);
xor XOR2 (N9739, N9730, N7717);
buf BUF1 (N9740, N9735);
nor NOR4 (N9741, N9734, N1047, N1130, N4123);
buf BUF1 (N9742, N9729);
xor XOR2 (N9743, N9719, N3227);
and AND2 (N9744, N9741, N720);
buf BUF1 (N9745, N9727);
xor XOR2 (N9746, N9743, N517);
or OR3 (N9747, N9710, N6545, N4701);
nand NAND2 (N9748, N9746, N2803);
or OR4 (N9749, N9738, N5455, N2200, N7120);
buf BUF1 (N9750, N9742);
xor XOR2 (N9751, N9747, N4093);
buf BUF1 (N9752, N9737);
or OR4 (N9753, N9745, N7269, N9155, N9530);
not NOT1 (N9754, N9740);
xor XOR2 (N9755, N9736, N2133);
or OR4 (N9756, N9754, N8261, N2550, N3402);
or OR4 (N9757, N9752, N2020, N8334, N7906);
buf BUF1 (N9758, N9756);
nand NAND3 (N9759, N9750, N3657, N7519);
nor NOR3 (N9760, N9749, N6994, N1373);
not NOT1 (N9761, N9760);
or OR3 (N9762, N9753, N8360, N419);
nor NOR3 (N9763, N9739, N8765, N8580);
not NOT1 (N9764, N9751);
nor NOR2 (N9765, N9755, N7487);
and AND4 (N9766, N9763, N16, N622, N7619);
buf BUF1 (N9767, N9748);
and AND3 (N9768, N9758, N3052, N5548);
nand NAND2 (N9769, N9764, N874);
and AND4 (N9770, N9759, N4063, N997, N1876);
nand NAND2 (N9771, N9767, N4408);
buf BUF1 (N9772, N9744);
and AND2 (N9773, N9757, N4810);
not NOT1 (N9774, N9768);
and AND2 (N9775, N9765, N4588);
nor NOR3 (N9776, N9771, N4922, N5593);
not NOT1 (N9777, N9773);
and AND3 (N9778, N9766, N4417, N5027);
not NOT1 (N9779, N9775);
nand NAND2 (N9780, N9761, N4030);
nand NAND4 (N9781, N9776, N6590, N7812, N2158);
nor NOR2 (N9782, N9781, N8439);
not NOT1 (N9783, N9770);
or OR2 (N9784, N9782, N202);
or OR3 (N9785, N9769, N6340, N6626);
nor NOR2 (N9786, N9784, N6510);
xor XOR2 (N9787, N9785, N4178);
not NOT1 (N9788, N9786);
xor XOR2 (N9789, N9762, N4062);
or OR3 (N9790, N9779, N1879, N176);
and AND4 (N9791, N9788, N3158, N7700, N5018);
nand NAND3 (N9792, N9789, N37, N2484);
xor XOR2 (N9793, N9774, N167);
or OR2 (N9794, N9778, N2846);
buf BUF1 (N9795, N9780);
buf BUF1 (N9796, N9783);
or OR4 (N9797, N9794, N9343, N6332, N2584);
buf BUF1 (N9798, N9777);
not NOT1 (N9799, N9790);
and AND2 (N9800, N9793, N7707);
or OR4 (N9801, N9799, N9416, N1228, N9475);
nand NAND3 (N9802, N9801, N1073, N191);
or OR3 (N9803, N9800, N7126, N3853);
or OR3 (N9804, N9802, N2065, N8025);
nand NAND2 (N9805, N9791, N2461);
and AND2 (N9806, N9804, N8814);
xor XOR2 (N9807, N9795, N5782);
nor NOR2 (N9808, N9787, N5455);
xor XOR2 (N9809, N9806, N892);
nand NAND4 (N9810, N9797, N1192, N5805, N669);
xor XOR2 (N9811, N9805, N3816);
nor NOR3 (N9812, N9808, N3026, N9439);
and AND2 (N9813, N9809, N177);
not NOT1 (N9814, N9798);
not NOT1 (N9815, N9796);
or OR2 (N9816, N9803, N6950);
not NOT1 (N9817, N9792);
and AND4 (N9818, N9772, N1021, N4888, N1010);
buf BUF1 (N9819, N9810);
nor NOR3 (N9820, N9819, N8565, N7245);
nand NAND2 (N9821, N9813, N4450);
not NOT1 (N9822, N9812);
buf BUF1 (N9823, N9818);
not NOT1 (N9824, N9817);
and AND2 (N9825, N9824, N1671);
or OR3 (N9826, N9820, N15, N6158);
and AND4 (N9827, N9814, N4395, N1197, N2698);
nor NOR3 (N9828, N9811, N3807, N814);
nor NOR2 (N9829, N9823, N1521);
not NOT1 (N9830, N9827);
nand NAND2 (N9831, N9830, N7471);
nand NAND3 (N9832, N9822, N5748, N7700);
buf BUF1 (N9833, N9826);
nor NOR2 (N9834, N9825, N3030);
xor XOR2 (N9835, N9815, N5462);
buf BUF1 (N9836, N9835);
or OR3 (N9837, N9836, N7826, N2877);
or OR3 (N9838, N9834, N8528, N5267);
buf BUF1 (N9839, N9838);
nor NOR3 (N9840, N9833, N3991, N5318);
nand NAND4 (N9841, N9816, N481, N7596, N2812);
nand NAND2 (N9842, N9832, N3390);
xor XOR2 (N9843, N9841, N4836);
not NOT1 (N9844, N9807);
and AND2 (N9845, N9831, N9710);
xor XOR2 (N9846, N9828, N728);
xor XOR2 (N9847, N9829, N88);
buf BUF1 (N9848, N9844);
nor NOR2 (N9849, N9840, N7860);
and AND4 (N9850, N9843, N2623, N6772, N1377);
and AND4 (N9851, N9850, N9079, N2124, N9115);
xor XOR2 (N9852, N9837, N2660);
xor XOR2 (N9853, N9849, N734);
buf BUF1 (N9854, N9821);
nor NOR2 (N9855, N9851, N5241);
nand NAND3 (N9856, N9842, N9417, N3094);
xor XOR2 (N9857, N9854, N4619);
not NOT1 (N9858, N9845);
or OR4 (N9859, N9847, N705, N5981, N1744);
nand NAND3 (N9860, N9858, N5724, N3557);
not NOT1 (N9861, N9853);
and AND3 (N9862, N9861, N4036, N4651);
buf BUF1 (N9863, N9862);
and AND4 (N9864, N9857, N9637, N6053, N7734);
buf BUF1 (N9865, N9839);
or OR3 (N9866, N9863, N9243, N3273);
and AND3 (N9867, N9856, N5034, N7736);
and AND3 (N9868, N9848, N4938, N2650);
xor XOR2 (N9869, N9860, N5735);
buf BUF1 (N9870, N9865);
and AND2 (N9871, N9867, N9730);
buf BUF1 (N9872, N9868);
nand NAND2 (N9873, N9872, N2852);
and AND2 (N9874, N9869, N5079);
nand NAND4 (N9875, N9864, N5239, N5371, N5292);
buf BUF1 (N9876, N9855);
buf BUF1 (N9877, N9876);
not NOT1 (N9878, N9866);
nand NAND2 (N9879, N9873, N2598);
or OR4 (N9880, N9877, N7348, N7427, N6078);
nor NOR3 (N9881, N9859, N9811, N6426);
buf BUF1 (N9882, N9874);
or OR2 (N9883, N9882, N1872);
nand NAND2 (N9884, N9875, N616);
xor XOR2 (N9885, N9871, N5888);
not NOT1 (N9886, N9880);
nand NAND4 (N9887, N9881, N5936, N5193, N7143);
nor NOR4 (N9888, N9884, N4751, N396, N8236);
nand NAND3 (N9889, N9846, N2730, N3608);
buf BUF1 (N9890, N9879);
and AND4 (N9891, N9887, N8720, N8007, N50);
and AND3 (N9892, N9852, N7343, N4454);
nor NOR4 (N9893, N9890, N8010, N8957, N8864);
nand NAND2 (N9894, N9870, N852);
buf BUF1 (N9895, N9894);
xor XOR2 (N9896, N9892, N9001);
and AND4 (N9897, N9888, N547, N7620, N7693);
or OR2 (N9898, N9895, N1740);
buf BUF1 (N9899, N9878);
xor XOR2 (N9900, N9885, N8889);
buf BUF1 (N9901, N9889);
not NOT1 (N9902, N9886);
xor XOR2 (N9903, N9902, N883);
nor NOR4 (N9904, N9898, N6285, N7379, N4495);
not NOT1 (N9905, N9904);
or OR4 (N9906, N9901, N5479, N1684, N8696);
not NOT1 (N9907, N9893);
buf BUF1 (N9908, N9899);
nand NAND3 (N9909, N9883, N7440, N1061);
or OR3 (N9910, N9905, N4657, N5132);
or OR3 (N9911, N9896, N5303, N585);
or OR2 (N9912, N9897, N9527);
nand NAND3 (N9913, N9907, N6165, N5877);
nand NAND4 (N9914, N9908, N3311, N85, N1233);
or OR4 (N9915, N9903, N768, N7343, N7444);
nor NOR4 (N9916, N9912, N1790, N2991, N5425);
or OR3 (N9917, N9915, N1250, N8475);
not NOT1 (N9918, N9917);
nand NAND4 (N9919, N9913, N7906, N2508, N6692);
not NOT1 (N9920, N9911);
nor NOR3 (N9921, N9906, N1506, N3759);
or OR3 (N9922, N9914, N7566, N2452);
or OR2 (N9923, N9919, N4836);
nor NOR4 (N9924, N9900, N5641, N6982, N7084);
nor NOR3 (N9925, N9923, N7388, N3221);
nand NAND3 (N9926, N9922, N7267, N4504);
xor XOR2 (N9927, N9924, N872);
or OR3 (N9928, N9891, N8950, N5084);
and AND3 (N9929, N9927, N1304, N7403);
buf BUF1 (N9930, N9921);
not NOT1 (N9931, N9916);
buf BUF1 (N9932, N9909);
or OR4 (N9933, N9910, N9779, N8332, N9130);
or OR2 (N9934, N9920, N3919);
nor NOR2 (N9935, N9932, N8087);
buf BUF1 (N9936, N9929);
xor XOR2 (N9937, N9926, N6399);
xor XOR2 (N9938, N9937, N9801);
nand NAND3 (N9939, N9925, N5174, N7899);
or OR3 (N9940, N9933, N5327, N7021);
nor NOR4 (N9941, N9939, N9480, N8660, N692);
buf BUF1 (N9942, N9930);
and AND3 (N9943, N9941, N4104, N7662);
nand NAND3 (N9944, N9935, N584, N1226);
not NOT1 (N9945, N9940);
not NOT1 (N9946, N9944);
and AND4 (N9947, N9945, N5048, N1860, N937);
nor NOR3 (N9948, N9934, N5342, N1592);
or OR2 (N9949, N9928, N8883);
nand NAND2 (N9950, N9938, N9391);
or OR2 (N9951, N9950, N9554);
xor XOR2 (N9952, N9947, N3012);
xor XOR2 (N9953, N9949, N5415);
nor NOR3 (N9954, N9918, N5257, N3399);
nor NOR4 (N9955, N9952, N6050, N5599, N138);
and AND3 (N9956, N9942, N6513, N7651);
xor XOR2 (N9957, N9948, N2692);
not NOT1 (N9958, N9954);
not NOT1 (N9959, N9957);
or OR3 (N9960, N9959, N5549, N8301);
not NOT1 (N9961, N9955);
nor NOR2 (N9962, N9953, N2977);
buf BUF1 (N9963, N9936);
buf BUF1 (N9964, N9956);
not NOT1 (N9965, N9931);
xor XOR2 (N9966, N9963, N8137);
nand NAND3 (N9967, N9964, N5231, N2174);
not NOT1 (N9968, N9943);
nand NAND4 (N9969, N9965, N9589, N4081, N5338);
xor XOR2 (N9970, N9946, N319);
xor XOR2 (N9971, N9966, N4201);
not NOT1 (N9972, N9960);
or OR4 (N9973, N9967, N7786, N5106, N3519);
and AND3 (N9974, N9961, N7651, N6474);
buf BUF1 (N9975, N9970);
buf BUF1 (N9976, N9951);
not NOT1 (N9977, N9971);
buf BUF1 (N9978, N9969);
nor NOR3 (N9979, N9958, N4662, N2490);
and AND3 (N9980, N9976, N5615, N29);
nor NOR4 (N9981, N9978, N6712, N9809, N7565);
not NOT1 (N9982, N9980);
or OR2 (N9983, N9975, N3378);
and AND2 (N9984, N9981, N6739);
not NOT1 (N9985, N9973);
xor XOR2 (N9986, N9982, N8926);
not NOT1 (N9987, N9972);
nand NAND3 (N9988, N9984, N6396, N4237);
nand NAND3 (N9989, N9985, N7500, N6739);
not NOT1 (N9990, N9983);
nor NOR4 (N9991, N9988, N6459, N4097, N2228);
nand NAND3 (N9992, N9979, N9533, N635);
or OR2 (N9993, N9962, N1178);
and AND3 (N9994, N9990, N940, N6011);
or OR2 (N9995, N9991, N6951);
buf BUF1 (N9996, N9992);
buf BUF1 (N9997, N9986);
nand NAND4 (N9998, N9989, N3757, N3147, N6094);
xor XOR2 (N9999, N9993, N8031);
nor NOR2 (N10000, N9998, N3931);
and AND3 (N10001, N9987, N330, N9243);
nor NOR4 (N10002, N9997, N2152, N977, N6268);
xor XOR2 (N10003, N9994, N4415);
buf BUF1 (N10004, N9999);
not NOT1 (N10005, N10002);
nand NAND3 (N10006, N9977, N231, N7691);
nor NOR2 (N10007, N9974, N6052);
xor XOR2 (N10008, N9995, N2413);
nand NAND3 (N10009, N10008, N7515, N9606);
and AND4 (N10010, N10007, N6728, N3518, N1671);
or OR2 (N10011, N9968, N5001);
nand NAND3 (N10012, N10010, N1691, N4973);
not NOT1 (N10013, N10000);
nor NOR3 (N10014, N9996, N1546, N2008);
not NOT1 (N10015, N10012);
xor XOR2 (N10016, N10011, N3074);
or OR3 (N10017, N10003, N6457, N6909);
nand NAND2 (N10018, N10016, N7419);
or OR2 (N10019, N10015, N2533);
buf BUF1 (N10020, N10019);
not NOT1 (N10021, N10005);
xor XOR2 (N10022, N10017, N706);
or OR3 (N10023, N10006, N2765, N8947);
not NOT1 (N10024, N10023);
nand NAND4 (N10025, N10024, N7708, N6026, N9842);
buf BUF1 (N10026, N10004);
or OR4 (N10027, N10018, N1048, N3893, N3142);
nand NAND2 (N10028, N10013, N2893);
and AND3 (N10029, N10026, N5104, N8154);
xor XOR2 (N10030, N10027, N6152);
nor NOR4 (N10031, N10009, N3130, N3119, N5902);
not NOT1 (N10032, N10014);
and AND2 (N10033, N10031, N7639);
xor XOR2 (N10034, N10030, N5886);
or OR4 (N10035, N10029, N9830, N5636, N3316);
nand NAND4 (N10036, N10028, N4665, N8509, N4086);
not NOT1 (N10037, N10022);
buf BUF1 (N10038, N10034);
buf BUF1 (N10039, N10032);
nor NOR3 (N10040, N10021, N1171, N9842);
nand NAND3 (N10041, N10020, N220, N8122);
and AND4 (N10042, N10038, N3527, N8915, N5751);
or OR2 (N10043, N10042, N7894);
buf BUF1 (N10044, N10040);
and AND3 (N10045, N10001, N190, N7419);
and AND3 (N10046, N10044, N38, N433);
not NOT1 (N10047, N10036);
and AND4 (N10048, N10039, N36, N8215, N2297);
or OR2 (N10049, N10043, N5336);
and AND3 (N10050, N10045, N3752, N519);
xor XOR2 (N10051, N10025, N7182);
or OR4 (N10052, N10051, N246, N9913, N3623);
nand NAND3 (N10053, N10050, N2103, N5517);
buf BUF1 (N10054, N10053);
and AND4 (N10055, N10035, N5114, N7428, N2852);
xor XOR2 (N10056, N10046, N6721);
buf BUF1 (N10057, N10056);
buf BUF1 (N10058, N10057);
xor XOR2 (N10059, N10048, N437);
buf BUF1 (N10060, N10047);
xor XOR2 (N10061, N10058, N3273);
not NOT1 (N10062, N10033);
nand NAND4 (N10063, N10059, N8036, N832, N1748);
xor XOR2 (N10064, N10049, N7930);
and AND4 (N10065, N10060, N1871, N2012, N4268);
buf BUF1 (N10066, N10062);
and AND2 (N10067, N10061, N8532);
nand NAND4 (N10068, N10055, N700, N720, N5893);
xor XOR2 (N10069, N10064, N8547);
not NOT1 (N10070, N10063);
xor XOR2 (N10071, N10041, N1783);
and AND4 (N10072, N10065, N7685, N8590, N4998);
not NOT1 (N10073, N10071);
not NOT1 (N10074, N10037);
not NOT1 (N10075, N10070);
and AND4 (N10076, N10054, N7576, N7201, N7729);
buf BUF1 (N10077, N10052);
nand NAND3 (N10078, N10067, N3421, N9717);
not NOT1 (N10079, N10077);
nand NAND4 (N10080, N10079, N9715, N1295, N5217);
not NOT1 (N10081, N10080);
or OR3 (N10082, N10074, N4414, N2993);
xor XOR2 (N10083, N10082, N81);
nor NOR3 (N10084, N10078, N6196, N7114);
or OR2 (N10085, N10069, N6132);
not NOT1 (N10086, N10068);
buf BUF1 (N10087, N10081);
and AND4 (N10088, N10072, N5497, N9179, N6058);
xor XOR2 (N10089, N10088, N6926);
xor XOR2 (N10090, N10087, N3345);
and AND4 (N10091, N10090, N8290, N9916, N5761);
nand NAND2 (N10092, N10083, N3899);
nand NAND4 (N10093, N10076, N9406, N9198, N2507);
nor NOR4 (N10094, N10073, N4331, N3118, N181);
nor NOR4 (N10095, N10093, N5978, N4235, N3775);
nor NOR3 (N10096, N10084, N1211, N4741);
xor XOR2 (N10097, N10095, N4770);
xor XOR2 (N10098, N10096, N3145);
nand NAND2 (N10099, N10094, N6018);
xor XOR2 (N10100, N10092, N2052);
nand NAND4 (N10101, N10089, N8503, N123, N9130);
nor NOR3 (N10102, N10066, N1216, N7301);
or OR2 (N10103, N10101, N7125);
nand NAND2 (N10104, N10100, N4104);
nand NAND2 (N10105, N10102, N8718);
not NOT1 (N10106, N10099);
and AND3 (N10107, N10105, N9229, N7798);
nand NAND4 (N10108, N10107, N2081, N4387, N8001);
and AND3 (N10109, N10085, N5276, N3433);
or OR3 (N10110, N10091, N8694, N2759);
or OR4 (N10111, N10104, N1008, N5145, N5189);
buf BUF1 (N10112, N10106);
not NOT1 (N10113, N10097);
buf BUF1 (N10114, N10098);
nand NAND3 (N10115, N10109, N1395, N1002);
and AND2 (N10116, N10111, N1327);
and AND2 (N10117, N10112, N2861);
or OR3 (N10118, N10116, N7513, N3157);
xor XOR2 (N10119, N10075, N467);
buf BUF1 (N10120, N10113);
nand NAND3 (N10121, N10108, N3802, N6818);
and AND4 (N10122, N10120, N8955, N2273, N3662);
xor XOR2 (N10123, N10118, N7314);
nor NOR2 (N10124, N10119, N3022);
xor XOR2 (N10125, N10103, N63);
and AND4 (N10126, N10123, N5572, N6847, N343);
not NOT1 (N10127, N10086);
and AND3 (N10128, N10125, N309, N1817);
xor XOR2 (N10129, N10122, N3447);
nor NOR4 (N10130, N10115, N6488, N3613, N4812);
not NOT1 (N10131, N10128);
xor XOR2 (N10132, N10129, N4292);
not NOT1 (N10133, N10117);
xor XOR2 (N10134, N10127, N8122);
or OR3 (N10135, N10121, N8511, N8069);
and AND2 (N10136, N10110, N8982);
xor XOR2 (N10137, N10132, N2009);
and AND3 (N10138, N10114, N8376, N7186);
nor NOR4 (N10139, N10130, N6905, N876, N5237);
nand NAND4 (N10140, N10131, N9579, N1024, N4284);
nor NOR4 (N10141, N10124, N7780, N6727, N7034);
xor XOR2 (N10142, N10140, N7139);
nand NAND4 (N10143, N10142, N1723, N2438, N8708);
xor XOR2 (N10144, N10138, N8535);
xor XOR2 (N10145, N10134, N5730);
or OR2 (N10146, N10133, N9905);
buf BUF1 (N10147, N10145);
and AND3 (N10148, N10144, N7646, N9714);
not NOT1 (N10149, N10143);
buf BUF1 (N10150, N10148);
buf BUF1 (N10151, N10137);
nand NAND3 (N10152, N10139, N5079, N3819);
or OR2 (N10153, N10151, N9877);
xor XOR2 (N10154, N10135, N1244);
nor NOR3 (N10155, N10141, N2102, N6100);
nor NOR4 (N10156, N10146, N7775, N8318, N3222);
not NOT1 (N10157, N10152);
nand NAND2 (N10158, N10150, N9749);
nand NAND3 (N10159, N10147, N1980, N1247);
or OR4 (N10160, N10158, N5341, N5354, N2379);
or OR2 (N10161, N10154, N8596);
or OR2 (N10162, N10157, N6094);
and AND4 (N10163, N10149, N6950, N6065, N7045);
not NOT1 (N10164, N10159);
buf BUF1 (N10165, N10156);
nand NAND4 (N10166, N10163, N7708, N9764, N640);
nor NOR3 (N10167, N10161, N7177, N6184);
or OR4 (N10168, N10136, N265, N6690, N4533);
not NOT1 (N10169, N10126);
not NOT1 (N10170, N10166);
nor NOR3 (N10171, N10169, N2331, N4735);
buf BUF1 (N10172, N10160);
and AND4 (N10173, N10155, N2419, N3594, N6541);
xor XOR2 (N10174, N10164, N2553);
buf BUF1 (N10175, N10167);
nand NAND2 (N10176, N10174, N910);
nand NAND2 (N10177, N10175, N1875);
and AND3 (N10178, N10162, N1235, N7688);
not NOT1 (N10179, N10173);
buf BUF1 (N10180, N10171);
buf BUF1 (N10181, N10165);
nand NAND3 (N10182, N10181, N4769, N1680);
nor NOR3 (N10183, N10180, N1676, N2478);
nand NAND4 (N10184, N10153, N8672, N8856, N5953);
buf BUF1 (N10185, N10172);
nand NAND3 (N10186, N10170, N9715, N320);
and AND4 (N10187, N10177, N10007, N8000, N6515);
not NOT1 (N10188, N10176);
nand NAND4 (N10189, N10179, N3303, N5825, N2361);
buf BUF1 (N10190, N10183);
buf BUF1 (N10191, N10188);
nor NOR4 (N10192, N10185, N2819, N7214, N713);
and AND2 (N10193, N10191, N4021);
nor NOR3 (N10194, N10187, N139, N4192);
and AND4 (N10195, N10189, N7532, N5718, N9365);
nor NOR4 (N10196, N10194, N7721, N4071, N7896);
nor NOR3 (N10197, N10192, N8525, N5836);
nand NAND3 (N10198, N10190, N6712, N3783);
buf BUF1 (N10199, N10168);
xor XOR2 (N10200, N10186, N9441);
xor XOR2 (N10201, N10182, N8216);
nand NAND2 (N10202, N10196, N4140);
or OR3 (N10203, N10199, N3509, N8473);
nand NAND4 (N10204, N10197, N9662, N1367, N953);
and AND3 (N10205, N10201, N5936, N8924);
and AND3 (N10206, N10205, N1864, N2565);
buf BUF1 (N10207, N10198);
nand NAND3 (N10208, N10204, N8604, N9295);
nand NAND4 (N10209, N10202, N6483, N1747, N5856);
not NOT1 (N10210, N10193);
buf BUF1 (N10211, N10210);
nand NAND2 (N10212, N10200, N6336);
buf BUF1 (N10213, N10208);
or OR3 (N10214, N10213, N10184, N7810);
not NOT1 (N10215, N2549);
or OR4 (N10216, N10212, N7572, N7592, N2177);
nor NOR2 (N10217, N10203, N5373);
nand NAND2 (N10218, N10207, N897);
not NOT1 (N10219, N10211);
nor NOR2 (N10220, N10206, N7832);
nand NAND2 (N10221, N10214, N6790);
buf BUF1 (N10222, N10220);
buf BUF1 (N10223, N10218);
or OR4 (N10224, N10215, N1493, N4066, N8917);
xor XOR2 (N10225, N10222, N2938);
buf BUF1 (N10226, N10178);
nor NOR2 (N10227, N10219, N2034);
or OR4 (N10228, N10195, N3520, N2572, N6814);
xor XOR2 (N10229, N10209, N383);
nor NOR3 (N10230, N10229, N7408, N9905);
and AND2 (N10231, N10226, N2838);
and AND2 (N10232, N10224, N1650);
and AND4 (N10233, N10230, N8887, N4234, N7168);
or OR4 (N10234, N10227, N3900, N5451, N1254);
nand NAND4 (N10235, N10232, N6821, N975, N2730);
or OR3 (N10236, N10216, N4026, N6991);
xor XOR2 (N10237, N10228, N3849);
or OR3 (N10238, N10234, N2862, N4069);
buf BUF1 (N10239, N10225);
and AND3 (N10240, N10233, N6156, N7894);
or OR4 (N10241, N10223, N2576, N3972, N72);
xor XOR2 (N10242, N10238, N7955);
and AND2 (N10243, N10240, N879);
xor XOR2 (N10244, N10231, N1326);
and AND2 (N10245, N10236, N7761);
nor NOR4 (N10246, N10237, N309, N2344, N7194);
buf BUF1 (N10247, N10235);
or OR3 (N10248, N10244, N4193, N8836);
not NOT1 (N10249, N10247);
xor XOR2 (N10250, N10242, N4182);
and AND4 (N10251, N10241, N6960, N6073, N7999);
buf BUF1 (N10252, N10249);
nor NOR4 (N10253, N10248, N3042, N4760, N1670);
nand NAND4 (N10254, N10221, N5635, N2042, N5444);
not NOT1 (N10255, N10217);
or OR3 (N10256, N10251, N7389, N7509);
not NOT1 (N10257, N10243);
nand NAND2 (N10258, N10246, N8087);
buf BUF1 (N10259, N10253);
not NOT1 (N10260, N10257);
or OR2 (N10261, N10256, N2046);
nor NOR4 (N10262, N10255, N9336, N1190, N1691);
nor NOR2 (N10263, N10262, N5345);
xor XOR2 (N10264, N10239, N2826);
not NOT1 (N10265, N10261);
nand NAND3 (N10266, N10252, N6392, N6076);
nand NAND3 (N10267, N10259, N412, N10062);
and AND2 (N10268, N10266, N7485);
nand NAND2 (N10269, N10265, N8900);
xor XOR2 (N10270, N10260, N2085);
xor XOR2 (N10271, N10269, N7548);
nor NOR2 (N10272, N10263, N7484);
or OR4 (N10273, N10250, N4115, N5381, N5202);
or OR3 (N10274, N10272, N4708, N2005);
and AND2 (N10275, N10270, N8783);
nor NOR2 (N10276, N10268, N7894);
and AND3 (N10277, N10258, N5515, N1487);
nand NAND2 (N10278, N10264, N3123);
nor NOR2 (N10279, N10254, N8982);
and AND4 (N10280, N10278, N216, N7338, N10051);
xor XOR2 (N10281, N10279, N8111);
buf BUF1 (N10282, N10274);
xor XOR2 (N10283, N10281, N1401);
nor NOR4 (N10284, N10283, N7867, N1406, N8215);
or OR2 (N10285, N10276, N2888);
nand NAND4 (N10286, N10284, N649, N1246, N4304);
and AND4 (N10287, N10285, N6275, N8460, N10253);
nor NOR2 (N10288, N10271, N3782);
not NOT1 (N10289, N10280);
nor NOR3 (N10290, N10277, N8716, N9822);
nor NOR3 (N10291, N10288, N2838, N8082);
and AND4 (N10292, N10290, N3781, N6343, N2912);
nand NAND3 (N10293, N10267, N4511, N534);
and AND3 (N10294, N10286, N565, N3482);
xor XOR2 (N10295, N10292, N9659);
or OR3 (N10296, N10275, N8756, N7986);
and AND2 (N10297, N10289, N25);
nand NAND2 (N10298, N10282, N2100);
nor NOR2 (N10299, N10296, N4306);
not NOT1 (N10300, N10287);
buf BUF1 (N10301, N10300);
and AND4 (N10302, N10245, N951, N10065, N2415);
buf BUF1 (N10303, N10295);
and AND3 (N10304, N10298, N1647, N54);
nand NAND2 (N10305, N10303, N8631);
nand NAND4 (N10306, N10302, N2715, N1621, N9555);
buf BUF1 (N10307, N10273);
xor XOR2 (N10308, N10299, N800);
xor XOR2 (N10309, N10297, N3696);
nor NOR3 (N10310, N10304, N8507, N1216);
nand NAND2 (N10311, N10294, N9523);
nor NOR3 (N10312, N10310, N9645, N807);
xor XOR2 (N10313, N10309, N423);
xor XOR2 (N10314, N10312, N10295);
or OR2 (N10315, N10301, N1587);
and AND3 (N10316, N10308, N3516, N3420);
or OR4 (N10317, N10311, N6465, N9006, N3163);
buf BUF1 (N10318, N10315);
or OR3 (N10319, N10307, N4778, N1372);
or OR4 (N10320, N10314, N8573, N3032, N9838);
xor XOR2 (N10321, N10316, N1356);
nor NOR2 (N10322, N10291, N1712);
or OR3 (N10323, N10317, N5343, N5594);
buf BUF1 (N10324, N10322);
xor XOR2 (N10325, N10321, N7851);
not NOT1 (N10326, N10325);
and AND2 (N10327, N10326, N1617);
or OR2 (N10328, N10305, N4742);
xor XOR2 (N10329, N10327, N4264);
and AND4 (N10330, N10306, N6223, N202, N1590);
xor XOR2 (N10331, N10330, N6761);
not NOT1 (N10332, N10319);
nor NOR2 (N10333, N10329, N7289);
not NOT1 (N10334, N10333);
not NOT1 (N10335, N10293);
and AND2 (N10336, N10323, N1203);
or OR3 (N10337, N10335, N2383, N1926);
not NOT1 (N10338, N10331);
and AND2 (N10339, N10332, N7837);
not NOT1 (N10340, N10339);
buf BUF1 (N10341, N10334);
or OR3 (N10342, N10328, N1542, N3219);
or OR2 (N10343, N10318, N3032);
or OR4 (N10344, N10320, N23, N4855, N2504);
xor XOR2 (N10345, N10340, N2201);
nor NOR2 (N10346, N10342, N2553);
or OR2 (N10347, N10338, N3783);
and AND2 (N10348, N10347, N6987);
nor NOR4 (N10349, N10345, N10064, N3976, N1101);
nor NOR4 (N10350, N10336, N3244, N92, N6218);
xor XOR2 (N10351, N10343, N1694);
or OR2 (N10352, N10350, N3000);
or OR4 (N10353, N10351, N9208, N6131, N9354);
nor NOR4 (N10354, N10346, N3177, N10268, N6450);
nand NAND3 (N10355, N10344, N7388, N2783);
and AND4 (N10356, N10349, N2747, N1287, N5815);
xor XOR2 (N10357, N10348, N2930);
nand NAND3 (N10358, N10337, N6515, N3826);
xor XOR2 (N10359, N10358, N9911);
not NOT1 (N10360, N10359);
xor XOR2 (N10361, N10313, N3602);
and AND2 (N10362, N10357, N656);
and AND4 (N10363, N10354, N7985, N9384, N8649);
nand NAND3 (N10364, N10363, N136, N6737);
not NOT1 (N10365, N10361);
or OR2 (N10366, N10355, N1026);
and AND2 (N10367, N10356, N2029);
and AND2 (N10368, N10367, N3305);
xor XOR2 (N10369, N10368, N6409);
and AND3 (N10370, N10352, N3696, N10208);
nand NAND4 (N10371, N10362, N2287, N732, N5298);
nand NAND4 (N10372, N10369, N1733, N1678, N6478);
nand NAND2 (N10373, N10353, N10338);
buf BUF1 (N10374, N10366);
buf BUF1 (N10375, N10371);
nor NOR4 (N10376, N10373, N3049, N9287, N6201);
and AND2 (N10377, N10324, N9823);
not NOT1 (N10378, N10377);
xor XOR2 (N10379, N10374, N6668);
and AND2 (N10380, N10365, N6925);
or OR4 (N10381, N10360, N1616, N10211, N4638);
or OR2 (N10382, N10370, N1749);
nor NOR3 (N10383, N10378, N3879, N3099);
not NOT1 (N10384, N10376);
and AND2 (N10385, N10372, N3658);
and AND2 (N10386, N10379, N8937);
not NOT1 (N10387, N10364);
xor XOR2 (N10388, N10387, N3294);
xor XOR2 (N10389, N10383, N4070);
and AND4 (N10390, N10341, N4377, N7789, N7293);
not NOT1 (N10391, N10389);
or OR3 (N10392, N10385, N4631, N4219);
nor NOR2 (N10393, N10382, N5906);
nor NOR4 (N10394, N10392, N3311, N4930, N9818);
buf BUF1 (N10395, N10386);
or OR3 (N10396, N10390, N933, N658);
nand NAND3 (N10397, N10394, N9697, N8102);
nor NOR2 (N10398, N10388, N9872);
xor XOR2 (N10399, N10384, N2680);
and AND3 (N10400, N10396, N6069, N860);
nor NOR3 (N10401, N10398, N3668, N9367);
nor NOR2 (N10402, N10391, N7443);
xor XOR2 (N10403, N10400, N8067);
or OR3 (N10404, N10395, N82, N165);
xor XOR2 (N10405, N10380, N3185);
xor XOR2 (N10406, N10397, N3216);
not NOT1 (N10407, N10401);
xor XOR2 (N10408, N10407, N2296);
not NOT1 (N10409, N10393);
nor NOR3 (N10410, N10403, N5686, N6906);
not NOT1 (N10411, N10405);
buf BUF1 (N10412, N10410);
and AND3 (N10413, N10406, N7756, N5200);
nor NOR4 (N10414, N10412, N7587, N5016, N9693);
xor XOR2 (N10415, N10414, N5513);
nor NOR4 (N10416, N10415, N7050, N3975, N3999);
or OR4 (N10417, N10399, N8641, N7259, N1240);
or OR3 (N10418, N10381, N5368, N6097);
buf BUF1 (N10419, N10413);
buf BUF1 (N10420, N10409);
nand NAND4 (N10421, N10408, N1249, N10302, N8175);
not NOT1 (N10422, N10419);
and AND2 (N10423, N10411, N2719);
nand NAND2 (N10424, N10402, N5804);
nand NAND4 (N10425, N10422, N5366, N6561, N5944);
buf BUF1 (N10426, N10424);
xor XOR2 (N10427, N10404, N9536);
or OR2 (N10428, N10375, N8804);
buf BUF1 (N10429, N10421);
and AND2 (N10430, N10429, N5657);
not NOT1 (N10431, N10427);
buf BUF1 (N10432, N10428);
nor NOR4 (N10433, N10426, N331, N1627, N3404);
nor NOR3 (N10434, N10423, N7026, N5698);
nor NOR4 (N10435, N10431, N10095, N837, N1630);
xor XOR2 (N10436, N10425, N6867);
and AND4 (N10437, N10436, N92, N9708, N7108);
and AND3 (N10438, N10418, N9990, N8750);
and AND2 (N10439, N10420, N4170);
xor XOR2 (N10440, N10430, N10324);
buf BUF1 (N10441, N10432);
not NOT1 (N10442, N10435);
buf BUF1 (N10443, N10416);
and AND4 (N10444, N10417, N564, N4425, N7666);
nand NAND3 (N10445, N10434, N3423, N9496);
not NOT1 (N10446, N10441);
buf BUF1 (N10447, N10444);
nand NAND4 (N10448, N10446, N9984, N3314, N4802);
xor XOR2 (N10449, N10433, N872);
and AND4 (N10450, N10438, N2800, N6262, N6018);
not NOT1 (N10451, N10439);
nor NOR4 (N10452, N10437, N4325, N3208, N5522);
buf BUF1 (N10453, N10440);
xor XOR2 (N10454, N10450, N9259);
xor XOR2 (N10455, N10445, N3059);
xor XOR2 (N10456, N10455, N5334);
and AND2 (N10457, N10442, N7063);
not NOT1 (N10458, N10454);
nand NAND2 (N10459, N10456, N2848);
nor NOR2 (N10460, N10447, N801);
nor NOR3 (N10461, N10452, N4764, N1540);
xor XOR2 (N10462, N10459, N4861);
and AND3 (N10463, N10448, N2187, N9764);
xor XOR2 (N10464, N10453, N5572);
and AND2 (N10465, N10457, N5180);
buf BUF1 (N10466, N10463);
and AND4 (N10467, N10460, N407, N2125, N186);
nor NOR4 (N10468, N10466, N7939, N4065, N10157);
or OR2 (N10469, N10458, N2443);
nor NOR2 (N10470, N10449, N1900);
not NOT1 (N10471, N10467);
nor NOR2 (N10472, N10462, N4472);
not NOT1 (N10473, N10469);
nand NAND2 (N10474, N10470, N492);
or OR4 (N10475, N10443, N8730, N7183, N3478);
not NOT1 (N10476, N10471);
xor XOR2 (N10477, N10468, N3086);
and AND2 (N10478, N10474, N3656);
nand NAND2 (N10479, N10476, N2996);
buf BUF1 (N10480, N10465);
or OR2 (N10481, N10475, N780);
not NOT1 (N10482, N10464);
buf BUF1 (N10483, N10479);
nor NOR3 (N10484, N10480, N606, N1591);
nor NOR2 (N10485, N10482, N3143);
nor NOR4 (N10486, N10477, N8003, N462, N9313);
not NOT1 (N10487, N10461);
nand NAND3 (N10488, N10451, N6411, N7148);
not NOT1 (N10489, N10481);
not NOT1 (N10490, N10489);
and AND4 (N10491, N10472, N3132, N6536, N3743);
or OR4 (N10492, N10488, N3168, N4120, N8508);
or OR4 (N10493, N10490, N3106, N9184, N4709);
buf BUF1 (N10494, N10491);
or OR2 (N10495, N10473, N1771);
nor NOR4 (N10496, N10494, N344, N3058, N9736);
or OR4 (N10497, N10496, N1755, N5755, N10089);
and AND4 (N10498, N10483, N5689, N3458, N6289);
not NOT1 (N10499, N10486);
and AND4 (N10500, N10497, N256, N1942, N7731);
xor XOR2 (N10501, N10499, N1025);
not NOT1 (N10502, N10501);
not NOT1 (N10503, N10493);
xor XOR2 (N10504, N10498, N8443);
or OR4 (N10505, N10504, N7432, N9716, N1827);
nor NOR3 (N10506, N10500, N7752, N3239);
not NOT1 (N10507, N10492);
nor NOR2 (N10508, N10505, N1172);
buf BUF1 (N10509, N10502);
nor NOR2 (N10510, N10485, N10402);
buf BUF1 (N10511, N10509);
buf BUF1 (N10512, N10508);
and AND3 (N10513, N10511, N5577, N6384);
nor NOR3 (N10514, N10507, N6860, N10401);
nor NOR2 (N10515, N10495, N7832);
or OR2 (N10516, N10510, N3420);
and AND3 (N10517, N10506, N770, N7349);
xor XOR2 (N10518, N10478, N10326);
and AND2 (N10519, N10513, N488);
not NOT1 (N10520, N10487);
buf BUF1 (N10521, N10520);
and AND3 (N10522, N10503, N3336, N3068);
not NOT1 (N10523, N10518);
nand NAND2 (N10524, N10512, N9856);
xor XOR2 (N10525, N10514, N2661);
nand NAND3 (N10526, N10484, N3291, N4733);
nand NAND4 (N10527, N10522, N7834, N3521, N7408);
and AND4 (N10528, N10523, N1057, N9458, N778);
buf BUF1 (N10529, N10521);
not NOT1 (N10530, N10527);
nor NOR3 (N10531, N10516, N5970, N3857);
or OR2 (N10532, N10515, N5890);
buf BUF1 (N10533, N10524);
or OR3 (N10534, N10528, N5031, N9007);
or OR4 (N10535, N10531, N3801, N2247, N5817);
buf BUF1 (N10536, N10517);
or OR4 (N10537, N10532, N8518, N4084, N2844);
nor NOR4 (N10538, N10534, N2337, N1265, N7128);
nor NOR2 (N10539, N10536, N1684);
nor NOR2 (N10540, N10526, N9791);
not NOT1 (N10541, N10540);
not NOT1 (N10542, N10533);
or OR4 (N10543, N10529, N3270, N5658, N3129);
nand NAND4 (N10544, N10535, N4617, N7657, N10255);
nand NAND2 (N10545, N10539, N5622);
xor XOR2 (N10546, N10542, N7154);
nand NAND2 (N10547, N10538, N8706);
nand NAND3 (N10548, N10544, N8491, N7122);
or OR2 (N10549, N10543, N2670);
xor XOR2 (N10550, N10530, N1686);
or OR3 (N10551, N10519, N10540, N1856);
xor XOR2 (N10552, N10549, N10301);
xor XOR2 (N10553, N10525, N3495);
xor XOR2 (N10554, N10547, N6109);
nand NAND2 (N10555, N10552, N3438);
buf BUF1 (N10556, N10555);
or OR4 (N10557, N10556, N7907, N7036, N7781);
nand NAND3 (N10558, N10548, N8075, N8538);
nand NAND3 (N10559, N10545, N1732, N3757);
or OR2 (N10560, N10551, N368);
or OR3 (N10561, N10541, N7909, N9142);
buf BUF1 (N10562, N10550);
buf BUF1 (N10563, N10559);
nor NOR2 (N10564, N10553, N10014);
nor NOR4 (N10565, N10561, N5745, N6342, N8131);
and AND2 (N10566, N10562, N5488);
nand NAND3 (N10567, N10546, N9976, N10048);
nor NOR3 (N10568, N10557, N7831, N4205);
nand NAND4 (N10569, N10554, N2560, N8984, N5572);
and AND2 (N10570, N10560, N177);
or OR3 (N10571, N10564, N7109, N4591);
or OR4 (N10572, N10558, N10088, N1864, N972);
and AND3 (N10573, N10568, N1991, N5846);
nand NAND2 (N10574, N10567, N9525);
nor NOR4 (N10575, N10537, N6846, N1041, N5953);
and AND4 (N10576, N10565, N8572, N6826, N1201);
and AND2 (N10577, N10576, N3857);
xor XOR2 (N10578, N10575, N7044);
nor NOR4 (N10579, N10563, N8738, N943, N1411);
buf BUF1 (N10580, N10577);
buf BUF1 (N10581, N10579);
not NOT1 (N10582, N10573);
or OR3 (N10583, N10571, N6995, N5616);
xor XOR2 (N10584, N10583, N8584);
xor XOR2 (N10585, N10572, N8370);
and AND3 (N10586, N10569, N9559, N3046);
not NOT1 (N10587, N10570);
and AND4 (N10588, N10566, N5427, N6570, N3917);
and AND2 (N10589, N10574, N9231);
xor XOR2 (N10590, N10578, N9142);
buf BUF1 (N10591, N10582);
buf BUF1 (N10592, N10589);
nand NAND3 (N10593, N10591, N3989, N9400);
or OR3 (N10594, N10584, N5257, N3787);
buf BUF1 (N10595, N10590);
or OR2 (N10596, N10586, N1844);
buf BUF1 (N10597, N10585);
and AND3 (N10598, N10587, N8501, N4466);
buf BUF1 (N10599, N10595);
and AND4 (N10600, N10581, N10222, N10401, N6320);
nand NAND4 (N10601, N10598, N2626, N7899, N355);
and AND3 (N10602, N10599, N544, N1084);
not NOT1 (N10603, N10588);
nor NOR3 (N10604, N10596, N5135, N5179);
not NOT1 (N10605, N10600);
and AND4 (N10606, N10593, N924, N8514, N1328);
xor XOR2 (N10607, N10597, N9780);
nor NOR4 (N10608, N10592, N4159, N5023, N7059);
or OR4 (N10609, N10602, N94, N603, N8189);
or OR2 (N10610, N10608, N4057);
and AND3 (N10611, N10610, N4055, N2098);
or OR4 (N10612, N10605, N9751, N7577, N9474);
and AND3 (N10613, N10594, N383, N4015);
and AND3 (N10614, N10601, N3167, N7817);
nand NAND3 (N10615, N10606, N5287, N1748);
xor XOR2 (N10616, N10607, N8564);
buf BUF1 (N10617, N10603);
and AND4 (N10618, N10613, N2721, N8503, N10564);
buf BUF1 (N10619, N10614);
nor NOR4 (N10620, N10612, N7710, N5396, N7387);
nor NOR2 (N10621, N10617, N7992);
xor XOR2 (N10622, N10621, N7347);
nand NAND4 (N10623, N10615, N2195, N9190, N7704);
nand NAND2 (N10624, N10604, N10226);
buf BUF1 (N10625, N10580);
nor NOR2 (N10626, N10623, N4518);
not NOT1 (N10627, N10618);
not NOT1 (N10628, N10616);
not NOT1 (N10629, N10624);
and AND4 (N10630, N10626, N1453, N9953, N7084);
nor NOR3 (N10631, N10628, N6959, N2060);
nand NAND2 (N10632, N10619, N4889);
and AND4 (N10633, N10631, N8255, N4356, N876);
not NOT1 (N10634, N10633);
or OR3 (N10635, N10620, N616, N9463);
and AND2 (N10636, N10632, N2264);
nand NAND4 (N10637, N10622, N5256, N5916, N2521);
nor NOR2 (N10638, N10637, N4087);
and AND4 (N10639, N10609, N640, N3112, N8965);
or OR2 (N10640, N10638, N2060);
xor XOR2 (N10641, N10639, N6615);
buf BUF1 (N10642, N10625);
xor XOR2 (N10643, N10611, N4237);
nand NAND4 (N10644, N10643, N10329, N8558, N5123);
buf BUF1 (N10645, N10642);
and AND4 (N10646, N10634, N1629, N9121, N1694);
nand NAND2 (N10647, N10635, N9284);
xor XOR2 (N10648, N10645, N3383);
or OR2 (N10649, N10641, N8749);
and AND4 (N10650, N10636, N5302, N6939, N6708);
not NOT1 (N10651, N10640);
or OR4 (N10652, N10627, N918, N5137, N9667);
or OR2 (N10653, N10647, N5428);
nor NOR2 (N10654, N10646, N4832);
xor XOR2 (N10655, N10650, N8221);
buf BUF1 (N10656, N10652);
not NOT1 (N10657, N10653);
not NOT1 (N10658, N10649);
xor XOR2 (N10659, N10654, N10411);
nor NOR3 (N10660, N10651, N5663, N9637);
not NOT1 (N10661, N10655);
not NOT1 (N10662, N10629);
or OR4 (N10663, N10660, N5925, N1422, N7689);
buf BUF1 (N10664, N10659);
or OR2 (N10665, N10656, N5523);
nand NAND3 (N10666, N10648, N6944, N4051);
nand NAND3 (N10667, N10662, N1806, N6110);
or OR4 (N10668, N10664, N3665, N10215, N4573);
and AND3 (N10669, N10665, N3663, N8641);
not NOT1 (N10670, N10669);
or OR3 (N10671, N10658, N9290, N7534);
and AND3 (N10672, N10668, N3205, N8859);
not NOT1 (N10673, N10661);
not NOT1 (N10674, N10671);
not NOT1 (N10675, N10672);
buf BUF1 (N10676, N10675);
and AND4 (N10677, N10670, N3063, N6280, N9270);
nand NAND3 (N10678, N10667, N5631, N3550);
or OR3 (N10679, N10677, N2282, N5183);
or OR4 (N10680, N10674, N1190, N5145, N4639);
nor NOR3 (N10681, N10673, N8260, N4846);
xor XOR2 (N10682, N10663, N602);
nand NAND2 (N10683, N10681, N7216);
and AND3 (N10684, N10680, N6419, N7280);
and AND2 (N10685, N10679, N1045);
nand NAND3 (N10686, N10630, N352, N2947);
not NOT1 (N10687, N10657);
or OR3 (N10688, N10683, N10266, N2803);
xor XOR2 (N10689, N10682, N7472);
xor XOR2 (N10690, N10685, N10680);
nor NOR4 (N10691, N10678, N8280, N6525, N199);
and AND4 (N10692, N10690, N9422, N10162, N4574);
buf BUF1 (N10693, N10692);
nor NOR4 (N10694, N10689, N4861, N8577, N2548);
or OR4 (N10695, N10684, N5876, N5111, N5471);
xor XOR2 (N10696, N10666, N1359);
buf BUF1 (N10697, N10695);
nand NAND2 (N10698, N10688, N8271);
nor NOR2 (N10699, N10686, N2651);
xor XOR2 (N10700, N10687, N7417);
or OR3 (N10701, N10697, N8097, N1381);
or OR4 (N10702, N10644, N8889, N52, N2167);
nand NAND3 (N10703, N10698, N2010, N2420);
or OR2 (N10704, N10694, N2750);
nor NOR3 (N10705, N10704, N10270, N6713);
not NOT1 (N10706, N10703);
or OR2 (N10707, N10702, N7644);
nor NOR4 (N10708, N10707, N8649, N8419, N1695);
not NOT1 (N10709, N10706);
buf BUF1 (N10710, N10676);
xor XOR2 (N10711, N10705, N4713);
and AND2 (N10712, N10701, N5268);
or OR4 (N10713, N10711, N1183, N10081, N9462);
buf BUF1 (N10714, N10712);
not NOT1 (N10715, N10700);
nor NOR3 (N10716, N10709, N8626, N4181);
buf BUF1 (N10717, N10699);
and AND4 (N10718, N10696, N5824, N7383, N4208);
xor XOR2 (N10719, N10693, N8918);
or OR4 (N10720, N10691, N1605, N3007, N989);
and AND4 (N10721, N10715, N3737, N6277, N1330);
not NOT1 (N10722, N10719);
or OR4 (N10723, N10718, N1333, N8787, N5018);
nand NAND4 (N10724, N10716, N8975, N4467, N8676);
nor NOR3 (N10725, N10722, N966, N5402);
not NOT1 (N10726, N10710);
buf BUF1 (N10727, N10725);
or OR4 (N10728, N10708, N9934, N131, N9836);
xor XOR2 (N10729, N10724, N7756);
not NOT1 (N10730, N10723);
nor NOR2 (N10731, N10730, N9654);
or OR3 (N10732, N10727, N4108, N739);
buf BUF1 (N10733, N10721);
xor XOR2 (N10734, N10733, N8544);
xor XOR2 (N10735, N10729, N2946);
buf BUF1 (N10736, N10728);
buf BUF1 (N10737, N10736);
buf BUF1 (N10738, N10732);
nand NAND3 (N10739, N10726, N6534, N445);
xor XOR2 (N10740, N10735, N9363);
not NOT1 (N10741, N10720);
and AND2 (N10742, N10717, N5844);
not NOT1 (N10743, N10713);
xor XOR2 (N10744, N10739, N2700);
xor XOR2 (N10745, N10734, N10019);
not NOT1 (N10746, N10738);
not NOT1 (N10747, N10743);
xor XOR2 (N10748, N10744, N8447);
not NOT1 (N10749, N10748);
xor XOR2 (N10750, N10742, N4072);
and AND3 (N10751, N10740, N2163, N9947);
nand NAND3 (N10752, N10750, N4312, N2026);
or OR3 (N10753, N10746, N6262, N6094);
buf BUF1 (N10754, N10747);
not NOT1 (N10755, N10737);
xor XOR2 (N10756, N10755, N1594);
nand NAND4 (N10757, N10749, N2721, N1248, N4071);
nor NOR3 (N10758, N10753, N1326, N6736);
or OR3 (N10759, N10756, N878, N129);
xor XOR2 (N10760, N10745, N8178);
and AND4 (N10761, N10754, N6988, N2734, N10193);
xor XOR2 (N10762, N10751, N4350);
not NOT1 (N10763, N10741);
buf BUF1 (N10764, N10759);
nor NOR3 (N10765, N10757, N9131, N2717);
and AND4 (N10766, N10731, N3386, N9243, N3981);
not NOT1 (N10767, N10766);
xor XOR2 (N10768, N10767, N3643);
not NOT1 (N10769, N10764);
not NOT1 (N10770, N10762);
buf BUF1 (N10771, N10763);
not NOT1 (N10772, N10752);
or OR3 (N10773, N10769, N7345, N7851);
not NOT1 (N10774, N10758);
nor NOR3 (N10775, N10773, N3680, N98);
nand NAND2 (N10776, N10774, N9862);
nand NAND4 (N10777, N10765, N6389, N10381, N4319);
xor XOR2 (N10778, N10768, N5902);
nand NAND3 (N10779, N10778, N4099, N813);
and AND2 (N10780, N10771, N8858);
and AND2 (N10781, N10760, N3302);
nand NAND4 (N10782, N10772, N8780, N686, N7652);
xor XOR2 (N10783, N10761, N7763);
nand NAND2 (N10784, N10714, N2897);
nand NAND4 (N10785, N10776, N3231, N6089, N8635);
buf BUF1 (N10786, N10777);
buf BUF1 (N10787, N10784);
nor NOR2 (N10788, N10779, N7068);
buf BUF1 (N10789, N10775);
not NOT1 (N10790, N10789);
nor NOR4 (N10791, N10790, N1064, N7130, N2052);
nor NOR3 (N10792, N10785, N5425, N4426);
buf BUF1 (N10793, N10787);
and AND2 (N10794, N10786, N10308);
and AND3 (N10795, N10782, N1017, N3696);
nand NAND4 (N10796, N10781, N9243, N8474, N9687);
nor NOR2 (N10797, N10794, N9112);
xor XOR2 (N10798, N10791, N5580);
nand NAND4 (N10799, N10798, N226, N7131, N5667);
xor XOR2 (N10800, N10788, N9438);
buf BUF1 (N10801, N10795);
not NOT1 (N10802, N10799);
nor NOR3 (N10803, N10793, N4658, N10360);
buf BUF1 (N10804, N10783);
xor XOR2 (N10805, N10804, N6281);
buf BUF1 (N10806, N10770);
nand NAND2 (N10807, N10801, N8615);
nand NAND2 (N10808, N10780, N9190);
nor NOR3 (N10809, N10792, N2995, N9507);
and AND3 (N10810, N10807, N7476, N235);
xor XOR2 (N10811, N10796, N3128);
not NOT1 (N10812, N10803);
xor XOR2 (N10813, N10797, N5373);
buf BUF1 (N10814, N10811);
xor XOR2 (N10815, N10814, N8101);
or OR4 (N10816, N10800, N7827, N9777, N171);
or OR3 (N10817, N10816, N9480, N10584);
or OR4 (N10818, N10808, N8693, N7165, N5352);
nand NAND3 (N10819, N10805, N10095, N6670);
nor NOR4 (N10820, N10817, N1462, N8143, N6958);
and AND2 (N10821, N10820, N6063);
buf BUF1 (N10822, N10806);
not NOT1 (N10823, N10819);
not NOT1 (N10824, N10809);
nor NOR4 (N10825, N10810, N2275, N4922, N6631);
not NOT1 (N10826, N10802);
or OR3 (N10827, N10822, N5217, N4488);
not NOT1 (N10828, N10824);
not NOT1 (N10829, N10813);
not NOT1 (N10830, N10828);
and AND2 (N10831, N10826, N6581);
xor XOR2 (N10832, N10815, N2579);
or OR2 (N10833, N10831, N5039);
nand NAND4 (N10834, N10825, N214, N6916, N8171);
nor NOR4 (N10835, N10830, N180, N4080, N2546);
xor XOR2 (N10836, N10821, N2284);
buf BUF1 (N10837, N10836);
not NOT1 (N10838, N10812);
nand NAND2 (N10839, N10818, N979);
xor XOR2 (N10840, N10827, N380);
buf BUF1 (N10841, N10823);
not NOT1 (N10842, N10840);
or OR4 (N10843, N10838, N4743, N859, N5784);
nand NAND2 (N10844, N10842, N7647);
not NOT1 (N10845, N10843);
xor XOR2 (N10846, N10844, N4126);
not NOT1 (N10847, N10846);
or OR2 (N10848, N10835, N4324);
buf BUF1 (N10849, N10839);
or OR4 (N10850, N10845, N1292, N5267, N7285);
buf BUF1 (N10851, N10833);
and AND3 (N10852, N10848, N4260, N6622);
xor XOR2 (N10853, N10847, N9682);
not NOT1 (N10854, N10829);
not NOT1 (N10855, N10837);
or OR2 (N10856, N10832, N6008);
buf BUF1 (N10857, N10854);
nand NAND4 (N10858, N10849, N7804, N4115, N855);
or OR4 (N10859, N10850, N3981, N6568, N3924);
nand NAND4 (N10860, N10857, N5974, N4746, N658);
xor XOR2 (N10861, N10860, N2270);
nand NAND2 (N10862, N10841, N3696);
and AND4 (N10863, N10834, N1028, N7916, N5508);
or OR4 (N10864, N10862, N9105, N4951, N6064);
buf BUF1 (N10865, N10853);
buf BUF1 (N10866, N10861);
buf BUF1 (N10867, N10856);
not NOT1 (N10868, N10866);
not NOT1 (N10869, N10863);
buf BUF1 (N10870, N10868);
buf BUF1 (N10871, N10855);
and AND3 (N10872, N10852, N8371, N4369);
nand NAND3 (N10873, N10864, N7851, N9170);
and AND3 (N10874, N10865, N9492, N10369);
buf BUF1 (N10875, N10874);
not NOT1 (N10876, N10870);
buf BUF1 (N10877, N10875);
nor NOR4 (N10878, N10876, N198, N744, N7867);
nor NOR4 (N10879, N10871, N740, N4207, N7494);
buf BUF1 (N10880, N10879);
buf BUF1 (N10881, N10878);
xor XOR2 (N10882, N10851, N5165);
not NOT1 (N10883, N10880);
or OR3 (N10884, N10869, N10609, N888);
nor NOR2 (N10885, N10858, N1321);
nand NAND4 (N10886, N10881, N6794, N5468, N3445);
xor XOR2 (N10887, N10882, N6416);
nand NAND2 (N10888, N10884, N3321);
xor XOR2 (N10889, N10872, N5926);
buf BUF1 (N10890, N10859);
nand NAND4 (N10891, N10867, N7670, N5972, N529);
and AND3 (N10892, N10873, N5603, N7914);
xor XOR2 (N10893, N10887, N4949);
not NOT1 (N10894, N10877);
or OR4 (N10895, N10894, N8455, N5597, N7860);
xor XOR2 (N10896, N10885, N1336);
and AND4 (N10897, N10892, N5871, N10276, N2664);
or OR2 (N10898, N10891, N4064);
and AND3 (N10899, N10896, N2225, N7144);
nand NAND2 (N10900, N10899, N10503);
not NOT1 (N10901, N10886);
and AND2 (N10902, N10890, N7117);
nand NAND4 (N10903, N10883, N2797, N4447, N7722);
nand NAND3 (N10904, N10889, N4411, N10761);
xor XOR2 (N10905, N10900, N10173);
and AND3 (N10906, N10888, N7391, N9304);
nor NOR4 (N10907, N10903, N877, N6371, N4540);
and AND4 (N10908, N10904, N4772, N8394, N10649);
nor NOR4 (N10909, N10908, N8230, N2519, N5582);
and AND3 (N10910, N10907, N6839, N7681);
not NOT1 (N10911, N10897);
or OR2 (N10912, N10902, N9794);
xor XOR2 (N10913, N10898, N8113);
nand NAND4 (N10914, N10895, N4479, N3755, N8336);
buf BUF1 (N10915, N10914);
and AND4 (N10916, N10905, N8143, N1289, N1804);
and AND4 (N10917, N10910, N2481, N6256, N5738);
nor NOR2 (N10918, N10917, N5185);
buf BUF1 (N10919, N10918);
and AND3 (N10920, N10901, N8993, N8716);
nor NOR4 (N10921, N10909, N3978, N3134, N4222);
not NOT1 (N10922, N10915);
buf BUF1 (N10923, N10913);
or OR2 (N10924, N10916, N1985);
or OR4 (N10925, N10921, N4537, N6759, N5899);
nand NAND4 (N10926, N10925, N303, N3946, N7518);
nand NAND3 (N10927, N10919, N10521, N6050);
nand NAND3 (N10928, N10906, N8719, N9393);
nand NAND4 (N10929, N10927, N9435, N7262, N10157);
or OR2 (N10930, N10922, N2751);
or OR4 (N10931, N10920, N9630, N5882, N735);
or OR2 (N10932, N10931, N2671);
nor NOR4 (N10933, N10924, N10842, N2040, N7291);
nand NAND2 (N10934, N10923, N2137);
not NOT1 (N10935, N10929);
nor NOR3 (N10936, N10893, N6671, N83);
or OR4 (N10937, N10932, N2363, N10608, N9976);
not NOT1 (N10938, N10937);
buf BUF1 (N10939, N10928);
or OR3 (N10940, N10939, N2339, N9313);
nand NAND3 (N10941, N10940, N733, N3996);
xor XOR2 (N10942, N10936, N3692);
nor NOR3 (N10943, N10930, N4981, N7756);
nor NOR3 (N10944, N10911, N3270, N5065);
xor XOR2 (N10945, N10935, N1517);
or OR2 (N10946, N10934, N860);
not NOT1 (N10947, N10926);
nor NOR2 (N10948, N10912, N5879);
xor XOR2 (N10949, N10942, N556);
and AND3 (N10950, N10946, N955, N10631);
xor XOR2 (N10951, N10945, N1703);
buf BUF1 (N10952, N10938);
xor XOR2 (N10953, N10950, N549);
and AND2 (N10954, N10951, N8501);
or OR2 (N10955, N10949, N9101);
and AND2 (N10956, N10955, N3346);
or OR2 (N10957, N10933, N5010);
not NOT1 (N10958, N10956);
buf BUF1 (N10959, N10944);
xor XOR2 (N10960, N10947, N1010);
and AND3 (N10961, N10948, N7497, N10608);
nand NAND2 (N10962, N10957, N9680);
or OR3 (N10963, N10941, N8058, N2484);
nand NAND3 (N10964, N10959, N6554, N6806);
buf BUF1 (N10965, N10960);
not NOT1 (N10966, N10958);
nand NAND2 (N10967, N10952, N3716);
buf BUF1 (N10968, N10962);
and AND2 (N10969, N10943, N10161);
buf BUF1 (N10970, N10953);
nor NOR4 (N10971, N10970, N4743, N1825, N388);
nor NOR4 (N10972, N10963, N3024, N5711, N10042);
buf BUF1 (N10973, N10964);
or OR4 (N10974, N10954, N520, N9388, N5938);
not NOT1 (N10975, N10965);
buf BUF1 (N10976, N10971);
buf BUF1 (N10977, N10961);
nor NOR2 (N10978, N10972, N601);
nor NOR4 (N10979, N10968, N6151, N2970, N8161);
not NOT1 (N10980, N10967);
or OR4 (N10981, N10976, N5008, N4716, N1102);
or OR2 (N10982, N10978, N4170);
not NOT1 (N10983, N10973);
nand NAND3 (N10984, N10974, N9153, N3985);
buf BUF1 (N10985, N10975);
not NOT1 (N10986, N10980);
xor XOR2 (N10987, N10981, N3367);
or OR3 (N10988, N10985, N8645, N10616);
nor NOR4 (N10989, N10988, N6264, N2291, N1620);
and AND3 (N10990, N10966, N9731, N1243);
or OR4 (N10991, N10989, N6882, N4719, N3162);
or OR2 (N10992, N10979, N8180);
or OR4 (N10993, N10990, N1536, N1464, N6677);
not NOT1 (N10994, N10983);
not NOT1 (N10995, N10994);
and AND4 (N10996, N10986, N7810, N6341, N2017);
buf BUF1 (N10997, N10993);
nand NAND2 (N10998, N10984, N6190);
and AND4 (N10999, N10987, N723, N7391, N3311);
xor XOR2 (N11000, N10969, N1159);
nand NAND3 (N11001, N10982, N3771, N8080);
and AND4 (N11002, N10997, N2858, N5457, N9919);
nand NAND2 (N11003, N10991, N9200);
xor XOR2 (N11004, N10995, N864);
nor NOR4 (N11005, N11000, N496, N9485, N378);
and AND3 (N11006, N10992, N6097, N7409);
and AND3 (N11007, N11004, N8063, N1650);
and AND4 (N11008, N10977, N8133, N10034, N4268);
buf BUF1 (N11009, N11007);
or OR3 (N11010, N10999, N9938, N7878);
nor NOR2 (N11011, N11003, N6055);
xor XOR2 (N11012, N11005, N8715);
nor NOR4 (N11013, N11006, N9525, N1847, N7968);
not NOT1 (N11014, N11013);
and AND4 (N11015, N11010, N3212, N4715, N5443);
not NOT1 (N11016, N10996);
xor XOR2 (N11017, N11001, N1182);
and AND4 (N11018, N11002, N7816, N6629, N4605);
not NOT1 (N11019, N11018);
not NOT1 (N11020, N10998);
xor XOR2 (N11021, N11009, N491);
nand NAND4 (N11022, N11008, N6986, N1474, N1241);
nand NAND2 (N11023, N11022, N8741);
nor NOR4 (N11024, N11017, N1878, N10929, N3912);
and AND4 (N11025, N11014, N123, N9209, N2867);
xor XOR2 (N11026, N11021, N10968);
nor NOR3 (N11027, N11012, N735, N7787);
and AND4 (N11028, N11020, N7584, N7403, N5170);
and AND2 (N11029, N11016, N5894);
nor NOR2 (N11030, N11024, N4916);
and AND3 (N11031, N11025, N4471, N5858);
buf BUF1 (N11032, N11031);
nor NOR2 (N11033, N11019, N9549);
xor XOR2 (N11034, N11028, N927);
buf BUF1 (N11035, N11027);
nand NAND3 (N11036, N11034, N2146, N5233);
and AND4 (N11037, N11032, N4839, N6694, N1311);
nand NAND3 (N11038, N11030, N1600, N3610);
buf BUF1 (N11039, N11026);
nand NAND2 (N11040, N11039, N1376);
not NOT1 (N11041, N11035);
nor NOR2 (N11042, N11029, N5088);
or OR2 (N11043, N11036, N7506);
nand NAND4 (N11044, N11040, N5647, N2246, N7296);
or OR2 (N11045, N11023, N464);
not NOT1 (N11046, N11015);
nand NAND3 (N11047, N11033, N5807, N7694);
xor XOR2 (N11048, N11011, N5126);
nor NOR2 (N11049, N11048, N2053);
nor NOR2 (N11050, N11038, N8963);
or OR3 (N11051, N11049, N6183, N8081);
and AND2 (N11052, N11037, N1547);
nor NOR3 (N11053, N11051, N3671, N684);
buf BUF1 (N11054, N11042);
nor NOR3 (N11055, N11041, N8178, N6628);
and AND4 (N11056, N11052, N3602, N925, N9369);
xor XOR2 (N11057, N11053, N9471);
or OR2 (N11058, N11045, N10261);
and AND2 (N11059, N11055, N10314);
nand NAND2 (N11060, N11044, N6392);
or OR2 (N11061, N11058, N6485);
xor XOR2 (N11062, N11050, N507);
not NOT1 (N11063, N11062);
xor XOR2 (N11064, N11063, N10361);
xor XOR2 (N11065, N11057, N2152);
nand NAND3 (N11066, N11061, N6394, N4191);
not NOT1 (N11067, N11059);
not NOT1 (N11068, N11056);
and AND2 (N11069, N11047, N8512);
nor NOR2 (N11070, N11068, N8495);
buf BUF1 (N11071, N11054);
nor NOR3 (N11072, N11046, N2048, N9936);
xor XOR2 (N11073, N11069, N1997);
xor XOR2 (N11074, N11067, N9536);
and AND3 (N11075, N11071, N10941, N4065);
nor NOR2 (N11076, N11065, N997);
and AND3 (N11077, N11070, N2733, N3356);
nor NOR3 (N11078, N11064, N1708, N7324);
nand NAND3 (N11079, N11066, N4797, N2159);
nor NOR2 (N11080, N11076, N2973);
and AND4 (N11081, N11078, N6658, N3245, N6234);
not NOT1 (N11082, N11079);
and AND2 (N11083, N11072, N5357);
nor NOR2 (N11084, N11074, N5345);
nor NOR3 (N11085, N11084, N9693, N5046);
xor XOR2 (N11086, N11085, N10811);
not NOT1 (N11087, N11043);
xor XOR2 (N11088, N11086, N5160);
xor XOR2 (N11089, N11060, N6798);
nor NOR4 (N11090, N11075, N6492, N3198, N274);
not NOT1 (N11091, N11089);
buf BUF1 (N11092, N11088);
buf BUF1 (N11093, N11077);
xor XOR2 (N11094, N11081, N8558);
not NOT1 (N11095, N11093);
and AND3 (N11096, N11092, N2293, N6510);
not NOT1 (N11097, N11094);
buf BUF1 (N11098, N11091);
nand NAND4 (N11099, N11073, N892, N915, N9068);
or OR4 (N11100, N11090, N6972, N5763, N7684);
buf BUF1 (N11101, N11082);
xor XOR2 (N11102, N11098, N7075);
nor NOR3 (N11103, N11100, N2793, N1763);
buf BUF1 (N11104, N11087);
buf BUF1 (N11105, N11103);
buf BUF1 (N11106, N11104);
or OR3 (N11107, N11101, N4326, N7670);
or OR4 (N11108, N11102, N4888, N10307, N57);
and AND3 (N11109, N11095, N3778, N10630);
or OR2 (N11110, N11099, N10503);
buf BUF1 (N11111, N11110);
buf BUF1 (N11112, N11097);
not NOT1 (N11113, N11083);
or OR3 (N11114, N11106, N10443, N2611);
nor NOR2 (N11115, N11111, N6739);
buf BUF1 (N11116, N11108);
or OR4 (N11117, N11114, N5522, N6414, N6853);
nand NAND4 (N11118, N11107, N6557, N4428, N3879);
not NOT1 (N11119, N11116);
buf BUF1 (N11120, N11113);
nor NOR2 (N11121, N11080, N3850);
xor XOR2 (N11122, N11117, N1244);
xor XOR2 (N11123, N11119, N7826);
and AND3 (N11124, N11120, N2143, N8733);
nand NAND2 (N11125, N11105, N4939);
xor XOR2 (N11126, N11121, N8045);
nor NOR3 (N11127, N11125, N5922, N7659);
or OR2 (N11128, N11123, N560);
or OR4 (N11129, N11112, N2016, N7881, N3048);
and AND4 (N11130, N11109, N1609, N1927, N3030);
nand NAND2 (N11131, N11096, N4546);
xor XOR2 (N11132, N11129, N636);
or OR2 (N11133, N11132, N1898);
nand NAND3 (N11134, N11124, N8350, N4449);
or OR4 (N11135, N11127, N1151, N1491, N5422);
xor XOR2 (N11136, N11135, N1489);
xor XOR2 (N11137, N11134, N8196);
and AND4 (N11138, N11133, N4624, N1332, N4614);
nor NOR3 (N11139, N11122, N10074, N9597);
or OR2 (N11140, N11139, N5353);
or OR3 (N11141, N11115, N6342, N7277);
not NOT1 (N11142, N11128);
not NOT1 (N11143, N11138);
nor NOR2 (N11144, N11141, N3850);
buf BUF1 (N11145, N11144);
or OR2 (N11146, N11143, N5184);
and AND3 (N11147, N11136, N8557, N2875);
nand NAND4 (N11148, N11130, N6732, N7182, N7931);
xor XOR2 (N11149, N11137, N6317);
or OR4 (N11150, N11140, N8436, N1908, N5692);
not NOT1 (N11151, N11145);
nor NOR4 (N11152, N11147, N1216, N5683, N781);
nand NAND3 (N11153, N11118, N8415, N9346);
and AND2 (N11154, N11149, N2389);
nor NOR4 (N11155, N11150, N652, N4865, N2306);
or OR3 (N11156, N11142, N9829, N493);
and AND3 (N11157, N11148, N11006, N4874);
xor XOR2 (N11158, N11156, N1904);
xor XOR2 (N11159, N11155, N7381);
not NOT1 (N11160, N11158);
nand NAND4 (N11161, N11153, N4699, N10598, N4395);
xor XOR2 (N11162, N11159, N1189);
buf BUF1 (N11163, N11162);
nand NAND2 (N11164, N11160, N5126);
and AND2 (N11165, N11157, N1221);
or OR3 (N11166, N11161, N954, N10877);
and AND4 (N11167, N11163, N4480, N3646, N8530);
buf BUF1 (N11168, N11152);
buf BUF1 (N11169, N11146);
xor XOR2 (N11170, N11164, N10804);
buf BUF1 (N11171, N11166);
or OR4 (N11172, N11151, N5207, N9855, N1823);
or OR4 (N11173, N11168, N3793, N9408, N5667);
and AND2 (N11174, N11170, N7839);
nor NOR4 (N11175, N11172, N8368, N3779, N1822);
or OR4 (N11176, N11175, N10000, N5747, N258);
and AND2 (N11177, N11165, N4907);
buf BUF1 (N11178, N11173);
nor NOR2 (N11179, N11176, N5099);
xor XOR2 (N11180, N11154, N7005);
and AND3 (N11181, N11126, N9563, N1850);
not NOT1 (N11182, N11174);
nand NAND3 (N11183, N11131, N8197, N8126);
or OR4 (N11184, N11177, N5527, N2199, N10786);
buf BUF1 (N11185, N11182);
xor XOR2 (N11186, N11181, N4377);
not NOT1 (N11187, N11179);
buf BUF1 (N11188, N11187);
or OR2 (N11189, N11188, N7679);
not NOT1 (N11190, N11186);
nor NOR4 (N11191, N11183, N9802, N5333, N1123);
nand NAND4 (N11192, N11169, N5401, N948, N6991);
nor NOR3 (N11193, N11192, N7910, N9151);
buf BUF1 (N11194, N11178);
not NOT1 (N11195, N11185);
xor XOR2 (N11196, N11191, N8050);
and AND3 (N11197, N11184, N2188, N4082);
xor XOR2 (N11198, N11167, N5093);
and AND4 (N11199, N11190, N6552, N544, N2876);
nand NAND3 (N11200, N11197, N2269, N1559);
or OR4 (N11201, N11171, N4997, N9156, N438);
and AND2 (N11202, N11201, N6334);
buf BUF1 (N11203, N11195);
buf BUF1 (N11204, N11200);
or OR4 (N11205, N11198, N4963, N2841, N926);
nor NOR2 (N11206, N11180, N4774);
or OR2 (N11207, N11193, N6109);
and AND4 (N11208, N11202, N3151, N245, N8690);
buf BUF1 (N11209, N11205);
buf BUF1 (N11210, N11199);
or OR3 (N11211, N11207, N7482, N1950);
or OR4 (N11212, N11206, N3716, N10578, N6812);
buf BUF1 (N11213, N11194);
xor XOR2 (N11214, N11213, N1611);
or OR2 (N11215, N11196, N6164);
or OR2 (N11216, N11209, N10471);
not NOT1 (N11217, N11216);
xor XOR2 (N11218, N11203, N7683);
not NOT1 (N11219, N11217);
not NOT1 (N11220, N11210);
nor NOR4 (N11221, N11208, N11141, N7678, N3190);
nand NAND3 (N11222, N11214, N6535, N2132);
or OR2 (N11223, N11219, N9546);
and AND2 (N11224, N11220, N3103);
or OR2 (N11225, N11224, N629);
nand NAND3 (N11226, N11212, N2266, N8789);
buf BUF1 (N11227, N11222);
not NOT1 (N11228, N11227);
and AND2 (N11229, N11226, N2281);
and AND2 (N11230, N11204, N6345);
xor XOR2 (N11231, N11223, N9158);
nand NAND4 (N11232, N11229, N3487, N5018, N8329);
nand NAND4 (N11233, N11189, N1420, N3136, N10934);
and AND4 (N11234, N11231, N4276, N6888, N9218);
nor NOR4 (N11235, N11221, N675, N1678, N1436);
nand NAND3 (N11236, N11211, N26, N2325);
nand NAND4 (N11237, N11228, N2920, N9640, N6299);
nor NOR4 (N11238, N11236, N10443, N7234, N2531);
nand NAND2 (N11239, N11237, N6322);
not NOT1 (N11240, N11215);
xor XOR2 (N11241, N11232, N3636);
nor NOR3 (N11242, N11235, N8793, N2463);
or OR4 (N11243, N11230, N8097, N5233, N5419);
nor NOR3 (N11244, N11241, N8837, N456);
or OR3 (N11245, N11225, N4907, N9167);
or OR4 (N11246, N11234, N3341, N3608, N862);
not NOT1 (N11247, N11244);
nor NOR3 (N11248, N11240, N5079, N436);
and AND4 (N11249, N11238, N9760, N1637, N8726);
nand NAND2 (N11250, N11246, N10467);
and AND3 (N11251, N11242, N8226, N4871);
nor NOR2 (N11252, N11239, N1437);
and AND3 (N11253, N11243, N6555, N660);
buf BUF1 (N11254, N11245);
nor NOR3 (N11255, N11248, N3364, N282);
nand NAND4 (N11256, N11249, N6235, N9523, N8737);
or OR3 (N11257, N11252, N3416, N3252);
not NOT1 (N11258, N11257);
nor NOR2 (N11259, N11255, N2908);
nand NAND3 (N11260, N11253, N7422, N5091);
or OR4 (N11261, N11258, N4981, N3442, N2572);
xor XOR2 (N11262, N11254, N8216);
and AND4 (N11263, N11218, N7738, N7629, N9205);
nand NAND3 (N11264, N11233, N3506, N4769);
not NOT1 (N11265, N11261);
not NOT1 (N11266, N11259);
buf BUF1 (N11267, N11262);
or OR4 (N11268, N11265, N622, N8789, N7354);
not NOT1 (N11269, N11260);
buf BUF1 (N11270, N11264);
buf BUF1 (N11271, N11269);
nand NAND3 (N11272, N11271, N1032, N11125);
xor XOR2 (N11273, N11270, N8682);
not NOT1 (N11274, N11268);
not NOT1 (N11275, N11256);
and AND2 (N11276, N11247, N2804);
not NOT1 (N11277, N11263);
nand NAND4 (N11278, N11251, N106, N5998, N4189);
nand NAND4 (N11279, N11275, N6622, N6830, N2695);
nor NOR4 (N11280, N11278, N5269, N2585, N520);
not NOT1 (N11281, N11250);
nor NOR2 (N11282, N11276, N3649);
buf BUF1 (N11283, N11279);
not NOT1 (N11284, N11273);
xor XOR2 (N11285, N11274, N9123);
and AND3 (N11286, N11281, N9977, N2407);
not NOT1 (N11287, N11284);
xor XOR2 (N11288, N11282, N4410);
nand NAND2 (N11289, N11277, N6188);
xor XOR2 (N11290, N11288, N10853);
buf BUF1 (N11291, N11290);
not NOT1 (N11292, N11289);
and AND2 (N11293, N11291, N2915);
nor NOR2 (N11294, N11286, N1236);
nor NOR4 (N11295, N11294, N3643, N949, N3359);
not NOT1 (N11296, N11287);
nor NOR2 (N11297, N11272, N5056);
nor NOR2 (N11298, N11295, N8881);
nor NOR3 (N11299, N11298, N5231, N454);
or OR3 (N11300, N11285, N432, N5523);
nand NAND3 (N11301, N11300, N7947, N2240);
nor NOR4 (N11302, N11297, N4204, N2442, N1406);
and AND4 (N11303, N11296, N10636, N8833, N3107);
and AND2 (N11304, N11293, N5674);
nand NAND4 (N11305, N11266, N971, N1053, N6702);
not NOT1 (N11306, N11305);
not NOT1 (N11307, N11280);
and AND4 (N11308, N11301, N9529, N3550, N1335);
not NOT1 (N11309, N11267);
nor NOR2 (N11310, N11303, N8098);
not NOT1 (N11311, N11306);
not NOT1 (N11312, N11310);
nor NOR3 (N11313, N11302, N9510, N1478);
nor NOR2 (N11314, N11283, N9773);
xor XOR2 (N11315, N11292, N5175);
buf BUF1 (N11316, N11315);
nand NAND2 (N11317, N11304, N8609);
buf BUF1 (N11318, N11309);
nor NOR3 (N11319, N11299, N3324, N2387);
nand NAND3 (N11320, N11311, N7683, N5525);
xor XOR2 (N11321, N11314, N1517);
xor XOR2 (N11322, N11316, N1719);
not NOT1 (N11323, N11322);
nor NOR2 (N11324, N11317, N538);
and AND2 (N11325, N11321, N6164);
xor XOR2 (N11326, N11318, N5776);
buf BUF1 (N11327, N11323);
or OR3 (N11328, N11326, N6212, N1379);
nand NAND3 (N11329, N11325, N380, N7613);
or OR4 (N11330, N11308, N562, N10277, N737);
nand NAND4 (N11331, N11307, N10915, N2380, N6528);
nand NAND4 (N11332, N11313, N8594, N341, N7099);
not NOT1 (N11333, N11319);
nor NOR2 (N11334, N11327, N6416);
xor XOR2 (N11335, N11332, N4566);
nand NAND4 (N11336, N11320, N1397, N8618, N3853);
not NOT1 (N11337, N11312);
nor NOR4 (N11338, N11331, N7225, N8539, N6720);
buf BUF1 (N11339, N11333);
nor NOR4 (N11340, N11334, N3898, N2104, N9445);
not NOT1 (N11341, N11330);
buf BUF1 (N11342, N11338);
nand NAND2 (N11343, N11340, N6706);
xor XOR2 (N11344, N11342, N6012);
or OR3 (N11345, N11336, N8417, N6037);
and AND3 (N11346, N11344, N6573, N5083);
or OR3 (N11347, N11345, N2222, N7660);
buf BUF1 (N11348, N11346);
nand NAND3 (N11349, N11328, N3487, N6031);
or OR2 (N11350, N11329, N312);
nand NAND2 (N11351, N11324, N1544);
not NOT1 (N11352, N11339);
nand NAND3 (N11353, N11352, N5654, N5745);
not NOT1 (N11354, N11343);
or OR4 (N11355, N11337, N7275, N356, N4341);
and AND2 (N11356, N11354, N2116);
buf BUF1 (N11357, N11347);
buf BUF1 (N11358, N11349);
nand NAND3 (N11359, N11357, N8924, N168);
not NOT1 (N11360, N11350);
not NOT1 (N11361, N11360);
xor XOR2 (N11362, N11335, N734);
not NOT1 (N11363, N11361);
nor NOR2 (N11364, N11359, N6927);
buf BUF1 (N11365, N11353);
and AND2 (N11366, N11363, N6918);
not NOT1 (N11367, N11362);
or OR4 (N11368, N11364, N6865, N9466, N9884);
and AND2 (N11369, N11351, N1985);
or OR2 (N11370, N11367, N1921);
nand NAND4 (N11371, N11355, N7873, N1593, N5);
xor XOR2 (N11372, N11341, N7971);
nand NAND3 (N11373, N11366, N8927, N8080);
nor NOR3 (N11374, N11368, N6781, N7844);
nor NOR2 (N11375, N11371, N1408);
xor XOR2 (N11376, N11369, N6964);
not NOT1 (N11377, N11372);
and AND3 (N11378, N11377, N2982, N11059);
and AND4 (N11379, N11374, N10454, N2903, N6295);
and AND3 (N11380, N11356, N10502, N2802);
buf BUF1 (N11381, N11380);
nand NAND4 (N11382, N11376, N146, N1049, N6238);
buf BUF1 (N11383, N11375);
nand NAND4 (N11384, N11382, N10035, N2892, N2917);
nor NOR2 (N11385, N11365, N768);
nor NOR4 (N11386, N11381, N10789, N10184, N5576);
and AND2 (N11387, N11379, N10332);
or OR2 (N11388, N11385, N2669);
or OR4 (N11389, N11378, N5579, N9256, N10099);
buf BUF1 (N11390, N11387);
nor NOR3 (N11391, N11348, N11329, N3759);
or OR3 (N11392, N11370, N7751, N7298);
not NOT1 (N11393, N11386);
and AND2 (N11394, N11391, N2285);
not NOT1 (N11395, N11358);
nand NAND4 (N11396, N11390, N3182, N6881, N9852);
nand NAND2 (N11397, N11393, N11068);
buf BUF1 (N11398, N11395);
nor NOR2 (N11399, N11389, N11012);
nand NAND4 (N11400, N11394, N3690, N2401, N3664);
or OR4 (N11401, N11397, N2690, N8629, N1031);
not NOT1 (N11402, N11383);
and AND2 (N11403, N11388, N7088);
or OR2 (N11404, N11396, N10033);
xor XOR2 (N11405, N11384, N7886);
buf BUF1 (N11406, N11405);
and AND3 (N11407, N11373, N1949, N9245);
nor NOR2 (N11408, N11392, N7307);
or OR3 (N11409, N11407, N9094, N4901);
nor NOR4 (N11410, N11400, N4864, N1438, N5211);
buf BUF1 (N11411, N11399);
not NOT1 (N11412, N11404);
xor XOR2 (N11413, N11403, N10174);
nor NOR2 (N11414, N11402, N3722);
nand NAND4 (N11415, N11414, N8986, N8755, N344);
buf BUF1 (N11416, N11398);
nand NAND2 (N11417, N11415, N7950);
xor XOR2 (N11418, N11401, N9402);
nand NAND3 (N11419, N11412, N1544, N8327);
buf BUF1 (N11420, N11417);
buf BUF1 (N11421, N11411);
buf BUF1 (N11422, N11406);
not NOT1 (N11423, N11418);
nand NAND3 (N11424, N11421, N3882, N3);
buf BUF1 (N11425, N11413);
xor XOR2 (N11426, N11409, N10909);
buf BUF1 (N11427, N11416);
and AND2 (N11428, N11425, N2922);
xor XOR2 (N11429, N11424, N1846);
nand NAND3 (N11430, N11427, N8292, N2884);
buf BUF1 (N11431, N11410);
xor XOR2 (N11432, N11422, N5478);
not NOT1 (N11433, N11432);
nor NOR2 (N11434, N11431, N6740);
and AND2 (N11435, N11423, N5472);
nor NOR2 (N11436, N11429, N8456);
xor XOR2 (N11437, N11430, N3712);
xor XOR2 (N11438, N11435, N1972);
nand NAND2 (N11439, N11428, N8420);
and AND2 (N11440, N11434, N1031);
and AND2 (N11441, N11440, N3135);
buf BUF1 (N11442, N11419);
not NOT1 (N11443, N11436);
or OR2 (N11444, N11437, N10772);
buf BUF1 (N11445, N11433);
nor NOR2 (N11446, N11426, N5854);
and AND3 (N11447, N11408, N796, N7663);
not NOT1 (N11448, N11446);
nor NOR3 (N11449, N11444, N8410, N60);
nand NAND3 (N11450, N11448, N531, N8176);
or OR2 (N11451, N11439, N7949);
nand NAND4 (N11452, N11420, N8715, N7305, N9673);
xor XOR2 (N11453, N11449, N3688);
or OR4 (N11454, N11438, N309, N4180, N7315);
buf BUF1 (N11455, N11445);
nor NOR2 (N11456, N11442, N6250);
buf BUF1 (N11457, N11447);
buf BUF1 (N11458, N11455);
not NOT1 (N11459, N11452);
or OR4 (N11460, N11454, N5169, N9728, N10833);
xor XOR2 (N11461, N11450, N3955);
nor NOR2 (N11462, N11460, N9769);
buf BUF1 (N11463, N11453);
not NOT1 (N11464, N11441);
nor NOR3 (N11465, N11464, N6737, N7253);
and AND2 (N11466, N11451, N9854);
or OR3 (N11467, N11461, N11157, N7688);
buf BUF1 (N11468, N11457);
nor NOR2 (N11469, N11467, N7242);
xor XOR2 (N11470, N11469, N3554);
or OR2 (N11471, N11463, N7073);
xor XOR2 (N11472, N11459, N5255);
buf BUF1 (N11473, N11443);
buf BUF1 (N11474, N11473);
xor XOR2 (N11475, N11462, N2839);
not NOT1 (N11476, N11470);
and AND3 (N11477, N11475, N5890, N10802);
and AND2 (N11478, N11474, N202);
and AND2 (N11479, N11472, N7834);
or OR4 (N11480, N11458, N9187, N7871, N3749);
buf BUF1 (N11481, N11466);
or OR3 (N11482, N11479, N11111, N504);
not NOT1 (N11483, N11478);
nand NAND3 (N11484, N11465, N9815, N10900);
buf BUF1 (N11485, N11481);
nand NAND2 (N11486, N11476, N777);
not NOT1 (N11487, N11485);
nor NOR2 (N11488, N11484, N6216);
xor XOR2 (N11489, N11482, N5195);
nand NAND3 (N11490, N11488, N7205, N3383);
nor NOR4 (N11491, N11490, N153, N8627, N1728);
not NOT1 (N11492, N11491);
and AND4 (N11493, N11489, N2381, N5491, N6783);
buf BUF1 (N11494, N11480);
buf BUF1 (N11495, N11456);
buf BUF1 (N11496, N11492);
buf BUF1 (N11497, N11468);
xor XOR2 (N11498, N11487, N8266);
or OR2 (N11499, N11494, N11012);
not NOT1 (N11500, N11497);
buf BUF1 (N11501, N11498);
xor XOR2 (N11502, N11499, N2146);
buf BUF1 (N11503, N11471);
or OR2 (N11504, N11486, N1343);
buf BUF1 (N11505, N11477);
not NOT1 (N11506, N11503);
buf BUF1 (N11507, N11496);
buf BUF1 (N11508, N11500);
or OR3 (N11509, N11506, N8343, N237);
and AND2 (N11510, N11502, N11366);
nand NAND4 (N11511, N11493, N3835, N8390, N6516);
not NOT1 (N11512, N11509);
and AND3 (N11513, N11501, N7902, N11487);
buf BUF1 (N11514, N11483);
nand NAND2 (N11515, N11504, N10281);
and AND4 (N11516, N11511, N9624, N9010, N6619);
xor XOR2 (N11517, N11508, N9578);
and AND3 (N11518, N11513, N6606, N9655);
nand NAND3 (N11519, N11517, N2406, N2220);
xor XOR2 (N11520, N11510, N11424);
xor XOR2 (N11521, N11520, N1680);
nand NAND4 (N11522, N11514, N7074, N1513, N3189);
buf BUF1 (N11523, N11521);
nor NOR2 (N11524, N11507, N8222);
buf BUF1 (N11525, N11505);
not NOT1 (N11526, N11512);
and AND2 (N11527, N11525, N4240);
xor XOR2 (N11528, N11523, N10192);
or OR2 (N11529, N11515, N7014);
and AND2 (N11530, N11524, N6644);
nand NAND3 (N11531, N11516, N846, N6994);
and AND4 (N11532, N11527, N891, N9702, N5683);
buf BUF1 (N11533, N11519);
xor XOR2 (N11534, N11528, N4423);
not NOT1 (N11535, N11533);
nor NOR3 (N11536, N11532, N453, N5136);
xor XOR2 (N11537, N11536, N769);
nor NOR2 (N11538, N11526, N7191);
buf BUF1 (N11539, N11538);
and AND3 (N11540, N11534, N1374, N10241);
nor NOR4 (N11541, N11530, N7861, N8673, N10923);
nor NOR4 (N11542, N11522, N3621, N4659, N2334);
nor NOR4 (N11543, N11537, N8378, N6440, N2532);
nor NOR2 (N11544, N11495, N5353);
and AND2 (N11545, N11535, N9392);
not NOT1 (N11546, N11540);
nand NAND4 (N11547, N11546, N9432, N3750, N3236);
and AND3 (N11548, N11542, N600, N609);
nor NOR3 (N11549, N11529, N10582, N6857);
and AND3 (N11550, N11544, N11192, N6814);
or OR4 (N11551, N11541, N10001, N7552, N7285);
nor NOR3 (N11552, N11545, N1710, N296);
xor XOR2 (N11553, N11518, N2328);
and AND4 (N11554, N11550, N4919, N1865, N7096);
not NOT1 (N11555, N11543);
nand NAND4 (N11556, N11548, N6858, N8970, N10622);
nor NOR4 (N11557, N11552, N293, N10394, N1623);
not NOT1 (N11558, N11549);
xor XOR2 (N11559, N11553, N540);
nor NOR3 (N11560, N11547, N3857, N10258);
buf BUF1 (N11561, N11558);
buf BUF1 (N11562, N11554);
or OR3 (N11563, N11557, N9070, N2358);
nand NAND2 (N11564, N11559, N9539);
buf BUF1 (N11565, N11555);
nor NOR3 (N11566, N11531, N10428, N8599);
not NOT1 (N11567, N11561);
nand NAND3 (N11568, N11563, N6866, N4353);
buf BUF1 (N11569, N11539);
nand NAND2 (N11570, N11556, N1098);
not NOT1 (N11571, N11562);
or OR4 (N11572, N11571, N2717, N312, N2622);
xor XOR2 (N11573, N11565, N10777);
and AND3 (N11574, N11570, N8098, N76);
xor XOR2 (N11575, N11566, N8544);
not NOT1 (N11576, N11572);
xor XOR2 (N11577, N11560, N404);
nand NAND4 (N11578, N11567, N9699, N7037, N7269);
or OR3 (N11579, N11569, N1125, N8522);
and AND4 (N11580, N11577, N4858, N5704, N499);
buf BUF1 (N11581, N11564);
nor NOR2 (N11582, N11580, N8837);
or OR4 (N11583, N11551, N2387, N63, N5961);
or OR2 (N11584, N11576, N11275);
and AND2 (N11585, N11583, N8201);
nand NAND2 (N11586, N11585, N3037);
buf BUF1 (N11587, N11573);
buf BUF1 (N11588, N11579);
nor NOR3 (N11589, N11586, N4671, N1005);
or OR4 (N11590, N11578, N9871, N7879, N629);
nor NOR3 (N11591, N11588, N8029, N1688);
xor XOR2 (N11592, N11587, N11134);
or OR2 (N11593, N11582, N124);
not NOT1 (N11594, N11591);
nand NAND2 (N11595, N11594, N9598);
xor XOR2 (N11596, N11574, N2968);
not NOT1 (N11597, N11581);
nand NAND2 (N11598, N11592, N1862);
nor NOR2 (N11599, N11595, N9153);
or OR2 (N11600, N11584, N8826);
buf BUF1 (N11601, N11568);
xor XOR2 (N11602, N11599, N648);
xor XOR2 (N11603, N11596, N2955);
not NOT1 (N11604, N11603);
buf BUF1 (N11605, N11590);
nor NOR3 (N11606, N11604, N10941, N8565);
and AND3 (N11607, N11601, N9393, N6686);
nor NOR4 (N11608, N11600, N11380, N2377, N6337);
nand NAND3 (N11609, N11602, N2031, N2626);
not NOT1 (N11610, N11597);
nand NAND4 (N11611, N11598, N9731, N1029, N10288);
not NOT1 (N11612, N11589);
not NOT1 (N11613, N11593);
and AND3 (N11614, N11612, N11445, N9864);
not NOT1 (N11615, N11606);
nand NAND3 (N11616, N11607, N11147, N7864);
or OR4 (N11617, N11611, N11252, N11239, N9597);
and AND4 (N11618, N11615, N788, N1116, N4827);
nand NAND4 (N11619, N11618, N5039, N9964, N2751);
or OR3 (N11620, N11575, N7640, N11197);
or OR4 (N11621, N11613, N2082, N681, N3967);
nand NAND4 (N11622, N11605, N10448, N4611, N9458);
and AND3 (N11623, N11622, N3593, N8675);
or OR3 (N11624, N11621, N339, N11405);
and AND2 (N11625, N11617, N3552);
buf BUF1 (N11626, N11623);
nand NAND2 (N11627, N11609, N3017);
buf BUF1 (N11628, N11616);
nand NAND2 (N11629, N11614, N3614);
nor NOR3 (N11630, N11628, N4635, N1883);
buf BUF1 (N11631, N11610);
nand NAND3 (N11632, N11608, N4035, N636);
not NOT1 (N11633, N11626);
nor NOR2 (N11634, N11632, N4709);
buf BUF1 (N11635, N11631);
and AND2 (N11636, N11619, N1786);
buf BUF1 (N11637, N11636);
not NOT1 (N11638, N11624);
not NOT1 (N11639, N11620);
buf BUF1 (N11640, N11625);
buf BUF1 (N11641, N11638);
nor NOR2 (N11642, N11629, N11047);
nand NAND3 (N11643, N11639, N9935, N1428);
nor NOR3 (N11644, N11635, N7624, N5824);
nand NAND3 (N11645, N11643, N4134, N8416);
nor NOR3 (N11646, N11627, N6675, N9850);
or OR3 (N11647, N11634, N4816, N5689);
nand NAND3 (N11648, N11644, N319, N5949);
and AND3 (N11649, N11633, N7899, N4594);
nand NAND4 (N11650, N11646, N11347, N4875, N5222);
xor XOR2 (N11651, N11648, N9749);
nor NOR4 (N11652, N11640, N10199, N7933, N6319);
nand NAND2 (N11653, N11645, N1475);
nor NOR4 (N11654, N11630, N10196, N6512, N1991);
nor NOR4 (N11655, N11649, N2072, N2766, N8668);
nor NOR3 (N11656, N11655, N8575, N9662);
or OR4 (N11657, N11651, N659, N6079, N9275);
nand NAND2 (N11658, N11637, N7764);
buf BUF1 (N11659, N11641);
nand NAND3 (N11660, N11647, N7601, N9586);
or OR4 (N11661, N11653, N5964, N4598, N2788);
nor NOR3 (N11662, N11654, N10354, N10115);
nand NAND4 (N11663, N11642, N974, N5387, N7397);
nand NAND2 (N11664, N11660, N10859);
or OR2 (N11665, N11663, N9482);
not NOT1 (N11666, N11659);
and AND4 (N11667, N11662, N4509, N3323, N3767);
nor NOR4 (N11668, N11666, N10235, N3890, N7405);
buf BUF1 (N11669, N11650);
and AND3 (N11670, N11667, N5242, N5006);
and AND3 (N11671, N11670, N4745, N7690);
xor XOR2 (N11672, N11668, N7698);
nor NOR2 (N11673, N11652, N126);
not NOT1 (N11674, N11661);
nand NAND2 (N11675, N11658, N1089);
nor NOR2 (N11676, N11665, N10295);
not NOT1 (N11677, N11675);
and AND2 (N11678, N11674, N3895);
and AND3 (N11679, N11669, N4333, N4554);
buf BUF1 (N11680, N11678);
and AND3 (N11681, N11657, N9236, N2021);
xor XOR2 (N11682, N11676, N5430);
or OR3 (N11683, N11677, N301, N5510);
xor XOR2 (N11684, N11656, N8032);
nor NOR4 (N11685, N11664, N1784, N4184, N8493);
buf BUF1 (N11686, N11680);
xor XOR2 (N11687, N11673, N481);
not NOT1 (N11688, N11683);
xor XOR2 (N11689, N11684, N7539);
not NOT1 (N11690, N11681);
and AND3 (N11691, N11679, N8049, N6615);
not NOT1 (N11692, N11682);
not NOT1 (N11693, N11688);
and AND3 (N11694, N11692, N6068, N11279);
not NOT1 (N11695, N11690);
nand NAND2 (N11696, N11695, N7488);
and AND2 (N11697, N11685, N3485);
nor NOR4 (N11698, N11672, N10308, N1845, N8874);
and AND4 (N11699, N11686, N9664, N10527, N11333);
or OR2 (N11700, N11699, N6120);
xor XOR2 (N11701, N11700, N1119);
not NOT1 (N11702, N11698);
or OR2 (N11703, N11694, N8583);
nor NOR3 (N11704, N11701, N2786, N9365);
nand NAND3 (N11705, N11687, N4678, N2133);
or OR2 (N11706, N11693, N3384);
nand NAND2 (N11707, N11702, N5627);
nor NOR4 (N11708, N11703, N1994, N3211, N2698);
nor NOR2 (N11709, N11707, N1036);
not NOT1 (N11710, N11696);
not NOT1 (N11711, N11709);
nand NAND2 (N11712, N11708, N899);
or OR4 (N11713, N11711, N7191, N11452, N2367);
not NOT1 (N11714, N11712);
nand NAND4 (N11715, N11714, N8530, N6746, N3959);
not NOT1 (N11716, N11705);
not NOT1 (N11717, N11704);
not NOT1 (N11718, N11697);
nand NAND3 (N11719, N11715, N305, N10299);
buf BUF1 (N11720, N11671);
buf BUF1 (N11721, N11710);
or OR3 (N11722, N11691, N9828, N1498);
nor NOR4 (N11723, N11706, N8369, N10798, N7366);
nand NAND2 (N11724, N11716, N11716);
buf BUF1 (N11725, N11724);
xor XOR2 (N11726, N11718, N7272);
nand NAND2 (N11727, N11719, N11610);
or OR2 (N11728, N11723, N529);
xor XOR2 (N11729, N11689, N4551);
not NOT1 (N11730, N11722);
xor XOR2 (N11731, N11720, N5979);
nor NOR2 (N11732, N11728, N4172);
and AND3 (N11733, N11725, N8537, N6397);
buf BUF1 (N11734, N11733);
nand NAND2 (N11735, N11729, N7310);
and AND4 (N11736, N11717, N3289, N10759, N10522);
xor XOR2 (N11737, N11736, N7644);
nand NAND3 (N11738, N11735, N7774, N2446);
or OR4 (N11739, N11731, N10382, N1632, N3518);
not NOT1 (N11740, N11739);
and AND4 (N11741, N11737, N6279, N1593, N1477);
xor XOR2 (N11742, N11721, N6397);
xor XOR2 (N11743, N11742, N11636);
nand NAND3 (N11744, N11730, N4789, N4884);
nand NAND2 (N11745, N11740, N2634);
nor NOR2 (N11746, N11744, N2141);
or OR2 (N11747, N11726, N3413);
not NOT1 (N11748, N11727);
nor NOR3 (N11749, N11741, N10041, N9339);
not NOT1 (N11750, N11743);
nor NOR2 (N11751, N11745, N7554);
and AND4 (N11752, N11748, N8410, N5886, N4314);
and AND4 (N11753, N11713, N538, N6362, N4168);
xor XOR2 (N11754, N11749, N9550);
and AND4 (N11755, N11738, N7773, N3037, N8804);
nor NOR3 (N11756, N11750, N859, N10289);
or OR2 (N11757, N11755, N5466);
nor NOR4 (N11758, N11753, N6372, N10071, N1981);
nor NOR3 (N11759, N11757, N10389, N3985);
nor NOR3 (N11760, N11752, N6604, N3509);
not NOT1 (N11761, N11754);
xor XOR2 (N11762, N11746, N11735);
nand NAND2 (N11763, N11747, N3187);
xor XOR2 (N11764, N11756, N6935);
nor NOR2 (N11765, N11758, N7094);
xor XOR2 (N11766, N11764, N10861);
and AND3 (N11767, N11759, N875, N5438);
xor XOR2 (N11768, N11765, N6242);
xor XOR2 (N11769, N11762, N10359);
xor XOR2 (N11770, N11769, N8330);
buf BUF1 (N11771, N11760);
not NOT1 (N11772, N11770);
xor XOR2 (N11773, N11767, N2128);
not NOT1 (N11774, N11763);
or OR3 (N11775, N11761, N8252, N877);
not NOT1 (N11776, N11771);
nor NOR2 (N11777, N11776, N6295);
xor XOR2 (N11778, N11775, N11097);
and AND3 (N11779, N11777, N1159, N7827);
buf BUF1 (N11780, N11774);
buf BUF1 (N11781, N11780);
buf BUF1 (N11782, N11773);
nand NAND2 (N11783, N11751, N2681);
xor XOR2 (N11784, N11781, N3228);
not NOT1 (N11785, N11768);
nor NOR2 (N11786, N11785, N5065);
xor XOR2 (N11787, N11779, N1993);
not NOT1 (N11788, N11782);
nand NAND3 (N11789, N11783, N7242, N4421);
nand NAND3 (N11790, N11772, N5644, N9901);
nor NOR4 (N11791, N11789, N10953, N5756, N8459);
xor XOR2 (N11792, N11732, N5127);
nand NAND4 (N11793, N11766, N3484, N5418, N5909);
not NOT1 (N11794, N11788);
buf BUF1 (N11795, N11786);
not NOT1 (N11796, N11787);
not NOT1 (N11797, N11793);
or OR2 (N11798, N11734, N7687);
and AND2 (N11799, N11784, N4908);
xor XOR2 (N11800, N11790, N5565);
nand NAND2 (N11801, N11791, N3485);
and AND3 (N11802, N11796, N11027, N11387);
and AND4 (N11803, N11802, N3216, N2767, N11780);
nand NAND2 (N11804, N11778, N3683);
not NOT1 (N11805, N11800);
and AND4 (N11806, N11803, N7817, N4160, N10134);
nor NOR2 (N11807, N11797, N7562);
nand NAND2 (N11808, N11795, N8197);
nor NOR3 (N11809, N11807, N10820, N2415);
buf BUF1 (N11810, N11801);
buf BUF1 (N11811, N11808);
and AND2 (N11812, N11809, N10027);
nand NAND2 (N11813, N11799, N2450);
not NOT1 (N11814, N11810);
and AND2 (N11815, N11813, N10656);
and AND4 (N11816, N11798, N10648, N4654, N9776);
xor XOR2 (N11817, N11815, N8649);
nor NOR3 (N11818, N11794, N10262, N761);
buf BUF1 (N11819, N11814);
and AND3 (N11820, N11805, N9148, N8356);
nand NAND3 (N11821, N11811, N1433, N8640);
xor XOR2 (N11822, N11818, N2276);
xor XOR2 (N11823, N11806, N2981);
nor NOR2 (N11824, N11821, N4107);
nand NAND4 (N11825, N11817, N933, N1460, N872);
nor NOR4 (N11826, N11820, N11384, N6305, N3406);
nor NOR3 (N11827, N11819, N3525, N1369);
or OR3 (N11828, N11804, N11447, N10825);
and AND3 (N11829, N11816, N9813, N8188);
and AND3 (N11830, N11824, N11555, N4722);
and AND4 (N11831, N11830, N6298, N1323, N492);
and AND4 (N11832, N11828, N6028, N5026, N10477);
xor XOR2 (N11833, N11832, N9349);
buf BUF1 (N11834, N11822);
nor NOR3 (N11835, N11829, N2715, N4013);
or OR2 (N11836, N11834, N8645);
nand NAND3 (N11837, N11835, N3293, N5569);
nor NOR2 (N11838, N11826, N3408);
and AND4 (N11839, N11825, N1229, N9739, N6429);
nor NOR4 (N11840, N11838, N3491, N3385, N5044);
xor XOR2 (N11841, N11839, N8831);
buf BUF1 (N11842, N11841);
nor NOR2 (N11843, N11842, N221);
or OR3 (N11844, N11823, N8966, N4689);
xor XOR2 (N11845, N11827, N5299);
buf BUF1 (N11846, N11833);
nor NOR4 (N11847, N11844, N7938, N4083, N2623);
nand NAND3 (N11848, N11836, N5220, N4349);
nand NAND2 (N11849, N11847, N7864);
xor XOR2 (N11850, N11845, N923);
xor XOR2 (N11851, N11846, N5953);
or OR2 (N11852, N11843, N9342);
or OR3 (N11853, N11851, N5863, N8843);
buf BUF1 (N11854, N11853);
or OR4 (N11855, N11812, N3151, N3486, N3997);
xor XOR2 (N11856, N11792, N11093);
buf BUF1 (N11857, N11848);
xor XOR2 (N11858, N11837, N9949);
or OR3 (N11859, N11831, N5021, N7565);
or OR4 (N11860, N11857, N6098, N3008, N4800);
or OR3 (N11861, N11854, N7120, N6302);
buf BUF1 (N11862, N11849);
not NOT1 (N11863, N11840);
nand NAND3 (N11864, N11862, N1639, N7731);
buf BUF1 (N11865, N11850);
buf BUF1 (N11866, N11858);
xor XOR2 (N11867, N11866, N8369);
xor XOR2 (N11868, N11852, N2759);
buf BUF1 (N11869, N11856);
nor NOR4 (N11870, N11861, N6551, N4100, N8743);
and AND4 (N11871, N11869, N207, N6892, N10938);
not NOT1 (N11872, N11870);
and AND4 (N11873, N11871, N9142, N5501, N1011);
and AND3 (N11874, N11859, N6744, N5837);
and AND2 (N11875, N11855, N1840);
nand NAND2 (N11876, N11867, N487);
buf BUF1 (N11877, N11864);
xor XOR2 (N11878, N11865, N11374);
buf BUF1 (N11879, N11874);
nor NOR3 (N11880, N11879, N2561, N4204);
and AND4 (N11881, N11880, N8327, N7209, N1887);
or OR2 (N11882, N11878, N1197);
and AND2 (N11883, N11882, N5020);
not NOT1 (N11884, N11860);
nand NAND4 (N11885, N11868, N9991, N7044, N5132);
nor NOR4 (N11886, N11873, N6483, N11570, N11651);
and AND3 (N11887, N11886, N9724, N1296);
nand NAND4 (N11888, N11881, N4219, N7226, N10597);
nor NOR2 (N11889, N11883, N4482);
buf BUF1 (N11890, N11887);
and AND2 (N11891, N11875, N9522);
nand NAND3 (N11892, N11876, N7079, N10787);
not NOT1 (N11893, N11889);
not NOT1 (N11894, N11890);
not NOT1 (N11895, N11894);
nand NAND4 (N11896, N11877, N7188, N7122, N6706);
not NOT1 (N11897, N11892);
or OR3 (N11898, N11896, N4023, N3494);
nand NAND3 (N11899, N11893, N11265, N11625);
not NOT1 (N11900, N11863);
nor NOR2 (N11901, N11897, N6129);
nand NAND4 (N11902, N11885, N3370, N3332, N2963);
or OR4 (N11903, N11902, N5575, N623, N6148);
nand NAND2 (N11904, N11901, N2540);
and AND2 (N11905, N11884, N11381);
xor XOR2 (N11906, N11898, N2416);
nor NOR2 (N11907, N11895, N7182);
buf BUF1 (N11908, N11903);
and AND4 (N11909, N11891, N1073, N6513, N1097);
buf BUF1 (N11910, N11904);
nand NAND4 (N11911, N11888, N7946, N7846, N8991);
xor XOR2 (N11912, N11907, N2449);
not NOT1 (N11913, N11910);
xor XOR2 (N11914, N11872, N1657);
nor NOR3 (N11915, N11914, N11689, N1312);
or OR2 (N11916, N11906, N9344);
not NOT1 (N11917, N11899);
or OR4 (N11918, N11912, N9330, N2958, N7600);
nand NAND4 (N11919, N11909, N9855, N6377, N6766);
buf BUF1 (N11920, N11911);
and AND4 (N11921, N11913, N6625, N1115, N5575);
buf BUF1 (N11922, N11900);
or OR2 (N11923, N11918, N3714);
not NOT1 (N11924, N11923);
buf BUF1 (N11925, N11924);
not NOT1 (N11926, N11908);
not NOT1 (N11927, N11917);
nor NOR2 (N11928, N11927, N931);
buf BUF1 (N11929, N11915);
and AND3 (N11930, N11929, N9096, N2253);
nor NOR2 (N11931, N11922, N7746);
not NOT1 (N11932, N11905);
xor XOR2 (N11933, N11931, N10050);
xor XOR2 (N11934, N11926, N10550);
or OR2 (N11935, N11928, N5366);
and AND3 (N11936, N11921, N7657, N8000);
nand NAND3 (N11937, N11933, N9838, N5074);
not NOT1 (N11938, N11925);
nor NOR2 (N11939, N11932, N11238);
xor XOR2 (N11940, N11938, N8200);
not NOT1 (N11941, N11920);
or OR3 (N11942, N11916, N4996, N7620);
xor XOR2 (N11943, N11919, N8660);
buf BUF1 (N11944, N11941);
and AND3 (N11945, N11937, N3811, N1294);
and AND3 (N11946, N11942, N1955, N2669);
nor NOR2 (N11947, N11936, N6300);
and AND4 (N11948, N11943, N10678, N1158, N7872);
nand NAND4 (N11949, N11935, N11830, N8153, N2538);
nor NOR2 (N11950, N11939, N4335);
nand NAND3 (N11951, N11946, N3702, N10913);
not NOT1 (N11952, N11944);
not NOT1 (N11953, N11930);
nor NOR4 (N11954, N11948, N5799, N10572, N1863);
buf BUF1 (N11955, N11953);
nand NAND4 (N11956, N11950, N6046, N7803, N10976);
or OR3 (N11957, N11951, N1512, N11861);
not NOT1 (N11958, N11945);
or OR2 (N11959, N11949, N9123);
xor XOR2 (N11960, N11955, N8843);
nand NAND2 (N11961, N11954, N8488);
not NOT1 (N11962, N11959);
or OR3 (N11963, N11934, N10893, N6448);
not NOT1 (N11964, N11947);
nand NAND3 (N11965, N11952, N11483, N4841);
xor XOR2 (N11966, N11960, N4146);
nor NOR4 (N11967, N11958, N753, N818, N11033);
nor NOR3 (N11968, N11940, N2197, N9891);
not NOT1 (N11969, N11963);
xor XOR2 (N11970, N11965, N7373);
not NOT1 (N11971, N11968);
or OR4 (N11972, N11964, N11747, N1206, N4669);
nor NOR4 (N11973, N11966, N621, N11682, N9758);
not NOT1 (N11974, N11967);
buf BUF1 (N11975, N11957);
xor XOR2 (N11976, N11973, N4606);
not NOT1 (N11977, N11974);
nor NOR3 (N11978, N11961, N10247, N7617);
nor NOR2 (N11979, N11956, N3470);
and AND2 (N11980, N11969, N6971);
and AND4 (N11981, N11979, N4962, N10675, N577);
not NOT1 (N11982, N11971);
buf BUF1 (N11983, N11976);
buf BUF1 (N11984, N11977);
nand NAND2 (N11985, N11983, N497);
and AND3 (N11986, N11972, N4117, N1099);
xor XOR2 (N11987, N11962, N128);
not NOT1 (N11988, N11985);
buf BUF1 (N11989, N11980);
nand NAND4 (N11990, N11984, N854, N5244, N8786);
nand NAND4 (N11991, N11986, N2155, N2966, N10072);
or OR3 (N11992, N11975, N8591, N47);
not NOT1 (N11993, N11991);
or OR2 (N11994, N11981, N5483);
nor NOR2 (N11995, N11970, N9792);
nand NAND3 (N11996, N11988, N1190, N10062);
xor XOR2 (N11997, N11996, N297);
xor XOR2 (N11998, N11993, N3089);
or OR4 (N11999, N11987, N72, N8544, N342);
and AND3 (N12000, N11998, N2115, N4495);
buf BUF1 (N12001, N11992);
not NOT1 (N12002, N11997);
not NOT1 (N12003, N11978);
buf BUF1 (N12004, N11990);
and AND2 (N12005, N11982, N11109);
xor XOR2 (N12006, N12000, N7290);
nand NAND3 (N12007, N11995, N7690, N11857);
not NOT1 (N12008, N12006);
buf BUF1 (N12009, N12003);
xor XOR2 (N12010, N11989, N9731);
and AND3 (N12011, N12009, N4542, N6312);
xor XOR2 (N12012, N12011, N7866);
and AND4 (N12013, N12012, N7707, N9090, N3977);
not NOT1 (N12014, N12004);
not NOT1 (N12015, N12001);
buf BUF1 (N12016, N12015);
or OR3 (N12017, N12013, N8682, N5768);
nor NOR2 (N12018, N12010, N8634);
not NOT1 (N12019, N12005);
xor XOR2 (N12020, N11999, N5267);
nor NOR3 (N12021, N12007, N11769, N10617);
nand NAND2 (N12022, N12016, N1346);
xor XOR2 (N12023, N12014, N5880);
buf BUF1 (N12024, N12022);
xor XOR2 (N12025, N11994, N10671);
buf BUF1 (N12026, N12021);
buf BUF1 (N12027, N12008);
or OR3 (N12028, N12025, N9928, N5881);
nand NAND3 (N12029, N12023, N10597, N8709);
nand NAND3 (N12030, N12018, N1882, N10110);
xor XOR2 (N12031, N12002, N4075);
nor NOR4 (N12032, N12028, N11936, N4524, N10324);
xor XOR2 (N12033, N12020, N7096);
nor NOR3 (N12034, N12031, N4992, N10983);
buf BUF1 (N12035, N12027);
not NOT1 (N12036, N12024);
nand NAND2 (N12037, N12033, N9316);
nand NAND2 (N12038, N12034, N8502);
xor XOR2 (N12039, N12019, N181);
and AND3 (N12040, N12017, N7501, N877);
buf BUF1 (N12041, N12037);
and AND3 (N12042, N12038, N1237, N5878);
and AND3 (N12043, N12036, N10867, N7257);
xor XOR2 (N12044, N12041, N11786);
or OR2 (N12045, N12040, N2948);
buf BUF1 (N12046, N12039);
nand NAND2 (N12047, N12035, N4518);
not NOT1 (N12048, N12026);
nand NAND2 (N12049, N12043, N469);
and AND4 (N12050, N12049, N12038, N10027, N10388);
xor XOR2 (N12051, N12042, N9244);
or OR2 (N12052, N12046, N2125);
and AND4 (N12053, N12045, N392, N6131, N3197);
buf BUF1 (N12054, N12047);
not NOT1 (N12055, N12052);
xor XOR2 (N12056, N12051, N2992);
nor NOR4 (N12057, N12055, N5079, N7103, N2212);
or OR4 (N12058, N12044, N8885, N3336, N6001);
nor NOR4 (N12059, N12029, N2036, N10564, N10682);
buf BUF1 (N12060, N12059);
not NOT1 (N12061, N12060);
nor NOR4 (N12062, N12048, N6274, N3154, N3973);
or OR4 (N12063, N12057, N5187, N2464, N4772);
or OR3 (N12064, N12062, N1398, N2924);
not NOT1 (N12065, N12064);
xor XOR2 (N12066, N12061, N57);
nand NAND2 (N12067, N12066, N10931);
xor XOR2 (N12068, N12050, N8562);
or OR2 (N12069, N12058, N3834);
or OR4 (N12070, N12063, N262, N3904, N6582);
or OR2 (N12071, N12067, N7035);
buf BUF1 (N12072, N12054);
not NOT1 (N12073, N12053);
or OR2 (N12074, N12073, N5593);
nor NOR3 (N12075, N12070, N11959, N933);
and AND4 (N12076, N12056, N9879, N10973, N6928);
or OR3 (N12077, N12072, N785, N1705);
or OR3 (N12078, N12032, N11418, N2197);
buf BUF1 (N12079, N12071);
nand NAND4 (N12080, N12075, N10076, N5175, N5382);
nor NOR3 (N12081, N12030, N5950, N3952);
nor NOR4 (N12082, N12074, N1008, N6164, N5999);
xor XOR2 (N12083, N12077, N9981);
and AND2 (N12084, N12078, N9212);
or OR4 (N12085, N12083, N9237, N2855, N528);
nor NOR4 (N12086, N12081, N3145, N9489, N7625);
and AND2 (N12087, N12069, N11862);
not NOT1 (N12088, N12084);
and AND3 (N12089, N12087, N3250, N7631);
buf BUF1 (N12090, N12065);
xor XOR2 (N12091, N12079, N5655);
nand NAND3 (N12092, N12076, N7685, N1017);
buf BUF1 (N12093, N12086);
nor NOR2 (N12094, N12085, N3008);
and AND3 (N12095, N12091, N390, N7949);
not NOT1 (N12096, N12093);
and AND3 (N12097, N12094, N10628, N10915);
and AND4 (N12098, N12080, N1926, N9257, N10220);
buf BUF1 (N12099, N12082);
nor NOR2 (N12100, N12088, N6952);
nor NOR3 (N12101, N12100, N2048, N5313);
buf BUF1 (N12102, N12099);
nand NAND2 (N12103, N12101, N9407);
or OR3 (N12104, N12097, N7973, N2301);
nand NAND2 (N12105, N12092, N8194);
nor NOR2 (N12106, N12068, N260);
and AND4 (N12107, N12095, N3566, N11794, N2069);
xor XOR2 (N12108, N12096, N9439);
xor XOR2 (N12109, N12104, N5393);
buf BUF1 (N12110, N12098);
nand NAND2 (N12111, N12110, N11227);
xor XOR2 (N12112, N12109, N6664);
or OR4 (N12113, N12105, N10188, N3915, N2407);
or OR3 (N12114, N12089, N2170, N2833);
or OR4 (N12115, N12102, N7623, N2409, N11426);
or OR4 (N12116, N12113, N11156, N6037, N1683);
not NOT1 (N12117, N12114);
not NOT1 (N12118, N12103);
or OR4 (N12119, N12106, N8438, N2674, N8013);
not NOT1 (N12120, N12112);
or OR4 (N12121, N12120, N8108, N1291, N1248);
nand NAND2 (N12122, N12115, N1026);
nor NOR3 (N12123, N12121, N10244, N636);
or OR2 (N12124, N12118, N2413);
nor NOR3 (N12125, N12123, N6138, N11884);
buf BUF1 (N12126, N12125);
and AND4 (N12127, N12126, N4968, N884, N2865);
or OR3 (N12128, N12127, N5858, N1416);
not NOT1 (N12129, N12119);
nor NOR4 (N12130, N12107, N6141, N5882, N7520);
nor NOR2 (N12131, N12117, N2624);
buf BUF1 (N12132, N12108);
nor NOR3 (N12133, N12130, N4564, N4707);
or OR2 (N12134, N12128, N8039);
xor XOR2 (N12135, N12132, N5840);
not NOT1 (N12136, N12116);
xor XOR2 (N12137, N12136, N3793);
nor NOR2 (N12138, N12124, N1130);
not NOT1 (N12139, N12134);
xor XOR2 (N12140, N12139, N10604);
xor XOR2 (N12141, N12129, N7498);
xor XOR2 (N12142, N12140, N10522);
buf BUF1 (N12143, N12142);
or OR3 (N12144, N12122, N345, N10030);
nand NAND4 (N12145, N12137, N1381, N7115, N1098);
not NOT1 (N12146, N12133);
and AND3 (N12147, N12143, N6504, N1335);
and AND4 (N12148, N12146, N5163, N8988, N5422);
or OR2 (N12149, N12138, N1053);
nor NOR3 (N12150, N12149, N450, N9307);
not NOT1 (N12151, N12090);
buf BUF1 (N12152, N12145);
nor NOR3 (N12153, N12152, N5482, N270);
nor NOR4 (N12154, N12141, N3645, N571, N9604);
buf BUF1 (N12155, N12151);
buf BUF1 (N12156, N12111);
and AND2 (N12157, N12155, N4511);
or OR2 (N12158, N12144, N4505);
nand NAND4 (N12159, N12153, N1642, N11579, N632);
not NOT1 (N12160, N12147);
and AND4 (N12161, N12148, N668, N1658, N4003);
not NOT1 (N12162, N12157);
xor XOR2 (N12163, N12150, N2074);
xor XOR2 (N12164, N12158, N1189);
and AND4 (N12165, N12156, N6172, N11355, N4753);
xor XOR2 (N12166, N12163, N5083);
and AND2 (N12167, N12135, N6590);
xor XOR2 (N12168, N12167, N8463);
buf BUF1 (N12169, N12165);
nand NAND4 (N12170, N12131, N2814, N11690, N10289);
xor XOR2 (N12171, N12168, N1690);
and AND2 (N12172, N12171, N8782);
or OR3 (N12173, N12164, N953, N10797);
or OR4 (N12174, N12160, N5278, N1441, N3802);
nand NAND3 (N12175, N12174, N7882, N2328);
xor XOR2 (N12176, N12169, N9778);
nor NOR2 (N12177, N12173, N3221);
nand NAND2 (N12178, N12166, N9350);
buf BUF1 (N12179, N12177);
and AND4 (N12180, N12170, N4645, N2475, N3166);
and AND3 (N12181, N12176, N5541, N7124);
and AND3 (N12182, N12178, N401, N11730);
or OR2 (N12183, N12182, N5936);
nor NOR4 (N12184, N12175, N8605, N6604, N7723);
and AND3 (N12185, N12183, N453, N10738);
xor XOR2 (N12186, N12184, N4187);
xor XOR2 (N12187, N12185, N9221);
and AND3 (N12188, N12162, N947, N5385);
and AND2 (N12189, N12161, N1234);
or OR4 (N12190, N12181, N11656, N11299, N86);
or OR4 (N12191, N12154, N757, N1981, N6486);
nor NOR4 (N12192, N12188, N7402, N583, N5385);
buf BUF1 (N12193, N12191);
or OR3 (N12194, N12190, N5982, N11423);
or OR2 (N12195, N12193, N10631);
xor XOR2 (N12196, N12194, N5190);
nand NAND3 (N12197, N12172, N5246, N7725);
not NOT1 (N12198, N12189);
buf BUF1 (N12199, N12196);
buf BUF1 (N12200, N12186);
buf BUF1 (N12201, N12200);
xor XOR2 (N12202, N12199, N435);
and AND3 (N12203, N12192, N921, N8544);
buf BUF1 (N12204, N12187);
buf BUF1 (N12205, N12202);
nand NAND4 (N12206, N12159, N183, N2712, N1684);
nor NOR4 (N12207, N12204, N2160, N1794, N9066);
not NOT1 (N12208, N12201);
not NOT1 (N12209, N12203);
and AND3 (N12210, N12195, N1091, N6549);
or OR4 (N12211, N12208, N10994, N5465, N7521);
not NOT1 (N12212, N12198);
nand NAND2 (N12213, N12209, N4965);
buf BUF1 (N12214, N12213);
or OR3 (N12215, N12205, N9253, N2402);
and AND3 (N12216, N12215, N7720, N10641);
buf BUF1 (N12217, N12206);
nor NOR3 (N12218, N12211, N4674, N9980);
buf BUF1 (N12219, N12180);
or OR2 (N12220, N12210, N76);
nand NAND2 (N12221, N12212, N1679);
or OR2 (N12222, N12221, N10341);
and AND4 (N12223, N12216, N7913, N3679, N1795);
or OR2 (N12224, N12207, N1612);
buf BUF1 (N12225, N12217);
and AND2 (N12226, N12224, N5610);
nor NOR2 (N12227, N12219, N3098);
nor NOR3 (N12228, N12197, N8157, N6270);
nor NOR2 (N12229, N12218, N3992);
nor NOR3 (N12230, N12228, N12025, N10272);
buf BUF1 (N12231, N12222);
xor XOR2 (N12232, N12231, N2623);
and AND2 (N12233, N12230, N2947);
and AND4 (N12234, N12214, N10339, N6126, N1010);
or OR2 (N12235, N12232, N3778);
or OR3 (N12236, N12233, N5317, N11415);
not NOT1 (N12237, N12223);
and AND2 (N12238, N12229, N3842);
buf BUF1 (N12239, N12225);
and AND4 (N12240, N12179, N12201, N7193, N6914);
xor XOR2 (N12241, N12220, N11123);
and AND2 (N12242, N12237, N11300);
not NOT1 (N12243, N12234);
or OR2 (N12244, N12242, N6686);
not NOT1 (N12245, N12227);
xor XOR2 (N12246, N12226, N1858);
or OR3 (N12247, N12235, N5196, N9114);
xor XOR2 (N12248, N12241, N7139);
nand NAND2 (N12249, N12244, N11877);
xor XOR2 (N12250, N12236, N1091);
not NOT1 (N12251, N12238);
xor XOR2 (N12252, N12245, N2627);
and AND2 (N12253, N12252, N6836);
or OR4 (N12254, N12251, N2499, N7536, N8133);
xor XOR2 (N12255, N12247, N12206);
or OR4 (N12256, N12240, N9765, N1655, N4464);
and AND2 (N12257, N12239, N3093);
nor NOR2 (N12258, N12250, N5960);
xor XOR2 (N12259, N12243, N6682);
not NOT1 (N12260, N12258);
not NOT1 (N12261, N12254);
and AND2 (N12262, N12246, N7515);
buf BUF1 (N12263, N12260);
not NOT1 (N12264, N12255);
buf BUF1 (N12265, N12249);
and AND4 (N12266, N12256, N9665, N10337, N6474);
nand NAND3 (N12267, N12253, N2751, N10705);
nand NAND3 (N12268, N12257, N8113, N7847);
xor XOR2 (N12269, N12262, N10643);
not NOT1 (N12270, N12268);
or OR2 (N12271, N12269, N5509);
buf BUF1 (N12272, N12265);
and AND3 (N12273, N12270, N7404, N9640);
xor XOR2 (N12274, N12261, N2790);
xor XOR2 (N12275, N12272, N8605);
xor XOR2 (N12276, N12273, N10431);
and AND3 (N12277, N12259, N520, N4955);
and AND2 (N12278, N12274, N11544);
nand NAND3 (N12279, N12248, N9986, N9924);
not NOT1 (N12280, N12279);
nor NOR4 (N12281, N12280, N3976, N11663, N2598);
nor NOR3 (N12282, N12266, N3694, N8674);
buf BUF1 (N12283, N12271);
buf BUF1 (N12284, N12267);
nand NAND3 (N12285, N12284, N2792, N268);
buf BUF1 (N12286, N12285);
nand NAND3 (N12287, N12281, N654, N8084);
or OR3 (N12288, N12275, N1939, N6636);
not NOT1 (N12289, N12287);
not NOT1 (N12290, N12278);
buf BUF1 (N12291, N12276);
nand NAND2 (N12292, N12264, N3656);
buf BUF1 (N12293, N12290);
not NOT1 (N12294, N12289);
and AND2 (N12295, N12292, N11441);
buf BUF1 (N12296, N12263);
or OR3 (N12297, N12286, N4665, N1150);
not NOT1 (N12298, N12283);
xor XOR2 (N12299, N12277, N9162);
xor XOR2 (N12300, N12298, N6523);
nor NOR4 (N12301, N12300, N8801, N1109, N6533);
xor XOR2 (N12302, N12297, N7211);
not NOT1 (N12303, N12288);
xor XOR2 (N12304, N12291, N812);
nand NAND2 (N12305, N12294, N10316);
nand NAND4 (N12306, N12299, N2355, N4540, N1187);
nor NOR4 (N12307, N12295, N8118, N7499, N11497);
and AND4 (N12308, N12303, N11508, N125, N7287);
nor NOR4 (N12309, N12296, N8645, N6194, N6658);
nand NAND2 (N12310, N12309, N2529);
xor XOR2 (N12311, N12305, N1187);
buf BUF1 (N12312, N12282);
xor XOR2 (N12313, N12293, N8961);
or OR4 (N12314, N12310, N10907, N8535, N11731);
xor XOR2 (N12315, N12302, N907);
nor NOR3 (N12316, N12313, N10021, N5741);
buf BUF1 (N12317, N12304);
not NOT1 (N12318, N12312);
nand NAND3 (N12319, N12308, N3972, N5656);
xor XOR2 (N12320, N12319, N1065);
nand NAND3 (N12321, N12318, N7690, N8995);
or OR2 (N12322, N12301, N6342);
and AND2 (N12323, N12315, N9676);
and AND2 (N12324, N12322, N6677);
nand NAND4 (N12325, N12307, N7076, N9094, N10031);
nand NAND3 (N12326, N12317, N9193, N974);
nor NOR4 (N12327, N12326, N6955, N9955, N100);
buf BUF1 (N12328, N12321);
not NOT1 (N12329, N12325);
nor NOR4 (N12330, N12329, N569, N8263, N11839);
nand NAND4 (N12331, N12328, N12212, N1787, N2048);
not NOT1 (N12332, N12306);
nand NAND3 (N12333, N12332, N7987, N5112);
nor NOR4 (N12334, N12324, N3665, N1252, N11857);
nor NOR4 (N12335, N12331, N5331, N8472, N2168);
nor NOR3 (N12336, N12311, N5406, N9738);
or OR4 (N12337, N12333, N5014, N6535, N4046);
not NOT1 (N12338, N12336);
nor NOR3 (N12339, N12323, N12232, N3531);
or OR3 (N12340, N12334, N3897, N1245);
not NOT1 (N12341, N12316);
nor NOR4 (N12342, N12330, N2332, N10906, N3175);
nor NOR4 (N12343, N12340, N304, N7320, N7590);
not NOT1 (N12344, N12314);
buf BUF1 (N12345, N12320);
or OR3 (N12346, N12342, N3834, N1120);
buf BUF1 (N12347, N12337);
nor NOR4 (N12348, N12346, N11991, N8896, N3604);
and AND2 (N12349, N12345, N12146);
and AND2 (N12350, N12339, N11616);
nand NAND2 (N12351, N12341, N8555);
xor XOR2 (N12352, N12327, N579);
nand NAND3 (N12353, N12351, N1400, N11145);
xor XOR2 (N12354, N12344, N1047);
nand NAND3 (N12355, N12335, N10145, N996);
buf BUF1 (N12356, N12347);
or OR3 (N12357, N12355, N6447, N11003);
or OR2 (N12358, N12353, N7575);
nand NAND2 (N12359, N12352, N11342);
nor NOR3 (N12360, N12357, N5831, N5676);
not NOT1 (N12361, N12360);
xor XOR2 (N12362, N12356, N4484);
buf BUF1 (N12363, N12338);
buf BUF1 (N12364, N12349);
nand NAND2 (N12365, N12361, N8212);
xor XOR2 (N12366, N12348, N3760);
nand NAND2 (N12367, N12343, N12293);
and AND4 (N12368, N12362, N3465, N9445, N5308);
xor XOR2 (N12369, N12365, N8336);
nand NAND2 (N12370, N12366, N10304);
and AND4 (N12371, N12368, N10218, N4591, N9214);
not NOT1 (N12372, N12363);
nand NAND2 (N12373, N12350, N11202);
or OR2 (N12374, N12367, N4505);
not NOT1 (N12375, N12372);
and AND4 (N12376, N12369, N9587, N10284, N11587);
xor XOR2 (N12377, N12354, N11043);
buf BUF1 (N12378, N12371);
and AND4 (N12379, N12358, N377, N8085, N250);
or OR2 (N12380, N12364, N1429);
xor XOR2 (N12381, N12370, N12216);
and AND4 (N12382, N12373, N9248, N4837, N10905);
nand NAND4 (N12383, N12374, N5989, N5105, N1365);
nor NOR4 (N12384, N12377, N487, N9068, N6314);
or OR2 (N12385, N12382, N9452);
buf BUF1 (N12386, N12380);
or OR3 (N12387, N12385, N1101, N5043);
xor XOR2 (N12388, N12386, N8502);
xor XOR2 (N12389, N12359, N8408);
and AND4 (N12390, N12375, N1064, N11990, N11747);
nor NOR3 (N12391, N12376, N10424, N11056);
xor XOR2 (N12392, N12379, N6713);
buf BUF1 (N12393, N12387);
buf BUF1 (N12394, N12391);
nor NOR4 (N12395, N12383, N2861, N1360, N12116);
buf BUF1 (N12396, N12390);
buf BUF1 (N12397, N12381);
buf BUF1 (N12398, N12388);
nand NAND4 (N12399, N12378, N5468, N6063, N11028);
nor NOR4 (N12400, N12398, N5221, N2064, N3093);
nand NAND2 (N12401, N12394, N4412);
not NOT1 (N12402, N12392);
not NOT1 (N12403, N12402);
nor NOR3 (N12404, N12384, N359, N11055);
buf BUF1 (N12405, N12389);
not NOT1 (N12406, N12401);
not NOT1 (N12407, N12396);
or OR3 (N12408, N12393, N2482, N12009);
or OR3 (N12409, N12404, N8934, N2415);
xor XOR2 (N12410, N12406, N11530);
xor XOR2 (N12411, N12395, N8741);
or OR3 (N12412, N12409, N10896, N11380);
xor XOR2 (N12413, N12408, N1452);
or OR4 (N12414, N12413, N8647, N2230, N1055);
nand NAND4 (N12415, N12399, N11031, N4065, N5429);
not NOT1 (N12416, N12410);
nand NAND3 (N12417, N12405, N7872, N3387);
or OR2 (N12418, N12411, N6781);
nor NOR3 (N12419, N12412, N4465, N10046);
nand NAND3 (N12420, N12419, N12290, N10468);
nor NOR3 (N12421, N12420, N8932, N7523);
not NOT1 (N12422, N12418);
buf BUF1 (N12423, N12397);
or OR2 (N12424, N12400, N3174);
buf BUF1 (N12425, N12416);
and AND3 (N12426, N12422, N6704, N10490);
and AND2 (N12427, N12417, N2877);
buf BUF1 (N12428, N12423);
xor XOR2 (N12429, N12426, N9269);
buf BUF1 (N12430, N12414);
nor NOR3 (N12431, N12425, N4051, N6470);
and AND2 (N12432, N12421, N3805);
or OR2 (N12433, N12415, N6613);
nand NAND2 (N12434, N12427, N4284);
nor NOR2 (N12435, N12432, N1095);
not NOT1 (N12436, N12403);
and AND3 (N12437, N12435, N2539, N6833);
buf BUF1 (N12438, N12433);
and AND2 (N12439, N12434, N6047);
buf BUF1 (N12440, N12438);
xor XOR2 (N12441, N12430, N932);
buf BUF1 (N12442, N12431);
and AND2 (N12443, N12442, N5049);
nand NAND2 (N12444, N12441, N8515);
xor XOR2 (N12445, N12443, N176);
nor NOR3 (N12446, N12429, N919, N5200);
nand NAND2 (N12447, N12445, N9411);
xor XOR2 (N12448, N12436, N7341);
nand NAND4 (N12449, N12446, N513, N5614, N2730);
not NOT1 (N12450, N12440);
or OR2 (N12451, N12444, N9048);
and AND4 (N12452, N12450, N211, N3309, N927);
buf BUF1 (N12453, N12437);
nor NOR4 (N12454, N12428, N6001, N8160, N8151);
xor XOR2 (N12455, N12449, N2687);
nor NOR2 (N12456, N12407, N8208);
and AND4 (N12457, N12448, N11715, N12322, N3382);
nand NAND2 (N12458, N12424, N11755);
nor NOR3 (N12459, N12452, N12199, N2974);
nand NAND3 (N12460, N12453, N7113, N10970);
xor XOR2 (N12461, N12458, N5193);
xor XOR2 (N12462, N12439, N11212);
not NOT1 (N12463, N12462);
buf BUF1 (N12464, N12456);
xor XOR2 (N12465, N12455, N4816);
nor NOR3 (N12466, N12447, N1498, N952);
and AND3 (N12467, N12457, N7017, N3604);
nand NAND3 (N12468, N12467, N7130, N3342);
not NOT1 (N12469, N12465);
and AND3 (N12470, N12451, N6143, N3473);
not NOT1 (N12471, N12468);
buf BUF1 (N12472, N12454);
or OR3 (N12473, N12470, N3905, N4463);
buf BUF1 (N12474, N12459);
xor XOR2 (N12475, N12474, N6329);
nor NOR2 (N12476, N12472, N7811);
and AND4 (N12477, N12473, N962, N2585, N12214);
nor NOR2 (N12478, N12471, N9500);
nand NAND3 (N12479, N12478, N11356, N11870);
or OR2 (N12480, N12464, N5985);
nor NOR4 (N12481, N12475, N3211, N6722, N7978);
and AND2 (N12482, N12463, N6548);
nand NAND2 (N12483, N12481, N1384);
nor NOR3 (N12484, N12479, N4829, N4560);
xor XOR2 (N12485, N12483, N4184);
xor XOR2 (N12486, N12469, N2412);
not NOT1 (N12487, N12486);
not NOT1 (N12488, N12480);
and AND4 (N12489, N12485, N8336, N6885, N2975);
or OR4 (N12490, N12482, N8733, N11833, N2247);
nor NOR3 (N12491, N12466, N2441, N6251);
and AND4 (N12492, N12489, N6921, N10339, N10562);
nand NAND4 (N12493, N12488, N169, N12451, N2099);
nor NOR4 (N12494, N12490, N5422, N1355, N12040);
and AND2 (N12495, N12461, N10571);
not NOT1 (N12496, N12494);
nand NAND2 (N12497, N12487, N9754);
not NOT1 (N12498, N12497);
nor NOR4 (N12499, N12484, N6547, N6668, N9893);
xor XOR2 (N12500, N12492, N58);
buf BUF1 (N12501, N12500);
xor XOR2 (N12502, N12476, N12019);
and AND3 (N12503, N12501, N5150, N7321);
or OR2 (N12504, N12498, N8487);
xor XOR2 (N12505, N12499, N11625);
not NOT1 (N12506, N12503);
nor NOR2 (N12507, N12506, N1611);
nor NOR4 (N12508, N12496, N12440, N11595, N6142);
nand NAND3 (N12509, N12505, N3609, N996);
or OR3 (N12510, N12477, N11157, N318);
xor XOR2 (N12511, N12502, N3765);
xor XOR2 (N12512, N12495, N4797);
xor XOR2 (N12513, N12504, N36);
xor XOR2 (N12514, N12508, N12510);
buf BUF1 (N12515, N10186);
nor NOR3 (N12516, N12515, N1511, N7361);
nor NOR2 (N12517, N12460, N2112);
not NOT1 (N12518, N12507);
xor XOR2 (N12519, N12518, N8148);
xor XOR2 (N12520, N12493, N11856);
not NOT1 (N12521, N12491);
not NOT1 (N12522, N12514);
xor XOR2 (N12523, N12520, N7135);
nand NAND4 (N12524, N12521, N6083, N9041, N11218);
xor XOR2 (N12525, N12512, N7930);
or OR3 (N12526, N12519, N9458, N6667);
xor XOR2 (N12527, N12513, N9172);
buf BUF1 (N12528, N12527);
or OR3 (N12529, N12509, N9187, N8011);
buf BUF1 (N12530, N12523);
xor XOR2 (N12531, N12526, N9122);
or OR4 (N12532, N12517, N11762, N3777, N3971);
nor NOR3 (N12533, N12511, N8162, N4129);
nand NAND4 (N12534, N12530, N12290, N8835, N5462);
not NOT1 (N12535, N12525);
xor XOR2 (N12536, N12524, N297);
buf BUF1 (N12537, N12534);
nor NOR4 (N12538, N12537, N795, N9997, N3139);
nand NAND4 (N12539, N12522, N1348, N11558, N2361);
nand NAND3 (N12540, N12539, N11586, N3191);
nor NOR2 (N12541, N12531, N4652);
or OR4 (N12542, N12533, N2114, N10604, N644);
or OR4 (N12543, N12541, N10444, N1511, N6979);
or OR4 (N12544, N12532, N5151, N11763, N7516);
buf BUF1 (N12545, N12540);
buf BUF1 (N12546, N12538);
or OR3 (N12547, N12529, N10095, N392);
buf BUF1 (N12548, N12543);
or OR2 (N12549, N12548, N6211);
and AND2 (N12550, N12549, N8556);
or OR2 (N12551, N12536, N11087);
xor XOR2 (N12552, N12535, N773);
nor NOR2 (N12553, N12542, N3635);
nand NAND4 (N12554, N12547, N7592, N693, N4410);
nand NAND4 (N12555, N12554, N7256, N3139, N1001);
buf BUF1 (N12556, N12553);
buf BUF1 (N12557, N12550);
not NOT1 (N12558, N12544);
not NOT1 (N12559, N12555);
or OR2 (N12560, N12552, N7920);
nand NAND3 (N12561, N12556, N803, N11036);
xor XOR2 (N12562, N12557, N4704);
nand NAND3 (N12563, N12559, N6366, N10639);
xor XOR2 (N12564, N12528, N8158);
not NOT1 (N12565, N12563);
buf BUF1 (N12566, N12551);
or OR3 (N12567, N12566, N10297, N6852);
or OR2 (N12568, N12558, N6026);
or OR2 (N12569, N12545, N10058);
nor NOR4 (N12570, N12564, N5246, N1005, N8032);
nor NOR2 (N12571, N12565, N10264);
not NOT1 (N12572, N12516);
and AND3 (N12573, N12567, N4219, N8128);
and AND2 (N12574, N12562, N4209);
buf BUF1 (N12575, N12560);
nor NOR3 (N12576, N12570, N4277, N3758);
buf BUF1 (N12577, N12573);
nand NAND2 (N12578, N12572, N8406);
not NOT1 (N12579, N12546);
nand NAND4 (N12580, N12569, N4880, N281, N8601);
xor XOR2 (N12581, N12577, N7098);
and AND2 (N12582, N12571, N5866);
xor XOR2 (N12583, N12578, N8107);
not NOT1 (N12584, N12568);
and AND4 (N12585, N12574, N7123, N8728, N11022);
and AND3 (N12586, N12581, N7969, N1317);
buf BUF1 (N12587, N12580);
and AND3 (N12588, N12561, N9726, N6646);
and AND2 (N12589, N12575, N10750);
nand NAND3 (N12590, N12579, N9405, N10404);
nand NAND2 (N12591, N12586, N11989);
xor XOR2 (N12592, N12589, N3295);
and AND2 (N12593, N12583, N5564);
nor NOR3 (N12594, N12588, N4001, N12473);
nor NOR2 (N12595, N12584, N2320);
nand NAND3 (N12596, N12585, N7036, N5284);
not NOT1 (N12597, N12592);
nand NAND2 (N12598, N12591, N4470);
buf BUF1 (N12599, N12593);
not NOT1 (N12600, N12599);
not NOT1 (N12601, N12576);
and AND3 (N12602, N12582, N711, N1229);
and AND4 (N12603, N12601, N3952, N8907, N8863);
buf BUF1 (N12604, N12597);
buf BUF1 (N12605, N12604);
nor NOR3 (N12606, N12598, N12473, N12275);
nand NAND2 (N12607, N12602, N2695);
buf BUF1 (N12608, N12587);
and AND3 (N12609, N12605, N10827, N8496);
xor XOR2 (N12610, N12595, N8511);
buf BUF1 (N12611, N12608);
buf BUF1 (N12612, N12610);
xor XOR2 (N12613, N12612, N4308);
nand NAND4 (N12614, N12611, N8894, N12547, N3575);
not NOT1 (N12615, N12609);
nand NAND4 (N12616, N12600, N11111, N3829, N955);
nand NAND4 (N12617, N12616, N488, N5855, N7134);
nand NAND4 (N12618, N12615, N5722, N176, N7586);
and AND3 (N12619, N12613, N10304, N8792);
or OR2 (N12620, N12590, N4600);
xor XOR2 (N12621, N12618, N3612);
or OR2 (N12622, N12621, N3151);
xor XOR2 (N12623, N12596, N10845);
buf BUF1 (N12624, N12620);
or OR2 (N12625, N12623, N11711);
and AND4 (N12626, N12603, N7851, N7612, N9091);
xor XOR2 (N12627, N12626, N4254);
buf BUF1 (N12628, N12606);
nor NOR4 (N12629, N12624, N8188, N11393, N5364);
not NOT1 (N12630, N12594);
buf BUF1 (N12631, N12628);
or OR3 (N12632, N12622, N8385, N1031);
and AND2 (N12633, N12619, N160);
not NOT1 (N12634, N12631);
buf BUF1 (N12635, N12617);
buf BUF1 (N12636, N12635);
or OR2 (N12637, N12633, N5001);
buf BUF1 (N12638, N12632);
buf BUF1 (N12639, N12630);
not NOT1 (N12640, N12637);
and AND3 (N12641, N12629, N4892, N4975);
not NOT1 (N12642, N12641);
or OR4 (N12643, N12607, N2473, N5561, N616);
nand NAND4 (N12644, N12640, N8482, N8123, N1465);
not NOT1 (N12645, N12639);
xor XOR2 (N12646, N12627, N11248);
xor XOR2 (N12647, N12646, N10752);
buf BUF1 (N12648, N12644);
buf BUF1 (N12649, N12643);
not NOT1 (N12650, N12649);
and AND2 (N12651, N12625, N9999);
nand NAND3 (N12652, N12636, N9710, N4376);
not NOT1 (N12653, N12650);
and AND2 (N12654, N12614, N10387);
or OR3 (N12655, N12651, N3097, N11020);
nand NAND2 (N12656, N12647, N8939);
or OR2 (N12657, N12634, N1362);
nand NAND4 (N12658, N12645, N5867, N4131, N4174);
nor NOR4 (N12659, N12657, N11114, N12219, N3982);
not NOT1 (N12660, N12652);
nor NOR3 (N12661, N12642, N527, N916);
or OR2 (N12662, N12661, N87);
not NOT1 (N12663, N12659);
xor XOR2 (N12664, N12655, N11939);
buf BUF1 (N12665, N12662);
and AND2 (N12666, N12654, N9356);
nor NOR3 (N12667, N12664, N1980, N8341);
not NOT1 (N12668, N12638);
and AND4 (N12669, N12665, N3364, N5740, N10027);
nor NOR4 (N12670, N12663, N1591, N4009, N2906);
not NOT1 (N12671, N12653);
and AND2 (N12672, N12667, N348);
nor NOR3 (N12673, N12666, N7812, N9077);
and AND2 (N12674, N12672, N12338);
and AND3 (N12675, N12660, N7089, N5586);
buf BUF1 (N12676, N12669);
nor NOR2 (N12677, N12671, N10776);
or OR2 (N12678, N12670, N6326);
nand NAND3 (N12679, N12678, N446, N3818);
nand NAND4 (N12680, N12676, N10242, N11294, N749);
nand NAND2 (N12681, N12648, N6775);
buf BUF1 (N12682, N12675);
nand NAND2 (N12683, N12674, N3275);
or OR2 (N12684, N12683, N12368);
nand NAND2 (N12685, N12684, N3698);
not NOT1 (N12686, N12658);
and AND3 (N12687, N12682, N6207, N6331);
or OR2 (N12688, N12668, N12487);
or OR4 (N12689, N12656, N7954, N7898, N10866);
nand NAND3 (N12690, N12680, N6879, N10407);
not NOT1 (N12691, N12689);
or OR2 (N12692, N12673, N1538);
nand NAND2 (N12693, N12686, N7385);
nand NAND2 (N12694, N12692, N7502);
not NOT1 (N12695, N12677);
nor NOR4 (N12696, N12688, N10491, N5795, N3333);
nor NOR3 (N12697, N12690, N5497, N12161);
and AND3 (N12698, N12695, N1815, N7870);
nor NOR4 (N12699, N12685, N7524, N7700, N3767);
not NOT1 (N12700, N12679);
nor NOR3 (N12701, N12699, N7062, N9344);
buf BUF1 (N12702, N12687);
nand NAND3 (N12703, N12697, N6592, N6583);
and AND4 (N12704, N12694, N6313, N11806, N2426);
not NOT1 (N12705, N12701);
or OR4 (N12706, N12693, N9437, N12476, N1283);
or OR3 (N12707, N12702, N11892, N9868);
or OR4 (N12708, N12700, N4820, N9676, N3950);
nand NAND2 (N12709, N12708, N275);
and AND4 (N12710, N12681, N12226, N4042, N102);
buf BUF1 (N12711, N12704);
not NOT1 (N12712, N12710);
buf BUF1 (N12713, N12711);
buf BUF1 (N12714, N12705);
and AND2 (N12715, N12714, N10856);
and AND4 (N12716, N12703, N9015, N8998, N8391);
nand NAND3 (N12717, N12716, N8812, N1393);
nand NAND3 (N12718, N12715, N444, N6650);
or OR4 (N12719, N12706, N12280, N3403, N7411);
xor XOR2 (N12720, N12718, N324);
or OR4 (N12721, N12696, N2759, N816, N6441);
xor XOR2 (N12722, N12691, N9509);
nand NAND2 (N12723, N12709, N12290);
not NOT1 (N12724, N12712);
xor XOR2 (N12725, N12721, N7352);
nand NAND2 (N12726, N12724, N279);
xor XOR2 (N12727, N12707, N6676);
xor XOR2 (N12728, N12723, N11866);
and AND3 (N12729, N12698, N3205, N11456);
nand NAND2 (N12730, N12720, N8215);
and AND3 (N12731, N12713, N6691, N10277);
and AND4 (N12732, N12726, N2343, N4336, N2510);
not NOT1 (N12733, N12731);
or OR2 (N12734, N12727, N1341);
nand NAND4 (N12735, N12732, N1824, N5132, N12419);
xor XOR2 (N12736, N12717, N9744);
nor NOR3 (N12737, N12729, N6440, N4129);
buf BUF1 (N12738, N12719);
nor NOR4 (N12739, N12735, N2494, N3261, N12112);
buf BUF1 (N12740, N12722);
and AND4 (N12741, N12738, N6802, N2182, N4820);
and AND2 (N12742, N12733, N3874);
xor XOR2 (N12743, N12739, N10478);
and AND3 (N12744, N12743, N9964, N5596);
xor XOR2 (N12745, N12742, N11535);
xor XOR2 (N12746, N12734, N2937);
nor NOR3 (N12747, N12745, N851, N7608);
buf BUF1 (N12748, N12736);
not NOT1 (N12749, N12737);
buf BUF1 (N12750, N12748);
not NOT1 (N12751, N12740);
not NOT1 (N12752, N12749);
or OR2 (N12753, N12744, N4381);
buf BUF1 (N12754, N12746);
nor NOR4 (N12755, N12725, N6856, N11466, N4677);
or OR3 (N12756, N12754, N11490, N4018);
xor XOR2 (N12757, N12730, N11006);
buf BUF1 (N12758, N12751);
nand NAND3 (N12759, N12757, N2071, N5912);
or OR3 (N12760, N12755, N12692, N7194);
xor XOR2 (N12761, N12752, N359);
and AND2 (N12762, N12747, N1807);
xor XOR2 (N12763, N12758, N1911);
or OR4 (N12764, N12762, N5952, N7729, N5158);
xor XOR2 (N12765, N12728, N3598);
buf BUF1 (N12766, N12761);
and AND3 (N12767, N12759, N4181, N2681);
or OR3 (N12768, N12753, N1961, N2216);
nor NOR2 (N12769, N12768, N3970);
xor XOR2 (N12770, N12750, N1941);
buf BUF1 (N12771, N12756);
and AND4 (N12772, N12770, N12093, N1532, N2672);
nand NAND3 (N12773, N12771, N8440, N1559);
buf BUF1 (N12774, N12763);
buf BUF1 (N12775, N12766);
buf BUF1 (N12776, N12764);
xor XOR2 (N12777, N12765, N825);
nor NOR4 (N12778, N12776, N6184, N11461, N2425);
not NOT1 (N12779, N12772);
nand NAND4 (N12780, N12767, N6686, N2316, N3170);
buf BUF1 (N12781, N12769);
and AND4 (N12782, N12773, N9683, N7228, N7756);
nand NAND2 (N12783, N12778, N1357);
and AND2 (N12784, N12777, N9140);
buf BUF1 (N12785, N12781);
nor NOR3 (N12786, N12780, N684, N11105);
buf BUF1 (N12787, N12741);
not NOT1 (N12788, N12786);
or OR2 (N12789, N12774, N1599);
nand NAND3 (N12790, N12782, N7879, N9297);
nor NOR2 (N12791, N12787, N1803);
not NOT1 (N12792, N12760);
nand NAND3 (N12793, N12791, N6737, N3119);
not NOT1 (N12794, N12790);
buf BUF1 (N12795, N12794);
nand NAND3 (N12796, N12793, N11956, N3568);
not NOT1 (N12797, N12779);
nor NOR2 (N12798, N12795, N8961);
and AND3 (N12799, N12792, N9206, N145);
nor NOR3 (N12800, N12798, N2044, N8011);
not NOT1 (N12801, N12788);
nand NAND3 (N12802, N12784, N3002, N8247);
and AND4 (N12803, N12775, N6443, N1546, N2869);
xor XOR2 (N12804, N12800, N10258);
xor XOR2 (N12805, N12785, N9217);
nor NOR2 (N12806, N12797, N9893);
buf BUF1 (N12807, N12796);
buf BUF1 (N12808, N12801);
xor XOR2 (N12809, N12799, N124);
or OR3 (N12810, N12783, N6710, N9240);
nor NOR4 (N12811, N12803, N9688, N4838, N8957);
nor NOR4 (N12812, N12807, N9357, N656, N2099);
nor NOR2 (N12813, N12812, N1581);
xor XOR2 (N12814, N12804, N9259);
buf BUF1 (N12815, N12814);
buf BUF1 (N12816, N12805);
not NOT1 (N12817, N12789);
nand NAND3 (N12818, N12809, N7340, N3028);
and AND4 (N12819, N12813, N778, N2677, N1863);
or OR3 (N12820, N12808, N1810, N9276);
nor NOR3 (N12821, N12819, N12046, N10413);
nor NOR4 (N12822, N12810, N3940, N2167, N1817);
and AND4 (N12823, N12817, N7036, N5386, N7303);
or OR4 (N12824, N12818, N9817, N4926, N6120);
xor XOR2 (N12825, N12816, N10678);
nand NAND2 (N12826, N12823, N9833);
and AND2 (N12827, N12825, N2713);
and AND3 (N12828, N12826, N10323, N10383);
nor NOR4 (N12829, N12821, N9236, N5478, N5900);
nor NOR2 (N12830, N12820, N5356);
nand NAND3 (N12831, N12815, N1, N5544);
nor NOR4 (N12832, N12831, N744, N12773, N8213);
and AND4 (N12833, N12832, N10900, N978, N1390);
nand NAND2 (N12834, N12833, N2525);
not NOT1 (N12835, N12806);
nand NAND4 (N12836, N12811, N6450, N11052, N1637);
not NOT1 (N12837, N12830);
or OR4 (N12838, N12827, N12258, N10315, N2040);
nand NAND4 (N12839, N12835, N4280, N12697, N2934);
buf BUF1 (N12840, N12836);
and AND4 (N12841, N12829, N282, N10300, N8894);
and AND2 (N12842, N12837, N6961);
not NOT1 (N12843, N12828);
not NOT1 (N12844, N12842);
and AND2 (N12845, N12841, N738);
and AND2 (N12846, N12802, N11765);
or OR3 (N12847, N12840, N7555, N8422);
and AND3 (N12848, N12843, N9745, N822);
buf BUF1 (N12849, N12838);
nor NOR3 (N12850, N12824, N9342, N5621);
not NOT1 (N12851, N12839);
buf BUF1 (N12852, N12847);
nand NAND2 (N12853, N12852, N11698);
buf BUF1 (N12854, N12822);
and AND4 (N12855, N12844, N3538, N10884, N10913);
and AND3 (N12856, N12851, N2439, N9792);
xor XOR2 (N12857, N12855, N2432);
and AND2 (N12858, N12848, N2474);
xor XOR2 (N12859, N12856, N11979);
not NOT1 (N12860, N12854);
nand NAND4 (N12861, N12860, N10889, N1702, N5923);
not NOT1 (N12862, N12850);
nor NOR4 (N12863, N12861, N4299, N564, N98);
or OR2 (N12864, N12845, N10851);
nor NOR4 (N12865, N12863, N1161, N742, N1664);
buf BUF1 (N12866, N12862);
buf BUF1 (N12867, N12846);
xor XOR2 (N12868, N12866, N3862);
nand NAND2 (N12869, N12868, N10349);
xor XOR2 (N12870, N12853, N10355);
nor NOR3 (N12871, N12864, N5246, N11645);
nor NOR2 (N12872, N12834, N4129);
and AND3 (N12873, N12869, N10115, N12628);
buf BUF1 (N12874, N12849);
buf BUF1 (N12875, N12872);
nand NAND3 (N12876, N12858, N9390, N7240);
xor XOR2 (N12877, N12875, N10895);
buf BUF1 (N12878, N12859);
not NOT1 (N12879, N12865);
xor XOR2 (N12880, N12878, N1974);
or OR4 (N12881, N12880, N8072, N8773, N2012);
nor NOR4 (N12882, N12874, N10112, N1288, N2558);
nor NOR3 (N12883, N12873, N4366, N6833);
and AND2 (N12884, N12871, N10406);
or OR3 (N12885, N12876, N10193, N7990);
nor NOR3 (N12886, N12882, N5644, N9321);
nand NAND4 (N12887, N12879, N1108, N10779, N8696);
buf BUF1 (N12888, N12867);
and AND3 (N12889, N12870, N8803, N2411);
and AND2 (N12890, N12889, N7472);
buf BUF1 (N12891, N12885);
nand NAND2 (N12892, N12857, N6322);
buf BUF1 (N12893, N12883);
xor XOR2 (N12894, N12891, N12876);
xor XOR2 (N12895, N12893, N11047);
nand NAND2 (N12896, N12881, N10925);
nor NOR4 (N12897, N12888, N11560, N4627, N8591);
and AND4 (N12898, N12896, N12340, N4024, N1461);
buf BUF1 (N12899, N12895);
not NOT1 (N12900, N12886);
nor NOR4 (N12901, N12887, N12106, N3558, N8181);
or OR3 (N12902, N12892, N8856, N9339);
or OR3 (N12903, N12898, N4809, N1756);
nor NOR2 (N12904, N12894, N12392);
buf BUF1 (N12905, N12901);
not NOT1 (N12906, N12904);
not NOT1 (N12907, N12903);
xor XOR2 (N12908, N12899, N10216);
or OR4 (N12909, N12897, N10933, N5122, N5784);
nor NOR3 (N12910, N12909, N9669, N2677);
nand NAND2 (N12911, N12890, N11484);
buf BUF1 (N12912, N12907);
or OR2 (N12913, N12902, N11548);
not NOT1 (N12914, N12910);
nor NOR3 (N12915, N12913, N349, N6917);
nand NAND2 (N12916, N12914, N12648);
or OR2 (N12917, N12908, N11148);
xor XOR2 (N12918, N12916, N10636);
not NOT1 (N12919, N12900);
buf BUF1 (N12920, N12911);
or OR3 (N12921, N12919, N9868, N2825);
nor NOR2 (N12922, N12912, N8874);
or OR4 (N12923, N12922, N6095, N11427, N9811);
nand NAND2 (N12924, N12921, N8354);
nor NOR4 (N12925, N12906, N486, N6134, N6225);
or OR2 (N12926, N12917, N1849);
nand NAND3 (N12927, N12915, N9494, N10339);
buf BUF1 (N12928, N12923);
not NOT1 (N12929, N12926);
xor XOR2 (N12930, N12927, N12229);
nor NOR2 (N12931, N12884, N8411);
nor NOR3 (N12932, N12925, N9122, N11100);
not NOT1 (N12933, N12932);
buf BUF1 (N12934, N12918);
nor NOR3 (N12935, N12877, N7073, N11000);
and AND4 (N12936, N12930, N5417, N7919, N1641);
not NOT1 (N12937, N12936);
xor XOR2 (N12938, N12937, N9197);
not NOT1 (N12939, N12935);
and AND2 (N12940, N12933, N1529);
xor XOR2 (N12941, N12939, N12484);
xor XOR2 (N12942, N12905, N4578);
nand NAND3 (N12943, N12934, N3344, N4516);
not NOT1 (N12944, N12942);
not NOT1 (N12945, N12928);
buf BUF1 (N12946, N12920);
nor NOR4 (N12947, N12929, N3664, N4351, N7040);
nand NAND2 (N12948, N12941, N2242);
and AND2 (N12949, N12948, N6704);
nor NOR2 (N12950, N12924, N4526);
or OR3 (N12951, N12945, N6935, N174);
and AND2 (N12952, N12931, N11149);
nor NOR4 (N12953, N12951, N143, N8926, N512);
nand NAND2 (N12954, N12940, N7087);
buf BUF1 (N12955, N12946);
xor XOR2 (N12956, N12938, N1269);
and AND2 (N12957, N12956, N1234);
nand NAND4 (N12958, N12947, N8189, N4129, N3631);
buf BUF1 (N12959, N12955);
xor XOR2 (N12960, N12957, N3872);
nand NAND2 (N12961, N12950, N1511);
nand NAND2 (N12962, N12960, N11539);
nor NOR2 (N12963, N12954, N11518);
nor NOR2 (N12964, N12959, N6394);
or OR4 (N12965, N12943, N12139, N10398, N438);
and AND2 (N12966, N12944, N7682);
xor XOR2 (N12967, N12958, N7882);
and AND2 (N12968, N12966, N9337);
and AND3 (N12969, N12963, N3754, N5027);
or OR3 (N12970, N12969, N7755, N8406);
xor XOR2 (N12971, N12961, N6594);
nor NOR2 (N12972, N12971, N7715);
not NOT1 (N12973, N12949);
or OR2 (N12974, N12967, N10073);
nand NAND3 (N12975, N12953, N2333, N12435);
or OR2 (N12976, N12970, N1389);
or OR4 (N12977, N12968, N6464, N4293, N6652);
nor NOR2 (N12978, N12964, N10245);
nand NAND3 (N12979, N12974, N3589, N4515);
nor NOR4 (N12980, N12976, N8460, N3374, N870);
xor XOR2 (N12981, N12962, N8555);
buf BUF1 (N12982, N12979);
nor NOR2 (N12983, N12972, N7918);
xor XOR2 (N12984, N12982, N9196);
buf BUF1 (N12985, N12978);
nor NOR3 (N12986, N12965, N8375, N4425);
xor XOR2 (N12987, N12973, N1703);
xor XOR2 (N12988, N12981, N6161);
xor XOR2 (N12989, N12977, N11515);
nor NOR2 (N12990, N12984, N8201);
and AND3 (N12991, N12987, N1679, N2829);
and AND3 (N12992, N12975, N4676, N10003);
nand NAND2 (N12993, N12988, N2033);
nand NAND3 (N12994, N12989, N8173, N8815);
nand NAND4 (N12995, N12993, N11907, N5677, N11523);
or OR2 (N12996, N12992, N3433);
and AND3 (N12997, N12985, N12106, N6924);
not NOT1 (N12998, N12996);
nor NOR4 (N12999, N12991, N194, N3935, N6220);
nor NOR2 (N13000, N12983, N12021);
not NOT1 (N13001, N12994);
or OR2 (N13002, N12990, N5575);
buf BUF1 (N13003, N12986);
nor NOR3 (N13004, N12999, N3565, N2442);
or OR4 (N13005, N13002, N8805, N3388, N10831);
xor XOR2 (N13006, N12997, N202);
or OR2 (N13007, N13000, N187);
or OR3 (N13008, N12952, N6699, N7789);
nand NAND4 (N13009, N13006, N9053, N5273, N718);
or OR4 (N13010, N13001, N4263, N5842, N4183);
buf BUF1 (N13011, N13009);
buf BUF1 (N13012, N12980);
or OR3 (N13013, N13012, N7856, N12338);
or OR2 (N13014, N13005, N9210);
not NOT1 (N13015, N12995);
nand NAND3 (N13016, N13003, N5615, N9138);
nand NAND2 (N13017, N12998, N8784);
nand NAND4 (N13018, N13015, N8376, N8008, N1552);
nand NAND2 (N13019, N13007, N7476);
buf BUF1 (N13020, N13013);
buf BUF1 (N13021, N13014);
and AND4 (N13022, N13004, N11949, N11689, N2250);
nor NOR2 (N13023, N13021, N12705);
xor XOR2 (N13024, N13019, N7555);
or OR4 (N13025, N13024, N1228, N12524, N2500);
nand NAND3 (N13026, N13018, N2977, N1453);
nand NAND4 (N13027, N13025, N3567, N6465, N10466);
not NOT1 (N13028, N13008);
or OR2 (N13029, N13027, N8434);
or OR4 (N13030, N13022, N12708, N862, N10728);
and AND2 (N13031, N13016, N297);
nand NAND2 (N13032, N13011, N7968);
and AND3 (N13033, N13017, N7907, N10315);
nand NAND3 (N13034, N13023, N3045, N9733);
xor XOR2 (N13035, N13028, N2449);
buf BUF1 (N13036, N13030);
and AND2 (N13037, N13031, N1690);
nor NOR4 (N13038, N13034, N11485, N12594, N8521);
nand NAND2 (N13039, N13036, N3559);
and AND2 (N13040, N13035, N10138);
nor NOR2 (N13041, N13010, N2355);
nand NAND2 (N13042, N13041, N9923);
nand NAND3 (N13043, N13020, N2, N2053);
not NOT1 (N13044, N13032);
nor NOR3 (N13045, N13038, N8048, N2060);
buf BUF1 (N13046, N13039);
nor NOR2 (N13047, N13043, N113);
or OR3 (N13048, N13029, N1238, N735);
nand NAND2 (N13049, N13046, N4084);
and AND2 (N13050, N13047, N7985);
or OR4 (N13051, N13048, N10195, N9836, N4211);
nand NAND3 (N13052, N13042, N8160, N5393);
buf BUF1 (N13053, N13051);
or OR3 (N13054, N13050, N12041, N7075);
nor NOR4 (N13055, N13045, N2670, N1865, N1714);
or OR3 (N13056, N13040, N7469, N2306);
and AND3 (N13057, N13054, N3112, N8691);
not NOT1 (N13058, N13037);
xor XOR2 (N13059, N13056, N10425);
nand NAND4 (N13060, N13055, N837, N9256, N3558);
not NOT1 (N13061, N13057);
xor XOR2 (N13062, N13058, N11169);
and AND4 (N13063, N13044, N10554, N3882, N1282);
not NOT1 (N13064, N13060);
nand NAND4 (N13065, N13053, N4306, N9572, N8420);
xor XOR2 (N13066, N13033, N12069);
xor XOR2 (N13067, N13064, N12984);
or OR3 (N13068, N13026, N3333, N4642);
or OR3 (N13069, N13049, N5281, N5079);
not NOT1 (N13070, N13067);
buf BUF1 (N13071, N13062);
buf BUF1 (N13072, N13071);
buf BUF1 (N13073, N13066);
and AND3 (N13074, N13052, N3497, N9031);
xor XOR2 (N13075, N13068, N9057);
not NOT1 (N13076, N13073);
or OR3 (N13077, N13063, N5002, N9047);
or OR4 (N13078, N13072, N2329, N2820, N7318);
not NOT1 (N13079, N13076);
nor NOR2 (N13080, N13078, N8089);
not NOT1 (N13081, N13061);
and AND3 (N13082, N13081, N11016, N8641);
or OR4 (N13083, N13082, N8396, N5745, N9391);
nor NOR3 (N13084, N13059, N3766, N661);
or OR3 (N13085, N13069, N1629, N10623);
not NOT1 (N13086, N13083);
nand NAND3 (N13087, N13077, N11146, N10266);
and AND4 (N13088, N13079, N10844, N11033, N4140);
and AND3 (N13089, N13070, N3085, N1838);
nor NOR3 (N13090, N13086, N8512, N9117);
and AND4 (N13091, N13080, N12112, N3556, N2357);
buf BUF1 (N13092, N13075);
nand NAND3 (N13093, N13074, N12133, N3511);
nor NOR2 (N13094, N13065, N5919);
nand NAND3 (N13095, N13087, N3589, N9118);
and AND2 (N13096, N13093, N6317);
nor NOR2 (N13097, N13089, N8210);
buf BUF1 (N13098, N13097);
buf BUF1 (N13099, N13090);
or OR2 (N13100, N13092, N11423);
or OR2 (N13101, N13096, N1460);
and AND4 (N13102, N13084, N11797, N12814, N10364);
or OR2 (N13103, N13088, N9837);
nor NOR2 (N13104, N13098, N6094);
and AND4 (N13105, N13099, N86, N4906, N9312);
and AND4 (N13106, N13095, N2492, N8511, N3720);
buf BUF1 (N13107, N13091);
or OR2 (N13108, N13105, N7265);
nor NOR4 (N13109, N13106, N443, N9423, N2051);
buf BUF1 (N13110, N13094);
or OR2 (N13111, N13107, N12581);
xor XOR2 (N13112, N13101, N3139);
nor NOR2 (N13113, N13103, N1971);
xor XOR2 (N13114, N13112, N7577);
xor XOR2 (N13115, N13108, N10505);
nor NOR3 (N13116, N13114, N8845, N102);
and AND4 (N13117, N13111, N5189, N2348, N4180);
and AND3 (N13118, N13110, N5959, N12173);
xor XOR2 (N13119, N13104, N1333);
and AND4 (N13120, N13113, N7109, N4384, N9323);
nor NOR2 (N13121, N13120, N6875);
xor XOR2 (N13122, N13115, N11317);
nand NAND3 (N13123, N13102, N758, N5017);
nand NAND3 (N13124, N13100, N7144, N2119);
nand NAND2 (N13125, N13119, N8363);
nor NOR2 (N13126, N13124, N177);
xor XOR2 (N13127, N13122, N2375);
or OR4 (N13128, N13125, N5479, N4055, N6939);
nor NOR3 (N13129, N13085, N4787, N3072);
buf BUF1 (N13130, N13129);
or OR2 (N13131, N13127, N1930);
nor NOR4 (N13132, N13118, N5500, N9943, N1843);
nor NOR3 (N13133, N13109, N7724, N9004);
not NOT1 (N13134, N13126);
not NOT1 (N13135, N13130);
nand NAND4 (N13136, N13123, N8163, N906, N7812);
nand NAND2 (N13137, N13132, N3606);
not NOT1 (N13138, N13137);
nor NOR4 (N13139, N13121, N9779, N9623, N8073);
or OR2 (N13140, N13128, N4223);
and AND4 (N13141, N13133, N839, N7082, N1034);
and AND2 (N13142, N13117, N4011);
nand NAND4 (N13143, N13135, N2128, N4199, N6679);
nand NAND3 (N13144, N13139, N3009, N12348);
buf BUF1 (N13145, N13144);
xor XOR2 (N13146, N13131, N5157);
buf BUF1 (N13147, N13134);
nor NOR3 (N13148, N13141, N5709, N4504);
and AND3 (N13149, N13147, N11014, N4741);
not NOT1 (N13150, N13142);
xor XOR2 (N13151, N13148, N3322);
buf BUF1 (N13152, N13146);
buf BUF1 (N13153, N13143);
nand NAND3 (N13154, N13151, N8570, N3045);
buf BUF1 (N13155, N13149);
nand NAND3 (N13156, N13145, N11084, N11316);
nand NAND2 (N13157, N13155, N5644);
nor NOR4 (N13158, N13153, N7534, N935, N6676);
xor XOR2 (N13159, N13136, N8344);
nor NOR2 (N13160, N13138, N12286);
xor XOR2 (N13161, N13150, N12289);
xor XOR2 (N13162, N13140, N6382);
nor NOR4 (N13163, N13116, N7775, N9187, N949);
xor XOR2 (N13164, N13156, N11730);
xor XOR2 (N13165, N13158, N8261);
nand NAND4 (N13166, N13154, N6499, N6232, N3476);
not NOT1 (N13167, N13164);
and AND3 (N13168, N13166, N11307, N2496);
not NOT1 (N13169, N13168);
or OR3 (N13170, N13169, N4391, N3909);
and AND3 (N13171, N13159, N12110, N6999);
nand NAND3 (N13172, N13165, N9944, N165);
nor NOR2 (N13173, N13161, N7257);
xor XOR2 (N13174, N13170, N5178);
buf BUF1 (N13175, N13167);
nand NAND3 (N13176, N13160, N11603, N6078);
nor NOR2 (N13177, N13152, N460);
or OR3 (N13178, N13173, N876, N12026);
nand NAND4 (N13179, N13178, N4313, N6934, N2019);
or OR3 (N13180, N13172, N11604, N9544);
nand NAND3 (N13181, N13162, N8089, N9953);
nand NAND2 (N13182, N13163, N7975);
or OR4 (N13183, N13175, N8347, N8842, N10794);
buf BUF1 (N13184, N13176);
and AND3 (N13185, N13179, N7162, N5636);
or OR3 (N13186, N13180, N6690, N6208);
buf BUF1 (N13187, N13184);
and AND2 (N13188, N13181, N10000);
buf BUF1 (N13189, N13177);
nand NAND3 (N13190, N13171, N10163, N12793);
and AND2 (N13191, N13182, N11960);
xor XOR2 (N13192, N13185, N10733);
nor NOR3 (N13193, N13174, N9577, N3802);
not NOT1 (N13194, N13191);
buf BUF1 (N13195, N13193);
buf BUF1 (N13196, N13183);
nand NAND3 (N13197, N13188, N12111, N5142);
not NOT1 (N13198, N13186);
xor XOR2 (N13199, N13192, N8695);
and AND2 (N13200, N13199, N5166);
or OR3 (N13201, N13190, N11647, N775);
not NOT1 (N13202, N13189);
nor NOR3 (N13203, N13200, N3566, N11008);
nor NOR3 (N13204, N13195, N7827, N11857);
buf BUF1 (N13205, N13202);
nor NOR3 (N13206, N13196, N2134, N299);
nor NOR3 (N13207, N13198, N6342, N628);
or OR3 (N13208, N13206, N1604, N12976);
buf BUF1 (N13209, N13157);
buf BUF1 (N13210, N13201);
nor NOR2 (N13211, N13204, N702);
xor XOR2 (N13212, N13211, N9932);
buf BUF1 (N13213, N13187);
and AND3 (N13214, N13209, N8454, N10513);
buf BUF1 (N13215, N13214);
not NOT1 (N13216, N13208);
and AND3 (N13217, N13212, N7942, N10832);
and AND2 (N13218, N13194, N7202);
or OR4 (N13219, N13203, N3241, N4781, N12304);
and AND2 (N13220, N13197, N11819);
and AND4 (N13221, N13210, N7245, N6854, N7820);
buf BUF1 (N13222, N13213);
xor XOR2 (N13223, N13207, N2318);
or OR2 (N13224, N13216, N2043);
buf BUF1 (N13225, N13218);
buf BUF1 (N13226, N13219);
and AND4 (N13227, N13220, N5154, N8487, N2700);
not NOT1 (N13228, N13226);
buf BUF1 (N13229, N13228);
nor NOR2 (N13230, N13217, N3053);
nor NOR4 (N13231, N13224, N4814, N7310, N4629);
not NOT1 (N13232, N13221);
buf BUF1 (N13233, N13222);
nor NOR4 (N13234, N13233, N10936, N2414, N9135);
and AND4 (N13235, N13231, N7063, N9207, N12997);
nor NOR3 (N13236, N13205, N3916, N6293);
or OR2 (N13237, N13236, N4308);
buf BUF1 (N13238, N13225);
or OR2 (N13239, N13227, N2352);
buf BUF1 (N13240, N13234);
or OR3 (N13241, N13229, N1569, N7740);
xor XOR2 (N13242, N13223, N10208);
or OR3 (N13243, N13232, N8044, N12515);
not NOT1 (N13244, N13215);
or OR2 (N13245, N13242, N3739);
or OR3 (N13246, N13243, N10455, N1222);
xor XOR2 (N13247, N13237, N5632);
or OR2 (N13248, N13240, N4238);
buf BUF1 (N13249, N13245);
xor XOR2 (N13250, N13241, N879);
nand NAND2 (N13251, N13230, N9429);
xor XOR2 (N13252, N13249, N8515);
not NOT1 (N13253, N13238);
nand NAND4 (N13254, N13252, N2077, N9581, N8212);
buf BUF1 (N13255, N13244);
nor NOR2 (N13256, N13247, N4604);
xor XOR2 (N13257, N13235, N2295);
nor NOR3 (N13258, N13257, N10177, N11648);
buf BUF1 (N13259, N13250);
xor XOR2 (N13260, N13253, N8185);
or OR2 (N13261, N13254, N3577);
and AND4 (N13262, N13256, N4010, N947, N449);
nor NOR2 (N13263, N13260, N10072);
nor NOR3 (N13264, N13239, N2627, N1470);
not NOT1 (N13265, N13255);
xor XOR2 (N13266, N13264, N7499);
buf BUF1 (N13267, N13246);
nand NAND4 (N13268, N13267, N8300, N5610, N6901);
nand NAND3 (N13269, N13265, N9834, N1097);
not NOT1 (N13270, N13258);
and AND3 (N13271, N13251, N7919, N10916);
nand NAND3 (N13272, N13268, N1070, N8550);
xor XOR2 (N13273, N13266, N3748);
nor NOR2 (N13274, N13248, N7629);
and AND3 (N13275, N13259, N8132, N7517);
or OR2 (N13276, N13270, N12844);
or OR3 (N13277, N13276, N1370, N13021);
nor NOR2 (N13278, N13277, N7408);
xor XOR2 (N13279, N13271, N7484);
buf BUF1 (N13280, N13278);
buf BUF1 (N13281, N13280);
or OR2 (N13282, N13275, N9449);
nand NAND3 (N13283, N13281, N3796, N3884);
nand NAND3 (N13284, N13283, N12608, N10727);
buf BUF1 (N13285, N13272);
and AND3 (N13286, N13262, N7486, N160);
nor NOR2 (N13287, N13261, N6678);
xor XOR2 (N13288, N13287, N2981);
or OR2 (N13289, N13288, N6945);
or OR4 (N13290, N13284, N7946, N2403, N5005);
buf BUF1 (N13291, N13285);
buf BUF1 (N13292, N13263);
not NOT1 (N13293, N13269);
nor NOR3 (N13294, N13292, N13109, N9265);
nand NAND2 (N13295, N13294, N13228);
nand NAND4 (N13296, N13273, N1632, N4057, N3329);
nand NAND4 (N13297, N13295, N9435, N1295, N9662);
and AND4 (N13298, N13296, N851, N5592, N383);
nand NAND4 (N13299, N13298, N1686, N7357, N7223);
or OR2 (N13300, N13279, N12009);
nand NAND4 (N13301, N13293, N4561, N4112, N5069);
or OR4 (N13302, N13289, N5544, N7777, N9569);
buf BUF1 (N13303, N13302);
not NOT1 (N13304, N13282);
buf BUF1 (N13305, N13286);
not NOT1 (N13306, N13297);
buf BUF1 (N13307, N13291);
and AND4 (N13308, N13301, N10102, N4037, N526);
or OR2 (N13309, N13308, N1925);
not NOT1 (N13310, N13303);
buf BUF1 (N13311, N13307);
or OR4 (N13312, N13300, N6037, N11401, N9685);
or OR2 (N13313, N13290, N4);
or OR2 (N13314, N13311, N299);
xor XOR2 (N13315, N13310, N7273);
or OR4 (N13316, N13304, N4457, N752, N5708);
nand NAND3 (N13317, N13309, N5878, N5724);
buf BUF1 (N13318, N13312);
nor NOR3 (N13319, N13306, N12144, N10137);
buf BUF1 (N13320, N13317);
xor XOR2 (N13321, N13274, N12452);
nor NOR3 (N13322, N13318, N11957, N12072);
not NOT1 (N13323, N13320);
or OR3 (N13324, N13299, N1907, N1859);
or OR4 (N13325, N13315, N3941, N1417, N7794);
not NOT1 (N13326, N13325);
buf BUF1 (N13327, N13323);
nor NOR4 (N13328, N13305, N2463, N9352, N2331);
buf BUF1 (N13329, N13324);
nand NAND3 (N13330, N13316, N7257, N4514);
not NOT1 (N13331, N13329);
nand NAND2 (N13332, N13330, N8666);
buf BUF1 (N13333, N13313);
not NOT1 (N13334, N13327);
xor XOR2 (N13335, N13319, N12008);
nand NAND3 (N13336, N13331, N6854, N5523);
nor NOR2 (N13337, N13328, N2837);
buf BUF1 (N13338, N13326);
not NOT1 (N13339, N13335);
or OR3 (N13340, N13322, N11547, N8502);
not NOT1 (N13341, N13336);
or OR2 (N13342, N13333, N10968);
not NOT1 (N13343, N13332);
or OR2 (N13344, N13343, N13254);
not NOT1 (N13345, N13340);
or OR3 (N13346, N13337, N12970, N2469);
or OR2 (N13347, N13346, N11877);
or OR4 (N13348, N13338, N10472, N934, N8085);
buf BUF1 (N13349, N13342);
and AND4 (N13350, N13349, N11322, N12952, N6897);
or OR3 (N13351, N13334, N9536, N4391);
xor XOR2 (N13352, N13350, N12284);
xor XOR2 (N13353, N13341, N2525);
buf BUF1 (N13354, N13351);
and AND3 (N13355, N13348, N2279, N10714);
or OR3 (N13356, N13339, N2133, N12046);
nand NAND3 (N13357, N13355, N4474, N2975);
and AND4 (N13358, N13357, N12183, N4235, N51);
nor NOR4 (N13359, N13344, N6092, N9507, N4610);
xor XOR2 (N13360, N13359, N11967);
nand NAND2 (N13361, N13360, N12364);
nor NOR2 (N13362, N13361, N3085);
and AND2 (N13363, N13354, N7944);
xor XOR2 (N13364, N13347, N2184);
buf BUF1 (N13365, N13362);
nor NOR4 (N13366, N13358, N11849, N719, N352);
nand NAND4 (N13367, N13356, N1539, N8373, N10613);
buf BUF1 (N13368, N13366);
nor NOR4 (N13369, N13345, N10064, N7702, N4756);
nor NOR3 (N13370, N13364, N6667, N7935);
nor NOR3 (N13371, N13370, N8238, N4658);
nor NOR3 (N13372, N13369, N10359, N4037);
not NOT1 (N13373, N13368);
and AND3 (N13374, N13352, N12187, N1751);
nand NAND2 (N13375, N13367, N976);
not NOT1 (N13376, N13372);
buf BUF1 (N13377, N13376);
buf BUF1 (N13378, N13373);
buf BUF1 (N13379, N13374);
or OR4 (N13380, N13321, N5020, N2528, N136);
buf BUF1 (N13381, N13365);
nor NOR3 (N13382, N13380, N1379, N2108);
nand NAND4 (N13383, N13363, N1411, N906, N8922);
xor XOR2 (N13384, N13375, N8666);
xor XOR2 (N13385, N13383, N9987);
nand NAND2 (N13386, N13384, N2515);
and AND2 (N13387, N13382, N9783);
buf BUF1 (N13388, N13385);
xor XOR2 (N13389, N13379, N2446);
not NOT1 (N13390, N13389);
xor XOR2 (N13391, N13371, N13057);
nor NOR4 (N13392, N13377, N117, N4420, N12694);
nor NOR2 (N13393, N13378, N4871);
and AND3 (N13394, N13390, N11785, N6688);
nor NOR4 (N13395, N13381, N3779, N2446, N5014);
xor XOR2 (N13396, N13391, N12720);
xor XOR2 (N13397, N13353, N6979);
xor XOR2 (N13398, N13394, N255);
and AND3 (N13399, N13386, N1330, N12947);
xor XOR2 (N13400, N13388, N10773);
nor NOR2 (N13401, N13392, N8975);
or OR3 (N13402, N13393, N446, N8384);
buf BUF1 (N13403, N13400);
buf BUF1 (N13404, N13314);
not NOT1 (N13405, N13387);
and AND3 (N13406, N13395, N6667, N6074);
and AND4 (N13407, N13403, N13315, N2160, N8985);
and AND2 (N13408, N13397, N6081);
buf BUF1 (N13409, N13404);
not NOT1 (N13410, N13398);
buf BUF1 (N13411, N13406);
nor NOR2 (N13412, N13408, N5945);
not NOT1 (N13413, N13409);
and AND4 (N13414, N13410, N11844, N2837, N2467);
buf BUF1 (N13415, N13407);
nand NAND2 (N13416, N13396, N4845);
nand NAND4 (N13417, N13399, N11984, N4270, N9729);
xor XOR2 (N13418, N13417, N5131);
nand NAND2 (N13419, N13418, N9430);
and AND2 (N13420, N13419, N8423);
buf BUF1 (N13421, N13413);
buf BUF1 (N13422, N13402);
nand NAND4 (N13423, N13401, N13385, N10660, N4729);
and AND4 (N13424, N13405, N2108, N7279, N11771);
not NOT1 (N13425, N13424);
buf BUF1 (N13426, N13421);
not NOT1 (N13427, N13411);
and AND3 (N13428, N13423, N5068, N10318);
not NOT1 (N13429, N13428);
not NOT1 (N13430, N13427);
xor XOR2 (N13431, N13422, N2521);
not NOT1 (N13432, N13426);
nor NOR4 (N13433, N13415, N8759, N6937, N7348);
and AND2 (N13434, N13432, N7126);
not NOT1 (N13435, N13412);
nor NOR4 (N13436, N13414, N7657, N2450, N4544);
not NOT1 (N13437, N13435);
or OR2 (N13438, N13429, N8454);
nor NOR4 (N13439, N13416, N10139, N12376, N2260);
nor NOR4 (N13440, N13431, N2978, N8659, N6483);
and AND4 (N13441, N13438, N10743, N7772, N2102);
nand NAND3 (N13442, N13433, N9222, N6272);
not NOT1 (N13443, N13441);
nand NAND2 (N13444, N13425, N12122);
and AND3 (N13445, N13442, N12836, N11105);
nand NAND4 (N13446, N13436, N6812, N4991, N13401);
nand NAND2 (N13447, N13440, N13411);
nand NAND4 (N13448, N13437, N10708, N10480, N5279);
nand NAND2 (N13449, N13420, N2138);
and AND4 (N13450, N13439, N7007, N836, N5271);
xor XOR2 (N13451, N13446, N9701);
nand NAND3 (N13452, N13443, N4465, N3123);
or OR2 (N13453, N13430, N11776);
buf BUF1 (N13454, N13453);
nand NAND2 (N13455, N13449, N12074);
nor NOR2 (N13456, N13447, N1206);
xor XOR2 (N13457, N13444, N5626);
buf BUF1 (N13458, N13454);
nand NAND2 (N13459, N13434, N10662);
nor NOR3 (N13460, N13459, N9531, N7304);
and AND3 (N13461, N13452, N9711, N12339);
buf BUF1 (N13462, N13450);
xor XOR2 (N13463, N13445, N11477);
not NOT1 (N13464, N13458);
and AND3 (N13465, N13461, N10470, N2137);
nor NOR4 (N13466, N13464, N7438, N12787, N1348);
xor XOR2 (N13467, N13451, N12901);
and AND4 (N13468, N13465, N9884, N13215, N2657);
nand NAND3 (N13469, N13463, N6877, N4149);
or OR3 (N13470, N13466, N7305, N3094);
not NOT1 (N13471, N13448);
buf BUF1 (N13472, N13456);
or OR3 (N13473, N13469, N3202, N3284);
buf BUF1 (N13474, N13468);
and AND4 (N13475, N13457, N1582, N2666, N4792);
and AND4 (N13476, N13473, N5261, N11921, N6118);
or OR4 (N13477, N13474, N3967, N6118, N7970);
nand NAND4 (N13478, N13472, N731, N10238, N9628);
nand NAND4 (N13479, N13455, N1695, N12174, N8446);
nor NOR2 (N13480, N13476, N13010);
nor NOR3 (N13481, N13471, N1431, N7580);
not NOT1 (N13482, N13470);
or OR2 (N13483, N13460, N4641);
buf BUF1 (N13484, N13475);
and AND4 (N13485, N13480, N7803, N12328, N8526);
not NOT1 (N13486, N13481);
buf BUF1 (N13487, N13486);
nand NAND3 (N13488, N13479, N6348, N6617);
and AND4 (N13489, N13482, N1976, N1973, N7276);
or OR2 (N13490, N13489, N6492);
xor XOR2 (N13491, N13484, N7556);
xor XOR2 (N13492, N13485, N10777);
nor NOR3 (N13493, N13491, N12364, N5996);
nor NOR3 (N13494, N13462, N11618, N2632);
xor XOR2 (N13495, N13483, N3573);
xor XOR2 (N13496, N13478, N5165);
or OR4 (N13497, N13490, N12250, N10224, N2647);
and AND4 (N13498, N13493, N2128, N2219, N7141);
or OR4 (N13499, N13496, N10922, N9499, N12503);
buf BUF1 (N13500, N13467);
buf BUF1 (N13501, N13495);
buf BUF1 (N13502, N13497);
nor NOR2 (N13503, N13488, N9862);
or OR4 (N13504, N13502, N8855, N4345, N5795);
not NOT1 (N13505, N13498);
nor NOR4 (N13506, N13504, N3655, N4534, N12978);
and AND3 (N13507, N13506, N4632, N12976);
and AND3 (N13508, N13505, N11534, N223);
xor XOR2 (N13509, N13500, N6902);
nand NAND2 (N13510, N13503, N12103);
xor XOR2 (N13511, N13499, N12491);
and AND2 (N13512, N13494, N12439);
or OR2 (N13513, N13507, N9758);
xor XOR2 (N13514, N13487, N12827);
and AND4 (N13515, N13513, N4539, N1361, N2651);
xor XOR2 (N13516, N13477, N7375);
buf BUF1 (N13517, N13510);
xor XOR2 (N13518, N13516, N8481);
nor NOR3 (N13519, N13515, N7545, N7400);
not NOT1 (N13520, N13492);
nor NOR2 (N13521, N13501, N1547);
not NOT1 (N13522, N13518);
xor XOR2 (N13523, N13514, N5390);
or OR2 (N13524, N13519, N2369);
nand NAND3 (N13525, N13512, N5132, N12727);
nor NOR3 (N13526, N13520, N4537, N13092);
and AND3 (N13527, N13509, N4784, N3516);
xor XOR2 (N13528, N13525, N1342);
nand NAND2 (N13529, N13517, N8724);
not NOT1 (N13530, N13523);
buf BUF1 (N13531, N13524);
and AND4 (N13532, N13508, N13142, N10306, N5291);
xor XOR2 (N13533, N13532, N5708);
xor XOR2 (N13534, N13521, N10133);
nor NOR3 (N13535, N13534, N9890, N587);
buf BUF1 (N13536, N13511);
buf BUF1 (N13537, N13527);
or OR2 (N13538, N13537, N1487);
xor XOR2 (N13539, N13531, N10855);
nor NOR4 (N13540, N13522, N6193, N2056, N3043);
xor XOR2 (N13541, N13539, N9599);
nand NAND3 (N13542, N13533, N11475, N1930);
or OR2 (N13543, N13526, N2221);
and AND4 (N13544, N13542, N10589, N3774, N11275);
and AND4 (N13545, N13528, N4680, N12218, N12566);
or OR2 (N13546, N13543, N6989);
buf BUF1 (N13547, N13538);
xor XOR2 (N13548, N13535, N10676);
or OR4 (N13549, N13536, N6729, N9388, N10267);
xor XOR2 (N13550, N13540, N8059);
buf BUF1 (N13551, N13546);
or OR4 (N13552, N13545, N11090, N11036, N9041);
xor XOR2 (N13553, N13552, N6231);
or OR4 (N13554, N13547, N658, N4899, N8996);
not NOT1 (N13555, N13541);
xor XOR2 (N13556, N13555, N4709);
buf BUF1 (N13557, N13549);
xor XOR2 (N13558, N13530, N7820);
nor NOR2 (N13559, N13551, N5061);
xor XOR2 (N13560, N13548, N2999);
not NOT1 (N13561, N13558);
and AND4 (N13562, N13553, N2045, N4140, N6575);
buf BUF1 (N13563, N13559);
xor XOR2 (N13564, N13554, N8875);
nor NOR3 (N13565, N13562, N7370, N6170);
nor NOR2 (N13566, N13563, N906);
xor XOR2 (N13567, N13529, N3782);
buf BUF1 (N13568, N13567);
buf BUF1 (N13569, N13560);
xor XOR2 (N13570, N13561, N12873);
nand NAND4 (N13571, N13565, N598, N8440, N4924);
or OR2 (N13572, N13556, N6755);
and AND4 (N13573, N13570, N2611, N9305, N11570);
and AND4 (N13574, N13571, N13421, N13134, N9209);
nor NOR3 (N13575, N13568, N969, N6577);
or OR2 (N13576, N13575, N13132);
not NOT1 (N13577, N13574);
xor XOR2 (N13578, N13572, N9234);
nand NAND2 (N13579, N13569, N9371);
not NOT1 (N13580, N13550);
buf BUF1 (N13581, N13573);
xor XOR2 (N13582, N13579, N5769);
nor NOR3 (N13583, N13544, N12364, N8867);
nand NAND4 (N13584, N13566, N3815, N5330, N8493);
nand NAND4 (N13585, N13584, N11846, N10756, N3369);
buf BUF1 (N13586, N13577);
buf BUF1 (N13587, N13583);
nand NAND4 (N13588, N13578, N7374, N8245, N12236);
not NOT1 (N13589, N13557);
and AND3 (N13590, N13586, N4747, N4825);
not NOT1 (N13591, N13564);
not NOT1 (N13592, N13590);
buf BUF1 (N13593, N13580);
nand NAND4 (N13594, N13581, N4807, N5663, N233);
or OR2 (N13595, N13592, N6638);
nand NAND3 (N13596, N13585, N13268, N3328);
xor XOR2 (N13597, N13582, N4320);
nand NAND2 (N13598, N13587, N1547);
nor NOR4 (N13599, N13595, N3259, N6998, N6092);
buf BUF1 (N13600, N13576);
buf BUF1 (N13601, N13594);
and AND3 (N13602, N13596, N9506, N8399);
xor XOR2 (N13603, N13597, N11842);
buf BUF1 (N13604, N13598);
nor NOR2 (N13605, N13589, N12792);
xor XOR2 (N13606, N13604, N4716);
not NOT1 (N13607, N13602);
or OR4 (N13608, N13603, N6975, N11157, N421);
nand NAND4 (N13609, N13593, N7867, N11206, N10080);
nand NAND3 (N13610, N13609, N10044, N1318);
or OR3 (N13611, N13605, N6340, N6370);
not NOT1 (N13612, N13606);
not NOT1 (N13613, N13599);
xor XOR2 (N13614, N13591, N9495);
not NOT1 (N13615, N13613);
nand NAND3 (N13616, N13615, N5514, N12230);
nor NOR3 (N13617, N13600, N83, N7386);
and AND2 (N13618, N13601, N11219);
xor XOR2 (N13619, N13610, N835);
buf BUF1 (N13620, N13617);
and AND3 (N13621, N13616, N6494, N12861);
buf BUF1 (N13622, N13611);
buf BUF1 (N13623, N13608);
nor NOR4 (N13624, N13619, N7059, N7797, N4648);
not NOT1 (N13625, N13622);
and AND2 (N13626, N13623, N1042);
nand NAND2 (N13627, N13626, N4968);
nand NAND3 (N13628, N13614, N5693, N13466);
not NOT1 (N13629, N13627);
or OR4 (N13630, N13629, N11761, N12797, N13037);
xor XOR2 (N13631, N13618, N9394);
xor XOR2 (N13632, N13621, N10431);
or OR4 (N13633, N13631, N1095, N1173, N516);
nand NAND3 (N13634, N13588, N6189, N12868);
nor NOR4 (N13635, N13624, N10750, N4776, N7212);
nor NOR4 (N13636, N13628, N356, N6846, N7672);
and AND3 (N13637, N13620, N9873, N1807);
not NOT1 (N13638, N13633);
nand NAND3 (N13639, N13607, N1921, N420);
or OR2 (N13640, N13630, N5598);
nor NOR4 (N13641, N13635, N7728, N3765, N402);
xor XOR2 (N13642, N13640, N1473);
and AND2 (N13643, N13638, N9450);
buf BUF1 (N13644, N13612);
xor XOR2 (N13645, N13636, N1346);
xor XOR2 (N13646, N13643, N6867);
buf BUF1 (N13647, N13634);
and AND2 (N13648, N13641, N12964);
nor NOR4 (N13649, N13637, N12163, N10131, N4494);
xor XOR2 (N13650, N13639, N12637);
or OR2 (N13651, N13647, N9583);
or OR2 (N13652, N13625, N13198);
buf BUF1 (N13653, N13632);
buf BUF1 (N13654, N13649);
or OR2 (N13655, N13642, N4296);
nor NOR3 (N13656, N13645, N1991, N6969);
not NOT1 (N13657, N13653);
nand NAND4 (N13658, N13655, N10276, N4957, N4729);
and AND2 (N13659, N13657, N643);
nor NOR3 (N13660, N13656, N12935, N13137);
and AND4 (N13661, N13660, N12678, N13257, N10405);
xor XOR2 (N13662, N13659, N5192);
not NOT1 (N13663, N13646);
nand NAND4 (N13664, N13661, N10576, N11314, N4971);
not NOT1 (N13665, N13644);
or OR2 (N13666, N13652, N11272);
and AND2 (N13667, N13651, N8504);
or OR2 (N13668, N13654, N4346);
xor XOR2 (N13669, N13658, N8053);
xor XOR2 (N13670, N13662, N9721);
or OR2 (N13671, N13668, N1189);
not NOT1 (N13672, N13648);
nand NAND2 (N13673, N13670, N23);
not NOT1 (N13674, N13666);
nand NAND3 (N13675, N13672, N7057, N5393);
or OR3 (N13676, N13664, N8441, N1998);
not NOT1 (N13677, N13650);
nor NOR3 (N13678, N13669, N12761, N3620);
buf BUF1 (N13679, N13677);
or OR4 (N13680, N13673, N3154, N3707, N3500);
nor NOR3 (N13681, N13676, N3715, N8072);
nand NAND2 (N13682, N13681, N10544);
buf BUF1 (N13683, N13671);
or OR3 (N13684, N13679, N13112, N10978);
not NOT1 (N13685, N13663);
nor NOR3 (N13686, N13682, N11935, N3030);
not NOT1 (N13687, N13674);
xor XOR2 (N13688, N13678, N4727);
xor XOR2 (N13689, N13688, N7396);
and AND2 (N13690, N13689, N2274);
and AND4 (N13691, N13685, N54, N7028, N12243);
nor NOR3 (N13692, N13691, N13250, N9073);
buf BUF1 (N13693, N13680);
buf BUF1 (N13694, N13690);
not NOT1 (N13695, N13684);
or OR3 (N13696, N13675, N12270, N1057);
not NOT1 (N13697, N13692);
not NOT1 (N13698, N13693);
nand NAND4 (N13699, N13697, N8962, N8125, N7816);
xor XOR2 (N13700, N13696, N1537);
xor XOR2 (N13701, N13700, N8058);
buf BUF1 (N13702, N13699);
and AND2 (N13703, N13686, N9997);
nor NOR4 (N13704, N13694, N1058, N6605, N9221);
or OR3 (N13705, N13701, N9616, N9120);
nand NAND4 (N13706, N13703, N5755, N11272, N5962);
buf BUF1 (N13707, N13687);
or OR3 (N13708, N13704, N5538, N8706);
and AND4 (N13709, N13698, N6498, N12537, N3772);
nor NOR4 (N13710, N13708, N8807, N2234, N8531);
nand NAND4 (N13711, N13710, N8950, N10384, N3479);
buf BUF1 (N13712, N13695);
nor NOR2 (N13713, N13709, N11192);
nand NAND4 (N13714, N13667, N2005, N4633, N9884);
and AND3 (N13715, N13714, N2271, N11468);
not NOT1 (N13716, N13713);
buf BUF1 (N13717, N13702);
and AND4 (N13718, N13665, N5319, N1324, N12765);
buf BUF1 (N13719, N13717);
nor NOR2 (N13720, N13683, N2558);
and AND3 (N13721, N13715, N44, N7409);
xor XOR2 (N13722, N13719, N3346);
nor NOR4 (N13723, N13705, N4121, N5880, N3230);
or OR3 (N13724, N13716, N12438, N11268);
nor NOR2 (N13725, N13722, N10449);
xor XOR2 (N13726, N13718, N7991);
and AND4 (N13727, N13711, N7171, N4826, N1254);
nand NAND2 (N13728, N13726, N5752);
and AND3 (N13729, N13728, N7225, N73);
buf BUF1 (N13730, N13707);
not NOT1 (N13731, N13724);
or OR2 (N13732, N13720, N13323);
not NOT1 (N13733, N13706);
nor NOR2 (N13734, N13731, N1295);
nor NOR2 (N13735, N13730, N4112);
and AND4 (N13736, N13721, N13135, N6473, N10754);
xor XOR2 (N13737, N13736, N2657);
xor XOR2 (N13738, N13737, N10874);
not NOT1 (N13739, N13727);
or OR3 (N13740, N13729, N11490, N392);
or OR3 (N13741, N13733, N12094, N8648);
nor NOR2 (N13742, N13725, N5729);
buf BUF1 (N13743, N13742);
buf BUF1 (N13744, N13735);
or OR4 (N13745, N13712, N2694, N7900, N1677);
buf BUF1 (N13746, N13739);
nand NAND3 (N13747, N13723, N5970, N3654);
xor XOR2 (N13748, N13746, N4764);
not NOT1 (N13749, N13748);
not NOT1 (N13750, N13732);
nand NAND3 (N13751, N13738, N1934, N5603);
buf BUF1 (N13752, N13740);
nand NAND2 (N13753, N13743, N978);
not NOT1 (N13754, N13749);
and AND4 (N13755, N13751, N9387, N3652, N10602);
xor XOR2 (N13756, N13752, N5494);
xor XOR2 (N13757, N13753, N3509);
not NOT1 (N13758, N13734);
nor NOR2 (N13759, N13756, N1053);
xor XOR2 (N13760, N13744, N1507);
nor NOR4 (N13761, N13750, N10599, N2365, N964);
and AND4 (N13762, N13761, N5280, N13436, N1422);
nor NOR4 (N13763, N13758, N8603, N3465, N11033);
buf BUF1 (N13764, N13762);
and AND3 (N13765, N13755, N2088, N11459);
nor NOR2 (N13766, N13765, N11485);
buf BUF1 (N13767, N13745);
buf BUF1 (N13768, N13760);
not NOT1 (N13769, N13766);
xor XOR2 (N13770, N13757, N9747);
nor NOR4 (N13771, N13754, N10545, N9192, N4246);
nand NAND3 (N13772, N13747, N5347, N9025);
xor XOR2 (N13773, N13763, N4745);
and AND2 (N13774, N13741, N1333);
nand NAND2 (N13775, N13764, N6602);
and AND3 (N13776, N13774, N3592, N11178);
or OR2 (N13777, N13770, N11082);
not NOT1 (N13778, N13771);
xor XOR2 (N13779, N13768, N5631);
nand NAND4 (N13780, N13775, N443, N10658, N8617);
nor NOR4 (N13781, N13777, N3793, N11723, N4807);
or OR3 (N13782, N13779, N7943, N6553);
buf BUF1 (N13783, N13769);
or OR2 (N13784, N13776, N13217);
or OR3 (N13785, N13782, N6095, N10412);
nor NOR2 (N13786, N13780, N1036);
nand NAND2 (N13787, N13786, N7008);
or OR4 (N13788, N13784, N4021, N10310, N12175);
nor NOR3 (N13789, N13759, N8478, N5056);
and AND4 (N13790, N13787, N10650, N9551, N5696);
or OR3 (N13791, N13772, N10697, N1768);
nor NOR2 (N13792, N13773, N6866);
nor NOR4 (N13793, N13781, N11823, N10135, N7293);
not NOT1 (N13794, N13791);
buf BUF1 (N13795, N13778);
buf BUF1 (N13796, N13795);
nor NOR4 (N13797, N13790, N1732, N4105, N11205);
nor NOR3 (N13798, N13794, N1796, N2391);
xor XOR2 (N13799, N13789, N12318);
buf BUF1 (N13800, N13785);
xor XOR2 (N13801, N13798, N13560);
or OR2 (N13802, N13801, N610);
and AND3 (N13803, N13793, N12117, N5314);
xor XOR2 (N13804, N13797, N12115);
and AND3 (N13805, N13792, N8302, N8811);
and AND2 (N13806, N13783, N5431);
or OR4 (N13807, N13800, N11208, N9110, N156);
not NOT1 (N13808, N13804);
xor XOR2 (N13809, N13788, N6937);
or OR2 (N13810, N13805, N7962);
and AND2 (N13811, N13767, N13242);
or OR3 (N13812, N13803, N4415, N4332);
buf BUF1 (N13813, N13796);
nor NOR2 (N13814, N13799, N204);
nand NAND3 (N13815, N13802, N11392, N8260);
or OR4 (N13816, N13808, N5092, N3954, N3843);
buf BUF1 (N13817, N13813);
nor NOR2 (N13818, N13816, N8452);
nand NAND2 (N13819, N13807, N12174);
xor XOR2 (N13820, N13819, N7887);
and AND4 (N13821, N13810, N13769, N11307, N12904);
buf BUF1 (N13822, N13821);
nor NOR3 (N13823, N13818, N11046, N11957);
nand NAND2 (N13824, N13806, N13304);
or OR4 (N13825, N13824, N2360, N12123, N11468);
not NOT1 (N13826, N13825);
xor XOR2 (N13827, N13812, N6590);
nand NAND4 (N13828, N13817, N12544, N1558, N11814);
buf BUF1 (N13829, N13815);
nor NOR3 (N13830, N13823, N12848, N3507);
nand NAND4 (N13831, N13811, N11449, N928, N12155);
buf BUF1 (N13832, N13827);
buf BUF1 (N13833, N13822);
xor XOR2 (N13834, N13833, N11334);
nand NAND4 (N13835, N13826, N7120, N9547, N4243);
nand NAND3 (N13836, N13834, N12456, N13643);
xor XOR2 (N13837, N13820, N6123);
buf BUF1 (N13838, N13836);
xor XOR2 (N13839, N13809, N8852);
nand NAND3 (N13840, N13832, N12790, N11147);
buf BUF1 (N13841, N13837);
nand NAND4 (N13842, N13840, N3343, N7307, N590);
xor XOR2 (N13843, N13831, N1950);
nor NOR2 (N13844, N13830, N3793);
xor XOR2 (N13845, N13844, N8811);
xor XOR2 (N13846, N13839, N6853);
and AND4 (N13847, N13814, N894, N2968, N3973);
buf BUF1 (N13848, N13828);
nor NOR4 (N13849, N13847, N9049, N6967, N6354);
not NOT1 (N13850, N13835);
not NOT1 (N13851, N13850);
nor NOR4 (N13852, N13843, N11531, N3399, N7229);
nor NOR4 (N13853, N13852, N995, N10529, N730);
not NOT1 (N13854, N13846);
and AND2 (N13855, N13849, N11031);
not NOT1 (N13856, N13854);
nor NOR4 (N13857, N13841, N11134, N12107, N3315);
and AND2 (N13858, N13853, N9458);
or OR4 (N13859, N13848, N9354, N6024, N12202);
nor NOR4 (N13860, N13829, N8450, N4267, N11788);
xor XOR2 (N13861, N13860, N7273);
nand NAND4 (N13862, N13858, N11844, N10725, N9213);
buf BUF1 (N13863, N13855);
or OR3 (N13864, N13861, N12541, N10286);
nand NAND3 (N13865, N13863, N8794, N4624);
and AND4 (N13866, N13845, N3774, N1869, N6494);
buf BUF1 (N13867, N13865);
or OR3 (N13868, N13851, N7135, N3827);
nand NAND2 (N13869, N13864, N10047);
buf BUF1 (N13870, N13857);
nor NOR3 (N13871, N13859, N10355, N9070);
and AND4 (N13872, N13868, N11557, N10412, N8794);
buf BUF1 (N13873, N13862);
xor XOR2 (N13874, N13856, N4011);
nand NAND2 (N13875, N13869, N797);
buf BUF1 (N13876, N13871);
nand NAND4 (N13877, N13875, N2326, N2510, N10556);
nand NAND3 (N13878, N13838, N220, N4959);
nand NAND2 (N13879, N13870, N1249);
nor NOR3 (N13880, N13866, N3359, N13532);
not NOT1 (N13881, N13867);
or OR4 (N13882, N13880, N3246, N2543, N293);
xor XOR2 (N13883, N13842, N7622);
nand NAND3 (N13884, N13874, N8528, N463);
buf BUF1 (N13885, N13872);
not NOT1 (N13886, N13885);
buf BUF1 (N13887, N13884);
buf BUF1 (N13888, N13877);
nand NAND2 (N13889, N13876, N10498);
and AND2 (N13890, N13883, N3845);
buf BUF1 (N13891, N13882);
buf BUF1 (N13892, N13873);
buf BUF1 (N13893, N13879);
not NOT1 (N13894, N13886);
buf BUF1 (N13895, N13881);
not NOT1 (N13896, N13890);
and AND4 (N13897, N13878, N8851, N12138, N12221);
buf BUF1 (N13898, N13888);
nand NAND4 (N13899, N13892, N9260, N12937, N552);
not NOT1 (N13900, N13897);
xor XOR2 (N13901, N13898, N10531);
nand NAND4 (N13902, N13896, N6245, N8576, N2434);
xor XOR2 (N13903, N13887, N6066);
buf BUF1 (N13904, N13902);
nand NAND4 (N13905, N13893, N4846, N6391, N7832);
or OR3 (N13906, N13899, N7803, N11370);
and AND3 (N13907, N13901, N8165, N12720);
not NOT1 (N13908, N13891);
nor NOR4 (N13909, N13894, N11594, N4853, N11491);
xor XOR2 (N13910, N13906, N6433);
xor XOR2 (N13911, N13900, N2679);
or OR3 (N13912, N13895, N4702, N651);
or OR3 (N13913, N13911, N12985, N12787);
nand NAND2 (N13914, N13889, N12139);
nor NOR2 (N13915, N13907, N9224);
not NOT1 (N13916, N13913);
not NOT1 (N13917, N13916);
nor NOR2 (N13918, N13915, N7675);
not NOT1 (N13919, N13908);
xor XOR2 (N13920, N13918, N8968);
nand NAND2 (N13921, N13904, N5426);
nor NOR4 (N13922, N13903, N3047, N13474, N9523);
or OR4 (N13923, N13921, N2503, N12702, N6019);
not NOT1 (N13924, N13909);
buf BUF1 (N13925, N13924);
xor XOR2 (N13926, N13922, N4362);
nand NAND4 (N13927, N13920, N517, N8829, N8842);
nand NAND2 (N13928, N13910, N488);
not NOT1 (N13929, N13914);
nand NAND2 (N13930, N13926, N783);
or OR4 (N13931, N13919, N9788, N2998, N4903);
xor XOR2 (N13932, N13929, N10711);
nor NOR4 (N13933, N13912, N2484, N7132, N12342);
nor NOR3 (N13934, N13931, N4708, N11518);
and AND3 (N13935, N13917, N4603, N12220);
xor XOR2 (N13936, N13925, N12513);
buf BUF1 (N13937, N13927);
xor XOR2 (N13938, N13934, N1363);
xor XOR2 (N13939, N13928, N122);
xor XOR2 (N13940, N13932, N3575);
or OR4 (N13941, N13938, N1089, N13247, N11178);
or OR3 (N13942, N13940, N1240, N10096);
not NOT1 (N13943, N13935);
nand NAND2 (N13944, N13941, N6555);
not NOT1 (N13945, N13930);
buf BUF1 (N13946, N13942);
or OR3 (N13947, N13944, N7240, N1191);
not NOT1 (N13948, N13939);
or OR2 (N13949, N13946, N3814);
nor NOR2 (N13950, N13945, N1255);
not NOT1 (N13951, N13923);
nor NOR4 (N13952, N13951, N218, N8795, N13577);
not NOT1 (N13953, N13947);
and AND4 (N13954, N13937, N7507, N11788, N3034);
nand NAND4 (N13955, N13936, N5407, N7976, N6106);
and AND4 (N13956, N13905, N11830, N10872, N13272);
nor NOR2 (N13957, N13950, N10381);
not NOT1 (N13958, N13949);
and AND4 (N13959, N13943, N2401, N12379, N157);
xor XOR2 (N13960, N13957, N4438);
and AND4 (N13961, N13933, N131, N8857, N9900);
buf BUF1 (N13962, N13961);
and AND2 (N13963, N13955, N2571);
nor NOR2 (N13964, N13960, N3338);
xor XOR2 (N13965, N13948, N909);
nor NOR2 (N13966, N13958, N1199);
xor XOR2 (N13967, N13953, N3004);
xor XOR2 (N13968, N13963, N5210);
or OR2 (N13969, N13962, N973);
buf BUF1 (N13970, N13968);
not NOT1 (N13971, N13952);
or OR4 (N13972, N13967, N13710, N6864, N1868);
nand NAND3 (N13973, N13972, N4813, N3618);
xor XOR2 (N13974, N13954, N1975);
buf BUF1 (N13975, N13974);
buf BUF1 (N13976, N13966);
not NOT1 (N13977, N13959);
not NOT1 (N13978, N13956);
and AND4 (N13979, N13976, N4189, N12929, N5374);
buf BUF1 (N13980, N13975);
nand NAND4 (N13981, N13965, N9986, N7437, N8911);
and AND2 (N13982, N13977, N5315);
not NOT1 (N13983, N13971);
nor NOR2 (N13984, N13981, N3569);
buf BUF1 (N13985, N13970);
not NOT1 (N13986, N13982);
buf BUF1 (N13987, N13984);
not NOT1 (N13988, N13980);
buf BUF1 (N13989, N13985);
nor NOR2 (N13990, N13973, N11154);
nor NOR4 (N13991, N13990, N3128, N12791, N8258);
and AND4 (N13992, N13991, N10015, N355, N12098);
and AND2 (N13993, N13989, N12425);
or OR4 (N13994, N13987, N10458, N11574, N7959);
or OR2 (N13995, N13988, N984);
nor NOR4 (N13996, N13969, N3773, N3162, N675);
or OR3 (N13997, N13995, N4507, N3875);
xor XOR2 (N13998, N13986, N11563);
xor XOR2 (N13999, N13979, N12584);
nand NAND3 (N14000, N13999, N6122, N13707);
nand NAND4 (N14001, N13964, N9268, N4033, N3416);
nand NAND4 (N14002, N13994, N7758, N1174, N1572);
not NOT1 (N14003, N13993);
and AND4 (N14004, N14001, N1951, N3179, N2535);
xor XOR2 (N14005, N13996, N898);
or OR3 (N14006, N14004, N1326, N2860);
nor NOR4 (N14007, N13978, N10454, N11825, N2338);
xor XOR2 (N14008, N13992, N11163);
nand NAND4 (N14009, N14000, N7425, N2401, N10225);
not NOT1 (N14010, N13998);
buf BUF1 (N14011, N14010);
nand NAND2 (N14012, N13983, N422);
xor XOR2 (N14013, N13997, N3825);
or OR3 (N14014, N14003, N12636, N7714);
or OR3 (N14015, N14009, N4164, N12318);
xor XOR2 (N14016, N14015, N10307);
nor NOR3 (N14017, N14014, N11761, N11445);
xor XOR2 (N14018, N14002, N1689);
nand NAND3 (N14019, N14012, N130, N8452);
buf BUF1 (N14020, N14017);
and AND4 (N14021, N14011, N12271, N12111, N13524);
nor NOR3 (N14022, N14018, N13228, N13315);
and AND2 (N14023, N14007, N5318);
and AND3 (N14024, N14020, N6700, N5043);
buf BUF1 (N14025, N14013);
or OR4 (N14026, N14016, N1265, N3006, N6023);
xor XOR2 (N14027, N14024, N2917);
nand NAND4 (N14028, N14022, N10493, N13199, N12030);
nand NAND3 (N14029, N14021, N4735, N11730);
buf BUF1 (N14030, N14006);
nor NOR2 (N14031, N14025, N93);
nand NAND2 (N14032, N14027, N4047);
nor NOR4 (N14033, N14030, N174, N7052, N10345);
and AND4 (N14034, N14032, N1504, N3472, N11468);
not NOT1 (N14035, N14028);
buf BUF1 (N14036, N14029);
nor NOR3 (N14037, N14005, N13274, N9098);
nand NAND2 (N14038, N14026, N3378);
and AND2 (N14039, N14037, N6058);
xor XOR2 (N14040, N14034, N8733);
xor XOR2 (N14041, N14038, N7150);
xor XOR2 (N14042, N14039, N7606);
xor XOR2 (N14043, N14040, N1071);
and AND2 (N14044, N14043, N10234);
or OR4 (N14045, N14008, N8756, N11478, N12391);
not NOT1 (N14046, N14035);
nand NAND3 (N14047, N14044, N7604, N3842);
nor NOR3 (N14048, N14041, N9239, N9688);
not NOT1 (N14049, N14042);
not NOT1 (N14050, N14036);
and AND2 (N14051, N14046, N8701);
not NOT1 (N14052, N14045);
buf BUF1 (N14053, N14049);
buf BUF1 (N14054, N14031);
not NOT1 (N14055, N14023);
or OR2 (N14056, N14048, N11947);
buf BUF1 (N14057, N14056);
nor NOR4 (N14058, N14019, N11696, N8370, N13861);
xor XOR2 (N14059, N14057, N7248);
nor NOR3 (N14060, N14059, N3892, N8577);
and AND4 (N14061, N14051, N998, N11902, N12915);
or OR4 (N14062, N14055, N3772, N11621, N3603);
and AND3 (N14063, N14052, N3750, N5560);
xor XOR2 (N14064, N14053, N1723);
xor XOR2 (N14065, N14058, N4275);
buf BUF1 (N14066, N14060);
not NOT1 (N14067, N14054);
xor XOR2 (N14068, N14066, N8643);
nor NOR2 (N14069, N14050, N10132);
buf BUF1 (N14070, N14068);
nand NAND3 (N14071, N14070, N9889, N13650);
and AND4 (N14072, N14063, N4633, N2807, N4571);
not NOT1 (N14073, N14047);
or OR2 (N14074, N14071, N5113);
nor NOR4 (N14075, N14062, N12875, N510, N1137);
xor XOR2 (N14076, N14067, N2513);
buf BUF1 (N14077, N14033);
xor XOR2 (N14078, N14064, N1823);
xor XOR2 (N14079, N14074, N12200);
or OR4 (N14080, N14072, N2092, N8927, N10043);
nand NAND3 (N14081, N14077, N12098, N11500);
nand NAND3 (N14082, N14065, N4759, N9714);
or OR2 (N14083, N14080, N11976);
not NOT1 (N14084, N14069);
buf BUF1 (N14085, N14073);
not NOT1 (N14086, N14082);
and AND3 (N14087, N14079, N2514, N2725);
or OR3 (N14088, N14085, N8151, N5507);
nand NAND2 (N14089, N14078, N2403);
nand NAND2 (N14090, N14084, N7645);
and AND4 (N14091, N14090, N13341, N4158, N1102);
xor XOR2 (N14092, N14088, N4133);
buf BUF1 (N14093, N14087);
buf BUF1 (N14094, N14089);
buf BUF1 (N14095, N14086);
nor NOR2 (N14096, N14092, N6730);
xor XOR2 (N14097, N14091, N7522);
not NOT1 (N14098, N14096);
nor NOR3 (N14099, N14097, N5919, N7857);
nor NOR4 (N14100, N14075, N6407, N4355, N11462);
nand NAND4 (N14101, N14061, N13602, N1409, N3892);
not NOT1 (N14102, N14095);
and AND2 (N14103, N14094, N7794);
buf BUF1 (N14104, N14076);
and AND4 (N14105, N14099, N12442, N10846, N7247);
buf BUF1 (N14106, N14102);
not NOT1 (N14107, N14100);
xor XOR2 (N14108, N14104, N9251);
xor XOR2 (N14109, N14106, N4937);
or OR2 (N14110, N14083, N540);
or OR4 (N14111, N14105, N11031, N9435, N2064);
nand NAND2 (N14112, N14107, N5369);
xor XOR2 (N14113, N14112, N7085);
xor XOR2 (N14114, N14093, N4177);
buf BUF1 (N14115, N14111);
xor XOR2 (N14116, N14108, N6681);
nand NAND3 (N14117, N14101, N10101, N3884);
nor NOR3 (N14118, N14109, N11844, N144);
not NOT1 (N14119, N14116);
not NOT1 (N14120, N14098);
or OR3 (N14121, N14115, N12734, N8952);
nor NOR4 (N14122, N14110, N10422, N12998, N3886);
or OR3 (N14123, N14081, N7405, N1910);
or OR2 (N14124, N14114, N11591);
xor XOR2 (N14125, N14122, N3173);
and AND3 (N14126, N14121, N4069, N952);
xor XOR2 (N14127, N14119, N2260);
not NOT1 (N14128, N14120);
buf BUF1 (N14129, N14128);
nor NOR2 (N14130, N14118, N10004);
nor NOR4 (N14131, N14129, N13495, N467, N455);
not NOT1 (N14132, N14130);
and AND3 (N14133, N14113, N5751, N6526);
buf BUF1 (N14134, N14124);
xor XOR2 (N14135, N14103, N8891);
xor XOR2 (N14136, N14117, N122);
and AND3 (N14137, N14131, N12479, N12195);
buf BUF1 (N14138, N14134);
xor XOR2 (N14139, N14135, N4212);
nand NAND2 (N14140, N14123, N2195);
buf BUF1 (N14141, N14125);
xor XOR2 (N14142, N14138, N6610);
buf BUF1 (N14143, N14127);
and AND4 (N14144, N14126, N3982, N1905, N7123);
buf BUF1 (N14145, N14133);
or OR4 (N14146, N14139, N6896, N10634, N9617);
not NOT1 (N14147, N14145);
nand NAND2 (N14148, N14132, N7717);
nor NOR3 (N14149, N14146, N943, N11060);
xor XOR2 (N14150, N14136, N7820);
and AND2 (N14151, N14141, N3913);
xor XOR2 (N14152, N14143, N55);
xor XOR2 (N14153, N14142, N3547);
nand NAND4 (N14154, N14137, N6246, N6643, N166);
nor NOR4 (N14155, N14152, N421, N8076, N6682);
nand NAND2 (N14156, N14150, N9008);
nor NOR2 (N14157, N14154, N2404);
nor NOR3 (N14158, N14155, N691, N389);
xor XOR2 (N14159, N14158, N5593);
not NOT1 (N14160, N14159);
xor XOR2 (N14161, N14147, N12261);
nand NAND4 (N14162, N14151, N5687, N12452, N5844);
nand NAND4 (N14163, N14144, N7432, N6924, N3624);
xor XOR2 (N14164, N14149, N10092);
or OR2 (N14165, N14148, N4819);
buf BUF1 (N14166, N14140);
and AND4 (N14167, N14153, N11733, N2812, N10118);
or OR2 (N14168, N14156, N10749);
or OR4 (N14169, N14167, N908, N8145, N5806);
nand NAND4 (N14170, N14157, N3327, N7484, N7402);
nand NAND2 (N14171, N14166, N4173);
not NOT1 (N14172, N14162);
buf BUF1 (N14173, N14171);
not NOT1 (N14174, N14169);
xor XOR2 (N14175, N14174, N5911);
xor XOR2 (N14176, N14161, N12464);
or OR4 (N14177, N14170, N6773, N6856, N11384);
or OR2 (N14178, N14177, N4157);
nand NAND3 (N14179, N14178, N12957, N4911);
nor NOR2 (N14180, N14179, N1717);
buf BUF1 (N14181, N14173);
or OR2 (N14182, N14181, N8611);
or OR4 (N14183, N14172, N2067, N13186, N8886);
nand NAND2 (N14184, N14176, N13593);
not NOT1 (N14185, N14180);
and AND4 (N14186, N14183, N13239, N11370, N7530);
not NOT1 (N14187, N14184);
nand NAND2 (N14188, N14182, N7476);
xor XOR2 (N14189, N14185, N2364);
or OR2 (N14190, N14186, N5531);
buf BUF1 (N14191, N14168);
not NOT1 (N14192, N14164);
xor XOR2 (N14193, N14190, N3692);
buf BUF1 (N14194, N14189);
and AND4 (N14195, N14194, N9162, N8902, N6405);
nor NOR3 (N14196, N14195, N6577, N11972);
not NOT1 (N14197, N14196);
not NOT1 (N14198, N14192);
nand NAND4 (N14199, N14160, N13814, N8702, N5584);
and AND4 (N14200, N14191, N3657, N3710, N6731);
xor XOR2 (N14201, N14175, N12819);
buf BUF1 (N14202, N14198);
buf BUF1 (N14203, N14193);
nor NOR2 (N14204, N14199, N1649);
not NOT1 (N14205, N14197);
nand NAND4 (N14206, N14203, N3892, N476, N7371);
or OR2 (N14207, N14206, N9328);
nor NOR4 (N14208, N14163, N12572, N5763, N13999);
nor NOR4 (N14209, N14204, N12848, N13757, N2525);
and AND3 (N14210, N14209, N5724, N13617);
and AND3 (N14211, N14202, N2741, N7665);
and AND3 (N14212, N14200, N14077, N7659);
and AND4 (N14213, N14201, N977, N2173, N4666);
buf BUF1 (N14214, N14210);
xor XOR2 (N14215, N14213, N6902);
and AND4 (N14216, N14215, N4014, N9829, N10194);
and AND2 (N14217, N14214, N7590);
and AND2 (N14218, N14187, N13101);
not NOT1 (N14219, N14207);
or OR4 (N14220, N14216, N9652, N535, N8751);
or OR2 (N14221, N14219, N6050);
xor XOR2 (N14222, N14218, N3562);
nor NOR4 (N14223, N14208, N13641, N411, N13405);
and AND4 (N14224, N14165, N11969, N2529, N1320);
and AND2 (N14225, N14217, N6365);
buf BUF1 (N14226, N14212);
nor NOR3 (N14227, N14224, N78, N4740);
nor NOR3 (N14228, N14220, N5075, N5210);
nor NOR4 (N14229, N14223, N12696, N13868, N6738);
and AND3 (N14230, N14222, N275, N1232);
nand NAND4 (N14231, N14225, N6718, N168, N11423);
buf BUF1 (N14232, N14226);
buf BUF1 (N14233, N14211);
and AND4 (N14234, N14221, N2747, N1487, N12110);
not NOT1 (N14235, N14231);
nand NAND4 (N14236, N14235, N4807, N13333, N9367);
buf BUF1 (N14237, N14188);
or OR2 (N14238, N14236, N10465);
or OR4 (N14239, N14232, N9894, N11206, N1576);
xor XOR2 (N14240, N14228, N3233);
or OR3 (N14241, N14239, N9383, N8811);
buf BUF1 (N14242, N14227);
not NOT1 (N14243, N14242);
nor NOR2 (N14244, N14230, N6474);
xor XOR2 (N14245, N14243, N4705);
or OR2 (N14246, N14233, N9344);
not NOT1 (N14247, N14245);
and AND2 (N14248, N14205, N11610);
nor NOR4 (N14249, N14234, N3414, N8751, N2525);
not NOT1 (N14250, N14247);
and AND2 (N14251, N14237, N13493);
buf BUF1 (N14252, N14244);
nand NAND2 (N14253, N14246, N2650);
not NOT1 (N14254, N14251);
nand NAND2 (N14255, N14238, N1015);
xor XOR2 (N14256, N14240, N9730);
and AND4 (N14257, N14249, N12271, N1689, N7887);
nor NOR4 (N14258, N14257, N3913, N11826, N4665);
nor NOR4 (N14259, N14250, N3635, N12292, N5858);
nor NOR3 (N14260, N14259, N634, N1981);
buf BUF1 (N14261, N14255);
not NOT1 (N14262, N14260);
or OR2 (N14263, N14248, N1914);
and AND2 (N14264, N14256, N11995);
buf BUF1 (N14265, N14252);
and AND4 (N14266, N14253, N12615, N13345, N9357);
nor NOR4 (N14267, N14229, N4613, N14110, N4710);
and AND3 (N14268, N14261, N2498, N6865);
not NOT1 (N14269, N14263);
nor NOR4 (N14270, N14265, N8271, N2022, N3480);
buf BUF1 (N14271, N14268);
not NOT1 (N14272, N14241);
xor XOR2 (N14273, N14264, N11485);
or OR3 (N14274, N14272, N11539, N12149);
and AND2 (N14275, N14262, N7928);
not NOT1 (N14276, N14275);
and AND2 (N14277, N14269, N13109);
and AND3 (N14278, N14273, N2165, N11943);
or OR4 (N14279, N14254, N10993, N10900, N9759);
xor XOR2 (N14280, N14277, N13871);
not NOT1 (N14281, N14274);
or OR3 (N14282, N14278, N8607, N10297);
or OR4 (N14283, N14266, N6595, N10194, N7504);
xor XOR2 (N14284, N14280, N9675);
not NOT1 (N14285, N14271);
nand NAND3 (N14286, N14279, N6163, N13130);
and AND3 (N14287, N14276, N7101, N12923);
nor NOR4 (N14288, N14282, N12308, N49, N9818);
buf BUF1 (N14289, N14283);
xor XOR2 (N14290, N14289, N6119);
nor NOR2 (N14291, N14286, N3069);
buf BUF1 (N14292, N14285);
nand NAND4 (N14293, N14291, N6752, N841, N11141);
nor NOR4 (N14294, N14281, N12408, N1291, N11435);
buf BUF1 (N14295, N14270);
and AND4 (N14296, N14292, N4059, N8082, N135);
or OR3 (N14297, N14267, N11526, N265);
and AND2 (N14298, N14297, N2210);
xor XOR2 (N14299, N14295, N9259);
not NOT1 (N14300, N14298);
nand NAND2 (N14301, N14290, N7511);
and AND4 (N14302, N14300, N9068, N6701, N11901);
buf BUF1 (N14303, N14293);
buf BUF1 (N14304, N14299);
xor XOR2 (N14305, N14303, N4878);
and AND2 (N14306, N14296, N9034);
and AND2 (N14307, N14302, N2786);
nand NAND2 (N14308, N14301, N1380);
and AND4 (N14309, N14258, N674, N8763, N7345);
nand NAND2 (N14310, N14287, N13254);
or OR2 (N14311, N14288, N12728);
buf BUF1 (N14312, N14305);
xor XOR2 (N14313, N14308, N490);
xor XOR2 (N14314, N14304, N7190);
buf BUF1 (N14315, N14294);
not NOT1 (N14316, N14307);
nand NAND4 (N14317, N14310, N11126, N2972, N6681);
nor NOR2 (N14318, N14317, N5516);
buf BUF1 (N14319, N14318);
and AND4 (N14320, N14316, N211, N11231, N7080);
nor NOR2 (N14321, N14320, N188);
buf BUF1 (N14322, N14284);
buf BUF1 (N14323, N14313);
nor NOR4 (N14324, N14322, N14174, N2993, N5744);
nand NAND4 (N14325, N14324, N6744, N11245, N11683);
and AND2 (N14326, N14309, N2762);
or OR4 (N14327, N14325, N4661, N7399, N8542);
xor XOR2 (N14328, N14319, N5274);
or OR2 (N14329, N14306, N4016);
and AND3 (N14330, N14315, N2725, N9778);
not NOT1 (N14331, N14330);
not NOT1 (N14332, N14311);
nor NOR2 (N14333, N14327, N9787);
xor XOR2 (N14334, N14332, N11696);
or OR4 (N14335, N14329, N8802, N2690, N8191);
xor XOR2 (N14336, N14314, N6905);
nor NOR4 (N14337, N14328, N6419, N4448, N362);
not NOT1 (N14338, N14333);
buf BUF1 (N14339, N14337);
xor XOR2 (N14340, N14321, N10795);
and AND3 (N14341, N14336, N3936, N9211);
buf BUF1 (N14342, N14340);
buf BUF1 (N14343, N14326);
or OR4 (N14344, N14341, N372, N2067, N3152);
not NOT1 (N14345, N14323);
and AND4 (N14346, N14335, N6158, N5022, N902);
buf BUF1 (N14347, N14346);
xor XOR2 (N14348, N14342, N8602);
or OR2 (N14349, N14331, N12442);
xor XOR2 (N14350, N14349, N9780);
xor XOR2 (N14351, N14312, N9914);
nand NAND3 (N14352, N14347, N12467, N8899);
nand NAND2 (N14353, N14352, N5589);
xor XOR2 (N14354, N14348, N13763);
buf BUF1 (N14355, N14344);
nand NAND3 (N14356, N14353, N8810, N10008);
xor XOR2 (N14357, N14351, N3185);
xor XOR2 (N14358, N14354, N9362);
not NOT1 (N14359, N14343);
buf BUF1 (N14360, N14339);
xor XOR2 (N14361, N14358, N9826);
buf BUF1 (N14362, N14356);
nand NAND4 (N14363, N14355, N11135, N12524, N13760);
nand NAND2 (N14364, N14334, N6542);
nor NOR3 (N14365, N14357, N5038, N6663);
and AND4 (N14366, N14365, N1969, N10556, N14179);
nor NOR4 (N14367, N14350, N11882, N9014, N12186);
nor NOR2 (N14368, N14338, N1180);
buf BUF1 (N14369, N14368);
or OR4 (N14370, N14360, N8107, N9078, N12650);
nor NOR4 (N14371, N14363, N7145, N2820, N8547);
not NOT1 (N14372, N14359);
and AND4 (N14373, N14345, N2618, N6100, N12667);
not NOT1 (N14374, N14371);
nand NAND3 (N14375, N14367, N13192, N14253);
or OR3 (N14376, N14372, N2798, N4017);
and AND2 (N14377, N14366, N5304);
or OR3 (N14378, N14373, N1135, N3792);
not NOT1 (N14379, N14374);
or OR3 (N14380, N14375, N10841, N8292);
xor XOR2 (N14381, N14370, N9362);
nor NOR2 (N14382, N14381, N6358);
nand NAND3 (N14383, N14376, N12869, N405);
or OR2 (N14384, N14364, N2332);
and AND4 (N14385, N14369, N11345, N424, N2003);
nand NAND2 (N14386, N14361, N6388);
nand NAND3 (N14387, N14382, N4459, N6990);
nand NAND3 (N14388, N14379, N13082, N5205);
nor NOR4 (N14389, N14362, N7166, N10292, N8510);
nand NAND4 (N14390, N14386, N1873, N14156, N4086);
nor NOR4 (N14391, N14388, N9693, N5536, N12571);
not NOT1 (N14392, N14377);
nand NAND2 (N14393, N14384, N2353);
nand NAND2 (N14394, N14387, N6384);
buf BUF1 (N14395, N14392);
and AND3 (N14396, N14390, N12708, N4371);
xor XOR2 (N14397, N14395, N1993);
nand NAND3 (N14398, N14397, N6495, N2507);
nor NOR2 (N14399, N14391, N3921);
or OR3 (N14400, N14385, N5229, N10499);
and AND3 (N14401, N14389, N2686, N10130);
and AND3 (N14402, N14401, N6934, N11106);
nand NAND2 (N14403, N14393, N2541);
or OR3 (N14404, N14396, N13726, N4148);
nand NAND3 (N14405, N14403, N9183, N10957);
or OR2 (N14406, N14383, N13235);
and AND2 (N14407, N14378, N3244);
buf BUF1 (N14408, N14400);
nand NAND4 (N14409, N14399, N9590, N8535, N11028);
or OR4 (N14410, N14394, N4560, N12007, N11716);
nor NOR4 (N14411, N14402, N1222, N3122, N13332);
and AND4 (N14412, N14405, N5902, N8689, N6498);
nand NAND3 (N14413, N14412, N2363, N11400);
not NOT1 (N14414, N14406);
or OR3 (N14415, N14411, N7784, N218);
nand NAND2 (N14416, N14408, N3244);
xor XOR2 (N14417, N14416, N4209);
nand NAND4 (N14418, N14398, N3986, N11598, N341);
xor XOR2 (N14419, N14415, N7306);
or OR4 (N14420, N14410, N10346, N14306, N7516);
buf BUF1 (N14421, N14409);
xor XOR2 (N14422, N14420, N5838);
and AND3 (N14423, N14417, N14421, N1541);
xor XOR2 (N14424, N4861, N5758);
nand NAND4 (N14425, N14422, N1842, N10830, N1205);
nor NOR4 (N14426, N14404, N1135, N8539, N4287);
nor NOR2 (N14427, N14419, N13461);
nand NAND2 (N14428, N14426, N3669);
or OR4 (N14429, N14413, N5310, N356, N916);
or OR2 (N14430, N14425, N8375);
buf BUF1 (N14431, N14407);
or OR2 (N14432, N14431, N976);
and AND4 (N14433, N14427, N8110, N2657, N6673);
nand NAND3 (N14434, N14433, N492, N13812);
xor XOR2 (N14435, N14432, N3841);
xor XOR2 (N14436, N14435, N8073);
or OR2 (N14437, N14414, N3298);
nor NOR3 (N14438, N14380, N3937, N10695);
nor NOR3 (N14439, N14424, N9125, N5195);
and AND3 (N14440, N14429, N10606, N10687);
nand NAND2 (N14441, N14438, N11492);
not NOT1 (N14442, N14437);
not NOT1 (N14443, N14440);
xor XOR2 (N14444, N14441, N662);
nor NOR4 (N14445, N14430, N8317, N10373, N12819);
or OR4 (N14446, N14434, N2199, N12942, N3724);
and AND3 (N14447, N14418, N13457, N10894);
or OR2 (N14448, N14428, N8260);
not NOT1 (N14449, N14448);
not NOT1 (N14450, N14436);
or OR3 (N14451, N14439, N4195, N1370);
or OR4 (N14452, N14445, N840, N8000, N9663);
buf BUF1 (N14453, N14451);
not NOT1 (N14454, N14423);
xor XOR2 (N14455, N14452, N13009);
buf BUF1 (N14456, N14446);
xor XOR2 (N14457, N14453, N7975);
and AND2 (N14458, N14443, N10913);
buf BUF1 (N14459, N14450);
buf BUF1 (N14460, N14454);
xor XOR2 (N14461, N14457, N6775);
nand NAND4 (N14462, N14455, N14241, N12491, N1400);
nand NAND2 (N14463, N14460, N4226);
nor NOR4 (N14464, N14442, N5100, N13030, N1564);
or OR2 (N14465, N14456, N4874);
nor NOR3 (N14466, N14463, N2594, N10473);
or OR3 (N14467, N14459, N1485, N7140);
and AND4 (N14468, N14458, N8311, N1455, N649);
not NOT1 (N14469, N14444);
and AND2 (N14470, N14447, N1641);
nor NOR2 (N14471, N14464, N2143);
xor XOR2 (N14472, N14467, N1288);
and AND4 (N14473, N14468, N11623, N2059, N13964);
and AND2 (N14474, N14466, N477);
buf BUF1 (N14475, N14471);
buf BUF1 (N14476, N14462);
xor XOR2 (N14477, N14470, N9119);
buf BUF1 (N14478, N14475);
not NOT1 (N14479, N14477);
not NOT1 (N14480, N14472);
or OR4 (N14481, N14449, N8963, N2006, N11625);
or OR4 (N14482, N14461, N5943, N4485, N7837);
xor XOR2 (N14483, N14479, N5389);
nand NAND3 (N14484, N14476, N2772, N10948);
xor XOR2 (N14485, N14480, N5043);
nor NOR3 (N14486, N14484, N9839, N773);
buf BUF1 (N14487, N14465);
nor NOR2 (N14488, N14474, N1681);
nand NAND2 (N14489, N14482, N9276);
xor XOR2 (N14490, N14488, N5524);
xor XOR2 (N14491, N14473, N9746);
and AND3 (N14492, N14481, N8366, N11633);
or OR3 (N14493, N14485, N1902, N9960);
not NOT1 (N14494, N14491);
nor NOR2 (N14495, N14493, N7270);
buf BUF1 (N14496, N14487);
nand NAND3 (N14497, N14495, N5963, N11746);
or OR3 (N14498, N14486, N10021, N14481);
or OR4 (N14499, N14489, N4499, N12843, N3380);
and AND4 (N14500, N14494, N5686, N1626, N11008);
nand NAND3 (N14501, N14478, N12190, N7413);
nor NOR2 (N14502, N14500, N12777);
buf BUF1 (N14503, N14501);
or OR4 (N14504, N14503, N5764, N4871, N13451);
or OR2 (N14505, N14499, N2615);
nand NAND3 (N14506, N14469, N4881, N11571);
nor NOR3 (N14507, N14504, N11515, N257);
buf BUF1 (N14508, N14497);
and AND4 (N14509, N14496, N8438, N3003, N3525);
xor XOR2 (N14510, N14508, N7659);
xor XOR2 (N14511, N14490, N6450);
nand NAND3 (N14512, N14492, N4373, N5647);
xor XOR2 (N14513, N14483, N1724);
or OR4 (N14514, N14509, N1920, N12201, N1298);
buf BUF1 (N14515, N14502);
or OR3 (N14516, N14513, N7005, N8207);
nand NAND3 (N14517, N14514, N3118, N10330);
not NOT1 (N14518, N14517);
nand NAND4 (N14519, N14498, N6627, N3789, N13967);
nand NAND3 (N14520, N14506, N4936, N499);
and AND4 (N14521, N14507, N8948, N10550, N9223);
not NOT1 (N14522, N14515);
nand NAND4 (N14523, N14511, N2810, N6476, N7623);
nand NAND4 (N14524, N14505, N11423, N3836, N3032);
or OR2 (N14525, N14512, N7929);
and AND3 (N14526, N14518, N4191, N1510);
or OR4 (N14527, N14522, N3798, N3085, N13080);
nand NAND3 (N14528, N14527, N9853, N9012);
buf BUF1 (N14529, N14526);
nand NAND4 (N14530, N14516, N13531, N8153, N12556);
nand NAND3 (N14531, N14510, N6984, N287);
not NOT1 (N14532, N14524);
buf BUF1 (N14533, N14523);
or OR2 (N14534, N14525, N10789);
and AND2 (N14535, N14531, N6225);
or OR3 (N14536, N14535, N4834, N7508);
nor NOR4 (N14537, N14530, N12436, N6460, N9876);
buf BUF1 (N14538, N14521);
or OR2 (N14539, N14534, N13278);
buf BUF1 (N14540, N14528);
not NOT1 (N14541, N14540);
or OR4 (N14542, N14539, N13334, N5355, N12371);
nand NAND3 (N14543, N14529, N4308, N5487);
xor XOR2 (N14544, N14537, N2547);
and AND3 (N14545, N14538, N3340, N11909);
nor NOR3 (N14546, N14532, N1882, N13845);
xor XOR2 (N14547, N14545, N12512);
xor XOR2 (N14548, N14546, N11835);
and AND3 (N14549, N14519, N3219, N11651);
buf BUF1 (N14550, N14543);
and AND4 (N14551, N14536, N2507, N12313, N6882);
and AND4 (N14552, N14544, N5121, N12116, N14428);
buf BUF1 (N14553, N14547);
nor NOR4 (N14554, N14553, N11697, N6550, N381);
xor XOR2 (N14555, N14551, N10459);
nor NOR4 (N14556, N14554, N12464, N6194, N9615);
or OR3 (N14557, N14548, N7498, N5401);
xor XOR2 (N14558, N14520, N9665);
not NOT1 (N14559, N14556);
and AND2 (N14560, N14558, N9079);
or OR4 (N14561, N14557, N4403, N13784, N10481);
and AND4 (N14562, N14552, N1363, N13307, N596);
or OR2 (N14563, N14549, N9911);
buf BUF1 (N14564, N14550);
or OR2 (N14565, N14555, N5491);
nor NOR3 (N14566, N14533, N7853, N11205);
or OR4 (N14567, N14541, N1495, N14444, N14406);
not NOT1 (N14568, N14564);
xor XOR2 (N14569, N14542, N14561);
or OR2 (N14570, N601, N3663);
and AND3 (N14571, N14566, N11205, N295);
or OR3 (N14572, N14560, N8040, N12234);
not NOT1 (N14573, N14572);
xor XOR2 (N14574, N14570, N5952);
nor NOR4 (N14575, N14573, N11198, N7773, N8769);
nor NOR2 (N14576, N14562, N2621);
and AND3 (N14577, N14569, N12748, N10505);
nand NAND4 (N14578, N14563, N515, N4741, N10490);
or OR4 (N14579, N14567, N14140, N10145, N14249);
nor NOR3 (N14580, N14575, N3453, N9015);
xor XOR2 (N14581, N14577, N8870);
buf BUF1 (N14582, N14571);
buf BUF1 (N14583, N14579);
or OR3 (N14584, N14581, N1647, N1153);
or OR2 (N14585, N14574, N10287);
buf BUF1 (N14586, N14568);
nand NAND3 (N14587, N14565, N7368, N12896);
buf BUF1 (N14588, N14559);
nand NAND4 (N14589, N14584, N10480, N14477, N6325);
xor XOR2 (N14590, N14589, N13494);
not NOT1 (N14591, N14588);
xor XOR2 (N14592, N14586, N14223);
nor NOR4 (N14593, N14580, N9674, N13250, N8833);
nand NAND3 (N14594, N14593, N860, N1124);
and AND2 (N14595, N14587, N44);
buf BUF1 (N14596, N14585);
buf BUF1 (N14597, N14591);
buf BUF1 (N14598, N14592);
nor NOR4 (N14599, N14576, N6358, N8237, N2597);
nor NOR3 (N14600, N14594, N13539, N5153);
buf BUF1 (N14601, N14583);
nor NOR4 (N14602, N14590, N6809, N2870, N4612);
not NOT1 (N14603, N14601);
and AND3 (N14604, N14598, N13869, N10067);
xor XOR2 (N14605, N14596, N6269);
nor NOR4 (N14606, N14600, N13504, N2355, N10638);
and AND2 (N14607, N14582, N10165);
xor XOR2 (N14608, N14599, N7049);
or OR4 (N14609, N14595, N5692, N1817, N4986);
or OR2 (N14610, N14607, N12413);
nand NAND4 (N14611, N14597, N6783, N2908, N9102);
or OR3 (N14612, N14609, N7939, N10728);
buf BUF1 (N14613, N14605);
or OR4 (N14614, N14612, N1549, N7340, N5035);
xor XOR2 (N14615, N14611, N11227);
xor XOR2 (N14616, N14613, N12313);
and AND4 (N14617, N14615, N1780, N11317, N7292);
or OR4 (N14618, N14604, N11629, N5126, N6371);
or OR3 (N14619, N14618, N10034, N1887);
buf BUF1 (N14620, N14603);
nor NOR2 (N14621, N14578, N4887);
or OR2 (N14622, N14621, N2915);
nand NAND3 (N14623, N14620, N13885, N7287);
buf BUF1 (N14624, N14616);
nand NAND4 (N14625, N14623, N4813, N8779, N4034);
nor NOR4 (N14626, N14622, N6616, N14057, N10919);
not NOT1 (N14627, N14602);
and AND2 (N14628, N14617, N9139);
not NOT1 (N14629, N14624);
and AND4 (N14630, N14629, N5990, N11037, N12303);
not NOT1 (N14631, N14626);
nor NOR3 (N14632, N14625, N368, N11060);
or OR3 (N14633, N14630, N7894, N9874);
not NOT1 (N14634, N14619);
nor NOR3 (N14635, N14631, N11642, N5656);
or OR3 (N14636, N14610, N355, N13368);
not NOT1 (N14637, N14635);
nand NAND4 (N14638, N14628, N9365, N4297, N7429);
nand NAND4 (N14639, N14634, N10263, N13153, N12331);
buf BUF1 (N14640, N14627);
or OR3 (N14641, N14606, N2804, N6895);
nand NAND4 (N14642, N14614, N1237, N7908, N557);
not NOT1 (N14643, N14642);
not NOT1 (N14644, N14633);
nor NOR3 (N14645, N14638, N13302, N8770);
nor NOR4 (N14646, N14639, N9091, N10763, N2955);
buf BUF1 (N14647, N14640);
nor NOR4 (N14648, N14646, N4313, N5320, N2535);
and AND3 (N14649, N14608, N7487, N2459);
nand NAND4 (N14650, N14632, N7478, N9121, N8524);
not NOT1 (N14651, N14648);
or OR2 (N14652, N14647, N1242);
and AND3 (N14653, N14636, N11625, N13747);
nand NAND2 (N14654, N14651, N7608);
not NOT1 (N14655, N14641);
nor NOR3 (N14656, N14652, N13217, N968);
xor XOR2 (N14657, N14650, N5202);
and AND2 (N14658, N14655, N5612);
or OR2 (N14659, N14656, N10328);
or OR2 (N14660, N14659, N14028);
and AND3 (N14661, N14657, N2609, N12330);
not NOT1 (N14662, N14645);
buf BUF1 (N14663, N14653);
or OR4 (N14664, N14637, N3398, N7786, N2722);
not NOT1 (N14665, N14662);
xor XOR2 (N14666, N14664, N2225);
or OR2 (N14667, N14644, N11800);
nor NOR4 (N14668, N14666, N11209, N3080, N12471);
or OR3 (N14669, N14668, N9878, N9567);
or OR2 (N14670, N14649, N12903);
buf BUF1 (N14671, N14661);
nand NAND3 (N14672, N14654, N7254, N6152);
and AND2 (N14673, N14671, N2614);
and AND3 (N14674, N14670, N12140, N14424);
nand NAND4 (N14675, N14660, N12355, N6767, N9903);
or OR2 (N14676, N14673, N2402);
nor NOR3 (N14677, N14672, N1528, N3172);
not NOT1 (N14678, N14676);
nor NOR4 (N14679, N14677, N10602, N7650, N12429);
xor XOR2 (N14680, N14658, N11079);
xor XOR2 (N14681, N14669, N1993);
or OR2 (N14682, N14663, N1652);
xor XOR2 (N14683, N14678, N12570);
not NOT1 (N14684, N14680);
nor NOR3 (N14685, N14667, N5606, N1492);
buf BUF1 (N14686, N14683);
and AND3 (N14687, N14674, N2450, N13616);
not NOT1 (N14688, N14643);
not NOT1 (N14689, N14684);
nand NAND4 (N14690, N14682, N11552, N12758, N11945);
nand NAND3 (N14691, N14688, N12597, N10258);
not NOT1 (N14692, N14675);
buf BUF1 (N14693, N14689);
buf BUF1 (N14694, N14665);
not NOT1 (N14695, N14691);
or OR4 (N14696, N14679, N5209, N223, N10404);
and AND3 (N14697, N14694, N1251, N14542);
not NOT1 (N14698, N14697);
buf BUF1 (N14699, N14692);
and AND2 (N14700, N14690, N8262);
and AND4 (N14701, N14695, N8098, N2172, N4351);
buf BUF1 (N14702, N14687);
and AND4 (N14703, N14686, N13300, N12460, N2867);
buf BUF1 (N14704, N14698);
and AND2 (N14705, N14700, N3276);
not NOT1 (N14706, N14701);
not NOT1 (N14707, N14704);
xor XOR2 (N14708, N14706, N4523);
nor NOR4 (N14709, N14705, N2809, N948, N5496);
xor XOR2 (N14710, N14685, N11979);
or OR2 (N14711, N14710, N12505);
xor XOR2 (N14712, N14702, N11657);
nor NOR4 (N14713, N14696, N10013, N2409, N8245);
xor XOR2 (N14714, N14693, N5086);
nor NOR2 (N14715, N14714, N2790);
xor XOR2 (N14716, N14709, N4637);
xor XOR2 (N14717, N14715, N5213);
xor XOR2 (N14718, N14707, N2207);
buf BUF1 (N14719, N14703);
nand NAND3 (N14720, N14713, N11892, N2500);
nand NAND2 (N14721, N14708, N5139);
not NOT1 (N14722, N14720);
or OR3 (N14723, N14719, N3554, N2774);
not NOT1 (N14724, N14716);
not NOT1 (N14725, N14722);
or OR4 (N14726, N14712, N2642, N6396, N3907);
xor XOR2 (N14727, N14723, N2597);
and AND3 (N14728, N14726, N11479, N6499);
not NOT1 (N14729, N14724);
or OR2 (N14730, N14699, N7485);
nor NOR4 (N14731, N14718, N1012, N10364, N10704);
buf BUF1 (N14732, N14730);
not NOT1 (N14733, N14711);
or OR4 (N14734, N14729, N4662, N10470, N13733);
nand NAND3 (N14735, N14734, N6858, N8534);
or OR4 (N14736, N14735, N8229, N12585, N6382);
not NOT1 (N14737, N14732);
not NOT1 (N14738, N14728);
not NOT1 (N14739, N14733);
not NOT1 (N14740, N14731);
and AND4 (N14741, N14739, N3697, N13830, N7781);
and AND4 (N14742, N14681, N8632, N11221, N1642);
xor XOR2 (N14743, N14741, N4255);
xor XOR2 (N14744, N14740, N1391);
buf BUF1 (N14745, N14736);
nor NOR4 (N14746, N14743, N12469, N13293, N13961);
xor XOR2 (N14747, N14717, N9774);
nand NAND4 (N14748, N14744, N1754, N1773, N6616);
nor NOR4 (N14749, N14746, N3079, N14061, N895);
not NOT1 (N14750, N14738);
or OR2 (N14751, N14747, N14098);
xor XOR2 (N14752, N14749, N4620);
nand NAND4 (N14753, N14752, N9421, N8377, N12454);
nand NAND3 (N14754, N14725, N3230, N1934);
or OR3 (N14755, N14751, N5165, N7069);
and AND4 (N14756, N14748, N12441, N4774, N13575);
and AND2 (N14757, N14742, N10192);
and AND2 (N14758, N14737, N2821);
buf BUF1 (N14759, N14721);
not NOT1 (N14760, N14755);
buf BUF1 (N14761, N14758);
nand NAND3 (N14762, N14750, N499, N8266);
and AND3 (N14763, N14760, N9583, N4033);
or OR3 (N14764, N14745, N14736, N9140);
nor NOR4 (N14765, N14761, N3477, N8559, N11192);
and AND4 (N14766, N14756, N6099, N9112, N8592);
not NOT1 (N14767, N14759);
or OR3 (N14768, N14766, N9461, N5949);
not NOT1 (N14769, N14764);
nand NAND4 (N14770, N14767, N9224, N12002, N13076);
or OR4 (N14771, N14762, N6777, N7952, N14145);
or OR4 (N14772, N14757, N12488, N3432, N6028);
and AND4 (N14773, N14771, N4586, N3939, N12819);
nor NOR4 (N14774, N14768, N6468, N10524, N2823);
nand NAND2 (N14775, N14770, N2829);
buf BUF1 (N14776, N14754);
nor NOR4 (N14777, N14765, N11022, N8786, N1457);
or OR4 (N14778, N14774, N6601, N10931, N10085);
nand NAND4 (N14779, N14727, N7641, N14527, N12354);
nand NAND4 (N14780, N14777, N13167, N4348, N8922);
nor NOR3 (N14781, N14780, N663, N7939);
buf BUF1 (N14782, N14775);
or OR4 (N14783, N14779, N14508, N2559, N11367);
xor XOR2 (N14784, N14772, N1862);
xor XOR2 (N14785, N14782, N1327);
buf BUF1 (N14786, N14778);
nor NOR4 (N14787, N14776, N7767, N5948, N2339);
not NOT1 (N14788, N14773);
nand NAND4 (N14789, N14787, N5298, N14106, N13322);
not NOT1 (N14790, N14763);
not NOT1 (N14791, N14769);
and AND3 (N14792, N14786, N11216, N3329);
nand NAND4 (N14793, N14789, N6186, N8071, N12078);
nor NOR3 (N14794, N14784, N6256, N11589);
buf BUF1 (N14795, N14793);
not NOT1 (N14796, N14790);
xor XOR2 (N14797, N14795, N12436);
xor XOR2 (N14798, N14794, N1137);
and AND4 (N14799, N14785, N10551, N9375, N4779);
or OR4 (N14800, N14781, N4710, N5664, N2665);
xor XOR2 (N14801, N14798, N3844);
nand NAND3 (N14802, N14796, N11562, N9039);
xor XOR2 (N14803, N14799, N12590);
and AND3 (N14804, N14788, N4127, N6642);
not NOT1 (N14805, N14801);
nand NAND3 (N14806, N14800, N7355, N499);
xor XOR2 (N14807, N14791, N2103);
xor XOR2 (N14808, N14803, N10034);
xor XOR2 (N14809, N14805, N8858);
not NOT1 (N14810, N14753);
nand NAND2 (N14811, N14806, N7927);
nor NOR3 (N14812, N14807, N693, N7367);
and AND2 (N14813, N14812, N2677);
not NOT1 (N14814, N14792);
buf BUF1 (N14815, N14804);
and AND2 (N14816, N14813, N9912);
and AND2 (N14817, N14808, N6092);
xor XOR2 (N14818, N14802, N10509);
nor NOR4 (N14819, N14815, N2190, N7223, N872);
xor XOR2 (N14820, N14817, N6362);
not NOT1 (N14821, N14818);
buf BUF1 (N14822, N14809);
and AND4 (N14823, N14810, N5288, N3151, N3571);
nand NAND2 (N14824, N14797, N6717);
nor NOR2 (N14825, N14816, N9520);
nor NOR2 (N14826, N14823, N82);
nand NAND2 (N14827, N14783, N1601);
or OR4 (N14828, N14814, N11941, N11400, N14051);
xor XOR2 (N14829, N14821, N13208);
or OR2 (N14830, N14811, N9159);
nand NAND3 (N14831, N14830, N3873, N12474);
xor XOR2 (N14832, N14828, N13757);
nand NAND4 (N14833, N14832, N483, N8665, N8346);
xor XOR2 (N14834, N14824, N4705);
xor XOR2 (N14835, N14829, N8374);
nand NAND2 (N14836, N14827, N10623);
and AND3 (N14837, N14833, N12120, N881);
and AND3 (N14838, N14835, N1442, N3376);
nor NOR3 (N14839, N14831, N7412, N13395);
not NOT1 (N14840, N14838);
and AND4 (N14841, N14837, N1664, N9941, N5763);
or OR4 (N14842, N14839, N1931, N10414, N5104);
and AND2 (N14843, N14825, N12084);
nor NOR2 (N14844, N14841, N5494);
nand NAND2 (N14845, N14834, N764);
or OR3 (N14846, N14822, N5663, N4680);
nand NAND2 (N14847, N14845, N4640);
nor NOR2 (N14848, N14826, N4561);
nand NAND2 (N14849, N14842, N5215);
and AND4 (N14850, N14847, N7791, N12975, N4307);
nand NAND4 (N14851, N14849, N7961, N6140, N10769);
buf BUF1 (N14852, N14840);
buf BUF1 (N14853, N14836);
and AND2 (N14854, N14853, N12342);
xor XOR2 (N14855, N14854, N12212);
and AND3 (N14856, N14855, N9203, N8242);
and AND2 (N14857, N14851, N8212);
nor NOR2 (N14858, N14857, N1601);
not NOT1 (N14859, N14852);
xor XOR2 (N14860, N14819, N9582);
nand NAND4 (N14861, N14858, N3721, N11905, N7508);
xor XOR2 (N14862, N14848, N3900);
or OR3 (N14863, N14820, N10038, N6788);
or OR4 (N14864, N14862, N9917, N1404, N3087);
buf BUF1 (N14865, N14843);
nor NOR4 (N14866, N14863, N11373, N6045, N1355);
nor NOR3 (N14867, N14864, N3060, N3010);
and AND4 (N14868, N14866, N946, N13980, N8098);
nor NOR4 (N14869, N14850, N10181, N11079, N4899);
nor NOR4 (N14870, N14859, N3426, N5762, N9100);
buf BUF1 (N14871, N14860);
xor XOR2 (N14872, N14868, N6772);
or OR3 (N14873, N14844, N14020, N13189);
or OR3 (N14874, N14870, N12203, N8963);
xor XOR2 (N14875, N14846, N7681);
nand NAND4 (N14876, N14871, N1698, N2336, N12155);
xor XOR2 (N14877, N14861, N11010);
or OR3 (N14878, N14876, N4475, N14459);
buf BUF1 (N14879, N14877);
and AND2 (N14880, N14856, N9387);
nand NAND4 (N14881, N14869, N10758, N6069, N5980);
and AND2 (N14882, N14878, N14113);
xor XOR2 (N14883, N14882, N12339);
and AND3 (N14884, N14873, N12279, N12902);
buf BUF1 (N14885, N14874);
and AND3 (N14886, N14880, N4500, N8965);
and AND3 (N14887, N14885, N11891, N3342);
or OR3 (N14888, N14875, N4917, N10234);
not NOT1 (N14889, N14887);
or OR4 (N14890, N14879, N10982, N4840, N2701);
xor XOR2 (N14891, N14881, N5086);
or OR3 (N14892, N14872, N3350, N5615);
or OR4 (N14893, N14883, N6843, N12265, N2161);
nand NAND3 (N14894, N14892, N3355, N9728);
and AND3 (N14895, N14893, N11367, N14199);
xor XOR2 (N14896, N14865, N2079);
nor NOR4 (N14897, N14895, N11544, N3389, N2745);
and AND3 (N14898, N14889, N12157, N13194);
not NOT1 (N14899, N14890);
not NOT1 (N14900, N14891);
buf BUF1 (N14901, N14888);
and AND2 (N14902, N14894, N10609);
buf BUF1 (N14903, N14899);
nand NAND4 (N14904, N14896, N1285, N12806, N6580);
and AND4 (N14905, N14902, N8436, N3200, N4983);
nand NAND4 (N14906, N14905, N9236, N5850, N2966);
not NOT1 (N14907, N14904);
nor NOR3 (N14908, N14886, N8101, N3864);
buf BUF1 (N14909, N14906);
buf BUF1 (N14910, N14900);
buf BUF1 (N14911, N14867);
not NOT1 (N14912, N14903);
and AND3 (N14913, N14912, N10210, N6713);
not NOT1 (N14914, N14898);
and AND4 (N14915, N14901, N12646, N7127, N10090);
not NOT1 (N14916, N14914);
nand NAND3 (N14917, N14909, N7537, N13028);
or OR4 (N14918, N14913, N6044, N6373, N9668);
not NOT1 (N14919, N14918);
nor NOR4 (N14920, N14897, N7442, N11628, N13810);
or OR2 (N14921, N14916, N10798);
nand NAND3 (N14922, N14908, N14829, N5440);
xor XOR2 (N14923, N14919, N4015);
and AND3 (N14924, N14921, N9529, N9837);
buf BUF1 (N14925, N14884);
or OR2 (N14926, N14920, N105);
nor NOR4 (N14927, N14923, N13053, N843, N3305);
and AND2 (N14928, N14922, N9535);
not NOT1 (N14929, N14917);
and AND2 (N14930, N14911, N8580);
buf BUF1 (N14931, N14926);
buf BUF1 (N14932, N14928);
nor NOR4 (N14933, N14925, N14566, N1131, N14431);
buf BUF1 (N14934, N14927);
not NOT1 (N14935, N14931);
and AND4 (N14936, N14929, N6155, N5902, N3798);
or OR4 (N14937, N14915, N3565, N9534, N4893);
not NOT1 (N14938, N14936);
nor NOR4 (N14939, N14937, N9173, N9183, N4900);
buf BUF1 (N14940, N14930);
and AND3 (N14941, N14938, N855, N10804);
nor NOR4 (N14942, N14933, N1115, N14883, N12914);
nand NAND4 (N14943, N14932, N2034, N10678, N11073);
or OR4 (N14944, N14910, N5712, N5451, N14935);
nor NOR3 (N14945, N11125, N9885, N12384);
nor NOR2 (N14946, N14942, N10523);
not NOT1 (N14947, N14907);
and AND4 (N14948, N14924, N8004, N733, N8620);
or OR4 (N14949, N14944, N8018, N11109, N8671);
xor XOR2 (N14950, N14945, N4137);
nand NAND2 (N14951, N14947, N14711);
nor NOR3 (N14952, N14946, N5502, N7941);
and AND4 (N14953, N14934, N10427, N4041, N14128);
xor XOR2 (N14954, N14943, N8718);
not NOT1 (N14955, N14940);
buf BUF1 (N14956, N14939);
not NOT1 (N14957, N14941);
or OR2 (N14958, N14950, N5441);
not NOT1 (N14959, N14949);
or OR3 (N14960, N14954, N12869, N3608);
or OR2 (N14961, N14959, N4954);
nor NOR2 (N14962, N14956, N9590);
buf BUF1 (N14963, N14952);
xor XOR2 (N14964, N14957, N6872);
or OR2 (N14965, N14961, N2457);
nand NAND2 (N14966, N14951, N6607);
or OR4 (N14967, N14965, N3419, N8664, N5554);
nor NOR4 (N14968, N14948, N1716, N528, N5337);
buf BUF1 (N14969, N14963);
nand NAND4 (N14970, N14969, N10195, N14469, N13459);
and AND2 (N14971, N14953, N13259);
not NOT1 (N14972, N14970);
and AND2 (N14973, N14960, N3132);
nand NAND4 (N14974, N14968, N9512, N8580, N6141);
xor XOR2 (N14975, N14967, N7970);
buf BUF1 (N14976, N14962);
not NOT1 (N14977, N14973);
and AND4 (N14978, N14976, N3286, N4456, N608);
xor XOR2 (N14979, N14955, N12125);
not NOT1 (N14980, N14958);
nor NOR4 (N14981, N14978, N8927, N13849, N12026);
nand NAND4 (N14982, N14980, N211, N4226, N11751);
and AND2 (N14983, N14977, N1518);
buf BUF1 (N14984, N14979);
buf BUF1 (N14985, N14971);
buf BUF1 (N14986, N14974);
or OR2 (N14987, N14983, N5490);
buf BUF1 (N14988, N14981);
or OR2 (N14989, N14985, N13376);
and AND2 (N14990, N14972, N13022);
nand NAND2 (N14991, N14966, N2380);
and AND3 (N14992, N14991, N10475, N10135);
nor NOR2 (N14993, N14987, N8017);
buf BUF1 (N14994, N14986);
or OR2 (N14995, N14993, N2767);
or OR4 (N14996, N14984, N8028, N8448, N14701);
not NOT1 (N14997, N14988);
nand NAND3 (N14998, N14990, N14258, N14647);
or OR2 (N14999, N14997, N12787);
buf BUF1 (N15000, N14982);
or OR2 (N15001, N14964, N12264);
buf BUF1 (N15002, N15000);
or OR4 (N15003, N15001, N10548, N8155, N14661);
not NOT1 (N15004, N15002);
nor NOR3 (N15005, N14994, N3823, N8033);
nand NAND4 (N15006, N14992, N175, N2124, N4612);
not NOT1 (N15007, N14989);
not NOT1 (N15008, N15003);
or OR2 (N15009, N15007, N9094);
or OR4 (N15010, N14996, N11413, N362, N1131);
nor NOR4 (N15011, N15009, N8480, N2114, N1737);
nor NOR2 (N15012, N15006, N8018);
not NOT1 (N15013, N14998);
not NOT1 (N15014, N15004);
buf BUF1 (N15015, N15005);
buf BUF1 (N15016, N15014);
buf BUF1 (N15017, N14995);
xor XOR2 (N15018, N15015, N4003);
and AND3 (N15019, N15011, N11029, N5474);
or OR4 (N15020, N15018, N13654, N14108, N13999);
nand NAND2 (N15021, N15008, N6906);
and AND4 (N15022, N15020, N4993, N8813, N14435);
or OR4 (N15023, N15021, N8683, N13580, N10898);
nand NAND3 (N15024, N15019, N2885, N4025);
or OR3 (N15025, N15024, N2524, N6589);
not NOT1 (N15026, N15012);
nand NAND3 (N15027, N15023, N8876, N3072);
nand NAND4 (N15028, N15026, N3641, N8681, N12322);
xor XOR2 (N15029, N15016, N3208);
nor NOR2 (N15030, N15022, N11847);
buf BUF1 (N15031, N15017);
nor NOR4 (N15032, N15031, N10209, N1375, N14139);
or OR3 (N15033, N15032, N7859, N1076);
and AND4 (N15034, N14975, N6023, N642, N186);
and AND4 (N15035, N15028, N317, N4426, N11945);
buf BUF1 (N15036, N15030);
nand NAND4 (N15037, N15035, N5469, N12740, N6117);
or OR4 (N15038, N15034, N1407, N11934, N11848);
nand NAND2 (N15039, N15033, N9939);
buf BUF1 (N15040, N15038);
xor XOR2 (N15041, N15013, N6396);
xor XOR2 (N15042, N15025, N11377);
buf BUF1 (N15043, N15037);
xor XOR2 (N15044, N15041, N811);
nor NOR4 (N15045, N15029, N1014, N5711, N4994);
xor XOR2 (N15046, N15039, N8327);
xor XOR2 (N15047, N15045, N12837);
xor XOR2 (N15048, N15040, N9650);
xor XOR2 (N15049, N15043, N13480);
nor NOR3 (N15050, N15046, N9347, N11660);
and AND4 (N15051, N15048, N7704, N9597, N4438);
or OR4 (N15052, N15044, N9149, N5126, N12777);
xor XOR2 (N15053, N15047, N1700);
xor XOR2 (N15054, N15036, N4823);
xor XOR2 (N15055, N15050, N14324);
nor NOR2 (N15056, N15053, N1643);
or OR2 (N15057, N15010, N2902);
nor NOR2 (N15058, N15054, N34);
not NOT1 (N15059, N15058);
xor XOR2 (N15060, N15049, N14186);
nand NAND4 (N15061, N15056, N12860, N14110, N11490);
buf BUF1 (N15062, N15059);
and AND2 (N15063, N15057, N6645);
xor XOR2 (N15064, N14999, N14822);
not NOT1 (N15065, N15064);
xor XOR2 (N15066, N15027, N3291);
nor NOR4 (N15067, N15052, N14870, N11087, N5698);
xor XOR2 (N15068, N15060, N9270);
xor XOR2 (N15069, N15055, N8734);
and AND3 (N15070, N15063, N11170, N7171);
or OR4 (N15071, N15062, N2675, N13539, N1163);
nand NAND4 (N15072, N15070, N3442, N5236, N1313);
not NOT1 (N15073, N15065);
not NOT1 (N15074, N15042);
or OR3 (N15075, N15074, N1888, N11071);
or OR3 (N15076, N15069, N7432, N8288);
xor XOR2 (N15077, N15072, N2623);
nand NAND3 (N15078, N15066, N8336, N11998);
not NOT1 (N15079, N15068);
or OR3 (N15080, N15076, N10515, N14470);
buf BUF1 (N15081, N15077);
nand NAND4 (N15082, N15079, N12885, N2734, N1882);
or OR3 (N15083, N15082, N13739, N416);
buf BUF1 (N15084, N15061);
not NOT1 (N15085, N15083);
nor NOR4 (N15086, N15051, N12829, N11567, N10475);
or OR3 (N15087, N15086, N8448, N7024);
and AND4 (N15088, N15075, N3660, N11672, N13653);
nor NOR3 (N15089, N15080, N11081, N2508);
nor NOR3 (N15090, N15081, N3325, N491);
or OR4 (N15091, N15078, N412, N12946, N10994);
nor NOR2 (N15092, N15085, N2324);
nand NAND3 (N15093, N15089, N5523, N13989);
buf BUF1 (N15094, N15091);
buf BUF1 (N15095, N15093);
nor NOR3 (N15096, N15084, N12370, N5141);
buf BUF1 (N15097, N15073);
nand NAND4 (N15098, N15071, N12278, N10582, N5969);
buf BUF1 (N15099, N15096);
nand NAND3 (N15100, N15090, N6439, N2136);
xor XOR2 (N15101, N15097, N13715);
buf BUF1 (N15102, N15099);
and AND2 (N15103, N15102, N4370);
not NOT1 (N15104, N15094);
xor XOR2 (N15105, N15104, N7199);
or OR3 (N15106, N15100, N7107, N427);
nor NOR2 (N15107, N15087, N14832);
and AND3 (N15108, N15092, N13416, N8981);
not NOT1 (N15109, N15105);
xor XOR2 (N15110, N15098, N8511);
nor NOR3 (N15111, N15107, N4374, N11453);
and AND4 (N15112, N15109, N11199, N8567, N5508);
nand NAND2 (N15113, N15108, N14697);
buf BUF1 (N15114, N15101);
and AND4 (N15115, N15067, N1443, N6426, N2833);
nor NOR4 (N15116, N15088, N667, N5501, N6649);
buf BUF1 (N15117, N15095);
xor XOR2 (N15118, N15112, N1255);
buf BUF1 (N15119, N15118);
or OR4 (N15120, N15111, N12585, N7663, N13508);
buf BUF1 (N15121, N15117);
xor XOR2 (N15122, N15115, N2092);
buf BUF1 (N15123, N15119);
nand NAND2 (N15124, N15110, N3427);
nor NOR4 (N15125, N15123, N10016, N959, N1670);
nand NAND2 (N15126, N15120, N7220);
or OR4 (N15127, N15113, N1807, N2626, N14989);
not NOT1 (N15128, N15116);
and AND3 (N15129, N15127, N1527, N8468);
nand NAND4 (N15130, N15103, N3075, N5272, N4415);
xor XOR2 (N15131, N15106, N13794);
not NOT1 (N15132, N15131);
nand NAND4 (N15133, N15125, N5269, N813, N6992);
and AND2 (N15134, N15128, N14239);
nand NAND2 (N15135, N15133, N5263);
nor NOR2 (N15136, N15121, N11346);
or OR3 (N15137, N15136, N7118, N4711);
buf BUF1 (N15138, N15122);
xor XOR2 (N15139, N15137, N12386);
not NOT1 (N15140, N15126);
not NOT1 (N15141, N15135);
nand NAND4 (N15142, N15139, N12894, N14592, N6371);
buf BUF1 (N15143, N15130);
buf BUF1 (N15144, N15134);
and AND3 (N15145, N15138, N1374, N14884);
nor NOR4 (N15146, N15143, N14639, N7197, N2865);
not NOT1 (N15147, N15141);
buf BUF1 (N15148, N15129);
nand NAND2 (N15149, N15145, N4833);
buf BUF1 (N15150, N15148);
and AND3 (N15151, N15149, N14539, N12717);
xor XOR2 (N15152, N15150, N3791);
and AND3 (N15153, N15124, N1864, N5314);
xor XOR2 (N15154, N15153, N7347);
nand NAND3 (N15155, N15144, N13336, N1444);
or OR2 (N15156, N15154, N11808);
and AND2 (N15157, N15147, N7399);
not NOT1 (N15158, N15140);
nor NOR2 (N15159, N15155, N5853);
or OR4 (N15160, N15132, N12931, N14928, N11720);
or OR3 (N15161, N15160, N9384, N11642);
and AND4 (N15162, N15161, N5575, N1902, N2739);
xor XOR2 (N15163, N15151, N14569);
xor XOR2 (N15164, N15162, N1635);
buf BUF1 (N15165, N15152);
buf BUF1 (N15166, N15164);
not NOT1 (N15167, N15163);
xor XOR2 (N15168, N15156, N6386);
xor XOR2 (N15169, N15166, N6902);
not NOT1 (N15170, N15157);
and AND2 (N15171, N15159, N6832);
not NOT1 (N15172, N15158);
and AND4 (N15173, N15165, N3761, N7421, N4596);
nand NAND4 (N15174, N15171, N6145, N13187, N8839);
buf BUF1 (N15175, N15168);
or OR2 (N15176, N15173, N9175);
nor NOR3 (N15177, N15169, N3681, N3005);
nand NAND3 (N15178, N15142, N13553, N11010);
not NOT1 (N15179, N15172);
not NOT1 (N15180, N15179);
nor NOR3 (N15181, N15177, N2192, N1709);
xor XOR2 (N15182, N15167, N8026);
nor NOR3 (N15183, N15181, N5182, N10152);
nor NOR3 (N15184, N15182, N1, N7909);
buf BUF1 (N15185, N15175);
nor NOR2 (N15186, N15114, N5547);
nand NAND3 (N15187, N15184, N6728, N9747);
buf BUF1 (N15188, N15183);
nand NAND4 (N15189, N15176, N1821, N10436, N8193);
and AND2 (N15190, N15187, N11381);
or OR2 (N15191, N15180, N6983);
not NOT1 (N15192, N15146);
and AND4 (N15193, N15189, N4410, N13296, N9398);
nor NOR2 (N15194, N15188, N11125);
xor XOR2 (N15195, N15190, N4149);
and AND2 (N15196, N15185, N204);
nand NAND2 (N15197, N15191, N5912);
xor XOR2 (N15198, N15193, N5742);
nand NAND3 (N15199, N15198, N11216, N2810);
or OR2 (N15200, N15196, N3615);
nor NOR3 (N15201, N15199, N12689, N348);
or OR4 (N15202, N15194, N10209, N13595, N4558);
and AND2 (N15203, N15186, N10774);
not NOT1 (N15204, N15195);
and AND3 (N15205, N15203, N13822, N9263);
nor NOR4 (N15206, N15178, N9592, N6647, N11267);
not NOT1 (N15207, N15202);
nand NAND2 (N15208, N15204, N7111);
xor XOR2 (N15209, N15174, N8254);
xor XOR2 (N15210, N15200, N10248);
and AND2 (N15211, N15210, N1194);
xor XOR2 (N15212, N15207, N10408);
or OR4 (N15213, N15211, N8665, N7764, N13519);
nand NAND3 (N15214, N15208, N12516, N12730);
xor XOR2 (N15215, N15213, N6391);
or OR4 (N15216, N15212, N4701, N4555, N1005);
or OR2 (N15217, N15201, N1632);
or OR3 (N15218, N15214, N260, N5199);
and AND4 (N15219, N15218, N2880, N1528, N6858);
and AND3 (N15220, N15216, N3345, N4527);
buf BUF1 (N15221, N15215);
not NOT1 (N15222, N15209);
and AND2 (N15223, N15220, N622);
or OR3 (N15224, N15222, N3828, N8954);
and AND4 (N15225, N15170, N5305, N13770, N10123);
not NOT1 (N15226, N15217);
nor NOR3 (N15227, N15225, N2028, N4472);
not NOT1 (N15228, N15205);
or OR2 (N15229, N15227, N7654);
or OR2 (N15230, N15224, N8351);
buf BUF1 (N15231, N15221);
or OR4 (N15232, N15228, N1398, N17, N13154);
and AND4 (N15233, N15206, N4359, N3567, N8331);
nor NOR2 (N15234, N15232, N13571);
or OR4 (N15235, N15192, N6362, N5006, N9799);
or OR3 (N15236, N15233, N8961, N7665);
nand NAND4 (N15237, N15230, N2786, N7033, N10495);
buf BUF1 (N15238, N15219);
nand NAND2 (N15239, N15236, N13431);
not NOT1 (N15240, N15229);
nor NOR2 (N15241, N15240, N5611);
and AND2 (N15242, N15237, N2844);
or OR4 (N15243, N15197, N4071, N13517, N7673);
buf BUF1 (N15244, N15234);
and AND4 (N15245, N15226, N9716, N13972, N10958);
buf BUF1 (N15246, N15241);
nor NOR4 (N15247, N15245, N3897, N12807, N10094);
nand NAND3 (N15248, N15239, N1997, N6882);
nand NAND4 (N15249, N15223, N6965, N2319, N8345);
not NOT1 (N15250, N15238);
or OR4 (N15251, N15248, N11231, N14257, N11536);
not NOT1 (N15252, N15242);
nand NAND2 (N15253, N15251, N6751);
buf BUF1 (N15254, N15244);
and AND4 (N15255, N15253, N2378, N13783, N10449);
and AND2 (N15256, N15235, N2077);
buf BUF1 (N15257, N15231);
or OR3 (N15258, N15246, N13650, N3734);
not NOT1 (N15259, N15255);
xor XOR2 (N15260, N15259, N8009);
xor XOR2 (N15261, N15247, N2380);
nand NAND3 (N15262, N15258, N1155, N3092);
buf BUF1 (N15263, N15256);
or OR4 (N15264, N15262, N8983, N2261, N11856);
and AND4 (N15265, N15254, N52, N12340, N8157);
nand NAND3 (N15266, N15243, N4531, N805);
xor XOR2 (N15267, N15260, N3834);
buf BUF1 (N15268, N15257);
and AND2 (N15269, N15267, N7377);
not NOT1 (N15270, N15261);
nor NOR2 (N15271, N15249, N11502);
buf BUF1 (N15272, N15263);
not NOT1 (N15273, N15269);
or OR3 (N15274, N15270, N8893, N7020);
or OR3 (N15275, N15250, N8507, N10982);
buf BUF1 (N15276, N15268);
or OR2 (N15277, N15264, N7820);
and AND2 (N15278, N15271, N11150);
xor XOR2 (N15279, N15265, N3724);
not NOT1 (N15280, N15272);
xor XOR2 (N15281, N15277, N749);
nand NAND4 (N15282, N15281, N6307, N14419, N9838);
and AND3 (N15283, N15274, N1231, N7813);
nand NAND3 (N15284, N15252, N7479, N15075);
nor NOR2 (N15285, N15284, N6091);
or OR3 (N15286, N15266, N5233, N3005);
or OR2 (N15287, N15282, N4303);
or OR2 (N15288, N15279, N8028);
and AND3 (N15289, N15285, N14709, N3682);
xor XOR2 (N15290, N15289, N10892);
and AND4 (N15291, N15278, N8580, N5320, N5594);
xor XOR2 (N15292, N15283, N8037);
nor NOR3 (N15293, N15292, N1865, N8414);
xor XOR2 (N15294, N15286, N4608);
xor XOR2 (N15295, N15288, N13923);
and AND4 (N15296, N15276, N11540, N7372, N7086);
nand NAND4 (N15297, N15293, N1927, N7248, N15135);
buf BUF1 (N15298, N15297);
not NOT1 (N15299, N15294);
nand NAND4 (N15300, N15295, N8034, N7394, N10980);
or OR3 (N15301, N15290, N10386, N3769);
and AND4 (N15302, N15280, N12302, N4609, N9355);
xor XOR2 (N15303, N15273, N6175);
not NOT1 (N15304, N15302);
and AND3 (N15305, N15299, N13671, N4993);
nor NOR2 (N15306, N15275, N10204);
or OR4 (N15307, N15296, N6399, N5287, N5679);
or OR4 (N15308, N15291, N7052, N7538, N9005);
or OR2 (N15309, N15298, N9301);
nand NAND4 (N15310, N15308, N13337, N11094, N6456);
not NOT1 (N15311, N15304);
and AND3 (N15312, N15307, N4710, N8093);
and AND3 (N15313, N15306, N8464, N12210);
xor XOR2 (N15314, N15313, N9948);
and AND4 (N15315, N15303, N1368, N12874, N11446);
not NOT1 (N15316, N15309);
buf BUF1 (N15317, N15316);
nor NOR3 (N15318, N15311, N7445, N15086);
buf BUF1 (N15319, N15317);
or OR2 (N15320, N15319, N1769);
nor NOR3 (N15321, N15305, N12261, N6882);
xor XOR2 (N15322, N15287, N3493);
xor XOR2 (N15323, N15312, N12579);
nor NOR4 (N15324, N15301, N276, N9793, N271);
xor XOR2 (N15325, N15318, N2304);
xor XOR2 (N15326, N15314, N1006);
nor NOR2 (N15327, N15324, N10408);
or OR4 (N15328, N15322, N11625, N4699, N8198);
xor XOR2 (N15329, N15323, N5309);
buf BUF1 (N15330, N15300);
buf BUF1 (N15331, N15326);
nor NOR3 (N15332, N15330, N5904, N8309);
and AND2 (N15333, N15310, N13854);
not NOT1 (N15334, N15333);
buf BUF1 (N15335, N15332);
nand NAND4 (N15336, N15328, N10797, N13309, N11794);
nand NAND4 (N15337, N15325, N1826, N6834, N12555);
nand NAND4 (N15338, N15334, N2055, N1390, N4572);
nor NOR4 (N15339, N15338, N1646, N10094, N13693);
or OR2 (N15340, N15335, N5270);
and AND4 (N15341, N15321, N5225, N12916, N12682);
buf BUF1 (N15342, N15315);
buf BUF1 (N15343, N15340);
nor NOR4 (N15344, N15336, N1632, N1065, N3707);
xor XOR2 (N15345, N15331, N4671);
and AND2 (N15346, N15342, N7963);
xor XOR2 (N15347, N15337, N13727);
not NOT1 (N15348, N15343);
xor XOR2 (N15349, N15345, N3065);
buf BUF1 (N15350, N15347);
nor NOR4 (N15351, N15327, N2916, N9318, N10932);
nand NAND3 (N15352, N15344, N13398, N12740);
nand NAND2 (N15353, N15339, N9476);
xor XOR2 (N15354, N15329, N312);
buf BUF1 (N15355, N15350);
buf BUF1 (N15356, N15355);
buf BUF1 (N15357, N15349);
or OR2 (N15358, N15357, N7230);
buf BUF1 (N15359, N15348);
nand NAND2 (N15360, N15346, N13653);
nor NOR3 (N15361, N15358, N5475, N10158);
nor NOR2 (N15362, N15356, N7593);
xor XOR2 (N15363, N15351, N14064);
xor XOR2 (N15364, N15354, N6914);
buf BUF1 (N15365, N15360);
xor XOR2 (N15366, N15365, N3738);
nand NAND4 (N15367, N15353, N1996, N959, N13973);
nor NOR3 (N15368, N15341, N14613, N718);
not NOT1 (N15369, N15366);
and AND3 (N15370, N15364, N12408, N5927);
xor XOR2 (N15371, N15363, N10483);
nor NOR2 (N15372, N15359, N14260);
buf BUF1 (N15373, N15320);
nor NOR3 (N15374, N15371, N3191, N9);
buf BUF1 (N15375, N15372);
nor NOR4 (N15376, N15367, N4961, N6650, N8008);
not NOT1 (N15377, N15361);
nand NAND2 (N15378, N15352, N11967);
and AND3 (N15379, N15368, N11705, N9113);
nand NAND3 (N15380, N15374, N7136, N5874);
xor XOR2 (N15381, N15373, N7033);
nor NOR2 (N15382, N15377, N11816);
and AND4 (N15383, N15376, N1909, N12194, N14629);
or OR4 (N15384, N15381, N6802, N13433, N1322);
xor XOR2 (N15385, N15369, N14201);
xor XOR2 (N15386, N15370, N5331);
buf BUF1 (N15387, N15379);
and AND2 (N15388, N15362, N12705);
nor NOR4 (N15389, N15380, N3112, N6395, N3671);
not NOT1 (N15390, N15378);
or OR2 (N15391, N15387, N1465);
and AND3 (N15392, N15391, N2390, N11948);
and AND4 (N15393, N15386, N5345, N1917, N2636);
nor NOR2 (N15394, N15384, N9655);
or OR2 (N15395, N15393, N447);
and AND3 (N15396, N15388, N12276, N14286);
buf BUF1 (N15397, N15390);
buf BUF1 (N15398, N15397);
or OR4 (N15399, N15392, N8757, N9429, N13836);
nor NOR3 (N15400, N15382, N14743, N14937);
xor XOR2 (N15401, N15399, N11947);
buf BUF1 (N15402, N15385);
nor NOR2 (N15403, N15398, N2530);
nor NOR2 (N15404, N15401, N7444);
buf BUF1 (N15405, N15394);
or OR3 (N15406, N15405, N11314, N6858);
nand NAND3 (N15407, N15395, N409, N5791);
buf BUF1 (N15408, N15407);
not NOT1 (N15409, N15403);
not NOT1 (N15410, N15396);
xor XOR2 (N15411, N15389, N1757);
nand NAND2 (N15412, N15406, N8238);
nor NOR3 (N15413, N15412, N3303, N11117);
nor NOR4 (N15414, N15411, N7518, N11985, N5009);
or OR3 (N15415, N15408, N9679, N6562);
or OR4 (N15416, N15400, N1657, N9777, N7515);
buf BUF1 (N15417, N15410);
nor NOR3 (N15418, N15375, N13334, N9219);
xor XOR2 (N15419, N15409, N3182);
or OR2 (N15420, N15416, N7262);
not NOT1 (N15421, N15418);
nor NOR2 (N15422, N15414, N9262);
nor NOR4 (N15423, N15402, N8501, N6571, N1791);
nor NOR4 (N15424, N15423, N2697, N7109, N10761);
not NOT1 (N15425, N15404);
xor XOR2 (N15426, N15420, N6064);
not NOT1 (N15427, N15421);
or OR2 (N15428, N15383, N6344);
or OR3 (N15429, N15413, N8984, N2023);
nand NAND4 (N15430, N15425, N10981, N11913, N9137);
nand NAND3 (N15431, N15417, N5845, N99);
xor XOR2 (N15432, N15424, N10199);
nor NOR4 (N15433, N15428, N10795, N5837, N12965);
buf BUF1 (N15434, N15432);
not NOT1 (N15435, N15415);
buf BUF1 (N15436, N15430);
not NOT1 (N15437, N15429);
not NOT1 (N15438, N15419);
nand NAND2 (N15439, N15435, N7900);
buf BUF1 (N15440, N15437);
not NOT1 (N15441, N15422);
nor NOR4 (N15442, N15427, N8047, N10669, N10912);
buf BUF1 (N15443, N15438);
xor XOR2 (N15444, N15436, N12379);
not NOT1 (N15445, N15426);
nor NOR3 (N15446, N15441, N14227, N1231);
or OR3 (N15447, N15444, N4406, N2059);
buf BUF1 (N15448, N15439);
xor XOR2 (N15449, N15446, N309);
nor NOR3 (N15450, N15448, N2501, N923);
buf BUF1 (N15451, N15440);
buf BUF1 (N15452, N15433);
xor XOR2 (N15453, N15451, N14491);
and AND4 (N15454, N15431, N11982, N2897, N7639);
not NOT1 (N15455, N15453);
nand NAND3 (N15456, N15449, N10882, N13311);
and AND4 (N15457, N15445, N5763, N6858, N130);
not NOT1 (N15458, N15434);
not NOT1 (N15459, N15458);
nand NAND2 (N15460, N15447, N1979);
nor NOR3 (N15461, N15443, N31, N9566);
nor NOR2 (N15462, N15460, N6297);
and AND2 (N15463, N15455, N7524);
xor XOR2 (N15464, N15462, N5450);
or OR2 (N15465, N15452, N11250);
nand NAND3 (N15466, N15442, N4983, N3328);
xor XOR2 (N15467, N15457, N11202);
or OR4 (N15468, N15464, N13337, N11000, N484);
and AND4 (N15469, N15468, N1088, N1682, N1407);
nor NOR2 (N15470, N15459, N4868);
and AND2 (N15471, N15456, N4545);
not NOT1 (N15472, N15471);
not NOT1 (N15473, N15454);
and AND3 (N15474, N15466, N8477, N3996);
xor XOR2 (N15475, N15470, N14519);
xor XOR2 (N15476, N15467, N13224);
and AND3 (N15477, N15476, N3222, N311);
nand NAND4 (N15478, N15473, N10482, N1598, N5618);
buf BUF1 (N15479, N15469);
nand NAND3 (N15480, N15461, N4723, N5778);
nor NOR4 (N15481, N15472, N13129, N8725, N7001);
or OR2 (N15482, N15479, N3593);
buf BUF1 (N15483, N15482);
nor NOR3 (N15484, N15480, N11159, N1924);
and AND3 (N15485, N15481, N6747, N1973);
nor NOR4 (N15486, N15465, N1787, N3583, N5433);
and AND3 (N15487, N15478, N2159, N1407);
or OR2 (N15488, N15475, N6767);
buf BUF1 (N15489, N15488);
not NOT1 (N15490, N15477);
nand NAND4 (N15491, N15484, N14652, N13776, N1263);
not NOT1 (N15492, N15483);
nand NAND3 (N15493, N15490, N1444, N10503);
nor NOR3 (N15494, N15489, N8562, N3728);
nand NAND3 (N15495, N15493, N6561, N6945);
or OR4 (N15496, N15491, N8446, N15402, N10524);
not NOT1 (N15497, N15485);
buf BUF1 (N15498, N15492);
buf BUF1 (N15499, N15495);
nand NAND4 (N15500, N15494, N13355, N438, N12010);
xor XOR2 (N15501, N15496, N5658);
and AND4 (N15502, N15487, N6354, N14492, N11838);
nor NOR4 (N15503, N15450, N5085, N10386, N608);
nand NAND3 (N15504, N15500, N8673, N3722);
not NOT1 (N15505, N15502);
nor NOR4 (N15506, N15486, N13038, N815, N7967);
nor NOR4 (N15507, N15501, N7530, N14878, N8006);
not NOT1 (N15508, N15507);
and AND3 (N15509, N15463, N5075, N3476);
nand NAND3 (N15510, N15497, N6572, N1069);
and AND4 (N15511, N15503, N3173, N10332, N768);
buf BUF1 (N15512, N15498);
nor NOR3 (N15513, N15510, N13728, N7532);
and AND4 (N15514, N15511, N547, N10616, N13537);
nor NOR3 (N15515, N15506, N12403, N14733);
nor NOR3 (N15516, N15512, N12723, N9738);
or OR3 (N15517, N15474, N10114, N10610);
nor NOR4 (N15518, N15515, N1137, N8301, N548);
buf BUF1 (N15519, N15509);
xor XOR2 (N15520, N15499, N1383);
buf BUF1 (N15521, N15517);
or OR4 (N15522, N15508, N8864, N102, N10028);
not NOT1 (N15523, N15518);
nand NAND4 (N15524, N15521, N14243, N1403, N13342);
buf BUF1 (N15525, N15519);
xor XOR2 (N15526, N15504, N2060);
xor XOR2 (N15527, N15516, N12225);
or OR4 (N15528, N15527, N8232, N11974, N7807);
and AND3 (N15529, N15522, N14832, N6493);
nand NAND3 (N15530, N15529, N10761, N2342);
or OR4 (N15531, N15525, N3658, N5407, N2817);
buf BUF1 (N15532, N15520);
xor XOR2 (N15533, N15528, N7066);
nand NAND4 (N15534, N15514, N4739, N10756, N10609);
buf BUF1 (N15535, N15533);
nand NAND4 (N15536, N15513, N9277, N5664, N1381);
or OR2 (N15537, N15531, N1649);
and AND2 (N15538, N15523, N4553);
not NOT1 (N15539, N15536);
buf BUF1 (N15540, N15537);
buf BUF1 (N15541, N15526);
or OR2 (N15542, N15524, N8914);
buf BUF1 (N15543, N15534);
buf BUF1 (N15544, N15538);
not NOT1 (N15545, N15505);
nand NAND2 (N15546, N15539, N13955);
buf BUF1 (N15547, N15530);
and AND3 (N15548, N15540, N7681, N6194);
not NOT1 (N15549, N15535);
nor NOR4 (N15550, N15542, N7014, N3340, N3197);
nor NOR2 (N15551, N15546, N13262);
nor NOR4 (N15552, N15544, N111, N11277, N1123);
and AND2 (N15553, N15545, N8004);
not NOT1 (N15554, N15547);
buf BUF1 (N15555, N15550);
or OR3 (N15556, N15551, N7613, N4456);
buf BUF1 (N15557, N15541);
or OR2 (N15558, N15557, N1211);
nand NAND2 (N15559, N15556, N899);
nor NOR3 (N15560, N15549, N3007, N1750);
or OR4 (N15561, N15548, N7776, N11098, N11700);
or OR4 (N15562, N15561, N14674, N1696, N4274);
xor XOR2 (N15563, N15555, N1494);
buf BUF1 (N15564, N15559);
nor NOR3 (N15565, N15532, N7380, N10238);
nor NOR4 (N15566, N15558, N4442, N9742, N10243);
xor XOR2 (N15567, N15554, N289);
and AND4 (N15568, N15563, N13136, N15168, N12775);
buf BUF1 (N15569, N15543);
buf BUF1 (N15570, N15562);
nand NAND3 (N15571, N15569, N12582, N12108);
not NOT1 (N15572, N15552);
xor XOR2 (N15573, N15572, N10269);
xor XOR2 (N15574, N15570, N5382);
and AND4 (N15575, N15571, N6591, N9892, N14022);
and AND2 (N15576, N15564, N8378);
nand NAND2 (N15577, N15568, N7153);
xor XOR2 (N15578, N15573, N3642);
nand NAND2 (N15579, N15553, N9789);
not NOT1 (N15580, N15575);
nor NOR4 (N15581, N15566, N1822, N1585, N12525);
or OR4 (N15582, N15565, N2596, N8773, N15291);
buf BUF1 (N15583, N15574);
nor NOR3 (N15584, N15577, N8232, N7075);
nor NOR2 (N15585, N15583, N7208);
or OR3 (N15586, N15581, N14092, N973);
xor XOR2 (N15587, N15584, N1920);
nor NOR4 (N15588, N15580, N11276, N14004, N3697);
xor XOR2 (N15589, N15588, N1713);
or OR4 (N15590, N15582, N14855, N5573, N14241);
xor XOR2 (N15591, N15576, N3900);
nor NOR4 (N15592, N15579, N195, N5382, N14386);
or OR4 (N15593, N15586, N11332, N13295, N10738);
and AND4 (N15594, N15587, N9360, N8921, N10997);
nand NAND2 (N15595, N15591, N12695);
or OR3 (N15596, N15589, N380, N2019);
nor NOR2 (N15597, N15578, N6100);
nand NAND3 (N15598, N15592, N1311, N11590);
and AND3 (N15599, N15594, N1891, N10991);
not NOT1 (N15600, N15590);
xor XOR2 (N15601, N15596, N14853);
nand NAND3 (N15602, N15601, N13230, N2316);
xor XOR2 (N15603, N15597, N13886);
or OR2 (N15604, N15595, N5362);
buf BUF1 (N15605, N15593);
nor NOR3 (N15606, N15598, N15433, N4285);
buf BUF1 (N15607, N15604);
nor NOR3 (N15608, N15600, N4890, N7387);
buf BUF1 (N15609, N15560);
xor XOR2 (N15610, N15608, N9446);
xor XOR2 (N15611, N15610, N3634);
buf BUF1 (N15612, N15611);
buf BUF1 (N15613, N15602);
or OR3 (N15614, N15612, N15192, N3273);
not NOT1 (N15615, N15599);
not NOT1 (N15616, N15603);
nand NAND2 (N15617, N15607, N5805);
nand NAND4 (N15618, N15614, N13767, N2198, N980);
not NOT1 (N15619, N15609);
nor NOR3 (N15620, N15618, N9282, N13746);
nor NOR3 (N15621, N15605, N4115, N12310);
not NOT1 (N15622, N15615);
not NOT1 (N15623, N15567);
xor XOR2 (N15624, N15617, N11560);
and AND2 (N15625, N15606, N5086);
and AND2 (N15626, N15622, N4065);
nand NAND2 (N15627, N15624, N5215);
not NOT1 (N15628, N15619);
buf BUF1 (N15629, N15628);
nor NOR3 (N15630, N15626, N7080, N9274);
not NOT1 (N15631, N15630);
nand NAND4 (N15632, N15616, N6901, N10460, N1142);
or OR4 (N15633, N15632, N7292, N2239, N5100);
buf BUF1 (N15634, N15627);
nand NAND3 (N15635, N15625, N12748, N13258);
or OR2 (N15636, N15635, N4590);
xor XOR2 (N15637, N15633, N4774);
nand NAND3 (N15638, N15621, N11416, N7786);
nand NAND4 (N15639, N15623, N2256, N5398, N15229);
xor XOR2 (N15640, N15636, N29);
buf BUF1 (N15641, N15638);
buf BUF1 (N15642, N15585);
not NOT1 (N15643, N15634);
and AND4 (N15644, N15639, N1028, N7012, N5724);
and AND4 (N15645, N15644, N5580, N12883, N8010);
not NOT1 (N15646, N15629);
and AND3 (N15647, N15640, N232, N2723);
or OR3 (N15648, N15643, N6824, N14925);
and AND3 (N15649, N15647, N1653, N343);
nor NOR4 (N15650, N15641, N12142, N1201, N14746);
not NOT1 (N15651, N15650);
and AND4 (N15652, N15631, N3500, N4018, N14989);
xor XOR2 (N15653, N15637, N4614);
nand NAND4 (N15654, N15620, N8920, N9084, N8505);
nand NAND2 (N15655, N15642, N6325);
and AND4 (N15656, N15648, N2217, N6987, N12234);
nor NOR4 (N15657, N15613, N6201, N8114, N6887);
nor NOR4 (N15658, N15646, N10251, N7392, N9143);
buf BUF1 (N15659, N15653);
and AND4 (N15660, N15651, N10536, N11324, N11968);
buf BUF1 (N15661, N15645);
buf BUF1 (N15662, N15661);
and AND3 (N15663, N15655, N10122, N1638);
buf BUF1 (N15664, N15656);
nor NOR4 (N15665, N15659, N19, N13784, N13299);
nand NAND4 (N15666, N15654, N6137, N5976, N14272);
xor XOR2 (N15667, N15662, N5873);
xor XOR2 (N15668, N15649, N11716);
nand NAND3 (N15669, N15664, N2060, N13016);
nor NOR4 (N15670, N15669, N1915, N7785, N9292);
nand NAND2 (N15671, N15668, N7290);
or OR2 (N15672, N15671, N8333);
or OR2 (N15673, N15665, N2064);
nand NAND3 (N15674, N15658, N1640, N3034);
or OR2 (N15675, N15672, N10309);
or OR2 (N15676, N15667, N4407);
nand NAND2 (N15677, N15657, N10413);
xor XOR2 (N15678, N15670, N14747);
or OR3 (N15679, N15660, N4983, N6508);
not NOT1 (N15680, N15663);
nor NOR2 (N15681, N15666, N11501);
xor XOR2 (N15682, N15680, N14513);
or OR4 (N15683, N15674, N3000, N4815, N7415);
not NOT1 (N15684, N15682);
nand NAND4 (N15685, N15652, N7290, N6413, N11060);
or OR3 (N15686, N15675, N11009, N1119);
not NOT1 (N15687, N15685);
xor XOR2 (N15688, N15683, N10658);
buf BUF1 (N15689, N15679);
nand NAND3 (N15690, N15678, N6365, N9902);
nand NAND3 (N15691, N15688, N7030, N9356);
nand NAND2 (N15692, N15676, N9849);
and AND4 (N15693, N15690, N10907, N9118, N9795);
xor XOR2 (N15694, N15684, N1788);
xor XOR2 (N15695, N15681, N13188);
nand NAND2 (N15696, N15689, N9194);
xor XOR2 (N15697, N15677, N2015);
not NOT1 (N15698, N15691);
xor XOR2 (N15699, N15697, N5019);
or OR2 (N15700, N15686, N8824);
nand NAND4 (N15701, N15694, N14478, N13900, N1362);
and AND3 (N15702, N15700, N13437, N11022);
nor NOR3 (N15703, N15698, N3920, N11650);
nor NOR2 (N15704, N15673, N11705);
nor NOR2 (N15705, N15693, N13866);
not NOT1 (N15706, N15703);
nor NOR2 (N15707, N15696, N1698);
buf BUF1 (N15708, N15707);
not NOT1 (N15709, N15705);
buf BUF1 (N15710, N15706);
buf BUF1 (N15711, N15704);
buf BUF1 (N15712, N15709);
nor NOR2 (N15713, N15687, N9678);
buf BUF1 (N15714, N15713);
xor XOR2 (N15715, N15712, N10799);
buf BUF1 (N15716, N15692);
and AND2 (N15717, N15716, N10933);
nand NAND4 (N15718, N15702, N3133, N12643, N540);
and AND2 (N15719, N15714, N14673);
buf BUF1 (N15720, N15710);
buf BUF1 (N15721, N15701);
and AND3 (N15722, N15699, N7514, N8025);
nor NOR3 (N15723, N15717, N4456, N10801);
buf BUF1 (N15724, N15718);
nand NAND4 (N15725, N15723, N5617, N3161, N5009);
or OR4 (N15726, N15724, N15354, N10444, N14951);
nor NOR3 (N15727, N15719, N10297, N2297);
or OR2 (N15728, N15715, N1607);
nor NOR2 (N15729, N15728, N6390);
buf BUF1 (N15730, N15727);
or OR3 (N15731, N15722, N12118, N986);
xor XOR2 (N15732, N15730, N5879);
xor XOR2 (N15733, N15732, N6814);
nor NOR4 (N15734, N15695, N195, N7260, N1966);
buf BUF1 (N15735, N15733);
nor NOR3 (N15736, N15720, N13749, N14486);
or OR3 (N15737, N15725, N2108, N5072);
nand NAND3 (N15738, N15726, N3871, N9784);
or OR2 (N15739, N15711, N9542);
not NOT1 (N15740, N15731);
not NOT1 (N15741, N15729);
nand NAND4 (N15742, N15740, N15440, N826, N12580);
nand NAND4 (N15743, N15721, N6653, N13667, N1607);
buf BUF1 (N15744, N15708);
buf BUF1 (N15745, N15735);
or OR2 (N15746, N15741, N12724);
and AND2 (N15747, N15737, N12610);
xor XOR2 (N15748, N15744, N9889);
and AND2 (N15749, N15742, N6751);
and AND2 (N15750, N15743, N1297);
buf BUF1 (N15751, N15748);
nand NAND2 (N15752, N15750, N15485);
nand NAND2 (N15753, N15752, N7947);
xor XOR2 (N15754, N15736, N14660);
or OR2 (N15755, N15753, N1098);
buf BUF1 (N15756, N15754);
buf BUF1 (N15757, N15746);
xor XOR2 (N15758, N15739, N2413);
nor NOR4 (N15759, N15758, N8255, N4886, N4233);
not NOT1 (N15760, N15749);
nand NAND4 (N15761, N15747, N8294, N13995, N13674);
and AND4 (N15762, N15757, N308, N10209, N9707);
or OR2 (N15763, N15734, N1990);
and AND4 (N15764, N15755, N10900, N11096, N13006);
nor NOR4 (N15765, N15751, N11889, N15251, N7818);
buf BUF1 (N15766, N15765);
or OR4 (N15767, N15762, N7169, N7697, N2103);
or OR2 (N15768, N15760, N10552);
not NOT1 (N15769, N15768);
xor XOR2 (N15770, N15761, N10138);
xor XOR2 (N15771, N15766, N12888);
nor NOR4 (N15772, N15756, N4347, N14789, N11799);
and AND3 (N15773, N15770, N5987, N7510);
nand NAND3 (N15774, N15745, N3635, N8137);
nand NAND3 (N15775, N15769, N10155, N9962);
nand NAND4 (N15776, N15774, N7204, N1169, N9960);
buf BUF1 (N15777, N15738);
nor NOR3 (N15778, N15759, N12265, N5970);
xor XOR2 (N15779, N15767, N3510);
and AND4 (N15780, N15771, N15139, N1871, N1453);
buf BUF1 (N15781, N15764);
buf BUF1 (N15782, N15778);
nor NOR2 (N15783, N15777, N8330);
xor XOR2 (N15784, N15783, N7590);
buf BUF1 (N15785, N15772);
and AND2 (N15786, N15780, N8989);
nand NAND4 (N15787, N15782, N2694, N14095, N6324);
nor NOR3 (N15788, N15781, N7352, N11419);
buf BUF1 (N15789, N15763);
buf BUF1 (N15790, N15787);
and AND4 (N15791, N15786, N14831, N10069, N5156);
xor XOR2 (N15792, N15788, N10354);
nand NAND3 (N15793, N15779, N6012, N4241);
xor XOR2 (N15794, N15790, N6737);
nand NAND4 (N15795, N15773, N5274, N4623, N723);
nand NAND2 (N15796, N15792, N3020);
xor XOR2 (N15797, N15793, N3568);
buf BUF1 (N15798, N15797);
nor NOR4 (N15799, N15796, N5828, N11102, N5420);
nor NOR4 (N15800, N15789, N6644, N10273, N9556);
nand NAND3 (N15801, N15798, N10478, N5164);
not NOT1 (N15802, N15801);
or OR2 (N15803, N15785, N2019);
nor NOR3 (N15804, N15799, N10311, N14310);
or OR2 (N15805, N15800, N1845);
xor XOR2 (N15806, N15795, N2557);
not NOT1 (N15807, N15805);
xor XOR2 (N15808, N15775, N9353);
and AND4 (N15809, N15776, N3198, N2682, N12283);
buf BUF1 (N15810, N15806);
xor XOR2 (N15811, N15808, N10201);
nor NOR3 (N15812, N15809, N13588, N10502);
nand NAND2 (N15813, N15791, N13565);
nor NOR2 (N15814, N15803, N4428);
xor XOR2 (N15815, N15812, N2262);
not NOT1 (N15816, N15807);
nand NAND2 (N15817, N15815, N12902);
not NOT1 (N15818, N15804);
or OR2 (N15819, N15784, N11127);
nand NAND3 (N15820, N15816, N4846, N6251);
or OR3 (N15821, N15811, N1228, N5423);
or OR4 (N15822, N15813, N5684, N70, N1696);
buf BUF1 (N15823, N15810);
and AND2 (N15824, N15821, N4575);
nor NOR2 (N15825, N15822, N3275);
not NOT1 (N15826, N15825);
and AND2 (N15827, N15814, N12488);
not NOT1 (N15828, N15794);
buf BUF1 (N15829, N15827);
nor NOR3 (N15830, N15823, N4049, N6770);
not NOT1 (N15831, N15829);
xor XOR2 (N15832, N15828, N14191);
not NOT1 (N15833, N15830);
buf BUF1 (N15834, N15818);
nor NOR4 (N15835, N15833, N3546, N11746, N1455);
nor NOR4 (N15836, N15826, N2798, N682, N14991);
not NOT1 (N15837, N15819);
or OR2 (N15838, N15817, N1438);
nand NAND4 (N15839, N15836, N11724, N2232, N6987);
not NOT1 (N15840, N15837);
nand NAND2 (N15841, N15802, N12867);
not NOT1 (N15842, N15835);
not NOT1 (N15843, N15831);
nand NAND2 (N15844, N15843, N14666);
nand NAND3 (N15845, N15841, N455, N240);
buf BUF1 (N15846, N15838);
buf BUF1 (N15847, N15844);
nand NAND4 (N15848, N15847, N96, N15232, N3831);
not NOT1 (N15849, N15846);
not NOT1 (N15850, N15820);
not NOT1 (N15851, N15849);
and AND3 (N15852, N15848, N14913, N7996);
nand NAND3 (N15853, N15839, N10898, N6868);
nand NAND2 (N15854, N15850, N12125);
xor XOR2 (N15855, N15832, N991);
not NOT1 (N15856, N15840);
or OR4 (N15857, N15834, N2830, N14818, N14240);
not NOT1 (N15858, N15857);
nor NOR3 (N15859, N15858, N8700, N14458);
buf BUF1 (N15860, N15853);
xor XOR2 (N15861, N15845, N14347);
not NOT1 (N15862, N15842);
nand NAND2 (N15863, N15851, N3065);
nor NOR4 (N15864, N15855, N12341, N5597, N2552);
and AND2 (N15865, N15824, N506);
xor XOR2 (N15866, N15861, N9986);
xor XOR2 (N15867, N15856, N6787);
and AND2 (N15868, N15859, N8673);
not NOT1 (N15869, N15863);
or OR2 (N15870, N15869, N9624);
nor NOR2 (N15871, N15867, N13142);
xor XOR2 (N15872, N15852, N13066);
nor NOR3 (N15873, N15865, N11843, N7369);
or OR4 (N15874, N15862, N12129, N647, N12122);
nand NAND2 (N15875, N15872, N5776);
nand NAND3 (N15876, N15864, N4460, N9215);
nor NOR3 (N15877, N15854, N1186, N8904);
not NOT1 (N15878, N15866);
buf BUF1 (N15879, N15877);
buf BUF1 (N15880, N15876);
not NOT1 (N15881, N15873);
and AND2 (N15882, N15875, N1618);
nand NAND2 (N15883, N15871, N3335);
buf BUF1 (N15884, N15881);
nor NOR4 (N15885, N15874, N11261, N12123, N10450);
nor NOR2 (N15886, N15868, N6947);
and AND3 (N15887, N15883, N2262, N7057);
and AND2 (N15888, N15860, N12730);
or OR4 (N15889, N15878, N1859, N2726, N14553);
xor XOR2 (N15890, N15879, N9758);
or OR4 (N15891, N15884, N1282, N9574, N9491);
nand NAND4 (N15892, N15880, N9844, N4334, N10590);
or OR2 (N15893, N15891, N15868);
not NOT1 (N15894, N15892);
buf BUF1 (N15895, N15887);
not NOT1 (N15896, N15886);
nand NAND2 (N15897, N15885, N6719);
or OR3 (N15898, N15888, N9975, N9733);
xor XOR2 (N15899, N15870, N7426);
or OR2 (N15900, N15899, N15150);
and AND4 (N15901, N15897, N7323, N6077, N11385);
or OR3 (N15902, N15894, N10448, N3942);
nand NAND3 (N15903, N15895, N13985, N3375);
buf BUF1 (N15904, N15893);
nor NOR2 (N15905, N15902, N5208);
not NOT1 (N15906, N15890);
nand NAND2 (N15907, N15903, N13750);
nor NOR2 (N15908, N15904, N9143);
not NOT1 (N15909, N15906);
buf BUF1 (N15910, N15889);
nor NOR4 (N15911, N15896, N4645, N13329, N6431);
not NOT1 (N15912, N15901);
and AND4 (N15913, N15882, N1834, N8294, N5085);
nand NAND3 (N15914, N15908, N8071, N9862);
xor XOR2 (N15915, N15909, N13277);
nor NOR3 (N15916, N15910, N15909, N3150);
and AND2 (N15917, N15916, N4005);
and AND4 (N15918, N15917, N12086, N7688, N14695);
xor XOR2 (N15919, N15915, N14017);
and AND4 (N15920, N15913, N407, N946, N12758);
or OR2 (N15921, N15920, N13559);
nor NOR4 (N15922, N15905, N7939, N13669, N1047);
and AND2 (N15923, N15918, N11413);
nor NOR2 (N15924, N15919, N14885);
nor NOR4 (N15925, N15922, N2987, N14947, N15229);
not NOT1 (N15926, N15924);
not NOT1 (N15927, N15914);
nand NAND4 (N15928, N15926, N2643, N5943, N12624);
nor NOR2 (N15929, N15928, N3462);
not NOT1 (N15930, N15923);
nor NOR2 (N15931, N15912, N1825);
and AND3 (N15932, N15900, N3238, N3265);
nand NAND3 (N15933, N15907, N4459, N14403);
buf BUF1 (N15934, N15921);
nand NAND2 (N15935, N15930, N15681);
not NOT1 (N15936, N15927);
nand NAND3 (N15937, N15925, N4149, N3918);
xor XOR2 (N15938, N15898, N6362);
or OR4 (N15939, N15911, N8501, N5848, N5533);
nand NAND2 (N15940, N15931, N7410);
or OR3 (N15941, N15938, N12745, N15744);
buf BUF1 (N15942, N15934);
nand NAND4 (N15943, N15939, N3145, N11024, N5843);
nor NOR2 (N15944, N15929, N9514);
nor NOR4 (N15945, N15941, N14341, N7290, N9576);
nand NAND3 (N15946, N15943, N7024, N5504);
xor XOR2 (N15947, N15937, N165);
xor XOR2 (N15948, N15932, N12595);
buf BUF1 (N15949, N15940);
buf BUF1 (N15950, N15948);
nand NAND2 (N15951, N15950, N11169);
buf BUF1 (N15952, N15933);
not NOT1 (N15953, N15947);
and AND4 (N15954, N15949, N12997, N4878, N14482);
not NOT1 (N15955, N15951);
buf BUF1 (N15956, N15954);
xor XOR2 (N15957, N15935, N2420);
nor NOR2 (N15958, N15953, N13230);
nor NOR4 (N15959, N15952, N9222, N2737, N8876);
buf BUF1 (N15960, N15942);
and AND3 (N15961, N15944, N13293, N3387);
or OR4 (N15962, N15958, N7225, N11016, N14842);
and AND4 (N15963, N15960, N8331, N6853, N12457);
or OR3 (N15964, N15955, N12050, N14862);
and AND4 (N15965, N15961, N5013, N1060, N12722);
not NOT1 (N15966, N15945);
not NOT1 (N15967, N15956);
nor NOR2 (N15968, N15963, N5070);
nand NAND4 (N15969, N15946, N7934, N11376, N7057);
not NOT1 (N15970, N15965);
nor NOR4 (N15971, N15968, N9196, N7224, N2239);
xor XOR2 (N15972, N15966, N12212);
nand NAND3 (N15973, N15964, N11203, N10708);
and AND4 (N15974, N15936, N5355, N5998, N13075);
nand NAND2 (N15975, N15962, N1371);
or OR2 (N15976, N15972, N348);
or OR4 (N15977, N15975, N7972, N5265, N890);
and AND3 (N15978, N15974, N3323, N2664);
buf BUF1 (N15979, N15971);
buf BUF1 (N15980, N15970);
buf BUF1 (N15981, N15959);
buf BUF1 (N15982, N15969);
not NOT1 (N15983, N15973);
and AND2 (N15984, N15977, N10914);
buf BUF1 (N15985, N15967);
buf BUF1 (N15986, N15978);
nor NOR4 (N15987, N15984, N14000, N5169, N4761);
nand NAND2 (N15988, N15981, N2792);
nor NOR3 (N15989, N15985, N12110, N15563);
and AND3 (N15990, N15986, N15665, N3546);
buf BUF1 (N15991, N15976);
buf BUF1 (N15992, N15982);
buf BUF1 (N15993, N15992);
buf BUF1 (N15994, N15983);
not NOT1 (N15995, N15979);
and AND4 (N15996, N15995, N2028, N13431, N5949);
nor NOR4 (N15997, N15994, N9912, N6419, N14235);
nand NAND2 (N15998, N15996, N4755);
buf BUF1 (N15999, N15987);
and AND2 (N16000, N15997, N5059);
and AND3 (N16001, N15980, N13380, N15598);
and AND3 (N16002, N15989, N7260, N11728);
buf BUF1 (N16003, N16002);
xor XOR2 (N16004, N16001, N11682);
not NOT1 (N16005, N16000);
not NOT1 (N16006, N15991);
and AND4 (N16007, N15957, N2866, N8550, N1537);
xor XOR2 (N16008, N16007, N10959);
buf BUF1 (N16009, N16004);
nor NOR2 (N16010, N15993, N7314);
nand NAND2 (N16011, N15988, N7379);
nor NOR3 (N16012, N15998, N9867, N13747);
not NOT1 (N16013, N16010);
xor XOR2 (N16014, N16013, N11380);
not NOT1 (N16015, N16014);
and AND2 (N16016, N16009, N3389);
nor NOR2 (N16017, N16011, N14022);
or OR2 (N16018, N16017, N10066);
nand NAND2 (N16019, N15990, N4458);
nor NOR3 (N16020, N15999, N12947, N8885);
and AND4 (N16021, N16016, N9866, N13293, N6944);
endmodule