// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16;

output N107,N94,N114,N109,N110,N100,N112,N115,N106,N116;

and AND4 (N17, N4, N14, N8, N9);
and AND2 (N18, N14, N4);
not NOT1 (N19, N10);
buf BUF1 (N20, N4);
and AND4 (N21, N5, N19, N6, N4);
nor NOR3 (N22, N2, N4, N5);
not NOT1 (N23, N19);
nor NOR2 (N24, N9, N18);
nor NOR2 (N25, N18, N4);
nor NOR2 (N26, N16, N2);
xor XOR2 (N27, N5, N15);
and AND3 (N28, N14, N9, N21);
nand NAND3 (N29, N24, N6, N1);
and AND4 (N30, N6, N27, N5, N6);
and AND2 (N31, N6, N6);
not NOT1 (N32, N29);
or OR4 (N33, N30, N9, N23, N9);
nand NAND2 (N34, N23, N13);
not NOT1 (N35, N25);
or OR4 (N36, N34, N23, N14, N32);
nand NAND4 (N37, N21, N31, N28, N33);
buf BUF1 (N38, N33);
nand NAND3 (N39, N36, N5, N31);
xor XOR2 (N40, N19, N35);
nor NOR3 (N41, N19, N5, N14);
nand NAND2 (N42, N41, N15);
not NOT1 (N43, N30);
or OR2 (N44, N26, N21);
and AND3 (N45, N39, N44, N22);
or OR3 (N46, N4, N23, N38);
nor NOR4 (N47, N1, N45, N34, N39);
or OR3 (N48, N36, N5, N45);
nor NOR3 (N49, N38, N40, N29);
nor NOR4 (N50, N37, N29, N25, N15);
buf BUF1 (N51, N26);
buf BUF1 (N52, N51);
nand NAND3 (N53, N47, N42, N8);
or OR3 (N54, N18, N36, N8);
nand NAND3 (N55, N53, N32, N50);
and AND3 (N56, N15, N32, N22);
and AND3 (N57, N54, N33, N40);
buf BUF1 (N58, N48);
nand NAND3 (N59, N52, N38, N38);
xor XOR2 (N60, N55, N10);
buf BUF1 (N61, N46);
and AND4 (N62, N20, N18, N47, N5);
xor XOR2 (N63, N62, N38);
or OR3 (N64, N43, N15, N51);
and AND2 (N65, N56, N7);
buf BUF1 (N66, N64);
or OR4 (N67, N57, N17, N14, N20);
not NOT1 (N68, N2);
nand NAND3 (N69, N68, N59, N40);
nand NAND3 (N70, N9, N20, N50);
nand NAND3 (N71, N65, N45, N12);
not NOT1 (N72, N67);
not NOT1 (N73, N71);
or OR3 (N74, N66, N59, N31);
nand NAND2 (N75, N49, N7);
nand NAND4 (N76, N63, N58, N49, N67);
not NOT1 (N77, N54);
nor NOR2 (N78, N72, N42);
xor XOR2 (N79, N75, N31);
not NOT1 (N80, N74);
not NOT1 (N81, N80);
not NOT1 (N82, N77);
buf BUF1 (N83, N69);
nor NOR3 (N84, N70, N55, N39);
or OR4 (N85, N61, N9, N6, N75);
nand NAND2 (N86, N85, N4);
buf BUF1 (N87, N60);
or OR3 (N88, N79, N70, N87);
not NOT1 (N89, N66);
and AND2 (N90, N81, N77);
not NOT1 (N91, N82);
buf BUF1 (N92, N84);
and AND3 (N93, N78, N56, N54);
not NOT1 (N94, N93);
not NOT1 (N95, N83);
nand NAND2 (N96, N88, N67);
or OR3 (N97, N91, N86, N36);
nand NAND3 (N98, N41, N92, N96);
or OR2 (N99, N45, N45);
nand NAND4 (N100, N46, N36, N79, N61);
or OR2 (N101, N97, N26);
xor XOR2 (N102, N95, N23);
buf BUF1 (N103, N102);
buf BUF1 (N104, N101);
xor XOR2 (N105, N76, N29);
not NOT1 (N106, N73);
and AND3 (N107, N90, N75, N53);
or OR4 (N108, N98, N84, N19, N79);
and AND2 (N109, N108, N97);
nor NOR2 (N110, N89, N25);
nor NOR3 (N111, N104, N75, N108);
or OR2 (N112, N105, N67);
nand NAND4 (N113, N99, N26, N34, N68);
buf BUF1 (N114, N103);
buf BUF1 (N115, N113);
and AND3 (N116, N111, N67, N10);
endmodule