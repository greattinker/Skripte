// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12;

output N2003,N2005,N1987,N2010,N2011,N2008,N2004,N2002,N1995,N2012;

xor XOR2 (N13, N8, N10);
nor NOR3 (N14, N7, N6, N13);
and AND4 (N15, N14, N4, N7, N3);
nand NAND3 (N16, N14, N8, N11);
nor NOR2 (N17, N14, N16);
nand NAND2 (N18, N11, N10);
or OR2 (N19, N8, N14);
not NOT1 (N20, N16);
buf BUF1 (N21, N11);
not NOT1 (N22, N7);
nand NAND2 (N23, N11, N12);
and AND3 (N24, N5, N10, N9);
or OR3 (N25, N21, N18, N15);
nand NAND3 (N26, N10, N9, N10);
not NOT1 (N27, N23);
nand NAND3 (N28, N16, N26, N17);
nor NOR4 (N29, N4, N3, N1, N12);
or OR4 (N30, N19, N27, N16, N22);
not NOT1 (N31, N15);
xor XOR2 (N32, N12, N1);
not NOT1 (N33, N30);
nand NAND4 (N34, N26, N15, N27, N20);
buf BUF1 (N35, N6);
nand NAND4 (N36, N6, N27, N3, N25);
not NOT1 (N37, N28);
nand NAND4 (N38, N15, N37, N26, N17);
or OR2 (N39, N29, N2);
and AND2 (N40, N12, N23);
xor XOR2 (N41, N31, N29);
not NOT1 (N42, N36);
or OR3 (N43, N42, N21, N24);
or OR3 (N44, N9, N35, N15);
or OR4 (N45, N12, N7, N22, N35);
buf BUF1 (N46, N40);
or OR4 (N47, N44, N8, N19, N41);
xor XOR2 (N48, N5, N9);
not NOT1 (N49, N48);
buf BUF1 (N50, N45);
and AND3 (N51, N50, N30, N19);
buf BUF1 (N52, N32);
and AND3 (N53, N43, N11, N51);
or OR3 (N54, N49, N26, N52);
nand NAND2 (N55, N41, N4);
nand NAND4 (N56, N18, N11, N19, N39);
and AND3 (N57, N16, N30, N44);
and AND4 (N58, N55, N56, N19, N17);
nor NOR4 (N59, N51, N15, N50, N48);
xor XOR2 (N60, N59, N44);
nor NOR3 (N61, N47, N37, N39);
or OR2 (N62, N53, N32);
nand NAND4 (N63, N62, N47, N21, N43);
xor XOR2 (N64, N63, N39);
nor NOR4 (N65, N58, N45, N54, N48);
not NOT1 (N66, N32);
not NOT1 (N67, N34);
not NOT1 (N68, N60);
not NOT1 (N69, N64);
xor XOR2 (N70, N61, N13);
xor XOR2 (N71, N57, N11);
or OR3 (N72, N67, N58, N50);
nand NAND3 (N73, N38, N26, N68);
nor NOR3 (N74, N25, N37, N38);
not NOT1 (N75, N74);
buf BUF1 (N76, N65);
and AND4 (N77, N73, N18, N21, N14);
not NOT1 (N78, N72);
nor NOR3 (N79, N33, N8, N33);
and AND4 (N80, N70, N77, N31, N64);
xor XOR2 (N81, N17, N30);
and AND3 (N82, N81, N42, N30);
and AND2 (N83, N46, N42);
or OR3 (N84, N79, N68, N63);
nand NAND2 (N85, N66, N37);
and AND4 (N86, N80, N25, N27, N20);
or OR2 (N87, N78, N85);
buf BUF1 (N88, N56);
or OR3 (N89, N76, N39, N24);
xor XOR2 (N90, N69, N82);
not NOT1 (N91, N51);
nor NOR4 (N92, N83, N34, N69, N51);
buf BUF1 (N93, N84);
nor NOR4 (N94, N71, N47, N83, N42);
not NOT1 (N95, N75);
nand NAND4 (N96, N91, N46, N65, N20);
not NOT1 (N97, N86);
or OR3 (N98, N93, N42, N49);
buf BUF1 (N99, N89);
nor NOR4 (N100, N95, N80, N99, N72);
buf BUF1 (N101, N71);
not NOT1 (N102, N92);
xor XOR2 (N103, N87, N88);
nor NOR2 (N104, N45, N7);
xor XOR2 (N105, N94, N66);
nand NAND4 (N106, N90, N6, N53, N54);
buf BUF1 (N107, N103);
nor NOR4 (N108, N102, N95, N89, N105);
and AND2 (N109, N57, N21);
buf BUF1 (N110, N96);
nand NAND4 (N111, N101, N34, N76, N6);
nand NAND2 (N112, N109, N97);
nand NAND3 (N113, N78, N4, N64);
or OR2 (N114, N100, N67);
and AND3 (N115, N106, N33, N13);
nor NOR2 (N116, N110, N33);
nand NAND3 (N117, N113, N20, N107);
or OR4 (N118, N98, N70, N28, N45);
xor XOR2 (N119, N44, N59);
or OR3 (N120, N115, N5, N6);
xor XOR2 (N121, N111, N96);
or OR4 (N122, N118, N70, N70, N117);
buf BUF1 (N123, N13);
and AND4 (N124, N108, N45, N45, N76);
not NOT1 (N125, N120);
xor XOR2 (N126, N112, N44);
nor NOR2 (N127, N104, N75);
and AND4 (N128, N126, N50, N105, N50);
nor NOR2 (N129, N114, N126);
nor NOR4 (N130, N119, N128, N22, N16);
nand NAND4 (N131, N30, N45, N122, N44);
or OR3 (N132, N63, N59, N76);
buf BUF1 (N133, N123);
not NOT1 (N134, N131);
and AND3 (N135, N121, N28, N37);
not NOT1 (N136, N130);
buf BUF1 (N137, N132);
nor NOR3 (N138, N125, N111, N27);
buf BUF1 (N139, N129);
xor XOR2 (N140, N133, N47);
not NOT1 (N141, N136);
nand NAND4 (N142, N141, N41, N88, N118);
not NOT1 (N143, N127);
xor XOR2 (N144, N124, N16);
xor XOR2 (N145, N139, N142);
nand NAND4 (N146, N89, N25, N56, N3);
and AND2 (N147, N137, N111);
and AND4 (N148, N116, N25, N100, N24);
or OR2 (N149, N144, N7);
not NOT1 (N150, N140);
and AND4 (N151, N149, N55, N15, N107);
and AND4 (N152, N138, N129, N100, N43);
and AND2 (N153, N135, N17);
buf BUF1 (N154, N134);
or OR3 (N155, N152, N101, N131);
xor XOR2 (N156, N143, N43);
or OR2 (N157, N150, N125);
and AND3 (N158, N145, N126, N35);
buf BUF1 (N159, N158);
xor XOR2 (N160, N159, N52);
and AND3 (N161, N156, N84, N48);
nor NOR4 (N162, N154, N42, N53, N18);
nand NAND2 (N163, N162, N117);
not NOT1 (N164, N160);
nor NOR2 (N165, N161, N94);
xor XOR2 (N166, N148, N79);
xor XOR2 (N167, N153, N68);
or OR4 (N168, N146, N92, N82, N139);
buf BUF1 (N169, N147);
xor XOR2 (N170, N165, N89);
and AND2 (N171, N167, N105);
buf BUF1 (N172, N163);
and AND3 (N173, N170, N93, N104);
not NOT1 (N174, N166);
nor NOR2 (N175, N169, N27);
or OR4 (N176, N164, N42, N77, N76);
nand NAND3 (N177, N168, N145, N26);
and AND3 (N178, N173, N146, N166);
or OR2 (N179, N175, N28);
not NOT1 (N180, N174);
nand NAND4 (N181, N179, N115, N9, N56);
nor NOR2 (N182, N181, N27);
nand NAND2 (N183, N176, N115);
buf BUF1 (N184, N178);
not NOT1 (N185, N184);
not NOT1 (N186, N183);
nand NAND4 (N187, N182, N125, N131, N63);
not NOT1 (N188, N186);
nand NAND2 (N189, N157, N72);
nand NAND3 (N190, N177, N77, N37);
nand NAND3 (N191, N185, N11, N9);
nand NAND4 (N192, N180, N121, N182, N180);
not NOT1 (N193, N192);
buf BUF1 (N194, N151);
or OR2 (N195, N187, N128);
nor NOR3 (N196, N195, N3, N27);
not NOT1 (N197, N193);
xor XOR2 (N198, N196, N106);
nand NAND4 (N199, N189, N169, N12, N69);
xor XOR2 (N200, N188, N107);
and AND2 (N201, N194, N177);
xor XOR2 (N202, N171, N61);
or OR4 (N203, N199, N85, N76, N149);
nand NAND2 (N204, N191, N121);
and AND3 (N205, N200, N200, N122);
buf BUF1 (N206, N197);
buf BUF1 (N207, N206);
nor NOR4 (N208, N205, N163, N55, N174);
buf BUF1 (N209, N208);
nor NOR2 (N210, N198, N150);
xor XOR2 (N211, N202, N59);
or OR2 (N212, N203, N11);
buf BUF1 (N213, N212);
or OR3 (N214, N213, N38, N176);
not NOT1 (N215, N155);
nand NAND4 (N216, N172, N129, N99, N76);
nand NAND4 (N217, N215, N48, N78, N123);
and AND2 (N218, N217, N42);
not NOT1 (N219, N218);
nand NAND2 (N220, N211, N141);
nor NOR2 (N221, N209, N52);
buf BUF1 (N222, N221);
nor NOR2 (N223, N216, N216);
xor XOR2 (N224, N222, N187);
and AND4 (N225, N210, N215, N47, N110);
buf BUF1 (N226, N214);
nor NOR2 (N227, N201, N219);
not NOT1 (N228, N103);
xor XOR2 (N229, N225, N166);
not NOT1 (N230, N227);
and AND3 (N231, N190, N97, N226);
nor NOR4 (N232, N3, N220, N46, N171);
nand NAND2 (N233, N130, N232);
nor NOR4 (N234, N47, N168, N144, N2);
nand NAND3 (N235, N231, N182, N213);
nand NAND4 (N236, N204, N20, N110, N88);
not NOT1 (N237, N223);
or OR3 (N238, N224, N135, N111);
nand NAND2 (N239, N233, N81);
or OR3 (N240, N228, N235, N20);
and AND4 (N241, N133, N217, N17, N96);
nand NAND4 (N242, N237, N166, N223, N17);
buf BUF1 (N243, N229);
or OR3 (N244, N238, N206, N135);
and AND4 (N245, N241, N209, N129, N95);
and AND4 (N246, N245, N191, N231, N76);
nand NAND2 (N247, N230, N61);
buf BUF1 (N248, N242);
or OR2 (N249, N240, N74);
nor NOR4 (N250, N236, N19, N56, N227);
buf BUF1 (N251, N207);
or OR3 (N252, N250, N4, N175);
and AND4 (N253, N252, N233, N147, N219);
not NOT1 (N254, N249);
xor XOR2 (N255, N253, N41);
nand NAND4 (N256, N244, N10, N224, N73);
nor NOR3 (N257, N243, N23, N108);
or OR4 (N258, N239, N129, N4, N17);
nor NOR3 (N259, N257, N78, N72);
not NOT1 (N260, N255);
nand NAND2 (N261, N254, N87);
or OR4 (N262, N246, N230, N7, N183);
xor XOR2 (N263, N234, N157);
and AND2 (N264, N248, N31);
and AND3 (N265, N261, N161, N64);
and AND2 (N266, N256, N5);
buf BUF1 (N267, N259);
buf BUF1 (N268, N264);
xor XOR2 (N269, N258, N200);
buf BUF1 (N270, N263);
and AND4 (N271, N247, N63, N89, N99);
or OR2 (N272, N262, N146);
xor XOR2 (N273, N251, N34);
nand NAND2 (N274, N260, N90);
buf BUF1 (N275, N272);
nand NAND2 (N276, N273, N211);
buf BUF1 (N277, N269);
or OR2 (N278, N266, N238);
buf BUF1 (N279, N275);
not NOT1 (N280, N265);
xor XOR2 (N281, N277, N204);
or OR4 (N282, N280, N98, N252, N136);
nor NOR4 (N283, N278, N48, N211, N84);
or OR2 (N284, N271, N270);
or OR3 (N285, N132, N262, N1);
buf BUF1 (N286, N267);
and AND2 (N287, N285, N103);
not NOT1 (N288, N282);
buf BUF1 (N289, N268);
not NOT1 (N290, N287);
and AND2 (N291, N289, N62);
xor XOR2 (N292, N279, N56);
nor NOR4 (N293, N290, N29, N63, N99);
buf BUF1 (N294, N286);
and AND2 (N295, N283, N135);
not NOT1 (N296, N293);
nor NOR2 (N297, N296, N67);
or OR4 (N298, N274, N45, N23, N114);
xor XOR2 (N299, N284, N269);
or OR2 (N300, N276, N181);
not NOT1 (N301, N288);
nand NAND4 (N302, N298, N260, N262, N225);
not NOT1 (N303, N281);
buf BUF1 (N304, N294);
nor NOR3 (N305, N301, N249, N95);
buf BUF1 (N306, N302);
nand NAND4 (N307, N305, N264, N148, N171);
buf BUF1 (N308, N303);
not NOT1 (N309, N308);
or OR4 (N310, N299, N130, N37, N128);
nor NOR3 (N311, N295, N174, N280);
nand NAND4 (N312, N307, N173, N147, N40);
nor NOR4 (N313, N309, N33, N308, N21);
not NOT1 (N314, N312);
not NOT1 (N315, N297);
not NOT1 (N316, N311);
and AND4 (N317, N315, N249, N137, N4);
nand NAND3 (N318, N306, N151, N297);
buf BUF1 (N319, N310);
buf BUF1 (N320, N300);
nor NOR3 (N321, N314, N150, N163);
and AND2 (N322, N291, N41);
buf BUF1 (N323, N318);
xor XOR2 (N324, N322, N47);
buf BUF1 (N325, N304);
buf BUF1 (N326, N325);
nor NOR4 (N327, N317, N159, N187, N7);
nor NOR2 (N328, N320, N285);
buf BUF1 (N329, N319);
buf BUF1 (N330, N326);
xor XOR2 (N331, N323, N54);
nor NOR3 (N332, N313, N320, N59);
nor NOR4 (N333, N324, N187, N13, N13);
or OR3 (N334, N321, N264, N128);
and AND3 (N335, N292, N59, N64);
or OR2 (N336, N329, N169);
or OR4 (N337, N333, N320, N218, N70);
nand NAND3 (N338, N332, N293, N293);
not NOT1 (N339, N330);
nor NOR3 (N340, N334, N44, N54);
not NOT1 (N341, N338);
nand NAND3 (N342, N316, N158, N323);
or OR2 (N343, N335, N191);
and AND3 (N344, N341, N139, N141);
or OR4 (N345, N327, N158, N59, N11);
not NOT1 (N346, N345);
xor XOR2 (N347, N331, N4);
not NOT1 (N348, N336);
xor XOR2 (N349, N343, N267);
buf BUF1 (N350, N339);
buf BUF1 (N351, N342);
or OR4 (N352, N346, N30, N90, N31);
buf BUF1 (N353, N340);
xor XOR2 (N354, N344, N180);
xor XOR2 (N355, N352, N290);
not NOT1 (N356, N348);
or OR3 (N357, N355, N297, N181);
or OR2 (N358, N356, N289);
not NOT1 (N359, N328);
buf BUF1 (N360, N353);
or OR4 (N361, N357, N175, N208, N11);
nor NOR4 (N362, N358, N201, N138, N120);
nor NOR3 (N363, N354, N9, N290);
buf BUF1 (N364, N363);
xor XOR2 (N365, N351, N113);
not NOT1 (N366, N337);
or OR2 (N367, N362, N79);
and AND2 (N368, N364, N63);
buf BUF1 (N369, N359);
or OR3 (N370, N368, N58, N342);
or OR2 (N371, N366, N218);
xor XOR2 (N372, N350, N33);
xor XOR2 (N373, N361, N116);
buf BUF1 (N374, N360);
and AND4 (N375, N372, N6, N128, N171);
or OR3 (N376, N369, N3, N362);
nor NOR2 (N377, N365, N51);
buf BUF1 (N378, N349);
buf BUF1 (N379, N376);
nor NOR2 (N380, N379, N336);
buf BUF1 (N381, N380);
xor XOR2 (N382, N374, N308);
xor XOR2 (N383, N375, N375);
not NOT1 (N384, N367);
and AND2 (N385, N377, N219);
nand NAND3 (N386, N378, N367, N102);
and AND4 (N387, N382, N228, N148, N20);
nand NAND4 (N388, N347, N381, N20, N96);
nand NAND2 (N389, N146, N291);
and AND2 (N390, N371, N344);
and AND3 (N391, N387, N44, N344);
buf BUF1 (N392, N385);
nor NOR4 (N393, N388, N321, N346, N68);
nand NAND3 (N394, N386, N87, N185);
nor NOR2 (N395, N390, N349);
nand NAND3 (N396, N384, N154, N349);
or OR3 (N397, N370, N139, N190);
or OR2 (N398, N389, N48);
nor NOR2 (N399, N396, N15);
nor NOR3 (N400, N398, N236, N141);
and AND4 (N401, N397, N359, N153, N307);
buf BUF1 (N402, N395);
and AND2 (N403, N399, N386);
or OR2 (N404, N393, N393);
xor XOR2 (N405, N400, N143);
nand NAND4 (N406, N392, N27, N289, N399);
nor NOR4 (N407, N383, N3, N237, N363);
nand NAND4 (N408, N394, N14, N234, N374);
nor NOR2 (N409, N407, N132);
nand NAND2 (N410, N404, N274);
or OR2 (N411, N410, N295);
and AND2 (N412, N409, N4);
or OR4 (N413, N408, N220, N393, N272);
nand NAND2 (N414, N406, N91);
xor XOR2 (N415, N412, N249);
xor XOR2 (N416, N405, N223);
buf BUF1 (N417, N416);
xor XOR2 (N418, N391, N283);
xor XOR2 (N419, N402, N24);
buf BUF1 (N420, N413);
or OR2 (N421, N418, N131);
buf BUF1 (N422, N417);
nor NOR2 (N423, N401, N378);
and AND4 (N424, N423, N99, N38, N189);
nand NAND3 (N425, N373, N245, N154);
nor NOR4 (N426, N419, N73, N66, N257);
nor NOR2 (N427, N420, N87);
not NOT1 (N428, N424);
or OR2 (N429, N428, N302);
not NOT1 (N430, N411);
buf BUF1 (N431, N422);
or OR2 (N432, N414, N47);
xor XOR2 (N433, N432, N26);
nand NAND2 (N434, N403, N29);
buf BUF1 (N435, N426);
xor XOR2 (N436, N429, N214);
not NOT1 (N437, N436);
buf BUF1 (N438, N431);
xor XOR2 (N439, N430, N198);
xor XOR2 (N440, N425, N360);
xor XOR2 (N441, N421, N230);
nor NOR2 (N442, N440, N18);
or OR2 (N443, N437, N13);
nor NOR2 (N444, N435, N287);
buf BUF1 (N445, N415);
nor NOR2 (N446, N445, N14);
nand NAND4 (N447, N444, N381, N403, N264);
not NOT1 (N448, N439);
nor NOR3 (N449, N447, N94, N176);
not NOT1 (N450, N427);
nor NOR3 (N451, N443, N431, N3);
nand NAND4 (N452, N451, N304, N284, N75);
nand NAND3 (N453, N442, N252, N86);
nand NAND2 (N454, N434, N220);
nor NOR2 (N455, N433, N181);
buf BUF1 (N456, N448);
buf BUF1 (N457, N449);
not NOT1 (N458, N457);
buf BUF1 (N459, N452);
or OR4 (N460, N446, N320, N228, N214);
nor NOR3 (N461, N460, N67, N163);
nand NAND3 (N462, N450, N379, N53);
xor XOR2 (N463, N455, N172);
not NOT1 (N464, N454);
xor XOR2 (N465, N463, N377);
nand NAND2 (N466, N441, N383);
not NOT1 (N467, N465);
and AND2 (N468, N456, N193);
or OR4 (N469, N467, N31, N269, N428);
not NOT1 (N470, N461);
nor NOR2 (N471, N464, N86);
or OR4 (N472, N468, N56, N176, N157);
xor XOR2 (N473, N458, N88);
nand NAND4 (N474, N466, N425, N470, N380);
xor XOR2 (N475, N443, N400);
xor XOR2 (N476, N459, N400);
nand NAND4 (N477, N462, N87, N436, N5);
buf BUF1 (N478, N474);
buf BUF1 (N479, N469);
buf BUF1 (N480, N476);
and AND3 (N481, N477, N240, N306);
not NOT1 (N482, N472);
xor XOR2 (N483, N471, N273);
and AND2 (N484, N473, N311);
or OR3 (N485, N479, N97, N160);
and AND2 (N486, N453, N78);
and AND3 (N487, N481, N467, N392);
nor NOR4 (N488, N482, N466, N29, N486);
xor XOR2 (N489, N201, N120);
and AND2 (N490, N480, N354);
xor XOR2 (N491, N438, N338);
xor XOR2 (N492, N478, N409);
nor NOR2 (N493, N475, N287);
and AND4 (N494, N487, N322, N352, N206);
nand NAND3 (N495, N483, N41, N403);
buf BUF1 (N496, N484);
xor XOR2 (N497, N491, N343);
or OR2 (N498, N489, N77);
nand NAND3 (N499, N485, N340, N171);
buf BUF1 (N500, N496);
xor XOR2 (N501, N499, N439);
and AND3 (N502, N494, N35, N3);
and AND3 (N503, N497, N222, N13);
and AND4 (N504, N493, N33, N264, N143);
and AND2 (N505, N498, N71);
nor NOR2 (N506, N505, N436);
not NOT1 (N507, N488);
nor NOR2 (N508, N504, N75);
nor NOR2 (N509, N501, N275);
or OR2 (N510, N490, N410);
nor NOR2 (N511, N503, N224);
not NOT1 (N512, N506);
nand NAND4 (N513, N510, N247, N127, N373);
xor XOR2 (N514, N507, N214);
nand NAND4 (N515, N512, N123, N321, N134);
and AND2 (N516, N515, N487);
nand NAND2 (N517, N514, N299);
or OR3 (N518, N500, N297, N380);
not NOT1 (N519, N495);
or OR3 (N520, N492, N517, N484);
nor NOR3 (N521, N63, N318, N438);
xor XOR2 (N522, N518, N168);
not NOT1 (N523, N522);
not NOT1 (N524, N520);
nor NOR2 (N525, N513, N121);
buf BUF1 (N526, N511);
and AND2 (N527, N525, N368);
buf BUF1 (N528, N523);
buf BUF1 (N529, N502);
not NOT1 (N530, N521);
buf BUF1 (N531, N529);
not NOT1 (N532, N527);
nor NOR4 (N533, N519, N336, N167, N152);
and AND3 (N534, N530, N298, N494);
not NOT1 (N535, N528);
or OR4 (N536, N534, N155, N510, N475);
buf BUF1 (N537, N509);
or OR3 (N538, N531, N432, N431);
buf BUF1 (N539, N532);
buf BUF1 (N540, N538);
not NOT1 (N541, N540);
nor NOR2 (N542, N536, N207);
or OR2 (N543, N537, N311);
nand NAND2 (N544, N508, N59);
xor XOR2 (N545, N533, N214);
nand NAND3 (N546, N526, N475, N124);
not NOT1 (N547, N539);
or OR3 (N548, N547, N47, N90);
and AND2 (N549, N535, N333);
nand NAND3 (N550, N524, N249, N513);
xor XOR2 (N551, N546, N260);
xor XOR2 (N552, N545, N159);
not NOT1 (N553, N551);
not NOT1 (N554, N544);
not NOT1 (N555, N548);
and AND4 (N556, N555, N138, N532, N287);
not NOT1 (N557, N554);
nand NAND3 (N558, N516, N502, N306);
or OR2 (N559, N552, N227);
nor NOR3 (N560, N550, N556, N283);
buf BUF1 (N561, N331);
not NOT1 (N562, N542);
not NOT1 (N563, N561);
nand NAND3 (N564, N549, N118, N386);
or OR3 (N565, N557, N404, N200);
and AND3 (N566, N562, N59, N141);
buf BUF1 (N567, N541);
nor NOR2 (N568, N560, N222);
or OR3 (N569, N558, N195, N528);
and AND4 (N570, N568, N78, N475, N174);
and AND2 (N571, N559, N172);
and AND3 (N572, N565, N165, N551);
not NOT1 (N573, N571);
nand NAND2 (N574, N553, N535);
xor XOR2 (N575, N563, N273);
nand NAND4 (N576, N569, N488, N255, N264);
and AND2 (N577, N564, N312);
nor NOR4 (N578, N572, N521, N405, N502);
and AND4 (N579, N543, N210, N38, N448);
not NOT1 (N580, N570);
buf BUF1 (N581, N580);
not NOT1 (N582, N581);
or OR4 (N583, N576, N493, N459, N550);
nor NOR3 (N584, N583, N130, N184);
nor NOR3 (N585, N577, N520, N453);
nand NAND4 (N586, N574, N476, N156, N212);
xor XOR2 (N587, N573, N480);
buf BUF1 (N588, N587);
buf BUF1 (N589, N584);
buf BUF1 (N590, N585);
xor XOR2 (N591, N586, N221);
nand NAND4 (N592, N588, N504, N278, N343);
or OR4 (N593, N578, N407, N66, N180);
nor NOR2 (N594, N589, N60);
or OR3 (N595, N575, N372, N473);
or OR2 (N596, N592, N238);
nand NAND4 (N597, N566, N286, N509, N564);
buf BUF1 (N598, N567);
nand NAND2 (N599, N598, N46);
nand NAND4 (N600, N596, N524, N166, N504);
buf BUF1 (N601, N600);
nor NOR3 (N602, N594, N599, N511);
or OR3 (N603, N64, N13, N431);
nand NAND2 (N604, N597, N476);
buf BUF1 (N605, N590);
or OR3 (N606, N601, N457, N173);
or OR3 (N607, N593, N33, N33);
xor XOR2 (N608, N602, N69);
not NOT1 (N609, N607);
or OR4 (N610, N591, N486, N429, N11);
not NOT1 (N611, N608);
not NOT1 (N612, N606);
nor NOR3 (N613, N610, N78, N377);
xor XOR2 (N614, N582, N218);
xor XOR2 (N615, N614, N263);
and AND3 (N616, N595, N213, N77);
buf BUF1 (N617, N615);
not NOT1 (N618, N617);
or OR3 (N619, N613, N450, N400);
xor XOR2 (N620, N609, N564);
not NOT1 (N621, N611);
not NOT1 (N622, N620);
or OR3 (N623, N579, N214, N257);
nor NOR2 (N624, N618, N348);
xor XOR2 (N625, N612, N87);
nand NAND3 (N626, N624, N83, N420);
or OR2 (N627, N603, N561);
not NOT1 (N628, N616);
nor NOR3 (N629, N621, N560, N144);
buf BUF1 (N630, N604);
not NOT1 (N631, N619);
not NOT1 (N632, N629);
and AND3 (N633, N632, N9, N163);
buf BUF1 (N634, N605);
and AND2 (N635, N622, N95);
or OR2 (N636, N623, N408);
buf BUF1 (N637, N636);
not NOT1 (N638, N625);
xor XOR2 (N639, N633, N246);
nor NOR4 (N640, N634, N225, N165, N291);
buf BUF1 (N641, N626);
nand NAND3 (N642, N630, N315, N8);
or OR2 (N643, N627, N603);
not NOT1 (N644, N637);
xor XOR2 (N645, N638, N395);
buf BUF1 (N646, N645);
nand NAND2 (N647, N628, N56);
and AND4 (N648, N639, N184, N342, N462);
or OR2 (N649, N642, N198);
nor NOR2 (N650, N649, N365);
not NOT1 (N651, N646);
and AND4 (N652, N640, N236, N611, N238);
nor NOR4 (N653, N643, N78, N573, N591);
not NOT1 (N654, N652);
not NOT1 (N655, N641);
not NOT1 (N656, N635);
nor NOR3 (N657, N654, N434, N606);
xor XOR2 (N658, N650, N164);
xor XOR2 (N659, N651, N648);
nor NOR2 (N660, N278, N176);
buf BUF1 (N661, N660);
buf BUF1 (N662, N647);
and AND2 (N663, N659, N88);
nand NAND4 (N664, N644, N439, N435, N118);
nand NAND4 (N665, N657, N250, N618, N517);
or OR4 (N666, N656, N259, N220, N117);
xor XOR2 (N667, N665, N628);
buf BUF1 (N668, N666);
nand NAND2 (N669, N655, N370);
nor NOR3 (N670, N669, N296, N83);
and AND2 (N671, N663, N587);
not NOT1 (N672, N662);
nand NAND4 (N673, N668, N337, N213, N157);
xor XOR2 (N674, N672, N61);
not NOT1 (N675, N631);
xor XOR2 (N676, N675, N492);
nand NAND3 (N677, N661, N196, N382);
and AND3 (N678, N676, N492, N488);
or OR4 (N679, N664, N417, N614, N31);
nand NAND2 (N680, N673, N309);
not NOT1 (N681, N680);
nand NAND2 (N682, N674, N98);
not NOT1 (N683, N677);
nand NAND2 (N684, N658, N202);
nor NOR2 (N685, N684, N466);
nand NAND4 (N686, N670, N320, N240, N244);
and AND3 (N687, N686, N499, N378);
buf BUF1 (N688, N685);
buf BUF1 (N689, N679);
and AND4 (N690, N688, N589, N224, N588);
and AND3 (N691, N671, N206, N377);
nand NAND4 (N692, N687, N430, N537, N111);
or OR4 (N693, N689, N382, N226, N171);
nor NOR3 (N694, N682, N640, N563);
buf BUF1 (N695, N667);
and AND2 (N696, N678, N655);
buf BUF1 (N697, N653);
and AND4 (N698, N696, N409, N181, N55);
and AND2 (N699, N693, N125);
not NOT1 (N700, N681);
and AND2 (N701, N698, N114);
buf BUF1 (N702, N700);
and AND3 (N703, N694, N690, N306);
nand NAND2 (N704, N642, N238);
or OR2 (N705, N703, N464);
not NOT1 (N706, N697);
nor NOR2 (N707, N692, N655);
not NOT1 (N708, N704);
buf BUF1 (N709, N699);
and AND2 (N710, N706, N25);
not NOT1 (N711, N705);
xor XOR2 (N712, N691, N698);
xor XOR2 (N713, N707, N406);
buf BUF1 (N714, N713);
nand NAND4 (N715, N714, N78, N208, N58);
not NOT1 (N716, N708);
and AND2 (N717, N709, N166);
or OR3 (N718, N717, N451, N673);
or OR4 (N719, N710, N356, N536, N146);
or OR4 (N720, N711, N310, N63, N251);
or OR4 (N721, N715, N127, N156, N397);
and AND3 (N722, N716, N60, N285);
nor NOR4 (N723, N695, N224, N469, N604);
nand NAND4 (N724, N721, N486, N644, N612);
or OR2 (N725, N702, N89);
xor XOR2 (N726, N683, N695);
buf BUF1 (N727, N720);
and AND2 (N728, N726, N196);
or OR2 (N729, N712, N417);
nand NAND4 (N730, N718, N693, N420, N122);
nand NAND4 (N731, N701, N506, N430, N634);
and AND2 (N732, N719, N185);
not NOT1 (N733, N723);
xor XOR2 (N734, N727, N203);
nor NOR2 (N735, N730, N37);
xor XOR2 (N736, N731, N623);
nand NAND3 (N737, N724, N428, N660);
not NOT1 (N738, N729);
and AND4 (N739, N734, N327, N439, N240);
buf BUF1 (N740, N739);
or OR3 (N741, N736, N587, N328);
nor NOR3 (N742, N737, N213, N406);
nor NOR4 (N743, N722, N60, N686, N188);
nor NOR4 (N744, N740, N273, N732, N197);
xor XOR2 (N745, N177, N265);
and AND3 (N746, N744, N132, N673);
nand NAND3 (N747, N735, N49, N63);
and AND2 (N748, N741, N418);
or OR4 (N749, N742, N742, N78, N373);
nor NOR4 (N750, N745, N115, N506, N617);
nor NOR4 (N751, N750, N117, N668, N114);
not NOT1 (N752, N746);
buf BUF1 (N753, N752);
xor XOR2 (N754, N733, N525);
buf BUF1 (N755, N749);
or OR3 (N756, N747, N183, N426);
nand NAND4 (N757, N753, N338, N430, N17);
not NOT1 (N758, N755);
or OR3 (N759, N728, N78, N241);
or OR4 (N760, N743, N31, N407, N113);
not NOT1 (N761, N756);
not NOT1 (N762, N751);
nor NOR3 (N763, N748, N2, N534);
nand NAND4 (N764, N757, N34, N287, N642);
nand NAND4 (N765, N761, N542, N47, N173);
buf BUF1 (N766, N759);
or OR4 (N767, N765, N673, N559, N86);
nand NAND3 (N768, N762, N657, N304);
buf BUF1 (N769, N768);
buf BUF1 (N770, N769);
xor XOR2 (N771, N770, N604);
and AND4 (N772, N767, N248, N250, N553);
nor NOR3 (N773, N758, N435, N572);
or OR2 (N774, N738, N537);
and AND4 (N775, N764, N534, N66, N473);
and AND3 (N776, N772, N567, N445);
buf BUF1 (N777, N766);
not NOT1 (N778, N776);
buf BUF1 (N779, N754);
and AND4 (N780, N779, N713, N647, N351);
nand NAND2 (N781, N763, N332);
nor NOR4 (N782, N771, N397, N611, N113);
nand NAND2 (N783, N778, N103);
not NOT1 (N784, N780);
nand NAND3 (N785, N725, N580, N596);
nor NOR4 (N786, N783, N413, N201, N121);
xor XOR2 (N787, N786, N773);
or OR2 (N788, N382, N233);
nand NAND4 (N789, N785, N431, N783, N652);
or OR3 (N790, N784, N237, N735);
xor XOR2 (N791, N787, N746);
nor NOR3 (N792, N789, N497, N153);
xor XOR2 (N793, N781, N733);
buf BUF1 (N794, N782);
and AND2 (N795, N793, N595);
or OR4 (N796, N792, N368, N548, N343);
and AND4 (N797, N788, N776, N700, N638);
or OR4 (N798, N796, N329, N241, N367);
nor NOR2 (N799, N797, N779);
and AND4 (N800, N774, N251, N469, N60);
buf BUF1 (N801, N760);
and AND3 (N802, N801, N9, N72);
nand NAND4 (N803, N798, N362, N689, N194);
not NOT1 (N804, N800);
nand NAND4 (N805, N802, N81, N169, N306);
xor XOR2 (N806, N790, N534);
or OR2 (N807, N794, N682);
nand NAND3 (N808, N806, N803, N364);
not NOT1 (N809, N751);
nand NAND2 (N810, N807, N471);
xor XOR2 (N811, N777, N665);
nor NOR4 (N812, N811, N155, N368, N23);
buf BUF1 (N813, N799);
buf BUF1 (N814, N791);
and AND2 (N815, N813, N254);
xor XOR2 (N816, N815, N313);
xor XOR2 (N817, N804, N366);
buf BUF1 (N818, N795);
nand NAND3 (N819, N818, N585, N222);
xor XOR2 (N820, N808, N733);
and AND4 (N821, N809, N427, N30, N484);
or OR3 (N822, N817, N572, N466);
nor NOR4 (N823, N775, N800, N308, N221);
nand NAND3 (N824, N823, N313, N436);
or OR4 (N825, N819, N449, N196, N39);
xor XOR2 (N826, N816, N91);
and AND3 (N827, N814, N201, N709);
buf BUF1 (N828, N825);
xor XOR2 (N829, N805, N777);
or OR2 (N830, N828, N497);
buf BUF1 (N831, N812);
not NOT1 (N832, N821);
or OR4 (N833, N820, N261, N68, N771);
not NOT1 (N834, N831);
xor XOR2 (N835, N834, N505);
not NOT1 (N836, N824);
or OR3 (N837, N836, N740, N168);
not NOT1 (N838, N830);
nor NOR3 (N839, N838, N332, N646);
not NOT1 (N840, N837);
buf BUF1 (N841, N810);
buf BUF1 (N842, N829);
nor NOR4 (N843, N827, N328, N529, N109);
nor NOR2 (N844, N832, N106);
not NOT1 (N845, N842);
xor XOR2 (N846, N826, N746);
buf BUF1 (N847, N835);
xor XOR2 (N848, N840, N555);
buf BUF1 (N849, N847);
and AND2 (N850, N844, N846);
xor XOR2 (N851, N670, N114);
nor NOR2 (N852, N849, N641);
buf BUF1 (N853, N843);
or OR3 (N854, N850, N440, N24);
nand NAND2 (N855, N839, N66);
and AND3 (N856, N853, N105, N274);
nor NOR4 (N857, N822, N276, N266, N527);
not NOT1 (N858, N841);
not NOT1 (N859, N833);
or OR4 (N860, N854, N818, N635, N429);
not NOT1 (N861, N857);
and AND2 (N862, N845, N615);
nand NAND3 (N863, N860, N528, N731);
buf BUF1 (N864, N852);
buf BUF1 (N865, N859);
buf BUF1 (N866, N861);
and AND2 (N867, N851, N641);
xor XOR2 (N868, N855, N432);
not NOT1 (N869, N856);
or OR3 (N870, N867, N376, N280);
and AND2 (N871, N868, N115);
nand NAND2 (N872, N862, N150);
buf BUF1 (N873, N872);
not NOT1 (N874, N848);
and AND3 (N875, N873, N644, N302);
nor NOR3 (N876, N865, N402, N852);
nor NOR3 (N877, N871, N763, N805);
nand NAND4 (N878, N864, N115, N617, N95);
or OR4 (N879, N878, N155, N215, N682);
or OR2 (N880, N877, N102);
xor XOR2 (N881, N866, N291);
buf BUF1 (N882, N879);
not NOT1 (N883, N880);
nand NAND4 (N884, N875, N117, N6, N401);
or OR2 (N885, N884, N221);
not NOT1 (N886, N876);
xor XOR2 (N887, N863, N564);
not NOT1 (N888, N870);
nand NAND3 (N889, N887, N299, N739);
buf BUF1 (N890, N881);
not NOT1 (N891, N886);
nor NOR2 (N892, N883, N610);
and AND4 (N893, N858, N592, N744, N590);
not NOT1 (N894, N888);
or OR3 (N895, N869, N389, N310);
nand NAND4 (N896, N874, N561, N600, N287);
not NOT1 (N897, N896);
xor XOR2 (N898, N882, N167);
not NOT1 (N899, N885);
and AND2 (N900, N898, N365);
not NOT1 (N901, N895);
nor NOR2 (N902, N892, N419);
or OR4 (N903, N902, N846, N28, N61);
xor XOR2 (N904, N889, N831);
not NOT1 (N905, N890);
not NOT1 (N906, N897);
not NOT1 (N907, N903);
xor XOR2 (N908, N906, N253);
and AND4 (N909, N899, N181, N751, N585);
and AND3 (N910, N901, N815, N732);
xor XOR2 (N911, N908, N130);
buf BUF1 (N912, N900);
nor NOR4 (N913, N910, N170, N545, N12);
or OR4 (N914, N909, N655, N787, N8);
buf BUF1 (N915, N914);
nand NAND4 (N916, N911, N94, N82, N167);
xor XOR2 (N917, N915, N70);
xor XOR2 (N918, N905, N357);
nand NAND4 (N919, N917, N415, N118, N81);
and AND2 (N920, N912, N32);
and AND2 (N921, N904, N396);
not NOT1 (N922, N891);
not NOT1 (N923, N918);
or OR4 (N924, N907, N47, N860, N315);
buf BUF1 (N925, N913);
buf BUF1 (N926, N924);
or OR4 (N927, N923, N696, N765, N691);
or OR3 (N928, N920, N847, N683);
buf BUF1 (N929, N928);
xor XOR2 (N930, N922, N139);
not NOT1 (N931, N916);
nor NOR2 (N932, N931, N300);
and AND4 (N933, N927, N364, N913, N743);
nand NAND4 (N934, N933, N365, N356, N448);
or OR4 (N935, N894, N548, N3, N482);
not NOT1 (N936, N926);
nor NOR2 (N937, N935, N788);
xor XOR2 (N938, N932, N92);
and AND4 (N939, N929, N453, N524, N184);
xor XOR2 (N940, N936, N551);
buf BUF1 (N941, N938);
nor NOR3 (N942, N937, N894, N325);
nor NOR4 (N943, N941, N172, N769, N899);
or OR3 (N944, N940, N551, N741);
buf BUF1 (N945, N921);
not NOT1 (N946, N934);
and AND3 (N947, N945, N659, N912);
nor NOR4 (N948, N919, N343, N78, N62);
or OR4 (N949, N947, N269, N600, N814);
buf BUF1 (N950, N946);
nor NOR3 (N951, N948, N614, N256);
nor NOR4 (N952, N942, N580, N239, N269);
buf BUF1 (N953, N925);
nor NOR3 (N954, N949, N487, N458);
not NOT1 (N955, N939);
not NOT1 (N956, N953);
or OR2 (N957, N954, N575);
xor XOR2 (N958, N951, N459);
xor XOR2 (N959, N950, N154);
not NOT1 (N960, N955);
and AND4 (N961, N943, N562, N861, N472);
nand NAND4 (N962, N957, N173, N294, N218);
xor XOR2 (N963, N930, N585);
xor XOR2 (N964, N961, N152);
and AND2 (N965, N956, N164);
nor NOR2 (N966, N952, N289);
nand NAND3 (N967, N960, N941, N685);
xor XOR2 (N968, N966, N408);
xor XOR2 (N969, N963, N725);
nor NOR2 (N970, N893, N225);
not NOT1 (N971, N944);
or OR2 (N972, N969, N258);
buf BUF1 (N973, N958);
buf BUF1 (N974, N964);
nor NOR3 (N975, N971, N48, N119);
nand NAND4 (N976, N968, N137, N229, N212);
nor NOR3 (N977, N962, N948, N260);
buf BUF1 (N978, N959);
or OR2 (N979, N976, N535);
and AND4 (N980, N978, N848, N547, N331);
or OR3 (N981, N975, N203, N747);
nand NAND3 (N982, N979, N52, N126);
not NOT1 (N983, N980);
not NOT1 (N984, N973);
buf BUF1 (N985, N983);
and AND2 (N986, N985, N232);
or OR4 (N987, N970, N80, N3, N370);
nand NAND2 (N988, N984, N900);
nor NOR3 (N989, N974, N755, N65);
and AND2 (N990, N988, N907);
or OR4 (N991, N965, N529, N148, N325);
buf BUF1 (N992, N972);
or OR3 (N993, N981, N630, N177);
and AND2 (N994, N991, N628);
buf BUF1 (N995, N967);
nand NAND3 (N996, N992, N488, N455);
xor XOR2 (N997, N993, N738);
buf BUF1 (N998, N994);
or OR3 (N999, N998, N710, N787);
nor NOR4 (N1000, N997, N937, N318, N751);
nand NAND3 (N1001, N989, N971, N31);
and AND3 (N1002, N990, N259, N73);
nand NAND2 (N1003, N1002, N44);
and AND2 (N1004, N1003, N960);
and AND3 (N1005, N1004, N795, N273);
nand NAND2 (N1006, N995, N193);
not NOT1 (N1007, N1001);
buf BUF1 (N1008, N999);
and AND2 (N1009, N987, N58);
not NOT1 (N1010, N1008);
nand NAND4 (N1011, N1009, N901, N724, N85);
buf BUF1 (N1012, N986);
xor XOR2 (N1013, N1005, N525);
nand NAND4 (N1014, N1010, N687, N249, N224);
nand NAND3 (N1015, N1011, N83, N953);
nand NAND2 (N1016, N977, N844);
nor NOR3 (N1017, N982, N350, N955);
or OR2 (N1018, N1006, N843);
nor NOR2 (N1019, N1018, N652);
or OR2 (N1020, N1014, N899);
xor XOR2 (N1021, N1015, N833);
and AND4 (N1022, N1012, N33, N417, N8);
nand NAND4 (N1023, N1013, N524, N783, N82);
and AND4 (N1024, N1023, N98, N957, N760);
nor NOR3 (N1025, N1007, N601, N251);
not NOT1 (N1026, N1021);
nand NAND2 (N1027, N1016, N968);
not NOT1 (N1028, N1019);
nor NOR2 (N1029, N1028, N855);
nand NAND4 (N1030, N1000, N527, N774, N34);
and AND2 (N1031, N1030, N966);
buf BUF1 (N1032, N1029);
or OR3 (N1033, N1027, N976, N569);
nand NAND3 (N1034, N1033, N569, N59);
or OR3 (N1035, N1017, N263, N730);
or OR4 (N1036, N1032, N905, N399, N320);
not NOT1 (N1037, N1036);
not NOT1 (N1038, N1022);
nor NOR2 (N1039, N1037, N316);
and AND4 (N1040, N996, N391, N630, N879);
xor XOR2 (N1041, N1035, N135);
xor XOR2 (N1042, N1038, N718);
nor NOR3 (N1043, N1034, N500, N263);
xor XOR2 (N1044, N1042, N590);
buf BUF1 (N1045, N1020);
buf BUF1 (N1046, N1045);
and AND2 (N1047, N1044, N116);
and AND3 (N1048, N1024, N724, N706);
not NOT1 (N1049, N1026);
nor NOR2 (N1050, N1049, N104);
not NOT1 (N1051, N1039);
nand NAND4 (N1052, N1051, N199, N859, N325);
or OR4 (N1053, N1040, N565, N1014, N947);
and AND3 (N1054, N1025, N667, N279);
xor XOR2 (N1055, N1050, N890);
or OR2 (N1056, N1031, N294);
or OR2 (N1057, N1055, N616);
nor NOR4 (N1058, N1054, N210, N204, N629);
not NOT1 (N1059, N1057);
nand NAND3 (N1060, N1046, N222, N774);
buf BUF1 (N1061, N1052);
buf BUF1 (N1062, N1048);
or OR3 (N1063, N1047, N420, N627);
or OR4 (N1064, N1041, N137, N809, N533);
nor NOR2 (N1065, N1062, N54);
or OR2 (N1066, N1064, N71);
not NOT1 (N1067, N1066);
and AND3 (N1068, N1058, N855, N540);
nand NAND2 (N1069, N1059, N94);
and AND4 (N1070, N1061, N274, N67, N688);
and AND3 (N1071, N1043, N634, N61);
and AND2 (N1072, N1060, N9);
and AND3 (N1073, N1056, N695, N684);
nand NAND3 (N1074, N1070, N291, N59);
buf BUF1 (N1075, N1065);
or OR3 (N1076, N1053, N770, N703);
not NOT1 (N1077, N1069);
and AND3 (N1078, N1068, N255, N605);
nor NOR3 (N1079, N1078, N552, N17);
not NOT1 (N1080, N1076);
or OR4 (N1081, N1079, N814, N283, N248);
xor XOR2 (N1082, N1067, N172);
buf BUF1 (N1083, N1080);
or OR4 (N1084, N1083, N896, N261, N985);
xor XOR2 (N1085, N1084, N489);
xor XOR2 (N1086, N1071, N398);
nand NAND2 (N1087, N1074, N59);
and AND3 (N1088, N1073, N315, N141);
and AND3 (N1089, N1086, N807, N28);
xor XOR2 (N1090, N1089, N303);
and AND3 (N1091, N1072, N898, N589);
nand NAND2 (N1092, N1087, N740);
or OR3 (N1093, N1081, N648, N689);
xor XOR2 (N1094, N1093, N790);
nor NOR3 (N1095, N1082, N1081, N187);
xor XOR2 (N1096, N1088, N415);
nor NOR2 (N1097, N1094, N515);
and AND3 (N1098, N1091, N934, N542);
nand NAND2 (N1099, N1075, N41);
or OR4 (N1100, N1063, N109, N626, N169);
not NOT1 (N1101, N1095);
buf BUF1 (N1102, N1092);
nand NAND3 (N1103, N1098, N18, N874);
buf BUF1 (N1104, N1101);
not NOT1 (N1105, N1104);
buf BUF1 (N1106, N1097);
and AND2 (N1107, N1077, N328);
nand NAND4 (N1108, N1105, N794, N162, N490);
nor NOR3 (N1109, N1096, N647, N573);
not NOT1 (N1110, N1090);
nor NOR4 (N1111, N1108, N704, N635, N496);
nand NAND2 (N1112, N1102, N816);
not NOT1 (N1113, N1109);
or OR2 (N1114, N1100, N1100);
nand NAND4 (N1115, N1110, N122, N1087, N499);
xor XOR2 (N1116, N1106, N888);
buf BUF1 (N1117, N1107);
or OR2 (N1118, N1115, N785);
nand NAND2 (N1119, N1085, N71);
nand NAND4 (N1120, N1119, N70, N287, N513);
and AND3 (N1121, N1118, N379, N122);
nor NOR2 (N1122, N1114, N645);
buf BUF1 (N1123, N1111);
xor XOR2 (N1124, N1116, N888);
or OR3 (N1125, N1123, N270, N875);
nor NOR4 (N1126, N1122, N368, N290, N410);
xor XOR2 (N1127, N1112, N265);
and AND2 (N1128, N1126, N223);
and AND2 (N1129, N1113, N590);
not NOT1 (N1130, N1099);
nor NOR2 (N1131, N1103, N255);
nor NOR3 (N1132, N1130, N911, N1111);
nor NOR2 (N1133, N1121, N573);
nand NAND2 (N1134, N1132, N306);
or OR3 (N1135, N1127, N841, N1039);
nor NOR2 (N1136, N1120, N247);
nor NOR2 (N1137, N1129, N696);
buf BUF1 (N1138, N1133);
buf BUF1 (N1139, N1131);
not NOT1 (N1140, N1134);
and AND2 (N1141, N1125, N313);
nand NAND3 (N1142, N1141, N226, N710);
and AND3 (N1143, N1142, N404, N114);
or OR4 (N1144, N1137, N286, N234, N398);
nand NAND2 (N1145, N1135, N892);
nor NOR3 (N1146, N1144, N78, N610);
buf BUF1 (N1147, N1138);
or OR3 (N1148, N1117, N15, N375);
nand NAND4 (N1149, N1148, N512, N706, N335);
and AND3 (N1150, N1147, N667, N931);
not NOT1 (N1151, N1124);
not NOT1 (N1152, N1139);
buf BUF1 (N1153, N1136);
nand NAND3 (N1154, N1146, N943, N671);
nor NOR4 (N1155, N1151, N262, N762, N532);
nor NOR3 (N1156, N1143, N475, N116);
nand NAND4 (N1157, N1145, N243, N691, N43);
not NOT1 (N1158, N1154);
nor NOR4 (N1159, N1152, N910, N191, N356);
nand NAND3 (N1160, N1149, N954, N817);
nand NAND4 (N1161, N1153, N612, N415, N670);
nor NOR3 (N1162, N1128, N1077, N192);
xor XOR2 (N1163, N1155, N104);
nor NOR2 (N1164, N1161, N1107);
xor XOR2 (N1165, N1158, N1098);
buf BUF1 (N1166, N1162);
nand NAND2 (N1167, N1166, N238);
not NOT1 (N1168, N1164);
or OR4 (N1169, N1163, N688, N1120, N556);
not NOT1 (N1170, N1169);
nand NAND3 (N1171, N1150, N852, N1129);
not NOT1 (N1172, N1170);
and AND2 (N1173, N1171, N4);
nand NAND2 (N1174, N1160, N361);
nor NOR3 (N1175, N1159, N340, N1102);
not NOT1 (N1176, N1140);
or OR2 (N1177, N1172, N589);
or OR2 (N1178, N1177, N229);
nor NOR2 (N1179, N1167, N13);
not NOT1 (N1180, N1174);
buf BUF1 (N1181, N1175);
nor NOR2 (N1182, N1179, N290);
nor NOR3 (N1183, N1156, N686, N718);
nor NOR3 (N1184, N1178, N930, N43);
or OR4 (N1185, N1168, N342, N566, N138);
buf BUF1 (N1186, N1184);
nor NOR2 (N1187, N1180, N1048);
xor XOR2 (N1188, N1185, N571);
not NOT1 (N1189, N1182);
nor NOR2 (N1190, N1183, N493);
not NOT1 (N1191, N1181);
xor XOR2 (N1192, N1190, N1089);
and AND3 (N1193, N1189, N647, N994);
not NOT1 (N1194, N1192);
not NOT1 (N1195, N1186);
buf BUF1 (N1196, N1173);
not NOT1 (N1197, N1187);
and AND4 (N1198, N1196, N45, N648, N1092);
and AND4 (N1199, N1176, N368, N895, N394);
xor XOR2 (N1200, N1188, N74);
or OR4 (N1201, N1165, N308, N587, N680);
nand NAND3 (N1202, N1201, N40, N548);
nor NOR4 (N1203, N1199, N347, N1145, N845);
nor NOR4 (N1204, N1193, N734, N631, N751);
xor XOR2 (N1205, N1198, N839);
and AND2 (N1206, N1191, N689);
xor XOR2 (N1207, N1200, N68);
xor XOR2 (N1208, N1194, N737);
buf BUF1 (N1209, N1203);
nand NAND4 (N1210, N1207, N82, N966, N855);
or OR3 (N1211, N1210, N724, N486);
and AND2 (N1212, N1209, N1167);
nand NAND2 (N1213, N1204, N707);
xor XOR2 (N1214, N1212, N119);
buf BUF1 (N1215, N1205);
buf BUF1 (N1216, N1157);
nor NOR2 (N1217, N1208, N620);
buf BUF1 (N1218, N1206);
not NOT1 (N1219, N1213);
and AND3 (N1220, N1219, N976, N172);
and AND3 (N1221, N1202, N403, N174);
not NOT1 (N1222, N1221);
xor XOR2 (N1223, N1211, N87);
not NOT1 (N1224, N1217);
or OR4 (N1225, N1224, N1013, N1022, N1051);
xor XOR2 (N1226, N1197, N932);
and AND4 (N1227, N1220, N1075, N330, N914);
or OR4 (N1228, N1218, N622, N604, N1193);
not NOT1 (N1229, N1228);
not NOT1 (N1230, N1216);
xor XOR2 (N1231, N1215, N483);
nand NAND2 (N1232, N1223, N619);
buf BUF1 (N1233, N1232);
not NOT1 (N1234, N1225);
xor XOR2 (N1235, N1226, N148);
or OR4 (N1236, N1229, N713, N26, N956);
xor XOR2 (N1237, N1214, N524);
xor XOR2 (N1238, N1227, N913);
and AND2 (N1239, N1230, N330);
not NOT1 (N1240, N1239);
buf BUF1 (N1241, N1236);
and AND3 (N1242, N1233, N809, N440);
nor NOR4 (N1243, N1234, N48, N148, N1062);
and AND2 (N1244, N1241, N1042);
xor XOR2 (N1245, N1222, N314);
nand NAND3 (N1246, N1237, N79, N602);
nor NOR4 (N1247, N1235, N222, N1144, N389);
nor NOR2 (N1248, N1231, N1100);
buf BUF1 (N1249, N1248);
nand NAND4 (N1250, N1246, N705, N857, N1238);
or OR3 (N1251, N154, N195, N255);
not NOT1 (N1252, N1242);
buf BUF1 (N1253, N1252);
or OR4 (N1254, N1240, N860, N111, N733);
nand NAND2 (N1255, N1243, N1100);
and AND4 (N1256, N1253, N534, N747, N764);
and AND2 (N1257, N1245, N226);
nor NOR4 (N1258, N1254, N40, N1065, N699);
xor XOR2 (N1259, N1251, N117);
or OR3 (N1260, N1257, N1081, N74);
buf BUF1 (N1261, N1195);
buf BUF1 (N1262, N1260);
xor XOR2 (N1263, N1262, N124);
and AND4 (N1264, N1250, N812, N559, N616);
nor NOR2 (N1265, N1255, N930);
or OR2 (N1266, N1258, N593);
not NOT1 (N1267, N1244);
or OR4 (N1268, N1259, N1261, N221, N276);
xor XOR2 (N1269, N871, N972);
nand NAND4 (N1270, N1269, N1244, N939, N809);
not NOT1 (N1271, N1266);
buf BUF1 (N1272, N1267);
or OR3 (N1273, N1271, N72, N735);
and AND4 (N1274, N1272, N1190, N176, N1185);
or OR2 (N1275, N1249, N1028);
not NOT1 (N1276, N1264);
buf BUF1 (N1277, N1276);
buf BUF1 (N1278, N1256);
nand NAND4 (N1279, N1273, N589, N468, N458);
xor XOR2 (N1280, N1277, N1010);
not NOT1 (N1281, N1247);
or OR4 (N1282, N1265, N798, N1216, N347);
or OR2 (N1283, N1278, N67);
not NOT1 (N1284, N1268);
not NOT1 (N1285, N1283);
or OR2 (N1286, N1284, N940);
buf BUF1 (N1287, N1263);
and AND4 (N1288, N1282, N3, N1067, N549);
buf BUF1 (N1289, N1281);
not NOT1 (N1290, N1270);
nor NOR2 (N1291, N1275, N861);
nor NOR4 (N1292, N1287, N1231, N1116, N321);
not NOT1 (N1293, N1285);
nor NOR3 (N1294, N1288, N131, N582);
not NOT1 (N1295, N1279);
or OR3 (N1296, N1291, N682, N133);
buf BUF1 (N1297, N1294);
and AND2 (N1298, N1280, N380);
nor NOR4 (N1299, N1290, N268, N272, N1018);
not NOT1 (N1300, N1292);
and AND4 (N1301, N1299, N567, N99, N936);
nor NOR2 (N1302, N1286, N671);
or OR2 (N1303, N1301, N1050);
buf BUF1 (N1304, N1289);
or OR4 (N1305, N1300, N281, N742, N408);
nand NAND4 (N1306, N1274, N992, N1037, N1248);
nand NAND3 (N1307, N1303, N322, N716);
and AND3 (N1308, N1295, N148, N1252);
xor XOR2 (N1309, N1298, N570);
not NOT1 (N1310, N1304);
buf BUF1 (N1311, N1308);
or OR2 (N1312, N1311, N133);
xor XOR2 (N1313, N1307, N306);
nor NOR3 (N1314, N1313, N805, N272);
buf BUF1 (N1315, N1293);
buf BUF1 (N1316, N1312);
not NOT1 (N1317, N1314);
buf BUF1 (N1318, N1297);
buf BUF1 (N1319, N1306);
xor XOR2 (N1320, N1316, N234);
buf BUF1 (N1321, N1315);
not NOT1 (N1322, N1305);
nor NOR2 (N1323, N1302, N1000);
and AND4 (N1324, N1318, N1276, N796, N339);
and AND3 (N1325, N1309, N1323, N1011);
xor XOR2 (N1326, N1002, N571);
nor NOR2 (N1327, N1322, N315);
xor XOR2 (N1328, N1327, N349);
and AND4 (N1329, N1321, N108, N426, N725);
not NOT1 (N1330, N1328);
xor XOR2 (N1331, N1329, N305);
buf BUF1 (N1332, N1319);
nand NAND2 (N1333, N1331, N2);
buf BUF1 (N1334, N1325);
nor NOR3 (N1335, N1310, N763, N647);
nor NOR2 (N1336, N1296, N749);
nand NAND4 (N1337, N1335, N891, N957, N1100);
nor NOR3 (N1338, N1330, N143, N144);
and AND2 (N1339, N1317, N36);
or OR4 (N1340, N1320, N337, N308, N75);
buf BUF1 (N1341, N1336);
buf BUF1 (N1342, N1337);
buf BUF1 (N1343, N1338);
buf BUF1 (N1344, N1333);
nor NOR3 (N1345, N1332, N727, N325);
or OR3 (N1346, N1342, N528, N1004);
xor XOR2 (N1347, N1341, N955);
nor NOR4 (N1348, N1344, N1285, N46, N562);
nor NOR4 (N1349, N1345, N687, N521, N675);
nand NAND4 (N1350, N1343, N211, N195, N999);
not NOT1 (N1351, N1348);
nand NAND3 (N1352, N1334, N729, N1214);
nor NOR2 (N1353, N1347, N214);
xor XOR2 (N1354, N1351, N915);
nor NOR4 (N1355, N1346, N1211, N696, N859);
or OR4 (N1356, N1355, N637, N482, N90);
not NOT1 (N1357, N1352);
or OR3 (N1358, N1349, N515, N540);
and AND4 (N1359, N1339, N536, N911, N103);
not NOT1 (N1360, N1358);
xor XOR2 (N1361, N1357, N1070);
nor NOR4 (N1362, N1324, N1203, N914, N585);
and AND4 (N1363, N1340, N252, N973, N1245);
and AND2 (N1364, N1350, N775);
not NOT1 (N1365, N1354);
xor XOR2 (N1366, N1363, N964);
nand NAND4 (N1367, N1365, N567, N68, N16);
and AND3 (N1368, N1367, N906, N127);
or OR2 (N1369, N1361, N396);
nand NAND2 (N1370, N1356, N191);
buf BUF1 (N1371, N1362);
buf BUF1 (N1372, N1326);
nand NAND2 (N1373, N1371, N862);
nand NAND2 (N1374, N1360, N192);
nand NAND4 (N1375, N1368, N399, N860, N662);
buf BUF1 (N1376, N1370);
nor NOR3 (N1377, N1366, N884, N719);
or OR2 (N1378, N1369, N1137);
xor XOR2 (N1379, N1374, N1210);
buf BUF1 (N1380, N1377);
not NOT1 (N1381, N1364);
nor NOR4 (N1382, N1378, N630, N295, N474);
and AND3 (N1383, N1382, N849, N151);
or OR3 (N1384, N1381, N1014, N900);
and AND4 (N1385, N1353, N313, N467, N421);
or OR2 (N1386, N1373, N1089);
xor XOR2 (N1387, N1359, N458);
buf BUF1 (N1388, N1383);
buf BUF1 (N1389, N1388);
and AND2 (N1390, N1376, N433);
xor XOR2 (N1391, N1385, N516);
and AND3 (N1392, N1389, N838, N19);
nand NAND2 (N1393, N1387, N951);
nand NAND4 (N1394, N1379, N229, N85, N1219);
or OR2 (N1395, N1386, N929);
xor XOR2 (N1396, N1394, N923);
and AND4 (N1397, N1393, N1222, N835, N1170);
buf BUF1 (N1398, N1380);
not NOT1 (N1399, N1390);
xor XOR2 (N1400, N1372, N1053);
not NOT1 (N1401, N1396);
and AND4 (N1402, N1392, N512, N1353, N1205);
buf BUF1 (N1403, N1375);
nand NAND2 (N1404, N1402, N119);
not NOT1 (N1405, N1400);
not NOT1 (N1406, N1391);
not NOT1 (N1407, N1404);
xor XOR2 (N1408, N1398, N1393);
nor NOR2 (N1409, N1395, N398);
xor XOR2 (N1410, N1384, N1053);
xor XOR2 (N1411, N1407, N1390);
and AND4 (N1412, N1405, N261, N195, N312);
not NOT1 (N1413, N1401);
and AND3 (N1414, N1397, N1157, N544);
and AND3 (N1415, N1403, N824, N1126);
and AND3 (N1416, N1412, N643, N194);
xor XOR2 (N1417, N1415, N1321);
nor NOR4 (N1418, N1417, N725, N1124, N258);
xor XOR2 (N1419, N1406, N1278);
not NOT1 (N1420, N1413);
or OR4 (N1421, N1399, N1174, N633, N254);
nand NAND4 (N1422, N1421, N150, N1231, N75);
and AND4 (N1423, N1409, N427, N1388, N721);
not NOT1 (N1424, N1408);
xor XOR2 (N1425, N1420, N598);
not NOT1 (N1426, N1419);
nor NOR3 (N1427, N1424, N854, N793);
xor XOR2 (N1428, N1411, N911);
buf BUF1 (N1429, N1428);
xor XOR2 (N1430, N1427, N1373);
nor NOR2 (N1431, N1426, N308);
xor XOR2 (N1432, N1410, N1072);
nor NOR4 (N1433, N1422, N1074, N1390, N1138);
or OR4 (N1434, N1431, N1167, N906, N14);
nand NAND3 (N1435, N1425, N226, N987);
or OR4 (N1436, N1435, N416, N299, N982);
buf BUF1 (N1437, N1430);
not NOT1 (N1438, N1436);
buf BUF1 (N1439, N1432);
buf BUF1 (N1440, N1423);
nand NAND4 (N1441, N1439, N587, N122, N872);
buf BUF1 (N1442, N1438);
and AND4 (N1443, N1437, N1269, N731, N422);
nor NOR3 (N1444, N1434, N1321, N458);
xor XOR2 (N1445, N1443, N271);
and AND3 (N1446, N1444, N1127, N212);
or OR2 (N1447, N1441, N374);
or OR4 (N1448, N1445, N166, N1313, N185);
xor XOR2 (N1449, N1442, N658);
not NOT1 (N1450, N1416);
not NOT1 (N1451, N1440);
nor NOR2 (N1452, N1446, N614);
buf BUF1 (N1453, N1414);
nor NOR4 (N1454, N1418, N9, N210, N251);
buf BUF1 (N1455, N1449);
nor NOR2 (N1456, N1429, N973);
nand NAND2 (N1457, N1452, N1041);
nand NAND3 (N1458, N1448, N747, N1142);
nand NAND2 (N1459, N1456, N622);
xor XOR2 (N1460, N1457, N110);
not NOT1 (N1461, N1451);
xor XOR2 (N1462, N1450, N1290);
nor NOR4 (N1463, N1459, N666, N648, N150);
nand NAND4 (N1464, N1461, N61, N532, N1230);
nand NAND2 (N1465, N1455, N997);
nand NAND4 (N1466, N1453, N1070, N244, N749);
nand NAND4 (N1467, N1433, N750, N1394, N693);
nand NAND3 (N1468, N1464, N1256, N174);
or OR4 (N1469, N1454, N266, N816, N117);
or OR4 (N1470, N1466, N9, N1459, N1397);
buf BUF1 (N1471, N1469);
or OR2 (N1472, N1467, N931);
buf BUF1 (N1473, N1465);
nor NOR3 (N1474, N1462, N1284, N1399);
buf BUF1 (N1475, N1458);
nor NOR2 (N1476, N1468, N1036);
buf BUF1 (N1477, N1463);
or OR2 (N1478, N1473, N744);
and AND3 (N1479, N1471, N1167, N421);
nand NAND2 (N1480, N1474, N278);
and AND2 (N1481, N1475, N1192);
xor XOR2 (N1482, N1480, N25);
or OR4 (N1483, N1477, N689, N61, N1109);
nand NAND3 (N1484, N1481, N344, N401);
xor XOR2 (N1485, N1460, N544);
or OR2 (N1486, N1447, N1387);
not NOT1 (N1487, N1470);
and AND2 (N1488, N1487, N590);
nor NOR3 (N1489, N1478, N699, N1269);
nor NOR2 (N1490, N1476, N391);
not NOT1 (N1491, N1485);
and AND4 (N1492, N1472, N662, N612, N501);
nand NAND3 (N1493, N1486, N148, N662);
or OR3 (N1494, N1479, N476, N807);
not NOT1 (N1495, N1488);
and AND4 (N1496, N1493, N5, N65, N39);
nor NOR2 (N1497, N1492, N1427);
nor NOR2 (N1498, N1490, N1247);
and AND4 (N1499, N1489, N1205, N21, N471);
buf BUF1 (N1500, N1494);
not NOT1 (N1501, N1484);
xor XOR2 (N1502, N1496, N523);
xor XOR2 (N1503, N1501, N525);
and AND3 (N1504, N1502, N228, N861);
or OR3 (N1505, N1497, N1232, N1275);
or OR3 (N1506, N1498, N1034, N252);
and AND3 (N1507, N1504, N735, N882);
buf BUF1 (N1508, N1499);
xor XOR2 (N1509, N1491, N698);
and AND4 (N1510, N1503, N1205, N794, N708);
xor XOR2 (N1511, N1495, N79);
nor NOR3 (N1512, N1507, N221, N1111);
nand NAND3 (N1513, N1500, N490, N855);
and AND4 (N1514, N1513, N180, N745, N33);
buf BUF1 (N1515, N1509);
xor XOR2 (N1516, N1506, N232);
and AND4 (N1517, N1482, N389, N211, N1454);
not NOT1 (N1518, N1514);
nor NOR3 (N1519, N1512, N1446, N1432);
buf BUF1 (N1520, N1519);
xor XOR2 (N1521, N1483, N797);
not NOT1 (N1522, N1518);
and AND3 (N1523, N1511, N1104, N545);
nand NAND3 (N1524, N1508, N1039, N1000);
and AND4 (N1525, N1517, N626, N1518, N657);
not NOT1 (N1526, N1525);
nand NAND4 (N1527, N1524, N645, N599, N486);
nor NOR3 (N1528, N1521, N319, N197);
nand NAND2 (N1529, N1523, N1012);
or OR2 (N1530, N1516, N616);
nand NAND2 (N1531, N1515, N1220);
not NOT1 (N1532, N1531);
not NOT1 (N1533, N1530);
nor NOR4 (N1534, N1529, N1105, N3, N988);
nand NAND4 (N1535, N1528, N587, N986, N891);
xor XOR2 (N1536, N1505, N554);
nand NAND4 (N1537, N1520, N345, N1374, N1262);
or OR2 (N1538, N1536, N1291);
xor XOR2 (N1539, N1526, N486);
nand NAND2 (N1540, N1535, N985);
or OR4 (N1541, N1539, N984, N524, N890);
xor XOR2 (N1542, N1534, N953);
nand NAND4 (N1543, N1540, N270, N411, N1322);
or OR4 (N1544, N1510, N1521, N874, N774);
nand NAND2 (N1545, N1543, N442);
or OR3 (N1546, N1532, N682, N3);
and AND3 (N1547, N1544, N1472, N425);
not NOT1 (N1548, N1547);
not NOT1 (N1549, N1546);
not NOT1 (N1550, N1541);
and AND4 (N1551, N1537, N179, N481, N219);
and AND2 (N1552, N1538, N1341);
xor XOR2 (N1553, N1550, N1179);
nor NOR3 (N1554, N1552, N426, N1120);
or OR3 (N1555, N1542, N346, N1148);
or OR4 (N1556, N1553, N1091, N353, N617);
nand NAND4 (N1557, N1545, N1342, N463, N849);
or OR3 (N1558, N1522, N498, N1303);
or OR2 (N1559, N1551, N1046);
xor XOR2 (N1560, N1556, N200);
not NOT1 (N1561, N1559);
and AND4 (N1562, N1557, N1555, N922, N1561);
or OR2 (N1563, N609, N85);
nor NOR3 (N1564, N1236, N7, N553);
xor XOR2 (N1565, N1560, N474);
nor NOR3 (N1566, N1558, N847, N176);
not NOT1 (N1567, N1565);
nor NOR2 (N1568, N1549, N13);
xor XOR2 (N1569, N1533, N205);
buf BUF1 (N1570, N1548);
nor NOR3 (N1571, N1566, N185, N20);
xor XOR2 (N1572, N1569, N1188);
xor XOR2 (N1573, N1567, N131);
nand NAND3 (N1574, N1573, N778, N67);
nor NOR4 (N1575, N1568, N1240, N1565, N372);
nor NOR2 (N1576, N1563, N809);
buf BUF1 (N1577, N1575);
or OR4 (N1578, N1562, N194, N1194, N1569);
xor XOR2 (N1579, N1572, N787);
buf BUF1 (N1580, N1527);
or OR4 (N1581, N1554, N1052, N1342, N991);
and AND2 (N1582, N1581, N751);
not NOT1 (N1583, N1576);
not NOT1 (N1584, N1571);
not NOT1 (N1585, N1584);
or OR2 (N1586, N1574, N50);
buf BUF1 (N1587, N1578);
not NOT1 (N1588, N1582);
nand NAND2 (N1589, N1564, N1055);
and AND2 (N1590, N1585, N85);
or OR2 (N1591, N1570, N317);
nor NOR4 (N1592, N1589, N353, N1125, N959);
not NOT1 (N1593, N1591);
xor XOR2 (N1594, N1587, N1121);
and AND4 (N1595, N1590, N596, N1220, N146);
nand NAND2 (N1596, N1595, N1224);
not NOT1 (N1597, N1586);
or OR2 (N1598, N1597, N813);
buf BUF1 (N1599, N1593);
and AND2 (N1600, N1580, N9);
not NOT1 (N1601, N1598);
nor NOR3 (N1602, N1583, N892, N585);
and AND3 (N1603, N1600, N216, N843);
nand NAND2 (N1604, N1588, N878);
nand NAND3 (N1605, N1602, N407, N1582);
or OR4 (N1606, N1599, N691, N479, N667);
or OR3 (N1607, N1592, N1559, N535);
and AND2 (N1608, N1601, N1512);
buf BUF1 (N1609, N1596);
xor XOR2 (N1610, N1577, N64);
xor XOR2 (N1611, N1610, N1211);
or OR3 (N1612, N1605, N859, N50);
or OR2 (N1613, N1603, N1222);
nand NAND4 (N1614, N1612, N17, N1118, N8);
nor NOR4 (N1615, N1609, N44, N753, N1061);
nand NAND3 (N1616, N1594, N188, N890);
nor NOR2 (N1617, N1616, N524);
nand NAND2 (N1618, N1614, N1585);
and AND3 (N1619, N1611, N869, N1009);
nor NOR2 (N1620, N1606, N279);
xor XOR2 (N1621, N1620, N389);
not NOT1 (N1622, N1613);
buf BUF1 (N1623, N1618);
or OR2 (N1624, N1617, N891);
nand NAND3 (N1625, N1604, N773, N1200);
nand NAND4 (N1626, N1619, N548, N25, N410);
or OR3 (N1627, N1624, N358, N1491);
xor XOR2 (N1628, N1621, N1062);
or OR2 (N1629, N1625, N1007);
nor NOR3 (N1630, N1615, N1327, N516);
nor NOR4 (N1631, N1608, N1560, N1357, N1440);
nor NOR3 (N1632, N1629, N1415, N59);
not NOT1 (N1633, N1626);
not NOT1 (N1634, N1622);
nor NOR4 (N1635, N1631, N1510, N1058, N1240);
xor XOR2 (N1636, N1633, N188);
xor XOR2 (N1637, N1607, N8);
xor XOR2 (N1638, N1634, N1136);
and AND2 (N1639, N1637, N406);
nand NAND3 (N1640, N1636, N1334, N1207);
not NOT1 (N1641, N1635);
buf BUF1 (N1642, N1638);
nand NAND3 (N1643, N1630, N290, N953);
xor XOR2 (N1644, N1627, N1170);
xor XOR2 (N1645, N1642, N458);
nor NOR3 (N1646, N1644, N1355, N185);
not NOT1 (N1647, N1623);
nor NOR4 (N1648, N1628, N712, N713, N298);
nor NOR3 (N1649, N1640, N952, N268);
nor NOR3 (N1650, N1647, N684, N897);
nor NOR2 (N1651, N1650, N713);
not NOT1 (N1652, N1639);
not NOT1 (N1653, N1652);
and AND2 (N1654, N1646, N27);
and AND4 (N1655, N1651, N441, N1122, N622);
not NOT1 (N1656, N1632);
xor XOR2 (N1657, N1649, N1402);
nand NAND4 (N1658, N1653, N1245, N642, N575);
and AND4 (N1659, N1658, N1216, N1394, N1308);
and AND4 (N1660, N1648, N257, N83, N4);
not NOT1 (N1661, N1643);
and AND2 (N1662, N1660, N231);
nor NOR3 (N1663, N1657, N524, N1532);
and AND3 (N1664, N1659, N289, N236);
or OR2 (N1665, N1654, N989);
nor NOR4 (N1666, N1645, N1037, N920, N870);
xor XOR2 (N1667, N1656, N1041);
buf BUF1 (N1668, N1655);
buf BUF1 (N1669, N1665);
buf BUF1 (N1670, N1666);
not NOT1 (N1671, N1641);
or OR4 (N1672, N1663, N1236, N488, N1634);
nand NAND4 (N1673, N1670, N380, N10, N540);
xor XOR2 (N1674, N1661, N155);
xor XOR2 (N1675, N1674, N945);
nor NOR3 (N1676, N1672, N115, N1545);
and AND3 (N1677, N1668, N1573, N1233);
and AND4 (N1678, N1664, N1661, N60, N715);
not NOT1 (N1679, N1676);
or OR3 (N1680, N1662, N1204, N1329);
xor XOR2 (N1681, N1671, N861);
not NOT1 (N1682, N1678);
and AND3 (N1683, N1677, N1093, N1657);
or OR4 (N1684, N1673, N1164, N674, N41);
nor NOR4 (N1685, N1667, N1310, N324, N836);
nand NAND3 (N1686, N1681, N1095, N131);
not NOT1 (N1687, N1685);
or OR4 (N1688, N1579, N1503, N93, N947);
not NOT1 (N1689, N1682);
nor NOR2 (N1690, N1679, N820);
and AND2 (N1691, N1689, N903);
or OR4 (N1692, N1680, N729, N722, N1077);
xor XOR2 (N1693, N1692, N309);
nand NAND4 (N1694, N1688, N1691, N742, N780);
and AND4 (N1695, N579, N1205, N1268, N1346);
or OR4 (N1696, N1695, N1648, N1424, N221);
or OR4 (N1697, N1690, N1643, N1401, N271);
nand NAND3 (N1698, N1675, N236, N1594);
not NOT1 (N1699, N1669);
or OR2 (N1700, N1684, N787);
xor XOR2 (N1701, N1700, N336);
buf BUF1 (N1702, N1699);
nor NOR2 (N1703, N1693, N18);
xor XOR2 (N1704, N1702, N1690);
not NOT1 (N1705, N1698);
or OR4 (N1706, N1687, N121, N847, N1381);
nor NOR2 (N1707, N1706, N979);
or OR3 (N1708, N1686, N1015, N189);
xor XOR2 (N1709, N1705, N1020);
buf BUF1 (N1710, N1704);
nand NAND3 (N1711, N1707, N1326, N1271);
and AND4 (N1712, N1683, N547, N1292, N1452);
buf BUF1 (N1713, N1701);
buf BUF1 (N1714, N1713);
or OR4 (N1715, N1703, N951, N192, N705);
or OR4 (N1716, N1696, N1641, N625, N1501);
buf BUF1 (N1717, N1712);
nor NOR2 (N1718, N1708, N1532);
nand NAND2 (N1719, N1717, N1441);
or OR3 (N1720, N1714, N874, N769);
nand NAND3 (N1721, N1711, N1423, N682);
buf BUF1 (N1722, N1697);
and AND3 (N1723, N1715, N125, N1612);
buf BUF1 (N1724, N1720);
or OR2 (N1725, N1724, N7);
and AND4 (N1726, N1719, N1268, N1197, N1390);
nand NAND3 (N1727, N1709, N1284, N386);
nand NAND3 (N1728, N1721, N1490, N405);
buf BUF1 (N1729, N1722);
not NOT1 (N1730, N1728);
and AND4 (N1731, N1718, N582, N1601, N158);
buf BUF1 (N1732, N1727);
nor NOR3 (N1733, N1725, N693, N746);
nor NOR2 (N1734, N1726, N58);
or OR2 (N1735, N1729, N1671);
nand NAND4 (N1736, N1716, N1117, N274, N25);
nand NAND3 (N1737, N1736, N626, N661);
nand NAND3 (N1738, N1732, N587, N1010);
buf BUF1 (N1739, N1733);
not NOT1 (N1740, N1738);
nand NAND3 (N1741, N1737, N255, N118);
and AND2 (N1742, N1710, N995);
xor XOR2 (N1743, N1730, N1551);
nor NOR4 (N1744, N1735, N85, N840, N1062);
and AND3 (N1745, N1734, N1410, N1005);
xor XOR2 (N1746, N1740, N789);
or OR3 (N1747, N1745, N518, N1720);
not NOT1 (N1748, N1747);
or OR2 (N1749, N1741, N49);
not NOT1 (N1750, N1744);
not NOT1 (N1751, N1746);
buf BUF1 (N1752, N1743);
nor NOR3 (N1753, N1723, N836, N424);
nand NAND4 (N1754, N1739, N1310, N370, N563);
or OR2 (N1755, N1751, N489);
nor NOR4 (N1756, N1694, N1387, N900, N523);
buf BUF1 (N1757, N1742);
or OR4 (N1758, N1755, N1453, N573, N227);
and AND4 (N1759, N1750, N429, N1748, N1094);
nor NOR3 (N1760, N923, N1175, N1263);
buf BUF1 (N1761, N1754);
not NOT1 (N1762, N1749);
xor XOR2 (N1763, N1756, N595);
nand NAND4 (N1764, N1759, N340, N1505, N756);
xor XOR2 (N1765, N1763, N1714);
and AND3 (N1766, N1762, N775, N177);
or OR2 (N1767, N1761, N1402);
not NOT1 (N1768, N1765);
buf BUF1 (N1769, N1768);
and AND2 (N1770, N1757, N1295);
nor NOR4 (N1771, N1753, N929, N88, N1284);
or OR2 (N1772, N1760, N658);
or OR3 (N1773, N1769, N843, N74);
buf BUF1 (N1774, N1752);
xor XOR2 (N1775, N1773, N241);
buf BUF1 (N1776, N1767);
and AND3 (N1777, N1758, N750, N1753);
or OR4 (N1778, N1731, N668, N1530, N198);
xor XOR2 (N1779, N1772, N1020);
or OR2 (N1780, N1779, N169);
and AND3 (N1781, N1780, N754, N1693);
and AND3 (N1782, N1764, N1561, N1328);
nor NOR4 (N1783, N1777, N1482, N1567, N128);
buf BUF1 (N1784, N1774);
nor NOR2 (N1785, N1776, N914);
and AND2 (N1786, N1766, N1145);
not NOT1 (N1787, N1785);
xor XOR2 (N1788, N1775, N1387);
or OR3 (N1789, N1770, N1008, N1137);
buf BUF1 (N1790, N1778);
buf BUF1 (N1791, N1789);
xor XOR2 (N1792, N1783, N259);
or OR3 (N1793, N1786, N163, N815);
nand NAND3 (N1794, N1793, N944, N541);
not NOT1 (N1795, N1781);
buf BUF1 (N1796, N1794);
not NOT1 (N1797, N1788);
nand NAND2 (N1798, N1790, N176);
nor NOR4 (N1799, N1771, N80, N434, N1357);
xor XOR2 (N1800, N1796, N1575);
xor XOR2 (N1801, N1798, N192);
not NOT1 (N1802, N1799);
and AND4 (N1803, N1782, N1494, N1802, N1677);
or OR2 (N1804, N484, N510);
or OR2 (N1805, N1801, N1248);
buf BUF1 (N1806, N1791);
nor NOR3 (N1807, N1784, N852, N505);
nor NOR4 (N1808, N1795, N758, N1647, N1786);
not NOT1 (N1809, N1807);
not NOT1 (N1810, N1787);
buf BUF1 (N1811, N1805);
nor NOR4 (N1812, N1792, N1216, N1681, N1544);
nand NAND2 (N1813, N1809, N276);
buf BUF1 (N1814, N1800);
nor NOR4 (N1815, N1806, N813, N260, N218);
buf BUF1 (N1816, N1811);
nor NOR4 (N1817, N1813, N1500, N1649, N217);
not NOT1 (N1818, N1797);
and AND2 (N1819, N1814, N314);
xor XOR2 (N1820, N1817, N52);
nor NOR2 (N1821, N1808, N1070);
nor NOR3 (N1822, N1820, N1317, N1338);
buf BUF1 (N1823, N1804);
or OR3 (N1824, N1810, N761, N649);
nand NAND4 (N1825, N1824, N908, N546, N500);
nand NAND2 (N1826, N1803, N1418);
xor XOR2 (N1827, N1825, N1792);
not NOT1 (N1828, N1819);
nor NOR3 (N1829, N1822, N1506, N1049);
nor NOR4 (N1830, N1828, N1735, N180, N225);
nor NOR2 (N1831, N1818, N1130);
or OR4 (N1832, N1812, N675, N965, N1314);
not NOT1 (N1833, N1829);
or OR2 (N1834, N1823, N1494);
xor XOR2 (N1835, N1833, N9);
not NOT1 (N1836, N1816);
not NOT1 (N1837, N1821);
not NOT1 (N1838, N1827);
and AND4 (N1839, N1836, N1569, N321, N734);
nor NOR3 (N1840, N1839, N427, N1735);
or OR4 (N1841, N1826, N1030, N383, N724);
buf BUF1 (N1842, N1840);
buf BUF1 (N1843, N1842);
buf BUF1 (N1844, N1843);
nor NOR2 (N1845, N1832, N1120);
nand NAND2 (N1846, N1835, N1634);
not NOT1 (N1847, N1834);
buf BUF1 (N1848, N1845);
not NOT1 (N1849, N1831);
nand NAND2 (N1850, N1838, N1566);
nand NAND4 (N1851, N1815, N1051, N1347, N1066);
buf BUF1 (N1852, N1846);
nand NAND3 (N1853, N1841, N1007, N650);
nand NAND3 (N1854, N1847, N1709, N1508);
and AND2 (N1855, N1851, N1232);
xor XOR2 (N1856, N1852, N901);
and AND4 (N1857, N1830, N1778, N549, N624);
not NOT1 (N1858, N1854);
nor NOR3 (N1859, N1855, N1470, N1351);
or OR2 (N1860, N1849, N206);
nor NOR3 (N1861, N1850, N7, N172);
buf BUF1 (N1862, N1858);
or OR4 (N1863, N1859, N1409, N1488, N215);
or OR4 (N1864, N1837, N948, N343, N1106);
xor XOR2 (N1865, N1862, N1422);
nor NOR2 (N1866, N1853, N45);
nand NAND4 (N1867, N1861, N1281, N1532, N318);
nand NAND3 (N1868, N1867, N768, N1303);
nor NOR2 (N1869, N1857, N1460);
or OR2 (N1870, N1868, N218);
not NOT1 (N1871, N1860);
xor XOR2 (N1872, N1870, N1405);
nand NAND3 (N1873, N1869, N1847, N1155);
nand NAND2 (N1874, N1865, N428);
xor XOR2 (N1875, N1873, N1156);
or OR3 (N1876, N1866, N122, N1192);
and AND4 (N1877, N1863, N1017, N1732, N1779);
and AND2 (N1878, N1876, N281);
not NOT1 (N1879, N1864);
nor NOR2 (N1880, N1844, N972);
xor XOR2 (N1881, N1872, N884);
nand NAND4 (N1882, N1881, N803, N454, N1745);
not NOT1 (N1883, N1882);
xor XOR2 (N1884, N1848, N1157);
buf BUF1 (N1885, N1877);
buf BUF1 (N1886, N1879);
not NOT1 (N1887, N1886);
xor XOR2 (N1888, N1874, N331);
buf BUF1 (N1889, N1871);
xor XOR2 (N1890, N1878, N1837);
not NOT1 (N1891, N1885);
buf BUF1 (N1892, N1891);
nand NAND3 (N1893, N1884, N157, N1177);
buf BUF1 (N1894, N1892);
and AND3 (N1895, N1889, N926, N495);
xor XOR2 (N1896, N1895, N1404);
or OR3 (N1897, N1887, N1667, N1143);
xor XOR2 (N1898, N1890, N596);
not NOT1 (N1899, N1856);
buf BUF1 (N1900, N1880);
nor NOR3 (N1901, N1900, N1841, N934);
buf BUF1 (N1902, N1893);
not NOT1 (N1903, N1898);
not NOT1 (N1904, N1903);
not NOT1 (N1905, N1875);
nand NAND3 (N1906, N1899, N1857, N349);
buf BUF1 (N1907, N1897);
or OR3 (N1908, N1907, N1448, N594);
or OR2 (N1909, N1883, N1897);
nand NAND4 (N1910, N1888, N534, N1592, N1453);
not NOT1 (N1911, N1896);
nand NAND3 (N1912, N1902, N776, N1857);
nor NOR3 (N1913, N1905, N1590, N1859);
or OR3 (N1914, N1894, N1371, N457);
and AND2 (N1915, N1911, N136);
and AND2 (N1916, N1909, N669);
nor NOR2 (N1917, N1916, N772);
buf BUF1 (N1918, N1914);
nand NAND4 (N1919, N1915, N444, N1690, N1343);
and AND4 (N1920, N1904, N876, N726, N450);
xor XOR2 (N1921, N1918, N312);
and AND3 (N1922, N1906, N62, N933);
and AND4 (N1923, N1921, N50, N1017, N142);
and AND4 (N1924, N1913, N351, N851, N82);
and AND3 (N1925, N1901, N1729, N18);
or OR4 (N1926, N1919, N1300, N846, N236);
buf BUF1 (N1927, N1920);
or OR3 (N1928, N1917, N1533, N608);
not NOT1 (N1929, N1912);
nor NOR4 (N1930, N1908, N974, N1518, N1382);
not NOT1 (N1931, N1930);
xor XOR2 (N1932, N1924, N337);
not NOT1 (N1933, N1923);
nand NAND2 (N1934, N1928, N690);
buf BUF1 (N1935, N1926);
nor NOR4 (N1936, N1922, N1355, N298, N784);
nor NOR4 (N1937, N1932, N1360, N160, N1546);
buf BUF1 (N1938, N1934);
xor XOR2 (N1939, N1933, N1374);
buf BUF1 (N1940, N1939);
xor XOR2 (N1941, N1936, N1517);
not NOT1 (N1942, N1941);
not NOT1 (N1943, N1925);
buf BUF1 (N1944, N1942);
buf BUF1 (N1945, N1931);
buf BUF1 (N1946, N1910);
and AND4 (N1947, N1943, N1895, N1706, N1015);
or OR2 (N1948, N1938, N668);
not NOT1 (N1949, N1947);
nand NAND2 (N1950, N1949, N444);
or OR2 (N1951, N1937, N1323);
nor NOR3 (N1952, N1935, N18, N159);
or OR2 (N1953, N1940, N947);
and AND2 (N1954, N1951, N1423);
nor NOR3 (N1955, N1950, N448, N1069);
nand NAND3 (N1956, N1945, N614, N716);
and AND4 (N1957, N1948, N1665, N966, N1410);
buf BUF1 (N1958, N1954);
nor NOR3 (N1959, N1953, N745, N755);
or OR2 (N1960, N1958, N1346);
nand NAND3 (N1961, N1946, N1894, N1043);
nand NAND2 (N1962, N1929, N1211);
not NOT1 (N1963, N1960);
xor XOR2 (N1964, N1957, N590);
or OR3 (N1965, N1962, N1058, N763);
nor NOR4 (N1966, N1952, N1128, N1063, N552);
nor NOR2 (N1967, N1927, N1588);
xor XOR2 (N1968, N1963, N1129);
buf BUF1 (N1969, N1968);
not NOT1 (N1970, N1967);
or OR2 (N1971, N1964, N905);
not NOT1 (N1972, N1955);
buf BUF1 (N1973, N1961);
nand NAND3 (N1974, N1971, N1605, N1940);
not NOT1 (N1975, N1959);
and AND2 (N1976, N1974, N1250);
nand NAND2 (N1977, N1975, N1624);
nand NAND4 (N1978, N1970, N545, N1463, N826);
xor XOR2 (N1979, N1969, N1224);
and AND2 (N1980, N1979, N1004);
nand NAND3 (N1981, N1965, N1377, N1282);
and AND4 (N1982, N1980, N700, N1059, N712);
nor NOR2 (N1983, N1982, N326);
nand NAND3 (N1984, N1944, N859, N1343);
and AND3 (N1985, N1977, N408, N742);
buf BUF1 (N1986, N1972);
nor NOR4 (N1987, N1983, N940, N1297, N1501);
nand NAND3 (N1988, N1978, N1581, N1436);
or OR4 (N1989, N1976, N1870, N302, N1447);
nand NAND4 (N1990, N1988, N770, N1696, N1048);
xor XOR2 (N1991, N1981, N883);
not NOT1 (N1992, N1973);
xor XOR2 (N1993, N1985, N1166);
buf BUF1 (N1994, N1956);
not NOT1 (N1995, N1992);
not NOT1 (N1996, N1993);
buf BUF1 (N1997, N1991);
nand NAND2 (N1998, N1989, N1844);
buf BUF1 (N1999, N1990);
and AND2 (N2000, N1994, N1142);
not NOT1 (N2001, N1997);
and AND2 (N2002, N1966, N1648);
buf BUF1 (N2003, N1986);
or OR3 (N2004, N1996, N620, N1500);
or OR2 (N2005, N1999, N158);
not NOT1 (N2006, N2001);
nand NAND3 (N2007, N1984, N221, N971);
buf BUF1 (N2008, N2000);
nor NOR3 (N2009, N1998, N1277, N1447);
and AND3 (N2010, N2009, N744, N953);
not NOT1 (N2011, N2007);
nand NAND4 (N2012, N2006, N888, N8, N1785);
endmodule