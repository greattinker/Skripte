// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;

output N12812,N12820,N12818,N12783,N12805,N12821,N12822,N12823,N12817,N12824;

xor XOR2 (N25, N21, N1);
nand NAND4 (N26, N3, N12, N19, N11);
or OR4 (N27, N16, N25, N22, N26);
not NOT1 (N28, N10);
nor NOR4 (N29, N23, N13, N12, N22);
xor XOR2 (N30, N20, N10);
not NOT1 (N31, N13);
and AND2 (N32, N31, N2);
and AND4 (N33, N13, N32, N11, N6);
and AND2 (N34, N23, N19);
nand NAND2 (N35, N4, N14);
nor NOR4 (N36, N5, N11, N13, N5);
nand NAND3 (N37, N5, N33, N18);
or OR4 (N38, N34, N36, N19, N27);
and AND3 (N39, N6, N25, N33);
and AND2 (N40, N8, N23);
not NOT1 (N41, N39);
xor XOR2 (N42, N10, N19);
or OR2 (N43, N23, N5);
xor XOR2 (N44, N38, N40);
xor XOR2 (N45, N16, N4);
xor XOR2 (N46, N28, N31);
nor NOR3 (N47, N42, N17, N16);
nand NAND2 (N48, N37, N1);
nand NAND4 (N49, N44, N10, N25, N30);
nor NOR3 (N50, N10, N14, N39);
xor XOR2 (N51, N50, N1);
and AND2 (N52, N49, N19);
not NOT1 (N53, N46);
buf BUF1 (N54, N52);
not NOT1 (N55, N53);
nand NAND2 (N56, N47, N26);
buf BUF1 (N57, N41);
or OR3 (N58, N43, N5, N6);
or OR2 (N59, N55, N25);
nand NAND4 (N60, N59, N21, N17, N55);
or OR3 (N61, N58, N1, N7);
nor NOR3 (N62, N57, N13, N35);
and AND4 (N63, N51, N46, N16, N59);
buf BUF1 (N64, N55);
buf BUF1 (N65, N60);
and AND3 (N66, N54, N60, N5);
not NOT1 (N67, N66);
nor NOR2 (N68, N67, N65);
nand NAND3 (N69, N67, N47, N19);
buf BUF1 (N70, N64);
nor NOR2 (N71, N68, N67);
not NOT1 (N72, N29);
and AND4 (N73, N70, N35, N31, N56);
xor XOR2 (N74, N29, N53);
not NOT1 (N75, N62);
not NOT1 (N76, N73);
and AND4 (N77, N48, N74, N8, N53);
and AND3 (N78, N35, N54, N44);
buf BUF1 (N79, N76);
not NOT1 (N80, N45);
and AND4 (N81, N77, N7, N5, N64);
xor XOR2 (N82, N69, N19);
and AND2 (N83, N80, N45);
not NOT1 (N84, N75);
nor NOR3 (N85, N78, N83, N57);
and AND2 (N86, N57, N41);
and AND3 (N87, N85, N19, N16);
xor XOR2 (N88, N72, N19);
buf BUF1 (N89, N81);
and AND4 (N90, N86, N29, N32, N32);
and AND4 (N91, N89, N62, N17, N44);
nor NOR2 (N92, N82, N11);
nor NOR3 (N93, N84, N32, N14);
nand NAND3 (N94, N87, N86, N43);
or OR3 (N95, N90, N35, N18);
nor NOR4 (N96, N71, N70, N79, N1);
buf BUF1 (N97, N25);
xor XOR2 (N98, N94, N38);
xor XOR2 (N99, N95, N31);
or OR4 (N100, N63, N41, N46, N28);
or OR3 (N101, N91, N42, N63);
and AND2 (N102, N97, N19);
and AND3 (N103, N88, N20, N57);
and AND3 (N104, N96, N88, N60);
nand NAND4 (N105, N104, N47, N36, N51);
not NOT1 (N106, N61);
xor XOR2 (N107, N93, N89);
and AND4 (N108, N106, N69, N86, N51);
or OR3 (N109, N107, N65, N3);
nor NOR3 (N110, N108, N23, N106);
or OR3 (N111, N98, N104, N29);
and AND4 (N112, N111, N80, N47, N20);
and AND4 (N113, N100, N17, N18, N11);
buf BUF1 (N114, N105);
not NOT1 (N115, N113);
nor NOR3 (N116, N102, N57, N75);
not NOT1 (N117, N116);
nor NOR2 (N118, N92, N31);
nor NOR3 (N119, N99, N29, N70);
nor NOR4 (N120, N117, N22, N112, N103);
nand NAND3 (N121, N75, N49, N26);
and AND4 (N122, N102, N117, N62, N120);
and AND3 (N123, N37, N87, N83);
xor XOR2 (N124, N119, N93);
nor NOR2 (N125, N115, N27);
buf BUF1 (N126, N118);
xor XOR2 (N127, N101, N117);
and AND4 (N128, N126, N75, N100, N51);
and AND4 (N129, N114, N97, N86, N89);
nor NOR2 (N130, N125, N49);
or OR4 (N131, N129, N74, N28, N48);
or OR4 (N132, N109, N45, N6, N86);
xor XOR2 (N133, N132, N24);
xor XOR2 (N134, N127, N61);
not NOT1 (N135, N123);
or OR4 (N136, N128, N91, N5, N51);
and AND4 (N137, N136, N13, N64, N132);
nand NAND4 (N138, N122, N11, N12, N81);
buf BUF1 (N139, N133);
not NOT1 (N140, N135);
xor XOR2 (N141, N139, N102);
nor NOR4 (N142, N124, N23, N22, N51);
or OR3 (N143, N121, N136, N47);
nor NOR4 (N144, N142, N120, N134, N140);
buf BUF1 (N145, N7);
nor NOR3 (N146, N80, N143, N25);
nand NAND2 (N147, N86, N110);
nand NAND2 (N148, N25, N147);
and AND3 (N149, N17, N52, N57);
xor XOR2 (N150, N131, N135);
nand NAND2 (N151, N149, N22);
and AND4 (N152, N148, N74, N144, N120);
buf BUF1 (N153, N60);
and AND3 (N154, N150, N120, N29);
xor XOR2 (N155, N152, N57);
or OR4 (N156, N145, N55, N130, N3);
and AND3 (N157, N17, N67, N74);
or OR3 (N158, N154, N96, N135);
nor NOR4 (N159, N153, N92, N145, N104);
nand NAND3 (N160, N155, N74, N133);
nand NAND3 (N161, N159, N22, N74);
not NOT1 (N162, N146);
or OR3 (N163, N137, N127, N114);
buf BUF1 (N164, N141);
and AND3 (N165, N161, N5, N129);
buf BUF1 (N166, N156);
nor NOR2 (N167, N158, N164);
xor XOR2 (N168, N128, N117);
xor XOR2 (N169, N162, N94);
xor XOR2 (N170, N163, N13);
xor XOR2 (N171, N165, N170);
or OR3 (N172, N157, N41, N160);
nand NAND4 (N173, N151, N64, N134, N149);
nor NOR2 (N174, N48, N105);
and AND3 (N175, N50, N128, N30);
and AND4 (N176, N169, N140, N7, N72);
nand NAND2 (N177, N173, N92);
or OR3 (N178, N176, N39, N38);
nand NAND4 (N179, N172, N71, N38, N147);
and AND2 (N180, N178, N135);
buf BUF1 (N181, N179);
and AND3 (N182, N175, N179, N156);
nand NAND2 (N183, N174, N148);
and AND2 (N184, N183, N101);
or OR2 (N185, N182, N132);
buf BUF1 (N186, N167);
and AND3 (N187, N138, N127, N185);
not NOT1 (N188, N11);
or OR2 (N189, N180, N131);
not NOT1 (N190, N188);
buf BUF1 (N191, N177);
xor XOR2 (N192, N187, N145);
buf BUF1 (N193, N192);
or OR2 (N194, N193, N154);
xor XOR2 (N195, N171, N40);
buf BUF1 (N196, N168);
or OR4 (N197, N191, N101, N139, N116);
and AND3 (N198, N197, N126, N187);
xor XOR2 (N199, N195, N53);
xor XOR2 (N200, N190, N137);
nor NOR4 (N201, N166, N81, N59, N42);
xor XOR2 (N202, N201, N108);
buf BUF1 (N203, N186);
nor NOR3 (N204, N198, N164, N62);
nand NAND2 (N205, N181, N138);
not NOT1 (N206, N196);
not NOT1 (N207, N189);
or OR4 (N208, N207, N61, N128, N23);
not NOT1 (N209, N203);
or OR2 (N210, N184, N108);
and AND2 (N211, N210, N153);
buf BUF1 (N212, N200);
xor XOR2 (N213, N199, N110);
and AND4 (N214, N206, N106, N59, N67);
and AND3 (N215, N204, N146, N213);
xor XOR2 (N216, N134, N174);
or OR2 (N217, N208, N186);
buf BUF1 (N218, N216);
buf BUF1 (N219, N209);
xor XOR2 (N220, N202, N123);
nand NAND2 (N221, N218, N58);
nand NAND4 (N222, N221, N37, N109, N191);
nand NAND3 (N223, N219, N101, N158);
nand NAND2 (N224, N215, N206);
buf BUF1 (N225, N222);
nor NOR2 (N226, N223, N41);
and AND3 (N227, N217, N222, N113);
nand NAND3 (N228, N214, N205, N81);
xor XOR2 (N229, N179, N138);
nand NAND3 (N230, N225, N101, N52);
not NOT1 (N231, N230);
nand NAND4 (N232, N226, N50, N229, N47);
and AND3 (N233, N13, N190, N166);
nor NOR2 (N234, N231, N167);
not NOT1 (N235, N233);
nor NOR2 (N236, N212, N54);
buf BUF1 (N237, N227);
nand NAND3 (N238, N235, N186, N108);
xor XOR2 (N239, N194, N187);
nand NAND4 (N240, N220, N83, N222, N71);
buf BUF1 (N241, N238);
nand NAND4 (N242, N241, N63, N144, N33);
nand NAND2 (N243, N240, N184);
or OR3 (N244, N236, N201, N180);
not NOT1 (N245, N211);
nor NOR4 (N246, N234, N110, N186, N237);
and AND3 (N247, N166, N87, N182);
nand NAND3 (N248, N244, N209, N147);
not NOT1 (N249, N242);
and AND2 (N250, N228, N41);
buf BUF1 (N251, N248);
and AND2 (N252, N243, N126);
buf BUF1 (N253, N252);
or OR2 (N254, N249, N77);
buf BUF1 (N255, N253);
not NOT1 (N256, N224);
xor XOR2 (N257, N232, N115);
or OR3 (N258, N245, N193, N112);
not NOT1 (N259, N246);
xor XOR2 (N260, N239, N252);
nand NAND4 (N261, N259, N73, N92, N137);
xor XOR2 (N262, N254, N192);
and AND2 (N263, N250, N36);
and AND4 (N264, N247, N177, N2, N55);
xor XOR2 (N265, N261, N130);
buf BUF1 (N266, N251);
not NOT1 (N267, N265);
and AND3 (N268, N258, N10, N124);
nor NOR4 (N269, N264, N229, N207, N211);
buf BUF1 (N270, N260);
buf BUF1 (N271, N263);
buf BUF1 (N272, N268);
nor NOR4 (N273, N266, N177, N180, N227);
not NOT1 (N274, N267);
nand NAND2 (N275, N255, N125);
xor XOR2 (N276, N272, N88);
not NOT1 (N277, N262);
nor NOR4 (N278, N270, N138, N230, N137);
nand NAND3 (N279, N275, N17, N214);
and AND2 (N280, N279, N120);
not NOT1 (N281, N269);
not NOT1 (N282, N274);
or OR2 (N283, N276, N136);
or OR4 (N284, N256, N130, N260, N97);
nand NAND4 (N285, N280, N278, N5, N29);
buf BUF1 (N286, N141);
buf BUF1 (N287, N286);
and AND2 (N288, N257, N112);
and AND3 (N289, N271, N12, N21);
not NOT1 (N290, N289);
buf BUF1 (N291, N285);
nand NAND3 (N292, N284, N106, N196);
buf BUF1 (N293, N291);
and AND4 (N294, N281, N129, N44, N36);
or OR2 (N295, N273, N84);
not NOT1 (N296, N283);
not NOT1 (N297, N282);
and AND3 (N298, N296, N86, N6);
not NOT1 (N299, N293);
not NOT1 (N300, N292);
not NOT1 (N301, N277);
xor XOR2 (N302, N297, N182);
buf BUF1 (N303, N300);
and AND3 (N304, N303, N17, N105);
or OR3 (N305, N287, N173, N300);
nand NAND4 (N306, N290, N196, N246, N53);
nor NOR2 (N307, N298, N27);
buf BUF1 (N308, N304);
nor NOR4 (N309, N294, N60, N45, N172);
or OR3 (N310, N299, N151, N146);
not NOT1 (N311, N288);
and AND2 (N312, N295, N116);
nor NOR2 (N313, N312, N210);
and AND4 (N314, N310, N37, N160, N68);
nor NOR2 (N315, N314, N70);
or OR4 (N316, N308, N181, N185, N29);
xor XOR2 (N317, N307, N83);
nor NOR2 (N318, N313, N211);
buf BUF1 (N319, N318);
buf BUF1 (N320, N319);
buf BUF1 (N321, N320);
nand NAND2 (N322, N316, N64);
nand NAND2 (N323, N309, N277);
not NOT1 (N324, N321);
buf BUF1 (N325, N323);
and AND3 (N326, N311, N123, N77);
or OR4 (N327, N322, N250, N288, N228);
not NOT1 (N328, N301);
not NOT1 (N329, N325);
or OR4 (N330, N328, N316, N268, N181);
and AND3 (N331, N324, N150, N143);
buf BUF1 (N332, N315);
or OR2 (N333, N330, N165);
nand NAND3 (N334, N317, N67, N87);
not NOT1 (N335, N333);
and AND2 (N336, N306, N96);
nand NAND4 (N337, N326, N322, N265, N208);
not NOT1 (N338, N302);
nand NAND4 (N339, N337, N265, N205, N153);
xor XOR2 (N340, N335, N290);
not NOT1 (N341, N339);
nand NAND4 (N342, N338, N77, N163, N70);
nand NAND3 (N343, N329, N307, N147);
and AND3 (N344, N340, N299, N51);
nor NOR2 (N345, N305, N338);
xor XOR2 (N346, N332, N149);
buf BUF1 (N347, N343);
not NOT1 (N348, N334);
or OR3 (N349, N331, N152, N175);
nor NOR2 (N350, N347, N116);
and AND3 (N351, N342, N246, N73);
nand NAND2 (N352, N327, N91);
buf BUF1 (N353, N350);
nand NAND4 (N354, N341, N258, N138, N258);
buf BUF1 (N355, N336);
nand NAND2 (N356, N353, N228);
nor NOR2 (N357, N348, N233);
nand NAND3 (N358, N355, N176, N54);
buf BUF1 (N359, N352);
or OR4 (N360, N349, N239, N214, N213);
or OR3 (N361, N345, N152, N272);
nand NAND4 (N362, N344, N60, N285, N355);
or OR3 (N363, N357, N108, N345);
or OR2 (N364, N360, N341);
nor NOR3 (N365, N354, N121, N295);
or OR2 (N366, N359, N97);
not NOT1 (N367, N366);
and AND4 (N368, N361, N366, N33, N153);
not NOT1 (N369, N363);
not NOT1 (N370, N364);
or OR3 (N371, N351, N109, N64);
buf BUF1 (N372, N356);
xor XOR2 (N373, N358, N171);
xor XOR2 (N374, N369, N291);
nand NAND2 (N375, N374, N14);
and AND3 (N376, N346, N193, N161);
nor NOR3 (N377, N370, N210, N129);
and AND4 (N378, N362, N202, N239, N321);
nor NOR4 (N379, N365, N102, N103, N212);
xor XOR2 (N380, N375, N57);
buf BUF1 (N381, N371);
xor XOR2 (N382, N372, N332);
nand NAND3 (N383, N380, N182, N66);
not NOT1 (N384, N381);
xor XOR2 (N385, N373, N37);
xor XOR2 (N386, N376, N159);
xor XOR2 (N387, N368, N255);
nor NOR4 (N388, N384, N231, N292, N78);
not NOT1 (N389, N385);
and AND2 (N390, N382, N104);
not NOT1 (N391, N390);
and AND2 (N392, N387, N204);
buf BUF1 (N393, N391);
buf BUF1 (N394, N379);
buf BUF1 (N395, N394);
xor XOR2 (N396, N377, N290);
not NOT1 (N397, N386);
nand NAND3 (N398, N388, N311, N70);
or OR4 (N399, N393, N323, N176, N258);
buf BUF1 (N400, N395);
xor XOR2 (N401, N383, N400);
xor XOR2 (N402, N212, N333);
xor XOR2 (N403, N367, N268);
not NOT1 (N404, N402);
and AND3 (N405, N401, N283, N287);
not NOT1 (N406, N396);
buf BUF1 (N407, N397);
nand NAND3 (N408, N389, N219, N338);
nor NOR3 (N409, N403, N123, N170);
buf BUF1 (N410, N392);
buf BUF1 (N411, N410);
xor XOR2 (N412, N411, N84);
or OR2 (N413, N405, N361);
and AND3 (N414, N406, N265, N107);
buf BUF1 (N415, N407);
xor XOR2 (N416, N414, N383);
and AND2 (N417, N416, N216);
nor NOR3 (N418, N417, N264, N327);
not NOT1 (N419, N418);
nor NOR3 (N420, N413, N73, N356);
xor XOR2 (N421, N412, N85);
or OR2 (N422, N408, N341);
buf BUF1 (N423, N421);
xor XOR2 (N424, N409, N316);
and AND2 (N425, N404, N131);
xor XOR2 (N426, N415, N70);
and AND4 (N427, N422, N115, N425, N282);
buf BUF1 (N428, N223);
buf BUF1 (N429, N424);
xor XOR2 (N430, N378, N359);
nor NOR3 (N431, N423, N325, N34);
not NOT1 (N432, N428);
xor XOR2 (N433, N429, N78);
nand NAND3 (N434, N420, N195, N247);
or OR2 (N435, N434, N96);
nand NAND2 (N436, N431, N117);
nand NAND2 (N437, N432, N293);
buf BUF1 (N438, N433);
xor XOR2 (N439, N399, N335);
xor XOR2 (N440, N398, N193);
or OR3 (N441, N435, N164, N185);
buf BUF1 (N442, N419);
buf BUF1 (N443, N437);
buf BUF1 (N444, N442);
nand NAND2 (N445, N430, N69);
xor XOR2 (N446, N438, N423);
xor XOR2 (N447, N443, N196);
buf BUF1 (N448, N436);
xor XOR2 (N449, N439, N398);
buf BUF1 (N450, N440);
xor XOR2 (N451, N427, N301);
or OR3 (N452, N426, N407, N126);
xor XOR2 (N453, N445, N68);
nand NAND2 (N454, N447, N279);
xor XOR2 (N455, N449, N136);
not NOT1 (N456, N450);
and AND4 (N457, N446, N137, N101, N344);
nand NAND3 (N458, N456, N191, N231);
buf BUF1 (N459, N448);
buf BUF1 (N460, N458);
nor NOR3 (N461, N444, N165, N321);
not NOT1 (N462, N460);
nand NAND2 (N463, N454, N330);
buf BUF1 (N464, N457);
or OR3 (N465, N459, N16, N299);
xor XOR2 (N466, N455, N426);
buf BUF1 (N467, N463);
nand NAND2 (N468, N462, N388);
buf BUF1 (N469, N465);
buf BUF1 (N470, N453);
buf BUF1 (N471, N466);
not NOT1 (N472, N468);
not NOT1 (N473, N469);
nor NOR4 (N474, N470, N425, N369, N342);
nor NOR2 (N475, N464, N161);
nand NAND4 (N476, N452, N323, N293, N150);
nor NOR4 (N477, N474, N422, N295, N453);
or OR2 (N478, N471, N111);
or OR3 (N479, N476, N36, N305);
nand NAND3 (N480, N473, N25, N238);
not NOT1 (N481, N479);
xor XOR2 (N482, N461, N446);
and AND2 (N483, N475, N136);
nand NAND2 (N484, N467, N474);
buf BUF1 (N485, N480);
buf BUF1 (N486, N481);
buf BUF1 (N487, N484);
xor XOR2 (N488, N485, N129);
not NOT1 (N489, N487);
nor NOR2 (N490, N483, N31);
xor XOR2 (N491, N441, N323);
nand NAND2 (N492, N482, N52);
and AND4 (N493, N478, N265, N68, N16);
nor NOR3 (N494, N492, N394, N243);
and AND3 (N495, N451, N377, N6);
buf BUF1 (N496, N490);
nor NOR4 (N497, N496, N40, N478, N169);
and AND4 (N498, N489, N282, N236, N276);
nor NOR4 (N499, N498, N8, N49, N221);
and AND3 (N500, N491, N295, N5);
nor NOR2 (N501, N499, N132);
not NOT1 (N502, N486);
nand NAND2 (N503, N497, N117);
xor XOR2 (N504, N503, N59);
or OR3 (N505, N495, N366, N208);
buf BUF1 (N506, N488);
nand NAND2 (N507, N494, N257);
not NOT1 (N508, N505);
buf BUF1 (N509, N493);
or OR3 (N510, N504, N11, N265);
nand NAND4 (N511, N507, N159, N456, N155);
xor XOR2 (N512, N511, N480);
xor XOR2 (N513, N500, N352);
xor XOR2 (N514, N512, N235);
nor NOR4 (N515, N472, N492, N67, N398);
not NOT1 (N516, N508);
not NOT1 (N517, N502);
xor XOR2 (N518, N513, N103);
nand NAND3 (N519, N506, N463, N422);
not NOT1 (N520, N517);
and AND3 (N521, N510, N247, N116);
buf BUF1 (N522, N509);
not NOT1 (N523, N519);
xor XOR2 (N524, N477, N334);
xor XOR2 (N525, N501, N279);
not NOT1 (N526, N521);
nor NOR3 (N527, N525, N77, N400);
nor NOR3 (N528, N527, N170, N464);
not NOT1 (N529, N514);
not NOT1 (N530, N524);
not NOT1 (N531, N526);
xor XOR2 (N532, N531, N388);
nor NOR4 (N533, N518, N520, N204, N439);
xor XOR2 (N534, N399, N524);
nand NAND4 (N535, N530, N139, N194, N445);
and AND2 (N536, N534, N156);
nand NAND3 (N537, N515, N480, N172);
nand NAND4 (N538, N532, N238, N453, N130);
nand NAND2 (N539, N522, N150);
nand NAND2 (N540, N538, N524);
buf BUF1 (N541, N540);
not NOT1 (N542, N528);
nor NOR4 (N543, N536, N5, N265, N286);
or OR3 (N544, N541, N153, N246);
or OR4 (N545, N529, N388, N353, N500);
nand NAND2 (N546, N545, N269);
nand NAND2 (N547, N535, N220);
xor XOR2 (N548, N542, N293);
nor NOR3 (N549, N547, N463, N453);
nor NOR4 (N550, N544, N161, N450, N520);
buf BUF1 (N551, N523);
nor NOR4 (N552, N516, N28, N351, N205);
xor XOR2 (N553, N543, N435);
nor NOR3 (N554, N549, N342, N483);
buf BUF1 (N555, N539);
xor XOR2 (N556, N554, N511);
xor XOR2 (N557, N548, N253);
xor XOR2 (N558, N550, N176);
nor NOR2 (N559, N533, N231);
nor NOR4 (N560, N558, N559, N388, N485);
xor XOR2 (N561, N551, N546);
not NOT1 (N562, N419);
nand NAND2 (N563, N49, N369);
nand NAND4 (N564, N563, N509, N101, N417);
nand NAND3 (N565, N557, N372, N124);
or OR4 (N566, N537, N264, N299, N278);
or OR3 (N567, N564, N539, N503);
nor NOR2 (N568, N561, N501);
not NOT1 (N569, N556);
not NOT1 (N570, N567);
buf BUF1 (N571, N562);
and AND2 (N572, N553, N433);
and AND3 (N573, N566, N105, N190);
or OR3 (N574, N560, N457, N199);
nor NOR2 (N575, N568, N453);
and AND2 (N576, N565, N47);
nor NOR2 (N577, N574, N452);
nor NOR2 (N578, N571, N342);
nor NOR4 (N579, N572, N349, N463, N115);
xor XOR2 (N580, N555, N333);
nand NAND3 (N581, N570, N466, N347);
and AND2 (N582, N581, N522);
xor XOR2 (N583, N578, N326);
and AND2 (N584, N575, N172);
or OR3 (N585, N584, N417, N93);
not NOT1 (N586, N585);
not NOT1 (N587, N580);
buf BUF1 (N588, N582);
nand NAND2 (N589, N583, N249);
xor XOR2 (N590, N552, N160);
not NOT1 (N591, N573);
or OR3 (N592, N569, N463, N202);
nand NAND4 (N593, N589, N261, N577, N376);
nor NOR3 (N594, N419, N230, N5);
xor XOR2 (N595, N586, N383);
nand NAND4 (N596, N594, N208, N277, N100);
nand NAND2 (N597, N595, N552);
xor XOR2 (N598, N579, N472);
or OR4 (N599, N590, N416, N111, N43);
nand NAND4 (N600, N599, N58, N10, N418);
nor NOR3 (N601, N596, N517, N375);
or OR4 (N602, N576, N392, N248, N303);
buf BUF1 (N603, N602);
and AND4 (N604, N587, N120, N81, N70);
nor NOR4 (N605, N603, N209, N533, N256);
nor NOR2 (N606, N588, N570);
not NOT1 (N607, N593);
and AND4 (N608, N597, N365, N215, N447);
buf BUF1 (N609, N600);
nand NAND4 (N610, N591, N387, N243, N413);
nand NAND2 (N611, N605, N147);
or OR3 (N612, N598, N52, N465);
and AND2 (N613, N604, N405);
not NOT1 (N614, N606);
and AND2 (N615, N614, N341);
or OR4 (N616, N615, N294, N570, N461);
buf BUF1 (N617, N609);
xor XOR2 (N618, N616, N206);
and AND4 (N619, N613, N579, N498, N475);
buf BUF1 (N620, N608);
nand NAND3 (N621, N607, N15, N222);
or OR3 (N622, N621, N272, N604);
buf BUF1 (N623, N619);
or OR4 (N624, N601, N303, N434, N181);
and AND2 (N625, N612, N494);
nor NOR3 (N626, N610, N450, N223);
not NOT1 (N627, N620);
buf BUF1 (N628, N625);
and AND4 (N629, N626, N132, N193, N336);
or OR2 (N630, N623, N106);
xor XOR2 (N631, N611, N449);
xor XOR2 (N632, N592, N538);
buf BUF1 (N633, N632);
or OR3 (N634, N617, N304, N144);
not NOT1 (N635, N629);
buf BUF1 (N636, N618);
nand NAND3 (N637, N631, N286, N85);
and AND4 (N638, N630, N622, N580, N58);
and AND4 (N639, N494, N466, N164, N74);
not NOT1 (N640, N638);
or OR3 (N641, N627, N25, N490);
and AND2 (N642, N635, N29);
buf BUF1 (N643, N641);
buf BUF1 (N644, N633);
nand NAND4 (N645, N643, N493, N213, N302);
not NOT1 (N646, N639);
and AND4 (N647, N634, N426, N622, N641);
nor NOR2 (N648, N647, N119);
buf BUF1 (N649, N642);
not NOT1 (N650, N640);
nor NOR2 (N651, N636, N249);
or OR4 (N652, N645, N606, N326, N208);
xor XOR2 (N653, N644, N254);
buf BUF1 (N654, N651);
or OR2 (N655, N650, N72);
nor NOR3 (N656, N628, N45, N244);
or OR3 (N657, N648, N656, N256);
buf BUF1 (N658, N204);
nor NOR2 (N659, N654, N20);
nand NAND4 (N660, N637, N588, N97, N633);
and AND3 (N661, N659, N271, N368);
or OR4 (N662, N658, N432, N521, N638);
buf BUF1 (N663, N660);
buf BUF1 (N664, N655);
or OR2 (N665, N646, N293);
buf BUF1 (N666, N665);
nor NOR2 (N667, N649, N104);
nand NAND2 (N668, N667, N435);
buf BUF1 (N669, N668);
not NOT1 (N670, N661);
buf BUF1 (N671, N653);
nand NAND3 (N672, N663, N327, N480);
buf BUF1 (N673, N666);
xor XOR2 (N674, N673, N428);
nor NOR3 (N675, N662, N204, N607);
xor XOR2 (N676, N664, N259);
nand NAND2 (N677, N652, N579);
and AND2 (N678, N676, N181);
or OR4 (N679, N678, N146, N636, N592);
xor XOR2 (N680, N671, N501);
buf BUF1 (N681, N624);
xor XOR2 (N682, N670, N366);
xor XOR2 (N683, N681, N202);
xor XOR2 (N684, N669, N568);
nor NOR4 (N685, N674, N290, N31, N574);
and AND3 (N686, N680, N328, N95);
buf BUF1 (N687, N672);
xor XOR2 (N688, N677, N234);
or OR2 (N689, N688, N257);
nor NOR2 (N690, N682, N370);
xor XOR2 (N691, N679, N520);
or OR4 (N692, N687, N123, N36, N49);
nor NOR4 (N693, N684, N412, N205, N341);
nand NAND4 (N694, N693, N677, N449, N629);
buf BUF1 (N695, N690);
nand NAND2 (N696, N683, N514);
xor XOR2 (N697, N686, N480);
nor NOR2 (N698, N685, N496);
nor NOR3 (N699, N675, N655, N673);
not NOT1 (N700, N698);
nor NOR2 (N701, N689, N341);
nor NOR3 (N702, N700, N134, N607);
or OR3 (N703, N701, N658, N274);
and AND3 (N704, N692, N692, N227);
or OR4 (N705, N703, N613, N668, N591);
and AND4 (N706, N704, N702, N648, N313);
nor NOR3 (N707, N68, N644, N371);
or OR4 (N708, N697, N552, N154, N107);
xor XOR2 (N709, N707, N396);
or OR2 (N710, N706, N534);
and AND2 (N711, N709, N247);
nor NOR2 (N712, N657, N155);
xor XOR2 (N713, N694, N555);
or OR2 (N714, N710, N649);
not NOT1 (N715, N695);
nand NAND2 (N716, N712, N441);
nor NOR2 (N717, N708, N406);
nand NAND4 (N718, N711, N247, N459, N630);
not NOT1 (N719, N716);
or OR4 (N720, N715, N275, N366, N647);
xor XOR2 (N721, N717, N365);
buf BUF1 (N722, N721);
and AND3 (N723, N718, N292, N428);
nor NOR3 (N724, N696, N100, N490);
nor NOR2 (N725, N719, N585);
buf BUF1 (N726, N714);
or OR3 (N727, N722, N80, N683);
xor XOR2 (N728, N726, N164);
and AND3 (N729, N725, N489, N16);
nor NOR3 (N730, N705, N361, N121);
or OR4 (N731, N699, N52, N704, N609);
nand NAND2 (N732, N729, N211);
xor XOR2 (N733, N731, N313);
nor NOR2 (N734, N733, N517);
or OR3 (N735, N691, N387, N321);
and AND3 (N736, N732, N209, N625);
not NOT1 (N737, N720);
not NOT1 (N738, N713);
nand NAND4 (N739, N723, N320, N302, N242);
xor XOR2 (N740, N724, N412);
not NOT1 (N741, N727);
xor XOR2 (N742, N740, N105);
buf BUF1 (N743, N739);
and AND2 (N744, N738, N468);
not NOT1 (N745, N744);
not NOT1 (N746, N743);
buf BUF1 (N747, N735);
and AND2 (N748, N741, N350);
xor XOR2 (N749, N748, N659);
nor NOR3 (N750, N737, N190, N419);
and AND4 (N751, N750, N346, N321, N693);
not NOT1 (N752, N749);
buf BUF1 (N753, N734);
nand NAND4 (N754, N742, N35, N664, N349);
or OR4 (N755, N752, N10, N585, N137);
or OR4 (N756, N747, N553, N606, N210);
not NOT1 (N757, N728);
nor NOR4 (N758, N753, N190, N16, N544);
buf BUF1 (N759, N758);
or OR3 (N760, N746, N562, N130);
xor XOR2 (N761, N751, N506);
buf BUF1 (N762, N736);
and AND3 (N763, N757, N150, N430);
nor NOR4 (N764, N745, N221, N593, N155);
nor NOR2 (N765, N756, N365);
xor XOR2 (N766, N762, N324);
not NOT1 (N767, N766);
nand NAND2 (N768, N764, N590);
not NOT1 (N769, N767);
buf BUF1 (N770, N755);
and AND2 (N771, N768, N468);
not NOT1 (N772, N761);
xor XOR2 (N773, N763, N507);
buf BUF1 (N774, N765);
buf BUF1 (N775, N773);
not NOT1 (N776, N759);
nand NAND4 (N777, N770, N548, N21, N611);
xor XOR2 (N778, N769, N687);
buf BUF1 (N779, N754);
or OR2 (N780, N779, N323);
not NOT1 (N781, N774);
nand NAND4 (N782, N780, N749, N404, N567);
buf BUF1 (N783, N772);
nor NOR3 (N784, N778, N153, N709);
buf BUF1 (N785, N775);
nor NOR4 (N786, N776, N742, N194, N782);
not NOT1 (N787, N462);
and AND3 (N788, N787, N392, N524);
buf BUF1 (N789, N783);
not NOT1 (N790, N730);
or OR3 (N791, N785, N63, N417);
xor XOR2 (N792, N784, N303);
or OR3 (N793, N781, N390, N62);
nand NAND2 (N794, N786, N573);
xor XOR2 (N795, N760, N304);
and AND2 (N796, N771, N574);
xor XOR2 (N797, N792, N746);
or OR3 (N798, N791, N126, N558);
and AND2 (N799, N795, N536);
or OR3 (N800, N797, N237, N62);
xor XOR2 (N801, N796, N680);
nor NOR2 (N802, N790, N691);
buf BUF1 (N803, N777);
not NOT1 (N804, N788);
xor XOR2 (N805, N799, N585);
buf BUF1 (N806, N804);
nor NOR4 (N807, N800, N694, N83, N615);
buf BUF1 (N808, N806);
or OR2 (N809, N805, N738);
nand NAND4 (N810, N801, N648, N253, N314);
or OR3 (N811, N808, N190, N299);
or OR2 (N812, N803, N769);
nand NAND3 (N813, N793, N591, N214);
not NOT1 (N814, N809);
not NOT1 (N815, N812);
and AND2 (N816, N798, N526);
nor NOR4 (N817, N794, N444, N194, N735);
xor XOR2 (N818, N817, N674);
not NOT1 (N819, N807);
not NOT1 (N820, N819);
and AND4 (N821, N820, N435, N381, N326);
xor XOR2 (N822, N818, N430);
xor XOR2 (N823, N811, N740);
or OR4 (N824, N810, N23, N493, N556);
buf BUF1 (N825, N821);
xor XOR2 (N826, N813, N442);
nor NOR3 (N827, N826, N756, N8);
and AND2 (N828, N802, N662);
buf BUF1 (N829, N816);
buf BUF1 (N830, N828);
nor NOR2 (N831, N829, N227);
nor NOR2 (N832, N827, N334);
or OR2 (N833, N823, N796);
xor XOR2 (N834, N825, N520);
or OR4 (N835, N834, N710, N161, N144);
or OR2 (N836, N832, N1);
buf BUF1 (N837, N789);
and AND2 (N838, N837, N62);
not NOT1 (N839, N815);
nor NOR2 (N840, N822, N204);
not NOT1 (N841, N831);
buf BUF1 (N842, N836);
nand NAND2 (N843, N835, N354);
buf BUF1 (N844, N839);
not NOT1 (N845, N824);
xor XOR2 (N846, N833, N688);
not NOT1 (N847, N846);
and AND2 (N848, N841, N288);
not NOT1 (N849, N845);
nor NOR3 (N850, N849, N755, N634);
nor NOR2 (N851, N814, N66);
nor NOR3 (N852, N838, N455, N536);
nand NAND4 (N853, N844, N106, N801, N402);
buf BUF1 (N854, N843);
not NOT1 (N855, N851);
or OR2 (N856, N854, N209);
and AND4 (N857, N840, N88, N109, N339);
xor XOR2 (N858, N830, N317);
nand NAND3 (N859, N858, N79, N656);
xor XOR2 (N860, N847, N612);
not NOT1 (N861, N848);
not NOT1 (N862, N857);
buf BUF1 (N863, N861);
or OR4 (N864, N859, N145, N574, N722);
xor XOR2 (N865, N856, N145);
nand NAND3 (N866, N860, N763, N26);
nor NOR3 (N867, N865, N537, N802);
xor XOR2 (N868, N852, N222);
not NOT1 (N869, N866);
xor XOR2 (N870, N855, N207);
nor NOR4 (N871, N864, N342, N449, N292);
not NOT1 (N872, N868);
nand NAND2 (N873, N853, N823);
nor NOR4 (N874, N850, N866, N864, N47);
not NOT1 (N875, N863);
and AND4 (N876, N875, N738, N437, N509);
nand NAND2 (N877, N842, N818);
nand NAND4 (N878, N869, N335, N474, N26);
buf BUF1 (N879, N870);
not NOT1 (N880, N879);
or OR4 (N881, N877, N255, N499, N310);
and AND3 (N882, N874, N475, N477);
xor XOR2 (N883, N881, N735);
nor NOR2 (N884, N878, N297);
nor NOR3 (N885, N873, N49, N769);
not NOT1 (N886, N872);
xor XOR2 (N887, N885, N822);
xor XOR2 (N888, N884, N292);
or OR3 (N889, N888, N597, N14);
nor NOR3 (N890, N889, N412, N378);
xor XOR2 (N891, N883, N818);
buf BUF1 (N892, N876);
xor XOR2 (N893, N890, N143);
buf BUF1 (N894, N862);
and AND2 (N895, N871, N548);
or OR4 (N896, N895, N887, N788, N406);
or OR3 (N897, N368, N45, N4);
nor NOR2 (N898, N893, N445);
or OR2 (N899, N896, N449);
and AND3 (N900, N894, N854, N691);
xor XOR2 (N901, N897, N22);
not NOT1 (N902, N882);
not NOT1 (N903, N899);
nand NAND3 (N904, N891, N175, N749);
not NOT1 (N905, N900);
or OR3 (N906, N867, N615, N449);
not NOT1 (N907, N892);
buf BUF1 (N908, N903);
xor XOR2 (N909, N904, N726);
nor NOR2 (N910, N907, N806);
or OR2 (N911, N901, N548);
buf BUF1 (N912, N911);
and AND2 (N913, N906, N870);
not NOT1 (N914, N912);
not NOT1 (N915, N886);
nor NOR4 (N916, N910, N332, N378, N656);
not NOT1 (N917, N908);
or OR2 (N918, N917, N595);
nor NOR3 (N919, N915, N452, N542);
and AND2 (N920, N913, N326);
buf BUF1 (N921, N918);
and AND4 (N922, N920, N275, N517, N339);
or OR3 (N923, N902, N395, N801);
or OR2 (N924, N923, N558);
nor NOR4 (N925, N905, N366, N637, N880);
or OR2 (N926, N66, N536);
not NOT1 (N927, N914);
xor XOR2 (N928, N898, N712);
not NOT1 (N929, N925);
xor XOR2 (N930, N919, N891);
nand NAND2 (N931, N930, N413);
buf BUF1 (N932, N928);
and AND2 (N933, N921, N860);
not NOT1 (N934, N931);
xor XOR2 (N935, N932, N281);
not NOT1 (N936, N935);
or OR4 (N937, N936, N246, N746, N168);
nand NAND2 (N938, N934, N635);
nor NOR4 (N939, N929, N16, N36, N354);
or OR3 (N940, N933, N890, N324);
nor NOR2 (N941, N922, N626);
not NOT1 (N942, N927);
nor NOR3 (N943, N940, N898, N765);
nand NAND4 (N944, N926, N729, N499, N40);
nor NOR2 (N945, N942, N70);
buf BUF1 (N946, N916);
or OR3 (N947, N938, N799, N388);
or OR2 (N948, N943, N783);
buf BUF1 (N949, N909);
nand NAND4 (N950, N939, N552, N625, N330);
not NOT1 (N951, N937);
not NOT1 (N952, N924);
and AND4 (N953, N950, N781, N664, N100);
nand NAND2 (N954, N948, N698);
nor NOR4 (N955, N952, N773, N338, N931);
and AND3 (N956, N946, N524, N203);
not NOT1 (N957, N944);
xor XOR2 (N958, N955, N930);
nor NOR4 (N959, N953, N224, N89, N163);
nand NAND2 (N960, N954, N886);
or OR3 (N961, N949, N21, N235);
not NOT1 (N962, N941);
and AND2 (N963, N951, N221);
or OR2 (N964, N960, N748);
not NOT1 (N965, N956);
nor NOR2 (N966, N945, N873);
nor NOR4 (N967, N965, N495, N591, N805);
not NOT1 (N968, N963);
xor XOR2 (N969, N964, N615);
or OR2 (N970, N967, N532);
buf BUF1 (N971, N957);
and AND4 (N972, N968, N359, N149, N900);
and AND3 (N973, N970, N635, N681);
not NOT1 (N974, N962);
and AND3 (N975, N959, N407, N354);
buf BUF1 (N976, N973);
or OR4 (N977, N971, N215, N251, N749);
and AND2 (N978, N977, N554);
nor NOR2 (N979, N975, N618);
not NOT1 (N980, N978);
not NOT1 (N981, N974);
nor NOR4 (N982, N972, N844, N306, N459);
or OR3 (N983, N947, N56, N605);
or OR3 (N984, N976, N669, N128);
nor NOR4 (N985, N980, N926, N526, N695);
not NOT1 (N986, N958);
or OR3 (N987, N961, N403, N771);
xor XOR2 (N988, N969, N496);
buf BUF1 (N989, N982);
xor XOR2 (N990, N979, N112);
not NOT1 (N991, N966);
xor XOR2 (N992, N983, N717);
xor XOR2 (N993, N987, N122);
xor XOR2 (N994, N986, N53);
not NOT1 (N995, N984);
and AND4 (N996, N992, N589, N905, N220);
or OR2 (N997, N994, N147);
not NOT1 (N998, N991);
xor XOR2 (N999, N997, N533);
and AND4 (N1000, N993, N290, N26, N678);
buf BUF1 (N1001, N995);
not NOT1 (N1002, N990);
nand NAND2 (N1003, N1000, N40);
not NOT1 (N1004, N1001);
not NOT1 (N1005, N985);
nand NAND4 (N1006, N996, N440, N939, N483);
nor NOR2 (N1007, N1003, N639);
buf BUF1 (N1008, N998);
xor XOR2 (N1009, N989, N590);
buf BUF1 (N1010, N1002);
nand NAND3 (N1011, N1004, N44, N908);
nor NOR4 (N1012, N1005, N756, N519, N730);
buf BUF1 (N1013, N1009);
buf BUF1 (N1014, N1007);
xor XOR2 (N1015, N1006, N426);
nand NAND3 (N1016, N1014, N154, N27);
nor NOR3 (N1017, N1010, N321, N587);
and AND4 (N1018, N1015, N516, N356, N661);
nand NAND2 (N1019, N999, N25);
and AND2 (N1020, N1012, N977);
xor XOR2 (N1021, N1018, N112);
or OR3 (N1022, N1011, N22, N515);
not NOT1 (N1023, N1013);
not NOT1 (N1024, N1021);
xor XOR2 (N1025, N1008, N17);
buf BUF1 (N1026, N1016);
not NOT1 (N1027, N988);
or OR3 (N1028, N1026, N580, N711);
or OR4 (N1029, N1027, N444, N340, N111);
or OR2 (N1030, N1020, N441);
or OR4 (N1031, N1019, N665, N8, N426);
or OR3 (N1032, N1024, N1003, N359);
nor NOR2 (N1033, N1022, N188);
nor NOR4 (N1034, N1023, N934, N680, N234);
or OR2 (N1035, N1033, N208);
xor XOR2 (N1036, N1029, N103);
buf BUF1 (N1037, N1036);
buf BUF1 (N1038, N1037);
nand NAND3 (N1039, N1034, N889, N730);
not NOT1 (N1040, N1031);
xor XOR2 (N1041, N981, N648);
or OR4 (N1042, N1030, N635, N319, N690);
buf BUF1 (N1043, N1032);
and AND3 (N1044, N1038, N615, N496);
not NOT1 (N1045, N1025);
xor XOR2 (N1046, N1040, N41);
xor XOR2 (N1047, N1045, N370);
nor NOR2 (N1048, N1044, N387);
and AND2 (N1049, N1043, N540);
nor NOR3 (N1050, N1049, N673, N84);
nand NAND3 (N1051, N1048, N120, N306);
nand NAND3 (N1052, N1046, N159, N108);
or OR3 (N1053, N1028, N694, N135);
nor NOR3 (N1054, N1050, N427, N529);
and AND3 (N1055, N1047, N584, N996);
or OR2 (N1056, N1054, N384);
or OR4 (N1057, N1017, N33, N166, N406);
nand NAND4 (N1058, N1052, N384, N72, N53);
and AND3 (N1059, N1041, N134, N844);
not NOT1 (N1060, N1056);
not NOT1 (N1061, N1035);
xor XOR2 (N1062, N1058, N844);
buf BUF1 (N1063, N1042);
or OR4 (N1064, N1039, N196, N155, N307);
nand NAND4 (N1065, N1051, N137, N400, N986);
not NOT1 (N1066, N1060);
not NOT1 (N1067, N1066);
and AND4 (N1068, N1059, N601, N306, N631);
and AND4 (N1069, N1064, N519, N725, N172);
nor NOR3 (N1070, N1068, N867, N442);
not NOT1 (N1071, N1055);
buf BUF1 (N1072, N1065);
and AND2 (N1073, N1069, N204);
and AND3 (N1074, N1053, N176, N199);
nand NAND3 (N1075, N1063, N335, N870);
nand NAND2 (N1076, N1067, N335);
or OR4 (N1077, N1075, N964, N317, N206);
and AND4 (N1078, N1072, N1040, N629, N761);
not NOT1 (N1079, N1076);
nor NOR2 (N1080, N1079, N913);
nor NOR3 (N1081, N1057, N811, N495);
nor NOR4 (N1082, N1061, N20, N772, N419);
or OR3 (N1083, N1082, N403, N223);
nor NOR3 (N1084, N1077, N569, N986);
nor NOR4 (N1085, N1062, N807, N933, N42);
not NOT1 (N1086, N1074);
and AND3 (N1087, N1070, N95, N366);
xor XOR2 (N1088, N1071, N66);
and AND4 (N1089, N1084, N69, N728, N694);
nor NOR3 (N1090, N1080, N669, N219);
nor NOR4 (N1091, N1078, N1068, N466, N477);
buf BUF1 (N1092, N1087);
buf BUF1 (N1093, N1073);
xor XOR2 (N1094, N1083, N1079);
nand NAND4 (N1095, N1090, N844, N781, N587);
xor XOR2 (N1096, N1092, N508);
xor XOR2 (N1097, N1091, N147);
nor NOR4 (N1098, N1094, N886, N567, N121);
nand NAND2 (N1099, N1085, N1);
not NOT1 (N1100, N1089);
not NOT1 (N1101, N1098);
or OR2 (N1102, N1096, N560);
not NOT1 (N1103, N1093);
nand NAND3 (N1104, N1088, N296, N800);
not NOT1 (N1105, N1103);
nand NAND2 (N1106, N1105, N562);
nand NAND2 (N1107, N1099, N179);
not NOT1 (N1108, N1086);
xor XOR2 (N1109, N1106, N551);
buf BUF1 (N1110, N1107);
or OR4 (N1111, N1104, N782, N561, N644);
not NOT1 (N1112, N1110);
or OR4 (N1113, N1111, N950, N485, N620);
buf BUF1 (N1114, N1097);
nor NOR3 (N1115, N1081, N609, N321);
or OR4 (N1116, N1113, N558, N870, N604);
not NOT1 (N1117, N1095);
xor XOR2 (N1118, N1109, N356);
not NOT1 (N1119, N1112);
not NOT1 (N1120, N1116);
and AND3 (N1121, N1119, N1048, N103);
nand NAND4 (N1122, N1118, N197, N998, N350);
nor NOR4 (N1123, N1108, N75, N1015, N1084);
not NOT1 (N1124, N1100);
nor NOR4 (N1125, N1102, N1082, N501, N876);
nor NOR3 (N1126, N1117, N216, N996);
and AND3 (N1127, N1122, N735, N287);
or OR4 (N1128, N1101, N145, N303, N403);
not NOT1 (N1129, N1127);
nor NOR4 (N1130, N1124, N77, N1029, N131);
nand NAND3 (N1131, N1125, N761, N69);
buf BUF1 (N1132, N1123);
buf BUF1 (N1133, N1115);
buf BUF1 (N1134, N1130);
xor XOR2 (N1135, N1129, N773);
or OR2 (N1136, N1135, N708);
xor XOR2 (N1137, N1120, N862);
or OR4 (N1138, N1134, N997, N979, N155);
and AND3 (N1139, N1136, N64, N1064);
xor XOR2 (N1140, N1133, N201);
or OR2 (N1141, N1121, N429);
and AND3 (N1142, N1139, N291, N670);
and AND4 (N1143, N1126, N470, N835, N376);
nand NAND4 (N1144, N1143, N595, N494, N1001);
not NOT1 (N1145, N1144);
xor XOR2 (N1146, N1145, N20);
buf BUF1 (N1147, N1131);
or OR3 (N1148, N1132, N569, N724);
and AND3 (N1149, N1141, N439, N671);
xor XOR2 (N1150, N1146, N319);
buf BUF1 (N1151, N1148);
nand NAND3 (N1152, N1151, N673, N805);
nor NOR3 (N1153, N1142, N186, N782);
xor XOR2 (N1154, N1149, N245);
buf BUF1 (N1155, N1153);
xor XOR2 (N1156, N1154, N9);
not NOT1 (N1157, N1152);
nor NOR3 (N1158, N1157, N410, N271);
xor XOR2 (N1159, N1114, N52);
buf BUF1 (N1160, N1128);
xor XOR2 (N1161, N1156, N928);
not NOT1 (N1162, N1160);
buf BUF1 (N1163, N1162);
nor NOR4 (N1164, N1147, N76, N687, N498);
xor XOR2 (N1165, N1164, N2);
buf BUF1 (N1166, N1137);
not NOT1 (N1167, N1161);
xor XOR2 (N1168, N1140, N760);
not NOT1 (N1169, N1166);
xor XOR2 (N1170, N1138, N1080);
xor XOR2 (N1171, N1158, N512);
not NOT1 (N1172, N1163);
not NOT1 (N1173, N1172);
xor XOR2 (N1174, N1169, N197);
nor NOR2 (N1175, N1165, N564);
and AND3 (N1176, N1170, N449, N274);
buf BUF1 (N1177, N1155);
or OR4 (N1178, N1177, N1024, N966, N916);
buf BUF1 (N1179, N1176);
and AND3 (N1180, N1171, N120, N1155);
and AND3 (N1181, N1175, N559, N431);
buf BUF1 (N1182, N1181);
or OR2 (N1183, N1174, N434);
and AND3 (N1184, N1167, N823, N62);
nor NOR4 (N1185, N1179, N680, N341, N503);
or OR3 (N1186, N1182, N953, N28);
nand NAND2 (N1187, N1184, N57);
nor NOR2 (N1188, N1187, N687);
and AND3 (N1189, N1188, N889, N1056);
buf BUF1 (N1190, N1186);
xor XOR2 (N1191, N1178, N653);
xor XOR2 (N1192, N1191, N817);
or OR3 (N1193, N1180, N629, N1149);
and AND4 (N1194, N1185, N553, N1025, N613);
nor NOR4 (N1195, N1168, N756, N607, N260);
nand NAND3 (N1196, N1189, N157, N7);
xor XOR2 (N1197, N1159, N182);
buf BUF1 (N1198, N1193);
xor XOR2 (N1199, N1194, N900);
nor NOR2 (N1200, N1196, N121);
not NOT1 (N1201, N1190);
buf BUF1 (N1202, N1192);
buf BUF1 (N1203, N1198);
nand NAND4 (N1204, N1173, N558, N151, N655);
nor NOR3 (N1205, N1201, N638, N380);
and AND2 (N1206, N1202, N1074);
nor NOR3 (N1207, N1206, N441, N672);
not NOT1 (N1208, N1195);
xor XOR2 (N1209, N1203, N651);
buf BUF1 (N1210, N1208);
xor XOR2 (N1211, N1204, N337);
nand NAND3 (N1212, N1199, N895, N528);
buf BUF1 (N1213, N1211);
buf BUF1 (N1214, N1207);
nor NOR2 (N1215, N1214, N724);
and AND2 (N1216, N1200, N350);
nor NOR4 (N1217, N1216, N1054, N390, N370);
or OR4 (N1218, N1217, N205, N118, N482);
not NOT1 (N1219, N1215);
xor XOR2 (N1220, N1197, N777);
buf BUF1 (N1221, N1218);
not NOT1 (N1222, N1220);
nor NOR4 (N1223, N1222, N49, N825, N1067);
or OR2 (N1224, N1223, N69);
buf BUF1 (N1225, N1209);
buf BUF1 (N1226, N1224);
or OR3 (N1227, N1226, N572, N42);
nand NAND2 (N1228, N1227, N651);
or OR3 (N1229, N1225, N100, N1132);
xor XOR2 (N1230, N1212, N1103);
or OR2 (N1231, N1210, N995);
xor XOR2 (N1232, N1221, N345);
xor XOR2 (N1233, N1231, N707);
nand NAND4 (N1234, N1228, N1204, N268, N539);
nand NAND4 (N1235, N1183, N122, N314, N417);
nand NAND4 (N1236, N1233, N1091, N663, N121);
and AND3 (N1237, N1219, N1023, N1008);
and AND3 (N1238, N1232, N809, N148);
and AND3 (N1239, N1238, N814, N230);
or OR2 (N1240, N1234, N597);
not NOT1 (N1241, N1240);
nand NAND2 (N1242, N1205, N762);
and AND3 (N1243, N1241, N502, N1204);
buf BUF1 (N1244, N1235);
not NOT1 (N1245, N1242);
or OR4 (N1246, N1243, N1065, N328, N1063);
nor NOR3 (N1247, N1239, N730, N632);
buf BUF1 (N1248, N1150);
nand NAND2 (N1249, N1248, N1151);
xor XOR2 (N1250, N1236, N161);
and AND4 (N1251, N1237, N557, N423, N966);
buf BUF1 (N1252, N1245);
not NOT1 (N1253, N1230);
buf BUF1 (N1254, N1249);
or OR4 (N1255, N1252, N563, N583, N266);
buf BUF1 (N1256, N1246);
buf BUF1 (N1257, N1229);
not NOT1 (N1258, N1247);
and AND2 (N1259, N1253, N371);
buf BUF1 (N1260, N1256);
or OR2 (N1261, N1257, N104);
nor NOR4 (N1262, N1244, N1126, N431, N1076);
xor XOR2 (N1263, N1262, N247);
buf BUF1 (N1264, N1213);
and AND4 (N1265, N1259, N331, N1258, N729);
and AND2 (N1266, N262, N485);
not NOT1 (N1267, N1266);
or OR4 (N1268, N1254, N466, N859, N1143);
not NOT1 (N1269, N1268);
or OR4 (N1270, N1255, N909, N456, N260);
nor NOR2 (N1271, N1269, N1111);
or OR3 (N1272, N1271, N340, N193);
not NOT1 (N1273, N1263);
or OR4 (N1274, N1272, N1189, N1049, N1147);
nor NOR3 (N1275, N1267, N648, N356);
buf BUF1 (N1276, N1260);
not NOT1 (N1277, N1261);
xor XOR2 (N1278, N1251, N884);
not NOT1 (N1279, N1250);
xor XOR2 (N1280, N1265, N521);
and AND4 (N1281, N1273, N267, N466, N1189);
nand NAND4 (N1282, N1280, N1142, N298, N1088);
and AND2 (N1283, N1278, N244);
nand NAND2 (N1284, N1270, N131);
nand NAND2 (N1285, N1283, N807);
nor NOR2 (N1286, N1285, N1083);
nand NAND4 (N1287, N1274, N517, N1194, N1020);
buf BUF1 (N1288, N1281);
or OR4 (N1289, N1279, N34, N523, N928);
xor XOR2 (N1290, N1264, N919);
nand NAND3 (N1291, N1289, N468, N393);
buf BUF1 (N1292, N1290);
and AND4 (N1293, N1288, N52, N339, N827);
xor XOR2 (N1294, N1292, N1272);
not NOT1 (N1295, N1286);
and AND3 (N1296, N1294, N315, N697);
nor NOR3 (N1297, N1295, N960, N1046);
buf BUF1 (N1298, N1293);
xor XOR2 (N1299, N1284, N75);
buf BUF1 (N1300, N1277);
nor NOR3 (N1301, N1275, N812, N657);
buf BUF1 (N1302, N1296);
and AND4 (N1303, N1276, N1187, N967, N1064);
and AND4 (N1304, N1300, N1242, N1276, N302);
xor XOR2 (N1305, N1298, N524);
nand NAND2 (N1306, N1291, N1043);
or OR4 (N1307, N1303, N418, N874, N997);
not NOT1 (N1308, N1307);
buf BUF1 (N1309, N1301);
xor XOR2 (N1310, N1302, N404);
nor NOR3 (N1311, N1297, N463, N867);
or OR4 (N1312, N1309, N88, N510, N543);
and AND3 (N1313, N1310, N128, N666);
nand NAND4 (N1314, N1282, N1037, N68, N1013);
or OR4 (N1315, N1304, N368, N999, N486);
not NOT1 (N1316, N1299);
xor XOR2 (N1317, N1316, N644);
nand NAND3 (N1318, N1308, N243, N940);
or OR4 (N1319, N1313, N664, N1081, N373);
nand NAND2 (N1320, N1312, N1201);
not NOT1 (N1321, N1311);
and AND4 (N1322, N1305, N826, N1241, N586);
nor NOR2 (N1323, N1322, N234);
nor NOR3 (N1324, N1323, N230, N552);
xor XOR2 (N1325, N1306, N31);
nand NAND4 (N1326, N1315, N548, N166, N672);
buf BUF1 (N1327, N1321);
not NOT1 (N1328, N1318);
nor NOR3 (N1329, N1327, N558, N112);
and AND2 (N1330, N1329, N1155);
not NOT1 (N1331, N1330);
xor XOR2 (N1332, N1320, N724);
nor NOR3 (N1333, N1317, N77, N234);
nor NOR4 (N1334, N1319, N138, N869, N553);
not NOT1 (N1335, N1332);
not NOT1 (N1336, N1334);
not NOT1 (N1337, N1336);
not NOT1 (N1338, N1324);
xor XOR2 (N1339, N1338, N1117);
xor XOR2 (N1340, N1287, N1306);
or OR3 (N1341, N1325, N656, N318);
buf BUF1 (N1342, N1337);
not NOT1 (N1343, N1326);
buf BUF1 (N1344, N1340);
nor NOR2 (N1345, N1314, N1259);
and AND4 (N1346, N1343, N428, N468, N994);
or OR2 (N1347, N1341, N86);
xor XOR2 (N1348, N1328, N941);
xor XOR2 (N1349, N1339, N1287);
nand NAND3 (N1350, N1335, N997, N46);
xor XOR2 (N1351, N1347, N925);
buf BUF1 (N1352, N1345);
nor NOR2 (N1353, N1351, N839);
xor XOR2 (N1354, N1353, N1168);
nand NAND2 (N1355, N1350, N318);
buf BUF1 (N1356, N1333);
not NOT1 (N1357, N1331);
buf BUF1 (N1358, N1355);
xor XOR2 (N1359, N1349, N581);
buf BUF1 (N1360, N1359);
nand NAND2 (N1361, N1358, N1092);
and AND4 (N1362, N1354, N616, N156, N200);
nor NOR3 (N1363, N1346, N971, N635);
or OR2 (N1364, N1352, N932);
nor NOR3 (N1365, N1364, N350, N1183);
nand NAND3 (N1366, N1360, N819, N1341);
nand NAND2 (N1367, N1365, N569);
buf BUF1 (N1368, N1356);
nand NAND2 (N1369, N1348, N761);
nor NOR3 (N1370, N1369, N1336, N748);
or OR4 (N1371, N1363, N840, N708, N645);
not NOT1 (N1372, N1368);
nor NOR3 (N1373, N1366, N947, N1155);
and AND2 (N1374, N1362, N239);
nor NOR2 (N1375, N1370, N419);
xor XOR2 (N1376, N1344, N1250);
and AND4 (N1377, N1367, N1307, N442, N943);
xor XOR2 (N1378, N1371, N281);
not NOT1 (N1379, N1361);
or OR2 (N1380, N1377, N1356);
xor XOR2 (N1381, N1375, N1057);
and AND4 (N1382, N1373, N498, N1340, N1276);
nor NOR4 (N1383, N1376, N989, N930, N456);
nor NOR2 (N1384, N1380, N34);
not NOT1 (N1385, N1378);
or OR3 (N1386, N1379, N822, N472);
buf BUF1 (N1387, N1383);
buf BUF1 (N1388, N1357);
or OR4 (N1389, N1382, N4, N1131, N843);
nand NAND3 (N1390, N1342, N166, N332);
nor NOR2 (N1391, N1386, N876);
nand NAND2 (N1392, N1391, N1305);
and AND2 (N1393, N1372, N48);
and AND4 (N1394, N1388, N953, N38, N670);
nor NOR2 (N1395, N1392, N1264);
not NOT1 (N1396, N1394);
xor XOR2 (N1397, N1374, N963);
not NOT1 (N1398, N1384);
and AND3 (N1399, N1390, N551, N1013);
xor XOR2 (N1400, N1397, N20);
nand NAND2 (N1401, N1395, N1088);
and AND3 (N1402, N1381, N803, N671);
nor NOR4 (N1403, N1398, N582, N1309, N284);
or OR3 (N1404, N1385, N1179, N1378);
not NOT1 (N1405, N1402);
not NOT1 (N1406, N1403);
and AND2 (N1407, N1404, N147);
or OR4 (N1408, N1406, N1333, N1085, N379);
nand NAND4 (N1409, N1389, N912, N924, N1361);
not NOT1 (N1410, N1401);
and AND3 (N1411, N1407, N522, N383);
and AND3 (N1412, N1408, N88, N411);
or OR2 (N1413, N1410, N532);
buf BUF1 (N1414, N1399);
not NOT1 (N1415, N1393);
and AND2 (N1416, N1411, N309);
not NOT1 (N1417, N1413);
nand NAND3 (N1418, N1415, N372, N841);
or OR4 (N1419, N1412, N748, N656, N698);
buf BUF1 (N1420, N1414);
or OR4 (N1421, N1405, N551, N425, N414);
not NOT1 (N1422, N1421);
buf BUF1 (N1423, N1420);
not NOT1 (N1424, N1419);
nor NOR3 (N1425, N1409, N1408, N1371);
not NOT1 (N1426, N1416);
or OR3 (N1427, N1426, N1242, N874);
nand NAND2 (N1428, N1417, N350);
nor NOR3 (N1429, N1428, N809, N1380);
not NOT1 (N1430, N1422);
buf BUF1 (N1431, N1423);
buf BUF1 (N1432, N1396);
or OR4 (N1433, N1425, N1313, N735, N279);
xor XOR2 (N1434, N1418, N532);
nor NOR4 (N1435, N1427, N795, N799, N1291);
nor NOR2 (N1436, N1433, N836);
and AND3 (N1437, N1434, N1131, N988);
xor XOR2 (N1438, N1430, N21);
and AND4 (N1439, N1435, N938, N1178, N1153);
not NOT1 (N1440, N1436);
buf BUF1 (N1441, N1440);
nand NAND4 (N1442, N1441, N102, N519, N248);
buf BUF1 (N1443, N1442);
or OR3 (N1444, N1387, N1388, N1063);
xor XOR2 (N1445, N1444, N1393);
not NOT1 (N1446, N1438);
and AND2 (N1447, N1446, N782);
nor NOR4 (N1448, N1431, N32, N666, N1083);
buf BUF1 (N1449, N1400);
xor XOR2 (N1450, N1448, N501);
or OR2 (N1451, N1439, N425);
nor NOR4 (N1452, N1450, N788, N645, N81);
xor XOR2 (N1453, N1447, N555);
nor NOR4 (N1454, N1445, N203, N634, N778);
not NOT1 (N1455, N1432);
not NOT1 (N1456, N1454);
or OR4 (N1457, N1449, N382, N310, N496);
and AND3 (N1458, N1451, N1336, N808);
nor NOR4 (N1459, N1452, N409, N685, N574);
not NOT1 (N1460, N1458);
not NOT1 (N1461, N1429);
not NOT1 (N1462, N1457);
nor NOR4 (N1463, N1459, N1063, N1271, N1330);
nand NAND2 (N1464, N1463, N506);
xor XOR2 (N1465, N1461, N583);
nor NOR3 (N1466, N1456, N304, N1202);
nand NAND3 (N1467, N1455, N399, N1048);
nand NAND2 (N1468, N1424, N851);
nor NOR4 (N1469, N1443, N559, N382, N819);
and AND4 (N1470, N1453, N106, N94, N1426);
or OR2 (N1471, N1464, N517);
nor NOR2 (N1472, N1467, N541);
and AND3 (N1473, N1472, N961, N138);
nor NOR4 (N1474, N1437, N1044, N653, N1377);
or OR2 (N1475, N1465, N1356);
xor XOR2 (N1476, N1470, N578);
and AND2 (N1477, N1462, N417);
or OR3 (N1478, N1477, N320, N174);
or OR4 (N1479, N1478, N1261, N1256, N444);
not NOT1 (N1480, N1460);
nand NAND2 (N1481, N1480, N590);
and AND4 (N1482, N1475, N300, N1385, N1192);
and AND3 (N1483, N1466, N97, N867);
xor XOR2 (N1484, N1476, N1449);
or OR4 (N1485, N1482, N1200, N1024, N1433);
not NOT1 (N1486, N1485);
or OR2 (N1487, N1483, N745);
xor XOR2 (N1488, N1473, N288);
nor NOR2 (N1489, N1481, N1207);
or OR3 (N1490, N1474, N161, N878);
xor XOR2 (N1491, N1488, N862);
and AND4 (N1492, N1486, N1169, N517, N752);
or OR4 (N1493, N1471, N1162, N547, N14);
nand NAND4 (N1494, N1492, N1176, N710, N391);
buf BUF1 (N1495, N1468);
nand NAND4 (N1496, N1489, N87, N1250, N1463);
or OR2 (N1497, N1469, N103);
and AND3 (N1498, N1491, N1146, N479);
nor NOR2 (N1499, N1479, N728);
or OR4 (N1500, N1495, N920, N1421, N962);
nor NOR2 (N1501, N1499, N1256);
buf BUF1 (N1502, N1490);
and AND3 (N1503, N1500, N219, N1027);
and AND3 (N1504, N1493, N1473, N439);
buf BUF1 (N1505, N1484);
nor NOR3 (N1506, N1496, N308, N163);
buf BUF1 (N1507, N1487);
nor NOR3 (N1508, N1507, N495, N1413);
nand NAND2 (N1509, N1506, N1290);
buf BUF1 (N1510, N1501);
buf BUF1 (N1511, N1497);
or OR2 (N1512, N1508, N1463);
not NOT1 (N1513, N1504);
not NOT1 (N1514, N1494);
nor NOR2 (N1515, N1498, N746);
xor XOR2 (N1516, N1514, N429);
nand NAND4 (N1517, N1515, N338, N1025, N1414);
not NOT1 (N1518, N1509);
buf BUF1 (N1519, N1503);
xor XOR2 (N1520, N1516, N50);
nand NAND3 (N1521, N1517, N581, N1351);
nand NAND4 (N1522, N1518, N4, N374, N856);
buf BUF1 (N1523, N1502);
and AND2 (N1524, N1505, N1395);
xor XOR2 (N1525, N1524, N88);
xor XOR2 (N1526, N1522, N1397);
and AND3 (N1527, N1525, N263, N1379);
and AND2 (N1528, N1520, N1106);
not NOT1 (N1529, N1528);
not NOT1 (N1530, N1510);
nor NOR3 (N1531, N1527, N440, N524);
xor XOR2 (N1532, N1529, N518);
buf BUF1 (N1533, N1523);
not NOT1 (N1534, N1519);
nor NOR3 (N1535, N1511, N284, N1180);
buf BUF1 (N1536, N1526);
xor XOR2 (N1537, N1530, N1269);
nor NOR3 (N1538, N1535, N1235, N268);
buf BUF1 (N1539, N1532);
or OR3 (N1540, N1537, N1532, N594);
nor NOR3 (N1541, N1540, N625, N996);
and AND4 (N1542, N1512, N800, N331, N1181);
or OR3 (N1543, N1536, N80, N404);
not NOT1 (N1544, N1541);
and AND4 (N1545, N1531, N145, N1520, N281);
nand NAND2 (N1546, N1521, N834);
nand NAND2 (N1547, N1544, N1104);
and AND2 (N1548, N1538, N1327);
nor NOR3 (N1549, N1546, N1308, N249);
and AND2 (N1550, N1549, N858);
and AND2 (N1551, N1542, N602);
nor NOR2 (N1552, N1513, N452);
not NOT1 (N1553, N1552);
buf BUF1 (N1554, N1551);
not NOT1 (N1555, N1534);
xor XOR2 (N1556, N1553, N1479);
xor XOR2 (N1557, N1548, N592);
xor XOR2 (N1558, N1539, N1465);
xor XOR2 (N1559, N1550, N352);
or OR4 (N1560, N1556, N1554, N424, N487);
buf BUF1 (N1561, N991);
buf BUF1 (N1562, N1558);
xor XOR2 (N1563, N1533, N1216);
xor XOR2 (N1564, N1563, N631);
xor XOR2 (N1565, N1547, N679);
nor NOR3 (N1566, N1545, N1456, N795);
buf BUF1 (N1567, N1562);
nand NAND2 (N1568, N1561, N1050);
not NOT1 (N1569, N1568);
buf BUF1 (N1570, N1567);
not NOT1 (N1571, N1555);
nor NOR4 (N1572, N1543, N1224, N1387, N1065);
and AND3 (N1573, N1569, N168, N1297);
buf BUF1 (N1574, N1566);
and AND2 (N1575, N1565, N1535);
xor XOR2 (N1576, N1575, N368);
nor NOR3 (N1577, N1564, N988, N924);
or OR2 (N1578, N1557, N81);
nor NOR3 (N1579, N1577, N1155, N857);
nor NOR4 (N1580, N1573, N577, N1294, N1041);
nor NOR2 (N1581, N1576, N596);
or OR3 (N1582, N1560, N103, N272);
or OR2 (N1583, N1582, N364);
nand NAND4 (N1584, N1574, N947, N1424, N500);
nand NAND4 (N1585, N1570, N625, N484, N1026);
not NOT1 (N1586, N1559);
buf BUF1 (N1587, N1581);
not NOT1 (N1588, N1585);
or OR2 (N1589, N1586, N1544);
not NOT1 (N1590, N1571);
or OR2 (N1591, N1590, N1056);
or OR2 (N1592, N1579, N499);
xor XOR2 (N1593, N1589, N1382);
nor NOR4 (N1594, N1583, N1448, N195, N1342);
and AND3 (N1595, N1588, N60, N1483);
buf BUF1 (N1596, N1594);
and AND2 (N1597, N1578, N625);
nand NAND2 (N1598, N1597, N846);
buf BUF1 (N1599, N1598);
buf BUF1 (N1600, N1584);
or OR4 (N1601, N1580, N804, N1417, N1223);
not NOT1 (N1602, N1595);
and AND2 (N1603, N1591, N603);
buf BUF1 (N1604, N1572);
nand NAND4 (N1605, N1592, N565, N126, N349);
xor XOR2 (N1606, N1593, N656);
xor XOR2 (N1607, N1606, N1014);
nor NOR3 (N1608, N1602, N408, N511);
xor XOR2 (N1609, N1599, N247);
nor NOR3 (N1610, N1596, N803, N1195);
buf BUF1 (N1611, N1601);
nand NAND2 (N1612, N1603, N443);
nor NOR3 (N1613, N1600, N459, N899);
nor NOR3 (N1614, N1608, N1129, N6);
nor NOR3 (N1615, N1610, N1568, N1593);
buf BUF1 (N1616, N1614);
xor XOR2 (N1617, N1612, N1453);
nor NOR4 (N1618, N1613, N14, N3, N235);
and AND4 (N1619, N1607, N394, N644, N257);
not NOT1 (N1620, N1618);
nor NOR4 (N1621, N1605, N438, N801, N539);
or OR3 (N1622, N1604, N284, N357);
xor XOR2 (N1623, N1621, N1550);
xor XOR2 (N1624, N1616, N919);
not NOT1 (N1625, N1587);
not NOT1 (N1626, N1622);
not NOT1 (N1627, N1625);
nand NAND4 (N1628, N1617, N1179, N924, N859);
nor NOR3 (N1629, N1615, N958, N961);
not NOT1 (N1630, N1629);
and AND2 (N1631, N1620, N834);
or OR3 (N1632, N1609, N944, N1225);
and AND2 (N1633, N1619, N1575);
nor NOR3 (N1634, N1626, N609, N693);
nor NOR2 (N1635, N1633, N494);
nor NOR4 (N1636, N1628, N941, N349, N363);
nand NAND3 (N1637, N1627, N1402, N932);
nand NAND4 (N1638, N1635, N586, N1212, N1618);
nand NAND4 (N1639, N1638, N1042, N1541, N672);
buf BUF1 (N1640, N1636);
and AND3 (N1641, N1631, N412, N167);
nand NAND2 (N1642, N1641, N988);
xor XOR2 (N1643, N1634, N435);
nor NOR4 (N1644, N1630, N838, N487, N1290);
xor XOR2 (N1645, N1644, N50);
not NOT1 (N1646, N1643);
and AND4 (N1647, N1632, N456, N257, N1189);
and AND2 (N1648, N1611, N1522);
not NOT1 (N1649, N1646);
and AND4 (N1650, N1649, N1504, N229, N1565);
nand NAND4 (N1651, N1648, N760, N1596, N494);
buf BUF1 (N1652, N1650);
not NOT1 (N1653, N1652);
not NOT1 (N1654, N1651);
buf BUF1 (N1655, N1642);
or OR3 (N1656, N1623, N149, N302);
nand NAND3 (N1657, N1654, N733, N1344);
and AND2 (N1658, N1640, N165);
and AND3 (N1659, N1657, N1376, N967);
xor XOR2 (N1660, N1656, N592);
buf BUF1 (N1661, N1659);
nand NAND4 (N1662, N1661, N1210, N1274, N1508);
or OR4 (N1663, N1647, N1388, N28, N1621);
and AND3 (N1664, N1663, N1200, N912);
xor XOR2 (N1665, N1645, N450);
buf BUF1 (N1666, N1658);
buf BUF1 (N1667, N1655);
xor XOR2 (N1668, N1660, N1431);
xor XOR2 (N1669, N1664, N40);
nor NOR3 (N1670, N1665, N748, N779);
nand NAND2 (N1671, N1668, N927);
nand NAND4 (N1672, N1653, N7, N171, N1146);
not NOT1 (N1673, N1671);
buf BUF1 (N1674, N1666);
buf BUF1 (N1675, N1670);
not NOT1 (N1676, N1662);
xor XOR2 (N1677, N1674, N1092);
buf BUF1 (N1678, N1677);
buf BUF1 (N1679, N1639);
xor XOR2 (N1680, N1676, N562);
xor XOR2 (N1681, N1624, N509);
not NOT1 (N1682, N1681);
nand NAND4 (N1683, N1673, N55, N1665, N299);
xor XOR2 (N1684, N1637, N960);
and AND4 (N1685, N1680, N1515, N1567, N954);
nor NOR4 (N1686, N1682, N1581, N907, N1427);
and AND4 (N1687, N1679, N1212, N1000, N1180);
nand NAND2 (N1688, N1686, N1496);
xor XOR2 (N1689, N1672, N1681);
or OR4 (N1690, N1687, N285, N280, N113);
or OR4 (N1691, N1684, N140, N1651, N964);
buf BUF1 (N1692, N1689);
xor XOR2 (N1693, N1683, N1229);
and AND2 (N1694, N1669, N668);
buf BUF1 (N1695, N1688);
xor XOR2 (N1696, N1692, N824);
or OR3 (N1697, N1693, N1496, N377);
not NOT1 (N1698, N1678);
buf BUF1 (N1699, N1698);
buf BUF1 (N1700, N1691);
and AND3 (N1701, N1696, N1022, N272);
nor NOR2 (N1702, N1675, N803);
or OR4 (N1703, N1695, N646, N1428, N479);
nand NAND3 (N1704, N1697, N700, N137);
nor NOR4 (N1705, N1701, N1144, N1349, N1132);
and AND4 (N1706, N1699, N185, N863, N816);
and AND4 (N1707, N1704, N1270, N846, N394);
buf BUF1 (N1708, N1690);
nand NAND2 (N1709, N1705, N224);
and AND2 (N1710, N1694, N1022);
not NOT1 (N1711, N1710);
or OR4 (N1712, N1711, N62, N941, N1623);
nor NOR2 (N1713, N1700, N657);
nand NAND3 (N1714, N1706, N1527, N1387);
not NOT1 (N1715, N1685);
not NOT1 (N1716, N1713);
nor NOR2 (N1717, N1709, N1417);
buf BUF1 (N1718, N1702);
buf BUF1 (N1719, N1708);
xor XOR2 (N1720, N1715, N162);
nor NOR3 (N1721, N1719, N77, N1193);
xor XOR2 (N1722, N1712, N1221);
or OR2 (N1723, N1714, N1139);
and AND2 (N1724, N1667, N1109);
and AND3 (N1725, N1703, N555, N414);
and AND3 (N1726, N1725, N1488, N100);
nand NAND3 (N1727, N1707, N1042, N482);
nand NAND3 (N1728, N1726, N894, N1162);
and AND4 (N1729, N1720, N1647, N684, N829);
nor NOR3 (N1730, N1716, N907, N753);
buf BUF1 (N1731, N1724);
not NOT1 (N1732, N1729);
buf BUF1 (N1733, N1721);
and AND4 (N1734, N1722, N1449, N1017, N1619);
nor NOR2 (N1735, N1728, N59);
not NOT1 (N1736, N1723);
or OR2 (N1737, N1736, N859);
nand NAND2 (N1738, N1730, N1219);
xor XOR2 (N1739, N1733, N856);
not NOT1 (N1740, N1739);
xor XOR2 (N1741, N1718, N47);
and AND4 (N1742, N1727, N1113, N580, N311);
xor XOR2 (N1743, N1731, N810);
not NOT1 (N1744, N1738);
buf BUF1 (N1745, N1741);
nand NAND2 (N1746, N1732, N1065);
not NOT1 (N1747, N1742);
or OR2 (N1748, N1745, N451);
buf BUF1 (N1749, N1748);
nand NAND4 (N1750, N1749, N675, N777, N512);
buf BUF1 (N1751, N1747);
buf BUF1 (N1752, N1737);
or OR4 (N1753, N1735, N1659, N655, N91);
buf BUF1 (N1754, N1750);
and AND2 (N1755, N1746, N529);
not NOT1 (N1756, N1754);
or OR3 (N1757, N1755, N1383, N1069);
xor XOR2 (N1758, N1756, N1351);
and AND4 (N1759, N1744, N655, N1164, N609);
nand NAND2 (N1760, N1751, N636);
and AND3 (N1761, N1740, N80, N777);
not NOT1 (N1762, N1717);
nor NOR3 (N1763, N1743, N1685, N1146);
nor NOR2 (N1764, N1753, N383);
not NOT1 (N1765, N1762);
not NOT1 (N1766, N1760);
xor XOR2 (N1767, N1758, N1724);
and AND2 (N1768, N1766, N1737);
nand NAND4 (N1769, N1761, N459, N842, N1323);
buf BUF1 (N1770, N1763);
not NOT1 (N1771, N1770);
nor NOR3 (N1772, N1764, N727, N460);
nor NOR4 (N1773, N1765, N1182, N1034, N1008);
or OR3 (N1774, N1772, N963, N1538);
and AND4 (N1775, N1774, N581, N626, N595);
nor NOR3 (N1776, N1771, N1523, N78);
xor XOR2 (N1777, N1775, N792);
and AND3 (N1778, N1776, N142, N498);
nand NAND2 (N1779, N1767, N1513);
or OR4 (N1780, N1777, N1242, N620, N87);
not NOT1 (N1781, N1757);
or OR3 (N1782, N1759, N1730, N1561);
or OR3 (N1783, N1752, N1027, N1663);
and AND2 (N1784, N1779, N552);
or OR4 (N1785, N1769, N1719, N1062, N1441);
xor XOR2 (N1786, N1768, N626);
and AND2 (N1787, N1780, N761);
nand NAND3 (N1788, N1781, N1590, N335);
nor NOR2 (N1789, N1782, N1650);
nor NOR4 (N1790, N1789, N640, N1473, N1736);
not NOT1 (N1791, N1790);
or OR4 (N1792, N1773, N314, N1085, N1725);
not NOT1 (N1793, N1792);
and AND2 (N1794, N1778, N1491);
or OR2 (N1795, N1786, N1334);
and AND3 (N1796, N1787, N1733, N623);
nor NOR4 (N1797, N1783, N894, N194, N1539);
not NOT1 (N1798, N1793);
buf BUF1 (N1799, N1734);
or OR3 (N1800, N1798, N618, N850);
buf BUF1 (N1801, N1797);
nor NOR3 (N1802, N1796, N1713, N12);
not NOT1 (N1803, N1799);
buf BUF1 (N1804, N1794);
buf BUF1 (N1805, N1784);
not NOT1 (N1806, N1804);
or OR4 (N1807, N1800, N492, N1663, N1266);
xor XOR2 (N1808, N1806, N1617);
or OR4 (N1809, N1788, N1697, N17, N1373);
xor XOR2 (N1810, N1791, N1656);
buf BUF1 (N1811, N1785);
buf BUF1 (N1812, N1807);
nand NAND2 (N1813, N1812, N1803);
buf BUF1 (N1814, N407);
or OR4 (N1815, N1805, N77, N1399, N893);
nand NAND4 (N1816, N1795, N734, N1434, N880);
or OR3 (N1817, N1815, N1530, N557);
not NOT1 (N1818, N1811);
nand NAND4 (N1819, N1810, N466, N852, N313);
and AND2 (N1820, N1808, N856);
or OR3 (N1821, N1809, N505, N678);
or OR2 (N1822, N1818, N580);
buf BUF1 (N1823, N1820);
buf BUF1 (N1824, N1814);
nor NOR2 (N1825, N1817, N130);
nor NOR2 (N1826, N1823, N1740);
nand NAND3 (N1827, N1822, N1600, N1170);
or OR4 (N1828, N1824, N1649, N90, N419);
nor NOR3 (N1829, N1828, N205, N593);
nor NOR4 (N1830, N1816, N1666, N1489, N604);
or OR4 (N1831, N1829, N1428, N1070, N1564);
buf BUF1 (N1832, N1831);
and AND2 (N1833, N1830, N1627);
not NOT1 (N1834, N1819);
or OR2 (N1835, N1801, N1205);
nand NAND3 (N1836, N1832, N643, N1601);
not NOT1 (N1837, N1836);
not NOT1 (N1838, N1813);
nor NOR2 (N1839, N1826, N1183);
xor XOR2 (N1840, N1839, N1201);
xor XOR2 (N1841, N1825, N1280);
xor XOR2 (N1842, N1835, N1402);
buf BUF1 (N1843, N1840);
buf BUF1 (N1844, N1842);
nor NOR4 (N1845, N1827, N238, N1221, N1449);
nor NOR4 (N1846, N1802, N414, N547, N1485);
or OR4 (N1847, N1843, N1084, N201, N209);
or OR3 (N1848, N1834, N1127, N45);
or OR4 (N1849, N1833, N1633, N422, N1083);
not NOT1 (N1850, N1845);
xor XOR2 (N1851, N1849, N611);
nor NOR4 (N1852, N1837, N1003, N1846, N1166);
and AND2 (N1853, N1698, N247);
and AND3 (N1854, N1850, N969, N1373);
nor NOR2 (N1855, N1847, N62);
nand NAND4 (N1856, N1838, N1562, N1749, N835);
xor XOR2 (N1857, N1851, N836);
buf BUF1 (N1858, N1857);
xor XOR2 (N1859, N1821, N1781);
and AND4 (N1860, N1859, N813, N1341, N1384);
or OR3 (N1861, N1844, N1260, N1664);
or OR2 (N1862, N1841, N120);
xor XOR2 (N1863, N1853, N262);
or OR3 (N1864, N1862, N1216, N543);
nor NOR3 (N1865, N1860, N453, N1682);
not NOT1 (N1866, N1861);
xor XOR2 (N1867, N1866, N1418);
or OR4 (N1868, N1854, N684, N711, N890);
and AND2 (N1869, N1858, N1322);
nand NAND4 (N1870, N1856, N1743, N566, N1605);
nor NOR4 (N1871, N1869, N1458, N1765, N95);
not NOT1 (N1872, N1865);
nand NAND3 (N1873, N1848, N1808, N1045);
and AND2 (N1874, N1867, N483);
or OR3 (N1875, N1872, N768, N934);
nor NOR3 (N1876, N1874, N1434, N30);
or OR2 (N1877, N1863, N211);
not NOT1 (N1878, N1870);
not NOT1 (N1879, N1868);
nor NOR4 (N1880, N1875, N1069, N946, N1315);
and AND2 (N1881, N1873, N1076);
buf BUF1 (N1882, N1864);
buf BUF1 (N1883, N1880);
and AND2 (N1884, N1883, N1719);
xor XOR2 (N1885, N1855, N777);
nand NAND4 (N1886, N1871, N1381, N1620, N248);
not NOT1 (N1887, N1877);
nor NOR4 (N1888, N1884, N93, N341, N125);
xor XOR2 (N1889, N1852, N133);
not NOT1 (N1890, N1887);
and AND2 (N1891, N1885, N1429);
buf BUF1 (N1892, N1879);
nand NAND4 (N1893, N1891, N1821, N1202, N909);
buf BUF1 (N1894, N1890);
nand NAND3 (N1895, N1881, N578, N276);
not NOT1 (N1896, N1895);
xor XOR2 (N1897, N1893, N515);
xor XOR2 (N1898, N1896, N1687);
not NOT1 (N1899, N1892);
nand NAND3 (N1900, N1878, N913, N1893);
not NOT1 (N1901, N1888);
buf BUF1 (N1902, N1882);
or OR4 (N1903, N1897, N276, N1812, N1084);
and AND4 (N1904, N1894, N1034, N759, N180);
and AND3 (N1905, N1898, N447, N950);
xor XOR2 (N1906, N1899, N1356);
not NOT1 (N1907, N1904);
buf BUF1 (N1908, N1886);
not NOT1 (N1909, N1903);
or OR2 (N1910, N1905, N1156);
nor NOR4 (N1911, N1900, N735, N977, N763);
and AND3 (N1912, N1911, N1442, N1042);
buf BUF1 (N1913, N1912);
or OR3 (N1914, N1901, N1152, N684);
nand NAND3 (N1915, N1906, N574, N1609);
nor NOR3 (N1916, N1889, N779, N1215);
not NOT1 (N1917, N1908);
not NOT1 (N1918, N1916);
and AND4 (N1919, N1914, N1354, N1884, N1899);
or OR2 (N1920, N1909, N1550);
buf BUF1 (N1921, N1918);
nor NOR4 (N1922, N1902, N1879, N1552, N1353);
nor NOR2 (N1923, N1915, N40);
nor NOR3 (N1924, N1910, N1110, N1587);
nand NAND3 (N1925, N1923, N546, N121);
or OR3 (N1926, N1913, N359, N1672);
xor XOR2 (N1927, N1907, N731);
not NOT1 (N1928, N1924);
xor XOR2 (N1929, N1927, N1497);
nor NOR2 (N1930, N1928, N344);
nor NOR4 (N1931, N1926, N311, N1286, N213);
not NOT1 (N1932, N1930);
xor XOR2 (N1933, N1919, N1499);
nor NOR2 (N1934, N1929, N1528);
or OR3 (N1935, N1931, N1480, N1871);
not NOT1 (N1936, N1876);
or OR3 (N1937, N1935, N1381, N633);
not NOT1 (N1938, N1921);
not NOT1 (N1939, N1934);
nor NOR3 (N1940, N1920, N1455, N1637);
buf BUF1 (N1941, N1939);
or OR3 (N1942, N1922, N390, N1068);
nand NAND2 (N1943, N1932, N185);
or OR2 (N1944, N1933, N506);
xor XOR2 (N1945, N1936, N1799);
not NOT1 (N1946, N1937);
xor XOR2 (N1947, N1938, N208);
not NOT1 (N1948, N1947);
xor XOR2 (N1949, N1943, N809);
buf BUF1 (N1950, N1942);
nand NAND4 (N1951, N1940, N1944, N100, N1160);
and AND3 (N1952, N913, N1404, N1420);
buf BUF1 (N1953, N1941);
nand NAND3 (N1954, N1949, N1459, N1823);
buf BUF1 (N1955, N1952);
xor XOR2 (N1956, N1946, N1895);
not NOT1 (N1957, N1951);
or OR4 (N1958, N1925, N1799, N969, N634);
buf BUF1 (N1959, N1955);
nand NAND3 (N1960, N1953, N452, N58);
nor NOR2 (N1961, N1954, N1567);
not NOT1 (N1962, N1945);
or OR3 (N1963, N1948, N891, N1959);
and AND4 (N1964, N902, N1331, N1504, N1653);
nor NOR2 (N1965, N1917, N187);
not NOT1 (N1966, N1958);
xor XOR2 (N1967, N1957, N267);
nor NOR3 (N1968, N1961, N585, N133);
nor NOR2 (N1969, N1962, N1402);
nor NOR4 (N1970, N1968, N972, N1146, N1529);
xor XOR2 (N1971, N1967, N77);
or OR2 (N1972, N1970, N734);
or OR4 (N1973, N1960, N181, N1078, N69);
xor XOR2 (N1974, N1963, N1500);
and AND4 (N1975, N1965, N1078, N619, N1637);
and AND3 (N1976, N1964, N396, N1961);
buf BUF1 (N1977, N1974);
nand NAND3 (N1978, N1976, N1465, N1867);
nand NAND2 (N1979, N1972, N1978);
or OR2 (N1980, N587, N888);
and AND2 (N1981, N1966, N154);
nand NAND4 (N1982, N1950, N810, N1181, N832);
not NOT1 (N1983, N1977);
not NOT1 (N1984, N1979);
or OR3 (N1985, N1956, N1069, N473);
or OR2 (N1986, N1975, N89);
and AND2 (N1987, N1969, N433);
not NOT1 (N1988, N1984);
nor NOR2 (N1989, N1985, N1095);
nor NOR4 (N1990, N1981, N1760, N1103, N909);
and AND3 (N1991, N1989, N1663, N1416);
and AND2 (N1992, N1987, N1725);
nor NOR2 (N1993, N1973, N1180);
nand NAND2 (N1994, N1990, N41);
nor NOR4 (N1995, N1988, N1703, N454, N6);
nor NOR2 (N1996, N1982, N1645);
not NOT1 (N1997, N1983);
nand NAND3 (N1998, N1991, N396, N1540);
nand NAND4 (N1999, N1998, N705, N85, N811);
nand NAND4 (N2000, N1997, N549, N1330, N477);
nor NOR2 (N2001, N1999, N416);
nand NAND2 (N2002, N1996, N1747);
xor XOR2 (N2003, N1992, N1349);
nor NOR2 (N2004, N1993, N1852);
xor XOR2 (N2005, N2001, N427);
not NOT1 (N2006, N2004);
and AND4 (N2007, N2002, N214, N1578, N704);
buf BUF1 (N2008, N2000);
or OR2 (N2009, N1986, N942);
or OR3 (N2010, N2008, N26, N338);
xor XOR2 (N2011, N2009, N1164);
not NOT1 (N2012, N2006);
nand NAND4 (N2013, N2005, N52, N1820, N317);
buf BUF1 (N2014, N2012);
xor XOR2 (N2015, N2013, N759);
nand NAND4 (N2016, N2010, N306, N773, N1464);
and AND3 (N2017, N2015, N1265, N112);
buf BUF1 (N2018, N2007);
buf BUF1 (N2019, N1971);
buf BUF1 (N2020, N1980);
not NOT1 (N2021, N2011);
xor XOR2 (N2022, N2018, N609);
not NOT1 (N2023, N2003);
or OR3 (N2024, N2020, N1717, N1579);
not NOT1 (N2025, N2022);
not NOT1 (N2026, N2021);
not NOT1 (N2027, N2017);
or OR3 (N2028, N2014, N359, N1888);
xor XOR2 (N2029, N1994, N291);
xor XOR2 (N2030, N2026, N642);
buf BUF1 (N2031, N2030);
not NOT1 (N2032, N2028);
or OR4 (N2033, N2031, N978, N394, N1970);
nand NAND2 (N2034, N1995, N248);
or OR4 (N2035, N2034, N622, N1744, N1646);
nor NOR4 (N2036, N2027, N149, N1795, N364);
and AND3 (N2037, N2033, N1734, N295);
and AND3 (N2038, N2016, N425, N1030);
nor NOR2 (N2039, N2019, N1634);
nand NAND3 (N2040, N2032, N50, N897);
and AND3 (N2041, N2024, N1005, N1830);
not NOT1 (N2042, N2035);
xor XOR2 (N2043, N2038, N283);
not NOT1 (N2044, N2039);
xor XOR2 (N2045, N2023, N109);
and AND3 (N2046, N2040, N1214, N81);
xor XOR2 (N2047, N2044, N511);
buf BUF1 (N2048, N2036);
buf BUF1 (N2049, N2041);
buf BUF1 (N2050, N2037);
or OR2 (N2051, N2045, N1597);
nand NAND4 (N2052, N2046, N1719, N971, N1331);
or OR3 (N2053, N2042, N1048, N1659);
not NOT1 (N2054, N2050);
and AND2 (N2055, N2053, N940);
and AND4 (N2056, N2047, N296, N722, N1122);
nor NOR2 (N2057, N2048, N921);
nor NOR4 (N2058, N2055, N1248, N1380, N737);
not NOT1 (N2059, N2058);
or OR2 (N2060, N2051, N2020);
buf BUF1 (N2061, N2056);
nor NOR4 (N2062, N2059, N1543, N1296, N1057);
nand NAND4 (N2063, N2054, N1890, N975, N1787);
not NOT1 (N2064, N2049);
nand NAND3 (N2065, N2062, N1075, N1852);
and AND3 (N2066, N2043, N1344, N186);
and AND3 (N2067, N2066, N1690, N1327);
nor NOR4 (N2068, N2029, N936, N139, N1548);
nand NAND3 (N2069, N2052, N796, N1755);
xor XOR2 (N2070, N2068, N2018);
buf BUF1 (N2071, N2065);
xor XOR2 (N2072, N2063, N1065);
and AND4 (N2073, N2071, N367, N1191, N1696);
and AND3 (N2074, N2060, N775, N1110);
buf BUF1 (N2075, N2025);
not NOT1 (N2076, N2069);
nand NAND3 (N2077, N2074, N1845, N698);
xor XOR2 (N2078, N2067, N533);
nand NAND3 (N2079, N2070, N764, N1027);
nor NOR3 (N2080, N2057, N1621, N1672);
and AND2 (N2081, N2072, N139);
nand NAND4 (N2082, N2080, N1253, N853, N597);
and AND4 (N2083, N2076, N1318, N1363, N209);
and AND2 (N2084, N2083, N534);
buf BUF1 (N2085, N2084);
nand NAND3 (N2086, N2078, N2052, N919);
xor XOR2 (N2087, N2077, N445);
nand NAND3 (N2088, N2082, N1932, N1876);
and AND3 (N2089, N2079, N1457, N1759);
and AND2 (N2090, N2086, N1498);
xor XOR2 (N2091, N2089, N693);
xor XOR2 (N2092, N2087, N1633);
not NOT1 (N2093, N2064);
nand NAND4 (N2094, N2091, N298, N1253, N278);
and AND3 (N2095, N2075, N241, N1723);
nand NAND4 (N2096, N2090, N1033, N616, N235);
or OR2 (N2097, N2081, N1951);
buf BUF1 (N2098, N2085);
nand NAND3 (N2099, N2098, N1339, N904);
or OR4 (N2100, N2097, N578, N2023, N1299);
nand NAND4 (N2101, N2099, N1646, N1169, N829);
not NOT1 (N2102, N2093);
and AND2 (N2103, N2101, N667);
nand NAND2 (N2104, N2095, N553);
not NOT1 (N2105, N2096);
or OR2 (N2106, N2105, N1293);
or OR2 (N2107, N2100, N2010);
and AND4 (N2108, N2103, N1299, N1115, N1563);
nand NAND3 (N2109, N2108, N182, N1994);
buf BUF1 (N2110, N2106);
nand NAND3 (N2111, N2073, N63, N311);
or OR4 (N2112, N2102, N1258, N1888, N952);
nand NAND4 (N2113, N2094, N1356, N1854, N727);
nand NAND4 (N2114, N2110, N2103, N774, N680);
or OR4 (N2115, N2061, N1225, N1543, N1729);
xor XOR2 (N2116, N2088, N1304);
xor XOR2 (N2117, N2111, N1267);
buf BUF1 (N2118, N2107);
buf BUF1 (N2119, N2104);
or OR2 (N2120, N2113, N422);
nand NAND3 (N2121, N2109, N916, N826);
or OR2 (N2122, N2112, N1693);
not NOT1 (N2123, N2122);
not NOT1 (N2124, N2120);
not NOT1 (N2125, N2115);
buf BUF1 (N2126, N2118);
and AND3 (N2127, N2123, N1409, N1012);
not NOT1 (N2128, N2121);
and AND3 (N2129, N2126, N1668, N1842);
not NOT1 (N2130, N2092);
not NOT1 (N2131, N2119);
nor NOR4 (N2132, N2124, N952, N1822, N752);
nor NOR3 (N2133, N2131, N934, N1989);
not NOT1 (N2134, N2114);
or OR4 (N2135, N2129, N627, N552, N334);
or OR4 (N2136, N2135, N775, N48, N383);
or OR4 (N2137, N2116, N249, N640, N1114);
xor XOR2 (N2138, N2128, N1973);
nor NOR4 (N2139, N2134, N1690, N143, N960);
buf BUF1 (N2140, N2130);
nand NAND2 (N2141, N2139, N2091);
buf BUF1 (N2142, N2127);
and AND3 (N2143, N2132, N1933, N1538);
buf BUF1 (N2144, N2141);
and AND3 (N2145, N2138, N1306, N250);
xor XOR2 (N2146, N2140, N1259);
xor XOR2 (N2147, N2137, N1745);
xor XOR2 (N2148, N2125, N173);
or OR3 (N2149, N2144, N1948, N1349);
buf BUF1 (N2150, N2142);
nand NAND3 (N2151, N2117, N1364, N2150);
xor XOR2 (N2152, N2013, N645);
xor XOR2 (N2153, N2146, N1067);
not NOT1 (N2154, N2152);
and AND2 (N2155, N2147, N266);
and AND4 (N2156, N2153, N595, N1669, N672);
nor NOR3 (N2157, N2145, N425, N1467);
xor XOR2 (N2158, N2143, N1416);
and AND2 (N2159, N2149, N198);
xor XOR2 (N2160, N2151, N608);
nor NOR4 (N2161, N2148, N42, N715, N1672);
nor NOR2 (N2162, N2136, N1483);
nand NAND3 (N2163, N2159, N1873, N439);
not NOT1 (N2164, N2162);
xor XOR2 (N2165, N2133, N1833);
nor NOR2 (N2166, N2160, N1419);
nor NOR3 (N2167, N2154, N882, N1170);
and AND4 (N2168, N2155, N1747, N2046, N118);
xor XOR2 (N2169, N2158, N1672);
nor NOR4 (N2170, N2165, N438, N108, N899);
and AND2 (N2171, N2156, N16);
not NOT1 (N2172, N2166);
or OR2 (N2173, N2167, N385);
and AND3 (N2174, N2168, N1372, N1913);
not NOT1 (N2175, N2161);
nor NOR4 (N2176, N2171, N1648, N221, N1392);
nand NAND4 (N2177, N2163, N44, N1093, N2027);
nand NAND4 (N2178, N2174, N264, N1824, N225);
xor XOR2 (N2179, N2170, N1236);
and AND2 (N2180, N2157, N1963);
not NOT1 (N2181, N2172);
not NOT1 (N2182, N2169);
nor NOR2 (N2183, N2180, N507);
and AND3 (N2184, N2179, N918, N1741);
and AND2 (N2185, N2164, N1643);
xor XOR2 (N2186, N2185, N526);
not NOT1 (N2187, N2178);
nand NAND3 (N2188, N2181, N2096, N438);
not NOT1 (N2189, N2186);
and AND4 (N2190, N2177, N1294, N1576, N1286);
nor NOR2 (N2191, N2190, N1126);
nand NAND2 (N2192, N2184, N1323);
or OR3 (N2193, N2192, N977, N1509);
nand NAND2 (N2194, N2182, N227);
and AND3 (N2195, N2187, N918, N102);
nand NAND4 (N2196, N2191, N1605, N1662, N238);
not NOT1 (N2197, N2188);
nor NOR3 (N2198, N2195, N1376, N306);
nor NOR3 (N2199, N2183, N1080, N1237);
nand NAND4 (N2200, N2198, N634, N763, N1311);
buf BUF1 (N2201, N2194);
or OR2 (N2202, N2199, N1274);
and AND2 (N2203, N2176, N1840);
nand NAND2 (N2204, N2189, N2027);
buf BUF1 (N2205, N2202);
not NOT1 (N2206, N2175);
not NOT1 (N2207, N2197);
and AND4 (N2208, N2207, N2056, N407, N2207);
nand NAND3 (N2209, N2206, N665, N2015);
and AND4 (N2210, N2205, N543, N154, N1841);
not NOT1 (N2211, N2196);
nand NAND3 (N2212, N2193, N1496, N1572);
and AND3 (N2213, N2203, N93, N532);
nor NOR4 (N2214, N2210, N1325, N219, N555);
not NOT1 (N2215, N2213);
buf BUF1 (N2216, N2214);
and AND3 (N2217, N2215, N1257, N168);
nand NAND3 (N2218, N2216, N2190, N103);
buf BUF1 (N2219, N2200);
or OR2 (N2220, N2217, N186);
or OR4 (N2221, N2209, N491, N1276, N2198);
or OR4 (N2222, N2212, N236, N1552, N1676);
nand NAND2 (N2223, N2208, N1159);
xor XOR2 (N2224, N2201, N628);
buf BUF1 (N2225, N2222);
or OR2 (N2226, N2204, N64);
nand NAND2 (N2227, N2221, N1030);
xor XOR2 (N2228, N2227, N128);
or OR3 (N2229, N2218, N1047, N868);
or OR4 (N2230, N2173, N1206, N1313, N1622);
nor NOR2 (N2231, N2220, N348);
nand NAND2 (N2232, N2228, N760);
nor NOR3 (N2233, N2226, N1161, N260);
buf BUF1 (N2234, N2230);
buf BUF1 (N2235, N2231);
xor XOR2 (N2236, N2225, N311);
or OR3 (N2237, N2229, N1642, N1185);
and AND2 (N2238, N2219, N2199);
buf BUF1 (N2239, N2236);
nor NOR3 (N2240, N2238, N2066, N56);
nand NAND3 (N2241, N2232, N2107, N1069);
buf BUF1 (N2242, N2240);
or OR2 (N2243, N2239, N2068);
not NOT1 (N2244, N2235);
buf BUF1 (N2245, N2244);
nor NOR3 (N2246, N2242, N1984, N1663);
nand NAND3 (N2247, N2237, N730, N74);
buf BUF1 (N2248, N2241);
or OR3 (N2249, N2247, N56, N1826);
xor XOR2 (N2250, N2223, N550);
buf BUF1 (N2251, N2234);
or OR2 (N2252, N2249, N2073);
not NOT1 (N2253, N2250);
nor NOR2 (N2254, N2233, N1678);
nand NAND2 (N2255, N2211, N987);
or OR4 (N2256, N2245, N28, N826, N2199);
not NOT1 (N2257, N2254);
or OR2 (N2258, N2243, N534);
xor XOR2 (N2259, N2258, N596);
buf BUF1 (N2260, N2252);
nor NOR2 (N2261, N2259, N1521);
not NOT1 (N2262, N2251);
nand NAND2 (N2263, N2256, N607);
nor NOR4 (N2264, N2246, N999, N1407, N58);
buf BUF1 (N2265, N2224);
xor XOR2 (N2266, N2253, N606);
not NOT1 (N2267, N2262);
buf BUF1 (N2268, N2257);
nand NAND4 (N2269, N2263, N396, N953, N1257);
and AND4 (N2270, N2269, N603, N785, N635);
nor NOR3 (N2271, N2265, N1436, N1193);
or OR4 (N2272, N2255, N947, N721, N178);
nor NOR3 (N2273, N2267, N1439, N1018);
not NOT1 (N2274, N2268);
buf BUF1 (N2275, N2248);
not NOT1 (N2276, N2273);
nor NOR4 (N2277, N2264, N1548, N2266, N1195);
nand NAND4 (N2278, N1372, N1415, N1074, N2275);
buf BUF1 (N2279, N992);
xor XOR2 (N2280, N2276, N1275);
nand NAND4 (N2281, N2270, N631, N918, N1314);
buf BUF1 (N2282, N2260);
nand NAND3 (N2283, N2274, N2250, N1294);
xor XOR2 (N2284, N2261, N1012);
buf BUF1 (N2285, N2278);
or OR2 (N2286, N2279, N2071);
xor XOR2 (N2287, N2281, N2106);
nand NAND4 (N2288, N2277, N1072, N101, N962);
nand NAND2 (N2289, N2280, N1280);
buf BUF1 (N2290, N2271);
nor NOR4 (N2291, N2286, N354, N1071, N1418);
not NOT1 (N2292, N2290);
buf BUF1 (N2293, N2287);
or OR3 (N2294, N2272, N1132, N393);
nor NOR2 (N2295, N2291, N1637);
nand NAND3 (N2296, N2295, N2292, N1205);
xor XOR2 (N2297, N205, N2238);
not NOT1 (N2298, N2288);
not NOT1 (N2299, N2293);
nand NAND4 (N2300, N2299, N1513, N1954, N181);
nand NAND4 (N2301, N2294, N1697, N496, N702);
nand NAND2 (N2302, N2284, N420);
buf BUF1 (N2303, N2301);
not NOT1 (N2304, N2296);
nand NAND4 (N2305, N2300, N1836, N671, N13);
nand NAND4 (N2306, N2303, N551, N2162, N1601);
not NOT1 (N2307, N2306);
nor NOR2 (N2308, N2283, N523);
or OR3 (N2309, N2289, N99, N1124);
nand NAND3 (N2310, N2298, N821, N883);
not NOT1 (N2311, N2302);
xor XOR2 (N2312, N2308, N1172);
nand NAND4 (N2313, N2309, N1717, N209, N1303);
buf BUF1 (N2314, N2307);
and AND3 (N2315, N2312, N1677, N450);
nor NOR3 (N2316, N2315, N1354, N2216);
or OR3 (N2317, N2314, N542, N726);
xor XOR2 (N2318, N2285, N1202);
nor NOR4 (N2319, N2313, N1220, N1150, N1727);
xor XOR2 (N2320, N2310, N261);
buf BUF1 (N2321, N2305);
buf BUF1 (N2322, N2321);
nand NAND2 (N2323, N2297, N396);
and AND4 (N2324, N2319, N1078, N2276, N2056);
nand NAND3 (N2325, N2320, N1315, N1950);
buf BUF1 (N2326, N2322);
buf BUF1 (N2327, N2324);
or OR4 (N2328, N2323, N1126, N2296, N547);
xor XOR2 (N2329, N2317, N1431);
nand NAND2 (N2330, N2329, N969);
or OR4 (N2331, N2304, N42, N804, N1873);
xor XOR2 (N2332, N2331, N1017);
not NOT1 (N2333, N2318);
nor NOR3 (N2334, N2326, N2150, N1298);
or OR2 (N2335, N2282, N261);
nor NOR4 (N2336, N2328, N2019, N1920, N1648);
and AND2 (N2337, N2330, N132);
nand NAND4 (N2338, N2327, N1088, N2209, N533);
nor NOR3 (N2339, N2335, N458, N1102);
and AND2 (N2340, N2325, N946);
buf BUF1 (N2341, N2339);
not NOT1 (N2342, N2334);
xor XOR2 (N2343, N2337, N345);
or OR2 (N2344, N2342, N1274);
not NOT1 (N2345, N2333);
or OR3 (N2346, N2344, N35, N187);
nand NAND4 (N2347, N2316, N906, N2252, N178);
and AND4 (N2348, N2346, N271, N581, N551);
nand NAND3 (N2349, N2345, N733, N146);
nor NOR3 (N2350, N2338, N973, N617);
buf BUF1 (N2351, N2311);
nor NOR4 (N2352, N2340, N2341, N1689, N1516);
buf BUF1 (N2353, N1704);
xor XOR2 (N2354, N2353, N2345);
xor XOR2 (N2355, N2336, N718);
nand NAND4 (N2356, N2351, N73, N127, N931);
not NOT1 (N2357, N2355);
buf BUF1 (N2358, N2354);
nor NOR3 (N2359, N2343, N1221, N410);
buf BUF1 (N2360, N2349);
or OR2 (N2361, N2356, N1976);
or OR4 (N2362, N2360, N2201, N1178, N778);
xor XOR2 (N2363, N2352, N2032);
nand NAND3 (N2364, N2357, N1645, N1998);
and AND4 (N2365, N2358, N1495, N449, N93);
or OR4 (N2366, N2365, N761, N1791, N1489);
nand NAND3 (N2367, N2361, N1315, N2128);
not NOT1 (N2368, N2348);
xor XOR2 (N2369, N2350, N1198);
not NOT1 (N2370, N2369);
and AND2 (N2371, N2370, N1620);
xor XOR2 (N2372, N2347, N1608);
xor XOR2 (N2373, N2364, N1721);
or OR3 (N2374, N2367, N14, N1023);
and AND2 (N2375, N2372, N1447);
nor NOR4 (N2376, N2362, N1585, N2111, N165);
xor XOR2 (N2377, N2363, N355);
not NOT1 (N2378, N2374);
or OR4 (N2379, N2332, N1520, N550, N1198);
buf BUF1 (N2380, N2371);
nand NAND3 (N2381, N2380, N529, N56);
or OR3 (N2382, N2376, N558, N472);
and AND4 (N2383, N2375, N1997, N2237, N266);
nand NAND2 (N2384, N2382, N1833);
or OR3 (N2385, N2381, N2011, N1770);
nor NOR2 (N2386, N2378, N2128);
nand NAND4 (N2387, N2377, N680, N1695, N801);
nor NOR2 (N2388, N2368, N441);
or OR4 (N2389, N2388, N1424, N1259, N2227);
not NOT1 (N2390, N2389);
or OR2 (N2391, N2387, N2272);
nand NAND2 (N2392, N2384, N537);
nor NOR3 (N2393, N2383, N488, N2141);
or OR4 (N2394, N2391, N523, N2358, N1719);
nand NAND2 (N2395, N2386, N1787);
xor XOR2 (N2396, N2379, N443);
nor NOR2 (N2397, N2390, N1550);
xor XOR2 (N2398, N2366, N14);
or OR3 (N2399, N2394, N446, N1208);
nand NAND3 (N2400, N2398, N761, N2235);
nor NOR2 (N2401, N2400, N2052);
nor NOR3 (N2402, N2373, N867, N2029);
nand NAND4 (N2403, N2396, N877, N430, N1231);
nor NOR4 (N2404, N2392, N2387, N2383, N1712);
nand NAND2 (N2405, N2395, N276);
xor XOR2 (N2406, N2403, N981);
and AND2 (N2407, N2393, N680);
buf BUF1 (N2408, N2401);
nand NAND4 (N2409, N2407, N2364, N1022, N549);
or OR4 (N2410, N2404, N753, N680, N1552);
and AND3 (N2411, N2399, N1151, N1980);
nand NAND4 (N2412, N2410, N1412, N440, N2016);
nor NOR4 (N2413, N2411, N2294, N2051, N726);
buf BUF1 (N2414, N2409);
xor XOR2 (N2415, N2413, N1741);
buf BUF1 (N2416, N2415);
not NOT1 (N2417, N2416);
nand NAND4 (N2418, N2385, N982, N893, N551);
buf BUF1 (N2419, N2414);
nand NAND3 (N2420, N2406, N112, N1001);
or OR4 (N2421, N2359, N807, N1503, N2336);
buf BUF1 (N2422, N2405);
buf BUF1 (N2423, N2421);
and AND2 (N2424, N2419, N1201);
buf BUF1 (N2425, N2418);
not NOT1 (N2426, N2423);
and AND2 (N2427, N2408, N137);
or OR4 (N2428, N2417, N366, N277, N779);
buf BUF1 (N2429, N2425);
nor NOR2 (N2430, N2397, N2415);
not NOT1 (N2431, N2426);
buf BUF1 (N2432, N2427);
buf BUF1 (N2433, N2402);
and AND3 (N2434, N2430, N1877, N1159);
xor XOR2 (N2435, N2429, N216);
not NOT1 (N2436, N2422);
nor NOR4 (N2437, N2433, N308, N555, N1086);
or OR3 (N2438, N2428, N310, N664);
buf BUF1 (N2439, N2436);
xor XOR2 (N2440, N2432, N2193);
nand NAND4 (N2441, N2412, N37, N1281, N753);
buf BUF1 (N2442, N2424);
and AND2 (N2443, N2439, N268);
xor XOR2 (N2444, N2434, N2293);
and AND3 (N2445, N2444, N859, N884);
nor NOR2 (N2446, N2431, N1096);
nor NOR3 (N2447, N2435, N2130, N2);
not NOT1 (N2448, N2420);
nor NOR3 (N2449, N2445, N2282, N1936);
nand NAND3 (N2450, N2448, N1433, N479);
nand NAND4 (N2451, N2446, N1884, N1942, N1120);
or OR4 (N2452, N2449, N1260, N373, N150);
and AND2 (N2453, N2450, N1431);
nor NOR3 (N2454, N2437, N1962, N1383);
buf BUF1 (N2455, N2442);
nand NAND2 (N2456, N2453, N780);
not NOT1 (N2457, N2441);
and AND2 (N2458, N2454, N2316);
and AND4 (N2459, N2438, N2135, N281, N1597);
and AND3 (N2460, N2456, N367, N676);
or OR4 (N2461, N2451, N947, N403, N1061);
or OR3 (N2462, N2460, N1104, N1612);
or OR3 (N2463, N2455, N2408, N1197);
nand NAND2 (N2464, N2461, N102);
xor XOR2 (N2465, N2452, N121);
and AND4 (N2466, N2443, N568, N930, N1572);
buf BUF1 (N2467, N2447);
and AND2 (N2468, N2465, N876);
and AND4 (N2469, N2468, N1444, N2141, N946);
nand NAND3 (N2470, N2466, N1004, N2261);
xor XOR2 (N2471, N2463, N1464);
or OR2 (N2472, N2467, N79);
nand NAND2 (N2473, N2470, N987);
not NOT1 (N2474, N2473);
not NOT1 (N2475, N2469);
xor XOR2 (N2476, N2462, N1060);
nor NOR3 (N2477, N2475, N1242, N544);
or OR2 (N2478, N2476, N1460);
nand NAND4 (N2479, N2464, N2338, N751, N709);
xor XOR2 (N2480, N2479, N1568);
nand NAND4 (N2481, N2471, N1929, N1172, N1373);
not NOT1 (N2482, N2458);
xor XOR2 (N2483, N2481, N365);
and AND2 (N2484, N2477, N884);
nand NAND4 (N2485, N2484, N796, N908, N683);
not NOT1 (N2486, N2472);
nor NOR2 (N2487, N2478, N19);
or OR2 (N2488, N2485, N1205);
buf BUF1 (N2489, N2482);
buf BUF1 (N2490, N2487);
xor XOR2 (N2491, N2490, N247);
or OR4 (N2492, N2491, N500, N1703, N595);
buf BUF1 (N2493, N2474);
and AND4 (N2494, N2493, N316, N966, N2199);
xor XOR2 (N2495, N2480, N1534);
and AND4 (N2496, N2494, N1817, N2363, N992);
nand NAND4 (N2497, N2496, N1025, N886, N805);
and AND3 (N2498, N2459, N726, N1419);
and AND3 (N2499, N2492, N2497, N1358);
or OR4 (N2500, N244, N469, N1679, N663);
nand NAND3 (N2501, N2457, N2454, N2396);
nand NAND2 (N2502, N2488, N2130);
not NOT1 (N2503, N2502);
and AND4 (N2504, N2486, N700, N346, N10);
nand NAND2 (N2505, N2499, N2189);
nor NOR4 (N2506, N2498, N2015, N765, N1605);
not NOT1 (N2507, N2500);
or OR4 (N2508, N2501, N491, N1381, N2251);
xor XOR2 (N2509, N2504, N2262);
nor NOR4 (N2510, N2489, N1281, N1789, N1731);
and AND4 (N2511, N2510, N38, N1339, N1110);
not NOT1 (N2512, N2503);
or OR2 (N2513, N2440, N298);
buf BUF1 (N2514, N2513);
xor XOR2 (N2515, N2514, N1676);
or OR4 (N2516, N2495, N501, N1726, N1192);
nor NOR3 (N2517, N2515, N767, N2400);
buf BUF1 (N2518, N2516);
xor XOR2 (N2519, N2483, N2099);
nor NOR4 (N2520, N2511, N149, N1754, N1144);
and AND4 (N2521, N2508, N2025, N472, N1942);
or OR4 (N2522, N2518, N2234, N1346, N2485);
buf BUF1 (N2523, N2520);
not NOT1 (N2524, N2521);
xor XOR2 (N2525, N2512, N2518);
nand NAND4 (N2526, N2507, N958, N696, N1426);
or OR4 (N2527, N2526, N2197, N2246, N985);
or OR3 (N2528, N2527, N543, N2371);
buf BUF1 (N2529, N2506);
nand NAND3 (N2530, N2524, N2384, N614);
or OR3 (N2531, N2522, N1801, N1617);
not NOT1 (N2532, N2505);
not NOT1 (N2533, N2517);
or OR2 (N2534, N2519, N1942);
or OR3 (N2535, N2533, N1017, N296);
nand NAND3 (N2536, N2528, N43, N238);
nand NAND2 (N2537, N2536, N2282);
or OR4 (N2538, N2535, N536, N1473, N1627);
xor XOR2 (N2539, N2525, N1560);
nand NAND3 (N2540, N2531, N717, N2496);
and AND2 (N2541, N2534, N2187);
or OR3 (N2542, N2540, N2480, N676);
and AND3 (N2543, N2539, N1915, N840);
nand NAND4 (N2544, N2509, N2247, N498, N273);
not NOT1 (N2545, N2541);
buf BUF1 (N2546, N2543);
xor XOR2 (N2547, N2530, N761);
nand NAND2 (N2548, N2546, N322);
buf BUF1 (N2549, N2544);
buf BUF1 (N2550, N2532);
nor NOR3 (N2551, N2548, N1843, N720);
not NOT1 (N2552, N2551);
nand NAND3 (N2553, N2550, N2256, N934);
nor NOR4 (N2554, N2547, N305, N116, N2501);
and AND3 (N2555, N2523, N1204, N1938);
nor NOR2 (N2556, N2554, N1077);
nor NOR4 (N2557, N2553, N2158, N1128, N924);
xor XOR2 (N2558, N2549, N2308);
nand NAND4 (N2559, N2558, N1907, N1029, N285);
xor XOR2 (N2560, N2555, N2157);
xor XOR2 (N2561, N2529, N2188);
not NOT1 (N2562, N2537);
buf BUF1 (N2563, N2561);
or OR2 (N2564, N2562, N531);
xor XOR2 (N2565, N2563, N235);
nor NOR4 (N2566, N2552, N2164, N2177, N817);
buf BUF1 (N2567, N2542);
nor NOR4 (N2568, N2560, N548, N511, N780);
and AND2 (N2569, N2559, N1320);
not NOT1 (N2570, N2565);
or OR4 (N2571, N2570, N1272, N1888, N754);
nand NAND4 (N2572, N2556, N197, N2357, N1744);
buf BUF1 (N2573, N2545);
and AND2 (N2574, N2567, N1345);
or OR2 (N2575, N2566, N1040);
xor XOR2 (N2576, N2538, N2244);
nor NOR3 (N2577, N2574, N714, N44);
nor NOR4 (N2578, N2564, N24, N1925, N2460);
nand NAND4 (N2579, N2573, N979, N1082, N1285);
xor XOR2 (N2580, N2579, N294);
and AND2 (N2581, N2576, N155);
nor NOR2 (N2582, N2580, N597);
not NOT1 (N2583, N2572);
and AND4 (N2584, N2557, N1922, N461, N435);
and AND2 (N2585, N2584, N244);
buf BUF1 (N2586, N2585);
and AND2 (N2587, N2583, N967);
and AND2 (N2588, N2575, N1388);
and AND3 (N2589, N2587, N1744, N501);
xor XOR2 (N2590, N2588, N802);
nand NAND3 (N2591, N2571, N1669, N813);
or OR3 (N2592, N2582, N75, N1286);
buf BUF1 (N2593, N2586);
or OR3 (N2594, N2569, N1453, N620);
nand NAND4 (N2595, N2581, N1200, N1933, N2164);
and AND2 (N2596, N2595, N1187);
xor XOR2 (N2597, N2590, N1113);
or OR2 (N2598, N2592, N808);
or OR3 (N2599, N2598, N1397, N1705);
nor NOR2 (N2600, N2591, N103);
buf BUF1 (N2601, N2577);
xor XOR2 (N2602, N2597, N408);
buf BUF1 (N2603, N2599);
nand NAND2 (N2604, N2600, N399);
buf BUF1 (N2605, N2601);
xor XOR2 (N2606, N2596, N1140);
nor NOR3 (N2607, N2605, N1716, N2448);
buf BUF1 (N2608, N2568);
xor XOR2 (N2609, N2603, N879);
nand NAND2 (N2610, N2594, N620);
nor NOR3 (N2611, N2610, N1219, N723);
xor XOR2 (N2612, N2589, N2074);
and AND2 (N2613, N2608, N213);
or OR3 (N2614, N2612, N385, N780);
and AND3 (N2615, N2613, N517, N1763);
buf BUF1 (N2616, N2602);
not NOT1 (N2617, N2614);
not NOT1 (N2618, N2609);
nand NAND3 (N2619, N2618, N68, N2002);
and AND3 (N2620, N2606, N1934, N304);
buf BUF1 (N2621, N2593);
nand NAND2 (N2622, N2621, N741);
not NOT1 (N2623, N2578);
buf BUF1 (N2624, N2617);
nand NAND2 (N2625, N2611, N1056);
and AND3 (N2626, N2604, N1947, N277);
not NOT1 (N2627, N2620);
or OR3 (N2628, N2607, N962, N951);
nor NOR4 (N2629, N2615, N1985, N83, N1606);
or OR4 (N2630, N2616, N1136, N1111, N10);
nor NOR2 (N2631, N2627, N2107);
xor XOR2 (N2632, N2623, N752);
nor NOR4 (N2633, N2628, N1162, N2370, N995);
xor XOR2 (N2634, N2626, N599);
nand NAND3 (N2635, N2633, N319, N276);
xor XOR2 (N2636, N2635, N2048);
not NOT1 (N2637, N2625);
not NOT1 (N2638, N2637);
and AND3 (N2639, N2630, N203, N1347);
nand NAND2 (N2640, N2638, N140);
xor XOR2 (N2641, N2622, N2380);
not NOT1 (N2642, N2636);
or OR3 (N2643, N2639, N2178, N1174);
buf BUF1 (N2644, N2632);
buf BUF1 (N2645, N2640);
xor XOR2 (N2646, N2634, N2498);
nand NAND4 (N2647, N2619, N2530, N2113, N735);
nand NAND4 (N2648, N2646, N2164, N2638, N914);
nand NAND3 (N2649, N2647, N1249, N405);
xor XOR2 (N2650, N2648, N1387);
and AND3 (N2651, N2629, N437, N2397);
xor XOR2 (N2652, N2650, N338);
or OR4 (N2653, N2631, N1799, N1759, N255);
buf BUF1 (N2654, N2644);
not NOT1 (N2655, N2624);
and AND4 (N2656, N2642, N222, N2023, N322);
and AND2 (N2657, N2641, N739);
buf BUF1 (N2658, N2654);
nor NOR3 (N2659, N2656, N1047, N37);
nor NOR4 (N2660, N2655, N421, N2473, N51);
buf BUF1 (N2661, N2659);
nand NAND3 (N2662, N2649, N1902, N1883);
nor NOR4 (N2663, N2661, N426, N1307, N296);
not NOT1 (N2664, N2662);
nor NOR3 (N2665, N2664, N1281, N2407);
nor NOR2 (N2666, N2660, N527);
or OR2 (N2667, N2657, N2300);
and AND3 (N2668, N2665, N1070, N504);
nor NOR3 (N2669, N2663, N1342, N2624);
or OR3 (N2670, N2669, N1843, N1691);
buf BUF1 (N2671, N2645);
xor XOR2 (N2672, N2668, N74);
not NOT1 (N2673, N2643);
or OR4 (N2674, N2671, N661, N433, N950);
and AND3 (N2675, N2670, N750, N1982);
xor XOR2 (N2676, N2666, N455);
buf BUF1 (N2677, N2667);
and AND4 (N2678, N2676, N2192, N2578, N247);
or OR2 (N2679, N2674, N2536);
and AND3 (N2680, N2672, N1855, N1352);
not NOT1 (N2681, N2652);
not NOT1 (N2682, N2653);
nand NAND4 (N2683, N2681, N865, N286, N2409);
nand NAND3 (N2684, N2675, N2420, N1579);
not NOT1 (N2685, N2679);
buf BUF1 (N2686, N2651);
buf BUF1 (N2687, N2658);
not NOT1 (N2688, N2680);
or OR3 (N2689, N2685, N135, N561);
buf BUF1 (N2690, N2673);
nor NOR4 (N2691, N2687, N640, N1787, N1819);
not NOT1 (N2692, N2677);
nand NAND3 (N2693, N2690, N2064, N2689);
buf BUF1 (N2694, N663);
not NOT1 (N2695, N2683);
nand NAND2 (N2696, N2682, N69);
or OR3 (N2697, N2692, N1711, N2269);
or OR3 (N2698, N2686, N1885, N2309);
not NOT1 (N2699, N2697);
not NOT1 (N2700, N2688);
not NOT1 (N2701, N2698);
xor XOR2 (N2702, N2684, N734);
and AND4 (N2703, N2694, N325, N1317, N1026);
not NOT1 (N2704, N2701);
nand NAND2 (N2705, N2696, N2389);
nand NAND3 (N2706, N2691, N2435, N2295);
not NOT1 (N2707, N2699);
not NOT1 (N2708, N2693);
nor NOR3 (N2709, N2706, N473, N555);
xor XOR2 (N2710, N2709, N2241);
nand NAND3 (N2711, N2707, N1488, N1724);
nor NOR2 (N2712, N2695, N1335);
or OR4 (N2713, N2712, N2174, N76, N977);
xor XOR2 (N2714, N2713, N2700);
or OR3 (N2715, N1936, N667, N733);
buf BUF1 (N2716, N2710);
nand NAND2 (N2717, N2678, N1609);
not NOT1 (N2718, N2703);
and AND3 (N2719, N2714, N119, N1264);
xor XOR2 (N2720, N2717, N1592);
not NOT1 (N2721, N2708);
not NOT1 (N2722, N2705);
not NOT1 (N2723, N2722);
xor XOR2 (N2724, N2720, N2147);
and AND2 (N2725, N2716, N622);
nor NOR2 (N2726, N2711, N175);
nand NAND4 (N2727, N2704, N419, N1540, N296);
not NOT1 (N2728, N2721);
and AND2 (N2729, N2715, N2533);
buf BUF1 (N2730, N2718);
or OR2 (N2731, N2724, N2431);
nor NOR3 (N2732, N2723, N1461, N1677);
xor XOR2 (N2733, N2730, N2419);
xor XOR2 (N2734, N2726, N1215);
and AND3 (N2735, N2732, N1249, N785);
or OR3 (N2736, N2719, N677, N902);
nor NOR4 (N2737, N2733, N344, N594, N665);
buf BUF1 (N2738, N2727);
or OR3 (N2739, N2725, N2556, N2038);
nor NOR3 (N2740, N2737, N2446, N1318);
and AND3 (N2741, N2739, N1628, N1862);
and AND3 (N2742, N2736, N777, N746);
or OR3 (N2743, N2735, N346, N725);
or OR3 (N2744, N2741, N890, N2255);
nor NOR3 (N2745, N2738, N1600, N2493);
not NOT1 (N2746, N2740);
nor NOR4 (N2747, N2734, N1656, N2259, N2306);
nand NAND3 (N2748, N2743, N98, N1765);
or OR4 (N2749, N2731, N2286, N815, N2322);
nand NAND4 (N2750, N2749, N2410, N165, N1277);
buf BUF1 (N2751, N2745);
not NOT1 (N2752, N2751);
nand NAND2 (N2753, N2742, N1808);
nor NOR4 (N2754, N2746, N933, N1987, N703);
buf BUF1 (N2755, N2750);
nor NOR2 (N2756, N2755, N1283);
xor XOR2 (N2757, N2728, N890);
and AND2 (N2758, N2756, N2119);
not NOT1 (N2759, N2753);
xor XOR2 (N2760, N2758, N582);
and AND2 (N2761, N2729, N865);
nand NAND4 (N2762, N2761, N718, N1900, N1317);
xor XOR2 (N2763, N2748, N1716);
nor NOR4 (N2764, N2760, N573, N2106, N1230);
or OR3 (N2765, N2757, N1906, N47);
and AND4 (N2766, N2702, N1710, N2278, N1286);
buf BUF1 (N2767, N2744);
not NOT1 (N2768, N2759);
buf BUF1 (N2769, N2766);
nor NOR3 (N2770, N2768, N733, N395);
xor XOR2 (N2771, N2770, N2396);
xor XOR2 (N2772, N2769, N1487);
or OR2 (N2773, N2765, N181);
nand NAND3 (N2774, N2772, N1014, N2032);
nand NAND4 (N2775, N2762, N304, N2222, N632);
xor XOR2 (N2776, N2775, N147);
or OR2 (N2777, N2774, N675);
xor XOR2 (N2778, N2764, N1321);
nand NAND4 (N2779, N2747, N169, N1632, N1816);
nand NAND4 (N2780, N2773, N1962, N1262, N2090);
xor XOR2 (N2781, N2780, N1289);
nor NOR4 (N2782, N2779, N2368, N2578, N1683);
xor XOR2 (N2783, N2767, N520);
not NOT1 (N2784, N2754);
or OR3 (N2785, N2783, N2360, N2691);
xor XOR2 (N2786, N2785, N2166);
xor XOR2 (N2787, N2752, N350);
nand NAND4 (N2788, N2784, N1179, N1503, N2104);
or OR2 (N2789, N2788, N2420);
nor NOR3 (N2790, N2787, N901, N2336);
nor NOR2 (N2791, N2786, N113);
nor NOR3 (N2792, N2790, N1970, N943);
buf BUF1 (N2793, N2782);
not NOT1 (N2794, N2781);
xor XOR2 (N2795, N2778, N2288);
nand NAND4 (N2796, N2793, N407, N1435, N2784);
xor XOR2 (N2797, N2777, N1547);
nand NAND2 (N2798, N2796, N1034);
buf BUF1 (N2799, N2776);
or OR4 (N2800, N2799, N274, N2498, N2432);
buf BUF1 (N2801, N2789);
and AND4 (N2802, N2792, N2474, N415, N645);
or OR2 (N2803, N2801, N1208);
nand NAND4 (N2804, N2771, N2785, N825, N969);
buf BUF1 (N2805, N2795);
or OR2 (N2806, N2797, N2108);
or OR2 (N2807, N2805, N1847);
and AND2 (N2808, N2791, N1074);
buf BUF1 (N2809, N2763);
nor NOR4 (N2810, N2798, N2403, N1735, N1558);
nor NOR2 (N2811, N2809, N2722);
nor NOR4 (N2812, N2802, N2278, N80, N1920);
nor NOR2 (N2813, N2810, N1396);
buf BUF1 (N2814, N2803);
nor NOR4 (N2815, N2794, N2313, N632, N679);
not NOT1 (N2816, N2813);
nor NOR4 (N2817, N2806, N2085, N2408, N909);
and AND2 (N2818, N2817, N2599);
not NOT1 (N2819, N2812);
not NOT1 (N2820, N2804);
nand NAND2 (N2821, N2814, N359);
xor XOR2 (N2822, N2811, N2619);
and AND2 (N2823, N2822, N1743);
xor XOR2 (N2824, N2816, N2330);
xor XOR2 (N2825, N2821, N1178);
xor XOR2 (N2826, N2807, N46);
nand NAND4 (N2827, N2818, N907, N126, N137);
or OR3 (N2828, N2826, N7, N203);
not NOT1 (N2829, N2825);
or OR3 (N2830, N2823, N39, N1490);
xor XOR2 (N2831, N2830, N128);
xor XOR2 (N2832, N2824, N1341);
and AND3 (N2833, N2827, N2376, N984);
nor NOR3 (N2834, N2815, N2298, N287);
not NOT1 (N2835, N2820);
nor NOR3 (N2836, N2800, N273, N271);
xor XOR2 (N2837, N2831, N1089);
not NOT1 (N2838, N2835);
buf BUF1 (N2839, N2834);
nor NOR4 (N2840, N2836, N1915, N2148, N2321);
nand NAND3 (N2841, N2839, N830, N2801);
buf BUF1 (N2842, N2828);
and AND3 (N2843, N2833, N2610, N1825);
and AND2 (N2844, N2843, N1686);
or OR2 (N2845, N2837, N654);
nor NOR2 (N2846, N2840, N1315);
xor XOR2 (N2847, N2846, N2337);
or OR2 (N2848, N2847, N2643);
or OR3 (N2849, N2832, N372, N2592);
xor XOR2 (N2850, N2842, N812);
nand NAND4 (N2851, N2849, N2156, N176, N223);
nand NAND4 (N2852, N2841, N302, N1924, N294);
not NOT1 (N2853, N2838);
buf BUF1 (N2854, N2808);
not NOT1 (N2855, N2852);
buf BUF1 (N2856, N2829);
nand NAND4 (N2857, N2845, N1284, N1465, N616);
not NOT1 (N2858, N2853);
xor XOR2 (N2859, N2858, N2047);
and AND3 (N2860, N2854, N2711, N2083);
and AND4 (N2861, N2856, N1495, N716, N1798);
nand NAND2 (N2862, N2819, N2072);
nand NAND3 (N2863, N2850, N1097, N700);
xor XOR2 (N2864, N2857, N840);
or OR2 (N2865, N2862, N2256);
buf BUF1 (N2866, N2851);
not NOT1 (N2867, N2864);
or OR3 (N2868, N2844, N1177, N2572);
and AND4 (N2869, N2866, N1092, N1604, N1282);
buf BUF1 (N2870, N2865);
xor XOR2 (N2871, N2859, N243);
buf BUF1 (N2872, N2860);
not NOT1 (N2873, N2869);
and AND3 (N2874, N2863, N1639, N1171);
or OR2 (N2875, N2848, N2403);
and AND3 (N2876, N2874, N1693, N1745);
nor NOR2 (N2877, N2855, N2227);
nor NOR3 (N2878, N2876, N1991, N1670);
nor NOR2 (N2879, N2861, N2455);
nor NOR4 (N2880, N2878, N2350, N208, N803);
buf BUF1 (N2881, N2879);
not NOT1 (N2882, N2875);
nor NOR3 (N2883, N2871, N1526, N2352);
nand NAND4 (N2884, N2868, N2344, N2150, N403);
or OR2 (N2885, N2881, N1947);
not NOT1 (N2886, N2870);
not NOT1 (N2887, N2867);
buf BUF1 (N2888, N2872);
xor XOR2 (N2889, N2880, N658);
buf BUF1 (N2890, N2885);
and AND3 (N2891, N2890, N2196, N204);
and AND2 (N2892, N2883, N815);
nand NAND4 (N2893, N2892, N861, N290, N411);
buf BUF1 (N2894, N2889);
xor XOR2 (N2895, N2894, N2862);
buf BUF1 (N2896, N2891);
nand NAND4 (N2897, N2888, N550, N2505, N1724);
nand NAND3 (N2898, N2895, N205, N1736);
not NOT1 (N2899, N2873);
buf BUF1 (N2900, N2896);
nand NAND2 (N2901, N2877, N520);
nand NAND3 (N2902, N2882, N591, N1626);
and AND2 (N2903, N2902, N1822);
or OR4 (N2904, N2893, N2862, N2230, N426);
or OR2 (N2905, N2904, N1402);
buf BUF1 (N2906, N2897);
and AND4 (N2907, N2886, N933, N2271, N830);
nor NOR4 (N2908, N2884, N684, N1700, N2703);
not NOT1 (N2909, N2887);
and AND2 (N2910, N2901, N2137);
xor XOR2 (N2911, N2910, N2586);
or OR3 (N2912, N2903, N1464, N2476);
and AND4 (N2913, N2907, N561, N1270, N568);
buf BUF1 (N2914, N2908);
not NOT1 (N2915, N2898);
and AND4 (N2916, N2911, N857, N850, N1265);
xor XOR2 (N2917, N2909, N491);
xor XOR2 (N2918, N2899, N1529);
xor XOR2 (N2919, N2918, N2718);
nor NOR3 (N2920, N2915, N1547, N2149);
nand NAND3 (N2921, N2916, N2771, N1037);
nand NAND3 (N2922, N2919, N1948, N224);
buf BUF1 (N2923, N2917);
nor NOR3 (N2924, N2921, N594, N2654);
xor XOR2 (N2925, N2924, N2162);
and AND3 (N2926, N2920, N1410, N365);
xor XOR2 (N2927, N2914, N597);
xor XOR2 (N2928, N2925, N1323);
nand NAND3 (N2929, N2923, N318, N2567);
or OR2 (N2930, N2922, N2149);
or OR2 (N2931, N2905, N1169);
or OR4 (N2932, N2912, N532, N1093, N2624);
nand NAND4 (N2933, N2930, N1686, N2166, N1762);
buf BUF1 (N2934, N2932);
and AND3 (N2935, N2900, N1035, N1328);
not NOT1 (N2936, N2933);
or OR2 (N2937, N2934, N2609);
xor XOR2 (N2938, N2937, N435);
not NOT1 (N2939, N2906);
or OR2 (N2940, N2926, N2733);
or OR4 (N2941, N2935, N1769, N1245, N858);
or OR4 (N2942, N2931, N2125, N2489, N1438);
or OR2 (N2943, N2942, N1449);
or OR3 (N2944, N2929, N2554, N1488);
buf BUF1 (N2945, N2943);
and AND4 (N2946, N2945, N2937, N1219, N1592);
not NOT1 (N2947, N2913);
buf BUF1 (N2948, N2947);
not NOT1 (N2949, N2944);
nand NAND3 (N2950, N2948, N1468, N722);
or OR4 (N2951, N2936, N1624, N983, N131);
or OR3 (N2952, N2939, N1691, N839);
xor XOR2 (N2953, N2950, N1278);
xor XOR2 (N2954, N2951, N2761);
buf BUF1 (N2955, N2946);
xor XOR2 (N2956, N2927, N2049);
not NOT1 (N2957, N2952);
nand NAND4 (N2958, N2928, N2788, N2256, N2291);
xor XOR2 (N2959, N2955, N2413);
or OR4 (N2960, N2938, N696, N908, N2481);
buf BUF1 (N2961, N2959);
not NOT1 (N2962, N2949);
nand NAND2 (N2963, N2954, N2075);
buf BUF1 (N2964, N2941);
not NOT1 (N2965, N2956);
buf BUF1 (N2966, N2963);
buf BUF1 (N2967, N2961);
and AND3 (N2968, N2965, N1608, N2623);
not NOT1 (N2969, N2962);
not NOT1 (N2970, N2958);
nor NOR2 (N2971, N2967, N21);
nand NAND4 (N2972, N2953, N488, N489, N2175);
nor NOR2 (N2973, N2957, N1416);
xor XOR2 (N2974, N2964, N1120);
or OR2 (N2975, N2940, N521);
xor XOR2 (N2976, N2974, N853);
nor NOR4 (N2977, N2966, N347, N334, N2390);
xor XOR2 (N2978, N2969, N289);
nor NOR4 (N2979, N2977, N542, N2797, N650);
nand NAND4 (N2980, N2971, N1839, N2609, N2482);
and AND2 (N2981, N2972, N702);
not NOT1 (N2982, N2978);
and AND3 (N2983, N2979, N2246, N1380);
nor NOR3 (N2984, N2973, N1333, N2378);
xor XOR2 (N2985, N2981, N1478);
or OR2 (N2986, N2984, N2350);
or OR2 (N2987, N2983, N235);
xor XOR2 (N2988, N2976, N408);
nand NAND4 (N2989, N2985, N856, N2072, N69);
nand NAND3 (N2990, N2989, N580, N1980);
xor XOR2 (N2991, N2960, N1632);
buf BUF1 (N2992, N2975);
nor NOR3 (N2993, N2980, N942, N2542);
or OR4 (N2994, N2988, N746, N1937, N143);
not NOT1 (N2995, N2968);
nor NOR2 (N2996, N2993, N54);
and AND4 (N2997, N2996, N2424, N157, N1244);
xor XOR2 (N2998, N2987, N1933);
or OR4 (N2999, N2991, N1386, N921, N2136);
nand NAND2 (N3000, N2998, N2556);
or OR3 (N3001, N2992, N1041, N252);
xor XOR2 (N3002, N2970, N785);
buf BUF1 (N3003, N2982);
or OR2 (N3004, N2986, N1641);
buf BUF1 (N3005, N3003);
xor XOR2 (N3006, N2995, N2497);
buf BUF1 (N3007, N3001);
buf BUF1 (N3008, N2994);
xor XOR2 (N3009, N2999, N1691);
buf BUF1 (N3010, N3000);
nand NAND2 (N3011, N3006, N883);
buf BUF1 (N3012, N3010);
nor NOR2 (N3013, N3005, N1849);
xor XOR2 (N3014, N3013, N872);
and AND4 (N3015, N3014, N1637, N2248, N1222);
or OR3 (N3016, N3009, N2509, N1660);
or OR3 (N3017, N3016, N285, N1369);
and AND3 (N3018, N3015, N2111, N2122);
and AND2 (N3019, N2990, N823);
nor NOR4 (N3020, N3004, N2267, N539, N2862);
and AND3 (N3021, N3008, N798, N2077);
and AND3 (N3022, N3012, N1942, N1709);
nor NOR4 (N3023, N3019, N1957, N1131, N369);
or OR2 (N3024, N3007, N1767);
xor XOR2 (N3025, N3023, N489);
xor XOR2 (N3026, N3011, N2710);
buf BUF1 (N3027, N3024);
nand NAND2 (N3028, N3018, N2952);
xor XOR2 (N3029, N3025, N3020);
and AND3 (N3030, N2828, N2007, N177);
xor XOR2 (N3031, N3030, N1081);
or OR2 (N3032, N3028, N2142);
or OR2 (N3033, N3002, N1578);
buf BUF1 (N3034, N3017);
and AND2 (N3035, N3033, N1307);
xor XOR2 (N3036, N3022, N2678);
xor XOR2 (N3037, N3031, N2966);
xor XOR2 (N3038, N3029, N995);
buf BUF1 (N3039, N3021);
not NOT1 (N3040, N3026);
and AND2 (N3041, N2997, N213);
nor NOR4 (N3042, N3034, N729, N1224, N128);
and AND3 (N3043, N3039, N1837, N2518);
or OR2 (N3044, N3041, N1542);
not NOT1 (N3045, N3043);
nor NOR4 (N3046, N3036, N1922, N2730, N142);
and AND2 (N3047, N3035, N843);
nor NOR3 (N3048, N3042, N698, N147);
nand NAND4 (N3049, N3044, N1439, N787, N2261);
nor NOR2 (N3050, N3049, N2975);
xor XOR2 (N3051, N3050, N2041);
buf BUF1 (N3052, N3051);
and AND3 (N3053, N3037, N887, N1719);
buf BUF1 (N3054, N3040);
nand NAND2 (N3055, N3047, N2917);
or OR2 (N3056, N3055, N1212);
buf BUF1 (N3057, N3038);
and AND3 (N3058, N3054, N676, N2926);
nand NAND4 (N3059, N3032, N3017, N1635, N1754);
not NOT1 (N3060, N3046);
nor NOR2 (N3061, N3053, N2233);
buf BUF1 (N3062, N3059);
xor XOR2 (N3063, N3061, N1075);
or OR2 (N3064, N3048, N1822);
and AND4 (N3065, N3052, N623, N2345, N2730);
buf BUF1 (N3066, N3057);
buf BUF1 (N3067, N3056);
buf BUF1 (N3068, N3027);
xor XOR2 (N3069, N3068, N1214);
not NOT1 (N3070, N3062);
xor XOR2 (N3071, N3063, N859);
not NOT1 (N3072, N3065);
or OR4 (N3073, N3072, N1099, N3056, N2691);
and AND2 (N3074, N3070, N1444);
not NOT1 (N3075, N3045);
xor XOR2 (N3076, N3075, N2712);
not NOT1 (N3077, N3071);
not NOT1 (N3078, N3067);
or OR2 (N3079, N3064, N2746);
or OR3 (N3080, N3078, N1561, N1717);
and AND4 (N3081, N3069, N2389, N1139, N2456);
or OR2 (N3082, N3066, N1203);
nor NOR4 (N3083, N3076, N138, N1459, N390);
buf BUF1 (N3084, N3080);
buf BUF1 (N3085, N3084);
buf BUF1 (N3086, N3083);
nor NOR4 (N3087, N3085, N2038, N1374, N1329);
and AND4 (N3088, N3074, N10, N801, N2175);
xor XOR2 (N3089, N3073, N2052);
not NOT1 (N3090, N3087);
xor XOR2 (N3091, N3079, N1045);
not NOT1 (N3092, N3081);
nand NAND3 (N3093, N3058, N270, N1150);
and AND3 (N3094, N3090, N788, N1610);
or OR2 (N3095, N3094, N2198);
nand NAND3 (N3096, N3095, N465, N910);
nor NOR4 (N3097, N3088, N1313, N12, N868);
and AND3 (N3098, N3082, N112, N1086);
nor NOR3 (N3099, N3089, N1498, N2543);
and AND4 (N3100, N3060, N1700, N736, N1431);
and AND4 (N3101, N3093, N1600, N921, N2595);
nor NOR2 (N3102, N3096, N1584);
not NOT1 (N3103, N3099);
nor NOR2 (N3104, N3077, N2438);
not NOT1 (N3105, N3086);
not NOT1 (N3106, N3097);
buf BUF1 (N3107, N3102);
xor XOR2 (N3108, N3091, N2637);
nor NOR2 (N3109, N3107, N1449);
buf BUF1 (N3110, N3106);
or OR4 (N3111, N3103, N500, N2659, N1423);
buf BUF1 (N3112, N3098);
buf BUF1 (N3113, N3104);
xor XOR2 (N3114, N3113, N750);
and AND3 (N3115, N3101, N2679, N2193);
nor NOR2 (N3116, N3111, N1983);
nor NOR2 (N3117, N3112, N2646);
nor NOR2 (N3118, N3105, N2063);
nor NOR4 (N3119, N3117, N757, N1204, N2313);
and AND3 (N3120, N3092, N2887, N2256);
buf BUF1 (N3121, N3109);
nand NAND2 (N3122, N3110, N2428);
nand NAND4 (N3123, N3118, N875, N578, N795);
buf BUF1 (N3124, N3122);
xor XOR2 (N3125, N3123, N1066);
xor XOR2 (N3126, N3121, N1634);
nand NAND4 (N3127, N3124, N1023, N7, N1973);
nor NOR2 (N3128, N3126, N2597);
not NOT1 (N3129, N3120);
not NOT1 (N3130, N3129);
buf BUF1 (N3131, N3119);
and AND4 (N3132, N3128, N1638, N1977, N1490);
xor XOR2 (N3133, N3116, N2410);
nand NAND4 (N3134, N3127, N1833, N1305, N432);
not NOT1 (N3135, N3115);
nand NAND3 (N3136, N3114, N1954, N3109);
buf BUF1 (N3137, N3134);
and AND3 (N3138, N3130, N2892, N2942);
nand NAND3 (N3139, N3125, N471, N1280);
nand NAND2 (N3140, N3135, N59);
nand NAND2 (N3141, N3133, N2454);
buf BUF1 (N3142, N3137);
not NOT1 (N3143, N3100);
nand NAND2 (N3144, N3142, N2799);
xor XOR2 (N3145, N3143, N1263);
nand NAND3 (N3146, N3136, N1043, N547);
nor NOR3 (N3147, N3108, N2757, N1680);
and AND3 (N3148, N3146, N1886, N2589);
not NOT1 (N3149, N3141);
or OR2 (N3150, N3144, N475);
xor XOR2 (N3151, N3150, N1583);
nor NOR2 (N3152, N3131, N2266);
nand NAND3 (N3153, N3145, N724, N2903);
xor XOR2 (N3154, N3153, N1618);
not NOT1 (N3155, N3151);
buf BUF1 (N3156, N3132);
buf BUF1 (N3157, N3140);
nand NAND2 (N3158, N3139, N899);
nor NOR4 (N3159, N3149, N628, N1490, N2909);
buf BUF1 (N3160, N3138);
and AND4 (N3161, N3152, N612, N1077, N59);
not NOT1 (N3162, N3159);
buf BUF1 (N3163, N3148);
xor XOR2 (N3164, N3160, N260);
xor XOR2 (N3165, N3162, N1973);
or OR3 (N3166, N3154, N2514, N2103);
or OR4 (N3167, N3161, N2294, N204, N2850);
nor NOR4 (N3168, N3167, N772, N542, N1039);
xor XOR2 (N3169, N3158, N799);
nor NOR3 (N3170, N3157, N382, N2454);
nand NAND3 (N3171, N3155, N2518, N2177);
xor XOR2 (N3172, N3171, N1478);
nor NOR3 (N3173, N3156, N1082, N2432);
nor NOR2 (N3174, N3164, N1682);
buf BUF1 (N3175, N3147);
nand NAND3 (N3176, N3165, N2084, N1740);
and AND2 (N3177, N3170, N354);
buf BUF1 (N3178, N3173);
or OR4 (N3179, N3174, N2743, N1335, N1854);
nand NAND3 (N3180, N3169, N1797, N1641);
nor NOR3 (N3181, N3172, N1978, N682);
buf BUF1 (N3182, N3177);
xor XOR2 (N3183, N3180, N382);
or OR3 (N3184, N3166, N1123, N2547);
nor NOR2 (N3185, N3179, N2617);
nand NAND2 (N3186, N3185, N150);
nor NOR4 (N3187, N3183, N1742, N1395, N2028);
or OR3 (N3188, N3178, N2549, N1853);
or OR2 (N3189, N3168, N1746);
buf BUF1 (N3190, N3182);
and AND4 (N3191, N3163, N2817, N1390, N1093);
buf BUF1 (N3192, N3175);
and AND4 (N3193, N3192, N697, N3133, N2116);
and AND4 (N3194, N3190, N2812, N2121, N1187);
nor NOR2 (N3195, N3193, N1059);
or OR2 (N3196, N3187, N582);
or OR3 (N3197, N3188, N640, N2902);
not NOT1 (N3198, N3181);
xor XOR2 (N3199, N3198, N211);
xor XOR2 (N3200, N3194, N2777);
buf BUF1 (N3201, N3189);
nor NOR2 (N3202, N3197, N2737);
xor XOR2 (N3203, N3200, N3068);
not NOT1 (N3204, N3201);
buf BUF1 (N3205, N3196);
not NOT1 (N3206, N3191);
and AND3 (N3207, N3199, N1769, N1530);
or OR3 (N3208, N3207, N2141, N3194);
and AND2 (N3209, N3186, N1722);
not NOT1 (N3210, N3203);
and AND3 (N3211, N3209, N3156, N1861);
xor XOR2 (N3212, N3208, N1891);
not NOT1 (N3213, N3211);
or OR2 (N3214, N3213, N2985);
or OR2 (N3215, N3176, N242);
and AND3 (N3216, N3184, N2755, N3012);
nor NOR4 (N3217, N3202, N2047, N72, N1563);
buf BUF1 (N3218, N3217);
nor NOR4 (N3219, N3206, N2497, N1225, N731);
and AND4 (N3220, N3210, N943, N2745, N43);
xor XOR2 (N3221, N3212, N2174);
nor NOR2 (N3222, N3205, N2727);
buf BUF1 (N3223, N3222);
buf BUF1 (N3224, N3215);
buf BUF1 (N3225, N3221);
buf BUF1 (N3226, N3195);
xor XOR2 (N3227, N3204, N3137);
xor XOR2 (N3228, N3224, N141);
not NOT1 (N3229, N3227);
nor NOR3 (N3230, N3228, N2851, N2889);
nand NAND2 (N3231, N3219, N2812);
buf BUF1 (N3232, N3218);
nor NOR3 (N3233, N3220, N1583, N2237);
nor NOR3 (N3234, N3225, N174, N2902);
buf BUF1 (N3235, N3232);
and AND3 (N3236, N3223, N1743, N2851);
nand NAND4 (N3237, N3233, N2393, N551, N120);
not NOT1 (N3238, N3230);
nor NOR3 (N3239, N3237, N149, N209);
not NOT1 (N3240, N3231);
not NOT1 (N3241, N3236);
nor NOR4 (N3242, N3240, N1319, N57, N560);
buf BUF1 (N3243, N3238);
buf BUF1 (N3244, N3235);
xor XOR2 (N3245, N3242, N1091);
not NOT1 (N3246, N3226);
or OR2 (N3247, N3245, N1234);
or OR3 (N3248, N3243, N644, N1305);
nand NAND3 (N3249, N3246, N715, N2107);
and AND3 (N3250, N3234, N279, N1071);
xor XOR2 (N3251, N3241, N485);
buf BUF1 (N3252, N3239);
and AND4 (N3253, N3244, N2014, N2733, N2525);
xor XOR2 (N3254, N3249, N2360);
nor NOR4 (N3255, N3216, N1338, N1289, N2959);
xor XOR2 (N3256, N3248, N2637);
buf BUF1 (N3257, N3250);
or OR2 (N3258, N3247, N2510);
nand NAND4 (N3259, N3254, N775, N262, N2428);
xor XOR2 (N3260, N3255, N2325);
not NOT1 (N3261, N3229);
or OR3 (N3262, N3259, N902, N487);
xor XOR2 (N3263, N3252, N74);
buf BUF1 (N3264, N3257);
nand NAND3 (N3265, N3214, N2525, N1107);
or OR3 (N3266, N3251, N2190, N1475);
nand NAND4 (N3267, N3265, N1872, N2488, N2103);
xor XOR2 (N3268, N3262, N2551);
not NOT1 (N3269, N3266);
xor XOR2 (N3270, N3256, N2302);
or OR4 (N3271, N3267, N2381, N174, N1591);
xor XOR2 (N3272, N3258, N71);
buf BUF1 (N3273, N3263);
and AND2 (N3274, N3268, N1499);
or OR4 (N3275, N3274, N1093, N3016, N813);
and AND4 (N3276, N3270, N2946, N1463, N150);
xor XOR2 (N3277, N3264, N2581);
nand NAND2 (N3278, N3272, N2113);
buf BUF1 (N3279, N3278);
or OR2 (N3280, N3269, N2259);
xor XOR2 (N3281, N3280, N2401);
nor NOR2 (N3282, N3253, N2543);
and AND4 (N3283, N3273, N2978, N710, N1131);
not NOT1 (N3284, N3271);
nor NOR3 (N3285, N3279, N939, N717);
nand NAND2 (N3286, N3276, N1648);
or OR2 (N3287, N3275, N2871);
and AND4 (N3288, N3260, N2584, N2504, N2079);
not NOT1 (N3289, N3286);
and AND2 (N3290, N3288, N782);
or OR2 (N3291, N3285, N856);
or OR3 (N3292, N3283, N475, N214);
nand NAND3 (N3293, N3292, N725, N972);
not NOT1 (N3294, N3290);
not NOT1 (N3295, N3294);
buf BUF1 (N3296, N3289);
buf BUF1 (N3297, N3296);
nand NAND3 (N3298, N3261, N2601, N2953);
or OR2 (N3299, N3287, N1927);
buf BUF1 (N3300, N3282);
and AND4 (N3301, N3281, N2097, N1879, N105);
buf BUF1 (N3302, N3299);
not NOT1 (N3303, N3291);
xor XOR2 (N3304, N3298, N672);
or OR2 (N3305, N3300, N2319);
or OR2 (N3306, N3293, N3282);
nor NOR4 (N3307, N3306, N1610, N2415, N1598);
buf BUF1 (N3308, N3297);
and AND2 (N3309, N3301, N540);
and AND2 (N3310, N3284, N3121);
nand NAND4 (N3311, N3307, N2327, N3225, N244);
not NOT1 (N3312, N3304);
not NOT1 (N3313, N3303);
nor NOR2 (N3314, N3302, N1411);
and AND4 (N3315, N3311, N1112, N382, N1503);
buf BUF1 (N3316, N3312);
buf BUF1 (N3317, N3309);
xor XOR2 (N3318, N3316, N518);
xor XOR2 (N3319, N3313, N60);
nor NOR4 (N3320, N3295, N2105, N1390, N1167);
xor XOR2 (N3321, N3305, N1507);
buf BUF1 (N3322, N3320);
or OR4 (N3323, N3310, N3090, N2294, N1767);
nand NAND4 (N3324, N3321, N2782, N706, N2534);
and AND3 (N3325, N3319, N385, N603);
nand NAND2 (N3326, N3314, N64);
not NOT1 (N3327, N3318);
or OR3 (N3328, N3326, N1933, N473);
xor XOR2 (N3329, N3322, N932);
not NOT1 (N3330, N3327);
xor XOR2 (N3331, N3328, N3183);
and AND3 (N3332, N3329, N1933, N2110);
nor NOR4 (N3333, N3331, N56, N2346, N3146);
buf BUF1 (N3334, N3315);
not NOT1 (N3335, N3334);
nand NAND3 (N3336, N3277, N672, N272);
or OR3 (N3337, N3323, N2752, N636);
xor XOR2 (N3338, N3332, N2088);
not NOT1 (N3339, N3325);
xor XOR2 (N3340, N3337, N391);
not NOT1 (N3341, N3336);
not NOT1 (N3342, N3338);
xor XOR2 (N3343, N3340, N3115);
and AND4 (N3344, N3317, N2277, N915, N3146);
and AND4 (N3345, N3330, N2137, N556, N1086);
and AND2 (N3346, N3333, N2182);
or OR3 (N3347, N3344, N2403, N511);
nand NAND2 (N3348, N3339, N2844);
nand NAND2 (N3349, N3348, N2727);
not NOT1 (N3350, N3347);
not NOT1 (N3351, N3343);
or OR4 (N3352, N3351, N1170, N2137, N2224);
and AND4 (N3353, N3341, N1681, N2996, N2848);
not NOT1 (N3354, N3353);
not NOT1 (N3355, N3352);
not NOT1 (N3356, N3345);
and AND3 (N3357, N3324, N487, N2398);
or OR3 (N3358, N3342, N2470, N2796);
xor XOR2 (N3359, N3358, N1643);
not NOT1 (N3360, N3355);
or OR4 (N3361, N3356, N816, N2383, N2315);
nand NAND3 (N3362, N3346, N1135, N416);
or OR2 (N3363, N3362, N827);
buf BUF1 (N3364, N3363);
nand NAND4 (N3365, N3364, N1146, N2922, N2231);
xor XOR2 (N3366, N3308, N1524);
not NOT1 (N3367, N3350);
or OR2 (N3368, N3365, N3054);
and AND4 (N3369, N3360, N2755, N1292, N603);
or OR3 (N3370, N3361, N2100, N1554);
buf BUF1 (N3371, N3357);
xor XOR2 (N3372, N3366, N1542);
buf BUF1 (N3373, N3335);
nor NOR4 (N3374, N3359, N3045, N1008, N863);
nand NAND4 (N3375, N3371, N2982, N2416, N2633);
not NOT1 (N3376, N3349);
xor XOR2 (N3377, N3370, N1601);
nand NAND2 (N3378, N3375, N77);
not NOT1 (N3379, N3376);
xor XOR2 (N3380, N3367, N3187);
xor XOR2 (N3381, N3372, N3047);
not NOT1 (N3382, N3374);
and AND3 (N3383, N3380, N309, N550);
and AND3 (N3384, N3373, N3077, N1003);
xor XOR2 (N3385, N3381, N877);
and AND3 (N3386, N3369, N2611, N55);
not NOT1 (N3387, N3377);
buf BUF1 (N3388, N3368);
not NOT1 (N3389, N3378);
and AND2 (N3390, N3383, N2050);
xor XOR2 (N3391, N3390, N1025);
and AND2 (N3392, N3391, N1699);
nand NAND2 (N3393, N3386, N1128);
nor NOR3 (N3394, N3379, N2602, N2703);
xor XOR2 (N3395, N3354, N2629);
not NOT1 (N3396, N3384);
and AND2 (N3397, N3388, N2260);
nand NAND4 (N3398, N3396, N2703, N680, N86);
and AND3 (N3399, N3382, N3111, N2255);
or OR3 (N3400, N3399, N1770, N1349);
not NOT1 (N3401, N3387);
not NOT1 (N3402, N3397);
and AND4 (N3403, N3395, N3042, N761, N879);
and AND3 (N3404, N3393, N1898, N466);
and AND2 (N3405, N3403, N1428);
nand NAND2 (N3406, N3398, N36);
and AND3 (N3407, N3392, N2798, N1691);
nor NOR4 (N3408, N3406, N173, N1043, N984);
not NOT1 (N3409, N3407);
buf BUF1 (N3410, N3389);
buf BUF1 (N3411, N3405);
buf BUF1 (N3412, N3385);
or OR3 (N3413, N3412, N1838, N2155);
nor NOR3 (N3414, N3401, N853, N18);
nor NOR2 (N3415, N3414, N2646);
not NOT1 (N3416, N3408);
or OR3 (N3417, N3400, N1577, N2824);
buf BUF1 (N3418, N3410);
or OR2 (N3419, N3415, N1834);
and AND3 (N3420, N3394, N2433, N3391);
nor NOR4 (N3421, N3413, N2107, N1142, N579);
xor XOR2 (N3422, N3402, N1185);
xor XOR2 (N3423, N3420, N3372);
nor NOR2 (N3424, N3418, N2304);
nand NAND2 (N3425, N3409, N520);
or OR3 (N3426, N3425, N3137, N2000);
or OR2 (N3427, N3411, N3150);
xor XOR2 (N3428, N3419, N1360);
nor NOR4 (N3429, N3404, N1827, N1662, N1643);
and AND4 (N3430, N3416, N3167, N1622, N1787);
not NOT1 (N3431, N3430);
nand NAND3 (N3432, N3427, N930, N2623);
xor XOR2 (N3433, N3429, N2178);
xor XOR2 (N3434, N3428, N3203);
nand NAND3 (N3435, N3433, N1722, N1273);
xor XOR2 (N3436, N3431, N720);
nand NAND3 (N3437, N3417, N305, N1136);
and AND4 (N3438, N3426, N1663, N2158, N169);
nor NOR4 (N3439, N3432, N556, N1482, N1441);
xor XOR2 (N3440, N3439, N880);
buf BUF1 (N3441, N3421);
and AND3 (N3442, N3422, N1032, N962);
not NOT1 (N3443, N3436);
nor NOR4 (N3444, N3443, N1844, N2962, N820);
and AND3 (N3445, N3435, N1229, N3211);
nand NAND4 (N3446, N3434, N1165, N1885, N1220);
not NOT1 (N3447, N3445);
xor XOR2 (N3448, N3423, N904);
or OR2 (N3449, N3448, N2671);
buf BUF1 (N3450, N3449);
xor XOR2 (N3451, N3441, N420);
and AND4 (N3452, N3442, N3433, N144, N1662);
xor XOR2 (N3453, N3437, N317);
or OR3 (N3454, N3450, N2581, N95);
nand NAND3 (N3455, N3438, N1305, N886);
not NOT1 (N3456, N3444);
nor NOR2 (N3457, N3452, N3396);
xor XOR2 (N3458, N3424, N2777);
and AND3 (N3459, N3451, N2576, N852);
nand NAND4 (N3460, N3447, N2946, N1209, N2251);
buf BUF1 (N3461, N3460);
xor XOR2 (N3462, N3457, N2353);
nand NAND3 (N3463, N3462, N3022, N2066);
not NOT1 (N3464, N3463);
and AND4 (N3465, N3455, N3232, N1080, N2415);
buf BUF1 (N3466, N3446);
and AND3 (N3467, N3465, N681, N2739);
not NOT1 (N3468, N3458);
not NOT1 (N3469, N3453);
nand NAND4 (N3470, N3456, N835, N582, N1005);
nand NAND4 (N3471, N3454, N2396, N2225, N1289);
nor NOR4 (N3472, N3459, N2885, N2642, N2458);
xor XOR2 (N3473, N3472, N1525);
nor NOR3 (N3474, N3468, N2899, N1922);
buf BUF1 (N3475, N3464);
not NOT1 (N3476, N3461);
not NOT1 (N3477, N3466);
xor XOR2 (N3478, N3467, N871);
not NOT1 (N3479, N3471);
nor NOR2 (N3480, N3473, N1716);
nor NOR3 (N3481, N3478, N733, N2375);
or OR4 (N3482, N3477, N3218, N2795, N1938);
xor XOR2 (N3483, N3481, N478);
buf BUF1 (N3484, N3482);
or OR4 (N3485, N3474, N418, N33, N2383);
and AND4 (N3486, N3479, N1546, N2636, N666);
or OR3 (N3487, N3486, N1564, N415);
nor NOR3 (N3488, N3469, N2952, N455);
nor NOR4 (N3489, N3485, N776, N2202, N2373);
buf BUF1 (N3490, N3476);
nand NAND3 (N3491, N3484, N3331, N347);
nand NAND2 (N3492, N3475, N377);
or OR3 (N3493, N3491, N2151, N2712);
buf BUF1 (N3494, N3487);
or OR2 (N3495, N3489, N950);
or OR2 (N3496, N3488, N184);
not NOT1 (N3497, N3492);
xor XOR2 (N3498, N3497, N3177);
and AND3 (N3499, N3493, N1688, N954);
nand NAND4 (N3500, N3494, N1009, N329, N3484);
nor NOR4 (N3501, N3490, N3112, N405, N126);
buf BUF1 (N3502, N3480);
buf BUF1 (N3503, N3483);
xor XOR2 (N3504, N3502, N1753);
or OR2 (N3505, N3498, N1503);
not NOT1 (N3506, N3440);
nor NOR3 (N3507, N3470, N2871, N1888);
xor XOR2 (N3508, N3499, N220);
nor NOR4 (N3509, N3505, N2342, N2938, N1600);
nor NOR2 (N3510, N3501, N2573);
nor NOR4 (N3511, N3504, N166, N122, N2200);
nor NOR3 (N3512, N3509, N2086, N3405);
xor XOR2 (N3513, N3508, N1001);
nor NOR4 (N3514, N3513, N2921, N283, N2695);
buf BUF1 (N3515, N3496);
nor NOR2 (N3516, N3514, N191);
nor NOR2 (N3517, N3511, N1312);
or OR2 (N3518, N3516, N2977);
or OR2 (N3519, N3506, N2936);
and AND4 (N3520, N3512, N357, N2839, N882);
nor NOR3 (N3521, N3503, N2344, N208);
nor NOR2 (N3522, N3500, N1910);
and AND3 (N3523, N3519, N929, N1084);
and AND2 (N3524, N3521, N3181);
or OR2 (N3525, N3515, N1233);
buf BUF1 (N3526, N3524);
xor XOR2 (N3527, N3525, N787);
nand NAND3 (N3528, N3526, N160, N2576);
and AND2 (N3529, N3523, N2180);
or OR3 (N3530, N3520, N1462, N3140);
nand NAND4 (N3531, N3522, N3126, N2397, N962);
and AND4 (N3532, N3527, N367, N1360, N2778);
or OR2 (N3533, N3532, N1720);
buf BUF1 (N3534, N3510);
nand NAND3 (N3535, N3529, N946, N3080);
xor XOR2 (N3536, N3518, N3228);
nand NAND3 (N3537, N3536, N1539, N546);
nand NAND4 (N3538, N3533, N1787, N2493, N2759);
nand NAND3 (N3539, N3530, N2726, N2096);
and AND3 (N3540, N3528, N3199, N168);
and AND3 (N3541, N3539, N222, N3408);
or OR4 (N3542, N3538, N2178, N2598, N412);
buf BUF1 (N3543, N3534);
or OR3 (N3544, N3517, N1265, N3399);
xor XOR2 (N3545, N3507, N2122);
not NOT1 (N3546, N3545);
or OR2 (N3547, N3542, N3179);
xor XOR2 (N3548, N3495, N939);
nor NOR3 (N3549, N3535, N1094, N1656);
buf BUF1 (N3550, N3546);
and AND2 (N3551, N3540, N745);
xor XOR2 (N3552, N3537, N1785);
xor XOR2 (N3553, N3531, N3457);
or OR4 (N3554, N3551, N526, N386, N2218);
nor NOR3 (N3555, N3548, N2564, N2018);
xor XOR2 (N3556, N3541, N1533);
nand NAND3 (N3557, N3543, N590, N2857);
nor NOR2 (N3558, N3549, N3444);
nand NAND4 (N3559, N3557, N1390, N2417, N625);
not NOT1 (N3560, N3550);
nor NOR4 (N3561, N3555, N1725, N934, N501);
nand NAND4 (N3562, N3554, N3426, N1831, N3053);
and AND2 (N3563, N3562, N2160);
nor NOR4 (N3564, N3561, N3342, N2435, N16);
not NOT1 (N3565, N3547);
and AND4 (N3566, N3565, N3559, N3450, N1423);
nor NOR4 (N3567, N653, N2158, N2003, N3291);
buf BUF1 (N3568, N3566);
xor XOR2 (N3569, N3567, N2876);
not NOT1 (N3570, N3544);
nand NAND4 (N3571, N3556, N2941, N1345, N101);
not NOT1 (N3572, N3570);
or OR2 (N3573, N3558, N592);
nand NAND3 (N3574, N3560, N3048, N2432);
xor XOR2 (N3575, N3574, N1524);
buf BUF1 (N3576, N3552);
buf BUF1 (N3577, N3568);
xor XOR2 (N3578, N3573, N1278);
not NOT1 (N3579, N3553);
nor NOR4 (N3580, N3576, N3361, N3132, N259);
xor XOR2 (N3581, N3569, N927);
nand NAND4 (N3582, N3577, N2137, N1598, N3256);
or OR4 (N3583, N3579, N2175, N1861, N3127);
xor XOR2 (N3584, N3580, N2025);
and AND2 (N3585, N3564, N1472);
nor NOR2 (N3586, N3578, N941);
nor NOR3 (N3587, N3584, N280, N1218);
xor XOR2 (N3588, N3563, N847);
not NOT1 (N3589, N3572);
or OR4 (N3590, N3589, N1693, N3062, N3446);
nand NAND2 (N3591, N3585, N3433);
not NOT1 (N3592, N3583);
and AND3 (N3593, N3588, N2451, N3219);
xor XOR2 (N3594, N3586, N1897);
or OR3 (N3595, N3575, N2939, N1012);
nor NOR3 (N3596, N3571, N2640, N833);
nand NAND2 (N3597, N3582, N2374);
and AND4 (N3598, N3597, N1019, N1329, N918);
nor NOR4 (N3599, N3596, N366, N2757, N1387);
or OR2 (N3600, N3590, N3101);
nor NOR2 (N3601, N3581, N1416);
buf BUF1 (N3602, N3591);
xor XOR2 (N3603, N3592, N2781);
and AND2 (N3604, N3601, N83);
and AND3 (N3605, N3593, N2112, N2621);
or OR2 (N3606, N3598, N2791);
nor NOR4 (N3607, N3587, N3226, N1390, N1599);
xor XOR2 (N3608, N3603, N1074);
not NOT1 (N3609, N3599);
not NOT1 (N3610, N3605);
or OR4 (N3611, N3594, N1109, N1015, N3553);
nor NOR4 (N3612, N3607, N1220, N3139, N1265);
nor NOR4 (N3613, N3606, N3582, N2318, N2772);
buf BUF1 (N3614, N3595);
buf BUF1 (N3615, N3600);
or OR3 (N3616, N3604, N685, N581);
or OR3 (N3617, N3613, N428, N2137);
nor NOR2 (N3618, N3610, N626);
nor NOR4 (N3619, N3609, N1524, N2649, N1213);
not NOT1 (N3620, N3618);
nand NAND4 (N3621, N3612, N279, N1414, N2750);
and AND2 (N3622, N3619, N2664);
buf BUF1 (N3623, N3611);
or OR2 (N3624, N3608, N1884);
not NOT1 (N3625, N3620);
or OR2 (N3626, N3615, N2427);
or OR3 (N3627, N3622, N2929, N56);
not NOT1 (N3628, N3623);
nor NOR3 (N3629, N3625, N2871, N2937);
not NOT1 (N3630, N3624);
and AND4 (N3631, N3617, N3329, N156, N2872);
not NOT1 (N3632, N3629);
and AND2 (N3633, N3627, N2664);
nor NOR3 (N3634, N3602, N2387, N2110);
nor NOR2 (N3635, N3631, N3218);
buf BUF1 (N3636, N3634);
or OR4 (N3637, N3614, N1261, N1709, N1264);
xor XOR2 (N3638, N3635, N2777);
and AND4 (N3639, N3636, N366, N1112, N2893);
nor NOR3 (N3640, N3639, N1347, N2032);
or OR4 (N3641, N3621, N2587, N604, N3268);
not NOT1 (N3642, N3630);
not NOT1 (N3643, N3638);
xor XOR2 (N3644, N3640, N2748);
not NOT1 (N3645, N3626);
nor NOR4 (N3646, N3645, N783, N934, N1697);
or OR3 (N3647, N3646, N788, N2297);
xor XOR2 (N3648, N3642, N1194);
nor NOR2 (N3649, N3616, N3581);
and AND3 (N3650, N3632, N427, N1180);
xor XOR2 (N3651, N3648, N1685);
buf BUF1 (N3652, N3641);
xor XOR2 (N3653, N3647, N101);
nand NAND4 (N3654, N3637, N3264, N1557, N1009);
buf BUF1 (N3655, N3650);
nor NOR3 (N3656, N3652, N270, N570);
and AND2 (N3657, N3628, N1911);
and AND3 (N3658, N3644, N481, N3187);
xor XOR2 (N3659, N3655, N2770);
and AND2 (N3660, N3651, N2941);
or OR4 (N3661, N3657, N1809, N2655, N2032);
nand NAND3 (N3662, N3658, N2936, N2408);
and AND4 (N3663, N3633, N2901, N2885, N1138);
not NOT1 (N3664, N3661);
or OR4 (N3665, N3660, N1586, N781, N2941);
or OR2 (N3666, N3654, N2695);
not NOT1 (N3667, N3643);
and AND2 (N3668, N3653, N2524);
nor NOR3 (N3669, N3656, N3629, N423);
not NOT1 (N3670, N3666);
nand NAND4 (N3671, N3649, N296, N3250, N1065);
or OR2 (N3672, N3671, N2269);
nand NAND2 (N3673, N3667, N1997);
buf BUF1 (N3674, N3664);
and AND4 (N3675, N3669, N769, N1620, N575);
buf BUF1 (N3676, N3663);
not NOT1 (N3677, N3665);
nand NAND4 (N3678, N3676, N571, N3409, N398);
buf BUF1 (N3679, N3673);
buf BUF1 (N3680, N3677);
xor XOR2 (N3681, N3659, N2017);
and AND3 (N3682, N3674, N1517, N731);
nand NAND4 (N3683, N3672, N941, N665, N2822);
buf BUF1 (N3684, N3678);
buf BUF1 (N3685, N3682);
buf BUF1 (N3686, N3679);
or OR4 (N3687, N3662, N2285, N406, N923);
not NOT1 (N3688, N3685);
xor XOR2 (N3689, N3680, N2766);
xor XOR2 (N3690, N3681, N3663);
and AND4 (N3691, N3689, N428, N1906, N1686);
xor XOR2 (N3692, N3684, N524);
or OR4 (N3693, N3675, N1530, N1075, N2532);
or OR4 (N3694, N3683, N1602, N1157, N3037);
xor XOR2 (N3695, N3694, N1374);
and AND3 (N3696, N3668, N2930, N2933);
xor XOR2 (N3697, N3690, N2124);
nor NOR3 (N3698, N3686, N2927, N1058);
nor NOR2 (N3699, N3698, N2501);
not NOT1 (N3700, N3688);
and AND2 (N3701, N3699, N2643);
and AND2 (N3702, N3701, N2555);
buf BUF1 (N3703, N3670);
and AND4 (N3704, N3687, N1957, N2164, N185);
xor XOR2 (N3705, N3697, N3380);
not NOT1 (N3706, N3703);
not NOT1 (N3707, N3705);
nand NAND4 (N3708, N3707, N2300, N2652, N3651);
not NOT1 (N3709, N3704);
or OR2 (N3710, N3692, N1618);
nand NAND4 (N3711, N3691, N2175, N2036, N1200);
xor XOR2 (N3712, N3710, N2659);
xor XOR2 (N3713, N3708, N2122);
and AND3 (N3714, N3700, N1730, N1521);
or OR2 (N3715, N3702, N100);
xor XOR2 (N3716, N3713, N2469);
nor NOR3 (N3717, N3712, N2765, N3527);
buf BUF1 (N3718, N3715);
and AND3 (N3719, N3706, N26, N1167);
and AND3 (N3720, N3716, N1999, N3132);
xor XOR2 (N3721, N3719, N822);
nor NOR4 (N3722, N3714, N3233, N1091, N72);
nand NAND3 (N3723, N3718, N3053, N425);
nor NOR3 (N3724, N3720, N1406, N324);
not NOT1 (N3725, N3709);
nor NOR2 (N3726, N3711, N964);
nand NAND2 (N3727, N3693, N3229);
buf BUF1 (N3728, N3727);
nand NAND4 (N3729, N3695, N3418, N391, N915);
and AND3 (N3730, N3723, N266, N3176);
buf BUF1 (N3731, N3728);
nor NOR4 (N3732, N3724, N3344, N1445, N1266);
or OR3 (N3733, N3732, N781, N2804);
xor XOR2 (N3734, N3721, N1865);
xor XOR2 (N3735, N3725, N3452);
nand NAND4 (N3736, N3717, N2249, N2180, N2730);
nand NAND2 (N3737, N3730, N2591);
nand NAND2 (N3738, N3726, N1401);
and AND3 (N3739, N3736, N42, N3227);
or OR2 (N3740, N3739, N1291);
and AND3 (N3741, N3733, N3426, N1196);
buf BUF1 (N3742, N3734);
not NOT1 (N3743, N3729);
xor XOR2 (N3744, N3696, N948);
not NOT1 (N3745, N3738);
or OR3 (N3746, N3742, N1908, N3368);
nor NOR3 (N3747, N3746, N3103, N2565);
xor XOR2 (N3748, N3737, N2977);
nor NOR4 (N3749, N3735, N1327, N542, N2973);
buf BUF1 (N3750, N3745);
not NOT1 (N3751, N3744);
or OR4 (N3752, N3743, N3487, N1057, N176);
and AND3 (N3753, N3740, N393, N718);
nor NOR2 (N3754, N3750, N1220);
xor XOR2 (N3755, N3749, N2246);
nand NAND3 (N3756, N3747, N2877, N3168);
nand NAND3 (N3757, N3754, N952, N2380);
nor NOR3 (N3758, N3757, N1847, N849);
or OR2 (N3759, N3752, N92);
or OR4 (N3760, N3748, N3243, N354, N250);
or OR2 (N3761, N3753, N3611);
and AND3 (N3762, N3759, N647, N3189);
not NOT1 (N3763, N3761);
not NOT1 (N3764, N3741);
nand NAND3 (N3765, N3751, N3452, N2952);
nor NOR2 (N3766, N3731, N2115);
nor NOR4 (N3767, N3764, N17, N1552, N945);
buf BUF1 (N3768, N3756);
not NOT1 (N3769, N3767);
nand NAND3 (N3770, N3722, N3304, N3065);
or OR4 (N3771, N3770, N2909, N3748, N3303);
buf BUF1 (N3772, N3771);
buf BUF1 (N3773, N3768);
nand NAND3 (N3774, N3758, N1209, N1629);
or OR4 (N3775, N3762, N92, N3663, N2819);
nand NAND2 (N3776, N3766, N429);
nor NOR3 (N3777, N3763, N1239, N3554);
xor XOR2 (N3778, N3765, N1205);
not NOT1 (N3779, N3777);
nand NAND3 (N3780, N3772, N3354, N2028);
and AND3 (N3781, N3774, N1630, N2354);
and AND4 (N3782, N3779, N1558, N2461, N851);
buf BUF1 (N3783, N3755);
and AND3 (N3784, N3775, N3034, N391);
not NOT1 (N3785, N3780);
nand NAND4 (N3786, N3776, N161, N1901, N3411);
nor NOR4 (N3787, N3785, N3454, N3747, N5);
nor NOR4 (N3788, N3782, N3462, N2942, N1066);
buf BUF1 (N3789, N3783);
nand NAND2 (N3790, N3786, N3068);
buf BUF1 (N3791, N3784);
or OR3 (N3792, N3781, N3273, N3011);
not NOT1 (N3793, N3760);
nand NAND2 (N3794, N3773, N2916);
nand NAND2 (N3795, N3778, N3781);
nand NAND2 (N3796, N3788, N3107);
nor NOR2 (N3797, N3791, N6);
nand NAND3 (N3798, N3793, N2006, N735);
nor NOR2 (N3799, N3797, N3150);
and AND4 (N3800, N3795, N2158, N2062, N3614);
nor NOR2 (N3801, N3792, N1712);
nor NOR4 (N3802, N3790, N977, N938, N3353);
nand NAND2 (N3803, N3789, N849);
or OR3 (N3804, N3802, N1547, N3289);
buf BUF1 (N3805, N3799);
buf BUF1 (N3806, N3800);
nand NAND2 (N3807, N3805, N983);
nor NOR2 (N3808, N3801, N494);
nor NOR4 (N3809, N3794, N2571, N206, N339);
not NOT1 (N3810, N3806);
nor NOR4 (N3811, N3804, N1890, N1742, N2952);
nand NAND4 (N3812, N3787, N2442, N3166, N2891);
buf BUF1 (N3813, N3811);
nand NAND4 (N3814, N3798, N874, N262, N2177);
or OR2 (N3815, N3769, N2626);
buf BUF1 (N3816, N3814);
or OR2 (N3817, N3816, N2755);
or OR4 (N3818, N3803, N986, N21, N1033);
buf BUF1 (N3819, N3807);
buf BUF1 (N3820, N3796);
nor NOR4 (N3821, N3818, N2184, N1786, N1349);
nand NAND4 (N3822, N3819, N1704, N99, N1231);
nor NOR2 (N3823, N3809, N3066);
not NOT1 (N3824, N3815);
buf BUF1 (N3825, N3808);
nor NOR3 (N3826, N3821, N3479, N2066);
not NOT1 (N3827, N3813);
buf BUF1 (N3828, N3822);
buf BUF1 (N3829, N3812);
nand NAND2 (N3830, N3825, N3810);
xor XOR2 (N3831, N1857, N3249);
xor XOR2 (N3832, N3827, N410);
buf BUF1 (N3833, N3832);
or OR3 (N3834, N3828, N1002, N875);
and AND3 (N3835, N3826, N706, N2974);
nand NAND4 (N3836, N3829, N73, N2239, N2625);
nor NOR2 (N3837, N3835, N2578);
not NOT1 (N3838, N3817);
or OR4 (N3839, N3823, N409, N2164, N3106);
xor XOR2 (N3840, N3831, N1603);
not NOT1 (N3841, N3830);
not NOT1 (N3842, N3837);
buf BUF1 (N3843, N3839);
nand NAND2 (N3844, N3842, N1139);
buf BUF1 (N3845, N3838);
nand NAND3 (N3846, N3834, N852, N2656);
and AND3 (N3847, N3845, N3242, N2346);
nor NOR2 (N3848, N3844, N2817);
nand NAND2 (N3849, N3833, N579);
xor XOR2 (N3850, N3849, N951);
not NOT1 (N3851, N3824);
nor NOR2 (N3852, N3851, N1437);
nor NOR3 (N3853, N3836, N2628, N2154);
and AND2 (N3854, N3847, N315);
nand NAND2 (N3855, N3841, N3029);
buf BUF1 (N3856, N3848);
nor NOR4 (N3857, N3840, N3490, N3128, N2980);
xor XOR2 (N3858, N3850, N2326);
and AND4 (N3859, N3852, N2909, N184, N3545);
and AND3 (N3860, N3853, N1245, N960);
xor XOR2 (N3861, N3857, N1762);
not NOT1 (N3862, N3854);
not NOT1 (N3863, N3856);
not NOT1 (N3864, N3863);
not NOT1 (N3865, N3843);
nand NAND4 (N3866, N3858, N903, N2630, N1519);
nand NAND2 (N3867, N3864, N721);
nor NOR2 (N3868, N3866, N875);
or OR4 (N3869, N3861, N328, N1391, N390);
nor NOR3 (N3870, N3855, N3700, N2108);
and AND2 (N3871, N3859, N3610);
not NOT1 (N3872, N3820);
nor NOR3 (N3873, N3871, N370, N403);
buf BUF1 (N3874, N3873);
nor NOR2 (N3875, N3868, N3795);
xor XOR2 (N3876, N3874, N2710);
not NOT1 (N3877, N3846);
not NOT1 (N3878, N3867);
and AND2 (N3879, N3877, N1692);
buf BUF1 (N3880, N3860);
nand NAND3 (N3881, N3878, N2004, N291);
buf BUF1 (N3882, N3872);
nand NAND2 (N3883, N3865, N1653);
buf BUF1 (N3884, N3883);
not NOT1 (N3885, N3884);
not NOT1 (N3886, N3875);
nand NAND4 (N3887, N3882, N2284, N3347, N980);
buf BUF1 (N3888, N3886);
xor XOR2 (N3889, N3870, N3601);
not NOT1 (N3890, N3881);
buf BUF1 (N3891, N3880);
and AND3 (N3892, N3862, N2038, N2280);
xor XOR2 (N3893, N3891, N1551);
nand NAND4 (N3894, N3887, N1452, N306, N656);
buf BUF1 (N3895, N3876);
buf BUF1 (N3896, N3888);
nand NAND2 (N3897, N3896, N3542);
nor NOR2 (N3898, N3879, N3430);
not NOT1 (N3899, N3897);
xor XOR2 (N3900, N3890, N1235);
nor NOR4 (N3901, N3885, N3720, N1767, N1080);
buf BUF1 (N3902, N3894);
and AND4 (N3903, N3902, N809, N2044, N1567);
buf BUF1 (N3904, N3892);
and AND3 (N3905, N3904, N617, N186);
not NOT1 (N3906, N3869);
and AND2 (N3907, N3895, N2990);
or OR3 (N3908, N3900, N1783, N2257);
not NOT1 (N3909, N3908);
nor NOR2 (N3910, N3909, N668);
buf BUF1 (N3911, N3889);
nor NOR3 (N3912, N3911, N1935, N1141);
buf BUF1 (N3913, N3910);
nor NOR3 (N3914, N3899, N2684, N529);
buf BUF1 (N3915, N3903);
not NOT1 (N3916, N3907);
and AND4 (N3917, N3905, N493, N2164, N1435);
nand NAND4 (N3918, N3912, N2018, N1278, N788);
xor XOR2 (N3919, N3913, N3788);
buf BUF1 (N3920, N3918);
or OR3 (N3921, N3915, N960, N1607);
buf BUF1 (N3922, N3917);
buf BUF1 (N3923, N3906);
and AND4 (N3924, N3916, N1418, N3870, N2387);
and AND4 (N3925, N3898, N1582, N307, N180);
buf BUF1 (N3926, N3922);
buf BUF1 (N3927, N3893);
nand NAND4 (N3928, N3901, N3499, N152, N3445);
buf BUF1 (N3929, N3928);
or OR3 (N3930, N3926, N2407, N2809);
or OR2 (N3931, N3929, N3482);
nor NOR4 (N3932, N3923, N1022, N1572, N2707);
xor XOR2 (N3933, N3921, N2602);
nor NOR2 (N3934, N3925, N2896);
buf BUF1 (N3935, N3920);
buf BUF1 (N3936, N3934);
or OR2 (N3937, N3931, N2397);
buf BUF1 (N3938, N3927);
xor XOR2 (N3939, N3914, N1768);
not NOT1 (N3940, N3939);
xor XOR2 (N3941, N3932, N1114);
and AND4 (N3942, N3937, N2822, N3441, N238);
nor NOR3 (N3943, N3924, N2041, N1550);
nor NOR4 (N3944, N3935, N1321, N2236, N378);
nand NAND4 (N3945, N3942, N425, N3520, N3507);
and AND3 (N3946, N3936, N1640, N739);
not NOT1 (N3947, N3941);
xor XOR2 (N3948, N3940, N780);
buf BUF1 (N3949, N3933);
buf BUF1 (N3950, N3943);
not NOT1 (N3951, N3944);
or OR2 (N3952, N3950, N2220);
nand NAND2 (N3953, N3948, N1423);
xor XOR2 (N3954, N3953, N1823);
buf BUF1 (N3955, N3930);
nand NAND3 (N3956, N3945, N1945, N2716);
buf BUF1 (N3957, N3949);
xor XOR2 (N3958, N3938, N1971);
and AND3 (N3959, N3919, N960, N1205);
xor XOR2 (N3960, N3946, N819);
and AND2 (N3961, N3954, N95);
or OR4 (N3962, N3960, N155, N317, N3838);
nor NOR4 (N3963, N3957, N964, N3034, N758);
buf BUF1 (N3964, N3952);
not NOT1 (N3965, N3958);
nor NOR2 (N3966, N3965, N1782);
not NOT1 (N3967, N3961);
and AND2 (N3968, N3951, N736);
not NOT1 (N3969, N3968);
xor XOR2 (N3970, N3963, N2699);
nand NAND2 (N3971, N3956, N3923);
or OR4 (N3972, N3971, N1849, N2539, N705);
or OR4 (N3973, N3964, N1971, N257, N1272);
buf BUF1 (N3974, N3966);
or OR3 (N3975, N3970, N1733, N1691);
nor NOR2 (N3976, N3955, N151);
nand NAND3 (N3977, N3967, N78, N134);
not NOT1 (N3978, N3976);
and AND4 (N3979, N3978, N1768, N681, N3484);
nand NAND2 (N3980, N3979, N3650);
and AND2 (N3981, N3973, N2721);
not NOT1 (N3982, N3959);
nand NAND3 (N3983, N3969, N2157, N3965);
nor NOR4 (N3984, N3983, N1258, N2095, N884);
xor XOR2 (N3985, N3947, N2601);
xor XOR2 (N3986, N3980, N1183);
not NOT1 (N3987, N3962);
not NOT1 (N3988, N3972);
not NOT1 (N3989, N3984);
buf BUF1 (N3990, N3989);
and AND2 (N3991, N3975, N247);
buf BUF1 (N3992, N3977);
buf BUF1 (N3993, N3982);
or OR2 (N3994, N3987, N2371);
or OR3 (N3995, N3988, N2772, N1457);
nand NAND4 (N3996, N3990, N2798, N2210, N3920);
or OR3 (N3997, N3974, N1866, N3499);
not NOT1 (N3998, N3994);
buf BUF1 (N3999, N3991);
not NOT1 (N4000, N3993);
not NOT1 (N4001, N3985);
or OR3 (N4002, N3995, N2457, N1571);
nand NAND2 (N4003, N3996, N508);
nand NAND4 (N4004, N3999, N2545, N2291, N2237);
and AND3 (N4005, N4002, N1979, N2697);
or OR2 (N4006, N3992, N1249);
buf BUF1 (N4007, N4005);
and AND2 (N4008, N4007, N3705);
and AND2 (N4009, N3981, N984);
or OR2 (N4010, N3997, N679);
xor XOR2 (N4011, N4006, N3861);
and AND2 (N4012, N4010, N3806);
xor XOR2 (N4013, N4008, N355);
and AND3 (N4014, N3986, N2608, N3081);
nand NAND3 (N4015, N4003, N2519, N3929);
or OR4 (N4016, N4011, N955, N3976, N3331);
and AND2 (N4017, N4009, N3478);
not NOT1 (N4018, N4012);
nand NAND2 (N4019, N4013, N1594);
or OR2 (N4020, N4004, N2867);
buf BUF1 (N4021, N4015);
not NOT1 (N4022, N4020);
and AND2 (N4023, N4001, N3909);
or OR3 (N4024, N4019, N64, N3717);
nand NAND4 (N4025, N4000, N2728, N880, N2456);
not NOT1 (N4026, N4018);
and AND3 (N4027, N4014, N329, N3813);
or OR2 (N4028, N4024, N2113);
or OR4 (N4029, N4028, N1444, N749, N3427);
nor NOR2 (N4030, N4027, N2393);
nand NAND4 (N4031, N4029, N1041, N50, N3333);
or OR3 (N4032, N4031, N229, N401);
nand NAND3 (N4033, N4017, N1939, N1098);
or OR2 (N4034, N3998, N1698);
xor XOR2 (N4035, N4033, N2812);
nand NAND2 (N4036, N4016, N3438);
not NOT1 (N4037, N4036);
xor XOR2 (N4038, N4026, N3220);
xor XOR2 (N4039, N4032, N2648);
not NOT1 (N4040, N4030);
not NOT1 (N4041, N4034);
or OR2 (N4042, N4037, N686);
and AND4 (N4043, N4022, N2536, N2781, N2929);
nand NAND4 (N4044, N4038, N3124, N3706, N1257);
or OR4 (N4045, N4023, N651, N2205, N1226);
and AND4 (N4046, N4040, N611, N3352, N2974);
xor XOR2 (N4047, N4044, N2181);
nor NOR4 (N4048, N4043, N603, N502, N1535);
buf BUF1 (N4049, N4025);
nor NOR2 (N4050, N4047, N1915);
and AND2 (N4051, N4021, N976);
not NOT1 (N4052, N4048);
nor NOR3 (N4053, N4052, N2442, N446);
not NOT1 (N4054, N4035);
nand NAND2 (N4055, N4045, N1492);
nand NAND3 (N4056, N4055, N950, N126);
nand NAND3 (N4057, N4054, N3919, N1520);
or OR2 (N4058, N4041, N797);
and AND4 (N4059, N4050, N1483, N2682, N1802);
nor NOR2 (N4060, N4049, N720);
and AND2 (N4061, N4057, N1154);
nor NOR2 (N4062, N4039, N3031);
xor XOR2 (N4063, N4056, N3605);
buf BUF1 (N4064, N4062);
and AND4 (N4065, N4046, N3974, N2741, N3881);
or OR4 (N4066, N4053, N3200, N1678, N3755);
nand NAND2 (N4067, N4060, N1357);
nand NAND2 (N4068, N4064, N1408);
not NOT1 (N4069, N4042);
not NOT1 (N4070, N4051);
and AND2 (N4071, N4070, N1165);
not NOT1 (N4072, N4067);
buf BUF1 (N4073, N4058);
and AND2 (N4074, N4059, N2201);
buf BUF1 (N4075, N4074);
nand NAND4 (N4076, N4068, N1901, N1730, N2315);
nand NAND3 (N4077, N4065, N2648, N112);
nand NAND2 (N4078, N4073, N1228);
buf BUF1 (N4079, N4063);
and AND3 (N4080, N4077, N2606, N1471);
nor NOR2 (N4081, N4071, N1875);
xor XOR2 (N4082, N4079, N2220);
and AND3 (N4083, N4078, N150, N1609);
or OR4 (N4084, N4066, N2766, N3141, N2754);
buf BUF1 (N4085, N4080);
buf BUF1 (N4086, N4085);
or OR4 (N4087, N4069, N204, N3792, N3567);
xor XOR2 (N4088, N4061, N2314);
not NOT1 (N4089, N4084);
or OR3 (N4090, N4087, N3235, N2008);
or OR4 (N4091, N4089, N2405, N71, N2450);
nor NOR3 (N4092, N4086, N2424, N769);
nor NOR2 (N4093, N4083, N4057);
buf BUF1 (N4094, N4092);
xor XOR2 (N4095, N4090, N3110);
buf BUF1 (N4096, N4082);
nor NOR2 (N4097, N4081, N3379);
buf BUF1 (N4098, N4076);
buf BUF1 (N4099, N4088);
xor XOR2 (N4100, N4096, N2581);
buf BUF1 (N4101, N4095);
buf BUF1 (N4102, N4094);
xor XOR2 (N4103, N4075, N2925);
not NOT1 (N4104, N4072);
xor XOR2 (N4105, N4100, N3797);
nor NOR4 (N4106, N4104, N1691, N1648, N107);
or OR3 (N4107, N4105, N2861, N1666);
and AND2 (N4108, N4101, N1732);
nor NOR4 (N4109, N4106, N2028, N2189, N178);
buf BUF1 (N4110, N4091);
xor XOR2 (N4111, N4093, N573);
xor XOR2 (N4112, N4107, N867);
nand NAND4 (N4113, N4109, N3736, N1225, N144);
and AND3 (N4114, N4099, N706, N3653);
not NOT1 (N4115, N4103);
buf BUF1 (N4116, N4111);
not NOT1 (N4117, N4102);
buf BUF1 (N4118, N4098);
not NOT1 (N4119, N4115);
not NOT1 (N4120, N4108);
buf BUF1 (N4121, N4120);
buf BUF1 (N4122, N4118);
or OR2 (N4123, N4121, N2868);
or OR3 (N4124, N4117, N1666, N2257);
or OR4 (N4125, N4122, N2029, N3592, N1477);
xor XOR2 (N4126, N4123, N3521);
buf BUF1 (N4127, N4110);
and AND4 (N4128, N4126, N706, N2714, N1414);
nand NAND2 (N4129, N4127, N3532);
not NOT1 (N4130, N4097);
nor NOR2 (N4131, N4116, N3022);
not NOT1 (N4132, N4114);
xor XOR2 (N4133, N4124, N3721);
nand NAND2 (N4134, N4130, N3882);
nand NAND3 (N4135, N4131, N252, N3062);
nor NOR2 (N4136, N4119, N293);
nor NOR3 (N4137, N4136, N3722, N3198);
buf BUF1 (N4138, N4137);
not NOT1 (N4139, N4125);
nand NAND3 (N4140, N4128, N727, N3495);
and AND3 (N4141, N4113, N3950, N3737);
nand NAND2 (N4142, N4141, N2956);
or OR4 (N4143, N4142, N2902, N786, N2091);
or OR2 (N4144, N4133, N945);
or OR2 (N4145, N4144, N3680);
nor NOR4 (N4146, N4138, N1413, N3981, N863);
or OR4 (N4147, N4145, N3837, N2338, N2811);
not NOT1 (N4148, N4140);
nand NAND3 (N4149, N4147, N3014, N4133);
xor XOR2 (N4150, N4112, N1990);
buf BUF1 (N4151, N4132);
not NOT1 (N4152, N4149);
or OR2 (N4153, N4148, N1938);
nand NAND4 (N4154, N4146, N1234, N1163, N1015);
xor XOR2 (N4155, N4139, N1106);
xor XOR2 (N4156, N4154, N2254);
xor XOR2 (N4157, N4135, N577);
nand NAND3 (N4158, N4156, N234, N2804);
not NOT1 (N4159, N4152);
and AND2 (N4160, N4129, N1954);
xor XOR2 (N4161, N4150, N2034);
or OR2 (N4162, N4134, N3666);
or OR4 (N4163, N4153, N3506, N2018, N2247);
buf BUF1 (N4164, N4162);
not NOT1 (N4165, N4164);
xor XOR2 (N4166, N4161, N2096);
and AND4 (N4167, N4166, N3171, N3254, N3858);
xor XOR2 (N4168, N4157, N1233);
and AND2 (N4169, N4155, N908);
buf BUF1 (N4170, N4160);
xor XOR2 (N4171, N4165, N2667);
not NOT1 (N4172, N4159);
buf BUF1 (N4173, N4151);
nand NAND3 (N4174, N4171, N3826, N1191);
not NOT1 (N4175, N4158);
nand NAND3 (N4176, N4163, N343, N3693);
buf BUF1 (N4177, N4172);
and AND4 (N4178, N4167, N1160, N2439, N3724);
nor NOR2 (N4179, N4174, N1387);
not NOT1 (N4180, N4173);
not NOT1 (N4181, N4179);
or OR4 (N4182, N4170, N3719, N3597, N2842);
xor XOR2 (N4183, N4175, N1569);
not NOT1 (N4184, N4143);
xor XOR2 (N4185, N4178, N1995);
nor NOR4 (N4186, N4168, N2303, N345, N3345);
not NOT1 (N4187, N4184);
nand NAND3 (N4188, N4181, N2637, N119);
nand NAND4 (N4189, N4185, N2879, N525, N3300);
or OR4 (N4190, N4169, N652, N3281, N1211);
xor XOR2 (N4191, N4189, N1242);
xor XOR2 (N4192, N4183, N2242);
xor XOR2 (N4193, N4186, N108);
nor NOR4 (N4194, N4182, N526, N4129, N1360);
buf BUF1 (N4195, N4180);
buf BUF1 (N4196, N4177);
and AND4 (N4197, N4187, N48, N649, N2127);
nand NAND3 (N4198, N4194, N3295, N1660);
xor XOR2 (N4199, N4192, N3678);
not NOT1 (N4200, N4197);
nand NAND2 (N4201, N4200, N232);
not NOT1 (N4202, N4199);
xor XOR2 (N4203, N4196, N382);
nand NAND3 (N4204, N4202, N1554, N3291);
nor NOR3 (N4205, N4195, N1520, N334);
xor XOR2 (N4206, N4191, N3933);
xor XOR2 (N4207, N4203, N15);
and AND3 (N4208, N4205, N74, N2795);
nand NAND2 (N4209, N4176, N1207);
xor XOR2 (N4210, N4208, N4120);
or OR3 (N4211, N4207, N3087, N1795);
and AND4 (N4212, N4201, N570, N2051, N2734);
not NOT1 (N4213, N4206);
nor NOR2 (N4214, N4188, N3869);
nor NOR4 (N4215, N4210, N1554, N4065, N1175);
nand NAND2 (N4216, N4211, N2567);
buf BUF1 (N4217, N4213);
buf BUF1 (N4218, N4209);
not NOT1 (N4219, N4204);
and AND4 (N4220, N4218, N179, N373, N4213);
not NOT1 (N4221, N4220);
nand NAND3 (N4222, N4217, N2155, N2072);
xor XOR2 (N4223, N4198, N1115);
nand NAND3 (N4224, N4223, N2266, N2781);
and AND4 (N4225, N4219, N928, N3870, N4121);
and AND2 (N4226, N4212, N615);
xor XOR2 (N4227, N4224, N2096);
nor NOR4 (N4228, N4221, N392, N3217, N387);
buf BUF1 (N4229, N4215);
nor NOR4 (N4230, N4190, N717, N2718, N312);
not NOT1 (N4231, N4216);
not NOT1 (N4232, N4229);
buf BUF1 (N4233, N4222);
nand NAND2 (N4234, N4228, N1928);
or OR2 (N4235, N4230, N1993);
nor NOR3 (N4236, N4227, N36, N2630);
nor NOR3 (N4237, N4235, N48, N3659);
xor XOR2 (N4238, N4232, N2287);
not NOT1 (N4239, N4214);
buf BUF1 (N4240, N4238);
buf BUF1 (N4241, N4236);
or OR2 (N4242, N4234, N4043);
nor NOR2 (N4243, N4239, N3611);
xor XOR2 (N4244, N4241, N2622);
xor XOR2 (N4245, N4231, N3011);
not NOT1 (N4246, N4225);
nor NOR3 (N4247, N4245, N2289, N2671);
or OR2 (N4248, N4240, N171);
and AND3 (N4249, N4237, N3260, N1991);
or OR3 (N4250, N4243, N2561, N2094);
and AND4 (N4251, N4246, N3168, N1264, N1820);
nor NOR4 (N4252, N4251, N414, N683, N885);
or OR3 (N4253, N4233, N2887, N3150);
buf BUF1 (N4254, N4248);
buf BUF1 (N4255, N4250);
or OR2 (N4256, N4254, N2701);
buf BUF1 (N4257, N4253);
and AND3 (N4258, N4193, N3494, N833);
nand NAND2 (N4259, N4256, N2701);
not NOT1 (N4260, N4257);
buf BUF1 (N4261, N4249);
nand NAND3 (N4262, N4226, N314, N422);
nor NOR3 (N4263, N4259, N1578, N4123);
nor NOR2 (N4264, N4260, N1684);
or OR4 (N4265, N4252, N1163, N1849, N951);
nor NOR3 (N4266, N4255, N258, N4068);
nand NAND2 (N4267, N4242, N970);
nor NOR3 (N4268, N4266, N1990, N3520);
or OR4 (N4269, N4258, N3407, N164, N3605);
and AND2 (N4270, N4268, N3620);
nor NOR2 (N4271, N4269, N1180);
not NOT1 (N4272, N4247);
and AND2 (N4273, N4261, N2659);
nor NOR2 (N4274, N4265, N3795);
xor XOR2 (N4275, N4244, N241);
and AND3 (N4276, N4273, N2109, N2425);
nor NOR3 (N4277, N4272, N3981, N2473);
not NOT1 (N4278, N4263);
nand NAND2 (N4279, N4276, N2191);
buf BUF1 (N4280, N4262);
xor XOR2 (N4281, N4274, N3583);
xor XOR2 (N4282, N4279, N909);
buf BUF1 (N4283, N4271);
not NOT1 (N4284, N4278);
and AND2 (N4285, N4280, N2728);
and AND4 (N4286, N4282, N1468, N120, N804);
nand NAND2 (N4287, N4277, N1959);
or OR3 (N4288, N4285, N2339, N1934);
buf BUF1 (N4289, N4286);
nand NAND4 (N4290, N4288, N3923, N1667, N3836);
or OR4 (N4291, N4287, N178, N3791, N2532);
not NOT1 (N4292, N4275);
or OR4 (N4293, N4289, N3349, N439, N3915);
nor NOR2 (N4294, N4270, N1011);
xor XOR2 (N4295, N4290, N2276);
not NOT1 (N4296, N4284);
nor NOR3 (N4297, N4264, N2487, N983);
buf BUF1 (N4298, N4292);
and AND4 (N4299, N4296, N2311, N13, N1363);
xor XOR2 (N4300, N4295, N884);
buf BUF1 (N4301, N4293);
and AND3 (N4302, N4299, N102, N2746);
buf BUF1 (N4303, N4294);
and AND4 (N4304, N4281, N869, N1862, N2431);
or OR2 (N4305, N4303, N1158);
and AND3 (N4306, N4297, N194, N1087);
xor XOR2 (N4307, N4283, N3690);
xor XOR2 (N4308, N4267, N1358);
nand NAND2 (N4309, N4305, N593);
nor NOR4 (N4310, N4308, N1351, N3578, N1113);
buf BUF1 (N4311, N4307);
nand NAND3 (N4312, N4304, N758, N941);
buf BUF1 (N4313, N4302);
and AND2 (N4314, N4298, N3374);
nor NOR4 (N4315, N4291, N4126, N103, N1407);
nand NAND3 (N4316, N4309, N1749, N2225);
xor XOR2 (N4317, N4311, N3191);
xor XOR2 (N4318, N4300, N2889);
buf BUF1 (N4319, N4318);
not NOT1 (N4320, N4310);
and AND4 (N4321, N4317, N2973, N2285, N577);
xor XOR2 (N4322, N4315, N3264);
not NOT1 (N4323, N4301);
nand NAND3 (N4324, N4312, N2778, N2334);
nor NOR3 (N4325, N4320, N483, N4136);
or OR2 (N4326, N4323, N3392);
or OR3 (N4327, N4316, N1231, N376);
nand NAND4 (N4328, N4313, N3889, N1428, N3155);
buf BUF1 (N4329, N4314);
and AND3 (N4330, N4321, N502, N2897);
xor XOR2 (N4331, N4322, N2235);
buf BUF1 (N4332, N4324);
buf BUF1 (N4333, N4327);
not NOT1 (N4334, N4326);
buf BUF1 (N4335, N4306);
and AND4 (N4336, N4330, N4166, N3585, N1758);
buf BUF1 (N4337, N4336);
nand NAND2 (N4338, N4325, N3095);
or OR3 (N4339, N4338, N4000, N991);
xor XOR2 (N4340, N4335, N623);
buf BUF1 (N4341, N4334);
nor NOR4 (N4342, N4319, N1604, N133, N757);
not NOT1 (N4343, N4339);
buf BUF1 (N4344, N4332);
not NOT1 (N4345, N4328);
xor XOR2 (N4346, N4333, N4050);
buf BUF1 (N4347, N4331);
and AND2 (N4348, N4341, N1553);
xor XOR2 (N4349, N4345, N3216);
or OR4 (N4350, N4348, N3504, N1389, N3244);
or OR3 (N4351, N4342, N1355, N2456);
xor XOR2 (N4352, N4344, N3874);
not NOT1 (N4353, N4337);
not NOT1 (N4354, N4346);
or OR2 (N4355, N4343, N526);
xor XOR2 (N4356, N4340, N1763);
not NOT1 (N4357, N4353);
buf BUF1 (N4358, N4352);
nand NAND4 (N4359, N4356, N3088, N1393, N3673);
nor NOR2 (N4360, N4329, N2708);
nand NAND3 (N4361, N4351, N3575, N4124);
nor NOR4 (N4362, N4354, N4309, N807, N3110);
buf BUF1 (N4363, N4360);
xor XOR2 (N4364, N4358, N4242);
not NOT1 (N4365, N4350);
buf BUF1 (N4366, N4355);
and AND3 (N4367, N4363, N1552, N3952);
nor NOR4 (N4368, N4349, N3153, N3430, N943);
xor XOR2 (N4369, N4368, N3996);
nor NOR3 (N4370, N4365, N2923, N1728);
or OR2 (N4371, N4359, N2874);
buf BUF1 (N4372, N4347);
nor NOR4 (N4373, N4372, N1410, N3873, N555);
or OR4 (N4374, N4367, N2147, N868, N2300);
nor NOR3 (N4375, N4357, N297, N3535);
nand NAND3 (N4376, N4373, N1150, N3264);
nand NAND3 (N4377, N4364, N1771, N1901);
nand NAND2 (N4378, N4361, N3953);
not NOT1 (N4379, N4376);
nor NOR2 (N4380, N4379, N2787);
nor NOR2 (N4381, N4378, N3369);
not NOT1 (N4382, N4371);
not NOT1 (N4383, N4377);
buf BUF1 (N4384, N4380);
and AND2 (N4385, N4382, N684);
nand NAND3 (N4386, N4384, N539, N309);
nor NOR4 (N4387, N4374, N2962, N568, N1896);
xor XOR2 (N4388, N4375, N3755);
nor NOR4 (N4389, N4388, N314, N2775, N2912);
nor NOR4 (N4390, N4381, N2569, N3033, N2378);
and AND2 (N4391, N4390, N724);
buf BUF1 (N4392, N4366);
buf BUF1 (N4393, N4391);
not NOT1 (N4394, N4386);
nand NAND4 (N4395, N4394, N366, N2613, N2759);
not NOT1 (N4396, N4383);
and AND4 (N4397, N4362, N1541, N2488, N28);
nand NAND3 (N4398, N4389, N3558, N3327);
nand NAND2 (N4399, N4369, N2209);
not NOT1 (N4400, N4398);
and AND3 (N4401, N4392, N3995, N2151);
nand NAND2 (N4402, N4400, N2893);
and AND2 (N4403, N4370, N3889);
nand NAND2 (N4404, N4399, N4181);
buf BUF1 (N4405, N4385);
and AND2 (N4406, N4387, N2738);
nor NOR3 (N4407, N4397, N1415, N4347);
or OR4 (N4408, N4407, N2104, N159, N1747);
buf BUF1 (N4409, N4401);
xor XOR2 (N4410, N4393, N4161);
buf BUF1 (N4411, N4409);
not NOT1 (N4412, N4411);
or OR2 (N4413, N4403, N1811);
not NOT1 (N4414, N4405);
and AND4 (N4415, N4404, N29, N4021, N2552);
xor XOR2 (N4416, N4412, N3013);
nand NAND3 (N4417, N4413, N107, N4019);
buf BUF1 (N4418, N4416);
nand NAND2 (N4419, N4410, N1994);
or OR2 (N4420, N4396, N3744);
and AND4 (N4421, N4406, N3561, N1057, N2070);
xor XOR2 (N4422, N4420, N4371);
xor XOR2 (N4423, N4418, N2753);
nor NOR2 (N4424, N4414, N1155);
nand NAND2 (N4425, N4424, N2331);
buf BUF1 (N4426, N4423);
or OR2 (N4427, N4408, N924);
not NOT1 (N4428, N4417);
and AND2 (N4429, N4415, N4081);
or OR2 (N4430, N4422, N1237);
or OR2 (N4431, N4425, N3787);
xor XOR2 (N4432, N4431, N469);
not NOT1 (N4433, N4430);
nor NOR4 (N4434, N4421, N3693, N2785, N765);
and AND4 (N4435, N4419, N2937, N2955, N584);
buf BUF1 (N4436, N4426);
not NOT1 (N4437, N4435);
nand NAND3 (N4438, N4436, N1507, N1471);
buf BUF1 (N4439, N4434);
not NOT1 (N4440, N4402);
buf BUF1 (N4441, N4428);
nor NOR3 (N4442, N4438, N56, N4335);
or OR3 (N4443, N4433, N4364, N1662);
nor NOR3 (N4444, N4437, N4271, N2260);
nand NAND4 (N4445, N4432, N2557, N3453, N4099);
buf BUF1 (N4446, N4440);
xor XOR2 (N4447, N4444, N2111);
buf BUF1 (N4448, N4447);
nor NOR2 (N4449, N4445, N3125);
buf BUF1 (N4450, N4427);
or OR4 (N4451, N4446, N2646, N2694, N1767);
and AND2 (N4452, N4395, N744);
or OR2 (N4453, N4441, N2637);
buf BUF1 (N4454, N4448);
buf BUF1 (N4455, N4449);
and AND3 (N4456, N4439, N207, N2718);
and AND4 (N4457, N4454, N3222, N1505, N3565);
nor NOR3 (N4458, N4429, N2078, N3354);
and AND4 (N4459, N4453, N4381, N3479, N2969);
and AND4 (N4460, N4452, N458, N2603, N2864);
not NOT1 (N4461, N4443);
nand NAND4 (N4462, N4442, N3092, N4203, N4131);
or OR4 (N4463, N4450, N3123, N847, N2472);
buf BUF1 (N4464, N4458);
xor XOR2 (N4465, N4463, N821);
nand NAND2 (N4466, N4459, N1733);
nor NOR4 (N4467, N4464, N3524, N2079, N3639);
nand NAND2 (N4468, N4461, N3845);
xor XOR2 (N4469, N4462, N957);
xor XOR2 (N4470, N4456, N3852);
xor XOR2 (N4471, N4470, N2058);
nor NOR4 (N4472, N4469, N1449, N2534, N650);
nor NOR3 (N4473, N4471, N1734, N3566);
not NOT1 (N4474, N4451);
or OR2 (N4475, N4467, N3823);
and AND2 (N4476, N4455, N1275);
xor XOR2 (N4477, N4473, N1808);
nor NOR4 (N4478, N4472, N185, N2941, N1687);
buf BUF1 (N4479, N4457);
and AND4 (N4480, N4466, N2836, N2937, N4254);
nand NAND2 (N4481, N4468, N2120);
and AND4 (N4482, N4477, N679, N1343, N2855);
not NOT1 (N4483, N4479);
nand NAND2 (N4484, N4481, N581);
and AND2 (N4485, N4465, N2427);
nor NOR3 (N4486, N4476, N2978, N2274);
nand NAND4 (N4487, N4482, N3807, N2978, N1674);
nor NOR4 (N4488, N4478, N1252, N1831, N3429);
buf BUF1 (N4489, N4486);
buf BUF1 (N4490, N4487);
buf BUF1 (N4491, N4485);
and AND2 (N4492, N4474, N877);
buf BUF1 (N4493, N4483);
not NOT1 (N4494, N4480);
not NOT1 (N4495, N4484);
or OR4 (N4496, N4460, N4182, N808, N1556);
nand NAND3 (N4497, N4495, N1640, N272);
nand NAND4 (N4498, N4492, N4092, N936, N1803);
or OR3 (N4499, N4497, N1673, N4173);
and AND2 (N4500, N4489, N875);
not NOT1 (N4501, N4496);
nand NAND3 (N4502, N4493, N671, N1837);
xor XOR2 (N4503, N4491, N354);
nand NAND3 (N4504, N4475, N589, N3417);
buf BUF1 (N4505, N4490);
xor XOR2 (N4506, N4501, N1514);
and AND2 (N4507, N4505, N1508);
nand NAND3 (N4508, N4503, N619, N2542);
not NOT1 (N4509, N4502);
or OR4 (N4510, N4488, N1523, N218, N4321);
nand NAND3 (N4511, N4509, N4463, N3918);
nor NOR4 (N4512, N4506, N432, N2060, N2866);
or OR4 (N4513, N4511, N2726, N1467, N3250);
not NOT1 (N4514, N4510);
and AND4 (N4515, N4500, N4001, N1445, N3377);
xor XOR2 (N4516, N4508, N2401);
nor NOR3 (N4517, N4499, N573, N582);
buf BUF1 (N4518, N4512);
or OR3 (N4519, N4498, N2103, N186);
nand NAND4 (N4520, N4494, N1340, N4366, N1048);
or OR4 (N4521, N4516, N1286, N1263, N3405);
nor NOR2 (N4522, N4513, N3190);
or OR2 (N4523, N4517, N2748);
buf BUF1 (N4524, N4520);
buf BUF1 (N4525, N4518);
buf BUF1 (N4526, N4523);
nor NOR2 (N4527, N4525, N1332);
and AND3 (N4528, N4515, N2251, N738);
nor NOR3 (N4529, N4521, N1129, N1518);
buf BUF1 (N4530, N4514);
xor XOR2 (N4531, N4504, N929);
not NOT1 (N4532, N4528);
or OR3 (N4533, N4532, N4125, N4503);
xor XOR2 (N4534, N4527, N3639);
xor XOR2 (N4535, N4533, N2408);
or OR2 (N4536, N4524, N2125);
xor XOR2 (N4537, N4534, N579);
nand NAND3 (N4538, N4536, N3699, N4173);
nor NOR4 (N4539, N4538, N683, N13, N2441);
not NOT1 (N4540, N4537);
and AND4 (N4541, N4530, N2383, N3721, N1399);
xor XOR2 (N4542, N4540, N1864);
buf BUF1 (N4543, N4526);
or OR4 (N4544, N4535, N2192, N941, N3568);
buf BUF1 (N4545, N4542);
and AND2 (N4546, N4543, N1627);
or OR2 (N4547, N4546, N2387);
nand NAND4 (N4548, N4545, N2438, N3975, N4359);
nor NOR2 (N4549, N4541, N3945);
or OR2 (N4550, N4539, N347);
nand NAND3 (N4551, N4531, N3925, N3329);
nor NOR4 (N4552, N4544, N3486, N2161, N1747);
and AND4 (N4553, N4549, N1886, N1489, N40);
nand NAND4 (N4554, N4550, N3910, N4353, N1508);
and AND4 (N4555, N4522, N1613, N1084, N2814);
xor XOR2 (N4556, N4529, N3633);
buf BUF1 (N4557, N4548);
or OR4 (N4558, N4557, N2981, N4001, N865);
and AND3 (N4559, N4519, N2955, N1903);
or OR2 (N4560, N4547, N3567);
nand NAND2 (N4561, N4554, N1288);
xor XOR2 (N4562, N4560, N142);
xor XOR2 (N4563, N4555, N1724);
not NOT1 (N4564, N4551);
buf BUF1 (N4565, N4559);
or OR4 (N4566, N4552, N3952, N2489, N2001);
or OR3 (N4567, N4565, N3216, N2416);
not NOT1 (N4568, N4561);
nor NOR3 (N4569, N4563, N4451, N2493);
or OR2 (N4570, N4507, N2901);
buf BUF1 (N4571, N4566);
not NOT1 (N4572, N4569);
nand NAND3 (N4573, N4567, N3772, N3617);
nand NAND4 (N4574, N4562, N1559, N3324, N3778);
nand NAND2 (N4575, N4558, N3783);
nand NAND3 (N4576, N4574, N1207, N2820);
not NOT1 (N4577, N4568);
not NOT1 (N4578, N4553);
not NOT1 (N4579, N4575);
or OR2 (N4580, N4576, N2059);
nor NOR2 (N4581, N4577, N966);
buf BUF1 (N4582, N4579);
or OR4 (N4583, N4573, N980, N1143, N4468);
nand NAND2 (N4584, N4578, N670);
buf BUF1 (N4585, N4571);
or OR2 (N4586, N4564, N488);
xor XOR2 (N4587, N4556, N1884);
not NOT1 (N4588, N4582);
not NOT1 (N4589, N4572);
buf BUF1 (N4590, N4584);
not NOT1 (N4591, N4581);
nand NAND4 (N4592, N4591, N934, N923, N3244);
not NOT1 (N4593, N4588);
buf BUF1 (N4594, N4587);
and AND2 (N4595, N4583, N2435);
or OR4 (N4596, N4570, N2760, N4123, N472);
and AND2 (N4597, N4592, N1607);
buf BUF1 (N4598, N4586);
nand NAND3 (N4599, N4590, N3546, N2761);
not NOT1 (N4600, N4585);
or OR3 (N4601, N4596, N1760, N4125);
and AND2 (N4602, N4600, N284);
nand NAND3 (N4603, N4598, N4045, N3797);
xor XOR2 (N4604, N4589, N3517);
not NOT1 (N4605, N4594);
buf BUF1 (N4606, N4604);
or OR4 (N4607, N4595, N2377, N3048, N1901);
and AND4 (N4608, N4593, N2596, N2332, N3612);
not NOT1 (N4609, N4606);
buf BUF1 (N4610, N4601);
buf BUF1 (N4611, N4580);
or OR4 (N4612, N4610, N3356, N4233, N2213);
nand NAND2 (N4613, N4611, N2294);
or OR3 (N4614, N4605, N2019, N4256);
and AND4 (N4615, N4602, N2884, N3393, N326);
xor XOR2 (N4616, N4612, N2583);
nand NAND2 (N4617, N4597, N2663);
nor NOR2 (N4618, N4607, N1302);
or OR3 (N4619, N4616, N3536, N4407);
or OR2 (N4620, N4599, N2870);
not NOT1 (N4621, N4618);
xor XOR2 (N4622, N4615, N3549);
buf BUF1 (N4623, N4609);
xor XOR2 (N4624, N4622, N260);
and AND3 (N4625, N4617, N4224, N160);
or OR4 (N4626, N4608, N434, N2440, N4625);
buf BUF1 (N4627, N2520);
or OR3 (N4628, N4613, N2759, N3142);
and AND2 (N4629, N4626, N3518);
nor NOR2 (N4630, N4603, N368);
xor XOR2 (N4631, N4627, N1175);
nand NAND4 (N4632, N4619, N472, N2742, N214);
or OR2 (N4633, N4620, N1399);
nand NAND4 (N4634, N4631, N2897, N2884, N4618);
or OR2 (N4635, N4630, N4485);
not NOT1 (N4636, N4624);
nand NAND4 (N4637, N4633, N137, N2422, N381);
and AND4 (N4638, N4629, N1035, N3027, N4040);
nand NAND2 (N4639, N4634, N3747);
xor XOR2 (N4640, N4637, N1040);
not NOT1 (N4641, N4635);
and AND3 (N4642, N4641, N1393, N2903);
buf BUF1 (N4643, N4623);
nor NOR3 (N4644, N4614, N3885, N2209);
not NOT1 (N4645, N4632);
xor XOR2 (N4646, N4645, N3680);
nor NOR3 (N4647, N4639, N3167, N4254);
or OR3 (N4648, N4621, N4575, N976);
buf BUF1 (N4649, N4628);
buf BUF1 (N4650, N4646);
xor XOR2 (N4651, N4649, N3926);
not NOT1 (N4652, N4647);
and AND4 (N4653, N4643, N3433, N1646, N1003);
buf BUF1 (N4654, N4652);
or OR3 (N4655, N4648, N1276, N884);
buf BUF1 (N4656, N4650);
buf BUF1 (N4657, N4640);
not NOT1 (N4658, N4655);
nor NOR4 (N4659, N4642, N2362, N1567, N874);
not NOT1 (N4660, N4651);
nand NAND3 (N4661, N4654, N2576, N1082);
and AND3 (N4662, N4653, N4342, N2535);
or OR4 (N4663, N4659, N2190, N4368, N3704);
or OR3 (N4664, N4657, N1591, N508);
or OR2 (N4665, N4656, N3782);
xor XOR2 (N4666, N4638, N749);
nand NAND3 (N4667, N4662, N3139, N4396);
buf BUF1 (N4668, N4664);
nor NOR2 (N4669, N4661, N3057);
nor NOR2 (N4670, N4666, N4566);
not NOT1 (N4671, N4636);
buf BUF1 (N4672, N4660);
nor NOR3 (N4673, N4665, N1406, N666);
not NOT1 (N4674, N4671);
buf BUF1 (N4675, N4644);
nand NAND2 (N4676, N4663, N4130);
not NOT1 (N4677, N4673);
not NOT1 (N4678, N4675);
nor NOR2 (N4679, N4672, N154);
or OR2 (N4680, N4676, N1263);
and AND4 (N4681, N4667, N931, N3311, N1877);
not NOT1 (N4682, N4677);
not NOT1 (N4683, N4674);
or OR2 (N4684, N4679, N4029);
and AND4 (N4685, N4681, N3090, N3970, N278);
and AND4 (N4686, N4684, N262, N873, N961);
or OR2 (N4687, N4686, N3787);
xor XOR2 (N4688, N4680, N3980);
not NOT1 (N4689, N4687);
nand NAND3 (N4690, N4685, N3485, N2908);
or OR3 (N4691, N4658, N631, N2745);
and AND2 (N4692, N4669, N4079);
xor XOR2 (N4693, N4692, N1335);
or OR4 (N4694, N4691, N3756, N3761, N1236);
and AND2 (N4695, N4694, N723);
buf BUF1 (N4696, N4695);
xor XOR2 (N4697, N4682, N284);
nand NAND3 (N4698, N4668, N3072, N730);
not NOT1 (N4699, N4696);
or OR3 (N4700, N4698, N3594, N3875);
nand NAND3 (N4701, N4683, N1926, N764);
nand NAND2 (N4702, N4700, N1396);
nor NOR4 (N4703, N4702, N1698, N913, N4207);
xor XOR2 (N4704, N4703, N1728);
and AND4 (N4705, N4697, N1381, N1531, N2674);
not NOT1 (N4706, N4690);
nor NOR3 (N4707, N4693, N3520, N3883);
and AND3 (N4708, N4705, N3039, N897);
not NOT1 (N4709, N4670);
or OR4 (N4710, N4678, N697, N2750, N986);
and AND2 (N4711, N4706, N4347);
xor XOR2 (N4712, N4708, N436);
nand NAND4 (N4713, N4704, N1640, N3021, N1254);
not NOT1 (N4714, N4688);
nand NAND2 (N4715, N4710, N3188);
or OR4 (N4716, N4699, N3732, N4479, N2106);
or OR2 (N4717, N4707, N491);
nor NOR2 (N4718, N4717, N3299);
or OR2 (N4719, N4712, N3149);
and AND2 (N4720, N4715, N4580);
buf BUF1 (N4721, N4720);
nand NAND3 (N4722, N4711, N4514, N1251);
nand NAND3 (N4723, N4722, N3314, N2095);
and AND2 (N4724, N4723, N2421);
xor XOR2 (N4725, N4724, N4697);
nor NOR4 (N4726, N4721, N4299, N1352, N2642);
nand NAND4 (N4727, N4701, N809, N2825, N712);
nor NOR2 (N4728, N4689, N280);
and AND3 (N4729, N4726, N3352, N4140);
xor XOR2 (N4730, N4725, N765);
and AND4 (N4731, N4730, N2819, N619, N1946);
not NOT1 (N4732, N4714);
not NOT1 (N4733, N4719);
not NOT1 (N4734, N4732);
not NOT1 (N4735, N4731);
and AND2 (N4736, N4735, N3017);
buf BUF1 (N4737, N4736);
xor XOR2 (N4738, N4713, N1677);
nor NOR2 (N4739, N4718, N3057);
or OR2 (N4740, N4737, N3063);
nor NOR4 (N4741, N4729, N1864, N3981, N2246);
buf BUF1 (N4742, N4738);
and AND4 (N4743, N4734, N4281, N2315, N3232);
nand NAND3 (N4744, N4741, N212, N2031);
xor XOR2 (N4745, N4733, N2548);
buf BUF1 (N4746, N4727);
not NOT1 (N4747, N4739);
or OR2 (N4748, N4742, N776);
and AND2 (N4749, N4747, N1481);
and AND3 (N4750, N4743, N4130, N3983);
xor XOR2 (N4751, N4746, N3810);
not NOT1 (N4752, N4751);
xor XOR2 (N4753, N4745, N2112);
nand NAND2 (N4754, N4709, N4293);
or OR4 (N4755, N4753, N4450, N2558, N3038);
buf BUF1 (N4756, N4748);
nor NOR3 (N4757, N4749, N4711, N462);
xor XOR2 (N4758, N4757, N203);
nor NOR4 (N4759, N4728, N759, N3171, N2786);
not NOT1 (N4760, N4754);
and AND2 (N4761, N4740, N2023);
and AND4 (N4762, N4744, N1497, N2603, N2178);
not NOT1 (N4763, N4750);
or OR4 (N4764, N4763, N1469, N4627, N303);
buf BUF1 (N4765, N4761);
nand NAND2 (N4766, N4760, N2507);
not NOT1 (N4767, N4766);
xor XOR2 (N4768, N4762, N2364);
and AND3 (N4769, N4764, N1997, N3121);
or OR2 (N4770, N4716, N4343);
xor XOR2 (N4771, N4769, N4454);
xor XOR2 (N4772, N4759, N4544);
xor XOR2 (N4773, N4768, N815);
buf BUF1 (N4774, N4770);
buf BUF1 (N4775, N4756);
nand NAND3 (N4776, N4774, N4527, N1546);
or OR2 (N4777, N4758, N4118);
xor XOR2 (N4778, N4777, N786);
nand NAND3 (N4779, N4778, N4056, N4450);
nand NAND2 (N4780, N4779, N2539);
or OR2 (N4781, N4771, N342);
not NOT1 (N4782, N4755);
nand NAND3 (N4783, N4772, N2523, N1917);
buf BUF1 (N4784, N4752);
nand NAND3 (N4785, N4776, N1371, N2065);
xor XOR2 (N4786, N4783, N1892);
nand NAND3 (N4787, N4780, N1235, N1145);
and AND2 (N4788, N4786, N4284);
nand NAND4 (N4789, N4788, N2017, N3063, N2837);
xor XOR2 (N4790, N4784, N534);
buf BUF1 (N4791, N4785);
or OR4 (N4792, N4791, N1465, N741, N3750);
not NOT1 (N4793, N4767);
xor XOR2 (N4794, N4775, N3518);
nand NAND2 (N4795, N4794, N746);
not NOT1 (N4796, N4781);
nor NOR4 (N4797, N4782, N3648, N2080, N4312);
and AND4 (N4798, N4789, N1913, N1546, N1328);
nand NAND3 (N4799, N4793, N2977, N3316);
nor NOR4 (N4800, N4787, N3497, N3562, N3519);
and AND4 (N4801, N4792, N1203, N4544, N1818);
nor NOR3 (N4802, N4790, N2052, N2872);
nand NAND3 (N4803, N4801, N519, N3557);
nor NOR4 (N4804, N4796, N1596, N2562, N1454);
xor XOR2 (N4805, N4804, N1348);
buf BUF1 (N4806, N4798);
nand NAND4 (N4807, N4803, N4090, N1435, N3888);
nand NAND4 (N4808, N4807, N982, N2287, N171);
buf BUF1 (N4809, N4806);
nand NAND4 (N4810, N4805, N1413, N2658, N2909);
not NOT1 (N4811, N4802);
nor NOR4 (N4812, N4765, N1179, N54, N831);
xor XOR2 (N4813, N4810, N1434);
and AND4 (N4814, N4811, N3551, N3107, N628);
xor XOR2 (N4815, N4797, N3290);
xor XOR2 (N4816, N4773, N4400);
nand NAND2 (N4817, N4816, N3529);
nor NOR3 (N4818, N4800, N1929, N2531);
nand NAND4 (N4819, N4795, N4796, N3224, N838);
and AND4 (N4820, N4813, N1484, N564, N1604);
nor NOR3 (N4821, N4815, N2431, N3069);
and AND3 (N4822, N4808, N2270, N136);
and AND2 (N4823, N4820, N4167);
nand NAND2 (N4824, N4812, N723);
or OR2 (N4825, N4822, N1119);
nor NOR2 (N4826, N4825, N254);
buf BUF1 (N4827, N4826);
buf BUF1 (N4828, N4809);
nor NOR2 (N4829, N4818, N4302);
nor NOR4 (N4830, N4814, N2432, N1339, N4543);
buf BUF1 (N4831, N4827);
and AND2 (N4832, N4821, N804);
xor XOR2 (N4833, N4832, N980);
or OR2 (N4834, N4831, N610);
not NOT1 (N4835, N4834);
and AND4 (N4836, N4830, N2968, N4533, N87);
xor XOR2 (N4837, N4828, N4553);
not NOT1 (N4838, N4837);
nor NOR2 (N4839, N4819, N3127);
not NOT1 (N4840, N4799);
or OR4 (N4841, N4817, N3331, N4031, N563);
buf BUF1 (N4842, N4833);
buf BUF1 (N4843, N4842);
buf BUF1 (N4844, N4829);
nor NOR2 (N4845, N4840, N1439);
buf BUF1 (N4846, N4844);
and AND3 (N4847, N4824, N3134, N1289);
or OR2 (N4848, N4838, N435);
nor NOR2 (N4849, N4836, N2786);
xor XOR2 (N4850, N4848, N1892);
or OR2 (N4851, N4847, N4363);
xor XOR2 (N4852, N4850, N2831);
nand NAND3 (N4853, N4843, N739, N613);
and AND3 (N4854, N4853, N573, N1017);
not NOT1 (N4855, N4841);
nand NAND4 (N4856, N4823, N2938, N3790, N1015);
and AND2 (N4857, N4835, N4652);
and AND3 (N4858, N4849, N1910, N2970);
nand NAND4 (N4859, N4855, N3428, N3915, N3841);
not NOT1 (N4860, N4839);
or OR4 (N4861, N4859, N345, N4432, N1272);
or OR3 (N4862, N4854, N357, N4443);
buf BUF1 (N4863, N4860);
buf BUF1 (N4864, N4846);
nand NAND3 (N4865, N4851, N2784, N621);
or OR4 (N4866, N4856, N952, N28, N2657);
or OR4 (N4867, N4865, N4058, N2650, N3719);
not NOT1 (N4868, N4852);
or OR4 (N4869, N4867, N3562, N3390, N2301);
xor XOR2 (N4870, N4861, N3272);
nand NAND4 (N4871, N4866, N2928, N227, N1904);
not NOT1 (N4872, N4869);
or OR3 (N4873, N4857, N2457, N3096);
and AND3 (N4874, N4872, N2938, N1960);
buf BUF1 (N4875, N4873);
xor XOR2 (N4876, N4863, N2561);
not NOT1 (N4877, N4875);
and AND3 (N4878, N4876, N529, N1324);
xor XOR2 (N4879, N4864, N1152);
xor XOR2 (N4880, N4862, N227);
and AND3 (N4881, N4880, N3627, N26);
or OR2 (N4882, N4868, N3102);
xor XOR2 (N4883, N4871, N2799);
nor NOR2 (N4884, N4874, N1692);
not NOT1 (N4885, N4877);
or OR3 (N4886, N4858, N2976, N1123);
nor NOR4 (N4887, N4878, N2553, N3084, N2688);
and AND3 (N4888, N4886, N610, N4794);
and AND4 (N4889, N4884, N2727, N3736, N3731);
buf BUF1 (N4890, N4888);
or OR2 (N4891, N4870, N973);
nor NOR2 (N4892, N4845, N772);
or OR3 (N4893, N4883, N1809, N867);
or OR3 (N4894, N4890, N4622, N1284);
buf BUF1 (N4895, N4894);
nand NAND2 (N4896, N4885, N2180);
or OR4 (N4897, N4893, N165, N306, N1505);
not NOT1 (N4898, N4897);
buf BUF1 (N4899, N4892);
or OR3 (N4900, N4895, N3313, N857);
or OR4 (N4901, N4882, N1607, N462, N4521);
not NOT1 (N4902, N4887);
and AND3 (N4903, N4889, N2529, N866);
nor NOR4 (N4904, N4901, N3054, N3140, N1594);
nand NAND3 (N4905, N4898, N4742, N1443);
nor NOR2 (N4906, N4905, N2858);
nand NAND3 (N4907, N4903, N2692, N533);
nand NAND3 (N4908, N4879, N3659, N4726);
nor NOR3 (N4909, N4902, N1709, N3301);
buf BUF1 (N4910, N4909);
or OR3 (N4911, N4899, N1362, N2299);
xor XOR2 (N4912, N4891, N1742);
or OR4 (N4913, N4910, N442, N1809, N3858);
xor XOR2 (N4914, N4907, N770);
or OR2 (N4915, N4912, N4853);
buf BUF1 (N4916, N4904);
xor XOR2 (N4917, N4900, N3280);
xor XOR2 (N4918, N4881, N3891);
not NOT1 (N4919, N4908);
buf BUF1 (N4920, N4919);
buf BUF1 (N4921, N4906);
buf BUF1 (N4922, N4920);
and AND4 (N4923, N4913, N4545, N4378, N4794);
or OR4 (N4924, N4923, N834, N2097, N213);
or OR2 (N4925, N4916, N55);
nand NAND4 (N4926, N4915, N1696, N2444, N3721);
or OR2 (N4927, N4925, N125);
buf BUF1 (N4928, N4921);
buf BUF1 (N4929, N4922);
and AND3 (N4930, N4928, N1170, N4871);
nand NAND3 (N4931, N4926, N1082, N1694);
xor XOR2 (N4932, N4917, N1276);
buf BUF1 (N4933, N4929);
nor NOR3 (N4934, N4927, N3365, N2421);
or OR4 (N4935, N4914, N2231, N229, N1876);
nand NAND2 (N4936, N4918, N2495);
nor NOR4 (N4937, N4936, N1963, N2729, N3542);
xor XOR2 (N4938, N4924, N4246);
not NOT1 (N4939, N4935);
nand NAND3 (N4940, N4930, N2645, N3300);
and AND2 (N4941, N4933, N2057);
nand NAND4 (N4942, N4940, N2612, N1561, N3538);
nand NAND3 (N4943, N4896, N1713, N481);
nand NAND2 (N4944, N4938, N1902);
buf BUF1 (N4945, N4937);
buf BUF1 (N4946, N4941);
nor NOR4 (N4947, N4945, N3778, N1326, N3399);
nand NAND2 (N4948, N4942, N2107);
xor XOR2 (N4949, N4944, N4223);
not NOT1 (N4950, N4934);
nand NAND4 (N4951, N4946, N4752, N3672, N1739);
buf BUF1 (N4952, N4943);
nand NAND4 (N4953, N4949, N2305, N2856, N939);
not NOT1 (N4954, N4951);
not NOT1 (N4955, N4953);
nor NOR3 (N4956, N4911, N2232, N4241);
nor NOR3 (N4957, N4948, N3992, N4135);
nand NAND4 (N4958, N4952, N1047, N273, N2210);
xor XOR2 (N4959, N4931, N908);
and AND4 (N4960, N4932, N2551, N2190, N326);
buf BUF1 (N4961, N4950);
buf BUF1 (N4962, N4960);
and AND3 (N4963, N4957, N2937, N3553);
buf BUF1 (N4964, N4956);
nand NAND3 (N4965, N4955, N1217, N2920);
nand NAND3 (N4966, N4958, N2373, N1072);
not NOT1 (N4967, N4939);
or OR3 (N4968, N4959, N2043, N4346);
not NOT1 (N4969, N4964);
nor NOR3 (N4970, N4963, N4468, N4041);
nor NOR4 (N4971, N4967, N1843, N1820, N4072);
or OR4 (N4972, N4970, N546, N206, N4456);
buf BUF1 (N4973, N4971);
buf BUF1 (N4974, N4961);
not NOT1 (N4975, N4968);
not NOT1 (N4976, N4965);
nor NOR3 (N4977, N4969, N4016, N3705);
and AND2 (N4978, N4972, N2191);
buf BUF1 (N4979, N4973);
or OR4 (N4980, N4975, N699, N1783, N778);
not NOT1 (N4981, N4976);
and AND3 (N4982, N4947, N3010, N1522);
xor XOR2 (N4983, N4966, N3091);
or OR3 (N4984, N4983, N1608, N2442);
or OR3 (N4985, N4984, N3696, N1521);
buf BUF1 (N4986, N4962);
nand NAND4 (N4987, N4980, N1587, N3120, N3900);
or OR3 (N4988, N4981, N4045, N1559);
nand NAND3 (N4989, N4974, N4764, N262);
nor NOR3 (N4990, N4978, N430, N3463);
xor XOR2 (N4991, N4954, N226);
xor XOR2 (N4992, N4988, N2323);
nand NAND4 (N4993, N4992, N1975, N744, N2966);
or OR2 (N4994, N4977, N2074);
and AND4 (N4995, N4987, N2022, N2299, N1295);
buf BUF1 (N4996, N4985);
nand NAND3 (N4997, N4993, N3220, N4062);
nand NAND3 (N4998, N4990, N367, N1694);
nor NOR2 (N4999, N4995, N3023);
not NOT1 (N5000, N4989);
or OR4 (N5001, N4986, N3216, N4055, N2360);
and AND4 (N5002, N4998, N2581, N1924, N1778);
nand NAND4 (N5003, N4991, N321, N2985, N1061);
buf BUF1 (N5004, N4979);
nor NOR2 (N5005, N5004, N4436);
buf BUF1 (N5006, N4999);
buf BUF1 (N5007, N5005);
not NOT1 (N5008, N5006);
nor NOR3 (N5009, N5003, N4985, N3822);
or OR4 (N5010, N4982, N4521, N3930, N4362);
not NOT1 (N5011, N5009);
nor NOR3 (N5012, N5010, N4676, N3108);
buf BUF1 (N5013, N4994);
xor XOR2 (N5014, N5012, N4802);
and AND2 (N5015, N5007, N4913);
or OR3 (N5016, N5013, N3515, N143);
or OR3 (N5017, N5008, N2526, N3114);
nor NOR2 (N5018, N5014, N1781);
nand NAND3 (N5019, N5016, N301, N3075);
buf BUF1 (N5020, N4996);
nand NAND2 (N5021, N5011, N2747);
or OR3 (N5022, N5018, N3245, N3119);
nor NOR3 (N5023, N5021, N3922, N3166);
nor NOR2 (N5024, N5015, N4682);
not NOT1 (N5025, N5001);
or OR2 (N5026, N5023, N3851);
and AND4 (N5027, N5024, N4009, N3510, N3280);
and AND4 (N5028, N5020, N1946, N1994, N2863);
nand NAND4 (N5029, N5028, N3293, N4151, N618);
not NOT1 (N5030, N5027);
nand NAND2 (N5031, N5002, N4088);
buf BUF1 (N5032, N5017);
nor NOR4 (N5033, N5031, N4673, N570, N2251);
buf BUF1 (N5034, N5022);
or OR3 (N5035, N5000, N662, N880);
xor XOR2 (N5036, N5019, N1942);
nor NOR3 (N5037, N5033, N4833, N3621);
or OR3 (N5038, N5034, N3071, N1678);
buf BUF1 (N5039, N5030);
nand NAND2 (N5040, N5026, N1905);
or OR3 (N5041, N5036, N4034, N3005);
not NOT1 (N5042, N5032);
nand NAND2 (N5043, N5029, N2264);
not NOT1 (N5044, N5040);
buf BUF1 (N5045, N5037);
buf BUF1 (N5046, N5035);
or OR2 (N5047, N5025, N3836);
or OR2 (N5048, N4997, N2373);
and AND4 (N5049, N5045, N3660, N2173, N2884);
and AND2 (N5050, N5044, N3214);
xor XOR2 (N5051, N5042, N311);
nor NOR2 (N5052, N5043, N4862);
xor XOR2 (N5053, N5052, N1751);
nor NOR2 (N5054, N5050, N1103);
buf BUF1 (N5055, N5046);
nor NOR4 (N5056, N5047, N1670, N4953, N390);
or OR2 (N5057, N5038, N73);
not NOT1 (N5058, N5053);
not NOT1 (N5059, N5056);
nor NOR3 (N5060, N5057, N4416, N3254);
nor NOR3 (N5061, N5054, N2742, N929);
buf BUF1 (N5062, N5048);
nand NAND3 (N5063, N5049, N1247, N1200);
buf BUF1 (N5064, N5051);
nand NAND2 (N5065, N5061, N643);
nor NOR4 (N5066, N5063, N2934, N3158, N3073);
and AND2 (N5067, N5041, N827);
nor NOR2 (N5068, N5060, N4115);
and AND2 (N5069, N5058, N492);
nor NOR2 (N5070, N5068, N455);
and AND3 (N5071, N5066, N171, N4878);
or OR2 (N5072, N5062, N2505);
buf BUF1 (N5073, N5065);
and AND3 (N5074, N5059, N836, N2830);
not NOT1 (N5075, N5071);
xor XOR2 (N5076, N5073, N2898);
buf BUF1 (N5077, N5039);
nand NAND2 (N5078, N5055, N2221);
or OR3 (N5079, N5070, N3721, N1532);
or OR3 (N5080, N5072, N3009, N3607);
not NOT1 (N5081, N5076);
not NOT1 (N5082, N5069);
nand NAND4 (N5083, N5078, N3844, N4821, N4304);
not NOT1 (N5084, N5064);
nand NAND2 (N5085, N5082, N4264);
nor NOR2 (N5086, N5077, N4472);
not NOT1 (N5087, N5075);
and AND3 (N5088, N5067, N2519, N864);
and AND4 (N5089, N5085, N1650, N1410, N1255);
nand NAND3 (N5090, N5080, N2540, N1334);
xor XOR2 (N5091, N5081, N912);
and AND4 (N5092, N5091, N1370, N1635, N3237);
and AND3 (N5093, N5092, N780, N971);
or OR4 (N5094, N5079, N4886, N4104, N1063);
nand NAND3 (N5095, N5090, N4395, N3427);
nor NOR4 (N5096, N5093, N1400, N94, N2112);
and AND3 (N5097, N5083, N3145, N4789);
nand NAND3 (N5098, N5089, N378, N4390);
not NOT1 (N5099, N5087);
nand NAND4 (N5100, N5084, N4093, N3099, N3127);
xor XOR2 (N5101, N5100, N2658);
buf BUF1 (N5102, N5095);
or OR3 (N5103, N5074, N5051, N3420);
and AND3 (N5104, N5101, N1285, N4900);
nand NAND2 (N5105, N5097, N2642);
or OR2 (N5106, N5086, N592);
or OR2 (N5107, N5105, N4148);
and AND3 (N5108, N5099, N2745, N2943);
xor XOR2 (N5109, N5096, N3302);
not NOT1 (N5110, N5098);
and AND3 (N5111, N5104, N3920, N926);
not NOT1 (N5112, N5106);
nand NAND2 (N5113, N5102, N4629);
or OR4 (N5114, N5110, N4149, N789, N3729);
xor XOR2 (N5115, N5107, N3846);
buf BUF1 (N5116, N5113);
xor XOR2 (N5117, N5116, N2841);
not NOT1 (N5118, N5094);
nor NOR2 (N5119, N5108, N4423);
nand NAND3 (N5120, N5117, N2673, N1641);
buf BUF1 (N5121, N5109);
and AND2 (N5122, N5114, N3962);
buf BUF1 (N5123, N5111);
xor XOR2 (N5124, N5120, N4178);
not NOT1 (N5125, N5121);
xor XOR2 (N5126, N5115, N4532);
not NOT1 (N5127, N5088);
nor NOR2 (N5128, N5126, N4522);
and AND4 (N5129, N5127, N1828, N445, N763);
nand NAND3 (N5130, N5112, N590, N2031);
xor XOR2 (N5131, N5103, N3999);
and AND4 (N5132, N5119, N2975, N3654, N4059);
and AND3 (N5133, N5129, N5063, N3110);
buf BUF1 (N5134, N5125);
nand NAND2 (N5135, N5131, N5025);
or OR2 (N5136, N5130, N4659);
xor XOR2 (N5137, N5134, N3575);
or OR2 (N5138, N5124, N4613);
and AND3 (N5139, N5123, N705, N3287);
not NOT1 (N5140, N5136);
not NOT1 (N5141, N5122);
and AND2 (N5142, N5135, N4196);
xor XOR2 (N5143, N5141, N4009);
or OR4 (N5144, N5118, N3184, N2919, N821);
not NOT1 (N5145, N5137);
and AND3 (N5146, N5139, N1473, N687);
not NOT1 (N5147, N5140);
and AND4 (N5148, N5138, N932, N4241, N1658);
nand NAND3 (N5149, N5143, N1223, N4476);
and AND2 (N5150, N5142, N2177);
nor NOR4 (N5151, N5144, N1131, N4199, N180);
buf BUF1 (N5152, N5146);
or OR2 (N5153, N5152, N4404);
nand NAND3 (N5154, N5128, N2444, N1304);
nor NOR4 (N5155, N5149, N365, N3178, N2324);
not NOT1 (N5156, N5153);
nand NAND4 (N5157, N5148, N4639, N915, N4311);
or OR2 (N5158, N5150, N4781);
or OR4 (N5159, N5151, N70, N1508, N2308);
nor NOR4 (N5160, N5157, N2390, N4115, N1797);
buf BUF1 (N5161, N5133);
and AND3 (N5162, N5158, N4374, N1922);
xor XOR2 (N5163, N5132, N4450);
nor NOR3 (N5164, N5161, N750, N2453);
not NOT1 (N5165, N5160);
xor XOR2 (N5166, N5156, N3622);
buf BUF1 (N5167, N5147);
buf BUF1 (N5168, N5162);
nand NAND3 (N5169, N5166, N4641, N1752);
and AND3 (N5170, N5145, N2301, N2552);
or OR2 (N5171, N5169, N3115);
or OR4 (N5172, N5159, N2789, N4972, N2946);
or OR2 (N5173, N5168, N3548);
xor XOR2 (N5174, N5170, N3742);
nor NOR4 (N5175, N5171, N1818, N419, N1014);
buf BUF1 (N5176, N5165);
nand NAND3 (N5177, N5163, N921, N1342);
nor NOR3 (N5178, N5174, N3760, N3601);
buf BUF1 (N5179, N5155);
or OR4 (N5180, N5164, N1185, N2703, N274);
nand NAND2 (N5181, N5167, N794);
xor XOR2 (N5182, N5172, N1142);
nor NOR4 (N5183, N5175, N1120, N5174, N2895);
nor NOR2 (N5184, N5176, N2047);
and AND4 (N5185, N5154, N1979, N4839, N4324);
and AND4 (N5186, N5182, N4999, N3624, N709);
not NOT1 (N5187, N5186);
not NOT1 (N5188, N5183);
or OR3 (N5189, N5188, N5074, N3686);
and AND2 (N5190, N5181, N1443);
not NOT1 (N5191, N5178);
buf BUF1 (N5192, N5180);
xor XOR2 (N5193, N5192, N2153);
xor XOR2 (N5194, N5187, N4033);
or OR4 (N5195, N5173, N1031, N3571, N3755);
or OR2 (N5196, N5193, N877);
buf BUF1 (N5197, N5177);
nand NAND2 (N5198, N5189, N2717);
xor XOR2 (N5199, N5185, N2812);
xor XOR2 (N5200, N5190, N2690);
or OR3 (N5201, N5199, N940, N5035);
and AND3 (N5202, N5184, N4734, N1155);
buf BUF1 (N5203, N5200);
not NOT1 (N5204, N5191);
or OR3 (N5205, N5202, N4044, N275);
buf BUF1 (N5206, N5197);
buf BUF1 (N5207, N5203);
and AND2 (N5208, N5206, N56);
not NOT1 (N5209, N5207);
nor NOR3 (N5210, N5198, N2356, N362);
xor XOR2 (N5211, N5210, N604);
nor NOR3 (N5212, N5204, N3938, N1177);
buf BUF1 (N5213, N5196);
buf BUF1 (N5214, N5212);
and AND3 (N5215, N5201, N4606, N463);
or OR3 (N5216, N5211, N2389, N5109);
not NOT1 (N5217, N5216);
buf BUF1 (N5218, N5179);
nand NAND4 (N5219, N5213, N3269, N428, N1104);
and AND2 (N5220, N5215, N843);
buf BUF1 (N5221, N5194);
not NOT1 (N5222, N5214);
nand NAND2 (N5223, N5218, N1406);
or OR3 (N5224, N5208, N1259, N1624);
xor XOR2 (N5225, N5221, N3562);
buf BUF1 (N5226, N5220);
not NOT1 (N5227, N5223);
nand NAND3 (N5228, N5227, N2331, N1559);
nor NOR2 (N5229, N5205, N664);
buf BUF1 (N5230, N5224);
nor NOR4 (N5231, N5225, N1252, N1266, N4672);
buf BUF1 (N5232, N5209);
nor NOR2 (N5233, N5217, N684);
and AND2 (N5234, N5226, N372);
xor XOR2 (N5235, N5229, N4049);
or OR4 (N5236, N5234, N1769, N3074, N3080);
buf BUF1 (N5237, N5230);
and AND2 (N5238, N5235, N1581);
and AND3 (N5239, N5231, N27, N3172);
nor NOR2 (N5240, N5236, N2996);
xor XOR2 (N5241, N5239, N960);
nand NAND2 (N5242, N5237, N3657);
and AND3 (N5243, N5238, N2723, N449);
or OR4 (N5244, N5240, N2074, N1615, N4365);
nor NOR4 (N5245, N5243, N3118, N1303, N1813);
and AND2 (N5246, N5228, N4734);
and AND3 (N5247, N5195, N3802, N4610);
or OR3 (N5248, N5233, N1967, N428);
not NOT1 (N5249, N5222);
and AND2 (N5250, N5245, N2487);
not NOT1 (N5251, N5232);
and AND3 (N5252, N5219, N1341, N1525);
buf BUF1 (N5253, N5241);
buf BUF1 (N5254, N5248);
nand NAND3 (N5255, N5250, N1103, N1909);
and AND2 (N5256, N5242, N4126);
not NOT1 (N5257, N5256);
xor XOR2 (N5258, N5254, N1682);
nand NAND4 (N5259, N5252, N178, N1911, N3013);
or OR3 (N5260, N5255, N2981, N4604);
not NOT1 (N5261, N5257);
nor NOR3 (N5262, N5261, N4008, N1640);
or OR2 (N5263, N5253, N435);
xor XOR2 (N5264, N5247, N1940);
nor NOR2 (N5265, N5246, N1107);
xor XOR2 (N5266, N5258, N3266);
nor NOR3 (N5267, N5265, N4562, N4898);
buf BUF1 (N5268, N5244);
buf BUF1 (N5269, N5251);
buf BUF1 (N5270, N5267);
nor NOR3 (N5271, N5264, N4771, N956);
or OR3 (N5272, N5260, N561, N2708);
or OR2 (N5273, N5259, N179);
nor NOR3 (N5274, N5249, N4125, N650);
nor NOR4 (N5275, N5273, N1166, N1779, N2750);
nor NOR2 (N5276, N5268, N3884);
xor XOR2 (N5277, N5262, N1994);
or OR3 (N5278, N5272, N3448, N3972);
nand NAND4 (N5279, N5266, N5192, N1761, N3484);
or OR2 (N5280, N5275, N4067);
not NOT1 (N5281, N5263);
and AND4 (N5282, N5278, N1322, N2415, N3695);
or OR2 (N5283, N5274, N1075);
or OR3 (N5284, N5283, N846, N5072);
nor NOR3 (N5285, N5270, N1909, N4158);
nor NOR2 (N5286, N5282, N4050);
xor XOR2 (N5287, N5285, N2841);
nor NOR2 (N5288, N5269, N4809);
and AND2 (N5289, N5279, N4554);
or OR3 (N5290, N5284, N522, N1223);
and AND2 (N5291, N5290, N1361);
nand NAND4 (N5292, N5271, N2806, N4600, N515);
xor XOR2 (N5293, N5287, N2404);
and AND4 (N5294, N5281, N2835, N4779, N3109);
buf BUF1 (N5295, N5294);
buf BUF1 (N5296, N5289);
or OR4 (N5297, N5288, N2262, N1828, N5277);
and AND4 (N5298, N4228, N3261, N144, N1419);
or OR2 (N5299, N5293, N3486);
or OR3 (N5300, N5286, N5048, N438);
and AND4 (N5301, N5296, N87, N2178, N802);
buf BUF1 (N5302, N5291);
or OR2 (N5303, N5276, N5138);
xor XOR2 (N5304, N5295, N967);
xor XOR2 (N5305, N5302, N2103);
or OR2 (N5306, N5300, N79);
or OR3 (N5307, N5297, N684, N1993);
or OR3 (N5308, N5305, N235, N4651);
not NOT1 (N5309, N5292);
nand NAND4 (N5310, N5280, N1879, N4757, N2217);
buf BUF1 (N5311, N5307);
xor XOR2 (N5312, N5301, N693);
nand NAND4 (N5313, N5298, N2011, N914, N5281);
and AND3 (N5314, N5304, N2076, N503);
and AND4 (N5315, N5306, N2799, N921, N789);
xor XOR2 (N5316, N5314, N2305);
and AND2 (N5317, N5309, N1305);
xor XOR2 (N5318, N5313, N1645);
nand NAND3 (N5319, N5310, N2558, N3336);
and AND2 (N5320, N5311, N4017);
nand NAND2 (N5321, N5308, N1376);
buf BUF1 (N5322, N5303);
not NOT1 (N5323, N5319);
or OR2 (N5324, N5323, N3439);
and AND4 (N5325, N5316, N1308, N2807, N668);
xor XOR2 (N5326, N5317, N308);
and AND3 (N5327, N5299, N1579, N2218);
buf BUF1 (N5328, N5318);
not NOT1 (N5329, N5315);
and AND2 (N5330, N5320, N4397);
nand NAND2 (N5331, N5328, N3670);
not NOT1 (N5332, N5324);
buf BUF1 (N5333, N5329);
buf BUF1 (N5334, N5331);
nand NAND3 (N5335, N5326, N2922, N4251);
buf BUF1 (N5336, N5325);
or OR3 (N5337, N5321, N2884, N1864);
not NOT1 (N5338, N5332);
nor NOR4 (N5339, N5322, N918, N3809, N4972);
or OR3 (N5340, N5330, N293, N2814);
buf BUF1 (N5341, N5333);
nor NOR3 (N5342, N5336, N2871, N2143);
nand NAND2 (N5343, N5334, N832);
and AND2 (N5344, N5343, N3284);
buf BUF1 (N5345, N5327);
not NOT1 (N5346, N5344);
and AND4 (N5347, N5341, N3641, N3236, N3105);
nor NOR3 (N5348, N5345, N155, N2047);
and AND2 (N5349, N5339, N4139);
or OR3 (N5350, N5335, N2830, N1165);
xor XOR2 (N5351, N5340, N5016);
or OR3 (N5352, N5350, N1405, N3742);
xor XOR2 (N5353, N5349, N4953);
or OR4 (N5354, N5351, N3891, N283, N1476);
nor NOR4 (N5355, N5353, N2829, N2909, N2851);
nor NOR3 (N5356, N5347, N4148, N34);
xor XOR2 (N5357, N5338, N3106);
xor XOR2 (N5358, N5342, N2930);
or OR2 (N5359, N5357, N2683);
nand NAND2 (N5360, N5358, N2563);
buf BUF1 (N5361, N5359);
buf BUF1 (N5362, N5356);
nand NAND2 (N5363, N5352, N326);
or OR4 (N5364, N5348, N4602, N2742, N220);
nor NOR2 (N5365, N5354, N5023);
not NOT1 (N5366, N5337);
buf BUF1 (N5367, N5361);
xor XOR2 (N5368, N5364, N1916);
nand NAND4 (N5369, N5365, N1976, N1861, N4135);
xor XOR2 (N5370, N5362, N1458);
buf BUF1 (N5371, N5355);
nand NAND3 (N5372, N5368, N2271, N723);
nor NOR4 (N5373, N5366, N1170, N1170, N1951);
or OR4 (N5374, N5346, N1348, N4416, N4104);
or OR2 (N5375, N5312, N4967);
xor XOR2 (N5376, N5367, N4653);
nand NAND2 (N5377, N5370, N2666);
nor NOR3 (N5378, N5377, N2810, N2953);
buf BUF1 (N5379, N5376);
not NOT1 (N5380, N5360);
buf BUF1 (N5381, N5372);
nand NAND3 (N5382, N5381, N4123, N4029);
or OR3 (N5383, N5363, N97, N2062);
nand NAND2 (N5384, N5373, N1617);
xor XOR2 (N5385, N5378, N1919);
buf BUF1 (N5386, N5383);
xor XOR2 (N5387, N5371, N1826);
xor XOR2 (N5388, N5374, N3890);
nor NOR3 (N5389, N5375, N4085, N4721);
and AND4 (N5390, N5380, N1955, N4695, N1990);
nand NAND4 (N5391, N5388, N3824, N3631, N5170);
not NOT1 (N5392, N5389);
nor NOR3 (N5393, N5385, N3954, N2922);
or OR3 (N5394, N5384, N2110, N1642);
or OR4 (N5395, N5386, N728, N1674, N4454);
not NOT1 (N5396, N5392);
and AND2 (N5397, N5382, N2653);
nor NOR2 (N5398, N5393, N1583);
nor NOR3 (N5399, N5395, N4175, N3845);
not NOT1 (N5400, N5398);
not NOT1 (N5401, N5390);
or OR2 (N5402, N5379, N1423);
nor NOR3 (N5403, N5402, N2279, N2719);
nor NOR2 (N5404, N5403, N4664);
xor XOR2 (N5405, N5404, N3869);
and AND4 (N5406, N5397, N1659, N3690, N2958);
or OR2 (N5407, N5406, N1255);
or OR3 (N5408, N5400, N4689, N4340);
not NOT1 (N5409, N5408);
nand NAND3 (N5410, N5369, N2273, N3049);
nand NAND4 (N5411, N5410, N339, N1257, N3055);
not NOT1 (N5412, N5399);
buf BUF1 (N5413, N5407);
buf BUF1 (N5414, N5405);
not NOT1 (N5415, N5396);
and AND4 (N5416, N5387, N4583, N3892, N3462);
nor NOR4 (N5417, N5391, N899, N4526, N2803);
and AND2 (N5418, N5417, N3525);
not NOT1 (N5419, N5409);
and AND3 (N5420, N5418, N4409, N2331);
xor XOR2 (N5421, N5415, N2844);
not NOT1 (N5422, N5394);
buf BUF1 (N5423, N5411);
nor NOR3 (N5424, N5401, N1556, N1559);
xor XOR2 (N5425, N5414, N4620);
nor NOR4 (N5426, N5413, N4078, N2742, N5241);
nor NOR3 (N5427, N5426, N2293, N3138);
buf BUF1 (N5428, N5419);
not NOT1 (N5429, N5427);
nor NOR2 (N5430, N5412, N4329);
and AND2 (N5431, N5421, N3557);
or OR4 (N5432, N5425, N4292, N4702, N1039);
or OR3 (N5433, N5423, N2138, N3595);
or OR3 (N5434, N5430, N1881, N34);
not NOT1 (N5435, N5416);
nand NAND4 (N5436, N5435, N5303, N2517, N5088);
and AND4 (N5437, N5429, N4940, N533, N4342);
buf BUF1 (N5438, N5431);
or OR2 (N5439, N5424, N2429);
and AND3 (N5440, N5438, N4084, N321);
buf BUF1 (N5441, N5428);
not NOT1 (N5442, N5420);
not NOT1 (N5443, N5437);
nand NAND3 (N5444, N5434, N3079, N1334);
and AND2 (N5445, N5433, N2526);
xor XOR2 (N5446, N5445, N3757);
nand NAND4 (N5447, N5442, N196, N2160, N3002);
nand NAND4 (N5448, N5447, N1867, N1487, N1474);
not NOT1 (N5449, N5443);
buf BUF1 (N5450, N5439);
nand NAND3 (N5451, N5441, N1824, N243);
nor NOR2 (N5452, N5449, N5156);
or OR4 (N5453, N5422, N477, N3065, N2229);
not NOT1 (N5454, N5432);
xor XOR2 (N5455, N5454, N3454);
buf BUF1 (N5456, N5448);
or OR4 (N5457, N5446, N4515, N3927, N3035);
not NOT1 (N5458, N5444);
buf BUF1 (N5459, N5436);
and AND2 (N5460, N5459, N3508);
buf BUF1 (N5461, N5456);
xor XOR2 (N5462, N5450, N1231);
buf BUF1 (N5463, N5452);
nand NAND4 (N5464, N5451, N4560, N5094, N1427);
nand NAND3 (N5465, N5460, N2038, N887);
buf BUF1 (N5466, N5458);
nor NOR2 (N5467, N5465, N2803);
and AND4 (N5468, N5462, N2168, N2783, N3066);
and AND3 (N5469, N5468, N4505, N3867);
nand NAND2 (N5470, N5453, N2164);
nor NOR2 (N5471, N5464, N1484);
not NOT1 (N5472, N5469);
and AND2 (N5473, N5461, N5229);
nand NAND2 (N5474, N5467, N4304);
nand NAND4 (N5475, N5472, N3548, N2345, N707);
nand NAND4 (N5476, N5470, N597, N2427, N3366);
and AND4 (N5477, N5455, N3231, N2057, N2176);
nand NAND2 (N5478, N5457, N3847);
buf BUF1 (N5479, N5463);
buf BUF1 (N5480, N5479);
nand NAND3 (N5481, N5474, N43, N3119);
buf BUF1 (N5482, N5440);
or OR4 (N5483, N5477, N2619, N1201, N1777);
nand NAND3 (N5484, N5480, N2950, N1870);
nor NOR4 (N5485, N5478, N3071, N4139, N3180);
nor NOR2 (N5486, N5466, N742);
nor NOR4 (N5487, N5481, N4837, N4032, N4729);
not NOT1 (N5488, N5484);
nor NOR2 (N5489, N5487, N3105);
buf BUF1 (N5490, N5489);
not NOT1 (N5491, N5475);
not NOT1 (N5492, N5483);
and AND3 (N5493, N5471, N378, N4553);
or OR2 (N5494, N5490, N624);
or OR2 (N5495, N5473, N2840);
xor XOR2 (N5496, N5485, N3374);
buf BUF1 (N5497, N5488);
nand NAND2 (N5498, N5496, N5467);
nand NAND3 (N5499, N5476, N1613, N4504);
nand NAND4 (N5500, N5486, N4659, N3238, N3725);
nor NOR4 (N5501, N5497, N1153, N955, N4044);
buf BUF1 (N5502, N5495);
buf BUF1 (N5503, N5494);
and AND3 (N5504, N5492, N210, N3213);
not NOT1 (N5505, N5503);
buf BUF1 (N5506, N5501);
buf BUF1 (N5507, N5482);
or OR2 (N5508, N5504, N5418);
nor NOR2 (N5509, N5491, N5020);
or OR4 (N5510, N5498, N1951, N5002, N5423);
nand NAND3 (N5511, N5500, N1080, N4242);
not NOT1 (N5512, N5508);
not NOT1 (N5513, N5499);
xor XOR2 (N5514, N5510, N1397);
nand NAND3 (N5515, N5493, N44, N2943);
nand NAND4 (N5516, N5511, N1157, N3062, N4154);
nor NOR3 (N5517, N5509, N657, N4740);
not NOT1 (N5518, N5514);
xor XOR2 (N5519, N5507, N3650);
nand NAND4 (N5520, N5506, N349, N1286, N2975);
buf BUF1 (N5521, N5512);
and AND3 (N5522, N5502, N4, N3668);
nor NOR2 (N5523, N5517, N3908);
or OR2 (N5524, N5522, N2534);
nor NOR4 (N5525, N5519, N4365, N5334, N671);
nor NOR4 (N5526, N5518, N410, N4451, N42);
not NOT1 (N5527, N5513);
buf BUF1 (N5528, N5505);
or OR2 (N5529, N5524, N3600);
not NOT1 (N5530, N5529);
buf BUF1 (N5531, N5527);
and AND2 (N5532, N5526, N400);
or OR3 (N5533, N5531, N2718, N1835);
xor XOR2 (N5534, N5521, N4146);
nor NOR3 (N5535, N5533, N4675, N3280);
not NOT1 (N5536, N5523);
not NOT1 (N5537, N5515);
nand NAND3 (N5538, N5532, N2477, N4277);
and AND2 (N5539, N5538, N3054);
nor NOR3 (N5540, N5525, N3397, N1808);
nand NAND4 (N5541, N5537, N587, N2615, N142);
or OR4 (N5542, N5528, N481, N1734, N572);
not NOT1 (N5543, N5534);
or OR4 (N5544, N5535, N839, N4539, N4049);
or OR3 (N5545, N5516, N3089, N1995);
nor NOR4 (N5546, N5543, N3701, N2235, N3797);
nand NAND3 (N5547, N5530, N3303, N4870);
or OR3 (N5548, N5536, N1224, N1828);
buf BUF1 (N5549, N5520);
and AND4 (N5550, N5539, N2654, N2881, N23);
buf BUF1 (N5551, N5545);
xor XOR2 (N5552, N5541, N5097);
not NOT1 (N5553, N5544);
nor NOR2 (N5554, N5540, N5051);
and AND4 (N5555, N5553, N4970, N412, N4848);
or OR3 (N5556, N5555, N4166, N3364);
xor XOR2 (N5557, N5556, N3904);
buf BUF1 (N5558, N5552);
not NOT1 (N5559, N5550);
and AND2 (N5560, N5542, N87);
buf BUF1 (N5561, N5558);
or OR2 (N5562, N5551, N1533);
xor XOR2 (N5563, N5546, N1481);
and AND4 (N5564, N5554, N1467, N4006, N1365);
or OR3 (N5565, N5562, N3279, N3360);
or OR4 (N5566, N5557, N2119, N716, N3530);
not NOT1 (N5567, N5559);
and AND3 (N5568, N5563, N118, N3276);
nor NOR2 (N5569, N5565, N847);
nor NOR2 (N5570, N5569, N4196);
xor XOR2 (N5571, N5568, N3003);
not NOT1 (N5572, N5561);
or OR4 (N5573, N5572, N2399, N5278, N1115);
not NOT1 (N5574, N5549);
or OR4 (N5575, N5571, N1616, N1840, N5156);
buf BUF1 (N5576, N5547);
nand NAND4 (N5577, N5567, N3206, N4171, N4098);
xor XOR2 (N5578, N5566, N5128);
xor XOR2 (N5579, N5576, N619);
and AND3 (N5580, N5573, N4218, N3594);
buf BUF1 (N5581, N5548);
xor XOR2 (N5582, N5581, N1181);
or OR2 (N5583, N5577, N1363);
nand NAND3 (N5584, N5570, N1125, N2040);
nand NAND2 (N5585, N5560, N3650);
nor NOR2 (N5586, N5584, N3399);
not NOT1 (N5587, N5574);
not NOT1 (N5588, N5587);
buf BUF1 (N5589, N5579);
or OR3 (N5590, N5588, N2682, N3600);
not NOT1 (N5591, N5578);
not NOT1 (N5592, N5583);
xor XOR2 (N5593, N5590, N1754);
buf BUF1 (N5594, N5593);
nand NAND4 (N5595, N5591, N2479, N1613, N1650);
xor XOR2 (N5596, N5595, N491);
nor NOR2 (N5597, N5582, N5275);
xor XOR2 (N5598, N5597, N3562);
or OR2 (N5599, N5580, N2687);
or OR3 (N5600, N5575, N3520, N1187);
and AND3 (N5601, N5586, N120, N4384);
and AND4 (N5602, N5592, N5167, N1473, N3056);
nand NAND4 (N5603, N5564, N3003, N2624, N2227);
or OR3 (N5604, N5594, N1902, N108);
or OR4 (N5605, N5589, N244, N312, N4887);
not NOT1 (N5606, N5600);
not NOT1 (N5607, N5596);
xor XOR2 (N5608, N5605, N524);
buf BUF1 (N5609, N5604);
nand NAND2 (N5610, N5607, N3391);
nor NOR4 (N5611, N5598, N3212, N3120, N1541);
nand NAND3 (N5612, N5611, N2691, N2192);
xor XOR2 (N5613, N5610, N4217);
not NOT1 (N5614, N5601);
and AND2 (N5615, N5599, N4963);
xor XOR2 (N5616, N5614, N1677);
buf BUF1 (N5617, N5603);
or OR4 (N5618, N5606, N3866, N1521, N748);
buf BUF1 (N5619, N5585);
not NOT1 (N5620, N5615);
or OR3 (N5621, N5618, N1452, N2398);
xor XOR2 (N5622, N5608, N3422);
and AND2 (N5623, N5620, N3087);
buf BUF1 (N5624, N5623);
nand NAND4 (N5625, N5622, N2880, N5108, N311);
or OR2 (N5626, N5621, N3244);
nand NAND4 (N5627, N5616, N4812, N385, N262);
nor NOR3 (N5628, N5617, N4853, N4821);
xor XOR2 (N5629, N5628, N2560);
or OR3 (N5630, N5625, N187, N602);
nand NAND2 (N5631, N5624, N5525);
buf BUF1 (N5632, N5602);
xor XOR2 (N5633, N5629, N97);
or OR4 (N5634, N5633, N3177, N3280, N776);
or OR3 (N5635, N5630, N2946, N2357);
not NOT1 (N5636, N5627);
and AND4 (N5637, N5619, N3728, N1498, N453);
and AND3 (N5638, N5609, N4930, N3970);
buf BUF1 (N5639, N5635);
buf BUF1 (N5640, N5639);
xor XOR2 (N5641, N5640, N3106);
buf BUF1 (N5642, N5612);
nor NOR2 (N5643, N5631, N3532);
nand NAND3 (N5644, N5637, N1993, N4322);
or OR3 (N5645, N5634, N4525, N4160);
xor XOR2 (N5646, N5644, N942);
buf BUF1 (N5647, N5642);
buf BUF1 (N5648, N5638);
not NOT1 (N5649, N5632);
nand NAND4 (N5650, N5646, N2423, N1072, N5376);
or OR2 (N5651, N5649, N3378);
not NOT1 (N5652, N5626);
nand NAND4 (N5653, N5648, N5297, N352, N4912);
not NOT1 (N5654, N5645);
xor XOR2 (N5655, N5653, N2207);
nand NAND4 (N5656, N5647, N1963, N4589, N1293);
buf BUF1 (N5657, N5641);
and AND3 (N5658, N5643, N3262, N2955);
nor NOR3 (N5659, N5655, N1790, N4908);
xor XOR2 (N5660, N5652, N1655);
buf BUF1 (N5661, N5636);
and AND3 (N5662, N5661, N4447, N3024);
not NOT1 (N5663, N5658);
xor XOR2 (N5664, N5657, N3646);
or OR3 (N5665, N5651, N3078, N3006);
buf BUF1 (N5666, N5654);
xor XOR2 (N5667, N5656, N3647);
buf BUF1 (N5668, N5659);
nand NAND4 (N5669, N5666, N2376, N585, N1161);
buf BUF1 (N5670, N5668);
and AND4 (N5671, N5663, N2092, N2908, N174);
or OR4 (N5672, N5670, N719, N2158, N2727);
nor NOR2 (N5673, N5613, N5489);
nand NAND4 (N5674, N5671, N2394, N3667, N3762);
nor NOR3 (N5675, N5674, N4039, N1609);
nor NOR3 (N5676, N5675, N2246, N3145);
buf BUF1 (N5677, N5650);
xor XOR2 (N5678, N5677, N1407);
nand NAND3 (N5679, N5664, N5539, N1825);
not NOT1 (N5680, N5665);
not NOT1 (N5681, N5676);
or OR2 (N5682, N5667, N163);
and AND3 (N5683, N5660, N4724, N1672);
nor NOR3 (N5684, N5680, N5504, N1171);
and AND4 (N5685, N5683, N3424, N2519, N3921);
nand NAND4 (N5686, N5669, N1977, N1182, N2733);
not NOT1 (N5687, N5662);
buf BUF1 (N5688, N5682);
nand NAND2 (N5689, N5681, N316);
buf BUF1 (N5690, N5684);
nand NAND2 (N5691, N5688, N1769);
not NOT1 (N5692, N5690);
not NOT1 (N5693, N5691);
nor NOR3 (N5694, N5685, N1510, N820);
and AND3 (N5695, N5692, N3631, N3714);
and AND2 (N5696, N5686, N2431);
buf BUF1 (N5697, N5696);
or OR2 (N5698, N5695, N40);
buf BUF1 (N5699, N5693);
not NOT1 (N5700, N5697);
nand NAND3 (N5701, N5700, N5482, N2789);
nand NAND2 (N5702, N5672, N213);
nand NAND4 (N5703, N5701, N219, N495, N906);
or OR2 (N5704, N5703, N1877);
nand NAND3 (N5705, N5698, N708, N930);
nor NOR4 (N5706, N5687, N5244, N5655, N3402);
or OR3 (N5707, N5705, N882, N3345);
buf BUF1 (N5708, N5678);
buf BUF1 (N5709, N5694);
or OR2 (N5710, N5679, N3356);
and AND4 (N5711, N5708, N812, N3869, N2739);
or OR2 (N5712, N5704, N2334);
not NOT1 (N5713, N5709);
nor NOR2 (N5714, N5713, N1742);
xor XOR2 (N5715, N5689, N928);
and AND3 (N5716, N5706, N2324, N3663);
buf BUF1 (N5717, N5711);
not NOT1 (N5718, N5673);
xor XOR2 (N5719, N5717, N4156);
buf BUF1 (N5720, N5715);
buf BUF1 (N5721, N5712);
not NOT1 (N5722, N5721);
nand NAND2 (N5723, N5719, N1418);
not NOT1 (N5724, N5722);
nand NAND4 (N5725, N5716, N2426, N3925, N537);
buf BUF1 (N5726, N5710);
and AND4 (N5727, N5726, N3679, N1730, N3295);
nand NAND4 (N5728, N5724, N2869, N2981, N5137);
or OR4 (N5729, N5707, N1659, N1961, N724);
nor NOR3 (N5730, N5728, N4876, N3578);
or OR2 (N5731, N5725, N3325);
or OR2 (N5732, N5727, N214);
buf BUF1 (N5733, N5729);
nand NAND3 (N5734, N5699, N359, N3957);
and AND2 (N5735, N5720, N3473);
xor XOR2 (N5736, N5734, N4042);
xor XOR2 (N5737, N5730, N4719);
xor XOR2 (N5738, N5723, N3763);
and AND3 (N5739, N5718, N5579, N2294);
or OR2 (N5740, N5702, N1516);
nor NOR3 (N5741, N5731, N5635, N3838);
nor NOR2 (N5742, N5732, N2568);
buf BUF1 (N5743, N5738);
and AND2 (N5744, N5735, N850);
or OR4 (N5745, N5744, N1543, N129, N2578);
xor XOR2 (N5746, N5740, N2948);
nor NOR4 (N5747, N5739, N2965, N750, N1003);
buf BUF1 (N5748, N5742);
buf BUF1 (N5749, N5748);
xor XOR2 (N5750, N5736, N653);
not NOT1 (N5751, N5745);
nand NAND3 (N5752, N5741, N2547, N2188);
not NOT1 (N5753, N5751);
nor NOR3 (N5754, N5737, N4856, N2997);
nand NAND2 (N5755, N5752, N1496);
buf BUF1 (N5756, N5750);
and AND4 (N5757, N5714, N2580, N2937, N736);
buf BUF1 (N5758, N5746);
not NOT1 (N5759, N5733);
or OR3 (N5760, N5755, N2158, N1653);
buf BUF1 (N5761, N5747);
or OR3 (N5762, N5761, N554, N4470);
and AND4 (N5763, N5757, N1108, N3474, N294);
buf BUF1 (N5764, N5759);
not NOT1 (N5765, N5756);
xor XOR2 (N5766, N5760, N4723);
buf BUF1 (N5767, N5766);
xor XOR2 (N5768, N5767, N917);
and AND4 (N5769, N5763, N1733, N3159, N387);
and AND3 (N5770, N5765, N3879, N37);
not NOT1 (N5771, N5743);
xor XOR2 (N5772, N5770, N4658);
not NOT1 (N5773, N5772);
buf BUF1 (N5774, N5762);
nor NOR3 (N5775, N5764, N1812, N4399);
and AND3 (N5776, N5753, N4911, N2306);
nor NOR3 (N5777, N5771, N3849, N4120);
and AND3 (N5778, N5758, N2742, N612);
buf BUF1 (N5779, N5749);
nand NAND4 (N5780, N5777, N4808, N1737, N5741);
nor NOR4 (N5781, N5775, N5041, N754, N3022);
not NOT1 (N5782, N5776);
or OR2 (N5783, N5778, N2644);
buf BUF1 (N5784, N5769);
nor NOR3 (N5785, N5784, N834, N1693);
or OR4 (N5786, N5785, N135, N3936, N279);
or OR4 (N5787, N5783, N4049, N1791, N2175);
nor NOR2 (N5788, N5787, N4295);
xor XOR2 (N5789, N5782, N2787);
or OR4 (N5790, N5789, N4300, N4227, N1297);
and AND3 (N5791, N5788, N2691, N3714);
xor XOR2 (N5792, N5779, N1221);
or OR3 (N5793, N5791, N1928, N4461);
and AND3 (N5794, N5780, N5793, N4820);
and AND2 (N5795, N4783, N2524);
and AND3 (N5796, N5795, N899, N992);
buf BUF1 (N5797, N5786);
and AND2 (N5798, N5773, N4641);
or OR2 (N5799, N5790, N242);
not NOT1 (N5800, N5799);
nor NOR4 (N5801, N5781, N5528, N178, N206);
nor NOR4 (N5802, N5754, N1442, N5453, N5692);
buf BUF1 (N5803, N5801);
and AND3 (N5804, N5792, N5200, N2172);
nor NOR2 (N5805, N5798, N5712);
xor XOR2 (N5806, N5804, N5324);
and AND2 (N5807, N5768, N3125);
nand NAND2 (N5808, N5796, N4894);
xor XOR2 (N5809, N5806, N2472);
not NOT1 (N5810, N5809);
and AND2 (N5811, N5810, N1597);
nor NOR4 (N5812, N5808, N1115, N2307, N903);
or OR4 (N5813, N5774, N4392, N3210, N4631);
nor NOR2 (N5814, N5794, N2456);
and AND3 (N5815, N5812, N1270, N1436);
xor XOR2 (N5816, N5797, N1848);
nor NOR3 (N5817, N5815, N2983, N3681);
xor XOR2 (N5818, N5816, N2522);
and AND3 (N5819, N5811, N4508, N4219);
xor XOR2 (N5820, N5803, N1736);
or OR4 (N5821, N5819, N872, N1994, N1200);
or OR4 (N5822, N5807, N3302, N1765, N5569);
not NOT1 (N5823, N5817);
buf BUF1 (N5824, N5820);
and AND3 (N5825, N5823, N3278, N1772);
buf BUF1 (N5826, N5821);
buf BUF1 (N5827, N5800);
and AND2 (N5828, N5802, N4831);
and AND4 (N5829, N5822, N3361, N2429, N861);
and AND3 (N5830, N5825, N5291, N2758);
nand NAND4 (N5831, N5813, N5526, N4462, N1052);
xor XOR2 (N5832, N5830, N5147);
nand NAND3 (N5833, N5826, N1087, N2014);
buf BUF1 (N5834, N5827);
buf BUF1 (N5835, N5831);
xor XOR2 (N5836, N5828, N1868);
or OR4 (N5837, N5836, N87, N4378, N5524);
or OR2 (N5838, N5814, N3967);
buf BUF1 (N5839, N5824);
buf BUF1 (N5840, N5818);
nor NOR2 (N5841, N5837, N4572);
nand NAND3 (N5842, N5832, N3466, N5674);
xor XOR2 (N5843, N5841, N1142);
and AND4 (N5844, N5840, N5278, N3712, N5192);
buf BUF1 (N5845, N5843);
xor XOR2 (N5846, N5839, N2906);
xor XOR2 (N5847, N5844, N4618);
xor XOR2 (N5848, N5834, N2930);
nor NOR2 (N5849, N5846, N2657);
and AND2 (N5850, N5842, N560);
or OR3 (N5851, N5835, N4209, N938);
and AND4 (N5852, N5838, N1875, N3904, N3833);
buf BUF1 (N5853, N5849);
or OR2 (N5854, N5829, N951);
nand NAND3 (N5855, N5845, N702, N366);
nand NAND3 (N5856, N5850, N689, N913);
xor XOR2 (N5857, N5853, N281);
nand NAND4 (N5858, N5847, N3123, N2800, N710);
nor NOR3 (N5859, N5848, N326, N3581);
buf BUF1 (N5860, N5856);
buf BUF1 (N5861, N5858);
and AND2 (N5862, N5859, N4984);
or OR2 (N5863, N5857, N271);
and AND2 (N5864, N5854, N2250);
or OR3 (N5865, N5851, N203, N3126);
nand NAND2 (N5866, N5805, N4463);
buf BUF1 (N5867, N5833);
buf BUF1 (N5868, N5852);
buf BUF1 (N5869, N5863);
not NOT1 (N5870, N5860);
nand NAND3 (N5871, N5855, N453, N4590);
and AND4 (N5872, N5870, N4849, N1138, N836);
or OR3 (N5873, N5861, N5457, N5601);
not NOT1 (N5874, N5867);
nand NAND4 (N5875, N5872, N919, N353, N5676);
buf BUF1 (N5876, N5875);
or OR3 (N5877, N5868, N1235, N5579);
xor XOR2 (N5878, N5877, N4195);
nor NOR2 (N5879, N5874, N126);
not NOT1 (N5880, N5862);
nand NAND2 (N5881, N5880, N4934);
or OR2 (N5882, N5869, N1309);
nand NAND4 (N5883, N5882, N1098, N888, N684);
nand NAND2 (N5884, N5883, N4972);
buf BUF1 (N5885, N5865);
not NOT1 (N5886, N5873);
nor NOR2 (N5887, N5878, N683);
nor NOR2 (N5888, N5866, N839);
nand NAND4 (N5889, N5884, N5037, N2420, N5300);
and AND4 (N5890, N5871, N901, N5068, N4992);
nand NAND4 (N5891, N5886, N3700, N842, N2700);
or OR4 (N5892, N5889, N4848, N5270, N4935);
xor XOR2 (N5893, N5887, N2457);
xor XOR2 (N5894, N5885, N2327);
xor XOR2 (N5895, N5891, N2212);
xor XOR2 (N5896, N5888, N5888);
buf BUF1 (N5897, N5892);
nor NOR3 (N5898, N5864, N4399, N5896);
nand NAND2 (N5899, N3463, N3618);
not NOT1 (N5900, N5898);
not NOT1 (N5901, N5893);
buf BUF1 (N5902, N5900);
buf BUF1 (N5903, N5901);
nor NOR4 (N5904, N5897, N4860, N1802, N241);
xor XOR2 (N5905, N5894, N374);
not NOT1 (N5906, N5876);
buf BUF1 (N5907, N5906);
and AND4 (N5908, N5907, N4614, N1723, N3552);
buf BUF1 (N5909, N5881);
buf BUF1 (N5910, N5905);
or OR4 (N5911, N5879, N5157, N1666, N1687);
not NOT1 (N5912, N5899);
xor XOR2 (N5913, N5911, N3293);
nand NAND3 (N5914, N5903, N1733, N109);
or OR2 (N5915, N5913, N1219);
nand NAND2 (N5916, N5915, N4944);
not NOT1 (N5917, N5914);
and AND4 (N5918, N5890, N4074, N1589, N3189);
buf BUF1 (N5919, N5895);
buf BUF1 (N5920, N5916);
or OR2 (N5921, N5904, N1332);
or OR3 (N5922, N5920, N3396, N1781);
or OR2 (N5923, N5918, N4079);
not NOT1 (N5924, N5921);
nand NAND3 (N5925, N5919, N5097, N2832);
and AND2 (N5926, N5925, N5772);
xor XOR2 (N5927, N5924, N5251);
nand NAND3 (N5928, N5927, N2640, N4720);
xor XOR2 (N5929, N5922, N5874);
or OR3 (N5930, N5928, N262, N5558);
nor NOR3 (N5931, N5909, N4366, N3751);
buf BUF1 (N5932, N5902);
nor NOR4 (N5933, N5908, N4417, N5090, N4660);
xor XOR2 (N5934, N5931, N782);
nand NAND3 (N5935, N5934, N185, N3022);
and AND3 (N5936, N5930, N3527, N1141);
nand NAND4 (N5937, N5935, N451, N5509, N4757);
xor XOR2 (N5938, N5936, N4313);
nor NOR4 (N5939, N5929, N4945, N4748, N5024);
nand NAND2 (N5940, N5926, N2228);
nor NOR4 (N5941, N5932, N3880, N2589, N5450);
xor XOR2 (N5942, N5939, N71);
nor NOR4 (N5943, N5938, N2428, N4840, N4721);
buf BUF1 (N5944, N5941);
and AND4 (N5945, N5943, N3842, N789, N5565);
xor XOR2 (N5946, N5940, N1370);
buf BUF1 (N5947, N5912);
nand NAND3 (N5948, N5910, N2145, N1441);
xor XOR2 (N5949, N5933, N1314);
not NOT1 (N5950, N5949);
not NOT1 (N5951, N5950);
nor NOR2 (N5952, N5946, N1243);
or OR3 (N5953, N5948, N1341, N4585);
and AND4 (N5954, N5953, N1172, N1795, N5718);
and AND4 (N5955, N5947, N2958, N3641, N5322);
not NOT1 (N5956, N5917);
nand NAND3 (N5957, N5942, N1646, N1603);
nand NAND4 (N5958, N5956, N332, N560, N2234);
not NOT1 (N5959, N5954);
xor XOR2 (N5960, N5944, N5942);
buf BUF1 (N5961, N5937);
xor XOR2 (N5962, N5945, N4389);
nand NAND2 (N5963, N5957, N5325);
nor NOR4 (N5964, N5955, N3944, N788, N5736);
nand NAND4 (N5965, N5923, N5432, N3269, N5213);
not NOT1 (N5966, N5965);
and AND3 (N5967, N5964, N5479, N1998);
buf BUF1 (N5968, N5962);
nor NOR2 (N5969, N5966, N91);
xor XOR2 (N5970, N5959, N1963);
or OR3 (N5971, N5967, N4244, N657);
or OR3 (N5972, N5963, N86, N4025);
nor NOR2 (N5973, N5958, N4934);
buf BUF1 (N5974, N5952);
and AND2 (N5975, N5971, N5118);
xor XOR2 (N5976, N5968, N791);
not NOT1 (N5977, N5972);
nand NAND2 (N5978, N5961, N1181);
not NOT1 (N5979, N5960);
buf BUF1 (N5980, N5951);
nor NOR3 (N5981, N5973, N581, N5418);
buf BUF1 (N5982, N5977);
nor NOR4 (N5983, N5974, N1502, N1795, N5830);
xor XOR2 (N5984, N5980, N5276);
not NOT1 (N5985, N5975);
nor NOR2 (N5986, N5982, N3656);
or OR4 (N5987, N5978, N5648, N4120, N3819);
and AND4 (N5988, N5976, N972, N3420, N228);
xor XOR2 (N5989, N5969, N403);
nor NOR4 (N5990, N5989, N1047, N3837, N3034);
and AND4 (N5991, N5990, N4585, N450, N5446);
not NOT1 (N5992, N5988);
or OR3 (N5993, N5983, N2274, N4541);
buf BUF1 (N5994, N5981);
nor NOR2 (N5995, N5994, N2594);
and AND3 (N5996, N5991, N5666, N4483);
nor NOR3 (N5997, N5970, N4045, N2485);
xor XOR2 (N5998, N5979, N4501);
nand NAND2 (N5999, N5984, N1364);
xor XOR2 (N6000, N5987, N4866);
nor NOR2 (N6001, N5999, N2414);
xor XOR2 (N6002, N5985, N3158);
buf BUF1 (N6003, N6001);
nand NAND3 (N6004, N5998, N3223, N3933);
or OR2 (N6005, N6004, N3067);
buf BUF1 (N6006, N6002);
and AND4 (N6007, N5996, N1586, N266, N945);
xor XOR2 (N6008, N5992, N933);
buf BUF1 (N6009, N5995);
or OR2 (N6010, N6007, N1278);
xor XOR2 (N6011, N5986, N5951);
xor XOR2 (N6012, N6011, N5646);
buf BUF1 (N6013, N6008);
or OR4 (N6014, N6000, N1234, N3714, N1791);
buf BUF1 (N6015, N6006);
nand NAND3 (N6016, N6003, N2461, N968);
nand NAND4 (N6017, N6005, N4435, N1900, N2771);
buf BUF1 (N6018, N6013);
xor XOR2 (N6019, N6015, N2242);
or OR2 (N6020, N6010, N1253);
xor XOR2 (N6021, N5997, N2436);
buf BUF1 (N6022, N6021);
or OR4 (N6023, N6012, N4049, N1140, N4527);
xor XOR2 (N6024, N5993, N2369);
buf BUF1 (N6025, N6017);
buf BUF1 (N6026, N6022);
nor NOR2 (N6027, N6018, N3392);
nand NAND2 (N6028, N6024, N3209);
xor XOR2 (N6029, N6020, N5077);
not NOT1 (N6030, N6016);
buf BUF1 (N6031, N6029);
nor NOR2 (N6032, N6031, N5460);
not NOT1 (N6033, N6009);
buf BUF1 (N6034, N6028);
or OR4 (N6035, N6032, N5517, N1224, N5405);
xor XOR2 (N6036, N6027, N3853);
not NOT1 (N6037, N6026);
not NOT1 (N6038, N6030);
nand NAND3 (N6039, N6038, N2205, N3483);
nand NAND2 (N6040, N6034, N3914);
nor NOR4 (N6041, N6036, N2767, N285, N3475);
or OR2 (N6042, N6033, N5805);
nand NAND2 (N6043, N6040, N2601);
xor XOR2 (N6044, N6035, N501);
not NOT1 (N6045, N6025);
and AND3 (N6046, N6041, N3315, N2758);
nor NOR3 (N6047, N6039, N692, N5513);
nor NOR2 (N6048, N6047, N3659);
and AND3 (N6049, N6014, N2323, N3169);
buf BUF1 (N6050, N6037);
buf BUF1 (N6051, N6023);
buf BUF1 (N6052, N6051);
and AND3 (N6053, N6045, N3660, N4343);
xor XOR2 (N6054, N6052, N4175);
or OR4 (N6055, N6043, N551, N2965, N56);
nand NAND2 (N6056, N6042, N2854);
and AND3 (N6057, N6019, N1145, N4591);
xor XOR2 (N6058, N6049, N5521);
not NOT1 (N6059, N6055);
buf BUF1 (N6060, N6054);
not NOT1 (N6061, N6046);
or OR2 (N6062, N6056, N2658);
xor XOR2 (N6063, N6048, N2543);
nand NAND3 (N6064, N6053, N4117, N1366);
or OR3 (N6065, N6061, N5272, N5485);
nor NOR3 (N6066, N6060, N1506, N2279);
and AND4 (N6067, N6050, N4455, N2223, N4428);
or OR2 (N6068, N6063, N2478);
nand NAND2 (N6069, N6057, N1483);
nor NOR3 (N6070, N6062, N770, N2734);
or OR3 (N6071, N6068, N3492, N4619);
buf BUF1 (N6072, N6069);
xor XOR2 (N6073, N6072, N1840);
or OR2 (N6074, N6059, N5146);
or OR3 (N6075, N6071, N5168, N199);
not NOT1 (N6076, N6075);
nand NAND3 (N6077, N6074, N1055, N2965);
or OR4 (N6078, N6064, N1266, N2433, N2713);
nand NAND3 (N6079, N6058, N4826, N5219);
nand NAND2 (N6080, N6066, N4615);
nor NOR3 (N6081, N6080, N1737, N3767);
xor XOR2 (N6082, N6070, N220);
or OR3 (N6083, N6078, N1910, N1988);
buf BUF1 (N6084, N6077);
and AND3 (N6085, N6083, N3758, N2567);
buf BUF1 (N6086, N6073);
xor XOR2 (N6087, N6082, N1035);
buf BUF1 (N6088, N6081);
and AND2 (N6089, N6087, N5317);
and AND4 (N6090, N6076, N5104, N1096, N1406);
not NOT1 (N6091, N6090);
nor NOR2 (N6092, N6089, N950);
nand NAND4 (N6093, N6067, N1475, N4954, N204);
xor XOR2 (N6094, N6084, N2972);
or OR3 (N6095, N6091, N1193, N2685);
xor XOR2 (N6096, N6086, N5549);
and AND4 (N6097, N6092, N2671, N5981, N5213);
xor XOR2 (N6098, N6044, N3705);
not NOT1 (N6099, N6065);
or OR3 (N6100, N6088, N3951, N5389);
or OR4 (N6101, N6093, N2281, N1767, N4360);
nor NOR3 (N6102, N6101, N4129, N4905);
not NOT1 (N6103, N6098);
nor NOR2 (N6104, N6095, N3153);
or OR3 (N6105, N6097, N74, N5806);
or OR3 (N6106, N6100, N4206, N3910);
or OR3 (N6107, N6094, N3427, N1537);
nand NAND2 (N6108, N6105, N4337);
not NOT1 (N6109, N6096);
nor NOR3 (N6110, N6085, N1913, N1429);
xor XOR2 (N6111, N6108, N4474);
nor NOR2 (N6112, N6109, N4213);
not NOT1 (N6113, N6102);
nand NAND3 (N6114, N6111, N2386, N1485);
or OR4 (N6115, N6114, N2924, N1774, N3243);
nor NOR2 (N6116, N6115, N2956);
xor XOR2 (N6117, N6107, N3484);
and AND3 (N6118, N6104, N3749, N2766);
buf BUF1 (N6119, N6113);
nor NOR3 (N6120, N6116, N2024, N3661);
and AND4 (N6121, N6119, N2080, N681, N3965);
and AND4 (N6122, N6117, N1964, N681, N4558);
and AND4 (N6123, N6110, N3232, N1954, N3973);
nand NAND4 (N6124, N6103, N126, N4695, N3605);
buf BUF1 (N6125, N6120);
xor XOR2 (N6126, N6121, N2804);
buf BUF1 (N6127, N6118);
not NOT1 (N6128, N6127);
not NOT1 (N6129, N6106);
nor NOR3 (N6130, N6124, N470, N5453);
nor NOR4 (N6131, N6099, N4286, N1748, N1154);
not NOT1 (N6132, N6079);
nor NOR2 (N6133, N6123, N5116);
not NOT1 (N6134, N6129);
nor NOR3 (N6135, N6128, N3021, N47);
and AND4 (N6136, N6131, N4594, N1009, N2592);
nor NOR4 (N6137, N6112, N930, N5228, N395);
or OR3 (N6138, N6125, N439, N2035);
nand NAND4 (N6139, N6126, N2489, N2126, N925);
and AND4 (N6140, N6138, N4742, N2298, N4388);
nand NAND4 (N6141, N6135, N4867, N2851, N3644);
and AND2 (N6142, N6137, N3913);
nor NOR2 (N6143, N6139, N2516);
buf BUF1 (N6144, N6133);
not NOT1 (N6145, N6122);
or OR2 (N6146, N6141, N1846);
and AND4 (N6147, N6142, N2337, N3467, N2452);
xor XOR2 (N6148, N6130, N4411);
not NOT1 (N6149, N6146);
nand NAND3 (N6150, N6144, N812, N5773);
nand NAND2 (N6151, N6140, N5648);
nor NOR2 (N6152, N6150, N4913);
buf BUF1 (N6153, N6149);
nor NOR3 (N6154, N6148, N5679, N1808);
or OR2 (N6155, N6151, N3489);
nor NOR4 (N6156, N6134, N4007, N1159, N2650);
buf BUF1 (N6157, N6132);
nor NOR4 (N6158, N6153, N1839, N2945, N3057);
not NOT1 (N6159, N6136);
xor XOR2 (N6160, N6147, N1627);
and AND2 (N6161, N6159, N6);
nand NAND2 (N6162, N6156, N3615);
not NOT1 (N6163, N6157);
nor NOR4 (N6164, N6163, N4712, N5125, N4972);
and AND2 (N6165, N6161, N217);
and AND4 (N6166, N6143, N3076, N4271, N4974);
xor XOR2 (N6167, N6154, N1678);
or OR3 (N6168, N6162, N2121, N1003);
not NOT1 (N6169, N6168);
or OR2 (N6170, N6164, N1965);
xor XOR2 (N6171, N6170, N1415);
nor NOR2 (N6172, N6155, N1979);
buf BUF1 (N6173, N6171);
nor NOR3 (N6174, N6166, N3999, N4812);
nand NAND3 (N6175, N6174, N2749, N405);
nand NAND4 (N6176, N6175, N5526, N2832, N303);
xor XOR2 (N6177, N6165, N1324);
not NOT1 (N6178, N6172);
or OR4 (N6179, N6167, N4783, N3744, N1536);
and AND3 (N6180, N6145, N2673, N1367);
not NOT1 (N6181, N6176);
nor NOR3 (N6182, N6173, N6076, N3781);
buf BUF1 (N6183, N6177);
not NOT1 (N6184, N6180);
nand NAND2 (N6185, N6160, N967);
or OR4 (N6186, N6184, N5607, N39, N4385);
buf BUF1 (N6187, N6186);
or OR4 (N6188, N6158, N2382, N4604, N4600);
and AND4 (N6189, N6182, N6176, N2032, N5223);
nor NOR3 (N6190, N6187, N3448, N1270);
nor NOR3 (N6191, N6179, N332, N1074);
or OR4 (N6192, N6185, N5852, N429, N1185);
nor NOR2 (N6193, N6152, N2361);
and AND3 (N6194, N6178, N428, N2204);
nand NAND2 (N6195, N6192, N5389);
not NOT1 (N6196, N6193);
nor NOR3 (N6197, N6194, N2219, N4190);
not NOT1 (N6198, N6188);
xor XOR2 (N6199, N6195, N5579);
nand NAND3 (N6200, N6181, N5657, N5649);
or OR2 (N6201, N6183, N2272);
not NOT1 (N6202, N6190);
xor XOR2 (N6203, N6197, N4410);
or OR3 (N6204, N6189, N3295, N4770);
not NOT1 (N6205, N6198);
xor XOR2 (N6206, N6205, N1289);
and AND4 (N6207, N6202, N1768, N901, N5764);
xor XOR2 (N6208, N6204, N3089);
not NOT1 (N6209, N6169);
buf BUF1 (N6210, N6203);
nor NOR3 (N6211, N6207, N500, N6067);
nor NOR2 (N6212, N6210, N2750);
xor XOR2 (N6213, N6200, N4526);
or OR4 (N6214, N6213, N4837, N5461, N3352);
nand NAND4 (N6215, N6214, N5416, N2980, N489);
buf BUF1 (N6216, N6199);
buf BUF1 (N6217, N6191);
and AND4 (N6218, N6215, N1359, N5483, N1864);
not NOT1 (N6219, N6218);
and AND3 (N6220, N6216, N2482, N5637);
nor NOR2 (N6221, N6217, N347);
or OR4 (N6222, N6206, N3806, N2830, N2347);
nor NOR2 (N6223, N6201, N971);
buf BUF1 (N6224, N6212);
and AND4 (N6225, N6220, N1523, N2719, N3866);
or OR2 (N6226, N6223, N3469);
nor NOR2 (N6227, N6225, N3049);
nor NOR3 (N6228, N6221, N4260, N5909);
or OR2 (N6229, N6196, N5879);
nand NAND3 (N6230, N6208, N5583, N5142);
or OR4 (N6231, N6209, N3219, N2592, N5154);
nand NAND2 (N6232, N6219, N1481);
xor XOR2 (N6233, N6224, N4522);
not NOT1 (N6234, N6229);
xor XOR2 (N6235, N6230, N2756);
or OR2 (N6236, N6233, N806);
nand NAND3 (N6237, N6236, N1800, N4187);
and AND3 (N6238, N6228, N182, N5338);
and AND4 (N6239, N6237, N4567, N392, N2741);
or OR2 (N6240, N6226, N5617);
buf BUF1 (N6241, N6238);
and AND3 (N6242, N6227, N904, N4118);
xor XOR2 (N6243, N6222, N2489);
nor NOR2 (N6244, N6235, N3283);
buf BUF1 (N6245, N6241);
buf BUF1 (N6246, N6244);
not NOT1 (N6247, N6246);
nor NOR3 (N6248, N6247, N5908, N1006);
xor XOR2 (N6249, N6242, N2831);
and AND2 (N6250, N6231, N4914);
or OR4 (N6251, N6248, N3095, N3607, N3570);
xor XOR2 (N6252, N6251, N4894);
or OR3 (N6253, N6232, N2935, N2681);
or OR3 (N6254, N6211, N3370, N4292);
buf BUF1 (N6255, N6234);
nand NAND3 (N6256, N6243, N2188, N1122);
xor XOR2 (N6257, N6254, N4949);
nand NAND3 (N6258, N6239, N1623, N6192);
buf BUF1 (N6259, N6253);
xor XOR2 (N6260, N6250, N3504);
and AND4 (N6261, N6257, N1488, N5865, N5723);
nand NAND2 (N6262, N6261, N6159);
nand NAND4 (N6263, N6260, N1327, N5304, N2707);
nor NOR2 (N6264, N6263, N2913);
buf BUF1 (N6265, N6255);
and AND4 (N6266, N6249, N3971, N3204, N1066);
not NOT1 (N6267, N6259);
nand NAND3 (N6268, N6264, N5510, N5087);
not NOT1 (N6269, N6256);
or OR4 (N6270, N6266, N4896, N67, N2277);
or OR2 (N6271, N6270, N5942);
nand NAND4 (N6272, N6271, N428, N5514, N86);
buf BUF1 (N6273, N6245);
or OR2 (N6274, N6272, N5094);
and AND4 (N6275, N6273, N5822, N1251, N2097);
not NOT1 (N6276, N6265);
nor NOR3 (N6277, N6258, N1172, N5543);
not NOT1 (N6278, N6276);
buf BUF1 (N6279, N6262);
nor NOR2 (N6280, N6278, N2268);
buf BUF1 (N6281, N6277);
nand NAND2 (N6282, N6267, N3072);
nor NOR3 (N6283, N6240, N1100, N4898);
or OR3 (N6284, N6274, N3594, N1710);
not NOT1 (N6285, N6283);
buf BUF1 (N6286, N6279);
nand NAND4 (N6287, N6286, N6161, N3842, N2346);
not NOT1 (N6288, N6287);
buf BUF1 (N6289, N6268);
nand NAND3 (N6290, N6275, N5721, N416);
not NOT1 (N6291, N6288);
and AND3 (N6292, N6291, N3505, N3276);
and AND3 (N6293, N6289, N3321, N5956);
and AND3 (N6294, N6282, N638, N2052);
nand NAND4 (N6295, N6280, N1751, N1380, N4455);
and AND4 (N6296, N6281, N5048, N4936, N2261);
xor XOR2 (N6297, N6290, N2119);
nor NOR4 (N6298, N6285, N3230, N3157, N3453);
not NOT1 (N6299, N6252);
xor XOR2 (N6300, N6284, N1769);
or OR3 (N6301, N6297, N5557, N1598);
nand NAND4 (N6302, N6296, N1129, N1048, N6121);
nor NOR4 (N6303, N6294, N5104, N498, N6166);
nand NAND4 (N6304, N6292, N4990, N4554, N228);
and AND3 (N6305, N6302, N4041, N452);
buf BUF1 (N6306, N6269);
buf BUF1 (N6307, N6304);
nand NAND4 (N6308, N6301, N4362, N2078, N2247);
buf BUF1 (N6309, N6298);
or OR2 (N6310, N6306, N1033);
not NOT1 (N6311, N6305);
xor XOR2 (N6312, N6311, N5659);
buf BUF1 (N6313, N6295);
nand NAND2 (N6314, N6300, N6216);
nor NOR3 (N6315, N6314, N3927, N3925);
nor NOR4 (N6316, N6313, N2120, N5081, N4616);
not NOT1 (N6317, N6308);
buf BUF1 (N6318, N6317);
or OR2 (N6319, N6309, N818);
buf BUF1 (N6320, N6315);
or OR3 (N6321, N6293, N2576, N4854);
or OR2 (N6322, N6318, N3246);
nand NAND3 (N6323, N6319, N5582, N3273);
or OR4 (N6324, N6310, N6260, N114, N3634);
nand NAND3 (N6325, N6323, N2284, N3371);
and AND3 (N6326, N6320, N4552, N1360);
nor NOR2 (N6327, N6322, N4895);
nand NAND4 (N6328, N6303, N5409, N1974, N4788);
not NOT1 (N6329, N6327);
nand NAND3 (N6330, N6326, N1448, N4104);
not NOT1 (N6331, N6324);
nand NAND3 (N6332, N6331, N341, N6116);
not NOT1 (N6333, N6316);
or OR4 (N6334, N6332, N127, N4655, N3943);
nand NAND2 (N6335, N6329, N5586);
not NOT1 (N6336, N6312);
nor NOR3 (N6337, N6336, N6247, N1107);
or OR2 (N6338, N6325, N4944);
xor XOR2 (N6339, N6307, N1783);
nor NOR3 (N6340, N6337, N5198, N122);
buf BUF1 (N6341, N6330);
and AND2 (N6342, N6340, N4848);
xor XOR2 (N6343, N6321, N2258);
or OR4 (N6344, N6343, N4375, N1783, N686);
buf BUF1 (N6345, N6335);
buf BUF1 (N6346, N6342);
xor XOR2 (N6347, N6299, N1143);
and AND3 (N6348, N6345, N1479, N1191);
not NOT1 (N6349, N6328);
xor XOR2 (N6350, N6348, N3613);
nor NOR2 (N6351, N6350, N5361);
nand NAND3 (N6352, N6347, N457, N1588);
xor XOR2 (N6353, N6333, N5648);
and AND4 (N6354, N6349, N3382, N77, N5270);
nand NAND4 (N6355, N6354, N5354, N4269, N2551);
not NOT1 (N6356, N6355);
nand NAND2 (N6357, N6334, N3905);
not NOT1 (N6358, N6344);
or OR2 (N6359, N6356, N3341);
or OR3 (N6360, N6338, N34, N4660);
and AND3 (N6361, N6358, N588, N4588);
not NOT1 (N6362, N6351);
not NOT1 (N6363, N6357);
xor XOR2 (N6364, N6353, N128);
and AND2 (N6365, N6363, N2389);
buf BUF1 (N6366, N6352);
or OR4 (N6367, N6364, N6270, N6046, N1522);
nand NAND4 (N6368, N6360, N5150, N3373, N4380);
not NOT1 (N6369, N6368);
nor NOR3 (N6370, N6367, N4321, N3739);
nor NOR4 (N6371, N6359, N3766, N1573, N1492);
or OR3 (N6372, N6362, N5237, N812);
buf BUF1 (N6373, N6346);
nor NOR2 (N6374, N6341, N452);
nor NOR4 (N6375, N6339, N693, N823, N2674);
nand NAND4 (N6376, N6365, N4145, N5795, N2877);
nand NAND3 (N6377, N6375, N6056, N5698);
buf BUF1 (N6378, N6371);
or OR2 (N6379, N6378, N2385);
nor NOR2 (N6380, N6361, N263);
or OR3 (N6381, N6376, N1183, N5938);
or OR3 (N6382, N6369, N1457, N975);
xor XOR2 (N6383, N6366, N1074);
nor NOR4 (N6384, N6379, N4614, N3848, N5504);
nor NOR4 (N6385, N6373, N3551, N5167, N6068);
nor NOR4 (N6386, N6374, N6252, N6190, N2275);
not NOT1 (N6387, N6386);
buf BUF1 (N6388, N6381);
nand NAND3 (N6389, N6383, N4060, N6097);
nor NOR4 (N6390, N6389, N4347, N5990, N5873);
buf BUF1 (N6391, N6377);
nor NOR3 (N6392, N6387, N1529, N238);
and AND3 (N6393, N6385, N3523, N4318);
xor XOR2 (N6394, N6372, N6150);
or OR4 (N6395, N6392, N6066, N2719, N5288);
nand NAND4 (N6396, N6394, N6017, N4017, N5517);
xor XOR2 (N6397, N6382, N5589);
or OR2 (N6398, N6395, N2437);
buf BUF1 (N6399, N6393);
and AND3 (N6400, N6384, N5165, N457);
and AND2 (N6401, N6396, N2834);
and AND2 (N6402, N6401, N3451);
not NOT1 (N6403, N6397);
buf BUF1 (N6404, N6370);
nand NAND4 (N6405, N6404, N2732, N6172, N3393);
xor XOR2 (N6406, N6399, N3010);
nor NOR2 (N6407, N6398, N2220);
and AND3 (N6408, N6403, N3874, N4444);
xor XOR2 (N6409, N6390, N5217);
buf BUF1 (N6410, N6406);
not NOT1 (N6411, N6400);
xor XOR2 (N6412, N6388, N4266);
nor NOR2 (N6413, N6411, N2050);
not NOT1 (N6414, N6402);
or OR4 (N6415, N6407, N3728, N1314, N5445);
and AND2 (N6416, N6391, N4308);
or OR4 (N6417, N6380, N3052, N1785, N1750);
not NOT1 (N6418, N6409);
buf BUF1 (N6419, N6417);
nor NOR3 (N6420, N6414, N3568, N286);
buf BUF1 (N6421, N6405);
nor NOR3 (N6422, N6410, N981, N433);
and AND4 (N6423, N6420, N4523, N5441, N2736);
not NOT1 (N6424, N6413);
xor XOR2 (N6425, N6422, N2061);
nor NOR3 (N6426, N6416, N12, N545);
nor NOR3 (N6427, N6418, N1871, N384);
and AND4 (N6428, N6427, N2093, N6295, N124);
buf BUF1 (N6429, N6419);
not NOT1 (N6430, N6428);
xor XOR2 (N6431, N6421, N2237);
nor NOR4 (N6432, N6430, N679, N1445, N1012);
not NOT1 (N6433, N6426);
xor XOR2 (N6434, N6432, N1182);
nand NAND2 (N6435, N6425, N2768);
nor NOR4 (N6436, N6435, N5061, N5380, N4164);
nand NAND2 (N6437, N6415, N5304);
not NOT1 (N6438, N6431);
or OR3 (N6439, N6408, N1652, N4684);
nor NOR2 (N6440, N6424, N5726);
not NOT1 (N6441, N6433);
xor XOR2 (N6442, N6436, N4359);
or OR4 (N6443, N6429, N269, N2484, N177);
or OR4 (N6444, N6434, N2119, N3636, N3956);
not NOT1 (N6445, N6438);
or OR2 (N6446, N6441, N1369);
nor NOR3 (N6447, N6446, N242, N3941);
buf BUF1 (N6448, N6443);
xor XOR2 (N6449, N6448, N944);
or OR2 (N6450, N6445, N4404);
and AND2 (N6451, N6412, N6203);
xor XOR2 (N6452, N6437, N4426);
or OR4 (N6453, N6452, N2700, N3429, N575);
nor NOR3 (N6454, N6439, N5568, N5838);
nand NAND4 (N6455, N6453, N6043, N2285, N6120);
buf BUF1 (N6456, N6423);
buf BUF1 (N6457, N6455);
buf BUF1 (N6458, N6456);
or OR2 (N6459, N6457, N6081);
nor NOR2 (N6460, N6450, N6077);
nand NAND4 (N6461, N6451, N5447, N99, N3931);
and AND3 (N6462, N6442, N1291, N6386);
nor NOR3 (N6463, N6460, N5086, N2188);
nor NOR3 (N6464, N6454, N5823, N4615);
not NOT1 (N6465, N6449);
nand NAND3 (N6466, N6461, N4480, N2480);
buf BUF1 (N6467, N6466);
nor NOR4 (N6468, N6459, N3681, N4373, N6060);
buf BUF1 (N6469, N6465);
buf BUF1 (N6470, N6440);
or OR3 (N6471, N6468, N3802, N5951);
nand NAND2 (N6472, N6467, N3225);
not NOT1 (N6473, N6463);
not NOT1 (N6474, N6458);
xor XOR2 (N6475, N6447, N755);
or OR4 (N6476, N6444, N4817, N4626, N4852);
or OR2 (N6477, N6476, N895);
or OR3 (N6478, N6475, N1335, N2600);
and AND3 (N6479, N6472, N5990, N1868);
nand NAND4 (N6480, N6469, N2269, N5382, N3264);
buf BUF1 (N6481, N6462);
xor XOR2 (N6482, N6473, N4785);
and AND2 (N6483, N6477, N2664);
xor XOR2 (N6484, N6471, N4092);
nor NOR2 (N6485, N6483, N6367);
and AND3 (N6486, N6478, N4100, N6440);
and AND3 (N6487, N6482, N4914, N740);
nand NAND4 (N6488, N6480, N4169, N1915, N5348);
and AND4 (N6489, N6484, N2883, N6335, N5320);
and AND2 (N6490, N6489, N2018);
and AND3 (N6491, N6481, N4395, N2112);
nor NOR2 (N6492, N6470, N4617);
and AND3 (N6493, N6479, N2297, N2071);
xor XOR2 (N6494, N6464, N1095);
nor NOR3 (N6495, N6487, N4800, N6029);
and AND2 (N6496, N6493, N98);
and AND3 (N6497, N6495, N2033, N681);
buf BUF1 (N6498, N6490);
not NOT1 (N6499, N6497);
and AND4 (N6500, N6492, N3267, N5819, N1018);
and AND3 (N6501, N6491, N2799, N4236);
xor XOR2 (N6502, N6496, N4445);
nand NAND2 (N6503, N6474, N4213);
nand NAND2 (N6504, N6494, N2690);
nand NAND2 (N6505, N6485, N3215);
buf BUF1 (N6506, N6505);
not NOT1 (N6507, N6498);
or OR4 (N6508, N6501, N2452, N162, N4337);
and AND3 (N6509, N6486, N3205, N1102);
nand NAND3 (N6510, N6503, N3034, N3179);
buf BUF1 (N6511, N6499);
and AND3 (N6512, N6508, N4344, N6444);
not NOT1 (N6513, N6500);
nor NOR3 (N6514, N6513, N6038, N4751);
buf BUF1 (N6515, N6511);
buf BUF1 (N6516, N6504);
xor XOR2 (N6517, N6512, N1375);
nand NAND4 (N6518, N6515, N5176, N6372, N5628);
or OR4 (N6519, N6518, N1284, N2457, N2058);
nor NOR2 (N6520, N6516, N3648);
xor XOR2 (N6521, N6520, N2155);
and AND4 (N6522, N6488, N4142, N2982, N4281);
and AND3 (N6523, N6502, N741, N3996);
xor XOR2 (N6524, N6506, N5589);
and AND4 (N6525, N6523, N2358, N6413, N1853);
buf BUF1 (N6526, N6522);
not NOT1 (N6527, N6521);
or OR3 (N6528, N6514, N683, N1977);
or OR2 (N6529, N6525, N1877);
not NOT1 (N6530, N6519);
or OR2 (N6531, N6530, N2806);
and AND4 (N6532, N6528, N3700, N4694, N6239);
and AND2 (N6533, N6517, N4876);
nand NAND4 (N6534, N6533, N2979, N5514, N3469);
buf BUF1 (N6535, N6532);
buf BUF1 (N6536, N6509);
not NOT1 (N6537, N6534);
and AND2 (N6538, N6524, N4017);
and AND3 (N6539, N6535, N2492, N325);
xor XOR2 (N6540, N6536, N3649);
or OR4 (N6541, N6539, N6161, N1053, N6);
not NOT1 (N6542, N6527);
or OR3 (N6543, N6537, N6493, N5955);
or OR4 (N6544, N6538, N5256, N2114, N1431);
nand NAND2 (N6545, N6543, N3816);
buf BUF1 (N6546, N6507);
buf BUF1 (N6547, N6529);
buf BUF1 (N6548, N6547);
nand NAND3 (N6549, N6544, N331, N658);
xor XOR2 (N6550, N6526, N3356);
or OR2 (N6551, N6540, N3344);
buf BUF1 (N6552, N6541);
buf BUF1 (N6553, N6546);
or OR4 (N6554, N6553, N6496, N2902, N4799);
xor XOR2 (N6555, N6510, N76);
xor XOR2 (N6556, N6552, N1336);
nand NAND3 (N6557, N6554, N3738, N1813);
xor XOR2 (N6558, N6556, N4368);
nor NOR2 (N6559, N6548, N6308);
nor NOR2 (N6560, N6555, N3922);
buf BUF1 (N6561, N6559);
xor XOR2 (N6562, N6542, N6093);
buf BUF1 (N6563, N6561);
buf BUF1 (N6564, N6558);
nor NOR2 (N6565, N6549, N1605);
or OR3 (N6566, N6551, N5613, N2193);
nor NOR3 (N6567, N6565, N3738, N4879);
buf BUF1 (N6568, N6566);
or OR4 (N6569, N6568, N6389, N3378, N2265);
nand NAND4 (N6570, N6560, N4302, N3419, N5912);
buf BUF1 (N6571, N6564);
xor XOR2 (N6572, N6571, N2360);
buf BUF1 (N6573, N6572);
not NOT1 (N6574, N6545);
xor XOR2 (N6575, N6563, N6050);
nand NAND3 (N6576, N6569, N600, N1348);
nor NOR4 (N6577, N6550, N6188, N889, N199);
nand NAND2 (N6578, N6562, N5192);
and AND3 (N6579, N6557, N1370, N3088);
or OR4 (N6580, N6575, N3064, N6040, N3545);
buf BUF1 (N6581, N6580);
not NOT1 (N6582, N6570);
nand NAND4 (N6583, N6579, N1400, N2313, N4629);
buf BUF1 (N6584, N6583);
nor NOR2 (N6585, N6531, N5116);
buf BUF1 (N6586, N6574);
or OR4 (N6587, N6577, N2469, N177, N5329);
nor NOR2 (N6588, N6567, N1362);
nand NAND2 (N6589, N6582, N1024);
nand NAND3 (N6590, N6586, N653, N3476);
or OR2 (N6591, N6576, N5688);
buf BUF1 (N6592, N6578);
xor XOR2 (N6593, N6591, N1640);
or OR4 (N6594, N6585, N4114, N3009, N6561);
buf BUF1 (N6595, N6593);
xor XOR2 (N6596, N6588, N619);
nand NAND2 (N6597, N6581, N680);
xor XOR2 (N6598, N6597, N3443);
nor NOR2 (N6599, N6584, N5568);
nand NAND3 (N6600, N6589, N5885, N1724);
not NOT1 (N6601, N6594);
not NOT1 (N6602, N6590);
not NOT1 (N6603, N6587);
or OR2 (N6604, N6595, N4140);
nand NAND4 (N6605, N6603, N1558, N3465, N404);
nor NOR3 (N6606, N6598, N969, N4051);
nor NOR4 (N6607, N6606, N3821, N1846, N6430);
and AND4 (N6608, N6602, N3231, N4118, N266);
nand NAND3 (N6609, N6600, N3734, N5355);
or OR4 (N6610, N6607, N1413, N658, N2205);
buf BUF1 (N6611, N6610);
and AND3 (N6612, N6599, N2166, N4948);
nor NOR2 (N6613, N6609, N2275);
buf BUF1 (N6614, N6605);
buf BUF1 (N6615, N6573);
not NOT1 (N6616, N6601);
buf BUF1 (N6617, N6614);
nand NAND4 (N6618, N6604, N2759, N1011, N4498);
buf BUF1 (N6619, N6617);
not NOT1 (N6620, N6612);
xor XOR2 (N6621, N6613, N315);
or OR4 (N6622, N6619, N3755, N3392, N2910);
not NOT1 (N6623, N6616);
and AND2 (N6624, N6615, N2658);
not NOT1 (N6625, N6621);
xor XOR2 (N6626, N6608, N4775);
or OR2 (N6627, N6611, N813);
buf BUF1 (N6628, N6627);
nor NOR4 (N6629, N6592, N1080, N1689, N2444);
and AND2 (N6630, N6624, N1823);
xor XOR2 (N6631, N6622, N2165);
or OR4 (N6632, N6628, N3666, N2457, N2927);
and AND2 (N6633, N6596, N4787);
nor NOR3 (N6634, N6632, N82, N4229);
and AND4 (N6635, N6626, N1824, N4311, N5085);
nor NOR4 (N6636, N6635, N3722, N267, N3711);
xor XOR2 (N6637, N6629, N5194);
buf BUF1 (N6638, N6623);
nor NOR2 (N6639, N6638, N2927);
xor XOR2 (N6640, N6633, N5269);
nand NAND3 (N6641, N6625, N6578, N4898);
nor NOR4 (N6642, N6639, N1721, N2983, N323);
nand NAND3 (N6643, N6642, N4971, N1636);
nor NOR3 (N6644, N6634, N2683, N5448);
or OR4 (N6645, N6637, N4850, N450, N1601);
not NOT1 (N6646, N6631);
nor NOR3 (N6647, N6641, N5535, N395);
xor XOR2 (N6648, N6640, N5326);
buf BUF1 (N6649, N6618);
xor XOR2 (N6650, N6646, N3434);
not NOT1 (N6651, N6645);
and AND4 (N6652, N6636, N5320, N362, N3984);
nor NOR3 (N6653, N6647, N671, N3855);
nand NAND3 (N6654, N6630, N5866, N3523);
nor NOR4 (N6655, N6651, N4964, N4898, N2992);
nand NAND2 (N6656, N6643, N2770);
nor NOR4 (N6657, N6652, N4125, N1516, N4440);
xor XOR2 (N6658, N6649, N4318);
buf BUF1 (N6659, N6648);
nand NAND2 (N6660, N6655, N3183);
nor NOR2 (N6661, N6620, N6322);
buf BUF1 (N6662, N6658);
xor XOR2 (N6663, N6660, N3670);
or OR3 (N6664, N6653, N5209, N1358);
nand NAND3 (N6665, N6662, N4509, N4215);
buf BUF1 (N6666, N6659);
nor NOR3 (N6667, N6666, N5200, N2500);
xor XOR2 (N6668, N6667, N2915);
nand NAND2 (N6669, N6663, N3698);
xor XOR2 (N6670, N6664, N5573);
or OR2 (N6671, N6657, N4903);
nor NOR3 (N6672, N6671, N6173, N578);
and AND2 (N6673, N6670, N5065);
nand NAND4 (N6674, N6668, N2270, N3096, N154);
nor NOR4 (N6675, N6656, N1422, N4105, N3728);
not NOT1 (N6676, N6650);
buf BUF1 (N6677, N6675);
and AND3 (N6678, N6665, N4573, N4844);
buf BUF1 (N6679, N6678);
buf BUF1 (N6680, N6673);
buf BUF1 (N6681, N6677);
not NOT1 (N6682, N6669);
xor XOR2 (N6683, N6674, N4212);
and AND3 (N6684, N6676, N131, N3993);
buf BUF1 (N6685, N6679);
xor XOR2 (N6686, N6680, N5395);
not NOT1 (N6687, N6685);
nand NAND3 (N6688, N6682, N4334, N4181);
or OR3 (N6689, N6683, N1299, N274);
buf BUF1 (N6690, N6644);
buf BUF1 (N6691, N6684);
or OR3 (N6692, N6681, N589, N2428);
and AND2 (N6693, N6692, N3401);
not NOT1 (N6694, N6689);
xor XOR2 (N6695, N6690, N2820);
nor NOR2 (N6696, N6672, N5187);
xor XOR2 (N6697, N6688, N2645);
buf BUF1 (N6698, N6697);
buf BUF1 (N6699, N6696);
not NOT1 (N6700, N6691);
buf BUF1 (N6701, N6698);
xor XOR2 (N6702, N6693, N5378);
nor NOR2 (N6703, N6700, N5355);
not NOT1 (N6704, N6699);
nand NAND2 (N6705, N6654, N6602);
nand NAND2 (N6706, N6703, N1034);
or OR2 (N6707, N6695, N3668);
not NOT1 (N6708, N6702);
buf BUF1 (N6709, N6686);
xor XOR2 (N6710, N6706, N3250);
nand NAND3 (N6711, N6710, N2508, N4209);
and AND4 (N6712, N6661, N3739, N2523, N1716);
and AND2 (N6713, N6705, N2734);
xor XOR2 (N6714, N6704, N549);
nand NAND3 (N6715, N6714, N3625, N5472);
nand NAND4 (N6716, N6711, N3568, N3630, N4052);
or OR2 (N6717, N6701, N5453);
or OR3 (N6718, N6716, N29, N1240);
not NOT1 (N6719, N6715);
not NOT1 (N6720, N6707);
buf BUF1 (N6721, N6712);
nand NAND4 (N6722, N6721, N6031, N4080, N2685);
not NOT1 (N6723, N6694);
not NOT1 (N6724, N6687);
xor XOR2 (N6725, N6723, N1452);
buf BUF1 (N6726, N6718);
xor XOR2 (N6727, N6726, N6270);
xor XOR2 (N6728, N6708, N5923);
xor XOR2 (N6729, N6719, N1541);
nor NOR2 (N6730, N6717, N4018);
nand NAND4 (N6731, N6713, N5823, N2329, N3893);
buf BUF1 (N6732, N6729);
buf BUF1 (N6733, N6728);
nand NAND2 (N6734, N6733, N2907);
buf BUF1 (N6735, N6731);
or OR2 (N6736, N6724, N4745);
and AND4 (N6737, N6722, N327, N3034, N5681);
and AND2 (N6738, N6725, N3922);
nor NOR3 (N6739, N6738, N6451, N4075);
buf BUF1 (N6740, N6736);
or OR2 (N6741, N6737, N3121);
not NOT1 (N6742, N6720);
or OR3 (N6743, N6740, N5216, N3840);
or OR3 (N6744, N6741, N4258, N4573);
nand NAND4 (N6745, N6730, N5906, N3477, N3515);
xor XOR2 (N6746, N6734, N2608);
nor NOR4 (N6747, N6732, N3973, N4616, N4023);
nor NOR2 (N6748, N6743, N525);
not NOT1 (N6749, N6727);
xor XOR2 (N6750, N6744, N3640);
xor XOR2 (N6751, N6742, N3128);
buf BUF1 (N6752, N6746);
not NOT1 (N6753, N6748);
not NOT1 (N6754, N6750);
xor XOR2 (N6755, N6735, N5351);
buf BUF1 (N6756, N6739);
not NOT1 (N6757, N6752);
xor XOR2 (N6758, N6757, N1099);
xor XOR2 (N6759, N6755, N4303);
buf BUF1 (N6760, N6753);
nor NOR3 (N6761, N6759, N1467, N3435);
not NOT1 (N6762, N6745);
or OR4 (N6763, N6762, N5980, N1248, N6098);
nand NAND2 (N6764, N6747, N1505);
nand NAND4 (N6765, N6763, N6186, N4673, N2516);
nor NOR3 (N6766, N6709, N5208, N1972);
xor XOR2 (N6767, N6749, N6439);
buf BUF1 (N6768, N6764);
and AND2 (N6769, N6768, N4732);
nor NOR2 (N6770, N6769, N1509);
and AND2 (N6771, N6756, N615);
xor XOR2 (N6772, N6760, N586);
nand NAND3 (N6773, N6767, N5060, N3361);
nor NOR4 (N6774, N6758, N1346, N669, N4954);
buf BUF1 (N6775, N6766);
and AND2 (N6776, N6754, N5880);
or OR2 (N6777, N6770, N1475);
nor NOR2 (N6778, N6751, N5764);
not NOT1 (N6779, N6777);
nor NOR2 (N6780, N6774, N1725);
buf BUF1 (N6781, N6761);
nand NAND4 (N6782, N6772, N5566, N3650, N6381);
buf BUF1 (N6783, N6782);
buf BUF1 (N6784, N6773);
buf BUF1 (N6785, N6784);
or OR3 (N6786, N6771, N3334, N5198);
nor NOR2 (N6787, N6786, N1745);
not NOT1 (N6788, N6775);
buf BUF1 (N6789, N6780);
buf BUF1 (N6790, N6788);
nor NOR4 (N6791, N6779, N2241, N3988, N1890);
buf BUF1 (N6792, N6778);
xor XOR2 (N6793, N6791, N1911);
not NOT1 (N6794, N6776);
or OR3 (N6795, N6787, N1088, N646);
nor NOR3 (N6796, N6789, N228, N1612);
not NOT1 (N6797, N6793);
buf BUF1 (N6798, N6790);
xor XOR2 (N6799, N6795, N400);
nor NOR2 (N6800, N6799, N6787);
and AND3 (N6801, N6798, N541, N6725);
buf BUF1 (N6802, N6796);
not NOT1 (N6803, N6802);
nor NOR4 (N6804, N6801, N2966, N4716, N6560);
buf BUF1 (N6805, N6781);
xor XOR2 (N6806, N6805, N240);
not NOT1 (N6807, N6785);
nor NOR4 (N6808, N6807, N118, N2958, N1238);
nand NAND4 (N6809, N6800, N5914, N2935, N4692);
xor XOR2 (N6810, N6809, N5830);
buf BUF1 (N6811, N6806);
xor XOR2 (N6812, N6804, N6016);
and AND4 (N6813, N6803, N3733, N1802, N4670);
or OR3 (N6814, N6783, N1576, N2423);
and AND3 (N6815, N6811, N861, N379);
or OR4 (N6816, N6794, N1448, N5425, N246);
or OR4 (N6817, N6814, N4145, N4936, N3474);
buf BUF1 (N6818, N6812);
xor XOR2 (N6819, N6808, N2204);
nand NAND4 (N6820, N6818, N1713, N4531, N2792);
xor XOR2 (N6821, N6817, N4753);
or OR3 (N6822, N6813, N596, N1487);
nand NAND2 (N6823, N6810, N457);
and AND3 (N6824, N6819, N3728, N4490);
not NOT1 (N6825, N6765);
and AND2 (N6826, N6821, N4058);
xor XOR2 (N6827, N6825, N2090);
buf BUF1 (N6828, N6826);
or OR2 (N6829, N6797, N1893);
buf BUF1 (N6830, N6823);
not NOT1 (N6831, N6816);
buf BUF1 (N6832, N6831);
not NOT1 (N6833, N6820);
nand NAND2 (N6834, N6832, N4897);
nor NOR4 (N6835, N6829, N4575, N1657, N2347);
nand NAND4 (N6836, N6824, N232, N6616, N2873);
nor NOR2 (N6837, N6828, N5407);
xor XOR2 (N6838, N6822, N1697);
and AND2 (N6839, N6833, N2848);
not NOT1 (N6840, N6838);
nand NAND2 (N6841, N6815, N2082);
xor XOR2 (N6842, N6835, N6721);
not NOT1 (N6843, N6830);
and AND3 (N6844, N6843, N4236, N5096);
buf BUF1 (N6845, N6827);
or OR3 (N6846, N6841, N1910, N2159);
buf BUF1 (N6847, N6846);
not NOT1 (N6848, N6792);
nor NOR2 (N6849, N6845, N4464);
and AND4 (N6850, N6839, N4886, N3655, N4639);
nor NOR4 (N6851, N6834, N2318, N1734, N5796);
nand NAND4 (N6852, N6842, N6647, N5279, N5617);
or OR3 (N6853, N6836, N3010, N5145);
and AND4 (N6854, N6840, N1125, N5720, N983);
nor NOR4 (N6855, N6852, N229, N2942, N6572);
nand NAND3 (N6856, N6853, N5926, N6720);
buf BUF1 (N6857, N6851);
nor NOR4 (N6858, N6837, N4640, N65, N3983);
or OR4 (N6859, N6858, N3024, N2189, N690);
not NOT1 (N6860, N6850);
or OR2 (N6861, N6848, N6440);
buf BUF1 (N6862, N6859);
nand NAND3 (N6863, N6847, N6592, N6156);
buf BUF1 (N6864, N6860);
xor XOR2 (N6865, N6855, N4971);
nand NAND2 (N6866, N6857, N2787);
nand NAND3 (N6867, N6856, N2713, N4157);
buf BUF1 (N6868, N6862);
xor XOR2 (N6869, N6854, N6224);
or OR2 (N6870, N6864, N305);
buf BUF1 (N6871, N6867);
or OR4 (N6872, N6844, N938, N762, N2227);
or OR2 (N6873, N6869, N1069);
and AND4 (N6874, N6866, N6222, N177, N2024);
buf BUF1 (N6875, N6865);
nor NOR4 (N6876, N6875, N5680, N5440, N1034);
buf BUF1 (N6877, N6863);
nand NAND2 (N6878, N6870, N3326);
nand NAND3 (N6879, N6871, N3494, N6184);
nor NOR4 (N6880, N6873, N6309, N6508, N5115);
or OR2 (N6881, N6878, N2236);
not NOT1 (N6882, N6868);
xor XOR2 (N6883, N6874, N1943);
xor XOR2 (N6884, N6882, N3879);
xor XOR2 (N6885, N6849, N1175);
nor NOR2 (N6886, N6881, N1800);
or OR3 (N6887, N6883, N6343, N3621);
and AND3 (N6888, N6884, N1839, N730);
xor XOR2 (N6889, N6877, N4699);
buf BUF1 (N6890, N6880);
nor NOR2 (N6891, N6886, N3033);
or OR3 (N6892, N6887, N1080, N3417);
or OR4 (N6893, N6885, N6883, N2354, N6429);
not NOT1 (N6894, N6888);
or OR4 (N6895, N6876, N6079, N1501, N469);
not NOT1 (N6896, N6879);
nand NAND2 (N6897, N6896, N5149);
buf BUF1 (N6898, N6890);
nor NOR3 (N6899, N6897, N2895, N624);
xor XOR2 (N6900, N6898, N3009);
not NOT1 (N6901, N6872);
not NOT1 (N6902, N6900);
not NOT1 (N6903, N6889);
not NOT1 (N6904, N6895);
or OR2 (N6905, N6899, N4716);
nor NOR2 (N6906, N6901, N2112);
nand NAND3 (N6907, N6903, N2302, N5561);
and AND2 (N6908, N6861, N1716);
xor XOR2 (N6909, N6905, N3591);
nor NOR3 (N6910, N6909, N932, N1538);
xor XOR2 (N6911, N6904, N2632);
and AND4 (N6912, N6908, N6082, N6403, N4573);
or OR3 (N6913, N6907, N3714, N4674);
and AND3 (N6914, N6891, N1888, N2824);
nand NAND2 (N6915, N6893, N2864);
or OR4 (N6916, N6911, N1186, N3127, N4096);
xor XOR2 (N6917, N6892, N3922);
xor XOR2 (N6918, N6914, N2144);
nand NAND2 (N6919, N6915, N5505);
nor NOR2 (N6920, N6916, N2412);
nor NOR3 (N6921, N6894, N5754, N4294);
or OR4 (N6922, N6910, N3061, N4812, N4634);
nand NAND4 (N6923, N6921, N2568, N5261, N4231);
and AND2 (N6924, N6918, N6696);
xor XOR2 (N6925, N6924, N6788);
buf BUF1 (N6926, N6912);
and AND4 (N6927, N6920, N2313, N4208, N17);
nand NAND2 (N6928, N6926, N175);
not NOT1 (N6929, N6923);
nor NOR4 (N6930, N6928, N2739, N1380, N4645);
buf BUF1 (N6931, N6902);
not NOT1 (N6932, N6913);
nand NAND2 (N6933, N6930, N3477);
not NOT1 (N6934, N6932);
and AND2 (N6935, N6919, N1996);
nand NAND4 (N6936, N6934, N2684, N228, N5664);
buf BUF1 (N6937, N6917);
and AND2 (N6938, N6922, N1286);
nand NAND4 (N6939, N6936, N4428, N1426, N791);
buf BUF1 (N6940, N6938);
or OR3 (N6941, N6925, N3531, N6678);
nor NOR3 (N6942, N6937, N3564, N525);
not NOT1 (N6943, N6939);
not NOT1 (N6944, N6933);
not NOT1 (N6945, N6943);
buf BUF1 (N6946, N6929);
nand NAND3 (N6947, N6931, N1078, N6751);
buf BUF1 (N6948, N6945);
nor NOR4 (N6949, N6942, N4639, N1397, N4285);
buf BUF1 (N6950, N6940);
nand NAND3 (N6951, N6941, N2011, N3537);
and AND3 (N6952, N6948, N2022, N6597);
and AND2 (N6953, N6949, N6118);
and AND3 (N6954, N6946, N4878, N6259);
not NOT1 (N6955, N6950);
buf BUF1 (N6956, N6955);
not NOT1 (N6957, N6947);
not NOT1 (N6958, N6927);
and AND2 (N6959, N6906, N2862);
not NOT1 (N6960, N6956);
or OR4 (N6961, N6944, N3484, N4988, N6493);
nor NOR4 (N6962, N6961, N470, N1024, N2051);
not NOT1 (N6963, N6957);
not NOT1 (N6964, N6952);
or OR3 (N6965, N6935, N6722, N5321);
xor XOR2 (N6966, N6953, N3967);
xor XOR2 (N6967, N6951, N66);
nand NAND3 (N6968, N6962, N3819, N963);
xor XOR2 (N6969, N6967, N1273);
nand NAND4 (N6970, N6969, N1110, N5113, N200);
not NOT1 (N6971, N6954);
buf BUF1 (N6972, N6968);
not NOT1 (N6973, N6963);
buf BUF1 (N6974, N6966);
not NOT1 (N6975, N6971);
nand NAND3 (N6976, N6965, N5617, N6010);
nand NAND3 (N6977, N6959, N6033, N6374);
xor XOR2 (N6978, N6973, N1562);
and AND2 (N6979, N6958, N1572);
nor NOR3 (N6980, N6975, N1495, N357);
buf BUF1 (N6981, N6979);
or OR2 (N6982, N6980, N3617);
and AND2 (N6983, N6981, N5620);
nor NOR3 (N6984, N6978, N1940, N879);
buf BUF1 (N6985, N6972);
nor NOR4 (N6986, N6982, N5187, N2627, N3948);
nor NOR2 (N6987, N6970, N3217);
xor XOR2 (N6988, N6964, N4131);
and AND2 (N6989, N6987, N4639);
nor NOR2 (N6990, N6983, N5928);
not NOT1 (N6991, N6990);
and AND3 (N6992, N6984, N5655, N2997);
nor NOR3 (N6993, N6977, N2168, N1260);
buf BUF1 (N6994, N6960);
and AND3 (N6995, N6992, N4616, N4826);
nor NOR3 (N6996, N6976, N777, N3326);
buf BUF1 (N6997, N6995);
and AND4 (N6998, N6974, N1523, N5465, N3302);
and AND3 (N6999, N6989, N600, N363);
nand NAND3 (N7000, N6993, N1826, N6763);
buf BUF1 (N7001, N6985);
buf BUF1 (N7002, N6996);
nor NOR3 (N7003, N6998, N1063, N3384);
buf BUF1 (N7004, N6991);
nand NAND3 (N7005, N6994, N6180, N4071);
and AND2 (N7006, N7004, N5421);
or OR3 (N7007, N6999, N997, N3654);
or OR2 (N7008, N7000, N1152);
or OR2 (N7009, N7007, N196);
nor NOR3 (N7010, N7009, N4465, N5351);
nor NOR3 (N7011, N7006, N3655, N2703);
and AND3 (N7012, N6986, N6411, N474);
not NOT1 (N7013, N6997);
xor XOR2 (N7014, N7012, N6980);
not NOT1 (N7015, N7005);
nand NAND4 (N7016, N6988, N276, N4063, N2964);
nand NAND4 (N7017, N7016, N5871, N6455, N5532);
buf BUF1 (N7018, N7002);
or OR4 (N7019, N7003, N5450, N2265, N4548);
xor XOR2 (N7020, N7015, N6199);
xor XOR2 (N7021, N7010, N3580);
xor XOR2 (N7022, N7014, N3208);
xor XOR2 (N7023, N7021, N6357);
buf BUF1 (N7024, N7013);
not NOT1 (N7025, N7008);
buf BUF1 (N7026, N7020);
or OR2 (N7027, N7019, N421);
nor NOR2 (N7028, N7011, N6628);
nor NOR4 (N7029, N7001, N2089, N5746, N2657);
and AND3 (N7030, N7022, N7015, N5662);
or OR4 (N7031, N7028, N4356, N3873, N1737);
nand NAND4 (N7032, N7030, N664, N369, N5402);
buf BUF1 (N7033, N7017);
not NOT1 (N7034, N7018);
xor XOR2 (N7035, N7031, N4984);
xor XOR2 (N7036, N7034, N2437);
not NOT1 (N7037, N7026);
nor NOR4 (N7038, N7033, N272, N2890, N4394);
nand NAND4 (N7039, N7029, N5585, N3787, N6488);
or OR2 (N7040, N7024, N5430);
not NOT1 (N7041, N7038);
and AND4 (N7042, N7027, N1343, N1647, N4247);
nor NOR3 (N7043, N7025, N1934, N6331);
xor XOR2 (N7044, N7036, N1568);
buf BUF1 (N7045, N7023);
not NOT1 (N7046, N7039);
nor NOR2 (N7047, N7045, N6887);
buf BUF1 (N7048, N7035);
not NOT1 (N7049, N7042);
and AND4 (N7050, N7048, N4222, N6670, N3496);
and AND3 (N7051, N7044, N998, N3576);
nand NAND2 (N7052, N7040, N5741);
or OR4 (N7053, N7051, N152, N3394, N4204);
nand NAND3 (N7054, N7041, N6886, N6117);
nand NAND3 (N7055, N7053, N6977, N4263);
xor XOR2 (N7056, N7046, N2859);
and AND2 (N7057, N7054, N606);
nand NAND4 (N7058, N7052, N6778, N3682, N5565);
not NOT1 (N7059, N7050);
and AND4 (N7060, N7057, N3173, N2617, N295);
nor NOR4 (N7061, N7032, N1427, N2571, N1770);
and AND2 (N7062, N7037, N2246);
nand NAND3 (N7063, N7043, N5773, N5599);
or OR2 (N7064, N7063, N5109);
xor XOR2 (N7065, N7064, N1529);
nand NAND2 (N7066, N7065, N2489);
xor XOR2 (N7067, N7066, N2090);
xor XOR2 (N7068, N7067, N2963);
xor XOR2 (N7069, N7056, N1751);
nand NAND3 (N7070, N7068, N4388, N5294);
nand NAND3 (N7071, N7069, N2682, N3707);
nand NAND4 (N7072, N7049, N4394, N4715, N3699);
nand NAND2 (N7073, N7055, N1813);
nor NOR4 (N7074, N7058, N225, N5389, N6863);
or OR2 (N7075, N7072, N4840);
buf BUF1 (N7076, N7073);
not NOT1 (N7077, N7075);
not NOT1 (N7078, N7074);
and AND3 (N7079, N7062, N786, N4565);
nand NAND2 (N7080, N7071, N2086);
nor NOR2 (N7081, N7079, N5544);
nor NOR2 (N7082, N7076, N3629);
and AND3 (N7083, N7078, N29, N2594);
and AND2 (N7084, N7047, N4888);
buf BUF1 (N7085, N7080);
buf BUF1 (N7086, N7085);
or OR2 (N7087, N7083, N4347);
or OR3 (N7088, N7087, N215, N3625);
or OR3 (N7089, N7086, N1958, N4263);
nand NAND4 (N7090, N7089, N3924, N6042, N4466);
xor XOR2 (N7091, N7081, N6525);
xor XOR2 (N7092, N7070, N6828);
buf BUF1 (N7093, N7082);
not NOT1 (N7094, N7091);
nand NAND2 (N7095, N7084, N834);
or OR2 (N7096, N7088, N6430);
buf BUF1 (N7097, N7094);
not NOT1 (N7098, N7093);
nand NAND2 (N7099, N7095, N1245);
xor XOR2 (N7100, N7061, N6822);
not NOT1 (N7101, N7098);
nor NOR3 (N7102, N7096, N4123, N6926);
or OR2 (N7103, N7059, N770);
xor XOR2 (N7104, N7060, N1122);
not NOT1 (N7105, N7104);
buf BUF1 (N7106, N7097);
or OR2 (N7107, N7100, N1132);
xor XOR2 (N7108, N7107, N6487);
buf BUF1 (N7109, N7108);
xor XOR2 (N7110, N7099, N6485);
not NOT1 (N7111, N7109);
not NOT1 (N7112, N7101);
xor XOR2 (N7113, N7110, N841);
nor NOR2 (N7114, N7077, N2265);
or OR2 (N7115, N7111, N4295);
nand NAND3 (N7116, N7106, N6227, N3614);
nor NOR2 (N7117, N7105, N3170);
xor XOR2 (N7118, N7092, N5650);
xor XOR2 (N7119, N7118, N1844);
not NOT1 (N7120, N7116);
not NOT1 (N7121, N7112);
not NOT1 (N7122, N7114);
xor XOR2 (N7123, N7090, N1509);
nor NOR3 (N7124, N7113, N4121, N5199);
nor NOR3 (N7125, N7117, N4418, N2270);
xor XOR2 (N7126, N7122, N6961);
nor NOR4 (N7127, N7102, N6003, N4963, N3602);
and AND2 (N7128, N7103, N3174);
or OR4 (N7129, N7119, N3482, N2152, N4617);
nand NAND3 (N7130, N7125, N1601, N7019);
buf BUF1 (N7131, N7126);
and AND4 (N7132, N7128, N6326, N4948, N1729);
or OR3 (N7133, N7129, N4695, N832);
nor NOR4 (N7134, N7123, N1826, N3549, N5447);
xor XOR2 (N7135, N7115, N5770);
not NOT1 (N7136, N7127);
buf BUF1 (N7137, N7133);
not NOT1 (N7138, N7132);
and AND3 (N7139, N7120, N3917, N2038);
or OR4 (N7140, N7124, N211, N1932, N4722);
buf BUF1 (N7141, N7139);
not NOT1 (N7142, N7131);
or OR2 (N7143, N7137, N4494);
not NOT1 (N7144, N7141);
nand NAND2 (N7145, N7142, N2122);
nand NAND3 (N7146, N7144, N4182, N6591);
nand NAND2 (N7147, N7130, N4379);
and AND2 (N7148, N7145, N2852);
xor XOR2 (N7149, N7143, N4983);
or OR2 (N7150, N7138, N1713);
xor XOR2 (N7151, N7146, N3502);
not NOT1 (N7152, N7135);
nand NAND2 (N7153, N7152, N2741);
or OR3 (N7154, N7150, N2695, N4205);
nor NOR4 (N7155, N7151, N870, N6982, N871);
not NOT1 (N7156, N7136);
buf BUF1 (N7157, N7148);
not NOT1 (N7158, N7140);
and AND3 (N7159, N7149, N671, N1165);
or OR2 (N7160, N7159, N5835);
and AND2 (N7161, N7155, N1112);
nor NOR3 (N7162, N7153, N6216, N5625);
xor XOR2 (N7163, N7147, N4260);
nand NAND4 (N7164, N7121, N7022, N1925, N3879);
or OR4 (N7165, N7161, N5489, N5730, N3249);
buf BUF1 (N7166, N7157);
not NOT1 (N7167, N7154);
or OR4 (N7168, N7160, N1186, N2312, N2173);
xor XOR2 (N7169, N7162, N5946);
xor XOR2 (N7170, N7165, N6202);
xor XOR2 (N7171, N7168, N132);
not NOT1 (N7172, N7171);
xor XOR2 (N7173, N7163, N6489);
xor XOR2 (N7174, N7158, N7155);
or OR3 (N7175, N7167, N405, N5790);
nand NAND4 (N7176, N7175, N5564, N7119, N1158);
not NOT1 (N7177, N7169);
buf BUF1 (N7178, N7166);
buf BUF1 (N7179, N7177);
not NOT1 (N7180, N7172);
nor NOR4 (N7181, N7173, N74, N4657, N5066);
nand NAND4 (N7182, N7156, N1748, N109, N7033);
not NOT1 (N7183, N7174);
and AND3 (N7184, N7180, N854, N4972);
and AND2 (N7185, N7164, N6748);
not NOT1 (N7186, N7183);
xor XOR2 (N7187, N7134, N1925);
or OR3 (N7188, N7184, N1734, N3294);
xor XOR2 (N7189, N7185, N2955);
and AND2 (N7190, N7186, N5485);
not NOT1 (N7191, N7170);
buf BUF1 (N7192, N7176);
not NOT1 (N7193, N7179);
or OR4 (N7194, N7191, N1730, N2368, N4989);
and AND4 (N7195, N7194, N500, N5767, N4976);
or OR2 (N7196, N7178, N2895);
not NOT1 (N7197, N7192);
nor NOR4 (N7198, N7182, N1507, N4709, N1159);
nand NAND4 (N7199, N7189, N3257, N3519, N6743);
and AND2 (N7200, N7197, N4308);
nor NOR2 (N7201, N7188, N4159);
xor XOR2 (N7202, N7201, N6449);
or OR3 (N7203, N7202, N4692, N4710);
buf BUF1 (N7204, N7195);
nand NAND2 (N7205, N7204, N4041);
and AND2 (N7206, N7198, N4267);
xor XOR2 (N7207, N7187, N6546);
not NOT1 (N7208, N7196);
nor NOR4 (N7209, N7205, N4575, N3467, N4804);
nor NOR3 (N7210, N7206, N5119, N2843);
not NOT1 (N7211, N7200);
nor NOR4 (N7212, N7208, N1652, N5755, N2813);
nand NAND4 (N7213, N7211, N1120, N718, N3463);
nand NAND2 (N7214, N7213, N159);
xor XOR2 (N7215, N7190, N6227);
or OR4 (N7216, N7209, N1509, N5400, N416);
not NOT1 (N7217, N7207);
buf BUF1 (N7218, N7216);
not NOT1 (N7219, N7214);
nor NOR2 (N7220, N7219, N777);
buf BUF1 (N7221, N7203);
not NOT1 (N7222, N7218);
or OR2 (N7223, N7199, N3933);
and AND4 (N7224, N7223, N3571, N7110, N2504);
nor NOR3 (N7225, N7212, N6253, N6034);
nand NAND3 (N7226, N7210, N3242, N3576);
or OR4 (N7227, N7224, N6228, N2925, N1139);
nor NOR2 (N7228, N7215, N4790);
nor NOR3 (N7229, N7221, N1547, N5841);
and AND2 (N7230, N7217, N7071);
nor NOR2 (N7231, N7226, N2812);
nor NOR4 (N7232, N7228, N1095, N6363, N3247);
nand NAND3 (N7233, N7227, N5694, N3223);
nor NOR3 (N7234, N7231, N5465, N6182);
and AND4 (N7235, N7220, N2078, N3334, N2555);
xor XOR2 (N7236, N7181, N3144);
or OR4 (N7237, N7233, N6015, N3154, N1774);
and AND3 (N7238, N7230, N1446, N5558);
or OR3 (N7239, N7236, N7116, N1654);
xor XOR2 (N7240, N7237, N6853);
not NOT1 (N7241, N7232);
xor XOR2 (N7242, N7235, N6210);
or OR3 (N7243, N7234, N5292, N1967);
or OR3 (N7244, N7225, N2527, N6816);
nand NAND3 (N7245, N7193, N414, N4814);
not NOT1 (N7246, N7238);
nand NAND4 (N7247, N7245, N4204, N1875, N4000);
xor XOR2 (N7248, N7242, N3272);
not NOT1 (N7249, N7241);
xor XOR2 (N7250, N7240, N1566);
and AND3 (N7251, N7250, N4072, N444);
xor XOR2 (N7252, N7239, N3999);
nor NOR4 (N7253, N7244, N2985, N5603, N1883);
nand NAND2 (N7254, N7251, N3711);
xor XOR2 (N7255, N7246, N5269);
not NOT1 (N7256, N7252);
buf BUF1 (N7257, N7253);
nand NAND4 (N7258, N7254, N3722, N6791, N2612);
nor NOR3 (N7259, N7222, N5703, N3034);
or OR4 (N7260, N7257, N6860, N3308, N2082);
xor XOR2 (N7261, N7248, N1213);
xor XOR2 (N7262, N7260, N4828);
or OR2 (N7263, N7247, N6962);
not NOT1 (N7264, N7263);
or OR4 (N7265, N7255, N2299, N4113, N1381);
and AND4 (N7266, N7249, N1314, N6495, N368);
buf BUF1 (N7267, N7243);
buf BUF1 (N7268, N7258);
or OR3 (N7269, N7261, N6999, N3104);
not NOT1 (N7270, N7268);
xor XOR2 (N7271, N7256, N3431);
not NOT1 (N7272, N7264);
nand NAND2 (N7273, N7265, N6769);
nand NAND2 (N7274, N7269, N782);
and AND3 (N7275, N7259, N956, N4067);
and AND2 (N7276, N7267, N7141);
xor XOR2 (N7277, N7275, N1859);
nand NAND2 (N7278, N7273, N1128);
or OR2 (N7279, N7271, N6189);
buf BUF1 (N7280, N7279);
xor XOR2 (N7281, N7266, N4196);
and AND3 (N7282, N7270, N985, N6576);
nor NOR4 (N7283, N7278, N1212, N6888, N122);
xor XOR2 (N7284, N7262, N3650);
not NOT1 (N7285, N7277);
nor NOR3 (N7286, N7272, N1569, N2629);
nand NAND4 (N7287, N7229, N1311, N5654, N4138);
buf BUF1 (N7288, N7284);
xor XOR2 (N7289, N7276, N4766);
nand NAND3 (N7290, N7287, N2331, N1829);
and AND3 (N7291, N7286, N1714, N2440);
not NOT1 (N7292, N7282);
not NOT1 (N7293, N7290);
buf BUF1 (N7294, N7280);
and AND2 (N7295, N7288, N5107);
xor XOR2 (N7296, N7295, N7140);
nor NOR3 (N7297, N7283, N4240, N4123);
or OR2 (N7298, N7292, N6119);
buf BUF1 (N7299, N7274);
or OR3 (N7300, N7289, N6923, N6958);
or OR3 (N7301, N7299, N5144, N4814);
buf BUF1 (N7302, N7296);
xor XOR2 (N7303, N7300, N3313);
buf BUF1 (N7304, N7297);
xor XOR2 (N7305, N7291, N3687);
xor XOR2 (N7306, N7285, N88);
or OR4 (N7307, N7304, N3756, N1572, N2129);
or OR4 (N7308, N7298, N3589, N6277, N2324);
not NOT1 (N7309, N7307);
and AND3 (N7310, N7303, N1155, N5585);
xor XOR2 (N7311, N7294, N680);
and AND2 (N7312, N7281, N1729);
nand NAND3 (N7313, N7312, N5727, N1225);
nor NOR2 (N7314, N7309, N5126);
nand NAND4 (N7315, N7305, N3481, N2575, N4940);
buf BUF1 (N7316, N7301);
not NOT1 (N7317, N7308);
not NOT1 (N7318, N7315);
not NOT1 (N7319, N7313);
nor NOR3 (N7320, N7319, N2659, N4094);
not NOT1 (N7321, N7320);
nor NOR4 (N7322, N7302, N6121, N1583, N6532);
nor NOR2 (N7323, N7321, N1264);
xor XOR2 (N7324, N7323, N1228);
nand NAND4 (N7325, N7314, N6354, N3077, N6771);
nand NAND2 (N7326, N7306, N6319);
buf BUF1 (N7327, N7316);
xor XOR2 (N7328, N7325, N6389);
xor XOR2 (N7329, N7327, N4673);
xor XOR2 (N7330, N7318, N3003);
not NOT1 (N7331, N7326);
or OR3 (N7332, N7328, N3068, N2308);
not NOT1 (N7333, N7331);
or OR2 (N7334, N7293, N5736);
not NOT1 (N7335, N7324);
buf BUF1 (N7336, N7334);
or OR2 (N7337, N7329, N1448);
nor NOR2 (N7338, N7336, N5886);
xor XOR2 (N7339, N7330, N2738);
nor NOR4 (N7340, N7310, N2171, N2421, N4318);
nor NOR2 (N7341, N7311, N5492);
buf BUF1 (N7342, N7337);
and AND4 (N7343, N7332, N4253, N4938, N5873);
buf BUF1 (N7344, N7341);
nand NAND3 (N7345, N7338, N3758, N6924);
or OR4 (N7346, N7322, N2200, N7293, N3907);
nor NOR2 (N7347, N7317, N1828);
nor NOR3 (N7348, N7339, N648, N6832);
and AND3 (N7349, N7335, N1773, N6529);
buf BUF1 (N7350, N7343);
or OR2 (N7351, N7347, N254);
buf BUF1 (N7352, N7333);
buf BUF1 (N7353, N7345);
not NOT1 (N7354, N7352);
and AND2 (N7355, N7350, N7219);
not NOT1 (N7356, N7353);
or OR4 (N7357, N7342, N2282, N248, N2751);
buf BUF1 (N7358, N7355);
or OR4 (N7359, N7340, N2432, N1644, N472);
nand NAND3 (N7360, N7344, N119, N6668);
not NOT1 (N7361, N7356);
buf BUF1 (N7362, N7346);
or OR4 (N7363, N7362, N5376, N2343, N3048);
nor NOR3 (N7364, N7359, N53, N4411);
not NOT1 (N7365, N7354);
or OR3 (N7366, N7358, N382, N1545);
buf BUF1 (N7367, N7366);
or OR4 (N7368, N7348, N6784, N6466, N2101);
and AND3 (N7369, N7367, N3200, N310);
not NOT1 (N7370, N7349);
xor XOR2 (N7371, N7365, N4955);
nand NAND2 (N7372, N7371, N3717);
not NOT1 (N7373, N7361);
buf BUF1 (N7374, N7368);
or OR4 (N7375, N7351, N2240, N6823, N5780);
nand NAND2 (N7376, N7363, N447);
or OR4 (N7377, N7369, N6942, N7342, N2440);
nand NAND2 (N7378, N7360, N5561);
nor NOR4 (N7379, N7377, N3345, N930, N6972);
xor XOR2 (N7380, N7378, N497);
buf BUF1 (N7381, N7375);
not NOT1 (N7382, N7374);
buf BUF1 (N7383, N7372);
and AND3 (N7384, N7379, N2863, N2978);
not NOT1 (N7385, N7373);
or OR2 (N7386, N7376, N1892);
not NOT1 (N7387, N7364);
xor XOR2 (N7388, N7387, N3192);
and AND3 (N7389, N7384, N1278, N1085);
not NOT1 (N7390, N7383);
nor NOR4 (N7391, N7389, N4691, N4123, N5123);
buf BUF1 (N7392, N7390);
nor NOR4 (N7393, N7357, N5935, N4141, N3050);
not NOT1 (N7394, N7380);
and AND3 (N7395, N7388, N2033, N170);
nor NOR4 (N7396, N7395, N6396, N3083, N5095);
or OR2 (N7397, N7385, N5986);
nor NOR4 (N7398, N7370, N254, N3152, N5103);
and AND2 (N7399, N7394, N2543);
buf BUF1 (N7400, N7393);
xor XOR2 (N7401, N7381, N6416);
or OR4 (N7402, N7386, N6047, N2396, N5998);
xor XOR2 (N7403, N7402, N388);
nand NAND3 (N7404, N7392, N2344, N661);
xor XOR2 (N7405, N7400, N4621);
xor XOR2 (N7406, N7401, N7153);
nand NAND4 (N7407, N7405, N3233, N601, N5534);
nand NAND3 (N7408, N7406, N1966, N3237);
buf BUF1 (N7409, N7399);
not NOT1 (N7410, N7396);
nor NOR4 (N7411, N7382, N6518, N530, N4964);
and AND2 (N7412, N7391, N1120);
nor NOR2 (N7413, N7411, N808);
nor NOR3 (N7414, N7410, N3319, N5724);
nand NAND3 (N7415, N7414, N2425, N3079);
or OR3 (N7416, N7407, N3263, N4554);
or OR3 (N7417, N7404, N2888, N2450);
xor XOR2 (N7418, N7417, N1593);
and AND4 (N7419, N7416, N829, N6961, N4426);
nor NOR3 (N7420, N7419, N4417, N3373);
nand NAND2 (N7421, N7397, N3552);
nand NAND3 (N7422, N7412, N1334, N2975);
nor NOR3 (N7423, N7398, N6488, N466);
buf BUF1 (N7424, N7409);
and AND2 (N7425, N7418, N6223);
nand NAND3 (N7426, N7420, N2662, N5738);
buf BUF1 (N7427, N7403);
or OR2 (N7428, N7425, N1550);
not NOT1 (N7429, N7415);
nand NAND4 (N7430, N7421, N6992, N3010, N6978);
and AND2 (N7431, N7428, N6694);
and AND2 (N7432, N7424, N2598);
xor XOR2 (N7433, N7429, N5830);
xor XOR2 (N7434, N7431, N2231);
xor XOR2 (N7435, N7413, N5365);
buf BUF1 (N7436, N7423);
not NOT1 (N7437, N7408);
xor XOR2 (N7438, N7433, N4465);
nand NAND2 (N7439, N7435, N6683);
nand NAND4 (N7440, N7439, N7170, N6696, N1474);
buf BUF1 (N7441, N7432);
nor NOR2 (N7442, N7436, N1627);
nor NOR2 (N7443, N7442, N3698);
and AND2 (N7444, N7426, N1729);
and AND2 (N7445, N7430, N6489);
nor NOR2 (N7446, N7444, N3075);
not NOT1 (N7447, N7445);
buf BUF1 (N7448, N7443);
or OR4 (N7449, N7437, N1414, N1457, N6847);
not NOT1 (N7450, N7434);
or OR2 (N7451, N7446, N4412);
or OR3 (N7452, N7451, N7172, N6499);
nand NAND3 (N7453, N7441, N4712, N2559);
nand NAND4 (N7454, N7422, N3622, N6152, N3342);
not NOT1 (N7455, N7453);
or OR3 (N7456, N7455, N5365, N3645);
not NOT1 (N7457, N7454);
buf BUF1 (N7458, N7427);
xor XOR2 (N7459, N7458, N5592);
nand NAND2 (N7460, N7440, N3173);
and AND4 (N7461, N7447, N1149, N7132, N3786);
or OR4 (N7462, N7450, N4397, N165, N7319);
not NOT1 (N7463, N7459);
or OR4 (N7464, N7457, N7412, N4293, N4474);
or OR3 (N7465, N7463, N6408, N4722);
xor XOR2 (N7466, N7462, N5439);
and AND2 (N7467, N7460, N2902);
nand NAND2 (N7468, N7449, N4122);
nor NOR2 (N7469, N7438, N1040);
nand NAND2 (N7470, N7465, N2917);
not NOT1 (N7471, N7461);
xor XOR2 (N7472, N7467, N5174);
and AND2 (N7473, N7464, N729);
not NOT1 (N7474, N7468);
xor XOR2 (N7475, N7474, N2500);
buf BUF1 (N7476, N7466);
or OR3 (N7477, N7472, N3286, N6234);
and AND3 (N7478, N7448, N5449, N4210);
xor XOR2 (N7479, N7456, N3316);
and AND3 (N7480, N7471, N2452, N4098);
and AND4 (N7481, N7470, N6602, N470, N1561);
not NOT1 (N7482, N7478);
nand NAND2 (N7483, N7480, N3595);
xor XOR2 (N7484, N7452, N5066);
nor NOR3 (N7485, N7473, N210, N393);
buf BUF1 (N7486, N7481);
xor XOR2 (N7487, N7469, N4873);
and AND2 (N7488, N7482, N3444);
and AND3 (N7489, N7479, N2166, N3809);
xor XOR2 (N7490, N7475, N2248);
or OR2 (N7491, N7486, N6868);
nand NAND3 (N7492, N7477, N3113, N2727);
xor XOR2 (N7493, N7489, N5694);
nor NOR2 (N7494, N7490, N5823);
or OR4 (N7495, N7483, N4689, N214, N5388);
buf BUF1 (N7496, N7493);
xor XOR2 (N7497, N7488, N2585);
nand NAND2 (N7498, N7496, N4629);
or OR3 (N7499, N7491, N6437, N6454);
nand NAND2 (N7500, N7498, N7179);
nand NAND3 (N7501, N7476, N566, N653);
xor XOR2 (N7502, N7497, N1392);
nor NOR3 (N7503, N7484, N3899, N6055);
and AND4 (N7504, N7502, N7483, N7230, N3600);
nor NOR3 (N7505, N7501, N4808, N5392);
xor XOR2 (N7506, N7505, N4697);
xor XOR2 (N7507, N7506, N3544);
not NOT1 (N7508, N7487);
not NOT1 (N7509, N7503);
or OR3 (N7510, N7494, N7198, N7149);
nor NOR3 (N7511, N7495, N256, N7166);
xor XOR2 (N7512, N7485, N6582);
and AND4 (N7513, N7511, N3944, N5820, N4798);
or OR2 (N7514, N7504, N601);
nor NOR2 (N7515, N7492, N6570);
not NOT1 (N7516, N7499);
nor NOR4 (N7517, N7510, N4505, N2379, N4374);
not NOT1 (N7518, N7512);
or OR2 (N7519, N7518, N7131);
nor NOR4 (N7520, N7509, N5037, N448, N5656);
buf BUF1 (N7521, N7513);
or OR3 (N7522, N7514, N7427, N1018);
and AND2 (N7523, N7517, N90);
or OR2 (N7524, N7522, N3216);
nand NAND4 (N7525, N7507, N1196, N5071, N4415);
nand NAND2 (N7526, N7519, N3336);
and AND3 (N7527, N7515, N5904, N950);
xor XOR2 (N7528, N7527, N4260);
or OR2 (N7529, N7500, N3655);
nand NAND4 (N7530, N7523, N3661, N2680, N6067);
xor XOR2 (N7531, N7516, N6315);
nor NOR2 (N7532, N7508, N4550);
buf BUF1 (N7533, N7531);
nand NAND3 (N7534, N7524, N4716, N1027);
xor XOR2 (N7535, N7525, N1323);
and AND2 (N7536, N7521, N59);
xor XOR2 (N7537, N7530, N5159);
nand NAND4 (N7538, N7529, N4220, N1491, N4619);
or OR3 (N7539, N7520, N2007, N6870);
xor XOR2 (N7540, N7539, N2091);
not NOT1 (N7541, N7528);
or OR4 (N7542, N7536, N5583, N2127, N6085);
nand NAND2 (N7543, N7542, N4301);
buf BUF1 (N7544, N7532);
buf BUF1 (N7545, N7543);
xor XOR2 (N7546, N7540, N1132);
xor XOR2 (N7547, N7526, N888);
nand NAND4 (N7548, N7547, N3195, N1939, N1542);
not NOT1 (N7549, N7534);
not NOT1 (N7550, N7533);
nor NOR4 (N7551, N7550, N1520, N4148, N6204);
not NOT1 (N7552, N7546);
or OR2 (N7553, N7541, N1153);
and AND3 (N7554, N7537, N2205, N1237);
buf BUF1 (N7555, N7551);
and AND3 (N7556, N7555, N5786, N696);
buf BUF1 (N7557, N7554);
buf BUF1 (N7558, N7552);
and AND3 (N7559, N7549, N1551, N6534);
xor XOR2 (N7560, N7545, N2163);
not NOT1 (N7561, N7557);
buf BUF1 (N7562, N7553);
nand NAND2 (N7563, N7558, N4833);
buf BUF1 (N7564, N7544);
and AND3 (N7565, N7556, N3032, N4353);
nor NOR2 (N7566, N7538, N3881);
nand NAND3 (N7567, N7566, N1540, N305);
nor NOR4 (N7568, N7560, N6525, N3075, N4698);
nor NOR2 (N7569, N7567, N2028);
nand NAND4 (N7570, N7535, N3752, N3246, N3893);
and AND2 (N7571, N7564, N2216);
or OR2 (N7572, N7561, N7355);
not NOT1 (N7573, N7570);
xor XOR2 (N7574, N7562, N4286);
or OR4 (N7575, N7571, N227, N2908, N5184);
and AND2 (N7576, N7572, N6658);
buf BUF1 (N7577, N7568);
buf BUF1 (N7578, N7563);
or OR4 (N7579, N7574, N2781, N3321, N1884);
nor NOR2 (N7580, N7559, N5692);
xor XOR2 (N7581, N7575, N6233);
xor XOR2 (N7582, N7569, N590);
buf BUF1 (N7583, N7565);
or OR3 (N7584, N7548, N5342, N2596);
and AND2 (N7585, N7583, N1788);
xor XOR2 (N7586, N7576, N2949);
nand NAND3 (N7587, N7584, N2171, N3532);
xor XOR2 (N7588, N7586, N3520);
or OR2 (N7589, N7587, N5119);
buf BUF1 (N7590, N7573);
nor NOR4 (N7591, N7585, N3336, N1153, N627);
and AND3 (N7592, N7580, N4150, N2202);
buf BUF1 (N7593, N7581);
or OR2 (N7594, N7578, N5611);
not NOT1 (N7595, N7577);
nand NAND2 (N7596, N7579, N6944);
xor XOR2 (N7597, N7593, N5074);
and AND2 (N7598, N7591, N98);
and AND2 (N7599, N7588, N4394);
and AND4 (N7600, N7598, N4155, N5343, N4139);
not NOT1 (N7601, N7594);
not NOT1 (N7602, N7595);
xor XOR2 (N7603, N7601, N5340);
xor XOR2 (N7604, N7582, N3616);
and AND4 (N7605, N7602, N2627, N5914, N2853);
nor NOR4 (N7606, N7604, N2359, N5753, N3131);
buf BUF1 (N7607, N7589);
or OR2 (N7608, N7607, N1482);
nor NOR3 (N7609, N7590, N661, N3517);
buf BUF1 (N7610, N7597);
nand NAND2 (N7611, N7596, N1302);
nor NOR2 (N7612, N7592, N2106);
xor XOR2 (N7613, N7605, N1624);
or OR4 (N7614, N7599, N1363, N3500, N21);
nand NAND3 (N7615, N7609, N4460, N1005);
nor NOR3 (N7616, N7608, N7240, N1453);
buf BUF1 (N7617, N7611);
nand NAND3 (N7618, N7614, N5260, N6292);
nand NAND3 (N7619, N7616, N3259, N2737);
or OR3 (N7620, N7610, N2219, N4132);
buf BUF1 (N7621, N7617);
nor NOR2 (N7622, N7613, N1278);
nand NAND3 (N7623, N7612, N812, N5212);
not NOT1 (N7624, N7603);
nor NOR2 (N7625, N7615, N5678);
or OR4 (N7626, N7625, N4720, N2902, N3938);
xor XOR2 (N7627, N7619, N5057);
or OR4 (N7628, N7600, N1251, N1248, N2721);
nand NAND4 (N7629, N7627, N7274, N1701, N3218);
xor XOR2 (N7630, N7623, N5857);
and AND3 (N7631, N7630, N6418, N7420);
buf BUF1 (N7632, N7618);
xor XOR2 (N7633, N7606, N7236);
buf BUF1 (N7634, N7632);
nand NAND2 (N7635, N7620, N107);
nor NOR3 (N7636, N7631, N517, N5831);
nand NAND4 (N7637, N7622, N6184, N4008, N2438);
not NOT1 (N7638, N7633);
nor NOR3 (N7639, N7636, N40, N273);
buf BUF1 (N7640, N7626);
nand NAND2 (N7641, N7634, N2762);
nand NAND2 (N7642, N7639, N867);
and AND3 (N7643, N7641, N2201, N3955);
or OR2 (N7644, N7635, N4551);
or OR3 (N7645, N7628, N2204, N1153);
nand NAND4 (N7646, N7642, N1104, N1422, N3395);
or OR4 (N7647, N7637, N6100, N3553, N1289);
buf BUF1 (N7648, N7643);
and AND3 (N7649, N7646, N4040, N4469);
nor NOR3 (N7650, N7648, N3064, N5910);
buf BUF1 (N7651, N7645);
nor NOR4 (N7652, N7651, N1207, N530, N862);
nor NOR4 (N7653, N7629, N5948, N5000, N307);
not NOT1 (N7654, N7649);
and AND4 (N7655, N7621, N6103, N7142, N5766);
nor NOR4 (N7656, N7655, N6275, N7532, N2845);
not NOT1 (N7657, N7653);
or OR2 (N7658, N7624, N7284);
nor NOR2 (N7659, N7658, N3724);
nor NOR2 (N7660, N7640, N7408);
xor XOR2 (N7661, N7657, N1356);
nor NOR3 (N7662, N7644, N2296, N1294);
and AND4 (N7663, N7660, N5813, N3734, N6528);
and AND2 (N7664, N7656, N7219);
or OR4 (N7665, N7661, N3781, N4497, N1325);
or OR2 (N7666, N7652, N667);
and AND3 (N7667, N7665, N7416, N703);
buf BUF1 (N7668, N7664);
not NOT1 (N7669, N7662);
or OR3 (N7670, N7666, N5023, N1637);
nor NOR3 (N7671, N7659, N3222, N2263);
nand NAND4 (N7672, N7650, N2342, N4191, N6064);
nand NAND3 (N7673, N7647, N3495, N843);
nand NAND2 (N7674, N7673, N7497);
not NOT1 (N7675, N7674);
nand NAND2 (N7676, N7667, N5530);
and AND4 (N7677, N7672, N4221, N606, N6795);
nand NAND4 (N7678, N7671, N3307, N2221, N5052);
nand NAND4 (N7679, N7678, N545, N6295, N6630);
xor XOR2 (N7680, N7669, N25);
nand NAND3 (N7681, N7670, N3387, N2875);
not NOT1 (N7682, N7680);
nand NAND2 (N7683, N7638, N2630);
buf BUF1 (N7684, N7679);
nor NOR3 (N7685, N7663, N2802, N5453);
and AND4 (N7686, N7684, N2236, N3589, N3654);
xor XOR2 (N7687, N7677, N3982);
xor XOR2 (N7688, N7654, N6483);
nand NAND2 (N7689, N7683, N3979);
and AND4 (N7690, N7668, N1906, N7484, N1925);
nor NOR3 (N7691, N7690, N4387, N1402);
and AND2 (N7692, N7691, N7247);
or OR2 (N7693, N7692, N3630);
xor XOR2 (N7694, N7675, N694);
or OR3 (N7695, N7681, N4211, N2490);
xor XOR2 (N7696, N7685, N3831);
and AND4 (N7697, N7682, N3915, N3504, N5669);
nand NAND4 (N7698, N7686, N2347, N4822, N1138);
and AND4 (N7699, N7689, N6651, N3672, N4607);
buf BUF1 (N7700, N7687);
buf BUF1 (N7701, N7676);
not NOT1 (N7702, N7693);
buf BUF1 (N7703, N7694);
and AND4 (N7704, N7701, N6071, N6056, N63);
xor XOR2 (N7705, N7697, N2534);
buf BUF1 (N7706, N7702);
or OR3 (N7707, N7703, N1221, N363);
not NOT1 (N7708, N7705);
not NOT1 (N7709, N7698);
nor NOR3 (N7710, N7706, N5248, N6067);
nand NAND4 (N7711, N7707, N1966, N7185, N2862);
buf BUF1 (N7712, N7711);
buf BUF1 (N7713, N7699);
nor NOR2 (N7714, N7700, N7299);
and AND4 (N7715, N7688, N389, N258, N5233);
nor NOR3 (N7716, N7696, N7224, N3760);
xor XOR2 (N7717, N7712, N6504);
not NOT1 (N7718, N7716);
buf BUF1 (N7719, N7709);
not NOT1 (N7720, N7708);
or OR4 (N7721, N7713, N3039, N7245, N816);
not NOT1 (N7722, N7710);
not NOT1 (N7723, N7722);
and AND4 (N7724, N7718, N1178, N4383, N3244);
xor XOR2 (N7725, N7721, N5325);
xor XOR2 (N7726, N7724, N7526);
nor NOR2 (N7727, N7704, N1423);
and AND4 (N7728, N7727, N4964, N7218, N2576);
or OR4 (N7729, N7723, N7706, N4763, N6708);
nor NOR4 (N7730, N7719, N5797, N4461, N5192);
xor XOR2 (N7731, N7726, N1395);
buf BUF1 (N7732, N7715);
not NOT1 (N7733, N7725);
not NOT1 (N7734, N7720);
not NOT1 (N7735, N7730);
or OR3 (N7736, N7729, N3685, N6128);
buf BUF1 (N7737, N7733);
and AND3 (N7738, N7734, N6075, N3498);
buf BUF1 (N7739, N7714);
not NOT1 (N7740, N7728);
not NOT1 (N7741, N7732);
xor XOR2 (N7742, N7739, N615);
buf BUF1 (N7743, N7737);
not NOT1 (N7744, N7695);
nand NAND2 (N7745, N7735, N1526);
and AND3 (N7746, N7741, N3992, N6179);
xor XOR2 (N7747, N7742, N1759);
or OR4 (N7748, N7738, N4737, N307, N2255);
or OR2 (N7749, N7731, N3699);
nand NAND4 (N7750, N7743, N1018, N3973, N3714);
or OR2 (N7751, N7746, N1745);
nor NOR2 (N7752, N7750, N4956);
and AND3 (N7753, N7740, N5966, N5663);
or OR4 (N7754, N7751, N3008, N6661, N6775);
and AND2 (N7755, N7753, N4826);
nand NAND4 (N7756, N7749, N5584, N3988, N4730);
buf BUF1 (N7757, N7752);
not NOT1 (N7758, N7748);
buf BUF1 (N7759, N7747);
or OR2 (N7760, N7759, N4403);
not NOT1 (N7761, N7744);
not NOT1 (N7762, N7760);
xor XOR2 (N7763, N7758, N7611);
not NOT1 (N7764, N7762);
or OR4 (N7765, N7764, N4189, N2216, N1126);
nand NAND3 (N7766, N7755, N67, N3699);
xor XOR2 (N7767, N7717, N2192);
nand NAND2 (N7768, N7761, N730);
and AND3 (N7769, N7757, N6081, N4864);
nand NAND3 (N7770, N7756, N6739, N5112);
or OR2 (N7771, N7736, N4050);
xor XOR2 (N7772, N7771, N754);
or OR2 (N7773, N7768, N1670);
or OR3 (N7774, N7772, N3815, N6958);
and AND4 (N7775, N7774, N1960, N2003, N7300);
buf BUF1 (N7776, N7767);
xor XOR2 (N7777, N7745, N4557);
not NOT1 (N7778, N7754);
nor NOR3 (N7779, N7763, N442, N3491);
not NOT1 (N7780, N7765);
buf BUF1 (N7781, N7777);
nor NOR2 (N7782, N7775, N1685);
and AND3 (N7783, N7781, N6733, N757);
xor XOR2 (N7784, N7766, N2247);
buf BUF1 (N7785, N7776);
xor XOR2 (N7786, N7779, N6021);
nor NOR3 (N7787, N7780, N2297, N1661);
and AND2 (N7788, N7782, N6927);
and AND3 (N7789, N7769, N1885, N5014);
and AND4 (N7790, N7778, N3649, N5744, N5485);
or OR2 (N7791, N7770, N4597);
nand NAND4 (N7792, N7787, N5341, N3341, N248);
or OR2 (N7793, N7791, N6926);
or OR3 (N7794, N7784, N7740, N2514);
nand NAND2 (N7795, N7773, N1064);
nor NOR4 (N7796, N7794, N5375, N27, N6686);
nor NOR4 (N7797, N7796, N3743, N4394, N2772);
and AND3 (N7798, N7795, N6236, N1493);
not NOT1 (N7799, N7790);
and AND4 (N7800, N7786, N3112, N7178, N5010);
buf BUF1 (N7801, N7799);
not NOT1 (N7802, N7783);
nor NOR3 (N7803, N7789, N956, N1497);
buf BUF1 (N7804, N7801);
not NOT1 (N7805, N7792);
buf BUF1 (N7806, N7804);
not NOT1 (N7807, N7797);
nand NAND4 (N7808, N7802, N4475, N1171, N1113);
not NOT1 (N7809, N7788);
or OR3 (N7810, N7808, N4534, N62);
or OR2 (N7811, N7785, N6055);
buf BUF1 (N7812, N7798);
or OR4 (N7813, N7803, N5972, N4488, N5652);
xor XOR2 (N7814, N7793, N2990);
and AND3 (N7815, N7814, N7091, N7434);
or OR2 (N7816, N7811, N7692);
and AND4 (N7817, N7807, N2943, N3936, N4881);
xor XOR2 (N7818, N7813, N5503);
nor NOR2 (N7819, N7806, N5181);
or OR4 (N7820, N7805, N6254, N4938, N1756);
and AND4 (N7821, N7800, N4072, N4513, N1092);
xor XOR2 (N7822, N7812, N2457);
xor XOR2 (N7823, N7822, N2113);
and AND3 (N7824, N7823, N3814, N5855);
not NOT1 (N7825, N7810);
and AND2 (N7826, N7820, N6709);
and AND4 (N7827, N7821, N824, N6166, N6308);
nor NOR4 (N7828, N7815, N5784, N5427, N4769);
xor XOR2 (N7829, N7818, N94);
not NOT1 (N7830, N7816);
nand NAND2 (N7831, N7824, N1626);
or OR4 (N7832, N7826, N5193, N1923, N1202);
and AND4 (N7833, N7828, N5304, N6180, N4945);
nand NAND2 (N7834, N7825, N3770);
nand NAND4 (N7835, N7817, N7250, N7339, N26);
nor NOR2 (N7836, N7809, N3851);
and AND2 (N7837, N7830, N3007);
buf BUF1 (N7838, N7827);
not NOT1 (N7839, N7829);
buf BUF1 (N7840, N7835);
not NOT1 (N7841, N7840);
xor XOR2 (N7842, N7841, N7075);
nor NOR2 (N7843, N7836, N2402);
or OR4 (N7844, N7838, N5633, N6997, N6845);
not NOT1 (N7845, N7834);
nand NAND3 (N7846, N7843, N4367, N1087);
and AND3 (N7847, N7846, N3104, N3642);
nand NAND2 (N7848, N7839, N6346);
nand NAND3 (N7849, N7831, N2644, N3764);
xor XOR2 (N7850, N7844, N7222);
or OR2 (N7851, N7837, N7129);
xor XOR2 (N7852, N7850, N5396);
nand NAND3 (N7853, N7847, N3676, N7115);
xor XOR2 (N7854, N7852, N5990);
and AND2 (N7855, N7845, N2900);
and AND4 (N7856, N7833, N1018, N4359, N7252);
nand NAND3 (N7857, N7848, N4906, N2976);
buf BUF1 (N7858, N7855);
nand NAND2 (N7859, N7832, N4579);
and AND2 (N7860, N7856, N6919);
and AND4 (N7861, N7849, N1376, N5010, N891);
xor XOR2 (N7862, N7858, N3249);
nand NAND2 (N7863, N7862, N206);
buf BUF1 (N7864, N7860);
buf BUF1 (N7865, N7842);
and AND2 (N7866, N7859, N2108);
not NOT1 (N7867, N7866);
and AND2 (N7868, N7863, N6439);
and AND4 (N7869, N7861, N7508, N122, N4498);
and AND3 (N7870, N7851, N4911, N4211);
not NOT1 (N7871, N7869);
buf BUF1 (N7872, N7865);
xor XOR2 (N7873, N7864, N6616);
xor XOR2 (N7874, N7867, N4007);
not NOT1 (N7875, N7854);
nand NAND2 (N7876, N7873, N3746);
xor XOR2 (N7877, N7872, N2766);
buf BUF1 (N7878, N7853);
buf BUF1 (N7879, N7868);
nand NAND4 (N7880, N7819, N5738, N1111, N4862);
xor XOR2 (N7881, N7874, N7153);
or OR3 (N7882, N7871, N3255, N6441);
xor XOR2 (N7883, N7881, N1546);
or OR2 (N7884, N7876, N7479);
nand NAND3 (N7885, N7878, N832, N3938);
or OR4 (N7886, N7877, N1766, N3446, N681);
or OR4 (N7887, N7879, N2209, N3216, N1152);
not NOT1 (N7888, N7880);
buf BUF1 (N7889, N7875);
and AND2 (N7890, N7887, N1717);
buf BUF1 (N7891, N7886);
buf BUF1 (N7892, N7884);
or OR4 (N7893, N7890, N6662, N423, N396);
not NOT1 (N7894, N7893);
buf BUF1 (N7895, N7883);
and AND4 (N7896, N7894, N2930, N2824, N6225);
nor NOR2 (N7897, N7857, N5127);
xor XOR2 (N7898, N7885, N3366);
xor XOR2 (N7899, N7896, N5936);
not NOT1 (N7900, N7898);
not NOT1 (N7901, N7888);
xor XOR2 (N7902, N7892, N1619);
xor XOR2 (N7903, N7870, N4281);
not NOT1 (N7904, N7903);
and AND4 (N7905, N7902, N2756, N462, N195);
or OR2 (N7906, N7891, N4552);
not NOT1 (N7907, N7889);
nor NOR4 (N7908, N7899, N5671, N7010, N2171);
buf BUF1 (N7909, N7901);
and AND2 (N7910, N7909, N3715);
xor XOR2 (N7911, N7904, N982);
nand NAND3 (N7912, N7897, N172, N3958);
not NOT1 (N7913, N7882);
nor NOR3 (N7914, N7895, N1486, N7491);
xor XOR2 (N7915, N7910, N3074);
xor XOR2 (N7916, N7907, N5900);
or OR2 (N7917, N7912, N6404);
not NOT1 (N7918, N7915);
buf BUF1 (N7919, N7900);
and AND3 (N7920, N7916, N5418, N5904);
nor NOR3 (N7921, N7920, N6199, N3753);
xor XOR2 (N7922, N7905, N5612);
nor NOR3 (N7923, N7917, N2149, N7671);
not NOT1 (N7924, N7921);
xor XOR2 (N7925, N7924, N6422);
and AND2 (N7926, N7918, N4387);
buf BUF1 (N7927, N7911);
nor NOR2 (N7928, N7925, N6884);
nor NOR2 (N7929, N7914, N349);
or OR3 (N7930, N7906, N4585, N4093);
and AND2 (N7931, N7930, N5121);
and AND3 (N7932, N7923, N5757, N4338);
or OR3 (N7933, N7932, N769, N7621);
nand NAND3 (N7934, N7922, N6281, N768);
and AND4 (N7935, N7929, N37, N4922, N3854);
or OR4 (N7936, N7927, N6799, N463, N2724);
or OR2 (N7937, N7928, N5203);
buf BUF1 (N7938, N7908);
nor NOR4 (N7939, N7933, N3811, N2146, N1312);
nor NOR4 (N7940, N7926, N7865, N1133, N3759);
buf BUF1 (N7941, N7934);
buf BUF1 (N7942, N7931);
nand NAND4 (N7943, N7939, N2379, N2657, N1236);
or OR4 (N7944, N7937, N411, N3898, N5282);
not NOT1 (N7945, N7943);
nor NOR4 (N7946, N7940, N6679, N4649, N5705);
or OR3 (N7947, N7938, N7005, N4314);
or OR4 (N7948, N7913, N5604, N3416, N1134);
or OR3 (N7949, N7947, N3049, N5885);
or OR3 (N7950, N7949, N376, N1436);
xor XOR2 (N7951, N7942, N1667);
and AND2 (N7952, N7936, N7097);
xor XOR2 (N7953, N7935, N4836);
and AND2 (N7954, N7953, N4114);
not NOT1 (N7955, N7954);
and AND4 (N7956, N7950, N6895, N4402, N2063);
buf BUF1 (N7957, N7951);
and AND4 (N7958, N7955, N7954, N1850, N944);
and AND2 (N7959, N7946, N7557);
buf BUF1 (N7960, N7952);
buf BUF1 (N7961, N7944);
nor NOR4 (N7962, N7941, N6239, N415, N5056);
nor NOR2 (N7963, N7960, N2677);
or OR3 (N7964, N7958, N6618, N1000);
nor NOR2 (N7965, N7959, N5943);
buf BUF1 (N7966, N7945);
buf BUF1 (N7967, N7966);
buf BUF1 (N7968, N7961);
nand NAND4 (N7969, N7919, N3488, N5295, N5077);
nand NAND2 (N7970, N7968, N216);
not NOT1 (N7971, N7965);
nor NOR2 (N7972, N7948, N7808);
nand NAND2 (N7973, N7963, N5345);
or OR4 (N7974, N7972, N4350, N1492, N6779);
nand NAND2 (N7975, N7964, N5603);
nand NAND4 (N7976, N7974, N7661, N1800, N7498);
xor XOR2 (N7977, N7962, N4512);
nor NOR2 (N7978, N7973, N4891);
and AND3 (N7979, N7970, N135, N1785);
nand NAND2 (N7980, N7976, N1982);
nand NAND4 (N7981, N7957, N5160, N5619, N4980);
buf BUF1 (N7982, N7981);
and AND2 (N7983, N7956, N5915);
nor NOR2 (N7984, N7971, N6672);
nand NAND4 (N7985, N7980, N3923, N4977, N3877);
or OR2 (N7986, N7979, N2299);
nor NOR4 (N7987, N7975, N6530, N7000, N2797);
buf BUF1 (N7988, N7983);
buf BUF1 (N7989, N7977);
xor XOR2 (N7990, N7985, N1125);
not NOT1 (N7991, N7969);
nand NAND3 (N7992, N7967, N5701, N7855);
nor NOR2 (N7993, N7989, N788);
or OR4 (N7994, N7986, N6065, N7301, N5121);
nor NOR4 (N7995, N7994, N4320, N7661, N6644);
nand NAND4 (N7996, N7990, N5415, N6141, N68);
xor XOR2 (N7997, N7992, N2098);
xor XOR2 (N7998, N7995, N5409);
and AND3 (N7999, N7996, N3046, N1132);
and AND4 (N8000, N7982, N1061, N4245, N6913);
xor XOR2 (N8001, N7998, N1301);
or OR2 (N8002, N7997, N5514);
xor XOR2 (N8003, N8001, N3955);
nand NAND4 (N8004, N7993, N3182, N4131, N5596);
nor NOR2 (N8005, N8000, N4166);
and AND3 (N8006, N8003, N3599, N5884);
or OR2 (N8007, N8005, N1300);
buf BUF1 (N8008, N8002);
nand NAND2 (N8009, N7984, N488);
xor XOR2 (N8010, N8007, N3883);
or OR3 (N8011, N8010, N2863, N7242);
buf BUF1 (N8012, N8006);
and AND3 (N8013, N8012, N788, N647);
buf BUF1 (N8014, N8008);
xor XOR2 (N8015, N8011, N1144);
nor NOR4 (N8016, N7991, N5655, N1862, N1160);
buf BUF1 (N8017, N7988);
and AND2 (N8018, N8014, N7714);
xor XOR2 (N8019, N7978, N3158);
nor NOR4 (N8020, N8015, N5404, N7301, N4623);
nor NOR4 (N8021, N7987, N5608, N7671, N671);
xor XOR2 (N8022, N8013, N3864);
not NOT1 (N8023, N8022);
nor NOR3 (N8024, N7999, N6805, N511);
xor XOR2 (N8025, N8018, N934);
not NOT1 (N8026, N8020);
buf BUF1 (N8027, N8021);
nor NOR3 (N8028, N8017, N2345, N1599);
not NOT1 (N8029, N8019);
nand NAND2 (N8030, N8027, N3354);
not NOT1 (N8031, N8023);
nand NAND3 (N8032, N8025, N6258, N228);
and AND2 (N8033, N8029, N154);
or OR2 (N8034, N8033, N706);
nor NOR2 (N8035, N8009, N946);
and AND4 (N8036, N8032, N820, N1956, N4859);
not NOT1 (N8037, N8024);
not NOT1 (N8038, N8037);
nor NOR4 (N8039, N8030, N5703, N3756, N1717);
nand NAND3 (N8040, N8004, N2115, N174);
and AND2 (N8041, N8034, N7463);
xor XOR2 (N8042, N8038, N6488);
nor NOR3 (N8043, N8028, N363, N6410);
nor NOR4 (N8044, N8035, N923, N6094, N7323);
nor NOR4 (N8045, N8044, N6172, N3730, N7139);
nor NOR3 (N8046, N8026, N7636, N5399);
nor NOR2 (N8047, N8045, N6131);
not NOT1 (N8048, N8046);
nand NAND2 (N8049, N8043, N6393);
nor NOR2 (N8050, N8036, N7773);
and AND3 (N8051, N8039, N2771, N3891);
nand NAND3 (N8052, N8016, N3909, N7150);
nor NOR3 (N8053, N8052, N2872, N1709);
or OR3 (N8054, N8047, N6500, N6733);
xor XOR2 (N8055, N8054, N4519);
buf BUF1 (N8056, N8040);
not NOT1 (N8057, N8031);
or OR4 (N8058, N8048, N2936, N738, N1248);
nand NAND2 (N8059, N8041, N7609);
nor NOR2 (N8060, N8057, N6476);
nand NAND3 (N8061, N8050, N2128, N1920);
nor NOR3 (N8062, N8053, N4028, N6964);
buf BUF1 (N8063, N8060);
and AND3 (N8064, N8062, N4177, N459);
xor XOR2 (N8065, N8055, N2274);
not NOT1 (N8066, N8065);
not NOT1 (N8067, N8061);
nor NOR2 (N8068, N8042, N3729);
not NOT1 (N8069, N8051);
not NOT1 (N8070, N8059);
or OR4 (N8071, N8056, N1640, N2118, N3653);
xor XOR2 (N8072, N8069, N3303);
nand NAND4 (N8073, N8063, N2602, N2743, N5704);
nor NOR4 (N8074, N8049, N1712, N5216, N6249);
and AND2 (N8075, N8072, N3749);
nand NAND2 (N8076, N8073, N4702);
and AND3 (N8077, N8066, N5137, N5835);
nand NAND3 (N8078, N8068, N332, N4740);
nand NAND4 (N8079, N8074, N601, N3639, N2326);
nor NOR2 (N8080, N8077, N2564);
not NOT1 (N8081, N8058);
nor NOR4 (N8082, N8070, N4769, N4892, N320);
xor XOR2 (N8083, N8078, N7247);
nand NAND2 (N8084, N8071, N657);
and AND3 (N8085, N8075, N4309, N173);
buf BUF1 (N8086, N8081);
buf BUF1 (N8087, N8076);
or OR3 (N8088, N8082, N608, N5124);
nand NAND3 (N8089, N8079, N2818, N6092);
not NOT1 (N8090, N8067);
not NOT1 (N8091, N8083);
and AND2 (N8092, N8085, N2654);
or OR3 (N8093, N8087, N380, N5936);
xor XOR2 (N8094, N8093, N6838);
and AND2 (N8095, N8080, N7171);
nand NAND4 (N8096, N8086, N3028, N7719, N7237);
or OR2 (N8097, N8096, N6756);
xor XOR2 (N8098, N8064, N3146);
or OR2 (N8099, N8092, N1177);
not NOT1 (N8100, N8098);
nand NAND2 (N8101, N8095, N3132);
and AND2 (N8102, N8094, N5237);
buf BUF1 (N8103, N8101);
nor NOR4 (N8104, N8091, N18, N1326, N2886);
nand NAND2 (N8105, N8103, N1660);
buf BUF1 (N8106, N8090);
not NOT1 (N8107, N8097);
and AND2 (N8108, N8100, N6360);
nand NAND3 (N8109, N8108, N7957, N461);
or OR2 (N8110, N8106, N855);
nand NAND2 (N8111, N8105, N2023);
and AND2 (N8112, N8099, N6691);
or OR2 (N8113, N8088, N7381);
nand NAND4 (N8114, N8089, N2867, N4086, N1041);
xor XOR2 (N8115, N8113, N3812);
and AND2 (N8116, N8114, N7744);
and AND2 (N8117, N8104, N5740);
not NOT1 (N8118, N8107);
nand NAND4 (N8119, N8084, N3719, N974, N2875);
or OR4 (N8120, N8112, N4853, N1925, N1528);
and AND4 (N8121, N8109, N6379, N1269, N6186);
nor NOR2 (N8122, N8115, N7527);
nand NAND2 (N8123, N8117, N1674);
xor XOR2 (N8124, N8121, N2836);
nand NAND3 (N8125, N8102, N3630, N7483);
and AND4 (N8126, N8111, N5640, N204, N2508);
and AND2 (N8127, N8123, N3544);
buf BUF1 (N8128, N8110);
or OR2 (N8129, N8126, N4638);
and AND4 (N8130, N8122, N2065, N6606, N1528);
nand NAND2 (N8131, N8119, N7596);
nor NOR4 (N8132, N8129, N2133, N8027, N3955);
and AND3 (N8133, N8132, N2294, N7774);
nand NAND4 (N8134, N8116, N1992, N115, N665);
buf BUF1 (N8135, N8134);
not NOT1 (N8136, N8118);
or OR3 (N8137, N8120, N6246, N6079);
nand NAND3 (N8138, N8133, N3608, N2551);
or OR4 (N8139, N8137, N3261, N4019, N2434);
buf BUF1 (N8140, N8125);
or OR3 (N8141, N8124, N1354, N3095);
nor NOR3 (N8142, N8135, N5594, N4737);
nand NAND2 (N8143, N8136, N543);
nor NOR2 (N8144, N8142, N4744);
or OR3 (N8145, N8130, N5016, N113);
not NOT1 (N8146, N8128);
buf BUF1 (N8147, N8131);
xor XOR2 (N8148, N8140, N2054);
nor NOR2 (N8149, N8147, N3092);
or OR3 (N8150, N8138, N2962, N6352);
buf BUF1 (N8151, N8150);
nor NOR2 (N8152, N8143, N3198);
xor XOR2 (N8153, N8139, N262);
xor XOR2 (N8154, N8151, N5311);
not NOT1 (N8155, N8141);
nor NOR4 (N8156, N8154, N5131, N5669, N5048);
buf BUF1 (N8157, N8127);
buf BUF1 (N8158, N8153);
or OR3 (N8159, N8148, N1947, N1764);
not NOT1 (N8160, N8159);
buf BUF1 (N8161, N8149);
nand NAND3 (N8162, N8158, N1795, N4619);
buf BUF1 (N8163, N8144);
xor XOR2 (N8164, N8152, N953);
nor NOR2 (N8165, N8157, N6000);
xor XOR2 (N8166, N8155, N6416);
buf BUF1 (N8167, N8146);
or OR2 (N8168, N8161, N1618);
xor XOR2 (N8169, N8165, N62);
nand NAND4 (N8170, N8145, N6739, N3169, N2305);
buf BUF1 (N8171, N8162);
buf BUF1 (N8172, N8169);
or OR4 (N8173, N8168, N1096, N3171, N5575);
nor NOR2 (N8174, N8160, N7965);
and AND3 (N8175, N8170, N14, N6475);
not NOT1 (N8176, N8173);
or OR4 (N8177, N8164, N3322, N7434, N7673);
nor NOR4 (N8178, N8167, N4106, N3447, N7098);
not NOT1 (N8179, N8156);
buf BUF1 (N8180, N8166);
and AND2 (N8181, N8172, N3488);
buf BUF1 (N8182, N8181);
or OR4 (N8183, N8175, N2762, N5319, N5607);
and AND4 (N8184, N8174, N2673, N7287, N2633);
buf BUF1 (N8185, N8183);
or OR3 (N8186, N8177, N3125, N3708);
buf BUF1 (N8187, N8182);
nand NAND3 (N8188, N8187, N8055, N8123);
xor XOR2 (N8189, N8180, N5559);
and AND4 (N8190, N8189, N2493, N1720, N5271);
nand NAND4 (N8191, N8171, N3613, N14, N113);
or OR2 (N8192, N8176, N5956);
or OR2 (N8193, N8163, N5707);
or OR3 (N8194, N8193, N5106, N1881);
and AND3 (N8195, N8186, N23, N5837);
not NOT1 (N8196, N8185);
and AND4 (N8197, N8191, N6567, N1602, N122);
and AND4 (N8198, N8178, N4264, N2889, N8094);
buf BUF1 (N8199, N8198);
and AND2 (N8200, N8179, N5185);
buf BUF1 (N8201, N8199);
nor NOR3 (N8202, N8201, N41, N4670);
buf BUF1 (N8203, N8192);
or OR3 (N8204, N8194, N3606, N8165);
nand NAND3 (N8205, N8196, N6626, N177);
xor XOR2 (N8206, N8197, N1833);
xor XOR2 (N8207, N8202, N1058);
buf BUF1 (N8208, N8206);
nor NOR2 (N8209, N8207, N8186);
nand NAND4 (N8210, N8208, N4946, N3918, N7440);
not NOT1 (N8211, N8203);
nand NAND2 (N8212, N8200, N6952);
buf BUF1 (N8213, N8205);
nor NOR4 (N8214, N8210, N6955, N2576, N5149);
nand NAND4 (N8215, N8212, N6884, N3647, N819);
xor XOR2 (N8216, N8190, N3747);
not NOT1 (N8217, N8204);
nand NAND3 (N8218, N8188, N5404, N2187);
nor NOR3 (N8219, N8209, N7208, N4279);
buf BUF1 (N8220, N8211);
nand NAND3 (N8221, N8217, N5073, N1846);
xor XOR2 (N8222, N8213, N334);
nor NOR4 (N8223, N8222, N476, N4372, N8023);
not NOT1 (N8224, N8221);
buf BUF1 (N8225, N8214);
not NOT1 (N8226, N8215);
not NOT1 (N8227, N8225);
buf BUF1 (N8228, N8216);
and AND4 (N8229, N8219, N2076, N1759, N4058);
nand NAND3 (N8230, N8229, N5623, N5285);
or OR4 (N8231, N8220, N1988, N96, N3596);
and AND3 (N8232, N8184, N4116, N1313);
or OR4 (N8233, N8228, N4725, N4796, N3644);
and AND4 (N8234, N8224, N6443, N2256, N1395);
nand NAND4 (N8235, N8230, N1781, N7948, N8044);
nand NAND4 (N8236, N8234, N5914, N6274, N6459);
nor NOR2 (N8237, N8235, N452);
not NOT1 (N8238, N8223);
nor NOR4 (N8239, N8227, N4632, N2718, N1157);
not NOT1 (N8240, N8232);
not NOT1 (N8241, N8237);
or OR2 (N8242, N8236, N2930);
not NOT1 (N8243, N8241);
and AND4 (N8244, N8231, N1742, N2289, N3279);
nor NOR4 (N8245, N8242, N4721, N1408, N2788);
xor XOR2 (N8246, N8243, N997);
xor XOR2 (N8247, N8240, N7106);
not NOT1 (N8248, N8195);
or OR4 (N8249, N8247, N6846, N7207, N86);
nand NAND3 (N8250, N8239, N2603, N2430);
nand NAND2 (N8251, N8250, N1025);
nand NAND2 (N8252, N8245, N2602);
nor NOR4 (N8253, N8218, N3733, N3779, N7330);
buf BUF1 (N8254, N8252);
nand NAND2 (N8255, N8226, N1299);
nand NAND2 (N8256, N8253, N1022);
buf BUF1 (N8257, N8256);
buf BUF1 (N8258, N8255);
not NOT1 (N8259, N8249);
or OR2 (N8260, N8257, N6841);
and AND2 (N8261, N8260, N2098);
nor NOR3 (N8262, N8254, N1918, N6945);
nand NAND2 (N8263, N8233, N8037);
and AND2 (N8264, N8263, N2078);
buf BUF1 (N8265, N8248);
nor NOR2 (N8266, N8244, N6911);
xor XOR2 (N8267, N8266, N7204);
xor XOR2 (N8268, N8265, N2585);
nand NAND3 (N8269, N8267, N7929, N1739);
or OR3 (N8270, N8262, N484, N6877);
not NOT1 (N8271, N8261);
nand NAND4 (N8272, N8246, N2001, N5909, N2114);
buf BUF1 (N8273, N8259);
nor NOR2 (N8274, N8238, N3486);
xor XOR2 (N8275, N8269, N603);
xor XOR2 (N8276, N8258, N6258);
xor XOR2 (N8277, N8270, N5939);
nor NOR3 (N8278, N8272, N1580, N409);
buf BUF1 (N8279, N8251);
nand NAND2 (N8280, N8268, N7970);
or OR4 (N8281, N8280, N281, N2856, N3169);
not NOT1 (N8282, N8264);
nand NAND3 (N8283, N8276, N6810, N5092);
buf BUF1 (N8284, N8273);
nor NOR2 (N8285, N8284, N494);
not NOT1 (N8286, N8274);
nand NAND4 (N8287, N8279, N1053, N190, N3860);
or OR4 (N8288, N8277, N6681, N7022, N3516);
xor XOR2 (N8289, N8286, N213);
nor NOR4 (N8290, N8288, N6666, N2661, N1068);
and AND2 (N8291, N8285, N4249);
buf BUF1 (N8292, N8271);
and AND4 (N8293, N8287, N7327, N2263, N2);
and AND3 (N8294, N8278, N2912, N5050);
nand NAND3 (N8295, N8291, N2750, N5399);
buf BUF1 (N8296, N8283);
nand NAND3 (N8297, N8296, N6764, N614);
xor XOR2 (N8298, N8295, N7466);
not NOT1 (N8299, N8298);
not NOT1 (N8300, N8281);
nand NAND3 (N8301, N8299, N4941, N3337);
and AND2 (N8302, N8300, N8079);
nand NAND3 (N8303, N8293, N5436, N4324);
not NOT1 (N8304, N8303);
or OR3 (N8305, N8282, N1126, N6325);
buf BUF1 (N8306, N8275);
buf BUF1 (N8307, N8292);
xor XOR2 (N8308, N8290, N4492);
nand NAND3 (N8309, N8306, N2401, N7340);
nor NOR4 (N8310, N8302, N2179, N7451, N2482);
buf BUF1 (N8311, N8297);
not NOT1 (N8312, N8308);
buf BUF1 (N8313, N8304);
not NOT1 (N8314, N8312);
nor NOR3 (N8315, N8313, N5404, N8040);
or OR4 (N8316, N8310, N540, N6811, N5918);
nor NOR3 (N8317, N8311, N7051, N85);
buf BUF1 (N8318, N8289);
xor XOR2 (N8319, N8301, N3169);
nand NAND3 (N8320, N8318, N7807, N868);
and AND2 (N8321, N8316, N6421);
not NOT1 (N8322, N8314);
buf BUF1 (N8323, N8307);
and AND4 (N8324, N8305, N4751, N3208, N4410);
nand NAND2 (N8325, N8309, N1652);
buf BUF1 (N8326, N8317);
and AND3 (N8327, N8294, N2625, N2681);
or OR4 (N8328, N8320, N4096, N5674, N704);
or OR3 (N8329, N8326, N4024, N2316);
nor NOR3 (N8330, N8321, N5084, N7223);
nand NAND3 (N8331, N8319, N211, N1813);
nand NAND2 (N8332, N8328, N4699);
not NOT1 (N8333, N8332);
xor XOR2 (N8334, N8325, N7876);
or OR3 (N8335, N8333, N2366, N3157);
nand NAND2 (N8336, N8330, N8272);
and AND2 (N8337, N8331, N738);
xor XOR2 (N8338, N8337, N6745);
xor XOR2 (N8339, N8338, N5688);
nand NAND2 (N8340, N8339, N7609);
not NOT1 (N8341, N8336);
or OR2 (N8342, N8322, N7993);
not NOT1 (N8343, N8342);
not NOT1 (N8344, N8323);
and AND4 (N8345, N8334, N8325, N3698, N4669);
not NOT1 (N8346, N8327);
or OR4 (N8347, N8346, N3478, N1703, N6587);
nand NAND3 (N8348, N8340, N6677, N2903);
nand NAND4 (N8349, N8344, N1712, N8176, N5878);
or OR4 (N8350, N8324, N2779, N4267, N6913);
and AND3 (N8351, N8347, N5796, N2793);
nor NOR2 (N8352, N8350, N1815);
nor NOR4 (N8353, N8349, N6298, N8105, N899);
or OR4 (N8354, N8329, N3447, N7324, N5923);
nand NAND4 (N8355, N8315, N265, N2963, N1990);
nor NOR2 (N8356, N8352, N6142);
nand NAND3 (N8357, N8355, N4221, N6615);
and AND4 (N8358, N8357, N241, N5577, N7883);
buf BUF1 (N8359, N8358);
nand NAND2 (N8360, N8335, N7143);
buf BUF1 (N8361, N8345);
buf BUF1 (N8362, N8354);
buf BUF1 (N8363, N8353);
xor XOR2 (N8364, N8343, N3229);
or OR3 (N8365, N8363, N1926, N1139);
nand NAND3 (N8366, N8364, N1628, N6098);
nand NAND2 (N8367, N8365, N6609);
nor NOR3 (N8368, N8359, N471, N1442);
not NOT1 (N8369, N8351);
nor NOR4 (N8370, N8362, N478, N2066, N2510);
nor NOR4 (N8371, N8361, N924, N2329, N3451);
nor NOR2 (N8372, N8356, N1760);
buf BUF1 (N8373, N8368);
buf BUF1 (N8374, N8366);
buf BUF1 (N8375, N8371);
or OR2 (N8376, N8374, N8193);
not NOT1 (N8377, N8341);
and AND3 (N8378, N8369, N1482, N7107);
not NOT1 (N8379, N8373);
nor NOR2 (N8380, N8372, N4047);
xor XOR2 (N8381, N8360, N4850);
nand NAND4 (N8382, N8377, N3752, N1655, N3416);
not NOT1 (N8383, N8375);
nor NOR3 (N8384, N8370, N3115, N3106);
xor XOR2 (N8385, N8348, N4075);
not NOT1 (N8386, N8385);
and AND3 (N8387, N8382, N6090, N4372);
and AND3 (N8388, N8384, N8105, N5308);
nor NOR2 (N8389, N8379, N2478);
xor XOR2 (N8390, N8388, N5502);
not NOT1 (N8391, N8383);
or OR4 (N8392, N8386, N3579, N3440, N4530);
or OR2 (N8393, N8392, N2945);
xor XOR2 (N8394, N8378, N4224);
not NOT1 (N8395, N8376);
buf BUF1 (N8396, N8380);
and AND2 (N8397, N8381, N2576);
nor NOR4 (N8398, N8387, N1277, N4029, N6225);
buf BUF1 (N8399, N8390);
not NOT1 (N8400, N8399);
buf BUF1 (N8401, N8395);
not NOT1 (N8402, N8401);
not NOT1 (N8403, N8398);
and AND2 (N8404, N8367, N3154);
nand NAND4 (N8405, N8404, N810, N3548, N4007);
nor NOR2 (N8406, N8394, N7085);
nand NAND3 (N8407, N8393, N1282, N533);
and AND4 (N8408, N8400, N311, N4440, N5396);
nor NOR4 (N8409, N8406, N1703, N1862, N529);
not NOT1 (N8410, N8407);
nor NOR2 (N8411, N8396, N5737);
and AND4 (N8412, N8411, N6287, N959, N4353);
or OR3 (N8413, N8412, N3061, N7876);
nor NOR2 (N8414, N8405, N7587);
and AND3 (N8415, N8408, N3825, N5153);
and AND3 (N8416, N8409, N5666, N8356);
not NOT1 (N8417, N8391);
nor NOR3 (N8418, N8402, N8305, N541);
nand NAND2 (N8419, N8403, N4583);
xor XOR2 (N8420, N8417, N4847);
xor XOR2 (N8421, N8397, N6043);
nor NOR4 (N8422, N8389, N4927, N578, N6621);
xor XOR2 (N8423, N8418, N8395);
or OR3 (N8424, N8419, N3879, N4818);
nor NOR4 (N8425, N8415, N2249, N7463, N7624);
xor XOR2 (N8426, N8414, N2090);
buf BUF1 (N8427, N8426);
or OR3 (N8428, N8425, N6089, N6541);
not NOT1 (N8429, N8420);
nand NAND3 (N8430, N8421, N6900, N7643);
buf BUF1 (N8431, N8428);
xor XOR2 (N8432, N8427, N2195);
or OR2 (N8433, N8429, N4241);
nor NOR4 (N8434, N8431, N7399, N4895, N3772);
nand NAND2 (N8435, N8432, N1062);
and AND2 (N8436, N8410, N5869);
and AND4 (N8437, N8436, N4204, N5674, N4413);
not NOT1 (N8438, N8437);
or OR3 (N8439, N8430, N7128, N3492);
nand NAND2 (N8440, N8416, N7667);
xor XOR2 (N8441, N8438, N2496);
nand NAND2 (N8442, N8424, N1211);
not NOT1 (N8443, N8442);
xor XOR2 (N8444, N8434, N5102);
and AND3 (N8445, N8413, N3086, N2944);
or OR3 (N8446, N8435, N8434, N1221);
buf BUF1 (N8447, N8433);
not NOT1 (N8448, N8423);
not NOT1 (N8449, N8439);
or OR4 (N8450, N8447, N3236, N6442, N68);
nand NAND3 (N8451, N8450, N3472, N6694);
xor XOR2 (N8452, N8451, N3404);
nor NOR2 (N8453, N8441, N4264);
not NOT1 (N8454, N8446);
or OR2 (N8455, N8452, N2275);
nand NAND4 (N8456, N8454, N3134, N6319, N5043);
or OR4 (N8457, N8453, N3462, N4593, N7226);
nand NAND2 (N8458, N8422, N8299);
and AND4 (N8459, N8458, N4942, N4746, N5454);
or OR2 (N8460, N8440, N1389);
and AND4 (N8461, N8444, N4120, N4045, N3561);
nor NOR3 (N8462, N8455, N885, N7233);
nand NAND2 (N8463, N8457, N5999);
and AND2 (N8464, N8459, N4772);
nor NOR3 (N8465, N8460, N7214, N5850);
nor NOR2 (N8466, N8443, N7721);
nor NOR3 (N8467, N8463, N7463, N6704);
nand NAND3 (N8468, N8448, N6133, N2996);
nor NOR2 (N8469, N8467, N1735);
nor NOR4 (N8470, N8468, N146, N2617, N1675);
or OR3 (N8471, N8456, N4032, N8057);
and AND4 (N8472, N8465, N6802, N4395, N4561);
or OR4 (N8473, N8462, N2068, N2268, N5925);
and AND4 (N8474, N8469, N2645, N7269, N7982);
nand NAND2 (N8475, N8464, N1386);
nand NAND4 (N8476, N8474, N5410, N4403, N6805);
not NOT1 (N8477, N8475);
nand NAND3 (N8478, N8449, N7047, N1652);
nand NAND4 (N8479, N8471, N3680, N2531, N7341);
nor NOR2 (N8480, N8470, N2498);
not NOT1 (N8481, N8480);
buf BUF1 (N8482, N8472);
not NOT1 (N8483, N8478);
xor XOR2 (N8484, N8473, N7251);
buf BUF1 (N8485, N8481);
buf BUF1 (N8486, N8484);
nand NAND3 (N8487, N8476, N940, N1421);
xor XOR2 (N8488, N8466, N284);
nand NAND2 (N8489, N8487, N5678);
buf BUF1 (N8490, N8486);
or OR3 (N8491, N8461, N7393, N3621);
not NOT1 (N8492, N8477);
nor NOR3 (N8493, N8490, N2450, N7348);
buf BUF1 (N8494, N8483);
nor NOR4 (N8495, N8489, N2627, N377, N6920);
and AND3 (N8496, N8495, N3131, N5496);
nand NAND4 (N8497, N8479, N447, N4609, N5362);
xor XOR2 (N8498, N8497, N7006);
nor NOR4 (N8499, N8494, N1388, N3268, N1117);
nand NAND4 (N8500, N8491, N8305, N1940, N190);
buf BUF1 (N8501, N8498);
or OR4 (N8502, N8492, N120, N351, N7580);
and AND3 (N8503, N8502, N2263, N2974);
buf BUF1 (N8504, N8503);
xor XOR2 (N8505, N8485, N4944);
xor XOR2 (N8506, N8482, N1062);
nand NAND4 (N8507, N8488, N5035, N3064, N7760);
and AND4 (N8508, N8507, N7877, N1306, N1261);
or OR2 (N8509, N8493, N1062);
nor NOR3 (N8510, N8504, N347, N7757);
and AND3 (N8511, N8505, N1358, N244);
or OR3 (N8512, N8499, N7999, N5703);
or OR3 (N8513, N8506, N8242, N7098);
and AND3 (N8514, N8512, N6034, N2839);
nor NOR2 (N8515, N8500, N4257);
xor XOR2 (N8516, N8510, N155);
buf BUF1 (N8517, N8501);
nand NAND2 (N8518, N8513, N5186);
xor XOR2 (N8519, N8511, N2776);
xor XOR2 (N8520, N8514, N6872);
not NOT1 (N8521, N8509);
nor NOR4 (N8522, N8508, N8130, N2145, N3810);
not NOT1 (N8523, N8515);
or OR4 (N8524, N8516, N4879, N772, N4699);
buf BUF1 (N8525, N8520);
not NOT1 (N8526, N8525);
nand NAND3 (N8527, N8526, N2121, N3352);
nor NOR3 (N8528, N8524, N5919, N8456);
nor NOR3 (N8529, N8527, N518, N438);
and AND4 (N8530, N8521, N1644, N6140, N7157);
and AND2 (N8531, N8445, N4378);
nand NAND3 (N8532, N8519, N4906, N963);
and AND4 (N8533, N8530, N1625, N1260, N3980);
nor NOR3 (N8534, N8532, N3596, N6751);
nand NAND2 (N8535, N8517, N8534);
or OR4 (N8536, N1387, N6904, N4447, N3617);
nand NAND3 (N8537, N8528, N33, N3982);
nor NOR3 (N8538, N8518, N4759, N422);
xor XOR2 (N8539, N8522, N6949);
and AND2 (N8540, N8529, N2204);
buf BUF1 (N8541, N8540);
xor XOR2 (N8542, N8531, N1550);
nand NAND2 (N8543, N8542, N3456);
nor NOR3 (N8544, N8538, N6531, N5977);
xor XOR2 (N8545, N8541, N3012);
not NOT1 (N8546, N8496);
or OR4 (N8547, N8544, N8323, N4208, N5334);
xor XOR2 (N8548, N8546, N6490);
or OR4 (N8549, N8533, N658, N5806, N6947);
xor XOR2 (N8550, N8549, N1438);
or OR2 (N8551, N8539, N3736);
nand NAND2 (N8552, N8551, N3350);
not NOT1 (N8553, N8552);
and AND3 (N8554, N8543, N4103, N2525);
and AND3 (N8555, N8523, N90, N7831);
nor NOR2 (N8556, N8537, N7726);
buf BUF1 (N8557, N8550);
nor NOR4 (N8558, N8548, N6008, N201, N7987);
buf BUF1 (N8559, N8535);
buf BUF1 (N8560, N8555);
not NOT1 (N8561, N8554);
and AND3 (N8562, N8553, N7421, N3794);
not NOT1 (N8563, N8562);
and AND2 (N8564, N8558, N6200);
xor XOR2 (N8565, N8560, N4812);
not NOT1 (N8566, N8565);
nand NAND4 (N8567, N8557, N6379, N5618, N5101);
nand NAND2 (N8568, N8566, N3321);
xor XOR2 (N8569, N8547, N4969);
and AND3 (N8570, N8561, N6476, N2230);
buf BUF1 (N8571, N8536);
and AND3 (N8572, N8564, N6173, N899);
xor XOR2 (N8573, N8563, N607);
nand NAND4 (N8574, N8572, N3345, N4834, N1662);
and AND4 (N8575, N8545, N5811, N3954, N4529);
xor XOR2 (N8576, N8567, N1718);
buf BUF1 (N8577, N8559);
buf BUF1 (N8578, N8575);
or OR4 (N8579, N8556, N2429, N1864, N2552);
xor XOR2 (N8580, N8570, N7437);
buf BUF1 (N8581, N8574);
not NOT1 (N8582, N8581);
and AND3 (N8583, N8576, N7062, N5797);
not NOT1 (N8584, N8583);
and AND3 (N8585, N8584, N4820, N3658);
or OR3 (N8586, N8582, N2516, N5493);
nor NOR4 (N8587, N8573, N2161, N1904, N1717);
buf BUF1 (N8588, N8571);
nor NOR2 (N8589, N8579, N3159);
buf BUF1 (N8590, N8577);
and AND4 (N8591, N8586, N1370, N5051, N4043);
nand NAND3 (N8592, N8585, N1758, N3060);
and AND4 (N8593, N8589, N8508, N4390, N1902);
or OR4 (N8594, N8588, N4373, N4041, N3343);
or OR3 (N8595, N8580, N4143, N1943);
and AND4 (N8596, N8569, N3891, N5359, N1445);
buf BUF1 (N8597, N8596);
nor NOR2 (N8598, N8595, N2271);
nand NAND2 (N8599, N8568, N497);
buf BUF1 (N8600, N8594);
and AND2 (N8601, N8587, N2306);
or OR2 (N8602, N8578, N5345);
not NOT1 (N8603, N8591);
nand NAND4 (N8604, N8590, N3299, N1255, N2177);
xor XOR2 (N8605, N8600, N2781);
or OR2 (N8606, N8601, N7899);
xor XOR2 (N8607, N8606, N1000);
xor XOR2 (N8608, N8605, N3530);
buf BUF1 (N8609, N8608);
xor XOR2 (N8610, N8603, N1832);
buf BUF1 (N8611, N8597);
xor XOR2 (N8612, N8610, N6922);
buf BUF1 (N8613, N8607);
or OR2 (N8614, N8602, N2940);
not NOT1 (N8615, N8599);
or OR2 (N8616, N8611, N3855);
buf BUF1 (N8617, N8613);
nand NAND3 (N8618, N8609, N4467, N914);
or OR4 (N8619, N8604, N7058, N5771, N6795);
and AND4 (N8620, N8614, N2184, N3187, N3799);
and AND3 (N8621, N8615, N4459, N7609);
not NOT1 (N8622, N8616);
and AND2 (N8623, N8612, N7932);
buf BUF1 (N8624, N8593);
not NOT1 (N8625, N8624);
not NOT1 (N8626, N8623);
nor NOR4 (N8627, N8622, N2855, N2512, N3852);
not NOT1 (N8628, N8592);
and AND2 (N8629, N8598, N5198);
or OR3 (N8630, N8629, N5255, N6259);
and AND2 (N8631, N8619, N2109);
nand NAND3 (N8632, N8625, N7260, N7175);
nand NAND2 (N8633, N8631, N8091);
or OR2 (N8634, N8618, N2712);
nand NAND2 (N8635, N8630, N7204);
not NOT1 (N8636, N8634);
buf BUF1 (N8637, N8620);
buf BUF1 (N8638, N8627);
xor XOR2 (N8639, N8621, N3437);
or OR3 (N8640, N8636, N257, N8108);
not NOT1 (N8641, N8632);
xor XOR2 (N8642, N8628, N5918);
or OR3 (N8643, N8635, N1285, N3691);
xor XOR2 (N8644, N8637, N6989);
not NOT1 (N8645, N8641);
and AND3 (N8646, N8626, N5257, N6748);
nor NOR3 (N8647, N8633, N8159, N4429);
nor NOR4 (N8648, N8643, N5608, N6846, N6091);
buf BUF1 (N8649, N8644);
and AND2 (N8650, N8647, N2930);
or OR3 (N8651, N8617, N2835, N6698);
xor XOR2 (N8652, N8651, N5873);
buf BUF1 (N8653, N8642);
not NOT1 (N8654, N8652);
not NOT1 (N8655, N8646);
nand NAND2 (N8656, N8638, N3625);
buf BUF1 (N8657, N8639);
nand NAND3 (N8658, N8649, N1379, N788);
nor NOR4 (N8659, N8658, N5857, N6384, N3122);
buf BUF1 (N8660, N8648);
nor NOR2 (N8661, N8650, N5496);
xor XOR2 (N8662, N8657, N2938);
nand NAND3 (N8663, N8655, N1710, N1498);
nand NAND4 (N8664, N8660, N6748, N6977, N6199);
nand NAND3 (N8665, N8664, N7274, N1646);
and AND3 (N8666, N8645, N7186, N8186);
xor XOR2 (N8667, N8662, N1973);
and AND4 (N8668, N8640, N7339, N7426, N6235);
or OR2 (N8669, N8666, N3267);
and AND3 (N8670, N8654, N7644, N3240);
xor XOR2 (N8671, N8670, N1444);
buf BUF1 (N8672, N8671);
nor NOR2 (N8673, N8668, N8120);
nand NAND3 (N8674, N8673, N2338, N7548);
or OR4 (N8675, N8669, N4175, N3972, N4486);
xor XOR2 (N8676, N8674, N4603);
or OR3 (N8677, N8661, N6748, N4509);
nand NAND3 (N8678, N8676, N8430, N2643);
and AND4 (N8679, N8653, N4260, N7891, N7172);
nand NAND3 (N8680, N8672, N5339, N2298);
nor NOR4 (N8681, N8665, N7534, N4584, N6795);
xor XOR2 (N8682, N8675, N1081);
not NOT1 (N8683, N8677);
buf BUF1 (N8684, N8663);
and AND3 (N8685, N8679, N7774, N5703);
or OR2 (N8686, N8678, N931);
or OR4 (N8687, N8682, N786, N77, N1309);
and AND2 (N8688, N8683, N3487);
nor NOR3 (N8689, N8680, N8310, N8000);
xor XOR2 (N8690, N8659, N6963);
not NOT1 (N8691, N8667);
and AND3 (N8692, N8681, N2495, N7632);
nor NOR4 (N8693, N8692, N7238, N5705, N3967);
buf BUF1 (N8694, N8688);
nor NOR4 (N8695, N8656, N3422, N5507, N1788);
or OR3 (N8696, N8686, N5458, N6552);
nor NOR4 (N8697, N8690, N4924, N7229, N7095);
and AND2 (N8698, N8696, N2038);
nor NOR4 (N8699, N8694, N2647, N8180, N7931);
nor NOR4 (N8700, N8691, N4379, N7987, N8256);
nand NAND2 (N8701, N8693, N3766);
not NOT1 (N8702, N8701);
nand NAND2 (N8703, N8695, N5910);
nor NOR2 (N8704, N8687, N5507);
or OR4 (N8705, N8700, N4343, N821, N6946);
and AND3 (N8706, N8699, N3023, N5428);
nor NOR2 (N8707, N8689, N2687);
and AND2 (N8708, N8685, N7578);
nor NOR3 (N8709, N8697, N6574, N8672);
not NOT1 (N8710, N8706);
buf BUF1 (N8711, N8707);
xor XOR2 (N8712, N8702, N1920);
or OR3 (N8713, N8684, N1261, N4983);
and AND2 (N8714, N8710, N4752);
xor XOR2 (N8715, N8713, N2418);
buf BUF1 (N8716, N8708);
not NOT1 (N8717, N8711);
buf BUF1 (N8718, N8703);
nor NOR3 (N8719, N8715, N2379, N1754);
buf BUF1 (N8720, N8716);
nor NOR4 (N8721, N8714, N2211, N3531, N4505);
nor NOR3 (N8722, N8704, N1266, N1569);
buf BUF1 (N8723, N8722);
or OR4 (N8724, N8709, N2719, N1122, N3311);
not NOT1 (N8725, N8720);
and AND4 (N8726, N8723, N3309, N3875, N566);
or OR2 (N8727, N8726, N7360);
xor XOR2 (N8728, N8721, N3299);
nor NOR3 (N8729, N8705, N828, N8128);
xor XOR2 (N8730, N8725, N3654);
and AND3 (N8731, N8730, N4979, N329);
xor XOR2 (N8732, N8727, N8119);
xor XOR2 (N8733, N8729, N4682);
not NOT1 (N8734, N8728);
nand NAND4 (N8735, N8719, N5216, N7182, N4852);
xor XOR2 (N8736, N8732, N3596);
or OR3 (N8737, N8731, N8000, N8391);
xor XOR2 (N8738, N8736, N8333);
nor NOR2 (N8739, N8737, N7701);
nor NOR3 (N8740, N8712, N2848, N1354);
buf BUF1 (N8741, N8698);
nand NAND4 (N8742, N8734, N7073, N1329, N6632);
and AND2 (N8743, N8738, N921);
xor XOR2 (N8744, N8724, N6165);
not NOT1 (N8745, N8739);
or OR3 (N8746, N8744, N5178, N7113);
buf BUF1 (N8747, N8741);
nor NOR3 (N8748, N8745, N4293, N7316);
buf BUF1 (N8749, N8718);
buf BUF1 (N8750, N8717);
nand NAND2 (N8751, N8746, N4352);
nor NOR2 (N8752, N8748, N5792);
and AND4 (N8753, N8743, N6268, N1964, N1217);
and AND4 (N8754, N8750, N3982, N5797, N4989);
or OR4 (N8755, N8735, N2459, N330, N7481);
nand NAND4 (N8756, N8733, N2123, N3583, N3744);
not NOT1 (N8757, N8756);
nor NOR2 (N8758, N8752, N5866);
xor XOR2 (N8759, N8758, N3143);
or OR3 (N8760, N8751, N2640, N126);
not NOT1 (N8761, N8749);
xor XOR2 (N8762, N8753, N479);
buf BUF1 (N8763, N8759);
xor XOR2 (N8764, N8762, N4199);
not NOT1 (N8765, N8747);
nand NAND2 (N8766, N8742, N8340);
and AND3 (N8767, N8754, N278, N698);
not NOT1 (N8768, N8764);
not NOT1 (N8769, N8768);
xor XOR2 (N8770, N8763, N1529);
nand NAND2 (N8771, N8766, N7778);
nand NAND3 (N8772, N8761, N1705, N7430);
xor XOR2 (N8773, N8757, N8501);
nand NAND3 (N8774, N8760, N4905, N2516);
not NOT1 (N8775, N8774);
xor XOR2 (N8776, N8772, N2116);
nand NAND4 (N8777, N8770, N5183, N6624, N2980);
nor NOR2 (N8778, N8771, N3264);
xor XOR2 (N8779, N8775, N3163);
nor NOR3 (N8780, N8777, N6291, N4367);
or OR3 (N8781, N8769, N8127, N5831);
not NOT1 (N8782, N8778);
buf BUF1 (N8783, N8782);
or OR4 (N8784, N8765, N2486, N977, N188);
nand NAND2 (N8785, N8784, N2758);
nor NOR4 (N8786, N8773, N3737, N2696, N4580);
xor XOR2 (N8787, N8755, N4424);
or OR3 (N8788, N8787, N146, N4838);
nor NOR3 (N8789, N8740, N121, N4627);
or OR3 (N8790, N8767, N1954, N5819);
not NOT1 (N8791, N8789);
not NOT1 (N8792, N8791);
or OR2 (N8793, N8781, N2018);
or OR4 (N8794, N8786, N5291, N2917, N2446);
not NOT1 (N8795, N8788);
buf BUF1 (N8796, N8776);
or OR2 (N8797, N8794, N2049);
buf BUF1 (N8798, N8792);
nand NAND4 (N8799, N8780, N6374, N1926, N5797);
xor XOR2 (N8800, N8798, N6644);
buf BUF1 (N8801, N8800);
not NOT1 (N8802, N8797);
or OR2 (N8803, N8795, N658);
nor NOR2 (N8804, N8802, N362);
nor NOR2 (N8805, N8790, N4335);
xor XOR2 (N8806, N8801, N7890);
nand NAND3 (N8807, N8804, N7661, N2683);
buf BUF1 (N8808, N8793);
or OR4 (N8809, N8808, N6442, N7265, N3057);
not NOT1 (N8810, N8785);
and AND3 (N8811, N8779, N7170, N524);
nor NOR2 (N8812, N8811, N4722);
buf BUF1 (N8813, N8807);
nor NOR3 (N8814, N8803, N2330, N793);
buf BUF1 (N8815, N8805);
nand NAND3 (N8816, N8810, N4989, N3226);
nor NOR4 (N8817, N8783, N5297, N8492, N2319);
nand NAND4 (N8818, N8799, N8199, N4009, N8331);
or OR3 (N8819, N8816, N6040, N4633);
nor NOR4 (N8820, N8796, N377, N6159, N8136);
buf BUF1 (N8821, N8813);
or OR2 (N8822, N8821, N4888);
buf BUF1 (N8823, N8822);
and AND3 (N8824, N8818, N6603, N3083);
nand NAND2 (N8825, N8817, N1135);
nor NOR4 (N8826, N8819, N8400, N2118, N956);
nor NOR4 (N8827, N8806, N4432, N2352, N7528);
and AND3 (N8828, N8820, N5394, N5805);
or OR3 (N8829, N8814, N6300, N1418);
not NOT1 (N8830, N8826);
not NOT1 (N8831, N8830);
nand NAND3 (N8832, N8828, N3884, N7375);
buf BUF1 (N8833, N8831);
nor NOR2 (N8834, N8833, N5979);
nand NAND2 (N8835, N8823, N5807);
buf BUF1 (N8836, N8809);
or OR4 (N8837, N8834, N214, N8125, N7237);
not NOT1 (N8838, N8837);
buf BUF1 (N8839, N8812);
not NOT1 (N8840, N8829);
not NOT1 (N8841, N8832);
nor NOR2 (N8842, N8836, N2747);
and AND2 (N8843, N8842, N4198);
nand NAND3 (N8844, N8843, N5001, N1753);
nand NAND4 (N8845, N8835, N1894, N107, N5432);
or OR3 (N8846, N8845, N5805, N2514);
xor XOR2 (N8847, N8839, N7483);
or OR3 (N8848, N8840, N8218, N4247);
or OR2 (N8849, N8844, N7582);
xor XOR2 (N8850, N8841, N6175);
nor NOR3 (N8851, N8815, N8251, N8600);
xor XOR2 (N8852, N8847, N7758);
not NOT1 (N8853, N8851);
not NOT1 (N8854, N8852);
and AND2 (N8855, N8853, N1672);
buf BUF1 (N8856, N8855);
buf BUF1 (N8857, N8827);
nand NAND2 (N8858, N8824, N5058);
nand NAND2 (N8859, N8848, N7185);
and AND2 (N8860, N8838, N268);
xor XOR2 (N8861, N8846, N1703);
not NOT1 (N8862, N8849);
nand NAND3 (N8863, N8856, N802, N3490);
xor XOR2 (N8864, N8859, N1254);
nand NAND4 (N8865, N8860, N5741, N2364, N1358);
and AND3 (N8866, N8850, N26, N1119);
not NOT1 (N8867, N8857);
buf BUF1 (N8868, N8854);
and AND2 (N8869, N8866, N1220);
nand NAND4 (N8870, N8868, N8455, N2120, N8109);
nand NAND3 (N8871, N8870, N5748, N6628);
and AND4 (N8872, N8862, N8791, N4144, N3371);
nand NAND2 (N8873, N8858, N7488);
xor XOR2 (N8874, N8865, N5790);
nor NOR2 (N8875, N8874, N3912);
and AND3 (N8876, N8864, N7174, N4238);
nor NOR2 (N8877, N8867, N5834);
nor NOR4 (N8878, N8869, N6737, N3924, N1581);
not NOT1 (N8879, N8873);
or OR3 (N8880, N8825, N6415, N2688);
buf BUF1 (N8881, N8877);
and AND3 (N8882, N8863, N2676, N2100);
and AND4 (N8883, N8875, N3614, N5668, N7895);
nor NOR3 (N8884, N8871, N3678, N8570);
nand NAND2 (N8885, N8872, N2537);
not NOT1 (N8886, N8861);
or OR4 (N8887, N8881, N1534, N5086, N5172);
and AND4 (N8888, N8886, N5015, N6124, N2110);
nand NAND3 (N8889, N8888, N6717, N6785);
nor NOR3 (N8890, N8880, N6381, N3241);
nand NAND2 (N8891, N8885, N1800);
nand NAND3 (N8892, N8889, N7936, N7094);
and AND3 (N8893, N8890, N7737, N7974);
or OR2 (N8894, N8883, N4438);
nand NAND3 (N8895, N8884, N3036, N427);
xor XOR2 (N8896, N8882, N6688);
nand NAND2 (N8897, N8892, N6701);
nand NAND3 (N8898, N8891, N6348, N308);
nand NAND4 (N8899, N8878, N3606, N5491, N487);
and AND2 (N8900, N8887, N6222);
xor XOR2 (N8901, N8879, N4917);
nor NOR2 (N8902, N8876, N6922);
nor NOR4 (N8903, N8893, N7156, N4702, N3903);
xor XOR2 (N8904, N8895, N7291);
and AND2 (N8905, N8897, N538);
buf BUF1 (N8906, N8894);
xor XOR2 (N8907, N8901, N2163);
nand NAND3 (N8908, N8903, N3271, N7995);
xor XOR2 (N8909, N8896, N257);
buf BUF1 (N8910, N8905);
nor NOR3 (N8911, N8899, N7900, N4909);
not NOT1 (N8912, N8909);
xor XOR2 (N8913, N8912, N2895);
and AND2 (N8914, N8911, N7662);
xor XOR2 (N8915, N8900, N924);
or OR4 (N8916, N8914, N1991, N3771, N8115);
not NOT1 (N8917, N8902);
nor NOR4 (N8918, N8917, N7870, N4677, N2442);
and AND2 (N8919, N8915, N4254);
buf BUF1 (N8920, N8913);
or OR4 (N8921, N8910, N1248, N6603, N4840);
or OR3 (N8922, N8898, N3861, N5413);
nor NOR3 (N8923, N8922, N5669, N8701);
or OR2 (N8924, N8919, N4307);
and AND3 (N8925, N8921, N7793, N7015);
and AND3 (N8926, N8918, N7669, N3032);
xor XOR2 (N8927, N8906, N7236);
or OR2 (N8928, N8925, N5544);
nand NAND4 (N8929, N8923, N6933, N5838, N6942);
buf BUF1 (N8930, N8924);
xor XOR2 (N8931, N8926, N7068);
buf BUF1 (N8932, N8927);
xor XOR2 (N8933, N8930, N5000);
nor NOR2 (N8934, N8920, N957);
nand NAND4 (N8935, N8916, N4552, N3993, N3284);
buf BUF1 (N8936, N8934);
xor XOR2 (N8937, N8907, N5547);
buf BUF1 (N8938, N8908);
or OR3 (N8939, N8931, N1366, N3909);
buf BUF1 (N8940, N8932);
buf BUF1 (N8941, N8928);
nand NAND2 (N8942, N8939, N2903);
and AND4 (N8943, N8933, N1752, N5616, N3938);
nor NOR2 (N8944, N8937, N7733);
buf BUF1 (N8945, N8929);
xor XOR2 (N8946, N8945, N3710);
and AND2 (N8947, N8940, N6549);
or OR3 (N8948, N8942, N2276, N5896);
or OR4 (N8949, N8904, N1302, N7349, N394);
nor NOR2 (N8950, N8936, N5592);
not NOT1 (N8951, N8938);
and AND4 (N8952, N8944, N7781, N8330, N1783);
xor XOR2 (N8953, N8949, N5642);
or OR3 (N8954, N8951, N7298, N1703);
and AND3 (N8955, N8943, N7940, N3368);
nor NOR4 (N8956, N8955, N3724, N1980, N3212);
nor NOR3 (N8957, N8950, N8833, N5366);
nand NAND2 (N8958, N8948, N95);
nor NOR4 (N8959, N8947, N5437, N1783, N4939);
nand NAND2 (N8960, N8957, N1113);
buf BUF1 (N8961, N8941);
nand NAND3 (N8962, N8935, N7141, N2291);
or OR4 (N8963, N8961, N7590, N3463, N4096);
nor NOR4 (N8964, N8954, N7865, N2261, N2267);
or OR4 (N8965, N8963, N3111, N3737, N4973);
nor NOR2 (N8966, N8964, N2893);
or OR4 (N8967, N8956, N3477, N4965, N492);
or OR2 (N8968, N8965, N4157);
xor XOR2 (N8969, N8952, N8167);
nand NAND3 (N8970, N8960, N1332, N6719);
nand NAND2 (N8971, N8958, N7907);
and AND3 (N8972, N8967, N2442, N967);
or OR4 (N8973, N8968, N8361, N6767, N670);
and AND2 (N8974, N8966, N4068);
not NOT1 (N8975, N8969);
xor XOR2 (N8976, N8962, N4557);
nand NAND2 (N8977, N8972, N406);
nor NOR4 (N8978, N8971, N2629, N4908, N8695);
not NOT1 (N8979, N8959);
not NOT1 (N8980, N8953);
or OR2 (N8981, N8979, N8182);
nand NAND3 (N8982, N8977, N5707, N3665);
buf BUF1 (N8983, N8970);
xor XOR2 (N8984, N8981, N2087);
xor XOR2 (N8985, N8976, N6070);
xor XOR2 (N8986, N8973, N8933);
and AND3 (N8987, N8982, N3133, N1736);
xor XOR2 (N8988, N8985, N1077);
nand NAND2 (N8989, N8988, N6530);
or OR3 (N8990, N8986, N640, N2084);
nand NAND4 (N8991, N8984, N8100, N1347, N5393);
not NOT1 (N8992, N8987);
or OR3 (N8993, N8978, N1712, N5367);
and AND4 (N8994, N8989, N2535, N7050, N855);
nor NOR3 (N8995, N8991, N3992, N116);
nor NOR2 (N8996, N8983, N5178);
nand NAND2 (N8997, N8974, N7086);
nor NOR2 (N8998, N8994, N3008);
not NOT1 (N8999, N8946);
and AND4 (N9000, N8975, N6179, N3156, N2564);
and AND2 (N9001, N8993, N2855);
nand NAND2 (N9002, N9001, N2564);
buf BUF1 (N9003, N8980);
nand NAND4 (N9004, N9002, N6699, N6366, N3849);
xor XOR2 (N9005, N9004, N6466);
or OR4 (N9006, N8995, N6233, N6948, N7703);
or OR2 (N9007, N8992, N3357);
and AND2 (N9008, N8999, N6452);
not NOT1 (N9009, N8996);
and AND2 (N9010, N8998, N6271);
xor XOR2 (N9011, N9010, N5141);
or OR2 (N9012, N9006, N6381);
buf BUF1 (N9013, N9011);
nand NAND3 (N9014, N9013, N7825, N5827);
xor XOR2 (N9015, N9000, N2560);
not NOT1 (N9016, N9008);
nand NAND3 (N9017, N8997, N1156, N1931);
and AND3 (N9018, N9009, N5803, N5177);
and AND2 (N9019, N9016, N6209);
and AND3 (N9020, N9007, N2599, N3032);
and AND2 (N9021, N9014, N289);
and AND3 (N9022, N9005, N3400, N1298);
not NOT1 (N9023, N9012);
and AND4 (N9024, N9023, N8131, N41, N6439);
buf BUF1 (N9025, N9022);
nand NAND2 (N9026, N9025, N5801);
nand NAND4 (N9027, N9003, N3099, N5344, N73);
nor NOR2 (N9028, N9018, N7355);
and AND3 (N9029, N9019, N7722, N7443);
or OR3 (N9030, N9017, N2375, N7881);
or OR4 (N9031, N9027, N1117, N4644, N407);
buf BUF1 (N9032, N8990);
buf BUF1 (N9033, N9020);
nand NAND2 (N9034, N9021, N6126);
or OR3 (N9035, N9028, N7159, N2297);
or OR3 (N9036, N9033, N3179, N3871);
nor NOR4 (N9037, N9034, N8890, N2605, N4762);
nand NAND3 (N9038, N9036, N110, N2038);
or OR2 (N9039, N9032, N4316);
buf BUF1 (N9040, N9024);
not NOT1 (N9041, N9035);
or OR2 (N9042, N9039, N1332);
nand NAND3 (N9043, N9041, N8075, N5343);
and AND2 (N9044, N9026, N3682);
or OR2 (N9045, N9037, N8624);
buf BUF1 (N9046, N9043);
xor XOR2 (N9047, N9038, N7182);
and AND3 (N9048, N9046, N900, N2989);
buf BUF1 (N9049, N9044);
xor XOR2 (N9050, N9045, N5326);
not NOT1 (N9051, N9049);
buf BUF1 (N9052, N9015);
not NOT1 (N9053, N9042);
xor XOR2 (N9054, N9051, N2454);
not NOT1 (N9055, N9048);
nand NAND4 (N9056, N9053, N151, N1458, N2437);
nand NAND2 (N9057, N9047, N2192);
buf BUF1 (N9058, N9054);
and AND2 (N9059, N9058, N6523);
not NOT1 (N9060, N9052);
buf BUF1 (N9061, N9030);
nand NAND3 (N9062, N9057, N4088, N8735);
xor XOR2 (N9063, N9061, N1141);
buf BUF1 (N9064, N9060);
buf BUF1 (N9065, N9056);
and AND2 (N9066, N9055, N6139);
not NOT1 (N9067, N9040);
or OR3 (N9068, N9059, N5311, N8416);
not NOT1 (N9069, N9031);
nand NAND2 (N9070, N9068, N8947);
xor XOR2 (N9071, N9067, N1826);
nand NAND4 (N9072, N9070, N64, N58, N2931);
or OR4 (N9073, N9071, N4217, N950, N5606);
and AND4 (N9074, N9065, N4162, N3487, N3477);
nand NAND3 (N9075, N9063, N8256, N6735);
nand NAND2 (N9076, N9069, N8682);
and AND2 (N9077, N9075, N1988);
xor XOR2 (N9078, N9074, N3229);
or OR2 (N9079, N9029, N5488);
and AND3 (N9080, N9062, N4860, N8255);
nor NOR3 (N9081, N9072, N7058, N1257);
nor NOR3 (N9082, N9077, N7531, N3510);
and AND4 (N9083, N9050, N3357, N4263, N1176);
buf BUF1 (N9084, N9078);
nand NAND3 (N9085, N9084, N5953, N2854);
not NOT1 (N9086, N9082);
and AND4 (N9087, N9080, N5186, N5182, N2734);
or OR4 (N9088, N9087, N832, N4599, N9021);
nand NAND4 (N9089, N9086, N8229, N1189, N3892);
buf BUF1 (N9090, N9089);
nor NOR2 (N9091, N9081, N4498);
or OR3 (N9092, N9066, N4483, N4390);
nand NAND3 (N9093, N9073, N4834, N1142);
and AND4 (N9094, N9085, N2547, N5102, N953);
or OR3 (N9095, N9092, N8340, N5975);
nand NAND4 (N9096, N9083, N4634, N3548, N3353);
or OR4 (N9097, N9095, N3046, N2070, N8038);
nor NOR4 (N9098, N9097, N3919, N4569, N3624);
and AND2 (N9099, N9093, N8999);
buf BUF1 (N9100, N9076);
nor NOR4 (N9101, N9064, N7875, N8387, N2490);
nand NAND3 (N9102, N9088, N5743, N7139);
nor NOR3 (N9103, N9091, N4574, N6485);
buf BUF1 (N9104, N9103);
nor NOR4 (N9105, N9090, N8019, N5075, N1674);
nor NOR3 (N9106, N9102, N6856, N774);
buf BUF1 (N9107, N9079);
nor NOR2 (N9108, N9098, N8831);
buf BUF1 (N9109, N9108);
nand NAND2 (N9110, N9101, N5654);
xor XOR2 (N9111, N9107, N4060);
xor XOR2 (N9112, N9099, N8428);
nand NAND4 (N9113, N9110, N8269, N463, N4512);
not NOT1 (N9114, N9094);
nand NAND4 (N9115, N9111, N1647, N5439, N2372);
nor NOR3 (N9116, N9109, N7894, N2801);
and AND2 (N9117, N9106, N4947);
or OR3 (N9118, N9096, N6194, N7544);
and AND2 (N9119, N9114, N6675);
and AND4 (N9120, N9104, N1668, N2919, N5907);
or OR4 (N9121, N9112, N8517, N8263, N1062);
or OR2 (N9122, N9116, N6949);
xor XOR2 (N9123, N9100, N2347);
buf BUF1 (N9124, N9122);
nand NAND3 (N9125, N9118, N5166, N1860);
or OR2 (N9126, N9120, N4858);
nor NOR3 (N9127, N9123, N3549, N916);
nor NOR3 (N9128, N9119, N2842, N9030);
nand NAND3 (N9129, N9128, N213, N3798);
or OR4 (N9130, N9129, N5226, N6578, N9051);
or OR3 (N9131, N9105, N871, N6762);
xor XOR2 (N9132, N9121, N7861);
buf BUF1 (N9133, N9117);
nand NAND3 (N9134, N9132, N4862, N4542);
and AND4 (N9135, N9126, N4412, N3515, N4942);
nand NAND3 (N9136, N9124, N2929, N9092);
and AND2 (N9137, N9125, N4863);
buf BUF1 (N9138, N9131);
nor NOR3 (N9139, N9138, N7835, N4902);
or OR4 (N9140, N9134, N7472, N3446, N8813);
buf BUF1 (N9141, N9136);
nand NAND2 (N9142, N9133, N6548);
not NOT1 (N9143, N9139);
and AND2 (N9144, N9115, N7557);
nand NAND2 (N9145, N9144, N7864);
not NOT1 (N9146, N9130);
or OR2 (N9147, N9140, N5182);
or OR4 (N9148, N9135, N694, N8460, N2783);
buf BUF1 (N9149, N9146);
xor XOR2 (N9150, N9147, N3195);
xor XOR2 (N9151, N9142, N3909);
nor NOR2 (N9152, N9145, N3198);
buf BUF1 (N9153, N9141);
nor NOR4 (N9154, N9149, N2127, N1825, N196);
not NOT1 (N9155, N9143);
not NOT1 (N9156, N9148);
nor NOR3 (N9157, N9113, N4723, N7547);
or OR4 (N9158, N9156, N3323, N2986, N1030);
xor XOR2 (N9159, N9153, N4404);
xor XOR2 (N9160, N9159, N4473);
and AND3 (N9161, N9127, N5469, N7785);
nand NAND2 (N9162, N9154, N6997);
not NOT1 (N9163, N9157);
or OR4 (N9164, N9151, N8109, N2166, N3040);
not NOT1 (N9165, N9155);
nand NAND3 (N9166, N9150, N8710, N3949);
nor NOR3 (N9167, N9137, N405, N2754);
nor NOR4 (N9168, N9160, N5986, N990, N2524);
and AND4 (N9169, N9165, N8858, N6167, N5918);
buf BUF1 (N9170, N9169);
nand NAND4 (N9171, N9158, N3934, N8062, N3289);
or OR4 (N9172, N9161, N8969, N3140, N3164);
not NOT1 (N9173, N9162);
or OR3 (N9174, N9168, N583, N9075);
not NOT1 (N9175, N9164);
nand NAND2 (N9176, N9172, N2388);
buf BUF1 (N9177, N9152);
buf BUF1 (N9178, N9167);
buf BUF1 (N9179, N9175);
nand NAND3 (N9180, N9179, N2228, N303);
and AND4 (N9181, N9171, N5947, N3915, N7751);
and AND2 (N9182, N9180, N7015);
not NOT1 (N9183, N9182);
or OR4 (N9184, N9178, N8893, N7584, N6657);
not NOT1 (N9185, N9177);
xor XOR2 (N9186, N9173, N3953);
not NOT1 (N9187, N9174);
or OR4 (N9188, N9183, N607, N3995, N2973);
and AND4 (N9189, N9166, N6267, N1680, N7858);
xor XOR2 (N9190, N9163, N4607);
nand NAND4 (N9191, N9185, N6236, N3065, N2957);
not NOT1 (N9192, N9187);
xor XOR2 (N9193, N9181, N7557);
nand NAND4 (N9194, N9184, N466, N824, N801);
nor NOR3 (N9195, N9191, N3847, N5647);
not NOT1 (N9196, N9192);
nor NOR2 (N9197, N9176, N6221);
buf BUF1 (N9198, N9190);
not NOT1 (N9199, N9195);
or OR2 (N9200, N9194, N8525);
xor XOR2 (N9201, N9197, N4953);
not NOT1 (N9202, N9188);
not NOT1 (N9203, N9186);
xor XOR2 (N9204, N9199, N6872);
and AND3 (N9205, N9201, N5353, N2285);
buf BUF1 (N9206, N9193);
not NOT1 (N9207, N9203);
buf BUF1 (N9208, N9196);
not NOT1 (N9209, N9170);
and AND3 (N9210, N9206, N8733, N7940);
not NOT1 (N9211, N9204);
buf BUF1 (N9212, N9211);
xor XOR2 (N9213, N9207, N6199);
not NOT1 (N9214, N9200);
not NOT1 (N9215, N9198);
or OR4 (N9216, N9213, N5795, N1302, N2184);
nand NAND2 (N9217, N9216, N4218);
or OR2 (N9218, N9205, N864);
and AND3 (N9219, N9217, N4250, N3796);
and AND4 (N9220, N9202, N7693, N3109, N3661);
not NOT1 (N9221, N9214);
xor XOR2 (N9222, N9215, N7590);
not NOT1 (N9223, N9208);
nand NAND2 (N9224, N9212, N1363);
nand NAND3 (N9225, N9209, N3372, N8621);
nor NOR2 (N9226, N9222, N7352);
not NOT1 (N9227, N9219);
xor XOR2 (N9228, N9218, N8162);
nor NOR3 (N9229, N9210, N652, N959);
or OR4 (N9230, N9223, N6150, N6778, N5673);
and AND3 (N9231, N9221, N3809, N1734);
nor NOR4 (N9232, N9226, N680, N263, N7991);
or OR4 (N9233, N9231, N4364, N7919, N3289);
xor XOR2 (N9234, N9189, N1950);
nand NAND4 (N9235, N9234, N8561, N3623, N7060);
nor NOR2 (N9236, N9220, N707);
not NOT1 (N9237, N9232);
xor XOR2 (N9238, N9224, N4700);
xor XOR2 (N9239, N9225, N4861);
xor XOR2 (N9240, N9230, N5432);
and AND3 (N9241, N9228, N6735, N4482);
nand NAND2 (N9242, N9240, N1301);
nand NAND3 (N9243, N9238, N6434, N8568);
and AND4 (N9244, N9236, N3739, N4850, N4376);
nor NOR3 (N9245, N9235, N2518, N5751);
or OR2 (N9246, N9241, N5224);
nand NAND3 (N9247, N9246, N3762, N4384);
nor NOR2 (N9248, N9245, N8893);
and AND2 (N9249, N9233, N9037);
or OR2 (N9250, N9248, N3614);
nor NOR2 (N9251, N9242, N4881);
and AND2 (N9252, N9251, N6515);
nand NAND3 (N9253, N9243, N1845, N7976);
xor XOR2 (N9254, N9237, N4223);
or OR4 (N9255, N9229, N1604, N4549, N7050);
xor XOR2 (N9256, N9255, N8125);
and AND2 (N9257, N9254, N3101);
buf BUF1 (N9258, N9244);
nand NAND3 (N9259, N9253, N903, N5278);
buf BUF1 (N9260, N9257);
xor XOR2 (N9261, N9256, N8416);
and AND3 (N9262, N9249, N5149, N6270);
buf BUF1 (N9263, N9259);
xor XOR2 (N9264, N9261, N5183);
and AND4 (N9265, N9227, N7584, N1902, N8254);
not NOT1 (N9266, N9262);
nor NOR4 (N9267, N9266, N7091, N3519, N2670);
and AND3 (N9268, N9258, N5093, N5614);
nor NOR3 (N9269, N9268, N7828, N2120);
xor XOR2 (N9270, N9260, N1753);
not NOT1 (N9271, N9264);
nand NAND3 (N9272, N9269, N2624, N1890);
nor NOR4 (N9273, N9252, N8620, N8615, N1570);
xor XOR2 (N9274, N9272, N7215);
nand NAND4 (N9275, N9274, N1521, N7034, N8825);
xor XOR2 (N9276, N9265, N3086);
and AND2 (N9277, N9270, N1288);
not NOT1 (N9278, N9247);
xor XOR2 (N9279, N9273, N3801);
and AND2 (N9280, N9267, N4896);
or OR4 (N9281, N9239, N5690, N2705, N1197);
nor NOR2 (N9282, N9281, N3411);
xor XOR2 (N9283, N9280, N53);
xor XOR2 (N9284, N9282, N836);
nor NOR3 (N9285, N9279, N8971, N4985);
or OR4 (N9286, N9263, N334, N7492, N5472);
nand NAND2 (N9287, N9277, N5162);
and AND2 (N9288, N9285, N3741);
buf BUF1 (N9289, N9286);
buf BUF1 (N9290, N9271);
nor NOR4 (N9291, N9250, N907, N2552, N1401);
buf BUF1 (N9292, N9284);
nand NAND4 (N9293, N9292, N7082, N1213, N4237);
xor XOR2 (N9294, N9288, N4328);
nor NOR2 (N9295, N9278, N7605);
buf BUF1 (N9296, N9275);
xor XOR2 (N9297, N9294, N8459);
xor XOR2 (N9298, N9291, N5052);
or OR3 (N9299, N9293, N1151, N2500);
nand NAND3 (N9300, N9298, N5773, N5021);
buf BUF1 (N9301, N9297);
or OR4 (N9302, N9290, N2898, N6104, N5333);
buf BUF1 (N9303, N9301);
xor XOR2 (N9304, N9295, N1946);
or OR2 (N9305, N9289, N8649);
and AND2 (N9306, N9283, N8969);
not NOT1 (N9307, N9303);
and AND2 (N9308, N9307, N2640);
xor XOR2 (N9309, N9306, N4122);
nand NAND2 (N9310, N9296, N3372);
xor XOR2 (N9311, N9304, N1066);
not NOT1 (N9312, N9276);
nor NOR2 (N9313, N9305, N7644);
or OR2 (N9314, N9309, N6599);
xor XOR2 (N9315, N9302, N760);
nor NOR3 (N9316, N9314, N5845, N1936);
nand NAND2 (N9317, N9308, N3467);
nand NAND2 (N9318, N9315, N3532);
buf BUF1 (N9319, N9318);
not NOT1 (N9320, N9310);
not NOT1 (N9321, N9287);
nor NOR2 (N9322, N9311, N5197);
xor XOR2 (N9323, N9322, N9192);
nor NOR2 (N9324, N9323, N1793);
and AND4 (N9325, N9317, N107, N8222, N1334);
buf BUF1 (N9326, N9300);
nor NOR2 (N9327, N9321, N609);
nand NAND3 (N9328, N9312, N6714, N6659);
not NOT1 (N9329, N9326);
or OR3 (N9330, N9319, N2953, N7798);
or OR3 (N9331, N9299, N7790, N7388);
nand NAND4 (N9332, N9324, N8680, N7031, N4017);
or OR4 (N9333, N9325, N5208, N3629, N6881);
nand NAND3 (N9334, N9330, N9237, N8510);
xor XOR2 (N9335, N9333, N7732);
nand NAND4 (N9336, N9328, N1355, N7743, N5207);
nor NOR3 (N9337, N9320, N5252, N4132);
nor NOR4 (N9338, N9335, N5847, N4874, N1241);
or OR2 (N9339, N9336, N6818);
not NOT1 (N9340, N9329);
nand NAND3 (N9341, N9316, N3522, N1777);
not NOT1 (N9342, N9340);
nor NOR3 (N9343, N9342, N8406, N9094);
buf BUF1 (N9344, N9339);
nor NOR3 (N9345, N9344, N4492, N8655);
nor NOR4 (N9346, N9327, N9310, N6855, N2993);
not NOT1 (N9347, N9313);
buf BUF1 (N9348, N9347);
xor XOR2 (N9349, N9338, N229);
nor NOR4 (N9350, N9346, N5215, N2141, N4776);
nand NAND4 (N9351, N9337, N3457, N6356, N6591);
xor XOR2 (N9352, N9351, N4088);
buf BUF1 (N9353, N9345);
xor XOR2 (N9354, N9348, N4743);
and AND2 (N9355, N9352, N1465);
nor NOR4 (N9356, N9334, N5487, N4951, N8909);
buf BUF1 (N9357, N9343);
nand NAND2 (N9358, N9353, N8798);
nor NOR2 (N9359, N9341, N2216);
and AND4 (N9360, N9358, N6056, N2757, N8494);
buf BUF1 (N9361, N9357);
or OR3 (N9362, N9359, N5229, N7641);
and AND4 (N9363, N9356, N1393, N4711, N4707);
xor XOR2 (N9364, N9363, N3624);
nand NAND4 (N9365, N9362, N1084, N3011, N5984);
and AND2 (N9366, N9355, N4434);
nor NOR2 (N9367, N9331, N1836);
or OR4 (N9368, N9367, N3461, N6542, N7278);
nor NOR4 (N9369, N9361, N698, N1809, N9071);
buf BUF1 (N9370, N9349);
xor XOR2 (N9371, N9365, N8178);
or OR2 (N9372, N9354, N3748);
or OR4 (N9373, N9350, N6657, N3681, N1045);
nand NAND3 (N9374, N9370, N9337, N4032);
nor NOR4 (N9375, N9360, N5004, N7871, N28);
nor NOR3 (N9376, N9364, N4371, N5109);
nor NOR3 (N9377, N9368, N3800, N6581);
buf BUF1 (N9378, N9374);
nand NAND4 (N9379, N9376, N2133, N6956, N8427);
buf BUF1 (N9380, N9373);
not NOT1 (N9381, N9378);
nor NOR2 (N9382, N9381, N2480);
nor NOR2 (N9383, N9332, N614);
or OR4 (N9384, N9375, N8763, N2021, N7586);
buf BUF1 (N9385, N9384);
buf BUF1 (N9386, N9371);
buf BUF1 (N9387, N9386);
and AND2 (N9388, N9369, N8862);
and AND2 (N9389, N9385, N7704);
not NOT1 (N9390, N9366);
and AND2 (N9391, N9382, N3271);
buf BUF1 (N9392, N9380);
and AND3 (N9393, N9390, N2555, N5858);
nand NAND2 (N9394, N9393, N4532);
and AND4 (N9395, N9389, N4563, N4319, N1557);
xor XOR2 (N9396, N9391, N9348);
nand NAND2 (N9397, N9372, N479);
nor NOR2 (N9398, N9383, N2209);
xor XOR2 (N9399, N9398, N4398);
and AND2 (N9400, N9399, N6918);
xor XOR2 (N9401, N9396, N1433);
xor XOR2 (N9402, N9401, N1749);
nor NOR3 (N9403, N9397, N3149, N871);
buf BUF1 (N9404, N9377);
buf BUF1 (N9405, N9404);
xor XOR2 (N9406, N9405, N4473);
buf BUF1 (N9407, N9394);
nor NOR2 (N9408, N9379, N7801);
nand NAND4 (N9409, N9406, N2298, N9152, N3348);
or OR4 (N9410, N9402, N9358, N8505, N9042);
buf BUF1 (N9411, N9403);
or OR3 (N9412, N9395, N62, N8229);
xor XOR2 (N9413, N9407, N1956);
xor XOR2 (N9414, N9400, N2284);
xor XOR2 (N9415, N9387, N6739);
buf BUF1 (N9416, N9392);
not NOT1 (N9417, N9413);
and AND3 (N9418, N9388, N4983, N6860);
nor NOR3 (N9419, N9410, N1919, N7845);
nand NAND3 (N9420, N9416, N5781, N587);
nor NOR2 (N9421, N9417, N3367);
nand NAND3 (N9422, N9408, N3431, N4394);
buf BUF1 (N9423, N9414);
not NOT1 (N9424, N9418);
and AND2 (N9425, N9411, N4338);
or OR4 (N9426, N9423, N79, N281, N6220);
buf BUF1 (N9427, N9424);
and AND3 (N9428, N9409, N2082, N4971);
nand NAND2 (N9429, N9420, N298);
and AND4 (N9430, N9427, N1515, N4896, N8208);
xor XOR2 (N9431, N9422, N7715);
xor XOR2 (N9432, N9426, N9250);
and AND2 (N9433, N9432, N6042);
nor NOR2 (N9434, N9433, N5410);
buf BUF1 (N9435, N9419);
nand NAND3 (N9436, N9415, N7700, N7800);
buf BUF1 (N9437, N9429);
xor XOR2 (N9438, N9436, N4435);
nand NAND2 (N9439, N9421, N8322);
xor XOR2 (N9440, N9434, N3195);
and AND3 (N9441, N9425, N3776, N508);
or OR4 (N9442, N9431, N6377, N4623, N9157);
buf BUF1 (N9443, N9430);
or OR4 (N9444, N9428, N1766, N3552, N3172);
and AND3 (N9445, N9442, N7236, N5377);
nor NOR3 (N9446, N9438, N7607, N7462);
nand NAND4 (N9447, N9446, N3037, N8907, N5171);
nand NAND2 (N9448, N9441, N4605);
not NOT1 (N9449, N9437);
or OR4 (N9450, N9443, N7129, N7118, N814);
nor NOR3 (N9451, N9412, N3947, N4052);
nand NAND3 (N9452, N9450, N4522, N3972);
and AND4 (N9453, N9440, N3552, N2370, N3308);
or OR4 (N9454, N9449, N6428, N7725, N5986);
nor NOR3 (N9455, N9439, N8895, N2131);
not NOT1 (N9456, N9453);
nand NAND2 (N9457, N9456, N5825);
and AND2 (N9458, N9452, N5835);
xor XOR2 (N9459, N9444, N2811);
nor NOR4 (N9460, N9448, N4897, N6767, N6603);
nor NOR2 (N9461, N9445, N8283);
buf BUF1 (N9462, N9458);
nand NAND4 (N9463, N9435, N7672, N8790, N6933);
nand NAND3 (N9464, N9463, N5756, N3956);
nand NAND3 (N9465, N9454, N4648, N7786);
not NOT1 (N9466, N9464);
or OR4 (N9467, N9451, N8456, N5921, N8711);
not NOT1 (N9468, N9460);
buf BUF1 (N9469, N9447);
not NOT1 (N9470, N9469);
xor XOR2 (N9471, N9462, N3183);
buf BUF1 (N9472, N9470);
buf BUF1 (N9473, N9468);
or OR4 (N9474, N9465, N429, N1581, N7534);
or OR3 (N9475, N9473, N8287, N3616);
and AND3 (N9476, N9472, N2858, N4677);
not NOT1 (N9477, N9461);
or OR2 (N9478, N9474, N3033);
buf BUF1 (N9479, N9457);
and AND4 (N9480, N9477, N4711, N8203, N3308);
and AND4 (N9481, N9475, N4302, N5778, N5575);
xor XOR2 (N9482, N9476, N3970);
buf BUF1 (N9483, N9466);
buf BUF1 (N9484, N9483);
nand NAND3 (N9485, N9471, N7513, N3939);
or OR2 (N9486, N9481, N1674);
and AND4 (N9487, N9478, N4674, N6828, N7649);
nand NAND4 (N9488, N9479, N3483, N4834, N8650);
not NOT1 (N9489, N9486);
not NOT1 (N9490, N9480);
nand NAND4 (N9491, N9467, N3640, N3930, N7852);
buf BUF1 (N9492, N9489);
nor NOR4 (N9493, N9487, N6641, N3731, N9048);
nor NOR4 (N9494, N9482, N7161, N3465, N8051);
buf BUF1 (N9495, N9488);
nand NAND2 (N9496, N9493, N4345);
nand NAND4 (N9497, N9459, N8621, N2300, N1273);
buf BUF1 (N9498, N9495);
nand NAND2 (N9499, N9455, N7579);
nor NOR4 (N9500, N9494, N6061, N2956, N6157);
nor NOR3 (N9501, N9492, N283, N4409);
or OR3 (N9502, N9496, N5893, N1646);
and AND2 (N9503, N9499, N4201);
nor NOR4 (N9504, N9502, N6681, N1605, N6170);
nand NAND4 (N9505, N9503, N7545, N7885, N104);
xor XOR2 (N9506, N9501, N4111);
nand NAND4 (N9507, N9497, N7346, N4710, N6649);
and AND4 (N9508, N9498, N5154, N4317, N4153);
not NOT1 (N9509, N9505);
buf BUF1 (N9510, N9506);
not NOT1 (N9511, N9510);
and AND2 (N9512, N9507, N2356);
or OR3 (N9513, N9509, N8861, N3055);
nor NOR2 (N9514, N9490, N1963);
not NOT1 (N9515, N9512);
nor NOR3 (N9516, N9511, N1737, N7825);
nor NOR3 (N9517, N9485, N4474, N3883);
nor NOR4 (N9518, N9513, N2613, N5356, N1955);
nor NOR3 (N9519, N9518, N7769, N4975);
xor XOR2 (N9520, N9508, N4925);
or OR4 (N9521, N9515, N4409, N7473, N3871);
buf BUF1 (N9522, N9514);
or OR3 (N9523, N9521, N2383, N1507);
nand NAND2 (N9524, N9484, N6189);
xor XOR2 (N9525, N9516, N4720);
nand NAND4 (N9526, N9500, N1991, N8437, N2814);
and AND4 (N9527, N9491, N6473, N6751, N7494);
not NOT1 (N9528, N9524);
or OR4 (N9529, N9525, N2512, N1233, N2046);
and AND4 (N9530, N9523, N4424, N2138, N3452);
nor NOR2 (N9531, N9517, N7768);
not NOT1 (N9532, N9531);
nand NAND4 (N9533, N9530, N5007, N7429, N8948);
xor XOR2 (N9534, N9528, N3856);
or OR3 (N9535, N9533, N5247, N2564);
or OR3 (N9536, N9534, N174, N8177);
or OR2 (N9537, N9522, N855);
nor NOR2 (N9538, N9519, N6376);
nor NOR4 (N9539, N9527, N3728, N9164, N245);
or OR2 (N9540, N9536, N6150);
nor NOR3 (N9541, N9539, N1265, N4379);
not NOT1 (N9542, N9504);
nor NOR3 (N9543, N9520, N1148, N7026);
nand NAND4 (N9544, N9526, N4015, N8506, N968);
buf BUF1 (N9545, N9538);
not NOT1 (N9546, N9529);
and AND2 (N9547, N9541, N5884);
buf BUF1 (N9548, N9540);
nor NOR2 (N9549, N9547, N9334);
not NOT1 (N9550, N9548);
nand NAND4 (N9551, N9543, N934, N7260, N6893);
nor NOR3 (N9552, N9532, N1254, N4029);
nand NAND4 (N9553, N9542, N1685, N8613, N1303);
buf BUF1 (N9554, N9550);
nand NAND4 (N9555, N9554, N744, N2313, N5733);
nand NAND2 (N9556, N9553, N6656);
buf BUF1 (N9557, N9552);
not NOT1 (N9558, N9535);
or OR3 (N9559, N9557, N1701, N611);
buf BUF1 (N9560, N9555);
nor NOR3 (N9561, N9560, N7814, N2846);
nor NOR3 (N9562, N9558, N6626, N8031);
nand NAND3 (N9563, N9559, N4114, N7225);
and AND4 (N9564, N9563, N5199, N7905, N5508);
and AND3 (N9565, N9546, N4450, N4767);
nor NOR4 (N9566, N9551, N8243, N5263, N1004);
nand NAND3 (N9567, N9544, N8836, N5756);
and AND4 (N9568, N9562, N2704, N2718, N5767);
nand NAND2 (N9569, N9565, N2990);
nor NOR2 (N9570, N9549, N5899);
nand NAND3 (N9571, N9566, N6131, N6392);
and AND3 (N9572, N9537, N8891, N924);
or OR3 (N9573, N9570, N7803, N1191);
and AND2 (N9574, N9561, N18);
nor NOR2 (N9575, N9573, N1806);
and AND2 (N9576, N9545, N8396);
not NOT1 (N9577, N9575);
xor XOR2 (N9578, N9576, N683);
buf BUF1 (N9579, N9577);
nand NAND2 (N9580, N9556, N1020);
or OR2 (N9581, N9574, N1667);
buf BUF1 (N9582, N9567);
not NOT1 (N9583, N9571);
nor NOR4 (N9584, N9564, N9421, N2104, N4116);
nor NOR3 (N9585, N9582, N1407, N2417);
nand NAND4 (N9586, N9581, N8695, N8078, N4753);
nand NAND2 (N9587, N9569, N1158);
xor XOR2 (N9588, N9585, N1763);
and AND2 (N9589, N9578, N3529);
or OR4 (N9590, N9587, N3521, N4547, N513);
not NOT1 (N9591, N9572);
xor XOR2 (N9592, N9568, N1445);
buf BUF1 (N9593, N9583);
and AND4 (N9594, N9589, N3466, N1195, N8823);
nor NOR3 (N9595, N9592, N8313, N8583);
nand NAND2 (N9596, N9591, N9275);
nand NAND3 (N9597, N9595, N6037, N8839);
nand NAND4 (N9598, N9580, N3924, N5441, N104);
nor NOR3 (N9599, N9584, N8284, N3843);
nand NAND4 (N9600, N9588, N3918, N39, N1977);
buf BUF1 (N9601, N9596);
or OR4 (N9602, N9590, N9004, N1979, N2176);
not NOT1 (N9603, N9598);
buf BUF1 (N9604, N9594);
buf BUF1 (N9605, N9600);
nand NAND2 (N9606, N9586, N8989);
buf BUF1 (N9607, N9605);
not NOT1 (N9608, N9607);
and AND3 (N9609, N9599, N2684, N8762);
not NOT1 (N9610, N9603);
nor NOR3 (N9611, N9608, N1057, N9409);
and AND4 (N9612, N9601, N3111, N734, N4339);
and AND2 (N9613, N9597, N7637);
and AND3 (N9614, N9604, N4462, N6283);
or OR3 (N9615, N9611, N8856, N2176);
and AND4 (N9616, N9614, N9131, N8703, N1904);
nor NOR4 (N9617, N9579, N2230, N6322, N7902);
and AND3 (N9618, N9613, N5031, N519);
nand NAND2 (N9619, N9606, N166);
not NOT1 (N9620, N9618);
buf BUF1 (N9621, N9602);
and AND3 (N9622, N9612, N6323, N477);
nand NAND3 (N9623, N9617, N8364, N3137);
nand NAND3 (N9624, N9610, N385, N2938);
buf BUF1 (N9625, N9619);
or OR4 (N9626, N9620, N8385, N4747, N2997);
nand NAND3 (N9627, N9624, N2295, N2674);
xor XOR2 (N9628, N9615, N1652);
and AND3 (N9629, N9623, N7861, N2246);
or OR3 (N9630, N9609, N3702, N3949);
and AND2 (N9631, N9626, N173);
nand NAND4 (N9632, N9629, N2977, N2427, N7021);
xor XOR2 (N9633, N9622, N5275);
nand NAND4 (N9634, N9633, N4857, N8564, N5407);
nand NAND4 (N9635, N9616, N9249, N7040, N1859);
and AND4 (N9636, N9630, N4837, N7083, N1039);
and AND3 (N9637, N9636, N7864, N4843);
nand NAND4 (N9638, N9627, N7759, N9062, N9407);
xor XOR2 (N9639, N9632, N2681);
and AND3 (N9640, N9637, N2073, N2319);
not NOT1 (N9641, N9631);
and AND3 (N9642, N9621, N7071, N4493);
nand NAND2 (N9643, N9635, N700);
xor XOR2 (N9644, N9628, N7718);
nand NAND4 (N9645, N9641, N6325, N9191, N7368);
or OR3 (N9646, N9644, N5209, N4682);
or OR4 (N9647, N9640, N5074, N1936, N2862);
xor XOR2 (N9648, N9643, N2214);
or OR4 (N9649, N9625, N5953, N462, N669);
buf BUF1 (N9650, N9645);
buf BUF1 (N9651, N9648);
and AND2 (N9652, N9634, N7203);
buf BUF1 (N9653, N9639);
buf BUF1 (N9654, N9647);
xor XOR2 (N9655, N9654, N3548);
nor NOR4 (N9656, N9638, N6872, N6618, N5032);
or OR4 (N9657, N9653, N6138, N6492, N4335);
and AND2 (N9658, N9651, N3460);
nand NAND2 (N9659, N9652, N2343);
or OR4 (N9660, N9655, N2108, N1229, N6376);
buf BUF1 (N9661, N9659);
xor XOR2 (N9662, N9657, N3369);
nand NAND2 (N9663, N9650, N7561);
and AND3 (N9664, N9642, N1903, N6002);
nor NOR3 (N9665, N9593, N3467, N4614);
nand NAND4 (N9666, N9663, N5466, N1269, N1436);
and AND4 (N9667, N9664, N8839, N8457, N5474);
not NOT1 (N9668, N9667);
nor NOR2 (N9669, N9661, N5585);
buf BUF1 (N9670, N9665);
or OR2 (N9671, N9660, N3182);
not NOT1 (N9672, N9669);
or OR2 (N9673, N9656, N7812);
buf BUF1 (N9674, N9670);
buf BUF1 (N9675, N9662);
buf BUF1 (N9676, N9668);
nor NOR4 (N9677, N9676, N2556, N2425, N6661);
or OR2 (N9678, N9666, N2680);
nand NAND2 (N9679, N9674, N1302);
and AND2 (N9680, N9673, N5505);
buf BUF1 (N9681, N9671);
not NOT1 (N9682, N9678);
buf BUF1 (N9683, N9646);
and AND3 (N9684, N9675, N2592, N3610);
and AND4 (N9685, N9658, N6557, N5920, N4436);
nand NAND2 (N9686, N9672, N3266);
or OR3 (N9687, N9649, N2903, N5673);
xor XOR2 (N9688, N9684, N829);
and AND4 (N9689, N9682, N2861, N6546, N9255);
not NOT1 (N9690, N9683);
or OR4 (N9691, N9685, N9010, N7588, N1740);
not NOT1 (N9692, N9680);
not NOT1 (N9693, N9691);
nor NOR4 (N9694, N9686, N6640, N1471, N8779);
buf BUF1 (N9695, N9690);
buf BUF1 (N9696, N9687);
not NOT1 (N9697, N9681);
nor NOR3 (N9698, N9697, N806, N5909);
nand NAND4 (N9699, N9689, N1712, N4357, N7979);
not NOT1 (N9700, N9677);
nand NAND2 (N9701, N9696, N3007);
nand NAND2 (N9702, N9692, N7351);
nand NAND3 (N9703, N9702, N599, N5332);
not NOT1 (N9704, N9695);
and AND3 (N9705, N9698, N9153, N6986);
not NOT1 (N9706, N9679);
buf BUF1 (N9707, N9699);
xor XOR2 (N9708, N9701, N9375);
nor NOR3 (N9709, N9706, N534, N7318);
nand NAND4 (N9710, N9688, N2221, N2720, N6917);
buf BUF1 (N9711, N9703);
buf BUF1 (N9712, N9705);
nand NAND4 (N9713, N9694, N6761, N9397, N558);
buf BUF1 (N9714, N9707);
nor NOR3 (N9715, N9708, N6561, N9688);
nor NOR4 (N9716, N9712, N4724, N472, N2332);
not NOT1 (N9717, N9704);
or OR2 (N9718, N9714, N4210);
or OR2 (N9719, N9713, N7282);
buf BUF1 (N9720, N9717);
nor NOR4 (N9721, N9716, N3761, N8572, N3674);
not NOT1 (N9722, N9720);
xor XOR2 (N9723, N9722, N5803);
and AND4 (N9724, N9693, N9483, N8923, N442);
nor NOR2 (N9725, N9718, N1836);
nor NOR4 (N9726, N9721, N7828, N3207, N8340);
buf BUF1 (N9727, N9711);
xor XOR2 (N9728, N9726, N7840);
not NOT1 (N9729, N9709);
buf BUF1 (N9730, N9723);
and AND3 (N9731, N9729, N7766, N6929);
nand NAND4 (N9732, N9724, N266, N8954, N1419);
xor XOR2 (N9733, N9731, N4039);
nor NOR3 (N9734, N9733, N418, N7641);
nand NAND3 (N9735, N9734, N6432, N4254);
and AND4 (N9736, N9710, N975, N5128, N1113);
and AND4 (N9737, N9730, N5081, N9667, N4872);
nor NOR4 (N9738, N9735, N9693, N3314, N4509);
xor XOR2 (N9739, N9737, N6785);
nand NAND3 (N9740, N9732, N3402, N9116);
nor NOR4 (N9741, N9725, N7844, N4974, N3005);
buf BUF1 (N9742, N9739);
not NOT1 (N9743, N9719);
and AND2 (N9744, N9738, N7747);
xor XOR2 (N9745, N9727, N9361);
not NOT1 (N9746, N9741);
and AND2 (N9747, N9728, N3138);
xor XOR2 (N9748, N9715, N8688);
nor NOR3 (N9749, N9745, N1313, N8647);
buf BUF1 (N9750, N9740);
buf BUF1 (N9751, N9747);
not NOT1 (N9752, N9748);
xor XOR2 (N9753, N9700, N1556);
buf BUF1 (N9754, N9752);
not NOT1 (N9755, N9750);
not NOT1 (N9756, N9751);
nand NAND2 (N9757, N9746, N2132);
or OR3 (N9758, N9755, N8978, N1059);
not NOT1 (N9759, N9743);
and AND2 (N9760, N9758, N3057);
xor XOR2 (N9761, N9754, N1520);
buf BUF1 (N9762, N9757);
xor XOR2 (N9763, N9753, N3898);
buf BUF1 (N9764, N9760);
nor NOR2 (N9765, N9736, N2730);
buf BUF1 (N9766, N9764);
and AND2 (N9767, N9744, N1529);
buf BUF1 (N9768, N9756);
xor XOR2 (N9769, N9768, N1328);
not NOT1 (N9770, N9763);
not NOT1 (N9771, N9769);
xor XOR2 (N9772, N9761, N9043);
nor NOR2 (N9773, N9742, N4280);
and AND2 (N9774, N9767, N1668);
xor XOR2 (N9775, N9762, N5946);
or OR3 (N9776, N9771, N8453, N2232);
not NOT1 (N9777, N9774);
xor XOR2 (N9778, N9773, N2287);
or OR3 (N9779, N9749, N2707, N8384);
or OR2 (N9780, N9759, N1799);
buf BUF1 (N9781, N9778);
nor NOR2 (N9782, N9777, N9125);
buf BUF1 (N9783, N9772);
nand NAND4 (N9784, N9776, N5510, N7324, N8618);
or OR4 (N9785, N9783, N3352, N2572, N1249);
nand NAND3 (N9786, N9784, N2212, N3497);
not NOT1 (N9787, N9785);
not NOT1 (N9788, N9781);
not NOT1 (N9789, N9766);
buf BUF1 (N9790, N9775);
and AND4 (N9791, N9780, N504, N6618, N4688);
nand NAND4 (N9792, N9789, N1559, N2525, N5787);
nand NAND3 (N9793, N9790, N6223, N3387);
nand NAND4 (N9794, N9787, N1310, N1929, N1871);
and AND3 (N9795, N9786, N6130, N8193);
nand NAND2 (N9796, N9793, N4548);
or OR3 (N9797, N9796, N2130, N3701);
xor XOR2 (N9798, N9797, N3502);
xor XOR2 (N9799, N9765, N251);
and AND2 (N9800, N9799, N7876);
xor XOR2 (N9801, N9788, N7960);
buf BUF1 (N9802, N9770);
nor NOR2 (N9803, N9795, N4417);
nand NAND3 (N9804, N9779, N4833, N5453);
nor NOR2 (N9805, N9804, N129);
not NOT1 (N9806, N9802);
nor NOR3 (N9807, N9806, N1506, N9071);
or OR4 (N9808, N9792, N5484, N7311, N4910);
xor XOR2 (N9809, N9805, N4480);
nand NAND2 (N9810, N9791, N2434);
or OR2 (N9811, N9808, N3574);
nand NAND4 (N9812, N9807, N4756, N5721, N4926);
nor NOR4 (N9813, N9810, N3082, N2323, N5066);
nor NOR2 (N9814, N9809, N1118);
buf BUF1 (N9815, N9798);
nand NAND4 (N9816, N9803, N1072, N4152, N223);
not NOT1 (N9817, N9812);
nor NOR2 (N9818, N9811, N1755);
nand NAND2 (N9819, N9815, N2991);
nand NAND3 (N9820, N9813, N5025, N2452);
nor NOR3 (N9821, N9818, N7587, N6470);
nor NOR4 (N9822, N9782, N8183, N1342, N1931);
nand NAND3 (N9823, N9819, N9288, N3624);
buf BUF1 (N9824, N9821);
or OR4 (N9825, N9794, N2970, N8900, N9677);
not NOT1 (N9826, N9814);
nor NOR3 (N9827, N9816, N2170, N4776);
and AND2 (N9828, N9825, N5585);
not NOT1 (N9829, N9827);
and AND4 (N9830, N9826, N2054, N390, N3601);
and AND3 (N9831, N9820, N7012, N2644);
nor NOR4 (N9832, N9800, N2830, N4917, N9520);
and AND4 (N9833, N9828, N8239, N9252, N7722);
xor XOR2 (N9834, N9832, N8833);
buf BUF1 (N9835, N9834);
and AND3 (N9836, N9833, N9637, N5529);
nand NAND3 (N9837, N9824, N9088, N8132);
xor XOR2 (N9838, N9823, N3620);
buf BUF1 (N9839, N9837);
and AND3 (N9840, N9831, N1337, N95);
and AND4 (N9841, N9839, N7649, N1912, N6885);
and AND3 (N9842, N9840, N556, N2707);
or OR2 (N9843, N9835, N285);
nand NAND2 (N9844, N9801, N8221);
not NOT1 (N9845, N9817);
not NOT1 (N9846, N9822);
nor NOR4 (N9847, N9836, N1278, N7573, N2879);
and AND4 (N9848, N9846, N9289, N1313, N1175);
xor XOR2 (N9849, N9843, N3154);
nor NOR4 (N9850, N9847, N2228, N3354, N1688);
not NOT1 (N9851, N9850);
xor XOR2 (N9852, N9851, N3168);
nand NAND2 (N9853, N9845, N3599);
nor NOR2 (N9854, N9844, N8606);
nand NAND4 (N9855, N9829, N6110, N5402, N6057);
xor XOR2 (N9856, N9854, N3574);
xor XOR2 (N9857, N9841, N493);
xor XOR2 (N9858, N9856, N3258);
or OR3 (N9859, N9842, N3372, N3583);
nor NOR4 (N9860, N9858, N2994, N794, N1384);
or OR3 (N9861, N9848, N2741, N7998);
and AND3 (N9862, N9861, N2128, N6129);
buf BUF1 (N9863, N9862);
nand NAND4 (N9864, N9855, N6820, N6711, N9794);
buf BUF1 (N9865, N9860);
not NOT1 (N9866, N9852);
buf BUF1 (N9867, N9857);
and AND3 (N9868, N9838, N4368, N7685);
or OR2 (N9869, N9867, N4855);
nand NAND2 (N9870, N9869, N912);
nand NAND3 (N9871, N9863, N3398, N4421);
nand NAND4 (N9872, N9871, N3746, N6544, N2174);
xor XOR2 (N9873, N9853, N2512);
nor NOR2 (N9874, N9866, N2587);
and AND4 (N9875, N9874, N4875, N6811, N10);
xor XOR2 (N9876, N9870, N7128);
xor XOR2 (N9877, N9865, N5378);
buf BUF1 (N9878, N9872);
xor XOR2 (N9879, N9878, N2426);
not NOT1 (N9880, N9875);
nor NOR2 (N9881, N9859, N3875);
nor NOR4 (N9882, N9864, N9791, N2014, N2872);
nand NAND2 (N9883, N9849, N2994);
or OR2 (N9884, N9880, N7475);
or OR4 (N9885, N9877, N9204, N166, N1426);
nand NAND4 (N9886, N9883, N3678, N303, N8448);
nor NOR2 (N9887, N9830, N9690);
nand NAND4 (N9888, N9886, N387, N1472, N3648);
xor XOR2 (N9889, N9882, N1003);
nor NOR2 (N9890, N9881, N7782);
xor XOR2 (N9891, N9879, N1552);
nor NOR4 (N9892, N9868, N7726, N7434, N6825);
not NOT1 (N9893, N9889);
nor NOR3 (N9894, N9888, N2425, N2199);
not NOT1 (N9895, N9891);
not NOT1 (N9896, N9876);
not NOT1 (N9897, N9873);
and AND3 (N9898, N9892, N3529, N8385);
or OR2 (N9899, N9897, N4933);
xor XOR2 (N9900, N9884, N7840);
nor NOR2 (N9901, N9898, N1451);
xor XOR2 (N9902, N9899, N391);
not NOT1 (N9903, N9887);
nor NOR3 (N9904, N9894, N8882, N2992);
buf BUF1 (N9905, N9896);
buf BUF1 (N9906, N9905);
xor XOR2 (N9907, N9893, N5568);
and AND3 (N9908, N9890, N9270, N2022);
and AND2 (N9909, N9904, N3722);
or OR3 (N9910, N9895, N4609, N2513);
and AND4 (N9911, N9906, N125, N5921, N2657);
not NOT1 (N9912, N9907);
or OR3 (N9913, N9902, N1079, N408);
nand NAND4 (N9914, N9910, N9292, N5956, N4830);
nand NAND3 (N9915, N9903, N8799, N6431);
nor NOR4 (N9916, N9915, N8, N2405, N2748);
xor XOR2 (N9917, N9901, N9429);
or OR4 (N9918, N9900, N6963, N4, N4805);
or OR2 (N9919, N9912, N8679);
and AND2 (N9920, N9918, N4850);
nand NAND4 (N9921, N9913, N2709, N8952, N5424);
or OR3 (N9922, N9909, N8100, N1529);
xor XOR2 (N9923, N9922, N1978);
buf BUF1 (N9924, N9923);
buf BUF1 (N9925, N9916);
xor XOR2 (N9926, N9919, N6833);
nor NOR2 (N9927, N9885, N5156);
or OR2 (N9928, N9925, N4351);
nor NOR2 (N9929, N9911, N5055);
nand NAND4 (N9930, N9928, N9029, N3404, N2636);
nor NOR3 (N9931, N9917, N4712, N4869);
nand NAND3 (N9932, N9926, N8296, N2848);
xor XOR2 (N9933, N9924, N5001);
not NOT1 (N9934, N9927);
nand NAND2 (N9935, N9933, N4008);
or OR2 (N9936, N9929, N9847);
or OR4 (N9937, N9931, N7997, N1493, N339);
buf BUF1 (N9938, N9920);
buf BUF1 (N9939, N9936);
or OR3 (N9940, N9921, N125, N211);
xor XOR2 (N9941, N9908, N7968);
xor XOR2 (N9942, N9930, N1183);
nor NOR2 (N9943, N9939, N7469);
buf BUF1 (N9944, N9914);
xor XOR2 (N9945, N9937, N5547);
buf BUF1 (N9946, N9943);
buf BUF1 (N9947, N9938);
xor XOR2 (N9948, N9941, N2776);
and AND4 (N9949, N9940, N8977, N5275, N1941);
and AND4 (N9950, N9945, N2233, N7156, N6080);
and AND3 (N9951, N9946, N2028, N7261);
nor NOR2 (N9952, N9948, N7622);
nor NOR4 (N9953, N9935, N1981, N3303, N5065);
nand NAND3 (N9954, N9949, N4726, N4944);
buf BUF1 (N9955, N9932);
xor XOR2 (N9956, N9954, N4818);
not NOT1 (N9957, N9956);
nand NAND2 (N9958, N9955, N3961);
buf BUF1 (N9959, N9958);
or OR2 (N9960, N9959, N5046);
or OR4 (N9961, N9942, N7433, N7092, N3788);
nor NOR4 (N9962, N9934, N284, N4953, N5787);
nor NOR3 (N9963, N9962, N3361, N603);
buf BUF1 (N9964, N9952);
nand NAND3 (N9965, N9950, N4260, N3896);
or OR2 (N9966, N9957, N245);
buf BUF1 (N9967, N9966);
nor NOR4 (N9968, N9967, N8112, N4659, N4788);
nor NOR2 (N9969, N9947, N5295);
xor XOR2 (N9970, N9960, N7361);
not NOT1 (N9971, N9965);
or OR4 (N9972, N9951, N1025, N2251, N9494);
xor XOR2 (N9973, N9972, N9329);
nor NOR4 (N9974, N9968, N6076, N3686, N4937);
not NOT1 (N9975, N9970);
buf BUF1 (N9976, N9971);
or OR3 (N9977, N9973, N904, N5848);
not NOT1 (N9978, N9974);
or OR4 (N9979, N9976, N808, N9628, N8909);
buf BUF1 (N9980, N9953);
or OR2 (N9981, N9980, N3251);
and AND4 (N9982, N9944, N3384, N3804, N988);
nor NOR3 (N9983, N9978, N2838, N6298);
nand NAND3 (N9984, N9977, N8764, N2376);
xor XOR2 (N9985, N9981, N5667);
and AND3 (N9986, N9975, N2218, N1734);
nor NOR2 (N9987, N9964, N6210);
nand NAND3 (N9988, N9979, N4806, N1927);
and AND4 (N9989, N9984, N8956, N2907, N9473);
buf BUF1 (N9990, N9983);
not NOT1 (N9991, N9961);
not NOT1 (N9992, N9987);
not NOT1 (N9993, N9963);
xor XOR2 (N9994, N9985, N2245);
nand NAND4 (N9995, N9991, N5157, N6910, N3564);
and AND3 (N9996, N9994, N2442, N662);
or OR3 (N9997, N9982, N7325, N1898);
or OR2 (N9998, N9995, N4864);
not NOT1 (N9999, N9998);
buf BUF1 (N10000, N9993);
not NOT1 (N10001, N9990);
buf BUF1 (N10002, N9969);
or OR4 (N10003, N9986, N1016, N4361, N9012);
not NOT1 (N10004, N10002);
nor NOR2 (N10005, N10001, N198);
and AND2 (N10006, N9999, N8409);
buf BUF1 (N10007, N10003);
nand NAND2 (N10008, N10004, N6277);
or OR2 (N10009, N9997, N8848);
nand NAND2 (N10010, N9992, N9255);
or OR2 (N10011, N10009, N4002);
xor XOR2 (N10012, N10011, N8679);
nor NOR3 (N10013, N9996, N9095, N6077);
xor XOR2 (N10014, N10013, N8909);
nand NAND3 (N10015, N9988, N3946, N4030);
not NOT1 (N10016, N10008);
not NOT1 (N10017, N10005);
xor XOR2 (N10018, N9989, N1294);
nand NAND2 (N10019, N10014, N2084);
nand NAND4 (N10020, N10018, N8240, N1778, N4843);
xor XOR2 (N10021, N10000, N1334);
buf BUF1 (N10022, N10012);
xor XOR2 (N10023, N10020, N736);
xor XOR2 (N10024, N10021, N3162);
or OR4 (N10025, N10007, N3189, N7252, N9675);
buf BUF1 (N10026, N10019);
not NOT1 (N10027, N10010);
nor NOR3 (N10028, N10006, N9883, N3966);
nand NAND3 (N10029, N10022, N6683, N4155);
and AND2 (N10030, N10016, N6165);
buf BUF1 (N10031, N10028);
not NOT1 (N10032, N10031);
xor XOR2 (N10033, N10015, N3423);
nor NOR2 (N10034, N10024, N1825);
not NOT1 (N10035, N10025);
nand NAND4 (N10036, N10032, N8500, N2934, N1005);
not NOT1 (N10037, N10035);
not NOT1 (N10038, N10017);
xor XOR2 (N10039, N10033, N8802);
or OR2 (N10040, N10034, N7033);
or OR2 (N10041, N10026, N2471);
and AND2 (N10042, N10027, N1789);
xor XOR2 (N10043, N10029, N8636);
not NOT1 (N10044, N10041);
buf BUF1 (N10045, N10043);
xor XOR2 (N10046, N10023, N3258);
or OR3 (N10047, N10044, N1938, N8755);
and AND2 (N10048, N10042, N9383);
or OR2 (N10049, N10045, N2336);
xor XOR2 (N10050, N10038, N1064);
not NOT1 (N10051, N10048);
buf BUF1 (N10052, N10051);
or OR2 (N10053, N10050, N3854);
not NOT1 (N10054, N10040);
or OR2 (N10055, N10053, N7756);
buf BUF1 (N10056, N10052);
nor NOR3 (N10057, N10046, N4290, N330);
and AND3 (N10058, N10030, N4861, N8406);
nor NOR3 (N10059, N10057, N7633, N86);
nor NOR4 (N10060, N10054, N650, N6604, N4438);
buf BUF1 (N10061, N10060);
nand NAND4 (N10062, N10061, N3175, N9994, N7079);
not NOT1 (N10063, N10059);
nand NAND3 (N10064, N10047, N9689, N2276);
nand NAND4 (N10065, N10036, N7876, N5759, N3670);
or OR2 (N10066, N10039, N5261);
or OR4 (N10067, N10049, N6517, N8909, N8184);
nor NOR3 (N10068, N10056, N9328, N4347);
not NOT1 (N10069, N10066);
not NOT1 (N10070, N10064);
not NOT1 (N10071, N10069);
nand NAND2 (N10072, N10055, N4534);
and AND2 (N10073, N10071, N5934);
nor NOR4 (N10074, N10058, N8382, N9809, N6009);
nand NAND3 (N10075, N10070, N1297, N7666);
buf BUF1 (N10076, N10074);
nor NOR3 (N10077, N10062, N7565, N7304);
xor XOR2 (N10078, N10037, N1813);
nand NAND3 (N10079, N10077, N7185, N4956);
nor NOR4 (N10080, N10067, N346, N8525, N5095);
nand NAND3 (N10081, N10072, N1071, N1332);
and AND2 (N10082, N10063, N2436);
and AND3 (N10083, N10078, N2765, N9884);
or OR4 (N10084, N10076, N8147, N7088, N3274);
nand NAND3 (N10085, N10065, N1869, N8127);
buf BUF1 (N10086, N10084);
nor NOR4 (N10087, N10075, N7018, N3522, N2350);
or OR2 (N10088, N10082, N6458);
xor XOR2 (N10089, N10068, N3026);
nand NAND3 (N10090, N10083, N4359, N2060);
and AND4 (N10091, N10087, N2613, N3771, N6603);
not NOT1 (N10092, N10079);
nand NAND4 (N10093, N10081, N289, N5953, N2091);
not NOT1 (N10094, N10085);
and AND2 (N10095, N10094, N1996);
and AND3 (N10096, N10093, N748, N9091);
buf BUF1 (N10097, N10095);
not NOT1 (N10098, N10088);
buf BUF1 (N10099, N10089);
or OR2 (N10100, N10098, N8810);
not NOT1 (N10101, N10086);
not NOT1 (N10102, N10080);
xor XOR2 (N10103, N10091, N9346);
and AND3 (N10104, N10102, N950, N6117);
buf BUF1 (N10105, N10104);
nand NAND2 (N10106, N10073, N4114);
or OR4 (N10107, N10099, N2887, N7965, N1060);
buf BUF1 (N10108, N10105);
not NOT1 (N10109, N10101);
not NOT1 (N10110, N10092);
and AND2 (N10111, N10109, N10057);
xor XOR2 (N10112, N10110, N3834);
and AND2 (N10113, N10100, N10027);
not NOT1 (N10114, N10106);
or OR2 (N10115, N10097, N65);
buf BUF1 (N10116, N10114);
or OR3 (N10117, N10116, N8732, N9261);
and AND3 (N10118, N10103, N4148, N1295);
nor NOR4 (N10119, N10113, N5907, N699, N1618);
nand NAND4 (N10120, N10115, N3602, N8129, N2701);
xor XOR2 (N10121, N10117, N9226);
nand NAND4 (N10122, N10108, N2214, N5611, N4107);
buf BUF1 (N10123, N10121);
nand NAND2 (N10124, N10107, N6226);
buf BUF1 (N10125, N10123);
nor NOR4 (N10126, N10096, N6447, N1021, N4867);
not NOT1 (N10127, N10120);
nor NOR2 (N10128, N10122, N8816);
nor NOR2 (N10129, N10124, N6022);
nand NAND3 (N10130, N10090, N4419, N795);
and AND2 (N10131, N10111, N6312);
or OR3 (N10132, N10129, N7794, N4095);
and AND3 (N10133, N10126, N8483, N8845);
nand NAND2 (N10134, N10128, N2207);
nand NAND2 (N10135, N10125, N6705);
or OR4 (N10136, N10133, N5977, N8179, N580);
nand NAND3 (N10137, N10118, N5632, N10105);
xor XOR2 (N10138, N10119, N8037);
nor NOR4 (N10139, N10131, N6158, N6136, N3611);
xor XOR2 (N10140, N10132, N3801);
nor NOR2 (N10141, N10134, N6195);
and AND2 (N10142, N10136, N8448);
nand NAND3 (N10143, N10130, N2429, N4484);
not NOT1 (N10144, N10127);
not NOT1 (N10145, N10135);
or OR4 (N10146, N10142, N6614, N7856, N3199);
xor XOR2 (N10147, N10146, N165);
buf BUF1 (N10148, N10144);
nand NAND3 (N10149, N10141, N3880, N4890);
nor NOR2 (N10150, N10138, N2064);
not NOT1 (N10151, N10145);
nor NOR2 (N10152, N10148, N4332);
buf BUF1 (N10153, N10143);
or OR3 (N10154, N10139, N6070, N2397);
nor NOR2 (N10155, N10150, N278);
not NOT1 (N10156, N10147);
nand NAND4 (N10157, N10155, N9075, N8717, N6454);
buf BUF1 (N10158, N10153);
nor NOR2 (N10159, N10158, N2965);
or OR3 (N10160, N10159, N6864, N8252);
xor XOR2 (N10161, N10156, N5070);
or OR4 (N10162, N10137, N6782, N1426, N3395);
or OR2 (N10163, N10161, N4265);
and AND4 (N10164, N10152, N9911, N898, N7614);
xor XOR2 (N10165, N10149, N503);
and AND4 (N10166, N10112, N4045, N9142, N6448);
nand NAND2 (N10167, N10164, N6735);
buf BUF1 (N10168, N10154);
and AND2 (N10169, N10163, N3521);
nor NOR2 (N10170, N10168, N3975);
nand NAND3 (N10171, N10165, N1973, N5616);
xor XOR2 (N10172, N10157, N9778);
nor NOR4 (N10173, N10151, N7462, N1456, N3585);
buf BUF1 (N10174, N10160);
nand NAND3 (N10175, N10174, N280, N6462);
or OR2 (N10176, N10169, N1859);
nor NOR4 (N10177, N10162, N3364, N7463, N380);
not NOT1 (N10178, N10171);
buf BUF1 (N10179, N10166);
nor NOR3 (N10180, N10178, N766, N6053);
nor NOR3 (N10181, N10175, N4877, N987);
not NOT1 (N10182, N10167);
and AND4 (N10183, N10176, N6694, N6317, N9305);
nand NAND2 (N10184, N10182, N2786);
or OR4 (N10185, N10173, N9578, N4682, N6597);
buf BUF1 (N10186, N10184);
and AND4 (N10187, N10170, N6736, N963, N1981);
and AND4 (N10188, N10177, N3322, N5018, N3702);
buf BUF1 (N10189, N10181);
buf BUF1 (N10190, N10172);
buf BUF1 (N10191, N10187);
or OR4 (N10192, N10190, N6564, N3915, N5055);
xor XOR2 (N10193, N10183, N4423);
not NOT1 (N10194, N10186);
buf BUF1 (N10195, N10188);
nand NAND3 (N10196, N10195, N7804, N2170);
not NOT1 (N10197, N10192);
not NOT1 (N10198, N10196);
xor XOR2 (N10199, N10193, N7461);
not NOT1 (N10200, N10191);
or OR2 (N10201, N10185, N7689);
or OR3 (N10202, N10194, N9299, N4429);
or OR4 (N10203, N10202, N1925, N671, N5050);
not NOT1 (N10204, N10201);
xor XOR2 (N10205, N10140, N6745);
or OR2 (N10206, N10197, N7191);
nor NOR3 (N10207, N10203, N4166, N6167);
nand NAND2 (N10208, N10206, N188);
or OR3 (N10209, N10207, N6845, N6321);
nor NOR3 (N10210, N10204, N7523, N9243);
nand NAND3 (N10211, N10210, N9060, N9287);
buf BUF1 (N10212, N10189);
nand NAND4 (N10213, N10179, N2011, N5944, N840);
and AND3 (N10214, N10198, N2526, N4245);
nor NOR3 (N10215, N10213, N7199, N9133);
nand NAND3 (N10216, N10212, N6902, N3719);
xor XOR2 (N10217, N10205, N2190);
nor NOR3 (N10218, N10217, N1678, N3373);
or OR3 (N10219, N10180, N336, N4568);
or OR3 (N10220, N10214, N9863, N5244);
nand NAND3 (N10221, N10216, N8232, N7291);
buf BUF1 (N10222, N10221);
and AND4 (N10223, N10220, N3017, N8583, N6998);
buf BUF1 (N10224, N10211);
nand NAND2 (N10225, N10215, N2924);
nand NAND4 (N10226, N10222, N8268, N2319, N1507);
or OR4 (N10227, N10199, N1442, N533, N5866);
buf BUF1 (N10228, N10227);
or OR4 (N10229, N10226, N5489, N7131, N3714);
or OR2 (N10230, N10200, N4729);
or OR3 (N10231, N10224, N1623, N7877);
not NOT1 (N10232, N10231);
nand NAND2 (N10233, N10232, N8851);
not NOT1 (N10234, N10219);
xor XOR2 (N10235, N10230, N518);
xor XOR2 (N10236, N10235, N5390);
nand NAND2 (N10237, N10223, N3706);
xor XOR2 (N10238, N10208, N1714);
and AND4 (N10239, N10209, N5557, N1487, N4943);
xor XOR2 (N10240, N10236, N8743);
or OR2 (N10241, N10229, N6017);
or OR4 (N10242, N10238, N2485, N3337, N1824);
nand NAND4 (N10243, N10237, N150, N2683, N7952);
buf BUF1 (N10244, N10239);
buf BUF1 (N10245, N10242);
nor NOR4 (N10246, N10244, N1776, N1086, N8666);
or OR2 (N10247, N10243, N9151);
xor XOR2 (N10248, N10234, N5884);
buf BUF1 (N10249, N10233);
not NOT1 (N10250, N10225);
xor XOR2 (N10251, N10241, N2423);
or OR4 (N10252, N10251, N5516, N615, N743);
and AND4 (N10253, N10240, N2073, N3977, N2296);
not NOT1 (N10254, N10245);
xor XOR2 (N10255, N10250, N6593);
and AND2 (N10256, N10228, N7606);
and AND4 (N10257, N10249, N4760, N8645, N781);
and AND4 (N10258, N10255, N7627, N10080, N5771);
xor XOR2 (N10259, N10254, N2867);
nor NOR4 (N10260, N10253, N2689, N5838, N7119);
buf BUF1 (N10261, N10260);
and AND2 (N10262, N10252, N268);
or OR4 (N10263, N10256, N561, N304, N9745);
xor XOR2 (N10264, N10259, N5641);
buf BUF1 (N10265, N10248);
or OR3 (N10266, N10264, N5983, N2756);
nand NAND4 (N10267, N10262, N3831, N1790, N907);
xor XOR2 (N10268, N10261, N1488);
not NOT1 (N10269, N10258);
and AND2 (N10270, N10268, N4006);
or OR2 (N10271, N10265, N9280);
and AND2 (N10272, N10247, N3064);
and AND3 (N10273, N10267, N6225, N388);
not NOT1 (N10274, N10272);
buf BUF1 (N10275, N10257);
nand NAND3 (N10276, N10275, N5866, N3675);
nor NOR4 (N10277, N10274, N990, N3102, N337);
or OR3 (N10278, N10263, N3408, N8252);
not NOT1 (N10279, N10278);
xor XOR2 (N10280, N10277, N9896);
xor XOR2 (N10281, N10270, N6793);
buf BUF1 (N10282, N10271);
xor XOR2 (N10283, N10246, N9003);
nor NOR2 (N10284, N10282, N6223);
xor XOR2 (N10285, N10284, N8099);
or OR2 (N10286, N10285, N8288);
and AND2 (N10287, N10280, N5330);
nor NOR2 (N10288, N10286, N2293);
nand NAND3 (N10289, N10276, N9100, N1777);
or OR4 (N10290, N10269, N2354, N3143, N6936);
buf BUF1 (N10291, N10273);
buf BUF1 (N10292, N10290);
not NOT1 (N10293, N10279);
xor XOR2 (N10294, N10218, N8622);
xor XOR2 (N10295, N10292, N4492);
and AND2 (N10296, N10291, N9124);
not NOT1 (N10297, N10296);
xor XOR2 (N10298, N10281, N8602);
nor NOR2 (N10299, N10295, N2124);
buf BUF1 (N10300, N10297);
and AND2 (N10301, N10266, N6919);
and AND2 (N10302, N10298, N6156);
nand NAND2 (N10303, N10300, N9653);
and AND2 (N10304, N10283, N8751);
and AND2 (N10305, N10301, N4462);
or OR4 (N10306, N10304, N3391, N152, N9217);
nand NAND3 (N10307, N10306, N2089, N4183);
buf BUF1 (N10308, N10287);
and AND4 (N10309, N10293, N6513, N4133, N2544);
buf BUF1 (N10310, N10288);
nand NAND2 (N10311, N10302, N4672);
nor NOR3 (N10312, N10311, N10123, N3779);
or OR3 (N10313, N10303, N3491, N8985);
xor XOR2 (N10314, N10299, N9963);
buf BUF1 (N10315, N10309);
nand NAND4 (N10316, N10305, N9338, N9229, N8429);
nor NOR4 (N10317, N10315, N8505, N6620, N6867);
nand NAND3 (N10318, N10317, N5586, N5027);
and AND4 (N10319, N10318, N2641, N1736, N4399);
not NOT1 (N10320, N10316);
or OR3 (N10321, N10319, N7775, N8547);
nand NAND4 (N10322, N10307, N1199, N3876, N5407);
nand NAND4 (N10323, N10308, N3780, N1645, N3089);
and AND4 (N10324, N10313, N5939, N8158, N8275);
or OR4 (N10325, N10320, N1187, N3972, N5462);
nand NAND3 (N10326, N10323, N51, N3539);
nand NAND3 (N10327, N10289, N6460, N6575);
or OR3 (N10328, N10325, N4979, N5513);
and AND2 (N10329, N10310, N851);
buf BUF1 (N10330, N10294);
nor NOR4 (N10331, N10314, N3181, N5301, N975);
not NOT1 (N10332, N10328);
or OR4 (N10333, N10330, N4078, N9861, N9370);
and AND4 (N10334, N10324, N5016, N8727, N9083);
xor XOR2 (N10335, N10331, N8286);
nor NOR3 (N10336, N10327, N1233, N10141);
buf BUF1 (N10337, N10329);
or OR2 (N10338, N10333, N6043);
or OR3 (N10339, N10337, N10189, N3167);
xor XOR2 (N10340, N10312, N7459);
xor XOR2 (N10341, N10339, N8270);
and AND2 (N10342, N10340, N1085);
nor NOR4 (N10343, N10342, N8065, N6479, N7071);
buf BUF1 (N10344, N10335);
buf BUF1 (N10345, N10322);
buf BUF1 (N10346, N10321);
not NOT1 (N10347, N10338);
and AND2 (N10348, N10343, N6150);
or OR2 (N10349, N10346, N1605);
and AND2 (N10350, N10348, N332);
nand NAND2 (N10351, N10332, N2936);
xor XOR2 (N10352, N10345, N9647);
and AND2 (N10353, N10341, N705);
nand NAND3 (N10354, N10349, N1150, N10156);
nor NOR4 (N10355, N10344, N5095, N8961, N4227);
buf BUF1 (N10356, N10353);
buf BUF1 (N10357, N10355);
nand NAND4 (N10358, N10350, N10280, N8319, N8807);
nor NOR2 (N10359, N10336, N2261);
or OR2 (N10360, N10356, N7435);
and AND3 (N10361, N10358, N5798, N8361);
not NOT1 (N10362, N10354);
nor NOR4 (N10363, N10334, N699, N4456, N5205);
nor NOR3 (N10364, N10326, N10053, N811);
not NOT1 (N10365, N10359);
nor NOR2 (N10366, N10351, N1215);
nand NAND4 (N10367, N10361, N9078, N9725, N1375);
or OR4 (N10368, N10365, N1179, N9757, N3187);
or OR4 (N10369, N10357, N4890, N7039, N7370);
nand NAND3 (N10370, N10369, N9541, N3468);
or OR4 (N10371, N10347, N5432, N5004, N6650);
nand NAND4 (N10372, N10368, N1607, N8796, N6957);
buf BUF1 (N10373, N10352);
xor XOR2 (N10374, N10366, N1224);
nor NOR3 (N10375, N10364, N34, N647);
xor XOR2 (N10376, N10371, N8572);
xor XOR2 (N10377, N10367, N2647);
and AND2 (N10378, N10363, N1947);
buf BUF1 (N10379, N10376);
or OR3 (N10380, N10360, N3043, N7675);
buf BUF1 (N10381, N10373);
nand NAND3 (N10382, N10377, N3723, N5431);
or OR2 (N10383, N10370, N3595);
nand NAND4 (N10384, N10380, N5174, N4028, N5089);
not NOT1 (N10385, N10383);
nand NAND3 (N10386, N10362, N2603, N9736);
not NOT1 (N10387, N10378);
buf BUF1 (N10388, N10375);
and AND3 (N10389, N10387, N479, N9028);
xor XOR2 (N10390, N10381, N1300);
nand NAND2 (N10391, N10389, N1148);
not NOT1 (N10392, N10386);
nor NOR3 (N10393, N10388, N6594, N7747);
buf BUF1 (N10394, N10374);
nor NOR4 (N10395, N10385, N5572, N7403, N5679);
and AND3 (N10396, N10395, N1727, N1136);
xor XOR2 (N10397, N10382, N4184);
not NOT1 (N10398, N10384);
or OR2 (N10399, N10394, N8604);
xor XOR2 (N10400, N10393, N3441);
and AND2 (N10401, N10379, N9570);
not NOT1 (N10402, N10397);
nand NAND3 (N10403, N10392, N3782, N8072);
buf BUF1 (N10404, N10399);
not NOT1 (N10405, N10401);
and AND4 (N10406, N10404, N7679, N5736, N8003);
or OR2 (N10407, N10372, N1092);
nor NOR3 (N10408, N10402, N5741, N9386);
xor XOR2 (N10409, N10398, N9544);
xor XOR2 (N10410, N10396, N8493);
xor XOR2 (N10411, N10390, N8158);
nand NAND2 (N10412, N10391, N4253);
and AND3 (N10413, N10406, N6581, N10120);
nor NOR2 (N10414, N10412, N4774);
nor NOR4 (N10415, N10407, N4366, N7611, N9246);
nor NOR4 (N10416, N10405, N7593, N3950, N637);
xor XOR2 (N10417, N10413, N4983);
or OR3 (N10418, N10403, N5991, N4542);
buf BUF1 (N10419, N10417);
xor XOR2 (N10420, N10415, N6463);
and AND2 (N10421, N10416, N1393);
nor NOR2 (N10422, N10419, N5672);
nor NOR3 (N10423, N10400, N6499, N958);
or OR4 (N10424, N10410, N9332, N8273, N2363);
buf BUF1 (N10425, N10411);
nor NOR4 (N10426, N10425, N181, N9900, N5665);
nand NAND3 (N10427, N10420, N8111, N3082);
nand NAND2 (N10428, N10418, N6309);
and AND4 (N10429, N10414, N9563, N9309, N5299);
nor NOR4 (N10430, N10426, N7469, N9543, N5529);
or OR3 (N10431, N10423, N2209, N1851);
or OR4 (N10432, N10430, N5626, N9271, N3906);
not NOT1 (N10433, N10427);
buf BUF1 (N10434, N10432);
not NOT1 (N10435, N10428);
or OR3 (N10436, N10424, N9214, N950);
xor XOR2 (N10437, N10429, N2615);
nand NAND3 (N10438, N10421, N7237, N4981);
nand NAND4 (N10439, N10408, N2752, N7804, N369);
or OR2 (N10440, N10437, N4948);
or OR4 (N10441, N10435, N1774, N5625, N9073);
nor NOR3 (N10442, N10436, N5081, N3431);
or OR4 (N10443, N10438, N423, N1437, N3906);
nor NOR2 (N10444, N10422, N6823);
and AND2 (N10445, N10433, N5465);
not NOT1 (N10446, N10431);
xor XOR2 (N10447, N10441, N9365);
or OR4 (N10448, N10409, N9195, N9357, N6148);
or OR2 (N10449, N10439, N7661);
not NOT1 (N10450, N10434);
xor XOR2 (N10451, N10442, N6024);
nor NOR4 (N10452, N10440, N3208, N2414, N9093);
xor XOR2 (N10453, N10450, N5624);
not NOT1 (N10454, N10446);
or OR4 (N10455, N10448, N4460, N1539, N8528);
nand NAND3 (N10456, N10445, N8702, N8527);
or OR3 (N10457, N10447, N5239, N6717);
nor NOR2 (N10458, N10449, N8532);
nand NAND4 (N10459, N10452, N3339, N4612, N3321);
nand NAND2 (N10460, N10455, N731);
buf BUF1 (N10461, N10454);
and AND2 (N10462, N10458, N6390);
and AND4 (N10463, N10451, N1018, N6711, N5244);
and AND3 (N10464, N10453, N8847, N7495);
buf BUF1 (N10465, N10463);
xor XOR2 (N10466, N10456, N857);
not NOT1 (N10467, N10461);
xor XOR2 (N10468, N10462, N9110);
or OR4 (N10469, N10443, N9223, N8147, N2481);
xor XOR2 (N10470, N10457, N10468);
nand NAND3 (N10471, N7063, N10410, N2148);
nand NAND4 (N10472, N10466, N1795, N6768, N9233);
xor XOR2 (N10473, N10470, N9470);
and AND3 (N10474, N10473, N1797, N2066);
xor XOR2 (N10475, N10460, N8116);
nor NOR2 (N10476, N10465, N9677);
nor NOR2 (N10477, N10472, N7665);
or OR4 (N10478, N10476, N3893, N5130, N4691);
xor XOR2 (N10479, N10444, N5351);
and AND4 (N10480, N10471, N8327, N7933, N4171);
buf BUF1 (N10481, N10474);
not NOT1 (N10482, N10480);
nor NOR2 (N10483, N10475, N6119);
nor NOR2 (N10484, N10469, N6269);
buf BUF1 (N10485, N10459);
not NOT1 (N10486, N10478);
or OR4 (N10487, N10479, N7277, N2006, N502);
buf BUF1 (N10488, N10486);
not NOT1 (N10489, N10467);
or OR2 (N10490, N10483, N7968);
or OR2 (N10491, N10485, N2933);
xor XOR2 (N10492, N10487, N3726);
nand NAND2 (N10493, N10477, N10005);
xor XOR2 (N10494, N10481, N5573);
and AND4 (N10495, N10482, N107, N3971, N5806);
not NOT1 (N10496, N10488);
or OR2 (N10497, N10492, N8156);
nor NOR2 (N10498, N10490, N5624);
nor NOR2 (N10499, N10491, N6984);
not NOT1 (N10500, N10495);
not NOT1 (N10501, N10484);
or OR2 (N10502, N10493, N4874);
xor XOR2 (N10503, N10502, N10051);
xor XOR2 (N10504, N10496, N6682);
buf BUF1 (N10505, N10497);
not NOT1 (N10506, N10501);
buf BUF1 (N10507, N10498);
nor NOR2 (N10508, N10503, N9802);
not NOT1 (N10509, N10489);
and AND4 (N10510, N10508, N9146, N9019, N7096);
nand NAND2 (N10511, N10500, N9178);
or OR4 (N10512, N10507, N1974, N2209, N3234);
and AND3 (N10513, N10512, N9513, N3547);
xor XOR2 (N10514, N10504, N8390);
nand NAND2 (N10515, N10499, N3576);
and AND3 (N10516, N10514, N3930, N2844);
not NOT1 (N10517, N10494);
and AND2 (N10518, N10505, N193);
or OR3 (N10519, N10513, N10262, N9192);
buf BUF1 (N10520, N10510);
xor XOR2 (N10521, N10520, N4722);
not NOT1 (N10522, N10464);
or OR4 (N10523, N10522, N1677, N2570, N4343);
and AND2 (N10524, N10518, N8664);
nand NAND4 (N10525, N10506, N2380, N4435, N8862);
not NOT1 (N10526, N10519);
not NOT1 (N10527, N10515);
nand NAND4 (N10528, N10517, N5217, N3354, N9218);
nor NOR3 (N10529, N10524, N6459, N9538);
nand NAND3 (N10530, N10527, N1925, N8122);
nor NOR4 (N10531, N10526, N4707, N1278, N6768);
buf BUF1 (N10532, N10516);
buf BUF1 (N10533, N10521);
xor XOR2 (N10534, N10528, N10009);
nor NOR3 (N10535, N10531, N10218, N5789);
or OR3 (N10536, N10534, N1485, N7390);
nor NOR3 (N10537, N10536, N2612, N3661);
not NOT1 (N10538, N10511);
xor XOR2 (N10539, N10530, N6871);
buf BUF1 (N10540, N10538);
xor XOR2 (N10541, N10532, N9759);
or OR2 (N10542, N10535, N3586);
not NOT1 (N10543, N10525);
or OR3 (N10544, N10529, N3700, N9633);
nand NAND3 (N10545, N10539, N1556, N10122);
nand NAND3 (N10546, N10543, N5986, N3743);
not NOT1 (N10547, N10542);
or OR3 (N10548, N10523, N613, N2083);
or OR4 (N10549, N10509, N9412, N3735, N4916);
nand NAND4 (N10550, N10540, N8497, N6086, N1376);
xor XOR2 (N10551, N10544, N4425);
not NOT1 (N10552, N10551);
or OR2 (N10553, N10537, N4364);
not NOT1 (N10554, N10553);
xor XOR2 (N10555, N10554, N9930);
not NOT1 (N10556, N10547);
xor XOR2 (N10557, N10546, N2360);
nand NAND4 (N10558, N10555, N7624, N1891, N3923);
nor NOR3 (N10559, N10533, N8378, N9253);
xor XOR2 (N10560, N10550, N7296);
nand NAND4 (N10561, N10549, N6731, N1890, N8405);
xor XOR2 (N10562, N10557, N9521);
buf BUF1 (N10563, N10541);
nor NOR2 (N10564, N10548, N2684);
or OR4 (N10565, N10564, N4858, N6042, N8810);
nand NAND4 (N10566, N10561, N1260, N9962, N4348);
and AND3 (N10567, N10545, N9795, N3142);
and AND4 (N10568, N10560, N7987, N142, N2323);
or OR3 (N10569, N10558, N2397, N7497);
nor NOR3 (N10570, N10563, N5357, N2768);
not NOT1 (N10571, N10562);
or OR3 (N10572, N10569, N8584, N8728);
nor NOR3 (N10573, N10570, N5834, N810);
buf BUF1 (N10574, N10566);
xor XOR2 (N10575, N10572, N7375);
buf BUF1 (N10576, N10565);
or OR4 (N10577, N10567, N9310, N7419, N5445);
buf BUF1 (N10578, N10571);
nor NOR3 (N10579, N10577, N8694, N5072);
xor XOR2 (N10580, N10575, N4288);
xor XOR2 (N10581, N10574, N2135);
xor XOR2 (N10582, N10552, N1724);
buf BUF1 (N10583, N10582);
and AND3 (N10584, N10583, N3932, N2192);
not NOT1 (N10585, N10584);
nand NAND3 (N10586, N10556, N8469, N1724);
xor XOR2 (N10587, N10585, N1353);
xor XOR2 (N10588, N10576, N7929);
or OR2 (N10589, N10586, N4363);
buf BUF1 (N10590, N10578);
or OR2 (N10591, N10587, N419);
or OR3 (N10592, N10589, N1999, N3433);
nand NAND3 (N10593, N10588, N5918, N6451);
buf BUF1 (N10594, N10593);
nand NAND2 (N10595, N10559, N1234);
nor NOR4 (N10596, N10592, N4736, N1184, N9349);
xor XOR2 (N10597, N10596, N9500);
xor XOR2 (N10598, N10591, N3979);
or OR2 (N10599, N10581, N5315);
nor NOR3 (N10600, N10595, N9057, N6826);
and AND4 (N10601, N10573, N6590, N4892, N3744);
and AND4 (N10602, N10568, N6680, N10454, N5053);
and AND4 (N10603, N10601, N10292, N2048, N6658);
nand NAND4 (N10604, N10580, N9123, N2185, N340);
buf BUF1 (N10605, N10602);
and AND4 (N10606, N10599, N1448, N4506, N5861);
not NOT1 (N10607, N10579);
xor XOR2 (N10608, N10603, N3828);
nand NAND4 (N10609, N10600, N9376, N6817, N6153);
and AND2 (N10610, N10597, N2516);
xor XOR2 (N10611, N10604, N2055);
not NOT1 (N10612, N10607);
nor NOR4 (N10613, N10594, N112, N8486, N1424);
buf BUF1 (N10614, N10606);
nand NAND4 (N10615, N10611, N2733, N4806, N3655);
xor XOR2 (N10616, N10605, N8900);
buf BUF1 (N10617, N10612);
nor NOR4 (N10618, N10609, N2455, N10300, N5523);
and AND2 (N10619, N10618, N2889);
nand NAND2 (N10620, N10608, N5189);
not NOT1 (N10621, N10613);
nand NAND2 (N10622, N10615, N5325);
nor NOR2 (N10623, N10598, N10172);
not NOT1 (N10624, N10622);
or OR3 (N10625, N10616, N344, N2533);
nor NOR3 (N10626, N10623, N4713, N2726);
not NOT1 (N10627, N10626);
not NOT1 (N10628, N10619);
nand NAND4 (N10629, N10610, N7170, N6982, N3268);
or OR2 (N10630, N10614, N9004);
not NOT1 (N10631, N10620);
nor NOR4 (N10632, N10625, N9495, N1638, N6821);
and AND2 (N10633, N10629, N9326);
and AND3 (N10634, N10624, N2227, N7498);
nand NAND3 (N10635, N10621, N5744, N8744);
nand NAND4 (N10636, N10635, N5965, N5638, N444);
not NOT1 (N10637, N10631);
xor XOR2 (N10638, N10637, N5528);
not NOT1 (N10639, N10633);
or OR2 (N10640, N10636, N9289);
or OR3 (N10641, N10634, N9743, N5372);
or OR4 (N10642, N10628, N9210, N8904, N3157);
nand NAND3 (N10643, N10630, N8736, N6756);
xor XOR2 (N10644, N10639, N1561);
nor NOR2 (N10645, N10617, N8652);
nand NAND2 (N10646, N10644, N565);
nand NAND2 (N10647, N10645, N9911);
nor NOR4 (N10648, N10642, N10303, N6563, N1068);
xor XOR2 (N10649, N10638, N6375);
xor XOR2 (N10650, N10641, N946);
nor NOR3 (N10651, N10647, N9078, N8142);
and AND3 (N10652, N10651, N6108, N6650);
not NOT1 (N10653, N10632);
xor XOR2 (N10654, N10643, N4703);
nor NOR3 (N10655, N10649, N9807, N1513);
nor NOR2 (N10656, N10627, N9745);
xor XOR2 (N10657, N10652, N4135);
xor XOR2 (N10658, N10648, N4187);
not NOT1 (N10659, N10655);
not NOT1 (N10660, N10590);
and AND4 (N10661, N10650, N2753, N6111, N9875);
and AND4 (N10662, N10661, N2006, N3463, N8600);
not NOT1 (N10663, N10662);
and AND3 (N10664, N10660, N5236, N2958);
xor XOR2 (N10665, N10659, N756);
and AND4 (N10666, N10664, N334, N1291, N5079);
or OR3 (N10667, N10657, N7081, N3255);
xor XOR2 (N10668, N10656, N1928);
nand NAND3 (N10669, N10646, N6220, N709);
not NOT1 (N10670, N10669);
nor NOR4 (N10671, N10663, N3544, N5487, N2743);
not NOT1 (N10672, N10671);
nor NOR3 (N10673, N10658, N1242, N9216);
not NOT1 (N10674, N10668);
nand NAND2 (N10675, N10673, N2083);
xor XOR2 (N10676, N10665, N8865);
not NOT1 (N10677, N10666);
not NOT1 (N10678, N10667);
or OR2 (N10679, N10653, N2752);
nor NOR3 (N10680, N10670, N10278, N2569);
and AND2 (N10681, N10674, N902);
not NOT1 (N10682, N10681);
buf BUF1 (N10683, N10672);
not NOT1 (N10684, N10640);
not NOT1 (N10685, N10654);
nor NOR4 (N10686, N10677, N8068, N10538, N6943);
xor XOR2 (N10687, N10679, N1409);
or OR4 (N10688, N10675, N8412, N8085, N10225);
buf BUF1 (N10689, N10686);
nor NOR2 (N10690, N10688, N3899);
and AND3 (N10691, N10685, N7747, N6748);
buf BUF1 (N10692, N10687);
not NOT1 (N10693, N10690);
buf BUF1 (N10694, N10692);
not NOT1 (N10695, N10684);
nand NAND3 (N10696, N10691, N10361, N387);
xor XOR2 (N10697, N10695, N3238);
xor XOR2 (N10698, N10694, N7657);
nand NAND4 (N10699, N10678, N3708, N7695, N2162);
or OR2 (N10700, N10680, N8640);
xor XOR2 (N10701, N10689, N7904);
or OR3 (N10702, N10700, N7363, N2343);
not NOT1 (N10703, N10701);
and AND3 (N10704, N10682, N2404, N5063);
not NOT1 (N10705, N10676);
buf BUF1 (N10706, N10704);
nand NAND4 (N10707, N10696, N5274, N2993, N3940);
xor XOR2 (N10708, N10707, N5043);
not NOT1 (N10709, N10683);
xor XOR2 (N10710, N10699, N5554);
or OR3 (N10711, N10693, N2900, N7549);
nor NOR4 (N10712, N10711, N4228, N2690, N10393);
nor NOR2 (N10713, N10705, N2151);
nor NOR3 (N10714, N10709, N1862, N8463);
or OR4 (N10715, N10706, N988, N1739, N8869);
nand NAND2 (N10716, N10710, N4451);
not NOT1 (N10717, N10714);
nand NAND3 (N10718, N10702, N828, N9528);
and AND4 (N10719, N10716, N10655, N398, N8420);
and AND2 (N10720, N10698, N8597);
and AND4 (N10721, N10713, N6658, N2736, N7727);
not NOT1 (N10722, N10720);
nor NOR2 (N10723, N10712, N7395);
buf BUF1 (N10724, N10722);
xor XOR2 (N10725, N10724, N349);
or OR2 (N10726, N10715, N3196);
or OR3 (N10727, N10723, N10602, N4334);
nand NAND4 (N10728, N10718, N8098, N7245, N7186);
or OR4 (N10729, N10719, N9337, N4346, N3240);
or OR2 (N10730, N10717, N10144);
xor XOR2 (N10731, N10727, N4912);
and AND3 (N10732, N10730, N1486, N9684);
not NOT1 (N10733, N10732);
and AND3 (N10734, N10725, N4847, N4506);
and AND3 (N10735, N10726, N4122, N8168);
and AND2 (N10736, N10735, N7103);
buf BUF1 (N10737, N10733);
xor XOR2 (N10738, N10736, N9782);
nor NOR4 (N10739, N10729, N834, N7225, N93);
and AND2 (N10740, N10737, N6610);
not NOT1 (N10741, N10731);
nor NOR4 (N10742, N10734, N5642, N9752, N515);
or OR3 (N10743, N10742, N7531, N9909);
nand NAND4 (N10744, N10697, N2770, N478, N3874);
nor NOR4 (N10745, N10738, N1025, N5668, N553);
nand NAND4 (N10746, N10741, N9217, N463, N1351);
and AND4 (N10747, N10746, N1000, N4973, N203);
and AND3 (N10748, N10745, N10499, N7844);
nor NOR4 (N10749, N10739, N5384, N1645, N1618);
not NOT1 (N10750, N10728);
not NOT1 (N10751, N10747);
buf BUF1 (N10752, N10721);
and AND2 (N10753, N10749, N3492);
xor XOR2 (N10754, N10703, N6429);
nor NOR3 (N10755, N10743, N1264, N1060);
buf BUF1 (N10756, N10751);
not NOT1 (N10757, N10752);
nor NOR2 (N10758, N10708, N2123);
or OR4 (N10759, N10755, N2024, N1562, N7257);
and AND4 (N10760, N10740, N5813, N9087, N6300);
nor NOR4 (N10761, N10753, N3263, N2612, N754);
not NOT1 (N10762, N10761);
nand NAND4 (N10763, N10750, N608, N2064, N8749);
buf BUF1 (N10764, N10744);
not NOT1 (N10765, N10758);
and AND3 (N10766, N10760, N6066, N10718);
buf BUF1 (N10767, N10763);
or OR2 (N10768, N10764, N3637);
xor XOR2 (N10769, N10759, N2702);
buf BUF1 (N10770, N10769);
nor NOR4 (N10771, N10770, N4582, N3604, N5983);
buf BUF1 (N10772, N10762);
not NOT1 (N10773, N10771);
not NOT1 (N10774, N10756);
and AND2 (N10775, N10757, N2885);
and AND2 (N10776, N10748, N649);
not NOT1 (N10777, N10774);
nand NAND3 (N10778, N10767, N580, N5925);
xor XOR2 (N10779, N10778, N2600);
xor XOR2 (N10780, N10765, N5072);
and AND4 (N10781, N10776, N1982, N3654, N8603);
buf BUF1 (N10782, N10754);
nor NOR2 (N10783, N10768, N10449);
buf BUF1 (N10784, N10775);
xor XOR2 (N10785, N10784, N2190);
nor NOR2 (N10786, N10783, N7928);
nand NAND2 (N10787, N10786, N8771);
not NOT1 (N10788, N10787);
and AND2 (N10789, N10780, N2846);
nor NOR3 (N10790, N10766, N9586, N7094);
or OR4 (N10791, N10789, N3191, N7328, N1347);
nand NAND3 (N10792, N10785, N3392, N5908);
nor NOR2 (N10793, N10788, N8259);
or OR2 (N10794, N10790, N6240);
nand NAND4 (N10795, N10777, N10684, N7479, N5944);
nand NAND2 (N10796, N10772, N8806);
xor XOR2 (N10797, N10782, N5372);
not NOT1 (N10798, N10797);
nand NAND4 (N10799, N10791, N5426, N4239, N4779);
buf BUF1 (N10800, N10794);
and AND4 (N10801, N10779, N3815, N1545, N4891);
nand NAND4 (N10802, N10796, N6699, N3143, N1044);
buf BUF1 (N10803, N10799);
or OR3 (N10804, N10801, N2963, N2451);
nand NAND4 (N10805, N10792, N10150, N246, N10776);
nand NAND3 (N10806, N10805, N5272, N6138);
xor XOR2 (N10807, N10800, N2249);
xor XOR2 (N10808, N10804, N4024);
buf BUF1 (N10809, N10793);
and AND4 (N10810, N10803, N8322, N300, N5417);
buf BUF1 (N10811, N10781);
nor NOR4 (N10812, N10802, N9210, N358, N5082);
and AND3 (N10813, N10812, N1587, N7470);
or OR3 (N10814, N10795, N8349, N4004);
nand NAND2 (N10815, N10808, N10719);
or OR2 (N10816, N10806, N3106);
or OR4 (N10817, N10813, N7955, N7335, N3778);
not NOT1 (N10818, N10798);
nor NOR3 (N10819, N10818, N3925, N2636);
or OR2 (N10820, N10819, N2452);
or OR4 (N10821, N10815, N1936, N9200, N1848);
nor NOR2 (N10822, N10816, N835);
nor NOR4 (N10823, N10811, N5236, N7835, N75);
xor XOR2 (N10824, N10810, N8774);
or OR2 (N10825, N10814, N4693);
nand NAND2 (N10826, N10773, N5046);
buf BUF1 (N10827, N10822);
or OR2 (N10828, N10809, N2540);
not NOT1 (N10829, N10827);
and AND2 (N10830, N10828, N6049);
buf BUF1 (N10831, N10824);
nand NAND3 (N10832, N10826, N551, N3719);
and AND4 (N10833, N10832, N2733, N2704, N8964);
not NOT1 (N10834, N10829);
buf BUF1 (N10835, N10830);
or OR4 (N10836, N10823, N3473, N5772, N2935);
buf BUF1 (N10837, N10835);
or OR4 (N10838, N10825, N9410, N6483, N7192);
nand NAND3 (N10839, N10834, N2419, N9409);
xor XOR2 (N10840, N10836, N7462);
and AND4 (N10841, N10821, N1412, N10264, N1846);
and AND4 (N10842, N10838, N2037, N5606, N5811);
or OR2 (N10843, N10833, N4413);
not NOT1 (N10844, N10841);
nor NOR3 (N10845, N10817, N3306, N4770);
nand NAND3 (N10846, N10842, N3474, N721);
buf BUF1 (N10847, N10845);
buf BUF1 (N10848, N10831);
or OR3 (N10849, N10820, N7738, N4839);
nor NOR3 (N10850, N10846, N1243, N3949);
not NOT1 (N10851, N10843);
and AND2 (N10852, N10837, N2630);
buf BUF1 (N10853, N10849);
nand NAND3 (N10854, N10853, N7440, N1011);
nor NOR3 (N10855, N10851, N8065, N8284);
nand NAND4 (N10856, N10852, N1153, N718, N1612);
nand NAND4 (N10857, N10856, N6945, N2040, N2700);
not NOT1 (N10858, N10850);
buf BUF1 (N10859, N10839);
nor NOR4 (N10860, N10807, N5196, N3853, N207);
xor XOR2 (N10861, N10857, N4170);
xor XOR2 (N10862, N10858, N4996);
xor XOR2 (N10863, N10844, N3866);
buf BUF1 (N10864, N10862);
or OR4 (N10865, N10854, N453, N8132, N998);
not NOT1 (N10866, N10864);
and AND2 (N10867, N10855, N9796);
buf BUF1 (N10868, N10865);
not NOT1 (N10869, N10840);
or OR3 (N10870, N10859, N3963, N7322);
buf BUF1 (N10871, N10847);
not NOT1 (N10872, N10861);
and AND2 (N10873, N10860, N1498);
not NOT1 (N10874, N10863);
nand NAND3 (N10875, N10866, N9782, N7774);
and AND3 (N10876, N10875, N1306, N6639);
or OR3 (N10877, N10868, N362, N1626);
nor NOR3 (N10878, N10877, N8926, N10727);
buf BUF1 (N10879, N10867);
and AND3 (N10880, N10871, N3709, N8448);
nor NOR2 (N10881, N10878, N2163);
nor NOR2 (N10882, N10869, N5969);
or OR3 (N10883, N10879, N4684, N1066);
not NOT1 (N10884, N10872);
nor NOR3 (N10885, N10873, N3495, N3178);
not NOT1 (N10886, N10883);
or OR3 (N10887, N10885, N4151, N929);
or OR4 (N10888, N10874, N2744, N6023, N4587);
not NOT1 (N10889, N10848);
nor NOR2 (N10890, N10888, N10400);
nand NAND3 (N10891, N10887, N3229, N7717);
and AND4 (N10892, N10870, N3649, N9699, N4748);
nor NOR2 (N10893, N10881, N2694);
buf BUF1 (N10894, N10880);
nor NOR3 (N10895, N10891, N7772, N4936);
or OR3 (N10896, N10882, N1783, N6907);
or OR4 (N10897, N10893, N9979, N2534, N1570);
or OR4 (N10898, N10884, N8658, N9628, N6630);
not NOT1 (N10899, N10889);
buf BUF1 (N10900, N10897);
not NOT1 (N10901, N10900);
buf BUF1 (N10902, N10894);
and AND2 (N10903, N10876, N10320);
xor XOR2 (N10904, N10898, N9636);
or OR2 (N10905, N10899, N5196);
xor XOR2 (N10906, N10890, N2658);
nor NOR3 (N10907, N10905, N7948, N5871);
or OR4 (N10908, N10903, N1287, N8210, N5373);
xor XOR2 (N10909, N10901, N8320);
or OR2 (N10910, N10895, N3884);
nand NAND4 (N10911, N10910, N3968, N4766, N3720);
and AND4 (N10912, N10911, N6152, N1802, N2330);
or OR2 (N10913, N10908, N3458);
or OR2 (N10914, N10904, N8863);
and AND2 (N10915, N10892, N7815);
and AND3 (N10916, N10902, N3492, N6433);
buf BUF1 (N10917, N10907);
nand NAND2 (N10918, N10896, N1545);
not NOT1 (N10919, N10912);
and AND2 (N10920, N10917, N240);
not NOT1 (N10921, N10919);
nor NOR2 (N10922, N10913, N633);
buf BUF1 (N10923, N10906);
or OR2 (N10924, N10909, N10435);
xor XOR2 (N10925, N10923, N1242);
nor NOR2 (N10926, N10925, N4248);
nand NAND4 (N10927, N10926, N3576, N4394, N3311);
nor NOR3 (N10928, N10916, N813, N6024);
buf BUF1 (N10929, N10920);
xor XOR2 (N10930, N10921, N7611);
buf BUF1 (N10931, N10929);
buf BUF1 (N10932, N10927);
xor XOR2 (N10933, N10918, N8588);
buf BUF1 (N10934, N10922);
or OR3 (N10935, N10930, N10729, N1760);
not NOT1 (N10936, N10932);
xor XOR2 (N10937, N10915, N8280);
or OR4 (N10938, N10928, N901, N1687, N6505);
and AND2 (N10939, N10935, N1726);
not NOT1 (N10940, N10936);
nor NOR2 (N10941, N10933, N1108);
not NOT1 (N10942, N10940);
nand NAND4 (N10943, N10937, N2871, N9390, N6952);
nor NOR2 (N10944, N10943, N4624);
buf BUF1 (N10945, N10938);
not NOT1 (N10946, N10934);
and AND2 (N10947, N10914, N6703);
buf BUF1 (N10948, N10945);
not NOT1 (N10949, N10924);
and AND2 (N10950, N10946, N4375);
nand NAND4 (N10951, N10931, N9880, N464, N2953);
or OR4 (N10952, N10944, N5651, N1529, N2608);
nand NAND4 (N10953, N10952, N8974, N9507, N200);
nand NAND3 (N10954, N10947, N1273, N10801);
nand NAND3 (N10955, N10950, N2559, N750);
not NOT1 (N10956, N10951);
buf BUF1 (N10957, N10939);
or OR3 (N10958, N10886, N9591, N6368);
buf BUF1 (N10959, N10941);
buf BUF1 (N10960, N10942);
not NOT1 (N10961, N10957);
nand NAND2 (N10962, N10956, N706);
nand NAND4 (N10963, N10955, N5723, N7340, N4537);
xor XOR2 (N10964, N10954, N5031);
nand NAND3 (N10965, N10959, N10833, N775);
nor NOR2 (N10966, N10964, N1202);
nor NOR3 (N10967, N10966, N8303, N3517);
xor XOR2 (N10968, N10965, N9338);
nor NOR4 (N10969, N10962, N10627, N10610, N9268);
buf BUF1 (N10970, N10969);
nor NOR2 (N10971, N10970, N5323);
not NOT1 (N10972, N10967);
buf BUF1 (N10973, N10948);
xor XOR2 (N10974, N10971, N5018);
nor NOR3 (N10975, N10963, N436, N8345);
nor NOR3 (N10976, N10958, N6745, N4364);
buf BUF1 (N10977, N10949);
and AND2 (N10978, N10953, N857);
nor NOR2 (N10979, N10961, N9969);
and AND4 (N10980, N10968, N1328, N10836, N5089);
nand NAND2 (N10981, N10977, N6240);
or OR3 (N10982, N10980, N8709, N960);
xor XOR2 (N10983, N10960, N6980);
xor XOR2 (N10984, N10978, N10576);
and AND2 (N10985, N10982, N5074);
buf BUF1 (N10986, N10975);
and AND2 (N10987, N10983, N1100);
nand NAND2 (N10988, N10974, N9330);
buf BUF1 (N10989, N10979);
buf BUF1 (N10990, N10973);
xor XOR2 (N10991, N10989, N2560);
and AND3 (N10992, N10981, N10385, N8121);
nand NAND2 (N10993, N10985, N2991);
xor XOR2 (N10994, N10988, N389);
buf BUF1 (N10995, N10976);
xor XOR2 (N10996, N10990, N4166);
nor NOR3 (N10997, N10991, N9945, N2010);
nand NAND2 (N10998, N10986, N9654);
buf BUF1 (N10999, N10992);
not NOT1 (N11000, N10997);
buf BUF1 (N11001, N10996);
and AND3 (N11002, N10987, N1894, N2946);
buf BUF1 (N11003, N11000);
and AND2 (N11004, N10984, N1365);
nor NOR3 (N11005, N10998, N600, N2871);
xor XOR2 (N11006, N11003, N7839);
buf BUF1 (N11007, N11005);
not NOT1 (N11008, N11001);
xor XOR2 (N11009, N11004, N10410);
xor XOR2 (N11010, N11007, N3579);
nand NAND2 (N11011, N10994, N3493);
not NOT1 (N11012, N10972);
xor XOR2 (N11013, N11009, N2167);
nand NAND4 (N11014, N11002, N10149, N4196, N5338);
not NOT1 (N11015, N10993);
buf BUF1 (N11016, N11011);
or OR2 (N11017, N10999, N785);
nand NAND4 (N11018, N11006, N8080, N4290, N2859);
or OR2 (N11019, N11017, N10491);
not NOT1 (N11020, N11018);
not NOT1 (N11021, N11013);
not NOT1 (N11022, N10995);
xor XOR2 (N11023, N11012, N6652);
nand NAND4 (N11024, N11019, N3535, N3777, N4785);
and AND2 (N11025, N11016, N2790);
nor NOR2 (N11026, N11023, N7818);
buf BUF1 (N11027, N11022);
xor XOR2 (N11028, N11010, N2381);
nor NOR3 (N11029, N11020, N9911, N10640);
not NOT1 (N11030, N11015);
nor NOR4 (N11031, N11021, N5040, N10635, N9053);
nor NOR4 (N11032, N11030, N4901, N9484, N4969);
buf BUF1 (N11033, N11025);
and AND2 (N11034, N11028, N4571);
or OR2 (N11035, N11029, N514);
nor NOR2 (N11036, N11034, N3567);
buf BUF1 (N11037, N11027);
and AND3 (N11038, N11024, N4643, N5417);
not NOT1 (N11039, N11033);
nor NOR3 (N11040, N11014, N2654, N10448);
or OR2 (N11041, N11008, N10634);
or OR2 (N11042, N11035, N2656);
not NOT1 (N11043, N11042);
not NOT1 (N11044, N11031);
xor XOR2 (N11045, N11044, N2590);
nor NOR3 (N11046, N11040, N9549, N9942);
not NOT1 (N11047, N11026);
nor NOR2 (N11048, N11043, N5102);
nor NOR3 (N11049, N11038, N1978, N3692);
or OR3 (N11050, N11039, N5932, N6406);
not NOT1 (N11051, N11048);
and AND2 (N11052, N11046, N3687);
nor NOR3 (N11053, N11032, N9442, N4596);
buf BUF1 (N11054, N11036);
or OR2 (N11055, N11041, N9299);
not NOT1 (N11056, N11045);
or OR3 (N11057, N11049, N10648, N8301);
or OR4 (N11058, N11057, N5960, N3754, N10510);
or OR4 (N11059, N11052, N1148, N565, N5244);
or OR4 (N11060, N11055, N2646, N5795, N4564);
and AND2 (N11061, N11060, N9981);
or OR4 (N11062, N11054, N7834, N7932, N1816);
xor XOR2 (N11063, N11058, N1356);
and AND4 (N11064, N11051, N1084, N1050, N8732);
buf BUF1 (N11065, N11062);
nor NOR3 (N11066, N11053, N4788, N5324);
and AND2 (N11067, N11037, N6417);
nor NOR4 (N11068, N11063, N7327, N7209, N5106);
nand NAND2 (N11069, N11068, N5714);
xor XOR2 (N11070, N11064, N9959);
buf BUF1 (N11071, N11047);
or OR2 (N11072, N11061, N2025);
nand NAND2 (N11073, N11072, N7725);
nor NOR2 (N11074, N11073, N4365);
and AND2 (N11075, N11065, N3172);
nand NAND3 (N11076, N11066, N6044, N9521);
buf BUF1 (N11077, N11074);
or OR4 (N11078, N11070, N394, N8274, N7939);
xor XOR2 (N11079, N11056, N8705);
not NOT1 (N11080, N11071);
not NOT1 (N11081, N11075);
nand NAND2 (N11082, N11067, N9854);
not NOT1 (N11083, N11082);
and AND4 (N11084, N11076, N2978, N5125, N1169);
and AND4 (N11085, N11081, N7, N7873, N7599);
buf BUF1 (N11086, N11079);
or OR2 (N11087, N11084, N10150);
not NOT1 (N11088, N11069);
nand NAND2 (N11089, N11086, N6063);
xor XOR2 (N11090, N11088, N6091);
and AND2 (N11091, N11089, N2068);
and AND2 (N11092, N11077, N3467);
and AND4 (N11093, N11080, N10633, N442, N5267);
not NOT1 (N11094, N11091);
or OR3 (N11095, N11087, N4589, N5531);
buf BUF1 (N11096, N11092);
not NOT1 (N11097, N11090);
nand NAND4 (N11098, N11096, N5640, N2416, N5680);
nor NOR3 (N11099, N11093, N5481, N7185);
not NOT1 (N11100, N11085);
xor XOR2 (N11101, N11097, N6857);
and AND3 (N11102, N11101, N3361, N4126);
nand NAND3 (N11103, N11050, N9039, N3243);
xor XOR2 (N11104, N11099, N3750);
nand NAND4 (N11105, N11102, N534, N5591, N1729);
nor NOR4 (N11106, N11083, N5992, N6200, N7465);
xor XOR2 (N11107, N11106, N7476);
or OR2 (N11108, N11100, N5684);
nand NAND3 (N11109, N11095, N2147, N5993);
xor XOR2 (N11110, N11059, N10005);
xor XOR2 (N11111, N11107, N2623);
and AND2 (N11112, N11109, N8159);
nor NOR3 (N11113, N11112, N5985, N2576);
xor XOR2 (N11114, N11078, N4234);
nand NAND2 (N11115, N11113, N9901);
or OR3 (N11116, N11104, N5430, N2744);
nand NAND4 (N11117, N11108, N736, N4364, N5073);
not NOT1 (N11118, N11114);
not NOT1 (N11119, N11111);
buf BUF1 (N11120, N11098);
not NOT1 (N11121, N11120);
nand NAND4 (N11122, N11118, N1339, N6383, N756);
nor NOR3 (N11123, N11094, N4949, N9214);
xor XOR2 (N11124, N11105, N501);
and AND3 (N11125, N11117, N5311, N3258);
nand NAND4 (N11126, N11110, N2278, N9030, N7941);
xor XOR2 (N11127, N11126, N6928);
not NOT1 (N11128, N11119);
and AND2 (N11129, N11115, N10762);
or OR3 (N11130, N11128, N536, N4886);
and AND2 (N11131, N11125, N5859);
xor XOR2 (N11132, N11124, N7795);
and AND3 (N11133, N11122, N6585, N6809);
not NOT1 (N11134, N11133);
or OR4 (N11135, N11134, N697, N8609, N7408);
or OR3 (N11136, N11103, N5453, N5721);
and AND2 (N11137, N11132, N4950);
nor NOR2 (N11138, N11129, N9448);
xor XOR2 (N11139, N11136, N6009);
not NOT1 (N11140, N11131);
and AND2 (N11141, N11130, N2619);
and AND2 (N11142, N11137, N9000);
or OR2 (N11143, N11142, N6356);
xor XOR2 (N11144, N11141, N3292);
and AND3 (N11145, N11138, N2557, N10754);
buf BUF1 (N11146, N11127);
or OR4 (N11147, N11144, N5996, N609, N7993);
or OR2 (N11148, N11146, N4960);
not NOT1 (N11149, N11139);
or OR2 (N11150, N11121, N6851);
xor XOR2 (N11151, N11148, N8401);
buf BUF1 (N11152, N11116);
or OR3 (N11153, N11135, N1616, N6408);
and AND2 (N11154, N11151, N6247);
nand NAND3 (N11155, N11152, N9708, N1068);
and AND4 (N11156, N11153, N163, N3978, N5659);
nor NOR4 (N11157, N11145, N6829, N7233, N9002);
and AND3 (N11158, N11123, N9358, N3931);
nand NAND4 (N11159, N11158, N555, N794, N5170);
or OR3 (N11160, N11140, N4930, N6128);
nand NAND2 (N11161, N11149, N2524);
or OR3 (N11162, N11150, N2514, N767);
or OR4 (N11163, N11156, N5814, N418, N10124);
buf BUF1 (N11164, N11162);
nor NOR4 (N11165, N11163, N8506, N7174, N5614);
nand NAND4 (N11166, N11160, N538, N6198, N4388);
buf BUF1 (N11167, N11165);
xor XOR2 (N11168, N11167, N4068);
not NOT1 (N11169, N11159);
nor NOR3 (N11170, N11168, N5555, N8735);
buf BUF1 (N11171, N11147);
or OR2 (N11172, N11166, N4252);
buf BUF1 (N11173, N11169);
or OR4 (N11174, N11173, N883, N2227, N2043);
xor XOR2 (N11175, N11154, N948);
nand NAND2 (N11176, N11174, N5672);
nand NAND3 (N11177, N11164, N4158, N10426);
xor XOR2 (N11178, N11175, N5213);
nand NAND4 (N11179, N11143, N1655, N6155, N5363);
not NOT1 (N11180, N11172);
or OR2 (N11181, N11180, N7432);
nand NAND3 (N11182, N11157, N10039, N10123);
xor XOR2 (N11183, N11161, N4427);
nand NAND3 (N11184, N11170, N970, N3126);
buf BUF1 (N11185, N11155);
or OR3 (N11186, N11179, N1362, N1206);
buf BUF1 (N11187, N11182);
not NOT1 (N11188, N11176);
or OR3 (N11189, N11178, N8420, N7662);
and AND2 (N11190, N11185, N5115);
buf BUF1 (N11191, N11183);
nand NAND3 (N11192, N11188, N5866, N7025);
nor NOR2 (N11193, N11191, N10880);
xor XOR2 (N11194, N11193, N10875);
buf BUF1 (N11195, N11177);
and AND3 (N11196, N11189, N8330, N10862);
or OR4 (N11197, N11196, N3997, N1732, N9705);
nor NOR4 (N11198, N11197, N5882, N8456, N1483);
xor XOR2 (N11199, N11198, N2004);
not NOT1 (N11200, N11171);
nor NOR4 (N11201, N11199, N7648, N10628, N10526);
buf BUF1 (N11202, N11184);
buf BUF1 (N11203, N11194);
or OR3 (N11204, N11201, N9947, N7486);
xor XOR2 (N11205, N11192, N8416);
not NOT1 (N11206, N11181);
nor NOR3 (N11207, N11203, N7587, N7513);
or OR3 (N11208, N11187, N7849, N3551);
xor XOR2 (N11209, N11204, N635);
buf BUF1 (N11210, N11200);
not NOT1 (N11211, N11209);
buf BUF1 (N11212, N11206);
buf BUF1 (N11213, N11202);
and AND3 (N11214, N11212, N3136, N5229);
nand NAND4 (N11215, N11195, N3701, N7502, N8463);
buf BUF1 (N11216, N11190);
or OR2 (N11217, N11213, N1098);
nand NAND3 (N11218, N11217, N3337, N6350);
not NOT1 (N11219, N11216);
or OR3 (N11220, N11219, N2678, N38);
not NOT1 (N11221, N11210);
xor XOR2 (N11222, N11211, N6038);
nor NOR3 (N11223, N11214, N4705, N363);
and AND4 (N11224, N11205, N2655, N7473, N5647);
not NOT1 (N11225, N11222);
nor NOR2 (N11226, N11208, N1958);
xor XOR2 (N11227, N11218, N10540);
and AND2 (N11228, N11186, N4970);
xor XOR2 (N11229, N11228, N10510);
buf BUF1 (N11230, N11215);
buf BUF1 (N11231, N11207);
nand NAND2 (N11232, N11223, N383);
and AND4 (N11233, N11229, N3123, N1117, N8992);
buf BUF1 (N11234, N11227);
xor XOR2 (N11235, N11230, N5791);
nor NOR2 (N11236, N11226, N1515);
not NOT1 (N11237, N11234);
buf BUF1 (N11238, N11221);
or OR2 (N11239, N11236, N1746);
or OR3 (N11240, N11225, N595, N4334);
xor XOR2 (N11241, N11232, N4308);
buf BUF1 (N11242, N11220);
nand NAND2 (N11243, N11233, N500);
and AND2 (N11244, N11241, N6142);
and AND2 (N11245, N11235, N3277);
nor NOR2 (N11246, N11237, N8053);
nor NOR3 (N11247, N11246, N3365, N1763);
nor NOR2 (N11248, N11239, N6056);
nand NAND4 (N11249, N11244, N1588, N85, N8623);
or OR2 (N11250, N11248, N7471);
or OR2 (N11251, N11247, N8386);
nand NAND3 (N11252, N11251, N7498, N6494);
nand NAND3 (N11253, N11224, N7535, N6132);
nand NAND4 (N11254, N11238, N3100, N5455, N10475);
not NOT1 (N11255, N11254);
not NOT1 (N11256, N11243);
nor NOR4 (N11257, N11242, N10033, N8709, N3781);
and AND4 (N11258, N11240, N9058, N5938, N11167);
buf BUF1 (N11259, N11256);
buf BUF1 (N11260, N11253);
nor NOR2 (N11261, N11257, N8382);
nand NAND4 (N11262, N11259, N9448, N3515, N9913);
nor NOR4 (N11263, N11250, N4697, N6245, N5177);
not NOT1 (N11264, N11261);
not NOT1 (N11265, N11258);
xor XOR2 (N11266, N11245, N3418);
buf BUF1 (N11267, N11249);
nand NAND3 (N11268, N11260, N5093, N1534);
buf BUF1 (N11269, N11262);
or OR2 (N11270, N11263, N4387);
buf BUF1 (N11271, N11252);
and AND3 (N11272, N11255, N185, N10127);
buf BUF1 (N11273, N11268);
nor NOR2 (N11274, N11264, N8078);
nand NAND4 (N11275, N11271, N11253, N6123, N933);
buf BUF1 (N11276, N11266);
nand NAND3 (N11277, N11231, N5036, N2705);
xor XOR2 (N11278, N11275, N9628);
xor XOR2 (N11279, N11277, N1559);
or OR2 (N11280, N11278, N9898);
and AND4 (N11281, N11279, N7447, N1324, N4600);
or OR2 (N11282, N11274, N1506);
or OR3 (N11283, N11269, N6968, N928);
buf BUF1 (N11284, N11283);
nand NAND3 (N11285, N11281, N9897, N2781);
xor XOR2 (N11286, N11284, N5124);
or OR2 (N11287, N11267, N2082);
xor XOR2 (N11288, N11265, N7323);
nor NOR2 (N11289, N11286, N7219);
or OR4 (N11290, N11289, N11261, N5205, N2612);
and AND2 (N11291, N11290, N6831);
nor NOR3 (N11292, N11282, N2970, N8053);
buf BUF1 (N11293, N11273);
not NOT1 (N11294, N11288);
xor XOR2 (N11295, N11292, N3124);
buf BUF1 (N11296, N11276);
xor XOR2 (N11297, N11270, N3910);
buf BUF1 (N11298, N11280);
nor NOR2 (N11299, N11294, N8709);
or OR2 (N11300, N11285, N4131);
nand NAND3 (N11301, N11298, N10547, N2645);
buf BUF1 (N11302, N11291);
not NOT1 (N11303, N11293);
nor NOR2 (N11304, N11295, N2824);
xor XOR2 (N11305, N11287, N1693);
or OR2 (N11306, N11297, N8533);
nor NOR3 (N11307, N11302, N8096, N3813);
xor XOR2 (N11308, N11303, N7737);
nand NAND3 (N11309, N11306, N9777, N8541);
or OR3 (N11310, N11301, N1138, N4800);
or OR4 (N11311, N11308, N5356, N2000, N2537);
nand NAND2 (N11312, N11310, N5663);
buf BUF1 (N11313, N11300);
nand NAND4 (N11314, N11307, N3992, N8896, N346);
xor XOR2 (N11315, N11304, N3539);
nand NAND3 (N11316, N11313, N1421, N2865);
and AND2 (N11317, N11299, N7067);
or OR2 (N11318, N11312, N4876);
or OR3 (N11319, N11318, N9673, N5179);
or OR4 (N11320, N11319, N6003, N1151, N8771);
nor NOR2 (N11321, N11309, N10911);
and AND3 (N11322, N11317, N9595, N3742);
nand NAND4 (N11323, N11296, N6065, N7671, N6277);
not NOT1 (N11324, N11305);
not NOT1 (N11325, N11323);
xor XOR2 (N11326, N11316, N9761);
nor NOR2 (N11327, N11311, N6971);
and AND4 (N11328, N11326, N807, N9236, N6002);
xor XOR2 (N11329, N11321, N3266);
and AND2 (N11330, N11325, N1736);
and AND4 (N11331, N11324, N11123, N2880, N9718);
or OR4 (N11332, N11329, N7077, N1873, N7495);
and AND4 (N11333, N11331, N8018, N4908, N6341);
not NOT1 (N11334, N11322);
or OR4 (N11335, N11332, N357, N6572, N6347);
xor XOR2 (N11336, N11314, N10570);
not NOT1 (N11337, N11315);
not NOT1 (N11338, N11336);
not NOT1 (N11339, N11272);
nor NOR2 (N11340, N11327, N393);
or OR4 (N11341, N11338, N5304, N1903, N4253);
not NOT1 (N11342, N11340);
nor NOR2 (N11343, N11337, N6522);
buf BUF1 (N11344, N11339);
not NOT1 (N11345, N11335);
not NOT1 (N11346, N11342);
or OR2 (N11347, N11328, N1562);
or OR3 (N11348, N11330, N9725, N9077);
or OR4 (N11349, N11344, N2980, N7300, N183);
xor XOR2 (N11350, N11341, N6070);
not NOT1 (N11351, N11346);
nor NOR2 (N11352, N11345, N8672);
and AND4 (N11353, N11351, N2746, N1712, N482);
nand NAND3 (N11354, N11343, N10253, N6414);
buf BUF1 (N11355, N11352);
buf BUF1 (N11356, N11347);
nand NAND3 (N11357, N11356, N7868, N10436);
not NOT1 (N11358, N11355);
and AND3 (N11359, N11349, N9141, N1162);
and AND2 (N11360, N11354, N6705);
or OR4 (N11361, N11357, N622, N823, N6122);
and AND3 (N11362, N11360, N2628, N4179);
not NOT1 (N11363, N11320);
nor NOR4 (N11364, N11348, N1338, N8088, N8033);
or OR2 (N11365, N11362, N1051);
and AND3 (N11366, N11359, N3706, N4701);
not NOT1 (N11367, N11334);
not NOT1 (N11368, N11358);
buf BUF1 (N11369, N11366);
xor XOR2 (N11370, N11369, N7188);
nor NOR2 (N11371, N11370, N10770);
buf BUF1 (N11372, N11364);
xor XOR2 (N11373, N11372, N9777);
and AND2 (N11374, N11373, N8096);
buf BUF1 (N11375, N11368);
xor XOR2 (N11376, N11375, N5427);
nand NAND4 (N11377, N11350, N8635, N849, N171);
buf BUF1 (N11378, N11374);
not NOT1 (N11379, N11377);
buf BUF1 (N11380, N11376);
buf BUF1 (N11381, N11363);
and AND4 (N11382, N11371, N6017, N8886, N9760);
buf BUF1 (N11383, N11382);
and AND4 (N11384, N11380, N8497, N2557, N2138);
not NOT1 (N11385, N11353);
or OR3 (N11386, N11384, N4197, N10009);
nand NAND2 (N11387, N11383, N7505);
buf BUF1 (N11388, N11365);
or OR4 (N11389, N11379, N2075, N7390, N3834);
nand NAND3 (N11390, N11387, N4872, N7841);
buf BUF1 (N11391, N11361);
not NOT1 (N11392, N11386);
and AND3 (N11393, N11388, N10432, N1507);
not NOT1 (N11394, N11381);
buf BUF1 (N11395, N11367);
or OR3 (N11396, N11389, N10140, N3041);
not NOT1 (N11397, N11333);
nand NAND4 (N11398, N11395, N9324, N6495, N8654);
or OR3 (N11399, N11392, N4262, N1400);
nor NOR3 (N11400, N11390, N5103, N4980);
and AND4 (N11401, N11393, N2511, N6433, N2178);
or OR3 (N11402, N11398, N3129, N915);
not NOT1 (N11403, N11397);
buf BUF1 (N11404, N11378);
nor NOR3 (N11405, N11401, N2973, N19);
not NOT1 (N11406, N11394);
nand NAND3 (N11407, N11404, N9888, N6460);
not NOT1 (N11408, N11385);
or OR4 (N11409, N11400, N1958, N1933, N6760);
xor XOR2 (N11410, N11409, N187);
or OR3 (N11411, N11391, N5344, N11141);
nor NOR4 (N11412, N11407, N9100, N8581, N1843);
xor XOR2 (N11413, N11402, N7586);
and AND2 (N11414, N11408, N3594);
nor NOR3 (N11415, N11414, N11405, N8550);
nand NAND3 (N11416, N4968, N7497, N11408);
buf BUF1 (N11417, N11399);
buf BUF1 (N11418, N11406);
xor XOR2 (N11419, N11412, N6136);
xor XOR2 (N11420, N11413, N10435);
nand NAND2 (N11421, N11417, N10583);
and AND4 (N11422, N11411, N768, N8764, N4591);
or OR2 (N11423, N11403, N3704);
nor NOR2 (N11424, N11418, N2270);
nor NOR2 (N11425, N11416, N3492);
not NOT1 (N11426, N11425);
and AND2 (N11427, N11396, N11101);
nor NOR3 (N11428, N11410, N8121, N5565);
nor NOR4 (N11429, N11427, N8088, N6137, N8104);
xor XOR2 (N11430, N11419, N3343);
or OR4 (N11431, N11430, N6142, N6195, N6739);
nor NOR2 (N11432, N11426, N9999);
nor NOR2 (N11433, N11415, N953);
xor XOR2 (N11434, N11423, N10781);
not NOT1 (N11435, N11431);
or OR3 (N11436, N11432, N4239, N4747);
xor XOR2 (N11437, N11428, N10173);
not NOT1 (N11438, N11422);
nor NOR2 (N11439, N11434, N4732);
or OR3 (N11440, N11437, N1043, N1761);
nand NAND2 (N11441, N11429, N1408);
and AND3 (N11442, N11441, N10146, N9927);
buf BUF1 (N11443, N11436);
and AND4 (N11444, N11421, N5288, N6957, N9277);
xor XOR2 (N11445, N11424, N1911);
and AND2 (N11446, N11443, N4714);
and AND2 (N11447, N11420, N9274);
nand NAND2 (N11448, N11439, N6796);
and AND2 (N11449, N11433, N5208);
nand NAND4 (N11450, N11448, N7592, N341, N1371);
xor XOR2 (N11451, N11447, N4946);
xor XOR2 (N11452, N11442, N8817);
or OR4 (N11453, N11446, N7495, N6506, N9158);
nor NOR4 (N11454, N11450, N3786, N6156, N10776);
buf BUF1 (N11455, N11453);
nand NAND3 (N11456, N11435, N9545, N6503);
xor XOR2 (N11457, N11440, N5814);
or OR3 (N11458, N11452, N3580, N9334);
and AND2 (N11459, N11455, N9875);
buf BUF1 (N11460, N11451);
and AND3 (N11461, N11456, N6513, N3851);
not NOT1 (N11462, N11449);
not NOT1 (N11463, N11461);
xor XOR2 (N11464, N11462, N6618);
or OR3 (N11465, N11454, N6030, N7457);
nand NAND2 (N11466, N11460, N6698);
xor XOR2 (N11467, N11445, N7519);
nand NAND3 (N11468, N11444, N776, N6603);
and AND3 (N11469, N11465, N6289, N9009);
or OR3 (N11470, N11468, N5243, N7269);
or OR3 (N11471, N11466, N10490, N3420);
or OR4 (N11472, N11463, N10674, N3848, N10457);
nand NAND3 (N11473, N11458, N6821, N2315);
not NOT1 (N11474, N11438);
nor NOR3 (N11475, N11472, N4099, N132);
nor NOR3 (N11476, N11467, N6814, N4366);
nand NAND3 (N11477, N11470, N5739, N6623);
not NOT1 (N11478, N11476);
not NOT1 (N11479, N11474);
or OR3 (N11480, N11477, N11219, N852);
nand NAND2 (N11481, N11478, N342);
nor NOR2 (N11482, N11475, N180);
xor XOR2 (N11483, N11473, N4498);
buf BUF1 (N11484, N11464);
or OR4 (N11485, N11457, N1217, N2438, N3580);
or OR3 (N11486, N11481, N9395, N8414);
xor XOR2 (N11487, N11471, N6563);
buf BUF1 (N11488, N11479);
or OR3 (N11489, N11484, N2695, N2812);
nor NOR3 (N11490, N11483, N9937, N2032);
nand NAND4 (N11491, N11490, N8726, N6225, N7891);
not NOT1 (N11492, N11459);
xor XOR2 (N11493, N11469, N637);
or OR2 (N11494, N11487, N9888);
buf BUF1 (N11495, N11482);
nand NAND4 (N11496, N11491, N7420, N2297, N3539);
and AND2 (N11497, N11494, N2935);
buf BUF1 (N11498, N11488);
or OR4 (N11499, N11485, N4779, N5304, N4865);
nand NAND4 (N11500, N11498, N1354, N3076, N7272);
nor NOR3 (N11501, N11495, N320, N7251);
buf BUF1 (N11502, N11501);
not NOT1 (N11503, N11497);
not NOT1 (N11504, N11480);
not NOT1 (N11505, N11493);
buf BUF1 (N11506, N11504);
and AND3 (N11507, N11503, N5212, N6732);
not NOT1 (N11508, N11492);
xor XOR2 (N11509, N11496, N11450);
nand NAND4 (N11510, N11507, N5259, N6945, N7507);
not NOT1 (N11511, N11500);
and AND4 (N11512, N11509, N10948, N6771, N8267);
buf BUF1 (N11513, N11499);
xor XOR2 (N11514, N11486, N3035);
and AND4 (N11515, N11510, N9723, N7257, N1470);
nand NAND4 (N11516, N11502, N4173, N9874, N797);
nor NOR3 (N11517, N11512, N9289, N8399);
nand NAND2 (N11518, N11506, N4792);
not NOT1 (N11519, N11513);
buf BUF1 (N11520, N11518);
nand NAND4 (N11521, N11505, N2533, N6446, N1967);
buf BUF1 (N11522, N11519);
or OR4 (N11523, N11516, N6364, N5951, N8186);
xor XOR2 (N11524, N11517, N164);
xor XOR2 (N11525, N11515, N6803);
nor NOR4 (N11526, N11524, N9651, N4746, N878);
not NOT1 (N11527, N11508);
xor XOR2 (N11528, N11489, N7816);
and AND4 (N11529, N11525, N7631, N4886, N9961);
not NOT1 (N11530, N11528);
or OR2 (N11531, N11529, N10778);
xor XOR2 (N11532, N11521, N5858);
xor XOR2 (N11533, N11531, N8636);
nor NOR4 (N11534, N11523, N5651, N10747, N3937);
or OR2 (N11535, N11534, N5693);
nand NAND4 (N11536, N11527, N4878, N629, N9227);
and AND3 (N11537, N11533, N2431, N9352);
not NOT1 (N11538, N11537);
buf BUF1 (N11539, N11514);
nand NAND2 (N11540, N11522, N9653);
xor XOR2 (N11541, N11532, N6410);
xor XOR2 (N11542, N11540, N9092);
nor NOR2 (N11543, N11539, N5736);
xor XOR2 (N11544, N11541, N3833);
nand NAND4 (N11545, N11542, N509, N8329, N3676);
nor NOR3 (N11546, N11530, N10624, N5220);
and AND2 (N11547, N11511, N8025);
buf BUF1 (N11548, N11544);
not NOT1 (N11549, N11535);
nor NOR2 (N11550, N11547, N776);
nand NAND2 (N11551, N11550, N5284);
and AND2 (N11552, N11551, N3863);
buf BUF1 (N11553, N11545);
xor XOR2 (N11554, N11552, N7341);
and AND3 (N11555, N11543, N6216, N7843);
xor XOR2 (N11556, N11536, N1520);
nand NAND3 (N11557, N11549, N10764, N10465);
xor XOR2 (N11558, N11548, N7770);
xor XOR2 (N11559, N11520, N7869);
not NOT1 (N11560, N11556);
or OR3 (N11561, N11559, N7143, N831);
buf BUF1 (N11562, N11538);
or OR4 (N11563, N11555, N377, N6630, N9486);
not NOT1 (N11564, N11562);
xor XOR2 (N11565, N11526, N3059);
or OR3 (N11566, N11546, N10769, N2960);
and AND4 (N11567, N11561, N7033, N4562, N2225);
and AND2 (N11568, N11565, N2515);
or OR3 (N11569, N11564, N8195, N2492);
and AND4 (N11570, N11563, N2653, N3714, N10318);
and AND2 (N11571, N11558, N2730);
and AND4 (N11572, N11569, N4631, N390, N9241);
nor NOR4 (N11573, N11566, N1709, N7151, N2884);
not NOT1 (N11574, N11567);
and AND4 (N11575, N11560, N5321, N7124, N5694);
nor NOR4 (N11576, N11568, N6183, N6694, N6251);
and AND4 (N11577, N11573, N3904, N3638, N634);
and AND3 (N11578, N11571, N3395, N4098);
or OR3 (N11579, N11575, N3411, N9892);
buf BUF1 (N11580, N11557);
xor XOR2 (N11581, N11574, N11539);
and AND2 (N11582, N11580, N4082);
and AND3 (N11583, N11577, N1221, N9488);
or OR4 (N11584, N11576, N8918, N1548, N10853);
not NOT1 (N11585, N11581);
and AND4 (N11586, N11583, N11228, N10202, N2232);
and AND4 (N11587, N11578, N6020, N2506, N7331);
nor NOR2 (N11588, N11586, N95);
buf BUF1 (N11589, N11587);
and AND2 (N11590, N11584, N9942);
and AND3 (N11591, N11585, N6573, N6527);
and AND2 (N11592, N11570, N10004);
or OR2 (N11593, N11553, N3522);
xor XOR2 (N11594, N11592, N3072);
buf BUF1 (N11595, N11591);
xor XOR2 (N11596, N11594, N6118);
or OR2 (N11597, N11589, N9701);
and AND4 (N11598, N11579, N9158, N4297, N5547);
and AND4 (N11599, N11595, N4124, N4927, N9679);
and AND4 (N11600, N11599, N11123, N2626, N6739);
xor XOR2 (N11601, N11572, N7256);
buf BUF1 (N11602, N11593);
buf BUF1 (N11603, N11590);
and AND3 (N11604, N11603, N3442, N5744);
and AND3 (N11605, N11597, N7271, N4411);
and AND3 (N11606, N11604, N9162, N6587);
nand NAND4 (N11607, N11588, N9225, N5274, N3989);
and AND4 (N11608, N11606, N3877, N4799, N5781);
nand NAND2 (N11609, N11602, N2059);
xor XOR2 (N11610, N11605, N5691);
xor XOR2 (N11611, N11609, N8190);
and AND3 (N11612, N11611, N3912, N1836);
xor XOR2 (N11613, N11608, N730);
or OR4 (N11614, N11554, N9684, N1954, N5904);
or OR3 (N11615, N11613, N679, N5906);
nor NOR2 (N11616, N11607, N9401);
not NOT1 (N11617, N11582);
xor XOR2 (N11618, N11600, N3713);
nand NAND3 (N11619, N11596, N10275, N2098);
nor NOR2 (N11620, N11617, N2619);
buf BUF1 (N11621, N11619);
xor XOR2 (N11622, N11612, N1120);
not NOT1 (N11623, N11598);
and AND3 (N11624, N11610, N2874, N7366);
buf BUF1 (N11625, N11618);
buf BUF1 (N11626, N11625);
nand NAND2 (N11627, N11614, N10038);
not NOT1 (N11628, N11615);
buf BUF1 (N11629, N11601);
buf BUF1 (N11630, N11623);
nand NAND2 (N11631, N11620, N6716);
and AND4 (N11632, N11621, N2580, N10982, N10736);
nor NOR3 (N11633, N11629, N7380, N2551);
and AND4 (N11634, N11630, N2149, N599, N4785);
or OR3 (N11635, N11634, N9667, N7168);
nand NAND4 (N11636, N11616, N8180, N11608, N10773);
nand NAND2 (N11637, N11628, N3124);
buf BUF1 (N11638, N11635);
or OR2 (N11639, N11626, N9968);
not NOT1 (N11640, N11636);
and AND2 (N11641, N11627, N7090);
nand NAND2 (N11642, N11631, N3580);
or OR4 (N11643, N11639, N7120, N7500, N1004);
nand NAND3 (N11644, N11632, N7015, N9501);
buf BUF1 (N11645, N11640);
or OR3 (N11646, N11624, N108, N4092);
xor XOR2 (N11647, N11643, N9473);
nand NAND2 (N11648, N11637, N2495);
buf BUF1 (N11649, N11641);
buf BUF1 (N11650, N11642);
xor XOR2 (N11651, N11645, N5958);
not NOT1 (N11652, N11644);
nand NAND4 (N11653, N11648, N3216, N4346, N5505);
nand NAND4 (N11654, N11651, N11489, N3283, N11212);
xor XOR2 (N11655, N11653, N11153);
nor NOR2 (N11656, N11647, N2221);
and AND3 (N11657, N11654, N2124, N8749);
nand NAND4 (N11658, N11649, N3451, N10368, N9123);
nor NOR4 (N11659, N11658, N5888, N815, N5700);
and AND4 (N11660, N11622, N7422, N4321, N10429);
buf BUF1 (N11661, N11633);
xor XOR2 (N11662, N11661, N10177);
not NOT1 (N11663, N11659);
and AND2 (N11664, N11662, N5381);
nand NAND2 (N11665, N11652, N5055);
not NOT1 (N11666, N11663);
and AND4 (N11667, N11665, N7131, N1080, N10181);
nand NAND3 (N11668, N11650, N5282, N9850);
nor NOR3 (N11669, N11655, N8322, N10158);
buf BUF1 (N11670, N11638);
and AND2 (N11671, N11664, N6008);
nor NOR2 (N11672, N11670, N9613);
or OR4 (N11673, N11656, N6950, N8769, N7082);
xor XOR2 (N11674, N11646, N7252);
buf BUF1 (N11675, N11671);
not NOT1 (N11676, N11667);
and AND3 (N11677, N11669, N8721, N7751);
xor XOR2 (N11678, N11672, N186);
and AND3 (N11679, N11675, N2820, N3129);
and AND3 (N11680, N11677, N6741, N1416);
nand NAND2 (N11681, N11678, N610);
or OR2 (N11682, N11660, N11073);
xor XOR2 (N11683, N11676, N11027);
or OR3 (N11684, N11668, N6196, N5628);
nor NOR4 (N11685, N11681, N3139, N4402, N6162);
not NOT1 (N11686, N11682);
nand NAND2 (N11687, N11673, N10436);
buf BUF1 (N11688, N11685);
or OR3 (N11689, N11688, N3775, N3059);
xor XOR2 (N11690, N11666, N4640);
buf BUF1 (N11691, N11687);
buf BUF1 (N11692, N11690);
buf BUF1 (N11693, N11657);
buf BUF1 (N11694, N11686);
nor NOR2 (N11695, N11679, N7835);
nor NOR2 (N11696, N11691, N6530);
nor NOR2 (N11697, N11689, N3482);
or OR3 (N11698, N11696, N8234, N2447);
nor NOR2 (N11699, N11697, N3762);
or OR4 (N11700, N11698, N2193, N3684, N3693);
or OR4 (N11701, N11694, N2926, N7970, N8301);
or OR3 (N11702, N11701, N7097, N8065);
and AND2 (N11703, N11683, N10290);
or OR3 (N11704, N11703, N1421, N10596);
nor NOR2 (N11705, N11700, N4933);
or OR2 (N11706, N11704, N7382);
nor NOR2 (N11707, N11706, N384);
and AND4 (N11708, N11707, N6207, N7481, N6340);
nor NOR4 (N11709, N11708, N10333, N881, N10342);
and AND2 (N11710, N11695, N6849);
and AND4 (N11711, N11699, N10025, N1610, N1657);
xor XOR2 (N11712, N11711, N1702);
and AND4 (N11713, N11710, N2316, N7455, N9696);
and AND4 (N11714, N11709, N1020, N10939, N3132);
xor XOR2 (N11715, N11693, N2470);
nor NOR2 (N11716, N11705, N9454);
nor NOR2 (N11717, N11674, N3165);
not NOT1 (N11718, N11692);
nand NAND4 (N11719, N11712, N5721, N5961, N4763);
not NOT1 (N11720, N11715);
not NOT1 (N11721, N11680);
not NOT1 (N11722, N11716);
buf BUF1 (N11723, N11719);
buf BUF1 (N11724, N11721);
xor XOR2 (N11725, N11702, N6000);
nand NAND4 (N11726, N11724, N1988, N2142, N4997);
buf BUF1 (N11727, N11713);
or OR3 (N11728, N11727, N9416, N776);
or OR4 (N11729, N11714, N8912, N11222, N8907);
xor XOR2 (N11730, N11723, N6091);
nand NAND3 (N11731, N11720, N10592, N1733);
and AND2 (N11732, N11718, N4691);
nor NOR2 (N11733, N11684, N867);
or OR2 (N11734, N11728, N8202);
or OR4 (N11735, N11729, N11300, N3191, N2239);
and AND4 (N11736, N11734, N213, N2441, N9628);
nor NOR4 (N11737, N11726, N5738, N7232, N3953);
or OR3 (N11738, N11735, N284, N5205);
and AND4 (N11739, N11730, N11161, N1683, N8660);
nor NOR4 (N11740, N11725, N6001, N2385, N2963);
nand NAND4 (N11741, N11740, N6478, N4049, N6330);
xor XOR2 (N11742, N11737, N601);
xor XOR2 (N11743, N11741, N5784);
and AND4 (N11744, N11739, N5586, N5400, N4096);
not NOT1 (N11745, N11733);
nand NAND2 (N11746, N11738, N8500);
not NOT1 (N11747, N11743);
buf BUF1 (N11748, N11746);
xor XOR2 (N11749, N11722, N8128);
nand NAND2 (N11750, N11748, N7500);
not NOT1 (N11751, N11732);
nand NAND2 (N11752, N11717, N2987);
buf BUF1 (N11753, N11752);
or OR3 (N11754, N11751, N7942, N1046);
or OR3 (N11755, N11747, N9764, N8994);
buf BUF1 (N11756, N11736);
xor XOR2 (N11757, N11731, N6803);
and AND4 (N11758, N11750, N4280, N193, N4015);
nand NAND3 (N11759, N11758, N256, N11079);
xor XOR2 (N11760, N11759, N8178);
not NOT1 (N11761, N11753);
and AND2 (N11762, N11749, N9922);
not NOT1 (N11763, N11761);
nor NOR3 (N11764, N11744, N4418, N11453);
nand NAND2 (N11765, N11755, N1945);
buf BUF1 (N11766, N11760);
nor NOR4 (N11767, N11762, N4415, N8826, N7154);
and AND3 (N11768, N11756, N9457, N7273);
nor NOR3 (N11769, N11765, N7692, N3175);
nor NOR2 (N11770, N11745, N4155);
or OR4 (N11771, N11766, N4292, N5790, N612);
and AND4 (N11772, N11742, N7452, N4634, N7440);
buf BUF1 (N11773, N11767);
and AND2 (N11774, N11770, N6226);
nand NAND2 (N11775, N11768, N3518);
buf BUF1 (N11776, N11764);
buf BUF1 (N11777, N11754);
nand NAND2 (N11778, N11775, N8319);
or OR4 (N11779, N11757, N11426, N5876, N10352);
and AND2 (N11780, N11773, N5567);
xor XOR2 (N11781, N11772, N752);
not NOT1 (N11782, N11769);
and AND4 (N11783, N11763, N6616, N5486, N1119);
nand NAND4 (N11784, N11771, N7589, N7132, N2294);
and AND4 (N11785, N11784, N1253, N7179, N7444);
nor NOR4 (N11786, N11776, N5314, N11486, N10873);
xor XOR2 (N11787, N11778, N4498);
not NOT1 (N11788, N11777);
not NOT1 (N11789, N11785);
nand NAND4 (N11790, N11781, N5569, N6464, N3498);
or OR2 (N11791, N11789, N4456);
not NOT1 (N11792, N11791);
and AND3 (N11793, N11788, N9434, N11604);
xor XOR2 (N11794, N11780, N490);
buf BUF1 (N11795, N11790);
nor NOR4 (N11796, N11794, N4309, N8102, N11749);
or OR2 (N11797, N11783, N8907);
buf BUF1 (N11798, N11779);
and AND2 (N11799, N11797, N9203);
nor NOR4 (N11800, N11795, N40, N609, N2901);
or OR4 (N11801, N11799, N1850, N5189, N8066);
nand NAND2 (N11802, N11796, N10747);
not NOT1 (N11803, N11798);
or OR4 (N11804, N11793, N10868, N6886, N2503);
nand NAND4 (N11805, N11786, N1663, N7618, N11047);
nor NOR2 (N11806, N11802, N2293);
xor XOR2 (N11807, N11803, N219);
xor XOR2 (N11808, N11774, N8511);
nor NOR4 (N11809, N11807, N7244, N11631, N9204);
and AND4 (N11810, N11782, N9018, N3872, N3162);
nand NAND3 (N11811, N11808, N1391, N3370);
and AND4 (N11812, N11806, N8464, N7552, N10564);
not NOT1 (N11813, N11801);
xor XOR2 (N11814, N11809, N117);
nand NAND2 (N11815, N11804, N3076);
nand NAND4 (N11816, N11814, N10559, N6108, N9324);
nor NOR2 (N11817, N11800, N3609);
nor NOR3 (N11818, N11816, N11387, N6586);
xor XOR2 (N11819, N11812, N4704);
and AND4 (N11820, N11819, N3399, N2638, N144);
nand NAND4 (N11821, N11805, N2834, N481, N8303);
xor XOR2 (N11822, N11813, N5525);
or OR3 (N11823, N11810, N10575, N9939);
nand NAND3 (N11824, N11787, N3771, N1351);
xor XOR2 (N11825, N11822, N2377);
buf BUF1 (N11826, N11818);
and AND3 (N11827, N11815, N9269, N9193);
and AND3 (N11828, N11820, N1360, N10733);
or OR4 (N11829, N11824, N1072, N3852, N4116);
or OR2 (N11830, N11825, N6387);
not NOT1 (N11831, N11817);
nand NAND4 (N11832, N11792, N11814, N5570, N3740);
or OR3 (N11833, N11823, N2187, N745);
not NOT1 (N11834, N11830);
and AND3 (N11835, N11828, N1280, N10140);
and AND4 (N11836, N11833, N6169, N10321, N7223);
not NOT1 (N11837, N11831);
or OR2 (N11838, N11835, N1364);
buf BUF1 (N11839, N11838);
nor NOR3 (N11840, N11827, N8763, N5255);
xor XOR2 (N11841, N11839, N5817);
buf BUF1 (N11842, N11836);
and AND2 (N11843, N11837, N8395);
nand NAND2 (N11844, N11840, N10177);
buf BUF1 (N11845, N11844);
buf BUF1 (N11846, N11829);
and AND3 (N11847, N11826, N5560, N10229);
or OR4 (N11848, N11842, N2779, N11133, N3376);
nand NAND2 (N11849, N11841, N983);
not NOT1 (N11850, N11846);
not NOT1 (N11851, N11821);
or OR4 (N11852, N11851, N4440, N5502, N10719);
or OR2 (N11853, N11834, N3037);
or OR4 (N11854, N11848, N8630, N816, N6415);
or OR3 (N11855, N11811, N147, N5759);
and AND4 (N11856, N11850, N8769, N5045, N10986);
or OR3 (N11857, N11854, N1513, N4921);
nor NOR4 (N11858, N11847, N8698, N1507, N10146);
buf BUF1 (N11859, N11856);
nand NAND4 (N11860, N11845, N5233, N7081, N7749);
nand NAND2 (N11861, N11857, N5926);
buf BUF1 (N11862, N11861);
and AND3 (N11863, N11855, N3894, N8243);
xor XOR2 (N11864, N11862, N5786);
and AND4 (N11865, N11863, N11646, N7291, N11377);
or OR2 (N11866, N11864, N2157);
buf BUF1 (N11867, N11865);
and AND3 (N11868, N11867, N2703, N843);
nand NAND3 (N11869, N11832, N369, N6918);
not NOT1 (N11870, N11869);
or OR4 (N11871, N11858, N6366, N9520, N4907);
and AND3 (N11872, N11852, N8784, N10991);
or OR4 (N11873, N11872, N6701, N8696, N1439);
nand NAND3 (N11874, N11866, N1713, N8036);
nor NOR4 (N11875, N11853, N9231, N10866, N11874);
not NOT1 (N11876, N3087);
nor NOR2 (N11877, N11875, N4492);
buf BUF1 (N11878, N11873);
not NOT1 (N11879, N11871);
nand NAND3 (N11880, N11877, N3578, N3459);
nand NAND3 (N11881, N11859, N11700, N4113);
and AND3 (N11882, N11881, N8566, N2413);
nor NOR4 (N11883, N11879, N141, N6351, N6305);
xor XOR2 (N11884, N11880, N2248);
and AND3 (N11885, N11870, N560, N5140);
not NOT1 (N11886, N11882);
nand NAND2 (N11887, N11885, N4043);
nor NOR4 (N11888, N11884, N924, N2550, N11697);
buf BUF1 (N11889, N11887);
buf BUF1 (N11890, N11868);
and AND3 (N11891, N11878, N351, N4839);
nor NOR4 (N11892, N11860, N10746, N5661, N11022);
and AND3 (N11893, N11890, N1629, N5548);
buf BUF1 (N11894, N11891);
xor XOR2 (N11895, N11883, N8686);
or OR4 (N11896, N11889, N10411, N7305, N10502);
or OR2 (N11897, N11843, N9054);
xor XOR2 (N11898, N11876, N3638);
nand NAND3 (N11899, N11893, N2305, N3986);
xor XOR2 (N11900, N11888, N735);
xor XOR2 (N11901, N11897, N1912);
not NOT1 (N11902, N11901);
or OR4 (N11903, N11898, N10220, N3444, N1139);
buf BUF1 (N11904, N11894);
nand NAND3 (N11905, N11886, N6620, N2512);
xor XOR2 (N11906, N11904, N9863);
nand NAND4 (N11907, N11849, N3251, N4483, N4738);
nand NAND2 (N11908, N11902, N8506);
nor NOR2 (N11909, N11905, N9119);
nand NAND4 (N11910, N11908, N4416, N5284, N11174);
xor XOR2 (N11911, N11907, N106);
buf BUF1 (N11912, N11896);
nor NOR4 (N11913, N11899, N2844, N528, N9156);
nor NOR4 (N11914, N11911, N4032, N6557, N8060);
or OR4 (N11915, N11913, N4602, N6792, N9957);
xor XOR2 (N11916, N11914, N4460);
or OR4 (N11917, N11900, N10657, N10397, N6773);
or OR2 (N11918, N11906, N3223);
and AND2 (N11919, N11910, N342);
nand NAND3 (N11920, N11917, N8669, N343);
buf BUF1 (N11921, N11909);
nand NAND2 (N11922, N11918, N11402);
buf BUF1 (N11923, N11895);
not NOT1 (N11924, N11923);
and AND2 (N11925, N11924, N2189);
nand NAND2 (N11926, N11922, N3440);
nand NAND4 (N11927, N11925, N2276, N3497, N4298);
and AND2 (N11928, N11927, N1373);
buf BUF1 (N11929, N11921);
nor NOR4 (N11930, N11926, N1368, N4373, N1832);
not NOT1 (N11931, N11903);
buf BUF1 (N11932, N11931);
or OR2 (N11933, N11919, N2855);
nand NAND2 (N11934, N11930, N4696);
nand NAND3 (N11935, N11912, N5394, N11323);
and AND3 (N11936, N11935, N4088, N9128);
and AND2 (N11937, N11892, N7039);
nand NAND3 (N11938, N11934, N3296, N6628);
nand NAND2 (N11939, N11929, N4685);
xor XOR2 (N11940, N11936, N6258);
nand NAND2 (N11941, N11939, N364);
not NOT1 (N11942, N11916);
xor XOR2 (N11943, N11940, N11260);
nand NAND4 (N11944, N11943, N2203, N3115, N10663);
and AND4 (N11945, N11933, N9728, N2042, N3583);
nand NAND2 (N11946, N11941, N4939);
nand NAND4 (N11947, N11932, N5137, N1719, N805);
not NOT1 (N11948, N11945);
nand NAND2 (N11949, N11937, N11871);
xor XOR2 (N11950, N11928, N9985);
and AND2 (N11951, N11946, N9596);
xor XOR2 (N11952, N11920, N4922);
xor XOR2 (N11953, N11947, N6091);
buf BUF1 (N11954, N11948);
not NOT1 (N11955, N11938);
xor XOR2 (N11956, N11954, N8449);
nand NAND2 (N11957, N11950, N11898);
nand NAND3 (N11958, N11915, N11483, N2824);
nand NAND4 (N11959, N11952, N8425, N7931, N9070);
not NOT1 (N11960, N11956);
buf BUF1 (N11961, N11953);
and AND4 (N11962, N11957, N7668, N8336, N10717);
or OR4 (N11963, N11949, N6687, N4572, N1740);
not NOT1 (N11964, N11942);
xor XOR2 (N11965, N11959, N5207);
nor NOR2 (N11966, N11951, N6738);
buf BUF1 (N11967, N11966);
not NOT1 (N11968, N11964);
not NOT1 (N11969, N11958);
or OR2 (N11970, N11963, N11059);
nor NOR3 (N11971, N11967, N6756, N4114);
and AND4 (N11972, N11960, N2743, N5620, N5449);
and AND2 (N11973, N11968, N531);
or OR3 (N11974, N11972, N5627, N2658);
and AND3 (N11975, N11955, N8466, N6984);
xor XOR2 (N11976, N11944, N4866);
nor NOR3 (N11977, N11970, N2302, N11320);
not NOT1 (N11978, N11961);
or OR3 (N11979, N11971, N3159, N1475);
nand NAND3 (N11980, N11977, N439, N7115);
xor XOR2 (N11981, N11974, N3370);
and AND3 (N11982, N11978, N5825, N11892);
xor XOR2 (N11983, N11965, N3271);
xor XOR2 (N11984, N11975, N6745);
nor NOR4 (N11985, N11969, N15, N7924, N11695);
or OR4 (N11986, N11984, N10184, N10736, N9839);
nand NAND3 (N11987, N11986, N10264, N4453);
buf BUF1 (N11988, N11980);
and AND3 (N11989, N11983, N2000, N1520);
xor XOR2 (N11990, N11987, N5850);
not NOT1 (N11991, N11982);
or OR4 (N11992, N11988, N6072, N4586, N4103);
not NOT1 (N11993, N11981);
or OR2 (N11994, N11962, N88);
or OR2 (N11995, N11973, N6232);
and AND3 (N11996, N11989, N9486, N4763);
buf BUF1 (N11997, N11985);
not NOT1 (N11998, N11992);
and AND4 (N11999, N11997, N9371, N10931, N10268);
nor NOR3 (N12000, N11996, N7564, N2226);
nor NOR4 (N12001, N11991, N4860, N2345, N7593);
buf BUF1 (N12002, N11999);
nand NAND2 (N12003, N11993, N7099);
nand NAND4 (N12004, N12000, N8779, N10939, N9127);
nor NOR3 (N12005, N12004, N9564, N768);
nor NOR2 (N12006, N11998, N8435);
and AND2 (N12007, N12006, N9004);
nand NAND4 (N12008, N12007, N2718, N204, N8468);
nor NOR4 (N12009, N12008, N10460, N3738, N1540);
buf BUF1 (N12010, N11994);
and AND2 (N12011, N12009, N5976);
nor NOR3 (N12012, N12003, N10222, N4485);
xor XOR2 (N12013, N11976, N1258);
or OR2 (N12014, N12002, N7606);
and AND3 (N12015, N12001, N7738, N11344);
and AND3 (N12016, N12012, N11255, N9402);
nor NOR4 (N12017, N11990, N8691, N7227, N6879);
nor NOR4 (N12018, N11995, N318, N10881, N2844);
nor NOR4 (N12019, N12017, N9454, N2908, N1940);
nor NOR3 (N12020, N12010, N7555, N11622);
or OR3 (N12021, N12018, N1417, N3277);
not NOT1 (N12022, N12020);
nor NOR2 (N12023, N12021, N6510);
or OR4 (N12024, N12005, N3486, N3586, N4185);
nand NAND4 (N12025, N12014, N307, N1882, N9771);
not NOT1 (N12026, N12013);
nor NOR3 (N12027, N12016, N946, N6370);
or OR3 (N12028, N12015, N9413, N7260);
nor NOR4 (N12029, N12024, N2789, N4205, N5232);
and AND4 (N12030, N12019, N9434, N863, N552);
or OR3 (N12031, N12022, N3713, N954);
or OR3 (N12032, N12029, N4222, N7162);
and AND2 (N12033, N11979, N10680);
not NOT1 (N12034, N12025);
nor NOR4 (N12035, N12033, N207, N4772, N4818);
buf BUF1 (N12036, N12027);
nand NAND4 (N12037, N12026, N6347, N5682, N9829);
buf BUF1 (N12038, N12036);
or OR2 (N12039, N12034, N6292);
buf BUF1 (N12040, N12032);
xor XOR2 (N12041, N12030, N7314);
nor NOR2 (N12042, N12023, N6132);
nor NOR2 (N12043, N12038, N9638);
nand NAND3 (N12044, N12043, N5599, N11481);
and AND2 (N12045, N12041, N5880);
nor NOR4 (N12046, N12042, N8016, N2133, N3828);
buf BUF1 (N12047, N12044);
not NOT1 (N12048, N12028);
not NOT1 (N12049, N12045);
and AND3 (N12050, N12035, N7049, N10023);
or OR4 (N12051, N12049, N11440, N11769, N9804);
nand NAND3 (N12052, N12047, N11119, N7775);
nand NAND4 (N12053, N12037, N7795, N4764, N6805);
nand NAND3 (N12054, N12046, N10151, N11041);
buf BUF1 (N12055, N12053);
xor XOR2 (N12056, N12055, N7554);
not NOT1 (N12057, N12039);
nor NOR3 (N12058, N12054, N9270, N6077);
not NOT1 (N12059, N12011);
and AND4 (N12060, N12051, N7039, N1244, N9268);
or OR4 (N12061, N12060, N4028, N11252, N9269);
nor NOR4 (N12062, N12050, N10202, N6430, N6088);
nand NAND2 (N12063, N12058, N10304);
or OR4 (N12064, N12048, N10218, N4334, N1243);
and AND3 (N12065, N12063, N4131, N489);
xor XOR2 (N12066, N12057, N1530);
xor XOR2 (N12067, N12040, N7450);
xor XOR2 (N12068, N12064, N9986);
and AND4 (N12069, N12062, N4668, N899, N7874);
xor XOR2 (N12070, N12066, N327);
buf BUF1 (N12071, N12065);
not NOT1 (N12072, N12059);
not NOT1 (N12073, N12067);
or OR2 (N12074, N12071, N11024);
not NOT1 (N12075, N12072);
not NOT1 (N12076, N12069);
or OR4 (N12077, N12070, N1761, N11836, N4105);
or OR3 (N12078, N12052, N7413, N4345);
or OR4 (N12079, N12078, N3143, N11126, N7294);
xor XOR2 (N12080, N12079, N8667);
xor XOR2 (N12081, N12076, N5101);
xor XOR2 (N12082, N12077, N9842);
nand NAND3 (N12083, N12081, N3239, N5862);
buf BUF1 (N12084, N12074);
or OR4 (N12085, N12068, N572, N135, N6476);
xor XOR2 (N12086, N12031, N3521);
not NOT1 (N12087, N12061);
nor NOR3 (N12088, N12084, N3797, N8825);
buf BUF1 (N12089, N12080);
nand NAND2 (N12090, N12088, N9173);
not NOT1 (N12091, N12085);
nor NOR4 (N12092, N12087, N8497, N10950, N4806);
xor XOR2 (N12093, N12090, N1336);
and AND2 (N12094, N12082, N9410);
nand NAND2 (N12095, N12089, N6217);
not NOT1 (N12096, N12092);
buf BUF1 (N12097, N12096);
xor XOR2 (N12098, N12083, N11161);
and AND4 (N12099, N12086, N4846, N8887, N10056);
or OR2 (N12100, N12093, N8761);
nor NOR3 (N12101, N12099, N8618, N4106);
nor NOR2 (N12102, N12094, N2795);
or OR4 (N12103, N12095, N3031, N11326, N7583);
xor XOR2 (N12104, N12075, N9216);
not NOT1 (N12105, N12091);
and AND4 (N12106, N12098, N1665, N1231, N7001);
nand NAND4 (N12107, N12097, N4352, N10300, N810);
or OR2 (N12108, N12101, N9556);
xor XOR2 (N12109, N12106, N2492);
xor XOR2 (N12110, N12102, N9137);
xor XOR2 (N12111, N12105, N4326);
buf BUF1 (N12112, N12111);
not NOT1 (N12113, N12073);
nand NAND3 (N12114, N12109, N7872, N10416);
xor XOR2 (N12115, N12056, N10135);
xor XOR2 (N12116, N12107, N1506);
or OR3 (N12117, N12108, N8055, N4119);
nand NAND2 (N12118, N12110, N2552);
nor NOR4 (N12119, N12100, N9183, N2918, N8582);
and AND2 (N12120, N12118, N8288);
nor NOR2 (N12121, N12116, N4860);
nor NOR3 (N12122, N12117, N10335, N9040);
nand NAND3 (N12123, N12113, N4925, N1612);
buf BUF1 (N12124, N12122);
or OR2 (N12125, N12104, N44);
xor XOR2 (N12126, N12123, N7331);
xor XOR2 (N12127, N12124, N7189);
or OR4 (N12128, N12115, N5719, N1134, N2862);
and AND4 (N12129, N12112, N9479, N4385, N9684);
nor NOR3 (N12130, N12129, N11217, N7261);
not NOT1 (N12131, N12121);
xor XOR2 (N12132, N12130, N3562);
or OR3 (N12133, N12127, N4141, N10831);
nor NOR2 (N12134, N12126, N487);
xor XOR2 (N12135, N12132, N3156);
not NOT1 (N12136, N12131);
buf BUF1 (N12137, N12114);
or OR4 (N12138, N12103, N2665, N6535, N6281);
or OR4 (N12139, N12125, N754, N11068, N475);
or OR3 (N12140, N12135, N7225, N10740);
or OR2 (N12141, N12128, N9614);
nor NOR3 (N12142, N12140, N4930, N5979);
or OR2 (N12143, N12142, N4701);
buf BUF1 (N12144, N12136);
buf BUF1 (N12145, N12139);
xor XOR2 (N12146, N12138, N11082);
nor NOR2 (N12147, N12137, N10874);
not NOT1 (N12148, N12134);
nand NAND2 (N12149, N12146, N8105);
not NOT1 (N12150, N12120);
buf BUF1 (N12151, N12145);
nand NAND2 (N12152, N12151, N2830);
xor XOR2 (N12153, N12119, N8370);
or OR3 (N12154, N12141, N11373, N11527);
and AND3 (N12155, N12150, N4514, N4011);
xor XOR2 (N12156, N12144, N11953);
nor NOR2 (N12157, N12154, N6328);
xor XOR2 (N12158, N12149, N3687);
xor XOR2 (N12159, N12158, N7629);
and AND4 (N12160, N12153, N10513, N1451, N7681);
or OR3 (N12161, N12152, N7760, N4997);
nand NAND4 (N12162, N12148, N4370, N1889, N10077);
nand NAND3 (N12163, N12156, N11771, N10371);
or OR3 (N12164, N12147, N4384, N11330);
and AND3 (N12165, N12143, N8927, N4084);
xor XOR2 (N12166, N12161, N1669);
and AND2 (N12167, N12155, N9842);
and AND3 (N12168, N12167, N4706, N10140);
or OR4 (N12169, N12160, N1566, N3011, N11061);
nand NAND2 (N12170, N12163, N5398);
buf BUF1 (N12171, N12166);
nand NAND3 (N12172, N12168, N9007, N11455);
not NOT1 (N12173, N12164);
xor XOR2 (N12174, N12159, N11935);
not NOT1 (N12175, N12165);
nand NAND3 (N12176, N12172, N8379, N9038);
nand NAND4 (N12177, N12169, N9747, N2746, N4914);
xor XOR2 (N12178, N12177, N8225);
nor NOR4 (N12179, N12173, N10003, N1057, N4413);
xor XOR2 (N12180, N12174, N2846);
buf BUF1 (N12181, N12133);
or OR2 (N12182, N12178, N11684);
or OR2 (N12183, N12162, N3148);
nand NAND3 (N12184, N12180, N667, N8843);
xor XOR2 (N12185, N12171, N327);
xor XOR2 (N12186, N12157, N5439);
nor NOR3 (N12187, N12186, N2810, N267);
buf BUF1 (N12188, N12184);
xor XOR2 (N12189, N12182, N3282);
or OR3 (N12190, N12185, N6643, N1999);
xor XOR2 (N12191, N12190, N10553);
and AND4 (N12192, N12179, N2428, N764, N2234);
and AND3 (N12193, N12188, N2048, N12145);
buf BUF1 (N12194, N12176);
nor NOR3 (N12195, N12187, N6009, N5026);
nand NAND2 (N12196, N12193, N1388);
xor XOR2 (N12197, N12196, N4115);
not NOT1 (N12198, N12191);
xor XOR2 (N12199, N12192, N8191);
or OR2 (N12200, N12170, N5987);
nand NAND2 (N12201, N12189, N8101);
buf BUF1 (N12202, N12195);
nand NAND3 (N12203, N12175, N7886, N7503);
nor NOR4 (N12204, N12203, N7245, N5864, N9895);
xor XOR2 (N12205, N12197, N10689);
nor NOR3 (N12206, N12198, N2168, N8195);
or OR3 (N12207, N12202, N10925, N415);
not NOT1 (N12208, N12199);
not NOT1 (N12209, N12200);
and AND3 (N12210, N12194, N4228, N5097);
not NOT1 (N12211, N12204);
not NOT1 (N12212, N12181);
not NOT1 (N12213, N12212);
and AND2 (N12214, N12213, N11062);
or OR2 (N12215, N12207, N11857);
nand NAND2 (N12216, N12210, N1283);
nor NOR2 (N12217, N12208, N708);
or OR2 (N12218, N12217, N4795);
nor NOR3 (N12219, N12206, N4993, N3081);
nand NAND3 (N12220, N12219, N9078, N10183);
not NOT1 (N12221, N12209);
not NOT1 (N12222, N12216);
nor NOR2 (N12223, N12211, N6717);
and AND3 (N12224, N12205, N10474, N863);
and AND4 (N12225, N12224, N4319, N8040, N6351);
nand NAND2 (N12226, N12225, N7228);
not NOT1 (N12227, N12183);
nor NOR2 (N12228, N12227, N6229);
or OR2 (N12229, N12220, N1638);
xor XOR2 (N12230, N12215, N11137);
xor XOR2 (N12231, N12226, N12128);
or OR3 (N12232, N12214, N2158, N10718);
xor XOR2 (N12233, N12223, N11248);
xor XOR2 (N12234, N12233, N9221);
or OR4 (N12235, N12232, N1521, N3671, N1837);
buf BUF1 (N12236, N12218);
nor NOR4 (N12237, N12221, N4132, N5198, N9805);
nor NOR2 (N12238, N12231, N6927);
nor NOR2 (N12239, N12201, N4389);
and AND2 (N12240, N12229, N45);
nand NAND2 (N12241, N12239, N11522);
or OR4 (N12242, N12240, N10579, N10474, N1434);
xor XOR2 (N12243, N12235, N9813);
nor NOR2 (N12244, N12234, N11247);
buf BUF1 (N12245, N12241);
nor NOR4 (N12246, N12228, N11621, N8184, N5886);
or OR2 (N12247, N12237, N11768);
buf BUF1 (N12248, N12238);
xor XOR2 (N12249, N12247, N8979);
nor NOR4 (N12250, N12248, N11013, N2966, N11349);
nand NAND2 (N12251, N12246, N6485);
not NOT1 (N12252, N12250);
and AND2 (N12253, N12236, N1605);
not NOT1 (N12254, N12245);
not NOT1 (N12255, N12249);
buf BUF1 (N12256, N12251);
buf BUF1 (N12257, N12222);
nor NOR2 (N12258, N12230, N754);
nor NOR2 (N12259, N12252, N4250);
nor NOR4 (N12260, N12244, N6036, N5077, N6262);
buf BUF1 (N12261, N12242);
nand NAND2 (N12262, N12257, N10254);
nand NAND3 (N12263, N12254, N8919, N9290);
buf BUF1 (N12264, N12256);
not NOT1 (N12265, N12243);
nand NAND4 (N12266, N12264, N10584, N4863, N12211);
and AND4 (N12267, N12261, N9617, N23, N268);
or OR4 (N12268, N12263, N11735, N8441, N149);
and AND2 (N12269, N12259, N7134);
and AND4 (N12270, N12253, N377, N1830, N7825);
not NOT1 (N12271, N12265);
nand NAND4 (N12272, N12262, N7426, N603, N1313);
and AND4 (N12273, N12268, N7895, N1943, N4085);
or OR2 (N12274, N12266, N11116);
or OR3 (N12275, N12270, N6294, N7547);
nand NAND3 (N12276, N12273, N6341, N8492);
nand NAND4 (N12277, N12267, N7243, N1383, N6957);
not NOT1 (N12278, N12274);
or OR2 (N12279, N12272, N11294);
or OR4 (N12280, N12277, N3412, N1437, N4414);
or OR4 (N12281, N12276, N1930, N1614, N5514);
xor XOR2 (N12282, N12255, N11716);
not NOT1 (N12283, N12258);
not NOT1 (N12284, N12281);
nor NOR3 (N12285, N12275, N9553, N9105);
and AND4 (N12286, N12280, N8960, N4320, N2324);
xor XOR2 (N12287, N12286, N1292);
nor NOR4 (N12288, N12271, N4750, N7334, N2487);
not NOT1 (N12289, N12282);
not NOT1 (N12290, N12288);
xor XOR2 (N12291, N12284, N11290);
xor XOR2 (N12292, N12279, N9713);
nand NAND2 (N12293, N12269, N9664);
nand NAND3 (N12294, N12287, N66, N8536);
xor XOR2 (N12295, N12294, N2780);
nor NOR2 (N12296, N12278, N8075);
not NOT1 (N12297, N12260);
buf BUF1 (N12298, N12292);
not NOT1 (N12299, N12297);
nor NOR4 (N12300, N12290, N2547, N12160, N7592);
buf BUF1 (N12301, N12298);
or OR2 (N12302, N12296, N5961);
nor NOR4 (N12303, N12302, N8173, N7956, N466);
not NOT1 (N12304, N12283);
nand NAND3 (N12305, N12304, N5285, N8826);
nand NAND4 (N12306, N12289, N3596, N8380, N7156);
nand NAND2 (N12307, N12291, N9194);
nand NAND3 (N12308, N12299, N219, N4882);
buf BUF1 (N12309, N12306);
or OR4 (N12310, N12285, N1439, N6153, N4584);
nand NAND3 (N12311, N12295, N5334, N9700);
not NOT1 (N12312, N12308);
or OR3 (N12313, N12307, N8167, N10878);
or OR4 (N12314, N12293, N2349, N7417, N8176);
not NOT1 (N12315, N12303);
and AND2 (N12316, N12314, N11224);
buf BUF1 (N12317, N12309);
or OR2 (N12318, N12300, N8824);
nand NAND2 (N12319, N12318, N10133);
nor NOR4 (N12320, N12311, N8084, N2930, N9796);
nand NAND2 (N12321, N12301, N8745);
nor NOR3 (N12322, N12317, N9428, N1744);
xor XOR2 (N12323, N12315, N12078);
xor XOR2 (N12324, N12319, N4899);
nor NOR4 (N12325, N12323, N428, N2528, N2937);
or OR4 (N12326, N12310, N1252, N1278, N9123);
nand NAND3 (N12327, N12312, N5335, N6109);
nor NOR2 (N12328, N12324, N11137);
buf BUF1 (N12329, N12328);
buf BUF1 (N12330, N12313);
xor XOR2 (N12331, N12320, N504);
nor NOR4 (N12332, N12326, N7189, N2760, N618);
and AND3 (N12333, N12322, N2850, N10495);
buf BUF1 (N12334, N12316);
nor NOR2 (N12335, N12329, N4900);
buf BUF1 (N12336, N12331);
xor XOR2 (N12337, N12330, N9982);
buf BUF1 (N12338, N12332);
or OR2 (N12339, N12327, N4135);
buf BUF1 (N12340, N12305);
nand NAND2 (N12341, N12336, N11606);
nor NOR2 (N12342, N12321, N58);
nor NOR2 (N12343, N12339, N8973);
nor NOR3 (N12344, N12338, N11830, N9821);
or OR4 (N12345, N12325, N3061, N5216, N2762);
and AND2 (N12346, N12335, N2363);
nor NOR2 (N12347, N12340, N3759);
or OR3 (N12348, N12337, N2822, N11169);
nand NAND3 (N12349, N12348, N7493, N11144);
xor XOR2 (N12350, N12334, N10374);
xor XOR2 (N12351, N12345, N9911);
buf BUF1 (N12352, N12342);
buf BUF1 (N12353, N12351);
xor XOR2 (N12354, N12333, N12029);
and AND2 (N12355, N12341, N11831);
and AND2 (N12356, N12346, N8558);
nand NAND3 (N12357, N12347, N10555, N265);
xor XOR2 (N12358, N12356, N1608);
and AND4 (N12359, N12349, N9310, N12149, N7322);
nor NOR2 (N12360, N12352, N3344);
buf BUF1 (N12361, N12358);
nor NOR2 (N12362, N12353, N11345);
nand NAND4 (N12363, N12359, N5111, N26, N5408);
or OR4 (N12364, N12361, N2964, N2910, N9678);
or OR3 (N12365, N12360, N5882, N948);
nor NOR4 (N12366, N12344, N5839, N9355, N11353);
and AND4 (N12367, N12363, N1813, N4745, N9097);
or OR4 (N12368, N12355, N7413, N3445, N3959);
nor NOR3 (N12369, N12362, N4039, N7624);
or OR3 (N12370, N12368, N6354, N4523);
xor XOR2 (N12371, N12354, N3429);
xor XOR2 (N12372, N12367, N5553);
or OR3 (N12373, N12357, N5629, N2148);
or OR4 (N12374, N12369, N4008, N10613, N139);
not NOT1 (N12375, N12371);
buf BUF1 (N12376, N12364);
buf BUF1 (N12377, N12372);
or OR4 (N12378, N12343, N6631, N3178, N2859);
nor NOR2 (N12379, N12370, N1113);
nor NOR4 (N12380, N12373, N8399, N6688, N5413);
buf BUF1 (N12381, N12379);
xor XOR2 (N12382, N12378, N6200);
xor XOR2 (N12383, N12382, N7449);
nor NOR4 (N12384, N12366, N3855, N1572, N7756);
or OR2 (N12385, N12380, N9585);
buf BUF1 (N12386, N12374);
or OR3 (N12387, N12350, N2555, N10565);
not NOT1 (N12388, N12386);
or OR2 (N12389, N12377, N7731);
xor XOR2 (N12390, N12376, N1381);
nand NAND4 (N12391, N12388, N11813, N8285, N7066);
nor NOR3 (N12392, N12390, N10388, N4281);
not NOT1 (N12393, N12385);
and AND2 (N12394, N12381, N6291);
not NOT1 (N12395, N12391);
nand NAND3 (N12396, N12387, N4839, N3450);
nand NAND4 (N12397, N12395, N3077, N2700, N12189);
xor XOR2 (N12398, N12393, N1951);
and AND2 (N12399, N12398, N12286);
buf BUF1 (N12400, N12397);
and AND4 (N12401, N12383, N3405, N8591, N1118);
nand NAND3 (N12402, N12365, N3485, N11171);
and AND3 (N12403, N12384, N5698, N6059);
xor XOR2 (N12404, N12394, N8137);
buf BUF1 (N12405, N12392);
or OR4 (N12406, N12403, N11931, N2625, N4662);
nor NOR3 (N12407, N12404, N5378, N4645);
xor XOR2 (N12408, N12405, N789);
nor NOR3 (N12409, N12396, N8257, N2860);
or OR3 (N12410, N12402, N2448, N11690);
and AND3 (N12411, N12400, N3895, N1951);
nand NAND2 (N12412, N12375, N11673);
or OR2 (N12413, N12401, N5499);
or OR3 (N12414, N12413, N10514, N4729);
or OR3 (N12415, N12411, N1313, N3686);
and AND3 (N12416, N12415, N883, N2227);
xor XOR2 (N12417, N12406, N5777);
nor NOR4 (N12418, N12410, N10693, N1107, N10063);
nor NOR3 (N12419, N12389, N2103, N485);
xor XOR2 (N12420, N12408, N4650);
xor XOR2 (N12421, N12399, N8927);
nor NOR3 (N12422, N12407, N105, N12008);
xor XOR2 (N12423, N12409, N5506);
and AND3 (N12424, N12418, N4424, N2841);
or OR4 (N12425, N12421, N1985, N5908, N11665);
not NOT1 (N12426, N12422);
or OR2 (N12427, N12419, N423);
xor XOR2 (N12428, N12427, N102);
xor XOR2 (N12429, N12412, N1707);
nand NAND3 (N12430, N12423, N7496, N1683);
and AND4 (N12431, N12417, N11653, N9042, N8899);
xor XOR2 (N12432, N12416, N8597);
nor NOR2 (N12433, N12414, N12074);
not NOT1 (N12434, N12433);
not NOT1 (N12435, N12428);
not NOT1 (N12436, N12430);
buf BUF1 (N12437, N12436);
not NOT1 (N12438, N12431);
and AND3 (N12439, N12438, N1606, N7962);
not NOT1 (N12440, N12429);
or OR2 (N12441, N12426, N1437);
buf BUF1 (N12442, N12420);
nand NAND2 (N12443, N12441, N12410);
not NOT1 (N12444, N12437);
or OR4 (N12445, N12435, N9614, N1778, N4084);
not NOT1 (N12446, N12443);
xor XOR2 (N12447, N12432, N745);
nor NOR3 (N12448, N12442, N5233, N11824);
not NOT1 (N12449, N12424);
buf BUF1 (N12450, N12440);
or OR2 (N12451, N12444, N8924);
nand NAND3 (N12452, N12445, N3029, N6088);
buf BUF1 (N12453, N12451);
and AND2 (N12454, N12446, N3548);
buf BUF1 (N12455, N12448);
or OR3 (N12456, N12453, N5335, N10059);
nor NOR2 (N12457, N12439, N6122);
xor XOR2 (N12458, N12450, N2567);
nand NAND3 (N12459, N12425, N3074, N6477);
and AND3 (N12460, N12458, N9981, N10141);
nor NOR3 (N12461, N12457, N5319, N7542);
or OR2 (N12462, N12455, N10892);
or OR4 (N12463, N12461, N1035, N8933, N1695);
xor XOR2 (N12464, N12460, N11992);
or OR3 (N12465, N12452, N1857, N6851);
not NOT1 (N12466, N12454);
buf BUF1 (N12467, N12463);
nor NOR4 (N12468, N12466, N10209, N12228, N7233);
xor XOR2 (N12469, N12434, N8589);
nor NOR2 (N12470, N12467, N11731);
not NOT1 (N12471, N12470);
nor NOR3 (N12472, N12468, N10923, N8689);
buf BUF1 (N12473, N12449);
not NOT1 (N12474, N12447);
nor NOR2 (N12475, N12472, N7360);
not NOT1 (N12476, N12462);
nor NOR4 (N12477, N12473, N806, N4670, N3650);
nand NAND2 (N12478, N12476, N5844);
and AND4 (N12479, N12464, N1943, N2142, N179);
not NOT1 (N12480, N12469);
nand NAND4 (N12481, N12474, N6068, N1249, N3685);
or OR4 (N12482, N12456, N3862, N10287, N82);
not NOT1 (N12483, N12481);
nor NOR4 (N12484, N12482, N3376, N8799, N12442);
nor NOR2 (N12485, N12477, N2876);
or OR4 (N12486, N12479, N4499, N2228, N6824);
nor NOR3 (N12487, N12480, N1108, N2522);
nand NAND2 (N12488, N12483, N9866);
not NOT1 (N12489, N12475);
buf BUF1 (N12490, N12484);
and AND2 (N12491, N12488, N6304);
nand NAND4 (N12492, N12491, N9174, N3314, N11214);
nor NOR4 (N12493, N12487, N2868, N5752, N9446);
not NOT1 (N12494, N12492);
nor NOR3 (N12495, N12471, N2341, N3065);
buf BUF1 (N12496, N12459);
xor XOR2 (N12497, N12485, N4501);
nor NOR4 (N12498, N12478, N8529, N12125, N12268);
buf BUF1 (N12499, N12465);
not NOT1 (N12500, N12494);
nor NOR4 (N12501, N12498, N6445, N1396, N9192);
xor XOR2 (N12502, N12489, N8237);
buf BUF1 (N12503, N12497);
or OR2 (N12504, N12499, N4894);
nand NAND2 (N12505, N12504, N9797);
nand NAND2 (N12506, N12501, N4530);
nand NAND2 (N12507, N12486, N8976);
not NOT1 (N12508, N12500);
buf BUF1 (N12509, N12496);
nor NOR4 (N12510, N12495, N11559, N9819, N8893);
buf BUF1 (N12511, N12510);
or OR4 (N12512, N12503, N258, N9895, N3735);
nand NAND4 (N12513, N12502, N3733, N10804, N9159);
or OR4 (N12514, N12505, N6494, N4391, N2300);
nor NOR4 (N12515, N12512, N10256, N11695, N1616);
and AND4 (N12516, N12507, N4695, N5506, N11518);
buf BUF1 (N12517, N12493);
not NOT1 (N12518, N12508);
xor XOR2 (N12519, N12490, N5125);
buf BUF1 (N12520, N12517);
xor XOR2 (N12521, N12515, N1545);
and AND3 (N12522, N12513, N2264, N6930);
nor NOR4 (N12523, N12506, N3217, N2573, N2779);
nor NOR3 (N12524, N12523, N6181, N3640);
and AND4 (N12525, N12511, N4184, N1755, N4210);
xor XOR2 (N12526, N12525, N2173);
buf BUF1 (N12527, N12520);
nor NOR3 (N12528, N12526, N4179, N12334);
or OR3 (N12529, N12522, N11714, N7893);
and AND3 (N12530, N12521, N11211, N7046);
not NOT1 (N12531, N12529);
buf BUF1 (N12532, N12527);
buf BUF1 (N12533, N12524);
not NOT1 (N12534, N12531);
buf BUF1 (N12535, N12534);
and AND4 (N12536, N12516, N8374, N5184, N3290);
nor NOR4 (N12537, N12519, N1729, N9754, N11893);
buf BUF1 (N12538, N12535);
not NOT1 (N12539, N12518);
and AND3 (N12540, N12533, N688, N7461);
and AND3 (N12541, N12514, N4175, N4845);
not NOT1 (N12542, N12532);
not NOT1 (N12543, N12539);
not NOT1 (N12544, N12537);
nor NOR2 (N12545, N12536, N11057);
not NOT1 (N12546, N12541);
nor NOR2 (N12547, N12546, N822);
nand NAND2 (N12548, N12509, N1788);
buf BUF1 (N12549, N12538);
nand NAND3 (N12550, N12543, N2811, N241);
nor NOR2 (N12551, N12549, N6181);
xor XOR2 (N12552, N12530, N8199);
xor XOR2 (N12553, N12550, N9555);
or OR3 (N12554, N12551, N3628, N8542);
xor XOR2 (N12555, N12553, N9794);
buf BUF1 (N12556, N12548);
nand NAND2 (N12557, N12552, N5206);
buf BUF1 (N12558, N12557);
nor NOR2 (N12559, N12540, N9455);
and AND4 (N12560, N12544, N9839, N771, N3081);
buf BUF1 (N12561, N12555);
and AND4 (N12562, N12528, N1800, N2883, N5268);
nand NAND2 (N12563, N12559, N9399);
xor XOR2 (N12564, N12556, N10065);
buf BUF1 (N12565, N12558);
nor NOR3 (N12566, N12560, N8654, N9726);
not NOT1 (N12567, N12547);
nand NAND4 (N12568, N12565, N2199, N8085, N6000);
nor NOR4 (N12569, N12563, N3052, N10865, N3298);
buf BUF1 (N12570, N12554);
buf BUF1 (N12571, N12561);
or OR3 (N12572, N12570, N7125, N4786);
nor NOR4 (N12573, N12569, N4015, N1205, N2115);
nor NOR4 (N12574, N12568, N3772, N10021, N1324);
or OR2 (N12575, N12574, N6731);
and AND4 (N12576, N12562, N10714, N8812, N2253);
not NOT1 (N12577, N12566);
or OR3 (N12578, N12542, N6613, N2312);
not NOT1 (N12579, N12545);
and AND2 (N12580, N12578, N3631);
nand NAND3 (N12581, N12567, N10505, N4776);
nand NAND2 (N12582, N12564, N2409);
nand NAND3 (N12583, N12575, N3017, N8758);
xor XOR2 (N12584, N12576, N4140);
nor NOR4 (N12585, N12577, N4946, N8173, N6022);
or OR3 (N12586, N12580, N11983, N6462);
nand NAND2 (N12587, N12579, N4979);
nor NOR2 (N12588, N12587, N3386);
xor XOR2 (N12589, N12584, N973);
xor XOR2 (N12590, N12582, N12577);
buf BUF1 (N12591, N12586);
nor NOR2 (N12592, N12585, N9727);
nand NAND2 (N12593, N12581, N1589);
nand NAND4 (N12594, N12571, N8223, N9591, N4789);
nor NOR4 (N12595, N12589, N2233, N9839, N613);
and AND2 (N12596, N12572, N8433);
buf BUF1 (N12597, N12591);
nand NAND4 (N12598, N12596, N8023, N5362, N9709);
not NOT1 (N12599, N12593);
or OR4 (N12600, N12597, N1325, N8979, N9645);
buf BUF1 (N12601, N12583);
and AND3 (N12602, N12601, N5082, N6711);
buf BUF1 (N12603, N12598);
nand NAND2 (N12604, N12592, N3616);
not NOT1 (N12605, N12594);
nand NAND4 (N12606, N12599, N1176, N592, N2774);
xor XOR2 (N12607, N12604, N6215);
nand NAND3 (N12608, N12602, N4989, N9834);
or OR2 (N12609, N12573, N1131);
or OR4 (N12610, N12605, N5186, N11205, N5532);
nor NOR3 (N12611, N12610, N4962, N8121);
and AND3 (N12612, N12611, N9490, N9376);
xor XOR2 (N12613, N12590, N9712);
nor NOR2 (N12614, N12612, N4128);
not NOT1 (N12615, N12606);
nand NAND3 (N12616, N12614, N10399, N2690);
nor NOR2 (N12617, N12588, N1436);
and AND2 (N12618, N12615, N7033);
not NOT1 (N12619, N12600);
xor XOR2 (N12620, N12618, N1303);
not NOT1 (N12621, N12619);
or OR2 (N12622, N12608, N7317);
or OR4 (N12623, N12595, N4557, N7211, N11513);
or OR2 (N12624, N12613, N6936);
buf BUF1 (N12625, N12623);
or OR3 (N12626, N12621, N12507, N579);
xor XOR2 (N12627, N12620, N1054);
or OR2 (N12628, N12607, N12287);
not NOT1 (N12629, N12622);
nor NOR4 (N12630, N12624, N170, N10967, N6546);
or OR2 (N12631, N12616, N10168);
buf BUF1 (N12632, N12617);
not NOT1 (N12633, N12628);
not NOT1 (N12634, N12631);
nand NAND3 (N12635, N12629, N3633, N1862);
buf BUF1 (N12636, N12609);
xor XOR2 (N12637, N12626, N12030);
or OR2 (N12638, N12627, N9678);
buf BUF1 (N12639, N12638);
nand NAND4 (N12640, N12630, N10125, N11551, N1091);
nor NOR3 (N12641, N12639, N10743, N87);
xor XOR2 (N12642, N12641, N3568);
not NOT1 (N12643, N12632);
nand NAND3 (N12644, N12625, N8184, N799);
buf BUF1 (N12645, N12603);
buf BUF1 (N12646, N12633);
not NOT1 (N12647, N12634);
not NOT1 (N12648, N12643);
xor XOR2 (N12649, N12647, N11072);
nor NOR4 (N12650, N12636, N6776, N6928, N3472);
not NOT1 (N12651, N12640);
not NOT1 (N12652, N12650);
xor XOR2 (N12653, N12646, N4675);
not NOT1 (N12654, N12644);
buf BUF1 (N12655, N12635);
xor XOR2 (N12656, N12645, N1926);
nor NOR4 (N12657, N12653, N12108, N10739, N6573);
not NOT1 (N12658, N12648);
or OR3 (N12659, N12654, N351, N3543);
and AND4 (N12660, N12649, N11993, N811, N10032);
buf BUF1 (N12661, N12637);
not NOT1 (N12662, N12659);
nand NAND2 (N12663, N12652, N9893);
xor XOR2 (N12664, N12661, N6196);
not NOT1 (N12665, N12658);
nor NOR3 (N12666, N12651, N11031, N4136);
nand NAND2 (N12667, N12642, N12101);
nand NAND4 (N12668, N12667, N528, N2555, N5483);
buf BUF1 (N12669, N12656);
or OR4 (N12670, N12664, N7096, N1963, N2521);
nor NOR4 (N12671, N12655, N10938, N11288, N1177);
not NOT1 (N12672, N12671);
nor NOR3 (N12673, N12666, N8265, N12045);
buf BUF1 (N12674, N12670);
and AND3 (N12675, N12663, N8746, N9008);
buf BUF1 (N12676, N12660);
buf BUF1 (N12677, N12657);
xor XOR2 (N12678, N12673, N3730);
nor NOR2 (N12679, N12675, N3770);
xor XOR2 (N12680, N12669, N7383);
or OR3 (N12681, N12678, N491, N9657);
not NOT1 (N12682, N12676);
or OR3 (N12683, N12680, N4200, N11950);
not NOT1 (N12684, N12662);
buf BUF1 (N12685, N12682);
xor XOR2 (N12686, N12672, N7837);
nand NAND3 (N12687, N12668, N10170, N2871);
buf BUF1 (N12688, N12684);
nand NAND3 (N12689, N12679, N6423, N9802);
or OR3 (N12690, N12689, N5862, N7176);
nor NOR2 (N12691, N12686, N10621);
or OR3 (N12692, N12691, N9393, N10379);
and AND3 (N12693, N12685, N4744, N2614);
and AND2 (N12694, N12692, N117);
or OR4 (N12695, N12688, N5927, N5625, N5793);
or OR2 (N12696, N12677, N801);
nor NOR2 (N12697, N12687, N7305);
and AND4 (N12698, N12674, N2913, N10507, N7293);
buf BUF1 (N12699, N12693);
nor NOR2 (N12700, N12690, N11267);
nor NOR2 (N12701, N12681, N1654);
nor NOR4 (N12702, N12700, N10130, N9344, N4292);
and AND2 (N12703, N12694, N10126);
xor XOR2 (N12704, N12698, N7206);
not NOT1 (N12705, N12701);
and AND2 (N12706, N12703, N7091);
or OR4 (N12707, N12697, N9656, N2124, N1518);
buf BUF1 (N12708, N12704);
buf BUF1 (N12709, N12699);
nand NAND3 (N12710, N12708, N8139, N4988);
buf BUF1 (N12711, N12706);
xor XOR2 (N12712, N12705, N2721);
nand NAND2 (N12713, N12711, N1253);
nor NOR2 (N12714, N12683, N427);
or OR2 (N12715, N12696, N10165);
and AND3 (N12716, N12712, N141, N8584);
and AND4 (N12717, N12713, N5369, N2215, N8180);
and AND4 (N12718, N12714, N8729, N2918, N619);
and AND3 (N12719, N12707, N12173, N12137);
or OR4 (N12720, N12695, N11948, N10294, N497);
xor XOR2 (N12721, N12719, N9834);
and AND2 (N12722, N12717, N10166);
not NOT1 (N12723, N12716);
or OR3 (N12724, N12709, N6837, N6363);
or OR2 (N12725, N12724, N4503);
buf BUF1 (N12726, N12665);
not NOT1 (N12727, N12702);
xor XOR2 (N12728, N12722, N1338);
xor XOR2 (N12729, N12715, N8882);
or OR3 (N12730, N12729, N8468, N12344);
nand NAND3 (N12731, N12723, N11756, N8248);
buf BUF1 (N12732, N12710);
or OR4 (N12733, N12721, N7370, N8849, N6124);
nor NOR2 (N12734, N12733, N9566);
xor XOR2 (N12735, N12718, N10492);
or OR2 (N12736, N12725, N3640);
not NOT1 (N12737, N12735);
nor NOR2 (N12738, N12728, N11021);
nor NOR2 (N12739, N12727, N8511);
not NOT1 (N12740, N12726);
and AND4 (N12741, N12736, N11509, N8349, N11476);
and AND3 (N12742, N12734, N6617, N9131);
nand NAND2 (N12743, N12739, N6728);
xor XOR2 (N12744, N12741, N4845);
not NOT1 (N12745, N12744);
nor NOR2 (N12746, N12731, N4928);
and AND3 (N12747, N12737, N10249, N2662);
nor NOR2 (N12748, N12730, N11592);
buf BUF1 (N12749, N12746);
nor NOR4 (N12750, N12738, N10142, N1993, N9963);
nand NAND4 (N12751, N12720, N1119, N6750, N11407);
nor NOR3 (N12752, N12745, N9474, N7690);
nor NOR2 (N12753, N12752, N1457);
nor NOR2 (N12754, N12750, N8928);
nor NOR4 (N12755, N12748, N11099, N8122, N2395);
or OR3 (N12756, N12751, N10221, N1873);
not NOT1 (N12757, N12743);
or OR2 (N12758, N12756, N6360);
and AND2 (N12759, N12749, N11855);
nand NAND3 (N12760, N12757, N2485, N3580);
or OR3 (N12761, N12742, N3492, N10614);
nand NAND2 (N12762, N12740, N9792);
not NOT1 (N12763, N12762);
not NOT1 (N12764, N12753);
nor NOR2 (N12765, N12761, N7771);
xor XOR2 (N12766, N12754, N12680);
nor NOR3 (N12767, N12765, N2860, N1784);
nor NOR3 (N12768, N12747, N9813, N4692);
nand NAND4 (N12769, N12763, N9441, N4009, N3082);
buf BUF1 (N12770, N12766);
or OR3 (N12771, N12768, N11584, N10977);
nor NOR3 (N12772, N12767, N1774, N1947);
nor NOR4 (N12773, N12759, N9738, N5945, N6528);
nand NAND4 (N12774, N12760, N1653, N8745, N4947);
or OR2 (N12775, N12772, N6534);
nor NOR2 (N12776, N12769, N8922);
and AND3 (N12777, N12764, N1554, N7662);
buf BUF1 (N12778, N12773);
not NOT1 (N12779, N12770);
buf BUF1 (N12780, N12758);
not NOT1 (N12781, N12755);
nand NAND4 (N12782, N12781, N6412, N9984, N9670);
nor NOR4 (N12783, N12779, N8645, N4062, N8655);
or OR3 (N12784, N12732, N7183, N5044);
nor NOR2 (N12785, N12776, N5791);
or OR2 (N12786, N12778, N5539);
or OR2 (N12787, N12785, N3794);
and AND3 (N12788, N12775, N4734, N4719);
xor XOR2 (N12789, N12787, N4618);
not NOT1 (N12790, N12789);
xor XOR2 (N12791, N12788, N328);
nor NOR3 (N12792, N12771, N6220, N7980);
nand NAND2 (N12793, N12780, N11187);
buf BUF1 (N12794, N12790);
nand NAND3 (N12795, N12784, N10853, N2872);
and AND4 (N12796, N12792, N9930, N5052, N3114);
xor XOR2 (N12797, N12795, N9223);
and AND3 (N12798, N12791, N620, N577);
or OR2 (N12799, N12786, N9409);
not NOT1 (N12800, N12798);
nor NOR4 (N12801, N12796, N8279, N168, N1603);
or OR4 (N12802, N12782, N1069, N5462, N4323);
nor NOR3 (N12803, N12794, N9988, N9039);
and AND2 (N12804, N12801, N771);
or OR2 (N12805, N12800, N2454);
or OR3 (N12806, N12793, N6967, N1739);
nor NOR4 (N12807, N12799, N9340, N8917, N9441);
xor XOR2 (N12808, N12806, N7865);
not NOT1 (N12809, N12797);
not NOT1 (N12810, N12808);
not NOT1 (N12811, N12804);
or OR3 (N12812, N12811, N4059, N3450);
or OR2 (N12813, N12809, N4953);
not NOT1 (N12814, N12774);
and AND2 (N12815, N12802, N713);
or OR4 (N12816, N12813, N1531, N12062, N5277);
or OR2 (N12817, N12807, N7469);
buf BUF1 (N12818, N12816);
and AND2 (N12819, N12810, N1592);
not NOT1 (N12820, N12803);
not NOT1 (N12821, N12815);
nand NAND4 (N12822, N12819, N8612, N6476, N11918);
or OR3 (N12823, N12814, N12529, N2099);
nand NAND3 (N12824, N12777, N10946, N12601);
endmodule