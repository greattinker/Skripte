// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16;

output N909,N914,N891,N910,N915,N905,N904,N903,N913,N916;

or OR3 (N17, N3, N3, N12);
and AND2 (N18, N3, N14);
nand NAND2 (N19, N4, N18);
not NOT1 (N20, N9);
or OR2 (N21, N20, N7);
not NOT1 (N22, N17);
nand NAND3 (N23, N22, N3, N3);
buf BUF1 (N24, N21);
buf BUF1 (N25, N22);
xor XOR2 (N26, N17, N13);
not NOT1 (N27, N12);
nor NOR4 (N28, N26, N10, N5, N1);
nor NOR4 (N29, N12, N5, N3, N22);
buf BUF1 (N30, N1);
not NOT1 (N31, N9);
nor NOR2 (N32, N20, N25);
xor XOR2 (N33, N8, N22);
xor XOR2 (N34, N32, N25);
not NOT1 (N35, N28);
nand NAND4 (N36, N23, N2, N28, N17);
xor XOR2 (N37, N24, N28);
nand NAND3 (N38, N30, N37, N5);
or OR3 (N39, N9, N14, N33);
and AND4 (N40, N19, N33, N32, N2);
not NOT1 (N41, N23);
or OR4 (N42, N34, N7, N5, N18);
and AND3 (N43, N42, N15, N14);
not NOT1 (N44, N39);
buf BUF1 (N45, N38);
not NOT1 (N46, N35);
nand NAND4 (N47, N41, N18, N36, N8);
nor NOR4 (N48, N14, N22, N4, N20);
or OR2 (N49, N31, N42);
xor XOR2 (N50, N27, N1);
nor NOR4 (N51, N45, N14, N10, N13);
or OR4 (N52, N51, N37, N43, N19);
or OR3 (N53, N47, N20, N50);
xor XOR2 (N54, N1, N51);
not NOT1 (N55, N25);
or OR2 (N56, N48, N28);
not NOT1 (N57, N55);
xor XOR2 (N58, N46, N52);
or OR4 (N59, N16, N10, N55, N39);
buf BUF1 (N60, N54);
nor NOR4 (N61, N40, N11, N26, N59);
nor NOR3 (N62, N31, N37, N31);
buf BUF1 (N63, N29);
xor XOR2 (N64, N58, N34);
nand NAND3 (N65, N64, N58, N11);
and AND2 (N66, N63, N25);
nand NAND2 (N67, N62, N5);
and AND3 (N68, N56, N15, N48);
or OR3 (N69, N44, N49, N58);
nand NAND3 (N70, N34, N57, N32);
buf BUF1 (N71, N30);
not NOT1 (N72, N53);
not NOT1 (N73, N66);
buf BUF1 (N74, N61);
xor XOR2 (N75, N69, N50);
xor XOR2 (N76, N75, N10);
nand NAND2 (N77, N73, N68);
xor XOR2 (N78, N5, N47);
or OR2 (N79, N70, N2);
and AND4 (N80, N79, N16, N29, N7);
buf BUF1 (N81, N67);
nand NAND3 (N82, N74, N15, N62);
buf BUF1 (N83, N65);
buf BUF1 (N84, N60);
or OR4 (N85, N80, N51, N45, N16);
not NOT1 (N86, N82);
or OR2 (N87, N72, N3);
or OR2 (N88, N83, N27);
and AND3 (N89, N81, N31, N88);
not NOT1 (N90, N64);
or OR4 (N91, N76, N1, N63, N21);
nor NOR4 (N92, N84, N44, N12, N6);
xor XOR2 (N93, N86, N67);
nand NAND2 (N94, N78, N3);
buf BUF1 (N95, N90);
or OR3 (N96, N91, N31, N12);
buf BUF1 (N97, N94);
nor NOR4 (N98, N77, N5, N17, N92);
not NOT1 (N99, N39);
nand NAND4 (N100, N89, N26, N43, N96);
buf BUF1 (N101, N2);
buf BUF1 (N102, N98);
nand NAND3 (N103, N101, N47, N65);
buf BUF1 (N104, N97);
or OR2 (N105, N87, N46);
nand NAND4 (N106, N104, N73, N4, N61);
and AND2 (N107, N93, N81);
nand NAND2 (N108, N100, N25);
nor NOR2 (N109, N107, N27);
not NOT1 (N110, N71);
nor NOR4 (N111, N85, N57, N100, N6);
buf BUF1 (N112, N109);
or OR3 (N113, N108, N13, N47);
buf BUF1 (N114, N105);
not NOT1 (N115, N112);
nor NOR3 (N116, N110, N21, N108);
nand NAND2 (N117, N115, N98);
and AND4 (N118, N113, N44, N16, N10);
and AND4 (N119, N116, N66, N40, N31);
nor NOR4 (N120, N111, N79, N1, N117);
nor NOR4 (N121, N112, N119, N74, N103);
buf BUF1 (N122, N58);
nor NOR4 (N123, N3, N13, N100, N98);
xor XOR2 (N124, N106, N119);
nor NOR3 (N125, N121, N83, N82);
nor NOR2 (N126, N122, N24);
nand NAND4 (N127, N125, N73, N60, N86);
not NOT1 (N128, N102);
and AND2 (N129, N124, N108);
and AND3 (N130, N123, N96, N128);
not NOT1 (N131, N113);
xor XOR2 (N132, N118, N130);
or OR2 (N133, N125, N95);
nor NOR3 (N134, N94, N118, N43);
xor XOR2 (N135, N126, N110);
nand NAND2 (N136, N133, N28);
or OR2 (N137, N99, N64);
nand NAND4 (N138, N114, N115, N99, N100);
nor NOR3 (N139, N132, N94, N69);
or OR2 (N140, N129, N65);
nor NOR3 (N141, N136, N126, N140);
or OR2 (N142, N3, N55);
nor NOR3 (N143, N141, N25, N13);
not NOT1 (N144, N135);
not NOT1 (N145, N120);
nor NOR3 (N146, N131, N126, N119);
nand NAND2 (N147, N138, N126);
buf BUF1 (N148, N143);
nor NOR3 (N149, N146, N10, N45);
nor NOR2 (N150, N148, N101);
and AND4 (N151, N144, N60, N113, N32);
and AND3 (N152, N137, N58, N147);
or OR3 (N153, N140, N33, N44);
nand NAND4 (N154, N145, N86, N26, N28);
not NOT1 (N155, N152);
not NOT1 (N156, N154);
xor XOR2 (N157, N127, N156);
nand NAND4 (N158, N52, N106, N47, N128);
xor XOR2 (N159, N155, N120);
buf BUF1 (N160, N142);
xor XOR2 (N161, N151, N157);
nand NAND2 (N162, N101, N81);
or OR2 (N163, N162, N146);
or OR4 (N164, N160, N7, N142, N127);
nand NAND2 (N165, N159, N134);
nor NOR4 (N166, N33, N95, N53, N160);
nor NOR3 (N167, N165, N68, N22);
xor XOR2 (N168, N167, N18);
nand NAND3 (N169, N163, N49, N100);
nand NAND2 (N170, N153, N62);
nand NAND2 (N171, N169, N16);
buf BUF1 (N172, N166);
not NOT1 (N173, N164);
xor XOR2 (N174, N158, N115);
nor NOR3 (N175, N168, N142, N17);
xor XOR2 (N176, N170, N125);
nand NAND3 (N177, N139, N144, N19);
or OR4 (N178, N174, N151, N105, N140);
buf BUF1 (N179, N178);
nor NOR4 (N180, N176, N73, N29, N36);
xor XOR2 (N181, N173, N122);
buf BUF1 (N182, N175);
nand NAND3 (N183, N181, N171, N147);
and AND4 (N184, N171, N14, N75, N167);
and AND4 (N185, N177, N180, N143, N41);
and AND2 (N186, N63, N110);
nor NOR4 (N187, N149, N182, N25, N108);
nor NOR4 (N188, N135, N128, N77, N4);
or OR3 (N189, N150, N107, N64);
nor NOR2 (N190, N185, N189);
nand NAND3 (N191, N148, N25, N47);
nor NOR4 (N192, N186, N89, N179, N18);
or OR4 (N193, N72, N118, N48, N47);
or OR4 (N194, N191, N35, N36, N156);
nor NOR4 (N195, N190, N18, N19, N134);
or OR4 (N196, N184, N59, N78, N56);
nand NAND2 (N197, N195, N14);
or OR4 (N198, N183, N169, N35, N31);
xor XOR2 (N199, N198, N133);
nand NAND2 (N200, N187, N104);
nand NAND3 (N201, N161, N11, N180);
nand NAND4 (N202, N193, N187, N10, N84);
not NOT1 (N203, N194);
nand NAND2 (N204, N172, N128);
xor XOR2 (N205, N202, N53);
xor XOR2 (N206, N196, N46);
buf BUF1 (N207, N203);
buf BUF1 (N208, N192);
nand NAND3 (N209, N199, N66, N28);
and AND3 (N210, N200, N159, N150);
nand NAND2 (N211, N210, N155);
nor NOR4 (N212, N201, N180, N50, N129);
nor NOR3 (N213, N197, N80, N141);
not NOT1 (N214, N209);
buf BUF1 (N215, N204);
and AND3 (N216, N205, N176, N103);
and AND2 (N217, N216, N175);
or OR4 (N218, N207, N47, N152, N150);
buf BUF1 (N219, N188);
nand NAND2 (N220, N213, N56);
and AND2 (N221, N212, N194);
and AND4 (N222, N215, N79, N180, N215);
buf BUF1 (N223, N218);
not NOT1 (N224, N206);
or OR3 (N225, N221, N203, N218);
buf BUF1 (N226, N217);
xor XOR2 (N227, N226, N177);
nor NOR3 (N228, N224, N60, N57);
nand NAND2 (N229, N227, N58);
nor NOR2 (N230, N229, N161);
and AND4 (N231, N211, N113, N166, N69);
nand NAND4 (N232, N214, N50, N110, N213);
nor NOR3 (N233, N219, N107, N109);
and AND3 (N234, N230, N229, N5);
nand NAND2 (N235, N228, N227);
or OR4 (N236, N220, N194, N108, N131);
xor XOR2 (N237, N208, N40);
nand NAND3 (N238, N235, N200, N143);
xor XOR2 (N239, N236, N236);
buf BUF1 (N240, N225);
or OR4 (N241, N223, N5, N42, N145);
and AND2 (N242, N239, N158);
and AND2 (N243, N222, N88);
buf BUF1 (N244, N243);
and AND2 (N245, N234, N207);
nand NAND2 (N246, N237, N11);
and AND4 (N247, N244, N70, N73, N107);
or OR2 (N248, N240, N3);
or OR4 (N249, N233, N43, N190, N15);
nand NAND3 (N250, N231, N9, N164);
nor NOR3 (N251, N238, N9, N32);
buf BUF1 (N252, N247);
not NOT1 (N253, N241);
nand NAND4 (N254, N253, N107, N20, N19);
nor NOR4 (N255, N242, N142, N230, N197);
nor NOR4 (N256, N232, N29, N72, N178);
not NOT1 (N257, N249);
and AND4 (N258, N246, N229, N26, N93);
or OR2 (N259, N255, N15);
buf BUF1 (N260, N254);
nand NAND3 (N261, N250, N99, N234);
buf BUF1 (N262, N261);
or OR2 (N263, N252, N125);
and AND2 (N264, N257, N78);
nand NAND2 (N265, N248, N104);
and AND2 (N266, N245, N101);
not NOT1 (N267, N260);
or OR4 (N268, N263, N176, N120, N103);
and AND3 (N269, N264, N9, N54);
nor NOR3 (N270, N259, N17, N263);
nor NOR4 (N271, N256, N140, N6, N267);
buf BUF1 (N272, N187);
or OR2 (N273, N266, N88);
or OR2 (N274, N273, N16);
or OR4 (N275, N271, N122, N47, N140);
not NOT1 (N276, N274);
buf BUF1 (N277, N269);
xor XOR2 (N278, N268, N192);
nand NAND2 (N279, N258, N172);
and AND2 (N280, N251, N16);
or OR3 (N281, N262, N136, N66);
and AND2 (N282, N272, N233);
nand NAND2 (N283, N281, N206);
buf BUF1 (N284, N265);
buf BUF1 (N285, N270);
not NOT1 (N286, N275);
xor XOR2 (N287, N276, N74);
or OR4 (N288, N282, N229, N144, N261);
xor XOR2 (N289, N287, N256);
nor NOR2 (N290, N280, N23);
nor NOR2 (N291, N290, N51);
not NOT1 (N292, N279);
not NOT1 (N293, N291);
or OR4 (N294, N283, N142, N223, N131);
not NOT1 (N295, N288);
or OR3 (N296, N292, N179, N285);
not NOT1 (N297, N163);
xor XOR2 (N298, N296, N277);
nand NAND2 (N299, N207, N205);
xor XOR2 (N300, N294, N13);
xor XOR2 (N301, N297, N39);
nor NOR3 (N302, N300, N104, N85);
buf BUF1 (N303, N295);
or OR3 (N304, N302, N228, N85);
nor NOR4 (N305, N289, N5, N160, N224);
or OR4 (N306, N299, N80, N248, N96);
and AND3 (N307, N298, N287, N101);
and AND4 (N308, N307, N90, N109, N100);
not NOT1 (N309, N305);
xor XOR2 (N310, N293, N46);
nor NOR2 (N311, N301, N221);
not NOT1 (N312, N304);
xor XOR2 (N313, N278, N132);
nand NAND4 (N314, N309, N284, N144, N204);
nor NOR3 (N315, N250, N204, N208);
and AND2 (N316, N314, N174);
nand NAND4 (N317, N315, N224, N90, N26);
xor XOR2 (N318, N286, N10);
not NOT1 (N319, N316);
nand NAND2 (N320, N318, N32);
and AND2 (N321, N313, N246);
or OR3 (N322, N312, N207, N215);
nand NAND3 (N323, N311, N289, N282);
not NOT1 (N324, N317);
nand NAND2 (N325, N303, N180);
and AND4 (N326, N321, N303, N6, N135);
not NOT1 (N327, N323);
nand NAND4 (N328, N308, N269, N15, N253);
or OR3 (N329, N320, N147, N27);
buf BUF1 (N330, N306);
nor NOR4 (N331, N310, N87, N216, N162);
nor NOR3 (N332, N327, N35, N192);
and AND2 (N333, N322, N165);
xor XOR2 (N334, N325, N171);
nand NAND3 (N335, N328, N82, N119);
buf BUF1 (N336, N335);
or OR3 (N337, N331, N316, N70);
buf BUF1 (N338, N329);
xor XOR2 (N339, N324, N103);
and AND4 (N340, N336, N291, N282, N45);
nor NOR2 (N341, N319, N127);
nor NOR3 (N342, N337, N182, N292);
buf BUF1 (N343, N338);
xor XOR2 (N344, N334, N116);
or OR4 (N345, N341, N138, N280, N27);
or OR4 (N346, N333, N242, N154, N268);
and AND4 (N347, N343, N26, N135, N197);
or OR3 (N348, N347, N279, N167);
nor NOR2 (N349, N348, N179);
buf BUF1 (N350, N326);
and AND2 (N351, N342, N238);
xor XOR2 (N352, N349, N302);
and AND2 (N353, N340, N89);
and AND3 (N354, N344, N246, N195);
xor XOR2 (N355, N351, N18);
xor XOR2 (N356, N350, N141);
or OR4 (N357, N330, N328, N44, N269);
nand NAND2 (N358, N352, N107);
nand NAND4 (N359, N339, N129, N46, N110);
not NOT1 (N360, N332);
nand NAND2 (N361, N356, N226);
nor NOR4 (N362, N355, N298, N7, N226);
nor NOR4 (N363, N357, N162, N190, N213);
nor NOR4 (N364, N358, N17, N89, N57);
not NOT1 (N365, N345);
or OR4 (N366, N362, N121, N126, N145);
nand NAND2 (N367, N363, N166);
and AND4 (N368, N360, N201, N217, N150);
or OR2 (N369, N367, N87);
not NOT1 (N370, N359);
buf BUF1 (N371, N353);
or OR3 (N372, N361, N211, N87);
not NOT1 (N373, N368);
nand NAND2 (N374, N365, N217);
nor NOR4 (N375, N372, N249, N83, N346);
and AND3 (N376, N233, N37, N59);
or OR4 (N377, N374, N41, N239, N4);
buf BUF1 (N378, N369);
or OR4 (N379, N370, N264, N288, N88);
nor NOR4 (N380, N366, N172, N148, N117);
xor XOR2 (N381, N379, N240);
and AND4 (N382, N376, N261, N279, N87);
nand NAND2 (N383, N371, N192);
nand NAND3 (N384, N354, N217, N372);
or OR2 (N385, N382, N335);
buf BUF1 (N386, N384);
buf BUF1 (N387, N378);
nor NOR2 (N388, N377, N74);
or OR3 (N389, N380, N205, N241);
not NOT1 (N390, N381);
xor XOR2 (N391, N388, N338);
and AND2 (N392, N375, N276);
nor NOR4 (N393, N389, N23, N3, N37);
nand NAND3 (N394, N387, N244, N149);
or OR2 (N395, N386, N135);
or OR3 (N396, N394, N122, N242);
or OR4 (N397, N392, N75, N143, N71);
nand NAND4 (N398, N385, N251, N138, N301);
xor XOR2 (N399, N383, N204);
buf BUF1 (N400, N395);
xor XOR2 (N401, N391, N185);
nand NAND2 (N402, N398, N229);
or OR4 (N403, N402, N63, N43, N339);
buf BUF1 (N404, N399);
and AND2 (N405, N404, N324);
xor XOR2 (N406, N397, N244);
or OR2 (N407, N401, N133);
xor XOR2 (N408, N393, N187);
and AND3 (N409, N407, N397, N204);
xor XOR2 (N410, N405, N50);
nor NOR3 (N411, N403, N324, N270);
nand NAND3 (N412, N400, N113, N333);
nor NOR2 (N413, N390, N367);
buf BUF1 (N414, N409);
not NOT1 (N415, N414);
nand NAND2 (N416, N373, N109);
nand NAND4 (N417, N413, N377, N1, N257);
or OR3 (N418, N364, N370, N128);
or OR3 (N419, N417, N193, N173);
and AND2 (N420, N419, N265);
xor XOR2 (N421, N412, N65);
and AND2 (N422, N411, N8);
xor XOR2 (N423, N410, N382);
xor XOR2 (N424, N396, N390);
and AND2 (N425, N408, N217);
and AND4 (N426, N415, N271, N71, N362);
nor NOR4 (N427, N422, N217, N187, N319);
not NOT1 (N428, N423);
and AND3 (N429, N427, N216, N364);
nand NAND4 (N430, N429, N353, N375, N63);
nand NAND4 (N431, N416, N373, N189, N39);
or OR4 (N432, N431, N400, N399, N212);
buf BUF1 (N433, N426);
buf BUF1 (N434, N428);
nor NOR3 (N435, N432, N370, N231);
and AND2 (N436, N406, N60);
buf BUF1 (N437, N436);
nor NOR2 (N438, N420, N319);
buf BUF1 (N439, N430);
nand NAND3 (N440, N424, N249, N117);
nand NAND2 (N441, N437, N44);
buf BUF1 (N442, N441);
xor XOR2 (N443, N435, N196);
buf BUF1 (N444, N433);
nor NOR4 (N445, N421, N113, N51, N420);
or OR4 (N446, N425, N194, N389, N65);
not NOT1 (N447, N439);
buf BUF1 (N448, N438);
xor XOR2 (N449, N418, N192);
and AND2 (N450, N446, N42);
not NOT1 (N451, N443);
and AND3 (N452, N442, N221, N298);
nand NAND3 (N453, N445, N25, N306);
xor XOR2 (N454, N444, N59);
not NOT1 (N455, N448);
not NOT1 (N456, N453);
and AND3 (N457, N447, N314, N411);
and AND4 (N458, N456, N334, N168, N309);
buf BUF1 (N459, N434);
nand NAND3 (N460, N459, N263, N53);
and AND4 (N461, N450, N234, N174, N339);
not NOT1 (N462, N460);
not NOT1 (N463, N452);
buf BUF1 (N464, N462);
buf BUF1 (N465, N451);
buf BUF1 (N466, N455);
or OR2 (N467, N464, N419);
or OR2 (N468, N465, N100);
xor XOR2 (N469, N461, N175);
not NOT1 (N470, N468);
xor XOR2 (N471, N454, N457);
nor NOR4 (N472, N186, N63, N352, N256);
buf BUF1 (N473, N449);
and AND3 (N474, N466, N229, N285);
buf BUF1 (N475, N470);
not NOT1 (N476, N472);
not NOT1 (N477, N469);
nor NOR2 (N478, N471, N81);
buf BUF1 (N479, N467);
or OR2 (N480, N474, N248);
xor XOR2 (N481, N440, N107);
buf BUF1 (N482, N476);
and AND2 (N483, N475, N29);
nor NOR3 (N484, N480, N177, N278);
nor NOR4 (N485, N484, N406, N268, N27);
xor XOR2 (N486, N481, N89);
not NOT1 (N487, N483);
nor NOR4 (N488, N458, N229, N368, N463);
nand NAND4 (N489, N347, N20, N393, N99);
xor XOR2 (N490, N478, N330);
xor XOR2 (N491, N487, N12);
nand NAND3 (N492, N489, N445, N20);
buf BUF1 (N493, N488);
or OR2 (N494, N492, N52);
and AND2 (N495, N485, N37);
xor XOR2 (N496, N477, N106);
not NOT1 (N497, N482);
buf BUF1 (N498, N490);
nor NOR4 (N499, N495, N146, N439, N1);
xor XOR2 (N500, N479, N146);
nor NOR2 (N501, N497, N219);
nor NOR4 (N502, N473, N240, N103, N423);
nor NOR4 (N503, N493, N314, N151, N15);
xor XOR2 (N504, N491, N334);
not NOT1 (N505, N496);
and AND2 (N506, N503, N13);
buf BUF1 (N507, N504);
and AND3 (N508, N501, N501, N192);
not NOT1 (N509, N507);
and AND3 (N510, N486, N507, N100);
or OR2 (N511, N509, N88);
buf BUF1 (N512, N511);
not NOT1 (N513, N508);
buf BUF1 (N514, N510);
and AND2 (N515, N494, N441);
nand NAND3 (N516, N515, N234, N235);
nor NOR3 (N517, N514, N405, N364);
or OR4 (N518, N506, N466, N294, N77);
not NOT1 (N519, N512);
and AND2 (N520, N505, N512);
nor NOR2 (N521, N518, N438);
and AND2 (N522, N498, N303);
buf BUF1 (N523, N519);
and AND4 (N524, N516, N36, N108, N197);
and AND2 (N525, N499, N309);
and AND3 (N526, N523, N12, N158);
xor XOR2 (N527, N522, N479);
or OR3 (N528, N500, N238, N500);
nor NOR2 (N529, N528, N20);
nand NAND3 (N530, N513, N478, N192);
xor XOR2 (N531, N530, N167);
and AND2 (N532, N520, N6);
buf BUF1 (N533, N502);
xor XOR2 (N534, N532, N469);
or OR3 (N535, N527, N514, N140);
nor NOR4 (N536, N517, N470, N88, N422);
or OR3 (N537, N521, N526, N40);
nor NOR2 (N538, N334, N198);
not NOT1 (N539, N534);
or OR2 (N540, N529, N266);
nor NOR4 (N541, N533, N174, N40, N254);
nand NAND2 (N542, N538, N85);
not NOT1 (N543, N536);
or OR4 (N544, N535, N106, N122, N428);
nor NOR4 (N545, N544, N540, N529, N516);
or OR3 (N546, N326, N174, N405);
nand NAND3 (N547, N524, N109, N419);
nor NOR2 (N548, N539, N38);
and AND4 (N549, N541, N545, N236, N119);
buf BUF1 (N550, N473);
and AND4 (N551, N547, N412, N414, N223);
and AND2 (N552, N550, N225);
and AND4 (N553, N552, N422, N61, N353);
and AND4 (N554, N542, N143, N529, N184);
xor XOR2 (N555, N551, N372);
not NOT1 (N556, N549);
buf BUF1 (N557, N553);
or OR3 (N558, N546, N271, N325);
or OR2 (N559, N525, N130);
buf BUF1 (N560, N531);
not NOT1 (N561, N559);
xor XOR2 (N562, N558, N179);
or OR3 (N563, N562, N52, N428);
nor NOR4 (N564, N537, N64, N266, N265);
nor NOR4 (N565, N557, N18, N158, N33);
nand NAND2 (N566, N561, N307);
or OR3 (N567, N566, N425, N448);
nand NAND2 (N568, N560, N91);
buf BUF1 (N569, N563);
and AND3 (N570, N565, N169, N445);
not NOT1 (N571, N555);
and AND4 (N572, N543, N463, N78, N317);
xor XOR2 (N573, N567, N57);
not NOT1 (N574, N568);
and AND2 (N575, N564, N475);
or OR2 (N576, N572, N497);
or OR4 (N577, N554, N506, N142, N313);
nand NAND3 (N578, N575, N84, N373);
or OR3 (N579, N576, N566, N480);
not NOT1 (N580, N548);
nand NAND2 (N581, N578, N248);
or OR4 (N582, N556, N451, N203, N318);
not NOT1 (N583, N582);
and AND2 (N584, N580, N461);
and AND3 (N585, N584, N241, N578);
not NOT1 (N586, N573);
or OR4 (N587, N574, N515, N34, N444);
nand NAND3 (N588, N577, N433, N188);
nor NOR4 (N589, N570, N578, N11, N369);
nand NAND2 (N590, N587, N161);
or OR4 (N591, N590, N27, N479, N12);
buf BUF1 (N592, N579);
or OR3 (N593, N589, N402, N557);
nor NOR4 (N594, N592, N269, N367, N287);
or OR3 (N595, N583, N130, N28);
and AND4 (N596, N591, N253, N287, N176);
and AND3 (N597, N581, N520, N530);
xor XOR2 (N598, N585, N442);
and AND2 (N599, N596, N38);
not NOT1 (N600, N569);
not NOT1 (N601, N595);
buf BUF1 (N602, N598);
nor NOR4 (N603, N602, N104, N383, N12);
not NOT1 (N604, N601);
and AND4 (N605, N597, N292, N436, N471);
xor XOR2 (N606, N588, N276);
not NOT1 (N607, N594);
xor XOR2 (N608, N586, N22);
and AND3 (N609, N606, N17, N544);
buf BUF1 (N610, N603);
nor NOR4 (N611, N607, N394, N168, N548);
nor NOR4 (N612, N604, N10, N189, N4);
nand NAND3 (N613, N593, N89, N92);
nor NOR3 (N614, N610, N57, N73);
nor NOR2 (N615, N571, N42);
or OR2 (N616, N608, N271);
buf BUF1 (N617, N613);
nor NOR2 (N618, N605, N215);
not NOT1 (N619, N611);
xor XOR2 (N620, N618, N462);
not NOT1 (N621, N617);
or OR4 (N622, N600, N617, N431, N203);
not NOT1 (N623, N599);
buf BUF1 (N624, N614);
and AND2 (N625, N609, N181);
not NOT1 (N626, N625);
nor NOR4 (N627, N612, N314, N400, N575);
and AND3 (N628, N627, N378, N456);
and AND2 (N629, N619, N43);
nor NOR3 (N630, N615, N287, N309);
or OR4 (N631, N630, N302, N396, N572);
not NOT1 (N632, N628);
and AND3 (N633, N621, N630, N453);
nand NAND2 (N634, N624, N606);
and AND4 (N635, N623, N434, N526, N224);
and AND2 (N636, N616, N606);
or OR3 (N637, N629, N228, N72);
not NOT1 (N638, N634);
nor NOR3 (N639, N622, N62, N327);
nor NOR4 (N640, N633, N226, N341, N468);
not NOT1 (N641, N638);
or OR3 (N642, N626, N479, N307);
xor XOR2 (N643, N632, N560);
not NOT1 (N644, N631);
nand NAND3 (N645, N643, N415, N517);
buf BUF1 (N646, N641);
or OR3 (N647, N645, N347, N115);
or OR2 (N648, N637, N500);
buf BUF1 (N649, N620);
and AND4 (N650, N636, N232, N527, N458);
nand NAND2 (N651, N635, N86);
or OR2 (N652, N646, N347);
or OR3 (N653, N648, N479, N505);
not NOT1 (N654, N639);
not NOT1 (N655, N652);
or OR3 (N656, N650, N162, N41);
not NOT1 (N657, N642);
and AND2 (N658, N647, N614);
nor NOR4 (N659, N654, N62, N427, N105);
and AND2 (N660, N653, N46);
not NOT1 (N661, N649);
not NOT1 (N662, N651);
and AND4 (N663, N656, N125, N235, N542);
xor XOR2 (N664, N663, N369);
nand NAND2 (N665, N657, N452);
not NOT1 (N666, N662);
buf BUF1 (N667, N644);
buf BUF1 (N668, N666);
xor XOR2 (N669, N660, N460);
or OR2 (N670, N655, N282);
nand NAND3 (N671, N664, N202, N653);
nand NAND3 (N672, N640, N566, N571);
not NOT1 (N673, N670);
xor XOR2 (N674, N661, N575);
not NOT1 (N675, N665);
nor NOR3 (N676, N673, N148, N501);
and AND2 (N677, N668, N315);
or OR2 (N678, N671, N86);
xor XOR2 (N679, N675, N80);
or OR4 (N680, N679, N10, N474, N101);
or OR4 (N681, N672, N634, N256, N662);
and AND2 (N682, N669, N71);
buf BUF1 (N683, N680);
nand NAND4 (N684, N681, N354, N452, N514);
or OR3 (N685, N682, N483, N226);
buf BUF1 (N686, N658);
buf BUF1 (N687, N674);
nor NOR4 (N688, N687, N297, N424, N81);
buf BUF1 (N689, N659);
and AND4 (N690, N667, N662, N325, N248);
xor XOR2 (N691, N676, N300);
or OR3 (N692, N689, N281, N405);
buf BUF1 (N693, N677);
nand NAND2 (N694, N685, N185);
nand NAND2 (N695, N694, N231);
xor XOR2 (N696, N678, N333);
buf BUF1 (N697, N696);
nor NOR2 (N698, N695, N148);
nor NOR3 (N699, N692, N58, N147);
nor NOR3 (N700, N693, N32, N335);
nand NAND2 (N701, N697, N442);
or OR4 (N702, N700, N700, N579, N333);
or OR2 (N703, N701, N23);
nor NOR4 (N704, N703, N484, N485, N243);
buf BUF1 (N705, N688);
nor NOR3 (N706, N699, N539, N205);
nor NOR3 (N707, N705, N145, N657);
nor NOR4 (N708, N704, N98, N72, N319);
buf BUF1 (N709, N708);
not NOT1 (N710, N706);
nor NOR4 (N711, N710, N619, N119, N85);
or OR2 (N712, N683, N447);
or OR3 (N713, N707, N138, N636);
nor NOR3 (N714, N691, N339, N13);
not NOT1 (N715, N702);
nor NOR2 (N716, N690, N159);
nor NOR2 (N717, N714, N330);
nor NOR2 (N718, N712, N345);
nand NAND2 (N719, N718, N212);
not NOT1 (N720, N719);
nand NAND3 (N721, N717, N641, N480);
nor NOR2 (N722, N713, N710);
and AND4 (N723, N686, N300, N207, N496);
nor NOR2 (N724, N722, N559);
not NOT1 (N725, N720);
not NOT1 (N726, N709);
nor NOR3 (N727, N711, N100, N605);
buf BUF1 (N728, N715);
not NOT1 (N729, N727);
not NOT1 (N730, N725);
or OR4 (N731, N721, N643, N323, N519);
and AND2 (N732, N723, N431);
xor XOR2 (N733, N729, N366);
nand NAND4 (N734, N698, N519, N109, N631);
buf BUF1 (N735, N728);
nand NAND3 (N736, N733, N88, N217);
or OR3 (N737, N726, N477, N494);
not NOT1 (N738, N684);
buf BUF1 (N739, N737);
or OR2 (N740, N730, N65);
not NOT1 (N741, N731);
or OR2 (N742, N734, N12);
buf BUF1 (N743, N741);
or OR4 (N744, N740, N244, N378, N106);
and AND4 (N745, N735, N661, N348, N391);
not NOT1 (N746, N732);
and AND4 (N747, N743, N153, N666, N248);
nor NOR4 (N748, N739, N434, N97, N519);
or OR3 (N749, N748, N378, N41);
nor NOR4 (N750, N744, N590, N508, N572);
xor XOR2 (N751, N738, N280);
and AND2 (N752, N736, N173);
xor XOR2 (N753, N752, N455);
not NOT1 (N754, N745);
nor NOR2 (N755, N749, N210);
not NOT1 (N756, N716);
buf BUF1 (N757, N754);
and AND3 (N758, N755, N645, N378);
not NOT1 (N759, N724);
buf BUF1 (N760, N746);
xor XOR2 (N761, N750, N754);
buf BUF1 (N762, N760);
not NOT1 (N763, N757);
and AND2 (N764, N761, N621);
nor NOR3 (N765, N756, N391, N428);
nand NAND2 (N766, N764, N646);
nand NAND4 (N767, N763, N593, N415, N630);
nor NOR3 (N768, N762, N521, N177);
or OR2 (N769, N753, N445);
nand NAND4 (N770, N747, N728, N304, N374);
nand NAND4 (N771, N768, N393, N501, N194);
not NOT1 (N772, N758);
buf BUF1 (N773, N751);
or OR2 (N774, N765, N592);
buf BUF1 (N775, N771);
and AND3 (N776, N742, N749, N514);
buf BUF1 (N777, N776);
buf BUF1 (N778, N777);
not NOT1 (N779, N767);
nor NOR2 (N780, N759, N260);
or OR4 (N781, N779, N636, N571, N437);
nor NOR2 (N782, N766, N415);
nor NOR3 (N783, N770, N4, N644);
buf BUF1 (N784, N783);
xor XOR2 (N785, N773, N24);
nand NAND4 (N786, N782, N140, N211, N146);
buf BUF1 (N787, N781);
buf BUF1 (N788, N772);
or OR4 (N789, N786, N369, N179, N418);
not NOT1 (N790, N778);
buf BUF1 (N791, N785);
xor XOR2 (N792, N774, N155);
nor NOR4 (N793, N780, N69, N109, N317);
or OR3 (N794, N784, N659, N117);
not NOT1 (N795, N793);
or OR3 (N796, N791, N648, N308);
nor NOR3 (N797, N792, N99, N455);
nand NAND2 (N798, N795, N391);
or OR3 (N799, N789, N175, N381);
buf BUF1 (N800, N799);
nand NAND3 (N801, N788, N196, N50);
nand NAND3 (N802, N801, N787, N729);
buf BUF1 (N803, N742);
nand NAND3 (N804, N769, N8, N60);
nand NAND3 (N805, N798, N155, N640);
and AND3 (N806, N775, N653, N335);
and AND3 (N807, N802, N783, N747);
and AND2 (N808, N807, N754);
and AND3 (N809, N794, N447, N598);
buf BUF1 (N810, N808);
buf BUF1 (N811, N797);
xor XOR2 (N812, N803, N399);
and AND3 (N813, N810, N735, N481);
not NOT1 (N814, N790);
or OR2 (N815, N811, N519);
xor XOR2 (N816, N813, N300);
and AND3 (N817, N809, N366, N157);
nor NOR2 (N818, N816, N123);
and AND2 (N819, N800, N379);
nand NAND3 (N820, N815, N728, N487);
not NOT1 (N821, N805);
nand NAND3 (N822, N819, N329, N210);
buf BUF1 (N823, N806);
xor XOR2 (N824, N796, N535);
and AND2 (N825, N804, N389);
not NOT1 (N826, N817);
not NOT1 (N827, N814);
not NOT1 (N828, N827);
nor NOR4 (N829, N828, N22, N399, N63);
not NOT1 (N830, N824);
not NOT1 (N831, N820);
xor XOR2 (N832, N812, N281);
xor XOR2 (N833, N829, N134);
nor NOR4 (N834, N833, N214, N88, N206);
not NOT1 (N835, N830);
or OR4 (N836, N832, N287, N162, N187);
buf BUF1 (N837, N822);
buf BUF1 (N838, N818);
buf BUF1 (N839, N821);
not NOT1 (N840, N838);
nor NOR4 (N841, N836, N268, N330, N115);
buf BUF1 (N842, N831);
and AND4 (N843, N835, N665, N9, N373);
not NOT1 (N844, N834);
or OR3 (N845, N826, N701, N41);
not NOT1 (N846, N837);
nand NAND4 (N847, N840, N279, N629, N211);
nand NAND2 (N848, N847, N733);
nor NOR2 (N849, N846, N235);
and AND4 (N850, N841, N376, N231, N551);
or OR3 (N851, N845, N642, N291);
or OR3 (N852, N823, N832, N720);
buf BUF1 (N853, N843);
buf BUF1 (N854, N839);
xor XOR2 (N855, N825, N425);
xor XOR2 (N856, N852, N66);
and AND3 (N857, N854, N260, N693);
nand NAND2 (N858, N855, N612);
nor NOR2 (N859, N842, N559);
xor XOR2 (N860, N848, N730);
xor XOR2 (N861, N851, N69);
buf BUF1 (N862, N857);
buf BUF1 (N863, N850);
nand NAND2 (N864, N853, N384);
or OR2 (N865, N858, N34);
xor XOR2 (N866, N864, N411);
nor NOR4 (N867, N862, N137, N782, N318);
and AND2 (N868, N844, N313);
not NOT1 (N869, N868);
buf BUF1 (N870, N866);
or OR4 (N871, N867, N250, N166, N685);
not NOT1 (N872, N863);
nand NAND4 (N873, N861, N262, N467, N227);
nor NOR4 (N874, N849, N350, N211, N218);
buf BUF1 (N875, N865);
buf BUF1 (N876, N874);
nand NAND3 (N877, N873, N468, N161);
nand NAND2 (N878, N860, N871);
buf BUF1 (N879, N791);
or OR2 (N880, N869, N23);
not NOT1 (N881, N878);
and AND4 (N882, N859, N671, N543, N637);
xor XOR2 (N883, N880, N663);
or OR3 (N884, N870, N472, N556);
nand NAND3 (N885, N876, N783, N875);
buf BUF1 (N886, N472);
and AND4 (N887, N856, N187, N428, N664);
buf BUF1 (N888, N884);
not NOT1 (N889, N886);
and AND3 (N890, N872, N386, N837);
nand NAND3 (N891, N885, N19, N231);
buf BUF1 (N892, N890);
nand NAND2 (N893, N888, N834);
buf BUF1 (N894, N893);
not NOT1 (N895, N881);
buf BUF1 (N896, N892);
buf BUF1 (N897, N883);
and AND4 (N898, N897, N784, N565, N587);
or OR3 (N899, N889, N324, N357);
not NOT1 (N900, N894);
xor XOR2 (N901, N898, N788);
or OR3 (N902, N896, N245, N76);
and AND2 (N903, N879, N351);
or OR4 (N904, N882, N622, N272, N36);
not NOT1 (N905, N902);
not NOT1 (N906, N895);
or OR4 (N907, N877, N39, N182, N274);
or OR4 (N908, N906, N799, N828, N594);
xor XOR2 (N909, N901, N544);
not NOT1 (N910, N908);
xor XOR2 (N911, N887, N466);
nand NAND4 (N912, N899, N169, N140, N167);
nor NOR3 (N913, N907, N11, N500);
nor NOR4 (N914, N900, N599, N10, N490);
or OR2 (N915, N912, N399);
or OR4 (N916, N911, N798, N631, N15);
endmodule