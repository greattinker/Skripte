// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17;

output N3006,N3011,N3013,N3000,N3014,N2994,N3001,N3015,N3007,N3017;

not NOT1 (N18, N7);
nand NAND4 (N19, N7, N16, N16, N8);
or OR2 (N20, N11, N15);
buf BUF1 (N21, N18);
and AND2 (N22, N6, N1);
or OR2 (N23, N12, N16);
not NOT1 (N24, N11);
or OR3 (N25, N3, N12, N10);
or OR3 (N26, N19, N22, N3);
or OR3 (N27, N7, N23, N24);
and AND4 (N28, N16, N9, N2, N18);
nor NOR2 (N29, N22, N1);
nand NAND4 (N30, N3, N18, N14, N25);
and AND4 (N31, N10, N3, N18, N30);
buf BUF1 (N32, N11);
or OR4 (N33, N14, N7, N22, N4);
and AND2 (N34, N26, N15);
buf BUF1 (N35, N16);
xor XOR2 (N36, N31, N31);
buf BUF1 (N37, N29);
and AND3 (N38, N28, N12, N29);
nor NOR3 (N39, N37, N9, N21);
nand NAND2 (N40, N28, N17);
or OR3 (N41, N34, N25, N22);
nor NOR3 (N42, N27, N4, N16);
nand NAND3 (N43, N38, N9, N29);
not NOT1 (N44, N36);
and AND2 (N45, N40, N27);
not NOT1 (N46, N43);
nor NOR3 (N47, N45, N44, N38);
not NOT1 (N48, N27);
xor XOR2 (N49, N48, N43);
nor NOR4 (N50, N20, N12, N14, N41);
or OR4 (N51, N35, N13, N30, N44);
and AND3 (N52, N13, N22, N40);
or OR4 (N53, N39, N25, N46, N13);
nor NOR3 (N54, N7, N33, N47);
not NOT1 (N55, N19);
nand NAND3 (N56, N17, N25, N26);
and AND4 (N57, N55, N1, N28, N56);
not NOT1 (N58, N28);
not NOT1 (N59, N42);
and AND2 (N60, N53, N26);
and AND2 (N61, N52, N32);
nor NOR3 (N62, N42, N16, N25);
or OR2 (N63, N62, N13);
not NOT1 (N64, N57);
buf BUF1 (N65, N51);
xor XOR2 (N66, N58, N17);
or OR4 (N67, N50, N25, N21, N55);
nor NOR2 (N68, N59, N39);
buf BUF1 (N69, N64);
nor NOR4 (N70, N66, N26, N53, N36);
xor XOR2 (N71, N68, N52);
xor XOR2 (N72, N54, N7);
xor XOR2 (N73, N63, N44);
nand NAND4 (N74, N72, N67, N55, N37);
buf BUF1 (N75, N28);
nor NOR3 (N76, N73, N41, N17);
nand NAND2 (N77, N75, N42);
not NOT1 (N78, N74);
or OR2 (N79, N77, N25);
nor NOR2 (N80, N69, N42);
buf BUF1 (N81, N71);
and AND3 (N82, N70, N75, N52);
xor XOR2 (N83, N65, N55);
buf BUF1 (N84, N78);
nor NOR3 (N85, N80, N69, N44);
and AND2 (N86, N81, N1);
buf BUF1 (N87, N82);
xor XOR2 (N88, N79, N78);
xor XOR2 (N89, N85, N83);
nand NAND4 (N90, N33, N6, N24, N6);
buf BUF1 (N91, N87);
buf BUF1 (N92, N89);
nor NOR3 (N93, N92, N31, N48);
nor NOR3 (N94, N61, N2, N13);
not NOT1 (N95, N91);
or OR2 (N96, N84, N52);
or OR2 (N97, N49, N23);
xor XOR2 (N98, N60, N4);
and AND2 (N99, N88, N31);
and AND3 (N100, N86, N85, N95);
xor XOR2 (N101, N100, N61);
not NOT1 (N102, N53);
or OR4 (N103, N96, N64, N8, N16);
nor NOR3 (N104, N98, N71, N84);
nor NOR2 (N105, N99, N68);
nand NAND3 (N106, N104, N45, N51);
or OR3 (N107, N101, N16, N48);
nand NAND3 (N108, N105, N89, N78);
or OR2 (N109, N106, N19);
and AND2 (N110, N76, N103);
and AND3 (N111, N45, N36, N31);
and AND2 (N112, N110, N55);
or OR4 (N113, N112, N106, N13, N33);
nor NOR3 (N114, N90, N18, N91);
not NOT1 (N115, N109);
and AND3 (N116, N108, N26, N91);
nand NAND4 (N117, N113, N2, N89, N41);
buf BUF1 (N118, N117);
nand NAND3 (N119, N107, N21, N42);
not NOT1 (N120, N114);
buf BUF1 (N121, N111);
or OR3 (N122, N121, N44, N44);
and AND4 (N123, N94, N91, N53, N39);
nor NOR4 (N124, N122, N24, N80, N18);
xor XOR2 (N125, N124, N41);
or OR4 (N126, N119, N9, N89, N88);
buf BUF1 (N127, N102);
not NOT1 (N128, N97);
xor XOR2 (N129, N125, N62);
not NOT1 (N130, N116);
nand NAND4 (N131, N115, N121, N122, N125);
xor XOR2 (N132, N128, N79);
not NOT1 (N133, N131);
xor XOR2 (N134, N133, N13);
or OR4 (N135, N134, N44, N82, N115);
buf BUF1 (N136, N129);
or OR4 (N137, N130, N67, N55, N103);
and AND2 (N138, N126, N135);
nor NOR2 (N139, N33, N13);
or OR4 (N140, N123, N16, N82, N40);
xor XOR2 (N141, N137, N18);
or OR4 (N142, N127, N27, N83, N105);
or OR3 (N143, N142, N16, N67);
buf BUF1 (N144, N143);
buf BUF1 (N145, N141);
and AND3 (N146, N132, N7, N41);
not NOT1 (N147, N120);
and AND2 (N148, N93, N141);
not NOT1 (N149, N138);
nor NOR2 (N150, N145, N141);
xor XOR2 (N151, N144, N98);
nor NOR2 (N152, N151, N66);
xor XOR2 (N153, N136, N86);
xor XOR2 (N154, N140, N39);
nor NOR2 (N155, N152, N112);
and AND2 (N156, N147, N12);
nor NOR3 (N157, N155, N125, N127);
xor XOR2 (N158, N157, N133);
and AND3 (N159, N154, N146, N157);
nor NOR2 (N160, N59, N73);
xor XOR2 (N161, N159, N59);
nor NOR2 (N162, N149, N152);
or OR3 (N163, N148, N50, N20);
nor NOR2 (N164, N162, N74);
xor XOR2 (N165, N118, N104);
xor XOR2 (N166, N156, N100);
and AND2 (N167, N150, N120);
nand NAND4 (N168, N167, N95, N156, N133);
xor XOR2 (N169, N160, N148);
nor NOR4 (N170, N161, N107, N37, N83);
and AND3 (N171, N170, N168, N46);
nor NOR2 (N172, N21, N1);
buf BUF1 (N173, N166);
and AND2 (N174, N139, N155);
nand NAND4 (N175, N174, N46, N28, N125);
nand NAND3 (N176, N171, N163, N66);
not NOT1 (N177, N113);
not NOT1 (N178, N176);
xor XOR2 (N179, N165, N58);
and AND4 (N180, N164, N141, N12, N110);
buf BUF1 (N181, N175);
xor XOR2 (N182, N179, N138);
and AND2 (N183, N178, N10);
nor NOR4 (N184, N158, N45, N67, N15);
and AND3 (N185, N173, N89, N34);
and AND3 (N186, N153, N107, N98);
nand NAND3 (N187, N184, N144, N78);
and AND2 (N188, N187, N10);
not NOT1 (N189, N181);
not NOT1 (N190, N183);
nor NOR3 (N191, N169, N98, N15);
not NOT1 (N192, N182);
and AND3 (N193, N192, N186, N167);
not NOT1 (N194, N27);
not NOT1 (N195, N194);
buf BUF1 (N196, N189);
or OR2 (N197, N180, N134);
nand NAND2 (N198, N196, N38);
and AND4 (N199, N188, N196, N198, N159);
and AND3 (N200, N157, N144, N53);
nor NOR2 (N201, N199, N142);
xor XOR2 (N202, N177, N133);
or OR4 (N203, N191, N191, N151, N60);
buf BUF1 (N204, N201);
nand NAND2 (N205, N204, N130);
or OR3 (N206, N202, N29, N125);
or OR3 (N207, N197, N82, N135);
not NOT1 (N208, N205);
nand NAND4 (N209, N203, N67, N128, N49);
not NOT1 (N210, N190);
buf BUF1 (N211, N200);
or OR3 (N212, N195, N45, N168);
nor NOR2 (N213, N193, N117);
or OR3 (N214, N206, N195, N39);
and AND4 (N215, N209, N108, N189, N48);
buf BUF1 (N216, N210);
nor NOR3 (N217, N172, N17, N130);
nor NOR4 (N218, N185, N41, N2, N142);
and AND4 (N219, N213, N58, N106, N204);
buf BUF1 (N220, N216);
nor NOR2 (N221, N220, N157);
and AND2 (N222, N212, N210);
nor NOR4 (N223, N217, N126, N90, N146);
and AND4 (N224, N208, N198, N7, N51);
xor XOR2 (N225, N219, N47);
nand NAND2 (N226, N221, N34);
nand NAND3 (N227, N222, N1, N61);
not NOT1 (N228, N224);
not NOT1 (N229, N223);
nor NOR2 (N230, N215, N12);
buf BUF1 (N231, N226);
buf BUF1 (N232, N230);
not NOT1 (N233, N218);
or OR3 (N234, N225, N157, N109);
buf BUF1 (N235, N228);
and AND3 (N236, N229, N6, N164);
not NOT1 (N237, N233);
or OR3 (N238, N234, N48, N187);
or OR4 (N239, N227, N115, N192, N48);
or OR4 (N240, N207, N98, N71, N180);
xor XOR2 (N241, N240, N223);
xor XOR2 (N242, N231, N225);
xor XOR2 (N243, N236, N63);
nand NAND4 (N244, N242, N66, N68, N47);
xor XOR2 (N245, N241, N146);
or OR4 (N246, N237, N72, N95, N173);
nor NOR4 (N247, N232, N78, N58, N227);
buf BUF1 (N248, N243);
and AND4 (N249, N214, N150, N28, N68);
xor XOR2 (N250, N211, N47);
buf BUF1 (N251, N235);
nand NAND2 (N252, N246, N14);
nor NOR4 (N253, N248, N143, N207, N3);
nand NAND4 (N254, N249, N224, N130, N247);
buf BUF1 (N255, N114);
not NOT1 (N256, N245);
nor NOR4 (N257, N256, N141, N211, N98);
nor NOR3 (N258, N252, N35, N224);
and AND3 (N259, N238, N145, N182);
not NOT1 (N260, N259);
nand NAND3 (N261, N258, N144, N234);
or OR2 (N262, N239, N89);
not NOT1 (N263, N254);
or OR2 (N264, N262, N111);
buf BUF1 (N265, N244);
or OR3 (N266, N251, N265, N31);
buf BUF1 (N267, N129);
or OR3 (N268, N264, N188, N141);
xor XOR2 (N269, N253, N120);
buf BUF1 (N270, N263);
or OR2 (N271, N269, N58);
buf BUF1 (N272, N267);
not NOT1 (N273, N255);
nand NAND2 (N274, N271, N228);
buf BUF1 (N275, N250);
not NOT1 (N276, N273);
nand NAND2 (N277, N276, N39);
and AND3 (N278, N260, N270, N7);
and AND2 (N279, N24, N268);
xor XOR2 (N280, N15, N180);
nor NOR4 (N281, N277, N31, N254, N240);
not NOT1 (N282, N261);
or OR2 (N283, N278, N110);
nand NAND3 (N284, N280, N100, N94);
nor NOR3 (N285, N279, N75, N184);
or OR4 (N286, N272, N245, N278, N256);
buf BUF1 (N287, N266);
or OR2 (N288, N274, N226);
not NOT1 (N289, N284);
and AND2 (N290, N257, N49);
not NOT1 (N291, N281);
nor NOR4 (N292, N289, N256, N252, N228);
nor NOR2 (N293, N288, N142);
xor XOR2 (N294, N290, N88);
nand NAND3 (N295, N285, N58, N25);
and AND3 (N296, N295, N168, N24);
or OR4 (N297, N275, N296, N5, N224);
nand NAND2 (N298, N20, N87);
nor NOR3 (N299, N286, N5, N97);
not NOT1 (N300, N299);
and AND2 (N301, N283, N74);
or OR4 (N302, N298, N219, N247, N183);
not NOT1 (N303, N300);
buf BUF1 (N304, N287);
nor NOR4 (N305, N303, N79, N85, N6);
buf BUF1 (N306, N294);
nor NOR3 (N307, N297, N127, N144);
xor XOR2 (N308, N304, N247);
or OR2 (N309, N282, N28);
nand NAND2 (N310, N309, N281);
not NOT1 (N311, N292);
and AND2 (N312, N301, N58);
buf BUF1 (N313, N306);
buf BUF1 (N314, N307);
and AND3 (N315, N311, N40, N310);
nand NAND2 (N316, N124, N238);
not NOT1 (N317, N316);
buf BUF1 (N318, N291);
buf BUF1 (N319, N313);
not NOT1 (N320, N317);
buf BUF1 (N321, N314);
nor NOR4 (N322, N315, N289, N34, N238);
nand NAND2 (N323, N305, N242);
nand NAND4 (N324, N320, N6, N323, N172);
nor NOR3 (N325, N324, N25, N21);
buf BUF1 (N326, N304);
or OR2 (N327, N325, N4);
xor XOR2 (N328, N322, N55);
and AND3 (N329, N321, N41, N206);
buf BUF1 (N330, N329);
not NOT1 (N331, N326);
or OR2 (N332, N319, N141);
or OR2 (N333, N308, N44);
nor NOR3 (N334, N331, N279, N239);
and AND3 (N335, N302, N281, N322);
buf BUF1 (N336, N293);
not NOT1 (N337, N330);
and AND4 (N338, N336, N156, N146, N111);
and AND2 (N339, N328, N259);
buf BUF1 (N340, N337);
buf BUF1 (N341, N339);
xor XOR2 (N342, N338, N205);
or OR2 (N343, N340, N226);
nand NAND3 (N344, N335, N74, N288);
buf BUF1 (N345, N341);
and AND4 (N346, N332, N22, N144, N111);
buf BUF1 (N347, N346);
and AND4 (N348, N312, N14, N85, N195);
buf BUF1 (N349, N348);
buf BUF1 (N350, N327);
xor XOR2 (N351, N333, N215);
nand NAND3 (N352, N342, N226, N130);
not NOT1 (N353, N351);
and AND2 (N354, N318, N274);
nand NAND3 (N355, N345, N96, N249);
not NOT1 (N356, N347);
or OR3 (N357, N354, N343, N112);
buf BUF1 (N358, N319);
nand NAND3 (N359, N357, N198, N347);
buf BUF1 (N360, N356);
nand NAND4 (N361, N352, N299, N116, N73);
nor NOR2 (N362, N353, N163);
buf BUF1 (N363, N355);
buf BUF1 (N364, N361);
and AND4 (N365, N358, N353, N145, N13);
xor XOR2 (N366, N349, N40);
or OR3 (N367, N334, N236, N143);
and AND2 (N368, N362, N92);
not NOT1 (N369, N359);
not NOT1 (N370, N365);
or OR3 (N371, N364, N283, N58);
and AND3 (N372, N360, N265, N319);
xor XOR2 (N373, N344, N211);
or OR3 (N374, N370, N345, N349);
not NOT1 (N375, N368);
or OR3 (N376, N372, N182, N150);
or OR3 (N377, N366, N28, N310);
buf BUF1 (N378, N375);
xor XOR2 (N379, N377, N217);
buf BUF1 (N380, N350);
and AND3 (N381, N376, N224, N216);
xor XOR2 (N382, N380, N100);
buf BUF1 (N383, N379);
not NOT1 (N384, N378);
or OR3 (N385, N381, N279, N241);
and AND2 (N386, N369, N319);
or OR4 (N387, N373, N359, N101, N193);
buf BUF1 (N388, N374);
not NOT1 (N389, N387);
nand NAND3 (N390, N367, N347, N286);
buf BUF1 (N391, N371);
nand NAND2 (N392, N389, N382);
buf BUF1 (N393, N7);
nor NOR2 (N394, N385, N22);
not NOT1 (N395, N383);
nor NOR3 (N396, N390, N214, N187);
nor NOR4 (N397, N393, N232, N240, N324);
and AND2 (N398, N386, N93);
nor NOR2 (N399, N384, N212);
or OR4 (N400, N388, N334, N87, N362);
or OR2 (N401, N398, N89);
not NOT1 (N402, N397);
or OR2 (N403, N363, N207);
and AND2 (N404, N396, N365);
and AND3 (N405, N404, N353, N366);
nand NAND3 (N406, N392, N169, N45);
nor NOR3 (N407, N406, N292, N174);
buf BUF1 (N408, N399);
and AND2 (N409, N400, N392);
xor XOR2 (N410, N409, N259);
not NOT1 (N411, N405);
nor NOR2 (N412, N395, N119);
nand NAND4 (N413, N401, N348, N339, N347);
not NOT1 (N414, N411);
nand NAND4 (N415, N408, N374, N254, N191);
not NOT1 (N416, N402);
nor NOR4 (N417, N407, N203, N228, N298);
buf BUF1 (N418, N415);
buf BUF1 (N419, N413);
nor NOR3 (N420, N416, N386, N247);
or OR2 (N421, N418, N274);
not NOT1 (N422, N419);
and AND2 (N423, N420, N62);
nor NOR2 (N424, N410, N9);
nand NAND4 (N425, N403, N274, N210, N212);
nand NAND2 (N426, N394, N119);
nor NOR4 (N427, N422, N285, N30, N285);
nor NOR2 (N428, N425, N407);
and AND4 (N429, N426, N180, N381, N38);
nor NOR4 (N430, N421, N286, N191, N261);
nor NOR4 (N431, N427, N179, N421, N46);
or OR4 (N432, N423, N352, N394, N228);
or OR4 (N433, N428, N256, N172, N49);
not NOT1 (N434, N433);
and AND2 (N435, N431, N392);
nor NOR2 (N436, N424, N400);
nand NAND2 (N437, N412, N74);
or OR2 (N438, N417, N143);
or OR3 (N439, N437, N187, N340);
nor NOR3 (N440, N439, N369, N173);
nor NOR4 (N441, N429, N333, N225, N434);
and AND2 (N442, N113, N16);
xor XOR2 (N443, N442, N302);
xor XOR2 (N444, N391, N60);
or OR4 (N445, N443, N289, N201, N47);
buf BUF1 (N446, N432);
or OR4 (N447, N446, N16, N167, N170);
buf BUF1 (N448, N447);
not NOT1 (N449, N444);
xor XOR2 (N450, N436, N290);
not NOT1 (N451, N435);
and AND4 (N452, N438, N170, N274, N187);
buf BUF1 (N453, N440);
or OR4 (N454, N448, N321, N333, N122);
and AND3 (N455, N450, N96, N421);
not NOT1 (N456, N454);
or OR3 (N457, N455, N81, N353);
not NOT1 (N458, N449);
not NOT1 (N459, N451);
xor XOR2 (N460, N414, N334);
or OR2 (N461, N457, N289);
buf BUF1 (N462, N460);
or OR2 (N463, N453, N346);
buf BUF1 (N464, N462);
nand NAND4 (N465, N456, N404, N27, N190);
buf BUF1 (N466, N463);
or OR4 (N467, N466, N190, N336, N428);
xor XOR2 (N468, N458, N409);
and AND4 (N469, N465, N311, N190, N125);
and AND2 (N470, N464, N243);
and AND2 (N471, N441, N341);
xor XOR2 (N472, N461, N299);
not NOT1 (N473, N467);
buf BUF1 (N474, N473);
and AND2 (N475, N474, N358);
nor NOR3 (N476, N452, N202, N180);
buf BUF1 (N477, N471);
xor XOR2 (N478, N445, N359);
nand NAND4 (N479, N478, N289, N388, N213);
and AND3 (N480, N469, N48, N171);
nor NOR2 (N481, N480, N71);
buf BUF1 (N482, N459);
nor NOR2 (N483, N476, N321);
nor NOR4 (N484, N482, N27, N470, N111);
or OR4 (N485, N352, N276, N72, N21);
or OR4 (N486, N477, N91, N120, N28);
not NOT1 (N487, N430);
and AND4 (N488, N479, N29, N263, N1);
xor XOR2 (N489, N484, N388);
and AND3 (N490, N485, N238, N84);
or OR3 (N491, N468, N349, N29);
and AND2 (N492, N483, N404);
not NOT1 (N493, N490);
nand NAND4 (N494, N488, N274, N470, N199);
not NOT1 (N495, N494);
nand NAND2 (N496, N472, N226);
buf BUF1 (N497, N489);
and AND2 (N498, N481, N289);
or OR2 (N499, N475, N283);
or OR3 (N500, N491, N386, N372);
nor NOR4 (N501, N495, N17, N368, N371);
and AND4 (N502, N500, N77, N173, N66);
and AND2 (N503, N492, N106);
and AND2 (N504, N499, N433);
nor NOR2 (N505, N496, N484);
xor XOR2 (N506, N493, N1);
xor XOR2 (N507, N486, N240);
xor XOR2 (N508, N503, N226);
or OR2 (N509, N505, N231);
and AND3 (N510, N507, N286, N280);
nand NAND4 (N511, N502, N408, N358, N204);
nor NOR4 (N512, N509, N111, N430, N191);
not NOT1 (N513, N510);
nor NOR3 (N514, N508, N505, N68);
not NOT1 (N515, N514);
nand NAND4 (N516, N501, N198, N438, N162);
nand NAND2 (N517, N506, N151);
buf BUF1 (N518, N511);
or OR2 (N519, N487, N155);
and AND2 (N520, N515, N56);
buf BUF1 (N521, N497);
nand NAND2 (N522, N513, N125);
or OR3 (N523, N517, N132, N150);
buf BUF1 (N524, N512);
nand NAND2 (N525, N522, N264);
and AND2 (N526, N498, N259);
or OR2 (N527, N504, N45);
nor NOR4 (N528, N520, N387, N264, N86);
xor XOR2 (N529, N516, N34);
not NOT1 (N530, N528);
xor XOR2 (N531, N530, N231);
not NOT1 (N532, N526);
and AND2 (N533, N519, N491);
not NOT1 (N534, N532);
and AND3 (N535, N518, N54, N79);
buf BUF1 (N536, N525);
buf BUF1 (N537, N523);
nand NAND4 (N538, N536, N416, N195, N64);
not NOT1 (N539, N535);
nand NAND2 (N540, N527, N123);
and AND4 (N541, N534, N257, N226, N484);
xor XOR2 (N542, N529, N367);
xor XOR2 (N543, N541, N354);
and AND2 (N544, N540, N139);
nand NAND3 (N545, N539, N137, N3);
xor XOR2 (N546, N543, N299);
xor XOR2 (N547, N542, N546);
buf BUF1 (N548, N427);
and AND2 (N549, N547, N433);
buf BUF1 (N550, N537);
not NOT1 (N551, N545);
not NOT1 (N552, N533);
not NOT1 (N553, N549);
or OR4 (N554, N553, N206, N144, N53);
nand NAND4 (N555, N548, N237, N257, N440);
nor NOR2 (N556, N521, N97);
or OR3 (N557, N538, N487, N452);
or OR4 (N558, N550, N432, N375, N360);
nand NAND2 (N559, N558, N83);
or OR3 (N560, N556, N298, N446);
or OR3 (N561, N557, N40, N289);
and AND2 (N562, N555, N398);
buf BUF1 (N563, N544);
or OR2 (N564, N551, N245);
and AND3 (N565, N559, N214, N76);
nor NOR4 (N566, N563, N552, N57, N465);
nand NAND4 (N567, N507, N30, N278, N449);
and AND3 (N568, N524, N243, N175);
nand NAND4 (N569, N560, N514, N397, N31);
and AND3 (N570, N569, N312, N459);
nand NAND2 (N571, N570, N429);
not NOT1 (N572, N571);
nand NAND3 (N573, N565, N148, N351);
xor XOR2 (N574, N567, N127);
xor XOR2 (N575, N554, N287);
not NOT1 (N576, N564);
nor NOR3 (N577, N561, N467, N84);
nor NOR4 (N578, N572, N543, N41, N39);
nand NAND3 (N579, N531, N143, N49);
buf BUF1 (N580, N576);
buf BUF1 (N581, N573);
or OR3 (N582, N579, N310, N309);
not NOT1 (N583, N581);
buf BUF1 (N584, N580);
or OR2 (N585, N578, N488);
nor NOR2 (N586, N583, N418);
not NOT1 (N587, N568);
not NOT1 (N588, N587);
nor NOR3 (N589, N566, N84, N208);
xor XOR2 (N590, N588, N580);
or OR3 (N591, N582, N443, N140);
or OR4 (N592, N586, N347, N484, N192);
or OR4 (N593, N590, N293, N97, N293);
buf BUF1 (N594, N577);
xor XOR2 (N595, N594, N465);
xor XOR2 (N596, N593, N464);
or OR3 (N597, N589, N580, N8);
or OR2 (N598, N575, N54);
not NOT1 (N599, N595);
nor NOR2 (N600, N574, N361);
nand NAND3 (N601, N591, N492, N434);
nand NAND3 (N602, N562, N532, N520);
buf BUF1 (N603, N601);
nor NOR3 (N604, N585, N308, N76);
nor NOR4 (N605, N584, N71, N498, N476);
nor NOR2 (N606, N599, N439);
nor NOR4 (N607, N598, N60, N383, N172);
or OR2 (N608, N605, N573);
nor NOR3 (N609, N603, N235, N226);
not NOT1 (N610, N604);
not NOT1 (N611, N600);
nand NAND2 (N612, N611, N323);
not NOT1 (N613, N592);
nor NOR4 (N614, N606, N61, N183, N591);
xor XOR2 (N615, N612, N365);
nand NAND3 (N616, N610, N282, N575);
nor NOR3 (N617, N609, N582, N227);
not NOT1 (N618, N607);
or OR3 (N619, N616, N355, N359);
nor NOR2 (N620, N596, N255);
or OR2 (N621, N597, N30);
nor NOR3 (N622, N618, N26, N477);
and AND3 (N623, N613, N406, N391);
buf BUF1 (N624, N620);
xor XOR2 (N625, N619, N11);
not NOT1 (N626, N625);
and AND3 (N627, N626, N307, N45);
xor XOR2 (N628, N615, N321);
nand NAND3 (N629, N602, N498, N259);
xor XOR2 (N630, N629, N193);
or OR3 (N631, N608, N397, N63);
or OR4 (N632, N614, N247, N595, N300);
nand NAND2 (N633, N617, N111);
xor XOR2 (N634, N621, N279);
buf BUF1 (N635, N633);
nand NAND2 (N636, N623, N177);
nand NAND4 (N637, N632, N501, N325, N399);
or OR3 (N638, N628, N247, N193);
xor XOR2 (N639, N634, N74);
or OR2 (N640, N639, N47);
nor NOR2 (N641, N637, N379);
nand NAND3 (N642, N636, N380, N38);
or OR3 (N643, N630, N543, N609);
nor NOR4 (N644, N643, N409, N290, N403);
xor XOR2 (N645, N622, N37);
nor NOR3 (N646, N641, N43, N443);
and AND3 (N647, N645, N587, N590);
or OR2 (N648, N627, N509);
or OR2 (N649, N631, N577);
xor XOR2 (N650, N640, N33);
nand NAND2 (N651, N646, N437);
nand NAND3 (N652, N635, N485, N30);
not NOT1 (N653, N650);
or OR4 (N654, N642, N26, N90, N632);
nand NAND3 (N655, N638, N276, N304);
not NOT1 (N656, N652);
xor XOR2 (N657, N649, N313);
not NOT1 (N658, N656);
not NOT1 (N659, N655);
buf BUF1 (N660, N657);
nand NAND2 (N661, N648, N310);
buf BUF1 (N662, N624);
and AND4 (N663, N654, N227, N288, N68);
not NOT1 (N664, N651);
nor NOR3 (N665, N653, N400, N237);
nand NAND4 (N666, N663, N327, N1, N115);
nand NAND3 (N667, N662, N33, N497);
and AND3 (N668, N658, N74, N159);
nor NOR2 (N669, N664, N541);
or OR2 (N670, N660, N122);
nand NAND4 (N671, N670, N461, N513, N388);
nor NOR3 (N672, N666, N527, N380);
and AND3 (N673, N661, N279, N231);
nor NOR2 (N674, N665, N85);
or OR2 (N675, N668, N350);
xor XOR2 (N676, N674, N625);
nand NAND3 (N677, N671, N631, N290);
and AND4 (N678, N676, N355, N241, N320);
xor XOR2 (N679, N678, N316);
and AND2 (N680, N669, N557);
not NOT1 (N681, N677);
and AND4 (N682, N644, N476, N493, N419);
nor NOR4 (N683, N647, N253, N336, N551);
buf BUF1 (N684, N681);
or OR2 (N685, N673, N292);
or OR4 (N686, N675, N102, N336, N535);
xor XOR2 (N687, N686, N132);
nand NAND3 (N688, N685, N629, N666);
not NOT1 (N689, N679);
buf BUF1 (N690, N667);
or OR2 (N691, N689, N14);
nand NAND2 (N692, N659, N581);
xor XOR2 (N693, N683, N124);
not NOT1 (N694, N672);
nand NAND3 (N695, N690, N626, N385);
xor XOR2 (N696, N694, N333);
buf BUF1 (N697, N680);
xor XOR2 (N698, N697, N324);
buf BUF1 (N699, N696);
xor XOR2 (N700, N691, N692);
buf BUF1 (N701, N239);
buf BUF1 (N702, N688);
buf BUF1 (N703, N701);
nand NAND3 (N704, N698, N562, N694);
or OR2 (N705, N702, N281);
xor XOR2 (N706, N695, N246);
and AND3 (N707, N703, N136, N397);
not NOT1 (N708, N682);
not NOT1 (N709, N707);
buf BUF1 (N710, N708);
or OR4 (N711, N704, N519, N330, N380);
or OR2 (N712, N710, N91);
nor NOR4 (N713, N711, N460, N273, N287);
buf BUF1 (N714, N699);
and AND3 (N715, N684, N556, N206);
xor XOR2 (N716, N687, N137);
not NOT1 (N717, N712);
nor NOR4 (N718, N714, N171, N250, N538);
buf BUF1 (N719, N693);
nand NAND3 (N720, N717, N122, N236);
and AND2 (N721, N700, N476);
xor XOR2 (N722, N713, N567);
nor NOR4 (N723, N705, N497, N358, N30);
not NOT1 (N724, N721);
nand NAND3 (N725, N719, N359, N113);
xor XOR2 (N726, N723, N183);
nand NAND3 (N727, N725, N259, N574);
and AND3 (N728, N727, N277, N255);
not NOT1 (N729, N722);
or OR4 (N730, N715, N654, N637, N391);
buf BUF1 (N731, N720);
or OR2 (N732, N728, N266);
xor XOR2 (N733, N706, N185);
nor NOR2 (N734, N718, N467);
not NOT1 (N735, N726);
or OR4 (N736, N732, N678, N647, N364);
and AND4 (N737, N724, N80, N10, N294);
nand NAND4 (N738, N736, N267, N158, N664);
and AND4 (N739, N738, N528, N415, N22);
and AND4 (N740, N735, N609, N416, N466);
nor NOR3 (N741, N740, N266, N527);
xor XOR2 (N742, N741, N123);
nand NAND2 (N743, N709, N246);
and AND2 (N744, N729, N723);
buf BUF1 (N745, N744);
xor XOR2 (N746, N716, N329);
not NOT1 (N747, N730);
xor XOR2 (N748, N742, N466);
nand NAND4 (N749, N731, N676, N301, N7);
nor NOR2 (N750, N745, N434);
nand NAND3 (N751, N743, N277, N203);
or OR3 (N752, N747, N724, N46);
nor NOR4 (N753, N737, N393, N99, N676);
not NOT1 (N754, N739);
and AND4 (N755, N746, N518, N529, N319);
nand NAND3 (N756, N753, N515, N467);
nor NOR2 (N757, N733, N286);
or OR3 (N758, N734, N271, N311);
or OR3 (N759, N750, N71, N151);
not NOT1 (N760, N758);
buf BUF1 (N761, N751);
nor NOR4 (N762, N761, N521, N435, N6);
xor XOR2 (N763, N760, N487);
and AND4 (N764, N754, N519, N596, N497);
nand NAND3 (N765, N763, N680, N601);
nand NAND2 (N766, N757, N654);
or OR2 (N767, N766, N410);
buf BUF1 (N768, N752);
xor XOR2 (N769, N765, N247);
nor NOR4 (N770, N762, N271, N169, N65);
or OR2 (N771, N756, N701);
nand NAND3 (N772, N767, N708, N748);
or OR2 (N773, N403, N165);
not NOT1 (N774, N769);
xor XOR2 (N775, N773, N465);
or OR4 (N776, N772, N104, N441, N304);
buf BUF1 (N777, N755);
or OR4 (N778, N764, N680, N764, N517);
nand NAND2 (N779, N771, N221);
and AND4 (N780, N768, N660, N7, N456);
not NOT1 (N781, N778);
xor XOR2 (N782, N775, N6);
and AND3 (N783, N782, N460, N196);
not NOT1 (N784, N776);
or OR4 (N785, N780, N360, N765, N108);
not NOT1 (N786, N783);
or OR3 (N787, N785, N138, N478);
and AND3 (N788, N770, N682, N325);
nand NAND3 (N789, N787, N273, N488);
or OR2 (N790, N779, N317);
nand NAND2 (N791, N774, N297);
not NOT1 (N792, N789);
nor NOR3 (N793, N759, N632, N402);
not NOT1 (N794, N786);
buf BUF1 (N795, N777);
nor NOR2 (N796, N794, N477);
and AND4 (N797, N795, N265, N600, N271);
not NOT1 (N798, N796);
nor NOR2 (N799, N793, N520);
and AND3 (N800, N797, N427, N348);
nand NAND3 (N801, N799, N211, N586);
nand NAND4 (N802, N791, N396, N795, N693);
nand NAND4 (N803, N801, N781, N716, N522);
or OR2 (N804, N131, N497);
or OR4 (N805, N784, N799, N174, N545);
nor NOR2 (N806, N800, N79);
or OR2 (N807, N802, N753);
and AND2 (N808, N805, N803);
nand NAND2 (N809, N361, N472);
or OR3 (N810, N804, N631, N636);
nand NAND4 (N811, N807, N676, N242, N667);
xor XOR2 (N812, N788, N315);
nor NOR2 (N813, N809, N34);
buf BUF1 (N814, N806);
nand NAND4 (N815, N808, N92, N254, N11);
not NOT1 (N816, N815);
nor NOR4 (N817, N812, N737, N79, N257);
nor NOR4 (N818, N811, N320, N753, N357);
nor NOR3 (N819, N798, N657, N812);
buf BUF1 (N820, N810);
nand NAND2 (N821, N790, N676);
buf BUF1 (N822, N817);
nand NAND4 (N823, N813, N231, N559, N345);
and AND2 (N824, N818, N794);
buf BUF1 (N825, N822);
and AND4 (N826, N820, N439, N132, N615);
nand NAND2 (N827, N816, N562);
and AND4 (N828, N821, N190, N115, N172);
xor XOR2 (N829, N828, N82);
nand NAND4 (N830, N814, N747, N347, N259);
not NOT1 (N831, N825);
nand NAND3 (N832, N792, N464, N217);
nor NOR2 (N833, N819, N147);
and AND4 (N834, N833, N210, N12, N265);
buf BUF1 (N835, N831);
buf BUF1 (N836, N826);
nand NAND4 (N837, N824, N765, N823, N758);
and AND2 (N838, N827, N482);
or OR3 (N839, N656, N42, N547);
buf BUF1 (N840, N836);
and AND3 (N841, N749, N679, N321);
and AND3 (N842, N840, N306, N255);
xor XOR2 (N843, N841, N150);
and AND2 (N844, N834, N341);
not NOT1 (N845, N837);
xor XOR2 (N846, N839, N59);
and AND2 (N847, N844, N265);
not NOT1 (N848, N846);
nand NAND4 (N849, N843, N508, N22, N483);
buf BUF1 (N850, N842);
xor XOR2 (N851, N850, N821);
or OR3 (N852, N829, N492, N753);
or OR3 (N853, N845, N826, N587);
or OR3 (N854, N832, N807, N181);
nor NOR3 (N855, N851, N143, N549);
xor XOR2 (N856, N849, N227);
and AND2 (N857, N838, N322);
buf BUF1 (N858, N855);
nand NAND4 (N859, N835, N432, N811, N432);
nor NOR2 (N860, N859, N402);
nand NAND3 (N861, N856, N335, N280);
buf BUF1 (N862, N853);
nand NAND4 (N863, N848, N103, N630, N5);
nor NOR4 (N864, N858, N37, N719, N854);
buf BUF1 (N865, N563);
nor NOR4 (N866, N861, N488, N77, N226);
nand NAND3 (N867, N857, N464, N36);
xor XOR2 (N868, N867, N185);
nor NOR4 (N869, N864, N347, N269, N352);
or OR2 (N870, N868, N788);
or OR3 (N871, N860, N599, N523);
and AND4 (N872, N847, N322, N723, N847);
or OR2 (N873, N872, N421);
or OR3 (N874, N852, N329, N429);
nand NAND4 (N875, N862, N442, N452, N410);
not NOT1 (N876, N875);
nor NOR2 (N877, N874, N207);
and AND4 (N878, N869, N795, N67, N582);
and AND3 (N879, N877, N323, N858);
buf BUF1 (N880, N866);
xor XOR2 (N881, N865, N263);
nand NAND3 (N882, N870, N305, N264);
nand NAND3 (N883, N863, N799, N313);
buf BUF1 (N884, N882);
xor XOR2 (N885, N871, N191);
not NOT1 (N886, N883);
not NOT1 (N887, N885);
and AND3 (N888, N878, N292, N594);
or OR4 (N889, N873, N636, N386, N43);
and AND4 (N890, N886, N140, N452, N450);
and AND4 (N891, N890, N232, N105, N588);
and AND4 (N892, N889, N164, N743, N343);
not NOT1 (N893, N888);
or OR2 (N894, N887, N838);
or OR4 (N895, N891, N854, N855, N112);
buf BUF1 (N896, N881);
nand NAND3 (N897, N879, N889, N58);
or OR3 (N898, N892, N536, N310);
not NOT1 (N899, N894);
xor XOR2 (N900, N897, N58);
nor NOR3 (N901, N898, N404, N750);
and AND2 (N902, N830, N5);
nor NOR2 (N903, N895, N647);
not NOT1 (N904, N899);
nand NAND4 (N905, N884, N195, N779, N205);
not NOT1 (N906, N896);
nand NAND2 (N907, N904, N158);
xor XOR2 (N908, N893, N837);
not NOT1 (N909, N905);
buf BUF1 (N910, N907);
nand NAND3 (N911, N880, N212, N20);
xor XOR2 (N912, N902, N493);
not NOT1 (N913, N876);
or OR2 (N914, N901, N53);
and AND2 (N915, N913, N554);
not NOT1 (N916, N915);
nand NAND2 (N917, N914, N320);
buf BUF1 (N918, N917);
or OR2 (N919, N909, N455);
xor XOR2 (N920, N919, N506);
xor XOR2 (N921, N920, N777);
nand NAND2 (N922, N906, N274);
nor NOR2 (N923, N918, N45);
nor NOR3 (N924, N923, N578, N744);
or OR2 (N925, N910, N421);
or OR4 (N926, N924, N350, N623, N72);
nor NOR2 (N927, N925, N268);
not NOT1 (N928, N926);
xor XOR2 (N929, N903, N256);
or OR4 (N930, N916, N402, N566, N258);
nand NAND2 (N931, N900, N360);
not NOT1 (N932, N911);
buf BUF1 (N933, N927);
or OR4 (N934, N930, N548, N616, N562);
not NOT1 (N935, N921);
nand NAND3 (N936, N933, N828, N168);
and AND4 (N937, N908, N769, N709, N663);
or OR4 (N938, N935, N223, N937, N824);
not NOT1 (N939, N415);
or OR3 (N940, N922, N95, N137);
or OR2 (N941, N938, N7);
nand NAND4 (N942, N912, N576, N755, N606);
nor NOR4 (N943, N934, N671, N378, N757);
buf BUF1 (N944, N928);
nand NAND2 (N945, N941, N100);
or OR3 (N946, N931, N329, N685);
buf BUF1 (N947, N929);
buf BUF1 (N948, N946);
nand NAND3 (N949, N945, N140, N391);
nand NAND3 (N950, N948, N284, N933);
not NOT1 (N951, N944);
or OR3 (N952, N950, N772, N142);
xor XOR2 (N953, N939, N496);
not NOT1 (N954, N947);
xor XOR2 (N955, N954, N249);
and AND3 (N956, N953, N723, N505);
xor XOR2 (N957, N955, N457);
buf BUF1 (N958, N936);
xor XOR2 (N959, N951, N171);
or OR4 (N960, N942, N826, N457, N124);
nand NAND2 (N961, N952, N761);
xor XOR2 (N962, N960, N149);
nand NAND4 (N963, N959, N312, N452, N854);
and AND3 (N964, N961, N926, N260);
xor XOR2 (N965, N940, N632);
nand NAND4 (N966, N949, N374, N613, N14);
and AND2 (N967, N966, N854);
nand NAND4 (N968, N967, N265, N541, N22);
xor XOR2 (N969, N956, N774);
buf BUF1 (N970, N965);
nor NOR3 (N971, N962, N785, N16);
not NOT1 (N972, N957);
nor NOR4 (N973, N932, N683, N380, N410);
buf BUF1 (N974, N958);
buf BUF1 (N975, N943);
nor NOR2 (N976, N972, N142);
not NOT1 (N977, N975);
buf BUF1 (N978, N970);
xor XOR2 (N979, N974, N880);
not NOT1 (N980, N978);
and AND2 (N981, N964, N15);
or OR4 (N982, N968, N388, N139, N396);
nand NAND4 (N983, N979, N757, N592, N274);
nor NOR3 (N984, N980, N838, N662);
nor NOR3 (N985, N984, N851, N687);
buf BUF1 (N986, N973);
and AND3 (N987, N969, N166, N518);
buf BUF1 (N988, N971);
nand NAND4 (N989, N986, N672, N264, N402);
and AND4 (N990, N988, N129, N537, N491);
not NOT1 (N991, N985);
nor NOR4 (N992, N976, N652, N601, N430);
or OR4 (N993, N981, N611, N914, N453);
nand NAND3 (N994, N977, N857, N173);
and AND2 (N995, N989, N16);
or OR4 (N996, N994, N562, N271, N102);
xor XOR2 (N997, N991, N183);
xor XOR2 (N998, N997, N485);
xor XOR2 (N999, N990, N997);
xor XOR2 (N1000, N983, N129);
buf BUF1 (N1001, N992);
nor NOR3 (N1002, N998, N564, N836);
buf BUF1 (N1003, N1001);
xor XOR2 (N1004, N995, N997);
buf BUF1 (N1005, N1003);
xor XOR2 (N1006, N1000, N164);
buf BUF1 (N1007, N1005);
not NOT1 (N1008, N982);
and AND3 (N1009, N987, N162, N744);
or OR3 (N1010, N1002, N698, N618);
xor XOR2 (N1011, N999, N660);
nand NAND4 (N1012, N1008, N843, N687, N919);
not NOT1 (N1013, N1009);
xor XOR2 (N1014, N1007, N409);
not NOT1 (N1015, N1004);
not NOT1 (N1016, N1006);
xor XOR2 (N1017, N1010, N751);
xor XOR2 (N1018, N1015, N540);
xor XOR2 (N1019, N996, N661);
not NOT1 (N1020, N1011);
and AND3 (N1021, N1019, N496, N270);
and AND2 (N1022, N1021, N759);
and AND4 (N1023, N1014, N366, N77, N651);
nor NOR2 (N1024, N1013, N55);
nand NAND2 (N1025, N1022, N850);
buf BUF1 (N1026, N993);
xor XOR2 (N1027, N1020, N981);
xor XOR2 (N1028, N1018, N719);
and AND4 (N1029, N1016, N479, N860, N55);
or OR4 (N1030, N1026, N225, N493, N315);
and AND3 (N1031, N1027, N769, N313);
nand NAND3 (N1032, N1028, N770, N27);
or OR4 (N1033, N1032, N657, N641, N267);
and AND2 (N1034, N1033, N793);
not NOT1 (N1035, N1024);
nand NAND3 (N1036, N1023, N224, N819);
not NOT1 (N1037, N1031);
buf BUF1 (N1038, N1037);
or OR2 (N1039, N1025, N277);
or OR4 (N1040, N1039, N784, N185, N269);
or OR3 (N1041, N1017, N630, N710);
nor NOR4 (N1042, N1041, N295, N855, N182);
nor NOR2 (N1043, N1030, N661);
and AND3 (N1044, N1043, N436, N918);
nand NAND3 (N1045, N1036, N409, N800);
or OR3 (N1046, N1034, N808, N718);
nand NAND2 (N1047, N1040, N82);
xor XOR2 (N1048, N1012, N896);
nor NOR4 (N1049, N1046, N754, N937, N1030);
nor NOR3 (N1050, N1045, N608, N660);
or OR4 (N1051, N1038, N330, N854, N340);
buf BUF1 (N1052, N1035);
not NOT1 (N1053, N1042);
xor XOR2 (N1054, N1044, N336);
nor NOR2 (N1055, N963, N918);
or OR3 (N1056, N1029, N632, N969);
nand NAND4 (N1057, N1054, N187, N45, N170);
buf BUF1 (N1058, N1056);
buf BUF1 (N1059, N1057);
xor XOR2 (N1060, N1049, N90);
nand NAND4 (N1061, N1058, N110, N781, N797);
and AND4 (N1062, N1060, N476, N1025, N389);
xor XOR2 (N1063, N1050, N535);
nand NAND4 (N1064, N1051, N356, N108, N947);
nand NAND4 (N1065, N1061, N775, N905, N922);
xor XOR2 (N1066, N1064, N190);
and AND3 (N1067, N1066, N369, N407);
buf BUF1 (N1068, N1053);
buf BUF1 (N1069, N1047);
nor NOR2 (N1070, N1055, N388);
xor XOR2 (N1071, N1062, N108);
not NOT1 (N1072, N1052);
nand NAND4 (N1073, N1068, N665, N971, N854);
or OR4 (N1074, N1072, N762, N92, N1021);
nor NOR4 (N1075, N1059, N815, N968, N1031);
or OR2 (N1076, N1067, N915);
xor XOR2 (N1077, N1063, N763);
buf BUF1 (N1078, N1076);
nor NOR2 (N1079, N1074, N501);
or OR2 (N1080, N1065, N362);
buf BUF1 (N1081, N1077);
and AND3 (N1082, N1080, N953, N545);
buf BUF1 (N1083, N1073);
or OR2 (N1084, N1070, N65);
not NOT1 (N1085, N1048);
and AND2 (N1086, N1078, N535);
not NOT1 (N1087, N1082);
or OR3 (N1088, N1079, N706, N669);
or OR3 (N1089, N1087, N815, N384);
not NOT1 (N1090, N1071);
buf BUF1 (N1091, N1081);
and AND2 (N1092, N1083, N667);
xor XOR2 (N1093, N1075, N410);
nand NAND2 (N1094, N1093, N104);
not NOT1 (N1095, N1084);
nand NAND2 (N1096, N1092, N1016);
or OR3 (N1097, N1090, N729, N821);
not NOT1 (N1098, N1096);
or OR2 (N1099, N1091, N121);
xor XOR2 (N1100, N1088, N704);
and AND3 (N1101, N1099, N116, N1019);
xor XOR2 (N1102, N1100, N25);
nor NOR2 (N1103, N1097, N406);
and AND4 (N1104, N1069, N59, N491, N1097);
buf BUF1 (N1105, N1103);
or OR3 (N1106, N1104, N338, N289);
or OR3 (N1107, N1105, N435, N77);
nand NAND4 (N1108, N1101, N958, N536, N820);
not NOT1 (N1109, N1106);
or OR3 (N1110, N1085, N837, N136);
and AND2 (N1111, N1095, N633);
and AND2 (N1112, N1102, N1066);
nor NOR4 (N1113, N1108, N1072, N940, N763);
nand NAND2 (N1114, N1094, N578);
not NOT1 (N1115, N1112);
or OR2 (N1116, N1086, N1058);
nor NOR4 (N1117, N1111, N466, N454, N1082);
or OR2 (N1118, N1114, N193);
or OR2 (N1119, N1109, N193);
buf BUF1 (N1120, N1107);
and AND4 (N1121, N1115, N507, N669, N558);
not NOT1 (N1122, N1119);
not NOT1 (N1123, N1113);
buf BUF1 (N1124, N1117);
xor XOR2 (N1125, N1121, N879);
or OR2 (N1126, N1110, N305);
and AND4 (N1127, N1098, N887, N203, N927);
not NOT1 (N1128, N1116);
nor NOR3 (N1129, N1124, N162, N405);
nor NOR2 (N1130, N1129, N914);
not NOT1 (N1131, N1123);
not NOT1 (N1132, N1128);
nand NAND3 (N1133, N1089, N754, N985);
xor XOR2 (N1134, N1131, N203);
or OR3 (N1135, N1127, N544, N968);
nand NAND4 (N1136, N1120, N630, N395, N83);
nand NAND2 (N1137, N1135, N638);
xor XOR2 (N1138, N1122, N1058);
nor NOR4 (N1139, N1126, N1090, N470, N113);
nand NAND4 (N1140, N1130, N448, N52, N4);
nand NAND4 (N1141, N1139, N1117, N376, N207);
nor NOR4 (N1142, N1133, N557, N260, N731);
xor XOR2 (N1143, N1138, N268);
nor NOR3 (N1144, N1134, N413, N299);
or OR3 (N1145, N1142, N194, N1031);
nor NOR2 (N1146, N1144, N615);
buf BUF1 (N1147, N1146);
nor NOR4 (N1148, N1140, N1073, N400, N756);
or OR4 (N1149, N1125, N878, N712, N347);
xor XOR2 (N1150, N1143, N872);
not NOT1 (N1151, N1150);
nand NAND4 (N1152, N1136, N1139, N1004, N152);
or OR4 (N1153, N1149, N725, N49, N633);
buf BUF1 (N1154, N1153);
nor NOR2 (N1155, N1151, N683);
nor NOR4 (N1156, N1155, N353, N982, N993);
or OR3 (N1157, N1118, N635, N515);
nor NOR4 (N1158, N1154, N1077, N605, N1126);
and AND4 (N1159, N1148, N975, N855, N495);
nand NAND4 (N1160, N1145, N145, N576, N329);
nand NAND4 (N1161, N1141, N842, N628, N34);
nor NOR3 (N1162, N1147, N55, N365);
or OR4 (N1163, N1161, N110, N372, N198);
nand NAND3 (N1164, N1156, N169, N677);
nor NOR2 (N1165, N1160, N123);
nand NAND3 (N1166, N1132, N728, N1030);
xor XOR2 (N1167, N1137, N804);
nand NAND2 (N1168, N1165, N498);
nor NOR3 (N1169, N1166, N43, N586);
xor XOR2 (N1170, N1169, N223);
and AND4 (N1171, N1152, N424, N781, N931);
or OR3 (N1172, N1159, N650, N1084);
or OR3 (N1173, N1167, N130, N410);
buf BUF1 (N1174, N1171);
nor NOR3 (N1175, N1170, N273, N99);
not NOT1 (N1176, N1173);
not NOT1 (N1177, N1158);
and AND4 (N1178, N1162, N77, N347, N987);
and AND3 (N1179, N1178, N793, N323);
not NOT1 (N1180, N1157);
and AND4 (N1181, N1175, N548, N225, N856);
buf BUF1 (N1182, N1180);
and AND4 (N1183, N1163, N87, N739, N1074);
and AND4 (N1184, N1168, N517, N272, N99);
not NOT1 (N1185, N1181);
nand NAND4 (N1186, N1182, N893, N626, N624);
buf BUF1 (N1187, N1177);
and AND3 (N1188, N1184, N772, N192);
not NOT1 (N1189, N1174);
or OR2 (N1190, N1187, N313);
and AND4 (N1191, N1164, N381, N1108, N840);
buf BUF1 (N1192, N1190);
nand NAND4 (N1193, N1186, N480, N1168, N794);
nand NAND2 (N1194, N1191, N701);
buf BUF1 (N1195, N1189);
not NOT1 (N1196, N1193);
not NOT1 (N1197, N1183);
nand NAND3 (N1198, N1179, N995, N668);
nor NOR2 (N1199, N1185, N312);
xor XOR2 (N1200, N1194, N255);
buf BUF1 (N1201, N1198);
or OR2 (N1202, N1196, N1135);
buf BUF1 (N1203, N1172);
nand NAND3 (N1204, N1201, N1134, N86);
or OR4 (N1205, N1192, N449, N1068, N614);
nor NOR4 (N1206, N1200, N1140, N63, N465);
nand NAND4 (N1207, N1188, N331, N942, N741);
not NOT1 (N1208, N1199);
nand NAND3 (N1209, N1208, N789, N1038);
buf BUF1 (N1210, N1197);
nor NOR2 (N1211, N1209, N123);
xor XOR2 (N1212, N1202, N1166);
or OR4 (N1213, N1211, N933, N1051, N803);
and AND2 (N1214, N1204, N684);
and AND3 (N1215, N1203, N1018, N1168);
not NOT1 (N1216, N1195);
or OR3 (N1217, N1214, N214, N404);
buf BUF1 (N1218, N1215);
nor NOR3 (N1219, N1213, N80, N216);
buf BUF1 (N1220, N1216);
nand NAND3 (N1221, N1176, N1199, N376);
not NOT1 (N1222, N1217);
nand NAND3 (N1223, N1222, N85, N241);
nor NOR4 (N1224, N1207, N29, N224, N1141);
not NOT1 (N1225, N1212);
or OR4 (N1226, N1219, N418, N256, N606);
buf BUF1 (N1227, N1224);
nand NAND2 (N1228, N1210, N1210);
and AND2 (N1229, N1220, N700);
xor XOR2 (N1230, N1225, N1113);
nand NAND2 (N1231, N1230, N175);
nor NOR2 (N1232, N1205, N172);
buf BUF1 (N1233, N1223);
not NOT1 (N1234, N1228);
xor XOR2 (N1235, N1221, N957);
or OR2 (N1236, N1227, N801);
nand NAND2 (N1237, N1226, N983);
or OR3 (N1238, N1231, N444, N1000);
nand NAND3 (N1239, N1236, N92, N582);
and AND4 (N1240, N1232, N197, N201, N417);
and AND3 (N1241, N1206, N965, N833);
and AND4 (N1242, N1235, N170, N707, N751);
not NOT1 (N1243, N1218);
and AND4 (N1244, N1238, N1094, N673, N952);
xor XOR2 (N1245, N1242, N1098);
and AND4 (N1246, N1237, N329, N313, N756);
and AND3 (N1247, N1233, N496, N127);
nor NOR3 (N1248, N1240, N1032, N380);
nor NOR2 (N1249, N1243, N345);
and AND4 (N1250, N1234, N933, N367, N729);
nor NOR2 (N1251, N1248, N482);
not NOT1 (N1252, N1246);
and AND3 (N1253, N1245, N942, N946);
or OR2 (N1254, N1251, N793);
not NOT1 (N1255, N1249);
or OR2 (N1256, N1239, N392);
xor XOR2 (N1257, N1247, N1140);
nand NAND2 (N1258, N1253, N610);
nor NOR3 (N1259, N1250, N817, N830);
xor XOR2 (N1260, N1257, N1179);
xor XOR2 (N1261, N1259, N324);
nor NOR2 (N1262, N1256, N51);
and AND2 (N1263, N1244, N500);
not NOT1 (N1264, N1255);
and AND3 (N1265, N1241, N406, N431);
xor XOR2 (N1266, N1265, N480);
not NOT1 (N1267, N1254);
or OR2 (N1268, N1252, N346);
not NOT1 (N1269, N1268);
and AND2 (N1270, N1269, N1265);
xor XOR2 (N1271, N1267, N13);
or OR4 (N1272, N1266, N498, N859, N539);
or OR3 (N1273, N1229, N996, N428);
and AND2 (N1274, N1270, N775);
not NOT1 (N1275, N1263);
nor NOR3 (N1276, N1264, N70, N258);
nand NAND3 (N1277, N1274, N456, N561);
or OR2 (N1278, N1272, N54);
and AND4 (N1279, N1278, N345, N74, N189);
nand NAND4 (N1280, N1262, N556, N756, N1251);
xor XOR2 (N1281, N1260, N1208);
buf BUF1 (N1282, N1271);
buf BUF1 (N1283, N1282);
and AND2 (N1284, N1277, N1035);
buf BUF1 (N1285, N1281);
buf BUF1 (N1286, N1258);
not NOT1 (N1287, N1273);
buf BUF1 (N1288, N1285);
or OR3 (N1289, N1283, N327, N44);
buf BUF1 (N1290, N1289);
xor XOR2 (N1291, N1280, N537);
xor XOR2 (N1292, N1288, N1116);
nand NAND3 (N1293, N1292, N885, N190);
buf BUF1 (N1294, N1287);
nand NAND2 (N1295, N1294, N1068);
xor XOR2 (N1296, N1286, N635);
buf BUF1 (N1297, N1296);
nand NAND4 (N1298, N1261, N806, N255, N1094);
and AND2 (N1299, N1291, N614);
and AND2 (N1300, N1295, N1135);
nor NOR4 (N1301, N1275, N7, N658, N1044);
buf BUF1 (N1302, N1293);
buf BUF1 (N1303, N1276);
buf BUF1 (N1304, N1284);
or OR2 (N1305, N1279, N771);
buf BUF1 (N1306, N1302);
xor XOR2 (N1307, N1305, N228);
nor NOR2 (N1308, N1307, N731);
and AND3 (N1309, N1300, N376, N464);
xor XOR2 (N1310, N1303, N1097);
and AND2 (N1311, N1310, N551);
and AND3 (N1312, N1301, N1237, N164);
and AND4 (N1313, N1308, N166, N147, N1112);
buf BUF1 (N1314, N1312);
buf BUF1 (N1315, N1297);
buf BUF1 (N1316, N1290);
and AND4 (N1317, N1315, N1278, N695, N636);
buf BUF1 (N1318, N1298);
nand NAND4 (N1319, N1306, N80, N1034, N797);
nor NOR2 (N1320, N1313, N1242);
or OR2 (N1321, N1314, N944);
not NOT1 (N1322, N1320);
or OR2 (N1323, N1318, N9);
and AND2 (N1324, N1311, N236);
not NOT1 (N1325, N1304);
xor XOR2 (N1326, N1299, N733);
and AND2 (N1327, N1319, N1008);
nand NAND3 (N1328, N1316, N500, N301);
nor NOR3 (N1329, N1325, N78, N653);
buf BUF1 (N1330, N1322);
buf BUF1 (N1331, N1327);
not NOT1 (N1332, N1328);
not NOT1 (N1333, N1329);
xor XOR2 (N1334, N1332, N462);
buf BUF1 (N1335, N1323);
xor XOR2 (N1336, N1321, N90);
nand NAND3 (N1337, N1334, N922, N645);
or OR2 (N1338, N1333, N460);
not NOT1 (N1339, N1338);
nor NOR4 (N1340, N1331, N1028, N925, N77);
or OR4 (N1341, N1326, N16, N918, N595);
nor NOR2 (N1342, N1339, N744);
buf BUF1 (N1343, N1342);
nor NOR2 (N1344, N1335, N1096);
nor NOR3 (N1345, N1337, N1011, N305);
buf BUF1 (N1346, N1344);
and AND4 (N1347, N1345, N709, N972, N54);
buf BUF1 (N1348, N1341);
nor NOR2 (N1349, N1324, N1010);
nand NAND2 (N1350, N1348, N1173);
xor XOR2 (N1351, N1349, N880);
not NOT1 (N1352, N1350);
buf BUF1 (N1353, N1352);
not NOT1 (N1354, N1309);
xor XOR2 (N1355, N1317, N189);
buf BUF1 (N1356, N1347);
and AND2 (N1357, N1355, N751);
and AND4 (N1358, N1346, N62, N1146, N1051);
buf BUF1 (N1359, N1354);
xor XOR2 (N1360, N1351, N1058);
nand NAND4 (N1361, N1353, N1034, N1190, N765);
xor XOR2 (N1362, N1361, N1136);
nor NOR2 (N1363, N1356, N1087);
xor XOR2 (N1364, N1330, N71);
buf BUF1 (N1365, N1340);
or OR3 (N1366, N1358, N890, N1178);
nor NOR3 (N1367, N1357, N1194, N485);
xor XOR2 (N1368, N1364, N620);
xor XOR2 (N1369, N1366, N885);
and AND2 (N1370, N1368, N1257);
nor NOR4 (N1371, N1369, N103, N220, N1001);
xor XOR2 (N1372, N1359, N431);
or OR4 (N1373, N1336, N1364, N1330, N859);
nand NAND2 (N1374, N1367, N452);
nor NOR2 (N1375, N1343, N1038);
xor XOR2 (N1376, N1373, N422);
not NOT1 (N1377, N1365);
and AND2 (N1378, N1377, N1254);
or OR3 (N1379, N1376, N1162, N951);
nor NOR4 (N1380, N1375, N792, N305, N626);
xor XOR2 (N1381, N1374, N374);
and AND2 (N1382, N1379, N307);
not NOT1 (N1383, N1382);
or OR4 (N1384, N1370, N395, N849, N666);
nand NAND3 (N1385, N1378, N37, N1138);
buf BUF1 (N1386, N1385);
not NOT1 (N1387, N1380);
or OR2 (N1388, N1381, N1143);
nand NAND2 (N1389, N1362, N323);
and AND4 (N1390, N1371, N410, N76, N910);
xor XOR2 (N1391, N1387, N1097);
buf BUF1 (N1392, N1372);
not NOT1 (N1393, N1392);
not NOT1 (N1394, N1363);
xor XOR2 (N1395, N1360, N349);
not NOT1 (N1396, N1393);
nor NOR4 (N1397, N1390, N468, N270, N715);
xor XOR2 (N1398, N1389, N1314);
or OR2 (N1399, N1394, N467);
or OR4 (N1400, N1398, N996, N915, N578);
and AND4 (N1401, N1397, N185, N923, N999);
xor XOR2 (N1402, N1388, N196);
or OR2 (N1403, N1401, N495);
or OR4 (N1404, N1386, N883, N1382, N223);
nor NOR3 (N1405, N1403, N247, N1303);
nand NAND3 (N1406, N1400, N814, N177);
buf BUF1 (N1407, N1399);
or OR3 (N1408, N1396, N937, N1301);
buf BUF1 (N1409, N1407);
not NOT1 (N1410, N1402);
nor NOR2 (N1411, N1409, N869);
and AND2 (N1412, N1404, N385);
or OR3 (N1413, N1410, N1135, N845);
not NOT1 (N1414, N1383);
or OR2 (N1415, N1412, N774);
or OR2 (N1416, N1395, N209);
and AND2 (N1417, N1411, N274);
buf BUF1 (N1418, N1408);
nand NAND4 (N1419, N1391, N552, N590, N1302);
and AND2 (N1420, N1417, N55);
nor NOR3 (N1421, N1413, N1203, N836);
buf BUF1 (N1422, N1421);
or OR4 (N1423, N1384, N631, N1381, N755);
not NOT1 (N1424, N1416);
not NOT1 (N1425, N1420);
not NOT1 (N1426, N1425);
nand NAND4 (N1427, N1422, N1256, N748, N1179);
not NOT1 (N1428, N1406);
and AND3 (N1429, N1418, N522, N544);
or OR3 (N1430, N1419, N1212, N378);
and AND2 (N1431, N1426, N688);
buf BUF1 (N1432, N1424);
not NOT1 (N1433, N1432);
or OR2 (N1434, N1415, N1232);
buf BUF1 (N1435, N1434);
not NOT1 (N1436, N1433);
or OR3 (N1437, N1429, N900, N1264);
or OR3 (N1438, N1427, N523, N1029);
nand NAND3 (N1439, N1437, N1247, N159);
nand NAND2 (N1440, N1431, N268);
buf BUF1 (N1441, N1428);
xor XOR2 (N1442, N1435, N392);
nor NOR2 (N1443, N1405, N1361);
xor XOR2 (N1444, N1414, N229);
nor NOR3 (N1445, N1430, N195, N770);
or OR2 (N1446, N1436, N197);
buf BUF1 (N1447, N1423);
not NOT1 (N1448, N1444);
buf BUF1 (N1449, N1439);
buf BUF1 (N1450, N1442);
nor NOR4 (N1451, N1438, N927, N1101, N627);
not NOT1 (N1452, N1451);
nand NAND3 (N1453, N1446, N232, N819);
buf BUF1 (N1454, N1452);
and AND3 (N1455, N1441, N910, N433);
buf BUF1 (N1456, N1445);
not NOT1 (N1457, N1455);
buf BUF1 (N1458, N1449);
nand NAND3 (N1459, N1443, N47, N891);
or OR3 (N1460, N1440, N6, N172);
and AND4 (N1461, N1447, N524, N328, N608);
and AND3 (N1462, N1448, N543, N1399);
not NOT1 (N1463, N1459);
nor NOR3 (N1464, N1463, N625, N1063);
not NOT1 (N1465, N1462);
xor XOR2 (N1466, N1464, N1451);
or OR3 (N1467, N1457, N931, N1194);
and AND2 (N1468, N1456, N1294);
nor NOR3 (N1469, N1453, N102, N234);
nor NOR2 (N1470, N1450, N890);
buf BUF1 (N1471, N1454);
xor XOR2 (N1472, N1465, N187);
not NOT1 (N1473, N1466);
buf BUF1 (N1474, N1460);
nand NAND2 (N1475, N1474, N194);
and AND2 (N1476, N1471, N1251);
or OR3 (N1477, N1473, N407, N833);
nor NOR4 (N1478, N1476, N290, N1096, N586);
and AND4 (N1479, N1469, N1458, N1, N761);
not NOT1 (N1480, N455);
xor XOR2 (N1481, N1477, N1254);
not NOT1 (N1482, N1479);
nor NOR3 (N1483, N1468, N832, N298);
nand NAND3 (N1484, N1482, N358, N715);
nand NAND4 (N1485, N1467, N852, N764, N969);
not NOT1 (N1486, N1478);
not NOT1 (N1487, N1485);
xor XOR2 (N1488, N1486, N1150);
nand NAND2 (N1489, N1472, N1138);
not NOT1 (N1490, N1480);
nand NAND2 (N1491, N1475, N1362);
or OR4 (N1492, N1487, N1346, N197, N1337);
not NOT1 (N1493, N1488);
and AND2 (N1494, N1461, N960);
buf BUF1 (N1495, N1489);
nor NOR4 (N1496, N1493, N1074, N677, N1224);
xor XOR2 (N1497, N1495, N251);
not NOT1 (N1498, N1490);
and AND3 (N1499, N1496, N238, N218);
not NOT1 (N1500, N1470);
xor XOR2 (N1501, N1497, N1462);
or OR4 (N1502, N1492, N89, N73, N100);
buf BUF1 (N1503, N1491);
not NOT1 (N1504, N1503);
nor NOR4 (N1505, N1481, N473, N1484, N588);
nor NOR4 (N1506, N339, N902, N882, N212);
nand NAND3 (N1507, N1500, N877, N1471);
nand NAND2 (N1508, N1504, N262);
xor XOR2 (N1509, N1498, N1424);
and AND2 (N1510, N1502, N438);
buf BUF1 (N1511, N1509);
xor XOR2 (N1512, N1505, N537);
xor XOR2 (N1513, N1511, N55);
nand NAND4 (N1514, N1508, N753, N450, N645);
buf BUF1 (N1515, N1512);
nand NAND2 (N1516, N1499, N450);
or OR2 (N1517, N1515, N836);
buf BUF1 (N1518, N1513);
not NOT1 (N1519, N1510);
not NOT1 (N1520, N1507);
and AND3 (N1521, N1483, N466, N381);
and AND4 (N1522, N1501, N339, N186, N1052);
xor XOR2 (N1523, N1516, N802);
buf BUF1 (N1524, N1523);
xor XOR2 (N1525, N1518, N283);
buf BUF1 (N1526, N1521);
not NOT1 (N1527, N1520);
and AND2 (N1528, N1517, N1112);
buf BUF1 (N1529, N1524);
nor NOR4 (N1530, N1529, N1386, N104, N425);
and AND2 (N1531, N1519, N102);
buf BUF1 (N1532, N1527);
and AND4 (N1533, N1531, N826, N1375, N561);
buf BUF1 (N1534, N1525);
xor XOR2 (N1535, N1534, N96);
nand NAND3 (N1536, N1522, N1156, N574);
and AND3 (N1537, N1514, N1188, N173);
nor NOR2 (N1538, N1494, N975);
and AND4 (N1539, N1526, N1456, N160, N258);
or OR3 (N1540, N1533, N841, N546);
nor NOR2 (N1541, N1537, N35);
nand NAND2 (N1542, N1539, N807);
nor NOR4 (N1543, N1538, N1523, N126, N41);
nand NAND2 (N1544, N1543, N830);
xor XOR2 (N1545, N1541, N697);
not NOT1 (N1546, N1544);
xor XOR2 (N1547, N1535, N412);
buf BUF1 (N1548, N1547);
nor NOR3 (N1549, N1548, N182, N582);
xor XOR2 (N1550, N1540, N1225);
or OR2 (N1551, N1542, N493);
not NOT1 (N1552, N1549);
and AND3 (N1553, N1530, N1371, N49);
or OR2 (N1554, N1532, N606);
and AND3 (N1555, N1552, N1296, N1017);
or OR3 (N1556, N1528, N412, N1455);
buf BUF1 (N1557, N1553);
and AND2 (N1558, N1550, N1350);
nand NAND3 (N1559, N1551, N1373, N1087);
nor NOR3 (N1560, N1506, N441, N922);
nor NOR2 (N1561, N1545, N80);
not NOT1 (N1562, N1556);
buf BUF1 (N1563, N1561);
and AND4 (N1564, N1546, N888, N739, N673);
buf BUF1 (N1565, N1563);
nor NOR3 (N1566, N1562, N504, N590);
nor NOR3 (N1567, N1565, N5, N172);
xor XOR2 (N1568, N1558, N607);
not NOT1 (N1569, N1554);
not NOT1 (N1570, N1557);
and AND3 (N1571, N1569, N856, N377);
nor NOR3 (N1572, N1536, N1523, N1449);
nor NOR4 (N1573, N1568, N105, N279, N978);
nand NAND2 (N1574, N1570, N1177);
nor NOR3 (N1575, N1555, N1126, N479);
xor XOR2 (N1576, N1559, N41);
not NOT1 (N1577, N1566);
nor NOR4 (N1578, N1574, N275, N569, N1467);
not NOT1 (N1579, N1578);
buf BUF1 (N1580, N1576);
or OR2 (N1581, N1560, N1429);
nand NAND3 (N1582, N1577, N273, N436);
xor XOR2 (N1583, N1571, N61);
buf BUF1 (N1584, N1580);
buf BUF1 (N1585, N1573);
buf BUF1 (N1586, N1583);
nand NAND2 (N1587, N1585, N1420);
and AND2 (N1588, N1587, N1188);
nor NOR2 (N1589, N1572, N656);
and AND2 (N1590, N1581, N1302);
nor NOR3 (N1591, N1584, N303, N833);
or OR4 (N1592, N1582, N295, N656, N423);
nor NOR4 (N1593, N1589, N1081, N1422, N1213);
and AND2 (N1594, N1593, N255);
not NOT1 (N1595, N1567);
and AND4 (N1596, N1588, N300, N1050, N961);
buf BUF1 (N1597, N1590);
and AND4 (N1598, N1597, N337, N1255, N928);
nor NOR4 (N1599, N1592, N1328, N854, N804);
and AND3 (N1600, N1595, N1321, N419);
nor NOR2 (N1601, N1564, N1053);
xor XOR2 (N1602, N1596, N709);
not NOT1 (N1603, N1602);
nand NAND2 (N1604, N1591, N1397);
nand NAND4 (N1605, N1601, N101, N829, N250);
or OR4 (N1606, N1604, N774, N496, N1171);
nand NAND3 (N1607, N1579, N860, N1545);
nor NOR2 (N1608, N1603, N466);
buf BUF1 (N1609, N1605);
nor NOR3 (N1610, N1598, N805, N1185);
nand NAND3 (N1611, N1607, N1229, N1382);
and AND2 (N1612, N1608, N240);
not NOT1 (N1613, N1610);
or OR3 (N1614, N1599, N1075, N1069);
buf BUF1 (N1615, N1594);
xor XOR2 (N1616, N1609, N673);
or OR2 (N1617, N1600, N1242);
or OR4 (N1618, N1611, N758, N1200, N661);
nor NOR4 (N1619, N1612, N573, N1315, N1507);
nand NAND4 (N1620, N1615, N195, N1020, N924);
xor XOR2 (N1621, N1618, N1047);
buf BUF1 (N1622, N1621);
not NOT1 (N1623, N1620);
and AND4 (N1624, N1619, N592, N1258, N49);
nand NAND4 (N1625, N1623, N1444, N836, N473);
or OR4 (N1626, N1622, N1573, N1608, N787);
xor XOR2 (N1627, N1575, N669);
nand NAND2 (N1628, N1617, N530);
buf BUF1 (N1629, N1628);
and AND2 (N1630, N1627, N1181);
buf BUF1 (N1631, N1613);
and AND4 (N1632, N1626, N1149, N8, N907);
not NOT1 (N1633, N1616);
or OR4 (N1634, N1606, N1616, N422, N460);
buf BUF1 (N1635, N1625);
and AND4 (N1636, N1631, N306, N434, N494);
buf BUF1 (N1637, N1614);
nand NAND2 (N1638, N1624, N1423);
not NOT1 (N1639, N1586);
or OR2 (N1640, N1632, N575);
nand NAND2 (N1641, N1634, N137);
not NOT1 (N1642, N1636);
nand NAND2 (N1643, N1638, N681);
xor XOR2 (N1644, N1629, N923);
buf BUF1 (N1645, N1630);
xor XOR2 (N1646, N1641, N148);
buf BUF1 (N1647, N1642);
xor XOR2 (N1648, N1637, N336);
xor XOR2 (N1649, N1633, N1511);
buf BUF1 (N1650, N1645);
not NOT1 (N1651, N1647);
not NOT1 (N1652, N1639);
xor XOR2 (N1653, N1635, N998);
not NOT1 (N1654, N1649);
buf BUF1 (N1655, N1646);
nand NAND2 (N1656, N1651, N183);
not NOT1 (N1657, N1650);
buf BUF1 (N1658, N1640);
or OR4 (N1659, N1655, N1231, N743, N1500);
nand NAND2 (N1660, N1653, N366);
not NOT1 (N1661, N1660);
buf BUF1 (N1662, N1661);
nor NOR3 (N1663, N1662, N777, N587);
xor XOR2 (N1664, N1659, N180);
nand NAND4 (N1665, N1644, N918, N294, N669);
and AND2 (N1666, N1665, N1221);
buf BUF1 (N1667, N1658);
buf BUF1 (N1668, N1657);
not NOT1 (N1669, N1668);
not NOT1 (N1670, N1643);
nand NAND3 (N1671, N1656, N411, N309);
not NOT1 (N1672, N1664);
or OR4 (N1673, N1671, N1074, N1147, N1650);
xor XOR2 (N1674, N1648, N1168);
and AND2 (N1675, N1669, N217);
buf BUF1 (N1676, N1675);
not NOT1 (N1677, N1676);
not NOT1 (N1678, N1654);
nand NAND3 (N1679, N1652, N260, N1218);
or OR2 (N1680, N1663, N973);
xor XOR2 (N1681, N1674, N1413);
xor XOR2 (N1682, N1667, N1457);
xor XOR2 (N1683, N1682, N1682);
nor NOR4 (N1684, N1681, N1069, N747, N484);
not NOT1 (N1685, N1670);
xor XOR2 (N1686, N1679, N424);
nand NAND4 (N1687, N1686, N76, N301, N988);
nand NAND4 (N1688, N1687, N1158, N1662, N1168);
nor NOR2 (N1689, N1683, N133);
nor NOR2 (N1690, N1689, N500);
or OR4 (N1691, N1685, N438, N1212, N1082);
or OR2 (N1692, N1672, N567);
nor NOR3 (N1693, N1666, N1108, N287);
buf BUF1 (N1694, N1678);
buf BUF1 (N1695, N1694);
buf BUF1 (N1696, N1684);
nand NAND3 (N1697, N1673, N1132, N1013);
nor NOR2 (N1698, N1697, N1149);
xor XOR2 (N1699, N1680, N958);
not NOT1 (N1700, N1677);
not NOT1 (N1701, N1698);
not NOT1 (N1702, N1688);
nor NOR4 (N1703, N1700, N754, N80, N329);
not NOT1 (N1704, N1699);
and AND4 (N1705, N1704, N244, N1332, N1549);
not NOT1 (N1706, N1695);
nand NAND3 (N1707, N1701, N770, N1195);
xor XOR2 (N1708, N1693, N975);
or OR2 (N1709, N1705, N1494);
or OR2 (N1710, N1703, N28);
not NOT1 (N1711, N1710);
nand NAND3 (N1712, N1691, N1457, N622);
or OR2 (N1713, N1711, N634);
nor NOR4 (N1714, N1712, N1656, N1295, N368);
and AND4 (N1715, N1708, N1502, N1332, N989);
not NOT1 (N1716, N1706);
not NOT1 (N1717, N1709);
xor XOR2 (N1718, N1702, N763);
not NOT1 (N1719, N1713);
nand NAND3 (N1720, N1696, N628, N91);
and AND3 (N1721, N1690, N505, N181);
not NOT1 (N1722, N1707);
xor XOR2 (N1723, N1692, N1463);
nor NOR2 (N1724, N1714, N1386);
or OR2 (N1725, N1715, N1641);
nor NOR2 (N1726, N1719, N880);
not NOT1 (N1727, N1724);
xor XOR2 (N1728, N1726, N1228);
nor NOR4 (N1729, N1716, N362, N19, N1365);
and AND2 (N1730, N1721, N388);
or OR4 (N1731, N1725, N1274, N1436, N587);
nor NOR3 (N1732, N1727, N27, N1120);
and AND4 (N1733, N1732, N870, N799, N1010);
nor NOR4 (N1734, N1730, N450, N649, N1112);
nand NAND4 (N1735, N1720, N1004, N268, N249);
nor NOR2 (N1736, N1718, N1577);
nand NAND3 (N1737, N1717, N252, N70);
nor NOR2 (N1738, N1736, N850);
or OR2 (N1739, N1722, N582);
not NOT1 (N1740, N1739);
or OR2 (N1741, N1738, N9);
xor XOR2 (N1742, N1723, N1186);
or OR3 (N1743, N1735, N260, N105);
xor XOR2 (N1744, N1733, N1223);
and AND2 (N1745, N1740, N10);
nand NAND3 (N1746, N1742, N854, N516);
nand NAND2 (N1747, N1746, N149);
nor NOR2 (N1748, N1745, N948);
and AND4 (N1749, N1748, N403, N541, N169);
nor NOR3 (N1750, N1737, N1008, N223);
buf BUF1 (N1751, N1728);
not NOT1 (N1752, N1731);
not NOT1 (N1753, N1750);
nand NAND3 (N1754, N1752, N376, N1332);
not NOT1 (N1755, N1749);
not NOT1 (N1756, N1754);
buf BUF1 (N1757, N1743);
nand NAND2 (N1758, N1744, N1521);
and AND3 (N1759, N1734, N1406, N1517);
buf BUF1 (N1760, N1747);
nand NAND4 (N1761, N1729, N1366, N653, N187);
and AND4 (N1762, N1755, N1364, N1501, N1510);
not NOT1 (N1763, N1757);
buf BUF1 (N1764, N1756);
not NOT1 (N1765, N1761);
or OR3 (N1766, N1762, N589, N393);
or OR2 (N1767, N1766, N1526);
not NOT1 (N1768, N1759);
xor XOR2 (N1769, N1767, N1686);
xor XOR2 (N1770, N1768, N105);
nor NOR2 (N1771, N1763, N734);
or OR4 (N1772, N1769, N1391, N326, N1264);
nor NOR2 (N1773, N1770, N341);
not NOT1 (N1774, N1772);
buf BUF1 (N1775, N1751);
not NOT1 (N1776, N1760);
xor XOR2 (N1777, N1765, N1568);
buf BUF1 (N1778, N1773);
nor NOR2 (N1779, N1758, N616);
not NOT1 (N1780, N1775);
or OR4 (N1781, N1776, N1669, N533, N1650);
or OR3 (N1782, N1771, N281, N1124);
nand NAND2 (N1783, N1774, N684);
nand NAND2 (N1784, N1779, N582);
not NOT1 (N1785, N1778);
buf BUF1 (N1786, N1777);
not NOT1 (N1787, N1782);
buf BUF1 (N1788, N1783);
buf BUF1 (N1789, N1785);
buf BUF1 (N1790, N1787);
nand NAND2 (N1791, N1741, N1564);
or OR2 (N1792, N1791, N1303);
nor NOR3 (N1793, N1789, N1723, N1209);
and AND4 (N1794, N1781, N936, N1275, N622);
buf BUF1 (N1795, N1786);
and AND4 (N1796, N1793, N1201, N1193, N1253);
and AND2 (N1797, N1795, N144);
and AND2 (N1798, N1792, N1000);
nand NAND3 (N1799, N1764, N1217, N1195);
and AND3 (N1800, N1794, N765, N521);
nor NOR2 (N1801, N1788, N875);
nor NOR4 (N1802, N1800, N1410, N322, N1010);
or OR4 (N1803, N1802, N1624, N1584, N377);
nand NAND2 (N1804, N1780, N1013);
nand NAND2 (N1805, N1753, N1554);
not NOT1 (N1806, N1805);
buf BUF1 (N1807, N1796);
nor NOR4 (N1808, N1806, N546, N222, N1234);
or OR4 (N1809, N1808, N265, N1680, N1401);
nor NOR2 (N1810, N1803, N1138);
nor NOR3 (N1811, N1784, N1769, N1727);
xor XOR2 (N1812, N1809, N593);
xor XOR2 (N1813, N1812, N1208);
not NOT1 (N1814, N1813);
not NOT1 (N1815, N1810);
nand NAND4 (N1816, N1801, N989, N1743, N1087);
nor NOR4 (N1817, N1797, N967, N294, N593);
xor XOR2 (N1818, N1816, N706);
nor NOR3 (N1819, N1798, N1182, N234);
nor NOR4 (N1820, N1819, N440, N320, N254);
xor XOR2 (N1821, N1811, N147);
xor XOR2 (N1822, N1799, N721);
nand NAND4 (N1823, N1815, N889, N1235, N1519);
buf BUF1 (N1824, N1817);
and AND2 (N1825, N1807, N1698);
xor XOR2 (N1826, N1823, N1634);
nor NOR4 (N1827, N1820, N665, N723, N665);
nor NOR2 (N1828, N1822, N1282);
nand NAND4 (N1829, N1814, N273, N1584, N1504);
or OR3 (N1830, N1825, N1564, N1212);
not NOT1 (N1831, N1790);
or OR4 (N1832, N1804, N607, N928, N789);
and AND2 (N1833, N1831, N747);
or OR3 (N1834, N1821, N1166, N110);
or OR2 (N1835, N1832, N993);
and AND3 (N1836, N1829, N455, N1128);
buf BUF1 (N1837, N1834);
xor XOR2 (N1838, N1828, N972);
nand NAND4 (N1839, N1838, N543, N1752, N1250);
nor NOR4 (N1840, N1839, N405, N878, N985);
nor NOR3 (N1841, N1840, N569, N1148);
xor XOR2 (N1842, N1841, N792);
or OR2 (N1843, N1842, N649);
and AND3 (N1844, N1827, N1101, N779);
nand NAND3 (N1845, N1837, N314, N80);
xor XOR2 (N1846, N1818, N544);
buf BUF1 (N1847, N1833);
not NOT1 (N1848, N1830);
or OR2 (N1849, N1847, N1829);
buf BUF1 (N1850, N1843);
buf BUF1 (N1851, N1845);
nor NOR2 (N1852, N1824, N1602);
buf BUF1 (N1853, N1851);
xor XOR2 (N1854, N1835, N728);
and AND3 (N1855, N1850, N1764, N487);
and AND4 (N1856, N1826, N982, N135, N1396);
nand NAND3 (N1857, N1855, N51, N1013);
and AND4 (N1858, N1846, N157, N143, N212);
xor XOR2 (N1859, N1858, N873);
buf BUF1 (N1860, N1856);
or OR2 (N1861, N1857, N104);
nor NOR4 (N1862, N1849, N6, N788, N1134);
and AND3 (N1863, N1862, N1017, N445);
or OR2 (N1864, N1836, N729);
not NOT1 (N1865, N1864);
nand NAND2 (N1866, N1865, N466);
not NOT1 (N1867, N1866);
or OR2 (N1868, N1860, N397);
buf BUF1 (N1869, N1867);
nand NAND2 (N1870, N1868, N1777);
nand NAND2 (N1871, N1848, N560);
or OR3 (N1872, N1871, N124, N1218);
buf BUF1 (N1873, N1854);
buf BUF1 (N1874, N1863);
nor NOR4 (N1875, N1844, N1715, N1497, N1688);
buf BUF1 (N1876, N1859);
buf BUF1 (N1877, N1853);
nor NOR2 (N1878, N1870, N14);
xor XOR2 (N1879, N1869, N688);
not NOT1 (N1880, N1876);
nor NOR4 (N1881, N1852, N1668, N743, N1280);
buf BUF1 (N1882, N1875);
nor NOR3 (N1883, N1872, N870, N1802);
nand NAND2 (N1884, N1880, N956);
or OR3 (N1885, N1879, N207, N418);
buf BUF1 (N1886, N1882);
nand NAND4 (N1887, N1881, N612, N1522, N425);
nor NOR3 (N1888, N1861, N311, N1364);
nor NOR4 (N1889, N1878, N954, N1068, N801);
nand NAND2 (N1890, N1883, N1083);
nor NOR2 (N1891, N1885, N1610);
not NOT1 (N1892, N1890);
xor XOR2 (N1893, N1884, N723);
or OR4 (N1894, N1873, N1459, N718, N1166);
or OR4 (N1895, N1888, N1019, N757, N186);
or OR4 (N1896, N1887, N1624, N599, N213);
nand NAND4 (N1897, N1895, N882, N302, N765);
and AND2 (N1898, N1892, N445);
buf BUF1 (N1899, N1886);
buf BUF1 (N1900, N1896);
buf BUF1 (N1901, N1891);
nor NOR4 (N1902, N1894, N797, N97, N1181);
nand NAND2 (N1903, N1899, N504);
and AND3 (N1904, N1897, N1796, N1850);
and AND4 (N1905, N1898, N1715, N1136, N580);
or OR3 (N1906, N1904, N439, N618);
buf BUF1 (N1907, N1905);
xor XOR2 (N1908, N1902, N1015);
xor XOR2 (N1909, N1907, N1384);
xor XOR2 (N1910, N1901, N37);
and AND4 (N1911, N1877, N1608, N1586, N345);
nand NAND3 (N1912, N1908, N690, N1533);
and AND3 (N1913, N1889, N1516, N958);
not NOT1 (N1914, N1911);
nor NOR2 (N1915, N1914, N519);
xor XOR2 (N1916, N1874, N1507);
not NOT1 (N1917, N1900);
nor NOR3 (N1918, N1906, N1487, N1520);
nand NAND4 (N1919, N1916, N293, N420, N1815);
xor XOR2 (N1920, N1918, N808);
nand NAND2 (N1921, N1915, N201);
nor NOR3 (N1922, N1903, N1302, N911);
or OR2 (N1923, N1909, N1267);
buf BUF1 (N1924, N1921);
and AND3 (N1925, N1919, N533, N703);
or OR3 (N1926, N1910, N1168, N191);
not NOT1 (N1927, N1912);
nor NOR2 (N1928, N1922, N366);
xor XOR2 (N1929, N1927, N1526);
nor NOR4 (N1930, N1924, N577, N1418, N912);
buf BUF1 (N1931, N1925);
and AND2 (N1932, N1893, N382);
nand NAND2 (N1933, N1923, N496);
nor NOR2 (N1934, N1929, N49);
or OR3 (N1935, N1913, N1150, N1916);
or OR2 (N1936, N1932, N335);
nand NAND2 (N1937, N1931, N441);
nand NAND3 (N1938, N1930, N727, N1737);
and AND3 (N1939, N1935, N447, N1806);
nor NOR4 (N1940, N1920, N1920, N1174, N1043);
nor NOR4 (N1941, N1936, N342, N1884, N1255);
and AND3 (N1942, N1917, N765, N1209);
nor NOR3 (N1943, N1942, N1308, N1704);
and AND4 (N1944, N1940, N569, N1395, N382);
and AND4 (N1945, N1926, N54, N1462, N212);
nor NOR2 (N1946, N1944, N90);
buf BUF1 (N1947, N1928);
nand NAND2 (N1948, N1947, N383);
or OR2 (N1949, N1934, N183);
nand NAND4 (N1950, N1945, N1593, N86, N527);
nor NOR2 (N1951, N1937, N1613);
nand NAND4 (N1952, N1951, N1101, N421, N216);
xor XOR2 (N1953, N1946, N782);
buf BUF1 (N1954, N1939);
xor XOR2 (N1955, N1948, N253);
buf BUF1 (N1956, N1938);
nand NAND3 (N1957, N1954, N882, N458);
buf BUF1 (N1958, N1949);
nor NOR3 (N1959, N1950, N477, N1447);
nand NAND3 (N1960, N1956, N298, N1327);
nand NAND2 (N1961, N1953, N284);
not NOT1 (N1962, N1952);
or OR2 (N1963, N1960, N1449);
buf BUF1 (N1964, N1955);
and AND2 (N1965, N1964, N1427);
nor NOR4 (N1966, N1965, N1407, N937, N1454);
nor NOR4 (N1967, N1962, N1456, N497, N1055);
xor XOR2 (N1968, N1959, N102);
not NOT1 (N1969, N1963);
and AND4 (N1970, N1969, N651, N1367, N935);
xor XOR2 (N1971, N1958, N1649);
and AND4 (N1972, N1968, N1066, N1303, N1688);
nor NOR3 (N1973, N1967, N971, N1644);
nand NAND3 (N1974, N1957, N670, N967);
nand NAND3 (N1975, N1974, N378, N541);
or OR2 (N1976, N1943, N549);
xor XOR2 (N1977, N1941, N760);
xor XOR2 (N1978, N1961, N291);
xor XOR2 (N1979, N1973, N717);
not NOT1 (N1980, N1975);
nand NAND2 (N1981, N1933, N94);
nand NAND3 (N1982, N1978, N465, N660);
nor NOR3 (N1983, N1979, N122, N1851);
not NOT1 (N1984, N1977);
xor XOR2 (N1985, N1972, N755);
nor NOR3 (N1986, N1971, N842, N892);
xor XOR2 (N1987, N1983, N1235);
and AND3 (N1988, N1985, N450, N422);
xor XOR2 (N1989, N1976, N953);
buf BUF1 (N1990, N1984);
nor NOR3 (N1991, N1982, N1072, N675);
nand NAND3 (N1992, N1966, N543, N1926);
buf BUF1 (N1993, N1986);
and AND2 (N1994, N1993, N1877);
or OR4 (N1995, N1989, N860, N1288, N993);
xor XOR2 (N1996, N1990, N513);
and AND2 (N1997, N1988, N1184);
nand NAND4 (N1998, N1997, N585, N1841, N1131);
buf BUF1 (N1999, N1992);
and AND2 (N2000, N1998, N245);
and AND4 (N2001, N1991, N1552, N368, N217);
not NOT1 (N2002, N1970);
or OR3 (N2003, N1996, N1945, N644);
buf BUF1 (N2004, N1980);
and AND4 (N2005, N1999, N997, N293, N1929);
nand NAND4 (N2006, N2000, N1556, N1452, N1926);
or OR4 (N2007, N1987, N261, N804, N981);
and AND4 (N2008, N1994, N338, N172, N1424);
nor NOR3 (N2009, N2002, N36, N45);
and AND3 (N2010, N2007, N717, N1084);
and AND4 (N2011, N1995, N385, N459, N382);
buf BUF1 (N2012, N2006);
buf BUF1 (N2013, N2012);
xor XOR2 (N2014, N2001, N431);
not NOT1 (N2015, N2008);
xor XOR2 (N2016, N2010, N863);
xor XOR2 (N2017, N2009, N974);
nor NOR4 (N2018, N2003, N1931, N1722, N1425);
not NOT1 (N2019, N2014);
nor NOR2 (N2020, N2005, N872);
and AND4 (N2021, N2016, N1904, N1849, N620);
buf BUF1 (N2022, N2021);
nand NAND3 (N2023, N2004, N1208, N1174);
nor NOR4 (N2024, N2022, N593, N1182, N628);
or OR2 (N2025, N1981, N1286);
nand NAND4 (N2026, N2015, N1740, N188, N1164);
or OR3 (N2027, N2018, N244, N179);
nand NAND3 (N2028, N2017, N977, N799);
buf BUF1 (N2029, N2028);
or OR2 (N2030, N2026, N1331);
nand NAND2 (N2031, N2023, N1833);
or OR3 (N2032, N2013, N1800, N677);
xor XOR2 (N2033, N2024, N868);
buf BUF1 (N2034, N2032);
or OR2 (N2035, N2031, N268);
not NOT1 (N2036, N2033);
not NOT1 (N2037, N2011);
and AND3 (N2038, N2037, N1126, N285);
nor NOR3 (N2039, N2019, N1089, N1218);
nand NAND3 (N2040, N2027, N1261, N305);
xor XOR2 (N2041, N2038, N546);
xor XOR2 (N2042, N2025, N286);
nand NAND2 (N2043, N2034, N835);
xor XOR2 (N2044, N2035, N1952);
xor XOR2 (N2045, N2042, N209);
xor XOR2 (N2046, N2041, N1748);
not NOT1 (N2047, N2030);
nor NOR2 (N2048, N2046, N677);
and AND2 (N2049, N2029, N851);
nand NAND3 (N2050, N2036, N639, N1341);
nor NOR2 (N2051, N2047, N1938);
xor XOR2 (N2052, N2044, N289);
not NOT1 (N2053, N2050);
or OR4 (N2054, N2039, N1928, N1640, N1653);
xor XOR2 (N2055, N2045, N1938);
nor NOR2 (N2056, N2043, N387);
not NOT1 (N2057, N2049);
buf BUF1 (N2058, N2040);
not NOT1 (N2059, N2052);
not NOT1 (N2060, N2057);
not NOT1 (N2061, N2020);
xor XOR2 (N2062, N2053, N1904);
not NOT1 (N2063, N2060);
nor NOR2 (N2064, N2062, N856);
nor NOR2 (N2065, N2051, N650);
nor NOR3 (N2066, N2063, N2038, N1576);
or OR3 (N2067, N2054, N1061, N1811);
not NOT1 (N2068, N2055);
nand NAND4 (N2069, N2059, N1410, N189, N1701);
nor NOR2 (N2070, N2056, N2057);
and AND2 (N2071, N2066, N1093);
or OR4 (N2072, N2065, N268, N2026, N617);
xor XOR2 (N2073, N2071, N110);
or OR2 (N2074, N2070, N1500);
or OR3 (N2075, N2068, N270, N437);
buf BUF1 (N2076, N2064);
xor XOR2 (N2077, N2073, N1601);
xor XOR2 (N2078, N2074, N1244);
xor XOR2 (N2079, N2069, N1276);
nor NOR4 (N2080, N2075, N968, N1830, N1851);
not NOT1 (N2081, N2079);
buf BUF1 (N2082, N2061);
or OR2 (N2083, N2080, N1998);
xor XOR2 (N2084, N2083, N1053);
not NOT1 (N2085, N2078);
nor NOR4 (N2086, N2085, N1955, N390, N437);
or OR4 (N2087, N2084, N1243, N1472, N774);
xor XOR2 (N2088, N2058, N1937);
nand NAND3 (N2089, N2086, N148, N488);
not NOT1 (N2090, N2089);
or OR4 (N2091, N2076, N401, N1231, N715);
or OR2 (N2092, N2091, N1369);
not NOT1 (N2093, N2087);
and AND3 (N2094, N2093, N1766, N1548);
xor XOR2 (N2095, N2088, N753);
nand NAND3 (N2096, N2072, N163, N1779);
or OR4 (N2097, N2094, N523, N809, N166);
buf BUF1 (N2098, N2082);
nor NOR4 (N2099, N2095, N197, N1262, N2095);
nand NAND2 (N2100, N2048, N581);
nand NAND3 (N2101, N2097, N1948, N106);
nor NOR2 (N2102, N2090, N1868);
xor XOR2 (N2103, N2098, N874);
and AND3 (N2104, N2101, N1464, N1946);
and AND2 (N2105, N2081, N814);
not NOT1 (N2106, N2077);
nand NAND3 (N2107, N2103, N354, N1108);
nor NOR3 (N2108, N2096, N86, N1565);
nor NOR3 (N2109, N2100, N1555, N162);
not NOT1 (N2110, N2108);
xor XOR2 (N2111, N2099, N90);
xor XOR2 (N2112, N2111, N24);
and AND4 (N2113, N2112, N628, N1456, N722);
not NOT1 (N2114, N2104);
not NOT1 (N2115, N2110);
and AND2 (N2116, N2092, N1647);
nor NOR4 (N2117, N2067, N1299, N1693, N2042);
buf BUF1 (N2118, N2102);
and AND2 (N2119, N2115, N1547);
and AND4 (N2120, N2116, N1721, N496, N107);
xor XOR2 (N2121, N2109, N800);
and AND4 (N2122, N2121, N551, N1947, N1872);
and AND3 (N2123, N2113, N2020, N390);
buf BUF1 (N2124, N2118);
and AND3 (N2125, N2106, N1536, N1738);
xor XOR2 (N2126, N2120, N2119);
nand NAND2 (N2127, N1047, N1443);
xor XOR2 (N2128, N2125, N315);
xor XOR2 (N2129, N2117, N905);
nand NAND4 (N2130, N2107, N1245, N650, N375);
or OR3 (N2131, N2130, N194, N757);
nand NAND3 (N2132, N2131, N630, N243);
buf BUF1 (N2133, N2126);
xor XOR2 (N2134, N2129, N146);
buf BUF1 (N2135, N2123);
or OR4 (N2136, N2122, N1783, N1380, N1761);
buf BUF1 (N2137, N2105);
and AND3 (N2138, N2137, N1066, N1103);
and AND2 (N2139, N2135, N376);
buf BUF1 (N2140, N2134);
buf BUF1 (N2141, N2138);
or OR4 (N2142, N2124, N1347, N1666, N1307);
xor XOR2 (N2143, N2142, N634);
nor NOR4 (N2144, N2141, N1423, N708, N973);
not NOT1 (N2145, N2136);
not NOT1 (N2146, N2143);
nor NOR2 (N2147, N2127, N563);
buf BUF1 (N2148, N2147);
nand NAND2 (N2149, N2146, N1415);
and AND4 (N2150, N2149, N1012, N1981, N1371);
buf BUF1 (N2151, N2133);
or OR3 (N2152, N2114, N872, N107);
and AND3 (N2153, N2150, N508, N1400);
buf BUF1 (N2154, N2128);
buf BUF1 (N2155, N2153);
nor NOR2 (N2156, N2145, N97);
nand NAND3 (N2157, N2132, N1906, N921);
nand NAND4 (N2158, N2156, N1583, N2094, N1775);
nand NAND3 (N2159, N2140, N1698, N989);
xor XOR2 (N2160, N2144, N1679);
not NOT1 (N2161, N2155);
and AND3 (N2162, N2161, N1483, N1646);
nor NOR2 (N2163, N2152, N1006);
buf BUF1 (N2164, N2148);
not NOT1 (N2165, N2160);
not NOT1 (N2166, N2159);
nand NAND2 (N2167, N2154, N1519);
and AND4 (N2168, N2157, N1760, N416, N1573);
buf BUF1 (N2169, N2163);
buf BUF1 (N2170, N2167);
or OR4 (N2171, N2164, N1472, N207, N22);
buf BUF1 (N2172, N2139);
or OR3 (N2173, N2172, N233, N2000);
not NOT1 (N2174, N2169);
nand NAND3 (N2175, N2162, N1725, N1822);
nand NAND3 (N2176, N2158, N2072, N208);
nor NOR2 (N2177, N2168, N2082);
and AND2 (N2178, N2174, N1436);
or OR4 (N2179, N2165, N8, N634, N1498);
or OR2 (N2180, N2175, N591);
or OR2 (N2181, N2173, N10);
xor XOR2 (N2182, N2177, N2076);
not NOT1 (N2183, N2181);
nand NAND3 (N2184, N2182, N1471, N745);
and AND4 (N2185, N2166, N1267, N894, N1316);
or OR4 (N2186, N2185, N1854, N1740, N742);
buf BUF1 (N2187, N2171);
not NOT1 (N2188, N2170);
nand NAND4 (N2189, N2184, N547, N1769, N571);
or OR3 (N2190, N2186, N1573, N1328);
not NOT1 (N2191, N2188);
or OR4 (N2192, N2176, N988, N1992, N1988);
nand NAND3 (N2193, N2190, N1804, N1561);
xor XOR2 (N2194, N2192, N1826);
or OR3 (N2195, N2151, N564, N1769);
buf BUF1 (N2196, N2179);
and AND4 (N2197, N2180, N326, N1422, N789);
or OR3 (N2198, N2189, N189, N2010);
nand NAND2 (N2199, N2198, N1702);
and AND4 (N2200, N2178, N1010, N1772, N1014);
or OR2 (N2201, N2187, N2084);
not NOT1 (N2202, N2193);
or OR4 (N2203, N2194, N1869, N8, N1136);
buf BUF1 (N2204, N2200);
or OR2 (N2205, N2191, N1558);
and AND3 (N2206, N2204, N430, N1597);
or OR4 (N2207, N2196, N962, N1471, N63);
buf BUF1 (N2208, N2207);
buf BUF1 (N2209, N2206);
not NOT1 (N2210, N2197);
nor NOR3 (N2211, N2203, N986, N171);
not NOT1 (N2212, N2210);
xor XOR2 (N2213, N2195, N573);
and AND4 (N2214, N2211, N625, N1747, N1946);
and AND2 (N2215, N2214, N1521);
xor XOR2 (N2216, N2205, N1235);
not NOT1 (N2217, N2215);
buf BUF1 (N2218, N2201);
not NOT1 (N2219, N2213);
and AND2 (N2220, N2219, N92);
xor XOR2 (N2221, N2217, N302);
and AND2 (N2222, N2216, N1237);
and AND4 (N2223, N2209, N162, N1304, N1507);
and AND4 (N2224, N2212, N32, N1373, N427);
buf BUF1 (N2225, N2221);
not NOT1 (N2226, N2218);
xor XOR2 (N2227, N2199, N919);
buf BUF1 (N2228, N2224);
and AND3 (N2229, N2222, N1235, N518);
not NOT1 (N2230, N2229);
buf BUF1 (N2231, N2183);
and AND4 (N2232, N2223, N1907, N2214, N2228);
xor XOR2 (N2233, N76, N1414);
buf BUF1 (N2234, N2233);
xor XOR2 (N2235, N2225, N477);
nand NAND2 (N2236, N2235, N183);
nor NOR2 (N2237, N2232, N655);
nor NOR3 (N2238, N2236, N19, N210);
not NOT1 (N2239, N2220);
and AND4 (N2240, N2231, N1662, N894, N752);
nor NOR4 (N2241, N2240, N1683, N79, N2053);
buf BUF1 (N2242, N2202);
nand NAND4 (N2243, N2238, N1561, N331, N1337);
or OR3 (N2244, N2241, N250, N1604);
buf BUF1 (N2245, N2208);
nor NOR3 (N2246, N2244, N696, N499);
nor NOR3 (N2247, N2234, N1376, N1883);
not NOT1 (N2248, N2239);
or OR3 (N2249, N2243, N55, N1783);
nor NOR4 (N2250, N2246, N1557, N1368, N818);
or OR4 (N2251, N2247, N1337, N293, N1945);
nand NAND4 (N2252, N2226, N1093, N1957, N1561);
xor XOR2 (N2253, N2237, N1065);
not NOT1 (N2254, N2230);
nand NAND3 (N2255, N2250, N941, N340);
nand NAND2 (N2256, N2242, N307);
nor NOR2 (N2257, N2255, N504);
buf BUF1 (N2258, N2253);
nor NOR4 (N2259, N2254, N50, N581, N919);
nor NOR2 (N2260, N2258, N1904);
xor XOR2 (N2261, N2252, N1671);
not NOT1 (N2262, N2260);
or OR3 (N2263, N2249, N121, N759);
nor NOR3 (N2264, N2257, N1123, N637);
or OR3 (N2265, N2245, N2084, N905);
xor XOR2 (N2266, N2227, N739);
and AND3 (N2267, N2251, N1537, N219);
or OR3 (N2268, N2263, N617, N1215);
buf BUF1 (N2269, N2256);
xor XOR2 (N2270, N2261, N2218);
nand NAND4 (N2271, N2266, N605, N1129, N904);
buf BUF1 (N2272, N2248);
not NOT1 (N2273, N2271);
buf BUF1 (N2274, N2259);
nand NAND2 (N2275, N2270, N1366);
buf BUF1 (N2276, N2268);
not NOT1 (N2277, N2264);
and AND3 (N2278, N2273, N1926, N1089);
nand NAND3 (N2279, N2275, N1311, N1762);
and AND2 (N2280, N2276, N2236);
not NOT1 (N2281, N2274);
buf BUF1 (N2282, N2269);
not NOT1 (N2283, N2265);
and AND3 (N2284, N2262, N708, N1207);
xor XOR2 (N2285, N2277, N349);
buf BUF1 (N2286, N2284);
and AND4 (N2287, N2281, N1357, N392, N1213);
nand NAND2 (N2288, N2282, N445);
nand NAND4 (N2289, N2280, N1013, N1704, N441);
or OR3 (N2290, N2289, N68, N1879);
or OR4 (N2291, N2267, N1646, N87, N2218);
nand NAND3 (N2292, N2279, N1684, N156);
or OR3 (N2293, N2286, N1359, N1636);
xor XOR2 (N2294, N2292, N1462);
nor NOR2 (N2295, N2285, N2109);
or OR2 (N2296, N2293, N360);
or OR2 (N2297, N2278, N1643);
nand NAND3 (N2298, N2296, N1539, N2163);
or OR2 (N2299, N2297, N370);
buf BUF1 (N2300, N2288);
xor XOR2 (N2301, N2294, N612);
nor NOR2 (N2302, N2290, N2091);
nor NOR4 (N2303, N2287, N1530, N1454, N170);
and AND3 (N2304, N2298, N1203, N2224);
and AND3 (N2305, N2283, N1128, N1394);
or OR4 (N2306, N2299, N735, N2091, N1535);
nand NAND3 (N2307, N2303, N338, N1889);
or OR3 (N2308, N2301, N1930, N123);
and AND4 (N2309, N2304, N71, N10, N2108);
nor NOR2 (N2310, N2300, N1726);
xor XOR2 (N2311, N2306, N1675);
not NOT1 (N2312, N2308);
buf BUF1 (N2313, N2309);
buf BUF1 (N2314, N2313);
buf BUF1 (N2315, N2311);
buf BUF1 (N2316, N2310);
or OR3 (N2317, N2307, N453, N826);
nand NAND2 (N2318, N2302, N1366);
and AND3 (N2319, N2312, N1209, N1338);
or OR3 (N2320, N2316, N2262, N676);
xor XOR2 (N2321, N2317, N1351);
not NOT1 (N2322, N2319);
nand NAND2 (N2323, N2315, N984);
nand NAND4 (N2324, N2295, N1560, N1958, N108);
not NOT1 (N2325, N2291);
not NOT1 (N2326, N2314);
nor NOR4 (N2327, N2272, N972, N1102, N1507);
and AND3 (N2328, N2318, N2324, N1597);
nand NAND4 (N2329, N1036, N813, N1231, N2303);
buf BUF1 (N2330, N2320);
xor XOR2 (N2331, N2305, N1018);
xor XOR2 (N2332, N2323, N1438);
and AND3 (N2333, N2321, N1909, N2270);
nand NAND2 (N2334, N2332, N1873);
xor XOR2 (N2335, N2325, N34);
nor NOR3 (N2336, N2334, N777, N2282);
buf BUF1 (N2337, N2330);
not NOT1 (N2338, N2328);
buf BUF1 (N2339, N2327);
or OR3 (N2340, N2333, N120, N2042);
buf BUF1 (N2341, N2339);
not NOT1 (N2342, N2335);
or OR4 (N2343, N2338, N1157, N1357, N1316);
nor NOR4 (N2344, N2337, N1403, N1204, N1117);
or OR3 (N2345, N2329, N524, N2086);
or OR2 (N2346, N2340, N2260);
buf BUF1 (N2347, N2341);
buf BUF1 (N2348, N2345);
xor XOR2 (N2349, N2326, N417);
xor XOR2 (N2350, N2336, N642);
and AND2 (N2351, N2344, N1946);
nand NAND2 (N2352, N2349, N1486);
nand NAND4 (N2353, N2331, N2235, N2259, N502);
xor XOR2 (N2354, N2353, N1528);
not NOT1 (N2355, N2343);
nor NOR2 (N2356, N2346, N876);
nand NAND3 (N2357, N2348, N112, N1437);
not NOT1 (N2358, N2322);
and AND3 (N2359, N2357, N1517, N815);
not NOT1 (N2360, N2358);
buf BUF1 (N2361, N2347);
and AND3 (N2362, N2354, N1191, N1245);
and AND3 (N2363, N2360, N1932, N1796);
not NOT1 (N2364, N2350);
nor NOR3 (N2365, N2359, N2157, N320);
and AND2 (N2366, N2355, N1345);
not NOT1 (N2367, N2352);
or OR4 (N2368, N2362, N2058, N1995, N436);
buf BUF1 (N2369, N2351);
nand NAND2 (N2370, N2367, N232);
not NOT1 (N2371, N2342);
nor NOR4 (N2372, N2364, N1261, N300, N358);
or OR3 (N2373, N2369, N819, N1822);
or OR2 (N2374, N2361, N1942);
or OR4 (N2375, N2371, N1950, N1135, N1776);
xor XOR2 (N2376, N2372, N2305);
not NOT1 (N2377, N2366);
nor NOR3 (N2378, N2363, N1088, N1495);
buf BUF1 (N2379, N2377);
or OR3 (N2380, N2356, N658, N345);
and AND4 (N2381, N2375, N1768, N1305, N1543);
nor NOR3 (N2382, N2365, N2288, N2333);
buf BUF1 (N2383, N2370);
buf BUF1 (N2384, N2381);
xor XOR2 (N2385, N2384, N1366);
nor NOR2 (N2386, N2376, N1612);
xor XOR2 (N2387, N2368, N2326);
not NOT1 (N2388, N2379);
nor NOR4 (N2389, N2382, N89, N729, N899);
not NOT1 (N2390, N2387);
xor XOR2 (N2391, N2386, N1555);
not NOT1 (N2392, N2385);
or OR2 (N2393, N2388, N1565);
nor NOR3 (N2394, N2391, N1734, N2259);
nor NOR2 (N2395, N2378, N2261);
or OR4 (N2396, N2373, N390, N2361, N1459);
not NOT1 (N2397, N2380);
xor XOR2 (N2398, N2383, N1054);
nor NOR4 (N2399, N2389, N95, N647, N226);
and AND4 (N2400, N2393, N2316, N1620, N1693);
and AND4 (N2401, N2392, N2088, N1036, N1064);
not NOT1 (N2402, N2397);
nand NAND3 (N2403, N2400, N2376, N469);
nor NOR3 (N2404, N2401, N1369, N998);
nor NOR2 (N2405, N2404, N233);
buf BUF1 (N2406, N2374);
not NOT1 (N2407, N2395);
and AND2 (N2408, N2398, N848);
or OR3 (N2409, N2408, N523, N1215);
or OR4 (N2410, N2407, N614, N2149, N1471);
or OR2 (N2411, N2406, N295);
and AND2 (N2412, N2402, N701);
buf BUF1 (N2413, N2396);
buf BUF1 (N2414, N2403);
nand NAND2 (N2415, N2413, N1363);
nand NAND2 (N2416, N2414, N2197);
nor NOR2 (N2417, N2405, N833);
buf BUF1 (N2418, N2390);
not NOT1 (N2419, N2399);
xor XOR2 (N2420, N2410, N1585);
and AND3 (N2421, N2416, N650, N1928);
buf BUF1 (N2422, N2421);
xor XOR2 (N2423, N2419, N2221);
nor NOR2 (N2424, N2422, N1679);
xor XOR2 (N2425, N2411, N1790);
not NOT1 (N2426, N2418);
buf BUF1 (N2427, N2426);
nor NOR4 (N2428, N2427, N1074, N1561, N841);
nand NAND3 (N2429, N2409, N2118, N1229);
and AND2 (N2430, N2423, N128);
buf BUF1 (N2431, N2412);
buf BUF1 (N2432, N2415);
nor NOR2 (N2433, N2417, N1815);
not NOT1 (N2434, N2431);
xor XOR2 (N2435, N2429, N1455);
not NOT1 (N2436, N2428);
not NOT1 (N2437, N2432);
not NOT1 (N2438, N2434);
and AND3 (N2439, N2438, N1033, N730);
or OR4 (N2440, N2420, N2403, N1436, N2291);
buf BUF1 (N2441, N2440);
and AND3 (N2442, N2436, N2328, N283);
and AND2 (N2443, N2441, N2013);
not NOT1 (N2444, N2437);
or OR2 (N2445, N2433, N1392);
nand NAND3 (N2446, N2435, N1861, N1596);
xor XOR2 (N2447, N2424, N989);
xor XOR2 (N2448, N2425, N166);
and AND3 (N2449, N2443, N236, N1847);
not NOT1 (N2450, N2430);
nand NAND2 (N2451, N2450, N2404);
xor XOR2 (N2452, N2448, N36);
and AND3 (N2453, N2444, N1682, N2208);
xor XOR2 (N2454, N2445, N1038);
or OR4 (N2455, N2442, N895, N2031, N222);
not NOT1 (N2456, N2394);
not NOT1 (N2457, N2451);
nand NAND2 (N2458, N2456, N599);
or OR3 (N2459, N2454, N1498, N1350);
buf BUF1 (N2460, N2452);
xor XOR2 (N2461, N2460, N1181);
xor XOR2 (N2462, N2458, N1297);
and AND3 (N2463, N2447, N13, N1387);
buf BUF1 (N2464, N2449);
or OR3 (N2465, N2457, N1139, N1187);
and AND3 (N2466, N2463, N2425, N370);
not NOT1 (N2467, N2462);
and AND3 (N2468, N2467, N526, N237);
or OR2 (N2469, N2465, N1035);
or OR2 (N2470, N2459, N77);
xor XOR2 (N2471, N2455, N1923);
and AND4 (N2472, N2446, N909, N1325, N1234);
and AND3 (N2473, N2461, N2066, N2423);
nor NOR3 (N2474, N2472, N1178, N713);
xor XOR2 (N2475, N2439, N1996);
or OR3 (N2476, N2464, N2197, N2183);
xor XOR2 (N2477, N2471, N1545);
nand NAND3 (N2478, N2475, N1283, N1307);
buf BUF1 (N2479, N2470);
buf BUF1 (N2480, N2477);
nor NOR3 (N2481, N2478, N2252, N1301);
buf BUF1 (N2482, N2466);
xor XOR2 (N2483, N2482, N2390);
not NOT1 (N2484, N2453);
nand NAND3 (N2485, N2479, N2211, N2460);
not NOT1 (N2486, N2484);
not NOT1 (N2487, N2476);
nor NOR4 (N2488, N2487, N1168, N650, N1175);
nand NAND2 (N2489, N2483, N1600);
and AND2 (N2490, N2480, N790);
nor NOR3 (N2491, N2486, N1668, N2079);
buf BUF1 (N2492, N2481);
nand NAND4 (N2493, N2492, N69, N925, N2038);
or OR2 (N2494, N2490, N52);
nand NAND4 (N2495, N2474, N1931, N1522, N38);
buf BUF1 (N2496, N2473);
not NOT1 (N2497, N2485);
xor XOR2 (N2498, N2493, N1201);
nand NAND3 (N2499, N2489, N1045, N135);
nand NAND2 (N2500, N2491, N1052);
buf BUF1 (N2501, N2468);
or OR2 (N2502, N2498, N506);
nand NAND2 (N2503, N2488, N2285);
nor NOR3 (N2504, N2499, N83, N1343);
not NOT1 (N2505, N2496);
nand NAND3 (N2506, N2497, N1349, N1363);
not NOT1 (N2507, N2503);
nand NAND2 (N2508, N2502, N164);
nor NOR2 (N2509, N2469, N1814);
or OR4 (N2510, N2501, N2045, N1938, N1360);
or OR3 (N2511, N2507, N1443, N1083);
xor XOR2 (N2512, N2505, N248);
or OR2 (N2513, N2510, N2241);
not NOT1 (N2514, N2508);
not NOT1 (N2515, N2513);
and AND2 (N2516, N2509, N1763);
not NOT1 (N2517, N2494);
buf BUF1 (N2518, N2516);
buf BUF1 (N2519, N2512);
nand NAND3 (N2520, N2518, N1014, N2071);
not NOT1 (N2521, N2511);
buf BUF1 (N2522, N2504);
buf BUF1 (N2523, N2520);
and AND2 (N2524, N2506, N282);
not NOT1 (N2525, N2522);
not NOT1 (N2526, N2514);
xor XOR2 (N2527, N2521, N1537);
not NOT1 (N2528, N2526);
buf BUF1 (N2529, N2515);
nand NAND4 (N2530, N2495, N2088, N777, N2026);
not NOT1 (N2531, N2530);
and AND4 (N2532, N2500, N259, N1499, N579);
nand NAND2 (N2533, N2532, N1673);
xor XOR2 (N2534, N2527, N2503);
nor NOR3 (N2535, N2525, N1820, N1161);
nor NOR4 (N2536, N2519, N863, N1220, N1034);
nor NOR4 (N2537, N2531, N1497, N903, N1064);
not NOT1 (N2538, N2534);
nand NAND3 (N2539, N2529, N1703, N2140);
buf BUF1 (N2540, N2535);
nand NAND2 (N2541, N2539, N2421);
buf BUF1 (N2542, N2538);
nand NAND4 (N2543, N2517, N1599, N1084, N2304);
not NOT1 (N2544, N2528);
not NOT1 (N2545, N2536);
nand NAND4 (N2546, N2541, N976, N171, N1648);
or OR2 (N2547, N2542, N2390);
not NOT1 (N2548, N2537);
and AND3 (N2549, N2544, N830, N1517);
xor XOR2 (N2550, N2545, N730);
buf BUF1 (N2551, N2546);
buf BUF1 (N2552, N2550);
and AND2 (N2553, N2540, N1738);
nand NAND4 (N2554, N2552, N2539, N2537, N2254);
buf BUF1 (N2555, N2553);
xor XOR2 (N2556, N2548, N1646);
nor NOR4 (N2557, N2556, N2033, N282, N2080);
buf BUF1 (N2558, N2555);
nand NAND3 (N2559, N2557, N696, N1653);
or OR2 (N2560, N2549, N1105);
xor XOR2 (N2561, N2558, N787);
nor NOR3 (N2562, N2551, N1229, N1543);
buf BUF1 (N2563, N2533);
nand NAND4 (N2564, N2523, N1721, N1992, N536);
nor NOR4 (N2565, N2560, N832, N1118, N1438);
and AND2 (N2566, N2564, N2264);
buf BUF1 (N2567, N2547);
nand NAND4 (N2568, N2562, N2479, N1189, N1238);
not NOT1 (N2569, N2567);
nand NAND4 (N2570, N2524, N151, N2279, N1909);
or OR4 (N2571, N2569, N2244, N1631, N2446);
or OR3 (N2572, N2543, N1530, N801);
nand NAND4 (N2573, N2572, N2247, N1006, N1601);
not NOT1 (N2574, N2554);
nand NAND2 (N2575, N2568, N1140);
and AND3 (N2576, N2559, N2345, N1036);
and AND2 (N2577, N2561, N1159);
and AND2 (N2578, N2574, N1346);
nor NOR4 (N2579, N2571, N1421, N1172, N694);
buf BUF1 (N2580, N2570);
and AND3 (N2581, N2563, N815, N1384);
or OR2 (N2582, N2565, N1866);
not NOT1 (N2583, N2580);
nand NAND2 (N2584, N2583, N59);
not NOT1 (N2585, N2575);
nand NAND2 (N2586, N2566, N127);
and AND2 (N2587, N2577, N1896);
or OR4 (N2588, N2585, N1346, N107, N2336);
buf BUF1 (N2589, N2573);
nand NAND2 (N2590, N2584, N571);
buf BUF1 (N2591, N2587);
and AND3 (N2592, N2581, N2473, N612);
and AND4 (N2593, N2579, N883, N686, N1034);
nand NAND4 (N2594, N2590, N1904, N238, N831);
xor XOR2 (N2595, N2578, N1346);
and AND3 (N2596, N2589, N1976, N762);
buf BUF1 (N2597, N2594);
nand NAND2 (N2598, N2586, N1104);
xor XOR2 (N2599, N2593, N1241);
and AND4 (N2600, N2592, N340, N2372, N799);
xor XOR2 (N2601, N2588, N136);
or OR4 (N2602, N2595, N2350, N339, N2298);
nand NAND2 (N2603, N2591, N1884);
and AND4 (N2604, N2576, N2367, N28, N468);
and AND4 (N2605, N2599, N161, N2344, N1100);
or OR3 (N2606, N2582, N2290, N140);
buf BUF1 (N2607, N2603);
xor XOR2 (N2608, N2596, N68);
buf BUF1 (N2609, N2598);
nor NOR3 (N2610, N2597, N2286, N704);
xor XOR2 (N2611, N2604, N754);
buf BUF1 (N2612, N2601);
not NOT1 (N2613, N2611);
nand NAND3 (N2614, N2600, N2407, N384);
not NOT1 (N2615, N2608);
buf BUF1 (N2616, N2615);
xor XOR2 (N2617, N2612, N1380);
not NOT1 (N2618, N2602);
nand NAND2 (N2619, N2617, N1977);
and AND4 (N2620, N2616, N2495, N1488, N2065);
xor XOR2 (N2621, N2606, N2430);
and AND2 (N2622, N2605, N818);
and AND3 (N2623, N2620, N19, N381);
or OR3 (N2624, N2610, N610, N2403);
buf BUF1 (N2625, N2607);
nand NAND2 (N2626, N2621, N1720);
xor XOR2 (N2627, N2623, N1434);
or OR2 (N2628, N2618, N45);
xor XOR2 (N2629, N2619, N2156);
nand NAND3 (N2630, N2627, N1364, N1522);
buf BUF1 (N2631, N2622);
xor XOR2 (N2632, N2624, N2493);
buf BUF1 (N2633, N2628);
not NOT1 (N2634, N2609);
or OR4 (N2635, N2614, N1744, N1314, N1470);
not NOT1 (N2636, N2630);
nand NAND2 (N2637, N2635, N246);
xor XOR2 (N2638, N2629, N297);
buf BUF1 (N2639, N2613);
xor XOR2 (N2640, N2632, N809);
not NOT1 (N2641, N2638);
buf BUF1 (N2642, N2625);
xor XOR2 (N2643, N2633, N1246);
xor XOR2 (N2644, N2626, N1832);
xor XOR2 (N2645, N2644, N1294);
or OR4 (N2646, N2637, N134, N2399, N730);
not NOT1 (N2647, N2643);
xor XOR2 (N2648, N2641, N2148);
buf BUF1 (N2649, N2634);
or OR2 (N2650, N2636, N1117);
nand NAND2 (N2651, N2639, N87);
and AND3 (N2652, N2647, N836, N431);
and AND3 (N2653, N2649, N1882, N878);
buf BUF1 (N2654, N2642);
xor XOR2 (N2655, N2652, N2556);
or OR4 (N2656, N2645, N1217, N1984, N1823);
and AND2 (N2657, N2650, N705);
not NOT1 (N2658, N2654);
and AND2 (N2659, N2646, N1770);
not NOT1 (N2660, N2640);
nor NOR4 (N2661, N2631, N876, N1156, N2250);
xor XOR2 (N2662, N2655, N1780);
and AND3 (N2663, N2656, N1274, N2633);
buf BUF1 (N2664, N2648);
xor XOR2 (N2665, N2664, N1981);
and AND2 (N2666, N2662, N914);
not NOT1 (N2667, N2653);
and AND2 (N2668, N2663, N2097);
nand NAND3 (N2669, N2659, N374, N356);
or OR3 (N2670, N2668, N525, N737);
nor NOR2 (N2671, N2651, N322);
not NOT1 (N2672, N2670);
buf BUF1 (N2673, N2667);
xor XOR2 (N2674, N2669, N1951);
or OR4 (N2675, N2658, N1914, N828, N1646);
or OR2 (N2676, N2673, N805);
xor XOR2 (N2677, N2674, N1195);
and AND3 (N2678, N2676, N2574, N215);
nand NAND4 (N2679, N2661, N1724, N1622, N568);
or OR4 (N2680, N2672, N2118, N1554, N2333);
nand NAND3 (N2681, N2660, N1623, N2112);
not NOT1 (N2682, N2680);
buf BUF1 (N2683, N2677);
xor XOR2 (N2684, N2681, N2354);
nor NOR2 (N2685, N2682, N1752);
or OR4 (N2686, N2666, N975, N1671, N135);
xor XOR2 (N2687, N2686, N2031);
or OR3 (N2688, N2665, N1258, N480);
nor NOR4 (N2689, N2687, N351, N944, N2244);
nor NOR4 (N2690, N2675, N1452, N2330, N2235);
nor NOR4 (N2691, N2685, N2436, N1141, N2565);
xor XOR2 (N2692, N2689, N54);
not NOT1 (N2693, N2671);
and AND3 (N2694, N2691, N1995, N70);
or OR4 (N2695, N2679, N278, N2639, N2360);
not NOT1 (N2696, N2695);
buf BUF1 (N2697, N2657);
or OR4 (N2698, N2696, N2360, N454, N158);
nand NAND4 (N2699, N2683, N545, N266, N1247);
nand NAND3 (N2700, N2684, N2128, N1080);
xor XOR2 (N2701, N2678, N2436);
or OR4 (N2702, N2697, N1327, N429, N1493);
nor NOR3 (N2703, N2692, N2351, N2549);
not NOT1 (N2704, N2694);
not NOT1 (N2705, N2688);
nand NAND4 (N2706, N2690, N1874, N115, N2178);
nand NAND4 (N2707, N2701, N2405, N836, N2582);
buf BUF1 (N2708, N2702);
nor NOR2 (N2709, N2698, N1100);
nand NAND4 (N2710, N2700, N1708, N2598, N4);
buf BUF1 (N2711, N2704);
xor XOR2 (N2712, N2699, N1053);
or OR4 (N2713, N2710, N2005, N307, N2329);
nand NAND4 (N2714, N2706, N650, N898, N1560);
and AND2 (N2715, N2714, N942);
nor NOR4 (N2716, N2711, N1928, N977, N1240);
nand NAND3 (N2717, N2715, N694, N1394);
nand NAND2 (N2718, N2707, N1115);
nor NOR2 (N2719, N2705, N1703);
not NOT1 (N2720, N2718);
nor NOR4 (N2721, N2713, N57, N504, N2264);
nand NAND3 (N2722, N2716, N605, N1320);
buf BUF1 (N2723, N2722);
xor XOR2 (N2724, N2709, N2344);
not NOT1 (N2725, N2712);
or OR4 (N2726, N2703, N1034, N463, N1417);
xor XOR2 (N2727, N2693, N1875);
nand NAND4 (N2728, N2719, N684, N1124, N359);
buf BUF1 (N2729, N2727);
and AND3 (N2730, N2721, N122, N1032);
and AND3 (N2731, N2730, N655, N1630);
nand NAND2 (N2732, N2708, N11);
buf BUF1 (N2733, N2728);
nand NAND4 (N2734, N2724, N1890, N890, N2727);
not NOT1 (N2735, N2734);
buf BUF1 (N2736, N2735);
buf BUF1 (N2737, N2736);
not NOT1 (N2738, N2737);
xor XOR2 (N2739, N2738, N1449);
nand NAND4 (N2740, N2725, N1631, N1496, N2014);
and AND4 (N2741, N2739, N1584, N122, N1846);
nand NAND3 (N2742, N2717, N2621, N2188);
nor NOR2 (N2743, N2723, N736);
and AND3 (N2744, N2743, N2084, N116);
buf BUF1 (N2745, N2729);
and AND4 (N2746, N2740, N2523, N2455, N117);
not NOT1 (N2747, N2746);
nor NOR3 (N2748, N2733, N1663, N1805);
not NOT1 (N2749, N2731);
not NOT1 (N2750, N2747);
not NOT1 (N2751, N2745);
not NOT1 (N2752, N2742);
or OR3 (N2753, N2744, N682, N30);
nor NOR2 (N2754, N2752, N1921);
buf BUF1 (N2755, N2751);
and AND3 (N2756, N2755, N1547, N1167);
and AND4 (N2757, N2749, N1966, N2532, N2522);
or OR4 (N2758, N2732, N268, N31, N2036);
not NOT1 (N2759, N2756);
xor XOR2 (N2760, N2758, N1475);
and AND4 (N2761, N2754, N2036, N783, N257);
nand NAND3 (N2762, N2748, N239, N2540);
not NOT1 (N2763, N2761);
or OR4 (N2764, N2720, N136, N1170, N1208);
not NOT1 (N2765, N2726);
nand NAND4 (N2766, N2753, N1021, N2295, N2487);
or OR3 (N2767, N2741, N234, N730);
nand NAND3 (N2768, N2757, N2330, N139);
or OR4 (N2769, N2750, N2072, N2754, N2090);
buf BUF1 (N2770, N2769);
nor NOR3 (N2771, N2767, N1288, N772);
xor XOR2 (N2772, N2759, N2561);
nor NOR4 (N2773, N2764, N202, N946, N2058);
nand NAND2 (N2774, N2760, N1820);
not NOT1 (N2775, N2772);
xor XOR2 (N2776, N2774, N60);
nor NOR3 (N2777, N2776, N425, N1121);
nand NAND3 (N2778, N2763, N2524, N214);
and AND4 (N2779, N2778, N2342, N471, N2002);
xor XOR2 (N2780, N2762, N1424);
and AND2 (N2781, N2777, N2473);
not NOT1 (N2782, N2771);
nand NAND3 (N2783, N2766, N2175, N1099);
xor XOR2 (N2784, N2780, N2270);
nand NAND3 (N2785, N2775, N1197, N680);
xor XOR2 (N2786, N2783, N1052);
nand NAND4 (N2787, N2768, N1845, N2430, N1593);
nand NAND3 (N2788, N2784, N1401, N698);
or OR2 (N2789, N2770, N75);
not NOT1 (N2790, N2781);
buf BUF1 (N2791, N2788);
buf BUF1 (N2792, N2789);
nor NOR2 (N2793, N2765, N2037);
nor NOR3 (N2794, N2792, N2577, N2127);
nand NAND3 (N2795, N2794, N1394, N1754);
or OR2 (N2796, N2790, N480);
nand NAND4 (N2797, N2785, N321, N1315, N1585);
nand NAND2 (N2798, N2782, N2080);
nand NAND2 (N2799, N2796, N2013);
and AND2 (N2800, N2786, N1603);
xor XOR2 (N2801, N2779, N1321);
buf BUF1 (N2802, N2791);
xor XOR2 (N2803, N2773, N772);
xor XOR2 (N2804, N2799, N152);
and AND3 (N2805, N2798, N1263, N2269);
nand NAND3 (N2806, N2797, N1831, N1165);
xor XOR2 (N2807, N2801, N2108);
buf BUF1 (N2808, N2802);
buf BUF1 (N2809, N2787);
xor XOR2 (N2810, N2803, N2308);
nor NOR2 (N2811, N2793, N320);
nor NOR4 (N2812, N2807, N417, N1352, N906);
not NOT1 (N2813, N2812);
or OR3 (N2814, N2811, N1933, N2059);
nand NAND4 (N2815, N2809, N1556, N979, N660);
not NOT1 (N2816, N2800);
nor NOR2 (N2817, N2804, N2025);
nand NAND3 (N2818, N2815, N2209, N1739);
nand NAND3 (N2819, N2806, N2025, N928);
or OR2 (N2820, N2814, N1622);
buf BUF1 (N2821, N2820);
and AND2 (N2822, N2813, N2626);
nor NOR2 (N2823, N2795, N347);
not NOT1 (N2824, N2816);
buf BUF1 (N2825, N2810);
and AND3 (N2826, N2825, N1423, N199);
and AND4 (N2827, N2823, N2506, N1550, N1506);
or OR3 (N2828, N2805, N200, N2444);
or OR4 (N2829, N2818, N450, N1558, N1731);
not NOT1 (N2830, N2819);
nand NAND3 (N2831, N2828, N2122, N2656);
and AND2 (N2832, N2829, N394);
buf BUF1 (N2833, N2827);
nand NAND3 (N2834, N2830, N578, N855);
nor NOR3 (N2835, N2808, N2379, N1871);
or OR4 (N2836, N2822, N2477, N1009, N574);
not NOT1 (N2837, N2832);
and AND3 (N2838, N2824, N2367, N662);
buf BUF1 (N2839, N2838);
not NOT1 (N2840, N2839);
xor XOR2 (N2841, N2821, N948);
or OR4 (N2842, N2836, N1946, N2772, N238);
xor XOR2 (N2843, N2826, N2261);
or OR3 (N2844, N2843, N2307, N83);
and AND4 (N2845, N2834, N1165, N2351, N570);
nand NAND3 (N2846, N2833, N2387, N2302);
and AND2 (N2847, N2835, N138);
buf BUF1 (N2848, N2840);
or OR2 (N2849, N2846, N2337);
buf BUF1 (N2850, N2842);
and AND2 (N2851, N2841, N1259);
or OR3 (N2852, N2844, N1857, N2737);
not NOT1 (N2853, N2852);
nor NOR3 (N2854, N2850, N2689, N593);
xor XOR2 (N2855, N2849, N636);
xor XOR2 (N2856, N2845, N1606);
buf BUF1 (N2857, N2854);
nor NOR4 (N2858, N2853, N808, N1800, N2175);
nor NOR2 (N2859, N2851, N432);
nor NOR2 (N2860, N2856, N1028);
xor XOR2 (N2861, N2847, N1399);
nand NAND4 (N2862, N2855, N985, N2738, N556);
or OR3 (N2863, N2859, N2463, N954);
nand NAND2 (N2864, N2858, N1650);
buf BUF1 (N2865, N2831);
or OR4 (N2866, N2862, N935, N1617, N2691);
nand NAND4 (N2867, N2866, N565, N627, N2539);
not NOT1 (N2868, N2857);
or OR2 (N2869, N2868, N287);
buf BUF1 (N2870, N2817);
or OR4 (N2871, N2863, N1283, N1722, N1651);
buf BUF1 (N2872, N2869);
nor NOR4 (N2873, N2870, N2841, N269, N630);
and AND2 (N2874, N2872, N1174);
not NOT1 (N2875, N2864);
nand NAND4 (N2876, N2875, N377, N2560, N52);
buf BUF1 (N2877, N2874);
or OR3 (N2878, N2837, N589, N46);
nor NOR3 (N2879, N2867, N2477, N215);
not NOT1 (N2880, N2878);
and AND4 (N2881, N2848, N721, N2765, N1542);
nor NOR4 (N2882, N2880, N2725, N228, N921);
buf BUF1 (N2883, N2871);
not NOT1 (N2884, N2881);
buf BUF1 (N2885, N2865);
nand NAND4 (N2886, N2885, N1087, N2654, N727);
and AND2 (N2887, N2876, N536);
nor NOR4 (N2888, N2879, N2403, N1984, N1043);
nand NAND2 (N2889, N2887, N1113);
or OR2 (N2890, N2861, N1852);
nor NOR2 (N2891, N2860, N1693);
nor NOR2 (N2892, N2883, N201);
nand NAND4 (N2893, N2890, N1706, N504, N1618);
and AND3 (N2894, N2889, N1374, N294);
or OR3 (N2895, N2886, N530, N1912);
and AND3 (N2896, N2884, N873, N1853);
nor NOR4 (N2897, N2873, N1978, N2442, N698);
and AND3 (N2898, N2892, N320, N152);
nand NAND2 (N2899, N2895, N1197);
and AND3 (N2900, N2882, N244, N1761);
buf BUF1 (N2901, N2897);
nand NAND3 (N2902, N2891, N61, N1841);
xor XOR2 (N2903, N2894, N250);
buf BUF1 (N2904, N2888);
not NOT1 (N2905, N2899);
not NOT1 (N2906, N2901);
buf BUF1 (N2907, N2904);
not NOT1 (N2908, N2905);
nand NAND2 (N2909, N2898, N1272);
or OR4 (N2910, N2908, N706, N243, N1778);
nor NOR4 (N2911, N2902, N478, N1563, N753);
or OR2 (N2912, N2877, N2805);
nor NOR4 (N2913, N2893, N595, N1609, N2178);
and AND3 (N2914, N2910, N2828, N1464);
nor NOR3 (N2915, N2907, N1886, N2688);
xor XOR2 (N2916, N2914, N1821);
not NOT1 (N2917, N2906);
and AND2 (N2918, N2917, N2536);
xor XOR2 (N2919, N2911, N1456);
not NOT1 (N2920, N2918);
not NOT1 (N2921, N2896);
buf BUF1 (N2922, N2916);
or OR3 (N2923, N2919, N1313, N170);
not NOT1 (N2924, N2922);
nor NOR3 (N2925, N2923, N1961, N943);
xor XOR2 (N2926, N2912, N1703);
not NOT1 (N2927, N2909);
not NOT1 (N2928, N2920);
and AND3 (N2929, N2925, N2311, N1036);
or OR4 (N2930, N2929, N63, N1433, N1099);
or OR2 (N2931, N2926, N1000);
nand NAND4 (N2932, N2915, N2617, N826, N2906);
xor XOR2 (N2933, N2930, N1812);
not NOT1 (N2934, N2903);
and AND3 (N2935, N2933, N1748, N621);
xor XOR2 (N2936, N2924, N2228);
or OR3 (N2937, N2921, N370, N1472);
nor NOR2 (N2938, N2932, N849);
nand NAND2 (N2939, N2928, N193);
or OR3 (N2940, N2936, N650, N1656);
xor XOR2 (N2941, N2927, N1024);
nand NAND3 (N2942, N2934, N2144, N1905);
and AND4 (N2943, N2931, N2238, N2256, N2542);
and AND3 (N2944, N2942, N1401, N376);
nand NAND4 (N2945, N2944, N1955, N2464, N2047);
nor NOR2 (N2946, N2940, N1487);
or OR4 (N2947, N2913, N475, N766, N1422);
or OR3 (N2948, N2943, N888, N1630);
nor NOR2 (N2949, N2939, N933);
nand NAND4 (N2950, N2946, N765, N1251, N887);
not NOT1 (N2951, N2937);
not NOT1 (N2952, N2935);
xor XOR2 (N2953, N2947, N2122);
xor XOR2 (N2954, N2949, N1057);
not NOT1 (N2955, N2950);
not NOT1 (N2956, N2938);
nor NOR4 (N2957, N2954, N2261, N1959, N804);
buf BUF1 (N2958, N2941);
buf BUF1 (N2959, N2948);
or OR4 (N2960, N2953, N152, N69, N361);
buf BUF1 (N2961, N2957);
or OR4 (N2962, N2951, N549, N796, N1460);
buf BUF1 (N2963, N2961);
not NOT1 (N2964, N2952);
not NOT1 (N2965, N2964);
xor XOR2 (N2966, N2963, N2185);
xor XOR2 (N2967, N2966, N164);
nand NAND2 (N2968, N2959, N1234);
and AND3 (N2969, N2967, N264, N1735);
and AND2 (N2970, N2960, N1287);
and AND4 (N2971, N2958, N139, N1851, N2292);
nand NAND3 (N2972, N2955, N784, N2066);
buf BUF1 (N2973, N2900);
nand NAND3 (N2974, N2970, N2418, N1709);
xor XOR2 (N2975, N2965, N2);
buf BUF1 (N2976, N2975);
nand NAND2 (N2977, N2974, N1518);
and AND3 (N2978, N2956, N2941, N1487);
or OR4 (N2979, N2978, N104, N278, N554);
not NOT1 (N2980, N2973);
or OR3 (N2981, N2979, N108, N1436);
not NOT1 (N2982, N2980);
xor XOR2 (N2983, N2976, N1282);
or OR3 (N2984, N2981, N332, N232);
xor XOR2 (N2985, N2971, N1689);
not NOT1 (N2986, N2984);
or OR4 (N2987, N2985, N1329, N271, N974);
nand NAND4 (N2988, N2986, N736, N700, N2708);
and AND2 (N2989, N2977, N1820);
or OR4 (N2990, N2983, N1276, N82, N2853);
buf BUF1 (N2991, N2962);
not NOT1 (N2992, N2968);
not NOT1 (N2993, N2987);
and AND2 (N2994, N2989, N946);
nor NOR2 (N2995, N2945, N2669);
buf BUF1 (N2996, N2992);
and AND4 (N2997, N2982, N894, N1184, N237);
xor XOR2 (N2998, N2988, N1800);
nand NAND2 (N2999, N2969, N168);
not NOT1 (N3000, N2972);
buf BUF1 (N3001, N2996);
buf BUF1 (N3002, N2999);
and AND4 (N3003, N2990, N2151, N2460, N902);
nor NOR3 (N3004, N2998, N1939, N113);
and AND2 (N3005, N2991, N543);
or OR2 (N3006, N3003, N885);
not NOT1 (N3007, N2997);
nor NOR3 (N3008, N2995, N457, N1791);
and AND2 (N3009, N2993, N138);
xor XOR2 (N3010, N3005, N2429);
and AND4 (N3011, N3010, N2115, N1659, N585);
not NOT1 (N3012, N3002);
nand NAND4 (N3013, N3004, N2445, N1204, N2399);
not NOT1 (N3014, N3009);
xor XOR2 (N3015, N3012, N1743);
not NOT1 (N3016, N3008);
or OR2 (N3017, N3016, N2812);
endmodule