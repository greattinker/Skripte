// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14;

output N3512,N3513,N3507,N3497,N3505,N3494,N3502,N3508,N3506,N3514;

nand NAND2 (N15, N3, N9);
nand NAND2 (N16, N4, N11);
and AND2 (N17, N10, N14);
nor NOR2 (N18, N6, N7);
nand NAND2 (N19, N12, N9);
not NOT1 (N20, N2);
nor NOR2 (N21, N16, N13);
or OR3 (N22, N1, N5, N2);
not NOT1 (N23, N12);
buf BUF1 (N24, N4);
buf BUF1 (N25, N22);
xor XOR2 (N26, N12, N10);
xor XOR2 (N27, N17, N1);
and AND3 (N28, N24, N23, N23);
nor NOR3 (N29, N12, N26, N26);
xor XOR2 (N30, N18, N17);
or OR2 (N31, N15, N21);
and AND3 (N32, N12, N25, N5);
nand NAND3 (N33, N18, N15, N7);
nor NOR2 (N34, N22, N33);
buf BUF1 (N35, N28);
not NOT1 (N36, N31);
nor NOR2 (N37, N16, N9);
buf BUF1 (N38, N20);
and AND2 (N39, N35, N10);
or OR4 (N40, N29, N8, N6, N6);
nand NAND3 (N41, N36, N10, N16);
buf BUF1 (N42, N30);
buf BUF1 (N43, N34);
xor XOR2 (N44, N43, N20);
buf BUF1 (N45, N37);
and AND3 (N46, N40, N28, N9);
nor NOR2 (N47, N41, N18);
nor NOR3 (N48, N47, N5, N44);
or OR4 (N49, N27, N10, N8, N34);
not NOT1 (N50, N32);
or OR2 (N51, N9, N33);
xor XOR2 (N52, N45, N24);
nor NOR3 (N53, N48, N38, N12);
nor NOR3 (N54, N36, N32, N26);
and AND3 (N55, N51, N7, N38);
or OR2 (N56, N42, N55);
nor NOR2 (N57, N6, N16);
or OR3 (N58, N50, N7, N33);
and AND3 (N59, N57, N42, N1);
and AND3 (N60, N53, N8, N6);
xor XOR2 (N61, N60, N31);
xor XOR2 (N62, N54, N42);
and AND4 (N63, N61, N60, N51, N33);
xor XOR2 (N64, N52, N15);
nor NOR4 (N65, N19, N56, N13, N32);
xor XOR2 (N66, N39, N17);
xor XOR2 (N67, N23, N64);
xor XOR2 (N68, N66, N47);
not NOT1 (N69, N54);
and AND3 (N70, N63, N59, N5);
not NOT1 (N71, N5);
and AND2 (N72, N62, N64);
not NOT1 (N73, N58);
and AND2 (N74, N71, N32);
xor XOR2 (N75, N72, N32);
and AND3 (N76, N67, N5, N6);
nand NAND2 (N77, N68, N20);
and AND3 (N78, N77, N39, N4);
or OR2 (N79, N75, N46);
or OR4 (N80, N28, N39, N44, N77);
or OR3 (N81, N79, N27, N74);
nand NAND4 (N82, N2, N49, N27, N63);
not NOT1 (N83, N37);
nor NOR2 (N84, N76, N46);
and AND4 (N85, N82, N35, N32, N67);
nor NOR2 (N86, N80, N60);
nor NOR2 (N87, N83, N2);
or OR3 (N88, N70, N58, N26);
nor NOR3 (N89, N86, N64, N70);
nor NOR2 (N90, N81, N16);
buf BUF1 (N91, N85);
nor NOR2 (N92, N84, N90);
nand NAND3 (N93, N40, N54, N34);
xor XOR2 (N94, N65, N27);
or OR4 (N95, N91, N31, N93, N19);
nor NOR3 (N96, N55, N57, N67);
nand NAND4 (N97, N73, N78, N52, N14);
and AND2 (N98, N34, N74);
xor XOR2 (N99, N98, N6);
and AND2 (N100, N92, N42);
or OR3 (N101, N95, N27, N54);
nand NAND4 (N102, N100, N19, N39, N76);
buf BUF1 (N103, N99);
or OR3 (N104, N96, N8, N9);
buf BUF1 (N105, N88);
or OR2 (N106, N69, N90);
or OR4 (N107, N102, N50, N22, N92);
or OR4 (N108, N87, N68, N52, N89);
nor NOR3 (N109, N95, N103, N21);
buf BUF1 (N110, N26);
xor XOR2 (N111, N109, N88);
buf BUF1 (N112, N105);
buf BUF1 (N113, N108);
nand NAND4 (N114, N106, N9, N7, N54);
or OR2 (N115, N107, N55);
buf BUF1 (N116, N97);
nor NOR3 (N117, N115, N87, N43);
and AND4 (N118, N117, N73, N9, N82);
nand NAND2 (N119, N118, N42);
or OR2 (N120, N104, N65);
and AND2 (N121, N120, N99);
or OR3 (N122, N114, N11, N87);
and AND3 (N123, N112, N5, N112);
or OR4 (N124, N122, N40, N49, N86);
nor NOR3 (N125, N121, N84, N108);
buf BUF1 (N126, N116);
or OR2 (N127, N119, N111);
or OR3 (N128, N64, N48, N124);
not NOT1 (N129, N64);
and AND4 (N130, N127, N109, N95, N32);
not NOT1 (N131, N130);
not NOT1 (N132, N123);
nor NOR3 (N133, N125, N109, N8);
nor NOR4 (N134, N94, N7, N20, N130);
xor XOR2 (N135, N131, N118);
xor XOR2 (N136, N129, N102);
nand NAND2 (N137, N133, N5);
nor NOR4 (N138, N110, N9, N62, N111);
and AND4 (N139, N135, N12, N131, N80);
nand NAND4 (N140, N136, N15, N4, N123);
buf BUF1 (N141, N138);
not NOT1 (N142, N139);
not NOT1 (N143, N128);
and AND3 (N144, N137, N80, N95);
or OR2 (N145, N143, N86);
buf BUF1 (N146, N113);
and AND4 (N147, N146, N49, N42, N84);
xor XOR2 (N148, N142, N128);
and AND4 (N149, N147, N60, N145, N2);
nand NAND3 (N150, N33, N149, N94);
nand NAND2 (N151, N64, N44);
or OR4 (N152, N151, N20, N99, N70);
xor XOR2 (N153, N141, N22);
and AND3 (N154, N140, N135, N111);
and AND4 (N155, N154, N105, N150, N13);
not NOT1 (N156, N37);
buf BUF1 (N157, N144);
buf BUF1 (N158, N101);
and AND4 (N159, N155, N30, N34, N142);
or OR2 (N160, N126, N30);
nand NAND3 (N161, N160, N65, N81);
nor NOR3 (N162, N148, N17, N16);
xor XOR2 (N163, N157, N86);
xor XOR2 (N164, N159, N68);
and AND2 (N165, N161, N90);
nand NAND4 (N166, N134, N38, N16, N30);
not NOT1 (N167, N162);
nor NOR4 (N168, N132, N102, N31, N136);
nand NAND2 (N169, N156, N139);
buf BUF1 (N170, N165);
buf BUF1 (N171, N158);
nand NAND4 (N172, N169, N164, N46, N23);
not NOT1 (N173, N133);
nand NAND2 (N174, N171, N63);
xor XOR2 (N175, N173, N24);
xor XOR2 (N176, N167, N171);
and AND4 (N177, N163, N59, N99, N107);
or OR2 (N178, N172, N1);
not NOT1 (N179, N152);
or OR3 (N180, N174, N76, N59);
or OR4 (N181, N179, N65, N39, N150);
and AND3 (N182, N168, N22, N132);
or OR3 (N183, N177, N39, N20);
xor XOR2 (N184, N183, N162);
nor NOR3 (N185, N175, N119, N119);
and AND4 (N186, N182, N126, N157, N171);
or OR4 (N187, N185, N141, N106, N117);
and AND3 (N188, N181, N71, N79);
xor XOR2 (N189, N153, N63);
nor NOR2 (N190, N166, N26);
xor XOR2 (N191, N178, N170);
or OR3 (N192, N48, N82, N64);
and AND2 (N193, N189, N16);
and AND2 (N194, N186, N116);
or OR2 (N195, N192, N102);
and AND4 (N196, N188, N144, N140, N144);
nand NAND3 (N197, N190, N10, N41);
or OR3 (N198, N191, N30, N140);
xor XOR2 (N199, N198, N18);
and AND4 (N200, N197, N23, N74, N52);
not NOT1 (N201, N199);
nor NOR4 (N202, N194, N1, N65, N1);
buf BUF1 (N203, N200);
not NOT1 (N204, N201);
nand NAND3 (N205, N203, N172, N84);
nor NOR2 (N206, N193, N81);
nand NAND4 (N207, N196, N186, N58, N63);
nor NOR3 (N208, N176, N201, N130);
nor NOR3 (N209, N204, N177, N83);
or OR3 (N210, N209, N167, N77);
and AND2 (N211, N202, N170);
buf BUF1 (N212, N187);
nor NOR2 (N213, N210, N137);
and AND2 (N214, N195, N65);
or OR2 (N215, N208, N169);
and AND3 (N216, N180, N126, N193);
or OR3 (N217, N214, N152, N65);
nand NAND3 (N218, N215, N87, N57);
xor XOR2 (N219, N218, N104);
nand NAND4 (N220, N217, N150, N166, N216);
nor NOR3 (N221, N185, N190, N86);
not NOT1 (N222, N211);
nor NOR3 (N223, N212, N106, N180);
nor NOR3 (N224, N213, N53, N221);
or OR3 (N225, N37, N146, N219);
xor XOR2 (N226, N125, N112);
and AND4 (N227, N205, N159, N175, N107);
nand NAND3 (N228, N222, N123, N186);
nand NAND3 (N229, N223, N204, N226);
not NOT1 (N230, N216);
nand NAND3 (N231, N220, N52, N228);
nor NOR4 (N232, N93, N126, N37, N40);
not NOT1 (N233, N224);
buf BUF1 (N234, N227);
nand NAND2 (N235, N233, N70);
nor NOR4 (N236, N184, N22, N117, N165);
buf BUF1 (N237, N230);
nor NOR4 (N238, N237, N165, N208, N217);
or OR3 (N239, N207, N209, N209);
xor XOR2 (N240, N229, N136);
xor XOR2 (N241, N225, N194);
xor XOR2 (N242, N240, N241);
nand NAND2 (N243, N173, N141);
nor NOR3 (N244, N242, N100, N24);
xor XOR2 (N245, N235, N192);
or OR3 (N246, N238, N135, N84);
xor XOR2 (N247, N234, N125);
nor NOR3 (N248, N243, N142, N180);
and AND2 (N249, N206, N215);
or OR2 (N250, N239, N5);
and AND4 (N251, N246, N94, N175, N49);
not NOT1 (N252, N249);
or OR4 (N253, N250, N57, N173, N235);
buf BUF1 (N254, N247);
nand NAND4 (N255, N252, N246, N88, N13);
or OR3 (N256, N236, N53, N212);
xor XOR2 (N257, N251, N15);
xor XOR2 (N258, N256, N96);
or OR3 (N259, N254, N128, N258);
or OR4 (N260, N223, N95, N194, N119);
and AND2 (N261, N232, N238);
nor NOR3 (N262, N255, N92, N77);
nor NOR3 (N263, N261, N149, N72);
not NOT1 (N264, N253);
not NOT1 (N265, N264);
nor NOR4 (N266, N259, N44, N28, N142);
xor XOR2 (N267, N248, N196);
nand NAND4 (N268, N263, N211, N262, N99);
and AND2 (N269, N63, N86);
not NOT1 (N270, N231);
xor XOR2 (N271, N268, N74);
not NOT1 (N272, N244);
not NOT1 (N273, N270);
or OR4 (N274, N245, N167, N8, N233);
and AND4 (N275, N260, N269, N178, N179);
not NOT1 (N276, N58);
buf BUF1 (N277, N265);
buf BUF1 (N278, N273);
not NOT1 (N279, N278);
not NOT1 (N280, N266);
and AND2 (N281, N279, N188);
nor NOR2 (N282, N272, N65);
buf BUF1 (N283, N280);
and AND3 (N284, N281, N5, N28);
xor XOR2 (N285, N276, N209);
or OR4 (N286, N284, N221, N137, N162);
and AND4 (N287, N257, N30, N170, N8);
or OR3 (N288, N274, N66, N115);
not NOT1 (N289, N277);
and AND2 (N290, N275, N102);
nor NOR4 (N291, N289, N195, N74, N108);
or OR4 (N292, N267, N167, N178, N201);
and AND4 (N293, N288, N24, N134, N264);
nor NOR3 (N294, N292, N45, N180);
buf BUF1 (N295, N293);
or OR3 (N296, N286, N59, N22);
nor NOR4 (N297, N285, N13, N106, N233);
not NOT1 (N298, N294);
nand NAND2 (N299, N298, N198);
not NOT1 (N300, N282);
and AND2 (N301, N297, N211);
not NOT1 (N302, N287);
xor XOR2 (N303, N271, N272);
buf BUF1 (N304, N295);
buf BUF1 (N305, N290);
xor XOR2 (N306, N300, N235);
nand NAND3 (N307, N296, N301, N95);
xor XOR2 (N308, N213, N154);
not NOT1 (N309, N302);
not NOT1 (N310, N304);
nand NAND4 (N311, N310, N112, N127, N60);
and AND2 (N312, N308, N50);
or OR3 (N313, N312, N53, N181);
or OR3 (N314, N307, N81, N203);
nor NOR4 (N315, N291, N203, N308, N296);
not NOT1 (N316, N313);
buf BUF1 (N317, N303);
buf BUF1 (N318, N305);
nand NAND4 (N319, N317, N305, N42, N172);
nor NOR3 (N320, N318, N28, N63);
not NOT1 (N321, N311);
or OR4 (N322, N316, N37, N180, N13);
not NOT1 (N323, N283);
nand NAND3 (N324, N315, N274, N136);
nor NOR3 (N325, N319, N95, N49);
nand NAND3 (N326, N314, N305, N187);
or OR2 (N327, N325, N272);
and AND3 (N328, N306, N214, N293);
nand NAND2 (N329, N320, N103);
nor NOR2 (N330, N322, N32);
or OR2 (N331, N321, N99);
or OR2 (N332, N329, N50);
not NOT1 (N333, N330);
and AND4 (N334, N309, N43, N243, N229);
not NOT1 (N335, N331);
buf BUF1 (N336, N335);
or OR3 (N337, N328, N310, N281);
nand NAND2 (N338, N337, N254);
not NOT1 (N339, N299);
buf BUF1 (N340, N339);
not NOT1 (N341, N334);
buf BUF1 (N342, N338);
not NOT1 (N343, N342);
buf BUF1 (N344, N327);
xor XOR2 (N345, N333, N249);
buf BUF1 (N346, N336);
not NOT1 (N347, N323);
nand NAND2 (N348, N324, N223);
or OR3 (N349, N348, N302, N228);
and AND4 (N350, N346, N111, N277, N96);
buf BUF1 (N351, N332);
not NOT1 (N352, N349);
buf BUF1 (N353, N350);
nor NOR2 (N354, N351, N35);
nand NAND4 (N355, N347, N125, N288, N208);
nor NOR2 (N356, N355, N107);
nand NAND4 (N357, N353, N270, N13, N171);
nand NAND3 (N358, N357, N294, N256);
or OR3 (N359, N343, N183, N78);
nor NOR2 (N360, N340, N349);
or OR4 (N361, N354, N356, N10, N204);
nor NOR4 (N362, N229, N20, N66, N355);
or OR2 (N363, N360, N257);
nor NOR4 (N364, N362, N194, N264, N48);
nor NOR2 (N365, N358, N113);
nor NOR4 (N366, N365, N290, N54, N165);
not NOT1 (N367, N326);
buf BUF1 (N368, N359);
or OR2 (N369, N366, N265);
nand NAND2 (N370, N364, N283);
nor NOR2 (N371, N344, N208);
nor NOR3 (N372, N370, N213, N99);
buf BUF1 (N373, N367);
nor NOR4 (N374, N368, N150, N16, N78);
xor XOR2 (N375, N361, N197);
buf BUF1 (N376, N345);
xor XOR2 (N377, N371, N111);
buf BUF1 (N378, N369);
buf BUF1 (N379, N374);
nand NAND3 (N380, N379, N112, N310);
and AND3 (N381, N341, N379, N174);
buf BUF1 (N382, N352);
nor NOR2 (N383, N363, N39);
nand NAND2 (N384, N372, N315);
xor XOR2 (N385, N373, N200);
nor NOR2 (N386, N380, N149);
nand NAND2 (N387, N386, N314);
nor NOR3 (N388, N381, N369, N261);
nand NAND2 (N389, N375, N346);
nand NAND4 (N390, N387, N229, N73, N86);
nand NAND2 (N391, N384, N381);
xor XOR2 (N392, N378, N192);
buf BUF1 (N393, N377);
buf BUF1 (N394, N391);
buf BUF1 (N395, N383);
buf BUF1 (N396, N388);
and AND4 (N397, N394, N81, N57, N123);
nand NAND3 (N398, N389, N275, N113);
or OR4 (N399, N376, N289, N125, N280);
not NOT1 (N400, N382);
nor NOR2 (N401, N396, N120);
and AND4 (N402, N392, N21, N32, N162);
xor XOR2 (N403, N398, N10);
nor NOR3 (N404, N393, N393, N283);
not NOT1 (N405, N385);
and AND3 (N406, N395, N101, N330);
nand NAND2 (N407, N397, N88);
buf BUF1 (N408, N404);
buf BUF1 (N409, N390);
or OR3 (N410, N407, N179, N222);
nand NAND2 (N411, N401, N49);
or OR2 (N412, N402, N351);
nor NOR2 (N413, N409, N321);
buf BUF1 (N414, N399);
nand NAND2 (N415, N413, N373);
or OR4 (N416, N408, N258, N392, N164);
or OR4 (N417, N412, N44, N274, N36);
not NOT1 (N418, N405);
not NOT1 (N419, N415);
xor XOR2 (N420, N416, N138);
xor XOR2 (N421, N410, N362);
and AND4 (N422, N400, N50, N208, N107);
and AND4 (N423, N418, N385, N137, N101);
nand NAND2 (N424, N419, N67);
xor XOR2 (N425, N421, N4);
xor XOR2 (N426, N423, N350);
and AND4 (N427, N403, N339, N173, N120);
xor XOR2 (N428, N417, N367);
xor XOR2 (N429, N406, N176);
nand NAND4 (N430, N424, N109, N95, N110);
nand NAND3 (N431, N429, N263, N196);
or OR2 (N432, N426, N282);
or OR2 (N433, N414, N275);
nor NOR4 (N434, N431, N89, N93, N103);
nand NAND3 (N435, N425, N272, N299);
not NOT1 (N436, N427);
xor XOR2 (N437, N428, N77);
or OR2 (N438, N432, N218);
xor XOR2 (N439, N420, N389);
buf BUF1 (N440, N435);
nand NAND2 (N441, N433, N190);
and AND4 (N442, N430, N39, N87, N424);
buf BUF1 (N443, N434);
buf BUF1 (N444, N422);
nor NOR2 (N445, N442, N313);
not NOT1 (N446, N444);
buf BUF1 (N447, N443);
not NOT1 (N448, N438);
buf BUF1 (N449, N441);
and AND2 (N450, N448, N137);
not NOT1 (N451, N449);
nor NOR2 (N452, N446, N81);
or OR4 (N453, N451, N11, N426, N436);
not NOT1 (N454, N97);
nor NOR2 (N455, N450, N86);
not NOT1 (N456, N437);
and AND3 (N457, N456, N2, N411);
and AND3 (N458, N271, N346, N34);
buf BUF1 (N459, N453);
not NOT1 (N460, N452);
nor NOR3 (N461, N457, N260, N341);
nand NAND4 (N462, N459, N53, N169, N201);
or OR2 (N463, N439, N68);
xor XOR2 (N464, N458, N146);
nand NAND4 (N465, N440, N330, N24, N206);
nand NAND3 (N466, N447, N366, N114);
not NOT1 (N467, N445);
nor NOR2 (N468, N465, N262);
nand NAND2 (N469, N454, N295);
not NOT1 (N470, N468);
or OR4 (N471, N461, N222, N201, N148);
or OR4 (N472, N463, N98, N146, N174);
not NOT1 (N473, N471);
xor XOR2 (N474, N460, N341);
or OR2 (N475, N474, N180);
and AND2 (N476, N472, N103);
buf BUF1 (N477, N466);
nor NOR4 (N478, N467, N427, N224, N159);
nor NOR2 (N479, N475, N355);
not NOT1 (N480, N470);
nand NAND3 (N481, N462, N236, N426);
nand NAND3 (N482, N479, N31, N280);
and AND3 (N483, N481, N447, N19);
or OR4 (N484, N483, N244, N168, N45);
and AND4 (N485, N478, N379, N347, N72);
buf BUF1 (N486, N484);
not NOT1 (N487, N473);
xor XOR2 (N488, N487, N268);
nand NAND3 (N489, N486, N147, N86);
or OR3 (N490, N485, N404, N248);
nand NAND3 (N491, N455, N90, N423);
and AND4 (N492, N490, N12, N456, N306);
and AND4 (N493, N464, N173, N442, N322);
and AND2 (N494, N482, N418);
nand NAND4 (N495, N488, N423, N265, N194);
xor XOR2 (N496, N489, N455);
xor XOR2 (N497, N477, N28);
not NOT1 (N498, N476);
buf BUF1 (N499, N492);
or OR4 (N500, N469, N180, N147, N264);
not NOT1 (N501, N497);
or OR2 (N502, N491, N59);
xor XOR2 (N503, N494, N211);
nor NOR3 (N504, N499, N484, N218);
xor XOR2 (N505, N495, N422);
nand NAND2 (N506, N502, N385);
buf BUF1 (N507, N496);
nor NOR3 (N508, N493, N234, N269);
or OR3 (N509, N505, N263, N228);
nand NAND4 (N510, N501, N61, N101, N128);
or OR2 (N511, N509, N255);
or OR4 (N512, N498, N140, N42, N152);
nand NAND4 (N513, N480, N232, N337, N125);
and AND2 (N514, N504, N111);
nand NAND3 (N515, N500, N374, N331);
nor NOR4 (N516, N510, N73, N11, N199);
and AND2 (N517, N513, N424);
buf BUF1 (N518, N506);
not NOT1 (N519, N518);
or OR4 (N520, N511, N383, N459, N61);
not NOT1 (N521, N507);
nand NAND3 (N522, N508, N315, N420);
nor NOR2 (N523, N520, N155);
not NOT1 (N524, N503);
not NOT1 (N525, N516);
xor XOR2 (N526, N515, N186);
xor XOR2 (N527, N526, N146);
nand NAND4 (N528, N524, N409, N348, N184);
not NOT1 (N529, N517);
and AND4 (N530, N519, N458, N370, N271);
and AND4 (N531, N529, N203, N485, N305);
not NOT1 (N532, N514);
xor XOR2 (N533, N525, N508);
buf BUF1 (N534, N532);
nor NOR3 (N535, N531, N459, N110);
nand NAND4 (N536, N534, N527, N234, N459);
nor NOR3 (N537, N187, N495, N405);
nor NOR4 (N538, N535, N341, N281, N49);
not NOT1 (N539, N522);
nand NAND2 (N540, N539, N434);
xor XOR2 (N541, N512, N328);
nor NOR3 (N542, N540, N346, N228);
or OR3 (N543, N538, N146, N183);
xor XOR2 (N544, N542, N492);
nor NOR2 (N545, N523, N534);
buf BUF1 (N546, N543);
and AND2 (N547, N546, N133);
nor NOR4 (N548, N537, N287, N461, N339);
not NOT1 (N549, N521);
buf BUF1 (N550, N544);
nand NAND3 (N551, N550, N15, N550);
nor NOR3 (N552, N541, N384, N125);
nor NOR2 (N553, N536, N234);
nor NOR4 (N554, N553, N189, N96, N530);
buf BUF1 (N555, N140);
and AND3 (N556, N552, N272, N372);
or OR2 (N557, N556, N539);
not NOT1 (N558, N549);
buf BUF1 (N559, N545);
and AND3 (N560, N559, N337, N121);
and AND4 (N561, N533, N148, N322, N237);
nor NOR4 (N562, N561, N18, N158, N216);
buf BUF1 (N563, N562);
and AND3 (N564, N548, N129, N443);
not NOT1 (N565, N554);
nor NOR3 (N566, N551, N199, N87);
xor XOR2 (N567, N558, N404);
and AND4 (N568, N563, N37, N152, N336);
or OR4 (N569, N528, N83, N91, N320);
or OR2 (N570, N557, N558);
xor XOR2 (N571, N564, N483);
not NOT1 (N572, N567);
not NOT1 (N573, N555);
nor NOR2 (N574, N547, N94);
not NOT1 (N575, N573);
not NOT1 (N576, N574);
nor NOR4 (N577, N560, N202, N430, N167);
and AND3 (N578, N569, N83, N57);
buf BUF1 (N579, N568);
buf BUF1 (N580, N575);
not NOT1 (N581, N579);
and AND3 (N582, N566, N254, N85);
nor NOR2 (N583, N578, N495);
or OR3 (N584, N580, N31, N125);
or OR2 (N585, N576, N447);
buf BUF1 (N586, N565);
and AND2 (N587, N586, N277);
buf BUF1 (N588, N585);
nor NOR2 (N589, N588, N266);
not NOT1 (N590, N570);
or OR4 (N591, N582, N174, N272, N240);
nor NOR4 (N592, N572, N436, N127, N423);
and AND3 (N593, N590, N426, N145);
or OR2 (N594, N589, N191);
or OR3 (N595, N594, N185, N291);
nand NAND2 (N596, N587, N312);
not NOT1 (N597, N577);
buf BUF1 (N598, N591);
or OR4 (N599, N595, N409, N455, N249);
and AND2 (N600, N596, N144);
buf BUF1 (N601, N599);
buf BUF1 (N602, N571);
nor NOR3 (N603, N583, N518, N50);
buf BUF1 (N604, N598);
buf BUF1 (N605, N600);
nor NOR2 (N606, N584, N342);
and AND4 (N607, N597, N267, N454, N473);
nor NOR2 (N608, N604, N329);
buf BUF1 (N609, N606);
nand NAND4 (N610, N608, N135, N387, N122);
nor NOR3 (N611, N610, N327, N564);
not NOT1 (N612, N609);
buf BUF1 (N613, N612);
nand NAND4 (N614, N605, N440, N286, N103);
xor XOR2 (N615, N593, N9);
buf BUF1 (N616, N601);
buf BUF1 (N617, N613);
and AND3 (N618, N615, N3, N285);
or OR4 (N619, N602, N126, N318, N564);
or OR3 (N620, N614, N76, N376);
nor NOR3 (N621, N611, N242, N441);
nor NOR2 (N622, N607, N36);
not NOT1 (N623, N617);
buf BUF1 (N624, N592);
buf BUF1 (N625, N620);
xor XOR2 (N626, N619, N90);
not NOT1 (N627, N618);
and AND4 (N628, N603, N289, N607, N163);
buf BUF1 (N629, N624);
nor NOR2 (N630, N621, N221);
buf BUF1 (N631, N622);
nand NAND3 (N632, N630, N297, N277);
and AND4 (N633, N626, N117, N420, N182);
nand NAND3 (N634, N629, N269, N103);
buf BUF1 (N635, N581);
buf BUF1 (N636, N616);
not NOT1 (N637, N628);
nand NAND4 (N638, N623, N385, N24, N146);
xor XOR2 (N639, N634, N332);
or OR2 (N640, N625, N152);
xor XOR2 (N641, N631, N144);
and AND2 (N642, N637, N56);
and AND3 (N643, N636, N58, N628);
nand NAND2 (N644, N638, N262);
nand NAND4 (N645, N640, N23, N431, N412);
nand NAND3 (N646, N627, N253, N100);
xor XOR2 (N647, N632, N337);
and AND2 (N648, N641, N216);
and AND3 (N649, N643, N559, N145);
or OR2 (N650, N649, N646);
not NOT1 (N651, N124);
nand NAND3 (N652, N642, N401, N43);
or OR4 (N653, N639, N626, N635, N26);
or OR2 (N654, N591, N153);
not NOT1 (N655, N653);
not NOT1 (N656, N644);
xor XOR2 (N657, N656, N65);
buf BUF1 (N658, N633);
nor NOR3 (N659, N657, N248, N495);
nor NOR3 (N660, N655, N238, N265);
nor NOR3 (N661, N648, N66, N148);
nand NAND2 (N662, N650, N588);
not NOT1 (N663, N659);
xor XOR2 (N664, N661, N170);
xor XOR2 (N665, N645, N253);
xor XOR2 (N666, N652, N160);
nand NAND4 (N667, N664, N397, N487, N603);
and AND2 (N668, N665, N565);
buf BUF1 (N669, N663);
buf BUF1 (N670, N669);
nor NOR3 (N671, N662, N247, N420);
buf BUF1 (N672, N667);
nor NOR2 (N673, N658, N168);
or OR2 (N674, N671, N480);
and AND3 (N675, N654, N631, N483);
not NOT1 (N676, N674);
xor XOR2 (N677, N673, N137);
buf BUF1 (N678, N675);
not NOT1 (N679, N668);
buf BUF1 (N680, N679);
or OR2 (N681, N670, N654);
or OR4 (N682, N681, N479, N655, N28);
buf BUF1 (N683, N682);
buf BUF1 (N684, N672);
buf BUF1 (N685, N684);
nor NOR3 (N686, N678, N371, N27);
or OR3 (N687, N686, N392, N260);
buf BUF1 (N688, N683);
xor XOR2 (N689, N688, N518);
nor NOR3 (N690, N647, N283, N209);
nand NAND3 (N691, N689, N510, N238);
and AND4 (N692, N685, N99, N513, N329);
buf BUF1 (N693, N651);
not NOT1 (N694, N691);
or OR4 (N695, N677, N1, N408, N14);
or OR2 (N696, N692, N450);
xor XOR2 (N697, N666, N441);
not NOT1 (N698, N695);
or OR2 (N699, N680, N291);
buf BUF1 (N700, N693);
buf BUF1 (N701, N694);
nand NAND2 (N702, N697, N165);
not NOT1 (N703, N702);
not NOT1 (N704, N701);
not NOT1 (N705, N660);
and AND3 (N706, N696, N32, N655);
nand NAND4 (N707, N687, N374, N676, N172);
nor NOR2 (N708, N673, N109);
and AND2 (N709, N699, N212);
and AND3 (N710, N704, N706, N489);
nor NOR3 (N711, N37, N19, N479);
nand NAND3 (N712, N705, N133, N600);
buf BUF1 (N713, N708);
nand NAND2 (N714, N710, N546);
not NOT1 (N715, N709);
xor XOR2 (N716, N690, N675);
and AND3 (N717, N703, N178, N107);
nor NOR2 (N718, N716, N476);
not NOT1 (N719, N718);
nand NAND3 (N720, N700, N344, N78);
and AND2 (N721, N720, N605);
xor XOR2 (N722, N714, N578);
or OR4 (N723, N717, N391, N409, N375);
not NOT1 (N724, N711);
not NOT1 (N725, N707);
buf BUF1 (N726, N724);
nor NOR4 (N727, N722, N308, N478, N6);
buf BUF1 (N728, N715);
buf BUF1 (N729, N728);
not NOT1 (N730, N719);
not NOT1 (N731, N712);
xor XOR2 (N732, N698, N711);
xor XOR2 (N733, N732, N417);
and AND3 (N734, N729, N577, N353);
and AND3 (N735, N725, N4, N679);
or OR4 (N736, N713, N88, N152, N426);
xor XOR2 (N737, N730, N52);
xor XOR2 (N738, N734, N58);
or OR2 (N739, N731, N31);
xor XOR2 (N740, N726, N273);
not NOT1 (N741, N721);
nand NAND2 (N742, N727, N341);
and AND3 (N743, N742, N148, N301);
or OR4 (N744, N740, N81, N728, N89);
nand NAND2 (N745, N735, N93);
nand NAND2 (N746, N737, N636);
nor NOR4 (N747, N733, N31, N236, N537);
or OR4 (N748, N747, N454, N296, N35);
or OR4 (N749, N736, N398, N515, N491);
nor NOR2 (N750, N744, N181);
or OR2 (N751, N739, N268);
and AND4 (N752, N746, N279, N23, N279);
buf BUF1 (N753, N749);
nor NOR2 (N754, N753, N41);
xor XOR2 (N755, N751, N537);
or OR2 (N756, N723, N641);
nand NAND2 (N757, N754, N117);
not NOT1 (N758, N756);
not NOT1 (N759, N743);
nor NOR2 (N760, N745, N348);
nand NAND2 (N761, N738, N543);
or OR2 (N762, N750, N44);
not NOT1 (N763, N755);
xor XOR2 (N764, N760, N337);
and AND3 (N765, N752, N127, N190);
and AND4 (N766, N762, N217, N384, N265);
nor NOR4 (N767, N748, N208, N131, N133);
or OR3 (N768, N761, N167, N655);
nor NOR4 (N769, N763, N262, N405, N313);
buf BUF1 (N770, N769);
and AND4 (N771, N764, N538, N688, N295);
nand NAND4 (N772, N767, N436, N767, N566);
xor XOR2 (N773, N771, N87);
nand NAND3 (N774, N741, N297, N652);
xor XOR2 (N775, N773, N149);
buf BUF1 (N776, N766);
nor NOR3 (N777, N758, N318, N720);
nor NOR3 (N778, N775, N400, N364);
xor XOR2 (N779, N777, N578);
not NOT1 (N780, N759);
nor NOR3 (N781, N780, N637, N675);
nand NAND4 (N782, N757, N71, N356, N360);
and AND3 (N783, N779, N355, N545);
or OR3 (N784, N768, N332, N120);
buf BUF1 (N785, N778);
not NOT1 (N786, N784);
and AND3 (N787, N786, N309, N503);
buf BUF1 (N788, N770);
nand NAND3 (N789, N782, N487, N267);
xor XOR2 (N790, N785, N80);
not NOT1 (N791, N783);
xor XOR2 (N792, N772, N6);
and AND2 (N793, N776, N155);
buf BUF1 (N794, N792);
nor NOR4 (N795, N781, N77, N184, N219);
xor XOR2 (N796, N790, N147);
or OR2 (N797, N793, N17);
xor XOR2 (N798, N796, N117);
or OR3 (N799, N787, N185, N649);
xor XOR2 (N800, N797, N365);
xor XOR2 (N801, N798, N298);
nor NOR2 (N802, N774, N230);
or OR4 (N803, N765, N258, N559, N359);
nand NAND2 (N804, N803, N681);
buf BUF1 (N805, N795);
or OR2 (N806, N799, N32);
nor NOR4 (N807, N788, N608, N411, N255);
buf BUF1 (N808, N804);
nand NAND4 (N809, N801, N675, N618, N210);
and AND2 (N810, N800, N571);
or OR3 (N811, N791, N397, N203);
and AND2 (N812, N806, N805);
or OR3 (N813, N267, N214, N340);
nand NAND3 (N814, N794, N224, N286);
buf BUF1 (N815, N789);
xor XOR2 (N816, N802, N445);
nand NAND4 (N817, N814, N539, N673, N362);
nor NOR2 (N818, N809, N349);
not NOT1 (N819, N815);
nand NAND4 (N820, N810, N514, N197, N614);
nor NOR3 (N821, N818, N463, N316);
and AND2 (N822, N812, N522);
not NOT1 (N823, N807);
or OR3 (N824, N817, N789, N251);
and AND2 (N825, N822, N403);
nor NOR4 (N826, N816, N645, N744, N170);
nand NAND2 (N827, N808, N282);
nor NOR3 (N828, N811, N627, N431);
or OR2 (N829, N821, N813);
not NOT1 (N830, N429);
not NOT1 (N831, N828);
xor XOR2 (N832, N824, N196);
buf BUF1 (N833, N831);
not NOT1 (N834, N825);
or OR4 (N835, N834, N499, N606, N513);
nand NAND4 (N836, N827, N702, N828, N579);
or OR3 (N837, N833, N788, N675);
and AND2 (N838, N823, N402);
buf BUF1 (N839, N826);
not NOT1 (N840, N820);
buf BUF1 (N841, N839);
buf BUF1 (N842, N837);
nor NOR3 (N843, N841, N762, N804);
nor NOR3 (N844, N842, N478, N810);
xor XOR2 (N845, N838, N54);
and AND3 (N846, N829, N134, N41);
or OR3 (N847, N830, N316, N474);
buf BUF1 (N848, N847);
buf BUF1 (N849, N844);
xor XOR2 (N850, N848, N157);
or OR4 (N851, N845, N641, N22, N475);
not NOT1 (N852, N846);
not NOT1 (N853, N835);
and AND2 (N854, N843, N177);
nor NOR2 (N855, N840, N369);
nand NAND2 (N856, N836, N223);
and AND2 (N857, N853, N577);
and AND3 (N858, N854, N837, N367);
or OR2 (N859, N858, N593);
and AND4 (N860, N850, N822, N178, N446);
and AND4 (N861, N855, N145, N315, N175);
or OR3 (N862, N851, N350, N841);
buf BUF1 (N863, N859);
not NOT1 (N864, N861);
xor XOR2 (N865, N849, N796);
xor XOR2 (N866, N832, N748);
and AND2 (N867, N862, N248);
xor XOR2 (N868, N864, N560);
buf BUF1 (N869, N867);
or OR4 (N870, N868, N765, N233, N572);
and AND2 (N871, N866, N387);
or OR4 (N872, N865, N836, N375, N765);
not NOT1 (N873, N857);
not NOT1 (N874, N871);
not NOT1 (N875, N869);
nand NAND4 (N876, N852, N519, N555, N805);
nor NOR4 (N877, N856, N308, N136, N825);
nand NAND2 (N878, N873, N332);
not NOT1 (N879, N877);
xor XOR2 (N880, N860, N509);
buf BUF1 (N881, N872);
not NOT1 (N882, N881);
nand NAND3 (N883, N819, N367, N359);
xor XOR2 (N884, N875, N760);
or OR3 (N885, N883, N559, N221);
not NOT1 (N886, N874);
nand NAND2 (N887, N863, N835);
or OR3 (N888, N887, N619, N389);
nor NOR3 (N889, N885, N566, N188);
not NOT1 (N890, N889);
nor NOR2 (N891, N870, N607);
nand NAND2 (N892, N886, N463);
xor XOR2 (N893, N879, N74);
or OR3 (N894, N890, N498, N806);
buf BUF1 (N895, N894);
not NOT1 (N896, N893);
not NOT1 (N897, N876);
and AND2 (N898, N897, N353);
nand NAND3 (N899, N898, N805, N145);
and AND4 (N900, N899, N150, N609, N577);
xor XOR2 (N901, N878, N774);
or OR2 (N902, N891, N498);
xor XOR2 (N903, N901, N406);
nor NOR3 (N904, N903, N16, N489);
not NOT1 (N905, N892);
or OR2 (N906, N882, N386);
or OR3 (N907, N902, N336, N875);
or OR3 (N908, N905, N657, N343);
or OR4 (N909, N884, N367, N355, N172);
buf BUF1 (N910, N895);
and AND4 (N911, N910, N381, N726, N432);
nand NAND4 (N912, N900, N669, N389, N720);
not NOT1 (N913, N907);
or OR2 (N914, N906, N101);
xor XOR2 (N915, N896, N893);
xor XOR2 (N916, N914, N485);
or OR2 (N917, N911, N385);
nand NAND4 (N918, N913, N538, N804, N693);
and AND4 (N919, N917, N658, N780, N808);
or OR4 (N920, N908, N519, N225, N365);
buf BUF1 (N921, N880);
buf BUF1 (N922, N916);
xor XOR2 (N923, N919, N808);
and AND2 (N924, N909, N288);
buf BUF1 (N925, N923);
or OR4 (N926, N925, N12, N323, N340);
not NOT1 (N927, N924);
or OR2 (N928, N915, N213);
or OR3 (N929, N926, N321, N168);
or OR3 (N930, N912, N454, N569);
nor NOR2 (N931, N930, N180);
not NOT1 (N932, N927);
nand NAND4 (N933, N888, N832, N822, N354);
buf BUF1 (N934, N922);
or OR3 (N935, N932, N466, N753);
nand NAND2 (N936, N918, N548);
not NOT1 (N937, N934);
buf BUF1 (N938, N933);
or OR3 (N939, N929, N254, N16);
or OR4 (N940, N904, N172, N19, N332);
not NOT1 (N941, N939);
nand NAND4 (N942, N935, N216, N534, N415);
not NOT1 (N943, N937);
nand NAND2 (N944, N921, N428);
nand NAND4 (N945, N920, N130, N775, N815);
not NOT1 (N946, N943);
and AND2 (N947, N931, N121);
nand NAND3 (N948, N928, N765, N68);
or OR2 (N949, N946, N568);
or OR4 (N950, N936, N63, N28, N628);
not NOT1 (N951, N938);
buf BUF1 (N952, N948);
and AND4 (N953, N942, N438, N434, N734);
xor XOR2 (N954, N953, N936);
nand NAND2 (N955, N951, N595);
not NOT1 (N956, N947);
nor NOR2 (N957, N941, N857);
xor XOR2 (N958, N944, N167);
xor XOR2 (N959, N955, N48);
nand NAND3 (N960, N950, N771, N921);
not NOT1 (N961, N960);
xor XOR2 (N962, N956, N780);
nor NOR2 (N963, N962, N215);
not NOT1 (N964, N940);
or OR2 (N965, N949, N836);
nand NAND2 (N966, N957, N130);
or OR3 (N967, N963, N572, N715);
nor NOR3 (N968, N961, N90, N823);
not NOT1 (N969, N968);
and AND3 (N970, N965, N637, N250);
not NOT1 (N971, N970);
not NOT1 (N972, N954);
not NOT1 (N973, N945);
nor NOR4 (N974, N952, N743, N23, N114);
buf BUF1 (N975, N972);
nand NAND3 (N976, N967, N877, N779);
and AND4 (N977, N959, N483, N707, N935);
nor NOR2 (N978, N974, N477);
nor NOR4 (N979, N976, N69, N596, N875);
xor XOR2 (N980, N969, N643);
nor NOR2 (N981, N958, N800);
and AND4 (N982, N980, N91, N539, N670);
xor XOR2 (N983, N982, N153);
buf BUF1 (N984, N966);
and AND2 (N985, N978, N754);
not NOT1 (N986, N981);
or OR3 (N987, N973, N643, N379);
xor XOR2 (N988, N985, N727);
not NOT1 (N989, N984);
buf BUF1 (N990, N986);
xor XOR2 (N991, N987, N187);
buf BUF1 (N992, N979);
nand NAND3 (N993, N983, N79, N242);
nor NOR4 (N994, N964, N938, N963, N391);
not NOT1 (N995, N989);
nand NAND4 (N996, N988, N651, N728, N446);
nand NAND2 (N997, N993, N817);
nor NOR2 (N998, N991, N786);
not NOT1 (N999, N995);
nand NAND2 (N1000, N994, N265);
not NOT1 (N1001, N992);
buf BUF1 (N1002, N998);
or OR2 (N1003, N977, N480);
not NOT1 (N1004, N997);
buf BUF1 (N1005, N971);
or OR3 (N1006, N999, N933, N488);
nand NAND2 (N1007, N1005, N547);
and AND2 (N1008, N1000, N814);
not NOT1 (N1009, N1008);
xor XOR2 (N1010, N1009, N968);
and AND3 (N1011, N1010, N719, N383);
nor NOR3 (N1012, N1004, N487, N584);
nand NAND4 (N1013, N1001, N511, N231, N154);
not NOT1 (N1014, N1011);
buf BUF1 (N1015, N1013);
or OR4 (N1016, N990, N393, N619, N242);
and AND2 (N1017, N1007, N248);
and AND2 (N1018, N975, N609);
nor NOR3 (N1019, N1002, N129, N626);
or OR4 (N1020, N1015, N247, N506, N127);
nor NOR2 (N1021, N1018, N484);
nor NOR2 (N1022, N1014, N130);
xor XOR2 (N1023, N1016, N321);
or OR3 (N1024, N1022, N633, N752);
or OR4 (N1025, N1024, N678, N612, N945);
and AND4 (N1026, N1021, N87, N955, N75);
nand NAND2 (N1027, N1026, N993);
not NOT1 (N1028, N1027);
not NOT1 (N1029, N1023);
not NOT1 (N1030, N1025);
nor NOR4 (N1031, N1030, N688, N538, N471);
xor XOR2 (N1032, N1017, N997);
or OR4 (N1033, N1029, N442, N240, N249);
nand NAND4 (N1034, N1028, N911, N211, N387);
xor XOR2 (N1035, N1020, N766);
not NOT1 (N1036, N1034);
or OR4 (N1037, N1032, N995, N516, N8);
nand NAND2 (N1038, N1031, N991);
and AND2 (N1039, N1006, N605);
not NOT1 (N1040, N1038);
xor XOR2 (N1041, N1033, N839);
buf BUF1 (N1042, N1037);
xor XOR2 (N1043, N1040, N984);
not NOT1 (N1044, N1039);
and AND2 (N1045, N1042, N764);
nand NAND3 (N1046, N1045, N242, N564);
and AND2 (N1047, N1012, N785);
not NOT1 (N1048, N1019);
buf BUF1 (N1049, N1044);
or OR3 (N1050, N1047, N388, N742);
buf BUF1 (N1051, N1049);
and AND2 (N1052, N1035, N797);
xor XOR2 (N1053, N1041, N359);
nor NOR4 (N1054, N1051, N219, N299, N746);
buf BUF1 (N1055, N1050);
xor XOR2 (N1056, N996, N380);
xor XOR2 (N1057, N1036, N831);
xor XOR2 (N1058, N1054, N462);
not NOT1 (N1059, N1043);
nor NOR3 (N1060, N1055, N721, N833);
xor XOR2 (N1061, N1046, N924);
and AND4 (N1062, N1061, N927, N912, N400);
and AND4 (N1063, N1058, N460, N58, N613);
nand NAND3 (N1064, N1063, N9, N77);
and AND3 (N1065, N1062, N496, N35);
buf BUF1 (N1066, N1060);
or OR4 (N1067, N1057, N1021, N354, N65);
and AND2 (N1068, N1064, N293);
not NOT1 (N1069, N1059);
buf BUF1 (N1070, N1052);
xor XOR2 (N1071, N1069, N410);
buf BUF1 (N1072, N1070);
xor XOR2 (N1073, N1071, N977);
xor XOR2 (N1074, N1056, N915);
nor NOR3 (N1075, N1053, N357, N146);
not NOT1 (N1076, N1065);
or OR2 (N1077, N1067, N172);
or OR2 (N1078, N1073, N964);
nor NOR2 (N1079, N1072, N957);
buf BUF1 (N1080, N1075);
buf BUF1 (N1081, N1080);
or OR3 (N1082, N1081, N211, N608);
not NOT1 (N1083, N1077);
buf BUF1 (N1084, N1079);
nand NAND2 (N1085, N1082, N412);
nand NAND3 (N1086, N1076, N699, N176);
not NOT1 (N1087, N1048);
nor NOR3 (N1088, N1085, N911, N542);
buf BUF1 (N1089, N1068);
xor XOR2 (N1090, N1088, N445);
or OR2 (N1091, N1087, N894);
or OR3 (N1092, N1084, N944, N887);
or OR4 (N1093, N1086, N487, N13, N81);
nor NOR4 (N1094, N1089, N15, N243, N1047);
not NOT1 (N1095, N1090);
or OR3 (N1096, N1094, N595, N333);
xor XOR2 (N1097, N1078, N277);
buf BUF1 (N1098, N1091);
not NOT1 (N1099, N1083);
nand NAND2 (N1100, N1066, N586);
and AND2 (N1101, N1074, N588);
not NOT1 (N1102, N1099);
and AND3 (N1103, N1097, N647, N704);
or OR3 (N1104, N1096, N46, N717);
and AND3 (N1105, N1095, N753, N1098);
xor XOR2 (N1106, N347, N460);
nor NOR4 (N1107, N1104, N1047, N25, N968);
nand NAND2 (N1108, N1105, N764);
buf BUF1 (N1109, N1100);
nand NAND3 (N1110, N1101, N636, N172);
not NOT1 (N1111, N1107);
or OR3 (N1112, N1103, N264, N80);
xor XOR2 (N1113, N1109, N408);
buf BUF1 (N1114, N1102);
not NOT1 (N1115, N1003);
buf BUF1 (N1116, N1108);
buf BUF1 (N1117, N1113);
buf BUF1 (N1118, N1111);
nor NOR2 (N1119, N1117, N1007);
xor XOR2 (N1120, N1106, N86);
or OR3 (N1121, N1112, N1028, N314);
and AND3 (N1122, N1116, N1025, N985);
xor XOR2 (N1123, N1119, N178);
xor XOR2 (N1124, N1122, N463);
nand NAND4 (N1125, N1093, N40, N76, N892);
not NOT1 (N1126, N1120);
and AND2 (N1127, N1115, N132);
buf BUF1 (N1128, N1127);
nor NOR3 (N1129, N1092, N341, N542);
nand NAND4 (N1130, N1129, N118, N51, N212);
nor NOR2 (N1131, N1123, N944);
not NOT1 (N1132, N1121);
buf BUF1 (N1133, N1126);
nand NAND2 (N1134, N1130, N378);
nand NAND4 (N1135, N1133, N557, N752, N1012);
or OR3 (N1136, N1134, N257, N480);
nor NOR4 (N1137, N1124, N856, N127, N1018);
not NOT1 (N1138, N1135);
and AND2 (N1139, N1110, N148);
nor NOR4 (N1140, N1114, N295, N697, N547);
nor NOR3 (N1141, N1128, N43, N161);
or OR4 (N1142, N1132, N599, N764, N179);
or OR4 (N1143, N1137, N810, N1100, N357);
buf BUF1 (N1144, N1118);
nand NAND4 (N1145, N1136, N917, N710, N1091);
or OR4 (N1146, N1143, N563, N114, N1125);
not NOT1 (N1147, N186);
not NOT1 (N1148, N1141);
nand NAND3 (N1149, N1144, N765, N1064);
buf BUF1 (N1150, N1145);
or OR3 (N1151, N1146, N859, N398);
xor XOR2 (N1152, N1151, N1094);
nand NAND2 (N1153, N1138, N984);
buf BUF1 (N1154, N1150);
not NOT1 (N1155, N1154);
or OR2 (N1156, N1140, N296);
buf BUF1 (N1157, N1149);
nor NOR2 (N1158, N1152, N244);
xor XOR2 (N1159, N1158, N547);
buf BUF1 (N1160, N1157);
nor NOR2 (N1161, N1153, N864);
not NOT1 (N1162, N1139);
xor XOR2 (N1163, N1155, N216);
nand NAND2 (N1164, N1162, N778);
nand NAND3 (N1165, N1164, N956, N1106);
not NOT1 (N1166, N1161);
or OR3 (N1167, N1165, N191, N847);
xor XOR2 (N1168, N1163, N1162);
buf BUF1 (N1169, N1168);
or OR4 (N1170, N1142, N794, N530, N1129);
xor XOR2 (N1171, N1160, N81);
nor NOR2 (N1172, N1166, N529);
and AND2 (N1173, N1170, N338);
and AND4 (N1174, N1148, N283, N71, N1014);
or OR3 (N1175, N1169, N255, N1052);
or OR4 (N1176, N1159, N54, N974, N703);
not NOT1 (N1177, N1167);
xor XOR2 (N1178, N1171, N974);
and AND3 (N1179, N1174, N759, N303);
nor NOR2 (N1180, N1178, N142);
nand NAND2 (N1181, N1173, N934);
xor XOR2 (N1182, N1175, N621);
nor NOR4 (N1183, N1182, N811, N918, N1133);
xor XOR2 (N1184, N1172, N595);
nor NOR4 (N1185, N1181, N50, N503, N1077);
xor XOR2 (N1186, N1156, N690);
nand NAND4 (N1187, N1147, N234, N569, N1075);
buf BUF1 (N1188, N1183);
nor NOR2 (N1189, N1131, N115);
nor NOR4 (N1190, N1189, N785, N643, N573);
or OR4 (N1191, N1177, N392, N891, N1154);
xor XOR2 (N1192, N1190, N1107);
xor XOR2 (N1193, N1191, N683);
not NOT1 (N1194, N1185);
not NOT1 (N1195, N1187);
xor XOR2 (N1196, N1195, N859);
nor NOR3 (N1197, N1186, N896, N10);
nor NOR4 (N1198, N1180, N296, N101, N58);
not NOT1 (N1199, N1197);
and AND3 (N1200, N1198, N593, N532);
xor XOR2 (N1201, N1196, N1043);
and AND3 (N1202, N1199, N235, N382);
or OR4 (N1203, N1176, N549, N815, N121);
xor XOR2 (N1204, N1193, N717);
xor XOR2 (N1205, N1179, N221);
xor XOR2 (N1206, N1184, N879);
not NOT1 (N1207, N1206);
nand NAND4 (N1208, N1207, N254, N174, N1071);
or OR3 (N1209, N1192, N630, N901);
or OR4 (N1210, N1209, N121, N45, N232);
nor NOR4 (N1211, N1194, N1184, N215, N1178);
not NOT1 (N1212, N1201);
xor XOR2 (N1213, N1204, N25);
buf BUF1 (N1214, N1210);
not NOT1 (N1215, N1208);
buf BUF1 (N1216, N1202);
nor NOR2 (N1217, N1200, N128);
and AND3 (N1218, N1216, N871, N1163);
xor XOR2 (N1219, N1215, N352);
xor XOR2 (N1220, N1214, N1209);
xor XOR2 (N1221, N1211, N1008);
nand NAND4 (N1222, N1205, N907, N686, N572);
not NOT1 (N1223, N1188);
not NOT1 (N1224, N1213);
nor NOR2 (N1225, N1223, N966);
xor XOR2 (N1226, N1222, N462);
and AND4 (N1227, N1220, N417, N422, N347);
buf BUF1 (N1228, N1226);
xor XOR2 (N1229, N1218, N1159);
nand NAND4 (N1230, N1203, N1061, N281, N644);
and AND3 (N1231, N1219, N1003, N574);
nor NOR3 (N1232, N1229, N519, N90);
or OR3 (N1233, N1228, N144, N1113);
xor XOR2 (N1234, N1232, N27);
nand NAND2 (N1235, N1227, N1124);
nor NOR3 (N1236, N1224, N1080, N613);
buf BUF1 (N1237, N1230);
or OR4 (N1238, N1234, N21, N225, N749);
nor NOR3 (N1239, N1231, N80, N959);
buf BUF1 (N1240, N1236);
xor XOR2 (N1241, N1212, N415);
xor XOR2 (N1242, N1241, N667);
buf BUF1 (N1243, N1233);
not NOT1 (N1244, N1235);
nand NAND2 (N1245, N1242, N1007);
and AND2 (N1246, N1244, N1154);
or OR2 (N1247, N1245, N1026);
and AND3 (N1248, N1225, N280, N1236);
buf BUF1 (N1249, N1246);
xor XOR2 (N1250, N1238, N191);
and AND2 (N1251, N1217, N593);
or OR2 (N1252, N1221, N967);
nor NOR2 (N1253, N1247, N1056);
not NOT1 (N1254, N1253);
nand NAND4 (N1255, N1243, N1179, N237, N56);
and AND2 (N1256, N1249, N129);
not NOT1 (N1257, N1239);
xor XOR2 (N1258, N1254, N6);
not NOT1 (N1259, N1240);
not NOT1 (N1260, N1258);
nand NAND3 (N1261, N1237, N730, N874);
not NOT1 (N1262, N1248);
and AND2 (N1263, N1256, N837);
buf BUF1 (N1264, N1252);
or OR3 (N1265, N1259, N359, N993);
or OR3 (N1266, N1264, N122, N882);
nand NAND2 (N1267, N1265, N1013);
buf BUF1 (N1268, N1255);
nor NOR4 (N1269, N1260, N1132, N492, N436);
xor XOR2 (N1270, N1262, N773);
not NOT1 (N1271, N1266);
or OR3 (N1272, N1271, N1176, N806);
xor XOR2 (N1273, N1269, N569);
xor XOR2 (N1274, N1270, N1125);
not NOT1 (N1275, N1267);
not NOT1 (N1276, N1268);
nor NOR2 (N1277, N1275, N861);
xor XOR2 (N1278, N1273, N43);
xor XOR2 (N1279, N1274, N666);
not NOT1 (N1280, N1263);
or OR2 (N1281, N1261, N766);
nor NOR4 (N1282, N1250, N626, N1134, N96);
nand NAND2 (N1283, N1279, N224);
not NOT1 (N1284, N1283);
nor NOR2 (N1285, N1272, N342);
nand NAND2 (N1286, N1257, N752);
xor XOR2 (N1287, N1281, N119);
nand NAND3 (N1288, N1278, N695, N1035);
nand NAND3 (N1289, N1280, N1228, N381);
or OR3 (N1290, N1276, N832, N51);
nand NAND4 (N1291, N1286, N204, N374, N812);
nand NAND2 (N1292, N1285, N323);
and AND4 (N1293, N1251, N137, N488, N1099);
and AND2 (N1294, N1291, N225);
and AND3 (N1295, N1293, N774, N1222);
not NOT1 (N1296, N1282);
nand NAND4 (N1297, N1294, N1123, N95, N50);
nor NOR2 (N1298, N1284, N1070);
not NOT1 (N1299, N1289);
nor NOR4 (N1300, N1287, N598, N1127, N486);
xor XOR2 (N1301, N1290, N934);
xor XOR2 (N1302, N1300, N1140);
buf BUF1 (N1303, N1277);
buf BUF1 (N1304, N1292);
nor NOR2 (N1305, N1304, N702);
not NOT1 (N1306, N1298);
xor XOR2 (N1307, N1306, N223);
and AND2 (N1308, N1299, N1202);
and AND2 (N1309, N1301, N898);
nor NOR4 (N1310, N1302, N178, N261, N144);
nand NAND3 (N1311, N1307, N685, N250);
buf BUF1 (N1312, N1311);
or OR3 (N1313, N1288, N115, N196);
xor XOR2 (N1314, N1303, N1009);
nor NOR3 (N1315, N1297, N1066, N843);
xor XOR2 (N1316, N1314, N783);
buf BUF1 (N1317, N1315);
or OR2 (N1318, N1316, N31);
buf BUF1 (N1319, N1317);
nor NOR4 (N1320, N1296, N401, N253, N338);
nand NAND3 (N1321, N1319, N1229, N1089);
buf BUF1 (N1322, N1321);
nor NOR4 (N1323, N1295, N517, N1188, N267);
and AND2 (N1324, N1312, N739);
xor XOR2 (N1325, N1322, N765);
and AND3 (N1326, N1320, N593, N748);
xor XOR2 (N1327, N1326, N1002);
buf BUF1 (N1328, N1310);
xor XOR2 (N1329, N1327, N1273);
nand NAND4 (N1330, N1329, N282, N585, N719);
buf BUF1 (N1331, N1309);
and AND3 (N1332, N1324, N758, N918);
and AND2 (N1333, N1318, N1076);
xor XOR2 (N1334, N1323, N952);
nor NOR3 (N1335, N1334, N82, N168);
xor XOR2 (N1336, N1305, N38);
nand NAND3 (N1337, N1330, N374, N327);
and AND3 (N1338, N1332, N700, N1180);
buf BUF1 (N1339, N1336);
nor NOR3 (N1340, N1338, N1004, N296);
or OR3 (N1341, N1325, N265, N1055);
nor NOR3 (N1342, N1340, N290, N295);
and AND4 (N1343, N1313, N716, N257, N1050);
xor XOR2 (N1344, N1331, N583);
nor NOR4 (N1345, N1333, N110, N1192, N726);
or OR4 (N1346, N1345, N199, N187, N1097);
buf BUF1 (N1347, N1342);
xor XOR2 (N1348, N1339, N1018);
or OR4 (N1349, N1348, N846, N711, N427);
nand NAND4 (N1350, N1328, N1190, N817, N789);
not NOT1 (N1351, N1308);
nor NOR3 (N1352, N1337, N354, N846);
and AND4 (N1353, N1352, N1026, N707, N573);
and AND2 (N1354, N1343, N269);
nand NAND3 (N1355, N1346, N1341, N727);
and AND4 (N1356, N778, N197, N339, N84);
nand NAND2 (N1357, N1335, N387);
xor XOR2 (N1358, N1357, N151);
not NOT1 (N1359, N1349);
nand NAND4 (N1360, N1358, N441, N1263, N368);
nor NOR3 (N1361, N1351, N504, N1329);
xor XOR2 (N1362, N1360, N726);
nand NAND4 (N1363, N1344, N329, N478, N195);
nor NOR2 (N1364, N1359, N481);
nor NOR2 (N1365, N1347, N930);
nand NAND2 (N1366, N1362, N1033);
xor XOR2 (N1367, N1363, N628);
or OR3 (N1368, N1366, N1252, N482);
xor XOR2 (N1369, N1368, N989);
xor XOR2 (N1370, N1364, N939);
xor XOR2 (N1371, N1353, N314);
not NOT1 (N1372, N1354);
buf BUF1 (N1373, N1355);
not NOT1 (N1374, N1361);
nand NAND4 (N1375, N1373, N1015, N1076, N248);
nand NAND4 (N1376, N1371, N1260, N641, N147);
and AND3 (N1377, N1356, N690, N557);
and AND2 (N1378, N1370, N403);
nor NOR2 (N1379, N1377, N1100);
or OR4 (N1380, N1378, N915, N1063, N1125);
buf BUF1 (N1381, N1380);
nor NOR4 (N1382, N1375, N834, N189, N1290);
or OR4 (N1383, N1382, N1253, N926, N49);
or OR2 (N1384, N1376, N1105);
buf BUF1 (N1385, N1372);
nor NOR2 (N1386, N1381, N705);
and AND3 (N1387, N1386, N990, N54);
buf BUF1 (N1388, N1369);
buf BUF1 (N1389, N1365);
nor NOR2 (N1390, N1350, N762);
buf BUF1 (N1391, N1389);
nor NOR2 (N1392, N1383, N88);
or OR3 (N1393, N1374, N187, N562);
not NOT1 (N1394, N1392);
and AND3 (N1395, N1390, N836, N501);
or OR4 (N1396, N1384, N528, N797, N178);
buf BUF1 (N1397, N1396);
and AND4 (N1398, N1367, N1342, N957, N1280);
and AND4 (N1399, N1387, N17, N1308, N683);
nand NAND3 (N1400, N1398, N216, N1297);
xor XOR2 (N1401, N1393, N1361);
and AND2 (N1402, N1397, N234);
not NOT1 (N1403, N1394);
not NOT1 (N1404, N1391);
and AND3 (N1405, N1400, N538, N1327);
buf BUF1 (N1406, N1385);
and AND2 (N1407, N1399, N1038);
nor NOR3 (N1408, N1404, N12, N461);
not NOT1 (N1409, N1407);
nand NAND3 (N1410, N1409, N570, N440);
and AND4 (N1411, N1402, N672, N1218, N1254);
nor NOR4 (N1412, N1411, N943, N982, N500);
and AND3 (N1413, N1412, N1347, N1061);
and AND4 (N1414, N1406, N207, N1232, N850);
or OR4 (N1415, N1388, N960, N454, N1221);
nand NAND4 (N1416, N1414, N1071, N1181, N566);
nor NOR3 (N1417, N1395, N553, N1245);
nand NAND3 (N1418, N1415, N1363, N378);
nor NOR3 (N1419, N1417, N1087, N1233);
nor NOR2 (N1420, N1379, N166);
nor NOR3 (N1421, N1418, N456, N868);
and AND2 (N1422, N1401, N114);
buf BUF1 (N1423, N1413);
not NOT1 (N1424, N1420);
xor XOR2 (N1425, N1422, N139);
not NOT1 (N1426, N1408);
or OR4 (N1427, N1416, N583, N1424, N227);
xor XOR2 (N1428, N802, N1054);
nand NAND4 (N1429, N1405, N166, N1189, N926);
nand NAND2 (N1430, N1419, N44);
not NOT1 (N1431, N1428);
xor XOR2 (N1432, N1426, N427);
and AND4 (N1433, N1423, N930, N1036, N1392);
and AND3 (N1434, N1421, N1018, N1401);
or OR4 (N1435, N1431, N732, N970, N30);
nor NOR2 (N1436, N1427, N651);
nor NOR3 (N1437, N1435, N973, N1035);
buf BUF1 (N1438, N1410);
nor NOR2 (N1439, N1434, N1017);
nand NAND4 (N1440, N1433, N613, N465, N268);
nor NOR2 (N1441, N1439, N954);
nand NAND3 (N1442, N1425, N243, N1022);
and AND3 (N1443, N1438, N651, N298);
or OR4 (N1444, N1429, N61, N11, N406);
nor NOR2 (N1445, N1441, N719);
xor XOR2 (N1446, N1437, N1117);
xor XOR2 (N1447, N1446, N148);
not NOT1 (N1448, N1432);
xor XOR2 (N1449, N1444, N1048);
nor NOR4 (N1450, N1442, N506, N515, N89);
nor NOR3 (N1451, N1449, N241, N1158);
not NOT1 (N1452, N1447);
xor XOR2 (N1453, N1430, N502);
xor XOR2 (N1454, N1440, N587);
xor XOR2 (N1455, N1403, N315);
nor NOR2 (N1456, N1451, N364);
nor NOR3 (N1457, N1436, N693, N1366);
or OR2 (N1458, N1454, N260);
and AND4 (N1459, N1450, N5, N1079, N649);
or OR2 (N1460, N1455, N463);
nor NOR4 (N1461, N1453, N514, N456, N44);
and AND3 (N1462, N1459, N621, N556);
not NOT1 (N1463, N1456);
nand NAND4 (N1464, N1460, N1224, N1402, N51);
xor XOR2 (N1465, N1458, N874);
and AND3 (N1466, N1463, N650, N70);
and AND4 (N1467, N1452, N1017, N751, N936);
and AND3 (N1468, N1445, N1064, N1349);
or OR2 (N1469, N1467, N1167);
not NOT1 (N1470, N1462);
nand NAND2 (N1471, N1464, N851);
and AND3 (N1472, N1468, N28, N894);
nand NAND3 (N1473, N1461, N1343, N1376);
buf BUF1 (N1474, N1471);
nand NAND2 (N1475, N1473, N482);
buf BUF1 (N1476, N1448);
xor XOR2 (N1477, N1443, N1472);
xor XOR2 (N1478, N1365, N743);
and AND2 (N1479, N1475, N436);
nor NOR3 (N1480, N1457, N696, N574);
and AND3 (N1481, N1476, N59, N1252);
nor NOR2 (N1482, N1477, N92);
buf BUF1 (N1483, N1480);
not NOT1 (N1484, N1478);
not NOT1 (N1485, N1466);
and AND4 (N1486, N1482, N1013, N765, N1300);
or OR4 (N1487, N1486, N1451, N261, N111);
not NOT1 (N1488, N1484);
and AND2 (N1489, N1469, N1131);
nor NOR4 (N1490, N1489, N919, N1325, N1319);
nand NAND2 (N1491, N1485, N233);
nor NOR2 (N1492, N1474, N93);
nand NAND2 (N1493, N1483, N1342);
buf BUF1 (N1494, N1487);
not NOT1 (N1495, N1491);
buf BUF1 (N1496, N1479);
not NOT1 (N1497, N1494);
and AND3 (N1498, N1470, N700, N1125);
or OR2 (N1499, N1498, N1352);
buf BUF1 (N1500, N1492);
buf BUF1 (N1501, N1495);
or OR2 (N1502, N1497, N160);
nand NAND2 (N1503, N1496, N1419);
not NOT1 (N1504, N1465);
nor NOR4 (N1505, N1501, N939, N1389, N216);
nor NOR3 (N1506, N1499, N735, N1498);
buf BUF1 (N1507, N1490);
buf BUF1 (N1508, N1493);
not NOT1 (N1509, N1505);
or OR3 (N1510, N1503, N186, N1352);
nor NOR3 (N1511, N1509, N531, N1482);
nand NAND4 (N1512, N1508, N379, N1436, N670);
xor XOR2 (N1513, N1500, N1437);
or OR2 (N1514, N1488, N1259);
and AND4 (N1515, N1514, N1074, N1249, N337);
xor XOR2 (N1516, N1511, N1210);
or OR2 (N1517, N1512, N1359);
not NOT1 (N1518, N1513);
xor XOR2 (N1519, N1504, N792);
not NOT1 (N1520, N1518);
nor NOR2 (N1521, N1516, N85);
nor NOR2 (N1522, N1502, N1393);
nor NOR3 (N1523, N1515, N948, N369);
nor NOR2 (N1524, N1510, N412);
or OR3 (N1525, N1521, N1018, N1361);
buf BUF1 (N1526, N1519);
nand NAND4 (N1527, N1523, N310, N765, N1500);
buf BUF1 (N1528, N1506);
or OR4 (N1529, N1520, N1044, N872, N1382);
nor NOR3 (N1530, N1526, N1215, N442);
or OR4 (N1531, N1529, N6, N697, N280);
or OR2 (N1532, N1517, N492);
and AND4 (N1533, N1525, N1119, N1347, N91);
or OR4 (N1534, N1532, N888, N1270, N81);
nand NAND3 (N1535, N1533, N482, N927);
nor NOR4 (N1536, N1524, N188, N924, N786);
or OR4 (N1537, N1536, N1072, N147, N703);
or OR4 (N1538, N1527, N1480, N51, N912);
or OR3 (N1539, N1538, N1247, N235);
xor XOR2 (N1540, N1535, N850);
nand NAND2 (N1541, N1531, N357);
or OR2 (N1542, N1541, N160);
or OR4 (N1543, N1540, N722, N100, N374);
and AND3 (N1544, N1481, N1031, N1260);
or OR4 (N1545, N1534, N1009, N13, N1326);
buf BUF1 (N1546, N1507);
and AND3 (N1547, N1545, N812, N309);
or OR4 (N1548, N1546, N1339, N160, N732);
nand NAND2 (N1549, N1528, N364);
and AND3 (N1550, N1542, N492, N1094);
xor XOR2 (N1551, N1530, N803);
or OR4 (N1552, N1544, N514, N593, N1195);
nand NAND2 (N1553, N1549, N1508);
or OR3 (N1554, N1553, N426, N1255);
and AND3 (N1555, N1551, N1457, N1400);
not NOT1 (N1556, N1543);
or OR3 (N1557, N1537, N1160, N118);
or OR3 (N1558, N1550, N778, N1046);
and AND2 (N1559, N1556, N137);
nand NAND2 (N1560, N1555, N1518);
buf BUF1 (N1561, N1554);
not NOT1 (N1562, N1558);
nand NAND4 (N1563, N1560, N856, N1559, N1060);
nor NOR2 (N1564, N673, N1521);
nor NOR3 (N1565, N1564, N700, N762);
and AND4 (N1566, N1563, N262, N554, N237);
nand NAND2 (N1567, N1561, N801);
and AND4 (N1568, N1566, N1376, N1079, N534);
nor NOR4 (N1569, N1565, N567, N361, N899);
or OR4 (N1570, N1547, N484, N113, N200);
nor NOR3 (N1571, N1562, N848, N66);
nor NOR2 (N1572, N1569, N1055);
nor NOR4 (N1573, N1568, N1158, N600, N112);
not NOT1 (N1574, N1567);
not NOT1 (N1575, N1572);
and AND2 (N1576, N1557, N1222);
nand NAND4 (N1577, N1570, N1251, N1520, N706);
buf BUF1 (N1578, N1539);
and AND3 (N1579, N1575, N911, N877);
xor XOR2 (N1580, N1578, N422);
xor XOR2 (N1581, N1577, N465);
nor NOR4 (N1582, N1579, N329, N520, N1468);
nand NAND2 (N1583, N1580, N1104);
nand NAND3 (N1584, N1583, N352, N1427);
nor NOR2 (N1585, N1574, N481);
and AND4 (N1586, N1573, N1157, N68, N1519);
nand NAND3 (N1587, N1548, N1318, N520);
buf BUF1 (N1588, N1587);
or OR3 (N1589, N1552, N590, N1356);
xor XOR2 (N1590, N1576, N898);
not NOT1 (N1591, N1590);
not NOT1 (N1592, N1571);
xor XOR2 (N1593, N1522, N344);
and AND3 (N1594, N1591, N345, N163);
or OR2 (N1595, N1592, N873);
xor XOR2 (N1596, N1582, N722);
not NOT1 (N1597, N1594);
or OR3 (N1598, N1581, N1269, N545);
buf BUF1 (N1599, N1585);
or OR2 (N1600, N1589, N841);
or OR2 (N1601, N1596, N581);
buf BUF1 (N1602, N1600);
xor XOR2 (N1603, N1599, N1057);
xor XOR2 (N1604, N1598, N1124);
or OR3 (N1605, N1601, N160, N383);
or OR4 (N1606, N1605, N1179, N980, N284);
nand NAND3 (N1607, N1604, N448, N1200);
buf BUF1 (N1608, N1606);
nor NOR2 (N1609, N1595, N1423);
nand NAND2 (N1610, N1597, N517);
nor NOR3 (N1611, N1586, N515, N1213);
nor NOR2 (N1612, N1609, N594);
and AND3 (N1613, N1603, N1430, N292);
nor NOR2 (N1614, N1607, N1393);
nor NOR3 (N1615, N1610, N1373, N707);
not NOT1 (N1616, N1584);
not NOT1 (N1617, N1616);
xor XOR2 (N1618, N1612, N980);
xor XOR2 (N1619, N1615, N1013);
nor NOR3 (N1620, N1602, N1070, N692);
nand NAND4 (N1621, N1593, N871, N1178, N221);
and AND3 (N1622, N1619, N708, N617);
xor XOR2 (N1623, N1621, N1564);
nor NOR2 (N1624, N1588, N1421);
not NOT1 (N1625, N1611);
nor NOR4 (N1626, N1624, N179, N1075, N1418);
not NOT1 (N1627, N1608);
and AND4 (N1628, N1614, N757, N1518, N1241);
buf BUF1 (N1629, N1628);
and AND3 (N1630, N1613, N315, N1478);
nor NOR4 (N1631, N1626, N641, N1622, N91);
buf BUF1 (N1632, N429);
or OR4 (N1633, N1629, N958, N514, N1099);
nor NOR2 (N1634, N1623, N601);
xor XOR2 (N1635, N1625, N1431);
xor XOR2 (N1636, N1634, N140);
nand NAND2 (N1637, N1633, N1271);
nand NAND2 (N1638, N1637, N1556);
nor NOR2 (N1639, N1618, N1316);
buf BUF1 (N1640, N1639);
nor NOR3 (N1641, N1630, N1392, N71);
and AND3 (N1642, N1635, N277, N427);
not NOT1 (N1643, N1638);
nor NOR2 (N1644, N1642, N937);
not NOT1 (N1645, N1640);
nor NOR2 (N1646, N1617, N91);
buf BUF1 (N1647, N1644);
buf BUF1 (N1648, N1636);
nor NOR2 (N1649, N1641, N449);
buf BUF1 (N1650, N1631);
xor XOR2 (N1651, N1647, N1078);
and AND3 (N1652, N1643, N322, N814);
xor XOR2 (N1653, N1645, N117);
nand NAND4 (N1654, N1652, N364, N626, N345);
and AND4 (N1655, N1632, N528, N1012, N1163);
not NOT1 (N1656, N1620);
and AND4 (N1657, N1655, N1503, N1318, N822);
and AND4 (N1658, N1656, N404, N800, N605);
nand NAND3 (N1659, N1646, N1658, N238);
xor XOR2 (N1660, N445, N301);
buf BUF1 (N1661, N1654);
nand NAND4 (N1662, N1649, N741, N1488, N266);
nand NAND4 (N1663, N1648, N1405, N1582, N533);
or OR3 (N1664, N1662, N610, N341);
or OR3 (N1665, N1627, N1563, N1607);
xor XOR2 (N1666, N1659, N1228);
and AND4 (N1667, N1661, N837, N1118, N865);
xor XOR2 (N1668, N1657, N1081);
not NOT1 (N1669, N1653);
or OR3 (N1670, N1669, N1195, N404);
buf BUF1 (N1671, N1660);
buf BUF1 (N1672, N1666);
nand NAND2 (N1673, N1650, N782);
not NOT1 (N1674, N1651);
nor NOR4 (N1675, N1665, N1529, N1307, N407);
not NOT1 (N1676, N1664);
not NOT1 (N1677, N1674);
and AND3 (N1678, N1671, N1408, N654);
nor NOR3 (N1679, N1673, N469, N810);
or OR4 (N1680, N1668, N938, N1490, N1304);
or OR2 (N1681, N1675, N246);
not NOT1 (N1682, N1679);
xor XOR2 (N1683, N1680, N484);
nand NAND3 (N1684, N1670, N161, N952);
buf BUF1 (N1685, N1667);
and AND4 (N1686, N1681, N586, N244, N1249);
buf BUF1 (N1687, N1686);
nand NAND2 (N1688, N1676, N552);
xor XOR2 (N1689, N1682, N1687);
nor NOR3 (N1690, N443, N988, N711);
and AND3 (N1691, N1683, N348, N17);
or OR3 (N1692, N1691, N835, N10);
nor NOR2 (N1693, N1690, N783);
nor NOR3 (N1694, N1693, N656, N131);
and AND2 (N1695, N1689, N1446);
nor NOR4 (N1696, N1688, N479, N369, N104);
nor NOR3 (N1697, N1696, N1597, N89);
nand NAND3 (N1698, N1672, N353, N830);
nor NOR4 (N1699, N1692, N961, N1190, N189);
or OR4 (N1700, N1694, N1481, N22, N1556);
not NOT1 (N1701, N1700);
not NOT1 (N1702, N1677);
or OR2 (N1703, N1695, N1551);
xor XOR2 (N1704, N1702, N786);
not NOT1 (N1705, N1698);
or OR4 (N1706, N1685, N947, N767, N1514);
not NOT1 (N1707, N1704);
or OR2 (N1708, N1678, N827);
not NOT1 (N1709, N1705);
nor NOR4 (N1710, N1707, N301, N1406, N590);
or OR2 (N1711, N1684, N770);
nand NAND3 (N1712, N1699, N190, N1192);
xor XOR2 (N1713, N1703, N1567);
and AND2 (N1714, N1708, N359);
buf BUF1 (N1715, N1714);
not NOT1 (N1716, N1697);
xor XOR2 (N1717, N1710, N240);
nand NAND4 (N1718, N1706, N357, N530, N1272);
or OR3 (N1719, N1709, N33, N535);
not NOT1 (N1720, N1719);
nor NOR3 (N1721, N1711, N1581, N370);
not NOT1 (N1722, N1701);
not NOT1 (N1723, N1663);
buf BUF1 (N1724, N1722);
nand NAND3 (N1725, N1716, N51, N1580);
xor XOR2 (N1726, N1712, N285);
buf BUF1 (N1727, N1725);
not NOT1 (N1728, N1723);
nand NAND3 (N1729, N1728, N401, N1060);
or OR2 (N1730, N1727, N188);
not NOT1 (N1731, N1717);
buf BUF1 (N1732, N1721);
xor XOR2 (N1733, N1718, N1246);
nor NOR4 (N1734, N1713, N865, N66, N644);
xor XOR2 (N1735, N1732, N1531);
not NOT1 (N1736, N1731);
not NOT1 (N1737, N1726);
and AND3 (N1738, N1735, N1308, N538);
xor XOR2 (N1739, N1730, N420);
and AND4 (N1740, N1739, N447, N56, N1219);
nor NOR4 (N1741, N1724, N77, N415, N524);
xor XOR2 (N1742, N1720, N805);
and AND3 (N1743, N1738, N592, N1092);
or OR4 (N1744, N1743, N464, N950, N140);
nand NAND2 (N1745, N1736, N1011);
nand NAND4 (N1746, N1715, N1583, N1576, N582);
not NOT1 (N1747, N1734);
not NOT1 (N1748, N1744);
buf BUF1 (N1749, N1746);
nor NOR2 (N1750, N1749, N654);
buf BUF1 (N1751, N1737);
and AND4 (N1752, N1729, N637, N1739, N589);
not NOT1 (N1753, N1751);
xor XOR2 (N1754, N1741, N658);
xor XOR2 (N1755, N1745, N36);
nor NOR2 (N1756, N1747, N1471);
xor XOR2 (N1757, N1733, N366);
nand NAND2 (N1758, N1740, N122);
nand NAND2 (N1759, N1757, N1046);
nor NOR4 (N1760, N1753, N537, N1551, N822);
xor XOR2 (N1761, N1742, N871);
and AND4 (N1762, N1755, N59, N1490, N1191);
buf BUF1 (N1763, N1762);
and AND2 (N1764, N1759, N358);
buf BUF1 (N1765, N1758);
and AND4 (N1766, N1756, N356, N831, N561);
not NOT1 (N1767, N1766);
or OR4 (N1768, N1752, N684, N1723, N1268);
and AND3 (N1769, N1768, N1018, N1549);
or OR3 (N1770, N1765, N909, N211);
and AND3 (N1771, N1767, N1622, N1437);
nand NAND3 (N1772, N1769, N1556, N169);
xor XOR2 (N1773, N1761, N1519);
nor NOR2 (N1774, N1764, N1674);
nor NOR2 (N1775, N1748, N1746);
not NOT1 (N1776, N1774);
nor NOR4 (N1777, N1772, N1195, N1415, N1569);
not NOT1 (N1778, N1760);
nor NOR3 (N1779, N1750, N373, N908);
or OR4 (N1780, N1754, N1614, N287, N27);
buf BUF1 (N1781, N1780);
not NOT1 (N1782, N1779);
nand NAND3 (N1783, N1763, N670, N1056);
buf BUF1 (N1784, N1783);
and AND2 (N1785, N1781, N1224);
buf BUF1 (N1786, N1771);
xor XOR2 (N1787, N1786, N959);
and AND2 (N1788, N1784, N347);
or OR4 (N1789, N1787, N621, N768, N581);
nor NOR2 (N1790, N1778, N988);
xor XOR2 (N1791, N1785, N1596);
nand NAND2 (N1792, N1770, N1170);
nor NOR2 (N1793, N1782, N1521);
buf BUF1 (N1794, N1773);
buf BUF1 (N1795, N1776);
nand NAND2 (N1796, N1795, N1486);
xor XOR2 (N1797, N1788, N178);
buf BUF1 (N1798, N1793);
or OR4 (N1799, N1794, N980, N407, N1044);
nor NOR3 (N1800, N1790, N202, N926);
and AND3 (N1801, N1775, N951, N1377);
nand NAND2 (N1802, N1799, N62);
and AND3 (N1803, N1777, N438, N1632);
buf BUF1 (N1804, N1789);
nor NOR2 (N1805, N1802, N167);
not NOT1 (N1806, N1804);
nand NAND2 (N1807, N1797, N1034);
not NOT1 (N1808, N1792);
not NOT1 (N1809, N1803);
nand NAND2 (N1810, N1801, N213);
nand NAND3 (N1811, N1805, N425, N1333);
not NOT1 (N1812, N1800);
xor XOR2 (N1813, N1809, N201);
xor XOR2 (N1814, N1808, N1190);
xor XOR2 (N1815, N1798, N1775);
or OR4 (N1816, N1811, N1366, N743, N1715);
buf BUF1 (N1817, N1791);
nand NAND2 (N1818, N1815, N580);
xor XOR2 (N1819, N1816, N773);
or OR2 (N1820, N1814, N1732);
nor NOR2 (N1821, N1819, N1656);
or OR4 (N1822, N1796, N145, N1190, N505);
nor NOR2 (N1823, N1813, N326);
nor NOR4 (N1824, N1812, N890, N1395, N697);
and AND4 (N1825, N1818, N200, N529, N350);
nor NOR3 (N1826, N1824, N12, N914);
and AND4 (N1827, N1823, N1651, N1378, N558);
not NOT1 (N1828, N1825);
nand NAND3 (N1829, N1820, N1522, N1790);
xor XOR2 (N1830, N1817, N649);
or OR2 (N1831, N1821, N183);
or OR3 (N1832, N1828, N1583, N228);
buf BUF1 (N1833, N1830);
buf BUF1 (N1834, N1826);
not NOT1 (N1835, N1833);
xor XOR2 (N1836, N1807, N1085);
buf BUF1 (N1837, N1822);
buf BUF1 (N1838, N1806);
nor NOR3 (N1839, N1835, N502, N1423);
buf BUF1 (N1840, N1829);
nand NAND4 (N1841, N1831, N1227, N1552, N70);
and AND4 (N1842, N1836, N703, N1649, N771);
buf BUF1 (N1843, N1842);
and AND3 (N1844, N1841, N489, N683);
or OR2 (N1845, N1838, N819);
and AND3 (N1846, N1832, N993, N556);
nand NAND4 (N1847, N1843, N1584, N775, N1617);
nand NAND2 (N1848, N1837, N511);
xor XOR2 (N1849, N1846, N25);
nor NOR4 (N1850, N1840, N527, N1328, N847);
nor NOR3 (N1851, N1845, N700, N1414);
and AND4 (N1852, N1839, N560, N1395, N202);
nor NOR4 (N1853, N1827, N1800, N1621, N1230);
not NOT1 (N1854, N1848);
xor XOR2 (N1855, N1850, N588);
buf BUF1 (N1856, N1847);
xor XOR2 (N1857, N1852, N1395);
nand NAND3 (N1858, N1849, N798, N1562);
not NOT1 (N1859, N1858);
nand NAND4 (N1860, N1854, N383, N1090, N845);
and AND3 (N1861, N1859, N276, N309);
xor XOR2 (N1862, N1851, N1311);
nor NOR2 (N1863, N1810, N1181);
buf BUF1 (N1864, N1844);
buf BUF1 (N1865, N1860);
nand NAND4 (N1866, N1853, N971, N474, N1763);
xor XOR2 (N1867, N1864, N269);
or OR3 (N1868, N1834, N1614, N1236);
and AND2 (N1869, N1867, N1737);
nor NOR2 (N1870, N1868, N124);
xor XOR2 (N1871, N1861, N1280);
and AND3 (N1872, N1862, N116, N1692);
nor NOR4 (N1873, N1872, N1805, N905, N1379);
nand NAND3 (N1874, N1869, N1391, N996);
xor XOR2 (N1875, N1856, N1577);
buf BUF1 (N1876, N1875);
or OR2 (N1877, N1871, N1685);
not NOT1 (N1878, N1866);
nand NAND3 (N1879, N1876, N639, N587);
xor XOR2 (N1880, N1870, N531);
buf BUF1 (N1881, N1878);
or OR2 (N1882, N1877, N635);
nand NAND4 (N1883, N1881, N566, N260, N1343);
nor NOR2 (N1884, N1865, N403);
and AND4 (N1885, N1863, N1350, N1482, N1088);
buf BUF1 (N1886, N1874);
and AND3 (N1887, N1885, N1876, N64);
xor XOR2 (N1888, N1855, N123);
nand NAND2 (N1889, N1882, N56);
nand NAND2 (N1890, N1883, N1);
not NOT1 (N1891, N1889);
xor XOR2 (N1892, N1886, N1068);
xor XOR2 (N1893, N1884, N1451);
and AND3 (N1894, N1892, N1312, N912);
nand NAND3 (N1895, N1880, N1797, N818);
nor NOR4 (N1896, N1887, N1048, N1720, N1);
buf BUF1 (N1897, N1896);
xor XOR2 (N1898, N1888, N996);
nand NAND4 (N1899, N1873, N867, N1375, N1292);
nand NAND4 (N1900, N1899, N741, N743, N1783);
and AND4 (N1901, N1897, N1104, N1732, N1687);
xor XOR2 (N1902, N1891, N47);
nor NOR2 (N1903, N1857, N249);
nand NAND4 (N1904, N1879, N1319, N1622, N1585);
and AND4 (N1905, N1903, N1651, N1450, N479);
and AND2 (N1906, N1902, N1790);
nor NOR3 (N1907, N1894, N1393, N164);
buf BUF1 (N1908, N1907);
not NOT1 (N1909, N1906);
not NOT1 (N1910, N1904);
and AND4 (N1911, N1901, N1246, N623, N692);
and AND3 (N1912, N1900, N171, N1034);
nor NOR4 (N1913, N1893, N474, N1693, N1671);
buf BUF1 (N1914, N1913);
or OR2 (N1915, N1905, N87);
nand NAND2 (N1916, N1914, N1873);
xor XOR2 (N1917, N1912, N557);
nand NAND2 (N1918, N1917, N760);
nor NOR4 (N1919, N1911, N72, N438, N1776);
buf BUF1 (N1920, N1919);
and AND4 (N1921, N1908, N665, N749, N1452);
xor XOR2 (N1922, N1910, N1046);
nand NAND4 (N1923, N1898, N1175, N138, N1273);
nand NAND3 (N1924, N1916, N80, N1811);
not NOT1 (N1925, N1915);
and AND3 (N1926, N1924, N1099, N1472);
nand NAND2 (N1927, N1920, N1034);
buf BUF1 (N1928, N1926);
or OR2 (N1929, N1890, N1315);
not NOT1 (N1930, N1922);
xor XOR2 (N1931, N1895, N1141);
and AND3 (N1932, N1909, N1621, N986);
xor XOR2 (N1933, N1925, N282);
nand NAND2 (N1934, N1932, N1697);
buf BUF1 (N1935, N1931);
buf BUF1 (N1936, N1933);
buf BUF1 (N1937, N1936);
and AND2 (N1938, N1930, N428);
or OR4 (N1939, N1929, N1659, N1570, N1757);
buf BUF1 (N1940, N1939);
nand NAND2 (N1941, N1923, N99);
buf BUF1 (N1942, N1941);
and AND3 (N1943, N1937, N1248, N700);
nand NAND3 (N1944, N1934, N599, N115);
nand NAND2 (N1945, N1944, N764);
nor NOR3 (N1946, N1928, N1565, N1274);
not NOT1 (N1947, N1940);
and AND4 (N1948, N1938, N958, N533, N1043);
or OR4 (N1949, N1946, N1149, N610, N355);
and AND3 (N1950, N1918, N1002, N111);
nand NAND2 (N1951, N1948, N1605);
xor XOR2 (N1952, N1945, N1353);
nor NOR4 (N1953, N1951, N1647, N570, N1811);
not NOT1 (N1954, N1953);
buf BUF1 (N1955, N1935);
buf BUF1 (N1956, N1921);
or OR3 (N1957, N1927, N1335, N607);
and AND4 (N1958, N1956, N21, N80, N661);
xor XOR2 (N1959, N1958, N1402);
xor XOR2 (N1960, N1950, N1481);
not NOT1 (N1961, N1955);
buf BUF1 (N1962, N1952);
or OR4 (N1963, N1943, N1742, N201, N1561);
xor XOR2 (N1964, N1961, N1885);
xor XOR2 (N1965, N1963, N1860);
xor XOR2 (N1966, N1954, N721);
nand NAND4 (N1967, N1966, N479, N458, N665);
buf BUF1 (N1968, N1947);
nor NOR4 (N1969, N1965, N1378, N632, N517);
nand NAND2 (N1970, N1959, N1225);
and AND2 (N1971, N1957, N809);
buf BUF1 (N1972, N1964);
xor XOR2 (N1973, N1967, N1748);
and AND4 (N1974, N1970, N644, N1594, N792);
and AND4 (N1975, N1962, N1947, N1064, N958);
not NOT1 (N1976, N1942);
xor XOR2 (N1977, N1971, N1949);
buf BUF1 (N1978, N1258);
nor NOR4 (N1979, N1977, N1354, N901, N1347);
nor NOR4 (N1980, N1978, N1810, N977, N11);
nand NAND4 (N1981, N1980, N340, N55, N387);
or OR4 (N1982, N1973, N65, N1103, N1341);
nor NOR3 (N1983, N1974, N1333, N819);
not NOT1 (N1984, N1969);
xor XOR2 (N1985, N1976, N1964);
and AND4 (N1986, N1982, N1654, N320, N503);
buf BUF1 (N1987, N1968);
and AND2 (N1988, N1986, N732);
nor NOR2 (N1989, N1988, N852);
not NOT1 (N1990, N1983);
not NOT1 (N1991, N1984);
not NOT1 (N1992, N1981);
buf BUF1 (N1993, N1985);
xor XOR2 (N1994, N1989, N1725);
not NOT1 (N1995, N1994);
or OR3 (N1996, N1993, N1646, N1781);
or OR2 (N1997, N1991, N1205);
and AND4 (N1998, N1979, N456, N1612, N344);
nand NAND3 (N1999, N1998, N414, N1510);
nor NOR3 (N2000, N1972, N1246, N46);
nor NOR4 (N2001, N1975, N1474, N149, N1911);
or OR3 (N2002, N2001, N1350, N360);
buf BUF1 (N2003, N2002);
xor XOR2 (N2004, N1995, N1994);
and AND3 (N2005, N1987, N955, N257);
buf BUF1 (N2006, N1999);
or OR4 (N2007, N2006, N1402, N1726, N907);
buf BUF1 (N2008, N2007);
nand NAND4 (N2009, N1960, N161, N729, N225);
xor XOR2 (N2010, N1990, N549);
or OR4 (N2011, N1996, N1901, N1419, N871);
nand NAND2 (N2012, N2004, N128);
buf BUF1 (N2013, N2008);
or OR3 (N2014, N2012, N883, N1735);
and AND3 (N2015, N2009, N1842, N1670);
and AND4 (N2016, N2010, N603, N977, N650);
not NOT1 (N2017, N2013);
xor XOR2 (N2018, N1997, N1689);
xor XOR2 (N2019, N2003, N185);
not NOT1 (N2020, N1992);
nand NAND4 (N2021, N2016, N1838, N636, N1599);
nand NAND3 (N2022, N2015, N1376, N670);
xor XOR2 (N2023, N2005, N607);
nand NAND3 (N2024, N2019, N489, N532);
xor XOR2 (N2025, N2017, N1244);
xor XOR2 (N2026, N2018, N4);
buf BUF1 (N2027, N2000);
and AND2 (N2028, N2023, N1233);
buf BUF1 (N2029, N2014);
nor NOR4 (N2030, N2029, N774, N192, N239);
and AND2 (N2031, N2028, N1956);
not NOT1 (N2032, N2020);
xor XOR2 (N2033, N2021, N264);
buf BUF1 (N2034, N2033);
buf BUF1 (N2035, N2030);
nand NAND4 (N2036, N2011, N1579, N1072, N1054);
or OR4 (N2037, N2035, N35, N1428, N1186);
and AND3 (N2038, N2026, N2023, N676);
or OR2 (N2039, N2024, N200);
or OR3 (N2040, N2022, N1804, N578);
nor NOR3 (N2041, N2039, N210, N1694);
not NOT1 (N2042, N2031);
xor XOR2 (N2043, N2040, N1007);
nor NOR4 (N2044, N2037, N1780, N772, N315);
not NOT1 (N2045, N2036);
nand NAND2 (N2046, N2043, N834);
buf BUF1 (N2047, N2046);
or OR3 (N2048, N2044, N275, N461);
not NOT1 (N2049, N2034);
xor XOR2 (N2050, N2041, N951);
and AND4 (N2051, N2038, N134, N1217, N856);
buf BUF1 (N2052, N2051);
and AND4 (N2053, N2027, N851, N773, N1585);
nor NOR4 (N2054, N2047, N1757, N169, N747);
xor XOR2 (N2055, N2053, N223);
buf BUF1 (N2056, N2055);
not NOT1 (N2057, N2056);
or OR4 (N2058, N2025, N1410, N1754, N30);
and AND2 (N2059, N2058, N83);
nor NOR3 (N2060, N2050, N374, N1694);
nand NAND4 (N2061, N2060, N950, N519, N223);
xor XOR2 (N2062, N2057, N1550);
buf BUF1 (N2063, N2032);
and AND2 (N2064, N2052, N1801);
or OR3 (N2065, N2045, N1390, N1887);
xor XOR2 (N2066, N2062, N938);
xor XOR2 (N2067, N2049, N1790);
nand NAND4 (N2068, N2067, N292, N458, N425);
or OR2 (N2069, N2042, N679);
not NOT1 (N2070, N2048);
and AND2 (N2071, N2054, N1609);
buf BUF1 (N2072, N2059);
nand NAND3 (N2073, N2065, N1282, N1518);
and AND2 (N2074, N2071, N1763);
and AND4 (N2075, N2072, N1042, N1830, N1787);
xor XOR2 (N2076, N2068, N1399);
not NOT1 (N2077, N2075);
or OR4 (N2078, N2069, N912, N170, N924);
not NOT1 (N2079, N2076);
not NOT1 (N2080, N2074);
xor XOR2 (N2081, N2080, N638);
nand NAND2 (N2082, N2081, N142);
xor XOR2 (N2083, N2079, N859);
and AND2 (N2084, N2083, N1416);
or OR3 (N2085, N2061, N625, N228);
and AND2 (N2086, N2070, N1514);
nor NOR2 (N2087, N2063, N1706);
buf BUF1 (N2088, N2077);
nand NAND2 (N2089, N2078, N1203);
buf BUF1 (N2090, N2085);
nand NAND2 (N2091, N2066, N1814);
and AND2 (N2092, N2091, N1762);
not NOT1 (N2093, N2082);
or OR2 (N2094, N2064, N654);
xor XOR2 (N2095, N2089, N245);
not NOT1 (N2096, N2087);
nand NAND4 (N2097, N2086, N1288, N246, N23);
nand NAND4 (N2098, N2090, N808, N182, N709);
not NOT1 (N2099, N2094);
and AND2 (N2100, N2093, N1455);
nand NAND3 (N2101, N2095, N146, N933);
or OR4 (N2102, N2084, N1242, N1982, N647);
nand NAND4 (N2103, N2101, N924, N860, N1459);
nor NOR4 (N2104, N2103, N371, N973, N1407);
xor XOR2 (N2105, N2092, N808);
nor NOR2 (N2106, N2099, N1720);
not NOT1 (N2107, N2096);
not NOT1 (N2108, N2073);
buf BUF1 (N2109, N2102);
and AND4 (N2110, N2107, N1192, N572, N1802);
and AND2 (N2111, N2104, N339);
xor XOR2 (N2112, N2106, N745);
not NOT1 (N2113, N2097);
not NOT1 (N2114, N2113);
buf BUF1 (N2115, N2100);
nor NOR4 (N2116, N2110, N200, N1857, N968);
nand NAND2 (N2117, N2109, N658);
not NOT1 (N2118, N2105);
and AND3 (N2119, N2114, N1980, N47);
not NOT1 (N2120, N2118);
nand NAND4 (N2121, N2117, N1416, N658, N1132);
xor XOR2 (N2122, N2116, N836);
nand NAND2 (N2123, N2120, N320);
not NOT1 (N2124, N2115);
nor NOR3 (N2125, N2119, N1072, N1160);
buf BUF1 (N2126, N2088);
not NOT1 (N2127, N2125);
or OR4 (N2128, N2122, N383, N113, N2102);
or OR3 (N2129, N2127, N1689, N1442);
buf BUF1 (N2130, N2124);
nand NAND4 (N2131, N2123, N1549, N508, N98);
buf BUF1 (N2132, N2131);
nand NAND2 (N2133, N2129, N1346);
buf BUF1 (N2134, N2108);
and AND4 (N2135, N2134, N2083, N13, N1289);
nor NOR3 (N2136, N2112, N1715, N236);
xor XOR2 (N2137, N2111, N1094);
buf BUF1 (N2138, N2136);
or OR3 (N2139, N2132, N1228, N856);
nor NOR4 (N2140, N2139, N531, N1295, N879);
not NOT1 (N2141, N2128);
nor NOR4 (N2142, N2133, N2123, N1613, N1446);
or OR2 (N2143, N2138, N149);
nand NAND4 (N2144, N2142, N1845, N339, N1589);
buf BUF1 (N2145, N2121);
not NOT1 (N2146, N2145);
nand NAND3 (N2147, N2144, N1606, N1115);
nor NOR4 (N2148, N2146, N1461, N1730, N609);
not NOT1 (N2149, N2141);
or OR3 (N2150, N2126, N1971, N929);
buf BUF1 (N2151, N2147);
xor XOR2 (N2152, N2151, N1785);
and AND2 (N2153, N2149, N419);
nor NOR3 (N2154, N2150, N1987, N1326);
nor NOR3 (N2155, N2152, N1296, N1515);
buf BUF1 (N2156, N2154);
buf BUF1 (N2157, N2137);
nand NAND3 (N2158, N2143, N2111, N988);
nand NAND3 (N2159, N2135, N2120, N2118);
nand NAND4 (N2160, N2158, N1629, N1107, N650);
or OR4 (N2161, N2157, N72, N1588, N1838);
and AND4 (N2162, N2153, N1342, N700, N1595);
not NOT1 (N2163, N2155);
nand NAND4 (N2164, N2148, N381, N729, N2023);
and AND2 (N2165, N2162, N882);
or OR2 (N2166, N2159, N1835);
nand NAND2 (N2167, N2166, N1015);
nor NOR3 (N2168, N2167, N1928, N969);
buf BUF1 (N2169, N2163);
or OR4 (N2170, N2156, N404, N1010, N150);
or OR2 (N2171, N2098, N1784);
nand NAND2 (N2172, N2130, N692);
buf BUF1 (N2173, N2165);
nand NAND4 (N2174, N2168, N2004, N2060, N1464);
and AND4 (N2175, N2172, N638, N1768, N833);
nand NAND3 (N2176, N2174, N817, N1583);
nor NOR4 (N2177, N2140, N332, N1808, N1571);
or OR2 (N2178, N2175, N259);
not NOT1 (N2179, N2178);
buf BUF1 (N2180, N2164);
and AND3 (N2181, N2160, N831, N269);
nor NOR2 (N2182, N2170, N1423);
buf BUF1 (N2183, N2176);
not NOT1 (N2184, N2169);
and AND4 (N2185, N2180, N275, N1123, N1265);
and AND4 (N2186, N2181, N1366, N1260, N1914);
and AND2 (N2187, N2173, N588);
nor NOR2 (N2188, N2179, N1284);
and AND2 (N2189, N2161, N554);
or OR4 (N2190, N2171, N1016, N1066, N553);
xor XOR2 (N2191, N2185, N1888);
or OR4 (N2192, N2177, N254, N1198, N1979);
not NOT1 (N2193, N2182);
and AND2 (N2194, N2192, N83);
xor XOR2 (N2195, N2191, N1143);
and AND4 (N2196, N2193, N1147, N1850, N204);
nand NAND4 (N2197, N2195, N531, N2162, N1749);
or OR3 (N2198, N2189, N122, N832);
not NOT1 (N2199, N2196);
buf BUF1 (N2200, N2187);
and AND4 (N2201, N2188, N1947, N1733, N1189);
buf BUF1 (N2202, N2201);
not NOT1 (N2203, N2194);
or OR2 (N2204, N2183, N1070);
xor XOR2 (N2205, N2197, N1416);
nor NOR3 (N2206, N2202, N2142, N544);
not NOT1 (N2207, N2206);
nor NOR3 (N2208, N2207, N1237, N1690);
nand NAND4 (N2209, N2200, N1841, N951, N582);
or OR2 (N2210, N2184, N2108);
xor XOR2 (N2211, N2186, N1509);
nor NOR4 (N2212, N2209, N1949, N1497, N516);
not NOT1 (N2213, N2190);
not NOT1 (N2214, N2212);
not NOT1 (N2215, N2205);
or OR2 (N2216, N2203, N876);
nor NOR4 (N2217, N2214, N671, N900, N2166);
or OR3 (N2218, N2211, N2162, N120);
and AND4 (N2219, N2218, N15, N990, N512);
xor XOR2 (N2220, N2204, N1515);
nor NOR3 (N2221, N2199, N176, N246);
nand NAND4 (N2222, N2215, N340, N311, N1655);
buf BUF1 (N2223, N2217);
not NOT1 (N2224, N2219);
or OR3 (N2225, N2223, N1089, N48);
buf BUF1 (N2226, N2216);
nor NOR2 (N2227, N2221, N1286);
and AND4 (N2228, N2198, N1617, N1640, N1847);
nor NOR4 (N2229, N2213, N23, N1425, N569);
or OR4 (N2230, N2226, N360, N1379, N313);
nand NAND2 (N2231, N2224, N351);
nor NOR3 (N2232, N2227, N1135, N109);
and AND2 (N2233, N2230, N627);
not NOT1 (N2234, N2222);
not NOT1 (N2235, N2231);
nor NOR3 (N2236, N2229, N1921, N1790);
not NOT1 (N2237, N2220);
buf BUF1 (N2238, N2228);
not NOT1 (N2239, N2225);
buf BUF1 (N2240, N2233);
and AND3 (N2241, N2239, N125, N1787);
nor NOR3 (N2242, N2210, N1231, N1777);
buf BUF1 (N2243, N2238);
buf BUF1 (N2244, N2237);
not NOT1 (N2245, N2234);
buf BUF1 (N2246, N2243);
buf BUF1 (N2247, N2244);
not NOT1 (N2248, N2245);
not NOT1 (N2249, N2240);
nor NOR4 (N2250, N2232, N1173, N2001, N1928);
nor NOR2 (N2251, N2208, N1486);
xor XOR2 (N2252, N2247, N947);
nor NOR4 (N2253, N2241, N353, N587, N996);
xor XOR2 (N2254, N2250, N1501);
nand NAND4 (N2255, N2251, N1530, N84, N2106);
not NOT1 (N2256, N2253);
or OR2 (N2257, N2252, N387);
buf BUF1 (N2258, N2257);
nor NOR3 (N2259, N2254, N835, N1308);
nor NOR4 (N2260, N2249, N1579, N1343, N495);
nand NAND2 (N2261, N2246, N2108);
nand NAND2 (N2262, N2258, N1300);
buf BUF1 (N2263, N2248);
and AND3 (N2264, N2242, N635, N39);
xor XOR2 (N2265, N2260, N954);
nand NAND3 (N2266, N2256, N1941, N618);
and AND2 (N2267, N2262, N1207);
or OR2 (N2268, N2236, N1599);
nand NAND2 (N2269, N2261, N712);
nor NOR3 (N2270, N2269, N2068, N100);
buf BUF1 (N2271, N2255);
nand NAND2 (N2272, N2259, N335);
nand NAND2 (N2273, N2266, N857);
xor XOR2 (N2274, N2264, N2198);
or OR2 (N2275, N2270, N512);
buf BUF1 (N2276, N2273);
nor NOR3 (N2277, N2235, N660, N1299);
buf BUF1 (N2278, N2265);
nor NOR3 (N2279, N2263, N6, N250);
nand NAND4 (N2280, N2275, N2155, N2, N190);
nand NAND3 (N2281, N2274, N866, N1844);
nand NAND4 (N2282, N2278, N1485, N1580, N841);
and AND4 (N2283, N2277, N52, N2112, N413);
buf BUF1 (N2284, N2279);
nand NAND2 (N2285, N2267, N1907);
or OR4 (N2286, N2284, N1354, N124, N1687);
xor XOR2 (N2287, N2282, N1619);
not NOT1 (N2288, N2285);
xor XOR2 (N2289, N2271, N674);
xor XOR2 (N2290, N2281, N1031);
nor NOR4 (N2291, N2289, N1766, N1899, N1);
xor XOR2 (N2292, N2268, N226);
or OR2 (N2293, N2286, N1016);
xor XOR2 (N2294, N2293, N339);
not NOT1 (N2295, N2276);
and AND4 (N2296, N2287, N1766, N1263, N1721);
buf BUF1 (N2297, N2290);
and AND3 (N2298, N2292, N1445, N202);
nand NAND3 (N2299, N2288, N196, N226);
nand NAND2 (N2300, N2291, N1521);
and AND3 (N2301, N2299, N10, N1089);
nor NOR3 (N2302, N2295, N900, N2030);
not NOT1 (N2303, N2283);
and AND4 (N2304, N2296, N1216, N826, N987);
xor XOR2 (N2305, N2294, N1227);
not NOT1 (N2306, N2305);
nor NOR2 (N2307, N2280, N1533);
buf BUF1 (N2308, N2301);
or OR2 (N2309, N2298, N75);
not NOT1 (N2310, N2302);
nor NOR4 (N2311, N2303, N149, N568, N1659);
nor NOR4 (N2312, N2272, N287, N1479, N669);
or OR4 (N2313, N2306, N374, N2312, N2180);
xor XOR2 (N2314, N1419, N510);
buf BUF1 (N2315, N2310);
xor XOR2 (N2316, N2309, N1644);
buf BUF1 (N2317, N2311);
not NOT1 (N2318, N2313);
xor XOR2 (N2319, N2318, N1309);
not NOT1 (N2320, N2308);
nand NAND2 (N2321, N2319, N277);
nor NOR4 (N2322, N2307, N2215, N1608, N1758);
buf BUF1 (N2323, N2320);
buf BUF1 (N2324, N2316);
or OR4 (N2325, N2315, N107, N81, N1636);
not NOT1 (N2326, N2304);
xor XOR2 (N2327, N2323, N382);
or OR3 (N2328, N2327, N1019, N1294);
nand NAND2 (N2329, N2317, N1270);
not NOT1 (N2330, N2314);
nand NAND4 (N2331, N2330, N2214, N656, N2297);
and AND4 (N2332, N1903, N1803, N365, N1143);
not NOT1 (N2333, N2326);
nor NOR3 (N2334, N2333, N308, N629);
nor NOR4 (N2335, N2322, N1302, N1113, N1683);
and AND2 (N2336, N2332, N787);
or OR4 (N2337, N2300, N1319, N2, N215);
nand NAND4 (N2338, N2337, N1247, N2045, N977);
or OR4 (N2339, N2331, N1108, N1197, N560);
not NOT1 (N2340, N2328);
buf BUF1 (N2341, N2335);
nand NAND4 (N2342, N2341, N1218, N282, N848);
nand NAND3 (N2343, N2336, N372, N1964);
nor NOR4 (N2344, N2338, N837, N1924, N469);
or OR4 (N2345, N2325, N1908, N666, N687);
nand NAND3 (N2346, N2321, N307, N1652);
not NOT1 (N2347, N2342);
buf BUF1 (N2348, N2345);
nand NAND3 (N2349, N2348, N524, N961);
or OR4 (N2350, N2329, N2132, N1375, N1241);
not NOT1 (N2351, N2347);
nand NAND4 (N2352, N2351, N1193, N1400, N978);
nor NOR2 (N2353, N2324, N2044);
xor XOR2 (N2354, N2339, N598);
nor NOR3 (N2355, N2350, N732, N1613);
xor XOR2 (N2356, N2354, N1734);
or OR4 (N2357, N2355, N1, N302, N1609);
and AND3 (N2358, N2356, N610, N287);
nor NOR3 (N2359, N2358, N90, N2221);
nor NOR3 (N2360, N2346, N621, N1017);
nand NAND4 (N2361, N2340, N1613, N81, N2200);
and AND4 (N2362, N2334, N1718, N983, N1332);
and AND4 (N2363, N2360, N2286, N1056, N1652);
buf BUF1 (N2364, N2362);
nor NOR4 (N2365, N2353, N1948, N907, N935);
not NOT1 (N2366, N2365);
or OR4 (N2367, N2359, N30, N2288, N2026);
buf BUF1 (N2368, N2349);
and AND3 (N2369, N2343, N1512, N667);
nand NAND3 (N2370, N2344, N2027, N1106);
buf BUF1 (N2371, N2368);
buf BUF1 (N2372, N2357);
xor XOR2 (N2373, N2363, N1425);
not NOT1 (N2374, N2367);
not NOT1 (N2375, N2374);
nor NOR4 (N2376, N2375, N568, N963, N363);
not NOT1 (N2377, N2373);
nor NOR2 (N2378, N2364, N1917);
buf BUF1 (N2379, N2376);
or OR3 (N2380, N2372, N2076, N1130);
and AND4 (N2381, N2379, N730, N1650, N986);
buf BUF1 (N2382, N2380);
nor NOR4 (N2383, N2352, N1811, N2123, N1308);
not NOT1 (N2384, N2383);
and AND4 (N2385, N2384, N719, N1761, N1895);
not NOT1 (N2386, N2382);
and AND4 (N2387, N2378, N1079, N607, N141);
and AND3 (N2388, N2377, N1483, N203);
or OR4 (N2389, N2387, N694, N453, N2238);
nor NOR2 (N2390, N2361, N1911);
xor XOR2 (N2391, N2385, N844);
and AND4 (N2392, N2370, N1251, N608, N2182);
nand NAND2 (N2393, N2386, N1412);
buf BUF1 (N2394, N2393);
nor NOR4 (N2395, N2371, N534, N1762, N1954);
and AND3 (N2396, N2366, N1713, N1568);
and AND4 (N2397, N2394, N2342, N934, N881);
buf BUF1 (N2398, N2389);
and AND4 (N2399, N2396, N1911, N1078, N1228);
or OR3 (N2400, N2392, N1842, N408);
or OR3 (N2401, N2381, N658, N1991);
not NOT1 (N2402, N2391);
nor NOR4 (N2403, N2388, N1798, N1092, N1073);
not NOT1 (N2404, N2403);
nand NAND2 (N2405, N2401, N1129);
or OR2 (N2406, N2369, N867);
xor XOR2 (N2407, N2390, N1144);
nor NOR3 (N2408, N2398, N464, N1484);
xor XOR2 (N2409, N2405, N1635);
not NOT1 (N2410, N2409);
buf BUF1 (N2411, N2402);
nand NAND2 (N2412, N2406, N462);
nor NOR4 (N2413, N2408, N359, N909, N1932);
nand NAND2 (N2414, N2407, N1491);
xor XOR2 (N2415, N2400, N744);
xor XOR2 (N2416, N2413, N2136);
buf BUF1 (N2417, N2411);
or OR3 (N2418, N2404, N2131, N1873);
buf BUF1 (N2419, N2418);
or OR2 (N2420, N2412, N2158);
nor NOR2 (N2421, N2420, N890);
not NOT1 (N2422, N2410);
nor NOR2 (N2423, N2416, N2154);
nor NOR2 (N2424, N2423, N1001);
and AND4 (N2425, N2421, N1551, N1454, N2211);
not NOT1 (N2426, N2397);
buf BUF1 (N2427, N2424);
nand NAND4 (N2428, N2395, N1748, N2052, N307);
and AND3 (N2429, N2426, N413, N1277);
and AND4 (N2430, N2427, N211, N203, N1718);
nand NAND4 (N2431, N2417, N115, N307, N2355);
buf BUF1 (N2432, N2419);
nor NOR4 (N2433, N2425, N1312, N1968, N338);
and AND4 (N2434, N2428, N867, N173, N53);
or OR4 (N2435, N2414, N1122, N479, N77);
or OR3 (N2436, N2432, N2240, N881);
and AND2 (N2437, N2415, N386);
not NOT1 (N2438, N2422);
xor XOR2 (N2439, N2436, N2051);
nand NAND4 (N2440, N2438, N1220, N134, N1868);
xor XOR2 (N2441, N2437, N679);
buf BUF1 (N2442, N2434);
nor NOR2 (N2443, N2430, N1484);
not NOT1 (N2444, N2440);
xor XOR2 (N2445, N2439, N1620);
or OR3 (N2446, N2435, N831, N1943);
and AND2 (N2447, N2429, N317);
buf BUF1 (N2448, N2443);
not NOT1 (N2449, N2431);
buf BUF1 (N2450, N2449);
and AND4 (N2451, N2446, N2152, N2403, N1733);
buf BUF1 (N2452, N2451);
and AND4 (N2453, N2444, N1832, N100, N1502);
nand NAND3 (N2454, N2433, N2074, N709);
not NOT1 (N2455, N2452);
nor NOR2 (N2456, N2441, N1068);
buf BUF1 (N2457, N2454);
and AND3 (N2458, N2455, N2045, N2211);
nor NOR3 (N2459, N2450, N1389, N581);
xor XOR2 (N2460, N2453, N782);
nor NOR2 (N2461, N2457, N1827);
or OR2 (N2462, N2448, N1170);
or OR3 (N2463, N2447, N1733, N2035);
not NOT1 (N2464, N2456);
nand NAND4 (N2465, N2463, N2381, N1597, N1341);
xor XOR2 (N2466, N2460, N314);
nand NAND4 (N2467, N2459, N1542, N1446, N776);
not NOT1 (N2468, N2461);
nand NAND4 (N2469, N2458, N1553, N797, N2313);
or OR2 (N2470, N2469, N2140);
buf BUF1 (N2471, N2445);
nor NOR4 (N2472, N2399, N1391, N1472, N1103);
xor XOR2 (N2473, N2470, N88);
buf BUF1 (N2474, N2473);
buf BUF1 (N2475, N2442);
nand NAND3 (N2476, N2474, N365, N335);
nor NOR2 (N2477, N2466, N1684);
and AND3 (N2478, N2462, N658, N1215);
buf BUF1 (N2479, N2465);
not NOT1 (N2480, N2479);
and AND2 (N2481, N2476, N445);
nor NOR4 (N2482, N2471, N323, N1736, N2372);
nor NOR4 (N2483, N2480, N1918, N906, N183);
nand NAND3 (N2484, N2481, N290, N2226);
not NOT1 (N2485, N2464);
buf BUF1 (N2486, N2472);
or OR3 (N2487, N2483, N1187, N1233);
nand NAND3 (N2488, N2482, N1273, N1180);
not NOT1 (N2489, N2487);
and AND4 (N2490, N2478, N657, N2354, N817);
buf BUF1 (N2491, N2485);
not NOT1 (N2492, N2490);
nand NAND4 (N2493, N2491, N18, N2074, N1535);
nor NOR2 (N2494, N2468, N1707);
not NOT1 (N2495, N2484);
and AND2 (N2496, N2492, N533);
and AND3 (N2497, N2496, N1721, N935);
nor NOR2 (N2498, N2486, N1692);
not NOT1 (N2499, N2475);
nand NAND4 (N2500, N2467, N2083, N1203, N1662);
nor NOR3 (N2501, N2498, N1455, N804);
not NOT1 (N2502, N2494);
or OR4 (N2503, N2493, N1702, N1069, N1389);
nor NOR2 (N2504, N2501, N1346);
nand NAND4 (N2505, N2499, N849, N2159, N1312);
or OR3 (N2506, N2488, N1406, N2285);
nand NAND3 (N2507, N2495, N1367, N1900);
or OR3 (N2508, N2497, N1265, N1898);
or OR4 (N2509, N2489, N530, N29, N141);
nand NAND3 (N2510, N2503, N2372, N2000);
not NOT1 (N2511, N2502);
nor NOR4 (N2512, N2510, N1548, N1151, N1893);
nor NOR4 (N2513, N2504, N1323, N2405, N2296);
xor XOR2 (N2514, N2505, N1318);
or OR3 (N2515, N2506, N1430, N2493);
or OR3 (N2516, N2500, N728, N1854);
nor NOR4 (N2517, N2509, N1617, N2063, N618);
not NOT1 (N2518, N2512);
and AND3 (N2519, N2508, N1656, N2444);
not NOT1 (N2520, N2513);
nand NAND2 (N2521, N2516, N763);
nand NAND3 (N2522, N2521, N1657, N594);
and AND2 (N2523, N2515, N1014);
and AND4 (N2524, N2520, N2262, N413, N568);
nor NOR2 (N2525, N2514, N2494);
xor XOR2 (N2526, N2477, N1630);
nor NOR4 (N2527, N2519, N2453, N1011, N949);
or OR4 (N2528, N2524, N458, N1000, N877);
not NOT1 (N2529, N2525);
nor NOR2 (N2530, N2528, N311);
or OR4 (N2531, N2529, N903, N2300, N1788);
and AND3 (N2532, N2517, N1540, N948);
nand NAND2 (N2533, N2507, N257);
nor NOR4 (N2534, N2511, N1258, N1278, N2379);
nor NOR2 (N2535, N2532, N1310);
not NOT1 (N2536, N2523);
buf BUF1 (N2537, N2536);
or OR2 (N2538, N2530, N2272);
nor NOR4 (N2539, N2527, N1910, N125, N535);
or OR4 (N2540, N2522, N2338, N2342, N2426);
not NOT1 (N2541, N2533);
xor XOR2 (N2542, N2541, N497);
nor NOR4 (N2543, N2531, N1602, N710, N1430);
and AND4 (N2544, N2543, N1828, N2137, N877);
nor NOR2 (N2545, N2518, N2483);
nor NOR3 (N2546, N2534, N1007, N2189);
buf BUF1 (N2547, N2544);
or OR4 (N2548, N2547, N355, N1764, N2217);
or OR4 (N2549, N2546, N1603, N1902, N2203);
nand NAND4 (N2550, N2545, N1512, N40, N1830);
or OR2 (N2551, N2539, N1515);
xor XOR2 (N2552, N2549, N2213);
nor NOR3 (N2553, N2542, N1307, N617);
xor XOR2 (N2554, N2535, N1937);
nor NOR2 (N2555, N2548, N680);
nor NOR2 (N2556, N2555, N315);
nor NOR3 (N2557, N2553, N121, N44);
or OR4 (N2558, N2552, N2399, N860, N260);
buf BUF1 (N2559, N2558);
nor NOR4 (N2560, N2538, N871, N1321, N673);
and AND4 (N2561, N2537, N1020, N1562, N1201);
xor XOR2 (N2562, N2540, N1986);
xor XOR2 (N2563, N2561, N1506);
nor NOR2 (N2564, N2554, N2385);
or OR3 (N2565, N2557, N2342, N633);
nor NOR2 (N2566, N2526, N396);
or OR2 (N2567, N2560, N1841);
nand NAND2 (N2568, N2567, N1912);
xor XOR2 (N2569, N2559, N2385);
not NOT1 (N2570, N2565);
nor NOR3 (N2571, N2562, N1649, N1301);
buf BUF1 (N2572, N2551);
nand NAND4 (N2573, N2556, N25, N2555, N200);
not NOT1 (N2574, N2571);
and AND2 (N2575, N2572, N1756);
or OR3 (N2576, N2564, N2290, N184);
nor NOR3 (N2577, N2569, N1134, N1285);
or OR2 (N2578, N2550, N1892);
nor NOR4 (N2579, N2563, N898, N224, N1775);
not NOT1 (N2580, N2568);
nor NOR4 (N2581, N2576, N2096, N306, N445);
or OR3 (N2582, N2575, N180, N1617);
and AND3 (N2583, N2582, N2523, N54);
nor NOR4 (N2584, N2573, N912, N2508, N1752);
xor XOR2 (N2585, N2566, N2041);
or OR2 (N2586, N2570, N2485);
buf BUF1 (N2587, N2584);
buf BUF1 (N2588, N2579);
buf BUF1 (N2589, N2580);
xor XOR2 (N2590, N2588, N653);
nor NOR4 (N2591, N2577, N1395, N1829, N1260);
and AND2 (N2592, N2591, N903);
or OR3 (N2593, N2585, N1888, N1329);
not NOT1 (N2594, N2590);
and AND4 (N2595, N2574, N805, N1239, N2349);
nor NOR3 (N2596, N2583, N1768, N1353);
buf BUF1 (N2597, N2589);
and AND2 (N2598, N2593, N336);
nand NAND3 (N2599, N2578, N2128, N103);
buf BUF1 (N2600, N2586);
nand NAND4 (N2601, N2595, N2142, N952, N2098);
xor XOR2 (N2602, N2599, N266);
or OR4 (N2603, N2597, N870, N2091, N2468);
and AND4 (N2604, N2600, N134, N73, N1750);
nand NAND4 (N2605, N2604, N514, N1839, N526);
nor NOR2 (N2606, N2592, N290);
nand NAND4 (N2607, N2581, N797, N1978, N828);
nor NOR2 (N2608, N2594, N305);
or OR4 (N2609, N2602, N1018, N1496, N1793);
buf BUF1 (N2610, N2598);
nor NOR4 (N2611, N2596, N1637, N534, N87);
nor NOR4 (N2612, N2606, N1435, N276, N602);
nor NOR4 (N2613, N2611, N571, N2059, N1576);
nor NOR3 (N2614, N2601, N2253, N853);
nor NOR3 (N2615, N2587, N559, N1405);
buf BUF1 (N2616, N2605);
xor XOR2 (N2617, N2610, N1727);
nand NAND2 (N2618, N2603, N1994);
xor XOR2 (N2619, N2617, N842);
or OR3 (N2620, N2616, N1234, N2258);
nand NAND3 (N2621, N2615, N393, N1023);
not NOT1 (N2622, N2619);
nand NAND4 (N2623, N2609, N322, N2559, N77);
nand NAND3 (N2624, N2612, N609, N1449);
not NOT1 (N2625, N2618);
xor XOR2 (N2626, N2608, N776);
xor XOR2 (N2627, N2621, N8);
or OR4 (N2628, N2626, N1332, N12, N1645);
buf BUF1 (N2629, N2625);
or OR2 (N2630, N2627, N541);
nand NAND3 (N2631, N2613, N1059, N489);
and AND3 (N2632, N2630, N1142, N1671);
nor NOR3 (N2633, N2623, N2248, N580);
not NOT1 (N2634, N2633);
nand NAND3 (N2635, N2634, N1254, N2269);
nor NOR3 (N2636, N2614, N1741, N2443);
nor NOR4 (N2637, N2635, N2450, N1890, N2468);
not NOT1 (N2638, N2631);
nand NAND3 (N2639, N2629, N269, N443);
or OR4 (N2640, N2632, N1170, N2045, N2068);
buf BUF1 (N2641, N2624);
nand NAND3 (N2642, N2622, N418, N399);
or OR3 (N2643, N2638, N2577, N457);
nor NOR2 (N2644, N2641, N2560);
nor NOR3 (N2645, N2639, N402, N533);
nor NOR3 (N2646, N2636, N1674, N2321);
nor NOR3 (N2647, N2607, N1961, N1888);
not NOT1 (N2648, N2645);
or OR3 (N2649, N2644, N2065, N967);
xor XOR2 (N2650, N2649, N2431);
nor NOR3 (N2651, N2648, N1776, N2151);
and AND3 (N2652, N2643, N2436, N2200);
nand NAND4 (N2653, N2646, N2413, N1530, N1956);
nor NOR3 (N2654, N2642, N2463, N2435);
or OR4 (N2655, N2650, N344, N1450, N540);
or OR2 (N2656, N2637, N2627);
buf BUF1 (N2657, N2647);
nor NOR3 (N2658, N2652, N1685, N1510);
xor XOR2 (N2659, N2655, N1414);
or OR4 (N2660, N2628, N2362, N339, N666);
nand NAND4 (N2661, N2640, N283, N1372, N183);
nor NOR4 (N2662, N2654, N1696, N2141, N1360);
nand NAND2 (N2663, N2661, N2348);
buf BUF1 (N2664, N2656);
xor XOR2 (N2665, N2651, N1474);
or OR2 (N2666, N2662, N1406);
nor NOR2 (N2667, N2658, N658);
nor NOR4 (N2668, N2657, N1929, N2079, N775);
or OR3 (N2669, N2665, N1167, N152);
or OR3 (N2670, N2664, N2357, N2309);
nor NOR3 (N2671, N2660, N1243, N2226);
or OR4 (N2672, N2669, N1051, N576, N645);
or OR2 (N2673, N2672, N362);
nor NOR2 (N2674, N2670, N1683);
nand NAND2 (N2675, N2663, N1781);
nor NOR2 (N2676, N2675, N1465);
and AND2 (N2677, N2620, N411);
xor XOR2 (N2678, N2668, N421);
not NOT1 (N2679, N2677);
nand NAND3 (N2680, N2678, N1052, N1148);
and AND3 (N2681, N2674, N686, N2507);
buf BUF1 (N2682, N2679);
not NOT1 (N2683, N2676);
nor NOR3 (N2684, N2653, N2541, N143);
or OR3 (N2685, N2684, N816, N847);
nor NOR2 (N2686, N2671, N612);
nor NOR3 (N2687, N2680, N1708, N2424);
buf BUF1 (N2688, N2683);
nor NOR3 (N2689, N2673, N119, N957);
not NOT1 (N2690, N2686);
buf BUF1 (N2691, N2659);
nor NOR4 (N2692, N2667, N219, N1636, N741);
or OR3 (N2693, N2681, N1360, N1457);
nor NOR2 (N2694, N2689, N492);
nand NAND4 (N2695, N2682, N1421, N1624, N1171);
xor XOR2 (N2696, N2692, N580);
nor NOR4 (N2697, N2695, N1336, N2112, N2143);
and AND2 (N2698, N2696, N2567);
xor XOR2 (N2699, N2691, N1335);
nor NOR4 (N2700, N2687, N439, N900, N752);
not NOT1 (N2701, N2688);
and AND4 (N2702, N2690, N930, N2338, N742);
buf BUF1 (N2703, N2702);
or OR3 (N2704, N2699, N739, N1985);
buf BUF1 (N2705, N2693);
buf BUF1 (N2706, N2701);
and AND4 (N2707, N2694, N1967, N2658, N356);
nand NAND2 (N2708, N2697, N1579);
nor NOR4 (N2709, N2706, N530, N556, N767);
or OR2 (N2710, N2708, N4);
not NOT1 (N2711, N2704);
not NOT1 (N2712, N2685);
buf BUF1 (N2713, N2712);
or OR3 (N2714, N2713, N608, N307);
xor XOR2 (N2715, N2700, N2318);
nor NOR4 (N2716, N2666, N1212, N192, N746);
nor NOR2 (N2717, N2705, N1894);
nand NAND4 (N2718, N2717, N2310, N235, N1525);
and AND4 (N2719, N2718, N1414, N361, N428);
buf BUF1 (N2720, N2711);
and AND2 (N2721, N2720, N829);
not NOT1 (N2722, N2715);
buf BUF1 (N2723, N2709);
xor XOR2 (N2724, N2714, N2270);
and AND2 (N2725, N2721, N245);
or OR4 (N2726, N2716, N127, N328, N608);
nor NOR4 (N2727, N2698, N823, N218, N895);
buf BUF1 (N2728, N2710);
xor XOR2 (N2729, N2728, N1425);
buf BUF1 (N2730, N2719);
nor NOR4 (N2731, N2725, N2149, N1471, N1811);
xor XOR2 (N2732, N2731, N839);
nor NOR4 (N2733, N2722, N695, N2104, N33);
and AND2 (N2734, N2733, N2512);
buf BUF1 (N2735, N2729);
buf BUF1 (N2736, N2724);
or OR4 (N2737, N2707, N1576, N244, N1569);
not NOT1 (N2738, N2732);
nor NOR4 (N2739, N2726, N1914, N2087, N5);
and AND3 (N2740, N2703, N320, N1449);
and AND3 (N2741, N2730, N242, N814);
and AND2 (N2742, N2738, N684);
nor NOR3 (N2743, N2727, N2676, N1472);
xor XOR2 (N2744, N2739, N140);
nor NOR4 (N2745, N2723, N2136, N1717, N1753);
nand NAND3 (N2746, N2736, N1050, N369);
nor NOR3 (N2747, N2744, N394, N76);
xor XOR2 (N2748, N2740, N1057);
buf BUF1 (N2749, N2745);
or OR4 (N2750, N2747, N2114, N1678, N290);
xor XOR2 (N2751, N2742, N1911);
or OR3 (N2752, N2750, N2426, N762);
not NOT1 (N2753, N2743);
or OR4 (N2754, N2746, N2673, N407, N1439);
nor NOR2 (N2755, N2753, N1564);
nor NOR4 (N2756, N2734, N337, N459, N131);
nand NAND3 (N2757, N2737, N101, N417);
not NOT1 (N2758, N2752);
nand NAND2 (N2759, N2741, N2630);
not NOT1 (N2760, N2759);
buf BUF1 (N2761, N2760);
nand NAND4 (N2762, N2751, N760, N1082, N133);
or OR4 (N2763, N2758, N2723, N1433, N633);
not NOT1 (N2764, N2755);
nor NOR3 (N2765, N2757, N2649, N1734);
and AND2 (N2766, N2756, N2282);
xor XOR2 (N2767, N2766, N1522);
buf BUF1 (N2768, N2767);
not NOT1 (N2769, N2748);
buf BUF1 (N2770, N2768);
nand NAND3 (N2771, N2735, N1364, N2449);
or OR4 (N2772, N2764, N652, N1428, N83);
not NOT1 (N2773, N2769);
xor XOR2 (N2774, N2749, N203);
and AND4 (N2775, N2774, N1203, N2506, N2384);
buf BUF1 (N2776, N2765);
nor NOR4 (N2777, N2776, N843, N354, N1831);
nand NAND3 (N2778, N2771, N905, N1372);
nand NAND4 (N2779, N2778, N101, N1495, N2572);
and AND2 (N2780, N2770, N827);
nand NAND2 (N2781, N2780, N1868);
buf BUF1 (N2782, N2773);
buf BUF1 (N2783, N2772);
or OR4 (N2784, N2763, N225, N79, N1760);
xor XOR2 (N2785, N2784, N2701);
buf BUF1 (N2786, N2781);
nor NOR2 (N2787, N2761, N2269);
and AND2 (N2788, N2783, N2601);
buf BUF1 (N2789, N2787);
buf BUF1 (N2790, N2762);
nand NAND3 (N2791, N2788, N1286, N2319);
nand NAND2 (N2792, N2782, N56);
nor NOR2 (N2793, N2779, N768);
nand NAND4 (N2794, N2790, N1966, N1612, N1412);
nand NAND3 (N2795, N2792, N1585, N7);
xor XOR2 (N2796, N2775, N2736);
nand NAND2 (N2797, N2785, N1669);
or OR2 (N2798, N2789, N1171);
and AND2 (N2799, N2777, N2762);
not NOT1 (N2800, N2786);
xor XOR2 (N2801, N2791, N1462);
or OR2 (N2802, N2794, N919);
and AND4 (N2803, N2802, N1027, N1001, N1515);
buf BUF1 (N2804, N2796);
nand NAND3 (N2805, N2804, N1791, N1472);
nor NOR2 (N2806, N2800, N984);
nor NOR4 (N2807, N2806, N868, N1453, N1588);
nor NOR2 (N2808, N2797, N842);
nand NAND3 (N2809, N2808, N427, N2358);
buf BUF1 (N2810, N2798);
buf BUF1 (N2811, N2801);
nand NAND2 (N2812, N2811, N1512);
not NOT1 (N2813, N2812);
buf BUF1 (N2814, N2795);
and AND3 (N2815, N2803, N2183, N1941);
buf BUF1 (N2816, N2754);
nor NOR4 (N2817, N2813, N1141, N817, N257);
nand NAND3 (N2818, N2816, N2224, N1292);
or OR3 (N2819, N2810, N1901, N1983);
nor NOR3 (N2820, N2793, N32, N1354);
nor NOR2 (N2821, N2807, N396);
xor XOR2 (N2822, N2809, N1661);
or OR4 (N2823, N2814, N2380, N1853, N1472);
not NOT1 (N2824, N2822);
xor XOR2 (N2825, N2824, N293);
not NOT1 (N2826, N2820);
nand NAND4 (N2827, N2815, N817, N1444, N1308);
nand NAND3 (N2828, N2817, N2683, N517);
not NOT1 (N2829, N2828);
nand NAND4 (N2830, N2823, N1065, N2776, N261);
nand NAND4 (N2831, N2827, N2557, N889, N2773);
and AND2 (N2832, N2818, N810);
and AND3 (N2833, N2821, N589, N331);
or OR3 (N2834, N2819, N2276, N275);
buf BUF1 (N2835, N2830);
nor NOR3 (N2836, N2826, N145, N1377);
nor NOR2 (N2837, N2805, N624);
buf BUF1 (N2838, N2836);
or OR2 (N2839, N2832, N1889);
nor NOR4 (N2840, N2833, N1960, N1818, N446);
not NOT1 (N2841, N2834);
or OR2 (N2842, N2841, N2127);
or OR2 (N2843, N2838, N1387);
nor NOR4 (N2844, N2829, N701, N908, N916);
or OR2 (N2845, N2840, N1163);
buf BUF1 (N2846, N2844);
xor XOR2 (N2847, N2837, N4);
buf BUF1 (N2848, N2843);
and AND3 (N2849, N2799, N344, N2206);
or OR3 (N2850, N2848, N819, N544);
nor NOR4 (N2851, N2835, N2338, N1592, N1486);
nor NOR4 (N2852, N2831, N419, N991, N64);
buf BUF1 (N2853, N2845);
xor XOR2 (N2854, N2825, N167);
and AND2 (N2855, N2839, N2447);
nand NAND3 (N2856, N2854, N2307, N697);
and AND4 (N2857, N2853, N2572, N1134, N1999);
and AND4 (N2858, N2851, N376, N512, N109);
xor XOR2 (N2859, N2852, N618);
or OR3 (N2860, N2859, N2467, N289);
nor NOR2 (N2861, N2860, N751);
buf BUF1 (N2862, N2858);
nor NOR3 (N2863, N2846, N1829, N734);
nand NAND2 (N2864, N2857, N310);
and AND2 (N2865, N2855, N2438);
not NOT1 (N2866, N2863);
nor NOR3 (N2867, N2856, N1640, N2719);
buf BUF1 (N2868, N2865);
and AND4 (N2869, N2842, N20, N2867, N473);
xor XOR2 (N2870, N2389, N773);
not NOT1 (N2871, N2866);
xor XOR2 (N2872, N2850, N1580);
xor XOR2 (N2873, N2868, N894);
and AND4 (N2874, N2872, N2740, N437, N25);
or OR4 (N2875, N2869, N2732, N97, N2027);
not NOT1 (N2876, N2849);
not NOT1 (N2877, N2874);
and AND2 (N2878, N2862, N1323);
or OR2 (N2879, N2876, N2572);
nor NOR4 (N2880, N2875, N2117, N1065, N335);
and AND4 (N2881, N2877, N1432, N2411, N2138);
buf BUF1 (N2882, N2871);
xor XOR2 (N2883, N2847, N2445);
xor XOR2 (N2884, N2882, N2254);
not NOT1 (N2885, N2878);
or OR3 (N2886, N2873, N2417, N2525);
xor XOR2 (N2887, N2864, N1476);
buf BUF1 (N2888, N2883);
nand NAND4 (N2889, N2880, N2530, N694, N768);
buf BUF1 (N2890, N2887);
xor XOR2 (N2891, N2881, N1113);
not NOT1 (N2892, N2886);
buf BUF1 (N2893, N2888);
nor NOR4 (N2894, N2861, N2026, N1937, N1091);
nor NOR2 (N2895, N2894, N1418);
xor XOR2 (N2896, N2891, N2601);
not NOT1 (N2897, N2884);
nand NAND3 (N2898, N2896, N1449, N1159);
not NOT1 (N2899, N2890);
or OR2 (N2900, N2895, N1193);
not NOT1 (N2901, N2898);
buf BUF1 (N2902, N2900);
not NOT1 (N2903, N2902);
or OR3 (N2904, N2885, N1216, N1710);
xor XOR2 (N2905, N2893, N1323);
nand NAND3 (N2906, N2889, N1571, N2770);
not NOT1 (N2907, N2879);
or OR4 (N2908, N2901, N936, N2370, N1742);
nand NAND2 (N2909, N2904, N2173);
nor NOR2 (N2910, N2892, N903);
not NOT1 (N2911, N2907);
not NOT1 (N2912, N2905);
and AND3 (N2913, N2908, N564, N2020);
nand NAND4 (N2914, N2913, N2746, N1504, N1263);
not NOT1 (N2915, N2870);
nand NAND2 (N2916, N2914, N2678);
xor XOR2 (N2917, N2916, N327);
nor NOR4 (N2918, N2912, N2698, N2267, N889);
not NOT1 (N2919, N2909);
nand NAND4 (N2920, N2917, N2562, N647, N1695);
and AND3 (N2921, N2911, N1333, N1900);
not NOT1 (N2922, N2899);
buf BUF1 (N2923, N2915);
nor NOR3 (N2924, N2903, N1877, N2426);
xor XOR2 (N2925, N2921, N2883);
not NOT1 (N2926, N2897);
buf BUF1 (N2927, N2924);
or OR2 (N2928, N2919, N544);
or OR3 (N2929, N2923, N945, N2796);
xor XOR2 (N2930, N2925, N1353);
or OR3 (N2931, N2922, N1583, N1440);
not NOT1 (N2932, N2918);
and AND2 (N2933, N2932, N1751);
buf BUF1 (N2934, N2929);
not NOT1 (N2935, N2910);
not NOT1 (N2936, N2931);
buf BUF1 (N2937, N2935);
not NOT1 (N2938, N2927);
nor NOR3 (N2939, N2920, N2146, N2558);
nand NAND4 (N2940, N2937, N246, N162, N2314);
or OR2 (N2941, N2934, N813);
nand NAND2 (N2942, N2938, N1186);
xor XOR2 (N2943, N2939, N1428);
buf BUF1 (N2944, N2928);
buf BUF1 (N2945, N2943);
or OR4 (N2946, N2945, N1154, N931, N1410);
nor NOR2 (N2947, N2940, N1255);
nor NOR2 (N2948, N2933, N2117);
xor XOR2 (N2949, N2942, N2629);
not NOT1 (N2950, N2948);
buf BUF1 (N2951, N2906);
xor XOR2 (N2952, N2941, N2096);
and AND4 (N2953, N2930, N2012, N1550, N435);
nand NAND3 (N2954, N2946, N2671, N969);
and AND2 (N2955, N2944, N1336);
xor XOR2 (N2956, N2949, N2944);
buf BUF1 (N2957, N2953);
nor NOR2 (N2958, N2955, N2937);
nand NAND4 (N2959, N2954, N2068, N2044, N2886);
buf BUF1 (N2960, N2950);
not NOT1 (N2961, N2952);
or OR2 (N2962, N2957, N2419);
buf BUF1 (N2963, N2962);
nand NAND2 (N2964, N2926, N59);
nand NAND3 (N2965, N2956, N2165, N254);
nor NOR4 (N2966, N2959, N1572, N615, N1439);
or OR2 (N2967, N2958, N1366);
buf BUF1 (N2968, N2936);
or OR4 (N2969, N2960, N841, N400, N2246);
and AND2 (N2970, N2968, N442);
nand NAND4 (N2971, N2951, N267, N2552, N1861);
xor XOR2 (N2972, N2961, N1209);
not NOT1 (N2973, N2963);
and AND4 (N2974, N2966, N708, N2049, N2151);
or OR3 (N2975, N2973, N2471, N2226);
and AND3 (N2976, N2971, N1327, N2270);
or OR3 (N2977, N2967, N2315, N2321);
not NOT1 (N2978, N2977);
buf BUF1 (N2979, N2974);
and AND2 (N2980, N2976, N1653);
nor NOR4 (N2981, N2975, N2158, N2368, N1914);
not NOT1 (N2982, N2965);
nor NOR3 (N2983, N2980, N1760, N2257);
or OR2 (N2984, N2964, N1196);
nor NOR2 (N2985, N2982, N454);
nand NAND2 (N2986, N2947, N2084);
not NOT1 (N2987, N2969);
nor NOR3 (N2988, N2983, N1137, N133);
nand NAND4 (N2989, N2981, N2517, N1314, N460);
or OR3 (N2990, N2988, N1777, N1966);
and AND3 (N2991, N2986, N1318, N352);
or OR2 (N2992, N2978, N1762);
nor NOR4 (N2993, N2984, N914, N767, N1457);
or OR2 (N2994, N2970, N101);
and AND4 (N2995, N2989, N757, N385, N2020);
xor XOR2 (N2996, N2995, N715);
not NOT1 (N2997, N2979);
nand NAND3 (N2998, N2997, N1230, N1685);
xor XOR2 (N2999, N2998, N494);
buf BUF1 (N3000, N2987);
nor NOR2 (N3001, N2993, N141);
and AND3 (N3002, N2985, N126, N1642);
nor NOR4 (N3003, N2991, N1877, N224, N284);
or OR3 (N3004, N2996, N2481, N1300);
not NOT1 (N3005, N3001);
nand NAND3 (N3006, N3000, N1174, N392);
buf BUF1 (N3007, N3004);
not NOT1 (N3008, N2992);
nand NAND2 (N3009, N2999, N973);
buf BUF1 (N3010, N2972);
and AND3 (N3011, N3008, N823, N3003);
not NOT1 (N3012, N2210);
buf BUF1 (N3013, N3006);
nor NOR4 (N3014, N3002, N970, N766, N2489);
nor NOR3 (N3015, N3014, N513, N2225);
or OR2 (N3016, N3013, N2152);
xor XOR2 (N3017, N3016, N1839);
nand NAND2 (N3018, N3005, N2006);
buf BUF1 (N3019, N3009);
not NOT1 (N3020, N2994);
and AND2 (N3021, N3019, N1391);
nor NOR4 (N3022, N3007, N1767, N2760, N1238);
not NOT1 (N3023, N3020);
buf BUF1 (N3024, N3010);
buf BUF1 (N3025, N3021);
nand NAND2 (N3026, N3025, N2572);
xor XOR2 (N3027, N3024, N371);
and AND3 (N3028, N3023, N2079, N2475);
or OR4 (N3029, N3027, N1144, N1013, N407);
buf BUF1 (N3030, N3011);
or OR2 (N3031, N3026, N2149);
nor NOR3 (N3032, N3029, N150, N2540);
xor XOR2 (N3033, N3022, N2059);
nor NOR4 (N3034, N3031, N708, N2375, N9);
xor XOR2 (N3035, N3018, N2343);
nand NAND3 (N3036, N3015, N2140, N732);
and AND4 (N3037, N3032, N1636, N848, N348);
buf BUF1 (N3038, N2990);
buf BUF1 (N3039, N3037);
nor NOR4 (N3040, N3030, N871, N1222, N1239);
nor NOR4 (N3041, N3028, N493, N2497, N2636);
nand NAND2 (N3042, N3033, N582);
and AND3 (N3043, N3041, N60, N1511);
buf BUF1 (N3044, N3035);
nand NAND3 (N3045, N3034, N235, N2452);
and AND4 (N3046, N3012, N2421, N2437, N1667);
or OR2 (N3047, N3040, N2577);
buf BUF1 (N3048, N3039);
and AND2 (N3049, N3046, N2124);
not NOT1 (N3050, N3036);
nand NAND4 (N3051, N3047, N2978, N1389, N556);
or OR4 (N3052, N3038, N841, N2257, N2945);
or OR2 (N3053, N3052, N2691);
not NOT1 (N3054, N3049);
xor XOR2 (N3055, N3050, N2438);
nand NAND3 (N3056, N3053, N1136, N2477);
or OR3 (N3057, N3051, N2078, N1454);
not NOT1 (N3058, N3044);
or OR2 (N3059, N3055, N2108);
nand NAND4 (N3060, N3017, N51, N1175, N1269);
and AND3 (N3061, N3042, N104, N1168);
or OR3 (N3062, N3059, N2173, N941);
or OR2 (N3063, N3054, N3039);
nor NOR3 (N3064, N3057, N2613, N1039);
xor XOR2 (N3065, N3045, N1288);
not NOT1 (N3066, N3063);
xor XOR2 (N3067, N3065, N2207);
buf BUF1 (N3068, N3056);
nand NAND3 (N3069, N3066, N2123, N2485);
and AND2 (N3070, N3058, N836);
or OR2 (N3071, N3060, N2054);
nor NOR4 (N3072, N3067, N49, N902, N1910);
xor XOR2 (N3073, N3071, N2605);
nor NOR3 (N3074, N3061, N2664, N1985);
xor XOR2 (N3075, N3043, N352);
not NOT1 (N3076, N3072);
nand NAND2 (N3077, N3074, N2790);
buf BUF1 (N3078, N3068);
and AND4 (N3079, N3073, N583, N2489, N32);
nor NOR4 (N3080, N3076, N2349, N1742, N794);
and AND3 (N3081, N3075, N1473, N1377);
and AND4 (N3082, N3062, N1757, N2722, N1240);
or OR3 (N3083, N3077, N2225, N561);
or OR2 (N3084, N3081, N1354);
nand NAND2 (N3085, N3078, N479);
not NOT1 (N3086, N3064);
nor NOR3 (N3087, N3080, N509, N2976);
or OR3 (N3088, N3087, N2842, N2558);
xor XOR2 (N3089, N3070, N1544);
not NOT1 (N3090, N3048);
buf BUF1 (N3091, N3088);
or OR4 (N3092, N3085, N2811, N2847, N1900);
or OR2 (N3093, N3092, N1436);
or OR2 (N3094, N3086, N2496);
buf BUF1 (N3095, N3090);
nand NAND4 (N3096, N3084, N926, N400, N2324);
and AND2 (N3097, N3079, N221);
xor XOR2 (N3098, N3082, N311);
xor XOR2 (N3099, N3069, N2654);
xor XOR2 (N3100, N3098, N944);
not NOT1 (N3101, N3094);
xor XOR2 (N3102, N3091, N2018);
xor XOR2 (N3103, N3099, N3088);
or OR4 (N3104, N3103, N3082, N1709, N2616);
buf BUF1 (N3105, N3102);
xor XOR2 (N3106, N3101, N2612);
and AND4 (N3107, N3089, N1828, N267, N1446);
xor XOR2 (N3108, N3093, N1970);
nor NOR4 (N3109, N3108, N803, N2137, N2784);
and AND4 (N3110, N3100, N2931, N349, N2427);
or OR3 (N3111, N3110, N157, N2832);
nand NAND2 (N3112, N3111, N3064);
xor XOR2 (N3113, N3107, N541);
or OR3 (N3114, N3113, N1499, N1118);
buf BUF1 (N3115, N3106);
nand NAND2 (N3116, N3104, N3055);
buf BUF1 (N3117, N3096);
not NOT1 (N3118, N3116);
xor XOR2 (N3119, N3114, N359);
nand NAND4 (N3120, N3097, N1736, N2860, N2836);
and AND2 (N3121, N3105, N1906);
nand NAND3 (N3122, N3118, N2552, N100);
or OR3 (N3123, N3117, N506, N711);
xor XOR2 (N3124, N3123, N59);
xor XOR2 (N3125, N3095, N1186);
not NOT1 (N3126, N3122);
nand NAND4 (N3127, N3109, N2940, N1305, N1104);
not NOT1 (N3128, N3115);
xor XOR2 (N3129, N3119, N990);
or OR4 (N3130, N3129, N445, N20, N1285);
nand NAND3 (N3131, N3112, N2220, N201);
nor NOR4 (N3132, N3130, N395, N1925, N2555);
xor XOR2 (N3133, N3124, N2302);
xor XOR2 (N3134, N3132, N2363);
and AND3 (N3135, N3127, N418, N1525);
xor XOR2 (N3136, N3131, N2284);
not NOT1 (N3137, N3125);
buf BUF1 (N3138, N3133);
nor NOR2 (N3139, N3138, N1089);
xor XOR2 (N3140, N3128, N2444);
buf BUF1 (N3141, N3140);
and AND2 (N3142, N3121, N1328);
buf BUF1 (N3143, N3137);
and AND4 (N3144, N3136, N2999, N1333, N1931);
nand NAND3 (N3145, N3143, N2963, N1208);
nor NOR2 (N3146, N3135, N2041);
nor NOR2 (N3147, N3142, N1850);
or OR3 (N3148, N3134, N2545, N3105);
or OR3 (N3149, N3145, N925, N2741);
xor XOR2 (N3150, N3144, N2436);
and AND3 (N3151, N3147, N1342, N401);
xor XOR2 (N3152, N3126, N2290);
nor NOR2 (N3153, N3152, N1851);
nor NOR3 (N3154, N3148, N1011, N1884);
nand NAND4 (N3155, N3139, N1707, N3119, N1780);
buf BUF1 (N3156, N3083);
or OR4 (N3157, N3151, N2649, N1803, N2628);
nand NAND4 (N3158, N3153, N2993, N1972, N2476);
xor XOR2 (N3159, N3158, N1117);
nor NOR3 (N3160, N3141, N2992, N1527);
not NOT1 (N3161, N3160);
buf BUF1 (N3162, N3149);
xor XOR2 (N3163, N3154, N2639);
or OR4 (N3164, N3157, N2007, N726, N2427);
xor XOR2 (N3165, N3164, N202);
nand NAND2 (N3166, N3155, N1174);
nand NAND4 (N3167, N3150, N2682, N319, N1845);
or OR2 (N3168, N3167, N1995);
xor XOR2 (N3169, N3159, N2556);
nand NAND2 (N3170, N3166, N2229);
or OR2 (N3171, N3165, N2222);
and AND2 (N3172, N3169, N3076);
not NOT1 (N3173, N3156);
buf BUF1 (N3174, N3171);
nor NOR4 (N3175, N3168, N869, N1032, N2032);
xor XOR2 (N3176, N3120, N1614);
nand NAND4 (N3177, N3161, N584, N2652, N2158);
buf BUF1 (N3178, N3173);
and AND4 (N3179, N3162, N1064, N2783, N828);
nand NAND2 (N3180, N3179, N379);
nor NOR2 (N3181, N3176, N1751);
buf BUF1 (N3182, N3181);
and AND2 (N3183, N3177, N272);
and AND2 (N3184, N3182, N2078);
not NOT1 (N3185, N3172);
not NOT1 (N3186, N3178);
nand NAND2 (N3187, N3175, N765);
or OR4 (N3188, N3187, N1782, N2274, N2638);
xor XOR2 (N3189, N3186, N531);
buf BUF1 (N3190, N3180);
not NOT1 (N3191, N3190);
xor XOR2 (N3192, N3183, N457);
nor NOR2 (N3193, N3191, N175);
or OR3 (N3194, N3192, N1213, N1810);
buf BUF1 (N3195, N3146);
nand NAND2 (N3196, N3185, N1300);
nand NAND4 (N3197, N3163, N889, N1750, N1812);
not NOT1 (N3198, N3193);
not NOT1 (N3199, N3195);
nand NAND3 (N3200, N3198, N2447, N182);
not NOT1 (N3201, N3197);
and AND3 (N3202, N3201, N669, N1342);
not NOT1 (N3203, N3170);
and AND4 (N3204, N3184, N1849, N1488, N282);
buf BUF1 (N3205, N3174);
not NOT1 (N3206, N3204);
xor XOR2 (N3207, N3194, N1774);
xor XOR2 (N3208, N3203, N1132);
and AND2 (N3209, N3199, N1336);
not NOT1 (N3210, N3200);
nand NAND4 (N3211, N3206, N977, N325, N2526);
not NOT1 (N3212, N3202);
not NOT1 (N3213, N3209);
buf BUF1 (N3214, N3210);
and AND4 (N3215, N3212, N2027, N2739, N437);
or OR2 (N3216, N3207, N1136);
not NOT1 (N3217, N3196);
xor XOR2 (N3218, N3217, N2400);
nor NOR3 (N3219, N3208, N2715, N1475);
xor XOR2 (N3220, N3219, N188);
and AND2 (N3221, N3215, N458);
not NOT1 (N3222, N3211);
and AND3 (N3223, N3218, N761, N2739);
and AND4 (N3224, N3214, N423, N351, N92);
nor NOR2 (N3225, N3205, N2021);
not NOT1 (N3226, N3221);
nor NOR3 (N3227, N3213, N3207, N717);
and AND2 (N3228, N3188, N1190);
not NOT1 (N3229, N3223);
nor NOR4 (N3230, N3222, N996, N309, N3070);
buf BUF1 (N3231, N3224);
not NOT1 (N3232, N3230);
not NOT1 (N3233, N3225);
buf BUF1 (N3234, N3231);
or OR4 (N3235, N3227, N1291, N1189, N485);
or OR4 (N3236, N3216, N1648, N1008, N2203);
not NOT1 (N3237, N3236);
nand NAND3 (N3238, N3228, N2264, N2915);
xor XOR2 (N3239, N3235, N174);
or OR2 (N3240, N3189, N2083);
or OR3 (N3241, N3229, N2550, N1366);
or OR4 (N3242, N3232, N257, N1216, N191);
not NOT1 (N3243, N3234);
buf BUF1 (N3244, N3238);
nand NAND3 (N3245, N3242, N3140, N2921);
not NOT1 (N3246, N3245);
buf BUF1 (N3247, N3241);
or OR3 (N3248, N3237, N1784, N604);
xor XOR2 (N3249, N3246, N2338);
or OR4 (N3250, N3244, N1887, N3069, N3158);
nor NOR2 (N3251, N3247, N2613);
buf BUF1 (N3252, N3239);
buf BUF1 (N3253, N3220);
not NOT1 (N3254, N3233);
nor NOR2 (N3255, N3240, N2361);
not NOT1 (N3256, N3243);
nor NOR3 (N3257, N3252, N2900, N1659);
and AND4 (N3258, N3256, N2623, N399, N1685);
and AND3 (N3259, N3249, N3048, N1218);
or OR2 (N3260, N3248, N1437);
and AND4 (N3261, N3226, N2089, N468, N102);
buf BUF1 (N3262, N3257);
nand NAND2 (N3263, N3261, N2825);
not NOT1 (N3264, N3262);
nand NAND3 (N3265, N3255, N1330, N102);
not NOT1 (N3266, N3254);
xor XOR2 (N3267, N3250, N682);
buf BUF1 (N3268, N3260);
not NOT1 (N3269, N3266);
xor XOR2 (N3270, N3269, N118);
buf BUF1 (N3271, N3268);
nand NAND3 (N3272, N3259, N1731, N1710);
and AND2 (N3273, N3265, N2091);
buf BUF1 (N3274, N3270);
xor XOR2 (N3275, N3273, N1379);
not NOT1 (N3276, N3274);
and AND4 (N3277, N3258, N2024, N1098, N111);
nand NAND4 (N3278, N3253, N229, N488, N2220);
not NOT1 (N3279, N3264);
buf BUF1 (N3280, N3277);
xor XOR2 (N3281, N3279, N524);
nand NAND4 (N3282, N3278, N2688, N2996, N2565);
xor XOR2 (N3283, N3272, N1267);
xor XOR2 (N3284, N3267, N1148);
buf BUF1 (N3285, N3263);
buf BUF1 (N3286, N3281);
nor NOR3 (N3287, N3283, N1320, N1301);
nor NOR3 (N3288, N3251, N416, N72);
or OR2 (N3289, N3287, N1214);
or OR3 (N3290, N3271, N113, N2391);
or OR3 (N3291, N3290, N413, N102);
or OR3 (N3292, N3282, N2641, N2895);
and AND4 (N3293, N3286, N2971, N2551, N480);
and AND3 (N3294, N3276, N1815, N1179);
xor XOR2 (N3295, N3280, N1510);
nand NAND3 (N3296, N3295, N486, N2773);
nand NAND4 (N3297, N3293, N1403, N181, N2263);
nand NAND4 (N3298, N3294, N70, N1084, N1855);
nor NOR3 (N3299, N3289, N2674, N2008);
and AND3 (N3300, N3288, N1744, N293);
and AND4 (N3301, N3291, N2102, N2623, N2645);
xor XOR2 (N3302, N3275, N2389);
not NOT1 (N3303, N3292);
xor XOR2 (N3304, N3303, N827);
xor XOR2 (N3305, N3298, N664);
and AND4 (N3306, N3285, N1866, N1709, N1913);
xor XOR2 (N3307, N3304, N2478);
and AND2 (N3308, N3307, N2733);
and AND3 (N3309, N3308, N514, N2451);
xor XOR2 (N3310, N3302, N1610);
or OR3 (N3311, N3284, N2654, N128);
xor XOR2 (N3312, N3296, N2457);
or OR3 (N3313, N3300, N2554, N1228);
nand NAND3 (N3314, N3310, N2369, N555);
nand NAND4 (N3315, N3312, N336, N1196, N810);
buf BUF1 (N3316, N3309);
buf BUF1 (N3317, N3313);
and AND2 (N3318, N3314, N1902);
xor XOR2 (N3319, N3297, N1235);
xor XOR2 (N3320, N3301, N490);
nor NOR4 (N3321, N3316, N1, N81, N1211);
nand NAND2 (N3322, N3311, N2449);
not NOT1 (N3323, N3319);
xor XOR2 (N3324, N3305, N2615);
not NOT1 (N3325, N3322);
xor XOR2 (N3326, N3324, N1516);
nor NOR4 (N3327, N3326, N1532, N1593, N2902);
nand NAND3 (N3328, N3317, N1283, N266);
nor NOR4 (N3329, N3328, N514, N2539, N536);
buf BUF1 (N3330, N3318);
and AND4 (N3331, N3323, N3260, N36, N1247);
nand NAND3 (N3332, N3299, N1605, N3008);
not NOT1 (N3333, N3325);
nand NAND3 (N3334, N3333, N1328, N1144);
or OR3 (N3335, N3332, N2887, N637);
xor XOR2 (N3336, N3335, N605);
and AND3 (N3337, N3330, N2757, N1486);
buf BUF1 (N3338, N3336);
buf BUF1 (N3339, N3315);
buf BUF1 (N3340, N3321);
not NOT1 (N3341, N3306);
xor XOR2 (N3342, N3320, N134);
or OR4 (N3343, N3340, N1218, N3322, N710);
nand NAND4 (N3344, N3331, N688, N2351, N570);
and AND3 (N3345, N3339, N2957, N2065);
not NOT1 (N3346, N3327);
nor NOR3 (N3347, N3343, N2144, N2058);
buf BUF1 (N3348, N3346);
nor NOR2 (N3349, N3338, N3081);
or OR3 (N3350, N3334, N2595, N28);
not NOT1 (N3351, N3329);
xor XOR2 (N3352, N3344, N1741);
and AND3 (N3353, N3348, N1414, N235);
xor XOR2 (N3354, N3342, N60);
xor XOR2 (N3355, N3349, N1763);
and AND3 (N3356, N3341, N33, N2041);
nand NAND3 (N3357, N3351, N2030, N2479);
nand NAND3 (N3358, N3345, N855, N2030);
or OR2 (N3359, N3357, N2115);
not NOT1 (N3360, N3337);
xor XOR2 (N3361, N3352, N1473);
nor NOR2 (N3362, N3359, N1040);
xor XOR2 (N3363, N3355, N2177);
nand NAND2 (N3364, N3347, N1256);
or OR4 (N3365, N3362, N2402, N3314, N2759);
xor XOR2 (N3366, N3358, N1674);
xor XOR2 (N3367, N3350, N1004);
and AND4 (N3368, N3354, N3077, N1242, N3354);
buf BUF1 (N3369, N3363);
nor NOR4 (N3370, N3360, N2231, N1369, N1351);
and AND2 (N3371, N3370, N3271);
nor NOR2 (N3372, N3353, N1593);
nand NAND4 (N3373, N3369, N937, N1338, N657);
and AND2 (N3374, N3368, N1350);
or OR3 (N3375, N3371, N1603, N2456);
buf BUF1 (N3376, N3373);
or OR4 (N3377, N3367, N1194, N3050, N2181);
not NOT1 (N3378, N3375);
nor NOR2 (N3379, N3365, N727);
and AND3 (N3380, N3378, N3312, N1433);
or OR4 (N3381, N3377, N1394, N2650, N2414);
xor XOR2 (N3382, N3364, N2963);
or OR3 (N3383, N3366, N1519, N1330);
nor NOR2 (N3384, N3356, N2269);
xor XOR2 (N3385, N3379, N3195);
buf BUF1 (N3386, N3380);
nand NAND2 (N3387, N3383, N12);
or OR4 (N3388, N3381, N828, N2982, N504);
or OR2 (N3389, N3372, N25);
or OR4 (N3390, N3385, N3111, N1477, N2950);
buf BUF1 (N3391, N3374);
and AND4 (N3392, N3361, N693, N2363, N1430);
or OR3 (N3393, N3384, N2579, N2261);
nor NOR2 (N3394, N3388, N1898);
not NOT1 (N3395, N3389);
nand NAND2 (N3396, N3390, N370);
buf BUF1 (N3397, N3387);
xor XOR2 (N3398, N3396, N2865);
nor NOR2 (N3399, N3386, N3049);
or OR4 (N3400, N3391, N967, N367, N3157);
xor XOR2 (N3401, N3399, N575);
buf BUF1 (N3402, N3400);
nor NOR2 (N3403, N3392, N385);
or OR2 (N3404, N3376, N1155);
nor NOR4 (N3405, N3382, N2329, N3121, N105);
buf BUF1 (N3406, N3402);
or OR4 (N3407, N3393, N950, N3250, N1681);
buf BUF1 (N3408, N3406);
nand NAND4 (N3409, N3397, N1659, N711, N695);
buf BUF1 (N3410, N3398);
nor NOR2 (N3411, N3405, N1731);
and AND4 (N3412, N3408, N316, N1635, N2319);
or OR3 (N3413, N3410, N1890, N737);
or OR2 (N3414, N3404, N2223);
and AND4 (N3415, N3407, N3296, N341, N1272);
and AND4 (N3416, N3412, N3113, N1864, N2116);
and AND4 (N3417, N3395, N2584, N905, N1559);
buf BUF1 (N3418, N3403);
nor NOR2 (N3419, N3415, N84);
or OR4 (N3420, N3414, N3270, N1373, N1184);
buf BUF1 (N3421, N3418);
and AND2 (N3422, N3401, N1078);
xor XOR2 (N3423, N3413, N527);
and AND4 (N3424, N3417, N3224, N637, N3132);
nor NOR4 (N3425, N3424, N1574, N2486, N2533);
nor NOR4 (N3426, N3416, N2243, N3048, N449);
nor NOR4 (N3427, N3425, N885, N1255, N2475);
nor NOR3 (N3428, N3419, N78, N2547);
nor NOR3 (N3429, N3409, N2501, N2666);
nor NOR2 (N3430, N3394, N2631);
buf BUF1 (N3431, N3422);
nor NOR2 (N3432, N3423, N337);
and AND3 (N3433, N3421, N3302, N2071);
and AND3 (N3434, N3430, N2257, N198);
and AND2 (N3435, N3426, N750);
nor NOR2 (N3436, N3420, N858);
xor XOR2 (N3437, N3429, N3038);
buf BUF1 (N3438, N3432);
nand NAND3 (N3439, N3428, N1051, N1858);
xor XOR2 (N3440, N3433, N1274);
or OR3 (N3441, N3434, N1696, N3379);
xor XOR2 (N3442, N3427, N1189);
and AND3 (N3443, N3437, N661, N1720);
nand NAND4 (N3444, N3431, N1072, N1529, N2116);
or OR4 (N3445, N3436, N1488, N3309, N3309);
nand NAND2 (N3446, N3441, N1736);
nand NAND4 (N3447, N3435, N1413, N1219, N1240);
xor XOR2 (N3448, N3440, N1660);
nor NOR3 (N3449, N3446, N1834, N342);
buf BUF1 (N3450, N3411);
or OR4 (N3451, N3444, N2282, N2988, N2000);
or OR3 (N3452, N3448, N3393, N1494);
xor XOR2 (N3453, N3438, N2500);
nand NAND4 (N3454, N3447, N3158, N1385, N3284);
xor XOR2 (N3455, N3443, N1896);
and AND3 (N3456, N3453, N179, N718);
and AND2 (N3457, N3449, N2508);
xor XOR2 (N3458, N3451, N2594);
nor NOR4 (N3459, N3458, N2992, N1762, N56);
nor NOR2 (N3460, N3456, N1294);
nand NAND2 (N3461, N3454, N1104);
buf BUF1 (N3462, N3442);
not NOT1 (N3463, N3445);
or OR3 (N3464, N3460, N2938, N1972);
and AND3 (N3465, N3439, N1694, N1993);
buf BUF1 (N3466, N3452);
xor XOR2 (N3467, N3465, N918);
and AND3 (N3468, N3462, N3295, N251);
not NOT1 (N3469, N3461);
and AND2 (N3470, N3464, N444);
not NOT1 (N3471, N3468);
not NOT1 (N3472, N3467);
nor NOR4 (N3473, N3455, N44, N588, N244);
buf BUF1 (N3474, N3463);
not NOT1 (N3475, N3471);
nand NAND2 (N3476, N3457, N3006);
nand NAND4 (N3477, N3472, N502, N403, N455);
buf BUF1 (N3478, N3477);
nand NAND2 (N3479, N3470, N827);
xor XOR2 (N3480, N3475, N662);
nor NOR3 (N3481, N3478, N1726, N1160);
or OR4 (N3482, N3481, N1651, N635, N715);
or OR3 (N3483, N3479, N2090, N1796);
not NOT1 (N3484, N3480);
nor NOR3 (N3485, N3476, N2937, N2300);
nand NAND2 (N3486, N3469, N2216);
xor XOR2 (N3487, N3486, N11);
buf BUF1 (N3488, N3482);
and AND4 (N3489, N3487, N2353, N2603, N2362);
not NOT1 (N3490, N3489);
or OR3 (N3491, N3473, N344, N857);
buf BUF1 (N3492, N3484);
and AND4 (N3493, N3483, N2147, N1340, N2011);
nor NOR2 (N3494, N3491, N1909);
xor XOR2 (N3495, N3485, N3479);
buf BUF1 (N3496, N3459);
xor XOR2 (N3497, N3490, N3337);
nand NAND4 (N3498, N3495, N2434, N3250, N620);
xor XOR2 (N3499, N3496, N2489);
buf BUF1 (N3500, N3498);
not NOT1 (N3501, N3466);
xor XOR2 (N3502, N3500, N348);
not NOT1 (N3503, N3474);
not NOT1 (N3504, N3493);
xor XOR2 (N3505, N3501, N2267);
nand NAND2 (N3506, N3504, N1306);
and AND3 (N3507, N3488, N2745, N2847);
not NOT1 (N3508, N3492);
nor NOR2 (N3509, N3450, N3212);
buf BUF1 (N3510, N3503);
xor XOR2 (N3511, N3509, N112);
or OR3 (N3512, N3499, N2631, N2748);
xor XOR2 (N3513, N3511, N2431);
xor XOR2 (N3514, N3510, N755);
endmodule