// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21;

output N2014,N2011,N2002,N2000,N2004,N2016,N2017,N2019,N1998,N2021;

buf BUF1 (N22, N17);
not NOT1 (N23, N1);
not NOT1 (N24, N22);
nor NOR2 (N25, N15, N1);
buf BUF1 (N26, N21);
nor NOR3 (N27, N24, N6, N2);
or OR4 (N28, N17, N26, N16, N27);
xor XOR2 (N29, N6, N10);
or OR2 (N30, N24, N21);
not NOT1 (N31, N9);
xor XOR2 (N32, N30, N28);
buf BUF1 (N33, N4);
or OR4 (N34, N12, N25, N29, N7);
or OR2 (N35, N8, N15);
nand NAND4 (N36, N27, N16, N27, N5);
xor XOR2 (N37, N6, N6);
xor XOR2 (N38, N21, N16);
buf BUF1 (N39, N30);
nor NOR4 (N40, N35, N37, N3, N4);
nand NAND2 (N41, N20, N32);
and AND4 (N42, N14, N28, N15, N32);
and AND2 (N43, N23, N14);
xor XOR2 (N44, N34, N16);
xor XOR2 (N45, N38, N37);
xor XOR2 (N46, N39, N42);
xor XOR2 (N47, N43, N14);
not NOT1 (N48, N46);
xor XOR2 (N49, N26, N26);
buf BUF1 (N50, N40);
nor NOR4 (N51, N44, N1, N29, N42);
or OR4 (N52, N47, N44, N44, N39);
and AND2 (N53, N41, N28);
nor NOR2 (N54, N36, N37);
nand NAND4 (N55, N50, N10, N4, N3);
not NOT1 (N56, N33);
nand NAND2 (N57, N55, N44);
not NOT1 (N58, N31);
nand NAND4 (N59, N57, N21, N10, N51);
and AND3 (N60, N26, N41, N22);
and AND3 (N61, N59, N38, N31);
not NOT1 (N62, N56);
or OR4 (N63, N60, N13, N3, N32);
not NOT1 (N64, N48);
buf BUF1 (N65, N49);
xor XOR2 (N66, N65, N19);
and AND4 (N67, N54, N26, N6, N36);
or OR3 (N68, N52, N38, N53);
buf BUF1 (N69, N47);
xor XOR2 (N70, N62, N8);
nor NOR3 (N71, N64, N20, N69);
xor XOR2 (N72, N24, N8);
buf BUF1 (N73, N58);
xor XOR2 (N74, N71, N5);
or OR3 (N75, N70, N19, N30);
xor XOR2 (N76, N66, N6);
nor NOR4 (N77, N61, N17, N62, N51);
not NOT1 (N78, N74);
nand NAND2 (N79, N45, N41);
nor NOR2 (N80, N75, N54);
nand NAND4 (N81, N78, N42, N40, N1);
not NOT1 (N82, N76);
nand NAND2 (N83, N80, N51);
buf BUF1 (N84, N68);
not NOT1 (N85, N81);
nor NOR4 (N86, N82, N51, N3, N62);
not NOT1 (N87, N83);
or OR2 (N88, N67, N46);
nor NOR3 (N89, N77, N80, N7);
not NOT1 (N90, N88);
nor NOR3 (N91, N79, N13, N72);
and AND2 (N92, N30, N26);
not NOT1 (N93, N73);
buf BUF1 (N94, N87);
nand NAND2 (N95, N92, N52);
buf BUF1 (N96, N93);
not NOT1 (N97, N95);
or OR3 (N98, N89, N40, N37);
nor NOR2 (N99, N96, N37);
nand NAND4 (N100, N84, N99, N77, N29);
buf BUF1 (N101, N13);
and AND2 (N102, N91, N97);
not NOT1 (N103, N88);
nor NOR3 (N104, N102, N32, N94);
buf BUF1 (N105, N64);
buf BUF1 (N106, N100);
nand NAND2 (N107, N105, N51);
xor XOR2 (N108, N63, N27);
nand NAND3 (N109, N106, N83, N24);
xor XOR2 (N110, N85, N27);
nand NAND3 (N111, N107, N81, N9);
nand NAND4 (N112, N86, N65, N106, N79);
and AND3 (N113, N103, N16, N26);
nor NOR3 (N114, N101, N111, N84);
not NOT1 (N115, N104);
and AND2 (N116, N113, N58);
nor NOR2 (N117, N81, N108);
or OR4 (N118, N36, N40, N96, N106);
buf BUF1 (N119, N118);
nor NOR4 (N120, N90, N87, N105, N114);
nor NOR2 (N121, N70, N106);
buf BUF1 (N122, N121);
and AND3 (N123, N122, N50, N38);
and AND3 (N124, N98, N107, N59);
and AND4 (N125, N116, N15, N45, N33);
xor XOR2 (N126, N112, N60);
not NOT1 (N127, N125);
nand NAND3 (N128, N109, N95, N35);
not NOT1 (N129, N117);
and AND4 (N130, N127, N104, N47, N121);
and AND2 (N131, N119, N127);
and AND2 (N132, N110, N61);
or OR3 (N133, N123, N45, N1);
xor XOR2 (N134, N128, N101);
buf BUF1 (N135, N120);
and AND3 (N136, N115, N110, N106);
buf BUF1 (N137, N126);
buf BUF1 (N138, N134);
nor NOR2 (N139, N131, N75);
buf BUF1 (N140, N130);
nor NOR4 (N141, N133, N134, N40, N135);
and AND4 (N142, N3, N121, N73, N76);
xor XOR2 (N143, N142, N70);
buf BUF1 (N144, N129);
xor XOR2 (N145, N143, N5);
or OR3 (N146, N144, N53, N38);
buf BUF1 (N147, N132);
buf BUF1 (N148, N124);
nor NOR2 (N149, N139, N137);
nand NAND4 (N150, N96, N140, N9, N133);
buf BUF1 (N151, N84);
or OR4 (N152, N151, N115, N19, N20);
buf BUF1 (N153, N138);
nor NOR2 (N154, N146, N16);
xor XOR2 (N155, N149, N60);
nand NAND4 (N156, N147, N59, N40, N154);
not NOT1 (N157, N154);
xor XOR2 (N158, N136, N18);
xor XOR2 (N159, N156, N93);
not NOT1 (N160, N150);
buf BUF1 (N161, N152);
nor NOR3 (N162, N157, N139, N66);
nor NOR3 (N163, N159, N136, N135);
or OR2 (N164, N145, N93);
nand NAND3 (N165, N153, N63, N83);
and AND3 (N166, N161, N128, N89);
and AND3 (N167, N141, N96, N155);
buf BUF1 (N168, N131);
xor XOR2 (N169, N163, N97);
xor XOR2 (N170, N165, N10);
or OR3 (N171, N167, N146, N123);
xor XOR2 (N172, N169, N153);
xor XOR2 (N173, N171, N128);
buf BUF1 (N174, N172);
or OR2 (N175, N168, N153);
and AND3 (N176, N148, N96, N35);
or OR3 (N177, N160, N16, N9);
not NOT1 (N178, N175);
buf BUF1 (N179, N158);
nor NOR4 (N180, N174, N144, N1, N103);
not NOT1 (N181, N180);
nor NOR2 (N182, N162, N165);
not NOT1 (N183, N176);
nor NOR3 (N184, N182, N68, N10);
not NOT1 (N185, N177);
nor NOR2 (N186, N166, N115);
nand NAND2 (N187, N164, N65);
buf BUF1 (N188, N179);
not NOT1 (N189, N181);
or OR2 (N190, N170, N112);
and AND3 (N191, N187, N132, N151);
nor NOR3 (N192, N185, N60, N116);
buf BUF1 (N193, N184);
and AND2 (N194, N186, N80);
buf BUF1 (N195, N188);
nor NOR2 (N196, N191, N149);
or OR3 (N197, N196, N71, N145);
and AND3 (N198, N183, N68, N26);
nor NOR3 (N199, N195, N100, N195);
not NOT1 (N200, N193);
xor XOR2 (N201, N199, N189);
not NOT1 (N202, N93);
and AND4 (N203, N197, N96, N22, N124);
xor XOR2 (N204, N192, N155);
or OR4 (N205, N178, N196, N201, N149);
and AND2 (N206, N149, N24);
nor NOR2 (N207, N204, N113);
xor XOR2 (N208, N198, N176);
nor NOR3 (N209, N202, N149, N57);
and AND2 (N210, N209, N146);
buf BUF1 (N211, N208);
nor NOR4 (N212, N205, N18, N142, N126);
nor NOR2 (N213, N203, N34);
nor NOR4 (N214, N206, N39, N26, N172);
nor NOR3 (N215, N200, N40, N107);
nand NAND4 (N216, N214, N176, N72, N95);
nand NAND4 (N217, N216, N118, N11, N105);
xor XOR2 (N218, N212, N191);
nor NOR2 (N219, N215, N25);
nor NOR3 (N220, N218, N206, N139);
not NOT1 (N221, N207);
or OR2 (N222, N220, N46);
buf BUF1 (N223, N217);
xor XOR2 (N224, N211, N181);
buf BUF1 (N225, N173);
or OR4 (N226, N225, N190, N201, N84);
nand NAND3 (N227, N58, N192, N47);
buf BUF1 (N228, N227);
buf BUF1 (N229, N224);
not NOT1 (N230, N226);
or OR2 (N231, N210, N52);
not NOT1 (N232, N213);
and AND2 (N233, N222, N225);
or OR3 (N234, N228, N121, N185);
or OR2 (N235, N221, N37);
xor XOR2 (N236, N223, N100);
not NOT1 (N237, N236);
not NOT1 (N238, N229);
buf BUF1 (N239, N235);
or OR3 (N240, N234, N151, N5);
nor NOR2 (N241, N230, N7);
buf BUF1 (N242, N240);
nor NOR3 (N243, N241, N143, N4);
nand NAND4 (N244, N237, N74, N22, N52);
or OR3 (N245, N219, N199, N190);
and AND3 (N246, N233, N121, N29);
or OR3 (N247, N238, N217, N168);
nand NAND3 (N248, N242, N148, N210);
or OR2 (N249, N245, N235);
buf BUF1 (N250, N243);
not NOT1 (N251, N250);
xor XOR2 (N252, N247, N44);
xor XOR2 (N253, N249, N5);
not NOT1 (N254, N248);
xor XOR2 (N255, N239, N39);
buf BUF1 (N256, N244);
nand NAND4 (N257, N252, N47, N112, N115);
and AND4 (N258, N257, N123, N5, N101);
nor NOR3 (N259, N253, N6, N32);
nand NAND3 (N260, N251, N159, N166);
nor NOR2 (N261, N259, N7);
nand NAND4 (N262, N246, N64, N52, N2);
and AND4 (N263, N255, N153, N50, N242);
and AND2 (N264, N262, N19);
nor NOR2 (N265, N194, N120);
xor XOR2 (N266, N261, N104);
buf BUF1 (N267, N260);
buf BUF1 (N268, N232);
nor NOR3 (N269, N268, N211, N13);
buf BUF1 (N270, N254);
or OR4 (N271, N270, N205, N92, N259);
xor XOR2 (N272, N267, N168);
not NOT1 (N273, N269);
nor NOR2 (N274, N258, N52);
or OR2 (N275, N274, N270);
not NOT1 (N276, N264);
not NOT1 (N277, N265);
and AND2 (N278, N263, N95);
nor NOR3 (N279, N276, N130, N248);
and AND3 (N280, N277, N55, N170);
nand NAND4 (N281, N272, N169, N47, N72);
xor XOR2 (N282, N275, N234);
nand NAND2 (N283, N279, N6);
and AND3 (N284, N271, N150, N70);
xor XOR2 (N285, N282, N114);
or OR2 (N286, N256, N275);
nand NAND4 (N287, N285, N49, N232, N199);
buf BUF1 (N288, N281);
not NOT1 (N289, N280);
nand NAND2 (N290, N283, N86);
not NOT1 (N291, N290);
and AND2 (N292, N278, N209);
nor NOR2 (N293, N288, N268);
xor XOR2 (N294, N292, N188);
not NOT1 (N295, N266);
nand NAND2 (N296, N293, N116);
xor XOR2 (N297, N286, N278);
xor XOR2 (N298, N296, N258);
buf BUF1 (N299, N273);
nor NOR2 (N300, N289, N148);
and AND4 (N301, N300, N228, N36, N4);
xor XOR2 (N302, N231, N73);
nand NAND3 (N303, N297, N176, N242);
nand NAND3 (N304, N284, N65, N93);
and AND2 (N305, N295, N220);
not NOT1 (N306, N287);
nor NOR2 (N307, N306, N288);
and AND3 (N308, N307, N250, N251);
nor NOR3 (N309, N308, N172, N135);
nor NOR2 (N310, N302, N279);
or OR3 (N311, N305, N291, N182);
not NOT1 (N312, N277);
or OR3 (N313, N303, N268, N172);
nor NOR2 (N314, N312, N101);
nand NAND3 (N315, N313, N145, N139);
buf BUF1 (N316, N315);
not NOT1 (N317, N301);
buf BUF1 (N318, N316);
nand NAND4 (N319, N309, N188, N125, N247);
xor XOR2 (N320, N311, N166);
xor XOR2 (N321, N319, N242);
and AND2 (N322, N320, N283);
or OR4 (N323, N304, N116, N142, N73);
or OR2 (N324, N314, N246);
or OR3 (N325, N317, N30, N10);
nand NAND4 (N326, N323, N152, N19, N54);
and AND2 (N327, N310, N168);
and AND2 (N328, N321, N22);
nor NOR3 (N329, N326, N41, N111);
not NOT1 (N330, N329);
not NOT1 (N331, N294);
nand NAND4 (N332, N327, N104, N35, N128);
buf BUF1 (N333, N299);
and AND2 (N334, N331, N170);
and AND3 (N335, N333, N170, N37);
nand NAND4 (N336, N328, N208, N310, N60);
and AND3 (N337, N325, N55, N64);
buf BUF1 (N338, N334);
nor NOR4 (N339, N337, N277, N128, N221);
not NOT1 (N340, N338);
or OR4 (N341, N324, N208, N93, N22);
nor NOR4 (N342, N330, N220, N275, N210);
not NOT1 (N343, N332);
nand NAND2 (N344, N343, N299);
xor XOR2 (N345, N342, N134);
buf BUF1 (N346, N345);
nand NAND2 (N347, N318, N238);
and AND2 (N348, N340, N80);
nor NOR4 (N349, N339, N150, N101, N167);
not NOT1 (N350, N341);
or OR3 (N351, N344, N257, N197);
nand NAND4 (N352, N348, N116, N172, N117);
and AND3 (N353, N347, N194, N135);
not NOT1 (N354, N346);
not NOT1 (N355, N350);
and AND4 (N356, N354, N17, N155, N67);
xor XOR2 (N357, N298, N76);
not NOT1 (N358, N335);
buf BUF1 (N359, N356);
or OR3 (N360, N352, N27, N195);
not NOT1 (N361, N357);
not NOT1 (N362, N358);
xor XOR2 (N363, N355, N279);
or OR3 (N364, N353, N328, N82);
nor NOR2 (N365, N362, N316);
nand NAND2 (N366, N359, N102);
xor XOR2 (N367, N365, N223);
and AND4 (N368, N366, N97, N299, N14);
nor NOR3 (N369, N367, N335, N264);
nand NAND2 (N370, N351, N9);
and AND3 (N371, N336, N345, N180);
not NOT1 (N372, N370);
not NOT1 (N373, N361);
nand NAND4 (N374, N364, N302, N12, N197);
or OR3 (N375, N373, N92, N14);
nor NOR2 (N376, N374, N158);
not NOT1 (N377, N376);
and AND2 (N378, N368, N362);
nor NOR4 (N379, N349, N163, N314, N340);
or OR2 (N380, N379, N343);
or OR4 (N381, N360, N24, N159, N60);
buf BUF1 (N382, N322);
not NOT1 (N383, N382);
nand NAND4 (N384, N378, N81, N82, N316);
xor XOR2 (N385, N371, N181);
not NOT1 (N386, N369);
nand NAND4 (N387, N372, N216, N88, N96);
buf BUF1 (N388, N377);
nor NOR3 (N389, N388, N186, N294);
nor NOR4 (N390, N385, N61, N115, N205);
nand NAND3 (N391, N380, N116, N109);
or OR4 (N392, N375, N338, N190, N243);
nand NAND4 (N393, N392, N262, N201, N264);
or OR4 (N394, N383, N171, N125, N86);
xor XOR2 (N395, N386, N101);
or OR3 (N396, N387, N195, N293);
or OR3 (N397, N391, N293, N343);
and AND4 (N398, N397, N226, N103, N350);
xor XOR2 (N399, N398, N132);
or OR4 (N400, N363, N235, N1, N132);
and AND3 (N401, N389, N296, N359);
xor XOR2 (N402, N394, N4);
nand NAND3 (N403, N393, N41, N117);
buf BUF1 (N404, N402);
and AND3 (N405, N381, N267, N251);
not NOT1 (N406, N384);
nand NAND3 (N407, N400, N159, N134);
not NOT1 (N408, N404);
buf BUF1 (N409, N405);
xor XOR2 (N410, N408, N300);
and AND3 (N411, N403, N68, N266);
and AND3 (N412, N401, N405, N353);
and AND4 (N413, N411, N30, N228, N246);
nand NAND2 (N414, N413, N376);
buf BUF1 (N415, N390);
nand NAND2 (N416, N399, N374);
nand NAND4 (N417, N395, N306, N45, N388);
not NOT1 (N418, N414);
xor XOR2 (N419, N410, N323);
nand NAND4 (N420, N417, N33, N15, N362);
nor NOR4 (N421, N420, N12, N195, N81);
and AND2 (N422, N421, N407);
nor NOR2 (N423, N169, N206);
nand NAND2 (N424, N422, N72);
not NOT1 (N425, N423);
not NOT1 (N426, N406);
or OR3 (N427, N418, N7, N250);
buf BUF1 (N428, N412);
nand NAND2 (N429, N425, N339);
xor XOR2 (N430, N426, N358);
and AND2 (N431, N409, N36);
nor NOR2 (N432, N424, N316);
buf BUF1 (N433, N431);
nor NOR4 (N434, N396, N208, N238, N112);
and AND2 (N435, N428, N350);
not NOT1 (N436, N419);
nor NOR2 (N437, N436, N277);
not NOT1 (N438, N435);
buf BUF1 (N439, N415);
nor NOR3 (N440, N430, N149, N257);
xor XOR2 (N441, N437, N417);
buf BUF1 (N442, N427);
xor XOR2 (N443, N429, N303);
nor NOR3 (N444, N434, N392, N155);
nand NAND3 (N445, N442, N165, N187);
xor XOR2 (N446, N432, N354);
nor NOR4 (N447, N441, N247, N81, N102);
nor NOR2 (N448, N433, N180);
xor XOR2 (N449, N438, N24);
nand NAND4 (N450, N447, N137, N112, N200);
nand NAND2 (N451, N448, N134);
nor NOR2 (N452, N451, N67);
nor NOR3 (N453, N416, N130, N402);
nor NOR4 (N454, N444, N441, N393, N230);
nand NAND3 (N455, N446, N93, N407);
nand NAND2 (N456, N453, N305);
buf BUF1 (N457, N439);
nor NOR2 (N458, N440, N221);
or OR3 (N459, N457, N76, N458);
nor NOR4 (N460, N225, N407, N53, N62);
buf BUF1 (N461, N449);
not NOT1 (N462, N455);
nand NAND4 (N463, N460, N188, N71, N22);
nand NAND2 (N464, N445, N88);
nor NOR2 (N465, N463, N20);
buf BUF1 (N466, N452);
not NOT1 (N467, N450);
xor XOR2 (N468, N462, N286);
or OR2 (N469, N467, N317);
or OR4 (N470, N466, N115, N324, N181);
or OR2 (N471, N464, N46);
or OR3 (N472, N469, N389, N110);
and AND3 (N473, N454, N169, N376);
nor NOR2 (N474, N465, N268);
or OR4 (N475, N456, N438, N49, N77);
and AND3 (N476, N459, N173, N17);
nand NAND3 (N477, N471, N116, N427);
nor NOR3 (N478, N477, N263, N67);
nor NOR3 (N479, N461, N39, N439);
and AND4 (N480, N474, N146, N187, N285);
buf BUF1 (N481, N443);
xor XOR2 (N482, N481, N154);
and AND2 (N483, N475, N390);
not NOT1 (N484, N470);
xor XOR2 (N485, N480, N151);
xor XOR2 (N486, N473, N354);
buf BUF1 (N487, N468);
or OR4 (N488, N487, N62, N261, N300);
not NOT1 (N489, N482);
and AND4 (N490, N489, N26, N139, N278);
buf BUF1 (N491, N476);
nand NAND4 (N492, N485, N376, N32, N9);
nand NAND4 (N493, N483, N64, N430, N289);
and AND4 (N494, N479, N432, N77, N325);
nor NOR4 (N495, N478, N236, N48, N198);
not NOT1 (N496, N491);
xor XOR2 (N497, N492, N158);
or OR2 (N498, N486, N381);
buf BUF1 (N499, N496);
xor XOR2 (N500, N472, N213);
not NOT1 (N501, N498);
buf BUF1 (N502, N494);
nand NAND3 (N503, N497, N82, N181);
xor XOR2 (N504, N490, N141);
xor XOR2 (N505, N499, N266);
or OR2 (N506, N484, N214);
and AND2 (N507, N504, N15);
and AND3 (N508, N502, N96, N79);
or OR3 (N509, N505, N462, N379);
nor NOR3 (N510, N493, N507, N325);
or OR2 (N511, N200, N415);
or OR4 (N512, N508, N411, N19, N183);
buf BUF1 (N513, N500);
or OR4 (N514, N488, N457, N96, N133);
buf BUF1 (N515, N511);
buf BUF1 (N516, N509);
nand NAND4 (N517, N516, N153, N458, N401);
nand NAND3 (N518, N514, N360, N460);
nand NAND3 (N519, N513, N34, N437);
nor NOR4 (N520, N515, N475, N512, N137);
xor XOR2 (N521, N406, N73);
nand NAND4 (N522, N501, N112, N81, N177);
nor NOR2 (N523, N519, N186);
and AND4 (N524, N510, N294, N471, N209);
and AND3 (N525, N495, N259, N134);
and AND3 (N526, N523, N100, N207);
nand NAND3 (N527, N503, N133, N461);
nor NOR2 (N528, N527, N380);
or OR3 (N529, N524, N279, N72);
not NOT1 (N530, N518);
not NOT1 (N531, N521);
not NOT1 (N532, N528);
and AND4 (N533, N526, N469, N106, N209);
not NOT1 (N534, N529);
nor NOR4 (N535, N520, N214, N242, N188);
nand NAND2 (N536, N534, N168);
nand NAND3 (N537, N535, N418, N483);
not NOT1 (N538, N537);
not NOT1 (N539, N522);
nor NOR3 (N540, N539, N210, N457);
nor NOR2 (N541, N506, N448);
buf BUF1 (N542, N531);
and AND3 (N543, N541, N152, N542);
nand NAND2 (N544, N88, N123);
not NOT1 (N545, N544);
xor XOR2 (N546, N533, N274);
xor XOR2 (N547, N543, N90);
nor NOR4 (N548, N545, N485, N199, N408);
not NOT1 (N549, N538);
buf BUF1 (N550, N548);
or OR3 (N551, N546, N434, N502);
not NOT1 (N552, N550);
nand NAND2 (N553, N540, N62);
and AND3 (N554, N517, N232, N144);
nor NOR2 (N555, N536, N506);
not NOT1 (N556, N552);
nor NOR3 (N557, N555, N451, N143);
not NOT1 (N558, N554);
nand NAND2 (N559, N557, N46);
nand NAND2 (N560, N559, N445);
xor XOR2 (N561, N532, N144);
or OR4 (N562, N560, N442, N405, N326);
and AND2 (N563, N547, N245);
buf BUF1 (N564, N525);
buf BUF1 (N565, N551);
xor XOR2 (N566, N558, N515);
or OR3 (N567, N564, N174, N226);
buf BUF1 (N568, N530);
xor XOR2 (N569, N567, N143);
buf BUF1 (N570, N565);
nand NAND2 (N571, N561, N472);
nor NOR2 (N572, N562, N392);
nand NAND2 (N573, N556, N153);
xor XOR2 (N574, N573, N16);
buf BUF1 (N575, N571);
buf BUF1 (N576, N572);
and AND3 (N577, N568, N434, N366);
xor XOR2 (N578, N577, N135);
xor XOR2 (N579, N553, N320);
or OR3 (N580, N578, N277, N47);
and AND2 (N581, N570, N566);
and AND3 (N582, N314, N19, N397);
and AND3 (N583, N576, N409, N498);
xor XOR2 (N584, N549, N6);
nor NOR4 (N585, N563, N449, N174, N351);
or OR3 (N586, N585, N381, N86);
xor XOR2 (N587, N583, N571);
nand NAND2 (N588, N584, N315);
nand NAND4 (N589, N579, N148, N163, N364);
and AND3 (N590, N588, N121, N394);
not NOT1 (N591, N582);
xor XOR2 (N592, N586, N37);
nand NAND2 (N593, N590, N99);
or OR4 (N594, N589, N10, N42, N123);
and AND3 (N595, N581, N314, N390);
nor NOR4 (N596, N580, N516, N96, N553);
or OR2 (N597, N594, N241);
nand NAND2 (N598, N574, N192);
or OR2 (N599, N596, N280);
xor XOR2 (N600, N598, N331);
nor NOR2 (N601, N575, N389);
or OR2 (N602, N600, N141);
nor NOR3 (N603, N569, N496, N371);
not NOT1 (N604, N597);
or OR2 (N605, N599, N502);
buf BUF1 (N606, N601);
or OR3 (N607, N602, N526, N533);
nor NOR4 (N608, N606, N35, N9, N281);
and AND4 (N609, N607, N155, N563, N293);
and AND4 (N610, N591, N2, N502, N54);
nor NOR3 (N611, N610, N109, N230);
or OR4 (N612, N608, N372, N10, N195);
or OR3 (N613, N587, N220, N547);
buf BUF1 (N614, N593);
xor XOR2 (N615, N613, N456);
nand NAND3 (N616, N605, N452, N581);
or OR3 (N617, N609, N497, N190);
nor NOR4 (N618, N614, N423, N153, N232);
xor XOR2 (N619, N616, N394);
xor XOR2 (N620, N619, N522);
nor NOR2 (N621, N603, N409);
xor XOR2 (N622, N618, N134);
xor XOR2 (N623, N611, N36);
buf BUF1 (N624, N612);
nand NAND2 (N625, N617, N283);
xor XOR2 (N626, N624, N584);
buf BUF1 (N627, N615);
xor XOR2 (N628, N621, N520);
and AND4 (N629, N623, N386, N360, N225);
nand NAND4 (N630, N627, N292, N164, N468);
not NOT1 (N631, N628);
xor XOR2 (N632, N592, N194);
and AND3 (N633, N620, N205, N110);
buf BUF1 (N634, N633);
buf BUF1 (N635, N625);
xor XOR2 (N636, N626, N179);
nand NAND4 (N637, N634, N519, N29, N490);
xor XOR2 (N638, N631, N495);
buf BUF1 (N639, N622);
nor NOR3 (N640, N629, N136, N33);
buf BUF1 (N641, N638);
and AND3 (N642, N630, N588, N42);
or OR3 (N643, N604, N470, N374);
nand NAND2 (N644, N640, N360);
or OR3 (N645, N632, N16, N387);
or OR3 (N646, N643, N539, N523);
or OR2 (N647, N646, N551);
buf BUF1 (N648, N645);
nand NAND2 (N649, N644, N409);
nor NOR4 (N650, N639, N444, N130, N160);
buf BUF1 (N651, N648);
buf BUF1 (N652, N650);
not NOT1 (N653, N642);
buf BUF1 (N654, N647);
and AND3 (N655, N651, N257, N537);
xor XOR2 (N656, N637, N109);
xor XOR2 (N657, N655, N526);
xor XOR2 (N658, N649, N488);
buf BUF1 (N659, N641);
and AND3 (N660, N654, N347, N451);
not NOT1 (N661, N635);
buf BUF1 (N662, N595);
and AND4 (N663, N636, N174, N491, N661);
xor XOR2 (N664, N144, N215);
and AND4 (N665, N662, N369, N148, N320);
or OR2 (N666, N660, N566);
and AND3 (N667, N666, N370, N46);
and AND4 (N668, N652, N346, N202, N76);
and AND2 (N669, N658, N225);
nand NAND3 (N670, N656, N139, N509);
and AND3 (N671, N669, N445, N666);
xor XOR2 (N672, N653, N381);
xor XOR2 (N673, N672, N211);
and AND3 (N674, N659, N256, N104);
buf BUF1 (N675, N663);
nor NOR4 (N676, N664, N471, N599, N271);
xor XOR2 (N677, N674, N443);
nand NAND2 (N678, N675, N647);
and AND4 (N679, N665, N39, N518, N26);
or OR2 (N680, N667, N647);
xor XOR2 (N681, N668, N99);
nand NAND2 (N682, N678, N625);
buf BUF1 (N683, N670);
or OR4 (N684, N680, N137, N201, N507);
xor XOR2 (N685, N677, N98);
nand NAND2 (N686, N683, N659);
not NOT1 (N687, N679);
or OR4 (N688, N673, N622, N224, N263);
not NOT1 (N689, N687);
xor XOR2 (N690, N657, N556);
buf BUF1 (N691, N676);
and AND2 (N692, N684, N291);
nor NOR2 (N693, N688, N513);
not NOT1 (N694, N686);
xor XOR2 (N695, N692, N566);
and AND2 (N696, N694, N429);
buf BUF1 (N697, N682);
and AND2 (N698, N689, N276);
xor XOR2 (N699, N685, N362);
xor XOR2 (N700, N699, N111);
nor NOR4 (N701, N696, N357, N322, N453);
and AND4 (N702, N671, N261, N112, N111);
buf BUF1 (N703, N690);
and AND3 (N704, N695, N316, N667);
not NOT1 (N705, N681);
xor XOR2 (N706, N703, N599);
xor XOR2 (N707, N691, N200);
xor XOR2 (N708, N707, N164);
nor NOR4 (N709, N698, N237, N418, N431);
or OR2 (N710, N702, N397);
and AND2 (N711, N705, N61);
xor XOR2 (N712, N701, N71);
and AND4 (N713, N700, N49, N645, N520);
nor NOR3 (N714, N712, N637, N445);
or OR2 (N715, N693, N314);
or OR2 (N716, N708, N440);
xor XOR2 (N717, N697, N444);
not NOT1 (N718, N714);
not NOT1 (N719, N710);
and AND4 (N720, N704, N106, N646, N367);
xor XOR2 (N721, N715, N698);
or OR2 (N722, N709, N82);
buf BUF1 (N723, N719);
or OR3 (N724, N706, N532, N400);
and AND3 (N725, N723, N288, N402);
nor NOR2 (N726, N720, N583);
nand NAND4 (N727, N724, N325, N341, N714);
buf BUF1 (N728, N725);
nor NOR2 (N729, N717, N525);
nor NOR2 (N730, N722, N499);
buf BUF1 (N731, N726);
xor XOR2 (N732, N727, N590);
or OR3 (N733, N711, N519, N430);
nand NAND3 (N734, N716, N265, N568);
buf BUF1 (N735, N713);
or OR2 (N736, N729, N311);
nand NAND4 (N737, N718, N478, N491, N507);
nand NAND3 (N738, N721, N535, N554);
or OR2 (N739, N732, N99);
or OR4 (N740, N734, N739, N497, N1);
nand NAND2 (N741, N625, N466);
xor XOR2 (N742, N731, N577);
nor NOR3 (N743, N740, N586, N220);
buf BUF1 (N744, N741);
not NOT1 (N745, N737);
or OR3 (N746, N738, N185, N635);
nor NOR4 (N747, N745, N621, N724, N463);
nor NOR2 (N748, N728, N28);
not NOT1 (N749, N742);
or OR2 (N750, N736, N290);
not NOT1 (N751, N747);
xor XOR2 (N752, N748, N633);
or OR2 (N753, N730, N229);
or OR3 (N754, N733, N77, N67);
nor NOR3 (N755, N735, N135, N402);
or OR4 (N756, N749, N639, N114, N606);
nor NOR2 (N757, N756, N94);
xor XOR2 (N758, N757, N316);
and AND2 (N759, N758, N403);
nand NAND2 (N760, N752, N659);
xor XOR2 (N761, N751, N341);
nand NAND2 (N762, N753, N345);
and AND4 (N763, N755, N270, N227, N431);
nor NOR4 (N764, N744, N693, N724, N246);
or OR3 (N765, N761, N102, N168);
or OR4 (N766, N754, N589, N179, N554);
xor XOR2 (N767, N762, N719);
or OR2 (N768, N746, N153);
and AND2 (N769, N764, N10);
and AND2 (N770, N769, N158);
not NOT1 (N771, N743);
or OR2 (N772, N763, N238);
nand NAND4 (N773, N770, N182, N692, N442);
or OR3 (N774, N760, N358, N623);
buf BUF1 (N775, N772);
or OR4 (N776, N775, N257, N212, N673);
nor NOR4 (N777, N776, N324, N226, N574);
or OR4 (N778, N768, N348, N292, N238);
or OR3 (N779, N771, N316, N523);
not NOT1 (N780, N767);
nand NAND2 (N781, N780, N370);
nand NAND2 (N782, N759, N571);
xor XOR2 (N783, N774, N622);
and AND2 (N784, N781, N430);
xor XOR2 (N785, N783, N696);
nand NAND4 (N786, N765, N348, N46, N137);
not NOT1 (N787, N786);
not NOT1 (N788, N777);
and AND2 (N789, N773, N341);
or OR2 (N790, N750, N785);
not NOT1 (N791, N496);
xor XOR2 (N792, N778, N355);
not NOT1 (N793, N766);
or OR2 (N794, N788, N159);
or OR3 (N795, N787, N232, N423);
or OR3 (N796, N791, N264, N195);
buf BUF1 (N797, N790);
or OR4 (N798, N795, N583, N23, N496);
or OR3 (N799, N798, N655, N700);
not NOT1 (N800, N793);
buf BUF1 (N801, N800);
buf BUF1 (N802, N784);
nor NOR2 (N803, N779, N454);
not NOT1 (N804, N799);
or OR4 (N805, N782, N441, N237, N54);
not NOT1 (N806, N803);
xor XOR2 (N807, N794, N387);
not NOT1 (N808, N805);
not NOT1 (N809, N802);
xor XOR2 (N810, N809, N737);
xor XOR2 (N811, N804, N581);
xor XOR2 (N812, N796, N794);
nor NOR4 (N813, N807, N343, N288, N419);
buf BUF1 (N814, N810);
nor NOR4 (N815, N808, N317, N335, N796);
or OR3 (N816, N792, N15, N289);
not NOT1 (N817, N811);
buf BUF1 (N818, N817);
buf BUF1 (N819, N801);
or OR4 (N820, N813, N568, N815, N267);
xor XOR2 (N821, N412, N153);
xor XOR2 (N822, N814, N48);
buf BUF1 (N823, N820);
or OR3 (N824, N819, N714, N32);
not NOT1 (N825, N823);
or OR4 (N826, N806, N489, N492, N24);
nand NAND4 (N827, N797, N400, N36, N478);
nand NAND3 (N828, N822, N747, N6);
nand NAND2 (N829, N827, N166);
and AND3 (N830, N825, N238, N97);
nand NAND2 (N831, N816, N285);
not NOT1 (N832, N812);
not NOT1 (N833, N824);
not NOT1 (N834, N826);
nor NOR3 (N835, N831, N581, N563);
xor XOR2 (N836, N835, N504);
not NOT1 (N837, N830);
not NOT1 (N838, N789);
not NOT1 (N839, N832);
xor XOR2 (N840, N829, N296);
buf BUF1 (N841, N828);
and AND4 (N842, N841, N442, N240, N197);
or OR3 (N843, N818, N454, N601);
or OR3 (N844, N834, N662, N649);
or OR2 (N845, N843, N211);
nor NOR4 (N846, N837, N649, N498, N73);
buf BUF1 (N847, N833);
or OR2 (N848, N836, N727);
nor NOR3 (N849, N845, N555, N680);
buf BUF1 (N850, N848);
nor NOR2 (N851, N840, N42);
nand NAND3 (N852, N849, N101, N286);
and AND4 (N853, N850, N506, N48, N22);
or OR3 (N854, N821, N77, N40);
not NOT1 (N855, N853);
not NOT1 (N856, N839);
xor XOR2 (N857, N855, N354);
nor NOR2 (N858, N857, N524);
not NOT1 (N859, N847);
buf BUF1 (N860, N842);
and AND3 (N861, N852, N502, N259);
buf BUF1 (N862, N858);
nand NAND2 (N863, N838, N132);
buf BUF1 (N864, N862);
not NOT1 (N865, N863);
nand NAND2 (N866, N844, N853);
not NOT1 (N867, N856);
nor NOR2 (N868, N851, N463);
buf BUF1 (N869, N866);
not NOT1 (N870, N854);
and AND3 (N871, N864, N566, N216);
nor NOR3 (N872, N869, N456, N503);
or OR2 (N873, N865, N137);
nor NOR3 (N874, N871, N385, N349);
and AND4 (N875, N874, N753, N414, N548);
nand NAND3 (N876, N868, N650, N72);
or OR3 (N877, N876, N39, N827);
xor XOR2 (N878, N870, N58);
nand NAND2 (N879, N872, N84);
nand NAND4 (N880, N873, N716, N262, N285);
and AND3 (N881, N860, N230, N643);
buf BUF1 (N882, N877);
buf BUF1 (N883, N878);
buf BUF1 (N884, N875);
buf BUF1 (N885, N880);
or OR4 (N886, N846, N731, N369, N389);
or OR3 (N887, N886, N47, N389);
or OR4 (N888, N883, N277, N690, N504);
nand NAND3 (N889, N888, N3, N335);
not NOT1 (N890, N867);
and AND3 (N891, N884, N174, N526);
buf BUF1 (N892, N879);
xor XOR2 (N893, N885, N832);
nor NOR3 (N894, N887, N470, N23);
not NOT1 (N895, N889);
not NOT1 (N896, N891);
or OR3 (N897, N892, N889, N19);
nor NOR2 (N898, N896, N452);
or OR3 (N899, N893, N447, N851);
nand NAND4 (N900, N897, N615, N365, N365);
and AND4 (N901, N859, N200, N498, N161);
or OR4 (N902, N882, N490, N445, N95);
or OR2 (N903, N902, N506);
nor NOR2 (N904, N901, N592);
not NOT1 (N905, N900);
xor XOR2 (N906, N890, N153);
xor XOR2 (N907, N903, N293);
nor NOR2 (N908, N898, N270);
nor NOR2 (N909, N904, N837);
or OR3 (N910, N895, N387, N550);
xor XOR2 (N911, N899, N152);
not NOT1 (N912, N894);
nor NOR3 (N913, N906, N633, N849);
nor NOR4 (N914, N907, N490, N738, N354);
nand NAND2 (N915, N909, N63);
buf BUF1 (N916, N908);
and AND3 (N917, N913, N13, N700);
buf BUF1 (N918, N912);
xor XOR2 (N919, N861, N476);
or OR2 (N920, N919, N758);
xor XOR2 (N921, N914, N674);
and AND2 (N922, N915, N304);
or OR2 (N923, N920, N159);
nand NAND4 (N924, N910, N618, N772, N501);
or OR2 (N925, N916, N779);
buf BUF1 (N926, N921);
not NOT1 (N927, N918);
xor XOR2 (N928, N917, N617);
nand NAND4 (N929, N905, N80, N866, N254);
xor XOR2 (N930, N925, N457);
xor XOR2 (N931, N929, N65);
buf BUF1 (N932, N923);
and AND3 (N933, N931, N154, N478);
nand NAND3 (N934, N922, N114, N101);
xor XOR2 (N935, N932, N877);
nand NAND4 (N936, N881, N254, N406, N209);
nand NAND3 (N937, N911, N583, N197);
or OR3 (N938, N936, N420, N377);
nor NOR4 (N939, N926, N920, N514, N505);
or OR3 (N940, N934, N336, N560);
xor XOR2 (N941, N933, N766);
xor XOR2 (N942, N927, N337);
nor NOR3 (N943, N937, N646, N91);
or OR3 (N944, N924, N821, N1);
or OR2 (N945, N941, N827);
buf BUF1 (N946, N935);
or OR2 (N947, N942, N702);
not NOT1 (N948, N947);
buf BUF1 (N949, N938);
nor NOR3 (N950, N944, N46, N826);
nand NAND3 (N951, N943, N675, N842);
not NOT1 (N952, N939);
buf BUF1 (N953, N950);
and AND2 (N954, N940, N78);
nor NOR4 (N955, N953, N411, N246, N792);
not NOT1 (N956, N952);
or OR4 (N957, N949, N397, N904, N128);
or OR4 (N958, N930, N59, N746, N539);
xor XOR2 (N959, N954, N351);
nand NAND4 (N960, N945, N554, N164, N591);
not NOT1 (N961, N958);
and AND2 (N962, N956, N64);
and AND4 (N963, N959, N146, N490, N902);
and AND3 (N964, N948, N298, N523);
or OR3 (N965, N960, N867, N69);
xor XOR2 (N966, N957, N927);
nand NAND3 (N967, N963, N206, N436);
not NOT1 (N968, N951);
not NOT1 (N969, N955);
nand NAND4 (N970, N962, N534, N475, N500);
or OR3 (N971, N969, N762, N897);
nand NAND2 (N972, N967, N478);
and AND3 (N973, N966, N140, N537);
or OR2 (N974, N961, N378);
xor XOR2 (N975, N928, N381);
buf BUF1 (N976, N970);
not NOT1 (N977, N975);
nor NOR2 (N978, N968, N46);
xor XOR2 (N979, N976, N65);
not NOT1 (N980, N965);
or OR3 (N981, N978, N608, N957);
xor XOR2 (N982, N981, N466);
xor XOR2 (N983, N946, N375);
not NOT1 (N984, N964);
buf BUF1 (N985, N974);
nor NOR2 (N986, N973, N126);
not NOT1 (N987, N979);
nand NAND3 (N988, N985, N434, N792);
and AND4 (N989, N987, N37, N866, N687);
or OR3 (N990, N977, N332, N785);
buf BUF1 (N991, N982);
and AND3 (N992, N990, N759, N377);
and AND4 (N993, N972, N707, N473, N889);
or OR2 (N994, N980, N2);
and AND3 (N995, N983, N2, N473);
buf BUF1 (N996, N991);
nand NAND2 (N997, N988, N876);
nand NAND2 (N998, N984, N814);
and AND2 (N999, N986, N926);
not NOT1 (N1000, N999);
and AND2 (N1001, N995, N554);
or OR4 (N1002, N1000, N404, N571, N704);
buf BUF1 (N1003, N997);
nor NOR2 (N1004, N998, N956);
nand NAND2 (N1005, N996, N671);
nor NOR2 (N1006, N993, N226);
nand NAND2 (N1007, N994, N815);
not NOT1 (N1008, N971);
or OR3 (N1009, N1003, N191, N293);
and AND2 (N1010, N992, N199);
or OR4 (N1011, N1004, N769, N413, N110);
not NOT1 (N1012, N1011);
nor NOR2 (N1013, N1006, N993);
not NOT1 (N1014, N1001);
or OR3 (N1015, N1010, N257, N319);
nor NOR4 (N1016, N1008, N399, N157, N758);
or OR3 (N1017, N1015, N845, N579);
nor NOR4 (N1018, N1012, N407, N820, N714);
not NOT1 (N1019, N1002);
not NOT1 (N1020, N1019);
xor XOR2 (N1021, N1007, N793);
nand NAND4 (N1022, N989, N240, N699, N74);
xor XOR2 (N1023, N1020, N969);
and AND3 (N1024, N1017, N696, N159);
not NOT1 (N1025, N1009);
or OR2 (N1026, N1005, N248);
xor XOR2 (N1027, N1018, N57);
xor XOR2 (N1028, N1014, N185);
or OR3 (N1029, N1025, N988, N500);
not NOT1 (N1030, N1028);
nand NAND3 (N1031, N1024, N736, N768);
nor NOR2 (N1032, N1027, N668);
xor XOR2 (N1033, N1030, N422);
nor NOR4 (N1034, N1033, N785, N238, N529);
nand NAND3 (N1035, N1021, N782, N995);
and AND4 (N1036, N1016, N138, N25, N685);
or OR2 (N1037, N1022, N129);
and AND3 (N1038, N1037, N464, N69);
buf BUF1 (N1039, N1034);
nor NOR3 (N1040, N1029, N869, N536);
and AND3 (N1041, N1032, N252, N970);
nor NOR4 (N1042, N1026, N35, N130, N703);
xor XOR2 (N1043, N1023, N300);
nor NOR4 (N1044, N1031, N502, N219, N778);
nor NOR3 (N1045, N1038, N356, N707);
xor XOR2 (N1046, N1035, N1003);
and AND3 (N1047, N1036, N732, N969);
nand NAND2 (N1048, N1047, N212);
nand NAND3 (N1049, N1041, N1024, N956);
buf BUF1 (N1050, N1039);
buf BUF1 (N1051, N1049);
nor NOR4 (N1052, N1040, N443, N580, N632);
not NOT1 (N1053, N1048);
or OR2 (N1054, N1045, N99);
nand NAND2 (N1055, N1043, N572);
nor NOR4 (N1056, N1044, N270, N292, N27);
or OR4 (N1057, N1054, N923, N746, N690);
not NOT1 (N1058, N1051);
or OR3 (N1059, N1052, N308, N601);
and AND4 (N1060, N1058, N14, N1007, N455);
buf BUF1 (N1061, N1042);
or OR3 (N1062, N1055, N114, N465);
or OR4 (N1063, N1057, N416, N524, N735);
buf BUF1 (N1064, N1053);
not NOT1 (N1065, N1062);
buf BUF1 (N1066, N1046);
xor XOR2 (N1067, N1056, N784);
or OR4 (N1068, N1013, N16, N180, N612);
xor XOR2 (N1069, N1050, N909);
and AND4 (N1070, N1066, N5, N332, N520);
nor NOR2 (N1071, N1064, N555);
or OR2 (N1072, N1070, N531);
and AND2 (N1073, N1069, N869);
not NOT1 (N1074, N1065);
nand NAND3 (N1075, N1068, N331, N905);
nand NAND3 (N1076, N1071, N879, N1001);
not NOT1 (N1077, N1072);
or OR2 (N1078, N1077, N141);
buf BUF1 (N1079, N1074);
and AND2 (N1080, N1073, N730);
or OR3 (N1081, N1078, N84, N1038);
or OR2 (N1082, N1080, N409);
not NOT1 (N1083, N1082);
or OR4 (N1084, N1063, N17, N670, N76);
buf BUF1 (N1085, N1079);
or OR2 (N1086, N1085, N98);
or OR3 (N1087, N1081, N590, N742);
not NOT1 (N1088, N1067);
and AND4 (N1089, N1060, N194, N224, N702);
nand NAND3 (N1090, N1076, N288, N319);
or OR4 (N1091, N1084, N579, N716, N184);
nor NOR2 (N1092, N1061, N570);
nor NOR2 (N1093, N1075, N124);
not NOT1 (N1094, N1087);
or OR2 (N1095, N1092, N441);
nor NOR3 (N1096, N1093, N158, N154);
nor NOR3 (N1097, N1090, N308, N309);
nand NAND3 (N1098, N1095, N443, N677);
nand NAND2 (N1099, N1083, N866);
nor NOR2 (N1100, N1088, N347);
xor XOR2 (N1101, N1100, N747);
nor NOR2 (N1102, N1089, N404);
xor XOR2 (N1103, N1101, N777);
not NOT1 (N1104, N1086);
buf BUF1 (N1105, N1059);
and AND2 (N1106, N1091, N472);
nor NOR3 (N1107, N1098, N639, N255);
not NOT1 (N1108, N1103);
nand NAND4 (N1109, N1102, N771, N806, N39);
and AND3 (N1110, N1106, N1031, N533);
buf BUF1 (N1111, N1094);
not NOT1 (N1112, N1110);
buf BUF1 (N1113, N1096);
nand NAND3 (N1114, N1108, N585, N1074);
not NOT1 (N1115, N1109);
not NOT1 (N1116, N1105);
not NOT1 (N1117, N1112);
buf BUF1 (N1118, N1104);
and AND2 (N1119, N1117, N1022);
or OR2 (N1120, N1119, N735);
and AND3 (N1121, N1097, N534, N1096);
or OR4 (N1122, N1113, N145, N1045, N785);
buf BUF1 (N1123, N1121);
xor XOR2 (N1124, N1115, N973);
nor NOR2 (N1125, N1107, N772);
and AND3 (N1126, N1120, N478, N544);
xor XOR2 (N1127, N1118, N551);
buf BUF1 (N1128, N1127);
xor XOR2 (N1129, N1111, N15);
nor NOR3 (N1130, N1128, N449, N1126);
not NOT1 (N1131, N224);
not NOT1 (N1132, N1129);
and AND4 (N1133, N1132, N1106, N134, N375);
nand NAND2 (N1134, N1133, N976);
and AND4 (N1135, N1116, N286, N961, N725);
buf BUF1 (N1136, N1130);
nor NOR4 (N1137, N1114, N411, N1041, N82);
buf BUF1 (N1138, N1122);
not NOT1 (N1139, N1123);
nand NAND4 (N1140, N1135, N387, N668, N656);
nor NOR3 (N1141, N1124, N177, N44);
not NOT1 (N1142, N1141);
nor NOR2 (N1143, N1140, N560);
or OR4 (N1144, N1142, N1047, N1140, N224);
nor NOR3 (N1145, N1125, N785, N266);
and AND2 (N1146, N1099, N17);
nand NAND3 (N1147, N1134, N157, N584);
xor XOR2 (N1148, N1138, N36);
nand NAND2 (N1149, N1137, N1031);
not NOT1 (N1150, N1136);
buf BUF1 (N1151, N1150);
buf BUF1 (N1152, N1147);
xor XOR2 (N1153, N1148, N591);
buf BUF1 (N1154, N1149);
or OR4 (N1155, N1144, N734, N672, N270);
and AND4 (N1156, N1139, N453, N683, N348);
and AND3 (N1157, N1146, N725, N391);
not NOT1 (N1158, N1157);
nor NOR3 (N1159, N1156, N796, N969);
nor NOR3 (N1160, N1152, N819, N216);
and AND3 (N1161, N1159, N741, N647);
xor XOR2 (N1162, N1160, N723);
and AND2 (N1163, N1131, N673);
not NOT1 (N1164, N1162);
and AND3 (N1165, N1163, N799, N1021);
xor XOR2 (N1166, N1153, N16);
or OR4 (N1167, N1164, N1063, N108, N1097);
xor XOR2 (N1168, N1155, N1099);
and AND2 (N1169, N1168, N302);
nor NOR3 (N1170, N1165, N73, N184);
buf BUF1 (N1171, N1151);
buf BUF1 (N1172, N1169);
or OR2 (N1173, N1166, N500);
buf BUF1 (N1174, N1170);
or OR3 (N1175, N1145, N272, N608);
or OR4 (N1176, N1175, N701, N907, N979);
nand NAND4 (N1177, N1176, N454, N25, N1129);
nor NOR3 (N1178, N1143, N270, N92);
or OR3 (N1179, N1158, N234, N98);
buf BUF1 (N1180, N1172);
nor NOR4 (N1181, N1167, N746, N719, N535);
nor NOR2 (N1182, N1154, N227);
xor XOR2 (N1183, N1177, N1087);
not NOT1 (N1184, N1182);
nor NOR2 (N1185, N1184, N905);
not NOT1 (N1186, N1161);
nand NAND2 (N1187, N1178, N449);
not NOT1 (N1188, N1183);
or OR4 (N1189, N1187, N523, N61, N730);
not NOT1 (N1190, N1181);
nor NOR2 (N1191, N1189, N911);
and AND2 (N1192, N1173, N281);
nor NOR2 (N1193, N1180, N692);
nand NAND4 (N1194, N1171, N193, N318, N332);
nor NOR2 (N1195, N1179, N799);
or OR4 (N1196, N1191, N297, N448, N1102);
xor XOR2 (N1197, N1188, N64);
and AND3 (N1198, N1190, N897, N660);
buf BUF1 (N1199, N1197);
not NOT1 (N1200, N1193);
buf BUF1 (N1201, N1174);
nand NAND3 (N1202, N1199, N328, N439);
nand NAND3 (N1203, N1194, N1189, N717);
nor NOR4 (N1204, N1202, N227, N296, N1116);
nor NOR4 (N1205, N1185, N631, N248, N1163);
or OR2 (N1206, N1186, N1146);
buf BUF1 (N1207, N1198);
nor NOR2 (N1208, N1196, N727);
buf BUF1 (N1209, N1206);
nand NAND3 (N1210, N1205, N145, N480);
nand NAND2 (N1211, N1195, N350);
buf BUF1 (N1212, N1210);
nor NOR4 (N1213, N1211, N617, N264, N802);
nor NOR4 (N1214, N1201, N120, N152, N1102);
and AND4 (N1215, N1200, N437, N206, N211);
nand NAND2 (N1216, N1207, N461);
and AND2 (N1217, N1192, N711);
buf BUF1 (N1218, N1208);
not NOT1 (N1219, N1218);
and AND4 (N1220, N1203, N867, N270, N847);
nor NOR2 (N1221, N1209, N960);
or OR4 (N1222, N1213, N357, N466, N117);
not NOT1 (N1223, N1220);
not NOT1 (N1224, N1219);
nor NOR4 (N1225, N1221, N576, N1116, N654);
and AND3 (N1226, N1216, N552, N690);
buf BUF1 (N1227, N1223);
nand NAND2 (N1228, N1212, N599);
buf BUF1 (N1229, N1226);
nand NAND3 (N1230, N1204, N949, N1205);
xor XOR2 (N1231, N1214, N835);
nand NAND4 (N1232, N1228, N1056, N1011, N649);
or OR2 (N1233, N1230, N866);
xor XOR2 (N1234, N1232, N296);
xor XOR2 (N1235, N1233, N840);
or OR4 (N1236, N1217, N604, N230, N1087);
nor NOR2 (N1237, N1229, N947);
xor XOR2 (N1238, N1222, N423);
nand NAND3 (N1239, N1238, N859, N924);
and AND3 (N1240, N1237, N218, N202);
not NOT1 (N1241, N1240);
nor NOR2 (N1242, N1241, N73);
nand NAND4 (N1243, N1215, N606, N936, N1055);
nand NAND3 (N1244, N1243, N878, N852);
buf BUF1 (N1245, N1231);
xor XOR2 (N1246, N1236, N135);
buf BUF1 (N1247, N1234);
nor NOR4 (N1248, N1235, N930, N961, N438);
nand NAND4 (N1249, N1248, N1108, N794, N943);
nor NOR2 (N1250, N1247, N137);
nand NAND3 (N1251, N1224, N226, N65);
nand NAND3 (N1252, N1244, N1218, N1249);
nor NOR3 (N1253, N505, N968, N253);
or OR4 (N1254, N1245, N309, N808, N311);
nand NAND4 (N1255, N1225, N152, N438, N256);
nor NOR3 (N1256, N1242, N22, N465);
or OR2 (N1257, N1251, N406);
not NOT1 (N1258, N1239);
and AND4 (N1259, N1253, N6, N1156, N601);
nor NOR3 (N1260, N1250, N565, N309);
or OR4 (N1261, N1252, N1240, N566, N326);
nor NOR3 (N1262, N1261, N1118, N957);
or OR3 (N1263, N1246, N616, N476);
buf BUF1 (N1264, N1263);
not NOT1 (N1265, N1262);
nor NOR2 (N1266, N1255, N1251);
xor XOR2 (N1267, N1265, N1046);
xor XOR2 (N1268, N1267, N401);
nor NOR3 (N1269, N1259, N1235, N80);
nor NOR3 (N1270, N1227, N67, N868);
or OR3 (N1271, N1268, N1033, N956);
buf BUF1 (N1272, N1258);
xor XOR2 (N1273, N1270, N621);
or OR4 (N1274, N1273, N82, N1035, N114);
nand NAND4 (N1275, N1257, N1166, N683, N1111);
or OR2 (N1276, N1260, N659);
nor NOR3 (N1277, N1272, N431, N265);
and AND2 (N1278, N1266, N929);
buf BUF1 (N1279, N1275);
xor XOR2 (N1280, N1269, N628);
nand NAND2 (N1281, N1278, N474);
and AND2 (N1282, N1274, N810);
nor NOR3 (N1283, N1276, N319, N159);
nand NAND4 (N1284, N1280, N936, N549, N312);
xor XOR2 (N1285, N1281, N241);
not NOT1 (N1286, N1256);
or OR2 (N1287, N1279, N562);
or OR4 (N1288, N1283, N590, N1019, N1102);
nand NAND4 (N1289, N1288, N352, N422, N1187);
xor XOR2 (N1290, N1286, N642);
or OR3 (N1291, N1282, N832, N1290);
buf BUF1 (N1292, N177);
xor XOR2 (N1293, N1287, N346);
buf BUF1 (N1294, N1277);
nor NOR2 (N1295, N1293, N311);
nor NOR2 (N1296, N1295, N4);
nand NAND2 (N1297, N1285, N1005);
and AND4 (N1298, N1292, N466, N1113, N521);
and AND3 (N1299, N1291, N846, N197);
nand NAND3 (N1300, N1271, N1003, N982);
buf BUF1 (N1301, N1296);
or OR3 (N1302, N1284, N645, N746);
nor NOR2 (N1303, N1302, N641);
nor NOR3 (N1304, N1294, N1095, N506);
buf BUF1 (N1305, N1298);
buf BUF1 (N1306, N1264);
or OR4 (N1307, N1301, N530, N418, N693);
or OR3 (N1308, N1303, N110, N190);
or OR2 (N1309, N1299, N1137);
xor XOR2 (N1310, N1289, N830);
or OR4 (N1311, N1305, N1121, N398, N742);
xor XOR2 (N1312, N1254, N763);
xor XOR2 (N1313, N1300, N1289);
xor XOR2 (N1314, N1312, N73);
buf BUF1 (N1315, N1313);
buf BUF1 (N1316, N1309);
buf BUF1 (N1317, N1310);
buf BUF1 (N1318, N1308);
buf BUF1 (N1319, N1306);
xor XOR2 (N1320, N1319, N609);
buf BUF1 (N1321, N1304);
xor XOR2 (N1322, N1314, N386);
nor NOR2 (N1323, N1311, N648);
or OR3 (N1324, N1321, N923, N68);
and AND3 (N1325, N1320, N707, N646);
or OR3 (N1326, N1317, N629, N1283);
nand NAND4 (N1327, N1297, N1223, N61, N175);
or OR4 (N1328, N1325, N146, N763, N65);
and AND4 (N1329, N1322, N165, N135, N950);
or OR2 (N1330, N1327, N900);
nor NOR3 (N1331, N1326, N1120, N91);
and AND4 (N1332, N1315, N1117, N1076, N625);
nor NOR3 (N1333, N1324, N68, N407);
not NOT1 (N1334, N1331);
xor XOR2 (N1335, N1318, N774);
not NOT1 (N1336, N1329);
buf BUF1 (N1337, N1330);
nor NOR3 (N1338, N1316, N237, N1306);
xor XOR2 (N1339, N1323, N770);
xor XOR2 (N1340, N1338, N1075);
buf BUF1 (N1341, N1328);
and AND2 (N1342, N1333, N386);
or OR3 (N1343, N1335, N1207, N1215);
buf BUF1 (N1344, N1342);
nor NOR4 (N1345, N1339, N653, N1248, N557);
xor XOR2 (N1346, N1334, N154);
xor XOR2 (N1347, N1345, N692);
nor NOR2 (N1348, N1332, N456);
not NOT1 (N1349, N1340);
nor NOR2 (N1350, N1343, N1086);
buf BUF1 (N1351, N1344);
or OR3 (N1352, N1341, N535, N873);
or OR3 (N1353, N1336, N1334, N241);
and AND3 (N1354, N1351, N1128, N723);
not NOT1 (N1355, N1352);
buf BUF1 (N1356, N1354);
or OR4 (N1357, N1350, N263, N461, N759);
nor NOR3 (N1358, N1353, N882, N919);
nor NOR4 (N1359, N1307, N541, N850, N687);
xor XOR2 (N1360, N1358, N381);
nand NAND4 (N1361, N1346, N203, N318, N1278);
or OR4 (N1362, N1357, N712, N503, N1071);
not NOT1 (N1363, N1355);
and AND4 (N1364, N1359, N538, N603, N1103);
nand NAND3 (N1365, N1360, N1262, N736);
not NOT1 (N1366, N1348);
not NOT1 (N1367, N1337);
buf BUF1 (N1368, N1365);
buf BUF1 (N1369, N1368);
or OR2 (N1370, N1369, N1261);
buf BUF1 (N1371, N1361);
buf BUF1 (N1372, N1366);
nor NOR2 (N1373, N1367, N718);
and AND2 (N1374, N1373, N1098);
nor NOR3 (N1375, N1371, N124, N310);
nand NAND3 (N1376, N1347, N1063, N1116);
or OR3 (N1377, N1364, N797, N929);
xor XOR2 (N1378, N1376, N334);
nand NAND2 (N1379, N1363, N63);
or OR2 (N1380, N1377, N1280);
or OR4 (N1381, N1370, N850, N685, N181);
buf BUF1 (N1382, N1374);
xor XOR2 (N1383, N1382, N509);
nand NAND3 (N1384, N1372, N160, N406);
nor NOR2 (N1385, N1362, N475);
and AND2 (N1386, N1356, N984);
nor NOR4 (N1387, N1375, N1122, N1314, N1236);
xor XOR2 (N1388, N1379, N307);
xor XOR2 (N1389, N1385, N1254);
and AND2 (N1390, N1349, N162);
and AND2 (N1391, N1380, N561);
nor NOR4 (N1392, N1378, N11, N330, N884);
and AND3 (N1393, N1381, N122, N124);
xor XOR2 (N1394, N1388, N1115);
not NOT1 (N1395, N1390);
and AND3 (N1396, N1389, N1392, N5);
xor XOR2 (N1397, N41, N799);
xor XOR2 (N1398, N1394, N816);
not NOT1 (N1399, N1396);
nand NAND2 (N1400, N1397, N1330);
buf BUF1 (N1401, N1399);
buf BUF1 (N1402, N1383);
and AND3 (N1403, N1393, N98, N236);
not NOT1 (N1404, N1401);
nor NOR2 (N1405, N1403, N324);
or OR4 (N1406, N1405, N125, N80, N415);
not NOT1 (N1407, N1391);
nand NAND2 (N1408, N1386, N737);
nand NAND2 (N1409, N1407, N229);
nor NOR4 (N1410, N1402, N609, N366, N1322);
and AND2 (N1411, N1408, N415);
or OR2 (N1412, N1410, N845);
not NOT1 (N1413, N1406);
buf BUF1 (N1414, N1404);
xor XOR2 (N1415, N1384, N977);
or OR2 (N1416, N1412, N1077);
not NOT1 (N1417, N1395);
nor NOR2 (N1418, N1411, N1126);
xor XOR2 (N1419, N1409, N213);
nand NAND2 (N1420, N1416, N104);
buf BUF1 (N1421, N1398);
and AND4 (N1422, N1417, N682, N1049, N151);
nor NOR4 (N1423, N1422, N58, N800, N7);
xor XOR2 (N1424, N1420, N964);
or OR4 (N1425, N1414, N238, N879, N1337);
not NOT1 (N1426, N1418);
nand NAND4 (N1427, N1419, N1056, N1140, N1351);
nand NAND3 (N1428, N1387, N199, N1085);
not NOT1 (N1429, N1425);
not NOT1 (N1430, N1400);
and AND3 (N1431, N1423, N918, N1321);
and AND2 (N1432, N1421, N962);
xor XOR2 (N1433, N1428, N692);
nand NAND2 (N1434, N1429, N49);
nand NAND2 (N1435, N1431, N897);
xor XOR2 (N1436, N1426, N265);
nor NOR4 (N1437, N1432, N716, N301, N1337);
and AND4 (N1438, N1424, N454, N174, N813);
nand NAND3 (N1439, N1436, N284, N944);
and AND4 (N1440, N1434, N704, N788, N1065);
not NOT1 (N1441, N1440);
or OR2 (N1442, N1433, N620);
nand NAND2 (N1443, N1438, N1034);
buf BUF1 (N1444, N1443);
or OR3 (N1445, N1437, N1119, N519);
and AND2 (N1446, N1435, N1408);
and AND2 (N1447, N1445, N816);
buf BUF1 (N1448, N1427);
nor NOR4 (N1449, N1446, N1342, N116, N395);
or OR4 (N1450, N1449, N335, N701, N1051);
nor NOR3 (N1451, N1442, N10, N228);
buf BUF1 (N1452, N1413);
and AND2 (N1453, N1448, N10);
nor NOR3 (N1454, N1439, N433, N702);
or OR4 (N1455, N1430, N613, N764, N525);
nand NAND2 (N1456, N1450, N82);
nand NAND2 (N1457, N1447, N1034);
nor NOR2 (N1458, N1457, N1239);
nor NOR2 (N1459, N1452, N886);
not NOT1 (N1460, N1453);
buf BUF1 (N1461, N1455);
or OR2 (N1462, N1441, N1213);
nand NAND4 (N1463, N1444, N311, N487, N782);
xor XOR2 (N1464, N1458, N1445);
buf BUF1 (N1465, N1462);
and AND3 (N1466, N1459, N360, N1099);
and AND4 (N1467, N1463, N909, N1048, N730);
not NOT1 (N1468, N1464);
xor XOR2 (N1469, N1454, N877);
buf BUF1 (N1470, N1461);
or OR3 (N1471, N1470, N1183, N1080);
buf BUF1 (N1472, N1466);
nand NAND2 (N1473, N1472, N1392);
nand NAND3 (N1474, N1460, N984, N1140);
nand NAND2 (N1475, N1467, N1443);
xor XOR2 (N1476, N1451, N1075);
xor XOR2 (N1477, N1476, N1009);
nand NAND3 (N1478, N1456, N948, N1322);
not NOT1 (N1479, N1477);
not NOT1 (N1480, N1475);
nand NAND4 (N1481, N1465, N858, N591, N246);
nand NAND2 (N1482, N1473, N26);
nor NOR3 (N1483, N1415, N107, N183);
or OR3 (N1484, N1469, N909, N684);
not NOT1 (N1485, N1483);
buf BUF1 (N1486, N1482);
nand NAND4 (N1487, N1481, N1313, N759, N1464);
nor NOR4 (N1488, N1485, N1405, N1087, N779);
and AND4 (N1489, N1484, N341, N1286, N1202);
nand NAND2 (N1490, N1479, N1198);
nor NOR3 (N1491, N1487, N385, N1224);
nor NOR2 (N1492, N1468, N1307);
or OR4 (N1493, N1478, N851, N9, N932);
or OR2 (N1494, N1480, N346);
buf BUF1 (N1495, N1490);
and AND3 (N1496, N1489, N621, N697);
and AND4 (N1497, N1496, N616, N342, N855);
nand NAND3 (N1498, N1474, N166, N292);
xor XOR2 (N1499, N1497, N16);
and AND2 (N1500, N1499, N992);
buf BUF1 (N1501, N1491);
not NOT1 (N1502, N1501);
xor XOR2 (N1503, N1502, N832);
or OR4 (N1504, N1492, N1299, N1475, N405);
and AND3 (N1505, N1495, N1351, N236);
or OR4 (N1506, N1486, N980, N907, N308);
buf BUF1 (N1507, N1504);
nand NAND2 (N1508, N1505, N728);
and AND4 (N1509, N1493, N1314, N1237, N219);
or OR4 (N1510, N1471, N1283, N1451, N1314);
xor XOR2 (N1511, N1500, N470);
not NOT1 (N1512, N1488);
not NOT1 (N1513, N1511);
buf BUF1 (N1514, N1513);
or OR4 (N1515, N1509, N993, N1266, N381);
buf BUF1 (N1516, N1512);
nor NOR4 (N1517, N1510, N1078, N890, N1145);
nor NOR4 (N1518, N1517, N1032, N284, N1406);
nor NOR4 (N1519, N1503, N1083, N448, N777);
nor NOR4 (N1520, N1506, N1055, N1418, N260);
nand NAND2 (N1521, N1494, N960);
xor XOR2 (N1522, N1498, N21);
or OR4 (N1523, N1507, N505, N367, N1124);
and AND2 (N1524, N1518, N109);
and AND2 (N1525, N1524, N1254);
nor NOR3 (N1526, N1514, N1312, N690);
nand NAND4 (N1527, N1508, N1098, N1022, N1321);
and AND2 (N1528, N1523, N1070);
and AND2 (N1529, N1520, N339);
nor NOR3 (N1530, N1516, N499, N1172);
buf BUF1 (N1531, N1526);
and AND4 (N1532, N1525, N139, N683, N937);
xor XOR2 (N1533, N1529, N713);
nand NAND4 (N1534, N1515, N187, N826, N1264);
nor NOR2 (N1535, N1528, N883);
and AND4 (N1536, N1530, N705, N475, N803);
nor NOR3 (N1537, N1536, N1131, N1397);
and AND4 (N1538, N1527, N1460, N695, N182);
nor NOR2 (N1539, N1522, N946);
nand NAND4 (N1540, N1533, N464, N863, N499);
xor XOR2 (N1541, N1535, N295);
nand NAND2 (N1542, N1540, N137);
nand NAND3 (N1543, N1532, N1351, N547);
or OR4 (N1544, N1538, N1255, N632, N145);
buf BUF1 (N1545, N1534);
or OR4 (N1546, N1545, N59, N1323, N408);
and AND3 (N1547, N1546, N611, N384);
and AND3 (N1548, N1547, N714, N310);
nor NOR2 (N1549, N1531, N526);
not NOT1 (N1550, N1537);
nand NAND4 (N1551, N1548, N1188, N1230, N1175);
nand NAND3 (N1552, N1519, N1309, N1086);
or OR2 (N1553, N1521, N180);
or OR3 (N1554, N1553, N675, N1479);
buf BUF1 (N1555, N1542);
nand NAND3 (N1556, N1555, N1517, N616);
not NOT1 (N1557, N1554);
nand NAND4 (N1558, N1543, N628, N340, N842);
and AND4 (N1559, N1544, N203, N771, N291);
xor XOR2 (N1560, N1539, N326);
not NOT1 (N1561, N1558);
or OR3 (N1562, N1561, N256, N165);
or OR2 (N1563, N1556, N51);
and AND3 (N1564, N1562, N1185, N519);
buf BUF1 (N1565, N1559);
or OR4 (N1566, N1541, N92, N588, N412);
and AND4 (N1567, N1565, N1142, N552, N1257);
not NOT1 (N1568, N1557);
nand NAND3 (N1569, N1567, N1280, N199);
not NOT1 (N1570, N1550);
not NOT1 (N1571, N1570);
or OR3 (N1572, N1569, N256, N281);
buf BUF1 (N1573, N1564);
and AND3 (N1574, N1551, N78, N1053);
xor XOR2 (N1575, N1568, N399);
buf BUF1 (N1576, N1552);
or OR2 (N1577, N1573, N1340);
nand NAND4 (N1578, N1563, N459, N239, N998);
nor NOR3 (N1579, N1572, N236, N751);
not NOT1 (N1580, N1574);
buf BUF1 (N1581, N1576);
nand NAND4 (N1582, N1577, N391, N355, N1058);
and AND2 (N1583, N1579, N669);
xor XOR2 (N1584, N1580, N661);
xor XOR2 (N1585, N1560, N1403);
buf BUF1 (N1586, N1549);
nand NAND4 (N1587, N1583, N1198, N129, N1117);
or OR3 (N1588, N1571, N1291, N116);
not NOT1 (N1589, N1587);
not NOT1 (N1590, N1582);
or OR3 (N1591, N1581, N1264, N1499);
nor NOR4 (N1592, N1591, N856, N906, N1107);
buf BUF1 (N1593, N1578);
nor NOR4 (N1594, N1566, N1311, N668, N285);
and AND2 (N1595, N1575, N605);
nand NAND3 (N1596, N1588, N337, N342);
xor XOR2 (N1597, N1584, N1472);
or OR4 (N1598, N1590, N580, N1301, N446);
xor XOR2 (N1599, N1596, N371);
or OR4 (N1600, N1586, N484, N1577, N260);
xor XOR2 (N1601, N1597, N1316);
nor NOR2 (N1602, N1594, N893);
xor XOR2 (N1603, N1602, N1073);
xor XOR2 (N1604, N1598, N932);
or OR2 (N1605, N1604, N92);
or OR2 (N1606, N1592, N848);
not NOT1 (N1607, N1601);
or OR4 (N1608, N1585, N1215, N38, N935);
and AND4 (N1609, N1603, N1346, N1034, N184);
nor NOR3 (N1610, N1593, N510, N1580);
or OR2 (N1611, N1589, N1161);
and AND3 (N1612, N1611, N1332, N1139);
buf BUF1 (N1613, N1610);
and AND2 (N1614, N1607, N1516);
nor NOR2 (N1615, N1595, N493);
xor XOR2 (N1616, N1606, N1241);
not NOT1 (N1617, N1600);
xor XOR2 (N1618, N1609, N90);
not NOT1 (N1619, N1614);
xor XOR2 (N1620, N1616, N848);
buf BUF1 (N1621, N1599);
xor XOR2 (N1622, N1612, N1443);
not NOT1 (N1623, N1605);
buf BUF1 (N1624, N1620);
and AND2 (N1625, N1623, N1203);
nand NAND2 (N1626, N1608, N210);
nand NAND3 (N1627, N1617, N618, N79);
nand NAND4 (N1628, N1619, N1416, N1567, N1209);
xor XOR2 (N1629, N1615, N654);
xor XOR2 (N1630, N1626, N1082);
nor NOR3 (N1631, N1628, N936, N662);
buf BUF1 (N1632, N1625);
not NOT1 (N1633, N1630);
not NOT1 (N1634, N1631);
or OR2 (N1635, N1633, N1035);
xor XOR2 (N1636, N1629, N237);
xor XOR2 (N1637, N1613, N511);
not NOT1 (N1638, N1621);
buf BUF1 (N1639, N1618);
and AND4 (N1640, N1639, N330, N211, N382);
or OR4 (N1641, N1640, N490, N1358, N1136);
buf BUF1 (N1642, N1622);
not NOT1 (N1643, N1627);
nor NOR4 (N1644, N1632, N660, N1096, N116);
nand NAND3 (N1645, N1638, N246, N1383);
xor XOR2 (N1646, N1637, N111);
not NOT1 (N1647, N1645);
xor XOR2 (N1648, N1646, N902);
xor XOR2 (N1649, N1647, N1314);
and AND2 (N1650, N1635, N1352);
and AND4 (N1651, N1642, N466, N1397, N1202);
xor XOR2 (N1652, N1634, N258);
buf BUF1 (N1653, N1643);
nand NAND2 (N1654, N1652, N185);
xor XOR2 (N1655, N1644, N1128);
xor XOR2 (N1656, N1649, N1108);
not NOT1 (N1657, N1650);
buf BUF1 (N1658, N1651);
xor XOR2 (N1659, N1624, N180);
nand NAND2 (N1660, N1653, N973);
buf BUF1 (N1661, N1655);
nor NOR2 (N1662, N1657, N1438);
xor XOR2 (N1663, N1641, N1135);
xor XOR2 (N1664, N1659, N397);
not NOT1 (N1665, N1660);
xor XOR2 (N1666, N1654, N1664);
and AND3 (N1667, N1276, N248, N226);
xor XOR2 (N1668, N1665, N351);
or OR3 (N1669, N1648, N827, N1544);
not NOT1 (N1670, N1667);
nand NAND3 (N1671, N1662, N792, N1005);
xor XOR2 (N1672, N1636, N1488);
not NOT1 (N1673, N1656);
xor XOR2 (N1674, N1658, N958);
or OR4 (N1675, N1673, N1153, N598, N15);
nor NOR2 (N1676, N1671, N987);
buf BUF1 (N1677, N1676);
and AND4 (N1678, N1663, N1089, N1093, N1130);
nor NOR4 (N1679, N1668, N1516, N1186, N527);
nand NAND3 (N1680, N1674, N189, N1171);
or OR4 (N1681, N1679, N718, N1494, N1362);
buf BUF1 (N1682, N1677);
and AND3 (N1683, N1670, N1207, N688);
buf BUF1 (N1684, N1681);
nand NAND4 (N1685, N1661, N508, N602, N525);
not NOT1 (N1686, N1680);
nor NOR2 (N1687, N1678, N760);
nand NAND3 (N1688, N1683, N1500, N1585);
xor XOR2 (N1689, N1687, N1219);
and AND2 (N1690, N1686, N1074);
nand NAND2 (N1691, N1688, N827);
nand NAND4 (N1692, N1691, N1317, N1156, N1036);
and AND4 (N1693, N1689, N991, N16, N606);
and AND2 (N1694, N1675, N756);
xor XOR2 (N1695, N1684, N1153);
xor XOR2 (N1696, N1694, N134);
xor XOR2 (N1697, N1685, N1464);
not NOT1 (N1698, N1695);
buf BUF1 (N1699, N1672);
nor NOR3 (N1700, N1697, N338, N502);
not NOT1 (N1701, N1690);
not NOT1 (N1702, N1682);
not NOT1 (N1703, N1698);
buf BUF1 (N1704, N1700);
not NOT1 (N1705, N1666);
xor XOR2 (N1706, N1669, N186);
xor XOR2 (N1707, N1702, N1664);
and AND2 (N1708, N1699, N849);
nor NOR3 (N1709, N1704, N1155, N900);
and AND3 (N1710, N1696, N1077, N743);
nand NAND4 (N1711, N1703, N569, N1323, N504);
nor NOR3 (N1712, N1708, N486, N920);
or OR2 (N1713, N1705, N1395);
or OR4 (N1714, N1693, N1296, N712, N1386);
not NOT1 (N1715, N1713);
and AND3 (N1716, N1715, N1559, N486);
not NOT1 (N1717, N1710);
buf BUF1 (N1718, N1714);
nor NOR4 (N1719, N1711, N223, N1646, N1085);
buf BUF1 (N1720, N1701);
not NOT1 (N1721, N1717);
and AND3 (N1722, N1718, N1300, N1154);
and AND3 (N1723, N1709, N55, N421);
nand NAND4 (N1724, N1721, N1686, N449, N1444);
and AND2 (N1725, N1720, N1294);
or OR2 (N1726, N1712, N1121);
buf BUF1 (N1727, N1719);
buf BUF1 (N1728, N1692);
xor XOR2 (N1729, N1706, N612);
nor NOR3 (N1730, N1726, N865, N536);
xor XOR2 (N1731, N1724, N1672);
and AND2 (N1732, N1723, N1405);
not NOT1 (N1733, N1725);
nor NOR3 (N1734, N1730, N816, N616);
not NOT1 (N1735, N1728);
nand NAND3 (N1736, N1731, N907, N929);
nor NOR2 (N1737, N1727, N65);
xor XOR2 (N1738, N1735, N164);
not NOT1 (N1739, N1734);
and AND4 (N1740, N1729, N447, N407, N1064);
not NOT1 (N1741, N1740);
or OR4 (N1742, N1722, N1523, N1700, N638);
and AND3 (N1743, N1737, N181, N1719);
or OR4 (N1744, N1733, N716, N1320, N771);
nand NAND2 (N1745, N1739, N908);
or OR3 (N1746, N1736, N947, N1672);
and AND4 (N1747, N1707, N582, N621, N1550);
or OR3 (N1748, N1732, N962, N360);
and AND2 (N1749, N1741, N1359);
xor XOR2 (N1750, N1747, N765);
or OR3 (N1751, N1750, N1153, N359);
xor XOR2 (N1752, N1738, N564);
not NOT1 (N1753, N1748);
nor NOR3 (N1754, N1753, N1115, N1272);
or OR3 (N1755, N1754, N319, N1715);
buf BUF1 (N1756, N1742);
nand NAND2 (N1757, N1745, N936);
and AND4 (N1758, N1756, N1591, N792, N137);
buf BUF1 (N1759, N1752);
and AND4 (N1760, N1759, N1598, N1200, N1150);
not NOT1 (N1761, N1760);
and AND2 (N1762, N1716, N1408);
or OR2 (N1763, N1761, N1513);
buf BUF1 (N1764, N1757);
nand NAND4 (N1765, N1746, N1358, N228, N1140);
or OR3 (N1766, N1758, N924, N1039);
nor NOR3 (N1767, N1751, N865, N1728);
nor NOR4 (N1768, N1763, N154, N179, N98);
not NOT1 (N1769, N1749);
nor NOR2 (N1770, N1766, N36);
or OR2 (N1771, N1743, N564);
nor NOR2 (N1772, N1744, N558);
not NOT1 (N1773, N1770);
xor XOR2 (N1774, N1764, N872);
nor NOR3 (N1775, N1762, N1487, N1534);
nor NOR3 (N1776, N1767, N879, N611);
buf BUF1 (N1777, N1769);
nand NAND3 (N1778, N1771, N237, N1163);
not NOT1 (N1779, N1765);
not NOT1 (N1780, N1774);
and AND4 (N1781, N1779, N768, N1150, N1241);
and AND4 (N1782, N1780, N985, N1217, N300);
xor XOR2 (N1783, N1777, N857);
and AND2 (N1784, N1775, N1635);
not NOT1 (N1785, N1776);
and AND4 (N1786, N1784, N388, N1539, N1544);
not NOT1 (N1787, N1783);
nand NAND2 (N1788, N1772, N1539);
buf BUF1 (N1789, N1788);
buf BUF1 (N1790, N1789);
xor XOR2 (N1791, N1787, N172);
xor XOR2 (N1792, N1781, N826);
nand NAND3 (N1793, N1755, N656, N746);
not NOT1 (N1794, N1786);
not NOT1 (N1795, N1773);
nor NOR4 (N1796, N1785, N1571, N1761, N1568);
or OR3 (N1797, N1791, N514, N234);
buf BUF1 (N1798, N1778);
and AND4 (N1799, N1798, N100, N986, N1758);
not NOT1 (N1800, N1796);
not NOT1 (N1801, N1793);
buf BUF1 (N1802, N1792);
nor NOR2 (N1803, N1782, N566);
or OR2 (N1804, N1801, N550);
buf BUF1 (N1805, N1790);
buf BUF1 (N1806, N1804);
buf BUF1 (N1807, N1768);
nand NAND2 (N1808, N1795, N1554);
not NOT1 (N1809, N1805);
buf BUF1 (N1810, N1800);
not NOT1 (N1811, N1797);
and AND4 (N1812, N1799, N409, N106, N722);
xor XOR2 (N1813, N1810, N1708);
nand NAND2 (N1814, N1808, N1333);
not NOT1 (N1815, N1807);
not NOT1 (N1816, N1812);
nor NOR4 (N1817, N1814, N871, N1151, N569);
not NOT1 (N1818, N1815);
not NOT1 (N1819, N1803);
nor NOR2 (N1820, N1813, N1142);
or OR2 (N1821, N1818, N38);
buf BUF1 (N1822, N1794);
or OR3 (N1823, N1819, N1140, N372);
or OR4 (N1824, N1817, N753, N1195, N1115);
or OR2 (N1825, N1820, N105);
or OR2 (N1826, N1811, N250);
or OR4 (N1827, N1826, N1571, N1162, N719);
nor NOR4 (N1828, N1823, N1767, N1156, N1336);
not NOT1 (N1829, N1816);
xor XOR2 (N1830, N1829, N1679);
buf BUF1 (N1831, N1809);
and AND3 (N1832, N1806, N1463, N1426);
buf BUF1 (N1833, N1822);
not NOT1 (N1834, N1832);
or OR3 (N1835, N1825, N1738, N1628);
nor NOR3 (N1836, N1802, N744, N1079);
nor NOR3 (N1837, N1830, N755, N691);
xor XOR2 (N1838, N1828, N1789);
nor NOR4 (N1839, N1821, N1332, N1589, N844);
xor XOR2 (N1840, N1824, N770);
buf BUF1 (N1841, N1834);
and AND4 (N1842, N1841, N1505, N668, N34);
or OR3 (N1843, N1833, N262, N294);
nand NAND2 (N1844, N1842, N959);
or OR3 (N1845, N1831, N792, N1288);
nor NOR4 (N1846, N1839, N1414, N1343, N1226);
not NOT1 (N1847, N1846);
xor XOR2 (N1848, N1827, N380);
nor NOR3 (N1849, N1837, N843, N1441);
xor XOR2 (N1850, N1843, N135);
and AND4 (N1851, N1835, N387, N1479, N753);
nor NOR2 (N1852, N1849, N349);
xor XOR2 (N1853, N1838, N1639);
not NOT1 (N1854, N1850);
or OR3 (N1855, N1844, N446, N1476);
nor NOR4 (N1856, N1853, N224, N1400, N37);
not NOT1 (N1857, N1845);
or OR3 (N1858, N1855, N72, N1250);
or OR2 (N1859, N1857, N323);
nand NAND2 (N1860, N1859, N284);
not NOT1 (N1861, N1840);
nor NOR2 (N1862, N1848, N1785);
or OR3 (N1863, N1856, N1738, N472);
nor NOR3 (N1864, N1863, N1402, N222);
nand NAND4 (N1865, N1864, N1490, N878, N1851);
or OR4 (N1866, N388, N306, N1006, N1020);
xor XOR2 (N1867, N1862, N1450);
nand NAND3 (N1868, N1858, N1023, N532);
or OR2 (N1869, N1865, N1492);
nor NOR2 (N1870, N1852, N1327);
nor NOR4 (N1871, N1869, N31, N979, N644);
xor XOR2 (N1872, N1847, N748);
buf BUF1 (N1873, N1861);
not NOT1 (N1874, N1860);
xor XOR2 (N1875, N1836, N1102);
and AND4 (N1876, N1868, N1701, N1508, N1645);
buf BUF1 (N1877, N1874);
and AND4 (N1878, N1867, N1727, N1520, N385);
nor NOR2 (N1879, N1854, N1660);
or OR2 (N1880, N1875, N1489);
buf BUF1 (N1881, N1880);
and AND3 (N1882, N1870, N1255, N577);
buf BUF1 (N1883, N1873);
nand NAND3 (N1884, N1881, N1541, N1270);
nand NAND2 (N1885, N1872, N1829);
not NOT1 (N1886, N1885);
and AND3 (N1887, N1886, N1453, N1202);
or OR2 (N1888, N1876, N1381);
and AND4 (N1889, N1866, N649, N352, N1440);
nand NAND2 (N1890, N1887, N434);
not NOT1 (N1891, N1890);
not NOT1 (N1892, N1871);
nand NAND3 (N1893, N1878, N518, N443);
or OR3 (N1894, N1892, N135, N12);
nand NAND3 (N1895, N1888, N617, N1047);
and AND4 (N1896, N1882, N1771, N439, N309);
buf BUF1 (N1897, N1879);
or OR4 (N1898, N1895, N1136, N475, N1881);
and AND4 (N1899, N1889, N864, N712, N119);
xor XOR2 (N1900, N1877, N1398);
not NOT1 (N1901, N1893);
and AND2 (N1902, N1897, N370);
or OR3 (N1903, N1894, N1508, N1862);
nand NAND4 (N1904, N1896, N24, N1144, N1097);
buf BUF1 (N1905, N1899);
and AND4 (N1906, N1900, N917, N1316, N431);
xor XOR2 (N1907, N1904, N530);
not NOT1 (N1908, N1883);
not NOT1 (N1909, N1902);
nor NOR2 (N1910, N1884, N1345);
nor NOR4 (N1911, N1898, N1793, N1045, N586);
nor NOR2 (N1912, N1905, N1087);
nand NAND2 (N1913, N1910, N1781);
or OR3 (N1914, N1907, N1640, N1660);
nor NOR4 (N1915, N1908, N79, N1003, N518);
nor NOR2 (N1916, N1903, N80);
nand NAND2 (N1917, N1909, N701);
xor XOR2 (N1918, N1911, N1607);
xor XOR2 (N1919, N1916, N953);
nor NOR3 (N1920, N1915, N887, N672);
nand NAND4 (N1921, N1913, N1802, N736, N1355);
buf BUF1 (N1922, N1920);
or OR2 (N1923, N1917, N1605);
buf BUF1 (N1924, N1914);
xor XOR2 (N1925, N1921, N1423);
nand NAND2 (N1926, N1901, N950);
nand NAND4 (N1927, N1925, N1569, N346, N150);
nor NOR3 (N1928, N1919, N1636, N1047);
nor NOR2 (N1929, N1926, N557);
or OR2 (N1930, N1912, N726);
and AND3 (N1931, N1930, N233, N1850);
xor XOR2 (N1932, N1931, N1499);
nand NAND4 (N1933, N1923, N1459, N1476, N831);
buf BUF1 (N1934, N1927);
and AND2 (N1935, N1924, N1605);
not NOT1 (N1936, N1933);
and AND3 (N1937, N1929, N902, N1135);
buf BUF1 (N1938, N1922);
nor NOR4 (N1939, N1928, N141, N1011, N1130);
not NOT1 (N1940, N1918);
or OR2 (N1941, N1936, N462);
buf BUF1 (N1942, N1941);
buf BUF1 (N1943, N1939);
xor XOR2 (N1944, N1943, N1673);
not NOT1 (N1945, N1932);
nand NAND2 (N1946, N1937, N546);
or OR4 (N1947, N1938, N88, N1796, N1360);
and AND3 (N1948, N1942, N576, N1516);
and AND3 (N1949, N1906, N1457, N1517);
nor NOR2 (N1950, N1949, N782);
buf BUF1 (N1951, N1950);
nor NOR3 (N1952, N1940, N277, N975);
nand NAND4 (N1953, N1946, N1005, N179, N1383);
or OR4 (N1954, N1947, N1907, N591, N839);
buf BUF1 (N1955, N1952);
xor XOR2 (N1956, N1948, N1249);
and AND4 (N1957, N1955, N65, N1697, N1494);
xor XOR2 (N1958, N1935, N386);
buf BUF1 (N1959, N1891);
and AND2 (N1960, N1954, N1634);
or OR2 (N1961, N1959, N1366);
and AND4 (N1962, N1956, N523, N1014, N380);
buf BUF1 (N1963, N1945);
not NOT1 (N1964, N1951);
xor XOR2 (N1965, N1963, N531);
nor NOR3 (N1966, N1962, N616, N369);
buf BUF1 (N1967, N1934);
not NOT1 (N1968, N1966);
nor NOR4 (N1969, N1953, N454, N1014, N1963);
nand NAND2 (N1970, N1961, N1800);
not NOT1 (N1971, N1967);
not NOT1 (N1972, N1970);
and AND2 (N1973, N1960, N862);
not NOT1 (N1974, N1964);
or OR2 (N1975, N1957, N501);
and AND3 (N1976, N1974, N1970, N1459);
nand NAND4 (N1977, N1976, N1506, N870, N1921);
or OR3 (N1978, N1975, N382, N393);
nor NOR4 (N1979, N1944, N1760, N1203, N190);
xor XOR2 (N1980, N1978, N1599);
nor NOR4 (N1981, N1968, N1752, N1715, N171);
buf BUF1 (N1982, N1971);
not NOT1 (N1983, N1972);
xor XOR2 (N1984, N1980, N692);
and AND4 (N1985, N1958, N804, N1129, N1251);
or OR2 (N1986, N1979, N937);
nand NAND4 (N1987, N1984, N858, N748, N1271);
nand NAND4 (N1988, N1981, N859, N1420, N243);
nor NOR3 (N1989, N1977, N719, N1352);
not NOT1 (N1990, N1989);
and AND3 (N1991, N1965, N1237, N1548);
nand NAND3 (N1992, N1991, N1470, N520);
and AND3 (N1993, N1988, N1794, N1887);
nor NOR2 (N1994, N1990, N1472);
xor XOR2 (N1995, N1994, N1565);
buf BUF1 (N1996, N1973);
nand NAND2 (N1997, N1987, N881);
buf BUF1 (N1998, N1992);
not NOT1 (N1999, N1996);
buf BUF1 (N2000, N1999);
and AND3 (N2001, N1969, N1460, N1958);
xor XOR2 (N2002, N1997, N1909);
or OR2 (N2003, N1995, N465);
not NOT1 (N2004, N1982);
buf BUF1 (N2005, N1986);
not NOT1 (N2006, N1993);
or OR4 (N2007, N1983, N1352, N613, N307);
nor NOR2 (N2008, N2005, N1116);
buf BUF1 (N2009, N2008);
buf BUF1 (N2010, N2007);
or OR2 (N2011, N1985, N1793);
xor XOR2 (N2012, N2009, N1133);
or OR4 (N2013, N2010, N63, N1705, N418);
nor NOR2 (N2014, N2001, N1668);
and AND4 (N2015, N2006, N228, N469, N634);
buf BUF1 (N2016, N2015);
buf BUF1 (N2017, N2012);
xor XOR2 (N2018, N2003, N790);
xor XOR2 (N2019, N2018, N1077);
nor NOR3 (N2020, N2013, N1627, N1620);
buf BUF1 (N2021, N2020);
endmodule