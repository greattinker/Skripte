// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17;

output N12803,N12815,N12813,N12807,N12812,N12816,N12798,N12808,N12800,N12817;

and AND4 (N18, N15, N10, N10, N15);
not NOT1 (N19, N10);
nand NAND2 (N20, N9, N7);
and AND4 (N21, N11, N18, N17, N13);
nand NAND4 (N22, N9, N15, N15, N10);
nand NAND4 (N23, N17, N18, N11, N17);
not NOT1 (N24, N18);
not NOT1 (N25, N9);
nor NOR4 (N26, N19, N25, N2, N6);
not NOT1 (N27, N11);
nand NAND2 (N28, N24, N1);
xor XOR2 (N29, N4, N12);
not NOT1 (N30, N24);
or OR3 (N31, N1, N29, N6);
and AND3 (N32, N12, N31, N14);
not NOT1 (N33, N30);
xor XOR2 (N34, N6, N6);
buf BUF1 (N35, N28);
not NOT1 (N36, N33);
or OR2 (N37, N36, N23);
buf BUF1 (N38, N1);
nand NAND3 (N39, N27, N2, N17);
nor NOR3 (N40, N39, N39, N9);
not NOT1 (N41, N34);
xor XOR2 (N42, N32, N21);
nand NAND3 (N43, N21, N11, N37);
xor XOR2 (N44, N23, N42);
buf BUF1 (N45, N9);
and AND4 (N46, N20, N28, N5, N30);
or OR2 (N47, N38, N23);
xor XOR2 (N48, N45, N22);
nor NOR3 (N49, N32, N19, N4);
xor XOR2 (N50, N44, N7);
nor NOR4 (N51, N47, N17, N34, N41);
not NOT1 (N52, N20);
not NOT1 (N53, N35);
or OR2 (N54, N52, N19);
or OR3 (N55, N51, N14, N21);
or OR3 (N56, N49, N50, N37);
buf BUF1 (N57, N51);
nand NAND3 (N58, N48, N31, N9);
nor NOR3 (N59, N43, N41, N38);
or OR3 (N60, N59, N19, N9);
nand NAND3 (N61, N60, N54, N24);
nor NOR3 (N62, N31, N24, N30);
buf BUF1 (N63, N62);
nand NAND3 (N64, N56, N56, N35);
nand NAND4 (N65, N61, N5, N61, N53);
and AND3 (N66, N8, N37, N18);
buf BUF1 (N67, N57);
and AND3 (N68, N67, N14, N7);
not NOT1 (N69, N66);
xor XOR2 (N70, N40, N22);
not NOT1 (N71, N58);
nor NOR4 (N72, N69, N57, N43, N2);
nand NAND2 (N73, N65, N11);
or OR3 (N74, N68, N16, N7);
nand NAND4 (N75, N72, N16, N31, N54);
and AND2 (N76, N64, N13);
buf BUF1 (N77, N76);
buf BUF1 (N78, N71);
xor XOR2 (N79, N55, N64);
nor NOR3 (N80, N46, N42, N32);
and AND4 (N81, N78, N30, N33, N40);
nor NOR4 (N82, N81, N49, N72, N17);
nand NAND4 (N83, N77, N78, N72, N10);
xor XOR2 (N84, N82, N73);
and AND4 (N85, N39, N38, N41, N43);
or OR3 (N86, N75, N45, N72);
xor XOR2 (N87, N74, N13);
or OR3 (N88, N85, N15, N2);
not NOT1 (N89, N86);
not NOT1 (N90, N87);
xor XOR2 (N91, N90, N34);
and AND2 (N92, N63, N48);
xor XOR2 (N93, N79, N22);
nor NOR3 (N94, N80, N49, N83);
nor NOR4 (N95, N82, N25, N14, N2);
buf BUF1 (N96, N95);
and AND4 (N97, N89, N49, N90, N64);
xor XOR2 (N98, N91, N47);
nand NAND4 (N99, N97, N25, N24, N50);
and AND3 (N100, N93, N35, N76);
and AND2 (N101, N92, N98);
xor XOR2 (N102, N51, N24);
nand NAND2 (N103, N26, N22);
or OR4 (N104, N99, N6, N18, N47);
buf BUF1 (N105, N84);
or OR4 (N106, N96, N63, N64, N69);
nand NAND3 (N107, N104, N5, N56);
not NOT1 (N108, N103);
not NOT1 (N109, N101);
nor NOR3 (N110, N109, N63, N63);
not NOT1 (N111, N94);
and AND3 (N112, N111, N91, N79);
and AND3 (N113, N88, N45, N34);
and AND3 (N114, N112, N68, N98);
buf BUF1 (N115, N105);
and AND2 (N116, N102, N39);
buf BUF1 (N117, N115);
or OR4 (N118, N107, N103, N39, N15);
nor NOR2 (N119, N117, N116);
nor NOR4 (N120, N116, N90, N77, N101);
or OR4 (N121, N108, N34, N4, N78);
xor XOR2 (N122, N118, N74);
nand NAND2 (N123, N106, N72);
nor NOR3 (N124, N70, N103, N19);
buf BUF1 (N125, N124);
nand NAND2 (N126, N100, N17);
not NOT1 (N127, N121);
buf BUF1 (N128, N120);
nor NOR4 (N129, N114, N1, N84, N32);
xor XOR2 (N130, N125, N87);
not NOT1 (N131, N122);
not NOT1 (N132, N131);
and AND2 (N133, N123, N123);
nor NOR3 (N134, N132, N12, N25);
nor NOR4 (N135, N128, N116, N7, N53);
nand NAND2 (N136, N135, N63);
nor NOR2 (N137, N127, N101);
xor XOR2 (N138, N129, N40);
not NOT1 (N139, N137);
nor NOR2 (N140, N110, N43);
nand NAND2 (N141, N126, N76);
not NOT1 (N142, N138);
xor XOR2 (N143, N130, N2);
buf BUF1 (N144, N142);
and AND2 (N145, N133, N53);
or OR2 (N146, N143, N81);
xor XOR2 (N147, N146, N54);
xor XOR2 (N148, N136, N40);
not NOT1 (N149, N147);
xor XOR2 (N150, N145, N109);
nand NAND3 (N151, N141, N19, N74);
or OR2 (N152, N134, N2);
not NOT1 (N153, N139);
xor XOR2 (N154, N119, N132);
not NOT1 (N155, N154);
not NOT1 (N156, N148);
buf BUF1 (N157, N152);
not NOT1 (N158, N153);
nand NAND4 (N159, N150, N52, N84, N64);
nand NAND4 (N160, N159, N149, N151, N1);
or OR3 (N161, N49, N66, N37);
buf BUF1 (N162, N120);
nor NOR2 (N163, N157, N25);
or OR3 (N164, N113, N37, N70);
nand NAND4 (N165, N161, N2, N6, N23);
nor NOR4 (N166, N144, N131, N61, N95);
xor XOR2 (N167, N164, N50);
nor NOR4 (N168, N166, N29, N44, N94);
nand NAND4 (N169, N165, N68, N144, N130);
or OR2 (N170, N163, N81);
buf BUF1 (N171, N168);
or OR4 (N172, N167, N104, N21, N159);
buf BUF1 (N173, N172);
not NOT1 (N174, N140);
xor XOR2 (N175, N169, N121);
or OR4 (N176, N173, N162, N153, N27);
and AND4 (N177, N47, N172, N36, N90);
and AND3 (N178, N158, N161, N126);
xor XOR2 (N179, N170, N59);
or OR3 (N180, N175, N72, N139);
xor XOR2 (N181, N177, N124);
buf BUF1 (N182, N179);
and AND4 (N183, N171, N66, N8, N81);
buf BUF1 (N184, N178);
and AND4 (N185, N155, N56, N90, N34);
or OR2 (N186, N183, N150);
buf BUF1 (N187, N156);
xor XOR2 (N188, N160, N70);
and AND3 (N189, N187, N17, N133);
or OR2 (N190, N186, N145);
or OR4 (N191, N185, N40, N69, N149);
or OR3 (N192, N191, N39, N5);
and AND2 (N193, N180, N192);
xor XOR2 (N194, N181, N185);
nor NOR3 (N195, N77, N50, N93);
buf BUF1 (N196, N194);
buf BUF1 (N197, N176);
not NOT1 (N198, N182);
and AND4 (N199, N184, N87, N99, N177);
nor NOR3 (N200, N189, N20, N123);
and AND4 (N201, N174, N13, N166, N117);
xor XOR2 (N202, N201, N139);
or OR2 (N203, N197, N133);
buf BUF1 (N204, N200);
or OR2 (N205, N188, N190);
nor NOR4 (N206, N15, N92, N33, N104);
xor XOR2 (N207, N205, N55);
xor XOR2 (N208, N206, N96);
xor XOR2 (N209, N204, N19);
buf BUF1 (N210, N193);
and AND2 (N211, N209, N147);
and AND3 (N212, N207, N162, N57);
xor XOR2 (N213, N195, N43);
buf BUF1 (N214, N196);
buf BUF1 (N215, N202);
nor NOR4 (N216, N203, N52, N57, N51);
and AND4 (N217, N213, N102, N80, N176);
nor NOR4 (N218, N211, N74, N143, N212);
xor XOR2 (N219, N213, N52);
not NOT1 (N220, N219);
or OR2 (N221, N214, N12);
nand NAND4 (N222, N215, N113, N155, N182);
or OR4 (N223, N217, N145, N12, N164);
and AND2 (N224, N210, N102);
and AND4 (N225, N224, N95, N193, N74);
xor XOR2 (N226, N221, N37);
not NOT1 (N227, N223);
buf BUF1 (N228, N218);
nand NAND4 (N229, N227, N110, N62, N219);
or OR4 (N230, N222, N162, N224, N24);
nand NAND4 (N231, N220, N210, N228, N113);
not NOT1 (N232, N200);
nor NOR3 (N233, N230, N80, N174);
nor NOR3 (N234, N199, N120, N51);
nand NAND3 (N235, N226, N83, N46);
nand NAND2 (N236, N229, N116);
xor XOR2 (N237, N198, N4);
or OR3 (N238, N236, N40, N153);
or OR2 (N239, N235, N215);
and AND2 (N240, N239, N173);
nand NAND3 (N241, N237, N132, N102);
not NOT1 (N242, N238);
not NOT1 (N243, N231);
buf BUF1 (N244, N234);
and AND3 (N245, N244, N157, N164);
or OR3 (N246, N216, N48, N79);
xor XOR2 (N247, N208, N105);
xor XOR2 (N248, N232, N106);
xor XOR2 (N249, N245, N205);
buf BUF1 (N250, N240);
nor NOR3 (N251, N241, N180, N41);
and AND2 (N252, N225, N221);
and AND2 (N253, N246, N78);
or OR4 (N254, N242, N114, N227, N175);
not NOT1 (N255, N251);
or OR4 (N256, N243, N227, N3, N53);
nand NAND4 (N257, N252, N16, N57, N123);
buf BUF1 (N258, N233);
xor XOR2 (N259, N249, N5);
nand NAND2 (N260, N255, N221);
buf BUF1 (N261, N250);
buf BUF1 (N262, N256);
nor NOR4 (N263, N260, N64, N68, N41);
and AND2 (N264, N263, N151);
nor NOR2 (N265, N258, N119);
and AND3 (N266, N259, N87, N146);
nor NOR2 (N267, N264, N129);
or OR3 (N268, N257, N151, N115);
xor XOR2 (N269, N254, N16);
or OR4 (N270, N248, N175, N26, N207);
not NOT1 (N271, N268);
not NOT1 (N272, N261);
or OR2 (N273, N253, N89);
xor XOR2 (N274, N247, N16);
not NOT1 (N275, N265);
nor NOR2 (N276, N271, N232);
nand NAND3 (N277, N267, N269, N9);
buf BUF1 (N278, N254);
or OR4 (N279, N274, N20, N208, N9);
nand NAND2 (N280, N273, N186);
not NOT1 (N281, N266);
and AND4 (N282, N277, N149, N46, N198);
nor NOR3 (N283, N272, N82, N100);
buf BUF1 (N284, N283);
not NOT1 (N285, N278);
nor NOR4 (N286, N270, N134, N164, N51);
nor NOR2 (N287, N285, N198);
and AND3 (N288, N279, N257, N148);
and AND3 (N289, N288, N169, N163);
and AND4 (N290, N262, N156, N168, N103);
nand NAND4 (N291, N286, N45, N241, N134);
nor NOR4 (N292, N282, N93, N99, N81);
nand NAND4 (N293, N290, N180, N130, N147);
not NOT1 (N294, N292);
or OR4 (N295, N293, N221, N284, N25);
buf BUF1 (N296, N88);
buf BUF1 (N297, N275);
buf BUF1 (N298, N297);
xor XOR2 (N299, N287, N109);
nand NAND2 (N300, N298, N154);
buf BUF1 (N301, N300);
buf BUF1 (N302, N301);
not NOT1 (N303, N296);
not NOT1 (N304, N281);
or OR2 (N305, N289, N216);
not NOT1 (N306, N276);
xor XOR2 (N307, N294, N38);
xor XOR2 (N308, N304, N175);
or OR3 (N309, N306, N124, N132);
buf BUF1 (N310, N308);
and AND2 (N311, N303, N64);
xor XOR2 (N312, N307, N187);
nor NOR3 (N313, N310, N173, N202);
nor NOR3 (N314, N302, N303, N201);
or OR4 (N315, N295, N249, N122, N154);
xor XOR2 (N316, N291, N159);
xor XOR2 (N317, N311, N79);
buf BUF1 (N318, N312);
not NOT1 (N319, N315);
or OR4 (N320, N319, N290, N105, N124);
xor XOR2 (N321, N280, N52);
nand NAND3 (N322, N299, N47, N52);
buf BUF1 (N323, N320);
xor XOR2 (N324, N316, N107);
nand NAND4 (N325, N323, N153, N173, N83);
or OR2 (N326, N324, N257);
buf BUF1 (N327, N314);
xor XOR2 (N328, N326, N317);
nor NOR4 (N329, N180, N104, N118, N115);
and AND3 (N330, N318, N168, N187);
nand NAND4 (N331, N327, N33, N107, N95);
nor NOR2 (N332, N313, N207);
not NOT1 (N333, N305);
nand NAND4 (N334, N331, N205, N64, N11);
or OR4 (N335, N325, N195, N129, N315);
not NOT1 (N336, N321);
nand NAND4 (N337, N309, N288, N90, N179);
and AND3 (N338, N322, N81, N226);
or OR4 (N339, N333, N95, N125, N174);
or OR4 (N340, N334, N104, N61, N315);
not NOT1 (N341, N332);
or OR2 (N342, N338, N38);
and AND2 (N343, N339, N19);
not NOT1 (N344, N341);
xor XOR2 (N345, N328, N320);
not NOT1 (N346, N344);
or OR2 (N347, N346, N328);
buf BUF1 (N348, N342);
nand NAND2 (N349, N345, N213);
xor XOR2 (N350, N347, N32);
nand NAND2 (N351, N329, N245);
and AND2 (N352, N337, N340);
buf BUF1 (N353, N208);
and AND4 (N354, N352, N256, N215, N119);
and AND2 (N355, N349, N350);
nand NAND2 (N356, N147, N350);
or OR3 (N357, N336, N164, N229);
or OR3 (N358, N356, N129, N127);
or OR2 (N359, N354, N355);
and AND4 (N360, N218, N41, N31, N328);
not NOT1 (N361, N343);
and AND4 (N362, N361, N11, N152, N332);
and AND2 (N363, N353, N169);
and AND3 (N364, N362, N241, N197);
buf BUF1 (N365, N359);
not NOT1 (N366, N363);
xor XOR2 (N367, N364, N151);
nand NAND3 (N368, N348, N107, N275);
or OR4 (N369, N366, N196, N257, N23);
xor XOR2 (N370, N365, N24);
and AND3 (N371, N358, N318, N178);
xor XOR2 (N372, N367, N53);
buf BUF1 (N373, N351);
nand NAND3 (N374, N360, N135, N233);
xor XOR2 (N375, N330, N345);
and AND2 (N376, N375, N16);
and AND3 (N377, N374, N375, N177);
xor XOR2 (N378, N373, N177);
and AND4 (N379, N368, N170, N84, N348);
or OR3 (N380, N378, N171, N300);
not NOT1 (N381, N335);
nor NOR3 (N382, N370, N252, N73);
not NOT1 (N383, N357);
nor NOR2 (N384, N376, N222);
buf BUF1 (N385, N379);
nor NOR3 (N386, N385, N170, N133);
nand NAND3 (N387, N383, N346, N244);
xor XOR2 (N388, N372, N72);
and AND4 (N389, N384, N341, N176, N239);
nor NOR3 (N390, N377, N23, N77);
not NOT1 (N391, N390);
and AND3 (N392, N381, N223, N30);
not NOT1 (N393, N388);
or OR3 (N394, N386, N365, N273);
and AND2 (N395, N389, N48);
not NOT1 (N396, N369);
and AND4 (N397, N382, N291, N251, N230);
or OR2 (N398, N392, N331);
nand NAND4 (N399, N394, N206, N233, N155);
nor NOR4 (N400, N380, N76, N108, N95);
xor XOR2 (N401, N393, N98);
and AND4 (N402, N391, N39, N24, N118);
or OR2 (N403, N397, N311);
not NOT1 (N404, N403);
nor NOR3 (N405, N371, N85, N201);
nor NOR4 (N406, N398, N256, N85, N35);
nor NOR4 (N407, N404, N335, N309, N279);
nand NAND4 (N408, N402, N78, N365, N39);
and AND4 (N409, N399, N269, N73, N47);
or OR3 (N410, N406, N264, N3);
not NOT1 (N411, N410);
nor NOR2 (N412, N387, N251);
xor XOR2 (N413, N400, N237);
buf BUF1 (N414, N411);
buf BUF1 (N415, N409);
buf BUF1 (N416, N395);
and AND2 (N417, N408, N278);
buf BUF1 (N418, N405);
buf BUF1 (N419, N414);
or OR3 (N420, N401, N286, N162);
buf BUF1 (N421, N420);
not NOT1 (N422, N418);
or OR2 (N423, N421, N240);
nor NOR2 (N424, N415, N59);
nor NOR2 (N425, N407, N177);
xor XOR2 (N426, N412, N361);
and AND3 (N427, N424, N88, N363);
xor XOR2 (N428, N423, N394);
and AND3 (N429, N416, N381, N385);
nor NOR4 (N430, N429, N40, N429, N326);
and AND4 (N431, N428, N53, N107, N47);
buf BUF1 (N432, N396);
nor NOR3 (N433, N430, N294, N10);
not NOT1 (N434, N432);
nand NAND2 (N435, N419, N291);
xor XOR2 (N436, N434, N113);
not NOT1 (N437, N426);
buf BUF1 (N438, N435);
nand NAND4 (N439, N433, N309, N422, N275);
not NOT1 (N440, N318);
nor NOR2 (N441, N436, N131);
xor XOR2 (N442, N431, N292);
and AND4 (N443, N425, N125, N437, N127);
nand NAND3 (N444, N290, N161, N390);
not NOT1 (N445, N442);
nand NAND2 (N446, N413, N87);
nor NOR4 (N447, N440, N11, N250, N94);
or OR2 (N448, N446, N293);
and AND4 (N449, N448, N125, N381, N306);
nor NOR2 (N450, N443, N224);
and AND4 (N451, N427, N141, N192, N351);
nor NOR3 (N452, N441, N7, N29);
nand NAND3 (N453, N444, N162, N41);
or OR3 (N454, N445, N139, N33);
and AND3 (N455, N450, N225, N73);
xor XOR2 (N456, N438, N265);
buf BUF1 (N457, N456);
xor XOR2 (N458, N447, N325);
buf BUF1 (N459, N458);
nor NOR3 (N460, N439, N411, N49);
or OR2 (N461, N457, N375);
nor NOR3 (N462, N417, N458, N264);
xor XOR2 (N463, N449, N173);
nor NOR4 (N464, N462, N226, N417, N237);
or OR3 (N465, N464, N224, N231);
nand NAND2 (N466, N451, N386);
buf BUF1 (N467, N454);
and AND3 (N468, N463, N376, N274);
and AND2 (N469, N466, N334);
xor XOR2 (N470, N452, N191);
and AND3 (N471, N461, N47, N245);
xor XOR2 (N472, N469, N138);
xor XOR2 (N473, N468, N440);
xor XOR2 (N474, N471, N169);
nand NAND2 (N475, N465, N15);
buf BUF1 (N476, N474);
and AND3 (N477, N470, N190, N35);
xor XOR2 (N478, N475, N257);
xor XOR2 (N479, N477, N387);
not NOT1 (N480, N478);
xor XOR2 (N481, N476, N301);
not NOT1 (N482, N479);
nor NOR3 (N483, N481, N90, N385);
xor XOR2 (N484, N480, N69);
and AND4 (N485, N467, N146, N135, N241);
or OR3 (N486, N483, N250, N269);
buf BUF1 (N487, N486);
buf BUF1 (N488, N472);
not NOT1 (N489, N460);
not NOT1 (N490, N487);
nand NAND2 (N491, N455, N218);
xor XOR2 (N492, N490, N463);
and AND2 (N493, N484, N102);
nor NOR3 (N494, N482, N248, N419);
or OR2 (N495, N473, N275);
nor NOR2 (N496, N492, N420);
xor XOR2 (N497, N496, N333);
not NOT1 (N498, N491);
xor XOR2 (N499, N494, N150);
not NOT1 (N500, N497);
nor NOR2 (N501, N500, N62);
nor NOR3 (N502, N495, N368, N123);
or OR2 (N503, N485, N171);
and AND4 (N504, N488, N125, N494, N161);
buf BUF1 (N505, N502);
not NOT1 (N506, N505);
or OR2 (N507, N504, N103);
nand NAND2 (N508, N506, N302);
not NOT1 (N509, N498);
or OR3 (N510, N493, N191, N452);
not NOT1 (N511, N501);
buf BUF1 (N512, N511);
buf BUF1 (N513, N507);
not NOT1 (N514, N509);
nand NAND4 (N515, N489, N353, N178, N473);
and AND2 (N516, N514, N66);
and AND4 (N517, N510, N420, N240, N13);
xor XOR2 (N518, N516, N343);
xor XOR2 (N519, N518, N422);
or OR2 (N520, N515, N342);
nor NOR3 (N521, N503, N141, N25);
nor NOR2 (N522, N499, N199);
and AND4 (N523, N459, N455, N77, N520);
nand NAND3 (N524, N129, N1, N205);
and AND2 (N525, N522, N148);
buf BUF1 (N526, N525);
xor XOR2 (N527, N524, N382);
nand NAND4 (N528, N521, N128, N194, N176);
or OR2 (N529, N508, N357);
or OR2 (N530, N513, N283);
nor NOR3 (N531, N523, N208, N268);
not NOT1 (N532, N529);
or OR3 (N533, N532, N194, N494);
nand NAND4 (N534, N528, N287, N82, N214);
nor NOR4 (N535, N527, N36, N471, N139);
and AND2 (N536, N530, N157);
nand NAND3 (N537, N534, N319, N502);
xor XOR2 (N538, N531, N370);
or OR3 (N539, N536, N58, N487);
xor XOR2 (N540, N537, N216);
buf BUF1 (N541, N512);
xor XOR2 (N542, N517, N189);
and AND4 (N543, N533, N378, N522, N384);
nor NOR4 (N544, N542, N461, N147, N218);
xor XOR2 (N545, N540, N234);
and AND2 (N546, N453, N129);
nor NOR2 (N547, N519, N90);
not NOT1 (N548, N535);
and AND4 (N549, N547, N300, N244, N380);
or OR4 (N550, N548, N529, N495, N57);
not NOT1 (N551, N539);
nor NOR4 (N552, N526, N198, N456, N535);
nor NOR3 (N553, N550, N379, N282);
or OR4 (N554, N538, N203, N475, N300);
nor NOR4 (N555, N545, N82, N176, N186);
nand NAND4 (N556, N549, N375, N551, N183);
or OR2 (N557, N552, N411);
or OR2 (N558, N191, N414);
not NOT1 (N559, N544);
nand NAND2 (N560, N553, N78);
xor XOR2 (N561, N556, N500);
nand NAND3 (N562, N543, N78, N243);
xor XOR2 (N563, N558, N391);
nand NAND2 (N564, N555, N331);
nand NAND3 (N565, N554, N237, N384);
xor XOR2 (N566, N557, N139);
and AND4 (N567, N565, N383, N390, N374);
xor XOR2 (N568, N560, N369);
buf BUF1 (N569, N567);
nand NAND3 (N570, N568, N62, N253);
not NOT1 (N571, N570);
xor XOR2 (N572, N571, N5);
nand NAND3 (N573, N541, N351, N68);
not NOT1 (N574, N573);
or OR4 (N575, N566, N317, N474, N144);
xor XOR2 (N576, N546, N298);
or OR2 (N577, N574, N534);
nand NAND3 (N578, N576, N92, N535);
or OR3 (N579, N564, N260, N413);
not NOT1 (N580, N563);
not NOT1 (N581, N575);
or OR3 (N582, N561, N390, N280);
and AND2 (N583, N559, N173);
buf BUF1 (N584, N581);
not NOT1 (N585, N583);
or OR2 (N586, N579, N469);
xor XOR2 (N587, N577, N42);
nand NAND2 (N588, N569, N475);
not NOT1 (N589, N586);
and AND2 (N590, N585, N157);
not NOT1 (N591, N580);
nor NOR2 (N592, N582, N463);
xor XOR2 (N593, N578, N5);
buf BUF1 (N594, N572);
or OR4 (N595, N592, N234, N160, N520);
buf BUF1 (N596, N588);
or OR3 (N597, N591, N173, N587);
not NOT1 (N598, N234);
xor XOR2 (N599, N597, N259);
xor XOR2 (N600, N596, N466);
nor NOR2 (N601, N595, N466);
not NOT1 (N602, N562);
and AND3 (N603, N601, N592, N187);
not NOT1 (N604, N590);
nand NAND3 (N605, N598, N57, N219);
buf BUF1 (N606, N605);
nor NOR4 (N607, N602, N404, N460, N465);
not NOT1 (N608, N600);
not NOT1 (N609, N594);
xor XOR2 (N610, N584, N515);
buf BUF1 (N611, N608);
xor XOR2 (N612, N593, N40);
nand NAND4 (N613, N589, N438, N408, N596);
nand NAND3 (N614, N603, N140, N196);
not NOT1 (N615, N610);
nor NOR2 (N616, N612, N606);
xor XOR2 (N617, N180, N368);
buf BUF1 (N618, N599);
nand NAND2 (N619, N604, N206);
buf BUF1 (N620, N618);
nand NAND3 (N621, N616, N564, N595);
buf BUF1 (N622, N620);
xor XOR2 (N623, N615, N130);
nand NAND2 (N624, N609, N520);
and AND2 (N625, N607, N306);
nor NOR4 (N626, N624, N119, N466, N289);
and AND4 (N627, N622, N304, N546, N254);
and AND2 (N628, N613, N577);
and AND2 (N629, N626, N567);
buf BUF1 (N630, N621);
nand NAND4 (N631, N628, N366, N174, N89);
nand NAND4 (N632, N619, N94, N327, N239);
xor XOR2 (N633, N632, N365);
nand NAND3 (N634, N631, N23, N537);
nor NOR4 (N635, N629, N527, N52, N215);
or OR4 (N636, N635, N105, N140, N112);
and AND4 (N637, N623, N625, N585, N486);
or OR2 (N638, N605, N349);
or OR3 (N639, N637, N544, N479);
nand NAND2 (N640, N630, N611);
nor NOR4 (N641, N41, N258, N281, N296);
nand NAND2 (N642, N614, N639);
nor NOR3 (N643, N407, N207, N224);
or OR3 (N644, N638, N615, N26);
and AND4 (N645, N617, N625, N613, N326);
or OR3 (N646, N636, N596, N132);
and AND3 (N647, N645, N608, N2);
buf BUF1 (N648, N643);
or OR3 (N649, N646, N636, N286);
nor NOR4 (N650, N642, N544, N19, N541);
buf BUF1 (N651, N641);
buf BUF1 (N652, N634);
not NOT1 (N653, N650);
not NOT1 (N654, N648);
buf BUF1 (N655, N627);
nand NAND3 (N656, N649, N604, N186);
buf BUF1 (N657, N640);
buf BUF1 (N658, N655);
and AND3 (N659, N647, N657, N409);
nand NAND4 (N660, N104, N117, N577, N465);
and AND2 (N661, N652, N105);
buf BUF1 (N662, N658);
buf BUF1 (N663, N656);
nor NOR3 (N664, N633, N241, N226);
or OR2 (N665, N664, N40);
buf BUF1 (N666, N653);
not NOT1 (N667, N660);
or OR2 (N668, N666, N492);
or OR3 (N669, N662, N534, N413);
nor NOR2 (N670, N663, N131);
xor XOR2 (N671, N659, N357);
xor XOR2 (N672, N651, N596);
xor XOR2 (N673, N665, N670);
xor XOR2 (N674, N578, N144);
nor NOR3 (N675, N654, N301, N276);
nand NAND4 (N676, N672, N590, N177, N153);
or OR4 (N677, N661, N248, N101, N608);
and AND4 (N678, N675, N610, N268, N454);
xor XOR2 (N679, N667, N133);
and AND4 (N680, N676, N529, N566, N495);
xor XOR2 (N681, N668, N44);
or OR3 (N682, N679, N437, N459);
xor XOR2 (N683, N677, N391);
and AND4 (N684, N683, N661, N599, N442);
and AND3 (N685, N673, N135, N164);
buf BUF1 (N686, N685);
nand NAND3 (N687, N681, N102, N139);
or OR2 (N688, N678, N661);
or OR2 (N689, N644, N553);
and AND2 (N690, N671, N404);
xor XOR2 (N691, N669, N66);
not NOT1 (N692, N686);
nand NAND3 (N693, N674, N200, N543);
nand NAND4 (N694, N680, N420, N477, N666);
nand NAND4 (N695, N687, N685, N83, N396);
nand NAND2 (N696, N694, N382);
or OR2 (N697, N688, N156);
nand NAND4 (N698, N691, N501, N87, N405);
nand NAND2 (N699, N698, N359);
xor XOR2 (N700, N697, N551);
nor NOR4 (N701, N693, N369, N410, N170);
and AND2 (N702, N690, N186);
nor NOR2 (N703, N700, N669);
nor NOR2 (N704, N702, N333);
buf BUF1 (N705, N701);
nor NOR2 (N706, N704, N654);
and AND2 (N707, N696, N323);
xor XOR2 (N708, N692, N650);
or OR4 (N709, N705, N288, N565, N409);
buf BUF1 (N710, N707);
buf BUF1 (N711, N699);
or OR4 (N712, N708, N614, N12, N653);
nand NAND4 (N713, N689, N469, N156, N125);
buf BUF1 (N714, N703);
not NOT1 (N715, N695);
not NOT1 (N716, N709);
buf BUF1 (N717, N714);
and AND2 (N718, N710, N600);
and AND3 (N719, N713, N547, N146);
xor XOR2 (N720, N719, N90);
or OR3 (N721, N711, N514, N415);
or OR3 (N722, N721, N433, N516);
xor XOR2 (N723, N720, N90);
nand NAND4 (N724, N715, N105, N652, N186);
or OR4 (N725, N723, N614, N279, N189);
xor XOR2 (N726, N712, N629);
nor NOR3 (N727, N718, N224, N525);
not NOT1 (N728, N706);
xor XOR2 (N729, N725, N391);
buf BUF1 (N730, N682);
or OR2 (N731, N722, N345);
or OR4 (N732, N730, N623, N727, N91);
xor XOR2 (N733, N626, N366);
xor XOR2 (N734, N731, N247);
not NOT1 (N735, N726);
or OR4 (N736, N684, N591, N334, N36);
not NOT1 (N737, N733);
nor NOR3 (N738, N732, N633, N612);
not NOT1 (N739, N717);
nand NAND4 (N740, N737, N186, N353, N159);
buf BUF1 (N741, N724);
and AND2 (N742, N739, N124);
not NOT1 (N743, N728);
and AND2 (N744, N716, N679);
nor NOR3 (N745, N744, N395, N348);
and AND2 (N746, N734, N600);
xor XOR2 (N747, N736, N550);
nand NAND3 (N748, N746, N497, N555);
and AND4 (N749, N743, N366, N380, N94);
buf BUF1 (N750, N729);
and AND3 (N751, N750, N97, N320);
nand NAND4 (N752, N749, N13, N446, N459);
and AND2 (N753, N752, N592);
xor XOR2 (N754, N738, N655);
nor NOR4 (N755, N742, N451, N452, N537);
buf BUF1 (N756, N755);
nand NAND3 (N757, N753, N421, N641);
nand NAND2 (N758, N757, N450);
not NOT1 (N759, N748);
and AND3 (N760, N754, N114, N489);
or OR3 (N761, N735, N184, N280);
buf BUF1 (N762, N747);
nor NOR3 (N763, N756, N747, N411);
xor XOR2 (N764, N762, N189);
nor NOR3 (N765, N764, N754, N534);
or OR2 (N766, N765, N203);
not NOT1 (N767, N759);
xor XOR2 (N768, N741, N277);
xor XOR2 (N769, N768, N332);
buf BUF1 (N770, N766);
nand NAND2 (N771, N740, N273);
not NOT1 (N772, N771);
xor XOR2 (N773, N769, N452);
xor XOR2 (N774, N760, N50);
xor XOR2 (N775, N745, N359);
nor NOR2 (N776, N770, N125);
or OR3 (N777, N775, N500, N126);
nor NOR3 (N778, N751, N758, N573);
buf BUF1 (N779, N259);
nand NAND4 (N780, N779, N657, N15, N422);
or OR3 (N781, N774, N498, N292);
xor XOR2 (N782, N767, N353);
buf BUF1 (N783, N772);
buf BUF1 (N784, N780);
buf BUF1 (N785, N778);
buf BUF1 (N786, N783);
and AND3 (N787, N782, N153, N42);
nor NOR3 (N788, N777, N611, N220);
xor XOR2 (N789, N763, N341);
and AND4 (N790, N785, N726, N378, N511);
xor XOR2 (N791, N776, N178);
or OR3 (N792, N791, N610, N353);
or OR3 (N793, N789, N187, N294);
not NOT1 (N794, N781);
or OR2 (N795, N786, N241);
or OR2 (N796, N784, N664);
and AND3 (N797, N795, N35, N221);
buf BUF1 (N798, N788);
not NOT1 (N799, N798);
xor XOR2 (N800, N794, N325);
nand NAND2 (N801, N797, N552);
xor XOR2 (N802, N800, N184);
or OR4 (N803, N792, N242, N161, N349);
not NOT1 (N804, N802);
nand NAND2 (N805, N796, N629);
or OR4 (N806, N803, N198, N279, N273);
xor XOR2 (N807, N806, N431);
buf BUF1 (N808, N773);
or OR2 (N809, N807, N412);
xor XOR2 (N810, N761, N431);
not NOT1 (N811, N808);
and AND2 (N812, N805, N341);
or OR2 (N813, N790, N56);
buf BUF1 (N814, N812);
xor XOR2 (N815, N811, N301);
xor XOR2 (N816, N813, N253);
and AND4 (N817, N814, N399, N657, N90);
nand NAND3 (N818, N817, N804, N381);
nor NOR3 (N819, N553, N300, N580);
buf BUF1 (N820, N816);
or OR4 (N821, N799, N119, N513, N646);
nand NAND4 (N822, N810, N166, N701, N788);
nand NAND2 (N823, N787, N408);
not NOT1 (N824, N815);
buf BUF1 (N825, N824);
nand NAND4 (N826, N823, N284, N277, N330);
buf BUF1 (N827, N809);
xor XOR2 (N828, N826, N193);
xor XOR2 (N829, N819, N30);
not NOT1 (N830, N825);
nand NAND4 (N831, N827, N377, N241, N448);
buf BUF1 (N832, N793);
buf BUF1 (N833, N821);
buf BUF1 (N834, N822);
buf BUF1 (N835, N801);
nor NOR4 (N836, N835, N467, N245, N538);
nand NAND4 (N837, N828, N573, N827, N619);
nor NOR2 (N838, N830, N704);
not NOT1 (N839, N832);
buf BUF1 (N840, N831);
xor XOR2 (N841, N834, N747);
and AND4 (N842, N837, N301, N599, N178);
or OR2 (N843, N839, N12);
xor XOR2 (N844, N838, N661);
buf BUF1 (N845, N841);
buf BUF1 (N846, N820);
or OR4 (N847, N836, N278, N754, N330);
or OR2 (N848, N818, N672);
nor NOR4 (N849, N843, N166, N371, N54);
and AND4 (N850, N840, N428, N806, N48);
and AND3 (N851, N848, N292, N660);
or OR3 (N852, N829, N395, N833);
and AND4 (N853, N249, N463, N65, N206);
and AND4 (N854, N852, N633, N819, N723);
nand NAND3 (N855, N851, N802, N677);
nand NAND2 (N856, N850, N536);
and AND4 (N857, N846, N794, N809, N806);
buf BUF1 (N858, N853);
nor NOR4 (N859, N856, N423, N201, N511);
buf BUF1 (N860, N858);
xor XOR2 (N861, N849, N225);
nor NOR2 (N862, N845, N80);
xor XOR2 (N863, N854, N861);
nor NOR4 (N864, N747, N618, N318, N535);
xor XOR2 (N865, N844, N572);
xor XOR2 (N866, N863, N425);
or OR2 (N867, N847, N475);
and AND4 (N868, N842, N338, N554, N287);
buf BUF1 (N869, N862);
nor NOR2 (N870, N869, N171);
and AND2 (N871, N859, N88);
not NOT1 (N872, N871);
xor XOR2 (N873, N866, N374);
buf BUF1 (N874, N873);
buf BUF1 (N875, N857);
xor XOR2 (N876, N855, N296);
xor XOR2 (N877, N864, N407);
and AND4 (N878, N875, N650, N135, N831);
and AND2 (N879, N860, N698);
buf BUF1 (N880, N865);
nor NOR4 (N881, N870, N435, N626, N391);
or OR2 (N882, N876, N129);
and AND4 (N883, N872, N309, N827, N233);
or OR4 (N884, N867, N831, N313, N718);
nand NAND3 (N885, N884, N701, N108);
and AND2 (N886, N881, N186);
or OR4 (N887, N874, N364, N699, N814);
not NOT1 (N888, N882);
nand NAND3 (N889, N887, N324, N860);
nor NOR2 (N890, N885, N177);
not NOT1 (N891, N878);
not NOT1 (N892, N889);
xor XOR2 (N893, N879, N262);
xor XOR2 (N894, N888, N67);
nor NOR2 (N895, N880, N238);
buf BUF1 (N896, N892);
and AND3 (N897, N883, N33, N335);
not NOT1 (N898, N894);
not NOT1 (N899, N893);
and AND2 (N900, N890, N306);
not NOT1 (N901, N899);
and AND3 (N902, N891, N661, N34);
xor XOR2 (N903, N877, N244);
and AND3 (N904, N897, N756, N857);
nor NOR3 (N905, N895, N378, N93);
not NOT1 (N906, N898);
buf BUF1 (N907, N903);
nor NOR4 (N908, N902, N429, N604, N390);
xor XOR2 (N909, N906, N784);
buf BUF1 (N910, N907);
nand NAND2 (N911, N908, N6);
and AND3 (N912, N900, N463, N204);
or OR3 (N913, N909, N906, N537);
nand NAND3 (N914, N904, N670, N529);
nand NAND4 (N915, N868, N735, N271, N325);
and AND3 (N916, N914, N271, N411);
and AND3 (N917, N913, N16, N90);
and AND2 (N918, N901, N808);
xor XOR2 (N919, N896, N393);
buf BUF1 (N920, N886);
and AND2 (N921, N917, N824);
buf BUF1 (N922, N918);
nand NAND4 (N923, N922, N341, N645, N174);
not NOT1 (N924, N912);
or OR4 (N925, N905, N350, N512, N526);
nand NAND3 (N926, N911, N184, N130);
not NOT1 (N927, N910);
not NOT1 (N928, N927);
nand NAND2 (N929, N919, N365);
xor XOR2 (N930, N921, N500);
buf BUF1 (N931, N926);
not NOT1 (N932, N931);
and AND3 (N933, N928, N241, N433);
nand NAND3 (N934, N929, N828, N344);
xor XOR2 (N935, N933, N915);
nor NOR4 (N936, N772, N287, N658, N527);
and AND4 (N937, N932, N51, N208, N908);
nor NOR2 (N938, N924, N565);
buf BUF1 (N939, N935);
xor XOR2 (N940, N920, N405);
not NOT1 (N941, N923);
nor NOR2 (N942, N937, N557);
nor NOR3 (N943, N934, N345, N256);
buf BUF1 (N944, N930);
xor XOR2 (N945, N936, N586);
buf BUF1 (N946, N939);
xor XOR2 (N947, N941, N99);
buf BUF1 (N948, N945);
and AND4 (N949, N948, N915, N806, N219);
xor XOR2 (N950, N916, N665);
xor XOR2 (N951, N950, N64);
buf BUF1 (N952, N946);
nor NOR4 (N953, N938, N510, N806, N124);
nor NOR4 (N954, N949, N698, N744, N822);
or OR3 (N955, N951, N352, N87);
or OR4 (N956, N943, N351, N478, N398);
nand NAND2 (N957, N953, N323);
or OR3 (N958, N940, N390, N805);
buf BUF1 (N959, N955);
nand NAND4 (N960, N958, N798, N699, N901);
not NOT1 (N961, N954);
and AND2 (N962, N959, N613);
and AND2 (N963, N957, N687);
buf BUF1 (N964, N942);
nand NAND3 (N965, N964, N736, N307);
nand NAND3 (N966, N952, N651, N312);
buf BUF1 (N967, N963);
nand NAND3 (N968, N961, N825, N458);
nand NAND3 (N969, N947, N637, N365);
or OR4 (N970, N965, N321, N846, N708);
nand NAND3 (N971, N944, N732, N503);
or OR4 (N972, N969, N779, N8, N693);
nor NOR2 (N973, N970, N237);
nor NOR3 (N974, N967, N971, N357);
and AND3 (N975, N893, N228, N701);
or OR3 (N976, N960, N47, N787);
buf BUF1 (N977, N973);
nor NOR4 (N978, N977, N470, N307, N855);
nor NOR3 (N979, N974, N90, N914);
or OR4 (N980, N968, N293, N967, N371);
or OR4 (N981, N978, N14, N399, N639);
or OR3 (N982, N956, N789, N719);
not NOT1 (N983, N982);
and AND4 (N984, N972, N180, N600, N71);
nor NOR2 (N985, N983, N31);
or OR3 (N986, N962, N407, N779);
or OR3 (N987, N985, N925, N702);
and AND4 (N988, N937, N326, N262, N688);
nor NOR2 (N989, N980, N440);
not NOT1 (N990, N986);
and AND2 (N991, N966, N116);
nand NAND4 (N992, N976, N297, N311, N446);
nand NAND3 (N993, N988, N49, N737);
buf BUF1 (N994, N979);
buf BUF1 (N995, N987);
xor XOR2 (N996, N990, N710);
xor XOR2 (N997, N994, N951);
nand NAND2 (N998, N984, N873);
nor NOR4 (N999, N981, N617, N458, N875);
buf BUF1 (N1000, N996);
and AND3 (N1001, N989, N240, N857);
or OR3 (N1002, N975, N337, N65);
nor NOR4 (N1003, N998, N499, N26, N575);
nand NAND2 (N1004, N1001, N422);
or OR3 (N1005, N992, N729, N29);
xor XOR2 (N1006, N991, N418);
buf BUF1 (N1007, N999);
nand NAND4 (N1008, N993, N132, N242, N178);
not NOT1 (N1009, N995);
and AND3 (N1010, N1000, N753, N999);
xor XOR2 (N1011, N1008, N389);
nand NAND3 (N1012, N1011, N915, N237);
or OR4 (N1013, N997, N442, N733, N78);
or OR2 (N1014, N1009, N907);
nand NAND3 (N1015, N1012, N717, N234);
not NOT1 (N1016, N1013);
nor NOR2 (N1017, N1004, N101);
xor XOR2 (N1018, N1015, N301);
nand NAND4 (N1019, N1016, N117, N359, N271);
buf BUF1 (N1020, N1010);
nand NAND2 (N1021, N1019, N575);
not NOT1 (N1022, N1006);
buf BUF1 (N1023, N1022);
nor NOR3 (N1024, N1014, N471, N310);
nand NAND4 (N1025, N1024, N357, N598, N507);
nand NAND3 (N1026, N1021, N202, N802);
buf BUF1 (N1027, N1005);
not NOT1 (N1028, N1018);
xor XOR2 (N1029, N1003, N920);
or OR4 (N1030, N1027, N412, N486, N615);
xor XOR2 (N1031, N1023, N570);
or OR4 (N1032, N1031, N41, N830, N221);
or OR3 (N1033, N1030, N735, N283);
nand NAND4 (N1034, N1033, N252, N441, N682);
and AND2 (N1035, N1032, N643);
not NOT1 (N1036, N1007);
xor XOR2 (N1037, N1020, N302);
or OR2 (N1038, N1037, N408);
or OR4 (N1039, N1038, N910, N829, N366);
xor XOR2 (N1040, N1039, N795);
and AND3 (N1041, N1026, N119, N890);
buf BUF1 (N1042, N1041);
and AND3 (N1043, N1035, N1026, N869);
xor XOR2 (N1044, N1043, N357);
xor XOR2 (N1045, N1017, N115);
not NOT1 (N1046, N1029);
nand NAND4 (N1047, N1034, N738, N526, N348);
or OR3 (N1048, N1040, N766, N153);
nand NAND4 (N1049, N1045, N263, N725, N818);
nand NAND2 (N1050, N1044, N284);
buf BUF1 (N1051, N1002);
buf BUF1 (N1052, N1051);
nor NOR2 (N1053, N1042, N373);
or OR3 (N1054, N1052, N353, N563);
or OR3 (N1055, N1025, N543, N134);
nand NAND2 (N1056, N1036, N329);
and AND2 (N1057, N1049, N962);
not NOT1 (N1058, N1046);
xor XOR2 (N1059, N1048, N724);
not NOT1 (N1060, N1028);
xor XOR2 (N1061, N1059, N312);
nand NAND3 (N1062, N1056, N247, N869);
or OR3 (N1063, N1047, N554, N468);
buf BUF1 (N1064, N1060);
nand NAND4 (N1065, N1055, N701, N54, N35);
buf BUF1 (N1066, N1063);
xor XOR2 (N1067, N1064, N381);
nand NAND4 (N1068, N1067, N379, N287, N959);
xor XOR2 (N1069, N1054, N642);
nor NOR4 (N1070, N1058, N589, N707, N720);
nor NOR4 (N1071, N1069, N785, N926, N710);
nor NOR3 (N1072, N1070, N279, N16);
not NOT1 (N1073, N1057);
nor NOR4 (N1074, N1065, N342, N126, N30);
nand NAND3 (N1075, N1072, N307, N450);
nand NAND2 (N1076, N1062, N725);
or OR4 (N1077, N1068, N903, N419, N678);
nand NAND3 (N1078, N1050, N620, N406);
buf BUF1 (N1079, N1053);
and AND2 (N1080, N1074, N320);
nand NAND2 (N1081, N1077, N691);
xor XOR2 (N1082, N1071, N573);
buf BUF1 (N1083, N1080);
buf BUF1 (N1084, N1078);
buf BUF1 (N1085, N1076);
buf BUF1 (N1086, N1075);
and AND2 (N1087, N1085, N397);
not NOT1 (N1088, N1084);
not NOT1 (N1089, N1066);
nand NAND2 (N1090, N1073, N637);
nor NOR3 (N1091, N1081, N967, N897);
nand NAND4 (N1092, N1088, N332, N792, N144);
nor NOR4 (N1093, N1089, N1055, N251, N228);
or OR2 (N1094, N1086, N854);
not NOT1 (N1095, N1082);
xor XOR2 (N1096, N1095, N437);
nand NAND4 (N1097, N1093, N77, N841, N531);
xor XOR2 (N1098, N1092, N128);
not NOT1 (N1099, N1096);
nor NOR3 (N1100, N1099, N382, N520);
xor XOR2 (N1101, N1083, N264);
or OR4 (N1102, N1087, N1031, N28, N692);
buf BUF1 (N1103, N1094);
and AND3 (N1104, N1091, N496, N59);
and AND3 (N1105, N1104, N492, N189);
buf BUF1 (N1106, N1102);
and AND2 (N1107, N1061, N515);
nor NOR3 (N1108, N1101, N761, N934);
xor XOR2 (N1109, N1097, N2);
or OR3 (N1110, N1103, N96, N57);
and AND3 (N1111, N1098, N721, N623);
or OR3 (N1112, N1079, N412, N255);
xor XOR2 (N1113, N1108, N469);
buf BUF1 (N1114, N1109);
or OR4 (N1115, N1107, N985, N993, N1053);
nor NOR4 (N1116, N1112, N1035, N1062, N883);
not NOT1 (N1117, N1111);
not NOT1 (N1118, N1105);
buf BUF1 (N1119, N1114);
or OR2 (N1120, N1116, N772);
and AND4 (N1121, N1106, N264, N260, N333);
nor NOR3 (N1122, N1118, N675, N356);
and AND3 (N1123, N1122, N12, N393);
nand NAND2 (N1124, N1110, N582);
xor XOR2 (N1125, N1090, N720);
xor XOR2 (N1126, N1121, N879);
not NOT1 (N1127, N1115);
nor NOR2 (N1128, N1123, N1102);
or OR2 (N1129, N1125, N248);
buf BUF1 (N1130, N1124);
nand NAND3 (N1131, N1128, N122, N615);
and AND3 (N1132, N1131, N44, N908);
not NOT1 (N1133, N1119);
and AND2 (N1134, N1120, N719);
nor NOR3 (N1135, N1134, N149, N65);
buf BUF1 (N1136, N1135);
nand NAND3 (N1137, N1117, N938, N999);
nor NOR2 (N1138, N1126, N863);
buf BUF1 (N1139, N1137);
and AND2 (N1140, N1132, N608);
nor NOR3 (N1141, N1133, N228, N651);
xor XOR2 (N1142, N1138, N220);
buf BUF1 (N1143, N1136);
or OR3 (N1144, N1141, N737, N698);
buf BUF1 (N1145, N1129);
xor XOR2 (N1146, N1139, N54);
nand NAND2 (N1147, N1130, N778);
not NOT1 (N1148, N1143);
or OR3 (N1149, N1145, N120, N715);
xor XOR2 (N1150, N1127, N81);
and AND4 (N1151, N1147, N545, N970, N652);
not NOT1 (N1152, N1148);
nor NOR3 (N1153, N1140, N674, N63);
or OR4 (N1154, N1142, N970, N41, N539);
buf BUF1 (N1155, N1113);
or OR3 (N1156, N1144, N387, N520);
buf BUF1 (N1157, N1155);
nand NAND3 (N1158, N1154, N76, N993);
nor NOR2 (N1159, N1156, N530);
and AND4 (N1160, N1149, N1136, N718, N404);
nand NAND2 (N1161, N1153, N652);
or OR2 (N1162, N1150, N730);
nor NOR2 (N1163, N1157, N883);
not NOT1 (N1164, N1160);
and AND2 (N1165, N1100, N71);
nand NAND3 (N1166, N1164, N1034, N1117);
or OR4 (N1167, N1159, N752, N925, N1072);
buf BUF1 (N1168, N1158);
xor XOR2 (N1169, N1167, N856);
or OR4 (N1170, N1165, N926, N180, N396);
or OR4 (N1171, N1170, N639, N920, N713);
nand NAND2 (N1172, N1152, N561);
nor NOR4 (N1173, N1162, N1135, N19, N804);
not NOT1 (N1174, N1151);
nand NAND2 (N1175, N1161, N1098);
nor NOR2 (N1176, N1169, N241);
nand NAND4 (N1177, N1163, N323, N431, N144);
or OR2 (N1178, N1175, N847);
not NOT1 (N1179, N1176);
xor XOR2 (N1180, N1168, N1001);
buf BUF1 (N1181, N1174);
nand NAND3 (N1182, N1146, N437, N965);
xor XOR2 (N1183, N1172, N1034);
buf BUF1 (N1184, N1166);
not NOT1 (N1185, N1183);
and AND2 (N1186, N1173, N386);
or OR4 (N1187, N1181, N147, N436, N1152);
or OR2 (N1188, N1178, N18);
and AND4 (N1189, N1188, N449, N598, N744);
not NOT1 (N1190, N1186);
and AND3 (N1191, N1179, N192, N366);
nand NAND2 (N1192, N1177, N1135);
and AND3 (N1193, N1185, N196, N529);
xor XOR2 (N1194, N1180, N619);
and AND4 (N1195, N1194, N876, N322, N977);
not NOT1 (N1196, N1191);
and AND2 (N1197, N1171, N70);
xor XOR2 (N1198, N1190, N1122);
not NOT1 (N1199, N1198);
nand NAND2 (N1200, N1195, N834);
not NOT1 (N1201, N1197);
buf BUF1 (N1202, N1182);
and AND4 (N1203, N1184, N12, N602, N692);
xor XOR2 (N1204, N1196, N1023);
and AND3 (N1205, N1199, N699, N724);
nor NOR2 (N1206, N1204, N585);
xor XOR2 (N1207, N1193, N1137);
not NOT1 (N1208, N1202);
and AND2 (N1209, N1205, N295);
xor XOR2 (N1210, N1207, N914);
or OR2 (N1211, N1206, N668);
xor XOR2 (N1212, N1208, N1197);
or OR2 (N1213, N1203, N164);
not NOT1 (N1214, N1189);
and AND4 (N1215, N1192, N1076, N399, N452);
and AND2 (N1216, N1214, N1111);
or OR2 (N1217, N1211, N977);
buf BUF1 (N1218, N1213);
nand NAND3 (N1219, N1210, N592, N1060);
and AND2 (N1220, N1219, N194);
nor NOR3 (N1221, N1212, N1118, N339);
not NOT1 (N1222, N1221);
nand NAND3 (N1223, N1222, N862, N394);
not NOT1 (N1224, N1223);
buf BUF1 (N1225, N1216);
or OR3 (N1226, N1217, N848, N1015);
buf BUF1 (N1227, N1220);
buf BUF1 (N1228, N1225);
or OR4 (N1229, N1209, N986, N248, N1120);
and AND2 (N1230, N1215, N223);
nor NOR4 (N1231, N1201, N1015, N652, N858);
nor NOR3 (N1232, N1224, N984, N1100);
not NOT1 (N1233, N1229);
xor XOR2 (N1234, N1228, N158);
buf BUF1 (N1235, N1234);
nor NOR3 (N1236, N1231, N1031, N409);
xor XOR2 (N1237, N1235, N616);
and AND4 (N1238, N1200, N990, N1007, N455);
nor NOR2 (N1239, N1236, N805);
nor NOR2 (N1240, N1230, N1016);
and AND3 (N1241, N1232, N882, N485);
not NOT1 (N1242, N1227);
and AND2 (N1243, N1238, N371);
nand NAND3 (N1244, N1241, N709, N538);
xor XOR2 (N1245, N1242, N346);
or OR4 (N1246, N1245, N964, N837, N296);
not NOT1 (N1247, N1244);
xor XOR2 (N1248, N1233, N1209);
buf BUF1 (N1249, N1218);
and AND2 (N1250, N1249, N905);
nor NOR4 (N1251, N1239, N1132, N711, N56);
or OR2 (N1252, N1247, N273);
nor NOR3 (N1253, N1248, N486, N243);
not NOT1 (N1254, N1253);
not NOT1 (N1255, N1187);
not NOT1 (N1256, N1240);
nor NOR2 (N1257, N1237, N736);
buf BUF1 (N1258, N1257);
nor NOR3 (N1259, N1250, N853, N889);
not NOT1 (N1260, N1258);
nand NAND2 (N1261, N1255, N938);
buf BUF1 (N1262, N1243);
buf BUF1 (N1263, N1256);
nor NOR4 (N1264, N1263, N857, N977, N828);
xor XOR2 (N1265, N1226, N1257);
nand NAND2 (N1266, N1260, N193);
not NOT1 (N1267, N1265);
and AND4 (N1268, N1254, N1093, N1003, N918);
buf BUF1 (N1269, N1267);
buf BUF1 (N1270, N1266);
or OR2 (N1271, N1259, N1186);
not NOT1 (N1272, N1268);
nand NAND4 (N1273, N1272, N888, N444, N291);
not NOT1 (N1274, N1270);
or OR4 (N1275, N1274, N1047, N1113, N774);
buf BUF1 (N1276, N1251);
nand NAND2 (N1277, N1275, N312);
nand NAND2 (N1278, N1262, N1056);
buf BUF1 (N1279, N1276);
nor NOR2 (N1280, N1269, N367);
or OR3 (N1281, N1252, N918, N770);
or OR2 (N1282, N1264, N1233);
buf BUF1 (N1283, N1281);
not NOT1 (N1284, N1278);
xor XOR2 (N1285, N1277, N1);
nand NAND3 (N1286, N1282, N972, N921);
nor NOR2 (N1287, N1284, N829);
and AND2 (N1288, N1287, N228);
and AND4 (N1289, N1286, N662, N305, N1136);
not NOT1 (N1290, N1283);
xor XOR2 (N1291, N1271, N111);
xor XOR2 (N1292, N1280, N940);
nor NOR2 (N1293, N1285, N801);
nand NAND3 (N1294, N1261, N723, N873);
and AND2 (N1295, N1290, N1244);
and AND3 (N1296, N1279, N1077, N432);
buf BUF1 (N1297, N1296);
nand NAND2 (N1298, N1295, N540);
buf BUF1 (N1299, N1294);
not NOT1 (N1300, N1291);
not NOT1 (N1301, N1246);
buf BUF1 (N1302, N1289);
nand NAND2 (N1303, N1301, N201);
and AND3 (N1304, N1298, N1138, N1277);
nand NAND4 (N1305, N1288, N315, N126, N1302);
nand NAND3 (N1306, N292, N1109, N219);
buf BUF1 (N1307, N1297);
and AND4 (N1308, N1300, N784, N725, N168);
buf BUF1 (N1309, N1307);
xor XOR2 (N1310, N1299, N134);
or OR2 (N1311, N1305, N390);
or OR4 (N1312, N1293, N132, N339, N1147);
nand NAND4 (N1313, N1312, N924, N368, N1125);
xor XOR2 (N1314, N1309, N975);
nor NOR4 (N1315, N1314, N928, N652, N499);
not NOT1 (N1316, N1311);
not NOT1 (N1317, N1304);
xor XOR2 (N1318, N1317, N416);
buf BUF1 (N1319, N1315);
nand NAND3 (N1320, N1273, N41, N224);
nand NAND2 (N1321, N1308, N332);
nor NOR2 (N1322, N1321, N19);
nor NOR3 (N1323, N1320, N205, N220);
nand NAND3 (N1324, N1310, N1158, N450);
nand NAND3 (N1325, N1318, N297, N980);
nand NAND4 (N1326, N1292, N723, N284, N709);
nand NAND4 (N1327, N1324, N608, N1142, N910);
nand NAND2 (N1328, N1327, N699);
nand NAND2 (N1329, N1319, N586);
nor NOR3 (N1330, N1303, N736, N78);
not NOT1 (N1331, N1313);
nand NAND2 (N1332, N1331, N1195);
xor XOR2 (N1333, N1316, N159);
or OR4 (N1334, N1328, N18, N1214, N498);
not NOT1 (N1335, N1334);
xor XOR2 (N1336, N1335, N930);
nor NOR4 (N1337, N1306, N787, N1163, N193);
nand NAND3 (N1338, N1323, N1293, N776);
nand NAND3 (N1339, N1329, N808, N845);
xor XOR2 (N1340, N1330, N45);
and AND4 (N1341, N1338, N1322, N840, N527);
nand NAND3 (N1342, N363, N485, N665);
nor NOR2 (N1343, N1332, N506);
nor NOR4 (N1344, N1336, N1330, N861, N919);
not NOT1 (N1345, N1337);
not NOT1 (N1346, N1340);
nand NAND3 (N1347, N1346, N611, N877);
not NOT1 (N1348, N1341);
not NOT1 (N1349, N1325);
or OR4 (N1350, N1345, N774, N286, N1038);
and AND4 (N1351, N1333, N116, N185, N241);
buf BUF1 (N1352, N1342);
and AND4 (N1353, N1326, N940, N571, N261);
buf BUF1 (N1354, N1343);
and AND3 (N1355, N1344, N1333, N820);
nor NOR3 (N1356, N1348, N904, N627);
or OR2 (N1357, N1349, N460);
buf BUF1 (N1358, N1351);
buf BUF1 (N1359, N1356);
nand NAND4 (N1360, N1358, N164, N665, N476);
buf BUF1 (N1361, N1354);
not NOT1 (N1362, N1352);
or OR3 (N1363, N1362, N567, N1150);
buf BUF1 (N1364, N1350);
buf BUF1 (N1365, N1353);
nor NOR4 (N1366, N1363, N1292, N437, N370);
and AND3 (N1367, N1364, N692, N755);
and AND3 (N1368, N1361, N180, N312);
and AND3 (N1369, N1366, N427, N509);
and AND2 (N1370, N1367, N1082);
buf BUF1 (N1371, N1368);
and AND3 (N1372, N1347, N403, N301);
xor XOR2 (N1373, N1371, N137);
and AND3 (N1374, N1373, N1192, N1102);
buf BUF1 (N1375, N1372);
xor XOR2 (N1376, N1365, N735);
or OR4 (N1377, N1357, N970, N418, N129);
or OR4 (N1378, N1374, N1085, N308, N443);
and AND2 (N1379, N1377, N227);
xor XOR2 (N1380, N1370, N303);
xor XOR2 (N1381, N1360, N280);
and AND3 (N1382, N1375, N831, N232);
or OR2 (N1383, N1339, N1161);
nor NOR4 (N1384, N1355, N1191, N724, N468);
not NOT1 (N1385, N1383);
or OR2 (N1386, N1380, N216);
xor XOR2 (N1387, N1369, N520);
nor NOR2 (N1388, N1385, N99);
or OR3 (N1389, N1384, N20, N662);
nand NAND2 (N1390, N1382, N657);
buf BUF1 (N1391, N1388);
or OR2 (N1392, N1381, N1326);
nand NAND4 (N1393, N1390, N957, N788, N639);
xor XOR2 (N1394, N1386, N393);
or OR4 (N1395, N1359, N667, N127, N294);
nand NAND4 (N1396, N1391, N212, N249, N1266);
and AND2 (N1397, N1394, N674);
nor NOR2 (N1398, N1389, N1358);
not NOT1 (N1399, N1398);
xor XOR2 (N1400, N1396, N479);
not NOT1 (N1401, N1400);
nor NOR2 (N1402, N1376, N628);
not NOT1 (N1403, N1387);
not NOT1 (N1404, N1392);
nor NOR4 (N1405, N1395, N970, N452, N77);
or OR3 (N1406, N1399, N660, N212);
buf BUF1 (N1407, N1397);
xor XOR2 (N1408, N1393, N168);
and AND3 (N1409, N1379, N755, N792);
or OR3 (N1410, N1378, N80, N1358);
nor NOR4 (N1411, N1402, N415, N684, N584);
not NOT1 (N1412, N1404);
or OR2 (N1413, N1410, N629);
nand NAND4 (N1414, N1408, N480, N378, N1188);
and AND2 (N1415, N1412, N1348);
nor NOR4 (N1416, N1414, N615, N749, N194);
xor XOR2 (N1417, N1415, N607);
nand NAND2 (N1418, N1416, N1275);
not NOT1 (N1419, N1418);
buf BUF1 (N1420, N1407);
or OR3 (N1421, N1419, N982, N404);
and AND3 (N1422, N1403, N1243, N994);
and AND2 (N1423, N1409, N243);
or OR2 (N1424, N1405, N1333);
or OR3 (N1425, N1421, N264, N798);
xor XOR2 (N1426, N1420, N1232);
nor NOR3 (N1427, N1413, N1249, N854);
or OR4 (N1428, N1401, N97, N1074, N521);
or OR2 (N1429, N1428, N1031);
or OR3 (N1430, N1424, N972, N364);
xor XOR2 (N1431, N1429, N1033);
or OR3 (N1432, N1411, N292, N424);
xor XOR2 (N1433, N1430, N73);
buf BUF1 (N1434, N1417);
not NOT1 (N1435, N1433);
nor NOR4 (N1436, N1423, N845, N527, N5);
not NOT1 (N1437, N1426);
buf BUF1 (N1438, N1436);
xor XOR2 (N1439, N1432, N477);
xor XOR2 (N1440, N1439, N255);
buf BUF1 (N1441, N1427);
xor XOR2 (N1442, N1434, N901);
xor XOR2 (N1443, N1406, N314);
nand NAND4 (N1444, N1437, N168, N339, N1431);
xor XOR2 (N1445, N968, N743);
not NOT1 (N1446, N1422);
nand NAND4 (N1447, N1445, N829, N1327, N667);
or OR2 (N1448, N1447, N1068);
buf BUF1 (N1449, N1438);
or OR4 (N1450, N1435, N33, N382, N878);
nor NOR3 (N1451, N1441, N213, N357);
nor NOR2 (N1452, N1451, N1264);
not NOT1 (N1453, N1425);
nand NAND2 (N1454, N1448, N5);
xor XOR2 (N1455, N1449, N513);
nor NOR2 (N1456, N1442, N1331);
buf BUF1 (N1457, N1456);
nand NAND2 (N1458, N1452, N465);
nand NAND3 (N1459, N1440, N275, N1019);
xor XOR2 (N1460, N1457, N429);
buf BUF1 (N1461, N1460);
buf BUF1 (N1462, N1454);
not NOT1 (N1463, N1458);
nor NOR4 (N1464, N1443, N181, N976, N1307);
nand NAND4 (N1465, N1444, N831, N520, N355);
nor NOR3 (N1466, N1464, N741, N363);
nor NOR2 (N1467, N1461, N1463);
nor NOR3 (N1468, N579, N625, N19);
nand NAND3 (N1469, N1467, N284, N336);
nor NOR4 (N1470, N1468, N1380, N1408, N588);
buf BUF1 (N1471, N1462);
nor NOR3 (N1472, N1455, N296, N119);
buf BUF1 (N1473, N1446);
nor NOR2 (N1474, N1465, N827);
or OR3 (N1475, N1471, N1320, N758);
xor XOR2 (N1476, N1459, N507);
nand NAND2 (N1477, N1466, N676);
xor XOR2 (N1478, N1472, N437);
not NOT1 (N1479, N1477);
and AND3 (N1480, N1453, N1451, N359);
and AND2 (N1481, N1450, N597);
nor NOR3 (N1482, N1480, N1354, N1466);
not NOT1 (N1483, N1474);
nor NOR4 (N1484, N1482, N603, N1089, N1036);
and AND2 (N1485, N1484, N251);
buf BUF1 (N1486, N1478);
or OR2 (N1487, N1469, N1013);
not NOT1 (N1488, N1481);
and AND4 (N1489, N1479, N1328, N776, N664);
xor XOR2 (N1490, N1475, N849);
buf BUF1 (N1491, N1483);
nor NOR2 (N1492, N1491, N1429);
or OR2 (N1493, N1489, N449);
or OR4 (N1494, N1486, N546, N10, N1417);
nor NOR4 (N1495, N1470, N1252, N854, N1201);
nor NOR3 (N1496, N1493, N975, N1186);
nor NOR4 (N1497, N1485, N823, N715, N568);
or OR4 (N1498, N1488, N733, N174, N510);
nand NAND2 (N1499, N1495, N523);
nor NOR3 (N1500, N1490, N635, N500);
or OR3 (N1501, N1499, N393, N706);
nor NOR3 (N1502, N1498, N1010, N1309);
not NOT1 (N1503, N1501);
and AND2 (N1504, N1503, N733);
buf BUF1 (N1505, N1497);
and AND3 (N1506, N1505, N1110, N244);
not NOT1 (N1507, N1473);
or OR4 (N1508, N1506, N212, N531, N1144);
or OR4 (N1509, N1496, N1479, N971, N753);
or OR2 (N1510, N1492, N1161);
buf BUF1 (N1511, N1487);
not NOT1 (N1512, N1476);
nand NAND4 (N1513, N1502, N1034, N571, N320);
and AND3 (N1514, N1513, N641, N1439);
nand NAND3 (N1515, N1511, N508, N1475);
nor NOR4 (N1516, N1494, N971, N860, N793);
or OR2 (N1517, N1510, N1070);
not NOT1 (N1518, N1504);
nand NAND2 (N1519, N1512, N268);
buf BUF1 (N1520, N1500);
not NOT1 (N1521, N1507);
not NOT1 (N1522, N1508);
or OR3 (N1523, N1516, N56, N1026);
nor NOR4 (N1524, N1509, N159, N469, N1032);
buf BUF1 (N1525, N1522);
not NOT1 (N1526, N1519);
buf BUF1 (N1527, N1523);
buf BUF1 (N1528, N1520);
and AND2 (N1529, N1525, N1399);
or OR2 (N1530, N1521, N1066);
and AND4 (N1531, N1517, N475, N1369, N73);
nand NAND4 (N1532, N1530, N1111, N264, N1022);
nand NAND3 (N1533, N1532, N204, N79);
or OR3 (N1534, N1526, N55, N99);
not NOT1 (N1535, N1518);
nand NAND4 (N1536, N1534, N1239, N893, N143);
nor NOR3 (N1537, N1533, N518, N587);
nand NAND4 (N1538, N1535, N1344, N489, N1146);
or OR4 (N1539, N1531, N1410, N1057, N1514);
or OR2 (N1540, N731, N790);
buf BUF1 (N1541, N1527);
or OR4 (N1542, N1537, N496, N1114, N146);
buf BUF1 (N1543, N1536);
and AND2 (N1544, N1541, N1434);
xor XOR2 (N1545, N1529, N583);
nor NOR2 (N1546, N1515, N331);
nor NOR4 (N1547, N1545, N332, N1227, N575);
and AND3 (N1548, N1546, N344, N508);
nand NAND4 (N1549, N1524, N835, N609, N545);
or OR4 (N1550, N1543, N750, N1038, N1049);
nor NOR3 (N1551, N1540, N1372, N410);
buf BUF1 (N1552, N1549);
nand NAND2 (N1553, N1551, N1139);
xor XOR2 (N1554, N1548, N547);
xor XOR2 (N1555, N1550, N186);
and AND4 (N1556, N1538, N46, N912, N1146);
or OR4 (N1557, N1556, N1272, N1148, N1273);
nand NAND3 (N1558, N1539, N185, N985);
and AND2 (N1559, N1547, N604);
xor XOR2 (N1560, N1558, N1279);
and AND2 (N1561, N1557, N1419);
buf BUF1 (N1562, N1544);
nor NOR4 (N1563, N1555, N147, N826, N935);
and AND4 (N1564, N1560, N1016, N630, N526);
buf BUF1 (N1565, N1552);
nand NAND4 (N1566, N1563, N433, N420, N1277);
not NOT1 (N1567, N1566);
or OR4 (N1568, N1565, N1280, N1333, N937);
or OR3 (N1569, N1528, N742, N982);
nor NOR3 (N1570, N1542, N1007, N749);
buf BUF1 (N1571, N1567);
buf BUF1 (N1572, N1553);
buf BUF1 (N1573, N1561);
not NOT1 (N1574, N1571);
xor XOR2 (N1575, N1564, N1292);
not NOT1 (N1576, N1559);
buf BUF1 (N1577, N1568);
nor NOR2 (N1578, N1572, N274);
xor XOR2 (N1579, N1554, N199);
nor NOR4 (N1580, N1576, N888, N316, N1560);
nand NAND2 (N1581, N1573, N367);
buf BUF1 (N1582, N1562);
and AND2 (N1583, N1582, N1410);
or OR4 (N1584, N1581, N652, N1276, N334);
not NOT1 (N1585, N1580);
not NOT1 (N1586, N1574);
buf BUF1 (N1587, N1578);
nor NOR2 (N1588, N1575, N434);
xor XOR2 (N1589, N1588, N1041);
and AND4 (N1590, N1583, N1135, N1434, N510);
not NOT1 (N1591, N1569);
buf BUF1 (N1592, N1577);
nor NOR4 (N1593, N1584, N1398, N798, N140);
nand NAND2 (N1594, N1585, N1285);
and AND4 (N1595, N1592, N307, N1193, N627);
not NOT1 (N1596, N1586);
buf BUF1 (N1597, N1591);
xor XOR2 (N1598, N1579, N1040);
xor XOR2 (N1599, N1587, N1159);
buf BUF1 (N1600, N1590);
not NOT1 (N1601, N1570);
nor NOR2 (N1602, N1597, N703);
nand NAND4 (N1603, N1600, N742, N616, N219);
nor NOR4 (N1604, N1599, N1218, N870, N345);
not NOT1 (N1605, N1602);
nand NAND4 (N1606, N1596, N654, N1500, N822);
and AND3 (N1607, N1601, N1131, N737);
nand NAND3 (N1608, N1603, N877, N1304);
nor NOR3 (N1609, N1595, N328, N1268);
xor XOR2 (N1610, N1607, N568);
buf BUF1 (N1611, N1604);
xor XOR2 (N1612, N1609, N375);
or OR2 (N1613, N1612, N162);
and AND4 (N1614, N1608, N629, N1402, N1360);
nand NAND3 (N1615, N1589, N1596, N445);
nand NAND3 (N1616, N1610, N227, N1146);
or OR2 (N1617, N1616, N123);
xor XOR2 (N1618, N1611, N1555);
nand NAND4 (N1619, N1594, N983, N1155, N800);
not NOT1 (N1620, N1593);
nor NOR4 (N1621, N1618, N289, N401, N514);
nand NAND2 (N1622, N1598, N169);
not NOT1 (N1623, N1605);
nor NOR4 (N1624, N1614, N558, N1578, N1312);
xor XOR2 (N1625, N1613, N241);
nand NAND4 (N1626, N1625, N1261, N1231, N71);
nand NAND4 (N1627, N1606, N1100, N1027, N809);
not NOT1 (N1628, N1626);
or OR3 (N1629, N1628, N1106, N973);
not NOT1 (N1630, N1620);
buf BUF1 (N1631, N1617);
not NOT1 (N1632, N1622);
nand NAND4 (N1633, N1619, N830, N208, N322);
xor XOR2 (N1634, N1631, N481);
not NOT1 (N1635, N1627);
or OR2 (N1636, N1623, N515);
or OR3 (N1637, N1624, N546, N1071);
nor NOR2 (N1638, N1621, N63);
or OR3 (N1639, N1635, N364, N983);
nand NAND3 (N1640, N1634, N522, N79);
xor XOR2 (N1641, N1629, N339);
not NOT1 (N1642, N1638);
nor NOR4 (N1643, N1615, N604, N208, N1356);
nand NAND3 (N1644, N1641, N1503, N1384);
nor NOR4 (N1645, N1640, N214, N342, N1027);
nand NAND3 (N1646, N1639, N134, N1113);
nor NOR2 (N1647, N1632, N1138);
xor XOR2 (N1648, N1637, N1020);
buf BUF1 (N1649, N1648);
not NOT1 (N1650, N1636);
buf BUF1 (N1651, N1642);
xor XOR2 (N1652, N1644, N1441);
buf BUF1 (N1653, N1643);
or OR2 (N1654, N1633, N267);
xor XOR2 (N1655, N1653, N475);
nor NOR4 (N1656, N1654, N1508, N347, N1329);
and AND2 (N1657, N1655, N861);
buf BUF1 (N1658, N1657);
xor XOR2 (N1659, N1646, N1630);
not NOT1 (N1660, N26);
not NOT1 (N1661, N1656);
nand NAND4 (N1662, N1652, N406, N1441, N1639);
and AND3 (N1663, N1649, N257, N9);
and AND4 (N1664, N1663, N1141, N1329, N718);
xor XOR2 (N1665, N1660, N1044);
or OR3 (N1666, N1664, N881, N1658);
not NOT1 (N1667, N558);
xor XOR2 (N1668, N1650, N929);
nor NOR4 (N1669, N1647, N1154, N676, N619);
or OR3 (N1670, N1645, N324, N1606);
not NOT1 (N1671, N1651);
xor XOR2 (N1672, N1666, N1110);
nand NAND2 (N1673, N1659, N773);
nand NAND4 (N1674, N1673, N1469, N44, N298);
buf BUF1 (N1675, N1661);
not NOT1 (N1676, N1669);
nand NAND3 (N1677, N1662, N1161, N1122);
and AND4 (N1678, N1665, N1509, N439, N393);
xor XOR2 (N1679, N1676, N1037);
and AND4 (N1680, N1668, N629, N1032, N396);
xor XOR2 (N1681, N1678, N1627);
xor XOR2 (N1682, N1671, N926);
nor NOR3 (N1683, N1674, N895, N992);
and AND4 (N1684, N1680, N1110, N1483, N1172);
xor XOR2 (N1685, N1683, N1051);
xor XOR2 (N1686, N1679, N796);
nor NOR2 (N1687, N1675, N1056);
and AND2 (N1688, N1681, N365);
nand NAND3 (N1689, N1687, N321, N1588);
nor NOR3 (N1690, N1677, N275, N1330);
or OR4 (N1691, N1672, N216, N417, N1195);
nand NAND2 (N1692, N1684, N1283);
and AND4 (N1693, N1688, N451, N176, N1594);
and AND4 (N1694, N1686, N1108, N146, N497);
nand NAND3 (N1695, N1692, N1335, N1640);
buf BUF1 (N1696, N1689);
xor XOR2 (N1697, N1670, N250);
nand NAND4 (N1698, N1667, N961, N753, N1006);
and AND3 (N1699, N1690, N955, N87);
buf BUF1 (N1700, N1694);
nor NOR4 (N1701, N1696, N1397, N200, N5);
or OR3 (N1702, N1691, N543, N1017);
not NOT1 (N1703, N1695);
nand NAND2 (N1704, N1693, N645);
and AND2 (N1705, N1702, N1002);
nand NAND4 (N1706, N1705, N49, N246, N594);
xor XOR2 (N1707, N1699, N337);
xor XOR2 (N1708, N1701, N1214);
or OR2 (N1709, N1700, N511);
xor XOR2 (N1710, N1707, N1675);
not NOT1 (N1711, N1697);
nand NAND3 (N1712, N1698, N910, N1267);
xor XOR2 (N1713, N1685, N732);
or OR4 (N1714, N1706, N834, N704, N1682);
buf BUF1 (N1715, N1389);
nor NOR3 (N1716, N1714, N411, N339);
buf BUF1 (N1717, N1708);
xor XOR2 (N1718, N1712, N41);
nand NAND2 (N1719, N1715, N1671);
and AND3 (N1720, N1718, N294, N690);
or OR4 (N1721, N1709, N351, N385, N451);
or OR3 (N1722, N1717, N1407, N933);
not NOT1 (N1723, N1720);
xor XOR2 (N1724, N1716, N1170);
and AND3 (N1725, N1704, N638, N113);
xor XOR2 (N1726, N1711, N1170);
and AND3 (N1727, N1722, N851, N1191);
nor NOR3 (N1728, N1703, N1085, N1292);
nor NOR4 (N1729, N1719, N837, N1080, N1493);
or OR3 (N1730, N1713, N1665, N1314);
not NOT1 (N1731, N1730);
and AND4 (N1732, N1729, N1213, N510, N107);
or OR3 (N1733, N1710, N880, N1533);
nand NAND2 (N1734, N1723, N1072);
or OR3 (N1735, N1728, N1571, N1337);
or OR4 (N1736, N1734, N326, N1124, N836);
xor XOR2 (N1737, N1721, N598);
or OR4 (N1738, N1727, N1449, N1165, N798);
nand NAND4 (N1739, N1733, N677, N1546, N886);
buf BUF1 (N1740, N1736);
nand NAND3 (N1741, N1735, N735, N1722);
buf BUF1 (N1742, N1741);
and AND3 (N1743, N1724, N871, N1454);
or OR3 (N1744, N1731, N1314, N1494);
buf BUF1 (N1745, N1740);
nand NAND4 (N1746, N1745, N312, N1391, N1065);
and AND4 (N1747, N1744, N1247, N1102, N1599);
xor XOR2 (N1748, N1737, N573);
nand NAND3 (N1749, N1732, N770, N1662);
nand NAND2 (N1750, N1746, N594);
nand NAND4 (N1751, N1725, N867, N1572, N742);
nor NOR4 (N1752, N1748, N434, N1210, N850);
nand NAND2 (N1753, N1750, N1641);
or OR2 (N1754, N1752, N735);
nand NAND3 (N1755, N1749, N32, N1637);
nand NAND4 (N1756, N1747, N789, N1064, N603);
nand NAND4 (N1757, N1726, N488, N88, N831);
not NOT1 (N1758, N1756);
nand NAND3 (N1759, N1758, N302, N1488);
or OR2 (N1760, N1743, N896);
xor XOR2 (N1761, N1759, N1697);
not NOT1 (N1762, N1760);
and AND4 (N1763, N1742, N1298, N70, N1300);
nor NOR2 (N1764, N1751, N523);
not NOT1 (N1765, N1755);
xor XOR2 (N1766, N1761, N750);
not NOT1 (N1767, N1762);
and AND3 (N1768, N1753, N903, N198);
nor NOR4 (N1769, N1763, N1734, N1690, N846);
not NOT1 (N1770, N1768);
nand NAND2 (N1771, N1764, N1490);
or OR3 (N1772, N1766, N1117, N282);
nand NAND4 (N1773, N1765, N1640, N251, N772);
nor NOR2 (N1774, N1769, N1471);
nand NAND2 (N1775, N1754, N790);
buf BUF1 (N1776, N1775);
and AND4 (N1777, N1739, N368, N9, N1408);
nand NAND4 (N1778, N1771, N1668, N453, N805);
buf BUF1 (N1779, N1773);
nand NAND3 (N1780, N1774, N792, N589);
nor NOR4 (N1781, N1770, N216, N1128, N969);
and AND3 (N1782, N1757, N1745, N1188);
not NOT1 (N1783, N1767);
nor NOR3 (N1784, N1781, N72, N1173);
nor NOR4 (N1785, N1772, N1144, N880, N982);
nand NAND3 (N1786, N1779, N44, N848);
buf BUF1 (N1787, N1777);
nor NOR3 (N1788, N1784, N663, N1712);
xor XOR2 (N1789, N1788, N72);
xor XOR2 (N1790, N1787, N1443);
nand NAND2 (N1791, N1785, N143);
not NOT1 (N1792, N1789);
xor XOR2 (N1793, N1782, N1694);
or OR2 (N1794, N1783, N1268);
xor XOR2 (N1795, N1790, N1090);
not NOT1 (N1796, N1738);
xor XOR2 (N1797, N1791, N1691);
buf BUF1 (N1798, N1786);
buf BUF1 (N1799, N1796);
nor NOR3 (N1800, N1778, N1626, N459);
nor NOR2 (N1801, N1799, N1589);
or OR3 (N1802, N1776, N1581, N691);
xor XOR2 (N1803, N1780, N134);
nand NAND4 (N1804, N1794, N324, N1444, N1206);
nand NAND2 (N1805, N1803, N977);
and AND4 (N1806, N1798, N396, N1627, N1147);
and AND4 (N1807, N1792, N1148, N1519, N1302);
buf BUF1 (N1808, N1805);
nor NOR2 (N1809, N1797, N1209);
not NOT1 (N1810, N1801);
or OR3 (N1811, N1810, N95, N1624);
xor XOR2 (N1812, N1806, N326);
and AND4 (N1813, N1800, N178, N1551, N157);
xor XOR2 (N1814, N1793, N1595);
or OR4 (N1815, N1814, N177, N1284, N1512);
nor NOR4 (N1816, N1811, N1602, N1387, N1719);
and AND3 (N1817, N1813, N1138, N95);
buf BUF1 (N1818, N1802);
nor NOR3 (N1819, N1809, N1194, N821);
nor NOR4 (N1820, N1807, N1417, N448, N898);
xor XOR2 (N1821, N1819, N662);
nand NAND4 (N1822, N1808, N662, N790, N645);
or OR2 (N1823, N1817, N357);
xor XOR2 (N1824, N1818, N145);
nor NOR4 (N1825, N1815, N911, N1254, N627);
nand NAND2 (N1826, N1823, N1557);
nor NOR2 (N1827, N1812, N468);
or OR2 (N1828, N1822, N173);
and AND4 (N1829, N1816, N1620, N1253, N1007);
and AND4 (N1830, N1824, N1647, N924, N390);
nand NAND4 (N1831, N1827, N638, N1753, N924);
and AND4 (N1832, N1830, N850, N1171, N1629);
xor XOR2 (N1833, N1795, N1640);
and AND4 (N1834, N1804, N786, N529, N943);
nand NAND2 (N1835, N1833, N1511);
xor XOR2 (N1836, N1825, N914);
not NOT1 (N1837, N1831);
not NOT1 (N1838, N1836);
not NOT1 (N1839, N1832);
buf BUF1 (N1840, N1839);
not NOT1 (N1841, N1835);
not NOT1 (N1842, N1841);
or OR2 (N1843, N1837, N1664);
or OR3 (N1844, N1829, N1811, N439);
xor XOR2 (N1845, N1838, N1590);
nor NOR2 (N1846, N1843, N644);
buf BUF1 (N1847, N1820);
and AND4 (N1848, N1847, N827, N1139, N1842);
and AND2 (N1849, N1274, N735);
nor NOR3 (N1850, N1821, N143, N704);
nor NOR3 (N1851, N1846, N238, N171);
nor NOR2 (N1852, N1844, N757);
buf BUF1 (N1853, N1848);
and AND3 (N1854, N1853, N971, N235);
xor XOR2 (N1855, N1849, N995);
buf BUF1 (N1856, N1851);
nand NAND4 (N1857, N1828, N1753, N1395, N1555);
or OR4 (N1858, N1845, N838, N704, N1677);
or OR4 (N1859, N1854, N771, N189, N1348);
or OR2 (N1860, N1840, N119);
xor XOR2 (N1861, N1826, N1624);
nor NOR3 (N1862, N1834, N1454, N398);
not NOT1 (N1863, N1850);
nor NOR4 (N1864, N1858, N1737, N1105, N377);
not NOT1 (N1865, N1855);
xor XOR2 (N1866, N1859, N532);
buf BUF1 (N1867, N1857);
not NOT1 (N1868, N1860);
nor NOR3 (N1869, N1861, N1439, N643);
and AND4 (N1870, N1862, N1496, N266, N1751);
xor XOR2 (N1871, N1865, N1307);
xor XOR2 (N1872, N1870, N17);
nor NOR3 (N1873, N1867, N1227, N1656);
not NOT1 (N1874, N1869);
not NOT1 (N1875, N1864);
buf BUF1 (N1876, N1873);
nor NOR3 (N1877, N1871, N774, N1110);
xor XOR2 (N1878, N1875, N6);
nand NAND4 (N1879, N1874, N1375, N1102, N896);
buf BUF1 (N1880, N1863);
or OR2 (N1881, N1866, N1730);
and AND4 (N1882, N1880, N326, N1017, N1327);
nor NOR2 (N1883, N1879, N493);
and AND3 (N1884, N1878, N416, N380);
and AND3 (N1885, N1876, N522, N1625);
and AND3 (N1886, N1884, N1184, N625);
and AND2 (N1887, N1856, N804);
buf BUF1 (N1888, N1886);
nor NOR4 (N1889, N1852, N1338, N1352, N1044);
nand NAND3 (N1890, N1883, N1055, N1804);
and AND3 (N1891, N1877, N82, N790);
nor NOR4 (N1892, N1882, N1434, N1765, N618);
not NOT1 (N1893, N1891);
not NOT1 (N1894, N1872);
nand NAND2 (N1895, N1868, N1128);
buf BUF1 (N1896, N1893);
or OR3 (N1897, N1889, N885, N830);
or OR2 (N1898, N1888, N1223);
nor NOR3 (N1899, N1890, N1329, N949);
and AND3 (N1900, N1885, N1436, N20);
and AND3 (N1901, N1887, N131, N318);
nand NAND2 (N1902, N1898, N870);
and AND3 (N1903, N1894, N900, N1457);
nand NAND3 (N1904, N1901, N1742, N248);
buf BUF1 (N1905, N1902);
buf BUF1 (N1906, N1892);
and AND4 (N1907, N1903, N1092, N1668, N890);
and AND3 (N1908, N1906, N1244, N1105);
nand NAND3 (N1909, N1908, N214, N813);
nor NOR3 (N1910, N1905, N554, N684);
not NOT1 (N1911, N1896);
and AND2 (N1912, N1895, N548);
and AND2 (N1913, N1881, N487);
buf BUF1 (N1914, N1909);
xor XOR2 (N1915, N1907, N1652);
nand NAND3 (N1916, N1912, N1068, N1415);
nand NAND3 (N1917, N1899, N766, N1648);
nand NAND4 (N1918, N1914, N571, N1315, N580);
buf BUF1 (N1919, N1904);
not NOT1 (N1920, N1918);
buf BUF1 (N1921, N1913);
nor NOR4 (N1922, N1921, N971, N824, N946);
xor XOR2 (N1923, N1919, N538);
nand NAND3 (N1924, N1911, N629, N1664);
nor NOR4 (N1925, N1897, N1596, N888, N961);
not NOT1 (N1926, N1900);
xor XOR2 (N1927, N1926, N1159);
not NOT1 (N1928, N1924);
xor XOR2 (N1929, N1915, N328);
nand NAND3 (N1930, N1928, N965, N164);
or OR4 (N1931, N1930, N236, N1501, N1210);
and AND4 (N1932, N1917, N438, N1678, N1863);
buf BUF1 (N1933, N1927);
and AND3 (N1934, N1916, N353, N1323);
not NOT1 (N1935, N1932);
and AND3 (N1936, N1929, N1332, N1564);
or OR4 (N1937, N1923, N1556, N597, N1389);
not NOT1 (N1938, N1934);
nand NAND2 (N1939, N1922, N1157);
nand NAND2 (N1940, N1925, N831);
and AND3 (N1941, N1937, N963, N583);
not NOT1 (N1942, N1938);
or OR4 (N1943, N1942, N1659, N103, N267);
xor XOR2 (N1944, N1910, N1134);
not NOT1 (N1945, N1943);
not NOT1 (N1946, N1935);
and AND4 (N1947, N1939, N1329, N1119, N416);
not NOT1 (N1948, N1941);
or OR3 (N1949, N1948, N429, N881);
and AND4 (N1950, N1940, N1764, N817, N278);
not NOT1 (N1951, N1920);
buf BUF1 (N1952, N1931);
xor XOR2 (N1953, N1952, N909);
or OR2 (N1954, N1949, N783);
nand NAND2 (N1955, N1945, N548);
and AND2 (N1956, N1953, N1451);
nor NOR2 (N1957, N1954, N1130);
and AND3 (N1958, N1957, N1765, N1874);
nand NAND3 (N1959, N1951, N1063, N1389);
nor NOR4 (N1960, N1956, N555, N1451, N1897);
and AND4 (N1961, N1955, N408, N704, N809);
xor XOR2 (N1962, N1944, N806);
and AND4 (N1963, N1960, N1688, N359, N960);
buf BUF1 (N1964, N1936);
xor XOR2 (N1965, N1963, N442);
xor XOR2 (N1966, N1946, N924);
or OR3 (N1967, N1959, N1782, N717);
nand NAND2 (N1968, N1964, N1824);
buf BUF1 (N1969, N1958);
nor NOR4 (N1970, N1966, N1058, N592, N1735);
nor NOR3 (N1971, N1947, N1793, N1491);
nor NOR2 (N1972, N1968, N1387);
or OR2 (N1973, N1971, N81);
nand NAND2 (N1974, N1965, N777);
nand NAND4 (N1975, N1950, N1101, N844, N1212);
xor XOR2 (N1976, N1969, N699);
not NOT1 (N1977, N1972);
buf BUF1 (N1978, N1967);
and AND4 (N1979, N1933, N722, N723, N810);
xor XOR2 (N1980, N1978, N583);
nand NAND2 (N1981, N1976, N372);
nand NAND4 (N1982, N1973, N544, N274, N1068);
not NOT1 (N1983, N1982);
or OR3 (N1984, N1977, N838, N385);
and AND3 (N1985, N1983, N223, N1817);
nor NOR3 (N1986, N1974, N832, N193);
and AND3 (N1987, N1980, N236, N158);
and AND4 (N1988, N1986, N501, N397, N668);
nor NOR4 (N1989, N1975, N156, N1106, N87);
nand NAND4 (N1990, N1979, N193, N1650, N1534);
nor NOR2 (N1991, N1984, N1392);
and AND2 (N1992, N1988, N919);
not NOT1 (N1993, N1985);
and AND3 (N1994, N1989, N252, N1856);
buf BUF1 (N1995, N1990);
not NOT1 (N1996, N1970);
not NOT1 (N1997, N1994);
xor XOR2 (N1998, N1991, N1179);
nand NAND4 (N1999, N1995, N1634, N1961, N417);
or OR3 (N2000, N1623, N328, N1436);
xor XOR2 (N2001, N1999, N1987);
or OR2 (N2002, N1506, N1882);
and AND4 (N2003, N1992, N1471, N806, N1547);
buf BUF1 (N2004, N2002);
xor XOR2 (N2005, N1962, N1401);
and AND2 (N2006, N1998, N1401);
xor XOR2 (N2007, N2005, N748);
xor XOR2 (N2008, N1993, N1457);
or OR2 (N2009, N2000, N619);
nand NAND2 (N2010, N2008, N436);
or OR3 (N2011, N2007, N984, N1623);
and AND4 (N2012, N1981, N410, N1885, N1900);
or OR4 (N2013, N2001, N1735, N1913, N1295);
not NOT1 (N2014, N2006);
or OR3 (N2015, N2011, N753, N1855);
or OR4 (N2016, N2012, N1671, N1223, N249);
and AND4 (N2017, N2003, N1817, N1416, N1290);
not NOT1 (N2018, N2010);
nor NOR4 (N2019, N2009, N1032, N1289, N838);
and AND3 (N2020, N1997, N981, N3);
and AND3 (N2021, N2018, N1555, N1510);
xor XOR2 (N2022, N2016, N321);
nor NOR2 (N2023, N1996, N1191);
xor XOR2 (N2024, N2017, N1118);
nand NAND2 (N2025, N2019, N1005);
and AND4 (N2026, N2020, N26, N1876, N1687);
nor NOR4 (N2027, N2015, N1187, N874, N1069);
and AND2 (N2028, N2025, N140);
and AND3 (N2029, N2004, N1611, N1727);
buf BUF1 (N2030, N2024);
not NOT1 (N2031, N2022);
xor XOR2 (N2032, N2030, N1586);
nor NOR3 (N2033, N2032, N856, N370);
buf BUF1 (N2034, N2031);
or OR4 (N2035, N2029, N712, N558, N1487);
buf BUF1 (N2036, N2028);
or OR4 (N2037, N2036, N116, N349, N711);
nand NAND2 (N2038, N2037, N637);
xor XOR2 (N2039, N2021, N350);
nand NAND4 (N2040, N2035, N1960, N1143, N911);
buf BUF1 (N2041, N2039);
and AND4 (N2042, N2027, N102, N1510, N943);
or OR2 (N2043, N2023, N1747);
nand NAND3 (N2044, N2014, N487, N1271);
buf BUF1 (N2045, N2042);
not NOT1 (N2046, N2045);
and AND2 (N2047, N2041, N1263);
nand NAND2 (N2048, N2026, N848);
or OR3 (N2049, N2033, N735, N484);
not NOT1 (N2050, N2047);
or OR2 (N2051, N2049, N1214);
or OR3 (N2052, N2048, N16, N1128);
xor XOR2 (N2053, N2046, N1235);
xor XOR2 (N2054, N2013, N1176);
and AND4 (N2055, N2053, N1820, N628, N1262);
nor NOR3 (N2056, N2052, N1377, N1602);
or OR4 (N2057, N2054, N189, N1197, N1685);
nand NAND2 (N2058, N2044, N827);
buf BUF1 (N2059, N2056);
nand NAND4 (N2060, N2050, N1612, N1481, N1391);
nand NAND2 (N2061, N2034, N1817);
not NOT1 (N2062, N2057);
or OR2 (N2063, N2060, N562);
xor XOR2 (N2064, N2055, N1890);
nor NOR3 (N2065, N2059, N1939, N1922);
nand NAND3 (N2066, N2051, N893, N1547);
xor XOR2 (N2067, N2062, N1466);
not NOT1 (N2068, N2066);
not NOT1 (N2069, N2063);
and AND3 (N2070, N2058, N1308, N1884);
nand NAND4 (N2071, N2038, N92, N904, N1140);
nor NOR2 (N2072, N2069, N948);
xor XOR2 (N2073, N2061, N1342);
buf BUF1 (N2074, N2070);
or OR2 (N2075, N2043, N861);
and AND3 (N2076, N2073, N600, N562);
not NOT1 (N2077, N2065);
nand NAND2 (N2078, N2067, N32);
buf BUF1 (N2079, N2076);
or OR2 (N2080, N2064, N558);
not NOT1 (N2081, N2080);
or OR2 (N2082, N2075, N1124);
and AND2 (N2083, N2072, N1543);
and AND2 (N2084, N2074, N1921);
not NOT1 (N2085, N2079);
nand NAND3 (N2086, N2083, N798, N588);
xor XOR2 (N2087, N2086, N656);
not NOT1 (N2088, N2081);
or OR3 (N2089, N2068, N1553, N556);
not NOT1 (N2090, N2082);
buf BUF1 (N2091, N2085);
nor NOR2 (N2092, N2089, N161);
and AND4 (N2093, N2090, N656, N117, N1388);
buf BUF1 (N2094, N2092);
xor XOR2 (N2095, N2093, N1513);
nand NAND4 (N2096, N2088, N275, N316, N2058);
or OR3 (N2097, N2071, N675, N496);
and AND4 (N2098, N2094, N2050, N493, N1019);
nor NOR2 (N2099, N2084, N1500);
nor NOR2 (N2100, N2097, N513);
nand NAND2 (N2101, N2077, N830);
nand NAND4 (N2102, N2091, N69, N380, N1236);
buf BUF1 (N2103, N2098);
nand NAND4 (N2104, N2095, N1798, N1291, N1663);
or OR2 (N2105, N2078, N763);
and AND2 (N2106, N2101, N794);
buf BUF1 (N2107, N2099);
or OR4 (N2108, N2103, N1044, N1709, N965);
and AND2 (N2109, N2107, N555);
not NOT1 (N2110, N2087);
or OR3 (N2111, N2106, N541, N14);
not NOT1 (N2112, N2102);
xor XOR2 (N2113, N2112, N1383);
nor NOR4 (N2114, N2110, N1405, N318, N595);
not NOT1 (N2115, N2111);
xor XOR2 (N2116, N2109, N1105);
nand NAND3 (N2117, N2114, N1893, N1559);
buf BUF1 (N2118, N2117);
buf BUF1 (N2119, N2116);
buf BUF1 (N2120, N2115);
buf BUF1 (N2121, N2108);
and AND2 (N2122, N2120, N407);
xor XOR2 (N2123, N2105, N827);
or OR3 (N2124, N2123, N301, N1769);
buf BUF1 (N2125, N2118);
buf BUF1 (N2126, N2096);
not NOT1 (N2127, N2113);
xor XOR2 (N2128, N2124, N1299);
nor NOR2 (N2129, N2121, N394);
or OR4 (N2130, N2127, N168, N1582, N2117);
nor NOR2 (N2131, N2119, N2095);
nand NAND2 (N2132, N2040, N869);
buf BUF1 (N2133, N2125);
buf BUF1 (N2134, N2128);
nand NAND2 (N2135, N2131, N410);
or OR2 (N2136, N2129, N1857);
buf BUF1 (N2137, N2132);
nand NAND2 (N2138, N2104, N1285);
nand NAND3 (N2139, N2133, N1033, N1730);
xor XOR2 (N2140, N2126, N2106);
nor NOR2 (N2141, N2134, N61);
nor NOR2 (N2142, N2136, N942);
and AND2 (N2143, N2130, N1970);
and AND3 (N2144, N2100, N1326, N983);
buf BUF1 (N2145, N2122);
or OR3 (N2146, N2145, N2118, N56);
nand NAND3 (N2147, N2143, N2145, N1068);
xor XOR2 (N2148, N2146, N16);
not NOT1 (N2149, N2147);
and AND3 (N2150, N2148, N797, N760);
nor NOR2 (N2151, N2142, N1468);
or OR2 (N2152, N2137, N2033);
or OR4 (N2153, N2139, N65, N1158, N1760);
or OR3 (N2154, N2138, N963, N1591);
nand NAND2 (N2155, N2151, N804);
buf BUF1 (N2156, N2135);
not NOT1 (N2157, N2156);
or OR2 (N2158, N2141, N1321);
buf BUF1 (N2159, N2157);
buf BUF1 (N2160, N2150);
buf BUF1 (N2161, N2140);
not NOT1 (N2162, N2152);
and AND3 (N2163, N2159, N1494, N482);
xor XOR2 (N2164, N2161, N1428);
xor XOR2 (N2165, N2153, N1077);
nor NOR3 (N2166, N2155, N128, N1797);
and AND4 (N2167, N2164, N925, N860, N1443);
nand NAND2 (N2168, N2166, N818);
buf BUF1 (N2169, N2149);
buf BUF1 (N2170, N2160);
buf BUF1 (N2171, N2169);
or OR3 (N2172, N2170, N907, N585);
xor XOR2 (N2173, N2154, N2033);
nand NAND4 (N2174, N2171, N2130, N1350, N1451);
nand NAND4 (N2175, N2173, N169, N598, N2167);
and AND3 (N2176, N1401, N125, N519);
and AND2 (N2177, N2174, N1463);
nor NOR3 (N2178, N2163, N210, N594);
buf BUF1 (N2179, N2158);
buf BUF1 (N2180, N2179);
or OR4 (N2181, N2144, N1165, N1864, N1141);
nand NAND3 (N2182, N2181, N106, N1436);
or OR4 (N2183, N2175, N2021, N1941, N1826);
buf BUF1 (N2184, N2162);
xor XOR2 (N2185, N2183, N27);
xor XOR2 (N2186, N2172, N1575);
nor NOR2 (N2187, N2168, N462);
xor XOR2 (N2188, N2186, N1593);
nor NOR3 (N2189, N2182, N219, N449);
nand NAND3 (N2190, N2187, N43, N337);
or OR4 (N2191, N2184, N1238, N219, N1110);
or OR4 (N2192, N2188, N68, N2167, N860);
nand NAND4 (N2193, N2185, N1093, N510, N1684);
nor NOR3 (N2194, N2190, N142, N1819);
and AND3 (N2195, N2189, N1144, N2169);
nand NAND3 (N2196, N2193, N1362, N971);
buf BUF1 (N2197, N2195);
buf BUF1 (N2198, N2177);
nand NAND3 (N2199, N2178, N2095, N1093);
xor XOR2 (N2200, N2194, N1226);
not NOT1 (N2201, N2191);
not NOT1 (N2202, N2165);
nor NOR4 (N2203, N2202, N1783, N1941, N1054);
xor XOR2 (N2204, N2180, N190);
nand NAND2 (N2205, N2204, N1514);
nand NAND4 (N2206, N2198, N2001, N869, N485);
not NOT1 (N2207, N2197);
not NOT1 (N2208, N2203);
xor XOR2 (N2209, N2206, N944);
or OR2 (N2210, N2209, N1291);
xor XOR2 (N2211, N2196, N1681);
and AND3 (N2212, N2192, N1509, N966);
nor NOR2 (N2213, N2205, N1878);
nor NOR4 (N2214, N2199, N890, N708, N2203);
or OR3 (N2215, N2200, N81, N156);
buf BUF1 (N2216, N2210);
nand NAND3 (N2217, N2201, N468, N1888);
and AND3 (N2218, N2208, N15, N1451);
nand NAND3 (N2219, N2214, N1832, N63);
nor NOR3 (N2220, N2219, N717, N1158);
buf BUF1 (N2221, N2176);
nor NOR2 (N2222, N2216, N1271);
xor XOR2 (N2223, N2221, N1154);
and AND2 (N2224, N2223, N2139);
buf BUF1 (N2225, N2224);
nor NOR2 (N2226, N2211, N345);
nand NAND3 (N2227, N2226, N2082, N1636);
nand NAND4 (N2228, N2225, N478, N965, N557);
and AND2 (N2229, N2218, N1967);
nor NOR4 (N2230, N2222, N1802, N1987, N1377);
and AND4 (N2231, N2207, N943, N1529, N2217);
nand NAND3 (N2232, N949, N1900, N1658);
not NOT1 (N2233, N2212);
or OR2 (N2234, N2228, N1294);
nand NAND4 (N2235, N2234, N509, N1132, N1702);
xor XOR2 (N2236, N2235, N168);
nor NOR2 (N2237, N2236, N699);
not NOT1 (N2238, N2227);
buf BUF1 (N2239, N2230);
buf BUF1 (N2240, N2220);
nand NAND4 (N2241, N2239, N1936, N1415, N564);
not NOT1 (N2242, N2231);
and AND3 (N2243, N2242, N2015, N2086);
and AND2 (N2244, N2237, N309);
xor XOR2 (N2245, N2244, N863);
buf BUF1 (N2246, N2238);
not NOT1 (N2247, N2240);
buf BUF1 (N2248, N2213);
buf BUF1 (N2249, N2248);
or OR3 (N2250, N2233, N284, N1011);
buf BUF1 (N2251, N2247);
xor XOR2 (N2252, N2249, N1292);
or OR4 (N2253, N2250, N1240, N62, N173);
not NOT1 (N2254, N2251);
and AND3 (N2255, N2245, N514, N1216);
nand NAND3 (N2256, N2229, N1918, N485);
and AND2 (N2257, N2232, N581);
xor XOR2 (N2258, N2255, N1389);
nor NOR4 (N2259, N2246, N1201, N1295, N599);
or OR4 (N2260, N2254, N982, N263, N1138);
buf BUF1 (N2261, N2253);
nand NAND3 (N2262, N2243, N201, N402);
buf BUF1 (N2263, N2260);
not NOT1 (N2264, N2252);
buf BUF1 (N2265, N2259);
not NOT1 (N2266, N2241);
and AND2 (N2267, N2261, N515);
and AND4 (N2268, N2257, N1412, N58, N1335);
nor NOR2 (N2269, N2265, N1740);
nor NOR3 (N2270, N2256, N2056, N859);
nor NOR3 (N2271, N2267, N902, N601);
nand NAND2 (N2272, N2215, N315);
nand NAND3 (N2273, N2270, N1576, N1897);
not NOT1 (N2274, N2269);
nand NAND3 (N2275, N2266, N1451, N782);
not NOT1 (N2276, N2274);
and AND3 (N2277, N2276, N1599, N908);
buf BUF1 (N2278, N2258);
xor XOR2 (N2279, N2278, N141);
nand NAND2 (N2280, N2277, N1608);
nand NAND3 (N2281, N2268, N769, N388);
buf BUF1 (N2282, N2264);
and AND2 (N2283, N2273, N1936);
or OR4 (N2284, N2279, N976, N1556, N197);
nand NAND3 (N2285, N2263, N2079, N475);
xor XOR2 (N2286, N2285, N225);
nand NAND3 (N2287, N2262, N1727, N824);
and AND2 (N2288, N2286, N1868);
buf BUF1 (N2289, N2275);
and AND4 (N2290, N2283, N1130, N1575, N464);
nor NOR2 (N2291, N2284, N3);
nand NAND4 (N2292, N2282, N1316, N1700, N1609);
not NOT1 (N2293, N2287);
nand NAND2 (N2294, N2291, N2256);
and AND2 (N2295, N2288, N1488);
xor XOR2 (N2296, N2295, N1230);
nand NAND2 (N2297, N2271, N694);
nand NAND2 (N2298, N2290, N1254);
or OR4 (N2299, N2294, N1599, N1596, N195);
and AND3 (N2300, N2299, N1798, N890);
nor NOR3 (N2301, N2292, N794, N846);
xor XOR2 (N2302, N2297, N1746);
and AND3 (N2303, N2301, N123, N1042);
xor XOR2 (N2304, N2302, N1658);
or OR2 (N2305, N2280, N813);
not NOT1 (N2306, N2296);
nand NAND4 (N2307, N2304, N1381, N567, N1688);
xor XOR2 (N2308, N2300, N1024);
nor NOR3 (N2309, N2306, N1944, N1371);
nor NOR2 (N2310, N2309, N620);
nor NOR4 (N2311, N2293, N755, N2181, N114);
nor NOR2 (N2312, N2303, N1094);
nand NAND3 (N2313, N2289, N1344, N701);
buf BUF1 (N2314, N2307);
not NOT1 (N2315, N2272);
not NOT1 (N2316, N2312);
nor NOR4 (N2317, N2310, N348, N2005, N95);
nand NAND2 (N2318, N2305, N322);
not NOT1 (N2319, N2318);
and AND2 (N2320, N2319, N911);
or OR4 (N2321, N2315, N2102, N1875, N1134);
xor XOR2 (N2322, N2314, N446);
and AND4 (N2323, N2308, N389, N2235, N1107);
xor XOR2 (N2324, N2298, N2007);
not NOT1 (N2325, N2323);
nand NAND2 (N2326, N2317, N1943);
and AND3 (N2327, N2316, N2179, N324);
and AND2 (N2328, N2321, N153);
nor NOR4 (N2329, N2326, N2004, N1536, N1215);
not NOT1 (N2330, N2313);
xor XOR2 (N2331, N2322, N266);
nor NOR3 (N2332, N2328, N2190, N1716);
or OR3 (N2333, N2320, N1974, N1318);
nor NOR4 (N2334, N2329, N1397, N991, N1055);
nand NAND2 (N2335, N2333, N703);
not NOT1 (N2336, N2324);
and AND2 (N2337, N2327, N1894);
nand NAND3 (N2338, N2325, N93, N440);
nor NOR4 (N2339, N2335, N700, N1433, N1772);
nand NAND2 (N2340, N2338, N764);
or OR2 (N2341, N2331, N130);
and AND2 (N2342, N2281, N1026);
nor NOR4 (N2343, N2341, N239, N233, N652);
nand NAND4 (N2344, N2334, N832, N810, N1940);
xor XOR2 (N2345, N2337, N599);
and AND2 (N2346, N2330, N57);
or OR2 (N2347, N2332, N2303);
buf BUF1 (N2348, N2342);
buf BUF1 (N2349, N2344);
not NOT1 (N2350, N2336);
nor NOR3 (N2351, N2346, N1310, N460);
xor XOR2 (N2352, N2351, N450);
xor XOR2 (N2353, N2348, N1107);
nand NAND4 (N2354, N2352, N1363, N1102, N1363);
or OR4 (N2355, N2345, N452, N831, N1862);
xor XOR2 (N2356, N2340, N2320);
and AND4 (N2357, N2343, N1981, N2101, N1557);
nand NAND4 (N2358, N2347, N298, N1203, N470);
nand NAND2 (N2359, N2339, N1713);
buf BUF1 (N2360, N2358);
or OR2 (N2361, N2356, N1787);
buf BUF1 (N2362, N2361);
xor XOR2 (N2363, N2353, N1128);
or OR3 (N2364, N2362, N1724, N1915);
xor XOR2 (N2365, N2363, N2331);
and AND3 (N2366, N2355, N611, N1868);
not NOT1 (N2367, N2366);
xor XOR2 (N2368, N2350, N2281);
buf BUF1 (N2369, N2311);
not NOT1 (N2370, N2365);
or OR3 (N2371, N2357, N808, N495);
not NOT1 (N2372, N2364);
buf BUF1 (N2373, N2360);
not NOT1 (N2374, N2371);
and AND4 (N2375, N2369, N1808, N1080, N2138);
nor NOR2 (N2376, N2372, N518);
not NOT1 (N2377, N2354);
nor NOR4 (N2378, N2377, N813, N1335, N542);
nand NAND4 (N2379, N2374, N2240, N1898, N994);
nand NAND4 (N2380, N2368, N885, N303, N101);
buf BUF1 (N2381, N2349);
and AND2 (N2382, N2378, N1440);
buf BUF1 (N2383, N2379);
or OR2 (N2384, N2376, N1040);
nand NAND3 (N2385, N2381, N2221, N1173);
not NOT1 (N2386, N2385);
not NOT1 (N2387, N2373);
buf BUF1 (N2388, N2384);
xor XOR2 (N2389, N2367, N346);
buf BUF1 (N2390, N2387);
or OR3 (N2391, N2389, N1810, N128);
nor NOR4 (N2392, N2380, N17, N623, N2338);
xor XOR2 (N2393, N2359, N31);
not NOT1 (N2394, N2375);
not NOT1 (N2395, N2393);
nand NAND2 (N2396, N2388, N1191);
or OR4 (N2397, N2386, N1906, N1366, N1473);
nor NOR2 (N2398, N2383, N1046);
not NOT1 (N2399, N2382);
not NOT1 (N2400, N2391);
or OR3 (N2401, N2399, N1980, N1928);
not NOT1 (N2402, N2395);
not NOT1 (N2403, N2394);
xor XOR2 (N2404, N2370, N1666);
not NOT1 (N2405, N2403);
xor XOR2 (N2406, N2405, N771);
and AND4 (N2407, N2398, N894, N1500, N773);
or OR3 (N2408, N2404, N760, N655);
nor NOR4 (N2409, N2400, N827, N1059, N196);
or OR3 (N2410, N2401, N813, N1434);
buf BUF1 (N2411, N2392);
or OR4 (N2412, N2407, N63, N2024, N1885);
nor NOR2 (N2413, N2397, N504);
nor NOR4 (N2414, N2406, N2110, N1376, N1867);
nor NOR3 (N2415, N2413, N2119, N1717);
not NOT1 (N2416, N2408);
nand NAND2 (N2417, N2410, N1326);
buf BUF1 (N2418, N2417);
and AND4 (N2419, N2414, N506, N2260, N1346);
buf BUF1 (N2420, N2409);
not NOT1 (N2421, N2416);
nor NOR4 (N2422, N2412, N277, N2048, N2115);
nand NAND4 (N2423, N2421, N2083, N1022, N702);
not NOT1 (N2424, N2402);
xor XOR2 (N2425, N2424, N1821);
buf BUF1 (N2426, N2396);
not NOT1 (N2427, N2423);
nor NOR3 (N2428, N2420, N36, N1335);
nor NOR2 (N2429, N2415, N1579);
nand NAND2 (N2430, N2411, N555);
not NOT1 (N2431, N2422);
nor NOR3 (N2432, N2431, N1534, N847);
xor XOR2 (N2433, N2428, N1283);
not NOT1 (N2434, N2429);
not NOT1 (N2435, N2433);
and AND4 (N2436, N2418, N784, N1971, N169);
or OR2 (N2437, N2434, N247);
buf BUF1 (N2438, N2390);
nand NAND2 (N2439, N2438, N136);
or OR3 (N2440, N2419, N1015, N116);
xor XOR2 (N2441, N2432, N157);
nand NAND3 (N2442, N2440, N1029, N385);
or OR4 (N2443, N2427, N1041, N978, N280);
buf BUF1 (N2444, N2442);
not NOT1 (N2445, N2437);
and AND2 (N2446, N2444, N954);
nor NOR3 (N2447, N2446, N737, N237);
buf BUF1 (N2448, N2426);
or OR4 (N2449, N2436, N220, N1576, N260);
nand NAND4 (N2450, N2430, N4, N686, N2396);
nand NAND3 (N2451, N2449, N87, N1294);
and AND2 (N2452, N2450, N579);
xor XOR2 (N2453, N2447, N1254);
or OR2 (N2454, N2435, N830);
nand NAND3 (N2455, N2425, N306, N1529);
and AND2 (N2456, N2441, N2123);
nor NOR2 (N2457, N2454, N25);
not NOT1 (N2458, N2457);
or OR3 (N2459, N2452, N192, N1895);
and AND3 (N2460, N2451, N986, N2001);
xor XOR2 (N2461, N2443, N2404);
buf BUF1 (N2462, N2456);
buf BUF1 (N2463, N2455);
nand NAND3 (N2464, N2463, N22, N585);
buf BUF1 (N2465, N2462);
not NOT1 (N2466, N2464);
xor XOR2 (N2467, N2466, N602);
nor NOR2 (N2468, N2453, N933);
xor XOR2 (N2469, N2468, N662);
buf BUF1 (N2470, N2460);
buf BUF1 (N2471, N2448);
nor NOR3 (N2472, N2467, N404, N244);
nand NAND3 (N2473, N2445, N76, N1234);
or OR3 (N2474, N2458, N1208, N757);
nor NOR4 (N2475, N2469, N508, N1549, N834);
buf BUF1 (N2476, N2471);
and AND3 (N2477, N2475, N2276, N731);
nor NOR2 (N2478, N2476, N630);
or OR4 (N2479, N2473, N1970, N1014, N393);
buf BUF1 (N2480, N2472);
not NOT1 (N2481, N2478);
nor NOR4 (N2482, N2470, N1696, N94, N2380);
buf BUF1 (N2483, N2465);
nor NOR3 (N2484, N2459, N1302, N365);
nand NAND4 (N2485, N2483, N1353, N1358, N1752);
nor NOR3 (N2486, N2477, N299, N1855);
xor XOR2 (N2487, N2474, N2466);
not NOT1 (N2488, N2480);
xor XOR2 (N2489, N2481, N1637);
buf BUF1 (N2490, N2485);
nor NOR4 (N2491, N2484, N1205, N2209, N643);
xor XOR2 (N2492, N2488, N429);
xor XOR2 (N2493, N2461, N1360);
buf BUF1 (N2494, N2490);
and AND4 (N2495, N2482, N1113, N399, N1362);
buf BUF1 (N2496, N2489);
xor XOR2 (N2497, N2496, N1245);
and AND3 (N2498, N2491, N2335, N923);
nand NAND3 (N2499, N2479, N222, N608);
not NOT1 (N2500, N2495);
not NOT1 (N2501, N2493);
not NOT1 (N2502, N2486);
or OR3 (N2503, N2497, N2370, N1553);
nand NAND3 (N2504, N2487, N1248, N897);
or OR2 (N2505, N2439, N955);
nor NOR4 (N2506, N2504, N1061, N2251, N334);
xor XOR2 (N2507, N2500, N1075);
not NOT1 (N2508, N2507);
or OR2 (N2509, N2501, N2266);
nand NAND4 (N2510, N2505, N484, N1436, N204);
not NOT1 (N2511, N2509);
nor NOR2 (N2512, N2502, N731);
or OR2 (N2513, N2503, N728);
nand NAND4 (N2514, N2499, N1383, N1324, N271);
or OR4 (N2515, N2506, N2451, N1295, N1291);
xor XOR2 (N2516, N2498, N354);
xor XOR2 (N2517, N2512, N2127);
nand NAND2 (N2518, N2517, N783);
or OR3 (N2519, N2508, N709, N393);
buf BUF1 (N2520, N2494);
or OR3 (N2521, N2520, N683, N25);
not NOT1 (N2522, N2519);
not NOT1 (N2523, N2516);
xor XOR2 (N2524, N2492, N1963);
buf BUF1 (N2525, N2510);
or OR2 (N2526, N2515, N1171);
nand NAND2 (N2527, N2513, N913);
xor XOR2 (N2528, N2526, N712);
nand NAND2 (N2529, N2528, N2482);
xor XOR2 (N2530, N2523, N925);
nand NAND3 (N2531, N2527, N1677, N2357);
buf BUF1 (N2532, N2530);
or OR3 (N2533, N2524, N1619, N2206);
and AND2 (N2534, N2514, N1596);
not NOT1 (N2535, N2511);
nor NOR2 (N2536, N2533, N667);
or OR3 (N2537, N2534, N18, N812);
xor XOR2 (N2538, N2522, N320);
not NOT1 (N2539, N2537);
and AND2 (N2540, N2532, N139);
buf BUF1 (N2541, N2536);
or OR4 (N2542, N2541, N95, N2103, N757);
xor XOR2 (N2543, N2540, N1300);
xor XOR2 (N2544, N2538, N719);
or OR3 (N2545, N2529, N1679, N1751);
buf BUF1 (N2546, N2535);
or OR3 (N2547, N2531, N1009, N1159);
buf BUF1 (N2548, N2545);
xor XOR2 (N2549, N2542, N979);
nor NOR4 (N2550, N2544, N1333, N2414, N254);
xor XOR2 (N2551, N2548, N761);
buf BUF1 (N2552, N2551);
xor XOR2 (N2553, N2539, N780);
buf BUF1 (N2554, N2547);
xor XOR2 (N2555, N2550, N76);
or OR2 (N2556, N2543, N2022);
xor XOR2 (N2557, N2518, N582);
xor XOR2 (N2558, N2555, N2480);
xor XOR2 (N2559, N2556, N2369);
not NOT1 (N2560, N2554);
and AND4 (N2561, N2560, N804, N1216, N1860);
nand NAND4 (N2562, N2559, N2436, N764, N1021);
and AND3 (N2563, N2561, N1905, N2549);
or OR4 (N2564, N2139, N2540, N2326, N44);
buf BUF1 (N2565, N2525);
nor NOR4 (N2566, N2565, N2294, N1605, N1995);
or OR4 (N2567, N2557, N1968, N293, N530);
nand NAND4 (N2568, N2567, N2395, N1251, N557);
xor XOR2 (N2569, N2552, N746);
not NOT1 (N2570, N2521);
xor XOR2 (N2571, N2558, N1346);
buf BUF1 (N2572, N2563);
nand NAND4 (N2573, N2568, N2491, N1205, N1824);
not NOT1 (N2574, N2564);
xor XOR2 (N2575, N2573, N163);
xor XOR2 (N2576, N2562, N1371);
nand NAND4 (N2577, N2569, N241, N561, N408);
nor NOR4 (N2578, N2575, N436, N565, N1463);
and AND4 (N2579, N2578, N44, N995, N946);
not NOT1 (N2580, N2546);
xor XOR2 (N2581, N2574, N1815);
xor XOR2 (N2582, N2579, N2366);
buf BUF1 (N2583, N2572);
xor XOR2 (N2584, N2583, N166);
nand NAND4 (N2585, N2576, N1808, N1321, N1919);
or OR3 (N2586, N2581, N1240, N1352);
and AND3 (N2587, N2585, N705, N1790);
not NOT1 (N2588, N2580);
or OR3 (N2589, N2571, N1316, N332);
not NOT1 (N2590, N2588);
not NOT1 (N2591, N2566);
nand NAND3 (N2592, N2553, N402, N2502);
and AND2 (N2593, N2570, N757);
and AND4 (N2594, N2590, N809, N457, N1283);
nor NOR3 (N2595, N2592, N120, N1731);
xor XOR2 (N2596, N2577, N2114);
buf BUF1 (N2597, N2582);
xor XOR2 (N2598, N2593, N754);
nor NOR3 (N2599, N2595, N626, N1221);
not NOT1 (N2600, N2598);
nand NAND2 (N2601, N2591, N2295);
or OR3 (N2602, N2597, N698, N310);
and AND4 (N2603, N2586, N2483, N2274, N2096);
or OR4 (N2604, N2600, N2293, N1728, N2391);
not NOT1 (N2605, N2602);
and AND4 (N2606, N2601, N985, N1539, N1300);
nand NAND3 (N2607, N2599, N1219, N190);
or OR2 (N2608, N2607, N1272);
nand NAND4 (N2609, N2594, N2527, N2408, N2567);
nor NOR2 (N2610, N2605, N2373);
xor XOR2 (N2611, N2610, N813);
nand NAND4 (N2612, N2589, N1059, N2503, N2201);
nand NAND3 (N2613, N2603, N1919, N617);
or OR2 (N2614, N2612, N151);
nand NAND3 (N2615, N2606, N765, N84);
and AND3 (N2616, N2615, N541, N598);
buf BUF1 (N2617, N2596);
nor NOR3 (N2618, N2617, N202, N1292);
and AND2 (N2619, N2584, N412);
xor XOR2 (N2620, N2616, N2133);
and AND4 (N2621, N2608, N1302, N1991, N1028);
xor XOR2 (N2622, N2620, N2436);
not NOT1 (N2623, N2618);
nor NOR4 (N2624, N2619, N1384, N646, N1448);
or OR3 (N2625, N2587, N1448, N2520);
nor NOR4 (N2626, N2622, N1028, N77, N377);
xor XOR2 (N2627, N2621, N1602);
nor NOR4 (N2628, N2627, N1562, N486, N2241);
not NOT1 (N2629, N2614);
nor NOR4 (N2630, N2628, N1864, N1806, N788);
xor XOR2 (N2631, N2625, N857);
xor XOR2 (N2632, N2630, N888);
nand NAND4 (N2633, N2632, N1678, N1989, N2290);
nand NAND3 (N2634, N2613, N106, N1552);
or OR2 (N2635, N2633, N718);
or OR2 (N2636, N2631, N2022);
not NOT1 (N2637, N2611);
or OR3 (N2638, N2635, N1828, N1970);
buf BUF1 (N2639, N2604);
and AND4 (N2640, N2609, N1939, N1526, N2244);
nand NAND3 (N2641, N2626, N2631, N1660);
buf BUF1 (N2642, N2640);
not NOT1 (N2643, N2623);
nand NAND4 (N2644, N2636, N203, N1040, N1249);
and AND2 (N2645, N2643, N2370);
xor XOR2 (N2646, N2624, N1931);
nand NAND4 (N2647, N2645, N2524, N1594, N238);
nor NOR3 (N2648, N2629, N1629, N631);
nor NOR4 (N2649, N2647, N536, N532, N2576);
not NOT1 (N2650, N2644);
buf BUF1 (N2651, N2649);
buf BUF1 (N2652, N2634);
nand NAND4 (N2653, N2651, N2287, N1188, N1188);
not NOT1 (N2654, N2641);
nor NOR2 (N2655, N2646, N1473);
xor XOR2 (N2656, N2642, N436);
nand NAND2 (N2657, N2637, N45);
xor XOR2 (N2658, N2650, N2369);
nand NAND3 (N2659, N2652, N233, N2367);
xor XOR2 (N2660, N2654, N12);
or OR4 (N2661, N2639, N2441, N1025, N1195);
buf BUF1 (N2662, N2658);
and AND2 (N2663, N2638, N84);
buf BUF1 (N2664, N2660);
nand NAND2 (N2665, N2662, N1185);
not NOT1 (N2666, N2663);
buf BUF1 (N2667, N2653);
or OR4 (N2668, N2656, N2392, N2064, N315);
and AND4 (N2669, N2667, N2661, N1008, N2549);
xor XOR2 (N2670, N1947, N155);
and AND3 (N2671, N2669, N1584, N1249);
not NOT1 (N2672, N2659);
nor NOR3 (N2673, N2666, N1762, N897);
and AND4 (N2674, N2664, N2387, N818, N806);
and AND2 (N2675, N2648, N787);
xor XOR2 (N2676, N2665, N548);
nand NAND2 (N2677, N2674, N2414);
xor XOR2 (N2678, N2670, N1280);
and AND3 (N2679, N2672, N1832, N27);
nand NAND2 (N2680, N2679, N398);
buf BUF1 (N2681, N2677);
xor XOR2 (N2682, N2655, N1521);
buf BUF1 (N2683, N2675);
not NOT1 (N2684, N2683);
nand NAND2 (N2685, N2680, N1791);
or OR2 (N2686, N2685, N1988);
not NOT1 (N2687, N2671);
and AND3 (N2688, N2673, N1937, N598);
or OR3 (N2689, N2682, N1940, N188);
not NOT1 (N2690, N2684);
nand NAND2 (N2691, N2678, N1396);
nand NAND2 (N2692, N2676, N2021);
and AND3 (N2693, N2689, N1734, N1118);
and AND3 (N2694, N2657, N298, N1776);
not NOT1 (N2695, N2681);
nor NOR4 (N2696, N2690, N1134, N2304, N1735);
buf BUF1 (N2697, N2695);
buf BUF1 (N2698, N2686);
or OR3 (N2699, N2692, N550, N949);
and AND3 (N2700, N2698, N1688, N2188);
not NOT1 (N2701, N2693);
and AND2 (N2702, N2697, N2692);
nor NOR4 (N2703, N2668, N904, N1188, N2434);
buf BUF1 (N2704, N2699);
and AND2 (N2705, N2691, N2030);
nor NOR3 (N2706, N2705, N163, N1501);
and AND3 (N2707, N2702, N369, N1770);
xor XOR2 (N2708, N2701, N638);
xor XOR2 (N2709, N2708, N1485);
xor XOR2 (N2710, N2688, N2430);
xor XOR2 (N2711, N2703, N1112);
nor NOR3 (N2712, N2707, N2514, N1788);
or OR4 (N2713, N2709, N73, N1094, N2390);
buf BUF1 (N2714, N2694);
xor XOR2 (N2715, N2696, N102);
not NOT1 (N2716, N2715);
and AND3 (N2717, N2704, N1064, N206);
xor XOR2 (N2718, N2717, N2595);
and AND2 (N2719, N2714, N379);
nor NOR3 (N2720, N2687, N1080, N58);
not NOT1 (N2721, N2706);
xor XOR2 (N2722, N2713, N1755);
xor XOR2 (N2723, N2710, N397);
buf BUF1 (N2724, N2712);
buf BUF1 (N2725, N2700);
not NOT1 (N2726, N2723);
or OR4 (N2727, N2722, N1680, N551, N2642);
and AND4 (N2728, N2726, N2532, N529, N1703);
xor XOR2 (N2729, N2718, N503);
and AND4 (N2730, N2724, N2186, N1186, N161);
and AND4 (N2731, N2728, N347, N910, N822);
and AND3 (N2732, N2729, N1158, N1691);
xor XOR2 (N2733, N2725, N915);
nor NOR3 (N2734, N2720, N547, N708);
buf BUF1 (N2735, N2733);
nor NOR2 (N2736, N2731, N1344);
nand NAND2 (N2737, N2711, N2364);
or OR2 (N2738, N2727, N2075);
buf BUF1 (N2739, N2732);
or OR4 (N2740, N2736, N1455, N1876, N648);
or OR4 (N2741, N2719, N1126, N2670, N1959);
xor XOR2 (N2742, N2735, N1091);
not NOT1 (N2743, N2742);
nor NOR2 (N2744, N2730, N92);
and AND4 (N2745, N2741, N1153, N2388, N995);
or OR2 (N2746, N2737, N646);
not NOT1 (N2747, N2721);
nor NOR2 (N2748, N2716, N1504);
nor NOR4 (N2749, N2743, N1031, N696, N962);
nor NOR4 (N2750, N2745, N2744, N48, N2339);
not NOT1 (N2751, N2148);
or OR2 (N2752, N2740, N1670);
buf BUF1 (N2753, N2750);
buf BUF1 (N2754, N2739);
and AND4 (N2755, N2748, N1433, N911, N2689);
xor XOR2 (N2756, N2738, N1757);
buf BUF1 (N2757, N2755);
nor NOR4 (N2758, N2734, N674, N2440, N650);
xor XOR2 (N2759, N2749, N1876);
buf BUF1 (N2760, N2746);
buf BUF1 (N2761, N2756);
nand NAND3 (N2762, N2753, N2418, N1974);
xor XOR2 (N2763, N2747, N1875);
and AND3 (N2764, N2762, N316, N2160);
or OR2 (N2765, N2760, N351);
nor NOR2 (N2766, N2754, N2579);
not NOT1 (N2767, N2752);
xor XOR2 (N2768, N2766, N975);
not NOT1 (N2769, N2759);
nor NOR3 (N2770, N2763, N1977, N2340);
not NOT1 (N2771, N2758);
xor XOR2 (N2772, N2761, N2424);
xor XOR2 (N2773, N2765, N962);
and AND4 (N2774, N2773, N70, N2325, N2249);
xor XOR2 (N2775, N2772, N892);
xor XOR2 (N2776, N2774, N714);
buf BUF1 (N2777, N2771);
or OR4 (N2778, N2764, N240, N2671, N2673);
not NOT1 (N2779, N2751);
buf BUF1 (N2780, N2775);
not NOT1 (N2781, N2780);
not NOT1 (N2782, N2770);
buf BUF1 (N2783, N2769);
or OR4 (N2784, N2783, N1246, N368, N1703);
nand NAND3 (N2785, N2779, N1152, N1782);
nor NOR2 (N2786, N2784, N1298);
xor XOR2 (N2787, N2757, N2085);
nor NOR3 (N2788, N2782, N1820, N625);
xor XOR2 (N2789, N2778, N82);
buf BUF1 (N2790, N2789);
not NOT1 (N2791, N2767);
or OR2 (N2792, N2790, N55);
buf BUF1 (N2793, N2786);
buf BUF1 (N2794, N2793);
xor XOR2 (N2795, N2777, N2254);
buf BUF1 (N2796, N2795);
not NOT1 (N2797, N2791);
nor NOR4 (N2798, N2788, N1167, N2702, N2702);
or OR3 (N2799, N2768, N2684, N1347);
nor NOR4 (N2800, N2799, N1047, N2426, N1294);
nor NOR3 (N2801, N2787, N1538, N308);
xor XOR2 (N2802, N2785, N1803);
buf BUF1 (N2803, N2776);
nor NOR3 (N2804, N2803, N75, N2473);
nor NOR2 (N2805, N2781, N296);
buf BUF1 (N2806, N2792);
not NOT1 (N2807, N2800);
nand NAND2 (N2808, N2798, N2649);
or OR4 (N2809, N2796, N2144, N2543, N688);
not NOT1 (N2810, N2802);
nand NAND3 (N2811, N2805, N2540, N2609);
buf BUF1 (N2812, N2811);
nor NOR4 (N2813, N2809, N2378, N2770, N2019);
nand NAND2 (N2814, N2801, N1214);
buf BUF1 (N2815, N2814);
not NOT1 (N2816, N2812);
buf BUF1 (N2817, N2810);
and AND4 (N2818, N2817, N286, N749, N370);
buf BUF1 (N2819, N2816);
not NOT1 (N2820, N2819);
nor NOR2 (N2821, N2807, N1178);
and AND3 (N2822, N2797, N2515, N2210);
buf BUF1 (N2823, N2804);
xor XOR2 (N2824, N2822, N1049);
or OR4 (N2825, N2806, N2325, N2434, N1064);
nor NOR2 (N2826, N2820, N2478);
and AND4 (N2827, N2815, N326, N1651, N2358);
not NOT1 (N2828, N2808);
not NOT1 (N2829, N2813);
xor XOR2 (N2830, N2818, N1074);
or OR4 (N2831, N2824, N647, N2488, N986);
and AND3 (N2832, N2830, N1488, N2124);
buf BUF1 (N2833, N2826);
xor XOR2 (N2834, N2823, N2390);
and AND3 (N2835, N2831, N716, N646);
buf BUF1 (N2836, N2821);
buf BUF1 (N2837, N2828);
buf BUF1 (N2838, N2834);
xor XOR2 (N2839, N2833, N1621);
or OR3 (N2840, N2839, N655, N2596);
nand NAND2 (N2841, N2794, N2756);
and AND3 (N2842, N2837, N676, N1757);
xor XOR2 (N2843, N2836, N1999);
nor NOR3 (N2844, N2835, N1315, N2071);
or OR3 (N2845, N2829, N503, N1773);
buf BUF1 (N2846, N2845);
not NOT1 (N2847, N2846);
nor NOR4 (N2848, N2827, N2634, N1598, N1277);
nand NAND2 (N2849, N2844, N206);
xor XOR2 (N2850, N2832, N506);
and AND4 (N2851, N2843, N418, N241, N1564);
not NOT1 (N2852, N2847);
or OR2 (N2853, N2848, N992);
nor NOR2 (N2854, N2853, N847);
xor XOR2 (N2855, N2854, N1181);
nor NOR3 (N2856, N2840, N1188, N837);
nor NOR2 (N2857, N2842, N287);
xor XOR2 (N2858, N2857, N996);
and AND2 (N2859, N2851, N864);
and AND3 (N2860, N2849, N2626, N1917);
nor NOR3 (N2861, N2841, N2055, N480);
and AND3 (N2862, N2838, N284, N1796);
nor NOR3 (N2863, N2856, N966, N2410);
buf BUF1 (N2864, N2850);
or OR4 (N2865, N2864, N917, N1611, N1831);
not NOT1 (N2866, N2825);
nand NAND3 (N2867, N2866, N277, N1246);
xor XOR2 (N2868, N2859, N1788);
nor NOR4 (N2869, N2858, N2308, N1154, N2101);
not NOT1 (N2870, N2867);
nor NOR4 (N2871, N2852, N2727, N1267, N483);
or OR2 (N2872, N2861, N2616);
xor XOR2 (N2873, N2860, N1264);
nor NOR2 (N2874, N2855, N1057);
nand NAND3 (N2875, N2862, N2797, N2081);
xor XOR2 (N2876, N2863, N3);
buf BUF1 (N2877, N2873);
and AND4 (N2878, N2874, N2847, N1694, N1001);
or OR2 (N2879, N2876, N2072);
not NOT1 (N2880, N2865);
nand NAND2 (N2881, N2869, N392);
and AND3 (N2882, N2872, N444, N2200);
nor NOR4 (N2883, N2875, N2582, N2840, N1639);
buf BUF1 (N2884, N2868);
xor XOR2 (N2885, N2881, N1263);
and AND4 (N2886, N2870, N712, N1210, N2052);
buf BUF1 (N2887, N2882);
or OR4 (N2888, N2879, N1313, N2525, N1787);
and AND4 (N2889, N2886, N212, N2650, N2148);
or OR3 (N2890, N2871, N1301, N1544);
or OR4 (N2891, N2885, N967, N649, N764);
buf BUF1 (N2892, N2887);
buf BUF1 (N2893, N2884);
buf BUF1 (N2894, N2883);
and AND2 (N2895, N2878, N1789);
not NOT1 (N2896, N2894);
nand NAND3 (N2897, N2891, N2762, N48);
nor NOR3 (N2898, N2893, N542, N2061);
xor XOR2 (N2899, N2897, N1718);
xor XOR2 (N2900, N2895, N2278);
and AND2 (N2901, N2900, N697);
and AND4 (N2902, N2896, N1300, N1052, N1427);
xor XOR2 (N2903, N2902, N1027);
xor XOR2 (N2904, N2889, N2133);
and AND2 (N2905, N2892, N487);
not NOT1 (N2906, N2880);
and AND3 (N2907, N2905, N1530, N2512);
and AND3 (N2908, N2898, N1126, N1576);
nand NAND3 (N2909, N2903, N2100, N785);
xor XOR2 (N2910, N2877, N1446);
and AND3 (N2911, N2901, N128, N340);
nor NOR3 (N2912, N2907, N600, N1163);
nand NAND4 (N2913, N2904, N1510, N1549, N2653);
xor XOR2 (N2914, N2906, N1270);
or OR3 (N2915, N2914, N778, N2379);
nand NAND2 (N2916, N2908, N1068);
and AND3 (N2917, N2913, N2607, N2175);
or OR3 (N2918, N2909, N1542, N1889);
nor NOR4 (N2919, N2918, N2373, N1672, N1540);
or OR2 (N2920, N2919, N597);
nor NOR4 (N2921, N2920, N2428, N905, N527);
nor NOR2 (N2922, N2916, N1655);
buf BUF1 (N2923, N2911);
and AND3 (N2924, N2923, N2457, N851);
nor NOR3 (N2925, N2899, N475, N2451);
xor XOR2 (N2926, N2910, N297);
nand NAND2 (N2927, N2915, N2588);
nor NOR2 (N2928, N2917, N739);
not NOT1 (N2929, N2890);
nor NOR2 (N2930, N2928, N179);
xor XOR2 (N2931, N2925, N287);
nor NOR2 (N2932, N2930, N2218);
buf BUF1 (N2933, N2912);
nor NOR3 (N2934, N2932, N682, N1426);
not NOT1 (N2935, N2931);
and AND2 (N2936, N2924, N406);
buf BUF1 (N2937, N2922);
xor XOR2 (N2938, N2888, N2449);
nand NAND4 (N2939, N2938, N404, N971, N522);
xor XOR2 (N2940, N2926, N1190);
nor NOR2 (N2941, N2929, N906);
buf BUF1 (N2942, N2937);
not NOT1 (N2943, N2939);
or OR4 (N2944, N2935, N1637, N2618, N511);
nor NOR4 (N2945, N2921, N385, N823, N393);
not NOT1 (N2946, N2934);
not NOT1 (N2947, N2944);
and AND2 (N2948, N2941, N1028);
xor XOR2 (N2949, N2947, N1337);
not NOT1 (N2950, N2946);
buf BUF1 (N2951, N2927);
xor XOR2 (N2952, N2951, N2460);
buf BUF1 (N2953, N2952);
or OR4 (N2954, N2949, N1061, N2158, N625);
and AND2 (N2955, N2933, N1134);
nand NAND2 (N2956, N2945, N873);
not NOT1 (N2957, N2950);
or OR2 (N2958, N2954, N1213);
or OR3 (N2959, N2936, N791, N547);
not NOT1 (N2960, N2955);
buf BUF1 (N2961, N2953);
or OR4 (N2962, N2940, N1032, N2015, N1222);
xor XOR2 (N2963, N2948, N418);
buf BUF1 (N2964, N2957);
and AND2 (N2965, N2942, N1535);
xor XOR2 (N2966, N2960, N1389);
xor XOR2 (N2967, N2963, N97);
nand NAND2 (N2968, N2966, N38);
and AND2 (N2969, N2959, N2414);
nor NOR4 (N2970, N2967, N626, N835, N2385);
nor NOR4 (N2971, N2968, N2019, N309, N288);
nor NOR2 (N2972, N2965, N2185);
or OR2 (N2973, N2962, N1257);
not NOT1 (N2974, N2958);
not NOT1 (N2975, N2973);
nor NOR2 (N2976, N2971, N2196);
or OR2 (N2977, N2972, N131);
nand NAND4 (N2978, N2970, N1280, N287, N2867);
xor XOR2 (N2979, N2956, N1066);
nor NOR4 (N2980, N2943, N545, N915, N1361);
nand NAND3 (N2981, N2979, N1423, N1501);
buf BUF1 (N2982, N2975);
not NOT1 (N2983, N2977);
not NOT1 (N2984, N2978);
xor XOR2 (N2985, N2981, N792);
not NOT1 (N2986, N2976);
or OR4 (N2987, N2983, N2902, N1017, N1131);
nor NOR4 (N2988, N2986, N1634, N775, N1392);
buf BUF1 (N2989, N2969);
nand NAND4 (N2990, N2989, N1614, N578, N2169);
and AND3 (N2991, N2985, N801, N2957);
buf BUF1 (N2992, N2984);
and AND2 (N2993, N2988, N535);
and AND4 (N2994, N2982, N2032, N1410, N1522);
nand NAND2 (N2995, N2964, N1879);
buf BUF1 (N2996, N2993);
and AND2 (N2997, N2991, N486);
xor XOR2 (N2998, N2995, N2401);
buf BUF1 (N2999, N2980);
nand NAND3 (N3000, N2997, N2024, N988);
nor NOR2 (N3001, N2987, N2183);
and AND3 (N3002, N3001, N2534, N1447);
xor XOR2 (N3003, N2999, N2866);
xor XOR2 (N3004, N2990, N1558);
nand NAND2 (N3005, N3000, N1862);
or OR4 (N3006, N2974, N1601, N2740, N1926);
and AND4 (N3007, N2998, N2373, N58, N2024);
buf BUF1 (N3008, N3005);
nor NOR4 (N3009, N2992, N146, N2466, N2430);
or OR2 (N3010, N3002, N1169);
not NOT1 (N3011, N2994);
nand NAND4 (N3012, N3003, N1243, N36, N2660);
nand NAND2 (N3013, N3004, N531);
nand NAND4 (N3014, N3007, N1920, N1091, N2374);
nor NOR2 (N3015, N3010, N26);
nand NAND4 (N3016, N3009, N1819, N1739, N1751);
and AND3 (N3017, N3016, N2983, N921);
buf BUF1 (N3018, N3006);
and AND4 (N3019, N3017, N2977, N1702, N1805);
nor NOR4 (N3020, N3019, N2165, N2287, N1370);
nand NAND4 (N3021, N3018, N825, N2332, N405);
not NOT1 (N3022, N3008);
not NOT1 (N3023, N3022);
not NOT1 (N3024, N2961);
nor NOR2 (N3025, N3023, N724);
or OR2 (N3026, N3012, N639);
not NOT1 (N3027, N3021);
nor NOR2 (N3028, N3011, N678);
or OR2 (N3029, N3015, N2795);
nand NAND3 (N3030, N3020, N1304, N2802);
nand NAND2 (N3031, N2996, N460);
buf BUF1 (N3032, N3029);
or OR4 (N3033, N3014, N1226, N2571, N1726);
xor XOR2 (N3034, N3032, N1741);
or OR2 (N3035, N3033, N475);
buf BUF1 (N3036, N3024);
nor NOR2 (N3037, N3026, N404);
and AND3 (N3038, N3035, N2418, N3011);
not NOT1 (N3039, N3037);
not NOT1 (N3040, N3030);
and AND3 (N3041, N3028, N1298, N439);
or OR2 (N3042, N3040, N1129);
or OR2 (N3043, N3027, N253);
and AND4 (N3044, N3042, N2842, N199, N2637);
and AND2 (N3045, N3025, N456);
nor NOR4 (N3046, N3038, N1451, N2450, N427);
and AND3 (N3047, N3044, N401, N1258);
xor XOR2 (N3048, N3041, N981);
buf BUF1 (N3049, N3031);
not NOT1 (N3050, N3043);
xor XOR2 (N3051, N3045, N3018);
buf BUF1 (N3052, N3051);
and AND2 (N3053, N3046, N2065);
not NOT1 (N3054, N3048);
nor NOR4 (N3055, N3049, N1441, N964, N1987);
nor NOR2 (N3056, N3050, N2707);
and AND2 (N3057, N3034, N222);
xor XOR2 (N3058, N3047, N2316);
buf BUF1 (N3059, N3058);
and AND3 (N3060, N3059, N1556, N169);
and AND2 (N3061, N3057, N210);
xor XOR2 (N3062, N3052, N1789);
nand NAND4 (N3063, N3061, N954, N2797, N524);
xor XOR2 (N3064, N3063, N2895);
and AND3 (N3065, N3039, N2391, N1406);
nand NAND4 (N3066, N3060, N77, N1437, N2700);
and AND3 (N3067, N3064, N2454, N718);
xor XOR2 (N3068, N3065, N2681);
nor NOR2 (N3069, N3036, N2056);
nand NAND3 (N3070, N3067, N2743, N986);
not NOT1 (N3071, N3068);
or OR4 (N3072, N3056, N2607, N248, N1900);
buf BUF1 (N3073, N3072);
buf BUF1 (N3074, N3071);
or OR3 (N3075, N3073, N825, N2591);
nor NOR3 (N3076, N3054, N425, N1267);
and AND4 (N3077, N3075, N1087, N977, N2807);
buf BUF1 (N3078, N3055);
or OR4 (N3079, N3077, N2379, N1506, N2796);
nand NAND2 (N3080, N3074, N1393);
and AND3 (N3081, N3076, N377, N2305);
xor XOR2 (N3082, N3079, N1173);
nand NAND3 (N3083, N3078, N789, N2430);
or OR4 (N3084, N3053, N1448, N1666, N2315);
nor NOR2 (N3085, N3083, N2849);
not NOT1 (N3086, N3013);
or OR3 (N3087, N3085, N2195, N2435);
or OR3 (N3088, N3087, N882, N2274);
buf BUF1 (N3089, N3066);
xor XOR2 (N3090, N3081, N2416);
and AND4 (N3091, N3082, N2000, N776, N871);
buf BUF1 (N3092, N3090);
xor XOR2 (N3093, N3069, N1489);
not NOT1 (N3094, N3062);
or OR2 (N3095, N3080, N18);
nand NAND4 (N3096, N3091, N3081, N2812, N341);
nor NOR2 (N3097, N3096, N1823);
not NOT1 (N3098, N3092);
not NOT1 (N3099, N3094);
nor NOR4 (N3100, N3086, N888, N2294, N2193);
nand NAND2 (N3101, N3093, N2191);
or OR4 (N3102, N3089, N1637, N71, N1632);
or OR2 (N3103, N3101, N1359);
xor XOR2 (N3104, N3084, N2371);
nor NOR3 (N3105, N3099, N2439, N1753);
not NOT1 (N3106, N3098);
nand NAND4 (N3107, N3102, N1697, N40, N207);
not NOT1 (N3108, N3103);
not NOT1 (N3109, N3070);
not NOT1 (N3110, N3106);
nand NAND4 (N3111, N3110, N2392, N747, N1695);
xor XOR2 (N3112, N3105, N2154);
nor NOR3 (N3113, N3112, N3085, N2123);
nor NOR3 (N3114, N3104, N2031, N60);
not NOT1 (N3115, N3114);
nand NAND4 (N3116, N3107, N2786, N1507, N2990);
xor XOR2 (N3117, N3100, N112);
not NOT1 (N3118, N3095);
nand NAND4 (N3119, N3118, N1799, N2110, N423);
and AND2 (N3120, N3113, N2648);
buf BUF1 (N3121, N3120);
nand NAND2 (N3122, N3108, N978);
or OR2 (N3123, N3111, N1451);
xor XOR2 (N3124, N3122, N1076);
or OR3 (N3125, N3123, N2001, N811);
buf BUF1 (N3126, N3124);
not NOT1 (N3127, N3126);
nand NAND3 (N3128, N3115, N2597, N402);
or OR3 (N3129, N3116, N1190, N750);
nand NAND3 (N3130, N3117, N33, N667);
buf BUF1 (N3131, N3127);
and AND4 (N3132, N3109, N195, N1067, N437);
xor XOR2 (N3133, N3128, N288);
nand NAND3 (N3134, N3088, N884, N2124);
xor XOR2 (N3135, N3119, N2544);
not NOT1 (N3136, N3129);
or OR3 (N3137, N3125, N474, N1757);
nor NOR4 (N3138, N3134, N942, N1547, N2473);
not NOT1 (N3139, N3121);
buf BUF1 (N3140, N3135);
buf BUF1 (N3141, N3136);
or OR4 (N3142, N3139, N873, N602, N670);
not NOT1 (N3143, N3138);
not NOT1 (N3144, N3141);
nand NAND4 (N3145, N3131, N2546, N2626, N996);
or OR2 (N3146, N3142, N547);
not NOT1 (N3147, N3097);
nand NAND2 (N3148, N3143, N650);
and AND3 (N3149, N3132, N876, N1697);
buf BUF1 (N3150, N3145);
xor XOR2 (N3151, N3130, N1279);
nor NOR3 (N3152, N3137, N2511, N1015);
buf BUF1 (N3153, N3144);
or OR4 (N3154, N3146, N2127, N1909, N1821);
or OR3 (N3155, N3151, N3122, N1442);
xor XOR2 (N3156, N3133, N916);
not NOT1 (N3157, N3148);
and AND3 (N3158, N3150, N84, N801);
or OR3 (N3159, N3158, N2058, N63);
nand NAND3 (N3160, N3153, N1998, N3048);
xor XOR2 (N3161, N3154, N2507);
not NOT1 (N3162, N3155);
and AND2 (N3163, N3157, N2971);
and AND3 (N3164, N3152, N1237, N803);
buf BUF1 (N3165, N3162);
nor NOR3 (N3166, N3160, N952, N437);
or OR3 (N3167, N3161, N622, N47);
or OR4 (N3168, N3164, N1509, N1186, N449);
nand NAND4 (N3169, N3147, N449, N1288, N766);
nor NOR2 (N3170, N3166, N2186);
xor XOR2 (N3171, N3159, N579);
nand NAND2 (N3172, N3168, N910);
nor NOR2 (N3173, N3169, N978);
and AND3 (N3174, N3170, N3146, N144);
nand NAND3 (N3175, N3172, N37, N1171);
xor XOR2 (N3176, N3156, N1733);
and AND4 (N3177, N3167, N1426, N2932, N1522);
buf BUF1 (N3178, N3173);
xor XOR2 (N3179, N3176, N509);
not NOT1 (N3180, N3179);
nand NAND4 (N3181, N3165, N2218, N1734, N1012);
xor XOR2 (N3182, N3171, N1858);
nor NOR2 (N3183, N3180, N2350);
nor NOR4 (N3184, N3178, N262, N904, N262);
nor NOR3 (N3185, N3182, N546, N2413);
and AND4 (N3186, N3183, N263, N3010, N168);
not NOT1 (N3187, N3163);
or OR2 (N3188, N3186, N356);
not NOT1 (N3189, N3177);
nor NOR3 (N3190, N3175, N2945, N2570);
nor NOR4 (N3191, N3181, N1619, N3151, N2127);
xor XOR2 (N3192, N3149, N1086);
xor XOR2 (N3193, N3140, N2592);
nand NAND2 (N3194, N3187, N886);
not NOT1 (N3195, N3188);
and AND4 (N3196, N3174, N2062, N56, N1009);
buf BUF1 (N3197, N3193);
nand NAND4 (N3198, N3197, N2973, N338, N108);
and AND4 (N3199, N3195, N795, N1516, N1251);
nand NAND3 (N3200, N3198, N2186, N526);
and AND3 (N3201, N3194, N1523, N894);
not NOT1 (N3202, N3190);
xor XOR2 (N3203, N3200, N752);
xor XOR2 (N3204, N3199, N801);
nor NOR2 (N3205, N3201, N699);
or OR2 (N3206, N3205, N2514);
nand NAND4 (N3207, N3192, N1472, N2581, N1406);
and AND2 (N3208, N3191, N3151);
not NOT1 (N3209, N3189);
buf BUF1 (N3210, N3209);
not NOT1 (N3211, N3208);
xor XOR2 (N3212, N3196, N2167);
or OR4 (N3213, N3204, N76, N436, N1799);
nand NAND4 (N3214, N3202, N757, N1564, N2977);
buf BUF1 (N3215, N3214);
or OR2 (N3216, N3184, N2289);
not NOT1 (N3217, N3211);
and AND4 (N3218, N3216, N1332, N121, N754);
not NOT1 (N3219, N3203);
and AND3 (N3220, N3217, N602, N1039);
and AND2 (N3221, N3215, N1520);
buf BUF1 (N3222, N3212);
nor NOR2 (N3223, N3218, N1997);
and AND4 (N3224, N3220, N531, N2132, N515);
not NOT1 (N3225, N3206);
nor NOR3 (N3226, N3210, N2101, N520);
or OR4 (N3227, N3213, N2883, N946, N3146);
nor NOR3 (N3228, N3221, N2615, N1113);
xor XOR2 (N3229, N3207, N1604);
and AND4 (N3230, N3228, N1206, N1474, N1154);
and AND2 (N3231, N3230, N1474);
and AND3 (N3232, N3231, N124, N1208);
xor XOR2 (N3233, N3219, N1521);
or OR2 (N3234, N3185, N3094);
nor NOR2 (N3235, N3222, N826);
buf BUF1 (N3236, N3233);
or OR3 (N3237, N3223, N3149, N2361);
or OR4 (N3238, N3226, N598, N2058, N1974);
xor XOR2 (N3239, N3237, N3191);
or OR3 (N3240, N3235, N35, N1606);
not NOT1 (N3241, N3225);
buf BUF1 (N3242, N3240);
not NOT1 (N3243, N3232);
not NOT1 (N3244, N3241);
and AND2 (N3245, N3229, N2645);
nor NOR4 (N3246, N3242, N896, N1796, N1484);
and AND2 (N3247, N3239, N1360);
nand NAND4 (N3248, N3245, N1373, N2863, N2149);
nand NAND4 (N3249, N3227, N175, N1841, N2290);
not NOT1 (N3250, N3243);
not NOT1 (N3251, N3249);
not NOT1 (N3252, N3238);
nand NAND3 (N3253, N3224, N349, N1621);
or OR2 (N3254, N3251, N1399);
xor XOR2 (N3255, N3248, N2443);
xor XOR2 (N3256, N3255, N2708);
xor XOR2 (N3257, N3250, N2200);
buf BUF1 (N3258, N3253);
buf BUF1 (N3259, N3247);
nor NOR2 (N3260, N3258, N2823);
nor NOR3 (N3261, N3246, N2128, N2226);
and AND2 (N3262, N3257, N1846);
not NOT1 (N3263, N3252);
buf BUF1 (N3264, N3236);
xor XOR2 (N3265, N3264, N1075);
not NOT1 (N3266, N3262);
buf BUF1 (N3267, N3259);
buf BUF1 (N3268, N3267);
nor NOR2 (N3269, N3254, N2591);
not NOT1 (N3270, N3256);
xor XOR2 (N3271, N3265, N2335);
or OR3 (N3272, N3244, N1381, N930);
nand NAND3 (N3273, N3269, N2526, N3161);
nand NAND3 (N3274, N3263, N2914, N1805);
not NOT1 (N3275, N3270);
and AND4 (N3276, N3275, N1559, N393, N894);
nor NOR3 (N3277, N3273, N1448, N1381);
nor NOR4 (N3278, N3266, N2515, N238, N2204);
not NOT1 (N3279, N3268);
nor NOR2 (N3280, N3272, N2101);
xor XOR2 (N3281, N3261, N1970);
xor XOR2 (N3282, N3274, N1299);
buf BUF1 (N3283, N3234);
buf BUF1 (N3284, N3280);
nor NOR3 (N3285, N3260, N3101, N627);
xor XOR2 (N3286, N3281, N1141);
or OR4 (N3287, N3285, N990, N1546, N325);
or OR4 (N3288, N3284, N1184, N259, N3077);
buf BUF1 (N3289, N3277);
not NOT1 (N3290, N3289);
xor XOR2 (N3291, N3283, N1653);
and AND4 (N3292, N3290, N398, N1967, N2821);
xor XOR2 (N3293, N3292, N670);
and AND3 (N3294, N3287, N1127, N1788);
nand NAND3 (N3295, N3278, N1221, N1898);
xor XOR2 (N3296, N3276, N301);
or OR4 (N3297, N3296, N2893, N2931, N1417);
not NOT1 (N3298, N3294);
buf BUF1 (N3299, N3271);
or OR2 (N3300, N3279, N2320);
not NOT1 (N3301, N3282);
or OR4 (N3302, N3293, N734, N2026, N643);
xor XOR2 (N3303, N3300, N3063);
xor XOR2 (N3304, N3299, N247);
not NOT1 (N3305, N3303);
or OR4 (N3306, N3286, N2081, N1856, N407);
buf BUF1 (N3307, N3301);
buf BUF1 (N3308, N3291);
and AND4 (N3309, N3304, N188, N874, N2413);
buf BUF1 (N3310, N3288);
xor XOR2 (N3311, N3305, N199);
and AND3 (N3312, N3311, N927, N1319);
buf BUF1 (N3313, N3307);
xor XOR2 (N3314, N3298, N1923);
and AND2 (N3315, N3306, N1729);
nand NAND2 (N3316, N3310, N377);
nand NAND2 (N3317, N3316, N1146);
or OR3 (N3318, N3309, N397, N3088);
buf BUF1 (N3319, N3297);
buf BUF1 (N3320, N3314);
xor XOR2 (N3321, N3317, N1895);
xor XOR2 (N3322, N3308, N308);
and AND2 (N3323, N3313, N1415);
nor NOR4 (N3324, N3302, N2886, N1521, N3033);
and AND4 (N3325, N3312, N3051, N1260, N1962);
and AND4 (N3326, N3325, N2417, N1144, N1665);
and AND3 (N3327, N3319, N1374, N2079);
and AND3 (N3328, N3318, N3219, N235);
nand NAND3 (N3329, N3323, N809, N316);
not NOT1 (N3330, N3322);
buf BUF1 (N3331, N3328);
xor XOR2 (N3332, N3327, N2054);
and AND4 (N3333, N3295, N2123, N261, N149);
xor XOR2 (N3334, N3329, N1525);
buf BUF1 (N3335, N3315);
or OR3 (N3336, N3331, N124, N2061);
nor NOR4 (N3337, N3320, N125, N2350, N1816);
nand NAND4 (N3338, N3334, N74, N1243, N2981);
not NOT1 (N3339, N3336);
nand NAND2 (N3340, N3326, N3277);
nor NOR2 (N3341, N3340, N1848);
and AND3 (N3342, N3339, N2242, N1924);
nor NOR4 (N3343, N3342, N2227, N1818, N1968);
not NOT1 (N3344, N3343);
not NOT1 (N3345, N3332);
xor XOR2 (N3346, N3338, N1350);
xor XOR2 (N3347, N3333, N3007);
not NOT1 (N3348, N3341);
and AND3 (N3349, N3324, N2604, N2697);
buf BUF1 (N3350, N3330);
buf BUF1 (N3351, N3344);
nor NOR4 (N3352, N3350, N3046, N1830, N346);
or OR2 (N3353, N3348, N2017);
not NOT1 (N3354, N3321);
and AND2 (N3355, N3353, N1972);
xor XOR2 (N3356, N3354, N2204);
buf BUF1 (N3357, N3356);
buf BUF1 (N3358, N3347);
not NOT1 (N3359, N3349);
nor NOR3 (N3360, N3352, N2434, N653);
xor XOR2 (N3361, N3359, N1641);
nand NAND4 (N3362, N3358, N2310, N691, N1106);
and AND4 (N3363, N3361, N2193, N95, N2360);
or OR3 (N3364, N3363, N240, N1314);
and AND4 (N3365, N3345, N3198, N1099, N2679);
nor NOR2 (N3366, N3355, N1264);
not NOT1 (N3367, N3364);
not NOT1 (N3368, N3367);
and AND3 (N3369, N3360, N1149, N3130);
or OR3 (N3370, N3337, N2511, N972);
and AND4 (N3371, N3370, N2047, N3197, N2269);
nor NOR3 (N3372, N3371, N1440, N2309);
or OR3 (N3373, N3346, N3258, N2941);
or OR4 (N3374, N3365, N2756, N3282, N1820);
nor NOR2 (N3375, N3357, N1430);
and AND2 (N3376, N3368, N3360);
buf BUF1 (N3377, N3369);
not NOT1 (N3378, N3375);
xor XOR2 (N3379, N3335, N331);
xor XOR2 (N3380, N3378, N2597);
not NOT1 (N3381, N3366);
buf BUF1 (N3382, N3380);
nor NOR2 (N3383, N3382, N2132);
not NOT1 (N3384, N3377);
xor XOR2 (N3385, N3372, N2540);
or OR2 (N3386, N3379, N2498);
nor NOR4 (N3387, N3362, N253, N2670, N3198);
nand NAND4 (N3388, N3383, N2002, N2993, N2739);
xor XOR2 (N3389, N3386, N1761);
not NOT1 (N3390, N3385);
nor NOR3 (N3391, N3388, N3010, N2204);
or OR2 (N3392, N3390, N1440);
buf BUF1 (N3393, N3351);
not NOT1 (N3394, N3393);
or OR4 (N3395, N3376, N2258, N1062, N69);
or OR4 (N3396, N3381, N570, N586, N1532);
and AND2 (N3397, N3392, N1070);
not NOT1 (N3398, N3384);
and AND4 (N3399, N3398, N1485, N2773, N864);
and AND3 (N3400, N3397, N1901, N1121);
nor NOR3 (N3401, N3395, N838, N1582);
or OR2 (N3402, N3373, N3214);
xor XOR2 (N3403, N3394, N532);
and AND4 (N3404, N3402, N2475, N629, N68);
not NOT1 (N3405, N3391);
not NOT1 (N3406, N3403);
and AND2 (N3407, N3399, N1173);
nor NOR4 (N3408, N3401, N870, N548, N64);
or OR3 (N3409, N3389, N2733, N2502);
nand NAND4 (N3410, N3408, N785, N3131, N2616);
nor NOR4 (N3411, N3400, N1884, N1201, N2701);
buf BUF1 (N3412, N3396);
or OR4 (N3413, N3374, N3302, N3075, N1315);
or OR4 (N3414, N3410, N2661, N1824, N2495);
or OR3 (N3415, N3414, N1478, N1985);
buf BUF1 (N3416, N3405);
or OR2 (N3417, N3411, N1679);
not NOT1 (N3418, N3407);
nand NAND3 (N3419, N3417, N2176, N2140);
buf BUF1 (N3420, N3416);
not NOT1 (N3421, N3419);
or OR3 (N3422, N3409, N1080, N3);
buf BUF1 (N3423, N3422);
nand NAND4 (N3424, N3413, N197, N3319, N2712);
not NOT1 (N3425, N3423);
xor XOR2 (N3426, N3418, N1099);
nand NAND4 (N3427, N3412, N1413, N1742, N1271);
and AND4 (N3428, N3406, N1126, N1770, N2160);
nor NOR4 (N3429, N3428, N2444, N2657, N1790);
nor NOR4 (N3430, N3424, N2180, N159, N2503);
nand NAND2 (N3431, N3421, N66);
xor XOR2 (N3432, N3415, N3218);
not NOT1 (N3433, N3430);
not NOT1 (N3434, N3427);
nand NAND3 (N3435, N3431, N471, N3207);
nand NAND3 (N3436, N3426, N1288, N1745);
and AND3 (N3437, N3387, N1304, N740);
not NOT1 (N3438, N3433);
and AND3 (N3439, N3434, N2451, N3195);
and AND2 (N3440, N3420, N2409);
nor NOR4 (N3441, N3404, N2149, N1655, N3112);
and AND4 (N3442, N3432, N1910, N1242, N2020);
not NOT1 (N3443, N3441);
not NOT1 (N3444, N3425);
or OR3 (N3445, N3442, N2947, N907);
buf BUF1 (N3446, N3438);
or OR2 (N3447, N3429, N364);
and AND4 (N3448, N3436, N25, N1254, N521);
nand NAND3 (N3449, N3437, N1481, N2725);
xor XOR2 (N3450, N3435, N1551);
nor NOR2 (N3451, N3450, N2982);
not NOT1 (N3452, N3444);
nand NAND2 (N3453, N3443, N2140);
and AND2 (N3454, N3452, N2441);
xor XOR2 (N3455, N3449, N2490);
nand NAND3 (N3456, N3440, N2551, N3216);
and AND4 (N3457, N3454, N1340, N3043, N3241);
nor NOR2 (N3458, N3439, N1152);
nor NOR2 (N3459, N3447, N53);
xor XOR2 (N3460, N3456, N1310);
xor XOR2 (N3461, N3455, N1789);
or OR4 (N3462, N3458, N1345, N1861, N1206);
and AND4 (N3463, N3459, N208, N2753, N2232);
buf BUF1 (N3464, N3462);
xor XOR2 (N3465, N3453, N620);
not NOT1 (N3466, N3464);
not NOT1 (N3467, N3463);
nor NOR2 (N3468, N3461, N272);
xor XOR2 (N3469, N3448, N2210);
buf BUF1 (N3470, N3445);
nand NAND4 (N3471, N3469, N2565, N1642, N615);
buf BUF1 (N3472, N3460);
not NOT1 (N3473, N3470);
not NOT1 (N3474, N3451);
nor NOR2 (N3475, N3465, N2664);
not NOT1 (N3476, N3474);
xor XOR2 (N3477, N3466, N2827);
nor NOR2 (N3478, N3446, N2638);
nand NAND3 (N3479, N3475, N228, N1956);
not NOT1 (N3480, N3467);
or OR2 (N3481, N3471, N1861);
not NOT1 (N3482, N3479);
xor XOR2 (N3483, N3476, N1860);
or OR3 (N3484, N3473, N161, N3068);
nor NOR2 (N3485, N3472, N7);
nand NAND3 (N3486, N3457, N943, N532);
not NOT1 (N3487, N3484);
nand NAND3 (N3488, N3483, N319, N1457);
buf BUF1 (N3489, N3478);
xor XOR2 (N3490, N3487, N3258);
or OR4 (N3491, N3490, N350, N2944, N648);
buf BUF1 (N3492, N3477);
and AND4 (N3493, N3488, N3225, N922, N2120);
nand NAND3 (N3494, N3468, N2361, N1587);
xor XOR2 (N3495, N3494, N2096);
xor XOR2 (N3496, N3481, N307);
nor NOR3 (N3497, N3493, N2466, N2960);
and AND4 (N3498, N3489, N221, N2713, N1407);
buf BUF1 (N3499, N3485);
buf BUF1 (N3500, N3495);
nand NAND4 (N3501, N3492, N1500, N2461, N1114);
or OR3 (N3502, N3501, N2378, N1012);
nand NAND3 (N3503, N3498, N1520, N133);
not NOT1 (N3504, N3499);
not NOT1 (N3505, N3491);
xor XOR2 (N3506, N3504, N2019);
nor NOR4 (N3507, N3502, N1042, N2129, N2445);
nand NAND3 (N3508, N3507, N763, N2258);
and AND3 (N3509, N3508, N2777, N340);
or OR2 (N3510, N3503, N2892);
nand NAND4 (N3511, N3510, N14, N488, N1694);
buf BUF1 (N3512, N3482);
not NOT1 (N3513, N3506);
buf BUF1 (N3514, N3512);
or OR4 (N3515, N3496, N265, N385, N2305);
nor NOR4 (N3516, N3486, N20, N2786, N1833);
nor NOR2 (N3517, N3505, N1273);
or OR2 (N3518, N3497, N782);
or OR2 (N3519, N3509, N2803);
buf BUF1 (N3520, N3518);
nor NOR3 (N3521, N3519, N3323, N2199);
not NOT1 (N3522, N3520);
xor XOR2 (N3523, N3522, N2663);
buf BUF1 (N3524, N3500);
nor NOR3 (N3525, N3513, N1114, N1172);
or OR2 (N3526, N3514, N1115);
nand NAND4 (N3527, N3525, N3028, N3455, N1163);
or OR4 (N3528, N3517, N2658, N294, N575);
buf BUF1 (N3529, N3527);
not NOT1 (N3530, N3528);
nand NAND4 (N3531, N3521, N1838, N1951, N1949);
or OR4 (N3532, N3523, N727, N3035, N3052);
or OR2 (N3533, N3529, N2351);
not NOT1 (N3534, N3524);
nor NOR4 (N3535, N3511, N641, N3358, N343);
xor XOR2 (N3536, N3534, N2953);
nor NOR2 (N3537, N3536, N2407);
not NOT1 (N3538, N3532);
xor XOR2 (N3539, N3531, N2505);
nand NAND4 (N3540, N3538, N397, N2443, N1090);
buf BUF1 (N3541, N3537);
or OR4 (N3542, N3540, N3088, N3360, N1963);
buf BUF1 (N3543, N3539);
and AND2 (N3544, N3533, N1584);
nor NOR2 (N3545, N3544, N712);
not NOT1 (N3546, N3542);
nor NOR2 (N3547, N3516, N2426);
buf BUF1 (N3548, N3543);
nand NAND3 (N3549, N3546, N1225, N2247);
not NOT1 (N3550, N3548);
and AND2 (N3551, N3515, N3000);
nor NOR3 (N3552, N3541, N3480, N1280);
xor XOR2 (N3553, N1837, N3225);
and AND4 (N3554, N3545, N3316, N1181, N1257);
not NOT1 (N3555, N3535);
and AND3 (N3556, N3547, N2509, N2409);
nor NOR4 (N3557, N3555, N697, N381, N1541);
or OR4 (N3558, N3557, N2876, N1783, N3195);
or OR3 (N3559, N3554, N2970, N1678);
and AND2 (N3560, N3553, N1445);
buf BUF1 (N3561, N3552);
buf BUF1 (N3562, N3530);
xor XOR2 (N3563, N3561, N448);
buf BUF1 (N3564, N3550);
nor NOR4 (N3565, N3559, N2456, N2688, N212);
not NOT1 (N3566, N3551);
xor XOR2 (N3567, N3565, N3276);
not NOT1 (N3568, N3562);
buf BUF1 (N3569, N3526);
nor NOR2 (N3570, N3566, N852);
nand NAND3 (N3571, N3568, N47, N1337);
nor NOR3 (N3572, N3567, N1145, N509);
xor XOR2 (N3573, N3560, N985);
nand NAND2 (N3574, N3558, N3440);
not NOT1 (N3575, N3571);
not NOT1 (N3576, N3549);
buf BUF1 (N3577, N3564);
buf BUF1 (N3578, N3570);
nand NAND3 (N3579, N3575, N1648, N2660);
nand NAND2 (N3580, N3579, N41);
buf BUF1 (N3581, N3580);
buf BUF1 (N3582, N3569);
nand NAND3 (N3583, N3563, N381, N2658);
buf BUF1 (N3584, N3556);
not NOT1 (N3585, N3581);
xor XOR2 (N3586, N3578, N305);
buf BUF1 (N3587, N3583);
nand NAND4 (N3588, N3585, N1307, N3139, N1073);
xor XOR2 (N3589, N3586, N2803);
xor XOR2 (N3590, N3572, N2767);
nand NAND4 (N3591, N3577, N2138, N1412, N3161);
buf BUF1 (N3592, N3582);
not NOT1 (N3593, N3591);
or OR4 (N3594, N3588, N878, N382, N3570);
and AND4 (N3595, N3576, N1488, N2247, N1649);
nand NAND4 (N3596, N3592, N2671, N2339, N794);
buf BUF1 (N3597, N3573);
xor XOR2 (N3598, N3590, N1627);
xor XOR2 (N3599, N3593, N1700);
nand NAND2 (N3600, N3595, N2729);
not NOT1 (N3601, N3584);
and AND2 (N3602, N3600, N1671);
buf BUF1 (N3603, N3598);
nand NAND2 (N3604, N3574, N3032);
buf BUF1 (N3605, N3602);
nand NAND3 (N3606, N3587, N1294, N1577);
and AND3 (N3607, N3606, N1122, N2704);
nor NOR3 (N3608, N3601, N2853, N2975);
and AND3 (N3609, N3594, N1204, N1104);
or OR2 (N3610, N3603, N3141);
or OR2 (N3611, N3604, N223);
buf BUF1 (N3612, N3610);
buf BUF1 (N3613, N3597);
or OR2 (N3614, N3599, N2291);
not NOT1 (N3615, N3607);
nand NAND4 (N3616, N3615, N1127, N374, N1417);
and AND3 (N3617, N3605, N529, N2741);
not NOT1 (N3618, N3611);
xor XOR2 (N3619, N3616, N3167);
nor NOR4 (N3620, N3618, N3011, N3251, N1763);
buf BUF1 (N3621, N3614);
not NOT1 (N3622, N3619);
or OR4 (N3623, N3622, N608, N2112, N3528);
or OR3 (N3624, N3623, N2305, N3588);
not NOT1 (N3625, N3624);
buf BUF1 (N3626, N3596);
buf BUF1 (N3627, N3589);
buf BUF1 (N3628, N3612);
not NOT1 (N3629, N3628);
and AND3 (N3630, N3621, N250, N120);
and AND4 (N3631, N3629, N2019, N2628, N1060);
xor XOR2 (N3632, N3630, N3379);
buf BUF1 (N3633, N3625);
nor NOR2 (N3634, N3632, N2762);
not NOT1 (N3635, N3633);
or OR2 (N3636, N3634, N1535);
not NOT1 (N3637, N3635);
xor XOR2 (N3638, N3617, N923);
and AND3 (N3639, N3627, N28, N160);
not NOT1 (N3640, N3608);
or OR2 (N3641, N3638, N915);
not NOT1 (N3642, N3613);
nor NOR2 (N3643, N3636, N2174);
buf BUF1 (N3644, N3641);
nand NAND2 (N3645, N3620, N1030);
buf BUF1 (N3646, N3626);
nor NOR4 (N3647, N3645, N2972, N1673, N3400);
and AND2 (N3648, N3643, N2002);
and AND2 (N3649, N3637, N990);
xor XOR2 (N3650, N3642, N1493);
nor NOR4 (N3651, N3649, N664, N3462, N3363);
nor NOR4 (N3652, N3644, N1551, N548, N52);
buf BUF1 (N3653, N3647);
not NOT1 (N3654, N3653);
nand NAND4 (N3655, N3609, N334, N889, N2368);
or OR2 (N3656, N3651, N1623);
not NOT1 (N3657, N3648);
or OR4 (N3658, N3640, N2041, N583, N2148);
not NOT1 (N3659, N3646);
xor XOR2 (N3660, N3639, N1397);
nand NAND2 (N3661, N3659, N3008);
nor NOR3 (N3662, N3631, N3180, N3046);
xor XOR2 (N3663, N3662, N759);
nor NOR4 (N3664, N3654, N1371, N209, N3022);
xor XOR2 (N3665, N3663, N2681);
not NOT1 (N3666, N3661);
or OR3 (N3667, N3656, N2371, N1774);
not NOT1 (N3668, N3652);
or OR2 (N3669, N3668, N419);
nor NOR4 (N3670, N3666, N2219, N750, N43);
nor NOR4 (N3671, N3655, N3634, N2262, N1617);
buf BUF1 (N3672, N3657);
not NOT1 (N3673, N3660);
or OR3 (N3674, N3658, N2522, N60);
nor NOR4 (N3675, N3673, N1982, N608, N1586);
not NOT1 (N3676, N3675);
not NOT1 (N3677, N3672);
not NOT1 (N3678, N3667);
nand NAND4 (N3679, N3665, N2863, N1625, N86);
and AND2 (N3680, N3670, N3371);
buf BUF1 (N3681, N3677);
nand NAND2 (N3682, N3671, N1571);
xor XOR2 (N3683, N3650, N370);
not NOT1 (N3684, N3680);
nor NOR2 (N3685, N3678, N959);
nor NOR4 (N3686, N3674, N229, N1102, N1652);
buf BUF1 (N3687, N3682);
xor XOR2 (N3688, N3687, N2080);
and AND4 (N3689, N3684, N2247, N830, N1989);
not NOT1 (N3690, N3669);
buf BUF1 (N3691, N3664);
nand NAND3 (N3692, N3688, N3361, N249);
not NOT1 (N3693, N3676);
xor XOR2 (N3694, N3685, N3059);
or OR4 (N3695, N3686, N1190, N286, N2187);
or OR4 (N3696, N3683, N934, N1372, N3012);
nand NAND2 (N3697, N3679, N2794);
buf BUF1 (N3698, N3692);
and AND4 (N3699, N3681, N1935, N1317, N2668);
not NOT1 (N3700, N3697);
buf BUF1 (N3701, N3696);
and AND3 (N3702, N3699, N567, N2479);
xor XOR2 (N3703, N3693, N2009);
buf BUF1 (N3704, N3702);
xor XOR2 (N3705, N3703, N423);
buf BUF1 (N3706, N3705);
or OR4 (N3707, N3691, N897, N689, N2516);
nand NAND2 (N3708, N3701, N2819);
xor XOR2 (N3709, N3689, N360);
or OR3 (N3710, N3695, N171, N294);
nor NOR3 (N3711, N3710, N1831, N1478);
xor XOR2 (N3712, N3704, N3074);
buf BUF1 (N3713, N3698);
buf BUF1 (N3714, N3707);
nor NOR3 (N3715, N3714, N2101, N2330);
and AND2 (N3716, N3690, N2492);
buf BUF1 (N3717, N3700);
or OR3 (N3718, N3708, N638, N128);
nor NOR4 (N3719, N3709, N3210, N3680, N2984);
xor XOR2 (N3720, N3706, N3504);
nor NOR2 (N3721, N3720, N2983);
nand NAND3 (N3722, N3713, N3410, N2459);
nand NAND4 (N3723, N3719, N3056, N1240, N941);
xor XOR2 (N3724, N3712, N1491);
nor NOR3 (N3725, N3724, N1362, N408);
nor NOR2 (N3726, N3722, N979);
or OR4 (N3727, N3715, N695, N547, N2775);
nor NOR4 (N3728, N3725, N2876, N342, N1843);
or OR4 (N3729, N3727, N2067, N3346, N1437);
and AND2 (N3730, N3728, N90);
or OR2 (N3731, N3717, N1184);
buf BUF1 (N3732, N3726);
xor XOR2 (N3733, N3723, N304);
not NOT1 (N3734, N3732);
nand NAND3 (N3735, N3716, N2371, N2434);
buf BUF1 (N3736, N3721);
nand NAND2 (N3737, N3711, N654);
or OR2 (N3738, N3731, N2445);
nand NAND3 (N3739, N3738, N880, N181);
or OR3 (N3740, N3730, N3510, N3672);
xor XOR2 (N3741, N3736, N1309);
xor XOR2 (N3742, N3718, N1479);
and AND2 (N3743, N3742, N2673);
buf BUF1 (N3744, N3740);
nand NAND4 (N3745, N3733, N2872, N3309, N1659);
nand NAND3 (N3746, N3734, N2829, N2892);
nor NOR4 (N3747, N3746, N840, N1193, N3274);
nand NAND4 (N3748, N3744, N1045, N1107, N83);
not NOT1 (N3749, N3735);
xor XOR2 (N3750, N3745, N3248);
or OR4 (N3751, N3741, N712, N3302, N1166);
or OR3 (N3752, N3747, N3247, N2115);
and AND3 (N3753, N3748, N3301, N3006);
and AND3 (N3754, N3737, N57, N414);
and AND3 (N3755, N3754, N2272, N3632);
or OR4 (N3756, N3749, N1068, N899, N2205);
and AND4 (N3757, N3753, N3000, N1251, N2581);
not NOT1 (N3758, N3757);
and AND2 (N3759, N3758, N1829);
and AND3 (N3760, N3755, N1579, N430);
xor XOR2 (N3761, N3760, N3395);
or OR3 (N3762, N3729, N3600, N124);
and AND3 (N3763, N3694, N2839, N1542);
nor NOR2 (N3764, N3762, N832);
nor NOR2 (N3765, N3763, N2939);
nor NOR3 (N3766, N3750, N2874, N929);
not NOT1 (N3767, N3752);
or OR2 (N3768, N3756, N1031);
nor NOR3 (N3769, N3767, N3060, N127);
nand NAND3 (N3770, N3739, N2623, N2156);
buf BUF1 (N3771, N3766);
or OR2 (N3772, N3764, N2143);
not NOT1 (N3773, N3759);
or OR3 (N3774, N3773, N945, N2245);
not NOT1 (N3775, N3765);
and AND3 (N3776, N3774, N399, N2902);
buf BUF1 (N3777, N3776);
or OR3 (N3778, N3777, N2547, N3717);
nor NOR2 (N3779, N3761, N1113);
nor NOR2 (N3780, N3771, N1113);
or OR3 (N3781, N3770, N1601, N2351);
and AND3 (N3782, N3743, N1171, N3725);
or OR2 (N3783, N3769, N2275);
buf BUF1 (N3784, N3775);
not NOT1 (N3785, N3772);
nor NOR4 (N3786, N3784, N367, N3250, N480);
or OR2 (N3787, N3786, N1479);
not NOT1 (N3788, N3779);
nor NOR3 (N3789, N3778, N2222, N1837);
not NOT1 (N3790, N3788);
or OR2 (N3791, N3780, N2901);
or OR3 (N3792, N3781, N688, N632);
nor NOR3 (N3793, N3791, N1350, N684);
not NOT1 (N3794, N3768);
buf BUF1 (N3795, N3793);
nand NAND2 (N3796, N3787, N1181);
or OR2 (N3797, N3751, N268);
or OR2 (N3798, N3795, N1852);
or OR3 (N3799, N3789, N430, N3397);
or OR4 (N3800, N3794, N2367, N2676, N2309);
nor NOR4 (N3801, N3799, N1252, N432, N1849);
nor NOR3 (N3802, N3800, N1279, N2071);
nor NOR2 (N3803, N3798, N1693);
and AND4 (N3804, N3801, N1925, N113, N1584);
or OR2 (N3805, N3802, N2276);
or OR2 (N3806, N3783, N2892);
or OR3 (N3807, N3796, N3003, N3087);
nand NAND3 (N3808, N3807, N1309, N403);
buf BUF1 (N3809, N3792);
and AND3 (N3810, N3797, N1539, N2799);
nand NAND4 (N3811, N3806, N3138, N3045, N2788);
buf BUF1 (N3812, N3804);
xor XOR2 (N3813, N3811, N57);
nand NAND4 (N3814, N3782, N2425, N2183, N1994);
nor NOR4 (N3815, N3790, N2097, N3388, N2077);
xor XOR2 (N3816, N3815, N3284);
nand NAND4 (N3817, N3808, N1242, N1207, N3429);
nor NOR2 (N3818, N3785, N2894);
xor XOR2 (N3819, N3803, N2932);
or OR2 (N3820, N3812, N1158);
nor NOR2 (N3821, N3814, N3665);
and AND3 (N3822, N3821, N3122, N1612);
and AND2 (N3823, N3805, N2478);
or OR2 (N3824, N3820, N718);
or OR2 (N3825, N3824, N239);
buf BUF1 (N3826, N3816);
xor XOR2 (N3827, N3818, N1091);
or OR3 (N3828, N3822, N1845, N2842);
not NOT1 (N3829, N3825);
xor XOR2 (N3830, N3819, N280);
buf BUF1 (N3831, N3809);
not NOT1 (N3832, N3827);
xor XOR2 (N3833, N3823, N474);
or OR3 (N3834, N3828, N3380, N531);
xor XOR2 (N3835, N3831, N1534);
not NOT1 (N3836, N3817);
xor XOR2 (N3837, N3835, N3173);
not NOT1 (N3838, N3829);
nand NAND4 (N3839, N3830, N70, N2342, N2414);
and AND2 (N3840, N3813, N747);
and AND2 (N3841, N3832, N1825);
buf BUF1 (N3842, N3810);
nand NAND4 (N3843, N3842, N3131, N2556, N522);
or OR2 (N3844, N3826, N3140);
nand NAND2 (N3845, N3844, N2153);
nand NAND3 (N3846, N3841, N1037, N1984);
xor XOR2 (N3847, N3839, N756);
or OR3 (N3848, N3846, N1767, N729);
not NOT1 (N3849, N3848);
nand NAND4 (N3850, N3838, N2820, N622, N2900);
or OR3 (N3851, N3849, N2380, N275);
and AND4 (N3852, N3840, N1942, N1116, N3210);
nand NAND2 (N3853, N3847, N184);
not NOT1 (N3854, N3843);
or OR4 (N3855, N3854, N3425, N830, N3255);
and AND4 (N3856, N3855, N3832, N1405, N2766);
not NOT1 (N3857, N3856);
or OR2 (N3858, N3857, N849);
or OR3 (N3859, N3852, N3633, N2113);
nor NOR3 (N3860, N3837, N3053, N2276);
and AND3 (N3861, N3860, N2153, N966);
not NOT1 (N3862, N3850);
not NOT1 (N3863, N3861);
and AND2 (N3864, N3851, N2891);
not NOT1 (N3865, N3863);
not NOT1 (N3866, N3833);
xor XOR2 (N3867, N3858, N1518);
not NOT1 (N3868, N3864);
nor NOR4 (N3869, N3845, N1502, N1877, N2804);
xor XOR2 (N3870, N3862, N1696);
xor XOR2 (N3871, N3853, N1134);
not NOT1 (N3872, N3868);
and AND3 (N3873, N3867, N2626, N3093);
nand NAND4 (N3874, N3834, N235, N1731, N2187);
nor NOR2 (N3875, N3865, N3144);
nor NOR2 (N3876, N3872, N1747);
nand NAND4 (N3877, N3866, N1107, N2616, N3140);
not NOT1 (N3878, N3876);
not NOT1 (N3879, N3878);
or OR3 (N3880, N3859, N1933, N1091);
buf BUF1 (N3881, N3836);
xor XOR2 (N3882, N3881, N286);
not NOT1 (N3883, N3880);
not NOT1 (N3884, N3874);
buf BUF1 (N3885, N3884);
not NOT1 (N3886, N3871);
buf BUF1 (N3887, N3869);
not NOT1 (N3888, N3875);
and AND2 (N3889, N3882, N365);
nand NAND4 (N3890, N3873, N1557, N1147, N3824);
nor NOR2 (N3891, N3886, N1448);
xor XOR2 (N3892, N3877, N3843);
or OR4 (N3893, N3888, N3310, N1677, N637);
xor XOR2 (N3894, N3887, N3784);
nor NOR2 (N3895, N3885, N1597);
not NOT1 (N3896, N3891);
nor NOR3 (N3897, N3890, N2262, N3329);
nor NOR2 (N3898, N3893, N3868);
not NOT1 (N3899, N3883);
or OR4 (N3900, N3898, N3075, N1459, N1828);
or OR3 (N3901, N3889, N2689, N2442);
nand NAND3 (N3902, N3870, N3850, N913);
or OR2 (N3903, N3902, N2949);
and AND2 (N3904, N3899, N417);
buf BUF1 (N3905, N3900);
nand NAND4 (N3906, N3894, N1375, N2357, N1918);
or OR3 (N3907, N3903, N1759, N976);
xor XOR2 (N3908, N3896, N1552);
nor NOR4 (N3909, N3906, N836, N714, N507);
buf BUF1 (N3910, N3909);
nor NOR2 (N3911, N3910, N1520);
xor XOR2 (N3912, N3904, N3092);
xor XOR2 (N3913, N3908, N250);
or OR4 (N3914, N3901, N647, N3526, N2328);
nand NAND4 (N3915, N3895, N3912, N1922, N2729);
nand NAND4 (N3916, N3286, N3015, N1589, N1194);
and AND2 (N3917, N3907, N2180);
or OR4 (N3918, N3915, N3535, N1079, N3510);
or OR4 (N3919, N3897, N3238, N3186, N589);
or OR2 (N3920, N3892, N2135);
nand NAND4 (N3921, N3914, N3329, N3423, N2947);
xor XOR2 (N3922, N3911, N2887);
or OR4 (N3923, N3913, N3610, N139, N264);
and AND3 (N3924, N3923, N382, N1656);
nand NAND2 (N3925, N3918, N1070);
nor NOR2 (N3926, N3925, N417);
not NOT1 (N3927, N3926);
not NOT1 (N3928, N3924);
nand NAND4 (N3929, N3916, N3119, N1972, N3392);
not NOT1 (N3930, N3919);
buf BUF1 (N3931, N3917);
not NOT1 (N3932, N3928);
nand NAND2 (N3933, N3920, N140);
and AND3 (N3934, N3922, N2164, N1809);
nor NOR4 (N3935, N3927, N3628, N1948, N2238);
nand NAND4 (N3936, N3930, N2547, N37, N3849);
and AND2 (N3937, N3935, N2189);
or OR4 (N3938, N3879, N3159, N3413, N1163);
and AND2 (N3939, N3905, N3202);
not NOT1 (N3940, N3931);
and AND3 (N3941, N3937, N951, N523);
not NOT1 (N3942, N3936);
and AND3 (N3943, N3933, N1202, N2571);
or OR4 (N3944, N3939, N1141, N3553, N770);
nand NAND3 (N3945, N3943, N1077, N1187);
nand NAND2 (N3946, N3944, N1646);
not NOT1 (N3947, N3938);
or OR3 (N3948, N3942, N2644, N3605);
buf BUF1 (N3949, N3934);
nand NAND2 (N3950, N3921, N2660);
nor NOR2 (N3951, N3932, N2575);
xor XOR2 (N3952, N3950, N3767);
or OR4 (N3953, N3951, N2077, N244, N1264);
buf BUF1 (N3954, N3952);
nor NOR3 (N3955, N3948, N3731, N133);
nor NOR2 (N3956, N3947, N2474);
nand NAND3 (N3957, N3954, N2518, N1003);
nand NAND4 (N3958, N3955, N2082, N795, N813);
not NOT1 (N3959, N3946);
or OR4 (N3960, N3953, N1101, N1945, N82);
xor XOR2 (N3961, N3940, N896);
and AND4 (N3962, N3949, N435, N1298, N2816);
or OR2 (N3963, N3945, N1770);
xor XOR2 (N3964, N3957, N3715);
and AND4 (N3965, N3941, N3623, N1157, N2345);
buf BUF1 (N3966, N3962);
buf BUF1 (N3967, N3929);
nor NOR4 (N3968, N3964, N2258, N2279, N3326);
nor NOR4 (N3969, N3965, N2741, N543, N3356);
not NOT1 (N3970, N3959);
nor NOR3 (N3971, N3960, N2627, N3113);
not NOT1 (N3972, N3969);
nor NOR4 (N3973, N3961, N1998, N1607, N3554);
nand NAND2 (N3974, N3973, N3296);
not NOT1 (N3975, N3974);
or OR2 (N3976, N3967, N2770);
xor XOR2 (N3977, N3976, N1331);
and AND2 (N3978, N3963, N1243);
buf BUF1 (N3979, N3972);
xor XOR2 (N3980, N3958, N3618);
not NOT1 (N3981, N3978);
buf BUF1 (N3982, N3970);
xor XOR2 (N3983, N3980, N232);
buf BUF1 (N3984, N3977);
buf BUF1 (N3985, N3975);
nor NOR3 (N3986, N3968, N2058, N2415);
nor NOR4 (N3987, N3956, N2441, N1795, N485);
buf BUF1 (N3988, N3986);
nand NAND3 (N3989, N3981, N3336, N2826);
xor XOR2 (N3990, N3982, N2261);
xor XOR2 (N3991, N3984, N2418);
and AND3 (N3992, N3987, N1383, N992);
xor XOR2 (N3993, N3992, N1502);
nand NAND2 (N3994, N3966, N2935);
and AND2 (N3995, N3979, N3386);
or OR2 (N3996, N3994, N1328);
and AND2 (N3997, N3995, N1137);
and AND3 (N3998, N3991, N1087, N1986);
xor XOR2 (N3999, N3993, N801);
buf BUF1 (N4000, N3998);
and AND3 (N4001, N3985, N2950, N2329);
nor NOR2 (N4002, N3990, N1812);
xor XOR2 (N4003, N3999, N2455);
not NOT1 (N4004, N3983);
not NOT1 (N4005, N3996);
buf BUF1 (N4006, N3989);
and AND3 (N4007, N4001, N10, N3933);
xor XOR2 (N4008, N3997, N55);
and AND4 (N4009, N4004, N1496, N1515, N2333);
or OR4 (N4010, N3971, N3155, N519, N1848);
not NOT1 (N4011, N3988);
nand NAND4 (N4012, N4009, N2883, N3036, N198);
or OR3 (N4013, N4006, N3610, N2754);
or OR3 (N4014, N4007, N2548, N3866);
nand NAND2 (N4015, N4010, N1295);
not NOT1 (N4016, N4015);
nor NOR2 (N4017, N4016, N919);
and AND3 (N4018, N4008, N2633, N1710);
buf BUF1 (N4019, N4005);
xor XOR2 (N4020, N4003, N3737);
and AND4 (N4021, N4018, N829, N1974, N2658);
xor XOR2 (N4022, N4002, N3011);
nand NAND4 (N4023, N4011, N3815, N3106, N3058);
not NOT1 (N4024, N4014);
nand NAND2 (N4025, N4020, N2545);
and AND3 (N4026, N4012, N3256, N2059);
buf BUF1 (N4027, N4024);
or OR2 (N4028, N4022, N2631);
xor XOR2 (N4029, N4021, N3447);
and AND2 (N4030, N4026, N1163);
nand NAND4 (N4031, N4027, N1969, N3000, N3144);
or OR2 (N4032, N4025, N2183);
xor XOR2 (N4033, N4031, N3271);
buf BUF1 (N4034, N4028);
nor NOR3 (N4035, N4029, N1358, N1327);
nor NOR3 (N4036, N4017, N3792, N1881);
not NOT1 (N4037, N4034);
nor NOR4 (N4038, N4035, N2527, N1673, N3587);
nor NOR3 (N4039, N4037, N3473, N1513);
nor NOR2 (N4040, N4013, N2053);
and AND4 (N4041, N4033, N939, N2133, N2146);
and AND2 (N4042, N4039, N3172);
nand NAND2 (N4043, N4041, N144);
buf BUF1 (N4044, N4042);
nand NAND2 (N4045, N4036, N1434);
not NOT1 (N4046, N4045);
not NOT1 (N4047, N4000);
nand NAND2 (N4048, N4032, N2243);
and AND3 (N4049, N4023, N2400, N649);
and AND3 (N4050, N4047, N534, N3015);
or OR3 (N4051, N4044, N290, N3334);
buf BUF1 (N4052, N4050);
buf BUF1 (N4053, N4048);
xor XOR2 (N4054, N4046, N300);
and AND2 (N4055, N4019, N1331);
nand NAND2 (N4056, N4052, N119);
not NOT1 (N4057, N4051);
or OR2 (N4058, N4040, N3989);
and AND3 (N4059, N4057, N1697, N2336);
xor XOR2 (N4060, N4059, N820);
nor NOR2 (N4061, N4049, N533);
buf BUF1 (N4062, N4043);
and AND2 (N4063, N4054, N2210);
not NOT1 (N4064, N4030);
not NOT1 (N4065, N4062);
nand NAND3 (N4066, N4058, N1830, N2318);
not NOT1 (N4067, N4065);
nand NAND3 (N4068, N4060, N2582, N2061);
or OR3 (N4069, N4066, N3503, N2357);
nor NOR2 (N4070, N4068, N2373);
nand NAND3 (N4071, N4064, N41, N413);
buf BUF1 (N4072, N4055);
xor XOR2 (N4073, N4067, N321);
nand NAND2 (N4074, N4061, N3680);
and AND3 (N4075, N4063, N2430, N630);
nor NOR2 (N4076, N4056, N3557);
xor XOR2 (N4077, N4070, N3212);
or OR4 (N4078, N4074, N1442, N797, N1769);
or OR2 (N4079, N4072, N3884);
not NOT1 (N4080, N4053);
and AND2 (N4081, N4079, N3659);
not NOT1 (N4082, N4073);
xor XOR2 (N4083, N4075, N1932);
nand NAND2 (N4084, N4083, N2118);
nand NAND3 (N4085, N4069, N2250, N2111);
xor XOR2 (N4086, N4078, N3325);
buf BUF1 (N4087, N4071);
nand NAND4 (N4088, N4077, N315, N1155, N1414);
nor NOR4 (N4089, N4082, N1259, N1763, N1743);
or OR4 (N4090, N4080, N1876, N360, N3954);
and AND3 (N4091, N4081, N1492, N1457);
nand NAND2 (N4092, N4088, N3985);
buf BUF1 (N4093, N4038);
nand NAND4 (N4094, N4089, N3374, N3446, N2302);
buf BUF1 (N4095, N4086);
or OR2 (N4096, N4094, N3553);
not NOT1 (N4097, N4090);
and AND4 (N4098, N4091, N3318, N1728, N652);
nand NAND3 (N4099, N4098, N3197, N2408);
not NOT1 (N4100, N4085);
not NOT1 (N4101, N4099);
nand NAND3 (N4102, N4095, N2137, N1775);
nor NOR4 (N4103, N4093, N386, N3694, N134);
nor NOR4 (N4104, N4084, N1468, N1966, N1209);
and AND4 (N4105, N4101, N3890, N2690, N2953);
or OR3 (N4106, N4097, N119, N1242);
or OR4 (N4107, N4100, N3614, N205, N3850);
not NOT1 (N4108, N4103);
nor NOR4 (N4109, N4102, N387, N2620, N2432);
buf BUF1 (N4110, N4092);
xor XOR2 (N4111, N4106, N2575);
buf BUF1 (N4112, N4109);
xor XOR2 (N4113, N4076, N1461);
or OR4 (N4114, N4105, N2304, N1587, N2709);
xor XOR2 (N4115, N4107, N3510);
nand NAND2 (N4116, N4110, N3902);
nor NOR4 (N4117, N4104, N1083, N850, N1210);
or OR3 (N4118, N4116, N3674, N441);
nor NOR3 (N4119, N4118, N921, N2826);
not NOT1 (N4120, N4119);
buf BUF1 (N4121, N4117);
nand NAND3 (N4122, N4087, N2054, N320);
nand NAND3 (N4123, N4112, N1310, N2159);
not NOT1 (N4124, N4115);
buf BUF1 (N4125, N4113);
nor NOR2 (N4126, N4124, N2866);
buf BUF1 (N4127, N4125);
xor XOR2 (N4128, N4108, N1389);
nand NAND2 (N4129, N4120, N890);
buf BUF1 (N4130, N4129);
xor XOR2 (N4131, N4127, N3210);
or OR2 (N4132, N4122, N2301);
and AND2 (N4133, N4130, N2805);
and AND4 (N4134, N4121, N2675, N1723, N3073);
xor XOR2 (N4135, N4096, N1076);
nor NOR4 (N4136, N4126, N2550, N1125, N3328);
or OR4 (N4137, N4114, N197, N673, N2986);
nand NAND2 (N4138, N4136, N2545);
or OR2 (N4139, N4111, N787);
xor XOR2 (N4140, N4138, N1393);
xor XOR2 (N4141, N4135, N3717);
nor NOR3 (N4142, N4123, N939, N543);
nand NAND3 (N4143, N4132, N1794, N79);
nor NOR3 (N4144, N4133, N1500, N4136);
nand NAND3 (N4145, N4140, N692, N602);
or OR2 (N4146, N4144, N2256);
nor NOR2 (N4147, N4131, N2368);
buf BUF1 (N4148, N4128);
or OR4 (N4149, N4147, N2436, N2461, N48);
not NOT1 (N4150, N4145);
buf BUF1 (N4151, N4134);
buf BUF1 (N4152, N4151);
not NOT1 (N4153, N4152);
or OR2 (N4154, N4148, N190);
and AND4 (N4155, N4150, N1170, N1987, N2553);
and AND2 (N4156, N4141, N2348);
nand NAND2 (N4157, N4149, N636);
or OR4 (N4158, N4142, N1922, N760, N3089);
nand NAND2 (N4159, N4146, N1045);
or OR3 (N4160, N4154, N4096, N2531);
not NOT1 (N4161, N4160);
buf BUF1 (N4162, N4153);
xor XOR2 (N4163, N4159, N585);
or OR3 (N4164, N4163, N1779, N2698);
and AND2 (N4165, N4143, N1274);
nand NAND3 (N4166, N4156, N1016, N3688);
buf BUF1 (N4167, N4137);
xor XOR2 (N4168, N4157, N3942);
and AND4 (N4169, N4168, N1686, N3706, N1538);
buf BUF1 (N4170, N4166);
not NOT1 (N4171, N4161);
buf BUF1 (N4172, N4169);
xor XOR2 (N4173, N4162, N262);
not NOT1 (N4174, N4171);
buf BUF1 (N4175, N4167);
nor NOR2 (N4176, N4172, N1501);
buf BUF1 (N4177, N4164);
buf BUF1 (N4178, N4173);
and AND3 (N4179, N4178, N769, N1000);
nand NAND3 (N4180, N4158, N1143, N1090);
nand NAND4 (N4181, N4179, N3623, N3918, N1181);
not NOT1 (N4182, N4174);
or OR3 (N4183, N4139, N1555, N1523);
xor XOR2 (N4184, N4177, N126);
not NOT1 (N4185, N4183);
and AND4 (N4186, N4175, N2497, N2114, N338);
or OR4 (N4187, N4181, N1027, N436, N2858);
and AND2 (N4188, N4180, N3731);
buf BUF1 (N4189, N4155);
buf BUF1 (N4190, N4188);
buf BUF1 (N4191, N4184);
nand NAND3 (N4192, N4182, N698, N399);
and AND3 (N4193, N4165, N3916, N4021);
nand NAND3 (N4194, N4193, N3011, N4140);
and AND3 (N4195, N4189, N2069, N941);
buf BUF1 (N4196, N4187);
nor NOR2 (N4197, N4186, N3318);
buf BUF1 (N4198, N4195);
and AND2 (N4199, N4192, N918);
nor NOR3 (N4200, N4185, N2577, N3930);
nand NAND3 (N4201, N4170, N3792, N3192);
nor NOR3 (N4202, N4200, N352, N3123);
nor NOR2 (N4203, N4197, N2310);
not NOT1 (N4204, N4194);
xor XOR2 (N4205, N4203, N1710);
nand NAND4 (N4206, N4205, N2757, N3646, N3595);
xor XOR2 (N4207, N4198, N3921);
or OR4 (N4208, N4206, N1486, N2183, N3327);
and AND3 (N4209, N4208, N682, N2765);
nor NOR4 (N4210, N4209, N2693, N3466, N4025);
not NOT1 (N4211, N4202);
not NOT1 (N4212, N4191);
nor NOR2 (N4213, N4204, N537);
xor XOR2 (N4214, N4207, N3483);
buf BUF1 (N4215, N4196);
buf BUF1 (N4216, N4212);
nor NOR4 (N4217, N4213, N1816, N3788, N1809);
xor XOR2 (N4218, N4210, N1935);
xor XOR2 (N4219, N4217, N75);
nor NOR4 (N4220, N4190, N865, N998, N3935);
nand NAND3 (N4221, N4211, N3296, N720);
or OR3 (N4222, N4214, N1686, N2499);
nor NOR2 (N4223, N4201, N483);
not NOT1 (N4224, N4176);
or OR2 (N4225, N4199, N308);
buf BUF1 (N4226, N4223);
not NOT1 (N4227, N4222);
xor XOR2 (N4228, N4215, N2794);
or OR2 (N4229, N4216, N2263);
and AND3 (N4230, N4218, N1484, N959);
xor XOR2 (N4231, N4220, N2515);
xor XOR2 (N4232, N4231, N303);
buf BUF1 (N4233, N4219);
or OR3 (N4234, N4229, N3425, N701);
or OR4 (N4235, N4226, N394, N3011, N1073);
nand NAND2 (N4236, N4228, N2530);
xor XOR2 (N4237, N4225, N1563);
xor XOR2 (N4238, N4224, N1893);
nor NOR2 (N4239, N4236, N3298);
or OR4 (N4240, N4235, N3191, N90, N3278);
or OR2 (N4241, N4240, N3137);
xor XOR2 (N4242, N4234, N2250);
nand NAND2 (N4243, N4242, N2861);
xor XOR2 (N4244, N4241, N3174);
nor NOR4 (N4245, N4237, N1632, N406, N3015);
nand NAND3 (N4246, N4244, N1601, N1624);
nor NOR2 (N4247, N4243, N772);
not NOT1 (N4248, N4238);
nand NAND4 (N4249, N4233, N1117, N1756, N338);
not NOT1 (N4250, N4227);
buf BUF1 (N4251, N4239);
and AND3 (N4252, N4248, N1583, N4160);
nand NAND3 (N4253, N4250, N516, N4027);
not NOT1 (N4254, N4251);
nand NAND3 (N4255, N4246, N2760, N72);
not NOT1 (N4256, N4255);
and AND3 (N4257, N4253, N2492, N4158);
buf BUF1 (N4258, N4232);
nand NAND3 (N4259, N4249, N1308, N4110);
nand NAND3 (N4260, N4245, N2605, N3091);
or OR3 (N4261, N4247, N2052, N670);
and AND2 (N4262, N4256, N448);
not NOT1 (N4263, N4254);
or OR3 (N4264, N4259, N2828, N226);
xor XOR2 (N4265, N4230, N1254);
nor NOR2 (N4266, N4258, N156);
xor XOR2 (N4267, N4252, N2933);
nand NAND3 (N4268, N4265, N2770, N2560);
not NOT1 (N4269, N4266);
nor NOR2 (N4270, N4257, N546);
nor NOR4 (N4271, N4264, N1486, N4072, N1042);
and AND2 (N4272, N4221, N2317);
xor XOR2 (N4273, N4270, N1715);
or OR2 (N4274, N4269, N2345);
nor NOR4 (N4275, N4263, N1967, N1250, N1533);
buf BUF1 (N4276, N4275);
nand NAND4 (N4277, N4260, N3240, N1839, N4038);
not NOT1 (N4278, N4273);
not NOT1 (N4279, N4261);
or OR4 (N4280, N4267, N3012, N1121, N2973);
nand NAND4 (N4281, N4278, N3036, N224, N1541);
buf BUF1 (N4282, N4277);
xor XOR2 (N4283, N4262, N2971);
buf BUF1 (N4284, N4274);
nor NOR4 (N4285, N4280, N4148, N409, N2827);
nand NAND4 (N4286, N4276, N3461, N2828, N212);
not NOT1 (N4287, N4271);
or OR4 (N4288, N4282, N2269, N2736, N1621);
nor NOR4 (N4289, N4287, N3603, N2194, N330);
not NOT1 (N4290, N4281);
nand NAND3 (N4291, N4285, N2462, N1863);
nand NAND4 (N4292, N4288, N1708, N3749, N482);
xor XOR2 (N4293, N4289, N4106);
and AND2 (N4294, N4286, N356);
or OR3 (N4295, N4284, N1066, N2241);
or OR4 (N4296, N4272, N5, N182, N1698);
and AND4 (N4297, N4292, N1633, N2969, N2390);
and AND3 (N4298, N4295, N3008, N2349);
nor NOR2 (N4299, N4291, N2312);
nand NAND4 (N4300, N4296, N1223, N3924, N2801);
nand NAND4 (N4301, N4299, N635, N3297, N4142);
nand NAND3 (N4302, N4294, N2574, N2842);
nand NAND4 (N4303, N4302, N4119, N3993, N1007);
not NOT1 (N4304, N4293);
nand NAND2 (N4305, N4279, N1871);
nand NAND3 (N4306, N4298, N3609, N254);
and AND2 (N4307, N4283, N1934);
buf BUF1 (N4308, N4306);
or OR4 (N4309, N4304, N3978, N3670, N2885);
nor NOR2 (N4310, N4300, N1728);
nor NOR4 (N4311, N4309, N1066, N1017, N1992);
nand NAND2 (N4312, N4303, N2847);
or OR4 (N4313, N4312, N3939, N2511, N2504);
xor XOR2 (N4314, N4297, N962);
and AND2 (N4315, N4311, N612);
nor NOR2 (N4316, N4315, N1763);
nand NAND4 (N4317, N4268, N631, N4239, N1746);
buf BUF1 (N4318, N4308);
or OR2 (N4319, N4313, N4269);
nor NOR2 (N4320, N4317, N1384);
nand NAND3 (N4321, N4310, N1636, N1283);
or OR4 (N4322, N4301, N1558, N1610, N1716);
buf BUF1 (N4323, N4290);
nand NAND2 (N4324, N4321, N2076);
buf BUF1 (N4325, N4318);
or OR2 (N4326, N4316, N3987);
nand NAND3 (N4327, N4326, N194, N2336);
xor XOR2 (N4328, N4325, N2601);
not NOT1 (N4329, N4322);
nand NAND2 (N4330, N4320, N30);
or OR2 (N4331, N4314, N2660);
nor NOR3 (N4332, N4330, N3695, N1369);
buf BUF1 (N4333, N4307);
and AND4 (N4334, N4323, N3995, N3506, N3543);
not NOT1 (N4335, N4305);
or OR3 (N4336, N4332, N142, N1158);
not NOT1 (N4337, N4329);
nor NOR3 (N4338, N4328, N2747, N1791);
buf BUF1 (N4339, N4331);
and AND2 (N4340, N4333, N2964);
buf BUF1 (N4341, N4335);
or OR3 (N4342, N4340, N464, N2743);
nand NAND3 (N4343, N4336, N589, N1422);
not NOT1 (N4344, N4341);
nand NAND2 (N4345, N4324, N4177);
and AND3 (N4346, N4319, N3264, N1667);
and AND4 (N4347, N4338, N2429, N3199, N4154);
not NOT1 (N4348, N4337);
buf BUF1 (N4349, N4327);
xor XOR2 (N4350, N4334, N973);
or OR2 (N4351, N4350, N1291);
buf BUF1 (N4352, N4349);
and AND3 (N4353, N4352, N1131, N2372);
or OR4 (N4354, N4339, N3435, N2504, N3852);
or OR4 (N4355, N4351, N155, N2738, N3435);
not NOT1 (N4356, N4353);
xor XOR2 (N4357, N4355, N1811);
xor XOR2 (N4358, N4347, N2950);
nor NOR2 (N4359, N4348, N3921);
nor NOR2 (N4360, N4344, N3933);
buf BUF1 (N4361, N4357);
or OR4 (N4362, N4342, N2289, N4270, N3016);
nor NOR3 (N4363, N4358, N3461, N1332);
not NOT1 (N4364, N4361);
nor NOR3 (N4365, N4362, N4360, N290);
xor XOR2 (N4366, N2063, N3034);
and AND2 (N4367, N4366, N3593);
xor XOR2 (N4368, N4346, N401);
xor XOR2 (N4369, N4368, N4006);
or OR4 (N4370, N4354, N3954, N53, N1858);
buf BUF1 (N4371, N4356);
nor NOR3 (N4372, N4370, N2880, N3693);
not NOT1 (N4373, N4365);
buf BUF1 (N4374, N4371);
nor NOR4 (N4375, N4343, N2227, N10, N2924);
nand NAND2 (N4376, N4374, N3864);
nand NAND3 (N4377, N4375, N334, N3352);
buf BUF1 (N4378, N4372);
buf BUF1 (N4379, N4359);
nand NAND2 (N4380, N4379, N500);
or OR2 (N4381, N4376, N547);
buf BUF1 (N4382, N4364);
nor NOR3 (N4383, N4363, N2728, N595);
or OR4 (N4384, N4377, N3307, N464, N3057);
buf BUF1 (N4385, N4369);
not NOT1 (N4386, N4383);
or OR3 (N4387, N4384, N572, N1657);
or OR3 (N4388, N4367, N2038, N1274);
nand NAND3 (N4389, N4378, N309, N2311);
buf BUF1 (N4390, N4373);
buf BUF1 (N4391, N4380);
or OR2 (N4392, N4381, N2060);
nand NAND3 (N4393, N4386, N2983, N2903);
buf BUF1 (N4394, N4385);
nor NOR4 (N4395, N4345, N164, N4138, N2083);
buf BUF1 (N4396, N4390);
nand NAND4 (N4397, N4389, N2873, N2914, N2966);
and AND3 (N4398, N4393, N2782, N4166);
or OR4 (N4399, N4398, N1060, N2848, N571);
xor XOR2 (N4400, N4399, N3928);
nor NOR2 (N4401, N4387, N578);
and AND2 (N4402, N4391, N485);
not NOT1 (N4403, N4382);
nand NAND3 (N4404, N4396, N2280, N1489);
or OR3 (N4405, N4403, N3728, N3093);
not NOT1 (N4406, N4388);
nor NOR2 (N4407, N4392, N3678);
nand NAND3 (N4408, N4405, N3228, N1997);
and AND2 (N4409, N4395, N1560);
nor NOR4 (N4410, N4407, N2775, N2205, N583);
and AND3 (N4411, N4397, N881, N272);
buf BUF1 (N4412, N4410);
not NOT1 (N4413, N4400);
xor XOR2 (N4414, N4411, N3757);
or OR3 (N4415, N4402, N1045, N93);
nor NOR2 (N4416, N4413, N2179);
nand NAND3 (N4417, N4401, N2021, N1597);
nor NOR2 (N4418, N4404, N2445);
not NOT1 (N4419, N4416);
nand NAND4 (N4420, N4418, N1440, N817, N969);
buf BUF1 (N4421, N4394);
buf BUF1 (N4422, N4409);
buf BUF1 (N4423, N4414);
xor XOR2 (N4424, N4421, N2591);
nor NOR2 (N4425, N4419, N3295);
buf BUF1 (N4426, N4423);
and AND4 (N4427, N4408, N3496, N2018, N1365);
and AND3 (N4428, N4425, N2955, N2560);
buf BUF1 (N4429, N4420);
or OR3 (N4430, N4412, N2714, N1438);
and AND4 (N4431, N4428, N3770, N4171, N1606);
nor NOR3 (N4432, N4424, N1184, N4216);
and AND3 (N4433, N4431, N2130, N1008);
xor XOR2 (N4434, N4430, N431);
and AND4 (N4435, N4406, N4009, N2400, N4222);
buf BUF1 (N4436, N4429);
buf BUF1 (N4437, N4435);
nand NAND3 (N4438, N4426, N4132, N3157);
nand NAND4 (N4439, N4427, N3980, N166, N1851);
nor NOR3 (N4440, N4434, N88, N1021);
nor NOR2 (N4441, N4440, N1695);
xor XOR2 (N4442, N4436, N3971);
and AND3 (N4443, N4432, N164, N4395);
and AND3 (N4444, N4433, N3352, N2395);
nand NAND3 (N4445, N4417, N3765, N3032);
or OR2 (N4446, N4422, N58);
xor XOR2 (N4447, N4415, N3327);
nand NAND3 (N4448, N4441, N774, N1730);
xor XOR2 (N4449, N4439, N1307);
or OR4 (N4450, N4449, N2984, N3674, N1600);
nand NAND3 (N4451, N4444, N3686, N2435);
not NOT1 (N4452, N4448);
not NOT1 (N4453, N4452);
nand NAND2 (N4454, N4438, N1821);
not NOT1 (N4455, N4453);
xor XOR2 (N4456, N4447, N3151);
not NOT1 (N4457, N4442);
nand NAND3 (N4458, N4445, N90, N3968);
nand NAND4 (N4459, N4450, N2572, N3870, N2133);
nor NOR2 (N4460, N4455, N1193);
buf BUF1 (N4461, N4443);
buf BUF1 (N4462, N4458);
buf BUF1 (N4463, N4454);
buf BUF1 (N4464, N4437);
not NOT1 (N4465, N4446);
nor NOR2 (N4466, N4457, N2662);
and AND3 (N4467, N4456, N566, N2992);
nand NAND3 (N4468, N4464, N3816, N594);
buf BUF1 (N4469, N4462);
nand NAND4 (N4470, N4463, N3102, N3440, N903);
buf BUF1 (N4471, N4466);
or OR3 (N4472, N4470, N2340, N4103);
xor XOR2 (N4473, N4468, N4139);
xor XOR2 (N4474, N4473, N2737);
not NOT1 (N4475, N4451);
nor NOR2 (N4476, N4461, N40);
and AND2 (N4477, N4467, N692);
and AND3 (N4478, N4471, N146, N373);
buf BUF1 (N4479, N4460);
nand NAND2 (N4480, N4476, N1865);
and AND4 (N4481, N4475, N2643, N671, N3798);
xor XOR2 (N4482, N4472, N1645);
and AND3 (N4483, N4469, N2781, N1308);
and AND2 (N4484, N4477, N146);
buf BUF1 (N4485, N4479);
xor XOR2 (N4486, N4485, N1158);
buf BUF1 (N4487, N4480);
nor NOR4 (N4488, N4483, N329, N928, N833);
or OR2 (N4489, N4486, N3083);
buf BUF1 (N4490, N4482);
not NOT1 (N4491, N4490);
nand NAND4 (N4492, N4487, N1486, N2043, N4383);
buf BUF1 (N4493, N4492);
and AND2 (N4494, N4493, N3969);
buf BUF1 (N4495, N4465);
buf BUF1 (N4496, N4489);
xor XOR2 (N4497, N4481, N3233);
not NOT1 (N4498, N4474);
and AND3 (N4499, N4478, N3896, N3080);
nand NAND4 (N4500, N4494, N3093, N4101, N2037);
nand NAND3 (N4501, N4495, N3574, N1815);
buf BUF1 (N4502, N4496);
or OR3 (N4503, N4500, N2107, N3473);
and AND3 (N4504, N4484, N3205, N1370);
or OR4 (N4505, N4459, N410, N1855, N4169);
and AND3 (N4506, N4501, N121, N4399);
or OR3 (N4507, N4497, N3004, N711);
nand NAND3 (N4508, N4507, N3982, N1453);
buf BUF1 (N4509, N4498);
or OR4 (N4510, N4488, N2245, N2718, N2776);
xor XOR2 (N4511, N4509, N1808);
nand NAND2 (N4512, N4502, N3530);
buf BUF1 (N4513, N4508);
or OR4 (N4514, N4510, N4193, N2289, N1132);
buf BUF1 (N4515, N4506);
nor NOR4 (N4516, N4511, N318, N4267, N4108);
xor XOR2 (N4517, N4514, N467);
or OR4 (N4518, N4517, N1303, N1249, N227);
nor NOR2 (N4519, N4516, N2805);
nor NOR2 (N4520, N4512, N1586);
nor NOR3 (N4521, N4513, N4015, N3514);
and AND2 (N4522, N4504, N3975);
xor XOR2 (N4523, N4505, N2807);
nand NAND4 (N4524, N4491, N1911, N3418, N3451);
xor XOR2 (N4525, N4524, N3952);
xor XOR2 (N4526, N4521, N1236);
buf BUF1 (N4527, N4525);
nor NOR4 (N4528, N4526, N1920, N619, N1910);
nor NOR4 (N4529, N4518, N309, N2567, N1823);
or OR4 (N4530, N4520, N2109, N1741, N3165);
or OR4 (N4531, N4530, N656, N1953, N1979);
or OR4 (N4532, N4531, N1293, N2087, N147);
not NOT1 (N4533, N4515);
nand NAND3 (N4534, N4519, N2628, N309);
or OR2 (N4535, N4503, N3588);
buf BUF1 (N4536, N4529);
or OR2 (N4537, N4528, N1474);
nor NOR4 (N4538, N4499, N4188, N2253, N4275);
nand NAND4 (N4539, N4535, N817, N2080, N3880);
xor XOR2 (N4540, N4522, N1771);
or OR2 (N4541, N4539, N3599);
nand NAND3 (N4542, N4527, N4, N2043);
or OR2 (N4543, N4523, N1722);
and AND4 (N4544, N4537, N2937, N3090, N866);
or OR2 (N4545, N4533, N3350);
buf BUF1 (N4546, N4541);
nor NOR3 (N4547, N4534, N3367, N3884);
nand NAND4 (N4548, N4543, N835, N2420, N1041);
or OR3 (N4549, N4548, N3297, N2289);
or OR2 (N4550, N4547, N1901);
or OR3 (N4551, N4545, N4478, N1769);
xor XOR2 (N4552, N4532, N3064);
and AND4 (N4553, N4544, N4079, N2439, N755);
and AND4 (N4554, N4536, N443, N3053, N2259);
and AND2 (N4555, N4554, N3693);
xor XOR2 (N4556, N4540, N2073);
buf BUF1 (N4557, N4549);
xor XOR2 (N4558, N4551, N1341);
not NOT1 (N4559, N4557);
or OR2 (N4560, N4553, N4033);
xor XOR2 (N4561, N4560, N3328);
not NOT1 (N4562, N4561);
nor NOR3 (N4563, N4546, N3678, N148);
buf BUF1 (N4564, N4542);
or OR2 (N4565, N4555, N1311);
xor XOR2 (N4566, N4558, N2183);
buf BUF1 (N4567, N4565);
nor NOR4 (N4568, N4552, N2990, N1506, N1047);
nor NOR2 (N4569, N4538, N4419);
and AND4 (N4570, N4566, N3998, N3393, N3783);
buf BUF1 (N4571, N4567);
nand NAND3 (N4572, N4568, N210, N3977);
and AND3 (N4573, N4569, N1190, N1803);
buf BUF1 (N4574, N4571);
not NOT1 (N4575, N4550);
nand NAND3 (N4576, N4573, N1199, N3242);
nand NAND3 (N4577, N4575, N1836, N3499);
buf BUF1 (N4578, N4577);
or OR4 (N4579, N4556, N80, N1314, N2749);
not NOT1 (N4580, N4562);
not NOT1 (N4581, N4570);
and AND3 (N4582, N4574, N207, N1659);
nor NOR2 (N4583, N4578, N2606);
buf BUF1 (N4584, N4576);
and AND4 (N4585, N4581, N4304, N4237, N2412);
nand NAND4 (N4586, N4572, N1715, N1963, N3332);
nand NAND2 (N4587, N4584, N1141);
buf BUF1 (N4588, N4587);
or OR4 (N4589, N4582, N984, N1923, N2508);
nor NOR4 (N4590, N4583, N653, N4311, N4495);
nor NOR2 (N4591, N4564, N2906);
nor NOR2 (N4592, N4579, N3014);
or OR4 (N4593, N4559, N1679, N3205, N3964);
not NOT1 (N4594, N4586);
nand NAND2 (N4595, N4588, N2579);
not NOT1 (N4596, N4589);
not NOT1 (N4597, N4596);
buf BUF1 (N4598, N4591);
nor NOR3 (N4599, N4580, N3332, N746);
and AND2 (N4600, N4598, N3509);
nor NOR4 (N4601, N4595, N2918, N3183, N2158);
or OR2 (N4602, N4594, N2776);
nand NAND4 (N4603, N4597, N3231, N609, N2518);
nand NAND3 (N4604, N4592, N2652, N926);
nand NAND2 (N4605, N4604, N2665);
and AND2 (N4606, N4593, N2120);
buf BUF1 (N4607, N4585);
and AND2 (N4608, N4590, N1744);
nor NOR3 (N4609, N4600, N4563, N2837);
xor XOR2 (N4610, N2967, N672);
buf BUF1 (N4611, N4608);
buf BUF1 (N4612, N4606);
nor NOR2 (N4613, N4605, N616);
xor XOR2 (N4614, N4609, N2770);
buf BUF1 (N4615, N4607);
nor NOR3 (N4616, N4603, N2220, N602);
xor XOR2 (N4617, N4599, N2723);
nand NAND4 (N4618, N4602, N3581, N2607, N2867);
or OR2 (N4619, N4618, N4539);
buf BUF1 (N4620, N4611);
or OR4 (N4621, N4619, N2026, N3057, N2508);
or OR2 (N4622, N4610, N1538);
or OR4 (N4623, N4622, N3641, N842, N3102);
and AND3 (N4624, N4601, N887, N4177);
nor NOR4 (N4625, N4613, N2813, N1522, N4346);
and AND3 (N4626, N4612, N1433, N1250);
buf BUF1 (N4627, N4621);
or OR3 (N4628, N4617, N733, N3104);
nand NAND4 (N4629, N4628, N1311, N2727, N394);
or OR3 (N4630, N4625, N4509, N2631);
buf BUF1 (N4631, N4626);
buf BUF1 (N4632, N4627);
xor XOR2 (N4633, N4631, N1828);
buf BUF1 (N4634, N4632);
nand NAND3 (N4635, N4623, N4564, N4069);
nand NAND2 (N4636, N4630, N2101);
xor XOR2 (N4637, N4636, N1405);
xor XOR2 (N4638, N4615, N3007);
and AND2 (N4639, N4635, N2530);
buf BUF1 (N4640, N4639);
buf BUF1 (N4641, N4633);
nand NAND4 (N4642, N4641, N1283, N887, N2196);
and AND2 (N4643, N4642, N1639);
or OR4 (N4644, N4643, N3948, N926, N3083);
not NOT1 (N4645, N4644);
not NOT1 (N4646, N4629);
not NOT1 (N4647, N4620);
buf BUF1 (N4648, N4624);
or OR2 (N4649, N4640, N587);
buf BUF1 (N4650, N4649);
nand NAND3 (N4651, N4637, N1543, N1513);
buf BUF1 (N4652, N4634);
or OR4 (N4653, N4614, N1295, N2790, N569);
not NOT1 (N4654, N4646);
nor NOR4 (N4655, N4616, N4231, N3749, N1130);
nor NOR2 (N4656, N4655, N2890);
or OR2 (N4657, N4648, N410);
nor NOR3 (N4658, N4651, N1741, N4257);
or OR3 (N4659, N4656, N3892, N2680);
xor XOR2 (N4660, N4658, N3049);
nand NAND3 (N4661, N4650, N280, N293);
and AND3 (N4662, N4661, N584, N3245);
not NOT1 (N4663, N4638);
nand NAND2 (N4664, N4652, N3790);
xor XOR2 (N4665, N4662, N99);
and AND3 (N4666, N4645, N2613, N3540);
buf BUF1 (N4667, N4657);
nor NOR4 (N4668, N4647, N2605, N4446, N2100);
and AND4 (N4669, N4663, N2097, N3322, N792);
xor XOR2 (N4670, N4668, N999);
or OR4 (N4671, N4664, N2658, N4529, N2891);
and AND3 (N4672, N4670, N708, N2688);
buf BUF1 (N4673, N4665);
buf BUF1 (N4674, N4653);
buf BUF1 (N4675, N4660);
and AND2 (N4676, N4667, N4075);
buf BUF1 (N4677, N4674);
nor NOR3 (N4678, N4666, N4609, N3186);
not NOT1 (N4679, N4672);
and AND2 (N4680, N4679, N2453);
or OR3 (N4681, N4676, N3615, N637);
xor XOR2 (N4682, N4678, N3999);
xor XOR2 (N4683, N4681, N2270);
and AND4 (N4684, N4673, N378, N3059, N1518);
not NOT1 (N4685, N4684);
and AND4 (N4686, N4680, N75, N769, N1282);
or OR4 (N4687, N4654, N2715, N1387, N1315);
nor NOR4 (N4688, N4687, N3180, N3931, N3802);
xor XOR2 (N4689, N4683, N1538);
not NOT1 (N4690, N4677);
and AND3 (N4691, N4669, N4424, N1777);
xor XOR2 (N4692, N4659, N4241);
nand NAND3 (N4693, N4689, N3243, N4231);
xor XOR2 (N4694, N4686, N3070);
not NOT1 (N4695, N4690);
not NOT1 (N4696, N4692);
nand NAND3 (N4697, N4675, N138, N2290);
and AND2 (N4698, N4682, N2734);
nor NOR4 (N4699, N4691, N1499, N776, N2960);
nand NAND3 (N4700, N4671, N1945, N4496);
nand NAND2 (N4701, N4688, N778);
not NOT1 (N4702, N4700);
and AND4 (N4703, N4693, N1785, N194, N139);
or OR3 (N4704, N4699, N4152, N1323);
and AND2 (N4705, N4701, N672);
xor XOR2 (N4706, N4702, N2243);
and AND3 (N4707, N4695, N1647, N1565);
or OR4 (N4708, N4697, N2890, N3808, N4038);
buf BUF1 (N4709, N4705);
or OR3 (N4710, N4704, N2912, N889);
not NOT1 (N4711, N4707);
or OR2 (N4712, N4696, N2554);
xor XOR2 (N4713, N4709, N4135);
nand NAND3 (N4714, N4713, N1219, N2770);
or OR4 (N4715, N4694, N2301, N1984, N2114);
not NOT1 (N4716, N4706);
nor NOR4 (N4717, N4708, N629, N360, N27);
xor XOR2 (N4718, N4711, N1283);
nand NAND4 (N4719, N4703, N2897, N2626, N1644);
xor XOR2 (N4720, N4710, N189);
xor XOR2 (N4721, N4717, N3506);
buf BUF1 (N4722, N4716);
nand NAND2 (N4723, N4712, N3039);
xor XOR2 (N4724, N4715, N3323);
buf BUF1 (N4725, N4698);
or OR3 (N4726, N4723, N1512, N3668);
nor NOR2 (N4727, N4725, N103);
nand NAND2 (N4728, N4727, N1244);
and AND4 (N4729, N4728, N3359, N658, N2441);
nand NAND2 (N4730, N4718, N364);
buf BUF1 (N4731, N4719);
nand NAND2 (N4732, N4685, N796);
nor NOR2 (N4733, N4721, N4146);
nor NOR2 (N4734, N4724, N3567);
nand NAND2 (N4735, N4729, N121);
nand NAND4 (N4736, N4732, N156, N2220, N2870);
buf BUF1 (N4737, N4731);
not NOT1 (N4738, N4737);
nor NOR4 (N4739, N4730, N2501, N1968, N1515);
buf BUF1 (N4740, N4738);
buf BUF1 (N4741, N4736);
and AND4 (N4742, N4733, N430, N3307, N4605);
xor XOR2 (N4743, N4726, N3761);
buf BUF1 (N4744, N4743);
buf BUF1 (N4745, N4741);
nand NAND2 (N4746, N4720, N3389);
xor XOR2 (N4747, N4714, N3904);
xor XOR2 (N4748, N4722, N1118);
not NOT1 (N4749, N4744);
buf BUF1 (N4750, N4747);
or OR4 (N4751, N4749, N837, N644, N2238);
or OR3 (N4752, N4735, N1344, N662);
nor NOR4 (N4753, N4752, N4140, N4148, N84);
xor XOR2 (N4754, N4751, N2099);
xor XOR2 (N4755, N4750, N2808);
xor XOR2 (N4756, N4746, N9);
buf BUF1 (N4757, N4745);
nor NOR2 (N4758, N4754, N3110);
not NOT1 (N4759, N4748);
and AND4 (N4760, N4757, N924, N1223, N869);
buf BUF1 (N4761, N4740);
buf BUF1 (N4762, N4761);
xor XOR2 (N4763, N4759, N202);
or OR2 (N4764, N4756, N2848);
and AND4 (N4765, N4742, N855, N1803, N2379);
and AND4 (N4766, N4739, N212, N4273, N2339);
buf BUF1 (N4767, N4734);
buf BUF1 (N4768, N4764);
nor NOR3 (N4769, N4767, N589, N209);
not NOT1 (N4770, N4760);
nor NOR2 (N4771, N4768, N4645);
buf BUF1 (N4772, N4766);
or OR2 (N4773, N4765, N4157);
nor NOR2 (N4774, N4770, N2478);
buf BUF1 (N4775, N4772);
nand NAND2 (N4776, N4755, N2934);
not NOT1 (N4777, N4771);
not NOT1 (N4778, N4777);
buf BUF1 (N4779, N4775);
not NOT1 (N4780, N4778);
nand NAND3 (N4781, N4776, N1456, N221);
nor NOR2 (N4782, N4779, N3410);
or OR4 (N4783, N4782, N1213, N4132, N2598);
buf BUF1 (N4784, N4763);
buf BUF1 (N4785, N4753);
buf BUF1 (N4786, N4783);
nand NAND2 (N4787, N4785, N4706);
not NOT1 (N4788, N4787);
buf BUF1 (N4789, N4788);
and AND2 (N4790, N4774, N77);
or OR3 (N4791, N4780, N1175, N1678);
nor NOR3 (N4792, N4784, N785, N2540);
xor XOR2 (N4793, N4781, N1223);
buf BUF1 (N4794, N4773);
or OR4 (N4795, N4769, N2528, N1734, N2245);
or OR2 (N4796, N4795, N3898);
xor XOR2 (N4797, N4789, N2741);
and AND4 (N4798, N4796, N4773, N1767, N4284);
buf BUF1 (N4799, N4790);
or OR3 (N4800, N4797, N1082, N2993);
not NOT1 (N4801, N4786);
buf BUF1 (N4802, N4793);
nand NAND2 (N4803, N4794, N2740);
nor NOR2 (N4804, N4762, N3757);
xor XOR2 (N4805, N4798, N632);
nor NOR4 (N4806, N4803, N1765, N4058, N2422);
or OR3 (N4807, N4806, N1120, N3741);
nand NAND4 (N4808, N4791, N3441, N4173, N3235);
nand NAND2 (N4809, N4804, N2698);
or OR4 (N4810, N4758, N423, N545, N4090);
buf BUF1 (N4811, N4799);
and AND4 (N4812, N4800, N3272, N1534, N4743);
buf BUF1 (N4813, N4801);
nor NOR4 (N4814, N4802, N3688, N2766, N2720);
not NOT1 (N4815, N4813);
nand NAND3 (N4816, N4792, N4252, N3258);
buf BUF1 (N4817, N4816);
nor NOR4 (N4818, N4807, N1206, N3087, N2086);
not NOT1 (N4819, N4814);
nor NOR2 (N4820, N4810, N2840);
nor NOR4 (N4821, N4817, N703, N4555, N920);
nor NOR2 (N4822, N4821, N1465);
buf BUF1 (N4823, N4808);
and AND2 (N4824, N4812, N3133);
and AND2 (N4825, N4815, N962);
nor NOR4 (N4826, N4823, N1903, N2627, N2231);
nor NOR3 (N4827, N4818, N72, N3347);
xor XOR2 (N4828, N4827, N1412);
xor XOR2 (N4829, N4820, N2481);
and AND2 (N4830, N4822, N4687);
buf BUF1 (N4831, N4825);
not NOT1 (N4832, N4824);
not NOT1 (N4833, N4829);
xor XOR2 (N4834, N4833, N1922);
nor NOR2 (N4835, N4834, N18);
nor NOR4 (N4836, N4830, N3732, N2105, N2430);
and AND2 (N4837, N4835, N1282);
nand NAND2 (N4838, N4832, N3045);
or OR2 (N4839, N4836, N1084);
nand NAND4 (N4840, N4828, N747, N3217, N1735);
nor NOR4 (N4841, N4809, N2374, N1085, N3409);
buf BUF1 (N4842, N4839);
and AND2 (N4843, N4837, N2600);
and AND4 (N4844, N4842, N2867, N4084, N4066);
buf BUF1 (N4845, N4841);
not NOT1 (N4846, N4826);
and AND4 (N4847, N4843, N3892, N2767, N297);
nor NOR3 (N4848, N4811, N1912, N3693);
buf BUF1 (N4849, N4844);
nor NOR3 (N4850, N4846, N570, N3953);
xor XOR2 (N4851, N4805, N3703);
buf BUF1 (N4852, N4850);
nand NAND3 (N4853, N4848, N351, N2687);
and AND3 (N4854, N4840, N1394, N2308);
nor NOR2 (N4855, N4845, N775);
or OR3 (N4856, N4838, N2170, N1814);
xor XOR2 (N4857, N4851, N3404);
buf BUF1 (N4858, N4856);
not NOT1 (N4859, N4852);
nor NOR2 (N4860, N4849, N818);
nor NOR3 (N4861, N4819, N380, N1457);
not NOT1 (N4862, N4859);
buf BUF1 (N4863, N4831);
nor NOR3 (N4864, N4858, N2350, N3598);
nand NAND4 (N4865, N4863, N1758, N3542, N1228);
nand NAND2 (N4866, N4860, N2163);
buf BUF1 (N4867, N4865);
buf BUF1 (N4868, N4853);
nor NOR3 (N4869, N4847, N734, N2061);
and AND4 (N4870, N4855, N1759, N2829, N3229);
xor XOR2 (N4871, N4869, N4836);
or OR2 (N4872, N4868, N4735);
buf BUF1 (N4873, N4866);
nor NOR2 (N4874, N4857, N1046);
nand NAND4 (N4875, N4872, N3935, N947, N4385);
not NOT1 (N4876, N4871);
not NOT1 (N4877, N4876);
nand NAND3 (N4878, N4874, N1415, N350);
or OR4 (N4879, N4877, N4702, N2383, N2203);
not NOT1 (N4880, N4875);
not NOT1 (N4881, N4867);
xor XOR2 (N4882, N4864, N1806);
xor XOR2 (N4883, N4878, N4622);
and AND3 (N4884, N4883, N822, N3979);
or OR3 (N4885, N4882, N1219, N3710);
and AND2 (N4886, N4880, N1286);
xor XOR2 (N4887, N4873, N3587);
not NOT1 (N4888, N4887);
nor NOR4 (N4889, N4862, N990, N3380, N518);
and AND2 (N4890, N4881, N4314);
nand NAND2 (N4891, N4885, N1837);
not NOT1 (N4892, N4870);
xor XOR2 (N4893, N4891, N1612);
or OR4 (N4894, N4884, N2816, N3744, N4528);
nor NOR2 (N4895, N4894, N1582);
not NOT1 (N4896, N4893);
nor NOR2 (N4897, N4861, N400);
buf BUF1 (N4898, N4890);
nand NAND4 (N4899, N4888, N4808, N1638, N1310);
xor XOR2 (N4900, N4895, N1922);
nand NAND3 (N4901, N4886, N1967, N2975);
not NOT1 (N4902, N4854);
not NOT1 (N4903, N4879);
and AND3 (N4904, N4889, N1273, N1148);
nor NOR2 (N4905, N4892, N395);
xor XOR2 (N4906, N4900, N3048);
xor XOR2 (N4907, N4896, N911);
xor XOR2 (N4908, N4905, N1046);
or OR2 (N4909, N4904, N2291);
not NOT1 (N4910, N4897);
not NOT1 (N4911, N4902);
nand NAND4 (N4912, N4899, N1703, N2796, N2426);
nor NOR3 (N4913, N4901, N3193, N619);
nor NOR3 (N4914, N4903, N4323, N2968);
and AND3 (N4915, N4914, N2049, N1357);
not NOT1 (N4916, N4913);
buf BUF1 (N4917, N4906);
buf BUF1 (N4918, N4911);
or OR3 (N4919, N4909, N3435, N37);
nor NOR2 (N4920, N4912, N2393);
nor NOR3 (N4921, N4917, N2489, N4422);
xor XOR2 (N4922, N4919, N219);
not NOT1 (N4923, N4908);
buf BUF1 (N4924, N4922);
buf BUF1 (N4925, N4921);
buf BUF1 (N4926, N4920);
not NOT1 (N4927, N4923);
or OR2 (N4928, N4927, N116);
xor XOR2 (N4929, N4928, N1731);
not NOT1 (N4930, N4898);
nand NAND2 (N4931, N4925, N1344);
buf BUF1 (N4932, N4926);
nand NAND4 (N4933, N4918, N4340, N611, N3248);
xor XOR2 (N4934, N4916, N328);
not NOT1 (N4935, N4930);
nor NOR4 (N4936, N4934, N4374, N2865, N892);
and AND2 (N4937, N4932, N325);
buf BUF1 (N4938, N4907);
and AND4 (N4939, N4915, N920, N2855, N3334);
or OR4 (N4940, N4933, N2516, N2452, N2422);
xor XOR2 (N4941, N4924, N2762);
xor XOR2 (N4942, N4935, N4295);
and AND4 (N4943, N4938, N4067, N3630, N3579);
and AND2 (N4944, N4943, N4821);
nor NOR2 (N4945, N4942, N1792);
buf BUF1 (N4946, N4931);
nor NOR4 (N4947, N4910, N3893, N3092, N1286);
nand NAND4 (N4948, N4947, N4358, N2885, N338);
or OR3 (N4949, N4948, N4534, N3414);
nand NAND3 (N4950, N4944, N1139, N2135);
xor XOR2 (N4951, N4950, N2689);
buf BUF1 (N4952, N4940);
and AND2 (N4953, N4946, N626);
nor NOR3 (N4954, N4953, N716, N3483);
xor XOR2 (N4955, N4939, N1219);
buf BUF1 (N4956, N4945);
nor NOR4 (N4957, N4956, N2058, N4925, N2312);
xor XOR2 (N4958, N4952, N2234);
buf BUF1 (N4959, N4958);
buf BUF1 (N4960, N4955);
buf BUF1 (N4961, N4936);
and AND4 (N4962, N4959, N1643, N2113, N2105);
not NOT1 (N4963, N4951);
not NOT1 (N4964, N4941);
xor XOR2 (N4965, N4954, N2194);
or OR3 (N4966, N4960, N4041, N4297);
and AND4 (N4967, N4957, N2153, N3092, N3041);
xor XOR2 (N4968, N4929, N3460);
and AND3 (N4969, N4949, N4032, N2712);
nand NAND4 (N4970, N4963, N3773, N4965, N2963);
and AND4 (N4971, N4509, N3872, N4447, N981);
nand NAND2 (N4972, N4968, N1770);
nand NAND2 (N4973, N4967, N576);
and AND3 (N4974, N4962, N3008, N2804);
nor NOR2 (N4975, N4974, N1522);
nor NOR3 (N4976, N4973, N2450, N3087);
and AND2 (N4977, N4971, N3428);
buf BUF1 (N4978, N4937);
xor XOR2 (N4979, N4964, N3419);
nand NAND3 (N4980, N4979, N2713, N4269);
or OR3 (N4981, N4977, N1971, N2488);
or OR2 (N4982, N4981, N1391);
nand NAND4 (N4983, N4975, N3764, N3654, N2261);
not NOT1 (N4984, N4982);
nor NOR3 (N4985, N4961, N2291, N2564);
xor XOR2 (N4986, N4978, N1005);
buf BUF1 (N4987, N4983);
buf BUF1 (N4988, N4972);
and AND4 (N4989, N4976, N4749, N4042, N3558);
nor NOR2 (N4990, N4989, N2672);
buf BUF1 (N4991, N4970);
not NOT1 (N4992, N4990);
and AND2 (N4993, N4992, N3947);
xor XOR2 (N4994, N4987, N3076);
xor XOR2 (N4995, N4994, N3575);
or OR2 (N4996, N4966, N578);
not NOT1 (N4997, N4995);
xor XOR2 (N4998, N4988, N3380);
nor NOR4 (N4999, N4993, N1653, N3356, N2230);
xor XOR2 (N5000, N4998, N4969);
xor XOR2 (N5001, N926, N1948);
not NOT1 (N5002, N4999);
not NOT1 (N5003, N4980);
and AND4 (N5004, N4991, N3574, N2122, N3384);
nor NOR3 (N5005, N4997, N4604, N4767);
buf BUF1 (N5006, N5000);
or OR4 (N5007, N5002, N835, N2287, N1726);
buf BUF1 (N5008, N4984);
and AND3 (N5009, N5007, N3927, N2065);
xor XOR2 (N5010, N5003, N1337);
xor XOR2 (N5011, N5006, N2190);
nor NOR2 (N5012, N5008, N704);
and AND4 (N5013, N5012, N2885, N3136, N2617);
nor NOR2 (N5014, N5011, N3765);
not NOT1 (N5015, N4985);
buf BUF1 (N5016, N5001);
nor NOR3 (N5017, N5015, N1237, N4924);
or OR3 (N5018, N5013, N2525, N718);
nor NOR4 (N5019, N5004, N3677, N4961, N4512);
buf BUF1 (N5020, N5014);
not NOT1 (N5021, N4986);
nand NAND4 (N5022, N4996, N1570, N187, N2961);
xor XOR2 (N5023, N5009, N862);
buf BUF1 (N5024, N5010);
or OR3 (N5025, N5020, N3704, N938);
xor XOR2 (N5026, N5022, N1211);
nand NAND2 (N5027, N5021, N869);
nor NOR2 (N5028, N5024, N4385);
nor NOR3 (N5029, N5023, N3590, N1679);
xor XOR2 (N5030, N5017, N4392);
not NOT1 (N5031, N5016);
buf BUF1 (N5032, N5029);
nor NOR2 (N5033, N5031, N3442);
nor NOR4 (N5034, N5032, N714, N2268, N3549);
not NOT1 (N5035, N5028);
and AND3 (N5036, N5019, N3960, N719);
not NOT1 (N5037, N5025);
or OR3 (N5038, N5027, N4440, N424);
not NOT1 (N5039, N5036);
nand NAND2 (N5040, N5034, N3669);
xor XOR2 (N5041, N5005, N4073);
buf BUF1 (N5042, N5018);
nor NOR2 (N5043, N5026, N2956);
xor XOR2 (N5044, N5039, N4846);
xor XOR2 (N5045, N5033, N1169);
xor XOR2 (N5046, N5043, N36);
xor XOR2 (N5047, N5030, N221);
or OR4 (N5048, N5045, N3045, N2095, N970);
xor XOR2 (N5049, N5047, N3168);
nor NOR3 (N5050, N5035, N1437, N828);
and AND4 (N5051, N5038, N4098, N781, N3574);
nor NOR2 (N5052, N5042, N3929);
nor NOR3 (N5053, N5048, N4879, N2853);
and AND3 (N5054, N5053, N763, N78);
not NOT1 (N5055, N5037);
nor NOR2 (N5056, N5049, N2110);
and AND4 (N5057, N5041, N744, N3179, N4514);
not NOT1 (N5058, N5056);
and AND4 (N5059, N5055, N2852, N609, N1968);
buf BUF1 (N5060, N5054);
not NOT1 (N5061, N5060);
nor NOR3 (N5062, N5044, N4767, N4788);
not NOT1 (N5063, N5062);
not NOT1 (N5064, N5059);
nand NAND4 (N5065, N5040, N796, N5035, N2370);
or OR2 (N5066, N5064, N2057);
nor NOR3 (N5067, N5051, N2540, N3467);
buf BUF1 (N5068, N5058);
and AND3 (N5069, N5067, N2027, N3988);
nand NAND3 (N5070, N5046, N945, N4186);
xor XOR2 (N5071, N5052, N55);
or OR2 (N5072, N5050, N2462);
xor XOR2 (N5073, N5063, N789);
nand NAND2 (N5074, N5071, N1795);
or OR3 (N5075, N5074, N3682, N2964);
nand NAND4 (N5076, N5068, N743, N1758, N1699);
buf BUF1 (N5077, N5073);
buf BUF1 (N5078, N5070);
and AND2 (N5079, N5076, N1545);
or OR2 (N5080, N5061, N817);
nand NAND3 (N5081, N5072, N4457, N2522);
or OR3 (N5082, N5078, N2017, N3201);
buf BUF1 (N5083, N5066);
xor XOR2 (N5084, N5082, N4794);
and AND3 (N5085, N5057, N4087, N1396);
nor NOR4 (N5086, N5080, N4836, N4031, N304);
xor XOR2 (N5087, N5081, N4317);
or OR2 (N5088, N5069, N814);
or OR3 (N5089, N5075, N1101, N1587);
nand NAND2 (N5090, N5079, N684);
and AND4 (N5091, N5086, N880, N56, N2575);
nor NOR2 (N5092, N5084, N4863);
nor NOR2 (N5093, N5089, N2807);
buf BUF1 (N5094, N5077);
buf BUF1 (N5095, N5091);
nor NOR2 (N5096, N5093, N2135);
nor NOR2 (N5097, N5092, N1313);
nor NOR3 (N5098, N5090, N271, N1798);
not NOT1 (N5099, N5094);
xor XOR2 (N5100, N5065, N4518);
xor XOR2 (N5101, N5100, N2649);
or OR2 (N5102, N5085, N5084);
xor XOR2 (N5103, N5097, N1725);
buf BUF1 (N5104, N5099);
or OR3 (N5105, N5083, N1072, N3194);
buf BUF1 (N5106, N5105);
nand NAND4 (N5107, N5106, N1733, N3243, N2123);
buf BUF1 (N5108, N5098);
buf BUF1 (N5109, N5101);
not NOT1 (N5110, N5102);
and AND2 (N5111, N5096, N1815);
xor XOR2 (N5112, N5109, N2741);
xor XOR2 (N5113, N5087, N3732);
nor NOR4 (N5114, N5113, N2090, N2268, N173);
and AND4 (N5115, N5110, N1100, N1186, N4631);
not NOT1 (N5116, N5088);
nand NAND2 (N5117, N5103, N2348);
xor XOR2 (N5118, N5107, N4561);
or OR4 (N5119, N5111, N4640, N3207, N1366);
or OR4 (N5120, N5116, N1596, N4674, N4401);
xor XOR2 (N5121, N5095, N4612);
and AND3 (N5122, N5118, N3090, N933);
not NOT1 (N5123, N5117);
buf BUF1 (N5124, N5122);
and AND3 (N5125, N5121, N4320, N2465);
nand NAND4 (N5126, N5104, N1307, N3083, N3748);
nor NOR3 (N5127, N5112, N1529, N3057);
buf BUF1 (N5128, N5108);
buf BUF1 (N5129, N5120);
nor NOR4 (N5130, N5126, N4566, N3353, N4428);
buf BUF1 (N5131, N5123);
buf BUF1 (N5132, N5125);
xor XOR2 (N5133, N5119, N1376);
and AND3 (N5134, N5115, N4103, N1816);
nand NAND2 (N5135, N5130, N1464);
xor XOR2 (N5136, N5135, N2657);
nor NOR3 (N5137, N5136, N349, N2886);
nor NOR3 (N5138, N5127, N2446, N3481);
or OR2 (N5139, N5128, N1193);
buf BUF1 (N5140, N5138);
buf BUF1 (N5141, N5133);
and AND3 (N5142, N5141, N3911, N4415);
not NOT1 (N5143, N5124);
buf BUF1 (N5144, N5142);
nor NOR4 (N5145, N5140, N4872, N3446, N4256);
and AND2 (N5146, N5132, N2387);
or OR3 (N5147, N5143, N217, N476);
buf BUF1 (N5148, N5147);
nand NAND4 (N5149, N5148, N3720, N4544, N3720);
or OR3 (N5150, N5114, N4740, N654);
buf BUF1 (N5151, N5150);
and AND2 (N5152, N5145, N3262);
nand NAND4 (N5153, N5149, N3559, N5027, N3521);
buf BUF1 (N5154, N5129);
or OR2 (N5155, N5137, N4244);
buf BUF1 (N5156, N5155);
or OR2 (N5157, N5146, N4476);
nor NOR4 (N5158, N5139, N562, N4812, N1242);
or OR4 (N5159, N5156, N883, N3036, N564);
or OR2 (N5160, N5151, N214);
and AND2 (N5161, N5134, N2846);
nor NOR4 (N5162, N5154, N4718, N1635, N4794);
or OR2 (N5163, N5131, N4534);
or OR4 (N5164, N5163, N1684, N4413, N318);
or OR2 (N5165, N5161, N1096);
xor XOR2 (N5166, N5158, N710);
not NOT1 (N5167, N5166);
buf BUF1 (N5168, N5144);
xor XOR2 (N5169, N5167, N5130);
nor NOR2 (N5170, N5164, N1959);
and AND2 (N5171, N5152, N4589);
and AND4 (N5172, N5171, N4234, N2548, N5095);
xor XOR2 (N5173, N5172, N473);
and AND3 (N5174, N5169, N1380, N2123);
and AND4 (N5175, N5173, N478, N4851, N1633);
buf BUF1 (N5176, N5174);
or OR3 (N5177, N5176, N2584, N852);
nand NAND3 (N5178, N5162, N802, N2894);
or OR2 (N5179, N5175, N1780);
nor NOR4 (N5180, N5179, N21, N3645, N3599);
nor NOR3 (N5181, N5178, N4245, N2003);
or OR2 (N5182, N5157, N3180);
nor NOR4 (N5183, N5153, N2922, N4489, N3329);
and AND4 (N5184, N5159, N3347, N4277, N351);
buf BUF1 (N5185, N5180);
or OR2 (N5186, N5165, N2870);
nand NAND3 (N5187, N5186, N63, N429);
xor XOR2 (N5188, N5168, N2530);
buf BUF1 (N5189, N5182);
nand NAND4 (N5190, N5177, N4892, N2396, N721);
nor NOR3 (N5191, N5170, N2098, N3833);
not NOT1 (N5192, N5160);
nor NOR2 (N5193, N5184, N1029);
xor XOR2 (N5194, N5190, N4976);
or OR2 (N5195, N5187, N854);
or OR2 (N5196, N5185, N428);
buf BUF1 (N5197, N5188);
not NOT1 (N5198, N5189);
nand NAND2 (N5199, N5198, N2334);
or OR4 (N5200, N5192, N1656, N1099, N2601);
or OR2 (N5201, N5191, N3150);
not NOT1 (N5202, N5197);
not NOT1 (N5203, N5199);
buf BUF1 (N5204, N5194);
buf BUF1 (N5205, N5196);
nor NOR2 (N5206, N5200, N502);
and AND4 (N5207, N5195, N3307, N505, N3765);
nand NAND3 (N5208, N5183, N560, N1084);
or OR4 (N5209, N5206, N1628, N846, N4173);
xor XOR2 (N5210, N5202, N3725);
or OR2 (N5211, N5210, N1604);
xor XOR2 (N5212, N5209, N2551);
xor XOR2 (N5213, N5181, N2830);
buf BUF1 (N5214, N5213);
nand NAND2 (N5215, N5205, N2837);
nor NOR2 (N5216, N5193, N3225);
and AND2 (N5217, N5207, N5092);
nand NAND4 (N5218, N5216, N1981, N3774, N3386);
buf BUF1 (N5219, N5208);
nand NAND3 (N5220, N5203, N3000, N2829);
nand NAND3 (N5221, N5215, N2771, N1506);
and AND2 (N5222, N5219, N3104);
and AND3 (N5223, N5218, N4775, N3237);
nor NOR2 (N5224, N5221, N2029);
and AND2 (N5225, N5224, N937);
not NOT1 (N5226, N5220);
buf BUF1 (N5227, N5222);
nand NAND4 (N5228, N5226, N4683, N452, N3140);
buf BUF1 (N5229, N5204);
and AND3 (N5230, N5212, N1937, N2969);
and AND2 (N5231, N5227, N1600);
xor XOR2 (N5232, N5223, N701);
not NOT1 (N5233, N5201);
buf BUF1 (N5234, N5229);
nand NAND2 (N5235, N5211, N828);
and AND3 (N5236, N5228, N2742, N2732);
not NOT1 (N5237, N5233);
buf BUF1 (N5238, N5231);
not NOT1 (N5239, N5232);
and AND4 (N5240, N5238, N1038, N4964, N2914);
and AND3 (N5241, N5239, N2691, N3954);
or OR2 (N5242, N5225, N237);
or OR3 (N5243, N5234, N3870, N4686);
nor NOR2 (N5244, N5242, N247);
not NOT1 (N5245, N5237);
buf BUF1 (N5246, N5241);
or OR2 (N5247, N5230, N3782);
xor XOR2 (N5248, N5246, N3797);
and AND2 (N5249, N5243, N832);
and AND3 (N5250, N5244, N2115, N712);
buf BUF1 (N5251, N5250);
nand NAND2 (N5252, N5235, N974);
xor XOR2 (N5253, N5240, N1676);
and AND4 (N5254, N5253, N4790, N5232, N2378);
or OR4 (N5255, N5254, N5213, N783, N3803);
not NOT1 (N5256, N5249);
nand NAND3 (N5257, N5214, N4513, N1763);
xor XOR2 (N5258, N5252, N375);
xor XOR2 (N5259, N5251, N2994);
and AND3 (N5260, N5258, N2818, N682);
xor XOR2 (N5261, N5255, N2590);
or OR4 (N5262, N5260, N1743, N153, N3247);
and AND4 (N5263, N5259, N2822, N3233, N664);
and AND2 (N5264, N5247, N3976);
or OR3 (N5265, N5264, N6, N4449);
or OR4 (N5266, N5263, N114, N1458, N1448);
or OR3 (N5267, N5217, N225, N613);
not NOT1 (N5268, N5262);
buf BUF1 (N5269, N5245);
or OR4 (N5270, N5256, N4075, N759, N881);
buf BUF1 (N5271, N5268);
xor XOR2 (N5272, N5266, N4662);
and AND3 (N5273, N5271, N4318, N995);
xor XOR2 (N5274, N5273, N1213);
nand NAND2 (N5275, N5265, N1275);
nand NAND4 (N5276, N5272, N5253, N2479, N3447);
and AND2 (N5277, N5270, N148);
and AND3 (N5278, N5275, N563, N2930);
nor NOR2 (N5279, N5257, N4293);
or OR3 (N5280, N5277, N2104, N2880);
or OR4 (N5281, N5278, N3563, N3840, N1417);
nor NOR2 (N5282, N5279, N1767);
not NOT1 (N5283, N5261);
nand NAND2 (N5284, N5283, N4279);
and AND3 (N5285, N5276, N3660, N441);
not NOT1 (N5286, N5281);
nor NOR2 (N5287, N5267, N43);
xor XOR2 (N5288, N5282, N187);
not NOT1 (N5289, N5236);
or OR3 (N5290, N5288, N2741, N18);
not NOT1 (N5291, N5287);
not NOT1 (N5292, N5280);
nor NOR3 (N5293, N5274, N3790, N3343);
buf BUF1 (N5294, N5286);
nand NAND3 (N5295, N5269, N1598, N3802);
not NOT1 (N5296, N5294);
and AND4 (N5297, N5291, N4807, N8, N2781);
nor NOR4 (N5298, N5295, N3234, N4347, N5198);
xor XOR2 (N5299, N5297, N157);
nand NAND3 (N5300, N5299, N4239, N314);
buf BUF1 (N5301, N5285);
or OR4 (N5302, N5289, N4024, N5266, N4379);
xor XOR2 (N5303, N5284, N3884);
not NOT1 (N5304, N5303);
nor NOR3 (N5305, N5301, N4302, N2296);
not NOT1 (N5306, N5293);
nor NOR3 (N5307, N5300, N937, N1862);
xor XOR2 (N5308, N5292, N1598);
nor NOR2 (N5309, N5296, N4636);
xor XOR2 (N5310, N5290, N238);
xor XOR2 (N5311, N5306, N3293);
and AND2 (N5312, N5308, N4514);
nand NAND3 (N5313, N5302, N2710, N4534);
buf BUF1 (N5314, N5304);
xor XOR2 (N5315, N5248, N1978);
nand NAND4 (N5316, N5312, N2224, N2310, N928);
buf BUF1 (N5317, N5313);
not NOT1 (N5318, N5307);
nor NOR4 (N5319, N5316, N1232, N5282, N3486);
or OR3 (N5320, N5315, N2617, N4425);
buf BUF1 (N5321, N5310);
or OR4 (N5322, N5311, N340, N2427, N5219);
nor NOR4 (N5323, N5322, N3762, N3102, N1419);
nor NOR4 (N5324, N5323, N980, N199, N45);
nand NAND2 (N5325, N5314, N3557);
xor XOR2 (N5326, N5325, N3813);
not NOT1 (N5327, N5305);
xor XOR2 (N5328, N5298, N263);
buf BUF1 (N5329, N5318);
not NOT1 (N5330, N5324);
or OR4 (N5331, N5320, N5003, N2879, N418);
buf BUF1 (N5332, N5321);
nand NAND3 (N5333, N5328, N5304, N2269);
nand NAND3 (N5334, N5317, N312, N1083);
not NOT1 (N5335, N5330);
xor XOR2 (N5336, N5333, N3275);
not NOT1 (N5337, N5329);
nor NOR4 (N5338, N5309, N2688, N2394, N4919);
nand NAND3 (N5339, N5327, N2048, N3895);
or OR4 (N5340, N5334, N3269, N4885, N3249);
xor XOR2 (N5341, N5337, N144);
and AND3 (N5342, N5326, N3700, N182);
buf BUF1 (N5343, N5319);
xor XOR2 (N5344, N5332, N3732);
xor XOR2 (N5345, N5331, N1397);
not NOT1 (N5346, N5340);
nor NOR4 (N5347, N5343, N4723, N2268, N2354);
not NOT1 (N5348, N5347);
not NOT1 (N5349, N5335);
xor XOR2 (N5350, N5348, N287);
nor NOR4 (N5351, N5350, N1879, N1593, N4863);
and AND3 (N5352, N5346, N1607, N1989);
xor XOR2 (N5353, N5339, N595);
nor NOR4 (N5354, N5353, N1358, N4834, N3809);
or OR2 (N5355, N5338, N1144);
xor XOR2 (N5356, N5341, N1208);
buf BUF1 (N5357, N5352);
xor XOR2 (N5358, N5344, N1384);
nand NAND4 (N5359, N5336, N4589, N842, N598);
or OR2 (N5360, N5349, N4895);
xor XOR2 (N5361, N5359, N3858);
buf BUF1 (N5362, N5361);
not NOT1 (N5363, N5362);
nand NAND4 (N5364, N5360, N2428, N2396, N941);
not NOT1 (N5365, N5363);
or OR3 (N5366, N5365, N5352, N709);
or OR3 (N5367, N5345, N3970, N5342);
or OR2 (N5368, N1936, N1898);
not NOT1 (N5369, N5356);
xor XOR2 (N5370, N5357, N4668);
not NOT1 (N5371, N5366);
not NOT1 (N5372, N5369);
xor XOR2 (N5373, N5351, N4427);
not NOT1 (N5374, N5355);
not NOT1 (N5375, N5354);
or OR2 (N5376, N5368, N2163);
not NOT1 (N5377, N5358);
not NOT1 (N5378, N5370);
not NOT1 (N5379, N5371);
and AND4 (N5380, N5367, N666, N2538, N2447);
nand NAND2 (N5381, N5372, N1517);
and AND4 (N5382, N5380, N2244, N4453, N3946);
nor NOR4 (N5383, N5376, N4754, N1867, N3033);
nand NAND2 (N5384, N5378, N3762);
nor NOR3 (N5385, N5374, N595, N4360);
not NOT1 (N5386, N5384);
not NOT1 (N5387, N5386);
buf BUF1 (N5388, N5385);
nor NOR4 (N5389, N5381, N703, N4204, N5291);
not NOT1 (N5390, N5373);
buf BUF1 (N5391, N5390);
buf BUF1 (N5392, N5364);
buf BUF1 (N5393, N5377);
xor XOR2 (N5394, N5388, N4859);
buf BUF1 (N5395, N5394);
xor XOR2 (N5396, N5393, N624);
nand NAND3 (N5397, N5382, N1954, N1709);
buf BUF1 (N5398, N5396);
nand NAND2 (N5399, N5375, N1532);
not NOT1 (N5400, N5399);
or OR2 (N5401, N5383, N3447);
or OR3 (N5402, N5398, N4290, N3717);
buf BUF1 (N5403, N5391);
and AND4 (N5404, N5379, N205, N2023, N2330);
or OR2 (N5405, N5400, N1916);
xor XOR2 (N5406, N5387, N3551);
xor XOR2 (N5407, N5395, N633);
xor XOR2 (N5408, N5403, N232);
and AND2 (N5409, N5402, N4829);
nor NOR2 (N5410, N5405, N3960);
buf BUF1 (N5411, N5407);
buf BUF1 (N5412, N5389);
and AND2 (N5413, N5397, N5148);
not NOT1 (N5414, N5412);
nand NAND3 (N5415, N5408, N5093, N1434);
buf BUF1 (N5416, N5406);
and AND4 (N5417, N5401, N43, N342, N793);
not NOT1 (N5418, N5411);
nor NOR2 (N5419, N5409, N2260);
buf BUF1 (N5420, N5413);
and AND4 (N5421, N5416, N694, N173, N3360);
or OR4 (N5422, N5415, N4661, N1838, N128);
xor XOR2 (N5423, N5417, N1075);
xor XOR2 (N5424, N5404, N4627);
or OR3 (N5425, N5414, N3760, N2939);
nor NOR3 (N5426, N5422, N4025, N2894);
buf BUF1 (N5427, N5392);
not NOT1 (N5428, N5423);
nor NOR3 (N5429, N5419, N5371, N2011);
xor XOR2 (N5430, N5410, N2314);
not NOT1 (N5431, N5418);
not NOT1 (N5432, N5420);
nand NAND3 (N5433, N5429, N1292, N1508);
xor XOR2 (N5434, N5432, N1837);
nor NOR2 (N5435, N5426, N4039);
buf BUF1 (N5436, N5428);
or OR2 (N5437, N5433, N232);
and AND4 (N5438, N5421, N1652, N486, N835);
or OR3 (N5439, N5425, N1971, N5158);
nand NAND3 (N5440, N5438, N1170, N3241);
and AND2 (N5441, N5436, N2885);
buf BUF1 (N5442, N5440);
xor XOR2 (N5443, N5442, N4826);
nor NOR4 (N5444, N5435, N3718, N4481, N4341);
not NOT1 (N5445, N5434);
buf BUF1 (N5446, N5443);
xor XOR2 (N5447, N5431, N2050);
nor NOR3 (N5448, N5437, N3817, N4190);
not NOT1 (N5449, N5441);
and AND2 (N5450, N5447, N2014);
nor NOR2 (N5451, N5448, N1333);
and AND2 (N5452, N5430, N557);
and AND2 (N5453, N5427, N688);
nand NAND4 (N5454, N5451, N2129, N1123, N3775);
or OR3 (N5455, N5449, N2494, N1132);
nor NOR3 (N5456, N5446, N3594, N1587);
buf BUF1 (N5457, N5455);
and AND3 (N5458, N5444, N4487, N3638);
or OR3 (N5459, N5458, N290, N3838);
xor XOR2 (N5460, N5457, N4807);
or OR3 (N5461, N5452, N5233, N3874);
and AND4 (N5462, N5456, N1279, N1396, N937);
nand NAND2 (N5463, N5461, N4106);
xor XOR2 (N5464, N5424, N330);
not NOT1 (N5465, N5460);
and AND2 (N5466, N5462, N5307);
nor NOR3 (N5467, N5450, N4680, N2543);
nor NOR4 (N5468, N5466, N4357, N2901, N4033);
or OR2 (N5469, N5467, N1686);
or OR2 (N5470, N5464, N2708);
nand NAND4 (N5471, N5463, N349, N3213, N1518);
or OR2 (N5472, N5471, N516);
nor NOR2 (N5473, N5469, N3665);
or OR2 (N5474, N5472, N2057);
buf BUF1 (N5475, N5470);
not NOT1 (N5476, N5474);
not NOT1 (N5477, N5476);
not NOT1 (N5478, N5468);
not NOT1 (N5479, N5459);
nand NAND4 (N5480, N5453, N2033, N2646, N5411);
nor NOR4 (N5481, N5465, N1653, N5304, N3842);
or OR3 (N5482, N5473, N5183, N1824);
nor NOR4 (N5483, N5480, N4935, N1264, N3494);
not NOT1 (N5484, N5482);
not NOT1 (N5485, N5445);
xor XOR2 (N5486, N5485, N2254);
xor XOR2 (N5487, N5484, N2934);
nor NOR2 (N5488, N5477, N1628);
not NOT1 (N5489, N5483);
nor NOR4 (N5490, N5479, N3568, N4453, N34);
and AND3 (N5491, N5490, N2527, N4071);
xor XOR2 (N5492, N5454, N5481);
buf BUF1 (N5493, N1938);
xor XOR2 (N5494, N5475, N5022);
not NOT1 (N5495, N5439);
and AND2 (N5496, N5486, N4050);
nor NOR3 (N5497, N5478, N2456, N3950);
and AND4 (N5498, N5487, N5325, N3318, N5275);
nor NOR2 (N5499, N5497, N1091);
nand NAND4 (N5500, N5488, N1668, N3576, N1955);
buf BUF1 (N5501, N5495);
xor XOR2 (N5502, N5501, N2637);
or OR2 (N5503, N5489, N5148);
and AND3 (N5504, N5502, N1252, N1);
nor NOR3 (N5505, N5503, N3228, N63);
or OR3 (N5506, N5494, N4125, N493);
buf BUF1 (N5507, N5493);
buf BUF1 (N5508, N5507);
xor XOR2 (N5509, N5498, N2294);
buf BUF1 (N5510, N5500);
nor NOR2 (N5511, N5506, N3677);
not NOT1 (N5512, N5492);
nand NAND2 (N5513, N5505, N3672);
nor NOR2 (N5514, N5499, N621);
nand NAND3 (N5515, N5513, N543, N4681);
not NOT1 (N5516, N5514);
buf BUF1 (N5517, N5496);
nor NOR4 (N5518, N5504, N2670, N565, N2597);
buf BUF1 (N5519, N5510);
buf BUF1 (N5520, N5517);
not NOT1 (N5521, N5519);
xor XOR2 (N5522, N5491, N2833);
xor XOR2 (N5523, N5515, N3314);
not NOT1 (N5524, N5523);
and AND2 (N5525, N5516, N607);
or OR3 (N5526, N5520, N3340, N4352);
xor XOR2 (N5527, N5525, N5216);
not NOT1 (N5528, N5521);
xor XOR2 (N5529, N5526, N642);
nand NAND2 (N5530, N5527, N151);
buf BUF1 (N5531, N5528);
xor XOR2 (N5532, N5529, N890);
buf BUF1 (N5533, N5524);
or OR2 (N5534, N5532, N4734);
buf BUF1 (N5535, N5518);
not NOT1 (N5536, N5522);
buf BUF1 (N5537, N5534);
buf BUF1 (N5538, N5537);
and AND4 (N5539, N5512, N4435, N1573, N1633);
and AND4 (N5540, N5531, N3379, N4576, N3218);
xor XOR2 (N5541, N5533, N162);
or OR4 (N5542, N5539, N4924, N2201, N4116);
buf BUF1 (N5543, N5508);
nor NOR2 (N5544, N5540, N3196);
nand NAND3 (N5545, N5535, N1607, N3650);
and AND2 (N5546, N5544, N799);
nand NAND2 (N5547, N5546, N2807);
nor NOR3 (N5548, N5511, N2059, N1097);
nor NOR3 (N5549, N5538, N2078, N1312);
or OR2 (N5550, N5548, N4487);
nand NAND4 (N5551, N5550, N655, N2390, N211);
and AND2 (N5552, N5541, N4727);
and AND3 (N5553, N5547, N4714, N4106);
and AND3 (N5554, N5542, N1598, N3747);
and AND4 (N5555, N5549, N186, N2770, N1978);
and AND4 (N5556, N5552, N2765, N4506, N987);
or OR4 (N5557, N5530, N812, N4268, N903);
and AND3 (N5558, N5554, N2311, N3341);
and AND2 (N5559, N5545, N1455);
not NOT1 (N5560, N5509);
and AND3 (N5561, N5559, N1999, N3386);
buf BUF1 (N5562, N5553);
or OR2 (N5563, N5536, N851);
xor XOR2 (N5564, N5558, N1104);
nand NAND3 (N5565, N5564, N3056, N1891);
or OR2 (N5566, N5556, N1345);
nor NOR4 (N5567, N5560, N2991, N3522, N758);
not NOT1 (N5568, N5557);
and AND2 (N5569, N5555, N1213);
or OR2 (N5570, N5567, N772);
xor XOR2 (N5571, N5543, N3487);
or OR2 (N5572, N5561, N1181);
and AND3 (N5573, N5571, N2798, N4252);
nor NOR2 (N5574, N5551, N2921);
buf BUF1 (N5575, N5570);
not NOT1 (N5576, N5563);
and AND2 (N5577, N5574, N4948);
and AND3 (N5578, N5576, N4390, N2854);
and AND3 (N5579, N5575, N4680, N3202);
and AND4 (N5580, N5568, N2928, N240, N5385);
not NOT1 (N5581, N5565);
buf BUF1 (N5582, N5569);
nand NAND3 (N5583, N5581, N2303, N3892);
or OR4 (N5584, N5582, N820, N3063, N2198);
buf BUF1 (N5585, N5579);
buf BUF1 (N5586, N5583);
buf BUF1 (N5587, N5572);
nand NAND4 (N5588, N5587, N39, N2581, N3888);
not NOT1 (N5589, N5566);
and AND2 (N5590, N5585, N3490);
xor XOR2 (N5591, N5573, N4730);
xor XOR2 (N5592, N5580, N3509);
xor XOR2 (N5593, N5578, N364);
not NOT1 (N5594, N5588);
not NOT1 (N5595, N5589);
not NOT1 (N5596, N5590);
not NOT1 (N5597, N5594);
or OR2 (N5598, N5597, N3119);
and AND3 (N5599, N5598, N3882, N5541);
and AND2 (N5600, N5584, N1138);
not NOT1 (N5601, N5591);
xor XOR2 (N5602, N5592, N2200);
or OR2 (N5603, N5596, N4319);
buf BUF1 (N5604, N5599);
nor NOR3 (N5605, N5600, N4132, N3499);
buf BUF1 (N5606, N5595);
buf BUF1 (N5607, N5603);
buf BUF1 (N5608, N5607);
nor NOR2 (N5609, N5608, N5035);
xor XOR2 (N5610, N5586, N5422);
nand NAND4 (N5611, N5604, N1689, N4633, N4515);
or OR3 (N5612, N5611, N4558, N3816);
xor XOR2 (N5613, N5610, N3514);
xor XOR2 (N5614, N5605, N4844);
or OR3 (N5615, N5614, N1581, N2750);
nand NAND3 (N5616, N5615, N4446, N79);
or OR4 (N5617, N5577, N3344, N3365, N5289);
nand NAND3 (N5618, N5616, N3097, N3102);
and AND2 (N5619, N5606, N364);
nor NOR2 (N5620, N5601, N623);
buf BUF1 (N5621, N5619);
not NOT1 (N5622, N5618);
buf BUF1 (N5623, N5613);
not NOT1 (N5624, N5621);
buf BUF1 (N5625, N5617);
buf BUF1 (N5626, N5612);
and AND4 (N5627, N5602, N1556, N3582, N3156);
nand NAND2 (N5628, N5625, N4478);
nor NOR3 (N5629, N5622, N72, N4070);
nor NOR4 (N5630, N5627, N130, N8, N5151);
not NOT1 (N5631, N5626);
nor NOR2 (N5632, N5631, N2655);
xor XOR2 (N5633, N5628, N3348);
and AND2 (N5634, N5562, N64);
or OR4 (N5635, N5633, N2473, N5624, N2047);
buf BUF1 (N5636, N778);
xor XOR2 (N5637, N5630, N2075);
not NOT1 (N5638, N5636);
nand NAND4 (N5639, N5637, N296, N3591, N3295);
nor NOR2 (N5640, N5634, N1135);
or OR4 (N5641, N5639, N5439, N3374, N1372);
or OR3 (N5642, N5632, N989, N5225);
nor NOR3 (N5643, N5620, N3453, N3586);
xor XOR2 (N5644, N5635, N2335);
nand NAND2 (N5645, N5640, N588);
or OR2 (N5646, N5629, N1307);
nor NOR4 (N5647, N5644, N3090, N519, N1809);
buf BUF1 (N5648, N5646);
nand NAND4 (N5649, N5647, N3840, N4393, N5344);
nor NOR2 (N5650, N5643, N499);
and AND2 (N5651, N5650, N5367);
and AND2 (N5652, N5648, N842);
buf BUF1 (N5653, N5593);
nand NAND2 (N5654, N5651, N4616);
and AND3 (N5655, N5638, N2924, N3125);
nor NOR3 (N5656, N5649, N2498, N3429);
nor NOR2 (N5657, N5623, N1272);
nor NOR3 (N5658, N5645, N5444, N1316);
xor XOR2 (N5659, N5653, N618);
nand NAND3 (N5660, N5659, N1154, N4974);
nand NAND3 (N5661, N5652, N722, N206);
or OR2 (N5662, N5656, N1784);
or OR4 (N5663, N5654, N4128, N930, N4475);
buf BUF1 (N5664, N5641);
or OR4 (N5665, N5660, N460, N2981, N2410);
or OR4 (N5666, N5663, N1769, N1648, N5121);
not NOT1 (N5667, N5609);
and AND4 (N5668, N5661, N3881, N2046, N1330);
nand NAND4 (N5669, N5666, N3454, N4740, N3170);
and AND4 (N5670, N5642, N2657, N1250, N5387);
or OR3 (N5671, N5664, N1469, N3462);
xor XOR2 (N5672, N5669, N3689);
buf BUF1 (N5673, N5662);
not NOT1 (N5674, N5657);
buf BUF1 (N5675, N5658);
nor NOR4 (N5676, N5667, N5450, N1214, N230);
buf BUF1 (N5677, N5655);
xor XOR2 (N5678, N5677, N1411);
nor NOR2 (N5679, N5673, N4815);
nor NOR2 (N5680, N5676, N2228);
buf BUF1 (N5681, N5675);
buf BUF1 (N5682, N5681);
buf BUF1 (N5683, N5670);
buf BUF1 (N5684, N5679);
nand NAND4 (N5685, N5668, N2620, N3093, N4806);
or OR2 (N5686, N5672, N5282);
and AND4 (N5687, N5665, N2457, N310, N3602);
buf BUF1 (N5688, N5685);
xor XOR2 (N5689, N5680, N4423);
or OR2 (N5690, N5678, N4299);
nand NAND4 (N5691, N5688, N4059, N2285, N2135);
nand NAND4 (N5692, N5671, N408, N4393, N5198);
nand NAND4 (N5693, N5686, N3026, N2864, N4351);
nand NAND3 (N5694, N5683, N2002, N4476);
not NOT1 (N5695, N5691);
nor NOR2 (N5696, N5674, N129);
nand NAND3 (N5697, N5692, N3731, N1198);
buf BUF1 (N5698, N5693);
or OR3 (N5699, N5684, N1536, N2848);
and AND3 (N5700, N5687, N1791, N5179);
buf BUF1 (N5701, N5697);
or OR3 (N5702, N5698, N983, N5653);
nor NOR4 (N5703, N5699, N1136, N4017, N4909);
and AND4 (N5704, N5701, N3041, N2232, N2463);
not NOT1 (N5705, N5700);
and AND3 (N5706, N5702, N148, N1014);
and AND4 (N5707, N5706, N3047, N4630, N5563);
not NOT1 (N5708, N5704);
buf BUF1 (N5709, N5707);
and AND3 (N5710, N5689, N2840, N2891);
not NOT1 (N5711, N5696);
and AND2 (N5712, N5710, N333);
or OR2 (N5713, N5703, N4774);
nor NOR4 (N5714, N5705, N2172, N453, N264);
or OR2 (N5715, N5690, N155);
not NOT1 (N5716, N5714);
nor NOR2 (N5717, N5709, N3298);
xor XOR2 (N5718, N5682, N3495);
buf BUF1 (N5719, N5695);
xor XOR2 (N5720, N5718, N4664);
xor XOR2 (N5721, N5712, N2230);
and AND2 (N5722, N5721, N70);
not NOT1 (N5723, N5719);
or OR4 (N5724, N5716, N4945, N4737, N3898);
xor XOR2 (N5725, N5715, N2960);
not NOT1 (N5726, N5694);
and AND2 (N5727, N5724, N5539);
and AND3 (N5728, N5717, N504, N4697);
or OR4 (N5729, N5723, N3302, N4679, N260);
xor XOR2 (N5730, N5720, N3823);
buf BUF1 (N5731, N5725);
xor XOR2 (N5732, N5722, N868);
or OR4 (N5733, N5732, N2470, N3594, N1024);
and AND4 (N5734, N5708, N3608, N3556, N3479);
xor XOR2 (N5735, N5713, N1583);
nand NAND2 (N5736, N5728, N4348);
not NOT1 (N5737, N5731);
nor NOR2 (N5738, N5729, N5260);
and AND2 (N5739, N5736, N3879);
xor XOR2 (N5740, N5734, N2052);
nor NOR3 (N5741, N5735, N5253, N5302);
xor XOR2 (N5742, N5737, N2999);
or OR2 (N5743, N5733, N5495);
and AND4 (N5744, N5740, N400, N2214, N4164);
nand NAND2 (N5745, N5739, N2513);
xor XOR2 (N5746, N5742, N1683);
and AND2 (N5747, N5738, N4558);
nor NOR4 (N5748, N5747, N1762, N2340, N1419);
or OR2 (N5749, N5727, N2570);
nor NOR3 (N5750, N5749, N1212, N3012);
not NOT1 (N5751, N5750);
nor NOR3 (N5752, N5744, N2763, N5473);
nand NAND2 (N5753, N5751, N2979);
nand NAND4 (N5754, N5726, N303, N4189, N3148);
nand NAND4 (N5755, N5741, N3198, N2167, N3011);
not NOT1 (N5756, N5743);
not NOT1 (N5757, N5752);
not NOT1 (N5758, N5748);
and AND3 (N5759, N5745, N620, N1161);
xor XOR2 (N5760, N5755, N4541);
not NOT1 (N5761, N5758);
buf BUF1 (N5762, N5759);
buf BUF1 (N5763, N5754);
nor NOR2 (N5764, N5760, N599);
not NOT1 (N5765, N5756);
nor NOR3 (N5766, N5765, N5224, N4451);
and AND4 (N5767, N5757, N557, N2170, N1629);
nand NAND2 (N5768, N5762, N856);
buf BUF1 (N5769, N5766);
xor XOR2 (N5770, N5768, N5269);
xor XOR2 (N5771, N5711, N1861);
not NOT1 (N5772, N5767);
not NOT1 (N5773, N5764);
nand NAND3 (N5774, N5773, N1110, N4715);
xor XOR2 (N5775, N5753, N4518);
xor XOR2 (N5776, N5774, N3454);
buf BUF1 (N5777, N5771);
nand NAND4 (N5778, N5770, N3161, N4685, N3165);
or OR2 (N5779, N5763, N2699);
buf BUF1 (N5780, N5769);
xor XOR2 (N5781, N5772, N2788);
and AND2 (N5782, N5780, N3000);
not NOT1 (N5783, N5761);
not NOT1 (N5784, N5777);
and AND3 (N5785, N5782, N2849, N4691);
nor NOR4 (N5786, N5746, N3261, N3430, N2618);
not NOT1 (N5787, N5781);
nor NOR2 (N5788, N5786, N4086);
or OR2 (N5789, N5778, N5303);
or OR3 (N5790, N5784, N378, N5530);
nor NOR3 (N5791, N5730, N890, N1454);
nand NAND2 (N5792, N5785, N1734);
not NOT1 (N5793, N5788);
and AND4 (N5794, N5776, N1901, N5147, N4981);
not NOT1 (N5795, N5793);
nor NOR4 (N5796, N5791, N3604, N4847, N961);
nand NAND2 (N5797, N5792, N1283);
nor NOR4 (N5798, N5796, N2102, N500, N4992);
not NOT1 (N5799, N5787);
and AND2 (N5800, N5775, N5743);
or OR3 (N5801, N5799, N3871, N4832);
not NOT1 (N5802, N5789);
nand NAND3 (N5803, N5797, N621, N3915);
buf BUF1 (N5804, N5783);
and AND4 (N5805, N5804, N4466, N2883, N5561);
not NOT1 (N5806, N5805);
xor XOR2 (N5807, N5795, N2403);
xor XOR2 (N5808, N5803, N38);
nor NOR2 (N5809, N5798, N2820);
buf BUF1 (N5810, N5808);
xor XOR2 (N5811, N5810, N4702);
or OR4 (N5812, N5790, N5736, N237, N5718);
nand NAND3 (N5813, N5800, N1346, N182);
not NOT1 (N5814, N5801);
nand NAND4 (N5815, N5794, N3708, N2041, N246);
nand NAND3 (N5816, N5813, N1741, N1137);
not NOT1 (N5817, N5802);
not NOT1 (N5818, N5806);
buf BUF1 (N5819, N5818);
nor NOR3 (N5820, N5779, N4574, N1111);
and AND4 (N5821, N5812, N4297, N3676, N2973);
buf BUF1 (N5822, N5815);
nand NAND4 (N5823, N5820, N954, N4600, N3982);
nand NAND2 (N5824, N5809, N1046);
nand NAND4 (N5825, N5824, N513, N1347, N4198);
xor XOR2 (N5826, N5822, N5060);
nand NAND3 (N5827, N5811, N3359, N2683);
nand NAND4 (N5828, N5807, N3900, N5422, N2407);
not NOT1 (N5829, N5827);
and AND3 (N5830, N5816, N4549, N2728);
not NOT1 (N5831, N5825);
nor NOR4 (N5832, N5830, N5575, N2515, N3669);
nor NOR2 (N5833, N5829, N4759);
not NOT1 (N5834, N5814);
not NOT1 (N5835, N5819);
not NOT1 (N5836, N5823);
xor XOR2 (N5837, N5834, N2877);
or OR4 (N5838, N5836, N2562, N1016, N4190);
nand NAND3 (N5839, N5835, N2343, N77);
nor NOR3 (N5840, N5828, N434, N4898);
and AND4 (N5841, N5840, N4687, N934, N5741);
not NOT1 (N5842, N5826);
and AND2 (N5843, N5838, N5373);
nor NOR4 (N5844, N5833, N2989, N716, N2645);
buf BUF1 (N5845, N5843);
buf BUF1 (N5846, N5817);
and AND4 (N5847, N5832, N1416, N3928, N639);
or OR4 (N5848, N5847, N762, N1290, N3527);
buf BUF1 (N5849, N5842);
xor XOR2 (N5850, N5821, N3515);
nor NOR2 (N5851, N5844, N4610);
nor NOR3 (N5852, N5837, N418, N5012);
and AND4 (N5853, N5848, N2305, N5684, N215);
nand NAND2 (N5854, N5839, N2972);
buf BUF1 (N5855, N5850);
and AND4 (N5856, N5854, N2459, N4683, N594);
nand NAND4 (N5857, N5852, N2749, N2887, N4250);
nor NOR3 (N5858, N5851, N2079, N3938);
xor XOR2 (N5859, N5841, N1762);
not NOT1 (N5860, N5845);
not NOT1 (N5861, N5849);
and AND4 (N5862, N5858, N99, N4148, N798);
and AND2 (N5863, N5861, N3704);
nor NOR2 (N5864, N5862, N4042);
and AND3 (N5865, N5863, N2012, N1677);
or OR3 (N5866, N5860, N2296, N4587);
nand NAND2 (N5867, N5859, N1025);
not NOT1 (N5868, N5846);
and AND2 (N5869, N5866, N3829);
nand NAND2 (N5870, N5853, N5404);
xor XOR2 (N5871, N5869, N4041);
and AND3 (N5872, N5864, N5142, N2680);
nand NAND4 (N5873, N5831, N5506, N524, N3537);
not NOT1 (N5874, N5872);
nor NOR2 (N5875, N5870, N667);
and AND3 (N5876, N5867, N1390, N2285);
buf BUF1 (N5877, N5876);
xor XOR2 (N5878, N5873, N4268);
not NOT1 (N5879, N5877);
nand NAND3 (N5880, N5878, N1059, N5010);
buf BUF1 (N5881, N5856);
xor XOR2 (N5882, N5857, N3235);
buf BUF1 (N5883, N5855);
buf BUF1 (N5884, N5879);
nor NOR2 (N5885, N5874, N1957);
buf BUF1 (N5886, N5868);
or OR3 (N5887, N5865, N2249, N2943);
nand NAND2 (N5888, N5882, N2883);
not NOT1 (N5889, N5885);
not NOT1 (N5890, N5881);
and AND4 (N5891, N5880, N70, N105, N48);
nor NOR4 (N5892, N5889, N1071, N4327, N5017);
nor NOR4 (N5893, N5884, N5754, N2222, N4569);
not NOT1 (N5894, N5875);
buf BUF1 (N5895, N5892);
buf BUF1 (N5896, N5883);
nor NOR2 (N5897, N5886, N4617);
buf BUF1 (N5898, N5871);
not NOT1 (N5899, N5895);
and AND3 (N5900, N5887, N24, N5209);
not NOT1 (N5901, N5891);
nor NOR2 (N5902, N5900, N297);
buf BUF1 (N5903, N5893);
buf BUF1 (N5904, N5902);
xor XOR2 (N5905, N5894, N218);
xor XOR2 (N5906, N5890, N969);
or OR4 (N5907, N5906, N4673, N377, N4024);
or OR4 (N5908, N5905, N3101, N1768, N952);
buf BUF1 (N5909, N5904);
or OR2 (N5910, N5897, N3790);
or OR4 (N5911, N5909, N251, N1591, N2398);
and AND4 (N5912, N5907, N1359, N4978, N4052);
and AND4 (N5913, N5912, N2363, N4484, N2814);
and AND3 (N5914, N5908, N5104, N5153);
nand NAND3 (N5915, N5899, N759, N5373);
buf BUF1 (N5916, N5898);
and AND3 (N5917, N5901, N265, N3964);
buf BUF1 (N5918, N5913);
or OR3 (N5919, N5888, N5646, N3093);
nor NOR4 (N5920, N5903, N3764, N3976, N3136);
nor NOR3 (N5921, N5919, N3192, N1417);
buf BUF1 (N5922, N5914);
nor NOR3 (N5923, N5916, N3195, N5602);
not NOT1 (N5924, N5910);
and AND3 (N5925, N5896, N4932, N5434);
and AND4 (N5926, N5911, N3328, N2480, N4126);
or OR2 (N5927, N5921, N1796);
not NOT1 (N5928, N5920);
not NOT1 (N5929, N5922);
not NOT1 (N5930, N5928);
not NOT1 (N5931, N5930);
nor NOR2 (N5932, N5917, N1577);
not NOT1 (N5933, N5931);
not NOT1 (N5934, N5923);
nor NOR2 (N5935, N5924, N1978);
nor NOR3 (N5936, N5926, N3765, N3052);
nand NAND4 (N5937, N5935, N1238, N2666, N125);
buf BUF1 (N5938, N5937);
nand NAND2 (N5939, N5934, N2499);
or OR2 (N5940, N5925, N1501);
not NOT1 (N5941, N5918);
and AND4 (N5942, N5938, N630, N987, N2391);
not NOT1 (N5943, N5929);
or OR4 (N5944, N5915, N2287, N5229, N550);
xor XOR2 (N5945, N5933, N690);
buf BUF1 (N5946, N5942);
and AND4 (N5947, N5945, N534, N3436, N1234);
and AND2 (N5948, N5943, N2004);
nor NOR4 (N5949, N5927, N1560, N5274, N1467);
or OR2 (N5950, N5948, N5434);
not NOT1 (N5951, N5936);
nor NOR4 (N5952, N5941, N171, N4025, N5566);
not NOT1 (N5953, N5949);
xor XOR2 (N5954, N5944, N1391);
and AND4 (N5955, N5953, N254, N1210, N3077);
nor NOR3 (N5956, N5952, N303, N1720);
not NOT1 (N5957, N5955);
nand NAND3 (N5958, N5957, N5532, N125);
xor XOR2 (N5959, N5947, N1521);
xor XOR2 (N5960, N5959, N3778);
buf BUF1 (N5961, N5940);
or OR2 (N5962, N5958, N5887);
xor XOR2 (N5963, N5950, N5205);
nor NOR2 (N5964, N5962, N988);
nor NOR4 (N5965, N5946, N2131, N1378, N5687);
buf BUF1 (N5966, N5963);
or OR2 (N5967, N5956, N3698);
buf BUF1 (N5968, N5939);
xor XOR2 (N5969, N5967, N1785);
or OR2 (N5970, N5964, N278);
xor XOR2 (N5971, N5932, N701);
nor NOR3 (N5972, N5960, N3976, N891);
nand NAND4 (N5973, N5961, N2829, N5093, N3141);
not NOT1 (N5974, N5969);
buf BUF1 (N5975, N5954);
nand NAND2 (N5976, N5974, N4041);
nand NAND3 (N5977, N5971, N2915, N4748);
xor XOR2 (N5978, N5973, N3267);
nor NOR3 (N5979, N5972, N5274, N2691);
and AND4 (N5980, N5951, N3395, N879, N1516);
xor XOR2 (N5981, N5976, N3906);
not NOT1 (N5982, N5978);
not NOT1 (N5983, N5979);
not NOT1 (N5984, N5982);
nand NAND4 (N5985, N5965, N2067, N798, N4259);
nor NOR3 (N5986, N5980, N3731, N1996);
buf BUF1 (N5987, N5975);
nand NAND3 (N5988, N5986, N2243, N2549);
buf BUF1 (N5989, N5983);
or OR4 (N5990, N5966, N1415, N3214, N2069);
nor NOR4 (N5991, N5970, N5088, N5338, N2021);
xor XOR2 (N5992, N5991, N5424);
or OR4 (N5993, N5981, N4027, N2666, N3851);
nand NAND4 (N5994, N5988, N4804, N2134, N2714);
nor NOR2 (N5995, N5992, N1574);
not NOT1 (N5996, N5995);
not NOT1 (N5997, N5987);
not NOT1 (N5998, N5968);
or OR4 (N5999, N5984, N2986, N3013, N3306);
xor XOR2 (N6000, N5996, N3320);
nor NOR2 (N6001, N5997, N2989);
buf BUF1 (N6002, N5999);
nor NOR2 (N6003, N5990, N1071);
and AND4 (N6004, N6003, N3524, N1127, N2007);
xor XOR2 (N6005, N5985, N33);
buf BUF1 (N6006, N5977);
xor XOR2 (N6007, N6002, N949);
nor NOR3 (N6008, N6004, N2121, N812);
nand NAND2 (N6009, N6007, N5375);
buf BUF1 (N6010, N6008);
nor NOR2 (N6011, N5993, N886);
and AND4 (N6012, N6001, N5177, N5832, N4131);
nor NOR3 (N6013, N6009, N1948, N1960);
and AND3 (N6014, N5998, N1051, N976);
and AND4 (N6015, N6011, N1283, N1779, N4920);
nand NAND2 (N6016, N6000, N1579);
not NOT1 (N6017, N5994);
or OR3 (N6018, N6010, N4006, N2413);
buf BUF1 (N6019, N5989);
xor XOR2 (N6020, N6014, N5927);
xor XOR2 (N6021, N6005, N2325);
and AND4 (N6022, N6021, N4113, N5717, N1346);
not NOT1 (N6023, N6022);
or OR4 (N6024, N6018, N2282, N830, N1427);
xor XOR2 (N6025, N6012, N2243);
buf BUF1 (N6026, N6025);
not NOT1 (N6027, N6017);
nor NOR3 (N6028, N6020, N5329, N3038);
nand NAND2 (N6029, N6016, N4919);
nand NAND3 (N6030, N6013, N2405, N2935);
nand NAND2 (N6031, N6026, N5486);
nor NOR4 (N6032, N6028, N3186, N2007, N3193);
buf BUF1 (N6033, N6031);
xor XOR2 (N6034, N6030, N1969);
not NOT1 (N6035, N6027);
not NOT1 (N6036, N6032);
nor NOR3 (N6037, N6033, N2028, N2304);
not NOT1 (N6038, N6023);
not NOT1 (N6039, N6029);
or OR4 (N6040, N6037, N4358, N3322, N318);
and AND3 (N6041, N6035, N1928, N4099);
xor XOR2 (N6042, N6024, N5492);
nand NAND3 (N6043, N6019, N289, N915);
buf BUF1 (N6044, N6036);
nand NAND4 (N6045, N6034, N3955, N4254, N1791);
nor NOR2 (N6046, N6038, N30);
nor NOR2 (N6047, N6015, N761);
not NOT1 (N6048, N6040);
and AND2 (N6049, N6043, N5330);
xor XOR2 (N6050, N6049, N2768);
nor NOR2 (N6051, N6041, N5395);
not NOT1 (N6052, N6051);
buf BUF1 (N6053, N6045);
buf BUF1 (N6054, N6050);
nand NAND4 (N6055, N6042, N2877, N868, N3208);
not NOT1 (N6056, N6044);
buf BUF1 (N6057, N6054);
nand NAND4 (N6058, N6048, N860, N4408, N445);
xor XOR2 (N6059, N6052, N3844);
buf BUF1 (N6060, N6059);
xor XOR2 (N6061, N6058, N2222);
not NOT1 (N6062, N6047);
nand NAND3 (N6063, N6053, N2205, N735);
buf BUF1 (N6064, N6061);
or OR3 (N6065, N6057, N2064, N920);
nor NOR3 (N6066, N6063, N3948, N3884);
nor NOR4 (N6067, N6006, N4622, N2938, N4616);
xor XOR2 (N6068, N6064, N5888);
nor NOR4 (N6069, N6065, N1954, N695, N371);
not NOT1 (N6070, N6060);
or OR4 (N6071, N6056, N3530, N2427, N5769);
or OR2 (N6072, N6062, N3909);
or OR2 (N6073, N6066, N5559);
not NOT1 (N6074, N6068);
nor NOR2 (N6075, N6071, N3162);
xor XOR2 (N6076, N6075, N649);
xor XOR2 (N6077, N6067, N5653);
not NOT1 (N6078, N6072);
and AND2 (N6079, N6074, N514);
and AND2 (N6080, N6070, N242);
nor NOR4 (N6081, N6077, N2479, N763, N3448);
nor NOR3 (N6082, N6081, N5699, N4420);
nand NAND2 (N6083, N6055, N1149);
xor XOR2 (N6084, N6073, N4324);
nor NOR2 (N6085, N6082, N214);
and AND2 (N6086, N6084, N4584);
or OR4 (N6087, N6085, N4369, N4565, N670);
and AND2 (N6088, N6080, N4905);
xor XOR2 (N6089, N6039, N1681);
nand NAND2 (N6090, N6078, N5884);
not NOT1 (N6091, N6090);
nor NOR3 (N6092, N6088, N5573, N3603);
xor XOR2 (N6093, N6092, N1238);
not NOT1 (N6094, N6089);
nor NOR3 (N6095, N6079, N3291, N178);
nand NAND3 (N6096, N6069, N100, N4193);
xor XOR2 (N6097, N6093, N161);
and AND4 (N6098, N6094, N4000, N4304, N3862);
not NOT1 (N6099, N6095);
not NOT1 (N6100, N6099);
nand NAND4 (N6101, N6087, N1092, N3286, N88);
nor NOR3 (N6102, N6100, N4349, N1666);
nand NAND3 (N6103, N6076, N3067, N2794);
nand NAND4 (N6104, N6102, N3498, N584, N2688);
not NOT1 (N6105, N6098);
xor XOR2 (N6106, N6083, N3705);
or OR4 (N6107, N6097, N1324, N1566, N4652);
buf BUF1 (N6108, N6101);
nand NAND3 (N6109, N6107, N5462, N3134);
and AND3 (N6110, N6103, N3538, N6008);
nand NAND3 (N6111, N6086, N3392, N4486);
buf BUF1 (N6112, N6046);
nor NOR3 (N6113, N6096, N4633, N4388);
xor XOR2 (N6114, N6109, N5030);
xor XOR2 (N6115, N6110, N3084);
buf BUF1 (N6116, N6113);
and AND4 (N6117, N6091, N2308, N3089, N330);
nor NOR2 (N6118, N6117, N5499);
xor XOR2 (N6119, N6115, N580);
not NOT1 (N6120, N6114);
nand NAND3 (N6121, N6116, N358, N780);
not NOT1 (N6122, N6119);
buf BUF1 (N6123, N6120);
not NOT1 (N6124, N6122);
or OR3 (N6125, N6108, N2491, N3268);
xor XOR2 (N6126, N6121, N2687);
buf BUF1 (N6127, N6126);
nand NAND2 (N6128, N6104, N768);
nor NOR4 (N6129, N6118, N4764, N1244, N1112);
or OR4 (N6130, N6105, N4255, N6044, N2239);
or OR2 (N6131, N6111, N4085);
or OR3 (N6132, N6124, N5096, N913);
nor NOR4 (N6133, N6127, N1416, N4112, N3007);
nor NOR4 (N6134, N6125, N4442, N2605, N3841);
and AND2 (N6135, N6128, N911);
nor NOR2 (N6136, N6134, N5064);
not NOT1 (N6137, N6132);
and AND4 (N6138, N6123, N545, N4449, N5742);
not NOT1 (N6139, N6135);
or OR4 (N6140, N6106, N4924, N1874, N742);
buf BUF1 (N6141, N6136);
and AND3 (N6142, N6112, N3900, N4684);
xor XOR2 (N6143, N6129, N3753);
xor XOR2 (N6144, N6133, N4319);
xor XOR2 (N6145, N6143, N2251);
buf BUF1 (N6146, N6130);
buf BUF1 (N6147, N6140);
not NOT1 (N6148, N6137);
not NOT1 (N6149, N6131);
not NOT1 (N6150, N6142);
nand NAND2 (N6151, N6149, N5311);
nand NAND3 (N6152, N6138, N3851, N4640);
buf BUF1 (N6153, N6151);
not NOT1 (N6154, N6146);
nor NOR2 (N6155, N6144, N4659);
buf BUF1 (N6156, N6139);
or OR3 (N6157, N6152, N1831, N5521);
nor NOR3 (N6158, N6156, N5367, N3333);
buf BUF1 (N6159, N6155);
nor NOR2 (N6160, N6157, N2118);
nand NAND4 (N6161, N6147, N4893, N3131, N4598);
and AND2 (N6162, N6154, N1607);
xor XOR2 (N6163, N6158, N950);
and AND3 (N6164, N6160, N3500, N3762);
not NOT1 (N6165, N6159);
nor NOR4 (N6166, N6148, N3249, N4972, N2183);
nor NOR3 (N6167, N6166, N695, N3749);
xor XOR2 (N6168, N6161, N576);
not NOT1 (N6169, N6163);
buf BUF1 (N6170, N6169);
xor XOR2 (N6171, N6165, N2157);
and AND3 (N6172, N6150, N3847, N4553);
nor NOR3 (N6173, N6172, N3097, N223);
or OR3 (N6174, N6145, N1377, N5035);
buf BUF1 (N6175, N6170);
nor NOR2 (N6176, N6141, N4445);
nand NAND4 (N6177, N6173, N4708, N3605, N429);
nor NOR2 (N6178, N6168, N218);
not NOT1 (N6179, N6176);
and AND2 (N6180, N6177, N1476);
and AND2 (N6181, N6167, N3057);
nor NOR2 (N6182, N6174, N141);
xor XOR2 (N6183, N6164, N2747);
nor NOR4 (N6184, N6171, N3590, N2168, N1077);
nand NAND2 (N6185, N6182, N4908);
or OR3 (N6186, N6179, N2920, N4130);
nor NOR4 (N6187, N6162, N2930, N970, N445);
or OR3 (N6188, N6180, N1284, N2956);
nand NAND3 (N6189, N6184, N359, N3114);
nand NAND3 (N6190, N6188, N1984, N353);
nand NAND3 (N6191, N6186, N3569, N3383);
nor NOR4 (N6192, N6189, N97, N1049, N3838);
or OR2 (N6193, N6178, N4388);
not NOT1 (N6194, N6181);
xor XOR2 (N6195, N6194, N5917);
and AND4 (N6196, N6183, N5948, N5554, N5323);
or OR3 (N6197, N6187, N3395, N4482);
and AND2 (N6198, N6192, N123);
or OR4 (N6199, N6197, N4614, N1037, N6153);
buf BUF1 (N6200, N3720);
xor XOR2 (N6201, N6200, N94);
or OR2 (N6202, N6199, N3776);
xor XOR2 (N6203, N6198, N596);
xor XOR2 (N6204, N6202, N5221);
nand NAND4 (N6205, N6193, N1628, N743, N967);
and AND2 (N6206, N6190, N664);
nand NAND4 (N6207, N6196, N170, N244, N1285);
xor XOR2 (N6208, N6175, N4398);
nand NAND4 (N6209, N6208, N3003, N273, N3493);
nor NOR4 (N6210, N6205, N1485, N581, N1511);
nor NOR4 (N6211, N6203, N3485, N2987, N4186);
nand NAND2 (N6212, N6204, N925);
not NOT1 (N6213, N6191);
buf BUF1 (N6214, N6210);
xor XOR2 (N6215, N6206, N2008);
not NOT1 (N6216, N6214);
xor XOR2 (N6217, N6216, N5207);
and AND4 (N6218, N6212, N3026, N6121, N1958);
nor NOR2 (N6219, N6201, N600);
nand NAND3 (N6220, N6185, N2793, N4322);
xor XOR2 (N6221, N6209, N62);
xor XOR2 (N6222, N6207, N3338);
or OR2 (N6223, N6195, N1493);
nand NAND3 (N6224, N6211, N770, N5329);
nand NAND2 (N6225, N6218, N797);
and AND4 (N6226, N6219, N1105, N4802, N5623);
nand NAND4 (N6227, N6217, N3800, N6058, N1162);
and AND3 (N6228, N6225, N3971, N2793);
xor XOR2 (N6229, N6226, N2315);
nand NAND4 (N6230, N6229, N3642, N1615, N1015);
nor NOR4 (N6231, N6224, N5106, N6205, N4654);
xor XOR2 (N6232, N6228, N384);
buf BUF1 (N6233, N6227);
nor NOR2 (N6234, N6231, N1326);
nor NOR3 (N6235, N6234, N1670, N4168);
and AND2 (N6236, N6233, N2982);
nand NAND2 (N6237, N6213, N3396);
or OR2 (N6238, N6223, N336);
nor NOR4 (N6239, N6215, N2246, N247, N5001);
buf BUF1 (N6240, N6236);
or OR3 (N6241, N6222, N1676, N5428);
and AND4 (N6242, N6230, N424, N5694, N5714);
not NOT1 (N6243, N6242);
nand NAND2 (N6244, N6235, N2596);
nor NOR3 (N6245, N6240, N895, N3296);
nor NOR4 (N6246, N6221, N2380, N5411, N5762);
or OR2 (N6247, N6245, N111);
nand NAND3 (N6248, N6241, N5282, N367);
buf BUF1 (N6249, N6220);
nor NOR2 (N6250, N6246, N4384);
buf BUF1 (N6251, N6232);
buf BUF1 (N6252, N6243);
buf BUF1 (N6253, N6247);
nor NOR2 (N6254, N6249, N5873);
and AND2 (N6255, N6254, N6228);
buf BUF1 (N6256, N6250);
and AND2 (N6257, N6255, N3453);
xor XOR2 (N6258, N6237, N882);
and AND2 (N6259, N6239, N1338);
and AND2 (N6260, N6253, N2657);
nand NAND3 (N6261, N6259, N2065, N941);
not NOT1 (N6262, N6251);
not NOT1 (N6263, N6257);
xor XOR2 (N6264, N6252, N5167);
or OR4 (N6265, N6248, N5857, N1963, N5774);
nand NAND2 (N6266, N6265, N2271);
nand NAND4 (N6267, N6238, N2264, N5207, N3394);
not NOT1 (N6268, N6258);
and AND4 (N6269, N6268, N5437, N3628, N521);
nor NOR2 (N6270, N6260, N3579);
and AND2 (N6271, N6256, N1748);
not NOT1 (N6272, N6270);
xor XOR2 (N6273, N6271, N4553);
or OR2 (N6274, N6264, N2606);
or OR4 (N6275, N6262, N2668, N3540, N1630);
and AND4 (N6276, N6266, N2410, N4617, N805);
buf BUF1 (N6277, N6273);
or OR3 (N6278, N6277, N2217, N4932);
nor NOR4 (N6279, N6269, N3868, N3343, N1318);
nor NOR4 (N6280, N6272, N5692, N979, N5777);
or OR4 (N6281, N6276, N5877, N2427, N2691);
buf BUF1 (N6282, N6263);
nand NAND3 (N6283, N6280, N4406, N5519);
xor XOR2 (N6284, N6261, N2108);
not NOT1 (N6285, N6274);
xor XOR2 (N6286, N6278, N2585);
nor NOR3 (N6287, N6275, N3129, N1571);
and AND2 (N6288, N6244, N2720);
nand NAND4 (N6289, N6281, N427, N4761, N2377);
or OR4 (N6290, N6284, N340, N3215, N345);
not NOT1 (N6291, N6286);
xor XOR2 (N6292, N6279, N1964);
and AND4 (N6293, N6287, N1933, N464, N1934);
buf BUF1 (N6294, N6282);
buf BUF1 (N6295, N6289);
and AND3 (N6296, N6267, N107, N2973);
not NOT1 (N6297, N6290);
or OR4 (N6298, N6296, N3862, N1373, N2873);
not NOT1 (N6299, N6298);
buf BUF1 (N6300, N6297);
nand NAND2 (N6301, N6293, N5030);
nor NOR2 (N6302, N6292, N314);
xor XOR2 (N6303, N6283, N5989);
xor XOR2 (N6304, N6294, N1005);
nand NAND3 (N6305, N6302, N906, N1450);
xor XOR2 (N6306, N6291, N4292);
nand NAND2 (N6307, N6300, N4822);
nor NOR2 (N6308, N6304, N1747);
or OR3 (N6309, N6307, N3907, N4688);
or OR4 (N6310, N6309, N2287, N4976, N1457);
not NOT1 (N6311, N6303);
buf BUF1 (N6312, N6299);
xor XOR2 (N6313, N6312, N940);
xor XOR2 (N6314, N6311, N326);
or OR4 (N6315, N6306, N4283, N5571, N5233);
nand NAND2 (N6316, N6295, N895);
buf BUF1 (N6317, N6285);
buf BUF1 (N6318, N6314);
buf BUF1 (N6319, N6316);
xor XOR2 (N6320, N6315, N4871);
xor XOR2 (N6321, N6301, N5844);
buf BUF1 (N6322, N6321);
xor XOR2 (N6323, N6318, N2123);
and AND3 (N6324, N6313, N2606, N4500);
and AND4 (N6325, N6320, N2073, N2290, N4957);
xor XOR2 (N6326, N6319, N154);
or OR4 (N6327, N6305, N499, N5992, N4582);
xor XOR2 (N6328, N6310, N1821);
buf BUF1 (N6329, N6323);
buf BUF1 (N6330, N6317);
buf BUF1 (N6331, N6322);
nand NAND3 (N6332, N6288, N5826, N1703);
nor NOR3 (N6333, N6331, N2099, N2099);
nor NOR4 (N6334, N6329, N944, N847, N2058);
nand NAND3 (N6335, N6326, N4131, N6072);
nor NOR2 (N6336, N6334, N6045);
and AND2 (N6337, N6333, N5855);
nor NOR4 (N6338, N6328, N24, N4127, N5357);
not NOT1 (N6339, N6327);
nand NAND4 (N6340, N6337, N5615, N4780, N791);
nand NAND3 (N6341, N6335, N6023, N882);
or OR4 (N6342, N6338, N1328, N3150, N6167);
not NOT1 (N6343, N6324);
and AND2 (N6344, N6308, N1826);
or OR3 (N6345, N6330, N2419, N1044);
nor NOR3 (N6346, N6339, N5464, N4525);
xor XOR2 (N6347, N6346, N5892);
and AND4 (N6348, N6336, N5643, N4534, N1836);
not NOT1 (N6349, N6325);
buf BUF1 (N6350, N6332);
xor XOR2 (N6351, N6345, N4630);
xor XOR2 (N6352, N6351, N2275);
buf BUF1 (N6353, N6341);
or OR4 (N6354, N6348, N4448, N5706, N3837);
or OR2 (N6355, N6340, N5869);
and AND2 (N6356, N6343, N1799);
not NOT1 (N6357, N6353);
not NOT1 (N6358, N6344);
nand NAND2 (N6359, N6355, N3184);
and AND3 (N6360, N6352, N2116, N1157);
not NOT1 (N6361, N6356);
nand NAND3 (N6362, N6347, N3118, N4340);
xor XOR2 (N6363, N6350, N1323);
xor XOR2 (N6364, N6349, N3371);
xor XOR2 (N6365, N6362, N5033);
buf BUF1 (N6366, N6365);
nor NOR4 (N6367, N6354, N2524, N2949, N2620);
nor NOR4 (N6368, N6366, N2394, N3827, N3529);
xor XOR2 (N6369, N6360, N2470);
xor XOR2 (N6370, N6357, N4085);
nor NOR2 (N6371, N6367, N6143);
buf BUF1 (N6372, N6358);
nand NAND2 (N6373, N6370, N3933);
and AND4 (N6374, N6364, N2937, N283, N748);
and AND2 (N6375, N6371, N880);
nand NAND3 (N6376, N6342, N1443, N1477);
nor NOR4 (N6377, N6359, N3676, N576, N3459);
not NOT1 (N6378, N6372);
or OR2 (N6379, N6377, N5202);
not NOT1 (N6380, N6373);
nor NOR2 (N6381, N6361, N1197);
nor NOR2 (N6382, N6379, N117);
nor NOR3 (N6383, N6380, N5301, N3392);
nand NAND2 (N6384, N6363, N6018);
xor XOR2 (N6385, N6381, N2114);
nor NOR3 (N6386, N6383, N550, N1411);
nor NOR3 (N6387, N6368, N5796, N2502);
buf BUF1 (N6388, N6385);
not NOT1 (N6389, N6386);
or OR2 (N6390, N6376, N5667);
xor XOR2 (N6391, N6382, N4932);
nor NOR2 (N6392, N6390, N6327);
and AND4 (N6393, N6378, N1362, N2360, N3017);
nor NOR3 (N6394, N6374, N1113, N372);
xor XOR2 (N6395, N6394, N1905);
buf BUF1 (N6396, N6375);
or OR4 (N6397, N6384, N2827, N5554, N6053);
nor NOR4 (N6398, N6389, N3184, N4417, N489);
and AND3 (N6399, N6395, N5815, N5796);
nor NOR3 (N6400, N6369, N1754, N3088);
nor NOR4 (N6401, N6392, N3437, N6219, N482);
nand NAND4 (N6402, N6391, N3607, N764, N3006);
buf BUF1 (N6403, N6396);
not NOT1 (N6404, N6402);
and AND4 (N6405, N6398, N4422, N4955, N2680);
xor XOR2 (N6406, N6405, N3357);
and AND3 (N6407, N6400, N3869, N4628);
nand NAND3 (N6408, N6404, N3924, N1173);
and AND2 (N6409, N6397, N2057);
or OR4 (N6410, N6406, N4912, N5580, N4458);
buf BUF1 (N6411, N6408);
nor NOR2 (N6412, N6403, N6323);
nor NOR2 (N6413, N6410, N6376);
buf BUF1 (N6414, N6407);
not NOT1 (N6415, N6413);
nor NOR2 (N6416, N6387, N1469);
not NOT1 (N6417, N6393);
and AND3 (N6418, N6415, N563, N1098);
nand NAND3 (N6419, N6401, N5781, N3629);
or OR3 (N6420, N6388, N5141, N4892);
and AND2 (N6421, N6417, N4778);
xor XOR2 (N6422, N6412, N690);
or OR2 (N6423, N6399, N5547);
and AND4 (N6424, N6420, N2428, N4067, N1330);
xor XOR2 (N6425, N6422, N1559);
xor XOR2 (N6426, N6411, N4894);
buf BUF1 (N6427, N6423);
or OR2 (N6428, N6424, N526);
buf BUF1 (N6429, N6409);
not NOT1 (N6430, N6429);
not NOT1 (N6431, N6414);
or OR4 (N6432, N6430, N2468, N2936, N2160);
or OR2 (N6433, N6426, N1147);
or OR3 (N6434, N6418, N3190, N4457);
nor NOR4 (N6435, N6427, N1586, N49, N1312);
buf BUF1 (N6436, N6434);
or OR2 (N6437, N6428, N3634);
xor XOR2 (N6438, N6421, N6279);
nand NAND4 (N6439, N6436, N1654, N3535, N1549);
and AND4 (N6440, N6437, N4359, N6049, N1527);
nor NOR3 (N6441, N6416, N928, N2417);
xor XOR2 (N6442, N6439, N4606);
not NOT1 (N6443, N6419);
or OR2 (N6444, N6441, N2739);
nor NOR4 (N6445, N6432, N3480, N4101, N3194);
buf BUF1 (N6446, N6445);
xor XOR2 (N6447, N6438, N3994);
nand NAND4 (N6448, N6435, N1170, N1930, N6300);
nand NAND3 (N6449, N6431, N397, N1343);
nor NOR3 (N6450, N6448, N3863, N3225);
xor XOR2 (N6451, N6433, N5850);
xor XOR2 (N6452, N6425, N6306);
nand NAND2 (N6453, N6449, N5173);
not NOT1 (N6454, N6443);
and AND3 (N6455, N6453, N5997, N3533);
or OR3 (N6456, N6440, N640, N3809);
not NOT1 (N6457, N6456);
or OR2 (N6458, N6457, N4178);
xor XOR2 (N6459, N6446, N4256);
or OR4 (N6460, N6455, N920, N3830, N4771);
or OR4 (N6461, N6454, N3953, N3711, N3992);
xor XOR2 (N6462, N6460, N177);
xor XOR2 (N6463, N6447, N1526);
nor NOR3 (N6464, N6452, N3218, N6262);
buf BUF1 (N6465, N6451);
or OR4 (N6466, N6444, N865, N2541, N5915);
and AND4 (N6467, N6442, N2896, N504, N2654);
nand NAND2 (N6468, N6465, N3500);
nor NOR4 (N6469, N6450, N712, N2353, N2381);
and AND2 (N6470, N6468, N3360);
nand NAND4 (N6471, N6470, N2290, N5659, N4983);
and AND4 (N6472, N6459, N297, N2385, N279);
not NOT1 (N6473, N6469);
buf BUF1 (N6474, N6458);
nand NAND4 (N6475, N6474, N124, N3637, N3125);
nand NAND4 (N6476, N6472, N5810, N580, N1500);
nor NOR4 (N6477, N6467, N3488, N6012, N1194);
buf BUF1 (N6478, N6476);
not NOT1 (N6479, N6464);
nor NOR2 (N6480, N6463, N4090);
not NOT1 (N6481, N6475);
or OR4 (N6482, N6473, N132, N4026, N5029);
not NOT1 (N6483, N6478);
buf BUF1 (N6484, N6483);
buf BUF1 (N6485, N6471);
not NOT1 (N6486, N6484);
buf BUF1 (N6487, N6480);
not NOT1 (N6488, N6461);
xor XOR2 (N6489, N6481, N1330);
nor NOR4 (N6490, N6488, N2576, N3109, N2141);
and AND4 (N6491, N6466, N4611, N6371, N4107);
not NOT1 (N6492, N6462);
not NOT1 (N6493, N6490);
or OR2 (N6494, N6489, N934);
xor XOR2 (N6495, N6487, N3937);
buf BUF1 (N6496, N6485);
xor XOR2 (N6497, N6492, N2433);
and AND2 (N6498, N6495, N3518);
buf BUF1 (N6499, N6486);
not NOT1 (N6500, N6499);
and AND3 (N6501, N6491, N5031, N3410);
not NOT1 (N6502, N6500);
nor NOR4 (N6503, N6477, N6026, N2134, N5882);
nand NAND2 (N6504, N6501, N4455);
xor XOR2 (N6505, N6482, N2338);
or OR2 (N6506, N6494, N1892);
xor XOR2 (N6507, N6479, N5588);
nor NOR4 (N6508, N6505, N1261, N156, N1194);
and AND2 (N6509, N6502, N4513);
nor NOR4 (N6510, N6508, N5928, N3896, N2505);
xor XOR2 (N6511, N6510, N5984);
nand NAND3 (N6512, N6507, N2137, N2166);
nor NOR4 (N6513, N6497, N839, N1491, N2263);
nand NAND2 (N6514, N6504, N5983);
nand NAND4 (N6515, N6511, N3733, N43, N5419);
nand NAND4 (N6516, N6509, N954, N2174, N2679);
xor XOR2 (N6517, N6506, N4088);
nand NAND2 (N6518, N6512, N926);
xor XOR2 (N6519, N6493, N4482);
not NOT1 (N6520, N6515);
buf BUF1 (N6521, N6514);
and AND2 (N6522, N6520, N1872);
not NOT1 (N6523, N6513);
not NOT1 (N6524, N6519);
buf BUF1 (N6525, N6516);
not NOT1 (N6526, N6523);
or OR3 (N6527, N6524, N5052, N3351);
and AND3 (N6528, N6498, N5517, N2591);
not NOT1 (N6529, N6503);
xor XOR2 (N6530, N6526, N2499);
nand NAND2 (N6531, N6529, N1650);
nor NOR3 (N6532, N6521, N5580, N3328);
nor NOR3 (N6533, N6525, N5391, N3752);
nor NOR3 (N6534, N6517, N3374, N4792);
not NOT1 (N6535, N6534);
nand NAND3 (N6536, N6522, N4022, N4296);
not NOT1 (N6537, N6496);
xor XOR2 (N6538, N6537, N3421);
xor XOR2 (N6539, N6527, N1515);
not NOT1 (N6540, N6535);
and AND3 (N6541, N6531, N1164, N6363);
or OR4 (N6542, N6530, N357, N5964, N820);
and AND2 (N6543, N6541, N1830);
and AND2 (N6544, N6528, N1634);
not NOT1 (N6545, N6532);
nor NOR3 (N6546, N6543, N1604, N1207);
and AND3 (N6547, N6545, N2588, N2408);
xor XOR2 (N6548, N6539, N2140);
xor XOR2 (N6549, N6547, N3736);
buf BUF1 (N6550, N6548);
not NOT1 (N6551, N6549);
nor NOR3 (N6552, N6533, N2687, N4257);
buf BUF1 (N6553, N6538);
and AND2 (N6554, N6546, N4905);
buf BUF1 (N6555, N6542);
not NOT1 (N6556, N6555);
or OR4 (N6557, N6556, N4697, N1643, N5522);
or OR2 (N6558, N6536, N1935);
or OR3 (N6559, N6553, N4222, N5);
nand NAND2 (N6560, N6540, N6489);
nand NAND2 (N6561, N6551, N1638);
nand NAND4 (N6562, N6518, N2867, N4981, N5809);
not NOT1 (N6563, N6557);
and AND3 (N6564, N6561, N3930, N4105);
and AND4 (N6565, N6563, N3159, N2820, N3146);
not NOT1 (N6566, N6550);
or OR3 (N6567, N6562, N5371, N3908);
xor XOR2 (N6568, N6552, N6227);
nand NAND4 (N6569, N6565, N3411, N2755, N5765);
nor NOR3 (N6570, N6559, N3092, N4195);
buf BUF1 (N6571, N6558);
nand NAND3 (N6572, N6568, N3274, N5643);
xor XOR2 (N6573, N6572, N3948);
or OR2 (N6574, N6566, N4995);
nand NAND2 (N6575, N6574, N1476);
xor XOR2 (N6576, N6571, N6562);
not NOT1 (N6577, N6573);
xor XOR2 (N6578, N6576, N5620);
nand NAND4 (N6579, N6544, N4176, N5906, N1597);
not NOT1 (N6580, N6567);
or OR2 (N6581, N6580, N182);
and AND4 (N6582, N6560, N4299, N3743, N5853);
buf BUF1 (N6583, N6554);
nand NAND4 (N6584, N6578, N3680, N4285, N2660);
nor NOR3 (N6585, N6564, N2488, N4329);
and AND4 (N6586, N6575, N474, N5974, N664);
not NOT1 (N6587, N6577);
buf BUF1 (N6588, N6569);
and AND2 (N6589, N6581, N1638);
and AND2 (N6590, N6583, N3503);
and AND3 (N6591, N6570, N1188, N2713);
xor XOR2 (N6592, N6589, N5892);
nor NOR2 (N6593, N6582, N5618);
nor NOR4 (N6594, N6587, N3244, N2062, N2655);
nor NOR4 (N6595, N6579, N3107, N5329, N2935);
nor NOR2 (N6596, N6588, N3589);
nand NAND4 (N6597, N6593, N6100, N2715, N779);
not NOT1 (N6598, N6595);
not NOT1 (N6599, N6598);
xor XOR2 (N6600, N6599, N2262);
buf BUF1 (N6601, N6592);
nand NAND4 (N6602, N6585, N1998, N4667, N6434);
nand NAND2 (N6603, N6590, N4898);
nand NAND2 (N6604, N6586, N2747);
nand NAND2 (N6605, N6594, N3406);
not NOT1 (N6606, N6591);
not NOT1 (N6607, N6606);
and AND2 (N6608, N6604, N403);
xor XOR2 (N6609, N6597, N3314);
not NOT1 (N6610, N6602);
not NOT1 (N6611, N6600);
xor XOR2 (N6612, N6601, N6604);
buf BUF1 (N6613, N6596);
xor XOR2 (N6614, N6609, N4772);
or OR3 (N6615, N6611, N5362, N5142);
buf BUF1 (N6616, N6610);
nand NAND3 (N6617, N6605, N1597, N5597);
not NOT1 (N6618, N6608);
nor NOR4 (N6619, N6616, N1859, N4515, N1076);
or OR2 (N6620, N6613, N6585);
or OR4 (N6621, N6603, N6588, N1407, N2411);
and AND2 (N6622, N6614, N611);
and AND4 (N6623, N6612, N1567, N563, N5372);
or OR4 (N6624, N6584, N5233, N846, N1797);
nor NOR2 (N6625, N6624, N536);
nand NAND2 (N6626, N6620, N1679);
nand NAND4 (N6627, N6615, N1401, N2283, N857);
not NOT1 (N6628, N6621);
and AND4 (N6629, N6617, N5893, N2231, N6148);
buf BUF1 (N6630, N6628);
nor NOR2 (N6631, N6625, N2172);
xor XOR2 (N6632, N6623, N1320);
not NOT1 (N6633, N6607);
nor NOR3 (N6634, N6633, N6456, N319);
and AND4 (N6635, N6629, N52, N4602, N3492);
or OR3 (N6636, N6619, N5369, N3480);
nand NAND4 (N6637, N6627, N3900, N1477, N6187);
nor NOR3 (N6638, N6634, N4141, N5970);
and AND3 (N6639, N6631, N1177, N1864);
xor XOR2 (N6640, N6639, N6316);
and AND4 (N6641, N6618, N2341, N4193, N4392);
or OR2 (N6642, N6637, N1985);
or OR4 (N6643, N6630, N3571, N1124, N3154);
or OR4 (N6644, N6636, N4724, N2824, N3708);
xor XOR2 (N6645, N6644, N4202);
nor NOR4 (N6646, N6645, N292, N3981, N3316);
or OR4 (N6647, N6638, N642, N4780, N1684);
not NOT1 (N6648, N6641);
not NOT1 (N6649, N6622);
and AND4 (N6650, N6632, N1383, N886, N5141);
nand NAND3 (N6651, N6643, N671, N2222);
and AND2 (N6652, N6647, N611);
nand NAND3 (N6653, N6650, N6505, N6046);
buf BUF1 (N6654, N6640);
xor XOR2 (N6655, N6654, N4709);
xor XOR2 (N6656, N6653, N1520);
buf BUF1 (N6657, N6646);
not NOT1 (N6658, N6656);
xor XOR2 (N6659, N6649, N2839);
nand NAND2 (N6660, N6657, N3167);
buf BUF1 (N6661, N6642);
buf BUF1 (N6662, N6660);
and AND2 (N6663, N6635, N4541);
nand NAND4 (N6664, N6626, N5348, N4434, N557);
not NOT1 (N6665, N6661);
xor XOR2 (N6666, N6659, N1101);
buf BUF1 (N6667, N6662);
not NOT1 (N6668, N6663);
buf BUF1 (N6669, N6667);
not NOT1 (N6670, N6655);
xor XOR2 (N6671, N6670, N6476);
xor XOR2 (N6672, N6648, N5348);
or OR2 (N6673, N6669, N643);
not NOT1 (N6674, N6658);
nor NOR4 (N6675, N6666, N3261, N3760, N3434);
nor NOR3 (N6676, N6651, N45, N2414);
nor NOR2 (N6677, N6675, N3431);
or OR2 (N6678, N6677, N3559);
buf BUF1 (N6679, N6665);
or OR4 (N6680, N6668, N1959, N1587, N4299);
nor NOR4 (N6681, N6678, N642, N4793, N2019);
and AND4 (N6682, N6681, N5324, N3321, N3466);
nand NAND4 (N6683, N6679, N6363, N3866, N4390);
buf BUF1 (N6684, N6683);
nand NAND4 (N6685, N6682, N3232, N1759, N4995);
not NOT1 (N6686, N6674);
or OR2 (N6687, N6684, N972);
xor XOR2 (N6688, N6687, N789);
not NOT1 (N6689, N6671);
nor NOR2 (N6690, N6672, N5357);
nand NAND3 (N6691, N6685, N1223, N108);
or OR3 (N6692, N6690, N1451, N3483);
xor XOR2 (N6693, N6692, N2717);
nand NAND4 (N6694, N6680, N3219, N5542, N1166);
nand NAND2 (N6695, N6688, N499);
nand NAND4 (N6696, N6689, N2004, N5406, N4830);
nand NAND3 (N6697, N6673, N808, N1974);
not NOT1 (N6698, N6696);
xor XOR2 (N6699, N6693, N3758);
and AND3 (N6700, N6676, N1631, N2452);
buf BUF1 (N6701, N6664);
or OR4 (N6702, N6694, N1435, N6649, N2798);
or OR3 (N6703, N6700, N803, N6116);
buf BUF1 (N6704, N6697);
nor NOR3 (N6705, N6701, N2793, N4157);
and AND4 (N6706, N6705, N1368, N5513, N6584);
nor NOR4 (N6707, N6702, N2737, N5048, N4984);
nor NOR2 (N6708, N6698, N5388);
nand NAND4 (N6709, N6706, N566, N5416, N5273);
nand NAND2 (N6710, N6707, N5748);
xor XOR2 (N6711, N6708, N3358);
buf BUF1 (N6712, N6691);
xor XOR2 (N6713, N6699, N3571);
nand NAND3 (N6714, N6695, N6578, N1771);
xor XOR2 (N6715, N6704, N5927);
nor NOR2 (N6716, N6713, N2448);
buf BUF1 (N6717, N6686);
nand NAND3 (N6718, N6715, N3206, N1821);
or OR3 (N6719, N6652, N4593, N5334);
nand NAND2 (N6720, N6717, N135);
nand NAND2 (N6721, N6711, N342);
nor NOR2 (N6722, N6710, N2794);
and AND2 (N6723, N6721, N1986);
not NOT1 (N6724, N6716);
xor XOR2 (N6725, N6720, N1254);
xor XOR2 (N6726, N6714, N4727);
or OR2 (N6727, N6709, N3456);
or OR2 (N6728, N6718, N2235);
and AND3 (N6729, N6725, N1066, N6130);
nor NOR3 (N6730, N6719, N3509, N1321);
xor XOR2 (N6731, N6726, N6313);
not NOT1 (N6732, N6731);
not NOT1 (N6733, N6728);
or OR3 (N6734, N6729, N2382, N3127);
or OR3 (N6735, N6733, N2057, N4808);
or OR3 (N6736, N6734, N631, N5368);
and AND2 (N6737, N6730, N2479);
nor NOR3 (N6738, N6723, N2295, N6223);
not NOT1 (N6739, N6735);
buf BUF1 (N6740, N6722);
and AND3 (N6741, N6712, N5160, N3816);
xor XOR2 (N6742, N6741, N3584);
nand NAND2 (N6743, N6703, N3394);
not NOT1 (N6744, N6724);
nand NAND4 (N6745, N6736, N117, N1637, N2792);
nor NOR2 (N6746, N6737, N6308);
not NOT1 (N6747, N6739);
or OR3 (N6748, N6747, N6016, N1655);
not NOT1 (N6749, N6738);
or OR4 (N6750, N6742, N1885, N4741, N87);
nand NAND2 (N6751, N6740, N1548);
buf BUF1 (N6752, N6748);
and AND4 (N6753, N6751, N2520, N4949, N6656);
buf BUF1 (N6754, N6749);
buf BUF1 (N6755, N6752);
not NOT1 (N6756, N6753);
buf BUF1 (N6757, N6746);
not NOT1 (N6758, N6744);
and AND2 (N6759, N6758, N5533);
nand NAND3 (N6760, N6750, N1502, N3611);
not NOT1 (N6761, N6745);
or OR4 (N6762, N6754, N5460, N1153, N3783);
not NOT1 (N6763, N6755);
not NOT1 (N6764, N6762);
buf BUF1 (N6765, N6743);
buf BUF1 (N6766, N6727);
not NOT1 (N6767, N6757);
nor NOR4 (N6768, N6767, N6203, N2097, N1278);
buf BUF1 (N6769, N6732);
nand NAND3 (N6770, N6763, N3682, N3035);
or OR3 (N6771, N6765, N2144, N1332);
nor NOR3 (N6772, N6756, N1540, N287);
nand NAND2 (N6773, N6768, N6197);
or OR2 (N6774, N6771, N422);
xor XOR2 (N6775, N6772, N222);
xor XOR2 (N6776, N6774, N5955);
not NOT1 (N6777, N6773);
nor NOR3 (N6778, N6761, N6392, N5724);
and AND3 (N6779, N6766, N1292, N3515);
not NOT1 (N6780, N6776);
nand NAND2 (N6781, N6780, N1905);
not NOT1 (N6782, N6770);
or OR4 (N6783, N6777, N928, N5204, N3473);
buf BUF1 (N6784, N6764);
xor XOR2 (N6785, N6760, N5999);
nor NOR2 (N6786, N6783, N2005);
xor XOR2 (N6787, N6781, N6081);
nor NOR4 (N6788, N6784, N4696, N3043, N5791);
or OR4 (N6789, N6779, N6272, N1857, N1416);
buf BUF1 (N6790, N6778);
or OR2 (N6791, N6788, N429);
xor XOR2 (N6792, N6775, N3225);
xor XOR2 (N6793, N6787, N2780);
nand NAND2 (N6794, N6782, N1678);
or OR3 (N6795, N6785, N6280, N382);
or OR2 (N6796, N6792, N525);
and AND2 (N6797, N6769, N2259);
nor NOR3 (N6798, N6793, N5510, N2202);
nand NAND2 (N6799, N6790, N1366);
nand NAND3 (N6800, N6786, N1306, N1559);
nand NAND2 (N6801, N6794, N2628);
nand NAND2 (N6802, N6799, N3285);
not NOT1 (N6803, N6801);
buf BUF1 (N6804, N6803);
and AND2 (N6805, N6798, N6133);
and AND2 (N6806, N6759, N2967);
and AND4 (N6807, N6791, N1937, N326, N1784);
not NOT1 (N6808, N6807);
nand NAND3 (N6809, N6805, N5835, N2321);
xor XOR2 (N6810, N6804, N6191);
nor NOR2 (N6811, N6802, N4440);
nor NOR2 (N6812, N6797, N414);
or OR3 (N6813, N6795, N6281, N3037);
not NOT1 (N6814, N6813);
nor NOR4 (N6815, N6800, N6275, N1045, N3290);
and AND3 (N6816, N6809, N2407, N6450);
not NOT1 (N6817, N6815);
and AND2 (N6818, N6812, N3548);
nor NOR2 (N6819, N6810, N2408);
buf BUF1 (N6820, N6818);
nand NAND3 (N6821, N6806, N6406, N3683);
buf BUF1 (N6822, N6814);
nand NAND2 (N6823, N6808, N6285);
xor XOR2 (N6824, N6819, N886);
nor NOR2 (N6825, N6816, N5406);
not NOT1 (N6826, N6789);
or OR2 (N6827, N6825, N2765);
xor XOR2 (N6828, N6817, N5400);
buf BUF1 (N6829, N6824);
not NOT1 (N6830, N6826);
buf BUF1 (N6831, N6830);
xor XOR2 (N6832, N6823, N6267);
xor XOR2 (N6833, N6831, N760);
or OR2 (N6834, N6828, N4571);
nor NOR2 (N6835, N6796, N3326);
not NOT1 (N6836, N6833);
and AND2 (N6837, N6835, N6782);
and AND2 (N6838, N6834, N94);
or OR4 (N6839, N6822, N2666, N2672, N726);
or OR3 (N6840, N6827, N5265, N2532);
or OR4 (N6841, N6836, N3771, N6048, N6451);
nor NOR2 (N6842, N6829, N5926);
nor NOR4 (N6843, N6841, N5193, N4471, N499);
not NOT1 (N6844, N6842);
buf BUF1 (N6845, N6843);
nor NOR3 (N6846, N6821, N4414, N735);
xor XOR2 (N6847, N6840, N6448);
nand NAND4 (N6848, N6837, N5356, N6366, N4997);
xor XOR2 (N6849, N6811, N756);
and AND3 (N6850, N6846, N4753, N958);
nand NAND2 (N6851, N6847, N4492);
nor NOR4 (N6852, N6832, N5294, N4975, N264);
nor NOR4 (N6853, N6844, N2082, N4571, N756);
nand NAND2 (N6854, N6853, N2249);
or OR3 (N6855, N6838, N4911, N5919);
and AND3 (N6856, N6839, N3826, N247);
or OR4 (N6857, N6851, N3527, N42, N5049);
or OR3 (N6858, N6856, N1202, N503);
buf BUF1 (N6859, N6855);
buf BUF1 (N6860, N6852);
or OR4 (N6861, N6858, N1799, N4210, N713);
nand NAND2 (N6862, N6859, N1488);
buf BUF1 (N6863, N6862);
xor XOR2 (N6864, N6849, N757);
not NOT1 (N6865, N6864);
nand NAND4 (N6866, N6861, N4996, N1393, N2208);
buf BUF1 (N6867, N6820);
or OR4 (N6868, N6863, N5648, N1673, N4251);
nand NAND3 (N6869, N6854, N6660, N4995);
xor XOR2 (N6870, N6857, N6040);
not NOT1 (N6871, N6870);
buf BUF1 (N6872, N6867);
or OR3 (N6873, N6866, N4678, N1366);
or OR2 (N6874, N6873, N4495);
nand NAND3 (N6875, N6874, N3005, N554);
not NOT1 (N6876, N6845);
and AND2 (N6877, N6868, N2190);
or OR4 (N6878, N6869, N1786, N6425, N5196);
nor NOR3 (N6879, N6876, N3267, N5469);
nand NAND3 (N6880, N6878, N3341, N6870);
and AND2 (N6881, N6871, N1392);
xor XOR2 (N6882, N6877, N2624);
and AND4 (N6883, N6881, N6489, N1278, N232);
not NOT1 (N6884, N6883);
xor XOR2 (N6885, N6882, N4365);
nor NOR4 (N6886, N6880, N2712, N3484, N5105);
not NOT1 (N6887, N6884);
buf BUF1 (N6888, N6879);
nor NOR2 (N6889, N6860, N5400);
buf BUF1 (N6890, N6886);
not NOT1 (N6891, N6865);
and AND3 (N6892, N6848, N3462, N1253);
nand NAND2 (N6893, N6890, N1593);
buf BUF1 (N6894, N6885);
not NOT1 (N6895, N6875);
nor NOR2 (N6896, N6850, N6540);
nand NAND2 (N6897, N6895, N706);
not NOT1 (N6898, N6892);
xor XOR2 (N6899, N6888, N2081);
xor XOR2 (N6900, N6891, N5513);
xor XOR2 (N6901, N6896, N5234);
buf BUF1 (N6902, N6889);
nor NOR4 (N6903, N6901, N4088, N2736, N1312);
buf BUF1 (N6904, N6897);
and AND2 (N6905, N6904, N4895);
nor NOR3 (N6906, N6902, N2617, N3161);
not NOT1 (N6907, N6887);
or OR2 (N6908, N6893, N5573);
or OR3 (N6909, N6894, N1931, N3103);
nand NAND3 (N6910, N6872, N3411, N6516);
and AND4 (N6911, N6908, N3519, N2447, N4212);
nor NOR4 (N6912, N6911, N6504, N4390, N4591);
xor XOR2 (N6913, N6899, N5803);
nand NAND3 (N6914, N6903, N4291, N2644);
nand NAND2 (N6915, N6913, N6572);
not NOT1 (N6916, N6910);
xor XOR2 (N6917, N6907, N3188);
nand NAND4 (N6918, N6915, N5099, N3510, N6860);
xor XOR2 (N6919, N6909, N1748);
and AND3 (N6920, N6906, N2484, N1757);
xor XOR2 (N6921, N6918, N2727);
and AND4 (N6922, N6898, N6652, N5852, N2626);
and AND2 (N6923, N6912, N2951);
buf BUF1 (N6924, N6919);
xor XOR2 (N6925, N6905, N4568);
not NOT1 (N6926, N6921);
nand NAND2 (N6927, N6922, N2529);
and AND4 (N6928, N6927, N2114, N6864, N6029);
buf BUF1 (N6929, N6914);
and AND3 (N6930, N6916, N5260, N4554);
not NOT1 (N6931, N6926);
nor NOR4 (N6932, N6917, N6107, N3175, N6856);
nor NOR4 (N6933, N6929, N5150, N6739, N3723);
xor XOR2 (N6934, N6932, N5554);
xor XOR2 (N6935, N6933, N4298);
buf BUF1 (N6936, N6900);
not NOT1 (N6937, N6930);
buf BUF1 (N6938, N6934);
buf BUF1 (N6939, N6931);
not NOT1 (N6940, N6925);
nor NOR3 (N6941, N6935, N5476, N6801);
and AND4 (N6942, N6939, N2489, N264, N1004);
or OR3 (N6943, N6923, N1446, N2426);
and AND4 (N6944, N6938, N1089, N2178, N2356);
nor NOR3 (N6945, N6941, N647, N4313);
buf BUF1 (N6946, N6945);
nand NAND4 (N6947, N6944, N52, N6458, N1826);
or OR4 (N6948, N6928, N6361, N1276, N829);
and AND3 (N6949, N6946, N6427, N1232);
not NOT1 (N6950, N6949);
or OR3 (N6951, N6924, N519, N1120);
not NOT1 (N6952, N6943);
nor NOR2 (N6953, N6936, N5093);
not NOT1 (N6954, N6952);
and AND3 (N6955, N6920, N1664, N6317);
buf BUF1 (N6956, N6940);
xor XOR2 (N6957, N6956, N6867);
not NOT1 (N6958, N6937);
and AND4 (N6959, N6954, N6230, N3678, N1946);
nand NAND4 (N6960, N6955, N1080, N3953, N671);
and AND4 (N6961, N6960, N1619, N4595, N5700);
nor NOR2 (N6962, N6961, N1616);
or OR3 (N6963, N6950, N2346, N3972);
nor NOR3 (N6964, N6942, N2349, N1176);
xor XOR2 (N6965, N6948, N4447);
nand NAND2 (N6966, N6963, N2560);
nand NAND2 (N6967, N6964, N3489);
buf BUF1 (N6968, N6953);
xor XOR2 (N6969, N6968, N5950);
and AND4 (N6970, N6966, N6524, N2346, N1764);
nor NOR3 (N6971, N6970, N3749, N5033);
or OR2 (N6972, N6958, N6644);
not NOT1 (N6973, N6972);
or OR3 (N6974, N6947, N5557, N6757);
buf BUF1 (N6975, N6951);
not NOT1 (N6976, N6973);
nor NOR3 (N6977, N6962, N5200, N6047);
nand NAND2 (N6978, N6974, N4128);
xor XOR2 (N6979, N6969, N6925);
nand NAND4 (N6980, N6979, N2241, N3620, N1333);
not NOT1 (N6981, N6975);
nand NAND3 (N6982, N6957, N6629, N867);
nand NAND3 (N6983, N6977, N6959, N3527);
and AND4 (N6984, N6854, N2542, N2112, N561);
buf BUF1 (N6985, N6984);
buf BUF1 (N6986, N6965);
buf BUF1 (N6987, N6986);
or OR3 (N6988, N6982, N815, N6630);
or OR4 (N6989, N6978, N1478, N2372, N6128);
xor XOR2 (N6990, N6967, N2193);
nand NAND2 (N6991, N6981, N1676);
not NOT1 (N6992, N6976);
or OR3 (N6993, N6983, N1564, N4259);
and AND3 (N6994, N6990, N2351, N6555);
or OR2 (N6995, N6992, N3732);
buf BUF1 (N6996, N6993);
nand NAND4 (N6997, N6980, N26, N3177, N3759);
not NOT1 (N6998, N6997);
not NOT1 (N6999, N6996);
buf BUF1 (N7000, N6985);
or OR2 (N7001, N6991, N2456);
and AND4 (N7002, N6989, N5119, N1813, N4533);
and AND4 (N7003, N6988, N6119, N3186, N1956);
or OR3 (N7004, N7000, N4150, N6109);
not NOT1 (N7005, N6971);
and AND2 (N7006, N6995, N2119);
nand NAND4 (N7007, N7004, N3554, N127, N1416);
nand NAND2 (N7008, N6998, N929);
or OR4 (N7009, N7003, N2656, N4646, N6326);
buf BUF1 (N7010, N7006);
not NOT1 (N7011, N7001);
not NOT1 (N7012, N7005);
and AND4 (N7013, N6999, N2640, N1399, N6928);
not NOT1 (N7014, N6994);
buf BUF1 (N7015, N7014);
not NOT1 (N7016, N7015);
xor XOR2 (N7017, N6987, N4953);
xor XOR2 (N7018, N7007, N5020);
xor XOR2 (N7019, N7012, N2378);
or OR4 (N7020, N7017, N1205, N6719, N1085);
xor XOR2 (N7021, N7010, N6767);
buf BUF1 (N7022, N7016);
buf BUF1 (N7023, N7022);
or OR2 (N7024, N7020, N3741);
not NOT1 (N7025, N7019);
or OR2 (N7026, N7008, N5256);
nand NAND3 (N7027, N7011, N1926, N4025);
nand NAND4 (N7028, N7027, N4873, N4779, N2715);
nor NOR3 (N7029, N7024, N2801, N3787);
nor NOR3 (N7030, N7002, N6188, N6876);
and AND4 (N7031, N7025, N6736, N5250, N2517);
buf BUF1 (N7032, N7021);
nand NAND3 (N7033, N7031, N6651, N5911);
buf BUF1 (N7034, N7029);
nor NOR4 (N7035, N7032, N6678, N1385, N345);
buf BUF1 (N7036, N7009);
not NOT1 (N7037, N7018);
not NOT1 (N7038, N7035);
and AND4 (N7039, N7030, N405, N1775, N3319);
buf BUF1 (N7040, N7037);
xor XOR2 (N7041, N7033, N4112);
and AND4 (N7042, N7026, N460, N1125, N6800);
xor XOR2 (N7043, N7023, N6408);
and AND3 (N7044, N7043, N6774, N4427);
not NOT1 (N7045, N7039);
xor XOR2 (N7046, N7040, N1054);
and AND3 (N7047, N7028, N6188, N2311);
nand NAND3 (N7048, N7034, N7036, N1624);
xor XOR2 (N7049, N5345, N4193);
nand NAND2 (N7050, N7044, N2179);
nor NOR4 (N7051, N7050, N509, N5382, N6153);
xor XOR2 (N7052, N7047, N1687);
nor NOR2 (N7053, N7046, N4858);
and AND3 (N7054, N7045, N3216, N6786);
or OR3 (N7055, N7042, N998, N6600);
and AND2 (N7056, N7051, N3076);
or OR3 (N7057, N7049, N2308, N7047);
or OR2 (N7058, N7056, N3765);
or OR4 (N7059, N7038, N5869, N4359, N5246);
buf BUF1 (N7060, N7055);
not NOT1 (N7061, N7052);
nand NAND2 (N7062, N7058, N5012);
buf BUF1 (N7063, N7053);
not NOT1 (N7064, N7013);
or OR4 (N7065, N7048, N2674, N3454, N3317);
or OR3 (N7066, N7065, N2440, N4983);
nor NOR2 (N7067, N7061, N5142);
nand NAND2 (N7068, N7041, N6701);
nor NOR2 (N7069, N7054, N4126);
xor XOR2 (N7070, N7066, N4506);
or OR4 (N7071, N7069, N2264, N1375, N388);
and AND3 (N7072, N7063, N546, N5777);
nand NAND4 (N7073, N7067, N6463, N5032, N1570);
nand NAND3 (N7074, N7060, N1499, N1294);
buf BUF1 (N7075, N7068);
or OR4 (N7076, N7059, N303, N4556, N5564);
nand NAND2 (N7077, N7076, N3117);
not NOT1 (N7078, N7071);
nand NAND3 (N7079, N7078, N39, N3661);
nor NOR4 (N7080, N7057, N1764, N3207, N2660);
not NOT1 (N7081, N7074);
nand NAND4 (N7082, N7081, N2378, N5618, N1607);
nand NAND2 (N7083, N7073, N4724);
and AND2 (N7084, N7064, N6238);
or OR2 (N7085, N7079, N5351);
nor NOR4 (N7086, N7077, N4343, N6625, N2772);
nand NAND4 (N7087, N7080, N1605, N6543, N562);
nor NOR4 (N7088, N7086, N1456, N1206, N6182);
nand NAND4 (N7089, N7072, N3899, N4250, N2384);
not NOT1 (N7090, N7075);
buf BUF1 (N7091, N7088);
nand NAND4 (N7092, N7070, N6921, N5868, N1165);
not NOT1 (N7093, N7084);
nand NAND3 (N7094, N7085, N6540, N5729);
not NOT1 (N7095, N7089);
nor NOR4 (N7096, N7087, N6128, N2401, N739);
buf BUF1 (N7097, N7094);
or OR3 (N7098, N7082, N6612, N4630);
not NOT1 (N7099, N7092);
and AND3 (N7100, N7098, N6765, N3262);
buf BUF1 (N7101, N7091);
xor XOR2 (N7102, N7101, N5371);
nor NOR2 (N7103, N7100, N6130);
not NOT1 (N7104, N7097);
and AND4 (N7105, N7093, N5731, N1279, N3187);
and AND2 (N7106, N7062, N2119);
or OR4 (N7107, N7090, N4341, N3775, N4215);
nor NOR4 (N7108, N7095, N3240, N1440, N6527);
or OR2 (N7109, N7104, N2112);
buf BUF1 (N7110, N7103);
or OR4 (N7111, N7106, N1668, N2326, N6313);
buf BUF1 (N7112, N7105);
not NOT1 (N7113, N7108);
buf BUF1 (N7114, N7112);
not NOT1 (N7115, N7107);
nand NAND4 (N7116, N7109, N6637, N2683, N6283);
xor XOR2 (N7117, N7099, N1960);
xor XOR2 (N7118, N7113, N6996);
or OR4 (N7119, N7118, N1895, N5900, N4467);
nor NOR2 (N7120, N7102, N1324);
buf BUF1 (N7121, N7083);
not NOT1 (N7122, N7119);
buf BUF1 (N7123, N7096);
xor XOR2 (N7124, N7111, N6548);
buf BUF1 (N7125, N7117);
nand NAND3 (N7126, N7116, N4033, N4170);
nor NOR3 (N7127, N7121, N2726, N3493);
nor NOR2 (N7128, N7127, N4107);
and AND3 (N7129, N7124, N459, N4581);
nand NAND4 (N7130, N7115, N4188, N4687, N4371);
or OR4 (N7131, N7128, N1536, N3488, N2962);
nor NOR2 (N7132, N7120, N5527);
buf BUF1 (N7133, N7130);
or OR2 (N7134, N7125, N2440);
buf BUF1 (N7135, N7131);
xor XOR2 (N7136, N7110, N253);
xor XOR2 (N7137, N7123, N1494);
not NOT1 (N7138, N7132);
or OR3 (N7139, N7138, N6090, N4262);
not NOT1 (N7140, N7126);
and AND4 (N7141, N7136, N4773, N6570, N3873);
nor NOR2 (N7142, N7114, N5589);
nand NAND3 (N7143, N7122, N5765, N2945);
xor XOR2 (N7144, N7140, N6182);
buf BUF1 (N7145, N7137);
buf BUF1 (N7146, N7133);
nand NAND2 (N7147, N7141, N1670);
not NOT1 (N7148, N7139);
not NOT1 (N7149, N7134);
buf BUF1 (N7150, N7148);
or OR4 (N7151, N7150, N4345, N1709, N2455);
nor NOR4 (N7152, N7143, N6246, N4639, N392);
xor XOR2 (N7153, N7144, N2450);
and AND2 (N7154, N7151, N6450);
or OR4 (N7155, N7153, N1619, N439, N6647);
xor XOR2 (N7156, N7129, N3855);
or OR3 (N7157, N7147, N4302, N1405);
or OR2 (N7158, N7154, N4512);
not NOT1 (N7159, N7158);
or OR2 (N7160, N7145, N786);
not NOT1 (N7161, N7159);
and AND2 (N7162, N7157, N2929);
nor NOR4 (N7163, N7135, N2760, N7082, N4858);
nor NOR4 (N7164, N7155, N4632, N4867, N5805);
nor NOR2 (N7165, N7142, N6130);
and AND2 (N7166, N7146, N2144);
buf BUF1 (N7167, N7161);
xor XOR2 (N7168, N7152, N1189);
or OR4 (N7169, N7166, N3450, N3651, N1097);
nand NAND4 (N7170, N7169, N5593, N180, N3784);
nand NAND2 (N7171, N7160, N1187);
or OR2 (N7172, N7168, N5460);
or OR2 (N7173, N7171, N1595);
buf BUF1 (N7174, N7164);
xor XOR2 (N7175, N7170, N1932);
xor XOR2 (N7176, N7173, N1826);
and AND2 (N7177, N7165, N1082);
or OR2 (N7178, N7172, N3928);
and AND3 (N7179, N7163, N2427, N1810);
and AND4 (N7180, N7167, N5033, N6630, N59);
not NOT1 (N7181, N7177);
and AND2 (N7182, N7174, N1776);
not NOT1 (N7183, N7181);
or OR2 (N7184, N7182, N5678);
or OR4 (N7185, N7179, N4419, N5092, N1403);
not NOT1 (N7186, N7183);
nand NAND4 (N7187, N7156, N1917, N5512, N1125);
buf BUF1 (N7188, N7186);
buf BUF1 (N7189, N7184);
or OR3 (N7190, N7188, N6431, N2848);
not NOT1 (N7191, N7162);
nor NOR4 (N7192, N7178, N2164, N781, N269);
nand NAND2 (N7193, N7176, N2878);
not NOT1 (N7194, N7185);
xor XOR2 (N7195, N7194, N3577);
nand NAND2 (N7196, N7189, N1725);
not NOT1 (N7197, N7180);
nor NOR2 (N7198, N7196, N3654);
not NOT1 (N7199, N7195);
not NOT1 (N7200, N7199);
and AND4 (N7201, N7192, N4610, N469, N5574);
and AND3 (N7202, N7187, N2283, N773);
nor NOR2 (N7203, N7198, N1030);
buf BUF1 (N7204, N7200);
nor NOR2 (N7205, N7193, N1794);
xor XOR2 (N7206, N7197, N3628);
buf BUF1 (N7207, N7203);
nand NAND2 (N7208, N7201, N1891);
and AND3 (N7209, N7205, N4182, N2464);
and AND3 (N7210, N7207, N2905, N3109);
and AND4 (N7211, N7204, N1171, N4156, N3082);
nand NAND2 (N7212, N7175, N2993);
and AND2 (N7213, N7190, N338);
not NOT1 (N7214, N7212);
not NOT1 (N7215, N7208);
nor NOR3 (N7216, N7206, N1126, N5826);
xor XOR2 (N7217, N7216, N3647);
nor NOR2 (N7218, N7191, N1899);
not NOT1 (N7219, N7217);
buf BUF1 (N7220, N7214);
or OR2 (N7221, N7220, N223);
nand NAND2 (N7222, N7219, N6398);
or OR4 (N7223, N7211, N4933, N6048, N3352);
and AND2 (N7224, N7209, N2582);
and AND4 (N7225, N7222, N6805, N1536, N5061);
buf BUF1 (N7226, N7149);
or OR3 (N7227, N7213, N2532, N5870);
nand NAND2 (N7228, N7215, N3738);
not NOT1 (N7229, N7221);
not NOT1 (N7230, N7218);
nor NOR2 (N7231, N7229, N1681);
buf BUF1 (N7232, N7230);
and AND2 (N7233, N7225, N5432);
nor NOR4 (N7234, N7227, N2841, N709, N7110);
and AND2 (N7235, N7233, N6602);
buf BUF1 (N7236, N7234);
or OR2 (N7237, N7210, N463);
not NOT1 (N7238, N7235);
and AND4 (N7239, N7202, N6031, N7194, N1640);
nor NOR3 (N7240, N7226, N3280, N2699);
nand NAND2 (N7241, N7239, N4313);
xor XOR2 (N7242, N7231, N5033);
not NOT1 (N7243, N7236);
not NOT1 (N7244, N7243);
xor XOR2 (N7245, N7238, N6770);
and AND3 (N7246, N7244, N7047, N446);
or OR2 (N7247, N7237, N6027);
buf BUF1 (N7248, N7228);
and AND3 (N7249, N7247, N3706, N4118);
buf BUF1 (N7250, N7240);
and AND2 (N7251, N7242, N1408);
buf BUF1 (N7252, N7232);
xor XOR2 (N7253, N7241, N4152);
not NOT1 (N7254, N7223);
not NOT1 (N7255, N7224);
not NOT1 (N7256, N7252);
xor XOR2 (N7257, N7253, N6287);
xor XOR2 (N7258, N7257, N1211);
or OR2 (N7259, N7258, N630);
not NOT1 (N7260, N7248);
nand NAND4 (N7261, N7255, N4995, N1138, N3347);
xor XOR2 (N7262, N7246, N4755);
not NOT1 (N7263, N7249);
not NOT1 (N7264, N7261);
xor XOR2 (N7265, N7254, N4250);
or OR4 (N7266, N7251, N365, N4467, N1209);
not NOT1 (N7267, N7262);
nand NAND2 (N7268, N7259, N1161);
xor XOR2 (N7269, N7268, N6097);
xor XOR2 (N7270, N7269, N832);
nor NOR4 (N7271, N7260, N6438, N4260, N446);
and AND2 (N7272, N7266, N4744);
nor NOR2 (N7273, N7245, N3097);
or OR4 (N7274, N7263, N522, N1589, N1198);
not NOT1 (N7275, N7272);
nand NAND4 (N7276, N7275, N4907, N3411, N1138);
nor NOR2 (N7277, N7273, N989);
buf BUF1 (N7278, N7276);
nand NAND3 (N7279, N7270, N388, N5143);
xor XOR2 (N7280, N7274, N3766);
and AND2 (N7281, N7280, N6754);
and AND2 (N7282, N7267, N4978);
and AND2 (N7283, N7279, N3762);
and AND3 (N7284, N7278, N3034, N868);
and AND4 (N7285, N7282, N388, N2802, N3672);
buf BUF1 (N7286, N7285);
xor XOR2 (N7287, N7284, N185);
buf BUF1 (N7288, N7265);
and AND4 (N7289, N7271, N5925, N4633, N1620);
not NOT1 (N7290, N7283);
nor NOR2 (N7291, N7250, N931);
or OR4 (N7292, N7277, N6174, N5706, N2930);
buf BUF1 (N7293, N7281);
xor XOR2 (N7294, N7286, N947);
and AND2 (N7295, N7287, N597);
or OR2 (N7296, N7290, N4771);
buf BUF1 (N7297, N7256);
nand NAND4 (N7298, N7297, N3982, N2251, N4053);
and AND2 (N7299, N7288, N3109);
nand NAND3 (N7300, N7298, N4631, N3501);
and AND2 (N7301, N7299, N4550);
buf BUF1 (N7302, N7264);
nand NAND3 (N7303, N7296, N4528, N2647);
xor XOR2 (N7304, N7294, N5637);
buf BUF1 (N7305, N7291);
nand NAND4 (N7306, N7301, N7275, N1890, N6582);
nor NOR4 (N7307, N7303, N268, N1047, N882);
nor NOR2 (N7308, N7300, N1203);
buf BUF1 (N7309, N7302);
xor XOR2 (N7310, N7308, N758);
or OR3 (N7311, N7293, N1059, N635);
nand NAND3 (N7312, N7309, N1985, N4204);
buf BUF1 (N7313, N7304);
nor NOR3 (N7314, N7292, N6353, N1925);
or OR4 (N7315, N7307, N6487, N3792, N371);
not NOT1 (N7316, N7295);
not NOT1 (N7317, N7314);
not NOT1 (N7318, N7289);
not NOT1 (N7319, N7305);
buf BUF1 (N7320, N7306);
nor NOR3 (N7321, N7310, N4601, N5172);
nand NAND2 (N7322, N7319, N4214);
not NOT1 (N7323, N7316);
or OR3 (N7324, N7318, N1442, N1244);
or OR2 (N7325, N7311, N6477);
nor NOR4 (N7326, N7325, N1522, N2148, N1422);
xor XOR2 (N7327, N7323, N4588);
xor XOR2 (N7328, N7315, N3289);
or OR2 (N7329, N7322, N566);
buf BUF1 (N7330, N7328);
buf BUF1 (N7331, N7327);
xor XOR2 (N7332, N7324, N2220);
xor XOR2 (N7333, N7313, N3941);
not NOT1 (N7334, N7317);
or OR2 (N7335, N7334, N6500);
buf BUF1 (N7336, N7326);
buf BUF1 (N7337, N7332);
nor NOR2 (N7338, N7331, N3768);
or OR3 (N7339, N7330, N3030, N3145);
xor XOR2 (N7340, N7336, N6155);
not NOT1 (N7341, N7339);
buf BUF1 (N7342, N7333);
not NOT1 (N7343, N7338);
buf BUF1 (N7344, N7312);
nor NOR2 (N7345, N7343, N2416);
buf BUF1 (N7346, N7321);
or OR3 (N7347, N7341, N3274, N1005);
nand NAND4 (N7348, N7344, N4254, N2378, N6492);
xor XOR2 (N7349, N7345, N1236);
not NOT1 (N7350, N7342);
xor XOR2 (N7351, N7320, N6732);
or OR2 (N7352, N7350, N3991);
nand NAND3 (N7353, N7351, N1115, N1528);
buf BUF1 (N7354, N7348);
nand NAND4 (N7355, N7335, N6850, N2184, N5365);
xor XOR2 (N7356, N7349, N3870);
and AND2 (N7357, N7337, N539);
not NOT1 (N7358, N7356);
buf BUF1 (N7359, N7357);
nor NOR4 (N7360, N7359, N1955, N312, N6131);
nand NAND2 (N7361, N7347, N2584);
and AND2 (N7362, N7353, N5196);
buf BUF1 (N7363, N7358);
buf BUF1 (N7364, N7362);
nand NAND2 (N7365, N7340, N3154);
and AND3 (N7366, N7365, N1446, N1358);
nand NAND3 (N7367, N7329, N6055, N5249);
nand NAND3 (N7368, N7346, N6416, N6951);
nor NOR3 (N7369, N7360, N487, N6451);
or OR2 (N7370, N7352, N2122);
xor XOR2 (N7371, N7370, N2508);
or OR2 (N7372, N7367, N997);
xor XOR2 (N7373, N7355, N6558);
nor NOR2 (N7374, N7368, N3779);
xor XOR2 (N7375, N7372, N2351);
buf BUF1 (N7376, N7363);
nor NOR3 (N7377, N7361, N1406, N4395);
and AND2 (N7378, N7354, N3500);
not NOT1 (N7379, N7373);
nor NOR2 (N7380, N7371, N2666);
or OR3 (N7381, N7369, N3692, N6459);
not NOT1 (N7382, N7364);
xor XOR2 (N7383, N7366, N2132);
not NOT1 (N7384, N7381);
not NOT1 (N7385, N7383);
nand NAND3 (N7386, N7380, N1823, N6550);
nand NAND2 (N7387, N7382, N2565);
nor NOR3 (N7388, N7377, N5386, N5215);
nor NOR4 (N7389, N7379, N2493, N5902, N7048);
nor NOR4 (N7390, N7374, N3150, N1235, N6640);
nand NAND3 (N7391, N7385, N4058, N7343);
nand NAND4 (N7392, N7389, N1396, N3777, N1113);
not NOT1 (N7393, N7388);
nand NAND3 (N7394, N7384, N4030, N140);
buf BUF1 (N7395, N7386);
nor NOR2 (N7396, N7387, N5835);
nand NAND4 (N7397, N7396, N4936, N6, N105);
or OR2 (N7398, N7390, N4643);
xor XOR2 (N7399, N7375, N3559);
or OR2 (N7400, N7393, N2506);
nor NOR4 (N7401, N7376, N6020, N192, N5230);
nor NOR3 (N7402, N7378, N233, N2012);
not NOT1 (N7403, N7394);
nor NOR2 (N7404, N7398, N1922);
buf BUF1 (N7405, N7401);
nor NOR2 (N7406, N7404, N5748);
or OR4 (N7407, N7402, N3934, N1393, N2890);
nor NOR2 (N7408, N7392, N7183);
buf BUF1 (N7409, N7391);
nor NOR4 (N7410, N7407, N559, N713, N6355);
and AND4 (N7411, N7399, N689, N375, N4607);
not NOT1 (N7412, N7406);
buf BUF1 (N7413, N7408);
xor XOR2 (N7414, N7397, N1941);
nand NAND3 (N7415, N7400, N3693, N2535);
nor NOR2 (N7416, N7413, N6900);
and AND2 (N7417, N7416, N6211);
not NOT1 (N7418, N7410);
nand NAND2 (N7419, N7412, N730);
xor XOR2 (N7420, N7395, N2693);
buf BUF1 (N7421, N7409);
nand NAND2 (N7422, N7415, N1460);
and AND2 (N7423, N7417, N2188);
nand NAND4 (N7424, N7418, N4334, N1611, N2147);
buf BUF1 (N7425, N7421);
nor NOR2 (N7426, N7405, N2053);
nor NOR4 (N7427, N7423, N2535, N4115, N54);
nand NAND3 (N7428, N7419, N1469, N5178);
nor NOR2 (N7429, N7411, N3670);
and AND3 (N7430, N7427, N1170, N3170);
not NOT1 (N7431, N7422);
and AND3 (N7432, N7431, N7190, N218);
nor NOR4 (N7433, N7429, N3313, N2975, N5562);
or OR2 (N7434, N7424, N4119);
buf BUF1 (N7435, N7430);
buf BUF1 (N7436, N7426);
or OR2 (N7437, N7436, N2973);
buf BUF1 (N7438, N7433);
buf BUF1 (N7439, N7414);
and AND4 (N7440, N7425, N6276, N1492, N6232);
not NOT1 (N7441, N7420);
or OR4 (N7442, N7439, N7330, N1254, N3275);
and AND2 (N7443, N7403, N6183);
buf BUF1 (N7444, N7432);
nand NAND3 (N7445, N7434, N3686, N4949);
buf BUF1 (N7446, N7445);
nor NOR2 (N7447, N7435, N5316);
and AND2 (N7448, N7437, N969);
nand NAND2 (N7449, N7448, N642);
nand NAND3 (N7450, N7444, N2050, N4033);
nand NAND2 (N7451, N7438, N4153);
and AND3 (N7452, N7443, N5420, N2355);
or OR3 (N7453, N7441, N5925, N5363);
buf BUF1 (N7454, N7442);
buf BUF1 (N7455, N7453);
or OR2 (N7456, N7452, N5995);
and AND4 (N7457, N7450, N6741, N7272, N331);
not NOT1 (N7458, N7455);
nor NOR3 (N7459, N7454, N7128, N5106);
not NOT1 (N7460, N7440);
and AND3 (N7461, N7447, N7437, N4805);
or OR4 (N7462, N7457, N5325, N2285, N3695);
nor NOR2 (N7463, N7456, N4605);
not NOT1 (N7464, N7446);
nand NAND2 (N7465, N7451, N5016);
or OR4 (N7466, N7458, N7223, N6027, N2418);
xor XOR2 (N7467, N7460, N2512);
buf BUF1 (N7468, N7466);
nor NOR3 (N7469, N7461, N6677, N5668);
buf BUF1 (N7470, N7464);
not NOT1 (N7471, N7463);
or OR2 (N7472, N7467, N1529);
not NOT1 (N7473, N7462);
or OR3 (N7474, N7465, N1715, N1673);
xor XOR2 (N7475, N7474, N5120);
nand NAND4 (N7476, N7473, N524, N3762, N3392);
nor NOR3 (N7477, N7428, N5349, N3924);
not NOT1 (N7478, N7472);
not NOT1 (N7479, N7477);
xor XOR2 (N7480, N7468, N252);
buf BUF1 (N7481, N7469);
xor XOR2 (N7482, N7449, N3591);
and AND4 (N7483, N7482, N299, N6752, N1680);
nor NOR3 (N7484, N7459, N2673, N6285);
nor NOR3 (N7485, N7471, N4933, N3676);
nor NOR3 (N7486, N7478, N915, N1487);
nand NAND2 (N7487, N7479, N4804);
and AND3 (N7488, N7476, N6870, N6918);
and AND3 (N7489, N7486, N6672, N2340);
nor NOR4 (N7490, N7483, N1342, N6582, N6894);
xor XOR2 (N7491, N7485, N3550);
nor NOR4 (N7492, N7481, N1237, N1783, N4438);
not NOT1 (N7493, N7489);
nand NAND3 (N7494, N7484, N4327, N1350);
nor NOR4 (N7495, N7491, N6806, N6955, N1669);
nor NOR2 (N7496, N7487, N7213);
or OR3 (N7497, N7490, N424, N3310);
not NOT1 (N7498, N7470);
xor XOR2 (N7499, N7496, N976);
buf BUF1 (N7500, N7493);
xor XOR2 (N7501, N7494, N7472);
nor NOR4 (N7502, N7495, N3000, N3045, N5461);
not NOT1 (N7503, N7502);
or OR4 (N7504, N7475, N743, N480, N2425);
and AND2 (N7505, N7498, N5466);
not NOT1 (N7506, N7501);
xor XOR2 (N7507, N7505, N5557);
not NOT1 (N7508, N7500);
buf BUF1 (N7509, N7492);
or OR4 (N7510, N7480, N6044, N3683, N1216);
not NOT1 (N7511, N7488);
not NOT1 (N7512, N7510);
or OR3 (N7513, N7508, N5256, N4100);
buf BUF1 (N7514, N7503);
nor NOR4 (N7515, N7497, N1199, N2254, N5493);
xor XOR2 (N7516, N7511, N6187);
buf BUF1 (N7517, N7514);
not NOT1 (N7518, N7504);
xor XOR2 (N7519, N7506, N226);
buf BUF1 (N7520, N7517);
nor NOR3 (N7521, N7518, N72, N1649);
xor XOR2 (N7522, N7507, N3560);
and AND3 (N7523, N7499, N4937, N6783);
nand NAND4 (N7524, N7513, N1834, N7350, N5132);
not NOT1 (N7525, N7523);
or OR4 (N7526, N7525, N418, N4294, N6807);
not NOT1 (N7527, N7515);
xor XOR2 (N7528, N7521, N5902);
nor NOR3 (N7529, N7520, N3025, N1506);
nor NOR2 (N7530, N7526, N2253);
buf BUF1 (N7531, N7527);
or OR4 (N7532, N7519, N307, N5010, N4499);
nor NOR3 (N7533, N7516, N7516, N1632);
and AND2 (N7534, N7530, N7095);
buf BUF1 (N7535, N7528);
not NOT1 (N7536, N7509);
not NOT1 (N7537, N7533);
and AND3 (N7538, N7537, N2265, N1610);
not NOT1 (N7539, N7529);
nand NAND2 (N7540, N7538, N4607);
or OR4 (N7541, N7540, N4369, N4328, N91);
not NOT1 (N7542, N7522);
or OR2 (N7543, N7536, N4119);
nor NOR2 (N7544, N7539, N2040);
not NOT1 (N7545, N7544);
nand NAND4 (N7546, N7535, N792, N6919, N4550);
buf BUF1 (N7547, N7545);
buf BUF1 (N7548, N7532);
xor XOR2 (N7549, N7524, N991);
and AND3 (N7550, N7512, N2609, N1256);
nand NAND2 (N7551, N7548, N4314);
nor NOR4 (N7552, N7542, N1934, N1534, N1418);
or OR3 (N7553, N7541, N4434, N2160);
and AND2 (N7554, N7546, N5892);
buf BUF1 (N7555, N7543);
and AND4 (N7556, N7550, N6331, N4739, N3804);
or OR2 (N7557, N7531, N7464);
buf BUF1 (N7558, N7554);
nor NOR3 (N7559, N7555, N5943, N2264);
not NOT1 (N7560, N7559);
xor XOR2 (N7561, N7549, N5692);
buf BUF1 (N7562, N7534);
and AND2 (N7563, N7547, N1874);
nor NOR4 (N7564, N7557, N7114, N4718, N2018);
or OR3 (N7565, N7553, N7450, N7533);
nor NOR4 (N7566, N7563, N2255, N2850, N4409);
xor XOR2 (N7567, N7562, N6902);
nand NAND3 (N7568, N7552, N7413, N5277);
buf BUF1 (N7569, N7561);
xor XOR2 (N7570, N7568, N4188);
and AND4 (N7571, N7569, N3490, N5506, N1315);
xor XOR2 (N7572, N7560, N4301);
buf BUF1 (N7573, N7565);
nand NAND2 (N7574, N7556, N918);
nor NOR2 (N7575, N7571, N4099);
buf BUF1 (N7576, N7570);
buf BUF1 (N7577, N7572);
and AND2 (N7578, N7564, N7569);
or OR3 (N7579, N7576, N678, N5143);
not NOT1 (N7580, N7578);
and AND2 (N7581, N7573, N7575);
and AND3 (N7582, N5670, N2993, N3665);
or OR3 (N7583, N7577, N6905, N2594);
not NOT1 (N7584, N7580);
and AND4 (N7585, N7584, N6170, N571, N1601);
xor XOR2 (N7586, N7583, N6221);
buf BUF1 (N7587, N7582);
not NOT1 (N7588, N7551);
nor NOR3 (N7589, N7567, N4315, N7350);
and AND4 (N7590, N7589, N1752, N7066, N46);
nor NOR4 (N7591, N7588, N1590, N138, N1436);
and AND3 (N7592, N7566, N1048, N2046);
xor XOR2 (N7593, N7586, N6228);
or OR4 (N7594, N7592, N3303, N541, N2156);
nor NOR3 (N7595, N7591, N5141, N714);
buf BUF1 (N7596, N7590);
and AND4 (N7597, N7585, N1223, N7245, N3885);
or OR3 (N7598, N7593, N3706, N6177);
buf BUF1 (N7599, N7587);
and AND2 (N7600, N7597, N6372);
or OR4 (N7601, N7594, N3967, N1972, N2486);
or OR4 (N7602, N7598, N841, N4721, N4015);
nor NOR3 (N7603, N7600, N2543, N6302);
xor XOR2 (N7604, N7558, N4297);
and AND4 (N7605, N7581, N746, N2625, N5801);
buf BUF1 (N7606, N7601);
nand NAND2 (N7607, N7599, N3477);
nor NOR4 (N7608, N7602, N349, N4024, N5162);
nand NAND4 (N7609, N7606, N5580, N5679, N817);
and AND3 (N7610, N7605, N6535, N1849);
not NOT1 (N7611, N7609);
nand NAND2 (N7612, N7596, N6912);
buf BUF1 (N7613, N7608);
not NOT1 (N7614, N7579);
or OR2 (N7615, N7611, N1892);
not NOT1 (N7616, N7607);
not NOT1 (N7617, N7610);
or OR2 (N7618, N7603, N5564);
nand NAND2 (N7619, N7616, N3425);
or OR4 (N7620, N7613, N3053, N6778, N7307);
not NOT1 (N7621, N7574);
and AND3 (N7622, N7604, N434, N5521);
nand NAND4 (N7623, N7614, N4227, N2060, N6095);
buf BUF1 (N7624, N7623);
or OR4 (N7625, N7595, N7347, N5112, N2330);
nand NAND2 (N7626, N7625, N948);
not NOT1 (N7627, N7615);
xor XOR2 (N7628, N7618, N1818);
nor NOR2 (N7629, N7619, N998);
xor XOR2 (N7630, N7617, N1002);
and AND2 (N7631, N7612, N3176);
xor XOR2 (N7632, N7627, N1648);
xor XOR2 (N7633, N7620, N3737);
nand NAND3 (N7634, N7633, N3716, N4657);
xor XOR2 (N7635, N7621, N2248);
not NOT1 (N7636, N7635);
or OR2 (N7637, N7632, N5564);
nor NOR3 (N7638, N7630, N383, N7532);
or OR4 (N7639, N7634, N4463, N3104, N4835);
and AND4 (N7640, N7626, N2291, N894, N379);
nor NOR2 (N7641, N7631, N6159);
and AND4 (N7642, N7641, N2431, N2944, N6342);
nand NAND3 (N7643, N7637, N21, N3155);
or OR2 (N7644, N7624, N6337);
or OR3 (N7645, N7636, N5231, N6186);
buf BUF1 (N7646, N7643);
and AND4 (N7647, N7646, N1223, N2907, N6653);
nor NOR4 (N7648, N7629, N7273, N3830, N3718);
and AND4 (N7649, N7645, N6257, N4818, N3674);
and AND3 (N7650, N7628, N6742, N610);
and AND4 (N7651, N7649, N4328, N5676, N7146);
xor XOR2 (N7652, N7644, N4272);
or OR4 (N7653, N7648, N64, N6264, N3311);
or OR3 (N7654, N7639, N4018, N638);
and AND2 (N7655, N7651, N4314);
xor XOR2 (N7656, N7655, N1001);
buf BUF1 (N7657, N7642);
buf BUF1 (N7658, N7640);
and AND4 (N7659, N7650, N1597, N942, N5351);
xor XOR2 (N7660, N7658, N5438);
nor NOR4 (N7661, N7654, N2647, N5698, N75);
xor XOR2 (N7662, N7653, N6644);
and AND2 (N7663, N7652, N5443);
buf BUF1 (N7664, N7661);
nand NAND2 (N7665, N7622, N1893);
xor XOR2 (N7666, N7663, N5477);
buf BUF1 (N7667, N7660);
buf BUF1 (N7668, N7664);
nand NAND4 (N7669, N7666, N3683, N2272, N5927);
nand NAND3 (N7670, N7638, N1230, N6718);
buf BUF1 (N7671, N7662);
nor NOR2 (N7672, N7647, N900);
buf BUF1 (N7673, N7671);
or OR2 (N7674, N7659, N2650);
xor XOR2 (N7675, N7657, N5693);
or OR2 (N7676, N7656, N1689);
not NOT1 (N7677, N7668);
not NOT1 (N7678, N7675);
buf BUF1 (N7679, N7674);
not NOT1 (N7680, N7676);
nand NAND4 (N7681, N7665, N5630, N2701, N5236);
nand NAND3 (N7682, N7673, N7466, N2098);
buf BUF1 (N7683, N7670);
buf BUF1 (N7684, N7679);
buf BUF1 (N7685, N7678);
nor NOR3 (N7686, N7677, N4170, N4788);
nand NAND4 (N7687, N7684, N2851, N5541, N6574);
and AND3 (N7688, N7669, N5296, N6532);
nand NAND4 (N7689, N7681, N6870, N4627, N1016);
and AND4 (N7690, N7687, N5130, N1706, N7492);
or OR4 (N7691, N7689, N3063, N1073, N5795);
nand NAND2 (N7692, N7686, N5109);
buf BUF1 (N7693, N7680);
not NOT1 (N7694, N7667);
nand NAND2 (N7695, N7692, N782);
xor XOR2 (N7696, N7682, N2881);
xor XOR2 (N7697, N7695, N5228);
nor NOR4 (N7698, N7697, N2276, N7679, N4962);
nand NAND3 (N7699, N7693, N1631, N1603);
nand NAND3 (N7700, N7685, N2699, N1023);
nand NAND4 (N7701, N7691, N4128, N2346, N6049);
buf BUF1 (N7702, N7694);
not NOT1 (N7703, N7688);
nor NOR3 (N7704, N7696, N159, N4667);
or OR4 (N7705, N7700, N7376, N4030, N6505);
xor XOR2 (N7706, N7690, N7091);
xor XOR2 (N7707, N7703, N3014);
nand NAND3 (N7708, N7704, N5990, N7291);
xor XOR2 (N7709, N7708, N3300);
buf BUF1 (N7710, N7702);
not NOT1 (N7711, N7683);
not NOT1 (N7712, N7699);
and AND2 (N7713, N7710, N1246);
and AND2 (N7714, N7705, N3299);
or OR2 (N7715, N7711, N3893);
or OR4 (N7716, N7706, N836, N5228, N445);
not NOT1 (N7717, N7713);
nand NAND4 (N7718, N7701, N240, N6991, N6280);
not NOT1 (N7719, N7717);
xor XOR2 (N7720, N7714, N6239);
buf BUF1 (N7721, N7718);
not NOT1 (N7722, N7707);
not NOT1 (N7723, N7720);
nand NAND4 (N7724, N7722, N1497, N5431, N429);
not NOT1 (N7725, N7672);
buf BUF1 (N7726, N7721);
xor XOR2 (N7727, N7723, N2574);
nand NAND4 (N7728, N7712, N1856, N1293, N3974);
not NOT1 (N7729, N7716);
buf BUF1 (N7730, N7728);
or OR4 (N7731, N7698, N5168, N5665, N1845);
not NOT1 (N7732, N7719);
nand NAND3 (N7733, N7709, N23, N5081);
and AND3 (N7734, N7724, N3166, N4474);
xor XOR2 (N7735, N7732, N1165);
and AND3 (N7736, N7733, N4416, N4142);
nor NOR4 (N7737, N7727, N4790, N7112, N3413);
buf BUF1 (N7738, N7737);
nor NOR2 (N7739, N7730, N7337);
xor XOR2 (N7740, N7715, N3616);
and AND4 (N7741, N7735, N2084, N6714, N5361);
nand NAND2 (N7742, N7726, N2220);
nor NOR3 (N7743, N7738, N3838, N382);
not NOT1 (N7744, N7742);
xor XOR2 (N7745, N7744, N1711);
nor NOR4 (N7746, N7731, N7283, N7566, N6925);
nand NAND3 (N7747, N7725, N7180, N555);
and AND4 (N7748, N7741, N5146, N6926, N5960);
buf BUF1 (N7749, N7748);
not NOT1 (N7750, N7749);
and AND3 (N7751, N7740, N2182, N860);
xor XOR2 (N7752, N7743, N7069);
and AND4 (N7753, N7734, N1880, N4069, N2296);
not NOT1 (N7754, N7753);
and AND3 (N7755, N7736, N4964, N702);
xor XOR2 (N7756, N7755, N4647);
nand NAND3 (N7757, N7756, N2388, N6175);
xor XOR2 (N7758, N7751, N2708);
or OR2 (N7759, N7739, N7313);
buf BUF1 (N7760, N7759);
and AND2 (N7761, N7752, N5954);
xor XOR2 (N7762, N7754, N3053);
nand NAND2 (N7763, N7746, N5184);
nand NAND3 (N7764, N7761, N4453, N6432);
buf BUF1 (N7765, N7747);
or OR2 (N7766, N7729, N3477);
not NOT1 (N7767, N7765);
nor NOR2 (N7768, N7757, N5321);
or OR4 (N7769, N7768, N4391, N2037, N1289);
not NOT1 (N7770, N7758);
nand NAND2 (N7771, N7769, N3319);
or OR2 (N7772, N7766, N884);
nor NOR2 (N7773, N7745, N1272);
buf BUF1 (N7774, N7763);
and AND4 (N7775, N7760, N4481, N3407, N6562);
not NOT1 (N7776, N7750);
buf BUF1 (N7777, N7775);
or OR4 (N7778, N7767, N2375, N6566, N1587);
not NOT1 (N7779, N7774);
nor NOR3 (N7780, N7770, N2384, N2397);
buf BUF1 (N7781, N7777);
not NOT1 (N7782, N7764);
nor NOR4 (N7783, N7772, N1439, N6105, N5174);
and AND4 (N7784, N7779, N5784, N7312, N6334);
nor NOR3 (N7785, N7773, N4499, N612);
not NOT1 (N7786, N7762);
nor NOR2 (N7787, N7785, N4812);
buf BUF1 (N7788, N7771);
not NOT1 (N7789, N7781);
xor XOR2 (N7790, N7780, N400);
and AND3 (N7791, N7776, N4899, N3541);
nand NAND4 (N7792, N7789, N1458, N6274, N7710);
or OR2 (N7793, N7783, N7574);
or OR2 (N7794, N7791, N5587);
xor XOR2 (N7795, N7790, N787);
xor XOR2 (N7796, N7794, N2504);
buf BUF1 (N7797, N7792);
not NOT1 (N7798, N7797);
buf BUF1 (N7799, N7786);
and AND2 (N7800, N7782, N6222);
or OR3 (N7801, N7793, N7628, N3174);
xor XOR2 (N7802, N7795, N1989);
not NOT1 (N7803, N7787);
nor NOR4 (N7804, N7799, N7516, N5864, N6357);
xor XOR2 (N7805, N7778, N4351);
nor NOR2 (N7806, N7802, N5682);
not NOT1 (N7807, N7803);
buf BUF1 (N7808, N7801);
nor NOR2 (N7809, N7807, N258);
xor XOR2 (N7810, N7808, N3430);
xor XOR2 (N7811, N7798, N7042);
nor NOR4 (N7812, N7810, N3160, N858, N2110);
or OR3 (N7813, N7806, N1856, N5055);
or OR3 (N7814, N7811, N4886, N6105);
or OR4 (N7815, N7800, N5432, N168, N1612);
buf BUF1 (N7816, N7788);
xor XOR2 (N7817, N7816, N5175);
buf BUF1 (N7818, N7815);
buf BUF1 (N7819, N7818);
not NOT1 (N7820, N7805);
xor XOR2 (N7821, N7812, N4978);
nor NOR3 (N7822, N7819, N6042, N1234);
or OR4 (N7823, N7813, N5149, N234, N605);
xor XOR2 (N7824, N7809, N4051);
nand NAND4 (N7825, N7796, N213, N6097, N1098);
not NOT1 (N7826, N7824);
nor NOR2 (N7827, N7822, N5846);
xor XOR2 (N7828, N7804, N7130);
nand NAND3 (N7829, N7814, N3832, N2503);
not NOT1 (N7830, N7826);
nand NAND3 (N7831, N7825, N5555, N2490);
buf BUF1 (N7832, N7830);
nor NOR4 (N7833, N7817, N6082, N4686, N3553);
not NOT1 (N7834, N7827);
or OR3 (N7835, N7834, N2595, N2461);
or OR4 (N7836, N7829, N5851, N741, N6880);
buf BUF1 (N7837, N7821);
nor NOR4 (N7838, N7833, N1037, N3092, N4923);
buf BUF1 (N7839, N7823);
and AND4 (N7840, N7838, N2278, N6860, N6694);
not NOT1 (N7841, N7832);
not NOT1 (N7842, N7828);
or OR3 (N7843, N7839, N5073, N679);
not NOT1 (N7844, N7835);
xor XOR2 (N7845, N7820, N6653);
and AND4 (N7846, N7837, N4346, N4666, N6599);
or OR3 (N7847, N7844, N3862, N5704);
nand NAND3 (N7848, N7784, N5563, N3660);
buf BUF1 (N7849, N7841);
buf BUF1 (N7850, N7836);
or OR4 (N7851, N7848, N7416, N4269, N3033);
buf BUF1 (N7852, N7842);
xor XOR2 (N7853, N7831, N2855);
nand NAND2 (N7854, N7851, N5371);
xor XOR2 (N7855, N7852, N6316);
and AND2 (N7856, N7840, N5670);
and AND2 (N7857, N7853, N2655);
nand NAND3 (N7858, N7847, N5158, N7631);
nor NOR3 (N7859, N7857, N696, N1696);
nand NAND4 (N7860, N7845, N307, N4516, N2022);
and AND3 (N7861, N7850, N170, N1950);
nor NOR4 (N7862, N7849, N2306, N3660, N7814);
and AND3 (N7863, N7843, N419, N2253);
not NOT1 (N7864, N7858);
buf BUF1 (N7865, N7855);
xor XOR2 (N7866, N7854, N1150);
xor XOR2 (N7867, N7859, N3013);
xor XOR2 (N7868, N7846, N1308);
xor XOR2 (N7869, N7860, N4774);
and AND2 (N7870, N7865, N5841);
nor NOR2 (N7871, N7867, N6341);
xor XOR2 (N7872, N7866, N4910);
xor XOR2 (N7873, N7869, N1139);
and AND2 (N7874, N7868, N1733);
not NOT1 (N7875, N7861);
not NOT1 (N7876, N7873);
buf BUF1 (N7877, N7856);
not NOT1 (N7878, N7864);
nand NAND3 (N7879, N7876, N159, N5813);
buf BUF1 (N7880, N7875);
and AND2 (N7881, N7879, N5618);
nand NAND4 (N7882, N7877, N5576, N2159, N5623);
or OR2 (N7883, N7878, N7379);
and AND3 (N7884, N7881, N3887, N1074);
xor XOR2 (N7885, N7883, N5092);
or OR2 (N7886, N7880, N1404);
nand NAND2 (N7887, N7886, N1525);
nor NOR3 (N7888, N7872, N5188, N885);
nor NOR3 (N7889, N7882, N4124, N3719);
and AND2 (N7890, N7888, N2804);
nor NOR4 (N7891, N7863, N6983, N4680, N6406);
not NOT1 (N7892, N7891);
not NOT1 (N7893, N7892);
not NOT1 (N7894, N7893);
xor XOR2 (N7895, N7862, N463);
not NOT1 (N7896, N7890);
buf BUF1 (N7897, N7871);
and AND3 (N7898, N7896, N560, N3204);
buf BUF1 (N7899, N7894);
and AND4 (N7900, N7874, N6913, N4222, N1099);
buf BUF1 (N7901, N7884);
not NOT1 (N7902, N7889);
nand NAND3 (N7903, N7902, N5307, N7484);
nand NAND3 (N7904, N7887, N2210, N1615);
nor NOR2 (N7905, N7895, N5299);
or OR4 (N7906, N7897, N468, N5331, N7366);
not NOT1 (N7907, N7903);
buf BUF1 (N7908, N7885);
nand NAND2 (N7909, N7899, N5730);
or OR2 (N7910, N7907, N7837);
or OR2 (N7911, N7898, N2978);
xor XOR2 (N7912, N7908, N1816);
and AND2 (N7913, N7910, N6969);
nand NAND2 (N7914, N7901, N2278);
and AND4 (N7915, N7911, N6080, N4133, N6328);
and AND2 (N7916, N7906, N3179);
or OR3 (N7917, N7870, N4018, N722);
nand NAND4 (N7918, N7909, N5865, N6145, N4304);
nand NAND4 (N7919, N7905, N3010, N4527, N7804);
buf BUF1 (N7920, N7918);
xor XOR2 (N7921, N7920, N3230);
buf BUF1 (N7922, N7917);
buf BUF1 (N7923, N7912);
and AND3 (N7924, N7904, N4438, N1666);
nor NOR3 (N7925, N7924, N246, N390);
and AND4 (N7926, N7915, N198, N795, N6625);
nor NOR2 (N7927, N7900, N3036);
nor NOR4 (N7928, N7926, N2585, N5012, N6192);
not NOT1 (N7929, N7913);
buf BUF1 (N7930, N7922);
buf BUF1 (N7931, N7925);
nor NOR3 (N7932, N7928, N2860, N2938);
nor NOR2 (N7933, N7916, N1581);
not NOT1 (N7934, N7923);
nand NAND3 (N7935, N7931, N6312, N2934);
or OR4 (N7936, N7935, N2926, N3740, N6855);
nand NAND4 (N7937, N7933, N6473, N5735, N2240);
not NOT1 (N7938, N7927);
nor NOR4 (N7939, N7929, N3018, N1206, N6252);
xor XOR2 (N7940, N7939, N7793);
buf BUF1 (N7941, N7932);
buf BUF1 (N7942, N7936);
not NOT1 (N7943, N7940);
buf BUF1 (N7944, N7930);
nand NAND4 (N7945, N7943, N5233, N771, N7542);
and AND3 (N7946, N7944, N2985, N3045);
or OR2 (N7947, N7921, N7133);
xor XOR2 (N7948, N7934, N904);
nor NOR2 (N7949, N7941, N5155);
xor XOR2 (N7950, N7942, N2049);
not NOT1 (N7951, N7919);
xor XOR2 (N7952, N7951, N6793);
buf BUF1 (N7953, N7945);
nand NAND4 (N7954, N7914, N346, N7346, N1694);
not NOT1 (N7955, N7949);
xor XOR2 (N7956, N7938, N3701);
nand NAND4 (N7957, N7947, N7240, N6330, N5758);
not NOT1 (N7958, N7937);
or OR3 (N7959, N7955, N1381, N7542);
xor XOR2 (N7960, N7954, N3565);
nor NOR3 (N7961, N7952, N483, N3416);
nand NAND2 (N7962, N7959, N662);
buf BUF1 (N7963, N7946);
or OR4 (N7964, N7950, N5906, N5293, N6085);
buf BUF1 (N7965, N7953);
or OR3 (N7966, N7965, N7840, N341);
buf BUF1 (N7967, N7957);
not NOT1 (N7968, N7964);
nand NAND4 (N7969, N7958, N1476, N3451, N3544);
not NOT1 (N7970, N7960);
nand NAND2 (N7971, N7970, N5434);
nor NOR4 (N7972, N7971, N2916, N3624, N6859);
buf BUF1 (N7973, N7961);
nand NAND2 (N7974, N7963, N6676);
or OR3 (N7975, N7967, N7568, N3654);
or OR4 (N7976, N7968, N4441, N673, N2722);
and AND3 (N7977, N7973, N3167, N7495);
nand NAND2 (N7978, N7962, N1596);
nor NOR2 (N7979, N7974, N1458);
and AND4 (N7980, N7976, N4759, N126, N5184);
xor XOR2 (N7981, N7966, N2930);
or OR4 (N7982, N7979, N6277, N4798, N6457);
xor XOR2 (N7983, N7980, N4191);
and AND3 (N7984, N7956, N822, N4184);
nand NAND4 (N7985, N7975, N1324, N7283, N719);
not NOT1 (N7986, N7985);
xor XOR2 (N7987, N7972, N1487);
or OR2 (N7988, N7984, N5872);
buf BUF1 (N7989, N7969);
not NOT1 (N7990, N7989);
xor XOR2 (N7991, N7986, N1623);
nand NAND3 (N7992, N7987, N637, N2804);
not NOT1 (N7993, N7992);
and AND4 (N7994, N7990, N7111, N3784, N1787);
or OR2 (N7995, N7983, N6037);
nand NAND3 (N7996, N7948, N7033, N635);
and AND4 (N7997, N7993, N7618, N535, N5896);
nand NAND2 (N7998, N7981, N2995);
nand NAND4 (N7999, N7995, N5641, N5261, N2249);
xor XOR2 (N8000, N7977, N6317);
and AND2 (N8001, N7998, N1685);
and AND3 (N8002, N8000, N5219, N5635);
xor XOR2 (N8003, N7997, N1910);
buf BUF1 (N8004, N7982);
not NOT1 (N8005, N8001);
and AND2 (N8006, N7999, N2592);
nand NAND4 (N8007, N8004, N3541, N6330, N2478);
xor XOR2 (N8008, N7996, N4784);
and AND3 (N8009, N8008, N509, N6345);
or OR2 (N8010, N8002, N3782);
nand NAND2 (N8011, N7991, N630);
not NOT1 (N8012, N7994);
and AND3 (N8013, N7978, N3004, N6389);
and AND3 (N8014, N8007, N4417, N5092);
nand NAND4 (N8015, N8011, N741, N3854, N2019);
or OR2 (N8016, N7988, N6806);
nand NAND2 (N8017, N8014, N2581);
nor NOR4 (N8018, N8013, N4086, N5056, N4463);
not NOT1 (N8019, N8016);
xor XOR2 (N8020, N8018, N4937);
buf BUF1 (N8021, N8009);
xor XOR2 (N8022, N8021, N678);
buf BUF1 (N8023, N8020);
and AND3 (N8024, N8006, N6746, N6288);
buf BUF1 (N8025, N8003);
and AND2 (N8026, N8024, N500);
nor NOR4 (N8027, N8026, N4098, N899, N1936);
and AND3 (N8028, N8010, N4898, N6856);
or OR4 (N8029, N8015, N6589, N26, N932);
not NOT1 (N8030, N8028);
nand NAND3 (N8031, N8023, N2442, N5255);
xor XOR2 (N8032, N8017, N7372);
nor NOR3 (N8033, N8030, N3544, N7284);
buf BUF1 (N8034, N8029);
xor XOR2 (N8035, N8027, N2324);
buf BUF1 (N8036, N8025);
or OR3 (N8037, N8033, N5115, N5972);
buf BUF1 (N8038, N8034);
nor NOR4 (N8039, N8037, N818, N184, N2069);
and AND4 (N8040, N8022, N7065, N1630, N4557);
nor NOR2 (N8041, N8038, N379);
xor XOR2 (N8042, N8035, N2120);
not NOT1 (N8043, N8019);
not NOT1 (N8044, N8031);
or OR2 (N8045, N8041, N3154);
not NOT1 (N8046, N8032);
buf BUF1 (N8047, N8036);
or OR4 (N8048, N8039, N6213, N6992, N2809);
and AND3 (N8049, N8045, N7367, N5801);
not NOT1 (N8050, N8044);
or OR2 (N8051, N8046, N7555);
or OR2 (N8052, N8047, N3865);
nor NOR4 (N8053, N8005, N2514, N6720, N7648);
or OR3 (N8054, N8049, N4853, N6701);
and AND4 (N8055, N8040, N5277, N1129, N1786);
buf BUF1 (N8056, N8042);
or OR4 (N8057, N8012, N557, N1637, N2521);
and AND4 (N8058, N8048, N5548, N2335, N1346);
not NOT1 (N8059, N8051);
or OR2 (N8060, N8043, N1162);
and AND4 (N8061, N8058, N2050, N3386, N5256);
or OR3 (N8062, N8052, N6497, N1766);
xor XOR2 (N8063, N8061, N1130);
nor NOR4 (N8064, N8060, N2701, N2855, N6356);
xor XOR2 (N8065, N8055, N7802);
buf BUF1 (N8066, N8054);
nor NOR3 (N8067, N8062, N1157, N3378);
or OR2 (N8068, N8056, N3542);
xor XOR2 (N8069, N8059, N5435);
or OR4 (N8070, N8053, N139, N1306, N5050);
not NOT1 (N8071, N8070);
and AND3 (N8072, N8067, N8029, N442);
and AND2 (N8073, N8065, N2784);
nor NOR3 (N8074, N8073, N3162, N6102);
nor NOR4 (N8075, N8057, N5650, N4793, N2193);
xor XOR2 (N8076, N8063, N306);
xor XOR2 (N8077, N8071, N6104);
nor NOR4 (N8078, N8077, N5343, N3859, N4193);
not NOT1 (N8079, N8064);
nor NOR4 (N8080, N8078, N6420, N6819, N5015);
buf BUF1 (N8081, N8079);
or OR3 (N8082, N8066, N7240, N3932);
and AND4 (N8083, N8069, N2348, N4485, N6391);
buf BUF1 (N8084, N8074);
xor XOR2 (N8085, N8080, N1023);
not NOT1 (N8086, N8085);
not NOT1 (N8087, N8081);
not NOT1 (N8088, N8075);
xor XOR2 (N8089, N8087, N50);
nor NOR3 (N8090, N8084, N7245, N6015);
or OR4 (N8091, N8072, N2411, N7935, N3809);
not NOT1 (N8092, N8076);
nor NOR3 (N8093, N8091, N2066, N4171);
and AND2 (N8094, N8068, N4337);
nor NOR2 (N8095, N8086, N4643);
nor NOR4 (N8096, N8093, N1478, N6835, N6607);
not NOT1 (N8097, N8088);
or OR3 (N8098, N8092, N2006, N4492);
nor NOR4 (N8099, N8089, N3342, N5818, N1358);
xor XOR2 (N8100, N8097, N5126);
not NOT1 (N8101, N8082);
xor XOR2 (N8102, N8096, N3197);
buf BUF1 (N8103, N8095);
not NOT1 (N8104, N8103);
nor NOR2 (N8105, N8094, N1624);
or OR4 (N8106, N8104, N5811, N6863, N7286);
buf BUF1 (N8107, N8102);
or OR2 (N8108, N8101, N1472);
or OR4 (N8109, N8099, N2834, N7113, N1121);
buf BUF1 (N8110, N8105);
nand NAND2 (N8111, N8110, N1699);
nand NAND3 (N8112, N8111, N5173, N4864);
nor NOR2 (N8113, N8050, N1803);
xor XOR2 (N8114, N8098, N4056);
and AND3 (N8115, N8108, N552, N5531);
not NOT1 (N8116, N8113);
xor XOR2 (N8117, N8112, N7851);
or OR3 (N8118, N8090, N1028, N6345);
xor XOR2 (N8119, N8106, N5469);
nor NOR4 (N8120, N8119, N779, N3912, N3185);
xor XOR2 (N8121, N8115, N5738);
or OR2 (N8122, N8117, N5214);
buf BUF1 (N8123, N8118);
not NOT1 (N8124, N8122);
nor NOR3 (N8125, N8083, N6543, N2683);
and AND2 (N8126, N8123, N7102);
xor XOR2 (N8127, N8125, N3371);
nand NAND4 (N8128, N8121, N5418, N7515, N6527);
nand NAND3 (N8129, N8107, N4805, N2269);
xor XOR2 (N8130, N8120, N6122);
xor XOR2 (N8131, N8130, N5262);
not NOT1 (N8132, N8131);
or OR4 (N8133, N8132, N7221, N663, N5354);
or OR3 (N8134, N8100, N5833, N7658);
xor XOR2 (N8135, N8129, N7354);
or OR3 (N8136, N8135, N4131, N2585);
nand NAND4 (N8137, N8114, N1218, N879, N5354);
xor XOR2 (N8138, N8116, N5660);
buf BUF1 (N8139, N8134);
buf BUF1 (N8140, N8124);
nand NAND4 (N8141, N8137, N6575, N389, N2571);
nand NAND2 (N8142, N8140, N919);
or OR2 (N8143, N8138, N3914);
not NOT1 (N8144, N8139);
not NOT1 (N8145, N8109);
or OR2 (N8146, N8126, N6998);
and AND4 (N8147, N8145, N1271, N2896, N7565);
and AND2 (N8148, N8128, N7992);
nand NAND4 (N8149, N8127, N246, N3167, N2350);
and AND3 (N8150, N8136, N5854, N4493);
and AND3 (N8151, N8147, N1425, N7228);
not NOT1 (N8152, N8144);
buf BUF1 (N8153, N8141);
xor XOR2 (N8154, N8153, N3659);
and AND2 (N8155, N8151, N7533);
and AND2 (N8156, N8152, N108);
nand NAND2 (N8157, N8148, N4832);
or OR3 (N8158, N8142, N611, N5463);
and AND3 (N8159, N8133, N7536, N3246);
and AND3 (N8160, N8146, N189, N5051);
nand NAND2 (N8161, N8149, N2202);
buf BUF1 (N8162, N8158);
or OR3 (N8163, N8160, N6158, N4570);
xor XOR2 (N8164, N8162, N4986);
buf BUF1 (N8165, N8164);
and AND3 (N8166, N8155, N7484, N2268);
not NOT1 (N8167, N8143);
and AND2 (N8168, N8167, N2326);
nor NOR4 (N8169, N8157, N2133, N7115, N2009);
nand NAND4 (N8170, N8156, N2306, N7112, N7839);
buf BUF1 (N8171, N8150);
buf BUF1 (N8172, N8154);
buf BUF1 (N8173, N8169);
xor XOR2 (N8174, N8161, N7363);
nand NAND4 (N8175, N8171, N2698, N3538, N4155);
not NOT1 (N8176, N8165);
or OR3 (N8177, N8173, N6633, N1062);
not NOT1 (N8178, N8168);
or OR3 (N8179, N8178, N4423, N6419);
not NOT1 (N8180, N8163);
not NOT1 (N8181, N8179);
and AND3 (N8182, N8177, N1203, N2587);
nand NAND4 (N8183, N8166, N2667, N5324, N5909);
xor XOR2 (N8184, N8170, N5178);
nand NAND3 (N8185, N8181, N6853, N6315);
and AND4 (N8186, N8180, N7088, N5048, N532);
nand NAND2 (N8187, N8184, N6976);
nor NOR2 (N8188, N8186, N2571);
or OR4 (N8189, N8172, N2448, N792, N6933);
not NOT1 (N8190, N8174);
not NOT1 (N8191, N8175);
not NOT1 (N8192, N8190);
nor NOR2 (N8193, N8176, N4188);
nor NOR3 (N8194, N8185, N194, N3178);
nor NOR4 (N8195, N8182, N5732, N5336, N7017);
xor XOR2 (N8196, N8192, N7281);
nor NOR2 (N8197, N8159, N4470);
nand NAND4 (N8198, N8191, N452, N4016, N1298);
xor XOR2 (N8199, N8188, N7391);
not NOT1 (N8200, N8198);
nand NAND4 (N8201, N8189, N1312, N7541, N3756);
nand NAND3 (N8202, N8196, N2920, N6616);
xor XOR2 (N8203, N8197, N7726);
and AND3 (N8204, N8195, N4963, N6436);
xor XOR2 (N8205, N8202, N4298);
not NOT1 (N8206, N8187);
nor NOR2 (N8207, N8193, N6553);
nor NOR2 (N8208, N8207, N7122);
not NOT1 (N8209, N8201);
not NOT1 (N8210, N8203);
xor XOR2 (N8211, N8200, N5391);
buf BUF1 (N8212, N8183);
nor NOR2 (N8213, N8212, N6499);
nor NOR3 (N8214, N8206, N4258, N5954);
nor NOR2 (N8215, N8214, N3678);
nor NOR2 (N8216, N8209, N6055);
and AND3 (N8217, N8204, N6887, N3736);
xor XOR2 (N8218, N8215, N7275);
not NOT1 (N8219, N8218);
and AND2 (N8220, N8194, N4719);
not NOT1 (N8221, N8220);
not NOT1 (N8222, N8217);
not NOT1 (N8223, N8216);
nand NAND2 (N8224, N8219, N6423);
buf BUF1 (N8225, N8211);
buf BUF1 (N8226, N8225);
not NOT1 (N8227, N8221);
nand NAND2 (N8228, N8213, N5654);
nor NOR2 (N8229, N8222, N2556);
nor NOR4 (N8230, N8224, N471, N6747, N1328);
buf BUF1 (N8231, N8229);
buf BUF1 (N8232, N8210);
nor NOR3 (N8233, N8205, N5531, N5840);
and AND4 (N8234, N8223, N3966, N7920, N1555);
buf BUF1 (N8235, N8228);
not NOT1 (N8236, N8235);
not NOT1 (N8237, N8234);
xor XOR2 (N8238, N8230, N3294);
and AND3 (N8239, N8199, N2351, N5357);
buf BUF1 (N8240, N8239);
nor NOR4 (N8241, N8236, N3699, N3637, N293);
buf BUF1 (N8242, N8226);
xor XOR2 (N8243, N8227, N6643);
or OR2 (N8244, N8231, N5137);
and AND3 (N8245, N8233, N5090, N7460);
buf BUF1 (N8246, N8237);
and AND3 (N8247, N8241, N6722, N248);
and AND2 (N8248, N8208, N7154);
buf BUF1 (N8249, N8247);
not NOT1 (N8250, N8245);
xor XOR2 (N8251, N8248, N4164);
buf BUF1 (N8252, N8232);
nor NOR3 (N8253, N8249, N5059, N2061);
xor XOR2 (N8254, N8252, N2724);
xor XOR2 (N8255, N8250, N2018);
or OR3 (N8256, N8246, N5267, N4836);
xor XOR2 (N8257, N8253, N5651);
and AND4 (N8258, N8242, N3694, N7550, N1828);
xor XOR2 (N8259, N8256, N5076);
nor NOR2 (N8260, N8255, N1908);
not NOT1 (N8261, N8257);
buf BUF1 (N8262, N8244);
nand NAND3 (N8263, N8261, N2305, N5726);
buf BUF1 (N8264, N8263);
and AND2 (N8265, N8240, N793);
not NOT1 (N8266, N8264);
buf BUF1 (N8267, N8243);
nand NAND2 (N8268, N8267, N2450);
xor XOR2 (N8269, N8259, N3698);
not NOT1 (N8270, N8260);
buf BUF1 (N8271, N8251);
or OR3 (N8272, N8270, N3073, N7076);
buf BUF1 (N8273, N8258);
nand NAND2 (N8274, N8265, N7591);
xor XOR2 (N8275, N8266, N4351);
xor XOR2 (N8276, N8275, N2440);
nor NOR4 (N8277, N8262, N2863, N3294, N5209);
xor XOR2 (N8278, N8269, N5245);
nand NAND4 (N8279, N8274, N3568, N3762, N4096);
and AND2 (N8280, N8278, N1548);
not NOT1 (N8281, N8277);
xor XOR2 (N8282, N8268, N3927);
or OR2 (N8283, N8254, N4295);
and AND3 (N8284, N8271, N4067, N8101);
nand NAND3 (N8285, N8281, N6886, N5761);
buf BUF1 (N8286, N8284);
nor NOR2 (N8287, N8279, N4754);
not NOT1 (N8288, N8272);
nor NOR2 (N8289, N8285, N8103);
not NOT1 (N8290, N8273);
and AND4 (N8291, N8290, N3516, N657, N1608);
and AND2 (N8292, N8287, N3832);
not NOT1 (N8293, N8282);
nor NOR3 (N8294, N8283, N4652, N5110);
buf BUF1 (N8295, N8238);
buf BUF1 (N8296, N8294);
buf BUF1 (N8297, N8280);
or OR3 (N8298, N8295, N1251, N7262);
and AND2 (N8299, N8288, N1780);
or OR2 (N8300, N8289, N6474);
buf BUF1 (N8301, N8293);
nand NAND2 (N8302, N8296, N7541);
or OR4 (N8303, N8292, N2127, N4292, N1238);
buf BUF1 (N8304, N8297);
or OR2 (N8305, N8303, N7558);
xor XOR2 (N8306, N8300, N249);
nand NAND2 (N8307, N8286, N6857);
not NOT1 (N8308, N8276);
buf BUF1 (N8309, N8304);
nand NAND2 (N8310, N8305, N1729);
not NOT1 (N8311, N8291);
nor NOR4 (N8312, N8310, N7021, N4925, N2828);
and AND2 (N8313, N8309, N5008);
or OR3 (N8314, N8308, N5482, N603);
nor NOR3 (N8315, N8306, N874, N5102);
xor XOR2 (N8316, N8312, N2115);
not NOT1 (N8317, N8313);
buf BUF1 (N8318, N8301);
or OR2 (N8319, N8299, N7527);
not NOT1 (N8320, N8316);
nor NOR2 (N8321, N8298, N1235);
xor XOR2 (N8322, N8319, N7045);
nor NOR4 (N8323, N8321, N6949, N6296, N7707);
or OR4 (N8324, N8320, N2719, N4749, N866);
or OR3 (N8325, N8314, N273, N3888);
buf BUF1 (N8326, N8302);
not NOT1 (N8327, N8307);
not NOT1 (N8328, N8324);
nand NAND2 (N8329, N8323, N684);
or OR4 (N8330, N8317, N1312, N480, N6218);
nor NOR2 (N8331, N8327, N5057);
buf BUF1 (N8332, N8330);
and AND3 (N8333, N8322, N5411, N7818);
not NOT1 (N8334, N8333);
not NOT1 (N8335, N8326);
xor XOR2 (N8336, N8315, N7187);
xor XOR2 (N8337, N8328, N7680);
xor XOR2 (N8338, N8337, N7411);
and AND2 (N8339, N8311, N33);
not NOT1 (N8340, N8318);
nor NOR4 (N8341, N8334, N2710, N3437, N7144);
not NOT1 (N8342, N8340);
buf BUF1 (N8343, N8329);
nor NOR3 (N8344, N8335, N6045, N365);
and AND4 (N8345, N8341, N1156, N2185, N5124);
nor NOR3 (N8346, N8342, N4604, N111);
nor NOR2 (N8347, N8331, N5645);
nand NAND4 (N8348, N8338, N5859, N6012, N1010);
or OR3 (N8349, N8339, N387, N192);
or OR3 (N8350, N8347, N1055, N5923);
nand NAND3 (N8351, N8349, N6387, N5900);
not NOT1 (N8352, N8350);
nand NAND2 (N8353, N8332, N5578);
buf BUF1 (N8354, N8352);
buf BUF1 (N8355, N8353);
nand NAND4 (N8356, N8343, N12, N4437, N7129);
and AND2 (N8357, N8351, N5726);
and AND4 (N8358, N8355, N2660, N3595, N1514);
buf BUF1 (N8359, N8358);
nor NOR2 (N8360, N8359, N5070);
nor NOR4 (N8361, N8356, N2827, N3485, N2610);
and AND4 (N8362, N8345, N7449, N8248, N5967);
or OR2 (N8363, N8362, N2685);
nand NAND2 (N8364, N8360, N2287);
nand NAND3 (N8365, N8364, N6572, N3143);
and AND4 (N8366, N8365, N5908, N8164, N3934);
buf BUF1 (N8367, N8354);
buf BUF1 (N8368, N8325);
not NOT1 (N8369, N8348);
nor NOR3 (N8370, N8336, N8185, N3137);
not NOT1 (N8371, N8369);
and AND3 (N8372, N8370, N4920, N4964);
buf BUF1 (N8373, N8357);
nor NOR3 (N8374, N8361, N5198, N5754);
not NOT1 (N8375, N8344);
not NOT1 (N8376, N8363);
or OR3 (N8377, N8367, N4731, N1554);
nor NOR4 (N8378, N8346, N1590, N7603, N8201);
and AND2 (N8379, N8376, N4809);
or OR2 (N8380, N8378, N1377);
not NOT1 (N8381, N8375);
nand NAND2 (N8382, N8372, N223);
or OR3 (N8383, N8381, N4558, N2726);
not NOT1 (N8384, N8383);
nor NOR4 (N8385, N8374, N2481, N2642, N3624);
or OR2 (N8386, N8379, N6577);
nor NOR3 (N8387, N8382, N7593, N1385);
and AND4 (N8388, N8385, N7289, N89, N1651);
buf BUF1 (N8389, N8384);
or OR3 (N8390, N8371, N6411, N7138);
xor XOR2 (N8391, N8386, N6072);
xor XOR2 (N8392, N8368, N7723);
nor NOR4 (N8393, N8392, N7355, N6367, N1763);
nor NOR4 (N8394, N8366, N5591, N6688, N4466);
and AND4 (N8395, N8377, N1529, N3334, N3243);
and AND2 (N8396, N8387, N8394);
xor XOR2 (N8397, N687, N5120);
buf BUF1 (N8398, N8396);
xor XOR2 (N8399, N8391, N2382);
not NOT1 (N8400, N8398);
xor XOR2 (N8401, N8397, N1455);
nand NAND4 (N8402, N8389, N2473, N4878, N1900);
buf BUF1 (N8403, N8380);
and AND4 (N8404, N8402, N3810, N7069, N1681);
not NOT1 (N8405, N8393);
buf BUF1 (N8406, N8405);
nand NAND2 (N8407, N8403, N7492);
nor NOR2 (N8408, N8390, N6171);
or OR2 (N8409, N8401, N6940);
buf BUF1 (N8410, N8406);
xor XOR2 (N8411, N8388, N3786);
or OR3 (N8412, N8395, N2561, N7139);
buf BUF1 (N8413, N8412);
nand NAND2 (N8414, N8400, N6061);
xor XOR2 (N8415, N8414, N4140);
not NOT1 (N8416, N8404);
not NOT1 (N8417, N8413);
xor XOR2 (N8418, N8409, N5147);
nand NAND4 (N8419, N8399, N6734, N7493, N4507);
or OR2 (N8420, N8373, N7255);
or OR2 (N8421, N8418, N8183);
nor NOR4 (N8422, N8407, N3071, N4807, N904);
buf BUF1 (N8423, N8415);
and AND3 (N8424, N8421, N5896, N1953);
and AND4 (N8425, N8424, N4189, N1006, N6051);
buf BUF1 (N8426, N8425);
and AND4 (N8427, N8422, N5774, N2764, N4119);
and AND3 (N8428, N8417, N1064, N6625);
xor XOR2 (N8429, N8420, N3886);
not NOT1 (N8430, N8428);
not NOT1 (N8431, N8423);
nor NOR2 (N8432, N8416, N6124);
not NOT1 (N8433, N8419);
nor NOR3 (N8434, N8426, N7493, N1016);
or OR3 (N8435, N8432, N299, N5742);
nor NOR2 (N8436, N8429, N1799);
nor NOR3 (N8437, N8430, N7880, N2235);
nand NAND3 (N8438, N8435, N2291, N6001);
and AND3 (N8439, N8437, N1528, N5268);
buf BUF1 (N8440, N8438);
or OR4 (N8441, N8434, N1352, N527, N5925);
buf BUF1 (N8442, N8431);
or OR4 (N8443, N8442, N7803, N397, N3249);
buf BUF1 (N8444, N8439);
not NOT1 (N8445, N8440);
buf BUF1 (N8446, N8436);
not NOT1 (N8447, N8444);
and AND3 (N8448, N8410, N7521, N3993);
xor XOR2 (N8449, N8433, N737);
nand NAND3 (N8450, N8446, N7986, N461);
nor NOR3 (N8451, N8408, N6076, N2117);
or OR4 (N8452, N8451, N1272, N3530, N286);
or OR2 (N8453, N8452, N3073);
and AND2 (N8454, N8448, N8361);
buf BUF1 (N8455, N8449);
or OR3 (N8456, N8453, N1871, N3525);
buf BUF1 (N8457, N8456);
and AND3 (N8458, N8443, N5379, N1433);
not NOT1 (N8459, N8447);
nand NAND2 (N8460, N8427, N46);
not NOT1 (N8461, N8457);
buf BUF1 (N8462, N8441);
xor XOR2 (N8463, N8454, N3442);
nor NOR2 (N8464, N8411, N7180);
and AND3 (N8465, N8458, N4959, N8268);
xor XOR2 (N8466, N8462, N5889);
or OR4 (N8467, N8459, N3665, N6564, N5926);
nand NAND4 (N8468, N8463, N6055, N4576, N2705);
not NOT1 (N8469, N8460);
or OR3 (N8470, N8465, N418, N7380);
xor XOR2 (N8471, N8464, N1885);
and AND3 (N8472, N8467, N5748, N7383);
not NOT1 (N8473, N8461);
and AND4 (N8474, N8473, N5847, N2243, N7008);
buf BUF1 (N8475, N8468);
or OR3 (N8476, N8474, N6224, N786);
and AND4 (N8477, N8471, N4813, N7991, N5587);
buf BUF1 (N8478, N8476);
xor XOR2 (N8479, N8475, N55);
and AND4 (N8480, N8445, N1284, N951, N167);
and AND2 (N8481, N8477, N508);
nand NAND4 (N8482, N8479, N5124, N7424, N5974);
buf BUF1 (N8483, N8472);
xor XOR2 (N8484, N8469, N4203);
or OR2 (N8485, N8470, N381);
buf BUF1 (N8486, N8482);
nand NAND3 (N8487, N8478, N7073, N1484);
not NOT1 (N8488, N8483);
nand NAND4 (N8489, N8455, N1871, N2199, N3686);
nor NOR3 (N8490, N8450, N4696, N4525);
buf BUF1 (N8491, N8490);
or OR2 (N8492, N8487, N5097);
buf BUF1 (N8493, N8491);
not NOT1 (N8494, N8492);
nand NAND3 (N8495, N8480, N4076, N682);
and AND2 (N8496, N8486, N6057);
or OR2 (N8497, N8496, N3889);
nand NAND4 (N8498, N8493, N5405, N1430, N915);
nor NOR3 (N8499, N8484, N8425, N4643);
not NOT1 (N8500, N8485);
or OR4 (N8501, N8466, N4272, N5625, N7601);
xor XOR2 (N8502, N8489, N8356);
not NOT1 (N8503, N8495);
buf BUF1 (N8504, N8498);
nand NAND2 (N8505, N8497, N1340);
or OR4 (N8506, N8505, N1759, N7820, N1490);
xor XOR2 (N8507, N8500, N2390);
and AND2 (N8508, N8503, N4934);
nand NAND3 (N8509, N8502, N3664, N3208);
not NOT1 (N8510, N8501);
or OR3 (N8511, N8508, N8481, N1962);
nor NOR2 (N8512, N4940, N741);
or OR3 (N8513, N8488, N6358, N1344);
nand NAND2 (N8514, N8510, N5723);
not NOT1 (N8515, N8504);
or OR3 (N8516, N8514, N1606, N4452);
or OR4 (N8517, N8516, N2877, N5863, N5595);
buf BUF1 (N8518, N8515);
nand NAND4 (N8519, N8507, N7387, N4657, N4408);
buf BUF1 (N8520, N8518);
and AND3 (N8521, N8499, N1452, N5936);
and AND3 (N8522, N8521, N4157, N2889);
not NOT1 (N8523, N8522);
buf BUF1 (N8524, N8494);
nand NAND2 (N8525, N8524, N248);
buf BUF1 (N8526, N8506);
xor XOR2 (N8527, N8520, N2346);
nor NOR2 (N8528, N8513, N320);
nand NAND2 (N8529, N8526, N3948);
or OR4 (N8530, N8525, N5861, N2642, N8490);
or OR3 (N8531, N8512, N1353, N336);
nand NAND2 (N8532, N8527, N3483);
or OR3 (N8533, N8509, N7592, N1979);
nor NOR3 (N8534, N8529, N367, N3676);
and AND4 (N8535, N8533, N7245, N332, N6984);
not NOT1 (N8536, N8523);
nand NAND3 (N8537, N8534, N4581, N271);
and AND2 (N8538, N8528, N4008);
and AND2 (N8539, N8530, N3343);
buf BUF1 (N8540, N8539);
not NOT1 (N8541, N8536);
or OR2 (N8542, N8511, N1874);
buf BUF1 (N8543, N8537);
xor XOR2 (N8544, N8538, N3756);
buf BUF1 (N8545, N8540);
xor XOR2 (N8546, N8544, N4103);
nor NOR3 (N8547, N8542, N6818, N7075);
and AND4 (N8548, N8543, N1768, N8527, N7338);
or OR4 (N8549, N8541, N1682, N431, N749);
buf BUF1 (N8550, N8535);
not NOT1 (N8551, N8549);
nand NAND4 (N8552, N8547, N957, N137, N6651);
and AND3 (N8553, N8546, N1966, N3456);
and AND4 (N8554, N8532, N1050, N8338, N6804);
xor XOR2 (N8555, N8554, N3139);
buf BUF1 (N8556, N8555);
nand NAND2 (N8557, N8552, N3561);
not NOT1 (N8558, N8553);
not NOT1 (N8559, N8557);
xor XOR2 (N8560, N8551, N1444);
or OR2 (N8561, N8556, N614);
nor NOR2 (N8562, N8545, N3508);
xor XOR2 (N8563, N8548, N1690);
nand NAND2 (N8564, N8531, N4738);
buf BUF1 (N8565, N8564);
nor NOR4 (N8566, N8519, N3421, N1423, N8045);
nand NAND2 (N8567, N8560, N7594);
not NOT1 (N8568, N8563);
not NOT1 (N8569, N8562);
and AND4 (N8570, N8559, N6911, N1929, N4891);
buf BUF1 (N8571, N8565);
nand NAND2 (N8572, N8567, N6389);
nor NOR2 (N8573, N8561, N8200);
buf BUF1 (N8574, N8573);
nor NOR2 (N8575, N8558, N5180);
nand NAND2 (N8576, N8571, N8306);
or OR2 (N8577, N8572, N4311);
not NOT1 (N8578, N8568);
or OR3 (N8579, N8574, N6973, N156);
or OR2 (N8580, N8550, N1927);
nand NAND4 (N8581, N8575, N1318, N754, N7429);
nand NAND3 (N8582, N8517, N1308, N1983);
xor XOR2 (N8583, N8566, N2293);
not NOT1 (N8584, N8581);
xor XOR2 (N8585, N8576, N4713);
nor NOR3 (N8586, N8583, N4151, N1263);
nor NOR3 (N8587, N8577, N4881, N4704);
xor XOR2 (N8588, N8580, N7630);
nor NOR4 (N8589, N8579, N7477, N1829, N2955);
nor NOR4 (N8590, N8588, N6153, N5055, N4980);
or OR4 (N8591, N8585, N6923, N5770, N8010);
xor XOR2 (N8592, N8587, N6526);
nor NOR3 (N8593, N8584, N8036, N4787);
xor XOR2 (N8594, N8589, N5906);
nand NAND3 (N8595, N8578, N5145, N4084);
or OR3 (N8596, N8590, N871, N6047);
not NOT1 (N8597, N8586);
nand NAND4 (N8598, N8594, N5120, N113, N132);
nand NAND2 (N8599, N8598, N6929);
nand NAND3 (N8600, N8582, N3553, N190);
and AND2 (N8601, N8592, N3186);
nor NOR4 (N8602, N8570, N8129, N4824, N7073);
nand NAND3 (N8603, N8593, N6592, N7193);
or OR2 (N8604, N8597, N8451);
nor NOR3 (N8605, N8599, N2693, N1771);
buf BUF1 (N8606, N8603);
not NOT1 (N8607, N8591);
nand NAND3 (N8608, N8605, N4197, N8190);
nand NAND4 (N8609, N8601, N2182, N7728, N5047);
and AND4 (N8610, N8607, N4886, N7326, N2902);
xor XOR2 (N8611, N8608, N5713);
and AND2 (N8612, N8611, N7790);
nand NAND2 (N8613, N8612, N1577);
not NOT1 (N8614, N8610);
nand NAND4 (N8615, N8609, N7734, N866, N2434);
nand NAND4 (N8616, N8569, N4605, N7907, N6900);
nand NAND4 (N8617, N8602, N5317, N3717, N251);
buf BUF1 (N8618, N8614);
nor NOR2 (N8619, N8596, N4771);
nand NAND4 (N8620, N8604, N3576, N6409, N6732);
buf BUF1 (N8621, N8600);
and AND4 (N8622, N8618, N2984, N188, N3701);
buf BUF1 (N8623, N8620);
not NOT1 (N8624, N8616);
and AND3 (N8625, N8622, N3276, N499);
or OR4 (N8626, N8624, N8126, N5519, N5198);
xor XOR2 (N8627, N8615, N2069);
buf BUF1 (N8628, N8625);
buf BUF1 (N8629, N8613);
not NOT1 (N8630, N8606);
or OR2 (N8631, N8629, N1572);
xor XOR2 (N8632, N8623, N4682);
buf BUF1 (N8633, N8621);
xor XOR2 (N8634, N8631, N8061);
or OR2 (N8635, N8630, N555);
buf BUF1 (N8636, N8634);
and AND2 (N8637, N8617, N3962);
or OR3 (N8638, N8633, N6886, N993);
or OR2 (N8639, N8638, N7098);
xor XOR2 (N8640, N8628, N7550);
and AND4 (N8641, N8637, N53, N7383, N5318);
nor NOR3 (N8642, N8626, N4155, N140);
nor NOR2 (N8643, N8636, N2281);
buf BUF1 (N8644, N8641);
not NOT1 (N8645, N8595);
xor XOR2 (N8646, N8644, N4995);
nor NOR3 (N8647, N8640, N6236, N6815);
nor NOR3 (N8648, N8639, N1088, N8084);
not NOT1 (N8649, N8627);
not NOT1 (N8650, N8649);
or OR4 (N8651, N8635, N462, N7905, N8609);
not NOT1 (N8652, N8648);
nor NOR2 (N8653, N8642, N5887);
xor XOR2 (N8654, N8632, N7421);
and AND3 (N8655, N8652, N4853, N4444);
nand NAND2 (N8656, N8619, N477);
nor NOR4 (N8657, N8646, N6838, N5657, N2415);
nor NOR2 (N8658, N8650, N2537);
nand NAND2 (N8659, N8654, N6629);
not NOT1 (N8660, N8647);
nor NOR3 (N8661, N8659, N2760, N6243);
buf BUF1 (N8662, N8645);
buf BUF1 (N8663, N8657);
buf BUF1 (N8664, N8663);
nor NOR2 (N8665, N8664, N6906);
not NOT1 (N8666, N8665);
nor NOR3 (N8667, N8658, N1926, N5145);
not NOT1 (N8668, N8651);
nor NOR2 (N8669, N8643, N7084);
and AND3 (N8670, N8661, N2925, N4111);
xor XOR2 (N8671, N8667, N133);
not NOT1 (N8672, N8660);
xor XOR2 (N8673, N8671, N172);
or OR3 (N8674, N8670, N2466, N8325);
xor XOR2 (N8675, N8666, N8220);
xor XOR2 (N8676, N8675, N1116);
and AND4 (N8677, N8655, N3389, N7457, N6741);
not NOT1 (N8678, N8674);
and AND2 (N8679, N8669, N4016);
nor NOR3 (N8680, N8653, N3545, N4141);
not NOT1 (N8681, N8680);
or OR2 (N8682, N8672, N3527);
nor NOR3 (N8683, N8679, N1719, N1239);
xor XOR2 (N8684, N8668, N2836);
nand NAND4 (N8685, N8678, N5420, N2725, N4264);
not NOT1 (N8686, N8683);
xor XOR2 (N8687, N8686, N2227);
buf BUF1 (N8688, N8687);
buf BUF1 (N8689, N8673);
not NOT1 (N8690, N8684);
or OR3 (N8691, N8656, N6386, N7734);
and AND4 (N8692, N8690, N6101, N2475, N6509);
nor NOR3 (N8693, N8685, N5760, N6445);
not NOT1 (N8694, N8688);
not NOT1 (N8695, N8693);
or OR4 (N8696, N8662, N7658, N3926, N5442);
and AND4 (N8697, N8696, N8497, N2363, N8559);
or OR3 (N8698, N8691, N7173, N560);
nor NOR4 (N8699, N8697, N5925, N4381, N7745);
and AND4 (N8700, N8681, N4510, N2117, N1201);
buf BUF1 (N8701, N8682);
or OR2 (N8702, N8689, N638);
nand NAND3 (N8703, N8701, N2171, N7996);
not NOT1 (N8704, N8677);
buf BUF1 (N8705, N8695);
and AND4 (N8706, N8702, N4487, N3606, N6532);
or OR2 (N8707, N8698, N26);
nand NAND2 (N8708, N8707, N7422);
and AND2 (N8709, N8700, N4417);
xor XOR2 (N8710, N8704, N3593);
not NOT1 (N8711, N8709);
nor NOR2 (N8712, N8676, N719);
xor XOR2 (N8713, N8692, N4074);
xor XOR2 (N8714, N8699, N6434);
buf BUF1 (N8715, N8710);
and AND4 (N8716, N8694, N8073, N6685, N4610);
or OR3 (N8717, N8706, N4087, N7448);
or OR4 (N8718, N8714, N1923, N1036, N6168);
xor XOR2 (N8719, N8715, N8520);
or OR3 (N8720, N8716, N7716, N254);
nand NAND2 (N8721, N8712, N3758);
nand NAND4 (N8722, N8713, N8341, N5181, N8239);
or OR3 (N8723, N8717, N5592, N1829);
nor NOR2 (N8724, N8705, N1866);
nand NAND3 (N8725, N8723, N296, N2655);
xor XOR2 (N8726, N8722, N2970);
and AND4 (N8727, N8724, N5198, N6636, N6510);
buf BUF1 (N8728, N8727);
or OR2 (N8729, N8726, N1581);
nor NOR2 (N8730, N8708, N5701);
buf BUF1 (N8731, N8720);
nand NAND4 (N8732, N8721, N1837, N555, N76);
not NOT1 (N8733, N8728);
nor NOR2 (N8734, N8732, N4010);
and AND3 (N8735, N8703, N11, N4015);
and AND2 (N8736, N8725, N2685);
or OR3 (N8737, N8719, N7795, N8566);
buf BUF1 (N8738, N8731);
xor XOR2 (N8739, N8737, N2909);
nand NAND4 (N8740, N8733, N4053, N3931, N7142);
or OR3 (N8741, N8711, N4875, N4601);
nor NOR2 (N8742, N8730, N4009);
and AND3 (N8743, N8735, N5514, N8598);
nor NOR2 (N8744, N8738, N6632);
xor XOR2 (N8745, N8729, N7648);
buf BUF1 (N8746, N8741);
and AND4 (N8747, N8718, N3307, N6050, N3631);
nand NAND2 (N8748, N8739, N4219);
nand NAND4 (N8749, N8736, N5143, N2389, N2326);
nor NOR4 (N8750, N8749, N121, N5352, N4710);
nor NOR3 (N8751, N8740, N4237, N5275);
nand NAND3 (N8752, N8746, N5885, N5723);
buf BUF1 (N8753, N8744);
not NOT1 (N8754, N8743);
xor XOR2 (N8755, N8747, N8215);
xor XOR2 (N8756, N8748, N3851);
and AND4 (N8757, N8753, N3498, N4455, N3540);
or OR4 (N8758, N8752, N7430, N4533, N8270);
nor NOR4 (N8759, N8750, N7518, N7405, N4298);
or OR3 (N8760, N8734, N2459, N6049);
xor XOR2 (N8761, N8742, N1987);
or OR4 (N8762, N8761, N1483, N8412, N3536);
xor XOR2 (N8763, N8751, N6477);
or OR4 (N8764, N8754, N6052, N2558, N4169);
and AND2 (N8765, N8760, N8501);
nor NOR2 (N8766, N8763, N840);
and AND3 (N8767, N8766, N3401, N6669);
nor NOR4 (N8768, N8755, N4144, N8724, N8675);
and AND4 (N8769, N8745, N7127, N3128, N8618);
or OR3 (N8770, N8757, N264, N5207);
nor NOR2 (N8771, N8765, N2371);
xor XOR2 (N8772, N8770, N5387);
nor NOR2 (N8773, N8767, N5869);
nand NAND2 (N8774, N8773, N4541);
and AND2 (N8775, N8758, N57);
nor NOR2 (N8776, N8759, N2647);
and AND4 (N8777, N8769, N5352, N6300, N3273);
and AND4 (N8778, N8772, N5115, N5378, N3834);
or OR2 (N8779, N8775, N6007);
not NOT1 (N8780, N8764);
or OR4 (N8781, N8777, N3984, N3015, N1547);
buf BUF1 (N8782, N8781);
nor NOR3 (N8783, N8782, N320, N3409);
nand NAND3 (N8784, N8776, N5225, N6389);
not NOT1 (N8785, N8771);
nand NAND2 (N8786, N8779, N8623);
nor NOR3 (N8787, N8786, N1769, N2891);
or OR2 (N8788, N8783, N7519);
buf BUF1 (N8789, N8778);
and AND2 (N8790, N8762, N7895);
or OR4 (N8791, N8788, N8503, N5575, N1073);
not NOT1 (N8792, N8768);
buf BUF1 (N8793, N8790);
not NOT1 (N8794, N8793);
nor NOR4 (N8795, N8789, N7753, N5004, N7684);
buf BUF1 (N8796, N8784);
or OR4 (N8797, N8794, N2037, N4444, N590);
buf BUF1 (N8798, N8792);
nand NAND4 (N8799, N8756, N5565, N4814, N7004);
and AND4 (N8800, N8787, N6771, N8745, N6483);
or OR4 (N8801, N8797, N2552, N7432, N1804);
nand NAND3 (N8802, N8801, N2701, N2300);
nand NAND3 (N8803, N8798, N7920, N2212);
and AND2 (N8804, N8791, N3931);
xor XOR2 (N8805, N8796, N7380);
xor XOR2 (N8806, N8774, N6500);
and AND3 (N8807, N8805, N4941, N4761);
nor NOR3 (N8808, N8780, N1737, N567);
nand NAND2 (N8809, N8799, N678);
or OR2 (N8810, N8806, N4764);
and AND3 (N8811, N8803, N6216, N3780);
xor XOR2 (N8812, N8785, N2189);
nor NOR2 (N8813, N8800, N8788);
nor NOR2 (N8814, N8808, N1379);
buf BUF1 (N8815, N8813);
buf BUF1 (N8816, N8804);
nor NOR2 (N8817, N8812, N3866);
buf BUF1 (N8818, N8817);
nor NOR2 (N8819, N8814, N1555);
xor XOR2 (N8820, N8815, N6725);
xor XOR2 (N8821, N8820, N3882);
and AND3 (N8822, N8810, N2617, N3924);
nor NOR3 (N8823, N8818, N784, N5319);
xor XOR2 (N8824, N8821, N2200);
xor XOR2 (N8825, N8795, N5670);
nor NOR4 (N8826, N8819, N7574, N4446, N8431);
nand NAND2 (N8827, N8822, N3816);
buf BUF1 (N8828, N8802);
and AND2 (N8829, N8825, N8420);
nor NOR4 (N8830, N8826, N3162, N283, N3807);
not NOT1 (N8831, N8828);
buf BUF1 (N8832, N8829);
xor XOR2 (N8833, N8831, N2163);
and AND3 (N8834, N8824, N909, N3115);
or OR2 (N8835, N8834, N4409);
nor NOR4 (N8836, N8835, N2608, N2149, N6619);
buf BUF1 (N8837, N8827);
xor XOR2 (N8838, N8809, N661);
or OR3 (N8839, N8823, N841, N7164);
not NOT1 (N8840, N8839);
buf BUF1 (N8841, N8836);
nor NOR3 (N8842, N8841, N7683, N7202);
not NOT1 (N8843, N8807);
and AND4 (N8844, N8816, N6251, N2559, N1158);
not NOT1 (N8845, N8844);
buf BUF1 (N8846, N8838);
nand NAND4 (N8847, N8846, N5874, N1461, N5466);
xor XOR2 (N8848, N8847, N6145);
not NOT1 (N8849, N8845);
buf BUF1 (N8850, N8840);
or OR2 (N8851, N8842, N5551);
or OR3 (N8852, N8811, N3663, N4061);
and AND2 (N8853, N8852, N4632);
not NOT1 (N8854, N8830);
buf BUF1 (N8855, N8849);
and AND3 (N8856, N8854, N7951, N3114);
xor XOR2 (N8857, N8855, N385);
not NOT1 (N8858, N8837);
nand NAND2 (N8859, N8853, N4184);
and AND2 (N8860, N8859, N3296);
nor NOR3 (N8861, N8832, N3485, N8780);
buf BUF1 (N8862, N8833);
or OR3 (N8863, N8848, N3741, N5442);
and AND3 (N8864, N8856, N1349, N2084);
nor NOR4 (N8865, N8850, N2656, N202, N5777);
not NOT1 (N8866, N8861);
nor NOR3 (N8867, N8857, N6012, N7812);
nor NOR2 (N8868, N8865, N3490);
and AND3 (N8869, N8866, N7663, N4623);
xor XOR2 (N8870, N8867, N5947);
xor XOR2 (N8871, N8864, N7874);
or OR4 (N8872, N8858, N7306, N4812, N4877);
buf BUF1 (N8873, N8868);
not NOT1 (N8874, N8871);
and AND4 (N8875, N8870, N4956, N2608, N851);
not NOT1 (N8876, N8843);
nor NOR2 (N8877, N8873, N6891);
buf BUF1 (N8878, N8862);
or OR3 (N8879, N8875, N3962, N7310);
xor XOR2 (N8880, N8874, N2021);
buf BUF1 (N8881, N8860);
not NOT1 (N8882, N8863);
nand NAND3 (N8883, N8876, N6178, N4613);
nor NOR4 (N8884, N8879, N5926, N4727, N379);
or OR3 (N8885, N8881, N1652, N6763);
buf BUF1 (N8886, N8872);
nor NOR4 (N8887, N8883, N2575, N125, N5856);
nand NAND2 (N8888, N8884, N3832);
not NOT1 (N8889, N8880);
and AND2 (N8890, N8885, N4004);
buf BUF1 (N8891, N8887);
and AND4 (N8892, N8889, N6831, N1015, N1524);
and AND4 (N8893, N8888, N3463, N1607, N7929);
or OR2 (N8894, N8886, N6503);
buf BUF1 (N8895, N8877);
nor NOR2 (N8896, N8894, N4523);
and AND4 (N8897, N8891, N2399, N1051, N6106);
and AND2 (N8898, N8890, N2349);
not NOT1 (N8899, N8896);
nor NOR2 (N8900, N8899, N4488);
nand NAND4 (N8901, N8878, N5295, N2228, N3040);
or OR4 (N8902, N8900, N4826, N8384, N769);
buf BUF1 (N8903, N8901);
or OR4 (N8904, N8898, N5851, N2107, N4148);
not NOT1 (N8905, N8892);
not NOT1 (N8906, N8893);
or OR3 (N8907, N8902, N3512, N2981);
nor NOR2 (N8908, N8906, N533);
nand NAND4 (N8909, N8903, N7709, N527, N4738);
or OR3 (N8910, N8904, N4832, N4277);
nand NAND3 (N8911, N8908, N5655, N3054);
nand NAND3 (N8912, N8905, N2423, N6773);
or OR3 (N8913, N8912, N4268, N2725);
or OR3 (N8914, N8897, N1811, N349);
nand NAND4 (N8915, N8895, N3185, N6053, N8451);
xor XOR2 (N8916, N8851, N1738);
not NOT1 (N8917, N8915);
nand NAND2 (N8918, N8911, N3185);
or OR3 (N8919, N8914, N8474, N1277);
nor NOR3 (N8920, N8907, N8644, N8077);
not NOT1 (N8921, N8920);
nor NOR3 (N8922, N8913, N4645, N5895);
and AND3 (N8923, N8916, N6306, N7537);
and AND4 (N8924, N8882, N6716, N3654, N7770);
or OR3 (N8925, N8918, N8852, N7917);
buf BUF1 (N8926, N8924);
not NOT1 (N8927, N8921);
and AND2 (N8928, N8922, N8212);
xor XOR2 (N8929, N8928, N5971);
nor NOR2 (N8930, N8909, N6929);
buf BUF1 (N8931, N8925);
or OR3 (N8932, N8929, N4390, N2672);
xor XOR2 (N8933, N8923, N7412);
nor NOR3 (N8934, N8931, N84, N7543);
nor NOR3 (N8935, N8910, N7614, N4733);
or OR4 (N8936, N8927, N970, N4831, N3343);
nor NOR3 (N8937, N8869, N6374, N7265);
not NOT1 (N8938, N8917);
nand NAND2 (N8939, N8938, N7152);
xor XOR2 (N8940, N8936, N6368);
or OR3 (N8941, N8919, N2685, N2339);
nor NOR3 (N8942, N8939, N6258, N8875);
nor NOR4 (N8943, N8933, N4998, N2101, N1774);
and AND2 (N8944, N8937, N1603);
nor NOR2 (N8945, N8944, N1986);
and AND2 (N8946, N8945, N3827);
not NOT1 (N8947, N8946);
and AND2 (N8948, N8940, N3326);
xor XOR2 (N8949, N8942, N595);
and AND4 (N8950, N8948, N3547, N368, N6894);
not NOT1 (N8951, N8941);
not NOT1 (N8952, N8930);
or OR2 (N8953, N8950, N8915);
nor NOR4 (N8954, N8943, N3215, N2352, N5075);
buf BUF1 (N8955, N8951);
buf BUF1 (N8956, N8949);
nand NAND2 (N8957, N8932, N5445);
xor XOR2 (N8958, N8956, N6092);
or OR4 (N8959, N8926, N5432, N8904, N1336);
xor XOR2 (N8960, N8947, N8674);
nand NAND2 (N8961, N8952, N536);
nor NOR4 (N8962, N8957, N1232, N3564, N1543);
or OR2 (N8963, N8934, N5933);
nand NAND4 (N8964, N8955, N4968, N1878, N8825);
buf BUF1 (N8965, N8961);
buf BUF1 (N8966, N8963);
nor NOR2 (N8967, N8959, N748);
and AND4 (N8968, N8965, N3673, N2465, N8094);
xor XOR2 (N8969, N8964, N1522);
xor XOR2 (N8970, N8958, N1073);
buf BUF1 (N8971, N8969);
buf BUF1 (N8972, N8967);
nand NAND4 (N8973, N8953, N6992, N6534, N3766);
and AND3 (N8974, N8972, N7155, N3665);
buf BUF1 (N8975, N8954);
not NOT1 (N8976, N8968);
or OR3 (N8977, N8974, N1875, N2938);
nand NAND4 (N8978, N8962, N3701, N3841, N4817);
xor XOR2 (N8979, N8975, N8082);
nand NAND4 (N8980, N8979, N4990, N5276, N5036);
buf BUF1 (N8981, N8980);
and AND4 (N8982, N8960, N2099, N1437, N1054);
nand NAND2 (N8983, N8978, N6258);
and AND2 (N8984, N8981, N6486);
or OR4 (N8985, N8970, N6607, N2145, N6429);
nand NAND4 (N8986, N8976, N3783, N4658, N6893);
not NOT1 (N8987, N8966);
buf BUF1 (N8988, N8985);
nand NAND4 (N8989, N8982, N4084, N1390, N3458);
not NOT1 (N8990, N8973);
or OR2 (N8991, N8983, N6253);
not NOT1 (N8992, N8989);
or OR4 (N8993, N8992, N6153, N8616, N8143);
buf BUF1 (N8994, N8990);
not NOT1 (N8995, N8988);
xor XOR2 (N8996, N8991, N4714);
buf BUF1 (N8997, N8986);
xor XOR2 (N8998, N8971, N3996);
and AND4 (N8999, N8935, N1904, N1176, N3329);
or OR2 (N9000, N8995, N2065);
xor XOR2 (N9001, N8999, N1159);
and AND2 (N9002, N9000, N3690);
nand NAND3 (N9003, N8993, N1922, N2974);
xor XOR2 (N9004, N9003, N4850);
not NOT1 (N9005, N8994);
nor NOR3 (N9006, N8984, N5159, N3688);
nand NAND3 (N9007, N8977, N559, N349);
buf BUF1 (N9008, N8996);
nor NOR2 (N9009, N9008, N7776);
buf BUF1 (N9010, N9002);
xor XOR2 (N9011, N9006, N1347);
xor XOR2 (N9012, N9004, N6375);
buf BUF1 (N9013, N9001);
not NOT1 (N9014, N9005);
or OR4 (N9015, N9012, N3899, N7731, N4534);
nand NAND2 (N9016, N8998, N4413);
and AND4 (N9017, N9013, N2926, N8300, N1466);
or OR4 (N9018, N8997, N1253, N2905, N815);
buf BUF1 (N9019, N9016);
nor NOR4 (N9020, N9014, N8356, N3853, N7222);
not NOT1 (N9021, N9018);
not NOT1 (N9022, N9020);
nand NAND3 (N9023, N8987, N2251, N3462);
or OR3 (N9024, N9009, N6318, N4471);
not NOT1 (N9025, N9019);
buf BUF1 (N9026, N9022);
not NOT1 (N9027, N9024);
nand NAND3 (N9028, N9026, N6546, N965);
xor XOR2 (N9029, N9017, N4273);
and AND2 (N9030, N9023, N6236);
nand NAND3 (N9031, N9007, N2777, N2349);
or OR4 (N9032, N9011, N3742, N5912, N5059);
or OR2 (N9033, N9028, N7304);
nand NAND4 (N9034, N9015, N2716, N7154, N4039);
buf BUF1 (N9035, N9033);
nor NOR4 (N9036, N9035, N6949, N4088, N1905);
and AND2 (N9037, N9031, N7172);
nor NOR3 (N9038, N9030, N7710, N5780);
nand NAND4 (N9039, N9032, N3229, N4490, N6670);
and AND2 (N9040, N9039, N7693);
nor NOR4 (N9041, N9036, N4274, N5361, N4451);
or OR3 (N9042, N9027, N1631, N3357);
not NOT1 (N9043, N9040);
or OR4 (N9044, N9042, N6470, N832, N4415);
xor XOR2 (N9045, N9041, N8772);
not NOT1 (N9046, N9021);
not NOT1 (N9047, N9010);
buf BUF1 (N9048, N9045);
and AND2 (N9049, N9044, N3484);
not NOT1 (N9050, N9038);
and AND3 (N9051, N9048, N2416, N5317);
not NOT1 (N9052, N9037);
nand NAND2 (N9053, N9046, N1894);
nand NAND2 (N9054, N9049, N1202);
buf BUF1 (N9055, N9029);
nor NOR3 (N9056, N9055, N5070, N1086);
not NOT1 (N9057, N9043);
nand NAND3 (N9058, N9057, N2753, N3596);
buf BUF1 (N9059, N9025);
or OR2 (N9060, N9056, N4088);
nand NAND3 (N9061, N9050, N7468, N7106);
not NOT1 (N9062, N9058);
or OR2 (N9063, N9052, N1110);
and AND3 (N9064, N9053, N8558, N8599);
and AND3 (N9065, N9063, N8764, N559);
or OR3 (N9066, N9034, N2978, N3049);
not NOT1 (N9067, N9060);
and AND4 (N9068, N9061, N4847, N4152, N2508);
xor XOR2 (N9069, N9067, N3899);
buf BUF1 (N9070, N9068);
not NOT1 (N9071, N9069);
xor XOR2 (N9072, N9064, N268);
not NOT1 (N9073, N9051);
xor XOR2 (N9074, N9073, N6623);
or OR2 (N9075, N9047, N755);
or OR3 (N9076, N9066, N476, N1376);
and AND3 (N9077, N9071, N2121, N974);
nand NAND4 (N9078, N9077, N4087, N398, N3655);
nor NOR2 (N9079, N9075, N212);
and AND2 (N9080, N9076, N1909);
and AND4 (N9081, N9080, N4968, N635, N5530);
and AND2 (N9082, N9079, N4041);
or OR3 (N9083, N9062, N8936, N5610);
not NOT1 (N9084, N9078);
buf BUF1 (N9085, N9083);
and AND4 (N9086, N9072, N6143, N231, N2808);
not NOT1 (N9087, N9081);
or OR3 (N9088, N9065, N2245, N8793);
not NOT1 (N9089, N9088);
nor NOR3 (N9090, N9084, N6482, N40);
and AND2 (N9091, N9090, N959);
nor NOR4 (N9092, N9082, N3232, N9023, N1072);
not NOT1 (N9093, N9085);
buf BUF1 (N9094, N9091);
xor XOR2 (N9095, N9089, N7873);
and AND3 (N9096, N9095, N5272, N3892);
or OR2 (N9097, N9092, N5264);
and AND3 (N9098, N9087, N5253, N796);
or OR4 (N9099, N9093, N5973, N7440, N6348);
not NOT1 (N9100, N9059);
nor NOR3 (N9101, N9054, N6458, N8045);
or OR4 (N9102, N9070, N1083, N8537, N7646);
or OR3 (N9103, N9086, N341, N5673);
buf BUF1 (N9104, N9103);
buf BUF1 (N9105, N9098);
and AND2 (N9106, N9096, N6810);
buf BUF1 (N9107, N9105);
nand NAND2 (N9108, N9102, N4018);
nor NOR2 (N9109, N9074, N6927);
and AND4 (N9110, N9101, N5637, N4818, N2801);
buf BUF1 (N9111, N9097);
nand NAND4 (N9112, N9104, N5116, N5632, N7250);
buf BUF1 (N9113, N9111);
nand NAND2 (N9114, N9110, N7440);
xor XOR2 (N9115, N9113, N4146);
xor XOR2 (N9116, N9106, N3568);
nand NAND2 (N9117, N9107, N1008);
or OR3 (N9118, N9112, N2801, N3860);
not NOT1 (N9119, N9100);
xor XOR2 (N9120, N9119, N5878);
buf BUF1 (N9121, N9108);
nand NAND2 (N9122, N9099, N3554);
nor NOR3 (N9123, N9118, N3947, N9062);
nor NOR2 (N9124, N9116, N4699);
and AND2 (N9125, N9121, N599);
not NOT1 (N9126, N9120);
nor NOR2 (N9127, N9122, N7876);
and AND2 (N9128, N9123, N2836);
and AND3 (N9129, N9125, N6325, N6782);
or OR2 (N9130, N9129, N5861);
nand NAND4 (N9131, N9114, N5747, N459, N2950);
xor XOR2 (N9132, N9109, N7743);
not NOT1 (N9133, N9131);
nand NAND3 (N9134, N9117, N1517, N3525);
not NOT1 (N9135, N9134);
and AND4 (N9136, N9133, N3953, N8583, N3692);
nor NOR4 (N9137, N9135, N502, N3457, N3389);
and AND2 (N9138, N9137, N8545);
not NOT1 (N9139, N9126);
and AND4 (N9140, N9094, N3706, N1102, N541);
nor NOR3 (N9141, N9130, N9018, N3922);
nor NOR2 (N9142, N9141, N6676);
buf BUF1 (N9143, N9128);
xor XOR2 (N9144, N9140, N8735);
nor NOR4 (N9145, N9144, N717, N2804, N6804);
or OR3 (N9146, N9143, N366, N908);
xor XOR2 (N9147, N9139, N3523);
nand NAND3 (N9148, N9142, N8811, N2418);
nor NOR2 (N9149, N9132, N4981);
buf BUF1 (N9150, N9149);
not NOT1 (N9151, N9138);
and AND4 (N9152, N9115, N406, N2920, N8329);
not NOT1 (N9153, N9136);
and AND3 (N9154, N9151, N4395, N2064);
or OR4 (N9155, N9148, N5125, N8475, N1036);
nand NAND4 (N9156, N9150, N4354, N8959, N3631);
buf BUF1 (N9157, N9146);
and AND4 (N9158, N9156, N7416, N367, N4205);
and AND3 (N9159, N9147, N3448, N3273);
not NOT1 (N9160, N9159);
or OR4 (N9161, N9153, N8357, N7994, N933);
not NOT1 (N9162, N9160);
nor NOR4 (N9163, N9155, N1822, N7054, N861);
nor NOR3 (N9164, N9157, N22, N614);
nand NAND2 (N9165, N9124, N7546);
not NOT1 (N9166, N9165);
xor XOR2 (N9167, N9161, N1660);
nand NAND4 (N9168, N9163, N7876, N5259, N3787);
and AND3 (N9169, N9152, N6222, N4983);
or OR4 (N9170, N9167, N2624, N2746, N7954);
not NOT1 (N9171, N9127);
buf BUF1 (N9172, N9171);
or OR4 (N9173, N9154, N7134, N6415, N8869);
xor XOR2 (N9174, N9145, N2587);
not NOT1 (N9175, N9162);
xor XOR2 (N9176, N9170, N4382);
and AND2 (N9177, N9168, N5408);
nor NOR3 (N9178, N9173, N5631, N3268);
and AND3 (N9179, N9158, N8002, N312);
xor XOR2 (N9180, N9177, N4407);
or OR3 (N9181, N9172, N7444, N8588);
and AND4 (N9182, N9164, N3411, N1650, N2895);
buf BUF1 (N9183, N9175);
nor NOR4 (N9184, N9182, N2285, N5309, N4319);
xor XOR2 (N9185, N9181, N4305);
or OR2 (N9186, N9166, N2314);
nand NAND3 (N9187, N9184, N3581, N2569);
xor XOR2 (N9188, N9179, N3941);
or OR2 (N9189, N9180, N4167);
nand NAND3 (N9190, N9187, N656, N633);
nand NAND4 (N9191, N9169, N8883, N7374, N8801);
nand NAND4 (N9192, N9183, N6965, N2163, N4883);
buf BUF1 (N9193, N9176);
xor XOR2 (N9194, N9178, N7027);
or OR4 (N9195, N9192, N4253, N6176, N1959);
or OR3 (N9196, N9193, N5090, N8432);
nand NAND3 (N9197, N9189, N4393, N2712);
nor NOR3 (N9198, N9174, N5758, N1144);
nand NAND3 (N9199, N9188, N2579, N4947);
buf BUF1 (N9200, N9198);
or OR3 (N9201, N9199, N8381, N1267);
nand NAND4 (N9202, N9191, N2637, N8829, N5320);
nor NOR4 (N9203, N9190, N4979, N4203, N7060);
buf BUF1 (N9204, N9203);
and AND4 (N9205, N9196, N9149, N3471, N8286);
nor NOR2 (N9206, N9195, N7802);
xor XOR2 (N9207, N9200, N9196);
xor XOR2 (N9208, N9206, N4125);
nor NOR4 (N9209, N9186, N3746, N6023, N3946);
nand NAND4 (N9210, N9204, N9117, N1166, N4675);
nor NOR3 (N9211, N9201, N825, N5912);
nand NAND4 (N9212, N9211, N424, N7345, N3244);
or OR2 (N9213, N9210, N2837);
nand NAND4 (N9214, N9205, N6282, N9117, N943);
buf BUF1 (N9215, N9207);
nand NAND4 (N9216, N9212, N7183, N1589, N4992);
nand NAND4 (N9217, N9213, N9037, N7295, N2741);
nor NOR3 (N9218, N9208, N4548, N7908);
or OR3 (N9219, N9214, N5350, N5557);
buf BUF1 (N9220, N9219);
or OR2 (N9221, N9209, N2158);
and AND3 (N9222, N9216, N5721, N3350);
buf BUF1 (N9223, N9220);
nand NAND4 (N9224, N9202, N7979, N3638, N9079);
nor NOR3 (N9225, N9185, N5533, N896);
not NOT1 (N9226, N9197);
not NOT1 (N9227, N9194);
and AND2 (N9228, N9218, N5904);
xor XOR2 (N9229, N9226, N7514);
buf BUF1 (N9230, N9224);
buf BUF1 (N9231, N9217);
xor XOR2 (N9232, N9231, N1078);
not NOT1 (N9233, N9227);
nand NAND2 (N9234, N9228, N9036);
buf BUF1 (N9235, N9234);
not NOT1 (N9236, N9221);
not NOT1 (N9237, N9222);
xor XOR2 (N9238, N9223, N2367);
nor NOR3 (N9239, N9235, N8997, N3417);
buf BUF1 (N9240, N9232);
or OR4 (N9241, N9237, N233, N761, N5802);
or OR3 (N9242, N9225, N3355, N4921);
or OR4 (N9243, N9239, N1569, N8682, N5831);
xor XOR2 (N9244, N9241, N8650);
buf BUF1 (N9245, N9229);
and AND3 (N9246, N9243, N6561, N3729);
buf BUF1 (N9247, N9244);
or OR2 (N9248, N9246, N3905);
and AND3 (N9249, N9215, N2164, N5235);
or OR4 (N9250, N9236, N142, N6006, N1503);
or OR3 (N9251, N9242, N1294, N2905);
and AND2 (N9252, N9247, N876);
not NOT1 (N9253, N9251);
or OR2 (N9254, N9238, N3397);
and AND4 (N9255, N9230, N1903, N5829, N1832);
and AND3 (N9256, N9250, N8857, N1558);
nand NAND3 (N9257, N9255, N9088, N785);
or OR4 (N9258, N9252, N7173, N322, N6406);
and AND4 (N9259, N9258, N6418, N7792, N4486);
nor NOR3 (N9260, N9253, N6142, N8744);
xor XOR2 (N9261, N9249, N5037);
buf BUF1 (N9262, N9240);
not NOT1 (N9263, N9233);
xor XOR2 (N9264, N9254, N3761);
buf BUF1 (N9265, N9248);
nor NOR2 (N9266, N9264, N8765);
and AND2 (N9267, N9263, N9159);
nor NOR3 (N9268, N9245, N5183, N4440);
xor XOR2 (N9269, N9261, N265);
nand NAND4 (N9270, N9269, N4791, N8649, N3924);
or OR4 (N9271, N9266, N5874, N113, N2831);
nand NAND2 (N9272, N9270, N4992);
buf BUF1 (N9273, N9265);
not NOT1 (N9274, N9260);
nand NAND4 (N9275, N9257, N6501, N3295, N147);
nor NOR2 (N9276, N9262, N1864);
buf BUF1 (N9277, N9275);
xor XOR2 (N9278, N9276, N7995);
or OR4 (N9279, N9278, N3315, N9031, N313);
xor XOR2 (N9280, N9272, N6693);
nor NOR4 (N9281, N9274, N7362, N6146, N7198);
not NOT1 (N9282, N9256);
and AND3 (N9283, N9271, N7247, N5019);
xor XOR2 (N9284, N9268, N853);
xor XOR2 (N9285, N9279, N2955);
not NOT1 (N9286, N9259);
not NOT1 (N9287, N9273);
nor NOR3 (N9288, N9287, N40, N1028);
buf BUF1 (N9289, N9285);
and AND2 (N9290, N9280, N6250);
buf BUF1 (N9291, N9289);
xor XOR2 (N9292, N9291, N5515);
not NOT1 (N9293, N9292);
nand NAND2 (N9294, N9290, N8092);
or OR3 (N9295, N9267, N9125, N5167);
or OR2 (N9296, N9284, N3747);
xor XOR2 (N9297, N9295, N8340);
not NOT1 (N9298, N9281);
nor NOR3 (N9299, N9283, N3123, N2764);
buf BUF1 (N9300, N9288);
or OR2 (N9301, N9296, N6460);
or OR2 (N9302, N9282, N3809);
or OR4 (N9303, N9298, N4922, N6807, N3660);
nand NAND2 (N9304, N9293, N7259);
not NOT1 (N9305, N9300);
buf BUF1 (N9306, N9277);
nand NAND4 (N9307, N9286, N3221, N1430, N5138);
not NOT1 (N9308, N9305);
nand NAND2 (N9309, N9302, N5785);
nand NAND2 (N9310, N9294, N5557);
buf BUF1 (N9311, N9308);
or OR4 (N9312, N9310, N2322, N3272, N6296);
not NOT1 (N9313, N9309);
not NOT1 (N9314, N9301);
buf BUF1 (N9315, N9299);
not NOT1 (N9316, N9297);
buf BUF1 (N9317, N9306);
xor XOR2 (N9318, N9316, N1497);
not NOT1 (N9319, N9303);
or OR2 (N9320, N9304, N1346);
buf BUF1 (N9321, N9317);
xor XOR2 (N9322, N9321, N4737);
not NOT1 (N9323, N9313);
nor NOR4 (N9324, N9307, N1032, N3642, N3934);
xor XOR2 (N9325, N9311, N4984);
not NOT1 (N9326, N9323);
and AND4 (N9327, N9325, N8230, N4126, N6514);
buf BUF1 (N9328, N9319);
nor NOR2 (N9329, N9312, N8293);
buf BUF1 (N9330, N9329);
and AND3 (N9331, N9326, N2935, N878);
nor NOR2 (N9332, N9331, N3274);
nor NOR4 (N9333, N9315, N8620, N5573, N1406);
nor NOR2 (N9334, N9332, N8633);
buf BUF1 (N9335, N9333);
nand NAND3 (N9336, N9322, N7103, N3224);
nand NAND2 (N9337, N9334, N3501);
nand NAND3 (N9338, N9330, N1855, N3997);
buf BUF1 (N9339, N9335);
and AND2 (N9340, N9327, N8390);
xor XOR2 (N9341, N9338, N5574);
or OR4 (N9342, N9328, N8064, N729, N4627);
not NOT1 (N9343, N9318);
nor NOR2 (N9344, N9342, N3083);
or OR4 (N9345, N9324, N1177, N6409, N6753);
and AND4 (N9346, N9345, N7768, N3413, N6523);
buf BUF1 (N9347, N9341);
nor NOR3 (N9348, N9344, N6143, N2749);
or OR2 (N9349, N9336, N6289);
xor XOR2 (N9350, N9339, N5306);
nand NAND4 (N9351, N9340, N1607, N5735, N1744);
nor NOR3 (N9352, N9320, N7820, N1742);
nand NAND2 (N9353, N9343, N1326);
not NOT1 (N9354, N9346);
buf BUF1 (N9355, N9352);
nor NOR4 (N9356, N9347, N6627, N6660, N5155);
or OR3 (N9357, N9337, N5194, N7023);
nor NOR2 (N9358, N9351, N844);
xor XOR2 (N9359, N9358, N6567);
or OR2 (N9360, N9353, N5770);
or OR2 (N9361, N9355, N2269);
nor NOR2 (N9362, N9359, N4273);
not NOT1 (N9363, N9360);
xor XOR2 (N9364, N9356, N6487);
nand NAND4 (N9365, N9350, N82, N8359, N3848);
not NOT1 (N9366, N9361);
xor XOR2 (N9367, N9366, N3774);
nor NOR2 (N9368, N9367, N6633);
and AND2 (N9369, N9354, N633);
not NOT1 (N9370, N9362);
buf BUF1 (N9371, N9365);
or OR4 (N9372, N9368, N8546, N7026, N1616);
or OR4 (N9373, N9357, N266, N6376, N5328);
not NOT1 (N9374, N9373);
buf BUF1 (N9375, N9348);
or OR4 (N9376, N9372, N2841, N1155, N6213);
nand NAND3 (N9377, N9370, N6254, N3178);
or OR3 (N9378, N9363, N8185, N7409);
and AND4 (N9379, N9314, N3319, N1069, N1965);
nand NAND4 (N9380, N9364, N2083, N1379, N449);
or OR2 (N9381, N9380, N8941);
nand NAND3 (N9382, N9377, N7303, N695);
nor NOR3 (N9383, N9381, N902, N5380);
xor XOR2 (N9384, N9382, N8203);
xor XOR2 (N9385, N9369, N7360);
not NOT1 (N9386, N9383);
not NOT1 (N9387, N9371);
nand NAND3 (N9388, N9386, N7107, N1011);
nor NOR2 (N9389, N9349, N4830);
not NOT1 (N9390, N9374);
buf BUF1 (N9391, N9388);
buf BUF1 (N9392, N9385);
and AND4 (N9393, N9378, N7245, N1721, N2364);
xor XOR2 (N9394, N9389, N7903);
nand NAND3 (N9395, N9394, N1134, N4342);
not NOT1 (N9396, N9387);
not NOT1 (N9397, N9393);
nand NAND3 (N9398, N9390, N4420, N6877);
or OR4 (N9399, N9376, N8995, N6964, N3854);
not NOT1 (N9400, N9375);
and AND2 (N9401, N9395, N1210);
nor NOR4 (N9402, N9398, N3750, N7902, N7970);
xor XOR2 (N9403, N9401, N6344);
xor XOR2 (N9404, N9391, N7243);
nor NOR3 (N9405, N9399, N7429, N8317);
nor NOR3 (N9406, N9404, N864, N5206);
not NOT1 (N9407, N9396);
xor XOR2 (N9408, N9402, N436);
not NOT1 (N9409, N9400);
not NOT1 (N9410, N9406);
nand NAND4 (N9411, N9405, N382, N8081, N5222);
nor NOR2 (N9412, N9408, N6546);
nand NAND3 (N9413, N9409, N7039, N2863);
not NOT1 (N9414, N9397);
buf BUF1 (N9415, N9414);
and AND4 (N9416, N9392, N2590, N4592, N7399);
buf BUF1 (N9417, N9384);
or OR4 (N9418, N9417, N3900, N435, N4497);
and AND4 (N9419, N9416, N3357, N2544, N3954);
nor NOR4 (N9420, N9419, N7627, N5419, N8245);
and AND4 (N9421, N9413, N705, N5843, N5140);
or OR2 (N9422, N9420, N8387);
nand NAND2 (N9423, N9412, N5820);
buf BUF1 (N9424, N9421);
not NOT1 (N9425, N9422);
and AND2 (N9426, N9379, N8258);
or OR3 (N9427, N9411, N4698, N1096);
not NOT1 (N9428, N9403);
and AND4 (N9429, N9415, N6744, N8496, N6502);
buf BUF1 (N9430, N9410);
and AND4 (N9431, N9430, N1694, N3701, N8982);
nand NAND2 (N9432, N9429, N3461);
buf BUF1 (N9433, N9428);
xor XOR2 (N9434, N9432, N5889);
buf BUF1 (N9435, N9418);
and AND3 (N9436, N9427, N1073, N2493);
and AND2 (N9437, N9426, N7170);
not NOT1 (N9438, N9435);
nor NOR2 (N9439, N9407, N6344);
not NOT1 (N9440, N9436);
and AND3 (N9441, N9439, N3326, N4945);
not NOT1 (N9442, N9438);
nand NAND3 (N9443, N9441, N6458, N6389);
or OR2 (N9444, N9437, N211);
xor XOR2 (N9445, N9424, N2746);
buf BUF1 (N9446, N9433);
xor XOR2 (N9447, N9440, N935);
nor NOR4 (N9448, N9444, N923, N7007, N4223);
xor XOR2 (N9449, N9443, N3788);
not NOT1 (N9450, N9448);
buf BUF1 (N9451, N9447);
or OR3 (N9452, N9451, N3019, N6256);
buf BUF1 (N9453, N9445);
xor XOR2 (N9454, N9446, N2408);
not NOT1 (N9455, N9431);
buf BUF1 (N9456, N9423);
or OR2 (N9457, N9450, N3227);
buf BUF1 (N9458, N9453);
nand NAND2 (N9459, N9449, N7045);
or OR2 (N9460, N9454, N7868);
nand NAND2 (N9461, N9452, N9226);
buf BUF1 (N9462, N9434);
not NOT1 (N9463, N9459);
not NOT1 (N9464, N9458);
xor XOR2 (N9465, N9460, N498);
and AND3 (N9466, N9425, N8350, N1110);
xor XOR2 (N9467, N9463, N4868);
xor XOR2 (N9468, N9464, N2128);
buf BUF1 (N9469, N9468);
xor XOR2 (N9470, N9457, N2489);
not NOT1 (N9471, N9465);
and AND4 (N9472, N9461, N5773, N6974, N4016);
and AND3 (N9473, N9456, N5632, N3728);
xor XOR2 (N9474, N9471, N3647);
nand NAND4 (N9475, N9472, N3704, N7683, N6766);
and AND4 (N9476, N9473, N8259, N5003, N922);
nand NAND3 (N9477, N9467, N5614, N9087);
xor XOR2 (N9478, N9466, N3058);
buf BUF1 (N9479, N9476);
not NOT1 (N9480, N9469);
or OR2 (N9481, N9477, N8780);
or OR4 (N9482, N9479, N4137, N9268, N2759);
and AND4 (N9483, N9470, N1056, N874, N3832);
and AND2 (N9484, N9442, N1841);
or OR3 (N9485, N9483, N4903, N2243);
or OR3 (N9486, N9462, N7063, N7097);
buf BUF1 (N9487, N9475);
nor NOR3 (N9488, N9482, N8897, N2482);
buf BUF1 (N9489, N9487);
nor NOR2 (N9490, N9484, N6781);
not NOT1 (N9491, N9488);
buf BUF1 (N9492, N9455);
not NOT1 (N9493, N9486);
nor NOR4 (N9494, N9478, N7726, N4030, N4107);
nor NOR3 (N9495, N9494, N2166, N8517);
not NOT1 (N9496, N9490);
not NOT1 (N9497, N9493);
buf BUF1 (N9498, N9495);
and AND4 (N9499, N9481, N6572, N385, N6099);
buf BUF1 (N9500, N9474);
xor XOR2 (N9501, N9500, N4408);
or OR4 (N9502, N9497, N4505, N2642, N7914);
not NOT1 (N9503, N9485);
xor XOR2 (N9504, N9492, N687);
nor NOR2 (N9505, N9502, N4953);
or OR3 (N9506, N9505, N1988, N6287);
or OR2 (N9507, N9506, N9112);
nor NOR4 (N9508, N9507, N4571, N7131, N2699);
not NOT1 (N9509, N9496);
or OR2 (N9510, N9491, N5941);
buf BUF1 (N9511, N9489);
buf BUF1 (N9512, N9510);
and AND3 (N9513, N9498, N4913, N7374);
and AND4 (N9514, N9501, N6229, N4589, N1069);
nand NAND4 (N9515, N9503, N2617, N1154, N857);
or OR2 (N9516, N9512, N1680);
nor NOR2 (N9517, N9514, N9186);
nor NOR3 (N9518, N9511, N8517, N577);
nand NAND2 (N9519, N9516, N7279);
nor NOR2 (N9520, N9508, N110);
not NOT1 (N9521, N9517);
buf BUF1 (N9522, N9521);
not NOT1 (N9523, N9519);
not NOT1 (N9524, N9499);
nor NOR4 (N9525, N9513, N8166, N4703, N7325);
nor NOR3 (N9526, N9520, N5231, N6814);
nor NOR4 (N9527, N9515, N2156, N4166, N6155);
nand NAND4 (N9528, N9526, N5636, N4325, N2494);
or OR2 (N9529, N9528, N8888);
nor NOR3 (N9530, N9480, N7095, N7598);
and AND2 (N9531, N9522, N3069);
and AND4 (N9532, N9509, N5056, N1880, N7449);
buf BUF1 (N9533, N9530);
buf BUF1 (N9534, N9523);
not NOT1 (N9535, N9534);
nor NOR2 (N9536, N9532, N1431);
xor XOR2 (N9537, N9524, N8336);
nor NOR4 (N9538, N9531, N1488, N7533, N5099);
xor XOR2 (N9539, N9533, N7818);
xor XOR2 (N9540, N9525, N249);
and AND2 (N9541, N9527, N219);
or OR4 (N9542, N9536, N3136, N4707, N2653);
or OR4 (N9543, N9504, N1942, N7468, N5402);
and AND2 (N9544, N9538, N2081);
not NOT1 (N9545, N9541);
or OR2 (N9546, N9539, N7980);
buf BUF1 (N9547, N9545);
or OR2 (N9548, N9535, N5925);
and AND4 (N9549, N9547, N2640, N7950, N807);
nor NOR2 (N9550, N9544, N3365);
and AND2 (N9551, N9518, N6790);
xor XOR2 (N9552, N9543, N3857);
nand NAND2 (N9553, N9529, N1670);
or OR3 (N9554, N9550, N1932, N6775);
nand NAND3 (N9555, N9553, N6346, N467);
xor XOR2 (N9556, N9542, N8864);
not NOT1 (N9557, N9549);
buf BUF1 (N9558, N9556);
xor XOR2 (N9559, N9540, N5695);
and AND3 (N9560, N9552, N1689, N3481);
xor XOR2 (N9561, N9548, N3108);
not NOT1 (N9562, N9558);
buf BUF1 (N9563, N9554);
xor XOR2 (N9564, N9561, N2157);
not NOT1 (N9565, N9551);
nand NAND3 (N9566, N9565, N384, N8256);
or OR3 (N9567, N9560, N274, N9552);
nor NOR4 (N9568, N9562, N8754, N5911, N1064);
not NOT1 (N9569, N9564);
nand NAND2 (N9570, N9557, N4465);
or OR2 (N9571, N9563, N8078);
buf BUF1 (N9572, N9569);
nand NAND4 (N9573, N9568, N2867, N8204, N6536);
buf BUF1 (N9574, N9555);
or OR3 (N9575, N9572, N5250, N632);
or OR3 (N9576, N9546, N5776, N4256);
buf BUF1 (N9577, N9567);
xor XOR2 (N9578, N9566, N1505);
nand NAND3 (N9579, N9571, N4419, N7665);
buf BUF1 (N9580, N9577);
xor XOR2 (N9581, N9576, N4455);
nand NAND4 (N9582, N9573, N5780, N8689, N7098);
xor XOR2 (N9583, N9580, N7440);
nand NAND3 (N9584, N9570, N3396, N6930);
nand NAND3 (N9585, N9583, N1339, N2802);
nand NAND3 (N9586, N9559, N4873, N362);
or OR3 (N9587, N9574, N2621, N8277);
xor XOR2 (N9588, N9584, N5950);
and AND2 (N9589, N9588, N6415);
or OR4 (N9590, N9585, N8903, N5563, N3371);
buf BUF1 (N9591, N9575);
or OR2 (N9592, N9590, N6866);
buf BUF1 (N9593, N9578);
nand NAND2 (N9594, N9582, N2042);
buf BUF1 (N9595, N9537);
buf BUF1 (N9596, N9579);
xor XOR2 (N9597, N9589, N4118);
not NOT1 (N9598, N9595);
not NOT1 (N9599, N9594);
xor XOR2 (N9600, N9593, N8459);
nor NOR4 (N9601, N9600, N7612, N6088, N57);
buf BUF1 (N9602, N9586);
and AND2 (N9603, N9598, N3992);
or OR3 (N9604, N9603, N4099, N1811);
not NOT1 (N9605, N9599);
or OR2 (N9606, N9605, N1908);
or OR2 (N9607, N9587, N5234);
nor NOR4 (N9608, N9581, N2855, N6398, N6960);
buf BUF1 (N9609, N9596);
xor XOR2 (N9610, N9607, N810);
nand NAND3 (N9611, N9606, N3665, N2506);
buf BUF1 (N9612, N9591);
nand NAND3 (N9613, N9601, N2408, N8712);
buf BUF1 (N9614, N9608);
nand NAND3 (N9615, N9614, N3761, N5837);
buf BUF1 (N9616, N9602);
and AND2 (N9617, N9609, N4002);
buf BUF1 (N9618, N9592);
and AND4 (N9619, N9597, N6319, N1027, N3202);
not NOT1 (N9620, N9619);
or OR2 (N9621, N9604, N4737);
xor XOR2 (N9622, N9618, N730);
nand NAND3 (N9623, N9616, N3688, N8198);
or OR3 (N9624, N9620, N7277, N7006);
nand NAND4 (N9625, N9624, N1215, N2472, N4440);
nand NAND3 (N9626, N9613, N6203, N528);
nand NAND2 (N9627, N9617, N2826);
xor XOR2 (N9628, N9623, N2709);
nand NAND4 (N9629, N9621, N9197, N6878, N2705);
nand NAND3 (N9630, N9629, N7717, N3790);
not NOT1 (N9631, N9628);
or OR2 (N9632, N9626, N2732);
nand NAND3 (N9633, N9622, N5974, N8586);
not NOT1 (N9634, N9615);
and AND4 (N9635, N9625, N5694, N2013, N4185);
and AND2 (N9636, N9634, N4047);
and AND3 (N9637, N9632, N3356, N8469);
and AND4 (N9638, N9637, N3931, N3000, N8946);
and AND2 (N9639, N9638, N6375);
nand NAND4 (N9640, N9639, N86, N7407, N5276);
nor NOR4 (N9641, N9640, N1179, N6879, N8806);
nor NOR4 (N9642, N9641, N7725, N5966, N7232);
nor NOR3 (N9643, N9627, N1614, N7958);
nand NAND4 (N9644, N9610, N283, N4390, N2796);
xor XOR2 (N9645, N9636, N962);
nand NAND4 (N9646, N9612, N5907, N2890, N1512);
and AND3 (N9647, N9635, N2765, N913);
and AND3 (N9648, N9646, N5147, N4107);
and AND2 (N9649, N9631, N1684);
and AND4 (N9650, N9645, N2232, N505, N6680);
not NOT1 (N9651, N9611);
nor NOR4 (N9652, N9649, N2786, N9055, N5896);
xor XOR2 (N9653, N9643, N4240);
xor XOR2 (N9654, N9651, N5862);
xor XOR2 (N9655, N9630, N1000);
xor XOR2 (N9656, N9648, N2701);
nor NOR4 (N9657, N9647, N6556, N7468, N2210);
buf BUF1 (N9658, N9652);
nor NOR4 (N9659, N9657, N1694, N7755, N5823);
nor NOR4 (N9660, N9633, N5697, N1068, N8524);
xor XOR2 (N9661, N9642, N3200);
and AND3 (N9662, N9660, N8383, N2414);
and AND4 (N9663, N9656, N6236, N4028, N5785);
xor XOR2 (N9664, N9653, N790);
nor NOR3 (N9665, N9658, N4292, N6536);
not NOT1 (N9666, N9664);
nand NAND4 (N9667, N9661, N5038, N178, N2160);
buf BUF1 (N9668, N9665);
and AND4 (N9669, N9654, N4184, N4998, N446);
and AND3 (N9670, N9644, N5520, N6711);
xor XOR2 (N9671, N9662, N5623);
nor NOR4 (N9672, N9650, N2984, N1357, N6315);
nand NAND4 (N9673, N9669, N2664, N1250, N4765);
nand NAND2 (N9674, N9663, N4710);
not NOT1 (N9675, N9672);
buf BUF1 (N9676, N9666);
buf BUF1 (N9677, N9670);
xor XOR2 (N9678, N9676, N3170);
and AND3 (N9679, N9674, N5174, N8200);
xor XOR2 (N9680, N9671, N5565);
or OR4 (N9681, N9673, N6428, N7308, N4106);
buf BUF1 (N9682, N9668);
buf BUF1 (N9683, N9667);
buf BUF1 (N9684, N9681);
and AND2 (N9685, N9682, N8062);
nand NAND3 (N9686, N9675, N2565, N5927);
nand NAND4 (N9687, N9659, N4747, N5802, N7777);
not NOT1 (N9688, N9684);
xor XOR2 (N9689, N9688, N3108);
nand NAND2 (N9690, N9686, N8105);
or OR3 (N9691, N9690, N4732, N7087);
xor XOR2 (N9692, N9679, N2951);
or OR4 (N9693, N9683, N9587, N8878, N6187);
xor XOR2 (N9694, N9685, N3032);
xor XOR2 (N9695, N9677, N6875);
and AND3 (N9696, N9693, N5414, N5253);
buf BUF1 (N9697, N9655);
not NOT1 (N9698, N9694);
buf BUF1 (N9699, N9698);
not NOT1 (N9700, N9687);
or OR3 (N9701, N9680, N8610, N4890);
not NOT1 (N9702, N9701);
and AND4 (N9703, N9678, N7149, N5724, N5463);
and AND3 (N9704, N9703, N4669, N7578);
or OR3 (N9705, N9689, N7527, N4804);
or OR3 (N9706, N9697, N3933, N7260);
nor NOR2 (N9707, N9702, N2857);
not NOT1 (N9708, N9700);
buf BUF1 (N9709, N9704);
and AND2 (N9710, N9696, N7487);
not NOT1 (N9711, N9706);
nand NAND4 (N9712, N9710, N2799, N4723, N3272);
buf BUF1 (N9713, N9708);
buf BUF1 (N9714, N9713);
nor NOR2 (N9715, N9707, N7192);
nor NOR3 (N9716, N9699, N6507, N6773);
nand NAND2 (N9717, N9715, N1972);
buf BUF1 (N9718, N9717);
nor NOR2 (N9719, N9714, N5977);
buf BUF1 (N9720, N9709);
nor NOR3 (N9721, N9705, N4270, N2240);
or OR2 (N9722, N9695, N2728);
buf BUF1 (N9723, N9716);
buf BUF1 (N9724, N9720);
nand NAND4 (N9725, N9712, N156, N6416, N7366);
not NOT1 (N9726, N9718);
or OR3 (N9727, N9721, N2864, N5956);
and AND4 (N9728, N9723, N6628, N7041, N6560);
buf BUF1 (N9729, N9722);
xor XOR2 (N9730, N9725, N8677);
or OR2 (N9731, N9692, N7270);
or OR2 (N9732, N9726, N5421);
not NOT1 (N9733, N9719);
not NOT1 (N9734, N9731);
and AND3 (N9735, N9727, N4730, N787);
nor NOR3 (N9736, N9734, N2972, N5328);
not NOT1 (N9737, N9711);
or OR2 (N9738, N9729, N2242);
buf BUF1 (N9739, N9737);
or OR3 (N9740, N9691, N8144, N5863);
nor NOR4 (N9741, N9728, N3476, N2804, N343);
nor NOR2 (N9742, N9735, N1940);
buf BUF1 (N9743, N9736);
buf BUF1 (N9744, N9740);
or OR2 (N9745, N9739, N1053);
not NOT1 (N9746, N9742);
and AND3 (N9747, N9733, N980, N2718);
xor XOR2 (N9748, N9732, N7532);
not NOT1 (N9749, N9743);
not NOT1 (N9750, N9730);
nand NAND4 (N9751, N9741, N6063, N8520, N9282);
or OR2 (N9752, N9748, N690);
not NOT1 (N9753, N9752);
nand NAND2 (N9754, N9749, N343);
nand NAND3 (N9755, N9745, N6080, N3686);
xor XOR2 (N9756, N9724, N2792);
nor NOR4 (N9757, N9753, N145, N6, N4338);
nor NOR2 (N9758, N9744, N112);
not NOT1 (N9759, N9738);
not NOT1 (N9760, N9751);
not NOT1 (N9761, N9759);
buf BUF1 (N9762, N9757);
or OR4 (N9763, N9762, N6098, N4973, N3821);
not NOT1 (N9764, N9750);
buf BUF1 (N9765, N9754);
and AND4 (N9766, N9764, N5188, N746, N5377);
nand NAND4 (N9767, N9763, N2080, N9534, N8794);
buf BUF1 (N9768, N9766);
or OR2 (N9769, N9767, N5372);
xor XOR2 (N9770, N9761, N3056);
or OR2 (N9771, N9758, N8674);
not NOT1 (N9772, N9755);
nor NOR4 (N9773, N9756, N2683, N8862, N2530);
or OR2 (N9774, N9769, N2806);
or OR3 (N9775, N9747, N5221, N5832);
nor NOR2 (N9776, N9746, N9114);
or OR3 (N9777, N9775, N9144, N2282);
not NOT1 (N9778, N9771);
xor XOR2 (N9779, N9770, N3300);
nor NOR3 (N9780, N9777, N9560, N2687);
and AND3 (N9781, N9768, N4190, N2325);
nor NOR4 (N9782, N9776, N3765, N8611, N1198);
or OR2 (N9783, N9760, N4937);
and AND2 (N9784, N9781, N3970);
nand NAND2 (N9785, N9778, N8527);
not NOT1 (N9786, N9774);
buf BUF1 (N9787, N9779);
buf BUF1 (N9788, N9783);
or OR2 (N9789, N9772, N883);
and AND2 (N9790, N9786, N5248);
or OR4 (N9791, N9789, N7528, N4562, N8852);
not NOT1 (N9792, N9788);
and AND3 (N9793, N9782, N5432, N3492);
nand NAND2 (N9794, N9780, N5507);
buf BUF1 (N9795, N9784);
nor NOR4 (N9796, N9795, N4527, N9431, N8686);
nor NOR2 (N9797, N9790, N5115);
xor XOR2 (N9798, N9794, N4895);
nand NAND3 (N9799, N9785, N2351, N3598);
nor NOR2 (N9800, N9796, N7356);
not NOT1 (N9801, N9799);
and AND3 (N9802, N9792, N4470, N4326);
or OR2 (N9803, N9773, N1669);
nor NOR2 (N9804, N9801, N2927);
buf BUF1 (N9805, N9797);
buf BUF1 (N9806, N9798);
xor XOR2 (N9807, N9800, N5457);
buf BUF1 (N9808, N9804);
or OR4 (N9809, N9803, N1074, N4743, N8873);
not NOT1 (N9810, N9791);
nor NOR4 (N9811, N9807, N2576, N4812, N5929);
buf BUF1 (N9812, N9765);
buf BUF1 (N9813, N9812);
not NOT1 (N9814, N9793);
buf BUF1 (N9815, N9808);
xor XOR2 (N9816, N9811, N2470);
and AND3 (N9817, N9813, N6421, N7020);
not NOT1 (N9818, N9814);
or OR2 (N9819, N9817, N8055);
not NOT1 (N9820, N9787);
or OR3 (N9821, N9809, N9338, N7319);
buf BUF1 (N9822, N9815);
nor NOR2 (N9823, N9816, N4302);
nand NAND3 (N9824, N9802, N4860, N4452);
or OR2 (N9825, N9810, N8568);
and AND4 (N9826, N9825, N113, N3295, N554);
buf BUF1 (N9827, N9826);
xor XOR2 (N9828, N9818, N8362);
and AND2 (N9829, N9822, N6475);
xor XOR2 (N9830, N9828, N7647);
nand NAND3 (N9831, N9823, N2722, N3200);
nand NAND2 (N9832, N9831, N2976);
nand NAND4 (N9833, N9832, N3662, N8064, N4461);
or OR4 (N9834, N9821, N3818, N2648, N3951);
nand NAND3 (N9835, N9819, N8612, N4711);
or OR4 (N9836, N9820, N5791, N8078, N480);
xor XOR2 (N9837, N9829, N1263);
nand NAND3 (N9838, N9835, N7877, N7522);
nor NOR4 (N9839, N9838, N2220, N9772, N9147);
buf BUF1 (N9840, N9834);
buf BUF1 (N9841, N9830);
xor XOR2 (N9842, N9840, N8879);
and AND2 (N9843, N9833, N951);
nor NOR4 (N9844, N9837, N9756, N3041, N8066);
buf BUF1 (N9845, N9806);
or OR2 (N9846, N9844, N5427);
xor XOR2 (N9847, N9839, N2417);
buf BUF1 (N9848, N9841);
or OR4 (N9849, N9843, N8320, N2838, N6293);
buf BUF1 (N9850, N9848);
buf BUF1 (N9851, N9836);
nand NAND3 (N9852, N9849, N4033, N9353);
and AND2 (N9853, N9824, N5502);
or OR2 (N9854, N9846, N1712);
nor NOR3 (N9855, N9847, N649, N943);
not NOT1 (N9856, N9805);
buf BUF1 (N9857, N9853);
or OR2 (N9858, N9852, N5603);
buf BUF1 (N9859, N9857);
xor XOR2 (N9860, N9859, N3326);
or OR4 (N9861, N9855, N6390, N9226, N6058);
nand NAND2 (N9862, N9842, N8035);
nor NOR4 (N9863, N9845, N9367, N6223, N5138);
or OR4 (N9864, N9862, N4638, N2915, N4759);
buf BUF1 (N9865, N9860);
or OR3 (N9866, N9827, N3487, N7144);
or OR3 (N9867, N9866, N3326, N4483);
nor NOR4 (N9868, N9863, N3110, N4010, N5002);
nand NAND4 (N9869, N9867, N3256, N2397, N4180);
xor XOR2 (N9870, N9850, N926);
xor XOR2 (N9871, N9870, N8847);
buf BUF1 (N9872, N9864);
or OR4 (N9873, N9869, N8209, N6627, N4929);
xor XOR2 (N9874, N9871, N3922);
and AND4 (N9875, N9861, N2232, N7370, N41);
nand NAND2 (N9876, N9865, N809);
nand NAND4 (N9877, N9868, N5518, N1532, N898);
and AND3 (N9878, N9856, N1839, N7052);
nand NAND4 (N9879, N9875, N9323, N5155, N3793);
xor XOR2 (N9880, N9877, N9403);
or OR2 (N9881, N9878, N616);
not NOT1 (N9882, N9876);
xor XOR2 (N9883, N9881, N1611);
buf BUF1 (N9884, N9882);
or OR2 (N9885, N9873, N6063);
and AND4 (N9886, N9851, N6039, N815, N1228);
xor XOR2 (N9887, N9858, N1492);
buf BUF1 (N9888, N9886);
nor NOR3 (N9889, N9885, N5584, N9287);
buf BUF1 (N9890, N9884);
buf BUF1 (N9891, N9887);
nand NAND3 (N9892, N9874, N8711, N7188);
not NOT1 (N9893, N9880);
nand NAND4 (N9894, N9888, N7718, N2324, N5397);
not NOT1 (N9895, N9890);
nor NOR3 (N9896, N9892, N3580, N4913);
xor XOR2 (N9897, N9889, N2551);
buf BUF1 (N9898, N9854);
nand NAND3 (N9899, N9883, N6714, N8771);
or OR3 (N9900, N9898, N4033, N893);
or OR2 (N9901, N9899, N2012);
buf BUF1 (N9902, N9872);
nor NOR3 (N9903, N9879, N4269, N6944);
or OR3 (N9904, N9893, N7196, N179);
xor XOR2 (N9905, N9891, N506);
or OR2 (N9906, N9903, N4567);
not NOT1 (N9907, N9896);
nor NOR3 (N9908, N9901, N1868, N9023);
buf BUF1 (N9909, N9906);
nand NAND2 (N9910, N9897, N7661);
and AND4 (N9911, N9895, N3805, N8799, N6070);
nor NOR4 (N9912, N9905, N3488, N6794, N5733);
and AND2 (N9913, N9904, N7410);
nor NOR3 (N9914, N9907, N9833, N3047);
not NOT1 (N9915, N9900);
and AND4 (N9916, N9914, N2741, N6675, N4623);
and AND3 (N9917, N9910, N1091, N7895);
nand NAND3 (N9918, N9894, N9194, N4806);
or OR2 (N9919, N9902, N9043);
nor NOR4 (N9920, N9919, N4812, N5820, N4015);
xor XOR2 (N9921, N9917, N56);
buf BUF1 (N9922, N9915);
or OR4 (N9923, N9911, N7992, N1749, N6269);
nand NAND2 (N9924, N9921, N8840);
or OR4 (N9925, N9912, N4464, N2021, N5741);
nand NAND4 (N9926, N9923, N7407, N4535, N6889);
xor XOR2 (N9927, N9918, N554);
or OR3 (N9928, N9926, N7123, N6689);
or OR4 (N9929, N9927, N6922, N6833, N960);
nand NAND4 (N9930, N9922, N215, N9382, N9412);
nand NAND3 (N9931, N9930, N6318, N418);
or OR4 (N9932, N9929, N7643, N6676, N8660);
buf BUF1 (N9933, N9913);
xor XOR2 (N9934, N9916, N6631);
and AND3 (N9935, N9933, N784, N5475);
and AND3 (N9936, N9935, N3166, N4371);
xor XOR2 (N9937, N9931, N9370);
nand NAND3 (N9938, N9937, N7029, N8051);
nand NAND3 (N9939, N9936, N3279, N4163);
nand NAND4 (N9940, N9934, N1369, N1801, N4365);
nor NOR2 (N9941, N9928, N1225);
and AND4 (N9942, N9908, N5254, N1741, N3586);
nand NAND4 (N9943, N9942, N504, N7812, N1486);
and AND3 (N9944, N9938, N5452, N5277);
nor NOR4 (N9945, N9940, N6141, N7746, N4945);
not NOT1 (N9946, N9945);
and AND2 (N9947, N9944, N7029);
nand NAND4 (N9948, N9924, N6706, N4926, N6749);
or OR3 (N9949, N9920, N9653, N4926);
buf BUF1 (N9950, N9939);
buf BUF1 (N9951, N9925);
nand NAND2 (N9952, N9948, N164);
xor XOR2 (N9953, N9943, N1033);
and AND2 (N9954, N9932, N6190);
xor XOR2 (N9955, N9954, N7792);
and AND3 (N9956, N9951, N412, N5472);
not NOT1 (N9957, N9950);
not NOT1 (N9958, N9957);
nand NAND3 (N9959, N9941, N1162, N4382);
xor XOR2 (N9960, N9959, N2703);
not NOT1 (N9961, N9947);
xor XOR2 (N9962, N9949, N2823);
or OR4 (N9963, N9955, N6315, N2204, N8406);
xor XOR2 (N9964, N9953, N9333);
nand NAND3 (N9965, N9961, N5789, N6835);
buf BUF1 (N9966, N9964);
or OR2 (N9967, N9966, N8806);
and AND2 (N9968, N9967, N2311);
and AND4 (N9969, N9946, N6868, N1516, N1863);
nand NAND2 (N9970, N9909, N879);
nand NAND3 (N9971, N9960, N4348, N1851);
not NOT1 (N9972, N9969);
or OR4 (N9973, N9956, N506, N3659, N6481);
and AND4 (N9974, N9972, N1823, N4212, N8387);
buf BUF1 (N9975, N9965);
xor XOR2 (N9976, N9975, N8333);
nand NAND4 (N9977, N9971, N387, N5727, N4523);
nor NOR4 (N9978, N9977, N6030, N9809, N1889);
and AND4 (N9979, N9974, N9424, N8973, N4613);
and AND3 (N9980, N9970, N3898, N2451);
buf BUF1 (N9981, N9962);
not NOT1 (N9982, N9979);
or OR4 (N9983, N9963, N7933, N4604, N5354);
buf BUF1 (N9984, N9982);
buf BUF1 (N9985, N9980);
not NOT1 (N9986, N9952);
xor XOR2 (N9987, N9983, N3900);
xor XOR2 (N9988, N9984, N1433);
nor NOR2 (N9989, N9973, N7785);
not NOT1 (N9990, N9968);
buf BUF1 (N9991, N9989);
buf BUF1 (N9992, N9990);
not NOT1 (N9993, N9991);
and AND2 (N9994, N9993, N9665);
nor NOR2 (N9995, N9958, N7234);
xor XOR2 (N9996, N9978, N4839);
xor XOR2 (N9997, N9976, N8469);
buf BUF1 (N9998, N9986);
nor NOR4 (N9999, N9988, N488, N3225, N2967);
nand NAND3 (N10000, N9992, N9666, N2676);
nor NOR2 (N10001, N9981, N9520);
nand NAND2 (N10002, N9985, N3221);
buf BUF1 (N10003, N9996);
xor XOR2 (N10004, N9998, N6019);
nor NOR2 (N10005, N9999, N274);
nor NOR3 (N10006, N9987, N6070, N9568);
or OR2 (N10007, N10004, N2601);
nand NAND4 (N10008, N10002, N3884, N2376, N3072);
and AND4 (N10009, N10000, N5059, N8177, N2357);
and AND3 (N10010, N9995, N5652, N6351);
and AND3 (N10011, N10003, N5853, N3027);
xor XOR2 (N10012, N10006, N1910);
nor NOR4 (N10013, N10005, N5634, N5361, N648);
buf BUF1 (N10014, N10007);
or OR2 (N10015, N10010, N6862);
nor NOR2 (N10016, N10012, N1495);
not NOT1 (N10017, N10016);
nand NAND4 (N10018, N10017, N6980, N4955, N5082);
not NOT1 (N10019, N10018);
not NOT1 (N10020, N9997);
not NOT1 (N10021, N10009);
buf BUF1 (N10022, N10019);
or OR3 (N10023, N10011, N3291, N8841);
xor XOR2 (N10024, N10023, N2145);
xor XOR2 (N10025, N10008, N5437);
and AND3 (N10026, N10025, N2259, N5316);
buf BUF1 (N10027, N10001);
and AND3 (N10028, N10014, N5862, N8317);
buf BUF1 (N10029, N9994);
nor NOR3 (N10030, N10026, N6804, N5573);
and AND2 (N10031, N10013, N9471);
xor XOR2 (N10032, N10015, N4929);
and AND3 (N10033, N10032, N1151, N5762);
nand NAND4 (N10034, N10027, N9673, N7129, N3262);
buf BUF1 (N10035, N10034);
or OR2 (N10036, N10021, N7878);
and AND4 (N10037, N10022, N9024, N1930, N5938);
buf BUF1 (N10038, N10028);
not NOT1 (N10039, N10036);
nand NAND4 (N10040, N10038, N8917, N9861, N4515);
buf BUF1 (N10041, N10040);
nor NOR3 (N10042, N10041, N5888, N5569);
buf BUF1 (N10043, N10030);
xor XOR2 (N10044, N10020, N9267);
not NOT1 (N10045, N10031);
not NOT1 (N10046, N10042);
or OR2 (N10047, N10033, N5634);
nand NAND3 (N10048, N10046, N7351, N7529);
or OR3 (N10049, N10045, N6159, N7445);
or OR4 (N10050, N10048, N6903, N5053, N6038);
not NOT1 (N10051, N10047);
or OR4 (N10052, N10051, N6397, N8823, N1047);
not NOT1 (N10053, N10050);
buf BUF1 (N10054, N10049);
and AND2 (N10055, N10037, N2101);
nand NAND4 (N10056, N10044, N8642, N4291, N3330);
buf BUF1 (N10057, N10029);
and AND4 (N10058, N10024, N1717, N1664, N9104);
nor NOR2 (N10059, N10043, N1755);
and AND2 (N10060, N10052, N7643);
not NOT1 (N10061, N10039);
buf BUF1 (N10062, N10061);
nand NAND4 (N10063, N10053, N2123, N1800, N2099);
not NOT1 (N10064, N10056);
not NOT1 (N10065, N10035);
and AND4 (N10066, N10054, N3402, N8595, N2636);
nor NOR2 (N10067, N10063, N9879);
nand NAND3 (N10068, N10064, N8261, N2082);
or OR4 (N10069, N10065, N8539, N8078, N8967);
buf BUF1 (N10070, N10057);
nand NAND3 (N10071, N10060, N6797, N4333);
and AND2 (N10072, N10068, N5778);
xor XOR2 (N10073, N10069, N3660);
and AND2 (N10074, N10058, N5461);
xor XOR2 (N10075, N10074, N4328);
or OR4 (N10076, N10062, N6973, N6684, N1610);
nor NOR2 (N10077, N10059, N8441);
or OR3 (N10078, N10067, N4906, N9922);
and AND2 (N10079, N10070, N1607);
buf BUF1 (N10080, N10076);
buf BUF1 (N10081, N10055);
xor XOR2 (N10082, N10066, N2977);
not NOT1 (N10083, N10077);
and AND4 (N10084, N10083, N7140, N9840, N9095);
nand NAND3 (N10085, N10082, N1832, N3715);
buf BUF1 (N10086, N10079);
buf BUF1 (N10087, N10081);
or OR2 (N10088, N10072, N6233);
or OR3 (N10089, N10075, N8266, N7285);
and AND2 (N10090, N10071, N9212);
or OR3 (N10091, N10080, N6092, N8835);
buf BUF1 (N10092, N10087);
and AND2 (N10093, N10091, N9475);
xor XOR2 (N10094, N10088, N6012);
nor NOR3 (N10095, N10073, N4863, N8547);
nand NAND4 (N10096, N10084, N9150, N6627, N4078);
nand NAND3 (N10097, N10089, N2999, N2503);
buf BUF1 (N10098, N10078);
and AND2 (N10099, N10097, N275);
buf BUF1 (N10100, N10093);
nor NOR2 (N10101, N10095, N385);
xor XOR2 (N10102, N10085, N8083);
nand NAND2 (N10103, N10100, N6183);
buf BUF1 (N10104, N10086);
nor NOR4 (N10105, N10092, N4152, N3052, N1038);
or OR3 (N10106, N10090, N3432, N5802);
and AND2 (N10107, N10096, N7292);
nor NOR4 (N10108, N10102, N4667, N7356, N4175);
xor XOR2 (N10109, N10103, N4010);
and AND3 (N10110, N10094, N6857, N8912);
or OR4 (N10111, N10108, N7571, N7366, N6791);
buf BUF1 (N10112, N10106);
nor NOR2 (N10113, N10111, N2413);
nor NOR3 (N10114, N10098, N9396, N8155);
buf BUF1 (N10115, N10112);
xor XOR2 (N10116, N10113, N3906);
nand NAND2 (N10117, N10105, N5864);
xor XOR2 (N10118, N10115, N1354);
or OR2 (N10119, N10114, N778);
or OR4 (N10120, N10104, N4173, N1419, N3970);
xor XOR2 (N10121, N10118, N9127);
not NOT1 (N10122, N10121);
and AND3 (N10123, N10122, N3488, N5273);
nor NOR2 (N10124, N10120, N2904);
not NOT1 (N10125, N10107);
not NOT1 (N10126, N10101);
nand NAND4 (N10127, N10123, N4541, N5658, N5104);
or OR4 (N10128, N10125, N4781, N7538, N3990);
or OR4 (N10129, N10124, N9964, N6039, N2305);
buf BUF1 (N10130, N10110);
or OR2 (N10131, N10128, N1610);
not NOT1 (N10132, N10117);
nor NOR3 (N10133, N10129, N4782, N5153);
or OR2 (N10134, N10119, N7697);
nand NAND3 (N10135, N10126, N8419, N6444);
and AND3 (N10136, N10109, N9149, N9328);
not NOT1 (N10137, N10136);
xor XOR2 (N10138, N10116, N659);
or OR2 (N10139, N10137, N3588);
nand NAND2 (N10140, N10139, N8601);
or OR2 (N10141, N10133, N6578);
and AND3 (N10142, N10138, N5200, N2096);
buf BUF1 (N10143, N10142);
and AND4 (N10144, N10130, N1970, N5487, N8854);
not NOT1 (N10145, N10143);
nor NOR4 (N10146, N10132, N4476, N7813, N3675);
nand NAND2 (N10147, N10145, N1820);
and AND4 (N10148, N10134, N2839, N1913, N1782);
buf BUF1 (N10149, N10131);
buf BUF1 (N10150, N10149);
not NOT1 (N10151, N10146);
nor NOR3 (N10152, N10150, N670, N1137);
not NOT1 (N10153, N10147);
nor NOR2 (N10154, N10152, N6863);
buf BUF1 (N10155, N10151);
or OR2 (N10156, N10127, N9025);
not NOT1 (N10157, N10156);
nand NAND3 (N10158, N10144, N1650, N8546);
buf BUF1 (N10159, N10135);
or OR2 (N10160, N10154, N4734);
or OR4 (N10161, N10160, N7531, N3606, N7807);
and AND3 (N10162, N10158, N5764, N7713);
and AND2 (N10163, N10157, N3444);
and AND2 (N10164, N10148, N7848);
buf BUF1 (N10165, N10140);
nand NAND4 (N10166, N10153, N2993, N4720, N1955);
buf BUF1 (N10167, N10161);
nor NOR4 (N10168, N10162, N709, N5772, N4111);
or OR4 (N10169, N10163, N1952, N739, N8589);
nor NOR2 (N10170, N10169, N4626);
or OR3 (N10171, N10155, N4082, N1492);
nor NOR2 (N10172, N10171, N10016);
buf BUF1 (N10173, N10168);
not NOT1 (N10174, N10159);
not NOT1 (N10175, N10174);
xor XOR2 (N10176, N10165, N9349);
or OR4 (N10177, N10166, N1839, N964, N279);
xor XOR2 (N10178, N10167, N6857);
not NOT1 (N10179, N10177);
nand NAND2 (N10180, N10175, N9123);
nor NOR3 (N10181, N10173, N6950, N9740);
nand NAND3 (N10182, N10164, N2768, N6513);
nor NOR2 (N10183, N10182, N6484);
and AND2 (N10184, N10099, N8355);
not NOT1 (N10185, N10172);
nor NOR2 (N10186, N10170, N6908);
buf BUF1 (N10187, N10180);
nand NAND4 (N10188, N10181, N4801, N1951, N3041);
xor XOR2 (N10189, N10178, N5219);
not NOT1 (N10190, N10184);
nor NOR3 (N10191, N10187, N2479, N5997);
or OR4 (N10192, N10190, N6732, N7568, N2668);
or OR2 (N10193, N10191, N4778);
not NOT1 (N10194, N10186);
xor XOR2 (N10195, N10185, N9893);
not NOT1 (N10196, N10193);
not NOT1 (N10197, N10141);
buf BUF1 (N10198, N10183);
xor XOR2 (N10199, N10197, N6978);
buf BUF1 (N10200, N10176);
buf BUF1 (N10201, N10179);
nor NOR3 (N10202, N10194, N4820, N5426);
and AND4 (N10203, N10196, N627, N6906, N9379);
buf BUF1 (N10204, N10201);
buf BUF1 (N10205, N10200);
buf BUF1 (N10206, N10192);
xor XOR2 (N10207, N10199, N4092);
not NOT1 (N10208, N10198);
and AND4 (N10209, N10206, N5540, N8903, N7098);
not NOT1 (N10210, N10195);
nor NOR4 (N10211, N10203, N7970, N4505, N3941);
buf BUF1 (N10212, N10210);
nand NAND3 (N10213, N10211, N5957, N4180);
not NOT1 (N10214, N10213);
buf BUF1 (N10215, N10207);
buf BUF1 (N10216, N10188);
nor NOR3 (N10217, N10202, N7317, N6553);
and AND2 (N10218, N10189, N5252);
xor XOR2 (N10219, N10216, N7270);
or OR4 (N10220, N10214, N6260, N7996, N1459);
nor NOR3 (N10221, N10208, N6409, N9474);
nor NOR3 (N10222, N10220, N2148, N1630);
nand NAND4 (N10223, N10219, N4546, N2260, N2933);
nor NOR3 (N10224, N10218, N1942, N669);
xor XOR2 (N10225, N10221, N4969);
and AND3 (N10226, N10209, N6358, N5437);
buf BUF1 (N10227, N10224);
nand NAND3 (N10228, N10227, N5760, N2634);
nand NAND4 (N10229, N10226, N9415, N6077, N2994);
not NOT1 (N10230, N10204);
nand NAND4 (N10231, N10230, N10110, N9388, N7273);
or OR3 (N10232, N10217, N2461, N7307);
or OR3 (N10233, N10212, N7715, N6133);
or OR4 (N10234, N10228, N9892, N3002, N2103);
nor NOR3 (N10235, N10223, N3848, N822);
buf BUF1 (N10236, N10205);
not NOT1 (N10237, N10233);
nor NOR4 (N10238, N10235, N7934, N8646, N7230);
nand NAND4 (N10239, N10231, N9331, N458, N7281);
and AND2 (N10240, N10238, N8386);
or OR2 (N10241, N10229, N2013);
buf BUF1 (N10242, N10225);
or OR3 (N10243, N10236, N3303, N9034);
or OR4 (N10244, N10234, N4103, N8482, N9757);
nor NOR2 (N10245, N10240, N2640);
nand NAND4 (N10246, N10232, N9097, N9782, N4749);
or OR3 (N10247, N10245, N3024, N6684);
not NOT1 (N10248, N10246);
xor XOR2 (N10249, N10244, N5591);
nor NOR3 (N10250, N10237, N8268, N9286);
not NOT1 (N10251, N10247);
and AND2 (N10252, N10215, N1492);
buf BUF1 (N10253, N10250);
xor XOR2 (N10254, N10253, N3333);
nor NOR3 (N10255, N10243, N2540, N775);
buf BUF1 (N10256, N10241);
buf BUF1 (N10257, N10255);
and AND4 (N10258, N10222, N1648, N5616, N9603);
not NOT1 (N10259, N10248);
nor NOR4 (N10260, N10239, N2273, N2953, N8528);
xor XOR2 (N10261, N10256, N9592);
and AND2 (N10262, N10257, N7685);
and AND2 (N10263, N10262, N7499);
not NOT1 (N10264, N10254);
xor XOR2 (N10265, N10252, N4545);
not NOT1 (N10266, N10258);
nor NOR3 (N10267, N10261, N9789, N10250);
nor NOR3 (N10268, N10249, N5060, N9558);
not NOT1 (N10269, N10242);
or OR3 (N10270, N10251, N4827, N6270);
not NOT1 (N10271, N10259);
nand NAND3 (N10272, N10264, N7494, N9053);
nand NAND4 (N10273, N10263, N6367, N187, N2321);
nor NOR2 (N10274, N10267, N9858);
or OR2 (N10275, N10272, N9688);
nand NAND3 (N10276, N10268, N10207, N7964);
buf BUF1 (N10277, N10260);
xor XOR2 (N10278, N10274, N7545);
not NOT1 (N10279, N10273);
xor XOR2 (N10280, N10275, N9593);
xor XOR2 (N10281, N10280, N1444);
xor XOR2 (N10282, N10276, N10134);
nand NAND2 (N10283, N10270, N6924);
nand NAND2 (N10284, N10278, N8364);
xor XOR2 (N10285, N10284, N9543);
nand NAND4 (N10286, N10283, N8545, N529, N7976);
and AND3 (N10287, N10282, N1114, N7523);
or OR2 (N10288, N10285, N6873);
and AND2 (N10289, N10288, N4520);
nand NAND4 (N10290, N10289, N2471, N1972, N4146);
nand NAND3 (N10291, N10279, N7268, N5298);
not NOT1 (N10292, N10291);
or OR3 (N10293, N10266, N6842, N6181);
or OR4 (N10294, N10269, N7758, N9274, N2742);
not NOT1 (N10295, N10277);
nor NOR4 (N10296, N10293, N2207, N6539, N141);
nor NOR4 (N10297, N10292, N3930, N5508, N5817);
nand NAND3 (N10298, N10271, N223, N9063);
or OR4 (N10299, N10287, N351, N2455, N1351);
not NOT1 (N10300, N10295);
buf BUF1 (N10301, N10286);
buf BUF1 (N10302, N10265);
buf BUF1 (N10303, N10298);
and AND3 (N10304, N10303, N6010, N7923);
not NOT1 (N10305, N10301);
nand NAND3 (N10306, N10294, N5322, N2666);
xor XOR2 (N10307, N10306, N3292);
and AND2 (N10308, N10290, N4139);
buf BUF1 (N10309, N10308);
xor XOR2 (N10310, N10297, N6345);
nand NAND2 (N10311, N10302, N3105);
nor NOR2 (N10312, N10300, N13);
or OR3 (N10313, N10310, N7906, N5865);
or OR2 (N10314, N10304, N2479);
nor NOR2 (N10315, N10311, N5974);
nor NOR2 (N10316, N10315, N6501);
nand NAND3 (N10317, N10316, N6499, N9059);
or OR3 (N10318, N10307, N4790, N7949);
nor NOR3 (N10319, N10281, N2120, N4847);
not NOT1 (N10320, N10312);
and AND3 (N10321, N10320, N8101, N6139);
xor XOR2 (N10322, N10299, N796);
nor NOR2 (N10323, N10313, N4955);
and AND4 (N10324, N10314, N6855, N3250, N3872);
not NOT1 (N10325, N10321);
buf BUF1 (N10326, N10322);
nor NOR2 (N10327, N10317, N4428);
xor XOR2 (N10328, N10318, N5656);
buf BUF1 (N10329, N10327);
not NOT1 (N10330, N10329);
xor XOR2 (N10331, N10309, N8138);
nand NAND3 (N10332, N10305, N5706, N2936);
buf BUF1 (N10333, N10326);
buf BUF1 (N10334, N10319);
nand NAND4 (N10335, N10325, N2820, N7467, N2983);
buf BUF1 (N10336, N10330);
buf BUF1 (N10337, N10331);
or OR2 (N10338, N10332, N7236);
nor NOR3 (N10339, N10338, N6620, N7933);
xor XOR2 (N10340, N10336, N4073);
nor NOR4 (N10341, N10335, N3098, N4125, N1855);
and AND2 (N10342, N10334, N647);
xor XOR2 (N10343, N10340, N4750);
nor NOR2 (N10344, N10339, N3154);
nand NAND4 (N10345, N10324, N2314, N3931, N6917);
buf BUF1 (N10346, N10333);
not NOT1 (N10347, N10345);
nand NAND2 (N10348, N10337, N4445);
and AND4 (N10349, N10323, N5868, N2652, N2133);
buf BUF1 (N10350, N10296);
nor NOR3 (N10351, N10347, N8172, N8785);
nand NAND2 (N10352, N10351, N1935);
nand NAND4 (N10353, N10348, N3864, N9566, N4084);
nand NAND4 (N10354, N10350, N1481, N930, N8354);
buf BUF1 (N10355, N10346);
and AND4 (N10356, N10355, N9781, N5472, N7797);
buf BUF1 (N10357, N10342);
buf BUF1 (N10358, N10343);
or OR4 (N10359, N10344, N1685, N1333, N8836);
not NOT1 (N10360, N10328);
buf BUF1 (N10361, N10349);
not NOT1 (N10362, N10356);
or OR4 (N10363, N10360, N2720, N1958, N4722);
or OR2 (N10364, N10361, N4971);
xor XOR2 (N10365, N10362, N1282);
nor NOR4 (N10366, N10352, N3391, N6805, N8669);
nand NAND2 (N10367, N10365, N3293);
not NOT1 (N10368, N10359);
nor NOR3 (N10369, N10341, N4703, N225);
nor NOR3 (N10370, N10357, N1967, N2194);
buf BUF1 (N10371, N10354);
nor NOR4 (N10372, N10367, N5749, N6012, N3121);
or OR2 (N10373, N10369, N28);
xor XOR2 (N10374, N10370, N10153);
nand NAND4 (N10375, N10374, N5348, N856, N3544);
buf BUF1 (N10376, N10371);
nor NOR3 (N10377, N10372, N4311, N6563);
or OR4 (N10378, N10363, N3960, N7760, N1768);
nor NOR2 (N10379, N10377, N6991);
and AND4 (N10380, N10353, N5954, N10169, N8279);
xor XOR2 (N10381, N10358, N1565);
nand NAND3 (N10382, N10375, N7187, N6515);
xor XOR2 (N10383, N10368, N3436);
buf BUF1 (N10384, N10373);
nor NOR3 (N10385, N10380, N8430, N7302);
and AND3 (N10386, N10384, N1993, N1523);
nand NAND3 (N10387, N10378, N8622, N1074);
and AND2 (N10388, N10379, N6658);
not NOT1 (N10389, N10385);
not NOT1 (N10390, N10383);
buf BUF1 (N10391, N10366);
nor NOR4 (N10392, N10387, N7217, N6958, N472);
nor NOR3 (N10393, N10381, N9162, N206);
nor NOR3 (N10394, N10388, N927, N3618);
xor XOR2 (N10395, N10394, N8459);
or OR2 (N10396, N10393, N4291);
nand NAND4 (N10397, N10376, N3175, N7710, N2216);
xor XOR2 (N10398, N10364, N5692);
nor NOR2 (N10399, N10396, N6559);
nor NOR2 (N10400, N10382, N4918);
nand NAND3 (N10401, N10397, N5105, N2839);
and AND3 (N10402, N10395, N3851, N2428);
nor NOR3 (N10403, N10391, N1420, N8990);
buf BUF1 (N10404, N10398);
not NOT1 (N10405, N10400);
and AND4 (N10406, N10402, N8745, N1661, N3843);
nor NOR3 (N10407, N10392, N6328, N3358);
xor XOR2 (N10408, N10406, N4217);
xor XOR2 (N10409, N10390, N903);
xor XOR2 (N10410, N10399, N1934);
not NOT1 (N10411, N10403);
xor XOR2 (N10412, N10411, N986);
nand NAND3 (N10413, N10409, N10078, N5051);
not NOT1 (N10414, N10407);
or OR2 (N10415, N10401, N7923);
and AND4 (N10416, N10410, N4819, N4341, N3900);
nand NAND3 (N10417, N10386, N8726, N10200);
and AND2 (N10418, N10416, N6519);
buf BUF1 (N10419, N10413);
or OR4 (N10420, N10414, N5126, N6177, N5090);
not NOT1 (N10421, N10419);
or OR2 (N10422, N10389, N418);
xor XOR2 (N10423, N10418, N7753);
and AND3 (N10424, N10408, N9486, N1892);
nand NAND4 (N10425, N10404, N8033, N6856, N8981);
nand NAND4 (N10426, N10425, N3741, N2408, N1017);
or OR4 (N10427, N10422, N6852, N4963, N4126);
xor XOR2 (N10428, N10415, N6335);
nand NAND3 (N10429, N10426, N4050, N7801);
nor NOR4 (N10430, N10429, N9587, N75, N7089);
nand NAND2 (N10431, N10424, N5913);
and AND2 (N10432, N10417, N7476);
nor NOR3 (N10433, N10423, N2335, N6756);
and AND4 (N10434, N10421, N8539, N2253, N494);
and AND2 (N10435, N10405, N7016);
nand NAND4 (N10436, N10427, N9506, N4326, N9329);
xor XOR2 (N10437, N10435, N3890);
not NOT1 (N10438, N10433);
nand NAND4 (N10439, N10434, N5733, N5175, N4555);
nor NOR2 (N10440, N10437, N4409);
nor NOR2 (N10441, N10431, N1717);
xor XOR2 (N10442, N10441, N6180);
or OR3 (N10443, N10430, N1253, N9400);
xor XOR2 (N10444, N10420, N5607);
nor NOR4 (N10445, N10412, N1393, N9597, N6411);
xor XOR2 (N10446, N10438, N4517);
xor XOR2 (N10447, N10445, N32);
xor XOR2 (N10448, N10436, N3842);
nor NOR2 (N10449, N10443, N9755);
xor XOR2 (N10450, N10447, N9804);
xor XOR2 (N10451, N10449, N3396);
or OR4 (N10452, N10442, N2647, N3035, N8294);
or OR3 (N10453, N10448, N583, N1052);
or OR4 (N10454, N10451, N5694, N6953, N1117);
or OR2 (N10455, N10428, N1897);
not NOT1 (N10456, N10432);
and AND3 (N10457, N10450, N7927, N3374);
xor XOR2 (N10458, N10444, N3948);
xor XOR2 (N10459, N10456, N5250);
buf BUF1 (N10460, N10440);
and AND2 (N10461, N10460, N34);
nor NOR4 (N10462, N10461, N493, N10321, N614);
nor NOR3 (N10463, N10457, N2699, N6539);
nor NOR3 (N10464, N10459, N4907, N2584);
and AND4 (N10465, N10458, N7623, N8421, N3167);
xor XOR2 (N10466, N10463, N7299);
not NOT1 (N10467, N10452);
nand NAND4 (N10468, N10455, N3194, N1737, N9100);
not NOT1 (N10469, N10466);
and AND2 (N10470, N10453, N324);
buf BUF1 (N10471, N10465);
nand NAND2 (N10472, N10471, N2786);
and AND3 (N10473, N10469, N9090, N4568);
and AND3 (N10474, N10464, N3543, N9501);
or OR3 (N10475, N10462, N935, N1590);
nand NAND3 (N10476, N10446, N4732, N8756);
nand NAND2 (N10477, N10470, N1116);
xor XOR2 (N10478, N10467, N9605);
and AND4 (N10479, N10472, N8767, N2870, N6254);
buf BUF1 (N10480, N10454);
or OR4 (N10481, N10477, N7173, N10097, N4742);
and AND2 (N10482, N10474, N1230);
or OR2 (N10483, N10480, N6485);
nand NAND2 (N10484, N10439, N1174);
nand NAND2 (N10485, N10478, N2021);
buf BUF1 (N10486, N10484);
not NOT1 (N10487, N10475);
and AND2 (N10488, N10486, N4607);
nor NOR4 (N10489, N10483, N10279, N2622, N6816);
not NOT1 (N10490, N10485);
xor XOR2 (N10491, N10489, N4776);
xor XOR2 (N10492, N10481, N6926);
and AND3 (N10493, N10492, N2587, N3375);
nor NOR4 (N10494, N10468, N1276, N4411, N6868);
nand NAND4 (N10495, N10476, N4011, N7805, N3123);
not NOT1 (N10496, N10495);
xor XOR2 (N10497, N10479, N647);
nand NAND4 (N10498, N10496, N1187, N6513, N8011);
xor XOR2 (N10499, N10482, N5745);
buf BUF1 (N10500, N10497);
and AND4 (N10501, N10473, N6563, N810, N5035);
xor XOR2 (N10502, N10490, N2597);
buf BUF1 (N10503, N10494);
not NOT1 (N10504, N10501);
xor XOR2 (N10505, N10502, N9417);
buf BUF1 (N10506, N10499);
nor NOR2 (N10507, N10500, N4405);
buf BUF1 (N10508, N10491);
not NOT1 (N10509, N10503);
or OR4 (N10510, N10505, N3848, N346, N1799);
xor XOR2 (N10511, N10507, N5098);
or OR4 (N10512, N10488, N5031, N10179, N9843);
nand NAND4 (N10513, N10511, N10262, N6774, N2842);
not NOT1 (N10514, N10504);
nand NAND3 (N10515, N10508, N9384, N2691);
nand NAND4 (N10516, N10506, N8527, N7965, N4956);
buf BUF1 (N10517, N10513);
nor NOR4 (N10518, N10487, N6730, N7524, N4343);
and AND3 (N10519, N10518, N10221, N9598);
buf BUF1 (N10520, N10498);
xor XOR2 (N10521, N10516, N4152);
or OR4 (N10522, N10515, N2929, N3268, N720);
buf BUF1 (N10523, N10521);
or OR2 (N10524, N10517, N10079);
nand NAND2 (N10525, N10493, N3727);
not NOT1 (N10526, N10509);
nor NOR4 (N10527, N10524, N3486, N4255, N7771);
or OR2 (N10528, N10519, N7173);
nand NAND2 (N10529, N10523, N2226);
and AND4 (N10530, N10514, N3708, N4766, N1688);
and AND2 (N10531, N10525, N3999);
and AND4 (N10532, N10527, N7867, N2798, N5854);
nor NOR2 (N10533, N10526, N1441);
nor NOR2 (N10534, N10510, N1490);
nor NOR2 (N10535, N10512, N4760);
xor XOR2 (N10536, N10529, N1258);
and AND2 (N10537, N10522, N2713);
nor NOR4 (N10538, N10534, N694, N2980, N4652);
and AND3 (N10539, N10537, N7929, N8079);
not NOT1 (N10540, N10531);
not NOT1 (N10541, N10530);
and AND3 (N10542, N10535, N9342, N5205);
nand NAND3 (N10543, N10528, N109, N7658);
nand NAND2 (N10544, N10538, N10127);
nor NOR3 (N10545, N10543, N10227, N4117);
buf BUF1 (N10546, N10542);
nand NAND2 (N10547, N10532, N8927);
and AND3 (N10548, N10541, N10445, N3111);
xor XOR2 (N10549, N10548, N846);
buf BUF1 (N10550, N10547);
or OR2 (N10551, N10545, N8498);
buf BUF1 (N10552, N10550);
xor XOR2 (N10553, N10520, N26);
nand NAND3 (N10554, N10533, N9783, N5090);
and AND3 (N10555, N10544, N6804, N9934);
nand NAND3 (N10556, N10552, N4628, N1655);
nand NAND3 (N10557, N10555, N2899, N7714);
xor XOR2 (N10558, N10556, N500);
not NOT1 (N10559, N10553);
nand NAND2 (N10560, N10554, N6546);
nor NOR4 (N10561, N10539, N4459, N6586, N7598);
and AND3 (N10562, N10551, N3701, N32);
not NOT1 (N10563, N10540);
buf BUF1 (N10564, N10559);
xor XOR2 (N10565, N10546, N6207);
or OR4 (N10566, N10561, N7822, N5309, N8927);
xor XOR2 (N10567, N10558, N7097);
nand NAND4 (N10568, N10549, N1939, N2399, N7016);
xor XOR2 (N10569, N10563, N1672);
buf BUF1 (N10570, N10568);
nand NAND3 (N10571, N10562, N104, N7559);
xor XOR2 (N10572, N10567, N5258);
not NOT1 (N10573, N10569);
nor NOR2 (N10574, N10573, N8360);
or OR3 (N10575, N10536, N6508, N5660);
nand NAND2 (N10576, N10566, N7481);
not NOT1 (N10577, N10565);
buf BUF1 (N10578, N10572);
nand NAND2 (N10579, N10557, N4337);
or OR4 (N10580, N10577, N242, N8227, N10230);
buf BUF1 (N10581, N10579);
nand NAND4 (N10582, N10580, N1683, N5229, N7405);
and AND2 (N10583, N10578, N9103);
buf BUF1 (N10584, N10564);
or OR4 (N10585, N10583, N5238, N10034, N10217);
nor NOR4 (N10586, N10585, N7925, N6597, N1193);
nor NOR2 (N10587, N10581, N4929);
nor NOR2 (N10588, N10587, N1720);
and AND4 (N10589, N10588, N4980, N889, N4013);
not NOT1 (N10590, N10575);
xor XOR2 (N10591, N10571, N6850);
nand NAND3 (N10592, N10574, N6598, N2689);
and AND3 (N10593, N10576, N9312, N1108);
xor XOR2 (N10594, N10570, N5664);
xor XOR2 (N10595, N10560, N8037);
xor XOR2 (N10596, N10591, N5291);
nor NOR2 (N10597, N10592, N7140);
nor NOR2 (N10598, N10586, N5722);
nand NAND4 (N10599, N10584, N7203, N6180, N10264);
xor XOR2 (N10600, N10590, N9773);
or OR2 (N10601, N10597, N5409);
nand NAND3 (N10602, N10589, N7458, N7893);
and AND4 (N10603, N10598, N1240, N9100, N6406);
or OR2 (N10604, N10595, N204);
buf BUF1 (N10605, N10604);
buf BUF1 (N10606, N10594);
or OR4 (N10607, N10596, N1592, N984, N3714);
buf BUF1 (N10608, N10602);
nand NAND3 (N10609, N10599, N8684, N3705);
nand NAND4 (N10610, N10605, N3934, N5401, N2011);
xor XOR2 (N10611, N10606, N9881);
not NOT1 (N10612, N10603);
nor NOR2 (N10613, N10610, N505);
not NOT1 (N10614, N10582);
nor NOR2 (N10615, N10593, N7935);
xor XOR2 (N10616, N10613, N7);
buf BUF1 (N10617, N10615);
nor NOR3 (N10618, N10617, N2091, N1377);
buf BUF1 (N10619, N10618);
and AND4 (N10620, N10607, N5327, N4279, N4261);
and AND3 (N10621, N10620, N5410, N1691);
xor XOR2 (N10622, N10619, N3822);
nor NOR2 (N10623, N10609, N2094);
not NOT1 (N10624, N10616);
or OR2 (N10625, N10624, N3273);
xor XOR2 (N10626, N10600, N6656);
or OR3 (N10627, N10601, N652, N4304);
xor XOR2 (N10628, N10625, N9202);
not NOT1 (N10629, N10622);
xor XOR2 (N10630, N10623, N750);
nor NOR2 (N10631, N10630, N8326);
nand NAND2 (N10632, N10614, N9280);
nor NOR4 (N10633, N10627, N7639, N8535, N817);
nand NAND2 (N10634, N10629, N8115);
nand NAND3 (N10635, N10634, N10583, N6249);
not NOT1 (N10636, N10608);
nand NAND4 (N10637, N10611, N6948, N8667, N3187);
not NOT1 (N10638, N10626);
xor XOR2 (N10639, N10633, N9759);
nor NOR4 (N10640, N10628, N4872, N1080, N5148);
and AND2 (N10641, N10639, N3825);
not NOT1 (N10642, N10638);
not NOT1 (N10643, N10636);
nor NOR4 (N10644, N10612, N9562, N2254, N1580);
nand NAND3 (N10645, N10621, N4691, N4316);
nand NAND3 (N10646, N10644, N9895, N1036);
buf BUF1 (N10647, N10646);
xor XOR2 (N10648, N10632, N8911);
nor NOR3 (N10649, N10640, N8004, N9181);
and AND4 (N10650, N10642, N8220, N8795, N5132);
nor NOR3 (N10651, N10635, N4288, N8049);
buf BUF1 (N10652, N10641);
xor XOR2 (N10653, N10649, N10056);
buf BUF1 (N10654, N10637);
nand NAND4 (N10655, N10654, N7644, N6547, N6485);
nand NAND3 (N10656, N10648, N10398, N8837);
nor NOR4 (N10657, N10653, N7920, N7761, N8946);
xor XOR2 (N10658, N10657, N4050);
or OR4 (N10659, N10643, N3978, N9419, N5752);
nand NAND3 (N10660, N10647, N7686, N669);
not NOT1 (N10661, N10660);
nor NOR3 (N10662, N10659, N4571, N5467);
buf BUF1 (N10663, N10645);
not NOT1 (N10664, N10661);
buf BUF1 (N10665, N10663);
and AND2 (N10666, N10658, N3098);
xor XOR2 (N10667, N10631, N10372);
and AND4 (N10668, N10665, N807, N7894, N1770);
not NOT1 (N10669, N10650);
xor XOR2 (N10670, N10667, N7525);
not NOT1 (N10671, N10670);
not NOT1 (N10672, N10662);
buf BUF1 (N10673, N10668);
not NOT1 (N10674, N10672);
xor XOR2 (N10675, N10652, N8952);
nand NAND3 (N10676, N10673, N3, N7252);
nand NAND4 (N10677, N10669, N10616, N671, N8356);
xor XOR2 (N10678, N10655, N10615);
xor XOR2 (N10679, N10656, N2936);
or OR3 (N10680, N10674, N3236, N8199);
and AND2 (N10681, N10675, N5362);
not NOT1 (N10682, N10679);
xor XOR2 (N10683, N10666, N7917);
and AND4 (N10684, N10676, N4518, N393, N10368);
buf BUF1 (N10685, N10671);
nor NOR3 (N10686, N10684, N3889, N5022);
not NOT1 (N10687, N10686);
buf BUF1 (N10688, N10683);
buf BUF1 (N10689, N10685);
xor XOR2 (N10690, N10682, N2115);
nor NOR3 (N10691, N10687, N4289, N7253);
nand NAND4 (N10692, N10681, N4209, N1046, N1292);
nor NOR2 (N10693, N10690, N4005);
nand NAND3 (N10694, N10651, N4337, N117);
buf BUF1 (N10695, N10691);
not NOT1 (N10696, N10689);
not NOT1 (N10697, N10696);
or OR4 (N10698, N10694, N8650, N4022, N5901);
xor XOR2 (N10699, N10697, N8735);
nand NAND2 (N10700, N10692, N6915);
buf BUF1 (N10701, N10700);
xor XOR2 (N10702, N10680, N4719);
nand NAND2 (N10703, N10678, N724);
and AND3 (N10704, N10677, N8538, N3421);
buf BUF1 (N10705, N10702);
and AND3 (N10706, N10698, N8755, N10129);
and AND4 (N10707, N10688, N2406, N7555, N1658);
or OR3 (N10708, N10705, N7333, N1418);
not NOT1 (N10709, N10664);
or OR4 (N10710, N10695, N876, N7184, N1718);
nor NOR3 (N10711, N10706, N5893, N6248);
not NOT1 (N10712, N10701);
or OR4 (N10713, N10712, N422, N9261, N4650);
or OR2 (N10714, N10710, N3618);
nor NOR2 (N10715, N10714, N3123);
nand NAND2 (N10716, N10704, N3349);
or OR2 (N10717, N10713, N7029);
and AND2 (N10718, N10715, N4948);
nor NOR2 (N10719, N10711, N565);
xor XOR2 (N10720, N10709, N8011);
nor NOR3 (N10721, N10699, N7350, N9538);
buf BUF1 (N10722, N10693);
or OR3 (N10723, N10717, N6492, N6730);
xor XOR2 (N10724, N10718, N2087);
xor XOR2 (N10725, N10708, N3764);
buf BUF1 (N10726, N10724);
and AND3 (N10727, N10720, N7694, N1717);
not NOT1 (N10728, N10725);
or OR2 (N10729, N10707, N2125);
nand NAND2 (N10730, N10727, N8183);
nand NAND4 (N10731, N10719, N10276, N9721, N9000);
nand NAND3 (N10732, N10728, N7498, N10264);
nand NAND2 (N10733, N10731, N8501);
and AND4 (N10734, N10733, N7268, N4231, N10529);
nand NAND4 (N10735, N10723, N7077, N6706, N2406);
buf BUF1 (N10736, N10729);
or OR3 (N10737, N10722, N3228, N8389);
and AND4 (N10738, N10721, N8658, N445, N2175);
buf BUF1 (N10739, N10738);
not NOT1 (N10740, N10703);
xor XOR2 (N10741, N10716, N9748);
buf BUF1 (N10742, N10735);
buf BUF1 (N10743, N10739);
and AND4 (N10744, N10740, N7734, N1007, N1797);
and AND2 (N10745, N10737, N5293);
and AND3 (N10746, N10743, N1769, N1315);
not NOT1 (N10747, N10741);
or OR3 (N10748, N10744, N599, N3722);
buf BUF1 (N10749, N10732);
nor NOR4 (N10750, N10742, N9477, N1397, N2853);
buf BUF1 (N10751, N10747);
xor XOR2 (N10752, N10736, N9812);
and AND2 (N10753, N10751, N7493);
xor XOR2 (N10754, N10753, N2684);
xor XOR2 (N10755, N10746, N8494);
nand NAND4 (N10756, N10748, N10121, N3404, N9458);
nor NOR3 (N10757, N10730, N10748, N8874);
and AND3 (N10758, N10757, N4296, N9011);
nor NOR3 (N10759, N10758, N7809, N4897);
xor XOR2 (N10760, N10754, N3298);
buf BUF1 (N10761, N10752);
and AND2 (N10762, N10750, N7168);
nand NAND2 (N10763, N10734, N6329);
nand NAND2 (N10764, N10761, N1147);
xor XOR2 (N10765, N10756, N8086);
not NOT1 (N10766, N10760);
buf BUF1 (N10767, N10762);
nor NOR4 (N10768, N10764, N8346, N6759, N5509);
or OR4 (N10769, N10745, N8544, N358, N10553);
nand NAND4 (N10770, N10767, N10372, N5613, N6299);
xor XOR2 (N10771, N10770, N7057);
nor NOR3 (N10772, N10771, N3363, N10274);
not NOT1 (N10773, N10763);
nor NOR4 (N10774, N10759, N729, N6122, N9956);
not NOT1 (N10775, N10768);
nor NOR4 (N10776, N10775, N1889, N10762, N5673);
or OR2 (N10777, N10766, N1558);
buf BUF1 (N10778, N10776);
or OR3 (N10779, N10755, N7037, N2580);
or OR3 (N10780, N10726, N9188, N9945);
nand NAND4 (N10781, N10765, N3957, N245, N1373);
buf BUF1 (N10782, N10749);
nand NAND3 (N10783, N10769, N1371, N584);
or OR2 (N10784, N10779, N4696);
or OR4 (N10785, N10777, N3675, N7183, N9890);
not NOT1 (N10786, N10785);
not NOT1 (N10787, N10786);
buf BUF1 (N10788, N10783);
buf BUF1 (N10789, N10788);
not NOT1 (N10790, N10780);
and AND3 (N10791, N10782, N15, N9173);
and AND2 (N10792, N10773, N1598);
and AND2 (N10793, N10772, N10269);
and AND2 (N10794, N10784, N369);
nor NOR3 (N10795, N10790, N7723, N10152);
not NOT1 (N10796, N10787);
not NOT1 (N10797, N10792);
and AND3 (N10798, N10774, N7591, N8942);
xor XOR2 (N10799, N10798, N1972);
xor XOR2 (N10800, N10793, N5283);
nor NOR2 (N10801, N10795, N3517);
xor XOR2 (N10802, N10799, N5568);
xor XOR2 (N10803, N10791, N8365);
or OR4 (N10804, N10801, N8668, N8643, N1905);
or OR3 (N10805, N10794, N1913, N7193);
not NOT1 (N10806, N10800);
xor XOR2 (N10807, N10804, N4783);
nor NOR3 (N10808, N10778, N5754, N1860);
or OR4 (N10809, N10802, N6998, N838, N2985);
nand NAND2 (N10810, N10806, N1881);
nand NAND3 (N10811, N10797, N6338, N928);
nand NAND4 (N10812, N10796, N7493, N4333, N398);
nand NAND2 (N10813, N10811, N9257);
and AND2 (N10814, N10809, N10303);
and AND2 (N10815, N10803, N7975);
nand NAND2 (N10816, N10813, N10083);
nor NOR3 (N10817, N10810, N3224, N1510);
nor NOR3 (N10818, N10815, N4298, N2437);
nand NAND2 (N10819, N10789, N8450);
nand NAND2 (N10820, N10816, N5813);
not NOT1 (N10821, N10808);
or OR3 (N10822, N10819, N1037, N8114);
nand NAND4 (N10823, N10805, N4044, N7735, N428);
xor XOR2 (N10824, N10781, N8908);
xor XOR2 (N10825, N10807, N2947);
and AND3 (N10826, N10823, N9044, N9391);
nand NAND4 (N10827, N10826, N10206, N4041, N10240);
not NOT1 (N10828, N10825);
not NOT1 (N10829, N10821);
and AND3 (N10830, N10814, N2032, N6120);
nor NOR3 (N10831, N10827, N926, N7115);
or OR4 (N10832, N10822, N10803, N10209, N10137);
nor NOR2 (N10833, N10832, N2345);
or OR3 (N10834, N10831, N6340, N9458);
xor XOR2 (N10835, N10820, N3841);
not NOT1 (N10836, N10834);
nand NAND4 (N10837, N10836, N1356, N5888, N6145);
or OR4 (N10838, N10812, N6432, N9298, N5043);
nor NOR4 (N10839, N10818, N7954, N1915, N10197);
or OR4 (N10840, N10830, N2305, N6828, N4638);
nand NAND2 (N10841, N10824, N10583);
not NOT1 (N10842, N10833);
buf BUF1 (N10843, N10837);
or OR4 (N10844, N10817, N2339, N6343, N8986);
not NOT1 (N10845, N10828);
xor XOR2 (N10846, N10842, N4441);
and AND3 (N10847, N10840, N10679, N746);
nand NAND4 (N10848, N10846, N10482, N1724, N7824);
nand NAND2 (N10849, N10848, N6790);
and AND2 (N10850, N10843, N7609);
nor NOR4 (N10851, N10849, N7963, N4447, N7920);
xor XOR2 (N10852, N10838, N10137);
not NOT1 (N10853, N10845);
buf BUF1 (N10854, N10829);
nand NAND4 (N10855, N10841, N8815, N1568, N10854);
nand NAND4 (N10856, N6706, N10001, N5005, N1443);
nand NAND2 (N10857, N10855, N3290);
or OR4 (N10858, N10856, N10261, N3841, N7549);
xor XOR2 (N10859, N10853, N5630);
nand NAND3 (N10860, N10850, N187, N7588);
not NOT1 (N10861, N10860);
xor XOR2 (N10862, N10861, N5530);
or OR2 (N10863, N10851, N687);
not NOT1 (N10864, N10857);
or OR3 (N10865, N10859, N6573, N5071);
and AND3 (N10866, N10847, N558, N10477);
or OR4 (N10867, N10852, N1140, N2602, N3343);
buf BUF1 (N10868, N10863);
or OR3 (N10869, N10865, N6470, N1541);
not NOT1 (N10870, N10866);
xor XOR2 (N10871, N10858, N733);
and AND2 (N10872, N10862, N4987);
nand NAND2 (N10873, N10868, N8605);
nand NAND2 (N10874, N10869, N6769);
buf BUF1 (N10875, N10872);
buf BUF1 (N10876, N10867);
not NOT1 (N10877, N10835);
buf BUF1 (N10878, N10871);
and AND3 (N10879, N10877, N5157, N6317);
not NOT1 (N10880, N10864);
xor XOR2 (N10881, N10875, N9523);
not NOT1 (N10882, N10870);
nor NOR4 (N10883, N10882, N7685, N7232, N6171);
xor XOR2 (N10884, N10881, N1446);
not NOT1 (N10885, N10879);
nor NOR2 (N10886, N10880, N7498);
not NOT1 (N10887, N10873);
and AND2 (N10888, N10886, N9266);
buf BUF1 (N10889, N10883);
xor XOR2 (N10890, N10888, N5045);
buf BUF1 (N10891, N10874);
buf BUF1 (N10892, N10889);
xor XOR2 (N10893, N10890, N7859);
not NOT1 (N10894, N10876);
nand NAND2 (N10895, N10884, N9435);
xor XOR2 (N10896, N10839, N10112);
buf BUF1 (N10897, N10887);
or OR2 (N10898, N10892, N9518);
not NOT1 (N10899, N10893);
or OR4 (N10900, N10885, N1921, N10327, N889);
or OR2 (N10901, N10844, N2901);
xor XOR2 (N10902, N10900, N4247);
or OR2 (N10903, N10902, N8365);
nand NAND4 (N10904, N10899, N4433, N10384, N2047);
or OR4 (N10905, N10904, N8991, N6420, N5087);
and AND2 (N10906, N10891, N8259);
xor XOR2 (N10907, N10901, N4726);
or OR3 (N10908, N10903, N1714, N2384);
nor NOR3 (N10909, N10878, N2258, N8850);
nor NOR3 (N10910, N10895, N9887, N1223);
not NOT1 (N10911, N10909);
xor XOR2 (N10912, N10898, N6172);
nor NOR3 (N10913, N10896, N5744, N7974);
not NOT1 (N10914, N10910);
and AND2 (N10915, N10913, N10071);
buf BUF1 (N10916, N10894);
buf BUF1 (N10917, N10911);
buf BUF1 (N10918, N10906);
nor NOR4 (N10919, N10907, N6350, N3754, N10890);
or OR2 (N10920, N10915, N7805);
and AND3 (N10921, N10920, N8738, N3349);
buf BUF1 (N10922, N10912);
buf BUF1 (N10923, N10914);
or OR3 (N10924, N10897, N3722, N7592);
xor XOR2 (N10925, N10919, N8135);
buf BUF1 (N10926, N10923);
or OR4 (N10927, N10926, N2649, N8165, N2370);
nor NOR2 (N10928, N10905, N10922);
nor NOR3 (N10929, N10193, N3514, N3874);
buf BUF1 (N10930, N10921);
buf BUF1 (N10931, N10916);
xor XOR2 (N10932, N10925, N938);
buf BUF1 (N10933, N10930);
not NOT1 (N10934, N10929);
nand NAND3 (N10935, N10932, N5091, N6802);
not NOT1 (N10936, N10924);
nand NAND3 (N10937, N10928, N2999, N4035);
and AND3 (N10938, N10935, N9127, N2312);
xor XOR2 (N10939, N10927, N4234);
and AND4 (N10940, N10917, N9276, N8154, N7835);
not NOT1 (N10941, N10918);
xor XOR2 (N10942, N10938, N1479);
nor NOR3 (N10943, N10941, N1773, N4488);
xor XOR2 (N10944, N10936, N1155);
not NOT1 (N10945, N10908);
nand NAND3 (N10946, N10934, N756, N4830);
buf BUF1 (N10947, N10939);
or OR2 (N10948, N10945, N6418);
nor NOR4 (N10949, N10943, N9435, N8708, N6901);
nor NOR2 (N10950, N10946, N6987);
nand NAND2 (N10951, N10950, N749);
xor XOR2 (N10952, N10940, N2022);
nand NAND4 (N10953, N10952, N10306, N865, N854);
xor XOR2 (N10954, N10933, N1922);
nor NOR2 (N10955, N10954, N5423);
buf BUF1 (N10956, N10951);
and AND3 (N10957, N10944, N5603, N9061);
nor NOR3 (N10958, N10942, N8873, N7933);
and AND4 (N10959, N10948, N6847, N5089, N9138);
not NOT1 (N10960, N10959);
nor NOR2 (N10961, N10956, N1145);
nor NOR2 (N10962, N10955, N902);
xor XOR2 (N10963, N10953, N8852);
nor NOR2 (N10964, N10949, N5903);
and AND4 (N10965, N10947, N3832, N3299, N1514);
xor XOR2 (N10966, N10965, N5010);
not NOT1 (N10967, N10964);
or OR3 (N10968, N10960, N1258, N3583);
or OR3 (N10969, N10968, N6090, N5006);
or OR2 (N10970, N10966, N7160);
nand NAND4 (N10971, N10969, N1634, N6865, N6506);
xor XOR2 (N10972, N10957, N5969);
buf BUF1 (N10973, N10958);
not NOT1 (N10974, N10931);
or OR2 (N10975, N10967, N813);
not NOT1 (N10976, N10962);
and AND3 (N10977, N10963, N6149, N3575);
nand NAND2 (N10978, N10974, N5047);
or OR3 (N10979, N10970, N8706, N8683);
and AND3 (N10980, N10973, N3713, N3223);
not NOT1 (N10981, N10961);
xor XOR2 (N10982, N10977, N10917);
nand NAND4 (N10983, N10971, N9500, N3590, N5102);
xor XOR2 (N10984, N10983, N3929);
buf BUF1 (N10985, N10972);
xor XOR2 (N10986, N10975, N8220);
nand NAND2 (N10987, N10986, N6062);
nand NAND3 (N10988, N10985, N5652, N9681);
or OR2 (N10989, N10976, N7239);
nand NAND2 (N10990, N10982, N10146);
nand NAND4 (N10991, N10984, N4845, N7858, N8622);
and AND3 (N10992, N10990, N521, N6925);
xor XOR2 (N10993, N10991, N9894);
nand NAND2 (N10994, N10978, N2622);
or OR2 (N10995, N10989, N9578);
nand NAND3 (N10996, N10988, N3585, N8632);
buf BUF1 (N10997, N10980);
xor XOR2 (N10998, N10997, N6137);
nor NOR4 (N10999, N10937, N6202, N5288, N8953);
buf BUF1 (N11000, N10998);
nor NOR3 (N11001, N10994, N9655, N2791);
nor NOR4 (N11002, N10992, N7472, N2707, N282);
not NOT1 (N11003, N11001);
not NOT1 (N11004, N11000);
and AND4 (N11005, N10999, N3691, N2526, N3069);
or OR3 (N11006, N10987, N9843, N2949);
buf BUF1 (N11007, N10979);
nor NOR2 (N11008, N11004, N2109);
nor NOR2 (N11009, N11002, N3080);
nor NOR3 (N11010, N10995, N833, N8947);
not NOT1 (N11011, N11003);
xor XOR2 (N11012, N10993, N1960);
not NOT1 (N11013, N11009);
xor XOR2 (N11014, N11010, N3301);
nor NOR2 (N11015, N10996, N10100);
nand NAND3 (N11016, N11007, N6624, N7749);
buf BUF1 (N11017, N11008);
buf BUF1 (N11018, N11005);
or OR2 (N11019, N11012, N10789);
or OR4 (N11020, N11016, N5903, N8270, N9392);
and AND4 (N11021, N11011, N5098, N7521, N598);
nor NOR4 (N11022, N11018, N8830, N724, N9145);
buf BUF1 (N11023, N11014);
or OR4 (N11024, N11017, N2510, N8909, N5298);
nand NAND3 (N11025, N11015, N10241, N3953);
nor NOR3 (N11026, N11022, N10931, N10722);
and AND3 (N11027, N11006, N7381, N9422);
not NOT1 (N11028, N11025);
not NOT1 (N11029, N11023);
and AND3 (N11030, N10981, N1714, N3439);
and AND4 (N11031, N11019, N6673, N202, N5409);
xor XOR2 (N11032, N11021, N10140);
buf BUF1 (N11033, N11028);
nor NOR4 (N11034, N11013, N8448, N3441, N5909);
and AND3 (N11035, N11034, N2308, N2781);
and AND2 (N11036, N11033, N10730);
not NOT1 (N11037, N11029);
nand NAND4 (N11038, N11036, N8838, N245, N8890);
and AND2 (N11039, N11037, N6085);
buf BUF1 (N11040, N11030);
xor XOR2 (N11041, N11026, N6001);
buf BUF1 (N11042, N11031);
or OR3 (N11043, N11040, N9490, N5184);
and AND3 (N11044, N11027, N613, N2140);
and AND2 (N11045, N11020, N6533);
xor XOR2 (N11046, N11032, N10814);
not NOT1 (N11047, N11039);
nor NOR2 (N11048, N11044, N1649);
nand NAND3 (N11049, N11046, N10268, N1637);
xor XOR2 (N11050, N11024, N2912);
and AND4 (N11051, N11041, N1928, N9887, N8671);
not NOT1 (N11052, N11043);
not NOT1 (N11053, N11038);
nand NAND2 (N11054, N11052, N2511);
not NOT1 (N11055, N11047);
or OR2 (N11056, N11042, N9439);
xor XOR2 (N11057, N11054, N4794);
and AND2 (N11058, N11056, N5438);
and AND3 (N11059, N11058, N3480, N9760);
not NOT1 (N11060, N11057);
buf BUF1 (N11061, N11049);
and AND4 (N11062, N11053, N7825, N6743, N8960);
buf BUF1 (N11063, N11062);
nor NOR2 (N11064, N11050, N7424);
nand NAND3 (N11065, N11045, N5368, N925);
and AND3 (N11066, N11051, N6445, N136);
nand NAND3 (N11067, N11064, N557, N1935);
and AND2 (N11068, N11059, N10655);
nand NAND2 (N11069, N11061, N1448);
nor NOR3 (N11070, N11060, N1331, N3229);
nand NAND2 (N11071, N11063, N7859);
or OR4 (N11072, N11067, N9274, N3904, N4119);
nor NOR2 (N11073, N11035, N5859);
buf BUF1 (N11074, N11071);
buf BUF1 (N11075, N11068);
and AND4 (N11076, N11070, N6864, N10978, N5940);
or OR2 (N11077, N11055, N9317);
buf BUF1 (N11078, N11066);
xor XOR2 (N11079, N11078, N7184);
xor XOR2 (N11080, N11069, N3362);
or OR2 (N11081, N11075, N1571);
nand NAND3 (N11082, N11076, N2152, N6647);
or OR4 (N11083, N11080, N5432, N8463, N2053);
xor XOR2 (N11084, N11081, N10209);
xor XOR2 (N11085, N11065, N9206);
and AND2 (N11086, N11048, N6471);
xor XOR2 (N11087, N11074, N10098);
buf BUF1 (N11088, N11084);
xor XOR2 (N11089, N11082, N8691);
buf BUF1 (N11090, N11079);
nand NAND2 (N11091, N11089, N9628);
nand NAND4 (N11092, N11086, N7004, N6342, N9557);
or OR4 (N11093, N11083, N6442, N7277, N7752);
xor XOR2 (N11094, N11085, N8535);
nor NOR4 (N11095, N11088, N1766, N10202, N448);
nor NOR4 (N11096, N11077, N4115, N1879, N6590);
and AND2 (N11097, N11096, N633);
buf BUF1 (N11098, N11090);
and AND4 (N11099, N11092, N4978, N1124, N10608);
nand NAND4 (N11100, N11072, N8747, N1667, N8726);
not NOT1 (N11101, N11099);
nand NAND2 (N11102, N11091, N10300);
not NOT1 (N11103, N11102);
nand NAND2 (N11104, N11098, N7529);
nand NAND2 (N11105, N11097, N10404);
nand NAND2 (N11106, N11087, N1658);
and AND4 (N11107, N11093, N1354, N5869, N3284);
and AND3 (N11108, N11105, N1748, N1573);
xor XOR2 (N11109, N11095, N2423);
xor XOR2 (N11110, N11101, N5478);
nand NAND4 (N11111, N11104, N8939, N8181, N7445);
and AND4 (N11112, N11106, N2101, N2636, N9012);
and AND3 (N11113, N11112, N9343, N6151);
or OR3 (N11114, N11103, N5064, N9019);
and AND4 (N11115, N11100, N2859, N783, N9775);
not NOT1 (N11116, N11114);
xor XOR2 (N11117, N11108, N4215);
xor XOR2 (N11118, N11107, N7827);
not NOT1 (N11119, N11116);
not NOT1 (N11120, N11113);
nor NOR2 (N11121, N11073, N749);
buf BUF1 (N11122, N11110);
nor NOR2 (N11123, N11094, N2564);
nand NAND2 (N11124, N11121, N10116);
buf BUF1 (N11125, N11117);
not NOT1 (N11126, N11111);
buf BUF1 (N11127, N11123);
nand NAND4 (N11128, N11120, N8592, N2451, N3793);
and AND3 (N11129, N11125, N10281, N10869);
or OR3 (N11130, N11128, N2462, N4021);
nor NOR2 (N11131, N11129, N10325);
and AND4 (N11132, N11118, N6789, N712, N3221);
nand NAND2 (N11133, N11119, N7228);
and AND4 (N11134, N11127, N2023, N3534, N4086);
buf BUF1 (N11135, N11132);
not NOT1 (N11136, N11122);
xor XOR2 (N11137, N11136, N3391);
nor NOR3 (N11138, N11109, N8612, N7335);
and AND2 (N11139, N11124, N7248);
buf BUF1 (N11140, N11134);
nand NAND2 (N11141, N11139, N11056);
nor NOR2 (N11142, N11135, N8600);
or OR3 (N11143, N11142, N9408, N5154);
and AND2 (N11144, N11140, N7657);
not NOT1 (N11145, N11141);
or OR4 (N11146, N11143, N2284, N9044, N719);
xor XOR2 (N11147, N11146, N7023);
and AND3 (N11148, N11130, N10944, N9806);
or OR3 (N11149, N11138, N10196, N2184);
xor XOR2 (N11150, N11148, N956);
nand NAND2 (N11151, N11137, N5989);
xor XOR2 (N11152, N11145, N9782);
nor NOR4 (N11153, N11151, N3489, N9884, N7615);
and AND2 (N11154, N11153, N7759);
or OR3 (N11155, N11154, N39, N1452);
xor XOR2 (N11156, N11155, N2392);
nand NAND2 (N11157, N11147, N10800);
xor XOR2 (N11158, N11156, N10470);
nor NOR3 (N11159, N11157, N2343, N10579);
nand NAND3 (N11160, N11131, N9238, N214);
buf BUF1 (N11161, N11158);
not NOT1 (N11162, N11159);
nand NAND4 (N11163, N11133, N4476, N3856, N7443);
xor XOR2 (N11164, N11144, N6992);
nor NOR4 (N11165, N11115, N4402, N10258, N7305);
and AND3 (N11166, N11149, N4059, N3308);
nor NOR4 (N11167, N11160, N653, N9865, N2063);
xor XOR2 (N11168, N11161, N1774);
or OR3 (N11169, N11166, N5222, N5596);
buf BUF1 (N11170, N11152);
nor NOR3 (N11171, N11165, N8035, N3557);
buf BUF1 (N11172, N11167);
nand NAND3 (N11173, N11172, N5531, N5261);
or OR3 (N11174, N11126, N9534, N1748);
nand NAND2 (N11175, N11170, N6593);
not NOT1 (N11176, N11173);
or OR2 (N11177, N11168, N4015);
and AND2 (N11178, N11171, N6241);
not NOT1 (N11179, N11174);
nand NAND4 (N11180, N11163, N2405, N1112, N567);
xor XOR2 (N11181, N11175, N10337);
and AND2 (N11182, N11169, N1928);
not NOT1 (N11183, N11181);
not NOT1 (N11184, N11182);
xor XOR2 (N11185, N11178, N6372);
buf BUF1 (N11186, N11183);
xor XOR2 (N11187, N11184, N9494);
nand NAND3 (N11188, N11179, N4574, N1576);
not NOT1 (N11189, N11186);
nor NOR3 (N11190, N11189, N6044, N2072);
not NOT1 (N11191, N11188);
nor NOR4 (N11192, N11176, N8016, N7703, N7787);
nand NAND3 (N11193, N11187, N2338, N6866);
or OR3 (N11194, N11190, N743, N2723);
nand NAND2 (N11195, N11177, N1826);
nor NOR3 (N11196, N11150, N3374, N835);
buf BUF1 (N11197, N11162);
or OR3 (N11198, N11194, N5317, N1418);
buf BUF1 (N11199, N11185);
buf BUF1 (N11200, N11180);
not NOT1 (N11201, N11199);
nor NOR2 (N11202, N11200, N9979);
and AND3 (N11203, N11201, N6991, N7228);
not NOT1 (N11204, N11193);
not NOT1 (N11205, N11192);
or OR3 (N11206, N11196, N6478, N1811);
or OR4 (N11207, N11164, N2507, N656, N7694);
nor NOR4 (N11208, N11205, N7583, N4070, N6409);
or OR3 (N11209, N11197, N7549, N1876);
buf BUF1 (N11210, N11207);
nand NAND4 (N11211, N11191, N7072, N9100, N500);
nor NOR4 (N11212, N11195, N10873, N3491, N3240);
and AND4 (N11213, N11208, N10811, N1134, N11201);
nor NOR4 (N11214, N11202, N7545, N9006, N636);
not NOT1 (N11215, N11213);
or OR3 (N11216, N11214, N10632, N494);
nor NOR4 (N11217, N11198, N7038, N2549, N10102);
nand NAND4 (N11218, N11211, N9800, N332, N3387);
or OR4 (N11219, N11203, N4091, N10245, N4658);
nor NOR2 (N11220, N11204, N6703);
or OR4 (N11221, N11215, N9665, N5860, N8590);
nor NOR2 (N11222, N11212, N10776);
and AND2 (N11223, N11210, N8744);
or OR3 (N11224, N11209, N8047, N3952);
and AND4 (N11225, N11216, N9573, N3075, N8806);
nor NOR4 (N11226, N11206, N4857, N6215, N10009);
nor NOR3 (N11227, N11219, N2774, N2379);
buf BUF1 (N11228, N11226);
not NOT1 (N11229, N11228);
or OR2 (N11230, N11223, N1651);
nand NAND2 (N11231, N11225, N6962);
and AND3 (N11232, N11231, N5105, N4785);
and AND4 (N11233, N11227, N3662, N6964, N6877);
nand NAND2 (N11234, N11229, N1584);
buf BUF1 (N11235, N11224);
nor NOR2 (N11236, N11233, N4574);
not NOT1 (N11237, N11236);
nand NAND4 (N11238, N11232, N6390, N2995, N6666);
buf BUF1 (N11239, N11235);
nand NAND2 (N11240, N11218, N1310);
xor XOR2 (N11241, N11221, N923);
or OR4 (N11242, N11230, N8456, N7539, N8054);
or OR2 (N11243, N11238, N6218);
or OR2 (N11244, N11234, N10673);
nand NAND3 (N11245, N11243, N10828, N4318);
buf BUF1 (N11246, N11220);
xor XOR2 (N11247, N11217, N1509);
nand NAND3 (N11248, N11246, N625, N8821);
not NOT1 (N11249, N11244);
xor XOR2 (N11250, N11241, N2548);
buf BUF1 (N11251, N11239);
not NOT1 (N11252, N11242);
nor NOR4 (N11253, N11247, N8828, N7738, N7491);
or OR3 (N11254, N11222, N10103, N939);
nand NAND4 (N11255, N11250, N6466, N9001, N540);
and AND3 (N11256, N11249, N5371, N6358);
nand NAND4 (N11257, N11256, N4076, N5935, N7676);
nor NOR2 (N11258, N11245, N8687);
nor NOR2 (N11259, N11251, N156);
and AND2 (N11260, N11240, N7572);
xor XOR2 (N11261, N11255, N6021);
buf BUF1 (N11262, N11257);
nand NAND3 (N11263, N11253, N7338, N7995);
nand NAND3 (N11264, N11252, N1667, N4532);
buf BUF1 (N11265, N11259);
nand NAND2 (N11266, N11260, N9412);
xor XOR2 (N11267, N11263, N4856);
or OR3 (N11268, N11262, N1474, N1460);
and AND3 (N11269, N11266, N9181, N4957);
not NOT1 (N11270, N11258);
not NOT1 (N11271, N11269);
xor XOR2 (N11272, N11270, N1826);
or OR3 (N11273, N11272, N5069, N7835);
buf BUF1 (N11274, N11261);
buf BUF1 (N11275, N11254);
not NOT1 (N11276, N11267);
not NOT1 (N11277, N11265);
and AND2 (N11278, N11275, N9022);
buf BUF1 (N11279, N11268);
nand NAND4 (N11280, N11237, N8060, N9217, N8103);
nor NOR4 (N11281, N11248, N10838, N9468, N1490);
buf BUF1 (N11282, N11276);
buf BUF1 (N11283, N11280);
not NOT1 (N11284, N11271);
nand NAND3 (N11285, N11281, N1097, N341);
not NOT1 (N11286, N11273);
buf BUF1 (N11287, N11286);
nand NAND2 (N11288, N11278, N942);
and AND4 (N11289, N11288, N8830, N6463, N7495);
and AND2 (N11290, N11277, N10758);
nand NAND3 (N11291, N11285, N5370, N7497);
nand NAND2 (N11292, N11289, N5394);
buf BUF1 (N11293, N11292);
not NOT1 (N11294, N11282);
xor XOR2 (N11295, N11293, N9979);
nor NOR2 (N11296, N11283, N10192);
xor XOR2 (N11297, N11290, N825);
or OR4 (N11298, N11284, N1460, N4933, N10340);
and AND3 (N11299, N11291, N5595, N5357);
or OR2 (N11300, N11296, N3936);
and AND3 (N11301, N11299, N2436, N9951);
xor XOR2 (N11302, N11264, N8548);
nor NOR4 (N11303, N11279, N8646, N10450, N4196);
buf BUF1 (N11304, N11298);
nand NAND2 (N11305, N11297, N4365);
buf BUF1 (N11306, N11302);
and AND3 (N11307, N11294, N5832, N9301);
nand NAND4 (N11308, N11303, N4543, N2767, N7063);
not NOT1 (N11309, N11287);
nor NOR2 (N11310, N11309, N2209);
xor XOR2 (N11311, N11304, N3269);
nand NAND4 (N11312, N11306, N887, N9795, N5669);
nor NOR2 (N11313, N11311, N3616);
nor NOR2 (N11314, N11301, N2471);
nand NAND3 (N11315, N11313, N454, N728);
xor XOR2 (N11316, N11308, N7486);
nand NAND4 (N11317, N11316, N2159, N4430, N4425);
and AND4 (N11318, N11315, N6500, N83, N1411);
and AND2 (N11319, N11274, N4164);
not NOT1 (N11320, N11319);
nor NOR2 (N11321, N11312, N5667);
not NOT1 (N11322, N11314);
buf BUF1 (N11323, N11322);
xor XOR2 (N11324, N11317, N10357);
buf BUF1 (N11325, N11318);
xor XOR2 (N11326, N11305, N4238);
buf BUF1 (N11327, N11300);
buf BUF1 (N11328, N11307);
not NOT1 (N11329, N11326);
and AND4 (N11330, N11321, N5126, N8397, N4395);
xor XOR2 (N11331, N11327, N687);
not NOT1 (N11332, N11329);
xor XOR2 (N11333, N11324, N3751);
not NOT1 (N11334, N11328);
buf BUF1 (N11335, N11295);
not NOT1 (N11336, N11330);
buf BUF1 (N11337, N11320);
and AND4 (N11338, N11336, N3189, N3668, N7727);
not NOT1 (N11339, N11333);
nor NOR3 (N11340, N11339, N10456, N3744);
nand NAND2 (N11341, N11310, N10528);
not NOT1 (N11342, N11340);
nor NOR4 (N11343, N11341, N6042, N46, N5174);
not NOT1 (N11344, N11343);
and AND2 (N11345, N11338, N7255);
not NOT1 (N11346, N11331);
or OR4 (N11347, N11325, N11173, N2915, N5296);
xor XOR2 (N11348, N11337, N8582);
or OR2 (N11349, N11342, N6330);
or OR3 (N11350, N11334, N794, N2691);
nor NOR2 (N11351, N11350, N1103);
nand NAND2 (N11352, N11335, N5361);
or OR3 (N11353, N11344, N4453, N1913);
and AND2 (N11354, N11352, N3836);
buf BUF1 (N11355, N11354);
and AND2 (N11356, N11345, N1452);
not NOT1 (N11357, N11323);
buf BUF1 (N11358, N11346);
and AND3 (N11359, N11332, N2672, N9315);
nand NAND4 (N11360, N11355, N1985, N4951, N3030);
or OR4 (N11361, N11353, N6011, N3589, N533);
buf BUF1 (N11362, N11347);
or OR4 (N11363, N11362, N5343, N8324, N6530);
and AND3 (N11364, N11349, N3383, N4);
or OR2 (N11365, N11364, N2020);
nand NAND4 (N11366, N11365, N6240, N10932, N5290);
or OR2 (N11367, N11356, N4734);
not NOT1 (N11368, N11359);
buf BUF1 (N11369, N11348);
and AND2 (N11370, N11363, N6456);
xor XOR2 (N11371, N11370, N2108);
buf BUF1 (N11372, N11369);
nand NAND3 (N11373, N11366, N5430, N838);
and AND3 (N11374, N11358, N2873, N9778);
or OR3 (N11375, N11357, N8713, N10766);
xor XOR2 (N11376, N11372, N2141);
or OR4 (N11377, N11376, N1641, N535, N11122);
or OR4 (N11378, N11360, N8683, N3345, N6470);
and AND4 (N11379, N11377, N6082, N7484, N4790);
and AND3 (N11380, N11371, N6008, N4887);
and AND3 (N11381, N11379, N335, N311);
not NOT1 (N11382, N11381);
buf BUF1 (N11383, N11382);
and AND2 (N11384, N11380, N8941);
not NOT1 (N11385, N11384);
buf BUF1 (N11386, N11385);
nand NAND3 (N11387, N11378, N5816, N627);
buf BUF1 (N11388, N11375);
and AND4 (N11389, N11374, N7539, N6672, N6664);
not NOT1 (N11390, N11389);
not NOT1 (N11391, N11387);
and AND4 (N11392, N11390, N142, N5525, N9107);
xor XOR2 (N11393, N11351, N9087);
and AND3 (N11394, N11391, N169, N7382);
not NOT1 (N11395, N11388);
or OR3 (N11396, N11373, N2678, N6633);
and AND2 (N11397, N11395, N11251);
nor NOR4 (N11398, N11396, N1052, N8184, N3939);
buf BUF1 (N11399, N11393);
and AND3 (N11400, N11383, N2737, N7160);
nor NOR2 (N11401, N11398, N10770);
xor XOR2 (N11402, N11367, N1610);
nand NAND3 (N11403, N11394, N9102, N11092);
buf BUF1 (N11404, N11402);
nand NAND3 (N11405, N11400, N8813, N4608);
buf BUF1 (N11406, N11405);
not NOT1 (N11407, N11406);
nor NOR3 (N11408, N11404, N395, N3678);
or OR2 (N11409, N11399, N1462);
nor NOR2 (N11410, N11386, N7423);
xor XOR2 (N11411, N11392, N7652);
and AND3 (N11412, N11408, N4578, N6372);
nor NOR4 (N11413, N11411, N3551, N5760, N4954);
or OR2 (N11414, N11397, N2846);
and AND3 (N11415, N11409, N6123, N3350);
not NOT1 (N11416, N11412);
not NOT1 (N11417, N11413);
not NOT1 (N11418, N11361);
buf BUF1 (N11419, N11368);
and AND4 (N11420, N11416, N6389, N6742, N5669);
nand NAND2 (N11421, N11420, N11343);
and AND4 (N11422, N11414, N6193, N6682, N1693);
nand NAND2 (N11423, N11422, N4511);
or OR4 (N11424, N11423, N4066, N8619, N6790);
xor XOR2 (N11425, N11424, N2044);
and AND4 (N11426, N11425, N1037, N8799, N11186);
nor NOR3 (N11427, N11410, N9048, N8836);
nor NOR2 (N11428, N11403, N2978);
or OR3 (N11429, N11426, N3500, N9239);
and AND2 (N11430, N11428, N2854);
and AND4 (N11431, N11407, N5178, N1290, N8898);
buf BUF1 (N11432, N11419);
nor NOR3 (N11433, N11430, N5338, N10844);
buf BUF1 (N11434, N11429);
nand NAND3 (N11435, N11433, N6337, N11065);
or OR4 (N11436, N11431, N1596, N1201, N7235);
nand NAND3 (N11437, N11417, N9071, N1354);
not NOT1 (N11438, N11401);
nor NOR3 (N11439, N11434, N1818, N10094);
or OR4 (N11440, N11432, N2898, N3282, N7046);
xor XOR2 (N11441, N11415, N7830);
and AND4 (N11442, N11439, N9629, N2363, N2509);
xor XOR2 (N11443, N11437, N4654);
and AND4 (N11444, N11441, N5441, N887, N3921);
not NOT1 (N11445, N11442);
and AND2 (N11446, N11440, N1383);
nand NAND3 (N11447, N11436, N9665, N7506);
or OR3 (N11448, N11444, N5147, N2600);
xor XOR2 (N11449, N11445, N4321);
and AND4 (N11450, N11447, N9952, N1709, N1248);
buf BUF1 (N11451, N11418);
buf BUF1 (N11452, N11427);
and AND2 (N11453, N11450, N10882);
nand NAND4 (N11454, N11443, N8942, N10671, N1236);
or OR4 (N11455, N11438, N1457, N5579, N4966);
not NOT1 (N11456, N11435);
nand NAND4 (N11457, N11456, N5429, N6629, N9129);
nor NOR3 (N11458, N11451, N6491, N5357);
xor XOR2 (N11459, N11453, N9778);
buf BUF1 (N11460, N11449);
and AND4 (N11461, N11454, N5216, N3520, N4161);
buf BUF1 (N11462, N11446);
nand NAND3 (N11463, N11461, N826, N8251);
not NOT1 (N11464, N11448);
nand NAND4 (N11465, N11462, N9687, N5417, N9794);
buf BUF1 (N11466, N11452);
buf BUF1 (N11467, N11466);
xor XOR2 (N11468, N11457, N7541);
nand NAND4 (N11469, N11465, N896, N10275, N2270);
or OR4 (N11470, N11421, N7035, N1533, N3736);
nand NAND4 (N11471, N11458, N775, N6717, N8531);
nor NOR3 (N11472, N11469, N4671, N4684);
or OR2 (N11473, N11468, N8783);
and AND3 (N11474, N11473, N5138, N2823);
buf BUF1 (N11475, N11455);
or OR4 (N11476, N11475, N9491, N4820, N11030);
not NOT1 (N11477, N11464);
nand NAND4 (N11478, N11476, N10006, N10464, N9051);
and AND2 (N11479, N11477, N9969);
nand NAND4 (N11480, N11463, N5, N2009, N9655);
xor XOR2 (N11481, N11472, N8920);
not NOT1 (N11482, N11479);
and AND3 (N11483, N11481, N2885, N6695);
not NOT1 (N11484, N11471);
nor NOR4 (N11485, N11478, N3941, N8262, N2393);
nand NAND4 (N11486, N11460, N2183, N9179, N11360);
and AND2 (N11487, N11467, N5900);
or OR2 (N11488, N11484, N3243);
buf BUF1 (N11489, N11486);
nand NAND4 (N11490, N11474, N7963, N7132, N7334);
nor NOR3 (N11491, N11480, N6322, N2685);
and AND2 (N11492, N11489, N2328);
nand NAND3 (N11493, N11487, N7937, N4573);
buf BUF1 (N11494, N11492);
not NOT1 (N11495, N11485);
and AND3 (N11496, N11459, N586, N11080);
nor NOR2 (N11497, N11493, N11064);
and AND4 (N11498, N11490, N6987, N4391, N1132);
nand NAND3 (N11499, N11498, N5895, N3346);
not NOT1 (N11500, N11488);
xor XOR2 (N11501, N11494, N5240);
xor XOR2 (N11502, N11491, N1624);
xor XOR2 (N11503, N11483, N7472);
not NOT1 (N11504, N11503);
and AND3 (N11505, N11497, N1191, N6042);
nand NAND3 (N11506, N11504, N9217, N1748);
nand NAND2 (N11507, N11500, N15);
xor XOR2 (N11508, N11501, N3815);
or OR2 (N11509, N11506, N777);
nand NAND4 (N11510, N11499, N11284, N4797, N6733);
xor XOR2 (N11511, N11507, N7161);
and AND2 (N11512, N11510, N9720);
nor NOR2 (N11513, N11495, N798);
not NOT1 (N11514, N11505);
nor NOR2 (N11515, N11511, N3963);
or OR3 (N11516, N11496, N2386, N10768);
not NOT1 (N11517, N11513);
and AND4 (N11518, N11512, N1197, N2707, N8956);
or OR3 (N11519, N11514, N9739, N8916);
nor NOR4 (N11520, N11517, N3207, N9861, N7812);
or OR4 (N11521, N11509, N7125, N646, N6663);
xor XOR2 (N11522, N11516, N7558);
buf BUF1 (N11523, N11521);
nand NAND3 (N11524, N11522, N2398, N7183);
not NOT1 (N11525, N11524);
buf BUF1 (N11526, N11518);
xor XOR2 (N11527, N11515, N4213);
nand NAND2 (N11528, N11519, N7790);
and AND2 (N11529, N11520, N11014);
xor XOR2 (N11530, N11525, N5890);
buf BUF1 (N11531, N11502);
or OR4 (N11532, N11523, N4140, N601, N10575);
nand NAND4 (N11533, N11482, N9029, N1089, N8984);
not NOT1 (N11534, N11526);
nor NOR4 (N11535, N11533, N10197, N8737, N11132);
or OR3 (N11536, N11532, N4692, N6288);
not NOT1 (N11537, N11536);
not NOT1 (N11538, N11534);
buf BUF1 (N11539, N11527);
or OR3 (N11540, N11470, N1567, N6490);
nand NAND3 (N11541, N11531, N4141, N9860);
xor XOR2 (N11542, N11528, N2630);
nand NAND2 (N11543, N11540, N10170);
not NOT1 (N11544, N11508);
buf BUF1 (N11545, N11544);
or OR3 (N11546, N11530, N2747, N1459);
not NOT1 (N11547, N11539);
or OR2 (N11548, N11538, N5958);
nand NAND4 (N11549, N11541, N5121, N4279, N6187);
xor XOR2 (N11550, N11535, N89);
xor XOR2 (N11551, N11543, N4703);
or OR4 (N11552, N11529, N10841, N2530, N7619);
buf BUF1 (N11553, N11542);
xor XOR2 (N11554, N11551, N255);
or OR3 (N11555, N11553, N529, N10510);
not NOT1 (N11556, N11547);
buf BUF1 (N11557, N11548);
and AND4 (N11558, N11545, N7078, N3359, N1139);
or OR3 (N11559, N11550, N1809, N6923);
and AND2 (N11560, N11559, N6720);
nand NAND3 (N11561, N11552, N9807, N8622);
or OR4 (N11562, N11560, N9230, N10164, N1443);
not NOT1 (N11563, N11549);
buf BUF1 (N11564, N11563);
or OR2 (N11565, N11554, N6244);
nand NAND4 (N11566, N11546, N9411, N4467, N789);
not NOT1 (N11567, N11537);
not NOT1 (N11568, N11566);
or OR3 (N11569, N11561, N11180, N3087);
and AND3 (N11570, N11562, N4416, N976);
nor NOR2 (N11571, N11568, N8612);
nand NAND4 (N11572, N11569, N11412, N6344, N5301);
xor XOR2 (N11573, N11570, N3202);
or OR2 (N11574, N11558, N5406);
nand NAND4 (N11575, N11574, N8271, N8720, N9947);
nand NAND4 (N11576, N11555, N9689, N3823, N2996);
nor NOR4 (N11577, N11572, N2757, N11265, N6142);
nor NOR2 (N11578, N11557, N749);
nor NOR2 (N11579, N11573, N7973);
buf BUF1 (N11580, N11556);
nor NOR2 (N11581, N11571, N8943);
buf BUF1 (N11582, N11567);
and AND2 (N11583, N11580, N339);
buf BUF1 (N11584, N11578);
and AND4 (N11585, N11582, N217, N3984, N151);
nand NAND4 (N11586, N11575, N4198, N3070, N4378);
buf BUF1 (N11587, N11583);
or OR2 (N11588, N11584, N1823);
xor XOR2 (N11589, N11588, N7155);
or OR4 (N11590, N11564, N4198, N8597, N6350);
or OR4 (N11591, N11587, N2930, N713, N10726);
nor NOR2 (N11592, N11577, N2172);
and AND4 (N11593, N11579, N9419, N11578, N5408);
not NOT1 (N11594, N11576);
or OR3 (N11595, N11593, N2866, N6727);
and AND4 (N11596, N11581, N2834, N5408, N7429);
nor NOR3 (N11597, N11596, N3292, N905);
buf BUF1 (N11598, N11591);
nand NAND3 (N11599, N11597, N4446, N7334);
and AND3 (N11600, N11592, N10878, N9795);
or OR4 (N11601, N11600, N4635, N1732, N4836);
and AND4 (N11602, N11599, N3052, N801, N4947);
xor XOR2 (N11603, N11589, N19);
or OR2 (N11604, N11565, N10992);
xor XOR2 (N11605, N11595, N1895);
buf BUF1 (N11606, N11585);
or OR3 (N11607, N11606, N2722, N3512);
buf BUF1 (N11608, N11598);
xor XOR2 (N11609, N11608, N1103);
nor NOR2 (N11610, N11586, N5892);
buf BUF1 (N11611, N11607);
not NOT1 (N11612, N11601);
or OR3 (N11613, N11603, N9025, N6850);
nor NOR2 (N11614, N11611, N7848);
xor XOR2 (N11615, N11613, N1222);
buf BUF1 (N11616, N11615);
xor XOR2 (N11617, N11610, N2015);
xor XOR2 (N11618, N11604, N6389);
not NOT1 (N11619, N11612);
xor XOR2 (N11620, N11590, N6313);
or OR4 (N11621, N11617, N3861, N876, N10526);
or OR4 (N11622, N11602, N2421, N2044, N10903);
xor XOR2 (N11623, N11622, N5082);
xor XOR2 (N11624, N11620, N4476);
xor XOR2 (N11625, N11594, N306);
buf BUF1 (N11626, N11605);
or OR2 (N11627, N11618, N6594);
buf BUF1 (N11628, N11609);
not NOT1 (N11629, N11625);
and AND4 (N11630, N11616, N6967, N4324, N3562);
or OR3 (N11631, N11628, N1198, N976);
buf BUF1 (N11632, N11624);
buf BUF1 (N11633, N11632);
buf BUF1 (N11634, N11633);
not NOT1 (N11635, N11627);
nand NAND3 (N11636, N11619, N3802, N6766);
xor XOR2 (N11637, N11614, N5590);
nor NOR2 (N11638, N11634, N6982);
not NOT1 (N11639, N11621);
not NOT1 (N11640, N11637);
buf BUF1 (N11641, N11640);
xor XOR2 (N11642, N11635, N7785);
and AND3 (N11643, N11631, N5504, N201);
not NOT1 (N11644, N11626);
xor XOR2 (N11645, N11641, N9514);
xor XOR2 (N11646, N11642, N11092);
or OR2 (N11647, N11629, N10101);
nor NOR3 (N11648, N11647, N7289, N949);
or OR2 (N11649, N11630, N2940);
or OR2 (N11650, N11643, N645);
buf BUF1 (N11651, N11649);
not NOT1 (N11652, N11650);
xor XOR2 (N11653, N11645, N7770);
nor NOR3 (N11654, N11653, N8847, N8437);
buf BUF1 (N11655, N11644);
and AND3 (N11656, N11655, N8007, N2171);
xor XOR2 (N11657, N11651, N2630);
buf BUF1 (N11658, N11623);
xor XOR2 (N11659, N11658, N8425);
and AND3 (N11660, N11636, N5369, N11432);
or OR2 (N11661, N11638, N2140);
nor NOR3 (N11662, N11656, N8246, N6251);
nand NAND4 (N11663, N11660, N2943, N8522, N3331);
xor XOR2 (N11664, N11646, N2960);
not NOT1 (N11665, N11661);
and AND4 (N11666, N11657, N3083, N3946, N9225);
not NOT1 (N11667, N11665);
buf BUF1 (N11668, N11666);
xor XOR2 (N11669, N11648, N5776);
nor NOR2 (N11670, N11659, N2953);
buf BUF1 (N11671, N11639);
or OR3 (N11672, N11664, N1045, N6564);
xor XOR2 (N11673, N11670, N5709);
not NOT1 (N11674, N11663);
or OR2 (N11675, N11667, N952);
nor NOR4 (N11676, N11673, N10075, N3096, N5044);
xor XOR2 (N11677, N11674, N7204);
not NOT1 (N11678, N11677);
nor NOR2 (N11679, N11654, N9571);
nand NAND2 (N11680, N11676, N81);
and AND4 (N11681, N11679, N4662, N10253, N8059);
xor XOR2 (N11682, N11662, N4006);
or OR4 (N11683, N11682, N8379, N7263, N9698);
nor NOR2 (N11684, N11678, N8604);
or OR2 (N11685, N11672, N650);
not NOT1 (N11686, N11683);
and AND2 (N11687, N11684, N8373);
and AND3 (N11688, N11675, N9302, N11440);
xor XOR2 (N11689, N11680, N848);
or OR2 (N11690, N11668, N1734);
xor XOR2 (N11691, N11687, N2684);
nor NOR2 (N11692, N11686, N9088);
or OR4 (N11693, N11685, N6016, N9560, N1304);
nand NAND4 (N11694, N11692, N5165, N2960, N6563);
not NOT1 (N11695, N11669);
nor NOR4 (N11696, N11694, N4114, N949, N11002);
or OR2 (N11697, N11652, N5152);
nand NAND2 (N11698, N11691, N1230);
xor XOR2 (N11699, N11696, N292);
xor XOR2 (N11700, N11697, N5461);
and AND2 (N11701, N11671, N93);
not NOT1 (N11702, N11681);
not NOT1 (N11703, N11701);
nand NAND2 (N11704, N11703, N4921);
not NOT1 (N11705, N11690);
buf BUF1 (N11706, N11698);
or OR4 (N11707, N11705, N7044, N4706, N5712);
xor XOR2 (N11708, N11699, N6522);
buf BUF1 (N11709, N11695);
buf BUF1 (N11710, N11689);
and AND4 (N11711, N11706, N10865, N7820, N4431);
xor XOR2 (N11712, N11708, N9428);
nand NAND4 (N11713, N11712, N2723, N6716, N7305);
and AND3 (N11714, N11713, N6990, N7048);
xor XOR2 (N11715, N11707, N4057);
or OR2 (N11716, N11702, N2115);
not NOT1 (N11717, N11710);
xor XOR2 (N11718, N11704, N7633);
xor XOR2 (N11719, N11718, N9800);
nor NOR2 (N11720, N11711, N7735);
or OR4 (N11721, N11709, N4419, N11613, N8404);
nand NAND3 (N11722, N11715, N4678, N8402);
nor NOR2 (N11723, N11719, N9308);
nand NAND3 (N11724, N11722, N627, N6553);
nor NOR4 (N11725, N11720, N6676, N3798, N5305);
nor NOR2 (N11726, N11700, N7557);
or OR2 (N11727, N11688, N230);
not NOT1 (N11728, N11717);
and AND3 (N11729, N11724, N11497, N5084);
buf BUF1 (N11730, N11721);
nor NOR3 (N11731, N11693, N5779, N4876);
xor XOR2 (N11732, N11727, N9191);
nor NOR2 (N11733, N11723, N10923);
not NOT1 (N11734, N11716);
nand NAND4 (N11735, N11731, N1619, N2227, N6428);
xor XOR2 (N11736, N11728, N6286);
nand NAND4 (N11737, N11735, N2394, N10589, N9215);
nor NOR2 (N11738, N11726, N7593);
not NOT1 (N11739, N11733);
nand NAND2 (N11740, N11730, N449);
xor XOR2 (N11741, N11725, N10010);
nor NOR4 (N11742, N11738, N9460, N2175, N4852);
buf BUF1 (N11743, N11732);
not NOT1 (N11744, N11734);
nor NOR4 (N11745, N11729, N19, N11655, N4814);
or OR3 (N11746, N11737, N260, N1774);
nand NAND3 (N11747, N11745, N11359, N7455);
not NOT1 (N11748, N11746);
and AND4 (N11749, N11743, N11102, N11367, N11644);
buf BUF1 (N11750, N11740);
nor NOR3 (N11751, N11742, N7777, N5888);
or OR4 (N11752, N11747, N5548, N3767, N10675);
nor NOR3 (N11753, N11741, N11204, N5907);
xor XOR2 (N11754, N11739, N10973);
not NOT1 (N11755, N11714);
nand NAND3 (N11756, N11753, N1716, N1785);
and AND2 (N11757, N11752, N9051);
not NOT1 (N11758, N11744);
buf BUF1 (N11759, N11756);
nor NOR4 (N11760, N11758, N9417, N1698, N3576);
not NOT1 (N11761, N11749);
nand NAND4 (N11762, N11757, N9423, N2238, N3686);
or OR3 (N11763, N11755, N3190, N7067);
or OR2 (N11764, N11763, N502);
buf BUF1 (N11765, N11750);
and AND3 (N11766, N11759, N4916, N6693);
not NOT1 (N11767, N11762);
and AND3 (N11768, N11760, N11579, N2978);
nand NAND3 (N11769, N11765, N5986, N4656);
nand NAND3 (N11770, N11748, N2664, N5546);
nor NOR4 (N11771, N11768, N3373, N2045, N9761);
buf BUF1 (N11772, N11770);
not NOT1 (N11773, N11761);
or OR3 (N11774, N11773, N1001, N1786);
or OR2 (N11775, N11769, N815);
or OR3 (N11776, N11751, N7634, N2585);
and AND2 (N11777, N11776, N3826);
and AND3 (N11778, N11772, N688, N1868);
buf BUF1 (N11779, N11774);
nand NAND2 (N11780, N11767, N7517);
xor XOR2 (N11781, N11780, N53);
xor XOR2 (N11782, N11764, N8659);
buf BUF1 (N11783, N11777);
nor NOR3 (N11784, N11775, N7142, N9793);
not NOT1 (N11785, N11783);
or OR3 (N11786, N11784, N4682, N7763);
and AND2 (N11787, N11786, N10759);
xor XOR2 (N11788, N11766, N9268);
buf BUF1 (N11789, N11785);
buf BUF1 (N11790, N11782);
and AND2 (N11791, N11771, N1231);
nor NOR3 (N11792, N11789, N1785, N2757);
xor XOR2 (N11793, N11787, N9397);
buf BUF1 (N11794, N11792);
or OR3 (N11795, N11793, N5389, N9828);
buf BUF1 (N11796, N11791);
nand NAND3 (N11797, N11779, N9531, N11317);
and AND3 (N11798, N11797, N443, N152);
and AND3 (N11799, N11794, N9799, N6780);
buf BUF1 (N11800, N11754);
xor XOR2 (N11801, N11798, N4551);
nor NOR3 (N11802, N11795, N4526, N8917);
nor NOR2 (N11803, N11796, N5892);
buf BUF1 (N11804, N11800);
and AND2 (N11805, N11778, N5617);
not NOT1 (N11806, N11803);
and AND4 (N11807, N11804, N3270, N1540, N3978);
nor NOR4 (N11808, N11736, N1595, N9952, N11430);
and AND2 (N11809, N11799, N3392);
xor XOR2 (N11810, N11788, N4355);
not NOT1 (N11811, N11806);
nand NAND4 (N11812, N11781, N1910, N1710, N635);
nand NAND4 (N11813, N11809, N4387, N7261, N2756);
or OR3 (N11814, N11807, N3282, N6721);
xor XOR2 (N11815, N11808, N7863);
and AND3 (N11816, N11790, N3901, N3888);
xor XOR2 (N11817, N11814, N7273);
nor NOR4 (N11818, N11815, N10277, N4385, N11292);
nand NAND4 (N11819, N11801, N5881, N1157, N10798);
nand NAND3 (N11820, N11816, N1011, N4083);
not NOT1 (N11821, N11805);
not NOT1 (N11822, N11820);
nand NAND3 (N11823, N11819, N221, N5806);
not NOT1 (N11824, N11812);
or OR4 (N11825, N11823, N4691, N573, N2571);
nand NAND3 (N11826, N11802, N10226, N124);
and AND4 (N11827, N11821, N10543, N489, N7981);
not NOT1 (N11828, N11818);
nand NAND2 (N11829, N11810, N5528);
nand NAND4 (N11830, N11829, N10483, N4750, N9616);
nand NAND4 (N11831, N11828, N5486, N2423, N1928);
and AND4 (N11832, N11827, N8225, N1391, N1614);
and AND4 (N11833, N11813, N10833, N10481, N454);
buf BUF1 (N11834, N11831);
or OR2 (N11835, N11834, N4057);
xor XOR2 (N11836, N11826, N3619);
not NOT1 (N11837, N11811);
or OR2 (N11838, N11835, N11760);
and AND2 (N11839, N11830, N7920);
nand NAND2 (N11840, N11825, N357);
and AND4 (N11841, N11833, N8062, N8138, N191);
nand NAND4 (N11842, N11824, N3718, N8442, N8279);
xor XOR2 (N11843, N11832, N4255);
buf BUF1 (N11844, N11838);
not NOT1 (N11845, N11839);
nand NAND2 (N11846, N11843, N4291);
or OR2 (N11847, N11836, N9539);
not NOT1 (N11848, N11841);
not NOT1 (N11849, N11848);
buf BUF1 (N11850, N11849);
nand NAND2 (N11851, N11847, N8170);
and AND3 (N11852, N11850, N11292, N518);
xor XOR2 (N11853, N11837, N8581);
buf BUF1 (N11854, N11852);
nand NAND2 (N11855, N11854, N4648);
buf BUF1 (N11856, N11853);
nor NOR2 (N11857, N11840, N4939);
nand NAND2 (N11858, N11856, N3550);
or OR2 (N11859, N11858, N6429);
nor NOR4 (N11860, N11846, N7099, N8250, N4297);
not NOT1 (N11861, N11855);
not NOT1 (N11862, N11857);
or OR3 (N11863, N11844, N2082, N3742);
and AND3 (N11864, N11845, N1682, N10501);
buf BUF1 (N11865, N11861);
or OR4 (N11866, N11851, N9342, N349, N4472);
xor XOR2 (N11867, N11817, N11619);
not NOT1 (N11868, N11866);
and AND2 (N11869, N11864, N3894);
not NOT1 (N11870, N11862);
nand NAND4 (N11871, N11822, N10160, N6647, N11842);
and AND3 (N11872, N71, N6007, N6089);
or OR4 (N11873, N11860, N8458, N7657, N10094);
and AND3 (N11874, N11871, N117, N4064);
not NOT1 (N11875, N11863);
xor XOR2 (N11876, N11872, N10967);
and AND3 (N11877, N11869, N4346, N8849);
buf BUF1 (N11878, N11868);
nor NOR4 (N11879, N11873, N1481, N1149, N3732);
nor NOR3 (N11880, N11867, N10543, N8508);
or OR4 (N11881, N11875, N1616, N11001, N4699);
xor XOR2 (N11882, N11865, N2164);
nor NOR2 (N11883, N11879, N739);
not NOT1 (N11884, N11883);
nand NAND2 (N11885, N11859, N1197);
xor XOR2 (N11886, N11877, N5477);
or OR2 (N11887, N11876, N2343);
xor XOR2 (N11888, N11882, N2364);
or OR3 (N11889, N11870, N9497, N163);
buf BUF1 (N11890, N11878);
or OR4 (N11891, N11888, N6713, N11196, N9824);
or OR4 (N11892, N11891, N2056, N6889, N5545);
or OR3 (N11893, N11884, N8021, N11437);
and AND3 (N11894, N11886, N7653, N308);
not NOT1 (N11895, N11893);
nand NAND2 (N11896, N11885, N10488);
not NOT1 (N11897, N11894);
or OR4 (N11898, N11881, N7128, N5360, N11162);
xor XOR2 (N11899, N11892, N6879);
nand NAND2 (N11900, N11895, N3961);
nand NAND3 (N11901, N11887, N6020, N7472);
xor XOR2 (N11902, N11901, N3659);
nor NOR4 (N11903, N11897, N788, N3377, N11466);
buf BUF1 (N11904, N11899);
nor NOR4 (N11905, N11902, N10884, N7657, N4376);
xor XOR2 (N11906, N11904, N1018);
and AND3 (N11907, N11900, N7093, N5800);
not NOT1 (N11908, N11907);
nor NOR2 (N11909, N11905, N5934);
nor NOR2 (N11910, N11874, N9814);
nand NAND4 (N11911, N11903, N8565, N8491, N9148);
not NOT1 (N11912, N11896);
and AND4 (N11913, N11911, N1741, N6689, N7560);
nor NOR2 (N11914, N11890, N2000);
nand NAND4 (N11915, N11912, N1439, N6615, N8365);
not NOT1 (N11916, N11910);
or OR4 (N11917, N11909, N11802, N4771, N7975);
xor XOR2 (N11918, N11916, N7976);
or OR3 (N11919, N11898, N541, N11712);
nand NAND4 (N11920, N11913, N951, N476, N8361);
buf BUF1 (N11921, N11917);
nor NOR2 (N11922, N11915, N9969);
xor XOR2 (N11923, N11906, N901);
buf BUF1 (N11924, N11889);
and AND3 (N11925, N11908, N10340, N9518);
or OR3 (N11926, N11922, N11500, N6543);
nor NOR4 (N11927, N11925, N9513, N2262, N3858);
and AND2 (N11928, N11920, N1182);
or OR4 (N11929, N11880, N3536, N4961, N8348);
not NOT1 (N11930, N11914);
not NOT1 (N11931, N11924);
nor NOR2 (N11932, N11929, N11595);
nor NOR2 (N11933, N11927, N2697);
or OR2 (N11934, N11923, N6868);
nand NAND2 (N11935, N11919, N6064);
and AND2 (N11936, N11918, N8631);
buf BUF1 (N11937, N11932);
not NOT1 (N11938, N11928);
and AND3 (N11939, N11934, N2508, N9512);
nand NAND3 (N11940, N11931, N10975, N8294);
or OR3 (N11941, N11930, N1261, N2786);
xor XOR2 (N11942, N11937, N2914);
or OR3 (N11943, N11942, N7258, N1161);
buf BUF1 (N11944, N11940);
buf BUF1 (N11945, N11941);
nand NAND3 (N11946, N11935, N190, N7722);
or OR4 (N11947, N11945, N6734, N1037, N8876);
nor NOR4 (N11948, N11921, N6226, N1167, N8478);
xor XOR2 (N11949, N11933, N4823);
nand NAND3 (N11950, N11949, N77, N6316);
nor NOR2 (N11951, N11943, N5552);
buf BUF1 (N11952, N11936);
nor NOR4 (N11953, N11950, N6545, N9144, N8321);
not NOT1 (N11954, N11944);
and AND4 (N11955, N11947, N4849, N1592, N8525);
buf BUF1 (N11956, N11952);
not NOT1 (N11957, N11953);
nor NOR3 (N11958, N11926, N297, N8758);
nand NAND3 (N11959, N11958, N6971, N1678);
nor NOR3 (N11960, N11959, N11337, N2909);
or OR2 (N11961, N11955, N8473);
or OR3 (N11962, N11961, N4975, N8702);
xor XOR2 (N11963, N11951, N4765);
and AND2 (N11964, N11962, N3486);
not NOT1 (N11965, N11964);
nand NAND2 (N11966, N11954, N4855);
and AND3 (N11967, N11939, N3657, N6445);
nor NOR3 (N11968, N11957, N7955, N3406);
and AND2 (N11969, N11967, N589);
and AND3 (N11970, N11938, N3023, N7399);
and AND2 (N11971, N11966, N9920);
nor NOR2 (N11972, N11969, N4080);
and AND4 (N11973, N11963, N234, N5202, N11219);
xor XOR2 (N11974, N11965, N1191);
nand NAND2 (N11975, N11971, N781);
xor XOR2 (N11976, N11970, N93);
nor NOR3 (N11977, N11972, N1749, N5625);
or OR2 (N11978, N11973, N8425);
nor NOR3 (N11979, N11948, N798, N5410);
xor XOR2 (N11980, N11946, N10789);
or OR2 (N11981, N11980, N11007);
nor NOR2 (N11982, N11956, N10857);
buf BUF1 (N11983, N11968);
and AND2 (N11984, N11979, N10765);
and AND2 (N11985, N11978, N7775);
nand NAND3 (N11986, N11974, N2648, N5262);
not NOT1 (N11987, N11975);
or OR4 (N11988, N11986, N5244, N5009, N6540);
or OR2 (N11989, N11985, N3484);
not NOT1 (N11990, N11987);
xor XOR2 (N11991, N11976, N11765);
xor XOR2 (N11992, N11988, N3156);
and AND3 (N11993, N11977, N11049, N11515);
or OR4 (N11994, N11991, N6930, N9865, N1292);
or OR4 (N11995, N11982, N10949, N302, N10938);
buf BUF1 (N11996, N11983);
not NOT1 (N11997, N11996);
not NOT1 (N11998, N11981);
nor NOR4 (N11999, N11960, N6090, N3038, N5250);
or OR3 (N12000, N11994, N10472, N11634);
buf BUF1 (N12001, N11992);
buf BUF1 (N12002, N11998);
and AND3 (N12003, N11997, N8706, N4775);
xor XOR2 (N12004, N11999, N10496);
buf BUF1 (N12005, N11993);
xor XOR2 (N12006, N12001, N3600);
or OR4 (N12007, N11989, N1396, N7240, N7041);
nand NAND2 (N12008, N12003, N9085);
nand NAND3 (N12009, N11995, N318, N7767);
nand NAND4 (N12010, N12006, N10566, N2226, N5860);
nor NOR3 (N12011, N12004, N3025, N3159);
xor XOR2 (N12012, N12011, N9454);
nor NOR3 (N12013, N12002, N261, N253);
not NOT1 (N12014, N12010);
xor XOR2 (N12015, N11990, N11833);
nor NOR4 (N12016, N11984, N1292, N10231, N325);
and AND3 (N12017, N12015, N5173, N1408);
xor XOR2 (N12018, N12013, N9623);
or OR4 (N12019, N12017, N1563, N10004, N4978);
or OR3 (N12020, N12018, N11348, N2169);
not NOT1 (N12021, N12016);
nor NOR4 (N12022, N12009, N8634, N11205, N7412);
buf BUF1 (N12023, N12005);
buf BUF1 (N12024, N12020);
not NOT1 (N12025, N12022);
not NOT1 (N12026, N12019);
xor XOR2 (N12027, N12008, N11736);
and AND3 (N12028, N12026, N1379, N7318);
xor XOR2 (N12029, N12023, N10502);
not NOT1 (N12030, N12025);
xor XOR2 (N12031, N12029, N2881);
nand NAND2 (N12032, N12012, N4309);
not NOT1 (N12033, N12014);
xor XOR2 (N12034, N12000, N10957);
xor XOR2 (N12035, N12034, N690);
buf BUF1 (N12036, N12035);
nor NOR3 (N12037, N12030, N7613, N7964);
buf BUF1 (N12038, N12031);
buf BUF1 (N12039, N12036);
not NOT1 (N12040, N12032);
and AND3 (N12041, N12021, N5570, N9355);
or OR2 (N12042, N12007, N926);
xor XOR2 (N12043, N12027, N6184);
buf BUF1 (N12044, N12039);
not NOT1 (N12045, N12043);
nor NOR3 (N12046, N12040, N7383, N11279);
buf BUF1 (N12047, N12037);
and AND3 (N12048, N12044, N4639, N8660);
nor NOR4 (N12049, N12048, N3376, N10260, N9261);
buf BUF1 (N12050, N12046);
xor XOR2 (N12051, N12038, N4158);
not NOT1 (N12052, N12024);
or OR4 (N12053, N12028, N3502, N2756, N953);
buf BUF1 (N12054, N12041);
nor NOR3 (N12055, N12049, N11966, N4466);
buf BUF1 (N12056, N12047);
and AND4 (N12057, N12056, N9021, N6221, N2774);
nor NOR2 (N12058, N12057, N6125);
nor NOR2 (N12059, N12052, N2596);
xor XOR2 (N12060, N12042, N9735);
nor NOR3 (N12061, N12053, N5865, N4689);
xor XOR2 (N12062, N12051, N2047);
and AND3 (N12063, N12062, N2944, N11924);
or OR2 (N12064, N12055, N9084);
not NOT1 (N12065, N12063);
nor NOR3 (N12066, N12045, N3750, N2505);
nor NOR3 (N12067, N12059, N10977, N1784);
nand NAND3 (N12068, N12054, N3981, N947);
buf BUF1 (N12069, N12050);
buf BUF1 (N12070, N12068);
buf BUF1 (N12071, N12070);
buf BUF1 (N12072, N12033);
or OR3 (N12073, N12058, N4552, N8303);
xor XOR2 (N12074, N12061, N224);
not NOT1 (N12075, N12071);
nor NOR2 (N12076, N12072, N4380);
nand NAND3 (N12077, N12074, N11563, N11455);
not NOT1 (N12078, N12067);
buf BUF1 (N12079, N12073);
buf BUF1 (N12080, N12076);
and AND3 (N12081, N12078, N11119, N2005);
nor NOR2 (N12082, N12079, N9415);
buf BUF1 (N12083, N12080);
xor XOR2 (N12084, N12082, N3726);
buf BUF1 (N12085, N12077);
nand NAND4 (N12086, N12083, N12041, N3997, N11677);
nor NOR3 (N12087, N12085, N265, N1845);
and AND3 (N12088, N12066, N8531, N1629);
buf BUF1 (N12089, N12086);
nor NOR2 (N12090, N12064, N4563);
xor XOR2 (N12091, N12087, N2809);
or OR4 (N12092, N12091, N2479, N417, N1310);
nand NAND2 (N12093, N12075, N800);
nand NAND3 (N12094, N12065, N9454, N10487);
and AND4 (N12095, N12088, N4231, N1335, N5025);
xor XOR2 (N12096, N12084, N11087);
or OR3 (N12097, N12089, N4615, N6060);
nor NOR3 (N12098, N12090, N4824, N4643);
not NOT1 (N12099, N12098);
not NOT1 (N12100, N12099);
xor XOR2 (N12101, N12060, N6862);
nor NOR2 (N12102, N12092, N2671);
buf BUF1 (N12103, N12095);
or OR3 (N12104, N12096, N5143, N422);
and AND2 (N12105, N12104, N737);
nand NAND4 (N12106, N12101, N10270, N10216, N6146);
buf BUF1 (N12107, N12103);
nand NAND3 (N12108, N12094, N6156, N6221);
nor NOR4 (N12109, N12100, N9808, N5359, N4689);
buf BUF1 (N12110, N12105);
or OR2 (N12111, N12106, N6548);
and AND2 (N12112, N12111, N4750);
or OR4 (N12113, N12097, N8311, N6178, N4621);
buf BUF1 (N12114, N12081);
xor XOR2 (N12115, N12112, N11237);
xor XOR2 (N12116, N12114, N10268);
or OR2 (N12117, N12107, N11226);
nand NAND4 (N12118, N12108, N9375, N8396, N9632);
or OR2 (N12119, N12116, N8996);
buf BUF1 (N12120, N12109);
xor XOR2 (N12121, N12102, N3202);
xor XOR2 (N12122, N12118, N2470);
and AND2 (N12123, N12119, N9962);
nor NOR2 (N12124, N12122, N7897);
or OR3 (N12125, N12110, N11689, N3717);
nand NAND3 (N12126, N12093, N3438, N6425);
buf BUF1 (N12127, N12115);
nor NOR4 (N12128, N12120, N11551, N8433, N7821);
buf BUF1 (N12129, N12128);
not NOT1 (N12130, N12126);
buf BUF1 (N12131, N12123);
not NOT1 (N12132, N12069);
nor NOR4 (N12133, N12124, N1255, N8623, N10904);
nand NAND4 (N12134, N12133, N9156, N5465, N3093);
and AND4 (N12135, N12117, N10573, N1314, N3078);
and AND4 (N12136, N12131, N3742, N5297, N1879);
buf BUF1 (N12137, N12129);
xor XOR2 (N12138, N12135, N8152);
buf BUF1 (N12139, N12138);
buf BUF1 (N12140, N12132);
not NOT1 (N12141, N12140);
buf BUF1 (N12142, N12136);
not NOT1 (N12143, N12134);
and AND3 (N12144, N12137, N11684, N3385);
not NOT1 (N12145, N12142);
not NOT1 (N12146, N12145);
or OR3 (N12147, N12144, N3326, N918);
buf BUF1 (N12148, N12141);
nand NAND2 (N12149, N12146, N10394);
not NOT1 (N12150, N12127);
xor XOR2 (N12151, N12139, N8561);
buf BUF1 (N12152, N12151);
and AND3 (N12153, N12121, N10304, N7816);
or OR3 (N12154, N12143, N2035, N2408);
nor NOR4 (N12155, N12125, N3065, N715, N7631);
not NOT1 (N12156, N12154);
nor NOR3 (N12157, N12152, N7750, N9534);
not NOT1 (N12158, N12153);
xor XOR2 (N12159, N12150, N11439);
buf BUF1 (N12160, N12149);
buf BUF1 (N12161, N12147);
xor XOR2 (N12162, N12155, N2693);
or OR2 (N12163, N12159, N6917);
xor XOR2 (N12164, N12161, N3830);
buf BUF1 (N12165, N12164);
buf BUF1 (N12166, N12148);
buf BUF1 (N12167, N12163);
not NOT1 (N12168, N12162);
nor NOR4 (N12169, N12168, N2368, N10248, N11600);
or OR3 (N12170, N12160, N10269, N11188);
nand NAND2 (N12171, N12169, N3950);
or OR2 (N12172, N12113, N8738);
not NOT1 (N12173, N12170);
xor XOR2 (N12174, N12165, N12112);
xor XOR2 (N12175, N12130, N6581);
and AND2 (N12176, N12167, N2570);
buf BUF1 (N12177, N12172);
xor XOR2 (N12178, N12166, N11818);
and AND2 (N12179, N12156, N9412);
nor NOR3 (N12180, N12178, N11959, N42);
nor NOR2 (N12181, N12176, N10604);
buf BUF1 (N12182, N12175);
nand NAND2 (N12183, N12158, N9608);
not NOT1 (N12184, N12183);
buf BUF1 (N12185, N12182);
and AND4 (N12186, N12173, N5121, N12012, N8163);
and AND2 (N12187, N12180, N1184);
xor XOR2 (N12188, N12185, N3747);
nor NOR4 (N12189, N12187, N9403, N4943, N6565);
xor XOR2 (N12190, N12171, N11138);
nor NOR2 (N12191, N12188, N7121);
or OR2 (N12192, N12181, N7884);
xor XOR2 (N12193, N12184, N1849);
nand NAND3 (N12194, N12179, N3432, N9008);
nor NOR2 (N12195, N12192, N1544);
not NOT1 (N12196, N12191);
nand NAND3 (N12197, N12195, N80, N64);
or OR4 (N12198, N12177, N1385, N3724, N6764);
nand NAND4 (N12199, N12174, N11057, N11623, N3315);
and AND3 (N12200, N12194, N5120, N5419);
buf BUF1 (N12201, N12197);
nand NAND3 (N12202, N12186, N3925, N1484);
xor XOR2 (N12203, N12190, N8970);
and AND3 (N12204, N12198, N9324, N4787);
or OR3 (N12205, N12204, N284, N35);
and AND2 (N12206, N12157, N11811);
nor NOR4 (N12207, N12206, N7901, N236, N10008);
xor XOR2 (N12208, N12189, N8310);
not NOT1 (N12209, N12200);
not NOT1 (N12210, N12207);
nand NAND2 (N12211, N12205, N2621);
nand NAND4 (N12212, N12193, N6916, N8655, N6632);
nor NOR2 (N12213, N12202, N10119);
buf BUF1 (N12214, N12209);
and AND4 (N12215, N12203, N10529, N11620, N12165);
not NOT1 (N12216, N12210);
or OR3 (N12217, N12211, N8071, N431);
buf BUF1 (N12218, N12215);
nand NAND3 (N12219, N12213, N2903, N2511);
or OR4 (N12220, N12199, N2451, N3006, N4391);
xor XOR2 (N12221, N12201, N9711);
or OR4 (N12222, N12217, N4123, N8462, N11747);
or OR3 (N12223, N12216, N5786, N1066);
xor XOR2 (N12224, N12218, N6609);
nor NOR3 (N12225, N12223, N2537, N8771);
xor XOR2 (N12226, N12220, N5753);
xor XOR2 (N12227, N12222, N5475);
or OR3 (N12228, N12226, N1995, N2213);
and AND3 (N12229, N12196, N66, N9050);
nor NOR2 (N12230, N12214, N6396);
nor NOR4 (N12231, N12230, N10438, N7612, N1943);
or OR4 (N12232, N12221, N8275, N6872, N3648);
xor XOR2 (N12233, N12219, N12065);
nor NOR3 (N12234, N12231, N4041, N4264);
or OR2 (N12235, N12234, N3314);
nor NOR3 (N12236, N12233, N809, N10361);
and AND3 (N12237, N12232, N3322, N10930);
or OR2 (N12238, N12228, N6826);
buf BUF1 (N12239, N12235);
or OR4 (N12240, N12212, N11184, N3561, N8903);
nor NOR4 (N12241, N12237, N8750, N8799, N8762);
xor XOR2 (N12242, N12208, N9214);
and AND3 (N12243, N12239, N8408, N1073);
or OR4 (N12244, N12240, N3580, N8283, N2097);
not NOT1 (N12245, N12229);
or OR3 (N12246, N12236, N1022, N11869);
buf BUF1 (N12247, N12225);
xor XOR2 (N12248, N12247, N2887);
buf BUF1 (N12249, N12238);
nor NOR3 (N12250, N12246, N8363, N406);
not NOT1 (N12251, N12245);
not NOT1 (N12252, N12248);
or OR2 (N12253, N12251, N11145);
not NOT1 (N12254, N12243);
nand NAND4 (N12255, N12252, N1299, N5532, N11812);
and AND4 (N12256, N12249, N8420, N12148, N11603);
and AND3 (N12257, N12227, N9855, N6402);
not NOT1 (N12258, N12250);
xor XOR2 (N12259, N12224, N717);
xor XOR2 (N12260, N12254, N11111);
and AND4 (N12261, N12259, N7874, N9996, N2594);
xor XOR2 (N12262, N12260, N3970);
buf BUF1 (N12263, N12261);
and AND4 (N12264, N12256, N209, N6618, N4820);
nand NAND4 (N12265, N12257, N7044, N10906, N10657);
xor XOR2 (N12266, N12244, N5923);
and AND3 (N12267, N12266, N8562, N4322);
nor NOR3 (N12268, N12263, N6191, N6185);
nand NAND4 (N12269, N12253, N2240, N10805, N7551);
not NOT1 (N12270, N12265);
xor XOR2 (N12271, N12264, N5295);
not NOT1 (N12272, N12258);
nor NOR4 (N12273, N12241, N7656, N11577, N3627);
nor NOR3 (N12274, N12271, N2119, N6819);
not NOT1 (N12275, N12274);
nand NAND2 (N12276, N12255, N6492);
not NOT1 (N12277, N12262);
not NOT1 (N12278, N12268);
buf BUF1 (N12279, N12272);
and AND3 (N12280, N12278, N2835, N1202);
nand NAND3 (N12281, N12273, N2923, N11119);
nor NOR4 (N12282, N12275, N2665, N3082, N4254);
not NOT1 (N12283, N12270);
nand NAND3 (N12284, N12277, N4771, N1501);
buf BUF1 (N12285, N12267);
not NOT1 (N12286, N12281);
nor NOR2 (N12287, N12280, N4236);
nor NOR4 (N12288, N12286, N3608, N4838, N10717);
nand NAND3 (N12289, N12269, N1212, N6640);
or OR3 (N12290, N12288, N3167, N2688);
not NOT1 (N12291, N12282);
and AND2 (N12292, N12284, N3453);
or OR3 (N12293, N12283, N5704, N5369);
and AND3 (N12294, N12287, N6617, N5449);
nor NOR2 (N12295, N12285, N657);
xor XOR2 (N12296, N12294, N6736);
and AND3 (N12297, N12292, N8527, N7730);
or OR4 (N12298, N12291, N1282, N899, N1854);
nor NOR3 (N12299, N12290, N8146, N3665);
not NOT1 (N12300, N12299);
nor NOR2 (N12301, N12297, N4932);
nand NAND3 (N12302, N12298, N12118, N1452);
not NOT1 (N12303, N12289);
xor XOR2 (N12304, N12296, N6159);
xor XOR2 (N12305, N12242, N2127);
nor NOR3 (N12306, N12304, N3624, N10966);
xor XOR2 (N12307, N12276, N11297);
buf BUF1 (N12308, N12295);
not NOT1 (N12309, N12279);
buf BUF1 (N12310, N12305);
nand NAND4 (N12311, N12310, N4500, N7142, N3524);
nand NAND4 (N12312, N12293, N11344, N297, N5300);
nand NAND2 (N12313, N12309, N8439);
buf BUF1 (N12314, N12308);
buf BUF1 (N12315, N12300);
buf BUF1 (N12316, N12302);
xor XOR2 (N12317, N12312, N2697);
nor NOR2 (N12318, N12314, N10211);
nand NAND3 (N12319, N12303, N3745, N2580);
nor NOR4 (N12320, N12317, N345, N2233, N5599);
nand NAND2 (N12321, N12306, N9410);
or OR2 (N12322, N12313, N7711);
xor XOR2 (N12323, N12322, N8540);
nand NAND3 (N12324, N12315, N1076, N10979);
buf BUF1 (N12325, N12323);
buf BUF1 (N12326, N12316);
xor XOR2 (N12327, N12324, N7624);
or OR3 (N12328, N12319, N7021, N12021);
and AND3 (N12329, N12307, N5504, N3089);
not NOT1 (N12330, N12301);
or OR3 (N12331, N12311, N4825, N4581);
xor XOR2 (N12332, N12329, N2087);
and AND3 (N12333, N12325, N4050, N4120);
nand NAND2 (N12334, N12333, N2085);
xor XOR2 (N12335, N12326, N6417);
not NOT1 (N12336, N12335);
and AND3 (N12337, N12328, N3849, N4723);
nand NAND3 (N12338, N12327, N1664, N11149);
nand NAND4 (N12339, N12334, N1360, N2134, N7810);
xor XOR2 (N12340, N12336, N3377);
nand NAND2 (N12341, N12338, N448);
xor XOR2 (N12342, N12337, N2292);
buf BUF1 (N12343, N12339);
buf BUF1 (N12344, N12321);
xor XOR2 (N12345, N12344, N4772);
not NOT1 (N12346, N12343);
nand NAND2 (N12347, N12318, N11910);
or OR2 (N12348, N12330, N6907);
or OR3 (N12349, N12347, N1810, N8693);
and AND3 (N12350, N12331, N6668, N5347);
and AND2 (N12351, N12346, N4144);
buf BUF1 (N12352, N12341);
buf BUF1 (N12353, N12348);
buf BUF1 (N12354, N12351);
nand NAND2 (N12355, N12350, N614);
not NOT1 (N12356, N12355);
not NOT1 (N12357, N12340);
buf BUF1 (N12358, N12332);
nand NAND4 (N12359, N12320, N11631, N1688, N1934);
nand NAND4 (N12360, N12354, N12221, N8823, N5748);
nor NOR3 (N12361, N12360, N2026, N8582);
and AND4 (N12362, N12345, N7720, N7712, N1330);
nor NOR4 (N12363, N12359, N1794, N2905, N3242);
not NOT1 (N12364, N12352);
nand NAND4 (N12365, N12364, N11801, N9923, N3482);
not NOT1 (N12366, N12362);
buf BUF1 (N12367, N12356);
or OR4 (N12368, N12353, N9994, N2110, N3946);
xor XOR2 (N12369, N12366, N9193);
not NOT1 (N12370, N12363);
or OR2 (N12371, N12357, N9430);
not NOT1 (N12372, N12370);
nand NAND4 (N12373, N12369, N9208, N8927, N6746);
or OR3 (N12374, N12373, N8714, N3215);
not NOT1 (N12375, N12342);
nor NOR4 (N12376, N12361, N8638, N1385, N10136);
or OR4 (N12377, N12365, N718, N8214, N956);
and AND2 (N12378, N12375, N8396);
nor NOR2 (N12379, N12371, N8394);
nand NAND3 (N12380, N12377, N12058, N7701);
nor NOR3 (N12381, N12367, N5468, N1000);
not NOT1 (N12382, N12380);
or OR3 (N12383, N12349, N10886, N6029);
and AND4 (N12384, N12381, N8390, N7384, N3904);
xor XOR2 (N12385, N12358, N5241);
and AND3 (N12386, N12379, N5836, N8134);
nand NAND2 (N12387, N12372, N694);
xor XOR2 (N12388, N12368, N4232);
xor XOR2 (N12389, N12376, N6788);
not NOT1 (N12390, N12385);
nand NAND3 (N12391, N12389, N11797, N3372);
xor XOR2 (N12392, N12390, N10293);
nand NAND4 (N12393, N12392, N179, N814, N5243);
or OR4 (N12394, N12384, N7335, N10492, N11450);
buf BUF1 (N12395, N12387);
xor XOR2 (N12396, N12382, N1534);
xor XOR2 (N12397, N12378, N12156);
buf BUF1 (N12398, N12386);
nand NAND3 (N12399, N12397, N11596, N6512);
nor NOR2 (N12400, N12394, N1698);
buf BUF1 (N12401, N12395);
or OR4 (N12402, N12400, N11843, N8564, N3369);
buf BUF1 (N12403, N12402);
xor XOR2 (N12404, N12374, N6240);
or OR2 (N12405, N12403, N11823);
buf BUF1 (N12406, N12404);
nor NOR3 (N12407, N12396, N1310, N8871);
not NOT1 (N12408, N12388);
and AND2 (N12409, N12391, N3139);
buf BUF1 (N12410, N12406);
not NOT1 (N12411, N12399);
nand NAND2 (N12412, N12393, N10138);
buf BUF1 (N12413, N12409);
or OR3 (N12414, N12401, N6901, N10566);
and AND2 (N12415, N12408, N7276);
nand NAND3 (N12416, N12411, N7730, N2811);
and AND4 (N12417, N12414, N8754, N10407, N7249);
or OR2 (N12418, N12407, N1064);
or OR2 (N12419, N12416, N11358);
buf BUF1 (N12420, N12415);
xor XOR2 (N12421, N12417, N38);
xor XOR2 (N12422, N12410, N9640);
buf BUF1 (N12423, N12418);
and AND2 (N12424, N12419, N1636);
nor NOR4 (N12425, N12383, N2409, N4071, N10547);
not NOT1 (N12426, N12424);
xor XOR2 (N12427, N12422, N4866);
nor NOR2 (N12428, N12412, N10439);
not NOT1 (N12429, N12426);
not NOT1 (N12430, N12413);
xor XOR2 (N12431, N12429, N7497);
not NOT1 (N12432, N12405);
xor XOR2 (N12433, N12432, N1724);
not NOT1 (N12434, N12430);
nand NAND2 (N12435, N12425, N4333);
not NOT1 (N12436, N12431);
not NOT1 (N12437, N12420);
nor NOR3 (N12438, N12421, N5748, N1436);
and AND2 (N12439, N12438, N1185);
or OR2 (N12440, N12437, N6295);
nand NAND4 (N12441, N12440, N4403, N7844, N4704);
xor XOR2 (N12442, N12423, N11389);
not NOT1 (N12443, N12436);
and AND3 (N12444, N12398, N12041, N8868);
and AND2 (N12445, N12434, N3875);
not NOT1 (N12446, N12445);
nand NAND2 (N12447, N12428, N9959);
buf BUF1 (N12448, N12435);
buf BUF1 (N12449, N12443);
not NOT1 (N12450, N12442);
or OR2 (N12451, N12444, N3177);
and AND3 (N12452, N12448, N998, N10732);
nand NAND4 (N12453, N12427, N1571, N2776, N3181);
buf BUF1 (N12454, N12450);
buf BUF1 (N12455, N12446);
nor NOR2 (N12456, N12439, N7202);
buf BUF1 (N12457, N12455);
nor NOR4 (N12458, N12451, N6514, N7255, N6467);
nor NOR4 (N12459, N12456, N1753, N11202, N1007);
nor NOR3 (N12460, N12458, N1975, N1240);
buf BUF1 (N12461, N12454);
not NOT1 (N12462, N12447);
xor XOR2 (N12463, N12433, N8670);
nor NOR2 (N12464, N12463, N1883);
not NOT1 (N12465, N12461);
nand NAND2 (N12466, N12452, N5158);
buf BUF1 (N12467, N12465);
not NOT1 (N12468, N12459);
and AND3 (N12469, N12449, N8160, N2503);
nand NAND3 (N12470, N12467, N5016, N3891);
or OR2 (N12471, N12470, N6148);
or OR4 (N12472, N12469, N3062, N3372, N12302);
nand NAND4 (N12473, N12460, N10675, N8649, N6373);
nand NAND4 (N12474, N12472, N7899, N6138, N11316);
nor NOR2 (N12475, N12468, N11991);
and AND3 (N12476, N12457, N9558, N4988);
xor XOR2 (N12477, N12473, N7750);
xor XOR2 (N12478, N12476, N10210);
nor NOR4 (N12479, N12441, N9841, N7488, N4651);
nor NOR4 (N12480, N12474, N6372, N12333, N6070);
xor XOR2 (N12481, N12477, N12103);
or OR4 (N12482, N12479, N1139, N8995, N1355);
or OR4 (N12483, N12475, N4185, N2656, N6495);
xor XOR2 (N12484, N12471, N8746);
nor NOR2 (N12485, N12481, N9093);
xor XOR2 (N12486, N12483, N5859);
xor XOR2 (N12487, N12464, N2485);
xor XOR2 (N12488, N12478, N8623);
xor XOR2 (N12489, N12480, N10185);
xor XOR2 (N12490, N12462, N4151);
not NOT1 (N12491, N12453);
not NOT1 (N12492, N12487);
xor XOR2 (N12493, N12485, N1405);
nor NOR3 (N12494, N12493, N6145, N5646);
nand NAND3 (N12495, N12494, N866, N5334);
not NOT1 (N12496, N12490);
buf BUF1 (N12497, N12482);
xor XOR2 (N12498, N12486, N2141);
buf BUF1 (N12499, N12496);
not NOT1 (N12500, N12498);
buf BUF1 (N12501, N12499);
not NOT1 (N12502, N12501);
nor NOR2 (N12503, N12500, N220);
nor NOR3 (N12504, N12491, N1847, N4967);
and AND4 (N12505, N12488, N11498, N2377, N12296);
nand NAND4 (N12506, N12495, N2914, N4081, N12439);
buf BUF1 (N12507, N12497);
xor XOR2 (N12508, N12489, N11724);
not NOT1 (N12509, N12466);
nor NOR4 (N12510, N12507, N5423, N2673, N11398);
or OR4 (N12511, N12492, N5947, N10012, N5052);
nor NOR4 (N12512, N12506, N3973, N4178, N5615);
nand NAND4 (N12513, N12484, N2179, N11784, N10336);
xor XOR2 (N12514, N12503, N12027);
buf BUF1 (N12515, N12502);
nor NOR2 (N12516, N12510, N11742);
nor NOR3 (N12517, N12509, N9992, N4371);
xor XOR2 (N12518, N12515, N1541);
buf BUF1 (N12519, N12517);
buf BUF1 (N12520, N12514);
nand NAND4 (N12521, N12519, N10509, N9435, N3507);
xor XOR2 (N12522, N12504, N7144);
nand NAND3 (N12523, N12511, N7516, N1645);
and AND3 (N12524, N12508, N6361, N4713);
and AND3 (N12525, N12521, N2842, N3845);
buf BUF1 (N12526, N12518);
nand NAND4 (N12527, N12524, N12235, N11244, N268);
or OR2 (N12528, N12522, N11505);
and AND2 (N12529, N12527, N876);
buf BUF1 (N12530, N12513);
buf BUF1 (N12531, N12505);
nand NAND2 (N12532, N12528, N4957);
xor XOR2 (N12533, N12525, N5386);
xor XOR2 (N12534, N12520, N11192);
or OR4 (N12535, N12533, N6288, N4805, N8457);
nand NAND3 (N12536, N12529, N3247, N3500);
or OR4 (N12537, N12516, N4651, N3960, N10188);
xor XOR2 (N12538, N12512, N9916);
and AND4 (N12539, N12537, N4268, N9292, N1243);
buf BUF1 (N12540, N12534);
buf BUF1 (N12541, N12540);
xor XOR2 (N12542, N12532, N5689);
nand NAND2 (N12543, N12526, N8778);
nand NAND3 (N12544, N12530, N8232, N12078);
xor XOR2 (N12545, N12536, N154);
xor XOR2 (N12546, N12523, N11829);
xor XOR2 (N12547, N12541, N508);
not NOT1 (N12548, N12539);
xor XOR2 (N12549, N12547, N4963);
nor NOR4 (N12550, N12545, N7593, N5828, N7840);
buf BUF1 (N12551, N12535);
buf BUF1 (N12552, N12542);
nor NOR2 (N12553, N12549, N9634);
nor NOR3 (N12554, N12531, N11286, N10866);
nor NOR4 (N12555, N12552, N10627, N4979, N5208);
nor NOR4 (N12556, N12548, N2507, N7158, N3193);
buf BUF1 (N12557, N12554);
buf BUF1 (N12558, N12551);
xor XOR2 (N12559, N12544, N11865);
not NOT1 (N12560, N12558);
or OR2 (N12561, N12556, N6450);
xor XOR2 (N12562, N12553, N6768);
nor NOR4 (N12563, N12559, N7134, N8978, N3212);
nand NAND2 (N12564, N12560, N5088);
buf BUF1 (N12565, N12563);
nand NAND4 (N12566, N12557, N12491, N3384, N11522);
xor XOR2 (N12567, N12555, N7668);
buf BUF1 (N12568, N12550);
xor XOR2 (N12569, N12562, N9980);
and AND3 (N12570, N12567, N1957, N8731);
nor NOR4 (N12571, N12538, N797, N6044, N3437);
nand NAND3 (N12572, N12565, N10393, N8594);
or OR2 (N12573, N12561, N12402);
and AND3 (N12574, N12572, N10176, N12456);
xor XOR2 (N12575, N12569, N4543);
or OR3 (N12576, N12574, N7104, N10190);
nor NOR4 (N12577, N12570, N7927, N1432, N903);
xor XOR2 (N12578, N12576, N8778);
and AND4 (N12579, N12568, N4084, N5953, N7991);
xor XOR2 (N12580, N12575, N4652);
nand NAND3 (N12581, N12580, N12478, N12106);
nor NOR2 (N12582, N12564, N2723);
not NOT1 (N12583, N12577);
xor XOR2 (N12584, N12566, N8854);
buf BUF1 (N12585, N12571);
xor XOR2 (N12586, N12579, N1989);
nand NAND2 (N12587, N12546, N9957);
buf BUF1 (N12588, N12585);
nor NOR4 (N12589, N12582, N11712, N8866, N8856);
nand NAND4 (N12590, N12578, N2627, N2798, N4189);
or OR4 (N12591, N12573, N9112, N4320, N12361);
not NOT1 (N12592, N12588);
buf BUF1 (N12593, N12586);
or OR2 (N12594, N12584, N879);
buf BUF1 (N12595, N12591);
not NOT1 (N12596, N12594);
xor XOR2 (N12597, N12590, N7511);
not NOT1 (N12598, N12583);
not NOT1 (N12599, N12587);
buf BUF1 (N12600, N12593);
buf BUF1 (N12601, N12543);
buf BUF1 (N12602, N12598);
xor XOR2 (N12603, N12596, N446);
buf BUF1 (N12604, N12597);
and AND4 (N12605, N12601, N893, N6642, N7293);
or OR2 (N12606, N12589, N6227);
and AND3 (N12607, N12606, N6479, N4570);
and AND2 (N12608, N12602, N10231);
buf BUF1 (N12609, N12595);
nor NOR3 (N12610, N12603, N6283, N2384);
or OR2 (N12611, N12604, N9797);
or OR4 (N12612, N12581, N3557, N9280, N1174);
nand NAND4 (N12613, N12610, N8759, N5421, N4813);
nor NOR3 (N12614, N12613, N7917, N2189);
xor XOR2 (N12615, N12605, N9089);
not NOT1 (N12616, N12609);
buf BUF1 (N12617, N12612);
or OR3 (N12618, N12615, N9077, N11611);
not NOT1 (N12619, N12592);
and AND4 (N12620, N12616, N3637, N9095, N6436);
not NOT1 (N12621, N12599);
nand NAND2 (N12622, N12614, N3247);
and AND4 (N12623, N12600, N10256, N7741, N6441);
buf BUF1 (N12624, N12623);
and AND2 (N12625, N12618, N5693);
nor NOR2 (N12626, N12625, N3091);
or OR4 (N12627, N12611, N3570, N4819, N4668);
not NOT1 (N12628, N12617);
and AND2 (N12629, N12619, N11508);
or OR4 (N12630, N12608, N10925, N4547, N639);
buf BUF1 (N12631, N12607);
not NOT1 (N12632, N12631);
or OR4 (N12633, N12627, N10991, N1691, N6608);
buf BUF1 (N12634, N12633);
xor XOR2 (N12635, N12621, N7717);
buf BUF1 (N12636, N12634);
xor XOR2 (N12637, N12626, N8703);
and AND3 (N12638, N12622, N8177, N8177);
and AND4 (N12639, N12638, N5899, N7904, N11137);
and AND3 (N12640, N12628, N9549, N8366);
buf BUF1 (N12641, N12624);
nand NAND3 (N12642, N12639, N8316, N8592);
nor NOR2 (N12643, N12641, N10785);
or OR4 (N12644, N12637, N2108, N3898, N8477);
and AND4 (N12645, N12642, N5318, N1816, N11703);
nand NAND3 (N12646, N12635, N2070, N2131);
or OR3 (N12647, N12645, N1811, N657);
and AND4 (N12648, N12620, N5514, N8533, N10506);
or OR3 (N12649, N12647, N4938, N2287);
nand NAND2 (N12650, N12646, N10954);
not NOT1 (N12651, N12644);
nand NAND2 (N12652, N12649, N1702);
xor XOR2 (N12653, N12643, N8790);
buf BUF1 (N12654, N12632);
buf BUF1 (N12655, N12648);
not NOT1 (N12656, N12650);
not NOT1 (N12657, N12640);
and AND4 (N12658, N12636, N9668, N6671, N796);
or OR2 (N12659, N12654, N7052);
or OR4 (N12660, N12657, N2148, N11052, N12021);
not NOT1 (N12661, N12652);
nand NAND3 (N12662, N12655, N6377, N6513);
and AND4 (N12663, N12656, N6752, N7075, N3906);
buf BUF1 (N12664, N12661);
nand NAND3 (N12665, N12664, N2173, N11986);
nor NOR4 (N12666, N12651, N586, N1547, N2286);
or OR4 (N12667, N12662, N9882, N11525, N2844);
buf BUF1 (N12668, N12660);
or OR3 (N12669, N12658, N11171, N1301);
xor XOR2 (N12670, N12669, N790);
or OR3 (N12671, N12629, N3567, N2823);
xor XOR2 (N12672, N12663, N2312);
not NOT1 (N12673, N12668);
nor NOR3 (N12674, N12653, N130, N6879);
not NOT1 (N12675, N12672);
nor NOR2 (N12676, N12665, N5577);
buf BUF1 (N12677, N12670);
and AND4 (N12678, N12673, N5707, N10719, N7259);
or OR2 (N12679, N12677, N676);
buf BUF1 (N12680, N12671);
buf BUF1 (N12681, N12680);
xor XOR2 (N12682, N12679, N1014);
nand NAND3 (N12683, N12666, N4591, N2032);
xor XOR2 (N12684, N12678, N8160);
or OR3 (N12685, N12667, N12527, N1438);
nand NAND2 (N12686, N12676, N4510);
nor NOR3 (N12687, N12685, N6612, N3190);
xor XOR2 (N12688, N12687, N5738);
nand NAND4 (N12689, N12675, N11806, N8988, N6891);
xor XOR2 (N12690, N12674, N4611);
buf BUF1 (N12691, N12689);
or OR2 (N12692, N12659, N11642);
and AND2 (N12693, N12690, N8167);
nand NAND2 (N12694, N12684, N4018);
or OR3 (N12695, N12682, N10724, N1229);
and AND2 (N12696, N12688, N2019);
or OR3 (N12697, N12630, N4587, N355);
and AND3 (N12698, N12692, N10633, N5346);
nor NOR3 (N12699, N12693, N6297, N9707);
xor XOR2 (N12700, N12686, N7189);
buf BUF1 (N12701, N12683);
not NOT1 (N12702, N12699);
xor XOR2 (N12703, N12702, N4038);
not NOT1 (N12704, N12697);
nand NAND2 (N12705, N12698, N3445);
and AND2 (N12706, N12694, N5702);
not NOT1 (N12707, N12695);
nor NOR2 (N12708, N12705, N4639);
buf BUF1 (N12709, N12706);
and AND3 (N12710, N12709, N3596, N10657);
and AND4 (N12711, N12681, N3567, N1781, N3131);
not NOT1 (N12712, N12710);
buf BUF1 (N12713, N12703);
nor NOR3 (N12714, N12700, N10565, N11526);
or OR3 (N12715, N12708, N6412, N2924);
or OR3 (N12716, N12713, N6675, N2495);
or OR3 (N12717, N12716, N10188, N8409);
not NOT1 (N12718, N12715);
and AND3 (N12719, N12701, N392, N1896);
not NOT1 (N12720, N12704);
buf BUF1 (N12721, N12696);
and AND4 (N12722, N12721, N7008, N145, N5694);
nor NOR4 (N12723, N12720, N664, N10834, N4335);
not NOT1 (N12724, N12723);
nor NOR2 (N12725, N12714, N7928);
and AND3 (N12726, N12707, N11141, N619);
nor NOR4 (N12727, N12717, N7127, N1839, N3716);
not NOT1 (N12728, N12712);
nand NAND4 (N12729, N12711, N10955, N3538, N6807);
nor NOR2 (N12730, N12725, N8406);
nor NOR4 (N12731, N12727, N2225, N1145, N5259);
nor NOR3 (N12732, N12691, N9496, N4220);
or OR3 (N12733, N12728, N11537, N1032);
xor XOR2 (N12734, N12718, N3475);
nor NOR3 (N12735, N12722, N10833, N9131);
not NOT1 (N12736, N12734);
xor XOR2 (N12737, N12729, N4805);
or OR3 (N12738, N12726, N1536, N6812);
nor NOR4 (N12739, N12737, N6470, N7986, N4486);
nor NOR3 (N12740, N12730, N9938, N6522);
buf BUF1 (N12741, N12732);
buf BUF1 (N12742, N12740);
or OR4 (N12743, N12736, N221, N9941, N485);
or OR4 (N12744, N12742, N9638, N2544, N1231);
and AND3 (N12745, N12735, N12599, N7568);
nand NAND4 (N12746, N12739, N12441, N4015, N1830);
buf BUF1 (N12747, N12719);
not NOT1 (N12748, N12746);
not NOT1 (N12749, N12748);
nand NAND3 (N12750, N12733, N11405, N9560);
xor XOR2 (N12751, N12747, N7016);
nand NAND4 (N12752, N12738, N2612, N9023, N2593);
and AND3 (N12753, N12744, N5594, N5153);
xor XOR2 (N12754, N12731, N7373);
or OR3 (N12755, N12754, N10058, N11574);
nand NAND2 (N12756, N12751, N11881);
xor XOR2 (N12757, N12749, N141);
or OR2 (N12758, N12741, N6928);
and AND2 (N12759, N12756, N167);
and AND2 (N12760, N12750, N12322);
nor NOR3 (N12761, N12724, N1262, N2831);
not NOT1 (N12762, N12743);
and AND4 (N12763, N12757, N2468, N9593, N1826);
buf BUF1 (N12764, N12753);
xor XOR2 (N12765, N12759, N5963);
nor NOR2 (N12766, N12765, N12424);
or OR2 (N12767, N12762, N2544);
xor XOR2 (N12768, N12760, N2114);
xor XOR2 (N12769, N12752, N669);
nand NAND4 (N12770, N12763, N9628, N2171, N11556);
not NOT1 (N12771, N12758);
and AND3 (N12772, N12767, N738, N422);
nor NOR4 (N12773, N12769, N9374, N9521, N5521);
xor XOR2 (N12774, N12745, N2727);
not NOT1 (N12775, N12770);
and AND4 (N12776, N12768, N1103, N1548, N4216);
or OR3 (N12777, N12755, N3839, N5515);
nand NAND2 (N12778, N12764, N6959);
and AND2 (N12779, N12773, N8176);
buf BUF1 (N12780, N12761);
nor NOR4 (N12781, N12778, N9394, N5770, N11354);
nor NOR2 (N12782, N12781, N917);
buf BUF1 (N12783, N12772);
nand NAND4 (N12784, N12766, N7068, N656, N3455);
nor NOR4 (N12785, N12784, N3487, N348, N12665);
xor XOR2 (N12786, N12783, N795);
buf BUF1 (N12787, N12782);
and AND3 (N12788, N12774, N8290, N3029);
nand NAND2 (N12789, N12788, N2878);
not NOT1 (N12790, N12780);
or OR2 (N12791, N12787, N11719);
xor XOR2 (N12792, N12789, N11953);
not NOT1 (N12793, N12775);
and AND4 (N12794, N12779, N2268, N2228, N6357);
not NOT1 (N12795, N12786);
or OR3 (N12796, N12794, N4755, N4573);
buf BUF1 (N12797, N12771);
not NOT1 (N12798, N12797);
not NOT1 (N12799, N12785);
nand NAND4 (N12800, N12792, N7966, N1621, N4800);
or OR4 (N12801, N12793, N5376, N1059, N11762);
or OR2 (N12802, N12777, N1295);
or OR4 (N12803, N12799, N10328, N2621, N10377);
nor NOR3 (N12804, N12791, N190, N6210);
and AND3 (N12805, N12796, N4603, N6668);
not NOT1 (N12806, N12795);
not NOT1 (N12807, N12801);
buf BUF1 (N12808, N12802);
and AND4 (N12809, N12805, N8372, N3785, N1320);
buf BUF1 (N12810, N12790);
buf BUF1 (N12811, N12804);
buf BUF1 (N12812, N12806);
xor XOR2 (N12813, N12811, N3671);
buf BUF1 (N12814, N12810);
nand NAND4 (N12815, N12814, N6188, N10848, N8712);
nor NOR2 (N12816, N12809, N12567);
and AND4 (N12817, N12776, N3077, N3807, N11349);
endmodule