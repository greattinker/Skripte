// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23;

output N3522,N3518,N3517,N3505,N3511,N3499,N3519,N3521,N3516,N3523;

xor XOR2 (N24, N23, N15);
and AND4 (N25, N15, N8, N17, N15);
nand NAND4 (N26, N23, N4, N4, N9);
and AND2 (N27, N3, N25);
nand NAND3 (N28, N21, N10, N24);
or OR2 (N29, N18, N1);
nor NOR2 (N30, N23, N1);
buf BUF1 (N31, N4);
nor NOR4 (N32, N30, N27, N30, N24);
nor NOR4 (N33, N17, N30, N26, N24);
or OR4 (N34, N21, N23, N30, N30);
xor XOR2 (N35, N25, N26);
xor XOR2 (N36, N25, N4);
nand NAND3 (N37, N12, N12, N14);
nor NOR4 (N38, N25, N16, N5, N18);
not NOT1 (N39, N37);
nand NAND2 (N40, N31, N26);
xor XOR2 (N41, N32, N10);
not NOT1 (N42, N41);
nor NOR2 (N43, N29, N31);
nand NAND3 (N44, N34, N37, N37);
xor XOR2 (N45, N39, N6);
nor NOR3 (N46, N36, N32, N18);
and AND4 (N47, N40, N3, N13, N6);
nor NOR3 (N48, N33, N38, N24);
xor XOR2 (N49, N23, N36);
and AND2 (N50, N46, N45);
nand NAND3 (N51, N44, N20, N14);
not NOT1 (N52, N3);
nor NOR3 (N53, N52, N34, N44);
nor NOR2 (N54, N53, N17);
nand NAND3 (N55, N43, N45, N34);
buf BUF1 (N56, N54);
buf BUF1 (N57, N47);
nor NOR4 (N58, N57, N48, N27, N8);
xor XOR2 (N59, N54, N17);
nand NAND4 (N60, N58, N49, N53, N23);
or OR4 (N61, N38, N2, N5, N13);
xor XOR2 (N62, N56, N23);
buf BUF1 (N63, N42);
not NOT1 (N64, N55);
nand NAND3 (N65, N28, N63, N14);
buf BUF1 (N66, N5);
nor NOR2 (N67, N51, N47);
not NOT1 (N68, N65);
xor XOR2 (N69, N67, N9);
nor NOR3 (N70, N35, N8, N32);
nor NOR3 (N71, N70, N18, N44);
xor XOR2 (N72, N68, N68);
or OR4 (N73, N62, N1, N35, N1);
or OR2 (N74, N66, N49);
buf BUF1 (N75, N60);
buf BUF1 (N76, N50);
nand NAND2 (N77, N76, N23);
or OR3 (N78, N73, N38, N41);
nor NOR3 (N79, N74, N35, N7);
nand NAND2 (N80, N64, N12);
nand NAND4 (N81, N61, N34, N8, N24);
nor NOR3 (N82, N71, N31, N42);
not NOT1 (N83, N79);
nor NOR3 (N84, N59, N30, N71);
nand NAND3 (N85, N78, N59, N55);
nor NOR3 (N86, N82, N80, N37);
nor NOR2 (N87, N82, N31);
nand NAND2 (N88, N72, N32);
nor NOR3 (N89, N88, N54, N72);
not NOT1 (N90, N83);
and AND3 (N91, N77, N14, N11);
buf BUF1 (N92, N86);
and AND3 (N93, N92, N14, N12);
or OR4 (N94, N89, N56, N49, N70);
or OR4 (N95, N90, N10, N91, N72);
buf BUF1 (N96, N5);
nor NOR2 (N97, N93, N59);
not NOT1 (N98, N84);
nor NOR2 (N99, N85, N93);
or OR3 (N100, N99, N62, N84);
and AND2 (N101, N94, N27);
nor NOR4 (N102, N81, N25, N58, N11);
buf BUF1 (N103, N75);
or OR2 (N104, N98, N9);
nor NOR4 (N105, N69, N61, N79, N34);
and AND4 (N106, N102, N94, N36, N73);
or OR4 (N107, N105, N8, N13, N30);
nor NOR4 (N108, N101, N68, N23, N68);
and AND3 (N109, N103, N48, N65);
or OR4 (N110, N97, N7, N76, N72);
or OR2 (N111, N95, N27);
or OR3 (N112, N104, N43, N64);
xor XOR2 (N113, N87, N23);
or OR2 (N114, N106, N41);
not NOT1 (N115, N107);
nand NAND3 (N116, N111, N66, N3);
or OR4 (N117, N113, N116, N109, N100);
buf BUF1 (N118, N37);
buf BUF1 (N119, N18);
or OR4 (N120, N7, N16, N93, N34);
nor NOR4 (N121, N118, N45, N6, N67);
xor XOR2 (N122, N108, N86);
and AND3 (N123, N96, N112, N112);
xor XOR2 (N124, N95, N102);
not NOT1 (N125, N123);
or OR3 (N126, N121, N83, N87);
xor XOR2 (N127, N124, N114);
or OR2 (N128, N4, N79);
or OR4 (N129, N122, N77, N62, N95);
nor NOR2 (N130, N126, N112);
nand NAND2 (N131, N117, N95);
and AND3 (N132, N110, N54, N90);
buf BUF1 (N133, N115);
buf BUF1 (N134, N131);
and AND2 (N135, N125, N37);
or OR3 (N136, N134, N124, N82);
not NOT1 (N137, N136);
not NOT1 (N138, N137);
and AND3 (N139, N119, N101, N47);
nand NAND4 (N140, N139, N79, N2, N6);
or OR4 (N141, N135, N111, N71, N41);
or OR3 (N142, N138, N87, N32);
nand NAND3 (N143, N129, N134, N76);
or OR3 (N144, N130, N100, N137);
buf BUF1 (N145, N140);
xor XOR2 (N146, N120, N31);
xor XOR2 (N147, N141, N63);
and AND4 (N148, N133, N87, N71, N38);
or OR3 (N149, N148, N141, N29);
xor XOR2 (N150, N147, N146);
not NOT1 (N151, N128);
not NOT1 (N152, N115);
not NOT1 (N153, N132);
nand NAND3 (N154, N145, N122, N92);
not NOT1 (N155, N154);
nand NAND4 (N156, N151, N58, N102, N140);
and AND3 (N157, N152, N17, N155);
nand NAND3 (N158, N19, N53, N9);
and AND4 (N159, N127, N100, N14, N41);
nand NAND3 (N160, N143, N1, N74);
or OR3 (N161, N157, N79, N39);
nand NAND4 (N162, N149, N77, N133, N152);
not NOT1 (N163, N153);
buf BUF1 (N164, N161);
xor XOR2 (N165, N158, N94);
not NOT1 (N166, N159);
not NOT1 (N167, N162);
not NOT1 (N168, N142);
and AND4 (N169, N144, N40, N136, N73);
nor NOR3 (N170, N156, N130, N94);
xor XOR2 (N171, N166, N63);
and AND3 (N172, N163, N148, N123);
xor XOR2 (N173, N160, N39);
nor NOR4 (N174, N170, N56, N160, N22);
buf BUF1 (N175, N164);
and AND3 (N176, N150, N173, N71);
nor NOR3 (N177, N2, N32, N47);
xor XOR2 (N178, N168, N164);
and AND2 (N179, N177, N18);
buf BUF1 (N180, N175);
xor XOR2 (N181, N171, N97);
or OR2 (N182, N167, N64);
nand NAND3 (N183, N174, N28, N5);
xor XOR2 (N184, N183, N27);
buf BUF1 (N185, N181);
xor XOR2 (N186, N176, N57);
buf BUF1 (N187, N172);
buf BUF1 (N188, N182);
nand NAND4 (N189, N185, N94, N27, N35);
xor XOR2 (N190, N186, N105);
xor XOR2 (N191, N165, N148);
not NOT1 (N192, N187);
nand NAND2 (N193, N169, N76);
and AND3 (N194, N188, N150, N40);
nand NAND4 (N195, N190, N93, N41, N51);
not NOT1 (N196, N184);
and AND2 (N197, N194, N48);
not NOT1 (N198, N197);
nand NAND2 (N199, N195, N51);
xor XOR2 (N200, N178, N139);
and AND2 (N201, N199, N172);
and AND4 (N202, N189, N42, N131, N76);
buf BUF1 (N203, N196);
not NOT1 (N204, N191);
buf BUF1 (N205, N198);
nor NOR4 (N206, N180, N170, N133, N136);
nand NAND2 (N207, N206, N69);
nor NOR4 (N208, N207, N83, N10, N135);
not NOT1 (N209, N205);
xor XOR2 (N210, N209, N180);
nor NOR4 (N211, N210, N19, N156, N141);
xor XOR2 (N212, N203, N167);
or OR4 (N213, N192, N120, N114, N193);
or OR4 (N214, N136, N87, N209, N4);
not NOT1 (N215, N201);
nor NOR3 (N216, N211, N205, N166);
not NOT1 (N217, N202);
not NOT1 (N218, N215);
or OR4 (N219, N218, N63, N210, N196);
not NOT1 (N220, N213);
not NOT1 (N221, N200);
buf BUF1 (N222, N221);
or OR2 (N223, N220, N52);
nor NOR3 (N224, N219, N67, N169);
nor NOR2 (N225, N204, N91);
or OR3 (N226, N223, N156, N148);
or OR3 (N227, N212, N141, N10);
xor XOR2 (N228, N179, N2);
nor NOR3 (N229, N224, N91, N205);
not NOT1 (N230, N226);
buf BUF1 (N231, N225);
not NOT1 (N232, N229);
not NOT1 (N233, N227);
nor NOR3 (N234, N222, N201, N190);
xor XOR2 (N235, N234, N191);
buf BUF1 (N236, N214);
nand NAND2 (N237, N217, N109);
xor XOR2 (N238, N235, N27);
nor NOR2 (N239, N230, N182);
nand NAND2 (N240, N239, N147);
and AND4 (N241, N228, N230, N54, N240);
xor XOR2 (N242, N112, N145);
buf BUF1 (N243, N236);
buf BUF1 (N244, N241);
or OR3 (N245, N208, N201, N182);
and AND4 (N246, N232, N65, N194, N186);
nand NAND3 (N247, N245, N230, N62);
xor XOR2 (N248, N233, N130);
nor NOR4 (N249, N237, N166, N62, N216);
or OR2 (N250, N49, N235);
xor XOR2 (N251, N242, N219);
nor NOR2 (N252, N250, N230);
nand NAND2 (N253, N238, N165);
buf BUF1 (N254, N246);
nor NOR3 (N255, N247, N37, N169);
nand NAND4 (N256, N252, N101, N120, N51);
not NOT1 (N257, N244);
or OR3 (N258, N231, N30, N227);
nand NAND4 (N259, N258, N20, N77, N58);
nor NOR4 (N260, N255, N196, N175, N162);
and AND3 (N261, N257, N31, N77);
buf BUF1 (N262, N243);
nor NOR4 (N263, N259, N11, N73, N19);
not NOT1 (N264, N249);
nand NAND3 (N265, N264, N251, N122);
buf BUF1 (N266, N238);
nor NOR3 (N267, N261, N10, N69);
nor NOR2 (N268, N262, N52);
not NOT1 (N269, N253);
or OR3 (N270, N265, N205, N127);
and AND4 (N271, N254, N247, N240, N114);
buf BUF1 (N272, N271);
and AND3 (N273, N248, N181, N261);
nor NOR4 (N274, N266, N236, N103, N8);
buf BUF1 (N275, N267);
and AND3 (N276, N270, N144, N127);
and AND4 (N277, N273, N165, N38, N11);
not NOT1 (N278, N263);
and AND3 (N279, N256, N267, N260);
or OR2 (N280, N44, N242);
or OR4 (N281, N268, N132, N46, N82);
nand NAND4 (N282, N274, N150, N139, N173);
nand NAND3 (N283, N275, N176, N112);
and AND4 (N284, N278, N179, N35, N269);
xor XOR2 (N285, N27, N148);
buf BUF1 (N286, N285);
or OR3 (N287, N277, N145, N192);
nand NAND4 (N288, N287, N238, N184, N171);
buf BUF1 (N289, N272);
or OR2 (N290, N282, N154);
and AND3 (N291, N286, N162, N41);
xor XOR2 (N292, N290, N231);
and AND2 (N293, N292, N92);
not NOT1 (N294, N283);
and AND4 (N295, N279, N41, N237, N172);
buf BUF1 (N296, N281);
nor NOR3 (N297, N294, N104, N134);
nor NOR3 (N298, N293, N84, N235);
buf BUF1 (N299, N284);
and AND3 (N300, N289, N19, N32);
buf BUF1 (N301, N299);
nand NAND2 (N302, N300, N194);
buf BUF1 (N303, N302);
xor XOR2 (N304, N303, N163);
nand NAND4 (N305, N297, N284, N8, N238);
nand NAND2 (N306, N291, N211);
not NOT1 (N307, N296);
buf BUF1 (N308, N301);
xor XOR2 (N309, N298, N122);
nor NOR2 (N310, N307, N126);
and AND2 (N311, N309, N250);
xor XOR2 (N312, N288, N175);
and AND4 (N313, N276, N39, N302, N118);
and AND2 (N314, N311, N36);
nor NOR4 (N315, N308, N202, N174, N92);
nor NOR2 (N316, N295, N126);
buf BUF1 (N317, N316);
buf BUF1 (N318, N315);
buf BUF1 (N319, N318);
not NOT1 (N320, N319);
or OR3 (N321, N305, N62, N249);
not NOT1 (N322, N310);
nand NAND4 (N323, N306, N308, N30, N253);
not NOT1 (N324, N314);
not NOT1 (N325, N321);
nor NOR3 (N326, N324, N306, N53);
xor XOR2 (N327, N322, N256);
or OR3 (N328, N325, N290, N113);
nor NOR2 (N329, N312, N174);
not NOT1 (N330, N304);
or OR3 (N331, N317, N32, N325);
xor XOR2 (N332, N326, N277);
nand NAND4 (N333, N280, N31, N237, N182);
buf BUF1 (N334, N313);
nor NOR4 (N335, N332, N245, N275, N246);
nor NOR2 (N336, N323, N177);
nor NOR2 (N337, N330, N29);
buf BUF1 (N338, N328);
not NOT1 (N339, N335);
or OR4 (N340, N336, N193, N261, N166);
buf BUF1 (N341, N334);
nand NAND2 (N342, N333, N316);
not NOT1 (N343, N340);
or OR4 (N344, N338, N324, N94, N224);
not NOT1 (N345, N320);
and AND3 (N346, N337, N242, N67);
or OR3 (N347, N341, N120, N306);
and AND3 (N348, N344, N225, N224);
not NOT1 (N349, N327);
and AND3 (N350, N331, N249, N290);
buf BUF1 (N351, N349);
and AND3 (N352, N343, N248, N294);
and AND4 (N353, N351, N346, N344, N184);
and AND3 (N354, N211, N246, N189);
xor XOR2 (N355, N339, N318);
not NOT1 (N356, N345);
nand NAND4 (N357, N353, N130, N209, N133);
xor XOR2 (N358, N357, N187);
xor XOR2 (N359, N347, N167);
xor XOR2 (N360, N329, N165);
nand NAND4 (N361, N348, N14, N302, N328);
nand NAND2 (N362, N356, N159);
xor XOR2 (N363, N355, N102);
nor NOR3 (N364, N362, N242, N310);
not NOT1 (N365, N361);
or OR2 (N366, N358, N98);
not NOT1 (N367, N359);
nor NOR2 (N368, N364, N313);
buf BUF1 (N369, N367);
buf BUF1 (N370, N352);
buf BUF1 (N371, N342);
nor NOR2 (N372, N368, N275);
not NOT1 (N373, N354);
not NOT1 (N374, N371);
xor XOR2 (N375, N350, N189);
or OR4 (N376, N370, N78, N89, N345);
not NOT1 (N377, N372);
nand NAND2 (N378, N374, N236);
and AND3 (N379, N369, N199, N339);
nand NAND2 (N380, N377, N305);
xor XOR2 (N381, N375, N355);
not NOT1 (N382, N365);
not NOT1 (N383, N366);
buf BUF1 (N384, N373);
not NOT1 (N385, N363);
nand NAND4 (N386, N383, N216, N253, N313);
buf BUF1 (N387, N384);
or OR2 (N388, N360, N35);
and AND2 (N389, N382, N152);
buf BUF1 (N390, N376);
or OR2 (N391, N381, N212);
buf BUF1 (N392, N379);
xor XOR2 (N393, N392, N114);
nand NAND4 (N394, N391, N54, N280, N184);
nand NAND2 (N395, N394, N195);
not NOT1 (N396, N395);
xor XOR2 (N397, N386, N64);
xor XOR2 (N398, N393, N282);
and AND3 (N399, N387, N21, N52);
xor XOR2 (N400, N396, N134);
nor NOR4 (N401, N400, N338, N129, N211);
buf BUF1 (N402, N399);
or OR2 (N403, N385, N6);
or OR2 (N404, N402, N121);
or OR2 (N405, N403, N88);
nand NAND2 (N406, N389, N31);
nand NAND2 (N407, N390, N389);
not NOT1 (N408, N388);
xor XOR2 (N409, N397, N163);
nor NOR3 (N410, N380, N279, N352);
not NOT1 (N411, N407);
nor NOR4 (N412, N404, N284, N239, N184);
nand NAND4 (N413, N410, N189, N205, N386);
nand NAND4 (N414, N378, N36, N44, N211);
nand NAND2 (N415, N411, N106);
and AND2 (N416, N413, N280);
xor XOR2 (N417, N409, N380);
and AND4 (N418, N414, N313, N240, N376);
or OR4 (N419, N417, N324, N6, N58);
or OR4 (N420, N408, N143, N242, N118);
and AND2 (N421, N420, N182);
nor NOR3 (N422, N401, N415, N58);
not NOT1 (N423, N104);
not NOT1 (N424, N412);
nor NOR2 (N425, N418, N390);
and AND4 (N426, N421, N70, N347, N163);
or OR4 (N427, N425, N337, N298, N183);
nor NOR2 (N428, N424, N358);
xor XOR2 (N429, N405, N90);
nand NAND3 (N430, N406, N39, N281);
nor NOR3 (N431, N422, N119, N359);
buf BUF1 (N432, N419);
buf BUF1 (N433, N429);
and AND4 (N434, N432, N223, N217, N329);
nand NAND3 (N435, N433, N377, N203);
or OR3 (N436, N431, N149, N50);
and AND2 (N437, N423, N101);
and AND4 (N438, N437, N51, N141, N391);
xor XOR2 (N439, N426, N127);
xor XOR2 (N440, N416, N113);
buf BUF1 (N441, N438);
not NOT1 (N442, N427);
xor XOR2 (N443, N441, N368);
not NOT1 (N444, N442);
nand NAND3 (N445, N444, N234, N315);
nor NOR3 (N446, N430, N195, N349);
and AND4 (N447, N440, N239, N22, N374);
or OR2 (N448, N443, N392);
and AND3 (N449, N398, N63, N137);
not NOT1 (N450, N435);
buf BUF1 (N451, N448);
or OR2 (N452, N434, N292);
and AND3 (N453, N436, N64, N231);
nor NOR2 (N454, N453, N449);
and AND3 (N455, N201, N321, N141);
nand NAND4 (N456, N447, N343, N358, N318);
and AND2 (N457, N439, N346);
nand NAND4 (N458, N451, N114, N33, N316);
not NOT1 (N459, N450);
and AND3 (N460, N459, N383, N328);
and AND3 (N461, N455, N344, N382);
nand NAND4 (N462, N452, N459, N93, N245);
not NOT1 (N463, N462);
nor NOR4 (N464, N463, N127, N206, N263);
nor NOR3 (N465, N461, N126, N307);
xor XOR2 (N466, N460, N63);
xor XOR2 (N467, N457, N284);
or OR4 (N468, N454, N187, N135, N108);
xor XOR2 (N469, N428, N427);
buf BUF1 (N470, N467);
and AND4 (N471, N458, N167, N35, N454);
nand NAND4 (N472, N456, N371, N246, N154);
xor XOR2 (N473, N446, N109);
and AND3 (N474, N464, N255, N251);
and AND2 (N475, N473, N295);
not NOT1 (N476, N445);
buf BUF1 (N477, N470);
xor XOR2 (N478, N471, N280);
buf BUF1 (N479, N466);
buf BUF1 (N480, N476);
xor XOR2 (N481, N468, N161);
buf BUF1 (N482, N465);
xor XOR2 (N483, N472, N121);
or OR4 (N484, N482, N73, N475, N353);
buf BUF1 (N485, N402);
buf BUF1 (N486, N485);
xor XOR2 (N487, N469, N21);
nand NAND3 (N488, N483, N306, N207);
nor NOR4 (N489, N477, N382, N257, N28);
xor XOR2 (N490, N479, N457);
nor NOR2 (N491, N488, N444);
xor XOR2 (N492, N481, N269);
nand NAND3 (N493, N491, N158, N43);
and AND4 (N494, N487, N55, N398, N31);
xor XOR2 (N495, N493, N421);
and AND3 (N496, N486, N292, N281);
buf BUF1 (N497, N478);
xor XOR2 (N498, N489, N196);
xor XOR2 (N499, N492, N321);
not NOT1 (N500, N497);
not NOT1 (N501, N494);
not NOT1 (N502, N501);
buf BUF1 (N503, N500);
or OR2 (N504, N499, N188);
nor NOR2 (N505, N504, N236);
nor NOR4 (N506, N505, N395, N216, N44);
and AND4 (N507, N498, N292, N254, N349);
nand NAND3 (N508, N495, N108, N258);
not NOT1 (N509, N503);
not NOT1 (N510, N502);
and AND4 (N511, N484, N311, N340, N51);
nor NOR4 (N512, N480, N180, N213, N282);
nor NOR4 (N513, N512, N72, N446, N314);
xor XOR2 (N514, N507, N2);
and AND2 (N515, N511, N257);
nor NOR3 (N516, N506, N5, N225);
xor XOR2 (N517, N516, N75);
or OR3 (N518, N514, N88, N42);
not NOT1 (N519, N513);
not NOT1 (N520, N496);
not NOT1 (N521, N490);
buf BUF1 (N522, N517);
xor XOR2 (N523, N515, N355);
or OR2 (N524, N522, N217);
not NOT1 (N525, N524);
buf BUF1 (N526, N521);
nor NOR2 (N527, N510, N476);
and AND4 (N528, N518, N26, N91, N460);
and AND3 (N529, N520, N20, N184);
buf BUF1 (N530, N529);
or OR3 (N531, N525, N264, N235);
not NOT1 (N532, N508);
nor NOR3 (N533, N474, N74, N386);
buf BUF1 (N534, N523);
or OR2 (N535, N528, N187);
and AND2 (N536, N531, N240);
or OR4 (N537, N533, N128, N2, N345);
xor XOR2 (N538, N537, N80);
and AND4 (N539, N532, N496, N291, N527);
nand NAND2 (N540, N417, N202);
buf BUF1 (N541, N539);
not NOT1 (N542, N535);
nand NAND3 (N543, N519, N510, N419);
and AND3 (N544, N538, N382, N297);
nand NAND3 (N545, N536, N302, N434);
or OR4 (N546, N545, N198, N294, N154);
nand NAND2 (N547, N540, N137);
not NOT1 (N548, N547);
or OR2 (N549, N548, N68);
nor NOR4 (N550, N541, N311, N227, N183);
nand NAND4 (N551, N542, N522, N449, N276);
nor NOR3 (N552, N551, N128, N508);
nor NOR4 (N553, N526, N404, N327, N188);
nor NOR4 (N554, N530, N175, N399, N418);
not NOT1 (N555, N546);
nor NOR4 (N556, N544, N175, N56, N525);
not NOT1 (N557, N534);
and AND3 (N558, N554, N296, N163);
nor NOR4 (N559, N557, N82, N172, N302);
and AND4 (N560, N543, N91, N479, N146);
nor NOR3 (N561, N556, N173, N87);
nand NAND2 (N562, N555, N400);
or OR2 (N563, N562, N553);
and AND2 (N564, N28, N154);
nor NOR4 (N565, N559, N121, N413, N474);
and AND3 (N566, N552, N411, N27);
nand NAND3 (N567, N561, N428, N220);
and AND3 (N568, N550, N24, N145);
nand NAND4 (N569, N564, N3, N234, N220);
or OR4 (N570, N568, N19, N485, N429);
nand NAND2 (N571, N563, N204);
and AND4 (N572, N560, N122, N125, N415);
nor NOR2 (N573, N549, N134);
xor XOR2 (N574, N509, N172);
and AND4 (N575, N569, N108, N244, N80);
nor NOR2 (N576, N566, N534);
nor NOR4 (N577, N573, N42, N575, N321);
or OR4 (N578, N336, N535, N23, N244);
xor XOR2 (N579, N571, N407);
nor NOR3 (N580, N558, N530, N552);
or OR4 (N581, N577, N438, N1, N521);
nor NOR3 (N582, N574, N501, N102);
not NOT1 (N583, N576);
buf BUF1 (N584, N565);
and AND4 (N585, N579, N229, N9, N562);
not NOT1 (N586, N572);
not NOT1 (N587, N584);
xor XOR2 (N588, N586, N539);
nor NOR4 (N589, N588, N440, N6, N417);
and AND4 (N590, N578, N3, N525, N368);
nor NOR4 (N591, N587, N250, N403, N441);
nand NAND3 (N592, N590, N177, N418);
buf BUF1 (N593, N580);
and AND3 (N594, N582, N26, N541);
nor NOR4 (N595, N592, N297, N160, N34);
nor NOR3 (N596, N581, N393, N574);
not NOT1 (N597, N596);
or OR4 (N598, N593, N373, N447, N194);
buf BUF1 (N599, N570);
buf BUF1 (N600, N595);
or OR4 (N601, N583, N600, N64, N347);
not NOT1 (N602, N431);
not NOT1 (N603, N567);
or OR4 (N604, N597, N446, N41, N418);
not NOT1 (N605, N601);
xor XOR2 (N606, N594, N344);
not NOT1 (N607, N605);
and AND4 (N608, N599, N80, N522, N115);
not NOT1 (N609, N598);
not NOT1 (N610, N604);
nand NAND2 (N611, N602, N542);
not NOT1 (N612, N606);
nor NOR4 (N613, N611, N402, N446, N244);
not NOT1 (N614, N589);
nor NOR4 (N615, N603, N87, N333, N325);
or OR2 (N616, N609, N404);
buf BUF1 (N617, N612);
or OR4 (N618, N617, N144, N219, N117);
nand NAND3 (N619, N615, N498, N131);
xor XOR2 (N620, N608, N336);
not NOT1 (N621, N614);
nor NOR2 (N622, N610, N402);
not NOT1 (N623, N591);
nand NAND4 (N624, N613, N607, N260, N137);
nand NAND4 (N625, N490, N263, N536, N378);
nand NAND2 (N626, N624, N402);
xor XOR2 (N627, N585, N570);
xor XOR2 (N628, N621, N290);
xor XOR2 (N629, N628, N487);
nor NOR4 (N630, N618, N588, N127, N258);
or OR2 (N631, N630, N561);
and AND4 (N632, N619, N404, N446, N542);
nand NAND3 (N633, N620, N94, N583);
nor NOR3 (N634, N633, N85, N73);
xor XOR2 (N635, N623, N360);
buf BUF1 (N636, N627);
nand NAND3 (N637, N616, N561, N138);
or OR3 (N638, N635, N278, N372);
xor XOR2 (N639, N625, N346);
not NOT1 (N640, N636);
and AND2 (N641, N639, N519);
nor NOR2 (N642, N629, N195);
xor XOR2 (N643, N641, N61);
nor NOR2 (N644, N637, N317);
and AND4 (N645, N634, N596, N161, N234);
buf BUF1 (N646, N644);
nand NAND2 (N647, N626, N181);
xor XOR2 (N648, N632, N549);
buf BUF1 (N649, N648);
buf BUF1 (N650, N638);
nor NOR2 (N651, N640, N215);
nor NOR4 (N652, N650, N285, N167, N557);
and AND2 (N653, N643, N590);
and AND3 (N654, N649, N505, N516);
and AND4 (N655, N653, N42, N4, N577);
xor XOR2 (N656, N655, N451);
or OR4 (N657, N656, N278, N646, N33);
not NOT1 (N658, N309);
and AND4 (N659, N647, N546, N442, N106);
nor NOR3 (N660, N654, N392, N160);
nor NOR3 (N661, N631, N533, N639);
buf BUF1 (N662, N645);
or OR2 (N663, N660, N528);
and AND4 (N664, N663, N6, N365, N502);
and AND3 (N665, N652, N655, N20);
not NOT1 (N666, N665);
nor NOR3 (N667, N662, N314, N44);
nor NOR2 (N668, N658, N334);
nand NAND2 (N669, N622, N541);
not NOT1 (N670, N659);
xor XOR2 (N671, N666, N362);
and AND2 (N672, N668, N368);
not NOT1 (N673, N657);
not NOT1 (N674, N661);
nand NAND2 (N675, N669, N224);
nor NOR3 (N676, N642, N385, N384);
or OR4 (N677, N674, N351, N220, N673);
nand NAND3 (N678, N169, N426, N546);
buf BUF1 (N679, N651);
not NOT1 (N680, N672);
xor XOR2 (N681, N676, N268);
or OR4 (N682, N675, N342, N395, N668);
nand NAND2 (N683, N679, N347);
xor XOR2 (N684, N682, N499);
nand NAND2 (N685, N684, N639);
nand NAND3 (N686, N683, N535, N516);
or OR4 (N687, N664, N547, N43, N364);
buf BUF1 (N688, N670);
or OR3 (N689, N686, N411, N355);
not NOT1 (N690, N667);
nand NAND4 (N691, N687, N292, N244, N365);
not NOT1 (N692, N691);
and AND3 (N693, N678, N573, N339);
buf BUF1 (N694, N671);
nor NOR3 (N695, N690, N63, N636);
or OR2 (N696, N692, N319);
buf BUF1 (N697, N677);
nand NAND4 (N698, N694, N225, N563, N353);
or OR3 (N699, N681, N51, N54);
xor XOR2 (N700, N696, N384);
and AND3 (N701, N695, N91, N596);
or OR3 (N702, N697, N394, N343);
not NOT1 (N703, N689);
xor XOR2 (N704, N702, N5);
nand NAND4 (N705, N699, N193, N573, N621);
or OR2 (N706, N685, N689);
buf BUF1 (N707, N701);
nand NAND4 (N708, N703, N668, N652, N231);
not NOT1 (N709, N704);
nor NOR4 (N710, N705, N254, N187, N377);
buf BUF1 (N711, N707);
nand NAND2 (N712, N709, N312);
and AND3 (N713, N708, N253, N572);
xor XOR2 (N714, N711, N192);
not NOT1 (N715, N713);
and AND3 (N716, N710, N10, N250);
nand NAND2 (N717, N715, N127);
or OR4 (N718, N693, N248, N58, N180);
not NOT1 (N719, N700);
buf BUF1 (N720, N712);
or OR3 (N721, N698, N635, N440);
or OR3 (N722, N718, N89, N676);
xor XOR2 (N723, N680, N89);
and AND4 (N724, N723, N153, N617, N314);
buf BUF1 (N725, N717);
and AND4 (N726, N721, N613, N635, N400);
nor NOR2 (N727, N720, N72);
not NOT1 (N728, N714);
nand NAND2 (N729, N726, N588);
and AND2 (N730, N728, N725);
xor XOR2 (N731, N623, N189);
nand NAND2 (N732, N688, N377);
xor XOR2 (N733, N706, N434);
xor XOR2 (N734, N731, N239);
not NOT1 (N735, N722);
buf BUF1 (N736, N729);
xor XOR2 (N737, N733, N116);
and AND4 (N738, N736, N198, N80, N270);
nor NOR2 (N739, N735, N124);
and AND4 (N740, N724, N529, N233, N259);
buf BUF1 (N741, N740);
buf BUF1 (N742, N734);
xor XOR2 (N743, N727, N19);
xor XOR2 (N744, N716, N20);
nand NAND2 (N745, N739, N186);
nand NAND2 (N746, N742, N533);
and AND2 (N747, N745, N403);
and AND2 (N748, N732, N417);
nand NAND2 (N749, N719, N190);
xor XOR2 (N750, N743, N505);
and AND3 (N751, N744, N172, N187);
xor XOR2 (N752, N738, N710);
buf BUF1 (N753, N747);
xor XOR2 (N754, N749, N305);
not NOT1 (N755, N752);
and AND3 (N756, N741, N391, N317);
or OR2 (N757, N755, N334);
not NOT1 (N758, N750);
nor NOR2 (N759, N737, N64);
xor XOR2 (N760, N746, N79);
not NOT1 (N761, N730);
buf BUF1 (N762, N760);
nand NAND4 (N763, N756, N500, N171, N649);
or OR3 (N764, N754, N683, N241);
not NOT1 (N765, N759);
not NOT1 (N766, N763);
buf BUF1 (N767, N748);
not NOT1 (N768, N767);
and AND3 (N769, N757, N517, N474);
nor NOR4 (N770, N765, N444, N577, N701);
and AND4 (N771, N761, N116, N174, N178);
nor NOR2 (N772, N766, N581);
and AND2 (N773, N770, N629);
not NOT1 (N774, N773);
xor XOR2 (N775, N762, N581);
not NOT1 (N776, N775);
not NOT1 (N777, N751);
xor XOR2 (N778, N777, N422);
nor NOR3 (N779, N778, N262, N488);
not NOT1 (N780, N769);
not NOT1 (N781, N780);
buf BUF1 (N782, N772);
xor XOR2 (N783, N782, N650);
not NOT1 (N784, N764);
and AND3 (N785, N781, N527, N489);
or OR3 (N786, N768, N361, N133);
xor XOR2 (N787, N753, N225);
not NOT1 (N788, N771);
or OR2 (N789, N774, N352);
and AND3 (N790, N787, N341, N84);
xor XOR2 (N791, N785, N636);
xor XOR2 (N792, N788, N318);
or OR4 (N793, N776, N739, N559, N135);
not NOT1 (N794, N793);
xor XOR2 (N795, N779, N531);
nand NAND3 (N796, N758, N303, N751);
buf BUF1 (N797, N791);
buf BUF1 (N798, N790);
and AND3 (N799, N795, N208, N17);
nand NAND3 (N800, N794, N712, N157);
and AND3 (N801, N796, N186, N349);
nor NOR4 (N802, N783, N309, N358, N516);
xor XOR2 (N803, N792, N133);
nand NAND4 (N804, N797, N113, N252, N305);
buf BUF1 (N805, N798);
xor XOR2 (N806, N803, N699);
not NOT1 (N807, N801);
not NOT1 (N808, N805);
nor NOR4 (N809, N804, N113, N371, N286);
buf BUF1 (N810, N808);
or OR4 (N811, N809, N123, N611, N540);
and AND4 (N812, N810, N534, N278, N467);
not NOT1 (N813, N806);
xor XOR2 (N814, N784, N473);
nand NAND4 (N815, N811, N717, N432, N206);
nand NAND2 (N816, N800, N712);
buf BUF1 (N817, N813);
and AND4 (N818, N807, N691, N499, N328);
buf BUF1 (N819, N815);
not NOT1 (N820, N786);
and AND4 (N821, N799, N337, N302, N626);
nor NOR2 (N822, N819, N212);
not NOT1 (N823, N820);
and AND2 (N824, N818, N187);
or OR2 (N825, N816, N740);
xor XOR2 (N826, N824, N813);
xor XOR2 (N827, N822, N409);
not NOT1 (N828, N825);
or OR2 (N829, N826, N72);
or OR3 (N830, N802, N503, N51);
xor XOR2 (N831, N812, N88);
not NOT1 (N832, N789);
xor XOR2 (N833, N814, N666);
xor XOR2 (N834, N823, N550);
buf BUF1 (N835, N834);
nand NAND4 (N836, N835, N493, N620, N9);
buf BUF1 (N837, N831);
not NOT1 (N838, N837);
nand NAND4 (N839, N827, N312, N628, N810);
or OR3 (N840, N828, N234, N581);
nor NOR4 (N841, N836, N297, N460, N156);
or OR3 (N842, N817, N290, N632);
xor XOR2 (N843, N821, N292);
xor XOR2 (N844, N843, N526);
nand NAND4 (N845, N844, N39, N20, N92);
not NOT1 (N846, N829);
or OR4 (N847, N841, N448, N487, N83);
not NOT1 (N848, N830);
xor XOR2 (N849, N840, N601);
and AND4 (N850, N842, N410, N113, N754);
and AND3 (N851, N832, N793, N351);
or OR4 (N852, N838, N251, N797, N301);
or OR4 (N853, N850, N93, N292, N641);
buf BUF1 (N854, N848);
nor NOR3 (N855, N849, N325, N672);
not NOT1 (N856, N853);
and AND4 (N857, N845, N443, N367, N160);
nor NOR4 (N858, N833, N593, N815, N201);
nand NAND2 (N859, N852, N706);
nor NOR3 (N860, N839, N118, N476);
nor NOR3 (N861, N854, N727, N803);
nand NAND2 (N862, N861, N795);
buf BUF1 (N863, N851);
xor XOR2 (N864, N858, N760);
nand NAND4 (N865, N847, N787, N557, N156);
and AND3 (N866, N864, N203, N653);
nor NOR2 (N867, N846, N390);
and AND3 (N868, N857, N843, N825);
or OR2 (N869, N860, N764);
not NOT1 (N870, N862);
buf BUF1 (N871, N867);
nor NOR3 (N872, N865, N870, N262);
nand NAND4 (N873, N706, N232, N44, N247);
or OR4 (N874, N871, N852, N217, N530);
nor NOR4 (N875, N866, N287, N229, N832);
nand NAND3 (N876, N875, N683, N65);
xor XOR2 (N877, N876, N803);
not NOT1 (N878, N872);
nor NOR4 (N879, N878, N145, N637, N644);
not NOT1 (N880, N856);
not NOT1 (N881, N879);
nor NOR2 (N882, N855, N278);
nand NAND3 (N883, N882, N12, N579);
or OR2 (N884, N877, N243);
buf BUF1 (N885, N873);
nand NAND4 (N886, N874, N481, N192, N299);
not NOT1 (N887, N863);
and AND3 (N888, N884, N372, N784);
not NOT1 (N889, N880);
nor NOR3 (N890, N868, N81, N574);
or OR2 (N891, N890, N38);
buf BUF1 (N892, N869);
nand NAND4 (N893, N885, N509, N432, N888);
nor NOR4 (N894, N76, N147, N343, N26);
not NOT1 (N895, N894);
nand NAND3 (N896, N883, N344, N234);
or OR4 (N897, N892, N34, N37, N150);
nand NAND3 (N898, N895, N92, N553);
or OR4 (N899, N896, N376, N482, N851);
nand NAND2 (N900, N891, N777);
nand NAND4 (N901, N859, N145, N582, N839);
and AND4 (N902, N899, N810, N750, N327);
nor NOR4 (N903, N901, N120, N249, N428);
not NOT1 (N904, N898);
buf BUF1 (N905, N900);
nor NOR3 (N906, N902, N293, N882);
and AND4 (N907, N897, N189, N652, N43);
nor NOR4 (N908, N906, N94, N581, N641);
nand NAND2 (N909, N887, N668);
xor XOR2 (N910, N908, N627);
buf BUF1 (N911, N893);
and AND2 (N912, N903, N857);
xor XOR2 (N913, N904, N694);
nand NAND2 (N914, N910, N660);
xor XOR2 (N915, N914, N645);
not NOT1 (N916, N907);
buf BUF1 (N917, N889);
nand NAND4 (N918, N913, N140, N638, N269);
or OR2 (N919, N917, N898);
nand NAND3 (N920, N909, N529, N118);
nor NOR4 (N921, N912, N176, N287, N1);
nand NAND3 (N922, N916, N540, N64);
buf BUF1 (N923, N881);
buf BUF1 (N924, N915);
and AND3 (N925, N922, N122, N369);
buf BUF1 (N926, N905);
nor NOR4 (N927, N923, N604, N666, N477);
nand NAND4 (N928, N926, N268, N345, N483);
nand NAND4 (N929, N919, N522, N132, N465);
buf BUF1 (N930, N911);
xor XOR2 (N931, N921, N753);
or OR2 (N932, N924, N137);
buf BUF1 (N933, N928);
not NOT1 (N934, N929);
and AND3 (N935, N918, N293, N575);
xor XOR2 (N936, N886, N578);
xor XOR2 (N937, N925, N509);
nor NOR2 (N938, N936, N804);
xor XOR2 (N939, N927, N788);
or OR2 (N940, N931, N665);
and AND4 (N941, N938, N409, N38, N413);
nor NOR2 (N942, N937, N517);
buf BUF1 (N943, N940);
or OR2 (N944, N930, N409);
not NOT1 (N945, N943);
or OR3 (N946, N941, N799, N638);
nand NAND4 (N947, N939, N946, N437, N388);
nor NOR4 (N948, N281, N802, N385, N16);
buf BUF1 (N949, N934);
not NOT1 (N950, N933);
and AND3 (N951, N948, N878, N589);
and AND4 (N952, N944, N760, N392, N71);
buf BUF1 (N953, N951);
not NOT1 (N954, N952);
and AND3 (N955, N920, N26, N615);
not NOT1 (N956, N942);
nand NAND3 (N957, N947, N257, N483);
xor XOR2 (N958, N953, N641);
or OR2 (N959, N935, N255);
buf BUF1 (N960, N945);
buf BUF1 (N961, N960);
not NOT1 (N962, N958);
nand NAND2 (N963, N957, N709);
not NOT1 (N964, N949);
or OR3 (N965, N932, N816, N882);
nor NOR4 (N966, N959, N53, N165, N440);
nand NAND2 (N967, N964, N792);
nand NAND2 (N968, N962, N878);
not NOT1 (N969, N968);
or OR2 (N970, N965, N57);
not NOT1 (N971, N955);
not NOT1 (N972, N961);
nor NOR4 (N973, N970, N224, N460, N279);
or OR3 (N974, N963, N796, N62);
buf BUF1 (N975, N956);
not NOT1 (N976, N954);
not NOT1 (N977, N974);
and AND2 (N978, N966, N962);
and AND2 (N979, N969, N624);
nand NAND2 (N980, N973, N218);
nor NOR2 (N981, N975, N115);
buf BUF1 (N982, N967);
or OR2 (N983, N980, N122);
xor XOR2 (N984, N982, N703);
nand NAND4 (N985, N979, N763, N661, N231);
not NOT1 (N986, N981);
or OR4 (N987, N983, N359, N898, N563);
xor XOR2 (N988, N976, N739);
and AND4 (N989, N977, N533, N712, N981);
and AND4 (N990, N950, N174, N821, N857);
buf BUF1 (N991, N984);
or OR4 (N992, N988, N366, N921, N470);
and AND4 (N993, N971, N12, N163, N260);
xor XOR2 (N994, N985, N973);
xor XOR2 (N995, N972, N37);
and AND2 (N996, N995, N117);
nor NOR3 (N997, N987, N884, N552);
and AND3 (N998, N990, N741, N600);
not NOT1 (N999, N986);
or OR2 (N1000, N999, N713);
nor NOR4 (N1001, N997, N346, N785, N929);
buf BUF1 (N1002, N998);
not NOT1 (N1003, N993);
xor XOR2 (N1004, N978, N35);
not NOT1 (N1005, N1002);
and AND3 (N1006, N994, N728, N980);
not NOT1 (N1007, N1005);
not NOT1 (N1008, N1006);
nand NAND4 (N1009, N992, N98, N680, N175);
and AND3 (N1010, N1004, N367, N63);
nor NOR2 (N1011, N989, N921);
buf BUF1 (N1012, N1008);
buf BUF1 (N1013, N1003);
xor XOR2 (N1014, N1000, N455);
nand NAND2 (N1015, N1007, N131);
not NOT1 (N1016, N1009);
not NOT1 (N1017, N996);
nor NOR2 (N1018, N991, N777);
buf BUF1 (N1019, N1016);
nand NAND2 (N1020, N1013, N137);
nor NOR2 (N1021, N1019, N50);
not NOT1 (N1022, N1012);
and AND3 (N1023, N1018, N663, N635);
xor XOR2 (N1024, N1022, N180);
and AND3 (N1025, N1017, N632, N403);
nor NOR4 (N1026, N1021, N271, N579, N384);
and AND4 (N1027, N1023, N556, N649, N745);
nor NOR3 (N1028, N1026, N577, N549);
xor XOR2 (N1029, N1028, N695);
nor NOR3 (N1030, N1029, N403, N424);
not NOT1 (N1031, N1020);
or OR3 (N1032, N1010, N627, N379);
xor XOR2 (N1033, N1025, N745);
nand NAND4 (N1034, N1014, N1002, N439, N283);
nor NOR4 (N1035, N1015, N282, N697, N351);
and AND3 (N1036, N1033, N331, N22);
nor NOR4 (N1037, N1035, N863, N745, N734);
buf BUF1 (N1038, N1011);
xor XOR2 (N1039, N1034, N330);
or OR4 (N1040, N1032, N79, N84, N590);
xor XOR2 (N1041, N1030, N743);
xor XOR2 (N1042, N1027, N725);
not NOT1 (N1043, N1001);
not NOT1 (N1044, N1037);
buf BUF1 (N1045, N1044);
not NOT1 (N1046, N1024);
nand NAND2 (N1047, N1036, N934);
or OR3 (N1048, N1042, N325, N435);
nand NAND3 (N1049, N1038, N839, N251);
and AND2 (N1050, N1031, N307);
nand NAND3 (N1051, N1040, N635, N702);
xor XOR2 (N1052, N1049, N299);
not NOT1 (N1053, N1048);
not NOT1 (N1054, N1045);
and AND4 (N1055, N1047, N851, N714, N197);
buf BUF1 (N1056, N1055);
nand NAND4 (N1057, N1046, N754, N604, N831);
nor NOR3 (N1058, N1053, N980, N975);
nor NOR2 (N1059, N1056, N136);
xor XOR2 (N1060, N1058, N6);
or OR2 (N1061, N1052, N528);
and AND2 (N1062, N1050, N530);
not NOT1 (N1063, N1057);
buf BUF1 (N1064, N1039);
nor NOR3 (N1065, N1041, N251, N2);
xor XOR2 (N1066, N1061, N636);
and AND4 (N1067, N1066, N596, N235, N116);
and AND3 (N1068, N1063, N45, N503);
nand NAND2 (N1069, N1054, N407);
not NOT1 (N1070, N1068);
xor XOR2 (N1071, N1070, N438);
nand NAND2 (N1072, N1064, N906);
buf BUF1 (N1073, N1069);
nor NOR4 (N1074, N1043, N569, N56, N428);
xor XOR2 (N1075, N1071, N332);
or OR3 (N1076, N1060, N593, N682);
nand NAND3 (N1077, N1073, N453, N843);
or OR3 (N1078, N1072, N768, N89);
nor NOR4 (N1079, N1065, N142, N748, N3);
not NOT1 (N1080, N1078);
nor NOR3 (N1081, N1080, N372, N288);
not NOT1 (N1082, N1062);
xor XOR2 (N1083, N1051, N949);
not NOT1 (N1084, N1074);
buf BUF1 (N1085, N1081);
xor XOR2 (N1086, N1059, N144);
or OR4 (N1087, N1079, N205, N413, N444);
xor XOR2 (N1088, N1076, N962);
nand NAND4 (N1089, N1087, N6, N460, N863);
and AND3 (N1090, N1086, N661, N1064);
or OR3 (N1091, N1077, N336, N1089);
nand NAND2 (N1092, N807, N914);
buf BUF1 (N1093, N1084);
or OR4 (N1094, N1085, N658, N286, N950);
or OR4 (N1095, N1082, N451, N1032, N444);
nand NAND3 (N1096, N1083, N615, N94);
buf BUF1 (N1097, N1093);
nor NOR3 (N1098, N1096, N436, N329);
not NOT1 (N1099, N1092);
and AND4 (N1100, N1075, N508, N995, N352);
or OR2 (N1101, N1094, N794);
or OR2 (N1102, N1067, N260);
nor NOR4 (N1103, N1102, N220, N172, N248);
nand NAND4 (N1104, N1099, N492, N426, N341);
or OR4 (N1105, N1095, N1028, N886, N1023);
xor XOR2 (N1106, N1100, N836);
nand NAND3 (N1107, N1097, N115, N451);
nor NOR2 (N1108, N1088, N637);
or OR2 (N1109, N1106, N227);
xor XOR2 (N1110, N1101, N464);
and AND2 (N1111, N1090, N388);
not NOT1 (N1112, N1103);
nand NAND3 (N1113, N1111, N837, N541);
and AND2 (N1114, N1107, N733);
nor NOR2 (N1115, N1114, N321);
nand NAND2 (N1116, N1091, N457);
nor NOR3 (N1117, N1116, N355, N527);
not NOT1 (N1118, N1105);
buf BUF1 (N1119, N1098);
or OR2 (N1120, N1119, N643);
xor XOR2 (N1121, N1117, N503);
buf BUF1 (N1122, N1108);
and AND4 (N1123, N1118, N125, N816, N733);
not NOT1 (N1124, N1120);
nor NOR3 (N1125, N1109, N511, N1105);
nand NAND4 (N1126, N1123, N105, N863, N747);
xor XOR2 (N1127, N1104, N855);
xor XOR2 (N1128, N1115, N365);
and AND3 (N1129, N1126, N662, N74);
and AND3 (N1130, N1112, N985, N1006);
not NOT1 (N1131, N1124);
and AND4 (N1132, N1131, N1076, N725, N565);
xor XOR2 (N1133, N1122, N724);
or OR3 (N1134, N1121, N485, N1061);
nand NAND2 (N1135, N1125, N299);
nor NOR4 (N1136, N1127, N190, N1028, N449);
xor XOR2 (N1137, N1130, N877);
nand NAND2 (N1138, N1129, N510);
xor XOR2 (N1139, N1113, N421);
nor NOR2 (N1140, N1110, N827);
xor XOR2 (N1141, N1140, N746);
xor XOR2 (N1142, N1141, N1015);
xor XOR2 (N1143, N1134, N310);
nand NAND3 (N1144, N1143, N200, N209);
buf BUF1 (N1145, N1135);
nor NOR2 (N1146, N1137, N442);
nand NAND3 (N1147, N1136, N206, N835);
not NOT1 (N1148, N1138);
or OR2 (N1149, N1148, N466);
and AND3 (N1150, N1146, N315, N289);
xor XOR2 (N1151, N1139, N329);
and AND3 (N1152, N1142, N951, N1006);
nand NAND4 (N1153, N1145, N141, N365, N58);
buf BUF1 (N1154, N1152);
or OR4 (N1155, N1149, N861, N958, N264);
nor NOR3 (N1156, N1155, N537, N692);
nand NAND2 (N1157, N1153, N903);
xor XOR2 (N1158, N1147, N391);
nand NAND3 (N1159, N1156, N322, N520);
not NOT1 (N1160, N1133);
buf BUF1 (N1161, N1132);
not NOT1 (N1162, N1157);
not NOT1 (N1163, N1128);
nor NOR2 (N1164, N1159, N333);
nor NOR2 (N1165, N1162, N279);
nand NAND3 (N1166, N1160, N569, N365);
xor XOR2 (N1167, N1144, N227);
xor XOR2 (N1168, N1154, N496);
not NOT1 (N1169, N1163);
nand NAND3 (N1170, N1166, N397, N1037);
not NOT1 (N1171, N1170);
xor XOR2 (N1172, N1169, N799);
and AND2 (N1173, N1151, N701);
not NOT1 (N1174, N1158);
buf BUF1 (N1175, N1168);
not NOT1 (N1176, N1150);
nor NOR2 (N1177, N1173, N685);
nand NAND3 (N1178, N1175, N791, N472);
buf BUF1 (N1179, N1177);
and AND2 (N1180, N1167, N84);
buf BUF1 (N1181, N1164);
and AND4 (N1182, N1171, N49, N19, N242);
and AND4 (N1183, N1178, N641, N161, N923);
xor XOR2 (N1184, N1183, N1123);
and AND3 (N1185, N1181, N1044, N110);
not NOT1 (N1186, N1184);
not NOT1 (N1187, N1174);
xor XOR2 (N1188, N1172, N1122);
xor XOR2 (N1189, N1161, N510);
or OR2 (N1190, N1185, N740);
not NOT1 (N1191, N1188);
nand NAND3 (N1192, N1187, N132, N1042);
nand NAND3 (N1193, N1179, N378, N1036);
and AND3 (N1194, N1191, N1071, N701);
xor XOR2 (N1195, N1186, N154);
not NOT1 (N1196, N1180);
xor XOR2 (N1197, N1176, N596);
not NOT1 (N1198, N1195);
and AND3 (N1199, N1190, N1023, N859);
or OR4 (N1200, N1197, N660, N361, N750);
xor XOR2 (N1201, N1194, N1065);
and AND2 (N1202, N1193, N809);
nor NOR3 (N1203, N1165, N833, N235);
nor NOR3 (N1204, N1196, N664, N316);
buf BUF1 (N1205, N1199);
and AND2 (N1206, N1205, N316);
buf BUF1 (N1207, N1198);
not NOT1 (N1208, N1200);
and AND3 (N1209, N1206, N817, N955);
buf BUF1 (N1210, N1182);
buf BUF1 (N1211, N1192);
xor XOR2 (N1212, N1202, N880);
buf BUF1 (N1213, N1210);
xor XOR2 (N1214, N1203, N673);
or OR4 (N1215, N1211, N834, N1038, N966);
and AND4 (N1216, N1213, N762, N68, N586);
buf BUF1 (N1217, N1215);
nand NAND3 (N1218, N1217, N386, N1209);
not NOT1 (N1219, N645);
not NOT1 (N1220, N1207);
nand NAND4 (N1221, N1219, N372, N991, N536);
nor NOR2 (N1222, N1214, N261);
nand NAND4 (N1223, N1204, N971, N973, N76);
not NOT1 (N1224, N1189);
not NOT1 (N1225, N1223);
buf BUF1 (N1226, N1220);
nor NOR4 (N1227, N1218, N836, N79, N580);
nand NAND3 (N1228, N1224, N290, N494);
nor NOR4 (N1229, N1201, N157, N633, N754);
xor XOR2 (N1230, N1221, N336);
nand NAND3 (N1231, N1229, N162, N928);
not NOT1 (N1232, N1212);
nor NOR4 (N1233, N1231, N308, N1086, N146);
xor XOR2 (N1234, N1227, N332);
buf BUF1 (N1235, N1234);
and AND3 (N1236, N1235, N10, N1129);
xor XOR2 (N1237, N1216, N651);
xor XOR2 (N1238, N1236, N934);
or OR3 (N1239, N1222, N918, N1233);
xor XOR2 (N1240, N588, N561);
buf BUF1 (N1241, N1228);
not NOT1 (N1242, N1226);
nor NOR4 (N1243, N1230, N152, N1187, N782);
nand NAND4 (N1244, N1208, N568, N217, N756);
nand NAND4 (N1245, N1243, N1034, N88, N332);
nand NAND2 (N1246, N1242, N179);
or OR2 (N1247, N1238, N417);
or OR2 (N1248, N1244, N141);
nand NAND3 (N1249, N1240, N987, N298);
xor XOR2 (N1250, N1237, N734);
not NOT1 (N1251, N1232);
nor NOR4 (N1252, N1241, N850, N921, N394);
nand NAND4 (N1253, N1252, N579, N512, N254);
not NOT1 (N1254, N1250);
and AND4 (N1255, N1251, N724, N830, N257);
nand NAND2 (N1256, N1254, N859);
buf BUF1 (N1257, N1249);
nand NAND4 (N1258, N1248, N333, N875, N460);
nand NAND3 (N1259, N1245, N54, N557);
nand NAND3 (N1260, N1225, N24, N492);
or OR2 (N1261, N1255, N1199);
not NOT1 (N1262, N1260);
and AND2 (N1263, N1246, N264);
not NOT1 (N1264, N1263);
xor XOR2 (N1265, N1239, N204);
not NOT1 (N1266, N1261);
and AND3 (N1267, N1265, N337, N425);
nor NOR2 (N1268, N1258, N493);
or OR2 (N1269, N1256, N771);
or OR3 (N1270, N1269, N1229, N1084);
or OR2 (N1271, N1268, N782);
not NOT1 (N1272, N1264);
nor NOR3 (N1273, N1271, N197, N865);
nor NOR3 (N1274, N1253, N389, N1231);
buf BUF1 (N1275, N1262);
buf BUF1 (N1276, N1273);
xor XOR2 (N1277, N1259, N82);
or OR2 (N1278, N1266, N196);
and AND4 (N1279, N1276, N1021, N459, N937);
and AND4 (N1280, N1272, N268, N47, N20);
nand NAND2 (N1281, N1274, N184);
or OR3 (N1282, N1275, N603, N202);
nand NAND2 (N1283, N1277, N1254);
and AND2 (N1284, N1257, N1204);
xor XOR2 (N1285, N1282, N1221);
xor XOR2 (N1286, N1281, N7);
buf BUF1 (N1287, N1267);
nor NOR3 (N1288, N1279, N435, N105);
xor XOR2 (N1289, N1280, N360);
not NOT1 (N1290, N1289);
buf BUF1 (N1291, N1270);
or OR3 (N1292, N1291, N727, N638);
nand NAND2 (N1293, N1286, N384);
nand NAND4 (N1294, N1288, N385, N1144, N441);
and AND4 (N1295, N1292, N646, N1139, N777);
nor NOR3 (N1296, N1247, N315, N632);
not NOT1 (N1297, N1295);
not NOT1 (N1298, N1283);
buf BUF1 (N1299, N1278);
not NOT1 (N1300, N1299);
and AND2 (N1301, N1297, N74);
not NOT1 (N1302, N1284);
nor NOR3 (N1303, N1301, N873, N229);
nor NOR3 (N1304, N1296, N1070, N537);
xor XOR2 (N1305, N1293, N245);
or OR4 (N1306, N1300, N1160, N977, N368);
xor XOR2 (N1307, N1305, N731);
or OR3 (N1308, N1302, N1155, N267);
or OR3 (N1309, N1307, N1112, N890);
not NOT1 (N1310, N1304);
and AND2 (N1311, N1303, N1047);
buf BUF1 (N1312, N1290);
nand NAND3 (N1313, N1312, N474, N1095);
buf BUF1 (N1314, N1309);
nor NOR4 (N1315, N1310, N1127, N70, N337);
nor NOR2 (N1316, N1315, N910);
or OR3 (N1317, N1294, N506, N580);
or OR2 (N1318, N1308, N754);
xor XOR2 (N1319, N1306, N1292);
not NOT1 (N1320, N1311);
nor NOR2 (N1321, N1316, N1050);
buf BUF1 (N1322, N1318);
nand NAND2 (N1323, N1319, N1010);
or OR3 (N1324, N1285, N675, N961);
nand NAND4 (N1325, N1324, N155, N506, N945);
not NOT1 (N1326, N1320);
and AND4 (N1327, N1323, N1132, N629, N432);
and AND2 (N1328, N1325, N133);
not NOT1 (N1329, N1321);
not NOT1 (N1330, N1314);
nand NAND3 (N1331, N1313, N1203, N856);
nor NOR4 (N1332, N1328, N1300, N1074, N1144);
or OR2 (N1333, N1287, N658);
and AND3 (N1334, N1331, N1020, N1056);
and AND3 (N1335, N1333, N440, N22);
buf BUF1 (N1336, N1322);
nand NAND3 (N1337, N1335, N13, N1041);
and AND4 (N1338, N1334, N221, N492, N1147);
nand NAND4 (N1339, N1327, N1125, N1002, N1269);
and AND3 (N1340, N1336, N1329, N892);
buf BUF1 (N1341, N336);
nor NOR4 (N1342, N1339, N1281, N1035, N962);
nand NAND3 (N1343, N1337, N803, N421);
buf BUF1 (N1344, N1326);
and AND4 (N1345, N1338, N1121, N797, N905);
not NOT1 (N1346, N1332);
or OR4 (N1347, N1298, N1321, N1087, N122);
nor NOR3 (N1348, N1317, N546, N223);
buf BUF1 (N1349, N1348);
buf BUF1 (N1350, N1343);
buf BUF1 (N1351, N1345);
buf BUF1 (N1352, N1341);
and AND4 (N1353, N1340, N597, N22, N999);
or OR3 (N1354, N1353, N519, N863);
nor NOR2 (N1355, N1342, N745);
nand NAND4 (N1356, N1349, N568, N279, N920);
buf BUF1 (N1357, N1350);
and AND2 (N1358, N1330, N1176);
or OR4 (N1359, N1346, N1236, N1113, N715);
or OR2 (N1360, N1357, N1126);
buf BUF1 (N1361, N1344);
nor NOR2 (N1362, N1358, N121);
nor NOR3 (N1363, N1347, N1259, N811);
not NOT1 (N1364, N1356);
not NOT1 (N1365, N1354);
and AND4 (N1366, N1364, N871, N748, N554);
not NOT1 (N1367, N1359);
buf BUF1 (N1368, N1366);
nand NAND3 (N1369, N1355, N527, N233);
nor NOR2 (N1370, N1362, N117);
buf BUF1 (N1371, N1370);
or OR2 (N1372, N1367, N530);
xor XOR2 (N1373, N1352, N1193);
or OR2 (N1374, N1363, N527);
xor XOR2 (N1375, N1361, N1256);
or OR3 (N1376, N1371, N1241, N1046);
nand NAND3 (N1377, N1351, N239, N1323);
not NOT1 (N1378, N1369);
or OR3 (N1379, N1360, N1049, N278);
or OR2 (N1380, N1365, N372);
xor XOR2 (N1381, N1379, N1034);
xor XOR2 (N1382, N1376, N819);
buf BUF1 (N1383, N1377);
nor NOR4 (N1384, N1382, N269, N1170, N1138);
or OR4 (N1385, N1381, N1195, N325, N1038);
not NOT1 (N1386, N1380);
buf BUF1 (N1387, N1374);
and AND3 (N1388, N1375, N380, N323);
not NOT1 (N1389, N1387);
nor NOR2 (N1390, N1385, N771);
xor XOR2 (N1391, N1368, N1332);
buf BUF1 (N1392, N1384);
not NOT1 (N1393, N1372);
xor XOR2 (N1394, N1378, N1165);
or OR4 (N1395, N1391, N532, N917, N1088);
or OR3 (N1396, N1394, N954, N127);
or OR2 (N1397, N1386, N1336);
and AND3 (N1398, N1393, N21, N1252);
not NOT1 (N1399, N1388);
not NOT1 (N1400, N1395);
or OR3 (N1401, N1400, N684, N1098);
and AND4 (N1402, N1389, N124, N963, N203);
xor XOR2 (N1403, N1402, N792);
not NOT1 (N1404, N1392);
and AND4 (N1405, N1396, N867, N645, N679);
nand NAND4 (N1406, N1405, N302, N802, N940);
and AND4 (N1407, N1404, N674, N555, N447);
and AND4 (N1408, N1406, N555, N471, N952);
and AND4 (N1409, N1401, N624, N760, N466);
xor XOR2 (N1410, N1383, N1330);
xor XOR2 (N1411, N1403, N103);
nand NAND4 (N1412, N1399, N1266, N107, N65);
xor XOR2 (N1413, N1412, N17);
nand NAND4 (N1414, N1398, N1241, N222, N1244);
buf BUF1 (N1415, N1408);
buf BUF1 (N1416, N1413);
or OR3 (N1417, N1416, N447, N635);
and AND4 (N1418, N1373, N440, N629, N649);
and AND2 (N1419, N1417, N816);
and AND2 (N1420, N1419, N249);
or OR2 (N1421, N1407, N265);
nand NAND3 (N1422, N1410, N265, N1188);
xor XOR2 (N1423, N1397, N817);
or OR2 (N1424, N1414, N1135);
nand NAND4 (N1425, N1421, N339, N664, N564);
and AND2 (N1426, N1390, N787);
or OR2 (N1427, N1409, N1129);
and AND3 (N1428, N1424, N63, N1380);
or OR4 (N1429, N1427, N967, N676, N1181);
not NOT1 (N1430, N1425);
not NOT1 (N1431, N1422);
not NOT1 (N1432, N1423);
nand NAND3 (N1433, N1432, N1140, N806);
or OR4 (N1434, N1415, N183, N1288, N446);
and AND4 (N1435, N1411, N725, N788, N300);
not NOT1 (N1436, N1426);
buf BUF1 (N1437, N1418);
not NOT1 (N1438, N1437);
or OR3 (N1439, N1435, N1378, N436);
or OR2 (N1440, N1434, N1328);
not NOT1 (N1441, N1433);
nor NOR4 (N1442, N1441, N760, N328, N1010);
or OR2 (N1443, N1431, N445);
buf BUF1 (N1444, N1438);
xor XOR2 (N1445, N1428, N1282);
nor NOR3 (N1446, N1429, N567, N698);
buf BUF1 (N1447, N1445);
buf BUF1 (N1448, N1446);
and AND3 (N1449, N1420, N1190, N1059);
buf BUF1 (N1450, N1439);
xor XOR2 (N1451, N1450, N235);
xor XOR2 (N1452, N1440, N816);
buf BUF1 (N1453, N1443);
not NOT1 (N1454, N1453);
xor XOR2 (N1455, N1449, N318);
nand NAND2 (N1456, N1447, N532);
or OR4 (N1457, N1448, N198, N216, N946);
xor XOR2 (N1458, N1442, N805);
nand NAND2 (N1459, N1451, N852);
or OR4 (N1460, N1456, N1415, N1326, N838);
xor XOR2 (N1461, N1457, N894);
nor NOR2 (N1462, N1436, N821);
nor NOR4 (N1463, N1430, N569, N988, N471);
nand NAND3 (N1464, N1462, N971, N485);
and AND2 (N1465, N1452, N681);
buf BUF1 (N1466, N1458);
buf BUF1 (N1467, N1464);
nand NAND2 (N1468, N1459, N371);
or OR4 (N1469, N1461, N1086, N1194, N1198);
nand NAND2 (N1470, N1455, N1152);
not NOT1 (N1471, N1460);
and AND2 (N1472, N1454, N1304);
nand NAND3 (N1473, N1470, N839, N560);
or OR4 (N1474, N1467, N1374, N1274, N598);
or OR4 (N1475, N1465, N86, N1188, N895);
xor XOR2 (N1476, N1471, N834);
nor NOR3 (N1477, N1469, N1012, N1255);
and AND4 (N1478, N1477, N1342, N878, N1285);
or OR4 (N1479, N1474, N1172, N113, N1043);
nand NAND2 (N1480, N1473, N11);
or OR2 (N1481, N1478, N112);
xor XOR2 (N1482, N1479, N322);
or OR2 (N1483, N1463, N696);
or OR3 (N1484, N1466, N1095, N981);
or OR4 (N1485, N1472, N650, N18, N945);
xor XOR2 (N1486, N1483, N270);
or OR3 (N1487, N1481, N108, N1485);
and AND4 (N1488, N291, N369, N1006, N1198);
or OR3 (N1489, N1487, N1255, N851);
nand NAND2 (N1490, N1482, N1021);
buf BUF1 (N1491, N1490);
nand NAND2 (N1492, N1491, N1482);
nand NAND2 (N1493, N1476, N1218);
nor NOR2 (N1494, N1492, N1149);
nand NAND3 (N1495, N1484, N1419, N497);
and AND3 (N1496, N1444, N945, N1148);
or OR2 (N1497, N1475, N928);
nor NOR3 (N1498, N1486, N972, N157);
nand NAND3 (N1499, N1494, N151, N437);
or OR3 (N1500, N1498, N706, N1499);
or OR4 (N1501, N1495, N871, N380, N242);
or OR4 (N1502, N1069, N1293, N445, N81);
xor XOR2 (N1503, N1489, N1454);
not NOT1 (N1504, N1480);
nor NOR3 (N1505, N1500, N33, N1485);
buf BUF1 (N1506, N1497);
buf BUF1 (N1507, N1502);
not NOT1 (N1508, N1507);
nand NAND2 (N1509, N1501, N838);
and AND4 (N1510, N1504, N383, N1046, N1151);
xor XOR2 (N1511, N1468, N1092);
not NOT1 (N1512, N1503);
nor NOR4 (N1513, N1509, N240, N320, N1432);
xor XOR2 (N1514, N1513, N1184);
buf BUF1 (N1515, N1511);
xor XOR2 (N1516, N1510, N871);
xor XOR2 (N1517, N1493, N1418);
and AND3 (N1518, N1516, N881, N1110);
nor NOR2 (N1519, N1518, N610);
not NOT1 (N1520, N1517);
buf BUF1 (N1521, N1520);
xor XOR2 (N1522, N1508, N380);
or OR2 (N1523, N1515, N822);
and AND4 (N1524, N1506, N1420, N1055, N1218);
nand NAND4 (N1525, N1519, N1206, N433, N976);
nand NAND3 (N1526, N1522, N478, N380);
nor NOR3 (N1527, N1496, N735, N929);
nand NAND2 (N1528, N1523, N205);
not NOT1 (N1529, N1524);
nand NAND4 (N1530, N1529, N831, N39, N150);
and AND3 (N1531, N1521, N262, N7);
nand NAND3 (N1532, N1530, N1079, N1193);
not NOT1 (N1533, N1525);
not NOT1 (N1534, N1532);
buf BUF1 (N1535, N1514);
or OR2 (N1536, N1528, N1267);
nor NOR2 (N1537, N1535, N839);
nor NOR2 (N1538, N1536, N1471);
nor NOR2 (N1539, N1527, N257);
or OR4 (N1540, N1533, N155, N437, N1136);
nor NOR3 (N1541, N1537, N340, N502);
nand NAND4 (N1542, N1538, N711, N1229, N1191);
xor XOR2 (N1543, N1488, N898);
nand NAND3 (N1544, N1539, N1360, N1061);
nor NOR2 (N1545, N1512, N59);
not NOT1 (N1546, N1505);
nor NOR2 (N1547, N1531, N1058);
nand NAND2 (N1548, N1540, N149);
not NOT1 (N1549, N1544);
nor NOR3 (N1550, N1549, N1540, N858);
not NOT1 (N1551, N1550);
nand NAND3 (N1552, N1548, N630, N600);
nand NAND4 (N1553, N1534, N950, N942, N1548);
xor XOR2 (N1554, N1546, N993);
not NOT1 (N1555, N1526);
not NOT1 (N1556, N1553);
nand NAND2 (N1557, N1556, N1181);
not NOT1 (N1558, N1541);
buf BUF1 (N1559, N1551);
nor NOR4 (N1560, N1542, N481, N1347, N665);
not NOT1 (N1561, N1559);
or OR2 (N1562, N1554, N842);
not NOT1 (N1563, N1560);
and AND2 (N1564, N1562, N274);
or OR2 (N1565, N1555, N1390);
nand NAND3 (N1566, N1565, N758, N1441);
not NOT1 (N1567, N1564);
xor XOR2 (N1568, N1557, N612);
or OR2 (N1569, N1563, N560);
not NOT1 (N1570, N1543);
xor XOR2 (N1571, N1561, N390);
nor NOR3 (N1572, N1552, N910, N901);
nand NAND4 (N1573, N1570, N400, N416, N747);
nand NAND3 (N1574, N1566, N1075, N537);
and AND3 (N1575, N1558, N371, N1047);
or OR3 (N1576, N1547, N1039, N1537);
xor XOR2 (N1577, N1571, N1446);
nand NAND4 (N1578, N1567, N1549, N1322, N381);
nor NOR2 (N1579, N1573, N1076);
xor XOR2 (N1580, N1575, N632);
nand NAND4 (N1581, N1578, N392, N705, N311);
not NOT1 (N1582, N1545);
nand NAND4 (N1583, N1574, N928, N691, N9);
not NOT1 (N1584, N1580);
xor XOR2 (N1585, N1579, N324);
and AND4 (N1586, N1576, N1455, N721, N160);
buf BUF1 (N1587, N1583);
buf BUF1 (N1588, N1585);
and AND2 (N1589, N1581, N762);
nor NOR3 (N1590, N1587, N940, N1514);
not NOT1 (N1591, N1590);
xor XOR2 (N1592, N1577, N419);
and AND2 (N1593, N1591, N1108);
buf BUF1 (N1594, N1589);
nor NOR2 (N1595, N1582, N1173);
buf BUF1 (N1596, N1592);
not NOT1 (N1597, N1593);
nand NAND3 (N1598, N1588, N413, N952);
buf BUF1 (N1599, N1594);
xor XOR2 (N1600, N1584, N667);
buf BUF1 (N1601, N1569);
not NOT1 (N1602, N1596);
nor NOR3 (N1603, N1598, N1504, N437);
xor XOR2 (N1604, N1599, N1085);
nor NOR4 (N1605, N1595, N559, N293, N778);
not NOT1 (N1606, N1601);
or OR2 (N1607, N1572, N1573);
nor NOR4 (N1608, N1600, N490, N763, N751);
nor NOR2 (N1609, N1605, N635);
nand NAND2 (N1610, N1604, N958);
or OR3 (N1611, N1602, N1424, N1075);
nand NAND4 (N1612, N1608, N994, N89, N612);
not NOT1 (N1613, N1607);
or OR2 (N1614, N1606, N1417);
and AND3 (N1615, N1613, N99, N1262);
xor XOR2 (N1616, N1609, N416);
not NOT1 (N1617, N1611);
not NOT1 (N1618, N1568);
nor NOR3 (N1619, N1615, N1323, N1353);
nor NOR3 (N1620, N1597, N1145, N297);
nor NOR2 (N1621, N1619, N696);
not NOT1 (N1622, N1617);
xor XOR2 (N1623, N1621, N592);
xor XOR2 (N1624, N1612, N1383);
or OR3 (N1625, N1620, N1333, N1265);
buf BUF1 (N1626, N1624);
buf BUF1 (N1627, N1603);
nor NOR2 (N1628, N1614, N465);
or OR4 (N1629, N1618, N810, N317, N1527);
and AND3 (N1630, N1586, N393, N571);
and AND4 (N1631, N1616, N1507, N891, N880);
buf BUF1 (N1632, N1631);
xor XOR2 (N1633, N1626, N630);
not NOT1 (N1634, N1622);
and AND4 (N1635, N1628, N716, N1249, N736);
nor NOR4 (N1636, N1633, N638, N926, N1433);
nand NAND3 (N1637, N1630, N132, N483);
not NOT1 (N1638, N1635);
or OR2 (N1639, N1627, N1224);
xor XOR2 (N1640, N1634, N893);
or OR2 (N1641, N1629, N114);
not NOT1 (N1642, N1639);
and AND4 (N1643, N1632, N410, N1282, N32);
nand NAND4 (N1644, N1641, N1623, N710, N1539);
not NOT1 (N1645, N203);
nor NOR4 (N1646, N1640, N1477, N1070, N77);
nor NOR3 (N1647, N1646, N872, N1502);
nand NAND4 (N1648, N1638, N566, N1104, N1118);
buf BUF1 (N1649, N1643);
nand NAND4 (N1650, N1645, N1035, N1150, N1289);
nand NAND2 (N1651, N1649, N812);
or OR3 (N1652, N1648, N836, N496);
or OR3 (N1653, N1647, N1391, N135);
nor NOR2 (N1654, N1644, N1232);
and AND4 (N1655, N1625, N1471, N192, N367);
nor NOR4 (N1656, N1637, N56, N137, N664);
buf BUF1 (N1657, N1636);
buf BUF1 (N1658, N1651);
not NOT1 (N1659, N1652);
nor NOR4 (N1660, N1654, N751, N1305, N1275);
xor XOR2 (N1661, N1653, N672);
buf BUF1 (N1662, N1657);
and AND3 (N1663, N1642, N330, N1335);
or OR3 (N1664, N1660, N1140, N730);
or OR3 (N1665, N1610, N1155, N1342);
nand NAND4 (N1666, N1663, N1109, N1382, N414);
buf BUF1 (N1667, N1661);
not NOT1 (N1668, N1650);
not NOT1 (N1669, N1664);
buf BUF1 (N1670, N1669);
nand NAND3 (N1671, N1665, N9, N920);
or OR3 (N1672, N1668, N1643, N966);
not NOT1 (N1673, N1671);
nor NOR2 (N1674, N1655, N1514);
nor NOR3 (N1675, N1672, N80, N805);
nand NAND3 (N1676, N1666, N244, N1436);
or OR4 (N1677, N1659, N1503, N1409, N1504);
xor XOR2 (N1678, N1675, N1217);
and AND4 (N1679, N1658, N1200, N310, N1332);
not NOT1 (N1680, N1673);
or OR3 (N1681, N1674, N1564, N1558);
or OR2 (N1682, N1667, N1035);
and AND2 (N1683, N1681, N1383);
nor NOR4 (N1684, N1656, N381, N477, N1587);
nand NAND4 (N1685, N1682, N481, N1123, N1175);
nand NAND3 (N1686, N1679, N246, N655);
and AND3 (N1687, N1676, N1094, N75);
and AND3 (N1688, N1677, N1556, N331);
nand NAND4 (N1689, N1670, N410, N395, N95);
and AND2 (N1690, N1685, N1171);
not NOT1 (N1691, N1687);
nor NOR4 (N1692, N1662, N521, N764, N1616);
nor NOR4 (N1693, N1686, N899, N829, N886);
xor XOR2 (N1694, N1690, N240);
nand NAND2 (N1695, N1691, N317);
or OR4 (N1696, N1692, N285, N1678, N753);
nor NOR4 (N1697, N1181, N606, N480, N111);
buf BUF1 (N1698, N1693);
buf BUF1 (N1699, N1684);
nand NAND4 (N1700, N1696, N673, N816, N1376);
not NOT1 (N1701, N1688);
not NOT1 (N1702, N1698);
not NOT1 (N1703, N1697);
or OR2 (N1704, N1689, N1626);
nand NAND4 (N1705, N1700, N791, N1646, N1130);
buf BUF1 (N1706, N1694);
nor NOR4 (N1707, N1683, N1072, N793, N1208);
and AND3 (N1708, N1706, N1348, N326);
or OR3 (N1709, N1705, N1306, N1567);
nand NAND4 (N1710, N1709, N1014, N920, N457);
nor NOR2 (N1711, N1704, N214);
xor XOR2 (N1712, N1710, N718);
buf BUF1 (N1713, N1680);
and AND2 (N1714, N1701, N1063);
nor NOR2 (N1715, N1711, N1308);
nand NAND2 (N1716, N1703, N640);
nand NAND2 (N1717, N1699, N1358);
and AND3 (N1718, N1695, N137, N1523);
and AND3 (N1719, N1713, N142, N405);
buf BUF1 (N1720, N1712);
or OR4 (N1721, N1719, N413, N242, N1189);
xor XOR2 (N1722, N1718, N67);
xor XOR2 (N1723, N1708, N246);
nand NAND2 (N1724, N1723, N395);
xor XOR2 (N1725, N1707, N1151);
nor NOR3 (N1726, N1716, N354, N954);
or OR3 (N1727, N1724, N1494, N982);
buf BUF1 (N1728, N1725);
buf BUF1 (N1729, N1715);
not NOT1 (N1730, N1717);
nor NOR2 (N1731, N1726, N216);
not NOT1 (N1732, N1730);
buf BUF1 (N1733, N1722);
nand NAND3 (N1734, N1721, N1659, N875);
or OR2 (N1735, N1727, N1113);
not NOT1 (N1736, N1720);
nor NOR4 (N1737, N1702, N642, N833, N338);
or OR2 (N1738, N1714, N469);
nor NOR2 (N1739, N1728, N1492);
not NOT1 (N1740, N1737);
buf BUF1 (N1741, N1736);
buf BUF1 (N1742, N1729);
not NOT1 (N1743, N1731);
not NOT1 (N1744, N1733);
or OR4 (N1745, N1735, N1371, N665, N564);
xor XOR2 (N1746, N1745, N362);
not NOT1 (N1747, N1740);
not NOT1 (N1748, N1739);
nand NAND4 (N1749, N1734, N222, N681, N544);
not NOT1 (N1750, N1738);
not NOT1 (N1751, N1749);
nand NAND3 (N1752, N1743, N117, N1052);
or OR2 (N1753, N1747, N431);
xor XOR2 (N1754, N1748, N1007);
or OR2 (N1755, N1752, N846);
and AND2 (N1756, N1751, N70);
not NOT1 (N1757, N1755);
xor XOR2 (N1758, N1754, N474);
not NOT1 (N1759, N1750);
or OR3 (N1760, N1753, N850, N438);
nand NAND2 (N1761, N1757, N110);
buf BUF1 (N1762, N1746);
nor NOR3 (N1763, N1756, N389, N1622);
nor NOR3 (N1764, N1741, N553, N1325);
not NOT1 (N1765, N1744);
nand NAND4 (N1766, N1758, N15, N1230, N1395);
nor NOR4 (N1767, N1765, N537, N1329, N1111);
xor XOR2 (N1768, N1764, N436);
buf BUF1 (N1769, N1767);
not NOT1 (N1770, N1760);
not NOT1 (N1771, N1762);
nor NOR4 (N1772, N1742, N1223, N119, N1173);
and AND3 (N1773, N1766, N1166, N801);
not NOT1 (N1774, N1769);
buf BUF1 (N1775, N1773);
nor NOR2 (N1776, N1772, N1030);
and AND3 (N1777, N1774, N779, N856);
xor XOR2 (N1778, N1776, N1379);
nand NAND4 (N1779, N1768, N919, N460, N1544);
not NOT1 (N1780, N1777);
and AND3 (N1781, N1778, N138, N1077);
nand NAND2 (N1782, N1770, N902);
nor NOR4 (N1783, N1781, N700, N1487, N1496);
nand NAND4 (N1784, N1771, N927, N1626, N840);
not NOT1 (N1785, N1732);
buf BUF1 (N1786, N1780);
nand NAND3 (N1787, N1786, N120, N727);
xor XOR2 (N1788, N1759, N515);
not NOT1 (N1789, N1783);
not NOT1 (N1790, N1761);
xor XOR2 (N1791, N1779, N722);
xor XOR2 (N1792, N1788, N727);
and AND4 (N1793, N1790, N506, N1364, N1182);
buf BUF1 (N1794, N1775);
and AND3 (N1795, N1784, N1198, N902);
nand NAND4 (N1796, N1791, N597, N1161, N480);
nor NOR2 (N1797, N1787, N1578);
nor NOR3 (N1798, N1796, N1381, N923);
buf BUF1 (N1799, N1785);
or OR4 (N1800, N1793, N1419, N332, N341);
nand NAND4 (N1801, N1789, N1499, N1666, N1526);
xor XOR2 (N1802, N1795, N1507);
nor NOR4 (N1803, N1763, N176, N515, N522);
not NOT1 (N1804, N1782);
buf BUF1 (N1805, N1803);
or OR3 (N1806, N1799, N428, N418);
nor NOR4 (N1807, N1806, N325, N176, N1102);
nor NOR4 (N1808, N1797, N803, N1573, N1683);
buf BUF1 (N1809, N1802);
and AND4 (N1810, N1805, N1163, N84, N1275);
nor NOR3 (N1811, N1809, N347, N1269);
not NOT1 (N1812, N1811);
not NOT1 (N1813, N1804);
not NOT1 (N1814, N1810);
not NOT1 (N1815, N1814);
not NOT1 (N1816, N1792);
nor NOR2 (N1817, N1807, N1778);
nor NOR4 (N1818, N1808, N346, N829, N10);
xor XOR2 (N1819, N1817, N1685);
xor XOR2 (N1820, N1812, N530);
nand NAND2 (N1821, N1800, N375);
buf BUF1 (N1822, N1801);
and AND2 (N1823, N1816, N700);
or OR2 (N1824, N1813, N864);
xor XOR2 (N1825, N1798, N85);
buf BUF1 (N1826, N1824);
or OR3 (N1827, N1815, N259, N1751);
nor NOR4 (N1828, N1818, N569, N1711, N1540);
and AND2 (N1829, N1823, N113);
not NOT1 (N1830, N1825);
not NOT1 (N1831, N1826);
nand NAND4 (N1832, N1830, N1583, N254, N1375);
buf BUF1 (N1833, N1820);
not NOT1 (N1834, N1831);
and AND2 (N1835, N1827, N488);
nor NOR4 (N1836, N1834, N1002, N1579, N1702);
and AND2 (N1837, N1794, N1428);
not NOT1 (N1838, N1835);
buf BUF1 (N1839, N1832);
not NOT1 (N1840, N1822);
nor NOR3 (N1841, N1819, N823, N1260);
nor NOR3 (N1842, N1839, N423, N1666);
or OR3 (N1843, N1821, N1469, N1018);
xor XOR2 (N1844, N1837, N247);
buf BUF1 (N1845, N1841);
nand NAND2 (N1846, N1840, N232);
not NOT1 (N1847, N1844);
not NOT1 (N1848, N1838);
or OR3 (N1849, N1847, N994, N1505);
buf BUF1 (N1850, N1848);
xor XOR2 (N1851, N1843, N132);
and AND2 (N1852, N1851, N1083);
or OR4 (N1853, N1849, N1469, N1509, N1306);
nand NAND2 (N1854, N1846, N726);
nand NAND3 (N1855, N1850, N1332, N1122);
and AND4 (N1856, N1852, N184, N497, N1779);
or OR4 (N1857, N1833, N1555, N135, N642);
or OR2 (N1858, N1829, N490);
nand NAND2 (N1859, N1854, N1768);
buf BUF1 (N1860, N1858);
nor NOR4 (N1861, N1853, N250, N1047, N631);
or OR2 (N1862, N1855, N135);
not NOT1 (N1863, N1836);
and AND4 (N1864, N1828, N1358, N1835, N366);
not NOT1 (N1865, N1857);
nand NAND2 (N1866, N1860, N529);
not NOT1 (N1867, N1859);
xor XOR2 (N1868, N1864, N1395);
not NOT1 (N1869, N1856);
and AND2 (N1870, N1867, N985);
nor NOR4 (N1871, N1868, N1718, N161, N283);
nor NOR2 (N1872, N1862, N650);
not NOT1 (N1873, N1861);
nor NOR2 (N1874, N1842, N1300);
and AND2 (N1875, N1874, N1006);
nor NOR2 (N1876, N1869, N993);
nor NOR4 (N1877, N1876, N1543, N1571, N1207);
not NOT1 (N1878, N1865);
buf BUF1 (N1879, N1872);
or OR3 (N1880, N1879, N897, N1610);
xor XOR2 (N1881, N1877, N470);
xor XOR2 (N1882, N1870, N1646);
nor NOR3 (N1883, N1866, N1842, N1085);
nor NOR3 (N1884, N1863, N133, N1876);
not NOT1 (N1885, N1884);
nor NOR2 (N1886, N1875, N469);
and AND4 (N1887, N1885, N1192, N1830, N1344);
buf BUF1 (N1888, N1881);
xor XOR2 (N1889, N1873, N179);
nor NOR4 (N1890, N1887, N1016, N1021, N1767);
nor NOR2 (N1891, N1886, N1201);
buf BUF1 (N1892, N1889);
nor NOR3 (N1893, N1882, N148, N169);
nand NAND4 (N1894, N1883, N373, N331, N340);
and AND4 (N1895, N1871, N130, N1645, N153);
not NOT1 (N1896, N1891);
nor NOR4 (N1897, N1893, N898, N1327, N1225);
or OR3 (N1898, N1878, N367, N236);
or OR2 (N1899, N1898, N1232);
nand NAND4 (N1900, N1880, N1206, N1230, N1768);
nand NAND4 (N1901, N1895, N750, N391, N1216);
xor XOR2 (N1902, N1888, N1846);
buf BUF1 (N1903, N1892);
nor NOR2 (N1904, N1894, N1686);
and AND2 (N1905, N1896, N418);
and AND3 (N1906, N1899, N1553, N1799);
nor NOR4 (N1907, N1845, N1511, N1450, N623);
nor NOR2 (N1908, N1900, N1853);
xor XOR2 (N1909, N1901, N451);
nand NAND4 (N1910, N1908, N503, N1052, N659);
nand NAND3 (N1911, N1897, N821, N1186);
nand NAND2 (N1912, N1906, N599);
not NOT1 (N1913, N1903);
or OR2 (N1914, N1890, N484);
nor NOR4 (N1915, N1909, N163, N1901, N1232);
not NOT1 (N1916, N1914);
nor NOR3 (N1917, N1905, N1033, N1172);
or OR2 (N1918, N1907, N828);
and AND3 (N1919, N1910, N782, N1652);
buf BUF1 (N1920, N1917);
buf BUF1 (N1921, N1915);
buf BUF1 (N1922, N1911);
and AND3 (N1923, N1912, N1842, N1633);
or OR4 (N1924, N1922, N35, N525, N972);
not NOT1 (N1925, N1904);
nand NAND2 (N1926, N1919, N192);
buf BUF1 (N1927, N1923);
nor NOR3 (N1928, N1925, N712, N721);
nor NOR3 (N1929, N1927, N16, N697);
nand NAND3 (N1930, N1929, N543, N353);
nor NOR2 (N1931, N1926, N660);
and AND3 (N1932, N1921, N461, N599);
or OR2 (N1933, N1932, N1694);
nor NOR4 (N1934, N1902, N1, N770, N819);
nand NAND4 (N1935, N1918, N986, N676, N315);
not NOT1 (N1936, N1930);
or OR3 (N1937, N1934, N792, N1935);
nor NOR2 (N1938, N614, N1663);
not NOT1 (N1939, N1913);
buf BUF1 (N1940, N1931);
or OR2 (N1941, N1936, N1356);
or OR3 (N1942, N1938, N1591, N1398);
or OR4 (N1943, N1924, N495, N1898, N912);
not NOT1 (N1944, N1928);
or OR2 (N1945, N1941, N758);
nor NOR4 (N1946, N1944, N27, N1044, N946);
xor XOR2 (N1947, N1937, N1367);
not NOT1 (N1948, N1942);
nand NAND4 (N1949, N1947, N1331, N1186, N683);
or OR2 (N1950, N1920, N503);
or OR4 (N1951, N1950, N710, N1469, N403);
xor XOR2 (N1952, N1939, N1047);
or OR2 (N1953, N1951, N149);
and AND4 (N1954, N1952, N42, N1829, N1155);
or OR2 (N1955, N1949, N504);
buf BUF1 (N1956, N1948);
nand NAND2 (N1957, N1946, N778);
nor NOR4 (N1958, N1953, N1229, N636, N140);
and AND3 (N1959, N1955, N1663, N1825);
not NOT1 (N1960, N1958);
not NOT1 (N1961, N1943);
not NOT1 (N1962, N1916);
and AND2 (N1963, N1962, N784);
or OR3 (N1964, N1963, N384, N465);
xor XOR2 (N1965, N1933, N481);
nand NAND2 (N1966, N1956, N278);
nor NOR4 (N1967, N1961, N1804, N700, N1353);
nor NOR3 (N1968, N1960, N1945, N497);
or OR3 (N1969, N1507, N1193, N743);
or OR3 (N1970, N1954, N1155, N592);
nand NAND2 (N1971, N1957, N27);
not NOT1 (N1972, N1964);
xor XOR2 (N1973, N1959, N36);
xor XOR2 (N1974, N1970, N1767);
xor XOR2 (N1975, N1965, N541);
buf BUF1 (N1976, N1966);
xor XOR2 (N1977, N1975, N1407);
buf BUF1 (N1978, N1968);
or OR3 (N1979, N1972, N1022, N1805);
buf BUF1 (N1980, N1978);
nor NOR3 (N1981, N1969, N299, N961);
or OR4 (N1982, N1979, N611, N916, N249);
buf BUF1 (N1983, N1971);
nor NOR2 (N1984, N1977, N1280);
and AND4 (N1985, N1976, N346, N1866, N1509);
or OR4 (N1986, N1967, N883, N231, N1940);
and AND4 (N1987, N1304, N1381, N135, N107);
nor NOR3 (N1988, N1986, N1368, N880);
buf BUF1 (N1989, N1984);
or OR3 (N1990, N1973, N795, N936);
xor XOR2 (N1991, N1988, N1353);
nand NAND4 (N1992, N1980, N175, N1042, N645);
xor XOR2 (N1993, N1992, N1151);
xor XOR2 (N1994, N1987, N304);
nand NAND2 (N1995, N1989, N1572);
nand NAND2 (N1996, N1974, N1070);
nor NOR4 (N1997, N1995, N554, N1203, N1889);
or OR4 (N1998, N1996, N391, N268, N1420);
buf BUF1 (N1999, N1991);
or OR2 (N2000, N1993, N1384);
or OR3 (N2001, N1985, N1765, N1342);
buf BUF1 (N2002, N1982);
nand NAND2 (N2003, N1998, N1408);
and AND4 (N2004, N2001, N821, N1625, N201);
and AND3 (N2005, N1983, N330, N1296);
nor NOR2 (N2006, N2005, N1296);
xor XOR2 (N2007, N2006, N688);
xor XOR2 (N2008, N1990, N1897);
nand NAND3 (N2009, N1981, N304, N1383);
xor XOR2 (N2010, N1999, N305);
not NOT1 (N2011, N2002);
or OR3 (N2012, N2010, N1251, N1816);
xor XOR2 (N2013, N2000, N480);
not NOT1 (N2014, N2008);
buf BUF1 (N2015, N2009);
nand NAND2 (N2016, N1997, N1037);
xor XOR2 (N2017, N2003, N546);
and AND4 (N2018, N2015, N620, N1248, N1940);
not NOT1 (N2019, N2017);
not NOT1 (N2020, N2018);
xor XOR2 (N2021, N2019, N513);
nor NOR2 (N2022, N2020, N1496);
xor XOR2 (N2023, N2021, N729);
nand NAND2 (N2024, N2013, N1575);
nand NAND2 (N2025, N1994, N1496);
not NOT1 (N2026, N2025);
xor XOR2 (N2027, N2004, N153);
not NOT1 (N2028, N2016);
or OR2 (N2029, N2014, N855);
nor NOR4 (N2030, N2011, N1182, N1695, N987);
and AND2 (N2031, N2030, N1688);
nand NAND3 (N2032, N2029, N499, N766);
not NOT1 (N2033, N2022);
nor NOR4 (N2034, N2028, N1793, N1852, N1642);
and AND4 (N2035, N2032, N456, N1214, N529);
buf BUF1 (N2036, N2012);
buf BUF1 (N2037, N2035);
buf BUF1 (N2038, N2026);
and AND2 (N2039, N2036, N1073);
and AND4 (N2040, N2023, N740, N1130, N218);
buf BUF1 (N2041, N2039);
buf BUF1 (N2042, N2033);
not NOT1 (N2043, N2041);
or OR4 (N2044, N2040, N838, N1268, N1248);
nor NOR3 (N2045, N2044, N1289, N1272);
buf BUF1 (N2046, N2037);
nor NOR3 (N2047, N2045, N435, N200);
not NOT1 (N2048, N2024);
or OR3 (N2049, N2034, N1678, N46);
and AND3 (N2050, N2031, N1646, N580);
or OR4 (N2051, N2027, N404, N1017, N1743);
nand NAND4 (N2052, N2050, N1268, N251, N271);
nor NOR4 (N2053, N2042, N908, N1842, N1706);
buf BUF1 (N2054, N2043);
or OR4 (N2055, N2038, N445, N354, N1714);
buf BUF1 (N2056, N2047);
and AND2 (N2057, N2051, N970);
or OR2 (N2058, N2053, N1827);
buf BUF1 (N2059, N2057);
buf BUF1 (N2060, N2054);
nor NOR3 (N2061, N2058, N1217, N617);
nand NAND3 (N2062, N2048, N1409, N2045);
nand NAND2 (N2063, N2056, N1604);
nand NAND3 (N2064, N2060, N1243, N266);
not NOT1 (N2065, N2052);
or OR3 (N2066, N2007, N411, N245);
nor NOR2 (N2067, N2061, N1051);
not NOT1 (N2068, N2065);
buf BUF1 (N2069, N2062);
and AND2 (N2070, N2046, N1302);
and AND4 (N2071, N2064, N871, N1855, N1020);
not NOT1 (N2072, N2059);
not NOT1 (N2073, N2049);
not NOT1 (N2074, N2071);
nor NOR2 (N2075, N2068, N488);
or OR2 (N2076, N2069, N412);
nor NOR4 (N2077, N2070, N384, N1783, N1696);
buf BUF1 (N2078, N2063);
buf BUF1 (N2079, N2072);
nor NOR2 (N2080, N2079, N412);
buf BUF1 (N2081, N2073);
nand NAND2 (N2082, N2081, N1342);
buf BUF1 (N2083, N2055);
nand NAND4 (N2084, N2083, N1057, N302, N669);
not NOT1 (N2085, N2084);
and AND4 (N2086, N2074, N1585, N1037, N438);
and AND4 (N2087, N2066, N528, N964, N1443);
or OR3 (N2088, N2086, N1602, N218);
and AND2 (N2089, N2088, N1857);
and AND3 (N2090, N2089, N2078, N2012);
not NOT1 (N2091, N1071);
nor NOR2 (N2092, N2076, N530);
nor NOR2 (N2093, N2082, N1325);
not NOT1 (N2094, N2067);
nor NOR4 (N2095, N2085, N1332, N1592, N1800);
buf BUF1 (N2096, N2090);
or OR2 (N2097, N2075, N2034);
xor XOR2 (N2098, N2093, N711);
nand NAND3 (N2099, N2080, N1873, N1611);
not NOT1 (N2100, N2096);
xor XOR2 (N2101, N2100, N642);
or OR3 (N2102, N2097, N295, N2086);
nor NOR4 (N2103, N2098, N1056, N484, N279);
nand NAND4 (N2104, N2094, N40, N1809, N912);
nand NAND2 (N2105, N2092, N1508);
buf BUF1 (N2106, N2105);
or OR2 (N2107, N2077, N1708);
nor NOR4 (N2108, N2099, N604, N1484, N1572);
or OR4 (N2109, N2104, N1510, N878, N99);
not NOT1 (N2110, N2101);
nor NOR4 (N2111, N2109, N1372, N1429, N1234);
nor NOR4 (N2112, N2087, N252, N1102, N568);
not NOT1 (N2113, N2108);
xor XOR2 (N2114, N2113, N535);
xor XOR2 (N2115, N2107, N1065);
nor NOR4 (N2116, N2111, N1098, N1585, N1312);
and AND4 (N2117, N2110, N314, N1170, N1464);
nor NOR3 (N2118, N2103, N1592, N412);
not NOT1 (N2119, N2114);
nand NAND2 (N2120, N2112, N929);
buf BUF1 (N2121, N2116);
or OR3 (N2122, N2121, N761, N2080);
buf BUF1 (N2123, N2102);
nor NOR2 (N2124, N2122, N1987);
nand NAND2 (N2125, N2106, N333);
xor XOR2 (N2126, N2117, N1550);
buf BUF1 (N2127, N2124);
xor XOR2 (N2128, N2095, N507);
and AND2 (N2129, N2119, N1694);
buf BUF1 (N2130, N2128);
not NOT1 (N2131, N2126);
xor XOR2 (N2132, N2115, N1434);
or OR4 (N2133, N2129, N1616, N1168, N615);
nor NOR4 (N2134, N2123, N1769, N73, N885);
or OR2 (N2135, N2125, N1147);
not NOT1 (N2136, N2118);
buf BUF1 (N2137, N2132);
xor XOR2 (N2138, N2120, N205);
or OR4 (N2139, N2137, N1051, N923, N1071);
nand NAND2 (N2140, N2091, N1361);
and AND2 (N2141, N2136, N1782);
not NOT1 (N2142, N2138);
and AND3 (N2143, N2127, N1614, N1778);
buf BUF1 (N2144, N2131);
buf BUF1 (N2145, N2139);
nor NOR2 (N2146, N2143, N711);
and AND2 (N2147, N2130, N1425);
or OR3 (N2148, N2142, N1318, N1564);
buf BUF1 (N2149, N2147);
nor NOR2 (N2150, N2148, N437);
nand NAND4 (N2151, N2145, N1860, N1357, N975);
nand NAND4 (N2152, N2151, N148, N1880, N172);
and AND3 (N2153, N2144, N1449, N1457);
and AND3 (N2154, N2149, N2041, N255);
buf BUF1 (N2155, N2150);
nand NAND4 (N2156, N2154, N1276, N2101, N1664);
nor NOR3 (N2157, N2155, N506, N2017);
not NOT1 (N2158, N2133);
nor NOR2 (N2159, N2156, N412);
nor NOR3 (N2160, N2134, N1889, N630);
nor NOR3 (N2161, N2135, N1577, N1826);
xor XOR2 (N2162, N2146, N66);
and AND3 (N2163, N2161, N1678, N2039);
buf BUF1 (N2164, N2162);
not NOT1 (N2165, N2158);
nor NOR2 (N2166, N2159, N1124);
nand NAND4 (N2167, N2160, N989, N1723, N1456);
nand NAND3 (N2168, N2157, N1941, N1583);
nand NAND3 (N2169, N2168, N1561, N39);
nand NAND4 (N2170, N2165, N288, N1753, N1773);
nor NOR4 (N2171, N2166, N1454, N603, N360);
xor XOR2 (N2172, N2153, N1899);
not NOT1 (N2173, N2164);
buf BUF1 (N2174, N2173);
not NOT1 (N2175, N2174);
not NOT1 (N2176, N2152);
buf BUF1 (N2177, N2175);
xor XOR2 (N2178, N2140, N1674);
nor NOR4 (N2179, N2178, N2017, N1264, N1658);
and AND2 (N2180, N2170, N1251);
and AND3 (N2181, N2163, N1974, N689);
xor XOR2 (N2182, N2176, N65);
buf BUF1 (N2183, N2167);
nand NAND3 (N2184, N2177, N840, N797);
buf BUF1 (N2185, N2184);
and AND2 (N2186, N2181, N1349);
nor NOR2 (N2187, N2179, N2158);
buf BUF1 (N2188, N2141);
or OR2 (N2189, N2182, N993);
not NOT1 (N2190, N2172);
buf BUF1 (N2191, N2190);
nor NOR3 (N2192, N2188, N279, N681);
buf BUF1 (N2193, N2180);
nor NOR4 (N2194, N2191, N541, N131, N747);
and AND2 (N2195, N2193, N245);
nor NOR4 (N2196, N2189, N1460, N582, N1691);
nand NAND3 (N2197, N2187, N1026, N1892);
xor XOR2 (N2198, N2185, N352);
and AND3 (N2199, N2192, N958, N1226);
nor NOR4 (N2200, N2183, N1887, N98, N29);
nor NOR2 (N2201, N2194, N21);
and AND3 (N2202, N2197, N116, N1040);
nor NOR4 (N2203, N2195, N2056, N341, N1793);
nor NOR3 (N2204, N2186, N1577, N1539);
or OR4 (N2205, N2171, N419, N456, N2147);
and AND2 (N2206, N2199, N107);
nor NOR3 (N2207, N2205, N1081, N213);
buf BUF1 (N2208, N2169);
nand NAND4 (N2209, N2200, N327, N1913, N1423);
nand NAND4 (N2210, N2209, N316, N414, N628);
buf BUF1 (N2211, N2202);
buf BUF1 (N2212, N2198);
nor NOR4 (N2213, N2204, N57, N2042, N1393);
or OR4 (N2214, N2207, N1588, N759, N615);
and AND4 (N2215, N2212, N1488, N1660, N2094);
buf BUF1 (N2216, N2215);
nor NOR4 (N2217, N2201, N15, N2160, N1261);
and AND2 (N2218, N2217, N2180);
and AND3 (N2219, N2206, N865, N2195);
buf BUF1 (N2220, N2211);
nand NAND3 (N2221, N2210, N2071, N379);
xor XOR2 (N2222, N2220, N111);
nand NAND2 (N2223, N2218, N824);
or OR2 (N2224, N2203, N1944);
buf BUF1 (N2225, N2221);
or OR3 (N2226, N2225, N670, N1991);
nor NOR3 (N2227, N2224, N635, N2190);
nor NOR2 (N2228, N2213, N1840);
nand NAND4 (N2229, N2223, N2068, N1439, N1765);
xor XOR2 (N2230, N2214, N462);
nor NOR4 (N2231, N2208, N1525, N557, N1911);
or OR2 (N2232, N2229, N581);
not NOT1 (N2233, N2232);
xor XOR2 (N2234, N2226, N831);
and AND4 (N2235, N2219, N287, N367, N712);
nor NOR3 (N2236, N2196, N1850, N1149);
not NOT1 (N2237, N2222);
not NOT1 (N2238, N2237);
and AND2 (N2239, N2238, N1539);
or OR4 (N2240, N2227, N2, N381, N1661);
buf BUF1 (N2241, N2230);
nand NAND3 (N2242, N2216, N2185, N1643);
and AND2 (N2243, N2231, N1992);
nor NOR3 (N2244, N2239, N520, N1385);
or OR3 (N2245, N2234, N1757, N653);
buf BUF1 (N2246, N2241);
and AND2 (N2247, N2233, N1228);
nor NOR3 (N2248, N2242, N1989, N396);
nor NOR3 (N2249, N2228, N213, N152);
or OR4 (N2250, N2243, N1608, N322, N266);
nor NOR2 (N2251, N2245, N1833);
nor NOR3 (N2252, N2250, N312, N1168);
xor XOR2 (N2253, N2251, N1443);
xor XOR2 (N2254, N2246, N1009);
or OR4 (N2255, N2236, N1442, N819, N411);
buf BUF1 (N2256, N2249);
or OR3 (N2257, N2255, N352, N335);
xor XOR2 (N2258, N2240, N1835);
xor XOR2 (N2259, N2252, N1155);
nand NAND4 (N2260, N2244, N605, N2021, N1929);
buf BUF1 (N2261, N2260);
or OR2 (N2262, N2253, N745);
buf BUF1 (N2263, N2256);
or OR3 (N2264, N2235, N960, N1207);
buf BUF1 (N2265, N2263);
or OR4 (N2266, N2247, N857, N931, N1498);
and AND3 (N2267, N2257, N381, N1447);
nor NOR2 (N2268, N2258, N1871);
or OR3 (N2269, N2259, N100, N1269);
nand NAND3 (N2270, N2269, N1784, N497);
nand NAND4 (N2271, N2266, N1504, N1762, N800);
buf BUF1 (N2272, N2268);
nand NAND4 (N2273, N2265, N291, N2035, N1012);
and AND4 (N2274, N2262, N156, N1087, N1770);
nor NOR3 (N2275, N2254, N849, N555);
or OR3 (N2276, N2273, N140, N1433);
or OR2 (N2277, N2270, N584);
nor NOR4 (N2278, N2276, N2234, N236, N1678);
not NOT1 (N2279, N2248);
buf BUF1 (N2280, N2275);
xor XOR2 (N2281, N2271, N1257);
buf BUF1 (N2282, N2261);
xor XOR2 (N2283, N2278, N411);
nor NOR3 (N2284, N2272, N1533, N1349);
and AND3 (N2285, N2279, N1116, N2099);
nand NAND3 (N2286, N2264, N1439, N824);
and AND2 (N2287, N2284, N1136);
or OR3 (N2288, N2277, N2233, N1317);
buf BUF1 (N2289, N2282);
not NOT1 (N2290, N2280);
not NOT1 (N2291, N2283);
not NOT1 (N2292, N2289);
not NOT1 (N2293, N2291);
and AND3 (N2294, N2288, N1213, N1168);
xor XOR2 (N2295, N2287, N1886);
xor XOR2 (N2296, N2295, N189);
nand NAND2 (N2297, N2286, N1188);
nand NAND3 (N2298, N2294, N2285, N1071);
xor XOR2 (N2299, N1921, N1985);
not NOT1 (N2300, N2296);
buf BUF1 (N2301, N2293);
nand NAND2 (N2302, N2274, N1944);
nor NOR3 (N2303, N2302, N1364, N1531);
or OR2 (N2304, N2281, N1332);
xor XOR2 (N2305, N2301, N464);
nor NOR4 (N2306, N2303, N1980, N487, N472);
xor XOR2 (N2307, N2292, N1856);
nor NOR4 (N2308, N2298, N2222, N317, N1695);
or OR3 (N2309, N2290, N1484, N455);
and AND4 (N2310, N2309, N602, N2301, N33);
not NOT1 (N2311, N2297);
nand NAND2 (N2312, N2304, N1586);
xor XOR2 (N2313, N2305, N1490);
xor XOR2 (N2314, N2310, N1862);
not NOT1 (N2315, N2299);
nor NOR2 (N2316, N2313, N1201);
buf BUF1 (N2317, N2312);
nand NAND4 (N2318, N2307, N2196, N1455, N205);
or OR3 (N2319, N2300, N2191, N761);
not NOT1 (N2320, N2306);
xor XOR2 (N2321, N2319, N473);
or OR2 (N2322, N2316, N281);
buf BUF1 (N2323, N2315);
not NOT1 (N2324, N2267);
nand NAND2 (N2325, N2320, N2321);
not NOT1 (N2326, N1165);
buf BUF1 (N2327, N2326);
and AND4 (N2328, N2318, N944, N1682, N1692);
buf BUF1 (N2329, N2317);
nor NOR2 (N2330, N2323, N344);
and AND3 (N2331, N2327, N282, N1765);
and AND4 (N2332, N2325, N1951, N1867, N1346);
nand NAND2 (N2333, N2308, N519);
nand NAND2 (N2334, N2328, N2084);
buf BUF1 (N2335, N2331);
or OR4 (N2336, N2314, N505, N1576, N1179);
xor XOR2 (N2337, N2334, N1593);
or OR4 (N2338, N2332, N1868, N182, N727);
and AND3 (N2339, N2330, N564, N1367);
nor NOR2 (N2340, N2329, N1917);
or OR4 (N2341, N2324, N2156, N207, N307);
or OR4 (N2342, N2337, N575, N264, N1525);
and AND2 (N2343, N2338, N922);
nor NOR3 (N2344, N2341, N298, N233);
xor XOR2 (N2345, N2333, N1545);
and AND4 (N2346, N2339, N107, N1688, N1801);
not NOT1 (N2347, N2346);
nand NAND4 (N2348, N2340, N1286, N1983, N2121);
nand NAND3 (N2349, N2322, N981, N662);
buf BUF1 (N2350, N2336);
not NOT1 (N2351, N2348);
buf BUF1 (N2352, N2343);
or OR4 (N2353, N2349, N2341, N1783, N338);
nor NOR4 (N2354, N2345, N892, N1815, N717);
not NOT1 (N2355, N2335);
not NOT1 (N2356, N2342);
nand NAND4 (N2357, N2353, N1379, N1705, N413);
nand NAND2 (N2358, N2344, N2294);
xor XOR2 (N2359, N2347, N1196);
buf BUF1 (N2360, N2356);
buf BUF1 (N2361, N2354);
not NOT1 (N2362, N2352);
or OR4 (N2363, N2358, N1735, N535, N2186);
or OR4 (N2364, N2355, N2152, N808, N966);
nand NAND2 (N2365, N2363, N1021);
xor XOR2 (N2366, N2360, N1574);
not NOT1 (N2367, N2351);
and AND4 (N2368, N2364, N2200, N1714, N1237);
not NOT1 (N2369, N2311);
xor XOR2 (N2370, N2368, N1386);
nor NOR3 (N2371, N2350, N2276, N1742);
not NOT1 (N2372, N2362);
nor NOR3 (N2373, N2366, N2370, N1827);
nor NOR2 (N2374, N1305, N830);
and AND2 (N2375, N2359, N592);
and AND2 (N2376, N2374, N1703);
and AND2 (N2377, N2369, N97);
not NOT1 (N2378, N2377);
not NOT1 (N2379, N2371);
not NOT1 (N2380, N2361);
not NOT1 (N2381, N2380);
buf BUF1 (N2382, N2378);
nand NAND4 (N2383, N2375, N420, N812, N683);
xor XOR2 (N2384, N2383, N267);
nor NOR2 (N2385, N2365, N304);
not NOT1 (N2386, N2376);
nand NAND2 (N2387, N2381, N1751);
and AND4 (N2388, N2379, N1286, N622, N1449);
nor NOR2 (N2389, N2372, N1134);
nand NAND2 (N2390, N2367, N1663);
nor NOR2 (N2391, N2384, N142);
not NOT1 (N2392, N2387);
nand NAND2 (N2393, N2386, N1166);
nor NOR3 (N2394, N2391, N1445, N969);
and AND2 (N2395, N2390, N1771);
nand NAND4 (N2396, N2385, N1497, N489, N2271);
buf BUF1 (N2397, N2395);
nor NOR2 (N2398, N2389, N70);
and AND2 (N2399, N2394, N574);
xor XOR2 (N2400, N2398, N1010);
or OR3 (N2401, N2373, N1142, N15);
nor NOR3 (N2402, N2397, N1439, N1211);
not NOT1 (N2403, N2402);
nor NOR2 (N2404, N2396, N1210);
and AND2 (N2405, N2400, N1712);
nor NOR3 (N2406, N2382, N2307, N46);
xor XOR2 (N2407, N2405, N387);
not NOT1 (N2408, N2403);
and AND3 (N2409, N2408, N1572, N1651);
nand NAND2 (N2410, N2404, N2262);
nor NOR2 (N2411, N2392, N1948);
and AND2 (N2412, N2407, N734);
or OR2 (N2413, N2411, N592);
nand NAND2 (N2414, N2406, N2147);
and AND4 (N2415, N2413, N1247, N1740, N1341);
nand NAND4 (N2416, N2401, N1703, N1854, N728);
xor XOR2 (N2417, N2393, N177);
nand NAND3 (N2418, N2417, N526, N675);
and AND4 (N2419, N2399, N1697, N949, N663);
xor XOR2 (N2420, N2416, N1117);
nor NOR4 (N2421, N2357, N1771, N2248, N1841);
buf BUF1 (N2422, N2409);
xor XOR2 (N2423, N2414, N636);
nor NOR3 (N2424, N2419, N1416, N585);
or OR4 (N2425, N2421, N223, N2258, N2134);
not NOT1 (N2426, N2422);
and AND3 (N2427, N2425, N393, N2340);
nor NOR2 (N2428, N2423, N965);
xor XOR2 (N2429, N2418, N563);
or OR2 (N2430, N2420, N29);
not NOT1 (N2431, N2412);
or OR4 (N2432, N2410, N1600, N1996, N1795);
or OR4 (N2433, N2431, N726, N212, N1644);
and AND4 (N2434, N2432, N536, N1337, N973);
nor NOR3 (N2435, N2427, N1431, N862);
nand NAND4 (N2436, N2428, N1891, N1438, N1638);
and AND3 (N2437, N2436, N1879, N1916);
buf BUF1 (N2438, N2437);
buf BUF1 (N2439, N2424);
and AND4 (N2440, N2430, N834, N755, N2431);
and AND2 (N2441, N2439, N2371);
nand NAND3 (N2442, N2441, N1941, N517);
or OR4 (N2443, N2415, N2420, N1296, N2279);
buf BUF1 (N2444, N2433);
xor XOR2 (N2445, N2444, N378);
xor XOR2 (N2446, N2435, N2419);
nor NOR3 (N2447, N2446, N1701, N1903);
or OR2 (N2448, N2426, N831);
not NOT1 (N2449, N2438);
nand NAND2 (N2450, N2429, N1917);
nor NOR4 (N2451, N2388, N1816, N1984, N446);
or OR2 (N2452, N2448, N562);
and AND3 (N2453, N2442, N1765, N663);
or OR2 (N2454, N2449, N957);
xor XOR2 (N2455, N2447, N1713);
buf BUF1 (N2456, N2445);
and AND2 (N2457, N2456, N1052);
xor XOR2 (N2458, N2455, N2291);
or OR3 (N2459, N2451, N895, N1505);
nand NAND4 (N2460, N2453, N1436, N1468, N571);
nor NOR2 (N2461, N2457, N550);
nor NOR3 (N2462, N2452, N1372, N2338);
nand NAND3 (N2463, N2459, N1675, N2246);
buf BUF1 (N2464, N2461);
xor XOR2 (N2465, N2462, N1191);
not NOT1 (N2466, N2440);
not NOT1 (N2467, N2458);
xor XOR2 (N2468, N2463, N1235);
nand NAND2 (N2469, N2460, N1659);
xor XOR2 (N2470, N2469, N865);
nor NOR2 (N2471, N2470, N790);
not NOT1 (N2472, N2464);
nand NAND4 (N2473, N2454, N39, N980, N340);
and AND2 (N2474, N2466, N2468);
buf BUF1 (N2475, N1061);
buf BUF1 (N2476, N2465);
nand NAND4 (N2477, N2476, N1892, N2045, N739);
xor XOR2 (N2478, N2471, N906);
and AND4 (N2479, N2467, N158, N1571, N175);
or OR4 (N2480, N2473, N172, N546, N934);
nand NAND3 (N2481, N2443, N1545, N1434);
or OR2 (N2482, N2474, N873);
or OR4 (N2483, N2480, N1134, N1210, N985);
and AND3 (N2484, N2477, N1281, N1287);
or OR3 (N2485, N2484, N94, N167);
xor XOR2 (N2486, N2485, N1875);
not NOT1 (N2487, N2481);
nand NAND2 (N2488, N2450, N1411);
buf BUF1 (N2489, N2488);
nand NAND3 (N2490, N2483, N2477, N1213);
nand NAND4 (N2491, N2490, N615, N2181, N1197);
and AND2 (N2492, N2482, N196);
and AND4 (N2493, N2434, N1738, N1639, N189);
nand NAND3 (N2494, N2486, N2087, N894);
not NOT1 (N2495, N2494);
or OR4 (N2496, N2489, N1521, N194, N1695);
not NOT1 (N2497, N2495);
nand NAND3 (N2498, N2492, N2307, N2095);
xor XOR2 (N2499, N2487, N396);
and AND3 (N2500, N2499, N952, N2135);
nor NOR4 (N2501, N2479, N2395, N127, N1934);
not NOT1 (N2502, N2475);
buf BUF1 (N2503, N2500);
xor XOR2 (N2504, N2472, N2150);
or OR4 (N2505, N2502, N320, N1662, N613);
nand NAND2 (N2506, N2504, N137);
xor XOR2 (N2507, N2478, N386);
buf BUF1 (N2508, N2506);
and AND3 (N2509, N2493, N641, N1498);
or OR3 (N2510, N2498, N1550, N1601);
not NOT1 (N2511, N2505);
or OR4 (N2512, N2511, N530, N1245, N637);
xor XOR2 (N2513, N2507, N423);
and AND4 (N2514, N2496, N1880, N2336, N2340);
or OR3 (N2515, N2508, N424, N501);
nor NOR4 (N2516, N2513, N1476, N408, N2037);
nor NOR3 (N2517, N2501, N1585, N1500);
nand NAND4 (N2518, N2510, N1133, N1504, N1590);
xor XOR2 (N2519, N2518, N2425);
nor NOR2 (N2520, N2515, N1750);
and AND3 (N2521, N2517, N1315, N2219);
buf BUF1 (N2522, N2514);
nand NAND2 (N2523, N2497, N918);
and AND4 (N2524, N2503, N1009, N1891, N453);
buf BUF1 (N2525, N2523);
nor NOR2 (N2526, N2516, N2044);
or OR3 (N2527, N2526, N2398, N746);
or OR3 (N2528, N2524, N1780, N1202);
nor NOR4 (N2529, N2491, N1718, N2025, N1128);
nand NAND3 (N2530, N2522, N446, N2137);
not NOT1 (N2531, N2525);
buf BUF1 (N2532, N2531);
buf BUF1 (N2533, N2529);
buf BUF1 (N2534, N2533);
or OR2 (N2535, N2521, N2500);
nand NAND4 (N2536, N2512, N954, N224, N821);
or OR4 (N2537, N2534, N1718, N2176, N475);
or OR2 (N2538, N2527, N1381);
nor NOR3 (N2539, N2528, N1024, N727);
xor XOR2 (N2540, N2530, N2206);
not NOT1 (N2541, N2537);
nand NAND3 (N2542, N2532, N1890, N621);
buf BUF1 (N2543, N2538);
and AND3 (N2544, N2540, N284, N2159);
nand NAND3 (N2545, N2536, N697, N970);
xor XOR2 (N2546, N2535, N525);
nand NAND4 (N2547, N2544, N2126, N2369, N1853);
nand NAND3 (N2548, N2546, N2524, N2215);
not NOT1 (N2549, N2520);
nor NOR2 (N2550, N2509, N1505);
nand NAND3 (N2551, N2545, N2338, N1283);
not NOT1 (N2552, N2541);
and AND4 (N2553, N2542, N2358, N2370, N238);
or OR4 (N2554, N2519, N860, N276, N1944);
buf BUF1 (N2555, N2548);
xor XOR2 (N2556, N2543, N546);
and AND3 (N2557, N2556, N2177, N749);
not NOT1 (N2558, N2555);
and AND2 (N2559, N2558, N2144);
and AND4 (N2560, N2547, N661, N1623, N53);
nor NOR4 (N2561, N2549, N1829, N822, N135);
nand NAND2 (N2562, N2554, N1988);
xor XOR2 (N2563, N2561, N1268);
and AND2 (N2564, N2552, N2062);
not NOT1 (N2565, N2539);
or OR4 (N2566, N2557, N1071, N1215, N2162);
buf BUF1 (N2567, N2564);
not NOT1 (N2568, N2550);
or OR3 (N2569, N2568, N2136, N888);
nor NOR3 (N2570, N2560, N782, N2295);
or OR4 (N2571, N2566, N1331, N360, N540);
xor XOR2 (N2572, N2563, N2084);
nand NAND4 (N2573, N2570, N1266, N723, N272);
buf BUF1 (N2574, N2571);
nand NAND3 (N2575, N2553, N1970, N535);
or OR4 (N2576, N2573, N1127, N363, N832);
nand NAND3 (N2577, N2551, N648, N1453);
xor XOR2 (N2578, N2559, N1615);
and AND4 (N2579, N2578, N735, N657, N769);
nor NOR3 (N2580, N2574, N316, N1899);
buf BUF1 (N2581, N2565);
xor XOR2 (N2582, N2580, N546);
or OR4 (N2583, N2577, N2397, N1400, N1193);
not NOT1 (N2584, N2579);
not NOT1 (N2585, N2567);
xor XOR2 (N2586, N2575, N892);
nand NAND3 (N2587, N2569, N342, N1371);
not NOT1 (N2588, N2584);
buf BUF1 (N2589, N2587);
buf BUF1 (N2590, N2585);
not NOT1 (N2591, N2590);
nor NOR3 (N2592, N2583, N39, N1424);
not NOT1 (N2593, N2576);
or OR3 (N2594, N2589, N86, N640);
not NOT1 (N2595, N2588);
buf BUF1 (N2596, N2595);
or OR3 (N2597, N2562, N95, N2086);
nand NAND4 (N2598, N2596, N483, N1688, N1394);
and AND3 (N2599, N2581, N1311, N1325);
nor NOR3 (N2600, N2599, N2235, N2198);
buf BUF1 (N2601, N2600);
or OR3 (N2602, N2598, N1622, N2406);
nor NOR2 (N2603, N2586, N2375);
and AND2 (N2604, N2602, N1661);
and AND2 (N2605, N2603, N1374);
nor NOR3 (N2606, N2591, N1621, N1921);
or OR3 (N2607, N2572, N565, N1460);
not NOT1 (N2608, N2597);
nor NOR3 (N2609, N2604, N2400, N409);
nor NOR4 (N2610, N2609, N382, N1511, N1021);
nor NOR2 (N2611, N2605, N2193);
or OR4 (N2612, N2601, N2077, N1215, N1162);
buf BUF1 (N2613, N2593);
nor NOR4 (N2614, N2608, N606, N625, N1769);
or OR2 (N2615, N2594, N946);
or OR4 (N2616, N2613, N2276, N1788, N651);
and AND2 (N2617, N2607, N1628);
and AND3 (N2618, N2611, N1688, N2298);
and AND3 (N2619, N2618, N2251, N1316);
buf BUF1 (N2620, N2592);
or OR3 (N2621, N2612, N904, N595);
nor NOR4 (N2622, N2582, N1218, N1980, N1122);
not NOT1 (N2623, N2616);
buf BUF1 (N2624, N2622);
or OR4 (N2625, N2606, N1042, N2068, N1418);
and AND2 (N2626, N2623, N1986);
and AND2 (N2627, N2617, N1553);
nor NOR4 (N2628, N2626, N582, N1308, N1817);
xor XOR2 (N2629, N2620, N764);
buf BUF1 (N2630, N2615);
nand NAND3 (N2631, N2610, N2356, N1373);
nand NAND3 (N2632, N2628, N1579, N1805);
and AND4 (N2633, N2614, N2119, N1585, N555);
not NOT1 (N2634, N2625);
nand NAND4 (N2635, N2634, N792, N2521, N1976);
or OR3 (N2636, N2621, N262, N1279);
buf BUF1 (N2637, N2633);
buf BUF1 (N2638, N2631);
nor NOR2 (N2639, N2636, N1730);
xor XOR2 (N2640, N2624, N33);
xor XOR2 (N2641, N2635, N1307);
or OR3 (N2642, N2629, N1461, N1784);
nor NOR4 (N2643, N2640, N407, N1541, N1979);
or OR2 (N2644, N2638, N2021);
or OR2 (N2645, N2643, N1042);
or OR4 (N2646, N2632, N1339, N1325, N852);
and AND2 (N2647, N2642, N436);
or OR4 (N2648, N2637, N106, N2222, N833);
buf BUF1 (N2649, N2619);
buf BUF1 (N2650, N2649);
nand NAND2 (N2651, N2644, N876);
or OR4 (N2652, N2645, N1304, N1246, N2115);
buf BUF1 (N2653, N2646);
and AND3 (N2654, N2630, N368, N279);
buf BUF1 (N2655, N2648);
buf BUF1 (N2656, N2627);
and AND2 (N2657, N2656, N684);
nand NAND3 (N2658, N2657, N2173, N1793);
xor XOR2 (N2659, N2641, N2057);
xor XOR2 (N2660, N2655, N1798);
nand NAND2 (N2661, N2639, N2593);
buf BUF1 (N2662, N2653);
xor XOR2 (N2663, N2659, N1899);
buf BUF1 (N2664, N2663);
nor NOR2 (N2665, N2662, N1462);
buf BUF1 (N2666, N2661);
nand NAND2 (N2667, N2647, N2142);
nor NOR3 (N2668, N2651, N864, N1087);
not NOT1 (N2669, N2652);
or OR4 (N2670, N2658, N1636, N1288, N1032);
and AND2 (N2671, N2668, N686);
nor NOR3 (N2672, N2670, N204, N2093);
or OR3 (N2673, N2672, N414, N1206);
xor XOR2 (N2674, N2666, N1217);
nand NAND2 (N2675, N2669, N919);
or OR2 (N2676, N2675, N1669);
not NOT1 (N2677, N2673);
not NOT1 (N2678, N2674);
nand NAND4 (N2679, N2677, N1458, N2364, N2198);
not NOT1 (N2680, N2650);
nor NOR3 (N2681, N2660, N1398, N2358);
nand NAND4 (N2682, N2676, N820, N1857, N810);
nand NAND2 (N2683, N2654, N2564);
nand NAND2 (N2684, N2679, N1836);
nor NOR2 (N2685, N2682, N1194);
and AND4 (N2686, N2667, N1336, N833, N2051);
xor XOR2 (N2687, N2680, N1549);
not NOT1 (N2688, N2685);
buf BUF1 (N2689, N2686);
nand NAND3 (N2690, N2683, N928, N348);
or OR3 (N2691, N2664, N92, N351);
or OR4 (N2692, N2689, N1155, N1048, N463);
and AND4 (N2693, N2687, N1555, N2494, N50);
xor XOR2 (N2694, N2692, N695);
and AND4 (N2695, N2688, N874, N2686, N1604);
buf BUF1 (N2696, N2691);
or OR4 (N2697, N2694, N1044, N151, N2542);
xor XOR2 (N2698, N2696, N1308);
or OR2 (N2699, N2697, N1402);
nand NAND2 (N2700, N2678, N1080);
or OR3 (N2701, N2699, N2408, N979);
buf BUF1 (N2702, N2665);
nand NAND3 (N2703, N2700, N2576, N110);
buf BUF1 (N2704, N2671);
buf BUF1 (N2705, N2695);
or OR3 (N2706, N2690, N2450, N61);
not NOT1 (N2707, N2706);
buf BUF1 (N2708, N2698);
and AND3 (N2709, N2708, N2419, N1198);
nor NOR2 (N2710, N2684, N566);
or OR2 (N2711, N2701, N1454);
or OR4 (N2712, N2704, N329, N1029, N2232);
not NOT1 (N2713, N2707);
nor NOR4 (N2714, N2693, N1440, N1736, N20);
and AND2 (N2715, N2714, N851);
xor XOR2 (N2716, N2705, N880);
nand NAND4 (N2717, N2716, N2203, N698, N1004);
and AND2 (N2718, N2711, N168);
nand NAND2 (N2719, N2710, N2237);
not NOT1 (N2720, N2702);
xor XOR2 (N2721, N2717, N2212);
and AND4 (N2722, N2721, N792, N2379, N372);
not NOT1 (N2723, N2720);
buf BUF1 (N2724, N2723);
and AND2 (N2725, N2703, N1519);
or OR3 (N2726, N2713, N1784, N78);
nor NOR3 (N2727, N2712, N8, N2454);
nor NOR3 (N2728, N2715, N2149, N1581);
xor XOR2 (N2729, N2724, N2064);
xor XOR2 (N2730, N2719, N1028);
or OR4 (N2731, N2709, N1499, N542, N2053);
buf BUF1 (N2732, N2728);
nand NAND3 (N2733, N2729, N2356, N1830);
not NOT1 (N2734, N2681);
and AND2 (N2735, N2726, N2176);
buf BUF1 (N2736, N2731);
buf BUF1 (N2737, N2734);
or OR3 (N2738, N2735, N861, N2445);
nand NAND2 (N2739, N2737, N945);
nand NAND2 (N2740, N2718, N1052);
not NOT1 (N2741, N2732);
nand NAND2 (N2742, N2739, N1622);
or OR3 (N2743, N2736, N958, N1308);
xor XOR2 (N2744, N2725, N792);
xor XOR2 (N2745, N2722, N660);
or OR3 (N2746, N2741, N2497, N2711);
nor NOR3 (N2747, N2740, N1594, N2447);
nor NOR2 (N2748, N2730, N2077);
buf BUF1 (N2749, N2747);
xor XOR2 (N2750, N2744, N2269);
nor NOR2 (N2751, N2749, N1424);
nor NOR3 (N2752, N2751, N2352, N2486);
nor NOR2 (N2753, N2743, N2448);
or OR4 (N2754, N2742, N2474, N2367, N38);
nor NOR4 (N2755, N2745, N2545, N1854, N983);
or OR3 (N2756, N2738, N1231, N159);
buf BUF1 (N2757, N2733);
xor XOR2 (N2758, N2753, N340);
buf BUF1 (N2759, N2758);
nor NOR3 (N2760, N2746, N1036, N1600);
and AND2 (N2761, N2756, N1730);
nor NOR2 (N2762, N2752, N1125);
nand NAND2 (N2763, N2748, N432);
not NOT1 (N2764, N2754);
and AND3 (N2765, N2755, N912, N1676);
and AND3 (N2766, N2764, N2646, N1038);
nand NAND3 (N2767, N2762, N1672, N160);
nand NAND4 (N2768, N2761, N502, N2633, N1697);
and AND4 (N2769, N2759, N265, N546, N475);
buf BUF1 (N2770, N2757);
not NOT1 (N2771, N2769);
xor XOR2 (N2772, N2765, N472);
nand NAND2 (N2773, N2767, N2170);
nor NOR4 (N2774, N2770, N1164, N1335, N2769);
or OR3 (N2775, N2763, N1802, N1050);
and AND4 (N2776, N2750, N1273, N1531, N862);
buf BUF1 (N2777, N2776);
not NOT1 (N2778, N2773);
xor XOR2 (N2779, N2775, N850);
not NOT1 (N2780, N2778);
nand NAND3 (N2781, N2774, N582, N1972);
not NOT1 (N2782, N2779);
nand NAND3 (N2783, N2782, N656, N1549);
xor XOR2 (N2784, N2780, N1325);
buf BUF1 (N2785, N2783);
nor NOR3 (N2786, N2727, N2011, N497);
or OR3 (N2787, N2786, N2512, N175);
or OR2 (N2788, N2777, N1966);
or OR3 (N2789, N2788, N152, N2690);
xor XOR2 (N2790, N2784, N2750);
not NOT1 (N2791, N2790);
buf BUF1 (N2792, N2789);
nand NAND3 (N2793, N2787, N2088, N1116);
not NOT1 (N2794, N2791);
not NOT1 (N2795, N2794);
buf BUF1 (N2796, N2795);
or OR3 (N2797, N2781, N110, N2677);
and AND2 (N2798, N2797, N2678);
and AND3 (N2799, N2792, N1590, N2414);
buf BUF1 (N2800, N2760);
buf BUF1 (N2801, N2771);
and AND3 (N2802, N2800, N2326, N580);
and AND4 (N2803, N2796, N287, N50, N1292);
nand NAND3 (N2804, N2803, N1224, N2588);
buf BUF1 (N2805, N2799);
xor XOR2 (N2806, N2768, N159);
and AND2 (N2807, N2793, N899);
and AND4 (N2808, N2798, N1704, N1590, N1);
and AND3 (N2809, N2766, N694, N465);
buf BUF1 (N2810, N2772);
nand NAND3 (N2811, N2804, N1408, N412);
xor XOR2 (N2812, N2806, N797);
xor XOR2 (N2813, N2810, N1869);
nand NAND2 (N2814, N2807, N1311);
or OR3 (N2815, N2814, N807, N1475);
buf BUF1 (N2816, N2785);
not NOT1 (N2817, N2813);
and AND2 (N2818, N2817, N29);
nand NAND2 (N2819, N2811, N222);
or OR4 (N2820, N2805, N584, N1114, N194);
not NOT1 (N2821, N2808);
buf BUF1 (N2822, N2812);
xor XOR2 (N2823, N2818, N1412);
xor XOR2 (N2824, N2819, N937);
or OR3 (N2825, N2802, N1873, N2065);
nand NAND3 (N2826, N2822, N2526, N2013);
buf BUF1 (N2827, N2823);
xor XOR2 (N2828, N2816, N42);
xor XOR2 (N2829, N2820, N953);
and AND4 (N2830, N2828, N2214, N943, N1234);
xor XOR2 (N2831, N2829, N2766);
not NOT1 (N2832, N2825);
xor XOR2 (N2833, N2815, N1770);
and AND3 (N2834, N2821, N877, N2138);
and AND4 (N2835, N2833, N1537, N37, N1665);
not NOT1 (N2836, N2831);
nor NOR2 (N2837, N2809, N1480);
or OR2 (N2838, N2830, N268);
and AND3 (N2839, N2835, N1287, N2705);
nand NAND3 (N2840, N2839, N1665, N167);
buf BUF1 (N2841, N2827);
xor XOR2 (N2842, N2824, N1433);
and AND2 (N2843, N2836, N2718);
not NOT1 (N2844, N2843);
nor NOR2 (N2845, N2838, N310);
or OR4 (N2846, N2837, N2016, N70, N2082);
nor NOR2 (N2847, N2826, N1362);
nand NAND2 (N2848, N2847, N2762);
or OR4 (N2849, N2845, N1302, N2585, N716);
xor XOR2 (N2850, N2801, N2558);
buf BUF1 (N2851, N2850);
or OR2 (N2852, N2846, N956);
nor NOR4 (N2853, N2852, N1092, N2101, N1934);
and AND2 (N2854, N2834, N165);
nand NAND3 (N2855, N2841, N1583, N596);
not NOT1 (N2856, N2842);
nor NOR2 (N2857, N2856, N942);
and AND4 (N2858, N2853, N1658, N1026, N1329);
xor XOR2 (N2859, N2844, N431);
and AND3 (N2860, N2855, N128, N2669);
nor NOR3 (N2861, N2859, N992, N1111);
and AND3 (N2862, N2851, N2516, N217);
or OR2 (N2863, N2861, N818);
nand NAND4 (N2864, N2849, N682, N1081, N42);
or OR3 (N2865, N2857, N758, N960);
or OR2 (N2866, N2848, N2426);
xor XOR2 (N2867, N2865, N2447);
not NOT1 (N2868, N2858);
nand NAND2 (N2869, N2863, N1780);
buf BUF1 (N2870, N2864);
or OR3 (N2871, N2860, N998, N2120);
not NOT1 (N2872, N2840);
and AND4 (N2873, N2869, N629, N2571, N888);
and AND2 (N2874, N2832, N1607);
nor NOR3 (N2875, N2872, N2391, N2773);
not NOT1 (N2876, N2868);
or OR3 (N2877, N2866, N1253, N1248);
not NOT1 (N2878, N2874);
nor NOR4 (N2879, N2877, N2377, N229, N805);
nor NOR4 (N2880, N2854, N317, N87, N1364);
nand NAND3 (N2881, N2870, N2129, N1334);
nor NOR3 (N2882, N2880, N2299, N2637);
buf BUF1 (N2883, N2876);
nand NAND4 (N2884, N2882, N2065, N2329, N1158);
buf BUF1 (N2885, N2879);
not NOT1 (N2886, N2881);
or OR3 (N2887, N2884, N802, N469);
xor XOR2 (N2888, N2871, N2395);
not NOT1 (N2889, N2887);
nand NAND3 (N2890, N2867, N1636, N606);
xor XOR2 (N2891, N2873, N340);
not NOT1 (N2892, N2885);
buf BUF1 (N2893, N2875);
buf BUF1 (N2894, N2886);
nand NAND4 (N2895, N2891, N2232, N135, N407);
not NOT1 (N2896, N2888);
or OR3 (N2897, N2883, N583, N2050);
buf BUF1 (N2898, N2890);
buf BUF1 (N2899, N2897);
nor NOR2 (N2900, N2878, N1657);
or OR3 (N2901, N2896, N2260, N2042);
and AND4 (N2902, N2895, N364, N2872, N559);
and AND3 (N2903, N2889, N2671, N2647);
nand NAND2 (N2904, N2901, N577);
xor XOR2 (N2905, N2898, N1152);
xor XOR2 (N2906, N2862, N1726);
buf BUF1 (N2907, N2902);
buf BUF1 (N2908, N2893);
nor NOR3 (N2909, N2903, N1830, N1696);
or OR2 (N2910, N2894, N2001);
nor NOR3 (N2911, N2892, N2522, N1011);
buf BUF1 (N2912, N2905);
not NOT1 (N2913, N2908);
or OR3 (N2914, N2911, N2720, N2321);
or OR4 (N2915, N2909, N1113, N1726, N1406);
nor NOR3 (N2916, N2914, N2909, N290);
xor XOR2 (N2917, N2906, N2423);
nor NOR2 (N2918, N2900, N2384);
and AND2 (N2919, N2917, N1520);
xor XOR2 (N2920, N2899, N360);
or OR3 (N2921, N2904, N1707, N1617);
or OR2 (N2922, N2916, N2184);
xor XOR2 (N2923, N2920, N2276);
not NOT1 (N2924, N2919);
nand NAND3 (N2925, N2922, N842, N1458);
nor NOR2 (N2926, N2921, N2174);
buf BUF1 (N2927, N2918);
or OR2 (N2928, N2907, N2347);
xor XOR2 (N2929, N2928, N1219);
and AND3 (N2930, N2925, N1249, N859);
nand NAND3 (N2931, N2929, N570, N824);
and AND3 (N2932, N2915, N1276, N2335);
or OR4 (N2933, N2924, N1644, N1393, N1622);
nor NOR4 (N2934, N2926, N121, N875, N2626);
nand NAND4 (N2935, N2923, N2422, N2796, N1845);
nor NOR3 (N2936, N2912, N1379, N512);
or OR3 (N2937, N2931, N2796, N25);
buf BUF1 (N2938, N2937);
nand NAND2 (N2939, N2938, N2887);
xor XOR2 (N2940, N2935, N947);
and AND3 (N2941, N2910, N1666, N2096);
and AND4 (N2942, N2939, N2642, N2681, N1937);
nor NOR3 (N2943, N2940, N231, N1110);
xor XOR2 (N2944, N2932, N1162);
xor XOR2 (N2945, N2942, N1037);
xor XOR2 (N2946, N2930, N2844);
or OR2 (N2947, N2913, N299);
or OR3 (N2948, N2927, N645, N1509);
and AND3 (N2949, N2941, N1980, N2142);
or OR2 (N2950, N2933, N2184);
nor NOR4 (N2951, N2949, N1016, N435, N2124);
and AND4 (N2952, N2936, N242, N2249, N1013);
buf BUF1 (N2953, N2934);
xor XOR2 (N2954, N2943, N937);
not NOT1 (N2955, N2948);
buf BUF1 (N2956, N2951);
buf BUF1 (N2957, N2954);
not NOT1 (N2958, N2952);
xor XOR2 (N2959, N2947, N1634);
nand NAND2 (N2960, N2950, N1633);
nand NAND2 (N2961, N2956, N2531);
nand NAND4 (N2962, N2944, N2468, N936, N188);
xor XOR2 (N2963, N2946, N129);
nor NOR4 (N2964, N2962, N2733, N2835, N2459);
xor XOR2 (N2965, N2963, N417);
and AND3 (N2966, N2959, N509, N737);
nand NAND4 (N2967, N2955, N1745, N2613, N1678);
buf BUF1 (N2968, N2960);
not NOT1 (N2969, N2967);
nor NOR4 (N2970, N2961, N731, N2594, N218);
or OR4 (N2971, N2965, N500, N977, N2184);
and AND4 (N2972, N2971, N2341, N1259, N2144);
or OR2 (N2973, N2970, N226);
nor NOR3 (N2974, N2958, N2432, N170);
and AND4 (N2975, N2973, N1055, N1335, N926);
nor NOR4 (N2976, N2972, N2498, N1603, N2010);
xor XOR2 (N2977, N2966, N2382);
xor XOR2 (N2978, N2968, N1465);
and AND2 (N2979, N2974, N286);
not NOT1 (N2980, N2977);
or OR3 (N2981, N2953, N1799, N1870);
not NOT1 (N2982, N2945);
buf BUF1 (N2983, N2978);
xor XOR2 (N2984, N2964, N331);
nor NOR4 (N2985, N2975, N1123, N2013, N2644);
nor NOR3 (N2986, N2981, N427, N1421);
or OR2 (N2987, N2986, N1378);
xor XOR2 (N2988, N2969, N93);
not NOT1 (N2989, N2984);
or OR4 (N2990, N2983, N2817, N40, N1773);
not NOT1 (N2991, N2979);
not NOT1 (N2992, N2991);
not NOT1 (N2993, N2980);
or OR4 (N2994, N2988, N935, N2330, N856);
not NOT1 (N2995, N2990);
not NOT1 (N2996, N2993);
nand NAND3 (N2997, N2957, N2239, N1829);
xor XOR2 (N2998, N2995, N37);
or OR2 (N2999, N2989, N763);
or OR3 (N3000, N2985, N2878, N1367);
nand NAND2 (N3001, N2987, N2458);
and AND3 (N3002, N2982, N619, N422);
and AND2 (N3003, N3000, N1341);
nor NOR4 (N3004, N2997, N144, N1760, N1036);
not NOT1 (N3005, N2992);
and AND2 (N3006, N2998, N1795);
and AND3 (N3007, N2999, N292, N391);
not NOT1 (N3008, N3007);
and AND3 (N3009, N3005, N68, N2176);
nand NAND3 (N3010, N3009, N2265, N2332);
nand NAND2 (N3011, N3001, N1174);
nor NOR3 (N3012, N3008, N631, N1856);
and AND4 (N3013, N3002, N1749, N1502, N3001);
xor XOR2 (N3014, N3012, N2760);
nand NAND2 (N3015, N2996, N371);
nand NAND4 (N3016, N3003, N1545, N1940, N694);
xor XOR2 (N3017, N3015, N144);
and AND4 (N3018, N2976, N1965, N2844, N2313);
not NOT1 (N3019, N3006);
and AND2 (N3020, N3016, N169);
not NOT1 (N3021, N3020);
and AND4 (N3022, N3019, N1251, N1750, N1914);
not NOT1 (N3023, N2994);
nor NOR4 (N3024, N3010, N2278, N363, N1597);
not NOT1 (N3025, N3021);
xor XOR2 (N3026, N3004, N191);
not NOT1 (N3027, N3018);
nand NAND2 (N3028, N3023, N1904);
not NOT1 (N3029, N3013);
buf BUF1 (N3030, N3011);
and AND3 (N3031, N3028, N371, N788);
or OR4 (N3032, N3026, N2241, N1181, N2298);
xor XOR2 (N3033, N3032, N1133);
or OR2 (N3034, N3014, N1377);
not NOT1 (N3035, N3017);
nor NOR2 (N3036, N3027, N2440);
buf BUF1 (N3037, N3024);
nand NAND2 (N3038, N3036, N2833);
or OR3 (N3039, N3025, N2635, N2080);
not NOT1 (N3040, N3039);
nor NOR2 (N3041, N3035, N2995);
xor XOR2 (N3042, N3041, N2346);
xor XOR2 (N3043, N3030, N839);
xor XOR2 (N3044, N3040, N41);
buf BUF1 (N3045, N3034);
or OR3 (N3046, N3037, N458, N943);
xor XOR2 (N3047, N3031, N2547);
nand NAND3 (N3048, N3033, N2259, N1489);
nand NAND3 (N3049, N3042, N2203, N2576);
nor NOR2 (N3050, N3044, N2751);
nand NAND3 (N3051, N3043, N2434, N623);
nor NOR3 (N3052, N3038, N83, N2835);
not NOT1 (N3053, N3048);
and AND4 (N3054, N3052, N1619, N1994, N2900);
xor XOR2 (N3055, N3047, N1859);
or OR3 (N3056, N3050, N186, N3025);
or OR2 (N3057, N3029, N1891);
nand NAND2 (N3058, N3057, N2141);
nand NAND3 (N3059, N3055, N2272, N152);
nor NOR2 (N3060, N3049, N1035);
nand NAND2 (N3061, N3053, N209);
xor XOR2 (N3062, N3054, N1755);
nand NAND3 (N3063, N3046, N874, N1143);
nor NOR4 (N3064, N3060, N1319, N2425, N2996);
or OR4 (N3065, N3058, N2253, N3015, N1401);
and AND2 (N3066, N3062, N261);
or OR2 (N3067, N3064, N886);
and AND3 (N3068, N3063, N936, N2354);
nor NOR2 (N3069, N3065, N1989);
nand NAND2 (N3070, N3067, N76);
xor XOR2 (N3071, N3045, N2270);
or OR4 (N3072, N3068, N1481, N2988, N922);
and AND2 (N3073, N3051, N2726);
nor NOR2 (N3074, N3073, N2292);
buf BUF1 (N3075, N3069);
not NOT1 (N3076, N3022);
nor NOR4 (N3077, N3070, N2813, N1263, N483);
or OR4 (N3078, N3071, N1461, N839, N1903);
and AND2 (N3079, N3066, N602);
nor NOR2 (N3080, N3076, N597);
nor NOR3 (N3081, N3072, N2383, N756);
nand NAND2 (N3082, N3081, N567);
xor XOR2 (N3083, N3056, N1387);
not NOT1 (N3084, N3079);
and AND2 (N3085, N3082, N836);
buf BUF1 (N3086, N3085);
nor NOR2 (N3087, N3078, N3064);
nor NOR2 (N3088, N3087, N2752);
not NOT1 (N3089, N3080);
xor XOR2 (N3090, N3084, N2493);
not NOT1 (N3091, N3086);
not NOT1 (N3092, N3090);
and AND3 (N3093, N3074, N1876, N2683);
xor XOR2 (N3094, N3075, N1305);
nand NAND2 (N3095, N3093, N128);
buf BUF1 (N3096, N3095);
xor XOR2 (N3097, N3077, N1244);
buf BUF1 (N3098, N3061);
or OR2 (N3099, N3098, N897);
nor NOR3 (N3100, N3088, N2900, N1686);
or OR3 (N3101, N3092, N1475, N1185);
buf BUF1 (N3102, N3101);
buf BUF1 (N3103, N3094);
nor NOR2 (N3104, N3059, N6);
nand NAND3 (N3105, N3091, N1530, N1373);
nor NOR4 (N3106, N3099, N658, N2753, N922);
and AND2 (N3107, N3102, N1714);
or OR2 (N3108, N3105, N2383);
xor XOR2 (N3109, N3107, N903);
xor XOR2 (N3110, N3103, N579);
and AND3 (N3111, N3110, N2903, N81);
buf BUF1 (N3112, N3108);
not NOT1 (N3113, N3100);
buf BUF1 (N3114, N3083);
buf BUF1 (N3115, N3113);
and AND3 (N3116, N3109, N1599, N1418);
nor NOR3 (N3117, N3096, N1087, N2642);
and AND2 (N3118, N3089, N270);
buf BUF1 (N3119, N3117);
buf BUF1 (N3120, N3111);
buf BUF1 (N3121, N3114);
and AND2 (N3122, N3106, N2448);
nor NOR4 (N3123, N3097, N3067, N1365, N2371);
buf BUF1 (N3124, N3119);
not NOT1 (N3125, N3122);
or OR3 (N3126, N3120, N2079, N605);
or OR3 (N3127, N3116, N1675, N646);
xor XOR2 (N3128, N3125, N2165);
nor NOR2 (N3129, N3112, N1682);
nand NAND3 (N3130, N3115, N2071, N1062);
nor NOR4 (N3131, N3124, N3118, N1325, N1400);
and AND2 (N3132, N1668, N493);
xor XOR2 (N3133, N3129, N145);
or OR2 (N3134, N3128, N2013);
and AND3 (N3135, N3104, N2880, N974);
and AND2 (N3136, N3126, N788);
nand NAND4 (N3137, N3131, N2734, N3127, N2852);
buf BUF1 (N3138, N1113);
nand NAND4 (N3139, N3136, N158, N1759, N2843);
nand NAND3 (N3140, N3121, N2359, N2242);
and AND3 (N3141, N3130, N2092, N3033);
buf BUF1 (N3142, N3134);
nand NAND3 (N3143, N3135, N834, N36);
and AND4 (N3144, N3143, N2138, N2046, N2586);
nor NOR2 (N3145, N3133, N1448);
buf BUF1 (N3146, N3123);
nor NOR4 (N3147, N3142, N2121, N1979, N2883);
or OR3 (N3148, N3144, N2707, N1591);
buf BUF1 (N3149, N3145);
buf BUF1 (N3150, N3132);
or OR2 (N3151, N3137, N1813);
nor NOR3 (N3152, N3149, N991, N2831);
not NOT1 (N3153, N3150);
not NOT1 (N3154, N3139);
nor NOR4 (N3155, N3138, N2109, N215, N3051);
or OR4 (N3156, N3141, N11, N494, N2122);
buf BUF1 (N3157, N3156);
not NOT1 (N3158, N3140);
nand NAND3 (N3159, N3147, N66, N1047);
xor XOR2 (N3160, N3159, N546);
xor XOR2 (N3161, N3158, N901);
nand NAND4 (N3162, N3155, N1157, N726, N2286);
nor NOR4 (N3163, N3153, N2228, N1280, N1842);
not NOT1 (N3164, N3157);
nand NAND4 (N3165, N3146, N339, N2777, N1252);
not NOT1 (N3166, N3165);
nand NAND3 (N3167, N3164, N52, N2835);
buf BUF1 (N3168, N3162);
nor NOR3 (N3169, N3154, N1441, N520);
buf BUF1 (N3170, N3161);
or OR4 (N3171, N3160, N1586, N2449, N1317);
nand NAND4 (N3172, N3168, N2123, N2392, N1703);
buf BUF1 (N3173, N3169);
nor NOR3 (N3174, N3170, N1644, N1705);
buf BUF1 (N3175, N3172);
nor NOR2 (N3176, N3166, N2428);
nand NAND3 (N3177, N3148, N2477, N527);
nand NAND4 (N3178, N3175, N2101, N1887, N922);
or OR3 (N3179, N3178, N2643, N198);
or OR4 (N3180, N3151, N676, N1175, N796);
buf BUF1 (N3181, N3177);
not NOT1 (N3182, N3173);
xor XOR2 (N3183, N3179, N107);
or OR2 (N3184, N3174, N3142);
buf BUF1 (N3185, N3184);
nor NOR4 (N3186, N3185, N2867, N2480, N1020);
buf BUF1 (N3187, N3183);
or OR2 (N3188, N3180, N2643);
nor NOR4 (N3189, N3186, N654, N2748, N1536);
xor XOR2 (N3190, N3182, N986);
or OR4 (N3191, N3187, N1105, N1611, N3104);
not NOT1 (N3192, N3176);
or OR2 (N3193, N3189, N3148);
buf BUF1 (N3194, N3190);
or OR2 (N3195, N3188, N1643);
or OR2 (N3196, N3167, N969);
buf BUF1 (N3197, N3194);
or OR4 (N3198, N3152, N181, N1650, N2370);
not NOT1 (N3199, N3163);
and AND3 (N3200, N3199, N1250, N1762);
not NOT1 (N3201, N3171);
and AND4 (N3202, N3193, N1672, N2989, N417);
buf BUF1 (N3203, N3198);
xor XOR2 (N3204, N3197, N68);
not NOT1 (N3205, N3191);
nand NAND3 (N3206, N3202, N964, N2398);
or OR2 (N3207, N3196, N632);
nor NOR4 (N3208, N3207, N3068, N3165, N40);
nor NOR3 (N3209, N3204, N2510, N1063);
xor XOR2 (N3210, N3203, N1046);
or OR3 (N3211, N3201, N3068, N2870);
not NOT1 (N3212, N3208);
nand NAND3 (N3213, N3205, N2538, N2020);
xor XOR2 (N3214, N3209, N2910);
not NOT1 (N3215, N3195);
nand NAND2 (N3216, N3181, N2893);
or OR3 (N3217, N3215, N2872, N2714);
buf BUF1 (N3218, N3213);
nor NOR4 (N3219, N3214, N232, N3138, N2996);
nor NOR3 (N3220, N3210, N2670, N2943);
nor NOR3 (N3221, N3218, N24, N2426);
nor NOR3 (N3222, N3211, N1736, N974);
nand NAND4 (N3223, N3220, N2736, N1893, N1703);
xor XOR2 (N3224, N3217, N1482);
or OR2 (N3225, N3222, N1779);
xor XOR2 (N3226, N3200, N2805);
and AND3 (N3227, N3224, N1495, N1115);
buf BUF1 (N3228, N3221);
and AND4 (N3229, N3212, N950, N1815, N3015);
xor XOR2 (N3230, N3223, N3046);
buf BUF1 (N3231, N3216);
nand NAND3 (N3232, N3230, N1512, N2576);
nand NAND3 (N3233, N3231, N2946, N990);
and AND4 (N3234, N3233, N381, N893, N2773);
not NOT1 (N3235, N3232);
xor XOR2 (N3236, N3192, N2788);
and AND4 (N3237, N3225, N1988, N560, N754);
nand NAND3 (N3238, N3228, N2894, N3003);
and AND4 (N3239, N3236, N1068, N1361, N2523);
and AND3 (N3240, N3234, N2141, N659);
or OR4 (N3241, N3237, N2064, N1367, N3040);
not NOT1 (N3242, N3206);
buf BUF1 (N3243, N3240);
xor XOR2 (N3244, N3238, N545);
buf BUF1 (N3245, N3243);
xor XOR2 (N3246, N3226, N1306);
xor XOR2 (N3247, N3239, N2370);
or OR4 (N3248, N3235, N772, N1204, N1461);
not NOT1 (N3249, N3241);
or OR2 (N3250, N3247, N1931);
nand NAND3 (N3251, N3229, N1753, N3108);
xor XOR2 (N3252, N3249, N2486);
xor XOR2 (N3253, N3227, N549);
nor NOR4 (N3254, N3246, N974, N2110, N1197);
xor XOR2 (N3255, N3251, N852);
and AND4 (N3256, N3253, N837, N1176, N2737);
xor XOR2 (N3257, N3219, N968);
nor NOR4 (N3258, N3252, N1329, N2757, N1148);
nand NAND2 (N3259, N3256, N2941);
nor NOR4 (N3260, N3254, N2152, N2701, N442);
and AND4 (N3261, N3257, N1926, N2802, N1683);
nor NOR2 (N3262, N3259, N3128);
nor NOR4 (N3263, N3262, N1183, N888, N3169);
and AND3 (N3264, N3244, N148, N2271);
not NOT1 (N3265, N3255);
xor XOR2 (N3266, N3242, N2640);
buf BUF1 (N3267, N3261);
or OR2 (N3268, N3260, N1718);
nor NOR3 (N3269, N3250, N408, N684);
nand NAND2 (N3270, N3264, N1770);
xor XOR2 (N3271, N3245, N1918);
xor XOR2 (N3272, N3248, N1153);
buf BUF1 (N3273, N3263);
or OR2 (N3274, N3268, N521);
or OR2 (N3275, N3266, N2277);
buf BUF1 (N3276, N3265);
not NOT1 (N3277, N3275);
nor NOR2 (N3278, N3274, N2331);
nor NOR2 (N3279, N3278, N739);
nor NOR4 (N3280, N3267, N2081, N1366, N1094);
not NOT1 (N3281, N3270);
nor NOR2 (N3282, N3276, N869);
xor XOR2 (N3283, N3281, N2065);
and AND4 (N3284, N3258, N1993, N2596, N2890);
nand NAND3 (N3285, N3284, N122, N1839);
buf BUF1 (N3286, N3272);
and AND2 (N3287, N3273, N1060);
nor NOR3 (N3288, N3279, N1298, N1471);
and AND4 (N3289, N3282, N236, N3263, N1636);
not NOT1 (N3290, N3289);
buf BUF1 (N3291, N3269);
xor XOR2 (N3292, N3286, N2505);
not NOT1 (N3293, N3290);
nor NOR2 (N3294, N3277, N3146);
or OR4 (N3295, N3285, N968, N3146, N2853);
buf BUF1 (N3296, N3287);
not NOT1 (N3297, N3295);
nor NOR3 (N3298, N3293, N3012, N2302);
and AND2 (N3299, N3298, N2679);
xor XOR2 (N3300, N3288, N1747);
xor XOR2 (N3301, N3292, N2714);
not NOT1 (N3302, N3294);
and AND3 (N3303, N3296, N934, N352);
nand NAND4 (N3304, N3280, N1613, N1936, N1268);
and AND2 (N3305, N3300, N2305);
nor NOR3 (N3306, N3297, N552, N241);
buf BUF1 (N3307, N3283);
not NOT1 (N3308, N3299);
nor NOR3 (N3309, N3271, N2610, N1684);
not NOT1 (N3310, N3304);
buf BUF1 (N3311, N3302);
buf BUF1 (N3312, N3309);
and AND3 (N3313, N3310, N1850, N45);
not NOT1 (N3314, N3306);
not NOT1 (N3315, N3307);
nand NAND2 (N3316, N3312, N1050);
nand NAND4 (N3317, N3311, N1008, N172, N1795);
not NOT1 (N3318, N3301);
nand NAND3 (N3319, N3318, N1919, N41);
nor NOR4 (N3320, N3319, N2163, N1224, N754);
not NOT1 (N3321, N3313);
and AND2 (N3322, N3303, N2886);
or OR2 (N3323, N3305, N3116);
not NOT1 (N3324, N3291);
nand NAND2 (N3325, N3322, N1183);
nand NAND4 (N3326, N3321, N2618, N1233, N2462);
xor XOR2 (N3327, N3325, N422);
not NOT1 (N3328, N3324);
buf BUF1 (N3329, N3326);
xor XOR2 (N3330, N3317, N3185);
buf BUF1 (N3331, N3328);
not NOT1 (N3332, N3314);
not NOT1 (N3333, N3329);
nand NAND4 (N3334, N3327, N1561, N221, N182);
buf BUF1 (N3335, N3330);
and AND4 (N3336, N3333, N1536, N803, N3219);
and AND2 (N3337, N3308, N3287);
xor XOR2 (N3338, N3337, N193);
and AND3 (N3339, N3336, N1874, N1276);
nand NAND4 (N3340, N3316, N2474, N1433, N51);
buf BUF1 (N3341, N3320);
not NOT1 (N3342, N3332);
or OR3 (N3343, N3339, N1932, N1604);
xor XOR2 (N3344, N3334, N59);
nand NAND2 (N3345, N3342, N2216);
and AND3 (N3346, N3341, N1052, N1818);
xor XOR2 (N3347, N3340, N594);
nor NOR2 (N3348, N3315, N3040);
and AND2 (N3349, N3347, N1393);
not NOT1 (N3350, N3323);
buf BUF1 (N3351, N3331);
and AND3 (N3352, N3351, N2968, N3116);
or OR4 (N3353, N3343, N3210, N2714, N1919);
buf BUF1 (N3354, N3335);
and AND2 (N3355, N3353, N400);
nor NOR2 (N3356, N3352, N10);
and AND4 (N3357, N3344, N1388, N1113, N1805);
not NOT1 (N3358, N3355);
buf BUF1 (N3359, N3357);
buf BUF1 (N3360, N3350);
nand NAND2 (N3361, N3346, N1298);
nand NAND4 (N3362, N3360, N994, N1244, N2105);
or OR2 (N3363, N3356, N1104);
nor NOR2 (N3364, N3349, N3226);
xor XOR2 (N3365, N3361, N95);
nor NOR2 (N3366, N3365, N448);
nand NAND3 (N3367, N3338, N926, N620);
and AND3 (N3368, N3367, N2307, N2848);
or OR4 (N3369, N3363, N808, N361, N196);
nor NOR3 (N3370, N3364, N453, N2534);
nand NAND4 (N3371, N3354, N3334, N3009, N1875);
nor NOR2 (N3372, N3362, N2434);
or OR3 (N3373, N3372, N3127, N3025);
or OR3 (N3374, N3366, N2682, N1905);
or OR4 (N3375, N3370, N2709, N595, N2086);
not NOT1 (N3376, N3373);
xor XOR2 (N3377, N3376, N2292);
xor XOR2 (N3378, N3374, N2435);
nand NAND2 (N3379, N3348, N1554);
or OR2 (N3380, N3345, N2980);
and AND3 (N3381, N3377, N2816, N3039);
buf BUF1 (N3382, N3378);
nand NAND4 (N3383, N3359, N343, N452, N1445);
buf BUF1 (N3384, N3371);
not NOT1 (N3385, N3381);
nand NAND3 (N3386, N3368, N599, N2248);
xor XOR2 (N3387, N3383, N3361);
nand NAND4 (N3388, N3380, N962, N2127, N1564);
nor NOR2 (N3389, N3388, N2047);
buf BUF1 (N3390, N3389);
or OR2 (N3391, N3387, N2195);
not NOT1 (N3392, N3391);
nand NAND2 (N3393, N3392, N2860);
nor NOR2 (N3394, N3384, N937);
and AND3 (N3395, N3382, N869, N2677);
buf BUF1 (N3396, N3395);
and AND4 (N3397, N3396, N536, N2748, N3082);
buf BUF1 (N3398, N3394);
and AND4 (N3399, N3375, N3275, N2942, N1704);
nand NAND3 (N3400, N3399, N2770, N1640);
nor NOR2 (N3401, N3385, N2138);
and AND4 (N3402, N3401, N3219, N662, N885);
nor NOR3 (N3403, N3369, N246, N2650);
or OR3 (N3404, N3398, N1579, N2538);
xor XOR2 (N3405, N3379, N946);
or OR2 (N3406, N3404, N2395);
nand NAND3 (N3407, N3358, N2612, N818);
nor NOR2 (N3408, N3397, N1283);
or OR3 (N3409, N3403, N313, N3301);
nand NAND3 (N3410, N3390, N1485, N337);
or OR4 (N3411, N3408, N1433, N1902, N1569);
not NOT1 (N3412, N3410);
xor XOR2 (N3413, N3407, N3411);
nand NAND2 (N3414, N3268, N2359);
or OR2 (N3415, N3413, N468);
and AND4 (N3416, N3412, N932, N1044, N476);
and AND4 (N3417, N3393, N2436, N635, N1244);
nor NOR2 (N3418, N3400, N1832);
nor NOR4 (N3419, N3414, N1151, N1504, N63);
nor NOR2 (N3420, N3418, N673);
not NOT1 (N3421, N3409);
buf BUF1 (N3422, N3415);
or OR2 (N3423, N3420, N330);
and AND3 (N3424, N3405, N1404, N2306);
buf BUF1 (N3425, N3424);
xor XOR2 (N3426, N3423, N2674);
and AND4 (N3427, N3406, N77, N3348, N2113);
nor NOR4 (N3428, N3402, N9, N2069, N2826);
nor NOR2 (N3429, N3419, N696);
or OR3 (N3430, N3428, N1107, N2935);
buf BUF1 (N3431, N3429);
nor NOR2 (N3432, N3416, N1215);
and AND2 (N3433, N3432, N1470);
xor XOR2 (N3434, N3427, N2401);
nor NOR3 (N3435, N3434, N1028, N947);
buf BUF1 (N3436, N3425);
buf BUF1 (N3437, N3431);
nand NAND2 (N3438, N3422, N2748);
xor XOR2 (N3439, N3430, N131);
nor NOR4 (N3440, N3386, N597, N3380, N2308);
and AND2 (N3441, N3439, N1163);
and AND3 (N3442, N3438, N1122, N1660);
and AND2 (N3443, N3421, N1729);
nor NOR4 (N3444, N3435, N3189, N785, N443);
xor XOR2 (N3445, N3433, N667);
buf BUF1 (N3446, N3417);
and AND4 (N3447, N3437, N2303, N2176, N3154);
nor NOR2 (N3448, N3447, N1433);
xor XOR2 (N3449, N3436, N1779);
buf BUF1 (N3450, N3442);
nor NOR2 (N3451, N3444, N1509);
nand NAND2 (N3452, N3443, N3379);
nand NAND3 (N3453, N3441, N290, N3031);
nor NOR4 (N3454, N3445, N859, N3121, N774);
or OR2 (N3455, N3451, N1217);
not NOT1 (N3456, N3455);
nand NAND3 (N3457, N3440, N1940, N264);
and AND3 (N3458, N3449, N2133, N1833);
buf BUF1 (N3459, N3426);
buf BUF1 (N3460, N3459);
nor NOR4 (N3461, N3458, N3027, N2030, N1237);
not NOT1 (N3462, N3453);
buf BUF1 (N3463, N3457);
or OR4 (N3464, N3462, N1633, N880, N2221);
xor XOR2 (N3465, N3464, N2005);
and AND3 (N3466, N3460, N685, N3125);
nor NOR3 (N3467, N3466, N2184, N890);
xor XOR2 (N3468, N3461, N1099);
nand NAND3 (N3469, N3454, N641, N2725);
xor XOR2 (N3470, N3468, N1352);
not NOT1 (N3471, N3448);
xor XOR2 (N3472, N3469, N1182);
nor NOR3 (N3473, N3467, N316, N2835);
xor XOR2 (N3474, N3446, N2886);
xor XOR2 (N3475, N3463, N2581);
and AND3 (N3476, N3450, N3088, N269);
nor NOR3 (N3477, N3474, N2762, N3200);
nor NOR2 (N3478, N3456, N2884);
and AND3 (N3479, N3475, N3232, N2375);
nor NOR3 (N3480, N3472, N2001, N1340);
or OR4 (N3481, N3473, N792, N1375, N1621);
nand NAND4 (N3482, N3470, N3422, N1008, N83);
buf BUF1 (N3483, N3481);
or OR4 (N3484, N3478, N2620, N894, N3448);
not NOT1 (N3485, N3480);
or OR2 (N3486, N3476, N2837);
buf BUF1 (N3487, N3483);
nand NAND4 (N3488, N3487, N4, N719, N2122);
nand NAND3 (N3489, N3488, N2938, N1224);
or OR4 (N3490, N3471, N908, N133, N330);
or OR3 (N3491, N3482, N1202, N2250);
and AND3 (N3492, N3477, N1019, N1714);
buf BUF1 (N3493, N3452);
nor NOR4 (N3494, N3493, N2141, N429, N834);
xor XOR2 (N3495, N3494, N584);
and AND2 (N3496, N3479, N1752);
nand NAND3 (N3497, N3491, N614, N1579);
or OR2 (N3498, N3496, N1592);
buf BUF1 (N3499, N3490);
buf BUF1 (N3500, N3485);
xor XOR2 (N3501, N3465, N627);
not NOT1 (N3502, N3497);
buf BUF1 (N3503, N3495);
nor NOR4 (N3504, N3501, N3285, N3387, N3437);
nor NOR4 (N3505, N3492, N1098, N3159, N272);
nand NAND3 (N3506, N3502, N3323, N2101);
and AND2 (N3507, N3506, N534);
buf BUF1 (N3508, N3504);
nor NOR3 (N3509, N3489, N2397, N719);
not NOT1 (N3510, N3507);
xor XOR2 (N3511, N3510, N1808);
buf BUF1 (N3512, N3484);
not NOT1 (N3513, N3512);
buf BUF1 (N3514, N3513);
not NOT1 (N3515, N3514);
and AND3 (N3516, N3486, N3140, N1145);
not NOT1 (N3517, N3498);
nor NOR4 (N3518, N3500, N1488, N1381, N2995);
nor NOR4 (N3519, N3508, N1255, N115, N3492);
xor XOR2 (N3520, N3515, N1305);
buf BUF1 (N3521, N3509);
buf BUF1 (N3522, N3520);
or OR2 (N3523, N3503, N1142);
endmodule