// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22;

output N16016,N15989,N15994,N16021,N16020,N16011,N16019,N16017,N16012,N16022;

nor NOR4 (N23, N15, N4, N20, N3);
buf BUF1 (N24, N13);
or OR3 (N25, N17, N11, N4);
buf BUF1 (N26, N10);
xor XOR2 (N27, N12, N4);
or OR2 (N28, N4, N22);
nand NAND4 (N29, N13, N10, N3, N15);
buf BUF1 (N30, N8);
nand NAND2 (N31, N3, N20);
nand NAND2 (N32, N31, N16);
nor NOR4 (N33, N16, N30, N6, N30);
buf BUF1 (N34, N4);
and AND2 (N35, N25, N13);
nand NAND4 (N36, N26, N32, N9, N27);
not NOT1 (N37, N33);
and AND4 (N38, N19, N1, N33, N4);
not NOT1 (N39, N15);
and AND3 (N40, N28, N3, N9);
buf BUF1 (N41, N37);
buf BUF1 (N42, N35);
xor XOR2 (N43, N39, N28);
nand NAND2 (N44, N34, N33);
xor XOR2 (N45, N40, N30);
or OR4 (N46, N24, N41, N4, N34);
and AND2 (N47, N44, N42);
buf BUF1 (N48, N3);
and AND2 (N49, N37, N40);
or OR3 (N50, N23, N32, N48);
nor NOR2 (N51, N32, N48);
nor NOR3 (N52, N47, N10, N26);
buf BUF1 (N53, N36);
buf BUF1 (N54, N52);
or OR4 (N55, N53, N22, N10, N7);
xor XOR2 (N56, N49, N13);
xor XOR2 (N57, N38, N25);
buf BUF1 (N58, N43);
buf BUF1 (N59, N55);
buf BUF1 (N60, N54);
xor XOR2 (N61, N46, N3);
or OR4 (N62, N51, N5, N24, N42);
or OR3 (N63, N61, N28, N54);
nand NAND4 (N64, N59, N27, N63, N53);
xor XOR2 (N65, N14, N8);
buf BUF1 (N66, N65);
and AND3 (N67, N29, N32, N2);
nor NOR4 (N68, N62, N8, N66, N8);
buf BUF1 (N69, N26);
not NOT1 (N70, N45);
buf BUF1 (N71, N69);
or OR3 (N72, N57, N33, N47);
nand NAND3 (N73, N56, N40, N17);
nand NAND4 (N74, N60, N16, N25, N12);
nor NOR2 (N75, N50, N9);
and AND4 (N76, N72, N17, N45, N42);
buf BUF1 (N77, N75);
nor NOR3 (N78, N74, N27, N70);
nand NAND3 (N79, N7, N41, N20);
not NOT1 (N80, N64);
not NOT1 (N81, N73);
buf BUF1 (N82, N67);
not NOT1 (N83, N58);
and AND4 (N84, N79, N1, N49, N6);
buf BUF1 (N85, N78);
nand NAND2 (N86, N82, N59);
buf BUF1 (N87, N81);
buf BUF1 (N88, N76);
not NOT1 (N89, N88);
or OR4 (N90, N86, N62, N87, N29);
and AND2 (N91, N72, N70);
nand NAND4 (N92, N80, N89, N45, N86);
xor XOR2 (N93, N76, N24);
and AND2 (N94, N77, N61);
and AND2 (N95, N94, N57);
xor XOR2 (N96, N92, N1);
and AND4 (N97, N95, N72, N96, N13);
or OR4 (N98, N86, N9, N6, N21);
nand NAND3 (N99, N84, N85, N37);
or OR2 (N100, N20, N31);
and AND3 (N101, N93, N10, N32);
or OR2 (N102, N71, N3);
xor XOR2 (N103, N83, N7);
xor XOR2 (N104, N100, N89);
nand NAND4 (N105, N102, N6, N86, N2);
nor NOR4 (N106, N101, N45, N3, N64);
or OR2 (N107, N97, N34);
or OR2 (N108, N99, N53);
and AND3 (N109, N105, N71, N84);
not NOT1 (N110, N107);
and AND3 (N111, N109, N71, N109);
xor XOR2 (N112, N110, N66);
nor NOR4 (N113, N98, N71, N101, N4);
nand NAND2 (N114, N68, N70);
buf BUF1 (N115, N113);
nor NOR2 (N116, N115, N10);
or OR4 (N117, N106, N113, N21, N52);
or OR3 (N118, N114, N12, N66);
or OR2 (N119, N116, N30);
nand NAND2 (N120, N117, N21);
nand NAND3 (N121, N120, N97, N3);
buf BUF1 (N122, N119);
xor XOR2 (N123, N103, N93);
not NOT1 (N124, N104);
xor XOR2 (N125, N91, N72);
and AND3 (N126, N111, N62, N40);
and AND2 (N127, N122, N20);
and AND4 (N128, N127, N100, N53, N18);
nand NAND2 (N129, N108, N38);
buf BUF1 (N130, N128);
nand NAND4 (N131, N129, N19, N127, N71);
nor NOR4 (N132, N112, N31, N79, N46);
nor NOR3 (N133, N118, N25, N95);
nor NOR3 (N134, N125, N115, N9);
not NOT1 (N135, N121);
buf BUF1 (N136, N124);
nand NAND2 (N137, N136, N88);
nor NOR3 (N138, N134, N20, N39);
nand NAND4 (N139, N135, N71, N116, N27);
nor NOR3 (N140, N126, N102, N133);
xor XOR2 (N141, N16, N121);
or OR3 (N142, N132, N39, N39);
not NOT1 (N143, N130);
not NOT1 (N144, N139);
nor NOR2 (N145, N141, N91);
buf BUF1 (N146, N137);
and AND2 (N147, N146, N130);
and AND3 (N148, N147, N146, N64);
nor NOR3 (N149, N123, N1, N125);
xor XOR2 (N150, N90, N23);
buf BUF1 (N151, N144);
not NOT1 (N152, N149);
xor XOR2 (N153, N138, N80);
buf BUF1 (N154, N142);
xor XOR2 (N155, N140, N19);
nor NOR4 (N156, N152, N120, N68, N6);
xor XOR2 (N157, N131, N46);
nand NAND2 (N158, N148, N17);
and AND3 (N159, N153, N118, N85);
nand NAND4 (N160, N151, N13, N31, N15);
and AND2 (N161, N150, N71);
nor NOR3 (N162, N160, N54, N104);
or OR3 (N163, N159, N149, N101);
and AND4 (N164, N143, N105, N129, N120);
and AND3 (N165, N158, N3, N36);
xor XOR2 (N166, N164, N29);
buf BUF1 (N167, N154);
or OR4 (N168, N156, N68, N67, N66);
nand NAND3 (N169, N165, N6, N67);
nor NOR4 (N170, N167, N96, N78, N159);
and AND2 (N171, N163, N106);
buf BUF1 (N172, N169);
nor NOR2 (N173, N171, N72);
and AND4 (N174, N161, N77, N46, N16);
or OR2 (N175, N155, N81);
or OR2 (N176, N170, N154);
buf BUF1 (N177, N172);
xor XOR2 (N178, N162, N134);
and AND4 (N179, N157, N23, N66, N140);
xor XOR2 (N180, N175, N98);
and AND2 (N181, N166, N136);
or OR2 (N182, N178, N21);
buf BUF1 (N183, N181);
nand NAND3 (N184, N145, N114, N1);
buf BUF1 (N185, N173);
buf BUF1 (N186, N184);
xor XOR2 (N187, N180, N168);
nand NAND4 (N188, N122, N174, N8, N97);
not NOT1 (N189, N160);
nand NAND4 (N190, N186, N143, N101, N37);
buf BUF1 (N191, N189);
buf BUF1 (N192, N183);
and AND4 (N193, N182, N66, N5, N188);
xor XOR2 (N194, N10, N132);
and AND2 (N195, N187, N170);
xor XOR2 (N196, N179, N35);
not NOT1 (N197, N177);
and AND2 (N198, N194, N75);
or OR4 (N199, N198, N129, N141, N19);
nor NOR2 (N200, N176, N116);
xor XOR2 (N201, N199, N60);
or OR2 (N202, N197, N198);
nand NAND4 (N203, N202, N192, N52, N143);
nand NAND2 (N204, N203, N125);
nand NAND2 (N205, N15, N171);
nand NAND3 (N206, N193, N125, N161);
nand NAND3 (N207, N205, N169, N89);
xor XOR2 (N208, N201, N104);
not NOT1 (N209, N204);
not NOT1 (N210, N207);
xor XOR2 (N211, N190, N3);
not NOT1 (N212, N195);
not NOT1 (N213, N196);
buf BUF1 (N214, N208);
nand NAND4 (N215, N206, N53, N196, N102);
not NOT1 (N216, N191);
nand NAND4 (N217, N200, N40, N129, N36);
buf BUF1 (N218, N185);
or OR2 (N219, N211, N134);
not NOT1 (N220, N216);
buf BUF1 (N221, N220);
and AND2 (N222, N219, N3);
nand NAND4 (N223, N217, N98, N156, N124);
not NOT1 (N224, N209);
nor NOR3 (N225, N222, N52, N114);
nand NAND4 (N226, N221, N154, N41, N14);
not NOT1 (N227, N223);
or OR4 (N228, N224, N17, N80, N146);
or OR4 (N229, N215, N158, N221, N92);
or OR3 (N230, N228, N166, N111);
nand NAND3 (N231, N212, N127, N27);
not NOT1 (N232, N226);
and AND3 (N233, N214, N156, N87);
xor XOR2 (N234, N233, N209);
and AND4 (N235, N213, N21, N14, N207);
and AND2 (N236, N234, N33);
xor XOR2 (N237, N236, N54);
nor NOR2 (N238, N231, N183);
xor XOR2 (N239, N235, N117);
nand NAND4 (N240, N237, N238, N187, N180);
and AND2 (N241, N134, N14);
not NOT1 (N242, N232);
nor NOR2 (N243, N229, N185);
and AND3 (N244, N225, N36, N132);
not NOT1 (N245, N242);
buf BUF1 (N246, N243);
nand NAND3 (N247, N240, N68, N155);
buf BUF1 (N248, N241);
nor NOR4 (N249, N247, N134, N35, N57);
xor XOR2 (N250, N218, N86);
or OR4 (N251, N248, N233, N70, N29);
nor NOR4 (N252, N239, N128, N24, N78);
or OR4 (N253, N246, N148, N129, N88);
or OR3 (N254, N227, N241, N178);
and AND3 (N255, N245, N99, N48);
nor NOR2 (N256, N250, N12);
nor NOR3 (N257, N210, N134, N222);
not NOT1 (N258, N249);
not NOT1 (N259, N256);
buf BUF1 (N260, N259);
and AND2 (N261, N253, N125);
buf BUF1 (N262, N258);
or OR3 (N263, N252, N250, N246);
xor XOR2 (N264, N255, N156);
xor XOR2 (N265, N263, N80);
and AND4 (N266, N262, N149, N263, N227);
buf BUF1 (N267, N254);
or OR4 (N268, N261, N165, N122, N36);
xor XOR2 (N269, N266, N233);
not NOT1 (N270, N257);
nand NAND4 (N271, N267, N142, N213, N131);
or OR2 (N272, N251, N111);
not NOT1 (N273, N271);
xor XOR2 (N274, N264, N260);
buf BUF1 (N275, N220);
nand NAND4 (N276, N265, N176, N174, N275);
buf BUF1 (N277, N264);
nor NOR3 (N278, N277, N22, N10);
not NOT1 (N279, N276);
xor XOR2 (N280, N268, N227);
and AND4 (N281, N244, N97, N277, N249);
and AND2 (N282, N269, N272);
not NOT1 (N283, N187);
nor NOR4 (N284, N274, N224, N138, N10);
xor XOR2 (N285, N230, N4);
nand NAND2 (N286, N281, N218);
or OR3 (N287, N286, N224, N109);
and AND4 (N288, N287, N280, N184, N32);
buf BUF1 (N289, N52);
and AND4 (N290, N288, N124, N65, N197);
and AND3 (N291, N278, N228, N2);
buf BUF1 (N292, N291);
and AND2 (N293, N279, N122);
nand NAND2 (N294, N285, N62);
buf BUF1 (N295, N270);
nor NOR4 (N296, N282, N23, N108, N179);
buf BUF1 (N297, N290);
nand NAND4 (N298, N289, N156, N82, N246);
not NOT1 (N299, N283);
not NOT1 (N300, N299);
nor NOR3 (N301, N300, N200, N93);
buf BUF1 (N302, N273);
buf BUF1 (N303, N296);
nor NOR2 (N304, N294, N213);
not NOT1 (N305, N284);
nand NAND4 (N306, N303, N51, N196, N219);
not NOT1 (N307, N293);
nor NOR2 (N308, N298, N35);
and AND3 (N309, N292, N33, N21);
or OR4 (N310, N302, N206, N131, N11);
xor XOR2 (N311, N306, N217);
xor XOR2 (N312, N297, N282);
not NOT1 (N313, N309);
or OR3 (N314, N307, N218, N65);
and AND4 (N315, N313, N171, N68, N248);
or OR3 (N316, N312, N167, N229);
or OR2 (N317, N315, N282);
buf BUF1 (N318, N311);
buf BUF1 (N319, N310);
or OR2 (N320, N301, N55);
and AND2 (N321, N308, N38);
xor XOR2 (N322, N305, N239);
and AND2 (N323, N322, N172);
xor XOR2 (N324, N304, N161);
nand NAND2 (N325, N316, N185);
or OR4 (N326, N321, N185, N69, N247);
nand NAND3 (N327, N323, N97, N232);
nor NOR2 (N328, N324, N149);
buf BUF1 (N329, N327);
nand NAND4 (N330, N320, N12, N226, N203);
buf BUF1 (N331, N317);
not NOT1 (N332, N331);
buf BUF1 (N333, N329);
and AND4 (N334, N325, N77, N47, N100);
nand NAND2 (N335, N332, N221);
xor XOR2 (N336, N328, N238);
and AND4 (N337, N326, N235, N42, N257);
nor NOR4 (N338, N330, N27, N22, N101);
and AND3 (N339, N319, N204, N21);
nand NAND3 (N340, N337, N148, N196);
nor NOR3 (N341, N295, N82, N104);
nor NOR2 (N342, N340, N216);
not NOT1 (N343, N318);
buf BUF1 (N344, N335);
xor XOR2 (N345, N342, N212);
nand NAND4 (N346, N338, N29, N166, N5);
nand NAND3 (N347, N344, N119, N335);
or OR3 (N348, N343, N9, N70);
nand NAND2 (N349, N341, N322);
and AND4 (N350, N314, N83, N72, N167);
not NOT1 (N351, N345);
xor XOR2 (N352, N350, N296);
and AND3 (N353, N347, N116, N22);
xor XOR2 (N354, N334, N61);
nor NOR4 (N355, N346, N294, N195, N192);
and AND3 (N356, N353, N63, N171);
xor XOR2 (N357, N354, N56);
xor XOR2 (N358, N357, N147);
nand NAND4 (N359, N349, N156, N44, N143);
nand NAND2 (N360, N351, N161);
nor NOR2 (N361, N359, N348);
and AND3 (N362, N62, N148, N74);
and AND2 (N363, N358, N167);
and AND4 (N364, N356, N220, N323, N312);
buf BUF1 (N365, N364);
not NOT1 (N366, N362);
buf BUF1 (N367, N336);
nand NAND2 (N368, N360, N70);
not NOT1 (N369, N355);
nand NAND4 (N370, N339, N86, N206, N217);
or OR4 (N371, N352, N214, N205, N176);
or OR3 (N372, N363, N161, N306);
and AND3 (N373, N367, N39, N247);
or OR3 (N374, N366, N50, N71);
not NOT1 (N375, N369);
buf BUF1 (N376, N365);
and AND4 (N377, N370, N15, N59, N279);
not NOT1 (N378, N373);
or OR2 (N379, N371, N195);
xor XOR2 (N380, N378, N244);
nor NOR3 (N381, N380, N187, N206);
nand NAND3 (N382, N372, N213, N187);
and AND3 (N383, N377, N230, N217);
nand NAND2 (N384, N379, N115);
nand NAND2 (N385, N383, N85);
or OR4 (N386, N376, N206, N299, N44);
not NOT1 (N387, N381);
and AND4 (N388, N382, N12, N364, N276);
or OR2 (N389, N384, N73);
nor NOR2 (N390, N333, N98);
xor XOR2 (N391, N361, N104);
buf BUF1 (N392, N375);
not NOT1 (N393, N374);
not NOT1 (N394, N393);
not NOT1 (N395, N390);
and AND3 (N396, N392, N390, N229);
buf BUF1 (N397, N389);
buf BUF1 (N398, N394);
or OR3 (N399, N368, N396, N295);
nand NAND4 (N400, N304, N346, N276, N310);
or OR3 (N401, N388, N127, N338);
or OR3 (N402, N385, N156, N81);
nand NAND3 (N403, N387, N264, N161);
nand NAND3 (N404, N400, N350, N359);
not NOT1 (N405, N386);
nand NAND4 (N406, N401, N211, N39, N110);
and AND3 (N407, N404, N164, N393);
not NOT1 (N408, N395);
nor NOR4 (N409, N399, N322, N381, N45);
xor XOR2 (N410, N408, N190);
and AND3 (N411, N407, N382, N269);
buf BUF1 (N412, N410);
xor XOR2 (N413, N409, N297);
and AND3 (N414, N397, N119, N32);
nand NAND4 (N415, N413, N80, N384, N155);
nand NAND2 (N416, N391, N188);
buf BUF1 (N417, N406);
nand NAND4 (N418, N417, N303, N401, N199);
not NOT1 (N419, N414);
not NOT1 (N420, N405);
not NOT1 (N421, N411);
nor NOR2 (N422, N419, N370);
or OR4 (N423, N420, N18, N339, N123);
nor NOR4 (N424, N402, N315, N136, N196);
not NOT1 (N425, N403);
or OR4 (N426, N422, N160, N143, N244);
nand NAND4 (N427, N423, N272, N294, N369);
xor XOR2 (N428, N415, N397);
nand NAND4 (N429, N427, N86, N9, N377);
or OR2 (N430, N426, N153);
not NOT1 (N431, N425);
or OR3 (N432, N421, N341, N12);
not NOT1 (N433, N432);
or OR4 (N434, N431, N433, N399, N117);
nor NOR3 (N435, N268, N6, N88);
xor XOR2 (N436, N398, N56);
xor XOR2 (N437, N412, N214);
and AND3 (N438, N428, N243, N222);
buf BUF1 (N439, N429);
not NOT1 (N440, N430);
buf BUF1 (N441, N435);
buf BUF1 (N442, N418);
nand NAND3 (N443, N436, N87, N291);
xor XOR2 (N444, N443, N108);
or OR4 (N445, N442, N434, N204, N23);
or OR3 (N446, N299, N391, N239);
nand NAND2 (N447, N446, N409);
buf BUF1 (N448, N445);
and AND2 (N449, N440, N370);
buf BUF1 (N450, N416);
xor XOR2 (N451, N444, N204);
nand NAND4 (N452, N448, N60, N380, N73);
and AND3 (N453, N451, N402, N147);
not NOT1 (N454, N441);
not NOT1 (N455, N447);
and AND2 (N456, N454, N9);
xor XOR2 (N457, N437, N439);
nor NOR4 (N458, N20, N145, N38, N38);
not NOT1 (N459, N457);
nor NOR3 (N460, N453, N305, N436);
nand NAND4 (N461, N456, N182, N412, N241);
nand NAND4 (N462, N450, N394, N58, N224);
and AND4 (N463, N449, N288, N202, N350);
nand NAND3 (N464, N462, N412, N412);
or OR2 (N465, N460, N462);
or OR3 (N466, N464, N153, N461);
or OR2 (N467, N216, N161);
not NOT1 (N468, N458);
and AND2 (N469, N424, N468);
buf BUF1 (N470, N37);
not NOT1 (N471, N470);
and AND3 (N472, N466, N196, N131);
nor NOR3 (N473, N452, N310, N54);
or OR4 (N474, N467, N470, N344, N283);
nor NOR3 (N475, N459, N422, N124);
and AND2 (N476, N455, N188);
and AND3 (N477, N472, N220, N9);
nand NAND2 (N478, N465, N401);
buf BUF1 (N479, N473);
nand NAND3 (N480, N475, N443, N52);
nand NAND3 (N481, N477, N52, N351);
and AND3 (N482, N474, N150, N324);
xor XOR2 (N483, N482, N48);
not NOT1 (N484, N471);
not NOT1 (N485, N483);
buf BUF1 (N486, N476);
buf BUF1 (N487, N486);
xor XOR2 (N488, N478, N303);
nand NAND2 (N489, N481, N454);
or OR3 (N490, N438, N405, N23);
and AND3 (N491, N490, N69, N300);
and AND2 (N492, N488, N405);
and AND3 (N493, N463, N95, N94);
or OR2 (N494, N485, N167);
buf BUF1 (N495, N494);
not NOT1 (N496, N480);
nor NOR2 (N497, N495, N374);
nor NOR3 (N498, N479, N54, N40);
xor XOR2 (N499, N492, N260);
not NOT1 (N500, N469);
nor NOR3 (N501, N493, N96, N494);
buf BUF1 (N502, N487);
not NOT1 (N503, N491);
not NOT1 (N504, N498);
or OR3 (N505, N500, N114, N286);
and AND3 (N506, N505, N345, N22);
or OR4 (N507, N502, N373, N83, N352);
and AND3 (N508, N484, N460, N80);
not NOT1 (N509, N496);
not NOT1 (N510, N489);
nor NOR2 (N511, N504, N504);
buf BUF1 (N512, N510);
or OR4 (N513, N506, N410, N475, N326);
buf BUF1 (N514, N503);
nand NAND4 (N515, N497, N304, N162, N286);
xor XOR2 (N516, N507, N369);
nor NOR3 (N517, N508, N421, N406);
and AND4 (N518, N512, N244, N175, N421);
buf BUF1 (N519, N511);
nand NAND2 (N520, N517, N99);
nor NOR2 (N521, N520, N121);
not NOT1 (N522, N518);
not NOT1 (N523, N515);
xor XOR2 (N524, N513, N146);
and AND4 (N525, N516, N471, N508, N143);
or OR2 (N526, N519, N437);
nand NAND2 (N527, N522, N267);
xor XOR2 (N528, N527, N266);
or OR3 (N529, N499, N169, N30);
or OR2 (N530, N514, N465);
nor NOR2 (N531, N525, N256);
or OR2 (N532, N523, N371);
buf BUF1 (N533, N530);
and AND4 (N534, N526, N173, N532, N67);
or OR3 (N535, N259, N433, N184);
not NOT1 (N536, N509);
xor XOR2 (N537, N501, N387);
not NOT1 (N538, N534);
nand NAND2 (N539, N521, N322);
buf BUF1 (N540, N537);
nand NAND4 (N541, N536, N393, N247, N174);
and AND3 (N542, N531, N397, N170);
nand NAND3 (N543, N542, N30, N154);
and AND2 (N544, N541, N35);
or OR3 (N545, N540, N26, N331);
nor NOR2 (N546, N544, N537);
nand NAND2 (N547, N528, N246);
xor XOR2 (N548, N546, N6);
nor NOR2 (N549, N533, N144);
or OR2 (N550, N545, N360);
or OR4 (N551, N538, N228, N211, N488);
buf BUF1 (N552, N547);
not NOT1 (N553, N539);
or OR3 (N554, N529, N412, N220);
not NOT1 (N555, N535);
or OR3 (N556, N548, N109, N157);
xor XOR2 (N557, N524, N191);
and AND4 (N558, N552, N300, N123, N261);
xor XOR2 (N559, N557, N330);
or OR4 (N560, N555, N89, N226, N393);
or OR3 (N561, N549, N228, N490);
nand NAND4 (N562, N556, N359, N210, N147);
buf BUF1 (N563, N553);
nand NAND4 (N564, N560, N418, N189, N90);
nand NAND4 (N565, N559, N7, N85, N384);
or OR4 (N566, N565, N327, N16, N355);
buf BUF1 (N567, N564);
not NOT1 (N568, N554);
nand NAND4 (N569, N563, N74, N292, N93);
buf BUF1 (N570, N562);
xor XOR2 (N571, N543, N235);
nand NAND2 (N572, N570, N359);
or OR2 (N573, N558, N11);
and AND4 (N574, N569, N141, N76, N243);
xor XOR2 (N575, N561, N214);
xor XOR2 (N576, N571, N549);
or OR3 (N577, N567, N159, N461);
nand NAND3 (N578, N573, N510, N154);
or OR3 (N579, N568, N497, N177);
nand NAND2 (N580, N578, N15);
and AND3 (N581, N566, N490, N510);
and AND4 (N582, N550, N556, N434, N93);
xor XOR2 (N583, N576, N470);
not NOT1 (N584, N575);
nor NOR4 (N585, N551, N524, N341, N579);
nor NOR4 (N586, N383, N117, N491, N336);
nor NOR2 (N587, N574, N132);
and AND3 (N588, N582, N247, N258);
or OR3 (N589, N580, N536, N368);
nor NOR4 (N590, N589, N561, N28, N104);
nand NAND2 (N591, N572, N172);
buf BUF1 (N592, N586);
and AND2 (N593, N591, N478);
nor NOR2 (N594, N581, N154);
and AND3 (N595, N583, N440, N98);
not NOT1 (N596, N587);
not NOT1 (N597, N594);
not NOT1 (N598, N590);
not NOT1 (N599, N595);
not NOT1 (N600, N593);
buf BUF1 (N601, N599);
nand NAND4 (N602, N585, N448, N49, N33);
or OR4 (N603, N588, N11, N499, N220);
not NOT1 (N604, N577);
nand NAND3 (N605, N601, N156, N50);
or OR3 (N606, N605, N236, N535);
xor XOR2 (N607, N596, N414);
and AND3 (N608, N603, N519, N422);
or OR2 (N609, N606, N169);
nand NAND4 (N610, N592, N444, N238, N36);
not NOT1 (N611, N598);
buf BUF1 (N612, N604);
xor XOR2 (N613, N607, N146);
and AND3 (N614, N608, N265, N367);
buf BUF1 (N615, N600);
not NOT1 (N616, N614);
nor NOR4 (N617, N615, N152, N49, N64);
xor XOR2 (N618, N584, N443);
or OR3 (N619, N611, N67, N527);
buf BUF1 (N620, N610);
or OR4 (N621, N616, N127, N464, N528);
nor NOR3 (N622, N597, N239, N568);
or OR2 (N623, N618, N531);
nand NAND4 (N624, N621, N384, N372, N30);
nor NOR4 (N625, N622, N305, N273, N591);
buf BUF1 (N626, N625);
nor NOR4 (N627, N609, N83, N569, N608);
buf BUF1 (N628, N612);
not NOT1 (N629, N626);
and AND3 (N630, N619, N153, N565);
nand NAND4 (N631, N620, N160, N441, N433);
nand NAND2 (N632, N630, N534);
nand NAND4 (N633, N602, N379, N497, N422);
buf BUF1 (N634, N628);
and AND4 (N635, N634, N389, N320, N9);
xor XOR2 (N636, N635, N49);
nor NOR4 (N637, N623, N81, N489, N300);
not NOT1 (N638, N617);
and AND4 (N639, N638, N401, N627, N527);
or OR2 (N640, N618, N522);
not NOT1 (N641, N629);
not NOT1 (N642, N631);
nand NAND4 (N643, N613, N253, N360, N415);
buf BUF1 (N644, N633);
xor XOR2 (N645, N644, N148);
not NOT1 (N646, N636);
not NOT1 (N647, N624);
xor XOR2 (N648, N639, N595);
nand NAND4 (N649, N632, N170, N229, N478);
buf BUF1 (N650, N637);
nor NOR2 (N651, N648, N393);
xor XOR2 (N652, N650, N133);
not NOT1 (N653, N643);
not NOT1 (N654, N646);
buf BUF1 (N655, N653);
nor NOR3 (N656, N645, N451, N264);
xor XOR2 (N657, N647, N474);
nand NAND4 (N658, N640, N10, N622, N511);
or OR3 (N659, N651, N593, N207);
not NOT1 (N660, N659);
nand NAND4 (N661, N652, N430, N121, N542);
and AND3 (N662, N641, N225, N187);
or OR2 (N663, N662, N648);
buf BUF1 (N664, N656);
not NOT1 (N665, N654);
and AND2 (N666, N657, N639);
or OR4 (N667, N661, N337, N366, N75);
not NOT1 (N668, N649);
nor NOR3 (N669, N668, N392, N545);
buf BUF1 (N670, N667);
nor NOR2 (N671, N665, N281);
nand NAND2 (N672, N670, N291);
and AND4 (N673, N663, N354, N466, N54);
nand NAND2 (N674, N660, N320);
nand NAND3 (N675, N672, N518, N78);
buf BUF1 (N676, N658);
xor XOR2 (N677, N675, N296);
or OR2 (N678, N677, N637);
nand NAND3 (N679, N673, N172, N665);
nor NOR3 (N680, N676, N252, N241);
buf BUF1 (N681, N642);
and AND2 (N682, N680, N525);
not NOT1 (N683, N682);
or OR3 (N684, N674, N82, N465);
xor XOR2 (N685, N679, N389);
and AND4 (N686, N683, N612, N362, N180);
or OR4 (N687, N684, N498, N17, N547);
xor XOR2 (N688, N671, N521);
and AND4 (N689, N686, N559, N269, N422);
buf BUF1 (N690, N688);
not NOT1 (N691, N664);
and AND4 (N692, N669, N375, N574, N380);
nor NOR3 (N693, N687, N27, N167);
xor XOR2 (N694, N678, N309);
and AND2 (N695, N694, N241);
nand NAND3 (N696, N690, N538, N492);
or OR3 (N697, N692, N537, N244);
not NOT1 (N698, N691);
nor NOR4 (N699, N681, N3, N658, N374);
nor NOR4 (N700, N689, N652, N461, N90);
xor XOR2 (N701, N655, N9);
or OR3 (N702, N700, N680, N536);
and AND4 (N703, N685, N542, N27, N195);
xor XOR2 (N704, N699, N444);
buf BUF1 (N705, N696);
buf BUF1 (N706, N703);
and AND4 (N707, N695, N90, N525, N677);
not NOT1 (N708, N698);
xor XOR2 (N709, N704, N332);
not NOT1 (N710, N707);
and AND2 (N711, N693, N577);
buf BUF1 (N712, N708);
nor NOR2 (N713, N710, N204);
and AND4 (N714, N705, N230, N293, N391);
xor XOR2 (N715, N713, N230);
not NOT1 (N716, N706);
or OR4 (N717, N697, N108, N127, N351);
buf BUF1 (N718, N716);
xor XOR2 (N719, N712, N594);
buf BUF1 (N720, N709);
and AND3 (N721, N714, N176, N701);
not NOT1 (N722, N516);
nand NAND4 (N723, N717, N717, N425, N296);
buf BUF1 (N724, N711);
nor NOR4 (N725, N715, N531, N586, N631);
xor XOR2 (N726, N722, N130);
or OR2 (N727, N726, N57);
and AND3 (N728, N725, N491, N14);
nand NAND2 (N729, N720, N84);
or OR3 (N730, N721, N407, N665);
or OR2 (N731, N724, N456);
not NOT1 (N732, N719);
nand NAND2 (N733, N723, N694);
nand NAND2 (N734, N731, N293);
and AND2 (N735, N728, N199);
or OR4 (N736, N718, N82, N23, N696);
or OR4 (N737, N735, N303, N385, N520);
nand NAND3 (N738, N734, N98, N195);
buf BUF1 (N739, N738);
nor NOR2 (N740, N732, N521);
not NOT1 (N741, N737);
not NOT1 (N742, N727);
and AND3 (N743, N739, N366, N146);
nand NAND2 (N744, N733, N604);
not NOT1 (N745, N702);
nor NOR2 (N746, N744, N403);
nand NAND3 (N747, N736, N650, N246);
xor XOR2 (N748, N741, N7);
or OR4 (N749, N747, N366, N520, N729);
buf BUF1 (N750, N711);
nand NAND4 (N751, N740, N548, N351, N701);
buf BUF1 (N752, N666);
and AND3 (N753, N748, N488, N361);
nand NAND2 (N754, N730, N598);
not NOT1 (N755, N745);
not NOT1 (N756, N742);
and AND3 (N757, N755, N315, N659);
or OR3 (N758, N746, N571, N236);
nor NOR3 (N759, N754, N132, N96);
buf BUF1 (N760, N753);
or OR2 (N761, N743, N683);
buf BUF1 (N762, N758);
not NOT1 (N763, N757);
xor XOR2 (N764, N759, N41);
buf BUF1 (N765, N763);
nor NOR2 (N766, N761, N36);
not NOT1 (N767, N766);
not NOT1 (N768, N764);
xor XOR2 (N769, N765, N523);
and AND3 (N770, N751, N659, N686);
nor NOR2 (N771, N760, N478);
buf BUF1 (N772, N767);
xor XOR2 (N773, N772, N527);
nor NOR2 (N774, N770, N481);
nand NAND4 (N775, N750, N471, N528, N243);
xor XOR2 (N776, N771, N222);
nand NAND4 (N777, N762, N27, N537, N62);
xor XOR2 (N778, N769, N391);
or OR3 (N779, N778, N599, N162);
not NOT1 (N780, N768);
nand NAND3 (N781, N777, N188, N323);
nor NOR2 (N782, N781, N609);
and AND3 (N783, N752, N3, N149);
or OR3 (N784, N780, N430, N430);
or OR3 (N785, N756, N478, N118);
nand NAND4 (N786, N776, N416, N65, N368);
nand NAND2 (N787, N786, N232);
nand NAND3 (N788, N783, N386, N159);
nand NAND2 (N789, N779, N334);
not NOT1 (N790, N785);
not NOT1 (N791, N782);
buf BUF1 (N792, N773);
buf BUF1 (N793, N774);
nor NOR3 (N794, N792, N108, N262);
and AND4 (N795, N793, N359, N697, N513);
xor XOR2 (N796, N794, N499);
or OR4 (N797, N749, N401, N283, N636);
nand NAND3 (N798, N797, N231, N526);
or OR2 (N799, N798, N762);
buf BUF1 (N800, N795);
xor XOR2 (N801, N775, N615);
nand NAND4 (N802, N790, N117, N757, N249);
nor NOR2 (N803, N799, N573);
or OR3 (N804, N788, N668, N687);
nand NAND4 (N805, N787, N266, N63, N505);
xor XOR2 (N806, N784, N79);
not NOT1 (N807, N805);
or OR4 (N808, N789, N736, N536, N374);
buf BUF1 (N809, N800);
or OR2 (N810, N808, N736);
buf BUF1 (N811, N791);
or OR3 (N812, N802, N621, N588);
buf BUF1 (N813, N801);
not NOT1 (N814, N812);
not NOT1 (N815, N804);
nor NOR3 (N816, N803, N91, N119);
buf BUF1 (N817, N815);
not NOT1 (N818, N806);
xor XOR2 (N819, N809, N484);
nor NOR3 (N820, N818, N326, N663);
not NOT1 (N821, N810);
nand NAND2 (N822, N819, N294);
xor XOR2 (N823, N816, N637);
nand NAND2 (N824, N811, N644);
nand NAND4 (N825, N814, N284, N146, N534);
not NOT1 (N826, N817);
xor XOR2 (N827, N807, N649);
nor NOR2 (N828, N827, N187);
or OR2 (N829, N822, N544);
nand NAND2 (N830, N821, N90);
nand NAND4 (N831, N829, N355, N511, N321);
nand NAND4 (N832, N830, N74, N125, N348);
buf BUF1 (N833, N826);
buf BUF1 (N834, N824);
nor NOR4 (N835, N828, N606, N55, N633);
nor NOR2 (N836, N833, N473);
nand NAND4 (N837, N820, N144, N350, N289);
or OR4 (N838, N836, N616, N710, N298);
nand NAND4 (N839, N838, N675, N363, N23);
or OR3 (N840, N834, N619, N659);
xor XOR2 (N841, N831, N687);
nand NAND2 (N842, N825, N279);
or OR3 (N843, N835, N154, N26);
buf BUF1 (N844, N823);
nand NAND3 (N845, N842, N83, N170);
nand NAND3 (N846, N813, N354, N787);
not NOT1 (N847, N796);
xor XOR2 (N848, N837, N800);
and AND4 (N849, N844, N13, N397, N336);
not NOT1 (N850, N840);
not NOT1 (N851, N850);
nor NOR4 (N852, N851, N265, N129, N720);
not NOT1 (N853, N839);
buf BUF1 (N854, N841);
or OR2 (N855, N852, N65);
buf BUF1 (N856, N853);
xor XOR2 (N857, N854, N393);
or OR2 (N858, N847, N608);
buf BUF1 (N859, N858);
or OR3 (N860, N832, N119, N644);
xor XOR2 (N861, N849, N221);
buf BUF1 (N862, N846);
not NOT1 (N863, N856);
or OR2 (N864, N860, N304);
and AND2 (N865, N863, N302);
buf BUF1 (N866, N859);
not NOT1 (N867, N855);
nor NOR4 (N868, N843, N410, N152, N397);
nand NAND2 (N869, N868, N119);
and AND4 (N870, N866, N147, N570, N741);
nand NAND2 (N871, N861, N89);
and AND3 (N872, N845, N130, N137);
and AND4 (N873, N848, N781, N277, N11);
buf BUF1 (N874, N862);
xor XOR2 (N875, N871, N117);
buf BUF1 (N876, N874);
xor XOR2 (N877, N870, N355);
or OR3 (N878, N877, N751, N648);
nor NOR4 (N879, N872, N293, N775, N775);
nand NAND2 (N880, N869, N662);
or OR2 (N881, N878, N421);
not NOT1 (N882, N881);
or OR4 (N883, N875, N569, N401, N447);
and AND2 (N884, N883, N494);
xor XOR2 (N885, N867, N44);
nand NAND3 (N886, N876, N196, N590);
nor NOR4 (N887, N882, N316, N618, N356);
or OR4 (N888, N873, N764, N186, N187);
nand NAND2 (N889, N888, N768);
and AND4 (N890, N857, N647, N342, N640);
and AND4 (N891, N890, N393, N227, N675);
or OR3 (N892, N865, N786, N692);
xor XOR2 (N893, N864, N702);
buf BUF1 (N894, N885);
nor NOR4 (N895, N892, N637, N548, N259);
nand NAND3 (N896, N879, N737, N176);
not NOT1 (N897, N894);
buf BUF1 (N898, N891);
and AND2 (N899, N897, N269);
not NOT1 (N900, N880);
xor XOR2 (N901, N887, N580);
nor NOR4 (N902, N900, N102, N601, N860);
not NOT1 (N903, N893);
and AND2 (N904, N902, N864);
not NOT1 (N905, N896);
not NOT1 (N906, N895);
and AND4 (N907, N905, N502, N248, N179);
buf BUF1 (N908, N889);
buf BUF1 (N909, N886);
or OR4 (N910, N908, N699, N731, N333);
buf BUF1 (N911, N903);
nand NAND3 (N912, N899, N596, N77);
and AND2 (N913, N906, N677);
or OR2 (N914, N912, N387);
not NOT1 (N915, N901);
not NOT1 (N916, N911);
nand NAND2 (N917, N916, N725);
xor XOR2 (N918, N914, N49);
nand NAND4 (N919, N918, N267, N768, N868);
or OR4 (N920, N904, N651, N667, N618);
nand NAND2 (N921, N920, N601);
or OR2 (N922, N915, N793);
xor XOR2 (N923, N909, N842);
buf BUF1 (N924, N898);
buf BUF1 (N925, N884);
nand NAND2 (N926, N922, N286);
buf BUF1 (N927, N924);
nor NOR4 (N928, N907, N332, N18, N97);
nand NAND2 (N929, N917, N691);
nor NOR2 (N930, N928, N534);
and AND3 (N931, N926, N440, N135);
not NOT1 (N932, N927);
nor NOR2 (N933, N923, N505);
and AND4 (N934, N933, N695, N467, N221);
or OR4 (N935, N910, N324, N327, N343);
nand NAND2 (N936, N930, N285);
not NOT1 (N937, N921);
and AND3 (N938, N919, N588, N484);
not NOT1 (N939, N929);
xor XOR2 (N940, N931, N115);
not NOT1 (N941, N934);
or OR4 (N942, N939, N694, N673, N360);
not NOT1 (N943, N935);
not NOT1 (N944, N936);
nor NOR3 (N945, N938, N422, N452);
or OR2 (N946, N937, N410);
or OR2 (N947, N944, N601);
or OR3 (N948, N940, N447, N561);
and AND2 (N949, N913, N565);
or OR3 (N950, N941, N14, N725);
buf BUF1 (N951, N943);
not NOT1 (N952, N951);
nor NOR4 (N953, N945, N814, N597, N39);
buf BUF1 (N954, N932);
buf BUF1 (N955, N952);
nand NAND2 (N956, N925, N371);
nand NAND4 (N957, N956, N45, N460, N652);
nor NOR4 (N958, N946, N56, N526, N745);
nor NOR3 (N959, N947, N78, N784);
nand NAND2 (N960, N949, N637);
not NOT1 (N961, N953);
or OR2 (N962, N955, N947);
nand NAND4 (N963, N950, N705, N713, N682);
nand NAND4 (N964, N963, N182, N913, N303);
buf BUF1 (N965, N961);
or OR3 (N966, N957, N793, N950);
nand NAND2 (N967, N958, N233);
not NOT1 (N968, N966);
and AND2 (N969, N965, N618);
and AND3 (N970, N959, N3, N524);
and AND3 (N971, N942, N426, N857);
or OR2 (N972, N964, N168);
or OR3 (N973, N971, N745, N177);
and AND4 (N974, N969, N873, N812, N50);
or OR3 (N975, N954, N592, N625);
xor XOR2 (N976, N970, N126);
xor XOR2 (N977, N973, N833);
or OR4 (N978, N975, N488, N459, N119);
or OR2 (N979, N972, N123);
and AND2 (N980, N962, N505);
not NOT1 (N981, N976);
not NOT1 (N982, N967);
not NOT1 (N983, N982);
not NOT1 (N984, N968);
buf BUF1 (N985, N948);
buf BUF1 (N986, N974);
buf BUF1 (N987, N985);
nand NAND3 (N988, N986, N275, N639);
and AND3 (N989, N979, N215, N447);
not NOT1 (N990, N977);
and AND2 (N991, N981, N587);
xor XOR2 (N992, N988, N361);
xor XOR2 (N993, N980, N738);
not NOT1 (N994, N993);
nor NOR4 (N995, N978, N605, N172, N992);
nand NAND4 (N996, N66, N664, N551, N911);
or OR2 (N997, N991, N730);
or OR4 (N998, N990, N468, N397, N877);
nand NAND4 (N999, N996, N76, N107, N108);
or OR2 (N1000, N994, N274);
xor XOR2 (N1001, N989, N92);
nand NAND2 (N1002, N1000, N117);
buf BUF1 (N1003, N984);
xor XOR2 (N1004, N999, N902);
nor NOR2 (N1005, N995, N314);
nand NAND2 (N1006, N960, N790);
and AND2 (N1007, N1002, N878);
nand NAND3 (N1008, N1001, N200, N487);
or OR4 (N1009, N997, N187, N602, N150);
and AND2 (N1010, N1003, N849);
xor XOR2 (N1011, N998, N425);
nand NAND3 (N1012, N983, N784, N89);
nand NAND2 (N1013, N1004, N572);
nand NAND4 (N1014, N1007, N1001, N75, N577);
not NOT1 (N1015, N1013);
not NOT1 (N1016, N1010);
or OR4 (N1017, N1012, N847, N137, N614);
xor XOR2 (N1018, N1005, N710);
nor NOR3 (N1019, N1009, N826, N281);
or OR3 (N1020, N1015, N305, N757);
and AND2 (N1021, N1014, N180);
and AND4 (N1022, N987, N49, N358, N484);
not NOT1 (N1023, N1017);
nor NOR3 (N1024, N1019, N849, N316);
or OR2 (N1025, N1023, N543);
not NOT1 (N1026, N1022);
buf BUF1 (N1027, N1025);
not NOT1 (N1028, N1021);
xor XOR2 (N1029, N1006, N1009);
or OR3 (N1030, N1027, N1017, N579);
xor XOR2 (N1031, N1028, N1016);
nor NOR3 (N1032, N743, N748, N750);
or OR3 (N1033, N1018, N896, N692);
or OR2 (N1034, N1026, N367);
nand NAND4 (N1035, N1031, N497, N564, N134);
and AND3 (N1036, N1008, N483, N276);
nor NOR4 (N1037, N1030, N742, N323, N255);
not NOT1 (N1038, N1020);
or OR4 (N1039, N1011, N312, N892, N82);
or OR4 (N1040, N1036, N473, N725, N301);
nor NOR3 (N1041, N1032, N422, N995);
buf BUF1 (N1042, N1040);
or OR4 (N1043, N1037, N142, N244, N86);
nor NOR4 (N1044, N1041, N504, N475, N491);
and AND4 (N1045, N1042, N500, N122, N40);
not NOT1 (N1046, N1029);
not NOT1 (N1047, N1038);
nor NOR2 (N1048, N1034, N828);
buf BUF1 (N1049, N1044);
nor NOR3 (N1050, N1024, N761, N175);
xor XOR2 (N1051, N1046, N778);
buf BUF1 (N1052, N1049);
or OR3 (N1053, N1050, N913, N546);
nor NOR2 (N1054, N1045, N26);
buf BUF1 (N1055, N1033);
and AND3 (N1056, N1035, N762, N267);
and AND4 (N1057, N1047, N558, N1043, N96);
nor NOR4 (N1058, N149, N1038, N838, N501);
or OR4 (N1059, N1057, N685, N147, N865);
nand NAND4 (N1060, N1059, N97, N595, N339);
not NOT1 (N1061, N1058);
not NOT1 (N1062, N1053);
nand NAND2 (N1063, N1055, N373);
buf BUF1 (N1064, N1060);
not NOT1 (N1065, N1062);
not NOT1 (N1066, N1052);
nor NOR2 (N1067, N1061, N110);
nand NAND3 (N1068, N1039, N194, N946);
xor XOR2 (N1069, N1065, N898);
nor NOR4 (N1070, N1066, N859, N1015, N447);
buf BUF1 (N1071, N1056);
and AND4 (N1072, N1067, N794, N586, N172);
buf BUF1 (N1073, N1070);
nand NAND4 (N1074, N1069, N686, N768, N322);
and AND2 (N1075, N1054, N400);
nand NAND4 (N1076, N1071, N252, N594, N270);
or OR4 (N1077, N1075, N283, N1050, N435);
nand NAND4 (N1078, N1077, N576, N276, N993);
buf BUF1 (N1079, N1076);
nand NAND4 (N1080, N1068, N880, N933, N47);
and AND4 (N1081, N1079, N378, N976, N156);
not NOT1 (N1082, N1080);
and AND2 (N1083, N1072, N741);
buf BUF1 (N1084, N1064);
and AND4 (N1085, N1063, N462, N609, N866);
or OR2 (N1086, N1082, N484);
nor NOR4 (N1087, N1084, N299, N206, N978);
nand NAND2 (N1088, N1086, N69);
buf BUF1 (N1089, N1073);
xor XOR2 (N1090, N1089, N106);
not NOT1 (N1091, N1090);
and AND2 (N1092, N1087, N626);
nor NOR2 (N1093, N1078, N55);
buf BUF1 (N1094, N1051);
xor XOR2 (N1095, N1093, N373);
nor NOR4 (N1096, N1095, N1028, N863, N1030);
buf BUF1 (N1097, N1088);
and AND4 (N1098, N1091, N499, N513, N57);
and AND4 (N1099, N1048, N1098, N733, N774);
not NOT1 (N1100, N597);
not NOT1 (N1101, N1100);
nor NOR2 (N1102, N1096, N242);
nor NOR4 (N1103, N1074, N1005, N360, N460);
nor NOR3 (N1104, N1101, N71, N430);
nor NOR3 (N1105, N1085, N653, N567);
nor NOR2 (N1106, N1102, N236);
xor XOR2 (N1107, N1103, N2);
buf BUF1 (N1108, N1106);
not NOT1 (N1109, N1094);
not NOT1 (N1110, N1081);
nand NAND4 (N1111, N1109, N906, N707, N364);
buf BUF1 (N1112, N1097);
nor NOR3 (N1113, N1110, N108, N413);
xor XOR2 (N1114, N1107, N751);
nor NOR4 (N1115, N1083, N645, N1079, N185);
nand NAND4 (N1116, N1108, N277, N757, N316);
or OR4 (N1117, N1114, N540, N1015, N932);
nand NAND4 (N1118, N1116, N1083, N66, N26);
or OR4 (N1119, N1118, N103, N951, N652);
xor XOR2 (N1120, N1115, N995);
xor XOR2 (N1121, N1113, N969);
or OR3 (N1122, N1111, N771, N942);
xor XOR2 (N1123, N1104, N845);
or OR2 (N1124, N1121, N1025);
or OR3 (N1125, N1124, N1040, N1015);
or OR4 (N1126, N1120, N1077, N194, N704);
and AND4 (N1127, N1119, N168, N45, N426);
or OR3 (N1128, N1122, N1098, N702);
not NOT1 (N1129, N1099);
not NOT1 (N1130, N1125);
not NOT1 (N1131, N1092);
buf BUF1 (N1132, N1112);
or OR2 (N1133, N1130, N312);
buf BUF1 (N1134, N1128);
xor XOR2 (N1135, N1117, N567);
xor XOR2 (N1136, N1123, N785);
or OR2 (N1137, N1105, N956);
nor NOR4 (N1138, N1127, N741, N166, N91);
not NOT1 (N1139, N1133);
and AND4 (N1140, N1134, N75, N346, N687);
or OR3 (N1141, N1140, N285, N631);
nand NAND2 (N1142, N1131, N175);
nand NAND4 (N1143, N1142, N54, N339, N194);
not NOT1 (N1144, N1141);
xor XOR2 (N1145, N1126, N457);
xor XOR2 (N1146, N1137, N461);
not NOT1 (N1147, N1143);
nand NAND2 (N1148, N1138, N272);
buf BUF1 (N1149, N1146);
xor XOR2 (N1150, N1139, N258);
nor NOR3 (N1151, N1147, N1032, N297);
nor NOR3 (N1152, N1151, N646, N915);
nor NOR4 (N1153, N1129, N163, N520, N873);
nand NAND3 (N1154, N1149, N161, N969);
not NOT1 (N1155, N1144);
nand NAND3 (N1156, N1154, N1122, N600);
xor XOR2 (N1157, N1136, N1108);
nand NAND4 (N1158, N1155, N432, N397, N592);
not NOT1 (N1159, N1148);
nor NOR4 (N1160, N1145, N468, N878, N170);
and AND3 (N1161, N1150, N323, N278);
buf BUF1 (N1162, N1135);
xor XOR2 (N1163, N1162, N828);
and AND4 (N1164, N1153, N1114, N723, N168);
not NOT1 (N1165, N1158);
or OR4 (N1166, N1159, N438, N644, N155);
xor XOR2 (N1167, N1165, N1067);
not NOT1 (N1168, N1160);
nand NAND2 (N1169, N1166, N321);
not NOT1 (N1170, N1168);
buf BUF1 (N1171, N1169);
xor XOR2 (N1172, N1170, N436);
not NOT1 (N1173, N1156);
buf BUF1 (N1174, N1172);
nand NAND4 (N1175, N1163, N434, N464, N463);
or OR4 (N1176, N1171, N142, N100, N1012);
xor XOR2 (N1177, N1132, N711);
not NOT1 (N1178, N1176);
nor NOR4 (N1179, N1175, N383, N509, N529);
nand NAND2 (N1180, N1177, N692);
or OR3 (N1181, N1164, N954, N756);
nor NOR2 (N1182, N1167, N744);
nor NOR3 (N1183, N1152, N289, N581);
and AND4 (N1184, N1157, N549, N786, N603);
not NOT1 (N1185, N1174);
or OR2 (N1186, N1184, N339);
not NOT1 (N1187, N1173);
nor NOR2 (N1188, N1183, N1129);
xor XOR2 (N1189, N1185, N988);
buf BUF1 (N1190, N1161);
nand NAND4 (N1191, N1180, N270, N483, N694);
buf BUF1 (N1192, N1191);
xor XOR2 (N1193, N1188, N303);
nor NOR4 (N1194, N1186, N581, N617, N598);
xor XOR2 (N1195, N1193, N1101);
buf BUF1 (N1196, N1194);
not NOT1 (N1197, N1178);
nor NOR2 (N1198, N1189, N988);
nand NAND3 (N1199, N1182, N1155, N1186);
nand NAND3 (N1200, N1195, N430, N258);
buf BUF1 (N1201, N1187);
and AND3 (N1202, N1199, N1144, N1121);
nand NAND3 (N1203, N1202, N470, N290);
not NOT1 (N1204, N1192);
not NOT1 (N1205, N1197);
xor XOR2 (N1206, N1201, N753);
buf BUF1 (N1207, N1206);
buf BUF1 (N1208, N1198);
buf BUF1 (N1209, N1200);
and AND3 (N1210, N1207, N860, N223);
buf BUF1 (N1211, N1204);
xor XOR2 (N1212, N1205, N999);
and AND4 (N1213, N1212, N843, N27, N1037);
nor NOR2 (N1214, N1190, N143);
buf BUF1 (N1215, N1181);
xor XOR2 (N1216, N1215, N139);
or OR2 (N1217, N1209, N193);
buf BUF1 (N1218, N1214);
nor NOR2 (N1219, N1218, N857);
not NOT1 (N1220, N1179);
nand NAND2 (N1221, N1220, N183);
and AND2 (N1222, N1216, N178);
nor NOR2 (N1223, N1217, N138);
nor NOR2 (N1224, N1208, N811);
or OR4 (N1225, N1213, N1090, N926, N712);
and AND3 (N1226, N1225, N214, N1055);
nand NAND4 (N1227, N1211, N448, N202, N515);
nor NOR3 (N1228, N1219, N914, N605);
or OR2 (N1229, N1222, N787);
nand NAND3 (N1230, N1228, N265, N1037);
or OR2 (N1231, N1227, N654);
not NOT1 (N1232, N1223);
not NOT1 (N1233, N1230);
not NOT1 (N1234, N1224);
buf BUF1 (N1235, N1232);
nand NAND3 (N1236, N1226, N289, N568);
nand NAND2 (N1237, N1235, N856);
nand NAND3 (N1238, N1203, N970, N58);
or OR3 (N1239, N1196, N1091, N501);
buf BUF1 (N1240, N1238);
nor NOR4 (N1241, N1229, N725, N1104, N1075);
or OR4 (N1242, N1239, N726, N1193, N1090);
and AND4 (N1243, N1233, N943, N239, N1054);
buf BUF1 (N1244, N1234);
not NOT1 (N1245, N1210);
buf BUF1 (N1246, N1243);
not NOT1 (N1247, N1241);
buf BUF1 (N1248, N1246);
and AND3 (N1249, N1242, N880, N93);
or OR4 (N1250, N1240, N415, N614, N891);
buf BUF1 (N1251, N1231);
nor NOR2 (N1252, N1251, N1021);
xor XOR2 (N1253, N1248, N97);
not NOT1 (N1254, N1250);
buf BUF1 (N1255, N1244);
and AND3 (N1256, N1254, N994, N1086);
xor XOR2 (N1257, N1256, N1180);
nand NAND4 (N1258, N1245, N490, N940, N295);
not NOT1 (N1259, N1249);
buf BUF1 (N1260, N1221);
nor NOR2 (N1261, N1237, N1209);
nand NAND3 (N1262, N1259, N775, N976);
or OR4 (N1263, N1236, N987, N476, N85);
xor XOR2 (N1264, N1263, N753);
or OR4 (N1265, N1260, N638, N550, N1060);
xor XOR2 (N1266, N1265, N1120);
buf BUF1 (N1267, N1247);
not NOT1 (N1268, N1266);
and AND4 (N1269, N1258, N20, N1046, N937);
not NOT1 (N1270, N1268);
not NOT1 (N1271, N1253);
and AND2 (N1272, N1264, N1210);
nand NAND4 (N1273, N1252, N240, N1208, N366);
xor XOR2 (N1274, N1271, N399);
and AND3 (N1275, N1272, N55, N835);
xor XOR2 (N1276, N1270, N702);
buf BUF1 (N1277, N1262);
buf BUF1 (N1278, N1276);
and AND3 (N1279, N1274, N399, N128);
nor NOR4 (N1280, N1277, N465, N373, N288);
nand NAND3 (N1281, N1278, N261, N89);
xor XOR2 (N1282, N1275, N211);
xor XOR2 (N1283, N1281, N818);
buf BUF1 (N1284, N1273);
and AND2 (N1285, N1269, N1207);
nand NAND4 (N1286, N1279, N1247, N630, N1259);
not NOT1 (N1287, N1255);
xor XOR2 (N1288, N1257, N428);
or OR3 (N1289, N1261, N233, N843);
not NOT1 (N1290, N1267);
nor NOR3 (N1291, N1282, N362, N1068);
nor NOR3 (N1292, N1291, N1143, N451);
not NOT1 (N1293, N1292);
buf BUF1 (N1294, N1287);
nand NAND2 (N1295, N1289, N873);
not NOT1 (N1296, N1294);
nor NOR3 (N1297, N1290, N50, N1131);
xor XOR2 (N1298, N1297, N879);
nand NAND3 (N1299, N1286, N598, N488);
nor NOR2 (N1300, N1284, N183);
nor NOR2 (N1301, N1280, N125);
nand NAND4 (N1302, N1288, N1079, N1026, N152);
xor XOR2 (N1303, N1302, N874);
not NOT1 (N1304, N1295);
not NOT1 (N1305, N1300);
nand NAND3 (N1306, N1285, N1177, N91);
xor XOR2 (N1307, N1303, N479);
or OR4 (N1308, N1301, N413, N859, N1075);
buf BUF1 (N1309, N1296);
and AND3 (N1310, N1304, N594, N1067);
buf BUF1 (N1311, N1298);
xor XOR2 (N1312, N1283, N852);
not NOT1 (N1313, N1310);
or OR4 (N1314, N1299, N545, N850, N177);
nor NOR4 (N1315, N1309, N815, N1103, N1308);
xor XOR2 (N1316, N495, N727);
xor XOR2 (N1317, N1311, N856);
nor NOR4 (N1318, N1315, N1193, N624, N1144);
nor NOR4 (N1319, N1317, N1069, N1052, N711);
nand NAND4 (N1320, N1319, N667, N706, N1207);
nand NAND2 (N1321, N1312, N946);
xor XOR2 (N1322, N1306, N442);
xor XOR2 (N1323, N1316, N643);
and AND4 (N1324, N1318, N726, N457, N1282);
or OR2 (N1325, N1322, N936);
nor NOR4 (N1326, N1307, N1324, N110, N1055);
buf BUF1 (N1327, N404);
nand NAND4 (N1328, N1321, N923, N300, N234);
xor XOR2 (N1329, N1328, N758);
nor NOR3 (N1330, N1325, N663, N324);
and AND4 (N1331, N1330, N1241, N456, N1162);
and AND2 (N1332, N1313, N149);
xor XOR2 (N1333, N1314, N8);
xor XOR2 (N1334, N1333, N63);
or OR3 (N1335, N1331, N1093, N47);
not NOT1 (N1336, N1326);
or OR4 (N1337, N1327, N1259, N440, N283);
nand NAND3 (N1338, N1335, N1190, N1);
or OR2 (N1339, N1323, N1105);
nand NAND4 (N1340, N1337, N1335, N1009, N926);
or OR3 (N1341, N1332, N542, N880);
and AND3 (N1342, N1341, N1034, N1150);
not NOT1 (N1343, N1293);
nand NAND4 (N1344, N1343, N60, N419, N68);
and AND3 (N1345, N1329, N1023, N318);
xor XOR2 (N1346, N1345, N792);
not NOT1 (N1347, N1344);
xor XOR2 (N1348, N1339, N721);
xor XOR2 (N1349, N1305, N1048);
not NOT1 (N1350, N1349);
nor NOR2 (N1351, N1338, N1119);
nand NAND4 (N1352, N1320, N1164, N888, N333);
buf BUF1 (N1353, N1340);
or OR2 (N1354, N1342, N909);
xor XOR2 (N1355, N1352, N364);
buf BUF1 (N1356, N1355);
xor XOR2 (N1357, N1353, N995);
xor XOR2 (N1358, N1334, N1346);
nor NOR3 (N1359, N644, N249, N1212);
nor NOR4 (N1360, N1356, N943, N976, N101);
or OR3 (N1361, N1360, N1102, N560);
and AND4 (N1362, N1357, N63, N557, N719);
buf BUF1 (N1363, N1350);
buf BUF1 (N1364, N1336);
buf BUF1 (N1365, N1362);
and AND3 (N1366, N1364, N369, N396);
not NOT1 (N1367, N1358);
not NOT1 (N1368, N1366);
nor NOR4 (N1369, N1367, N690, N322, N76);
or OR4 (N1370, N1363, N630, N1097, N392);
xor XOR2 (N1371, N1347, N621);
not NOT1 (N1372, N1371);
buf BUF1 (N1373, N1368);
or OR3 (N1374, N1373, N613, N1057);
not NOT1 (N1375, N1354);
nand NAND2 (N1376, N1374, N1359);
buf BUF1 (N1377, N1080);
nand NAND4 (N1378, N1375, N60, N1026, N1060);
nor NOR2 (N1379, N1351, N1328);
buf BUF1 (N1380, N1348);
buf BUF1 (N1381, N1361);
xor XOR2 (N1382, N1379, N996);
nor NOR2 (N1383, N1370, N1243);
xor XOR2 (N1384, N1378, N881);
nor NOR2 (N1385, N1381, N337);
nor NOR4 (N1386, N1369, N1265, N367, N1120);
nand NAND3 (N1387, N1386, N780, N1086);
and AND4 (N1388, N1377, N650, N408, N804);
nand NAND4 (N1389, N1380, N269, N1184, N670);
or OR3 (N1390, N1389, N372, N749);
nand NAND3 (N1391, N1382, N429, N1066);
xor XOR2 (N1392, N1385, N863);
xor XOR2 (N1393, N1390, N166);
xor XOR2 (N1394, N1372, N654);
not NOT1 (N1395, N1365);
not NOT1 (N1396, N1383);
nand NAND4 (N1397, N1393, N397, N1, N206);
xor XOR2 (N1398, N1376, N251);
nand NAND3 (N1399, N1397, N675, N373);
xor XOR2 (N1400, N1387, N1134);
nor NOR4 (N1401, N1400, N425, N1125, N273);
not NOT1 (N1402, N1394);
nor NOR4 (N1403, N1399, N716, N440, N120);
and AND2 (N1404, N1402, N582);
not NOT1 (N1405, N1404);
nand NAND3 (N1406, N1384, N644, N1374);
xor XOR2 (N1407, N1391, N285);
nand NAND2 (N1408, N1401, N866);
and AND4 (N1409, N1392, N789, N641, N632);
nor NOR4 (N1410, N1398, N1141, N788, N563);
nand NAND3 (N1411, N1409, N210, N604);
buf BUF1 (N1412, N1405);
and AND2 (N1413, N1411, N378);
buf BUF1 (N1414, N1406);
buf BUF1 (N1415, N1410);
buf BUF1 (N1416, N1414);
buf BUF1 (N1417, N1395);
buf BUF1 (N1418, N1416);
not NOT1 (N1419, N1412);
nor NOR3 (N1420, N1418, N283, N762);
nand NAND2 (N1421, N1407, N819);
nand NAND2 (N1422, N1421, N179);
or OR2 (N1423, N1413, N1177);
nand NAND2 (N1424, N1388, N1091);
xor XOR2 (N1425, N1423, N1232);
not NOT1 (N1426, N1396);
xor XOR2 (N1427, N1408, N1405);
or OR3 (N1428, N1426, N98, N1325);
nor NOR4 (N1429, N1427, N1223, N82, N829);
and AND4 (N1430, N1403, N1017, N1348, N1136);
or OR4 (N1431, N1429, N79, N200, N1321);
nand NAND2 (N1432, N1422, N942);
or OR3 (N1433, N1424, N1007, N735);
or OR2 (N1434, N1415, N710);
nand NAND3 (N1435, N1432, N979, N606);
and AND2 (N1436, N1417, N326);
xor XOR2 (N1437, N1428, N894);
xor XOR2 (N1438, N1430, N1117);
and AND3 (N1439, N1433, N837, N1428);
not NOT1 (N1440, N1438);
nand NAND4 (N1441, N1437, N128, N87, N755);
xor XOR2 (N1442, N1441, N153);
or OR3 (N1443, N1419, N425, N853);
nor NOR3 (N1444, N1425, N9, N1115);
nor NOR2 (N1445, N1444, N555);
and AND4 (N1446, N1442, N719, N1100, N950);
nand NAND4 (N1447, N1435, N129, N8, N1316);
not NOT1 (N1448, N1445);
nand NAND2 (N1449, N1443, N538);
or OR2 (N1450, N1434, N827);
not NOT1 (N1451, N1420);
nor NOR3 (N1452, N1446, N828, N1308);
xor XOR2 (N1453, N1440, N822);
xor XOR2 (N1454, N1449, N373);
nand NAND2 (N1455, N1453, N1371);
xor XOR2 (N1456, N1439, N926);
xor XOR2 (N1457, N1450, N785);
xor XOR2 (N1458, N1451, N84);
buf BUF1 (N1459, N1448);
not NOT1 (N1460, N1456);
or OR2 (N1461, N1460, N636);
nor NOR4 (N1462, N1454, N925, N1141, N1235);
nand NAND3 (N1463, N1436, N367, N1045);
nand NAND3 (N1464, N1457, N576, N731);
buf BUF1 (N1465, N1461);
not NOT1 (N1466, N1463);
xor XOR2 (N1467, N1452, N893);
nor NOR2 (N1468, N1464, N855);
nand NAND3 (N1469, N1467, N903, N1268);
not NOT1 (N1470, N1458);
xor XOR2 (N1471, N1455, N1175);
not NOT1 (N1472, N1468);
or OR3 (N1473, N1471, N827, N163);
and AND2 (N1474, N1465, N287);
nor NOR3 (N1475, N1459, N120, N838);
nor NOR3 (N1476, N1474, N1085, N639);
buf BUF1 (N1477, N1466);
xor XOR2 (N1478, N1475, N1017);
nor NOR4 (N1479, N1431, N137, N86, N668);
xor XOR2 (N1480, N1472, N1212);
and AND2 (N1481, N1480, N1257);
and AND4 (N1482, N1478, N796, N814, N1437);
buf BUF1 (N1483, N1473);
or OR4 (N1484, N1476, N411, N852, N1036);
or OR4 (N1485, N1477, N760, N36, N469);
nand NAND3 (N1486, N1481, N252, N1041);
xor XOR2 (N1487, N1482, N732);
nor NOR3 (N1488, N1470, N578, N338);
nand NAND3 (N1489, N1487, N291, N262);
xor XOR2 (N1490, N1484, N1396);
or OR2 (N1491, N1483, N1040);
nand NAND3 (N1492, N1462, N130, N213);
or OR4 (N1493, N1492, N445, N819, N1460);
xor XOR2 (N1494, N1491, N137);
nand NAND2 (N1495, N1447, N380);
nand NAND3 (N1496, N1469, N755, N422);
buf BUF1 (N1497, N1495);
or OR3 (N1498, N1497, N242, N1130);
nand NAND3 (N1499, N1490, N1072, N1279);
not NOT1 (N1500, N1489);
and AND4 (N1501, N1499, N445, N1274, N246);
buf BUF1 (N1502, N1501);
not NOT1 (N1503, N1486);
and AND4 (N1504, N1485, N528, N64, N1486);
or OR4 (N1505, N1502, N681, N349, N1333);
or OR4 (N1506, N1503, N50, N908, N1354);
and AND4 (N1507, N1505, N621, N503, N897);
not NOT1 (N1508, N1506);
not NOT1 (N1509, N1498);
or OR2 (N1510, N1488, N613);
nand NAND4 (N1511, N1504, N1120, N667, N1035);
nor NOR2 (N1512, N1496, N588);
nor NOR4 (N1513, N1508, N793, N863, N61);
nor NOR2 (N1514, N1512, N743);
xor XOR2 (N1515, N1510, N1386);
nand NAND2 (N1516, N1511, N376);
not NOT1 (N1517, N1494);
not NOT1 (N1518, N1500);
or OR3 (N1519, N1518, N1265, N553);
not NOT1 (N1520, N1519);
nor NOR3 (N1521, N1509, N999, N1175);
or OR4 (N1522, N1493, N696, N1116, N205);
buf BUF1 (N1523, N1507);
nand NAND3 (N1524, N1520, N1451, N222);
or OR3 (N1525, N1513, N992, N661);
nor NOR3 (N1526, N1514, N538, N628);
buf BUF1 (N1527, N1525);
nand NAND3 (N1528, N1523, N993, N960);
or OR2 (N1529, N1528, N273);
nor NOR3 (N1530, N1517, N711, N579);
not NOT1 (N1531, N1529);
nand NAND4 (N1532, N1526, N483, N981, N147);
and AND2 (N1533, N1532, N231);
xor XOR2 (N1534, N1515, N237);
xor XOR2 (N1535, N1533, N329);
buf BUF1 (N1536, N1521);
or OR3 (N1537, N1531, N786, N42);
and AND4 (N1538, N1530, N387, N145, N1520);
not NOT1 (N1539, N1527);
or OR3 (N1540, N1534, N1507, N157);
and AND3 (N1541, N1516, N140, N573);
nor NOR2 (N1542, N1539, N1105);
xor XOR2 (N1543, N1479, N65);
nor NOR4 (N1544, N1541, N1372, N846, N798);
or OR4 (N1545, N1537, N917, N404, N65);
or OR3 (N1546, N1522, N1385, N212);
or OR4 (N1547, N1524, N433, N763, N1306);
xor XOR2 (N1548, N1540, N535);
xor XOR2 (N1549, N1546, N670);
nand NAND2 (N1550, N1548, N1194);
nand NAND2 (N1551, N1547, N714);
and AND2 (N1552, N1550, N1457);
and AND3 (N1553, N1538, N506, N660);
xor XOR2 (N1554, N1553, N938);
or OR3 (N1555, N1535, N223, N1282);
xor XOR2 (N1556, N1542, N806);
buf BUF1 (N1557, N1543);
nor NOR3 (N1558, N1544, N526, N1527);
nand NAND3 (N1559, N1554, N1361, N1287);
or OR4 (N1560, N1551, N269, N836, N22);
or OR2 (N1561, N1552, N24);
nor NOR4 (N1562, N1558, N586, N116, N74);
buf BUF1 (N1563, N1556);
not NOT1 (N1564, N1545);
nand NAND4 (N1565, N1559, N556, N440, N498);
buf BUF1 (N1566, N1564);
or OR3 (N1567, N1562, N280, N1299);
buf BUF1 (N1568, N1565);
buf BUF1 (N1569, N1568);
buf BUF1 (N1570, N1567);
not NOT1 (N1571, N1536);
and AND3 (N1572, N1557, N1410, N316);
xor XOR2 (N1573, N1566, N58);
not NOT1 (N1574, N1573);
not NOT1 (N1575, N1555);
buf BUF1 (N1576, N1571);
or OR3 (N1577, N1574, N1016, N37);
xor XOR2 (N1578, N1575, N185);
nor NOR4 (N1579, N1578, N1009, N645, N655);
nand NAND3 (N1580, N1570, N1064, N1302);
buf BUF1 (N1581, N1579);
xor XOR2 (N1582, N1549, N575);
not NOT1 (N1583, N1572);
nor NOR3 (N1584, N1569, N1148, N1223);
not NOT1 (N1585, N1560);
nand NAND3 (N1586, N1577, N205, N312);
xor XOR2 (N1587, N1586, N520);
xor XOR2 (N1588, N1576, N232);
buf BUF1 (N1589, N1563);
or OR2 (N1590, N1588, N694);
and AND2 (N1591, N1561, N1003);
xor XOR2 (N1592, N1581, N795);
or OR2 (N1593, N1590, N745);
buf BUF1 (N1594, N1585);
buf BUF1 (N1595, N1592);
or OR3 (N1596, N1583, N1132, N1187);
buf BUF1 (N1597, N1595);
nand NAND2 (N1598, N1591, N339);
or OR2 (N1599, N1584, N1283);
xor XOR2 (N1600, N1596, N695);
or OR3 (N1601, N1598, N150, N1559);
xor XOR2 (N1602, N1599, N670);
buf BUF1 (N1603, N1602);
nand NAND3 (N1604, N1597, N1503, N1381);
nor NOR2 (N1605, N1604, N1411);
and AND3 (N1606, N1593, N1346, N528);
buf BUF1 (N1607, N1606);
nor NOR4 (N1608, N1582, N580, N1450, N1225);
or OR4 (N1609, N1608, N1540, N142, N709);
buf BUF1 (N1610, N1587);
and AND4 (N1611, N1601, N698, N703, N660);
not NOT1 (N1612, N1589);
not NOT1 (N1613, N1600);
nand NAND4 (N1614, N1605, N420, N178, N114);
nand NAND4 (N1615, N1614, N367, N656, N127);
nand NAND3 (N1616, N1611, N433, N1401);
nor NOR2 (N1617, N1613, N1225);
nand NAND2 (N1618, N1580, N1141);
xor XOR2 (N1619, N1615, N456);
xor XOR2 (N1620, N1607, N918);
or OR3 (N1621, N1619, N77, N1389);
xor XOR2 (N1622, N1621, N874);
nand NAND2 (N1623, N1609, N799);
nor NOR4 (N1624, N1594, N745, N879, N1024);
buf BUF1 (N1625, N1603);
nor NOR4 (N1626, N1620, N692, N729, N1126);
nand NAND3 (N1627, N1616, N881, N167);
nand NAND3 (N1628, N1617, N523, N493);
and AND3 (N1629, N1623, N800, N649);
or OR4 (N1630, N1625, N994, N667, N328);
xor XOR2 (N1631, N1622, N1411);
buf BUF1 (N1632, N1612);
xor XOR2 (N1633, N1624, N1473);
xor XOR2 (N1634, N1618, N412);
or OR3 (N1635, N1610, N1428, N788);
or OR4 (N1636, N1631, N1556, N1008, N785);
not NOT1 (N1637, N1636);
xor XOR2 (N1638, N1633, N1099);
nand NAND4 (N1639, N1629, N864, N158, N22);
nand NAND4 (N1640, N1628, N372, N301, N460);
not NOT1 (N1641, N1639);
not NOT1 (N1642, N1626);
or OR4 (N1643, N1637, N1066, N1217, N180);
or OR4 (N1644, N1638, N1172, N1223, N192);
not NOT1 (N1645, N1644);
buf BUF1 (N1646, N1642);
or OR2 (N1647, N1646, N635);
not NOT1 (N1648, N1647);
xor XOR2 (N1649, N1643, N1020);
nor NOR4 (N1650, N1640, N1055, N806, N1505);
nand NAND3 (N1651, N1648, N343, N709);
or OR4 (N1652, N1651, N206, N774, N624);
buf BUF1 (N1653, N1650);
and AND3 (N1654, N1635, N833, N994);
or OR2 (N1655, N1652, N374);
buf BUF1 (N1656, N1641);
xor XOR2 (N1657, N1627, N10);
buf BUF1 (N1658, N1649);
buf BUF1 (N1659, N1655);
and AND4 (N1660, N1656, N1563, N1134, N214);
buf BUF1 (N1661, N1645);
nand NAND4 (N1662, N1658, N1140, N22, N488);
and AND4 (N1663, N1657, N1453, N147, N936);
not NOT1 (N1664, N1662);
buf BUF1 (N1665, N1632);
xor XOR2 (N1666, N1630, N928);
not NOT1 (N1667, N1661);
or OR4 (N1668, N1659, N805, N808, N669);
nor NOR2 (N1669, N1664, N250);
not NOT1 (N1670, N1666);
and AND2 (N1671, N1670, N667);
or OR4 (N1672, N1663, N1058, N1502, N918);
not NOT1 (N1673, N1668);
nand NAND2 (N1674, N1667, N301);
and AND3 (N1675, N1672, N1277, N931);
not NOT1 (N1676, N1675);
nor NOR3 (N1677, N1673, N1131, N285);
and AND3 (N1678, N1634, N222, N77);
xor XOR2 (N1679, N1660, N212);
xor XOR2 (N1680, N1674, N657);
nor NOR2 (N1681, N1677, N66);
nor NOR3 (N1682, N1676, N414, N1051);
and AND2 (N1683, N1678, N125);
or OR3 (N1684, N1669, N253, N1130);
nand NAND4 (N1685, N1671, N999, N895, N36);
or OR2 (N1686, N1665, N1522);
or OR2 (N1687, N1684, N921);
nand NAND2 (N1688, N1683, N574);
xor XOR2 (N1689, N1679, N626);
xor XOR2 (N1690, N1654, N1010);
buf BUF1 (N1691, N1685);
not NOT1 (N1692, N1653);
buf BUF1 (N1693, N1691);
or OR2 (N1694, N1689, N1471);
buf BUF1 (N1695, N1694);
xor XOR2 (N1696, N1688, N1148);
nand NAND2 (N1697, N1680, N1424);
nor NOR2 (N1698, N1695, N1049);
nand NAND2 (N1699, N1681, N972);
xor XOR2 (N1700, N1692, N63);
nor NOR2 (N1701, N1693, N899);
or OR3 (N1702, N1699, N310, N1124);
not NOT1 (N1703, N1690);
not NOT1 (N1704, N1700);
or OR3 (N1705, N1686, N674, N1232);
nand NAND3 (N1706, N1696, N842, N988);
or OR2 (N1707, N1702, N271);
and AND2 (N1708, N1701, N760);
or OR2 (N1709, N1697, N1238);
nand NAND4 (N1710, N1698, N1332, N442, N1658);
buf BUF1 (N1711, N1707);
and AND3 (N1712, N1709, N394, N228);
xor XOR2 (N1713, N1687, N706);
nor NOR2 (N1714, N1682, N512);
and AND3 (N1715, N1713, N506, N800);
or OR2 (N1716, N1715, N597);
xor XOR2 (N1717, N1712, N1235);
buf BUF1 (N1718, N1716);
and AND4 (N1719, N1704, N80, N1238, N1479);
nand NAND3 (N1720, N1714, N150, N95);
or OR4 (N1721, N1711, N2, N1002, N883);
or OR3 (N1722, N1706, N765, N1516);
and AND2 (N1723, N1720, N440);
and AND3 (N1724, N1708, N1235, N1271);
not NOT1 (N1725, N1723);
nor NOR4 (N1726, N1718, N142, N715, N543);
xor XOR2 (N1727, N1721, N138);
buf BUF1 (N1728, N1717);
not NOT1 (N1729, N1710);
nor NOR2 (N1730, N1725, N1239);
nor NOR2 (N1731, N1729, N820);
xor XOR2 (N1732, N1728, N286);
and AND3 (N1733, N1722, N1411, N1424);
nand NAND2 (N1734, N1727, N65);
nor NOR4 (N1735, N1724, N1471, N1187, N1605);
buf BUF1 (N1736, N1732);
xor XOR2 (N1737, N1734, N432);
not NOT1 (N1738, N1735);
not NOT1 (N1739, N1719);
not NOT1 (N1740, N1705);
nor NOR2 (N1741, N1731, N181);
not NOT1 (N1742, N1740);
xor XOR2 (N1743, N1738, N3);
nor NOR4 (N1744, N1737, N1274, N1062, N673);
and AND4 (N1745, N1743, N1487, N913, N1028);
and AND2 (N1746, N1730, N587);
nor NOR3 (N1747, N1745, N733, N1153);
not NOT1 (N1748, N1703);
and AND2 (N1749, N1748, N1258);
and AND2 (N1750, N1726, N318);
and AND2 (N1751, N1749, N1349);
or OR3 (N1752, N1750, N164, N595);
buf BUF1 (N1753, N1752);
not NOT1 (N1754, N1736);
nand NAND2 (N1755, N1733, N1339);
nand NAND3 (N1756, N1746, N77, N839);
and AND3 (N1757, N1753, N859, N1089);
not NOT1 (N1758, N1756);
nor NOR3 (N1759, N1739, N1257, N1370);
nand NAND3 (N1760, N1747, N1738, N596);
or OR4 (N1761, N1754, N363, N495, N303);
not NOT1 (N1762, N1758);
nor NOR4 (N1763, N1757, N720, N347, N1361);
buf BUF1 (N1764, N1761);
nand NAND4 (N1765, N1744, N122, N1019, N669);
nand NAND3 (N1766, N1741, N1679, N1361);
nor NOR4 (N1767, N1759, N1495, N976, N459);
not NOT1 (N1768, N1765);
xor XOR2 (N1769, N1764, N630);
and AND2 (N1770, N1760, N1569);
buf BUF1 (N1771, N1769);
xor XOR2 (N1772, N1770, N671);
and AND3 (N1773, N1768, N447, N1517);
buf BUF1 (N1774, N1742);
or OR3 (N1775, N1774, N638, N851);
and AND3 (N1776, N1767, N1067, N315);
nor NOR4 (N1777, N1773, N1671, N623, N68);
xor XOR2 (N1778, N1763, N1554);
not NOT1 (N1779, N1775);
xor XOR2 (N1780, N1751, N1748);
and AND4 (N1781, N1780, N13, N963, N770);
nor NOR3 (N1782, N1762, N1593, N1416);
buf BUF1 (N1783, N1777);
not NOT1 (N1784, N1783);
xor XOR2 (N1785, N1782, N78);
nand NAND3 (N1786, N1771, N679, N183);
xor XOR2 (N1787, N1776, N1423);
nand NAND3 (N1788, N1779, N1210, N461);
nor NOR2 (N1789, N1781, N740);
nor NOR3 (N1790, N1789, N805, N882);
and AND4 (N1791, N1784, N1617, N339, N582);
nor NOR2 (N1792, N1788, N290);
xor XOR2 (N1793, N1791, N219);
or OR4 (N1794, N1793, N1278, N1154, N1549);
not NOT1 (N1795, N1786);
or OR4 (N1796, N1785, N1729, N602, N1768);
or OR4 (N1797, N1766, N554, N1133, N330);
not NOT1 (N1798, N1778);
xor XOR2 (N1799, N1792, N345);
not NOT1 (N1800, N1787);
buf BUF1 (N1801, N1799);
buf BUF1 (N1802, N1798);
xor XOR2 (N1803, N1755, N1518);
not NOT1 (N1804, N1800);
or OR2 (N1805, N1797, N156);
not NOT1 (N1806, N1772);
xor XOR2 (N1807, N1803, N133);
and AND2 (N1808, N1796, N1245);
or OR3 (N1809, N1804, N1028, N410);
not NOT1 (N1810, N1802);
buf BUF1 (N1811, N1805);
nand NAND2 (N1812, N1806, N230);
xor XOR2 (N1813, N1812, N558);
not NOT1 (N1814, N1807);
not NOT1 (N1815, N1794);
or OR4 (N1816, N1808, N177, N1123, N1777);
nor NOR3 (N1817, N1795, N1068, N1476);
not NOT1 (N1818, N1810);
nor NOR2 (N1819, N1814, N270);
xor XOR2 (N1820, N1815, N1776);
nor NOR2 (N1821, N1790, N741);
xor XOR2 (N1822, N1817, N171);
nand NAND3 (N1823, N1816, N525, N1268);
buf BUF1 (N1824, N1811);
and AND3 (N1825, N1819, N1183, N1516);
xor XOR2 (N1826, N1801, N1384);
xor XOR2 (N1827, N1822, N751);
xor XOR2 (N1828, N1827, N1681);
or OR3 (N1829, N1820, N1458, N1461);
not NOT1 (N1830, N1824);
nand NAND4 (N1831, N1826, N449, N1553, N1476);
nor NOR3 (N1832, N1821, N1083, N215);
nand NAND2 (N1833, N1825, N456);
nand NAND3 (N1834, N1809, N1711, N1222);
or OR2 (N1835, N1830, N1195);
not NOT1 (N1836, N1831);
or OR4 (N1837, N1818, N1519, N127, N1550);
nor NOR3 (N1838, N1832, N733, N1254);
and AND3 (N1839, N1836, N668, N1536);
xor XOR2 (N1840, N1829, N347);
buf BUF1 (N1841, N1833);
nand NAND4 (N1842, N1838, N1624, N1638, N1766);
nor NOR4 (N1843, N1828, N1317, N756, N1572);
and AND4 (N1844, N1837, N943, N563, N1158);
and AND4 (N1845, N1835, N793, N393, N1604);
xor XOR2 (N1846, N1813, N1128);
xor XOR2 (N1847, N1841, N925);
nand NAND2 (N1848, N1842, N129);
xor XOR2 (N1849, N1848, N502);
nor NOR2 (N1850, N1847, N412);
nor NOR4 (N1851, N1844, N291, N131, N1409);
nand NAND2 (N1852, N1849, N355);
xor XOR2 (N1853, N1840, N234);
buf BUF1 (N1854, N1846);
not NOT1 (N1855, N1839);
and AND4 (N1856, N1834, N709, N1787, N710);
buf BUF1 (N1857, N1856);
nand NAND3 (N1858, N1843, N6, N1730);
buf BUF1 (N1859, N1850);
xor XOR2 (N1860, N1854, N562);
not NOT1 (N1861, N1858);
buf BUF1 (N1862, N1859);
buf BUF1 (N1863, N1851);
or OR3 (N1864, N1845, N144, N1190);
xor XOR2 (N1865, N1861, N432);
nor NOR4 (N1866, N1864, N1805, N1116, N1531);
nand NAND4 (N1867, N1865, N1108, N349, N1046);
not NOT1 (N1868, N1852);
and AND4 (N1869, N1823, N1399, N205, N325);
and AND4 (N1870, N1869, N1084, N1680, N965);
or OR3 (N1871, N1853, N1795, N338);
nor NOR3 (N1872, N1863, N385, N814);
not NOT1 (N1873, N1857);
nand NAND3 (N1874, N1862, N1681, N1746);
nand NAND4 (N1875, N1866, N487, N356, N1254);
xor XOR2 (N1876, N1872, N532);
nand NAND4 (N1877, N1867, N984, N56, N700);
not NOT1 (N1878, N1855);
buf BUF1 (N1879, N1873);
nor NOR4 (N1880, N1870, N526, N1031, N1773);
and AND2 (N1881, N1860, N810);
not NOT1 (N1882, N1878);
nor NOR2 (N1883, N1875, N560);
buf BUF1 (N1884, N1881);
and AND2 (N1885, N1882, N549);
nor NOR3 (N1886, N1876, N204, N120);
nand NAND2 (N1887, N1884, N1067);
or OR3 (N1888, N1871, N739, N1595);
or OR3 (N1889, N1887, N523, N1602);
xor XOR2 (N1890, N1886, N1563);
nand NAND2 (N1891, N1879, N798);
nor NOR2 (N1892, N1890, N246);
nand NAND3 (N1893, N1885, N120, N1643);
nor NOR4 (N1894, N1892, N705, N400, N268);
buf BUF1 (N1895, N1891);
xor XOR2 (N1896, N1893, N1721);
nand NAND2 (N1897, N1868, N1483);
not NOT1 (N1898, N1889);
buf BUF1 (N1899, N1874);
nor NOR2 (N1900, N1877, N1466);
buf BUF1 (N1901, N1883);
buf BUF1 (N1902, N1897);
nand NAND2 (N1903, N1901, N367);
nor NOR2 (N1904, N1880, N438);
buf BUF1 (N1905, N1896);
xor XOR2 (N1906, N1898, N1093);
nand NAND2 (N1907, N1900, N665);
xor XOR2 (N1908, N1902, N810);
xor XOR2 (N1909, N1904, N1341);
xor XOR2 (N1910, N1908, N1540);
or OR4 (N1911, N1888, N491, N1380, N1781);
and AND2 (N1912, N1910, N1239);
buf BUF1 (N1913, N1906);
buf BUF1 (N1914, N1903);
or OR4 (N1915, N1895, N1015, N221, N1607);
not NOT1 (N1916, N1894);
not NOT1 (N1917, N1914);
buf BUF1 (N1918, N1905);
nand NAND2 (N1919, N1917, N608);
and AND3 (N1920, N1911, N1098, N1829);
and AND2 (N1921, N1920, N532);
and AND3 (N1922, N1913, N1716, N1244);
or OR3 (N1923, N1916, N1459, N1096);
xor XOR2 (N1924, N1922, N454);
nand NAND4 (N1925, N1921, N600, N950, N1120);
nand NAND2 (N1926, N1919, N1726);
and AND4 (N1927, N1924, N811, N850, N1340);
or OR3 (N1928, N1915, N165, N100);
nor NOR3 (N1929, N1909, N329, N432);
xor XOR2 (N1930, N1929, N657);
nand NAND3 (N1931, N1918, N217, N1678);
and AND4 (N1932, N1928, N434, N745, N526);
nand NAND4 (N1933, N1925, N889, N1882, N1622);
or OR2 (N1934, N1927, N309);
and AND3 (N1935, N1926, N866, N614);
xor XOR2 (N1936, N1907, N153);
xor XOR2 (N1937, N1923, N28);
buf BUF1 (N1938, N1935);
or OR2 (N1939, N1936, N187);
buf BUF1 (N1940, N1912);
nor NOR4 (N1941, N1940, N1357, N1333, N1777);
buf BUF1 (N1942, N1930);
or OR4 (N1943, N1941, N509, N1054, N510);
xor XOR2 (N1944, N1943, N1510);
buf BUF1 (N1945, N1934);
or OR4 (N1946, N1945, N827, N504, N696);
or OR2 (N1947, N1937, N1131);
not NOT1 (N1948, N1944);
not NOT1 (N1949, N1931);
and AND4 (N1950, N1942, N231, N1026, N902);
buf BUF1 (N1951, N1899);
or OR4 (N1952, N1949, N209, N1034, N179);
buf BUF1 (N1953, N1950);
not NOT1 (N1954, N1939);
buf BUF1 (N1955, N1932);
and AND4 (N1956, N1953, N308, N1181, N884);
xor XOR2 (N1957, N1948, N1148);
xor XOR2 (N1958, N1951, N1452);
buf BUF1 (N1959, N1954);
buf BUF1 (N1960, N1946);
not NOT1 (N1961, N1960);
xor XOR2 (N1962, N1956, N176);
buf BUF1 (N1963, N1952);
not NOT1 (N1964, N1955);
not NOT1 (N1965, N1957);
nor NOR3 (N1966, N1963, N917, N509);
not NOT1 (N1967, N1962);
xor XOR2 (N1968, N1958, N520);
not NOT1 (N1969, N1968);
nor NOR2 (N1970, N1969, N1914);
nor NOR2 (N1971, N1947, N1540);
and AND4 (N1972, N1964, N353, N1710, N1386);
or OR3 (N1973, N1938, N440, N1815);
xor XOR2 (N1974, N1933, N968);
nor NOR3 (N1975, N1966, N1319, N1188);
not NOT1 (N1976, N1972);
buf BUF1 (N1977, N1965);
xor XOR2 (N1978, N1959, N1425);
and AND2 (N1979, N1971, N88);
not NOT1 (N1980, N1976);
or OR4 (N1981, N1961, N623, N1744, N464);
nor NOR2 (N1982, N1980, N569);
and AND4 (N1983, N1977, N349, N479, N809);
or OR2 (N1984, N1978, N1532);
buf BUF1 (N1985, N1979);
and AND3 (N1986, N1982, N1495, N1711);
xor XOR2 (N1987, N1981, N1575);
nor NOR3 (N1988, N1984, N1142, N1276);
nor NOR3 (N1989, N1967, N1780, N248);
buf BUF1 (N1990, N1975);
not NOT1 (N1991, N1983);
nand NAND2 (N1992, N1973, N1031);
xor XOR2 (N1993, N1992, N1821);
nor NOR3 (N1994, N1990, N169, N886);
and AND3 (N1995, N1988, N1790, N1093);
or OR2 (N1996, N1986, N260);
or OR3 (N1997, N1974, N1469, N1062);
buf BUF1 (N1998, N1994);
nor NOR3 (N1999, N1996, N536, N1581);
nand NAND4 (N2000, N1970, N949, N1633, N1836);
xor XOR2 (N2001, N1999, N1968);
or OR2 (N2002, N1993, N779);
not NOT1 (N2003, N2000);
xor XOR2 (N2004, N1995, N1687);
nor NOR3 (N2005, N2002, N391, N996);
xor XOR2 (N2006, N1989, N560);
or OR2 (N2007, N1991, N1798);
nor NOR3 (N2008, N2004, N98, N1856);
not NOT1 (N2009, N2007);
or OR4 (N2010, N2009, N1311, N1017, N498);
nand NAND4 (N2011, N1987, N1857, N363, N1962);
and AND4 (N2012, N2010, N1909, N1484, N618);
buf BUF1 (N2013, N2012);
or OR3 (N2014, N2011, N1999, N1777);
nor NOR2 (N2015, N1998, N1485);
nand NAND3 (N2016, N2008, N998, N177);
and AND4 (N2017, N1997, N552, N990, N620);
xor XOR2 (N2018, N2003, N1447);
or OR4 (N2019, N2001, N319, N596, N1982);
and AND2 (N2020, N2005, N364);
buf BUF1 (N2021, N1985);
xor XOR2 (N2022, N2017, N1576);
or OR4 (N2023, N2015, N1772, N216, N2001);
xor XOR2 (N2024, N2006, N1943);
not NOT1 (N2025, N2022);
nor NOR3 (N2026, N2016, N372, N948);
and AND3 (N2027, N2026, N6, N42);
and AND2 (N2028, N2018, N64);
buf BUF1 (N2029, N2019);
or OR4 (N2030, N2027, N258, N1514, N21);
xor XOR2 (N2031, N2020, N861);
buf BUF1 (N2032, N2029);
nor NOR2 (N2033, N2032, N205);
nand NAND2 (N2034, N2028, N1996);
not NOT1 (N2035, N2030);
or OR3 (N2036, N2034, N113, N1599);
xor XOR2 (N2037, N2025, N921);
xor XOR2 (N2038, N2023, N1217);
and AND2 (N2039, N2014, N1344);
buf BUF1 (N2040, N2035);
buf BUF1 (N2041, N2024);
nor NOR2 (N2042, N2039, N1622);
nand NAND4 (N2043, N2036, N174, N1124, N1086);
not NOT1 (N2044, N2040);
buf BUF1 (N2045, N2037);
buf BUF1 (N2046, N2045);
nor NOR4 (N2047, N2046, N608, N1725, N572);
or OR3 (N2048, N2044, N1746, N56);
buf BUF1 (N2049, N2033);
nor NOR4 (N2050, N2049, N1602, N308, N2035);
xor XOR2 (N2051, N2048, N1447);
not NOT1 (N2052, N2021);
buf BUF1 (N2053, N2050);
buf BUF1 (N2054, N2053);
not NOT1 (N2055, N2038);
or OR3 (N2056, N2055, N1912, N183);
or OR3 (N2057, N2041, N310, N833);
nand NAND3 (N2058, N2031, N579, N236);
nor NOR3 (N2059, N2013, N1758, N1889);
nand NAND2 (N2060, N2051, N1111);
nand NAND2 (N2061, N2054, N1724);
nor NOR4 (N2062, N2056, N348, N271, N974);
and AND4 (N2063, N2047, N1544, N1006, N199);
and AND4 (N2064, N2058, N1158, N1034, N134);
and AND4 (N2065, N2062, N785, N1305, N1971);
and AND4 (N2066, N2059, N100, N953, N1303);
xor XOR2 (N2067, N2065, N267);
nor NOR3 (N2068, N2042, N1911, N346);
nand NAND3 (N2069, N2068, N1355, N917);
nor NOR4 (N2070, N2063, N1265, N1877, N210);
nor NOR4 (N2071, N2061, N460, N1752, N1796);
xor XOR2 (N2072, N2070, N671);
or OR2 (N2073, N2072, N433);
or OR4 (N2074, N2057, N350, N1150, N1112);
xor XOR2 (N2075, N2060, N37);
or OR3 (N2076, N2066, N1096, N1953);
nand NAND2 (N2077, N2073, N394);
buf BUF1 (N2078, N2071);
nand NAND4 (N2079, N2064, N1490, N1484, N776);
xor XOR2 (N2080, N2077, N807);
not NOT1 (N2081, N2069);
nand NAND4 (N2082, N2076, N999, N477, N1009);
not NOT1 (N2083, N2082);
and AND3 (N2084, N2078, N1410, N918);
or OR2 (N2085, N2081, N2058);
or OR4 (N2086, N2085, N850, N1437, N679);
or OR3 (N2087, N2067, N600, N62);
buf BUF1 (N2088, N2052);
or OR3 (N2089, N2080, N1489, N182);
and AND3 (N2090, N2088, N341, N824);
xor XOR2 (N2091, N2084, N1052);
or OR3 (N2092, N2043, N670, N495);
or OR2 (N2093, N2090, N1628);
or OR2 (N2094, N2086, N386);
buf BUF1 (N2095, N2094);
xor XOR2 (N2096, N2095, N955);
buf BUF1 (N2097, N2093);
not NOT1 (N2098, N2079);
buf BUF1 (N2099, N2074);
and AND2 (N2100, N2096, N88);
nand NAND2 (N2101, N2100, N1679);
not NOT1 (N2102, N2091);
nor NOR2 (N2103, N2097, N1569);
and AND4 (N2104, N2098, N1635, N841, N123);
nand NAND4 (N2105, N2104, N1477, N556, N12);
xor XOR2 (N2106, N2102, N336);
xor XOR2 (N2107, N2083, N114);
nor NOR3 (N2108, N2101, N1083, N2050);
nor NOR2 (N2109, N2103, N119);
nand NAND2 (N2110, N2089, N1058);
nand NAND2 (N2111, N2108, N1129);
buf BUF1 (N2112, N2075);
nand NAND2 (N2113, N2111, N1413);
not NOT1 (N2114, N2106);
or OR3 (N2115, N2109, N1603, N1372);
not NOT1 (N2116, N2110);
not NOT1 (N2117, N2114);
buf BUF1 (N2118, N2107);
buf BUF1 (N2119, N2113);
or OR3 (N2120, N2117, N628, N782);
and AND3 (N2121, N2087, N1033, N382);
nor NOR4 (N2122, N2118, N814, N1114, N261);
and AND3 (N2123, N2115, N12, N1550);
xor XOR2 (N2124, N2120, N1011);
or OR3 (N2125, N2123, N803, N1829);
and AND3 (N2126, N2119, N1254, N1806);
or OR2 (N2127, N2126, N1293);
nand NAND2 (N2128, N2116, N1532);
xor XOR2 (N2129, N2121, N852);
xor XOR2 (N2130, N2127, N1766);
or OR2 (N2131, N2125, N749);
nand NAND4 (N2132, N2128, N856, N120, N2125);
and AND3 (N2133, N2092, N1308, N1246);
xor XOR2 (N2134, N2112, N687);
not NOT1 (N2135, N2130);
buf BUF1 (N2136, N2132);
or OR4 (N2137, N2131, N850, N1806, N1464);
buf BUF1 (N2138, N2099);
not NOT1 (N2139, N2138);
buf BUF1 (N2140, N2139);
xor XOR2 (N2141, N2140, N992);
buf BUF1 (N2142, N2133);
buf BUF1 (N2143, N2105);
nor NOR4 (N2144, N2137, N1316, N1524, N1586);
buf BUF1 (N2145, N2124);
xor XOR2 (N2146, N2135, N556);
buf BUF1 (N2147, N2144);
and AND2 (N2148, N2142, N1283);
not NOT1 (N2149, N2136);
and AND4 (N2150, N2149, N1106, N444, N766);
nor NOR3 (N2151, N2122, N1167, N822);
or OR3 (N2152, N2151, N703, N810);
xor XOR2 (N2153, N2145, N52);
or OR4 (N2154, N2146, N611, N1060, N1311);
nand NAND2 (N2155, N2153, N450);
not NOT1 (N2156, N2154);
buf BUF1 (N2157, N2150);
buf BUF1 (N2158, N2152);
xor XOR2 (N2159, N2155, N1243);
or OR2 (N2160, N2129, N256);
not NOT1 (N2161, N2148);
nand NAND4 (N2162, N2160, N313, N1908, N281);
and AND3 (N2163, N2157, N1559, N131);
nor NOR4 (N2164, N2143, N540, N1345, N1264);
not NOT1 (N2165, N2156);
not NOT1 (N2166, N2163);
not NOT1 (N2167, N2134);
and AND4 (N2168, N2161, N1724, N1149, N1633);
nor NOR2 (N2169, N2147, N1630);
and AND4 (N2170, N2166, N526, N808, N1707);
xor XOR2 (N2171, N2170, N167);
nor NOR2 (N2172, N2164, N1135);
not NOT1 (N2173, N2141);
buf BUF1 (N2174, N2167);
buf BUF1 (N2175, N2174);
not NOT1 (N2176, N2165);
nand NAND3 (N2177, N2173, N1137, N1826);
or OR2 (N2178, N2168, N464);
nor NOR3 (N2179, N2158, N266, N173);
or OR3 (N2180, N2171, N1615, N466);
nand NAND3 (N2181, N2180, N621, N727);
xor XOR2 (N2182, N2178, N637);
xor XOR2 (N2183, N2159, N1672);
nand NAND4 (N2184, N2183, N2056, N914, N370);
nor NOR4 (N2185, N2162, N1923, N288, N1582);
xor XOR2 (N2186, N2177, N697);
or OR3 (N2187, N2172, N1169, N614);
nand NAND4 (N2188, N2184, N174, N1187, N1535);
xor XOR2 (N2189, N2185, N1104);
nand NAND4 (N2190, N2181, N150, N160, N1376);
nor NOR3 (N2191, N2188, N1383, N204);
buf BUF1 (N2192, N2191);
xor XOR2 (N2193, N2192, N862);
nor NOR3 (N2194, N2193, N984, N1926);
or OR4 (N2195, N2176, N1855, N1049, N535);
and AND2 (N2196, N2195, N736);
buf BUF1 (N2197, N2189);
and AND4 (N2198, N2197, N927, N1157, N467);
and AND2 (N2199, N2179, N1552);
buf BUF1 (N2200, N2199);
xor XOR2 (N2201, N2200, N1400);
or OR3 (N2202, N2196, N1227, N829);
xor XOR2 (N2203, N2182, N1995);
not NOT1 (N2204, N2175);
buf BUF1 (N2205, N2204);
nand NAND3 (N2206, N2190, N1030, N599);
nand NAND4 (N2207, N2201, N336, N926, N1125);
and AND3 (N2208, N2194, N194, N2036);
xor XOR2 (N2209, N2198, N1719);
and AND4 (N2210, N2209, N2073, N1409, N885);
xor XOR2 (N2211, N2205, N535);
and AND2 (N2212, N2207, N1905);
nand NAND2 (N2213, N2203, N52);
and AND2 (N2214, N2206, N1868);
and AND3 (N2215, N2187, N346, N909);
xor XOR2 (N2216, N2208, N1526);
and AND2 (N2217, N2212, N390);
xor XOR2 (N2218, N2202, N2125);
nor NOR3 (N2219, N2218, N335, N1709);
xor XOR2 (N2220, N2211, N2044);
buf BUF1 (N2221, N2217);
nand NAND4 (N2222, N2169, N793, N1204, N402);
nor NOR2 (N2223, N2215, N2197);
nand NAND3 (N2224, N2223, N3, N147);
not NOT1 (N2225, N2221);
not NOT1 (N2226, N2214);
buf BUF1 (N2227, N2213);
or OR4 (N2228, N2226, N623, N607, N1141);
nand NAND4 (N2229, N2186, N908, N15, N583);
nand NAND3 (N2230, N2216, N168, N1577);
xor XOR2 (N2231, N2230, N1815);
nand NAND3 (N2232, N2228, N2171, N1988);
or OR4 (N2233, N2227, N617, N1388, N164);
or OR2 (N2234, N2233, N124);
and AND2 (N2235, N2210, N220);
not NOT1 (N2236, N2229);
xor XOR2 (N2237, N2224, N620);
buf BUF1 (N2238, N2222);
or OR4 (N2239, N2236, N2185, N1741, N938);
not NOT1 (N2240, N2234);
xor XOR2 (N2241, N2225, N211);
xor XOR2 (N2242, N2232, N377);
nand NAND3 (N2243, N2220, N1498, N276);
and AND3 (N2244, N2239, N1522, N1146);
nor NOR4 (N2245, N2241, N813, N723, N892);
not NOT1 (N2246, N2243);
nor NOR2 (N2247, N2242, N2052);
or OR2 (N2248, N2238, N15);
not NOT1 (N2249, N2219);
nand NAND4 (N2250, N2240, N820, N424, N457);
and AND4 (N2251, N2247, N927, N2238, N39);
nor NOR3 (N2252, N2246, N181, N1569);
xor XOR2 (N2253, N2231, N1087);
nor NOR3 (N2254, N2249, N646, N94);
xor XOR2 (N2255, N2253, N1003);
nor NOR3 (N2256, N2244, N1011, N60);
or OR4 (N2257, N2255, N1024, N1000, N808);
buf BUF1 (N2258, N2250);
or OR3 (N2259, N2235, N2123, N2089);
and AND2 (N2260, N2259, N965);
not NOT1 (N2261, N2237);
or OR3 (N2262, N2258, N561, N1034);
nor NOR4 (N2263, N2245, N2080, N506, N1875);
nor NOR4 (N2264, N2248, N2112, N1747, N1313);
not NOT1 (N2265, N2262);
buf BUF1 (N2266, N2256);
xor XOR2 (N2267, N2265, N1517);
buf BUF1 (N2268, N2257);
or OR4 (N2269, N2254, N1196, N467, N60);
buf BUF1 (N2270, N2264);
and AND4 (N2271, N2269, N1577, N967, N1994);
and AND3 (N2272, N2266, N1729, N1063);
not NOT1 (N2273, N2260);
buf BUF1 (N2274, N2268);
nand NAND3 (N2275, N2267, N1417, N111);
not NOT1 (N2276, N2252);
xor XOR2 (N2277, N2263, N819);
or OR2 (N2278, N2275, N1977);
nand NAND3 (N2279, N2276, N1122, N1813);
buf BUF1 (N2280, N2251);
nor NOR3 (N2281, N2280, N1033, N1346);
or OR2 (N2282, N2281, N559);
xor XOR2 (N2283, N2278, N1091);
buf BUF1 (N2284, N2274);
or OR4 (N2285, N2270, N266, N1632, N1562);
xor XOR2 (N2286, N2273, N1212);
not NOT1 (N2287, N2271);
not NOT1 (N2288, N2279);
not NOT1 (N2289, N2285);
nand NAND2 (N2290, N2286, N1463);
and AND2 (N2291, N2284, N830);
not NOT1 (N2292, N2288);
nand NAND2 (N2293, N2291, N2018);
nand NAND2 (N2294, N2293, N181);
not NOT1 (N2295, N2272);
or OR3 (N2296, N2295, N681, N515);
or OR3 (N2297, N2261, N1400, N39);
and AND4 (N2298, N2282, N1816, N270, N908);
or OR4 (N2299, N2296, N705, N2254, N1492);
or OR4 (N2300, N2297, N100, N1312, N554);
buf BUF1 (N2301, N2298);
and AND3 (N2302, N2299, N1136, N1241);
nand NAND2 (N2303, N2287, N1504);
not NOT1 (N2304, N2277);
nor NOR3 (N2305, N2303, N693, N483);
and AND4 (N2306, N2300, N2304, N815, N93);
not NOT1 (N2307, N1134);
not NOT1 (N2308, N2292);
xor XOR2 (N2309, N2290, N244);
and AND3 (N2310, N2289, N1192, N1239);
xor XOR2 (N2311, N2306, N146);
buf BUF1 (N2312, N2308);
nand NAND4 (N2313, N2294, N1841, N1947, N366);
or OR4 (N2314, N2312, N899, N572, N2257);
and AND2 (N2315, N2302, N174);
nor NOR3 (N2316, N2311, N1356, N988);
buf BUF1 (N2317, N2315);
nand NAND2 (N2318, N2310, N2136);
not NOT1 (N2319, N2316);
xor XOR2 (N2320, N2313, N1433);
nor NOR2 (N2321, N2314, N1651);
or OR3 (N2322, N2319, N592, N293);
not NOT1 (N2323, N2301);
or OR2 (N2324, N2307, N200);
or OR4 (N2325, N2309, N1759, N677, N291);
nand NAND2 (N2326, N2324, N2255);
and AND2 (N2327, N2321, N1398);
nor NOR4 (N2328, N2305, N699, N469, N481);
buf BUF1 (N2329, N2322);
xor XOR2 (N2330, N2328, N2229);
xor XOR2 (N2331, N2317, N2030);
nor NOR2 (N2332, N2327, N1737);
xor XOR2 (N2333, N2318, N2263);
buf BUF1 (N2334, N2333);
nor NOR3 (N2335, N2325, N251, N513);
xor XOR2 (N2336, N2320, N2309);
nor NOR2 (N2337, N2326, N2008);
not NOT1 (N2338, N2283);
nor NOR4 (N2339, N2332, N240, N120, N805);
and AND3 (N2340, N2331, N509, N2203);
nand NAND2 (N2341, N2338, N417);
buf BUF1 (N2342, N2334);
and AND4 (N2343, N2340, N477, N406, N1811);
and AND4 (N2344, N2335, N1599, N1865, N806);
nor NOR3 (N2345, N2342, N1639, N2283);
buf BUF1 (N2346, N2343);
xor XOR2 (N2347, N2339, N1137);
or OR4 (N2348, N2336, N1812, N1599, N1799);
buf BUF1 (N2349, N2341);
nand NAND2 (N2350, N2345, N714);
or OR4 (N2351, N2349, N1906, N1534, N700);
xor XOR2 (N2352, N2348, N2067);
nand NAND4 (N2353, N2330, N505, N1580, N750);
and AND3 (N2354, N2344, N242, N1985);
or OR4 (N2355, N2323, N1251, N438, N1078);
and AND2 (N2356, N2354, N1528);
nor NOR4 (N2357, N2350, N464, N413, N1336);
and AND4 (N2358, N2353, N306, N2201, N1047);
or OR4 (N2359, N2358, N1951, N2211, N489);
xor XOR2 (N2360, N2352, N1268);
nor NOR4 (N2361, N2360, N604, N2008, N287);
nor NOR3 (N2362, N2357, N1314, N309);
nor NOR4 (N2363, N2337, N123, N1389, N629);
nand NAND4 (N2364, N2346, N234, N1223, N1805);
nand NAND3 (N2365, N2329, N2005, N1109);
xor XOR2 (N2366, N2365, N1531);
and AND2 (N2367, N2361, N269);
or OR2 (N2368, N2359, N1126);
and AND2 (N2369, N2368, N1886);
nor NOR2 (N2370, N2347, N1244);
or OR3 (N2371, N2364, N1012, N405);
not NOT1 (N2372, N2370);
nor NOR2 (N2373, N2369, N898);
xor XOR2 (N2374, N2371, N231);
xor XOR2 (N2375, N2367, N2100);
nand NAND2 (N2376, N2372, N1934);
nor NOR3 (N2377, N2366, N2287, N1554);
xor XOR2 (N2378, N2375, N707);
or OR3 (N2379, N2351, N960, N43);
buf BUF1 (N2380, N2363);
xor XOR2 (N2381, N2378, N987);
nand NAND4 (N2382, N2374, N877, N111, N2299);
xor XOR2 (N2383, N2380, N1190);
not NOT1 (N2384, N2382);
nor NOR4 (N2385, N2355, N238, N1193, N2052);
not NOT1 (N2386, N2381);
nand NAND3 (N2387, N2386, N2202, N1972);
nor NOR3 (N2388, N2373, N2290, N154);
buf BUF1 (N2389, N2383);
and AND4 (N2390, N2376, N1334, N568, N1656);
not NOT1 (N2391, N2388);
nor NOR2 (N2392, N2387, N457);
xor XOR2 (N2393, N2384, N155);
buf BUF1 (N2394, N2377);
buf BUF1 (N2395, N2356);
nor NOR2 (N2396, N2389, N264);
buf BUF1 (N2397, N2390);
or OR4 (N2398, N2397, N2338, N77, N2109);
not NOT1 (N2399, N2362);
xor XOR2 (N2400, N2395, N82);
nor NOR2 (N2401, N2396, N603);
xor XOR2 (N2402, N2401, N412);
nand NAND4 (N2403, N2392, N694, N1099, N1104);
or OR3 (N2404, N2402, N1235, N33);
or OR2 (N2405, N2393, N2223);
nand NAND4 (N2406, N2398, N2002, N33, N400);
buf BUF1 (N2407, N2394);
nor NOR3 (N2408, N2379, N2028, N1079);
not NOT1 (N2409, N2391);
not NOT1 (N2410, N2408);
not NOT1 (N2411, N2406);
not NOT1 (N2412, N2404);
buf BUF1 (N2413, N2409);
and AND4 (N2414, N2399, N1146, N1749, N1291);
nand NAND3 (N2415, N2412, N1526, N701);
nand NAND2 (N2416, N2405, N350);
and AND2 (N2417, N2414, N77);
or OR3 (N2418, N2413, N2131, N1491);
nor NOR4 (N2419, N2411, N2361, N1787, N2143);
xor XOR2 (N2420, N2417, N760);
nand NAND3 (N2421, N2420, N2389, N2102);
or OR2 (N2422, N2410, N1220);
not NOT1 (N2423, N2418);
not NOT1 (N2424, N2416);
nand NAND4 (N2425, N2415, N1375, N378, N601);
nand NAND3 (N2426, N2421, N1721, N1677);
xor XOR2 (N2427, N2423, N1888);
nand NAND3 (N2428, N2403, N1726, N953);
not NOT1 (N2429, N2426);
or OR3 (N2430, N2422, N493, N1372);
and AND2 (N2431, N2424, N588);
or OR4 (N2432, N2407, N2307, N1001, N1169);
and AND2 (N2433, N2431, N1221);
nor NOR2 (N2434, N2428, N1858);
not NOT1 (N2435, N2429);
buf BUF1 (N2436, N2425);
and AND2 (N2437, N2400, N1402);
and AND2 (N2438, N2437, N2090);
nor NOR4 (N2439, N2419, N1327, N462, N2188);
and AND4 (N2440, N2439, N2222, N1850, N1539);
not NOT1 (N2441, N2438);
xor XOR2 (N2442, N2436, N898);
buf BUF1 (N2443, N2441);
buf BUF1 (N2444, N2385);
nor NOR2 (N2445, N2434, N1453);
nand NAND2 (N2446, N2427, N1387);
xor XOR2 (N2447, N2443, N2220);
nor NOR2 (N2448, N2435, N1438);
not NOT1 (N2449, N2430);
nor NOR2 (N2450, N2445, N1157);
or OR2 (N2451, N2446, N339);
xor XOR2 (N2452, N2447, N1509);
and AND2 (N2453, N2449, N152);
nor NOR4 (N2454, N2450, N1985, N1346, N800);
xor XOR2 (N2455, N2451, N2149);
not NOT1 (N2456, N2454);
buf BUF1 (N2457, N2442);
buf BUF1 (N2458, N2455);
nor NOR2 (N2459, N2453, N1931);
or OR3 (N2460, N2458, N590, N499);
buf BUF1 (N2461, N2432);
nor NOR4 (N2462, N2459, N1788, N1795, N1273);
or OR2 (N2463, N2457, N716);
buf BUF1 (N2464, N2462);
or OR3 (N2465, N2452, N1502, N132);
or OR3 (N2466, N2465, N1590, N1535);
and AND3 (N2467, N2466, N2059, N1901);
and AND2 (N2468, N2464, N1219);
nor NOR4 (N2469, N2467, N894, N827, N2106);
not NOT1 (N2470, N2440);
xor XOR2 (N2471, N2469, N258);
and AND2 (N2472, N2470, N2436);
xor XOR2 (N2473, N2444, N282);
xor XOR2 (N2474, N2463, N1222);
buf BUF1 (N2475, N2461);
nor NOR2 (N2476, N2475, N271);
nor NOR3 (N2477, N2468, N1571, N1255);
or OR4 (N2478, N2476, N2120, N1799, N1368);
xor XOR2 (N2479, N2474, N1942);
nor NOR4 (N2480, N2473, N2384, N1677, N1);
not NOT1 (N2481, N2471);
and AND3 (N2482, N2478, N222, N2132);
xor XOR2 (N2483, N2456, N197);
and AND4 (N2484, N2480, N2115, N2091, N2062);
nor NOR3 (N2485, N2483, N728, N796);
or OR2 (N2486, N2433, N99);
xor XOR2 (N2487, N2482, N1266);
nand NAND3 (N2488, N2479, N2139, N2383);
buf BUF1 (N2489, N2485);
nand NAND4 (N2490, N2460, N2111, N685, N445);
and AND2 (N2491, N2488, N25);
nor NOR4 (N2492, N2486, N1887, N1032, N1257);
or OR4 (N2493, N2490, N36, N356, N254);
and AND4 (N2494, N2491, N224, N902, N1708);
or OR3 (N2495, N2492, N1500, N2298);
not NOT1 (N2496, N2489);
xor XOR2 (N2497, N2487, N653);
nand NAND2 (N2498, N2481, N1360);
nand NAND3 (N2499, N2484, N1028, N1780);
or OR2 (N2500, N2477, N591);
xor XOR2 (N2501, N2499, N818);
not NOT1 (N2502, N2496);
xor XOR2 (N2503, N2501, N312);
and AND4 (N2504, N2497, N744, N1678, N415);
xor XOR2 (N2505, N2503, N2464);
buf BUF1 (N2506, N2505);
xor XOR2 (N2507, N2506, N110);
nand NAND3 (N2508, N2498, N415, N2037);
and AND2 (N2509, N2472, N278);
and AND4 (N2510, N2495, N2316, N614, N2476);
not NOT1 (N2511, N2510);
or OR4 (N2512, N2493, N18, N1694, N1872);
nor NOR4 (N2513, N2500, N2069, N454, N182);
xor XOR2 (N2514, N2502, N981);
not NOT1 (N2515, N2494);
nand NAND4 (N2516, N2513, N1134, N1781, N895);
or OR3 (N2517, N2516, N254, N919);
or OR3 (N2518, N2509, N1791, N1711);
not NOT1 (N2519, N2512);
buf BUF1 (N2520, N2508);
buf BUF1 (N2521, N2519);
buf BUF1 (N2522, N2518);
and AND3 (N2523, N2517, N803, N701);
nand NAND2 (N2524, N2521, N2492);
or OR2 (N2525, N2522, N675);
xor XOR2 (N2526, N2448, N393);
nand NAND2 (N2527, N2507, N1148);
nor NOR4 (N2528, N2520, N2480, N298, N2390);
or OR4 (N2529, N2523, N1298, N1252, N19);
or OR2 (N2530, N2524, N1597);
or OR2 (N2531, N2514, N2182);
buf BUF1 (N2532, N2515);
buf BUF1 (N2533, N2529);
nand NAND2 (N2534, N2526, N1172);
nand NAND3 (N2535, N2534, N1752, N413);
and AND3 (N2536, N2532, N1770, N1344);
or OR4 (N2537, N2528, N469, N676, N789);
or OR4 (N2538, N2530, N210, N884, N2396);
not NOT1 (N2539, N2531);
xor XOR2 (N2540, N2539, N692);
nor NOR4 (N2541, N2540, N2136, N574, N2290);
nand NAND3 (N2542, N2533, N1757, N601);
and AND2 (N2543, N2538, N1069);
nand NAND2 (N2544, N2537, N1112);
buf BUF1 (N2545, N2541);
nor NOR3 (N2546, N2545, N1, N1706);
or OR4 (N2547, N2504, N27, N1784, N1872);
nand NAND4 (N2548, N2543, N284, N1325, N2093);
xor XOR2 (N2549, N2544, N1932);
not NOT1 (N2550, N2536);
and AND3 (N2551, N2548, N321, N787);
and AND3 (N2552, N2546, N1970, N2328);
buf BUF1 (N2553, N2549);
and AND4 (N2554, N2552, N644, N404, N606);
not NOT1 (N2555, N2554);
or OR4 (N2556, N2525, N922, N2187, N1545);
xor XOR2 (N2557, N2547, N746);
and AND3 (N2558, N2542, N1897, N358);
xor XOR2 (N2559, N2551, N1362);
nor NOR3 (N2560, N2553, N85, N1519);
xor XOR2 (N2561, N2560, N323);
buf BUF1 (N2562, N2535);
buf BUF1 (N2563, N2511);
nand NAND3 (N2564, N2550, N2070, N1949);
nor NOR3 (N2565, N2557, N2129, N819);
nor NOR2 (N2566, N2565, N1664);
xor XOR2 (N2567, N2563, N26);
or OR2 (N2568, N2555, N241);
nor NOR3 (N2569, N2567, N16, N924);
or OR4 (N2570, N2568, N1792, N1914, N1590);
nand NAND4 (N2571, N2562, N172, N1920, N254);
not NOT1 (N2572, N2566);
buf BUF1 (N2573, N2561);
nor NOR4 (N2574, N2570, N644, N465, N2284);
buf BUF1 (N2575, N2558);
xor XOR2 (N2576, N2573, N662);
xor XOR2 (N2577, N2527, N711);
xor XOR2 (N2578, N2577, N1383);
or OR4 (N2579, N2564, N838, N668, N2144);
nor NOR2 (N2580, N2572, N1889);
not NOT1 (N2581, N2575);
nor NOR2 (N2582, N2576, N2385);
nor NOR3 (N2583, N2574, N2030, N1985);
buf BUF1 (N2584, N2581);
xor XOR2 (N2585, N2584, N391);
or OR2 (N2586, N2571, N190);
nor NOR2 (N2587, N2559, N1072);
nand NAND4 (N2588, N2556, N2467, N1440, N1990);
or OR3 (N2589, N2585, N1772, N151);
and AND4 (N2590, N2586, N1243, N28, N1994);
and AND2 (N2591, N2579, N597);
nor NOR4 (N2592, N2569, N1898, N2129, N335);
or OR3 (N2593, N2578, N1816, N1544);
buf BUF1 (N2594, N2587);
buf BUF1 (N2595, N2582);
or OR2 (N2596, N2595, N1455);
nor NOR2 (N2597, N2593, N2067);
not NOT1 (N2598, N2596);
or OR3 (N2599, N2592, N333, N1502);
not NOT1 (N2600, N2583);
or OR4 (N2601, N2589, N1836, N1939, N467);
buf BUF1 (N2602, N2591);
xor XOR2 (N2603, N2599, N1324);
and AND3 (N2604, N2600, N2037, N1789);
and AND3 (N2605, N2590, N137, N424);
xor XOR2 (N2606, N2598, N2015);
xor XOR2 (N2607, N2601, N1599);
nand NAND3 (N2608, N2607, N1155, N124);
nand NAND4 (N2609, N2604, N303, N2537, N535);
and AND3 (N2610, N2597, N830, N2454);
xor XOR2 (N2611, N2610, N535);
and AND2 (N2612, N2608, N1796);
nor NOR4 (N2613, N2603, N952, N624, N610);
and AND4 (N2614, N2605, N812, N1888, N90);
buf BUF1 (N2615, N2580);
nor NOR4 (N2616, N2606, N1146, N1520, N342);
buf BUF1 (N2617, N2613);
not NOT1 (N2618, N2617);
buf BUF1 (N2619, N2618);
nand NAND2 (N2620, N2616, N1292);
not NOT1 (N2621, N2588);
not NOT1 (N2622, N2612);
nand NAND2 (N2623, N2594, N838);
nor NOR3 (N2624, N2622, N1178, N642);
buf BUF1 (N2625, N2611);
nand NAND4 (N2626, N2625, N1905, N684, N737);
or OR4 (N2627, N2609, N915, N2116, N1931);
xor XOR2 (N2628, N2624, N676);
not NOT1 (N2629, N2619);
xor XOR2 (N2630, N2614, N2509);
not NOT1 (N2631, N2623);
buf BUF1 (N2632, N2620);
xor XOR2 (N2633, N2621, N1828);
nor NOR3 (N2634, N2627, N92, N375);
nand NAND4 (N2635, N2615, N1077, N1356, N1033);
and AND3 (N2636, N2632, N625, N1732);
not NOT1 (N2637, N2635);
and AND3 (N2638, N2637, N576, N677);
nor NOR2 (N2639, N2630, N203);
nand NAND4 (N2640, N2628, N983, N1299, N60);
xor XOR2 (N2641, N2602, N482);
or OR3 (N2642, N2634, N673, N1448);
or OR3 (N2643, N2638, N1332, N644);
and AND2 (N2644, N2639, N2225);
or OR2 (N2645, N2629, N415);
or OR4 (N2646, N2643, N2088, N1998, N2054);
not NOT1 (N2647, N2636);
and AND2 (N2648, N2631, N767);
or OR2 (N2649, N2645, N674);
buf BUF1 (N2650, N2649);
nor NOR2 (N2651, N2633, N112);
nor NOR4 (N2652, N2644, N638, N1112, N2163);
nor NOR4 (N2653, N2626, N447, N1002, N971);
buf BUF1 (N2654, N2641);
buf BUF1 (N2655, N2646);
and AND3 (N2656, N2655, N1534, N2096);
buf BUF1 (N2657, N2652);
buf BUF1 (N2658, N2654);
nor NOR4 (N2659, N2657, N396, N2453, N1222);
nor NOR3 (N2660, N2658, N2429, N1210);
and AND2 (N2661, N2659, N1601);
xor XOR2 (N2662, N2647, N46);
nand NAND4 (N2663, N2648, N660, N1009, N1651);
buf BUF1 (N2664, N2663);
nand NAND3 (N2665, N2653, N1374, N2339);
not NOT1 (N2666, N2660);
or OR2 (N2667, N2651, N1568);
nand NAND4 (N2668, N2642, N686, N1488, N880);
xor XOR2 (N2669, N2665, N913);
and AND2 (N2670, N2667, N2054);
and AND2 (N2671, N2640, N2335);
nor NOR3 (N2672, N2664, N409, N595);
nand NAND4 (N2673, N2656, N289, N2284, N136);
nor NOR2 (N2674, N2668, N2627);
and AND2 (N2675, N2672, N1303);
nand NAND3 (N2676, N2674, N1837, N1279);
not NOT1 (N2677, N2650);
and AND3 (N2678, N2661, N2407, N2204);
nor NOR2 (N2679, N2677, N1302);
and AND4 (N2680, N2662, N133, N371, N390);
or OR2 (N2681, N2666, N1221);
buf BUF1 (N2682, N2681);
or OR2 (N2683, N2676, N208);
buf BUF1 (N2684, N2682);
not NOT1 (N2685, N2678);
not NOT1 (N2686, N2684);
nor NOR3 (N2687, N2671, N1905, N2633);
nor NOR2 (N2688, N2686, N605);
or OR3 (N2689, N2670, N2549, N1660);
or OR2 (N2690, N2689, N1781);
and AND2 (N2691, N2683, N2100);
xor XOR2 (N2692, N2691, N2081);
buf BUF1 (N2693, N2692);
not NOT1 (N2694, N2687);
xor XOR2 (N2695, N2690, N252);
or OR4 (N2696, N2675, N118, N1654, N354);
and AND3 (N2697, N2680, N2443, N905);
or OR3 (N2698, N2673, N706, N1721);
nor NOR3 (N2699, N2693, N2315, N429);
xor XOR2 (N2700, N2669, N1485);
and AND3 (N2701, N2688, N1427, N1203);
and AND4 (N2702, N2697, N1408, N490, N553);
buf BUF1 (N2703, N2698);
xor XOR2 (N2704, N2701, N1079);
and AND3 (N2705, N2703, N1935, N2219);
or OR3 (N2706, N2695, N2436, N2616);
nand NAND4 (N2707, N2679, N2615, N637, N1143);
and AND2 (N2708, N2685, N2413);
buf BUF1 (N2709, N2699);
and AND2 (N2710, N2694, N790);
nand NAND4 (N2711, N2700, N2035, N1990, N2031);
or OR4 (N2712, N2711, N2276, N1700, N1733);
nand NAND4 (N2713, N2705, N2219, N2406, N2435);
buf BUF1 (N2714, N2696);
or OR3 (N2715, N2713, N1523, N928);
buf BUF1 (N2716, N2706);
buf BUF1 (N2717, N2708);
nor NOR2 (N2718, N2702, N298);
nand NAND4 (N2719, N2704, N2224, N1733, N1864);
and AND4 (N2720, N2714, N1043, N2097, N1069);
or OR2 (N2721, N2710, N1300);
nand NAND2 (N2722, N2719, N1420);
buf BUF1 (N2723, N2715);
buf BUF1 (N2724, N2723);
nand NAND4 (N2725, N2718, N2389, N2150, N787);
nand NAND4 (N2726, N2716, N2361, N2447, N2335);
not NOT1 (N2727, N2722);
and AND3 (N2728, N2727, N40, N190);
buf BUF1 (N2729, N2726);
not NOT1 (N2730, N2729);
nand NAND3 (N2731, N2717, N1180, N467);
not NOT1 (N2732, N2730);
xor XOR2 (N2733, N2728, N2610);
xor XOR2 (N2734, N2721, N1491);
nor NOR4 (N2735, N2712, N1339, N2238, N835);
nand NAND3 (N2736, N2720, N1519, N2109);
or OR3 (N2737, N2734, N106, N2524);
xor XOR2 (N2738, N2733, N1238);
or OR4 (N2739, N2709, N1115, N1461, N1673);
or OR2 (N2740, N2732, N1641);
buf BUF1 (N2741, N2736);
xor XOR2 (N2742, N2724, N2458);
nand NAND2 (N2743, N2740, N2693);
or OR4 (N2744, N2743, N2634, N825, N567);
nor NOR4 (N2745, N2725, N2049, N323, N678);
xor XOR2 (N2746, N2731, N893);
buf BUF1 (N2747, N2744);
or OR3 (N2748, N2742, N314, N1318);
nand NAND3 (N2749, N2748, N973, N1512);
nor NOR2 (N2750, N2735, N2380);
not NOT1 (N2751, N2739);
buf BUF1 (N2752, N2745);
xor XOR2 (N2753, N2707, N1389);
nor NOR3 (N2754, N2746, N39, N248);
not NOT1 (N2755, N2753);
or OR2 (N2756, N2755, N2598);
buf BUF1 (N2757, N2751);
or OR3 (N2758, N2752, N161, N1002);
not NOT1 (N2759, N2747);
nor NOR4 (N2760, N2757, N470, N1422, N63);
not NOT1 (N2761, N2756);
not NOT1 (N2762, N2761);
not NOT1 (N2763, N2760);
or OR3 (N2764, N2758, N632, N1322);
nand NAND2 (N2765, N2763, N2462);
or OR3 (N2766, N2737, N2079, N2692);
nand NAND3 (N2767, N2749, N2731, N1911);
nand NAND3 (N2768, N2762, N404, N2265);
xor XOR2 (N2769, N2750, N918);
or OR2 (N2770, N2767, N269);
xor XOR2 (N2771, N2768, N1442);
nor NOR2 (N2772, N2765, N1615);
nor NOR2 (N2773, N2770, N2346);
nor NOR4 (N2774, N2759, N834, N1166, N1926);
and AND2 (N2775, N2774, N528);
nor NOR2 (N2776, N2772, N438);
xor XOR2 (N2777, N2766, N392);
nand NAND3 (N2778, N2741, N1577, N173);
buf BUF1 (N2779, N2778);
or OR2 (N2780, N2769, N1122);
nand NAND4 (N2781, N2771, N2169, N304, N10);
nor NOR3 (N2782, N2777, N1434, N1487);
or OR4 (N2783, N2780, N2339, N811, N1949);
buf BUF1 (N2784, N2775);
nand NAND3 (N2785, N2754, N2778, N1045);
and AND2 (N2786, N2738, N402);
and AND2 (N2787, N2781, N1472);
not NOT1 (N2788, N2779);
nor NOR2 (N2789, N2782, N2775);
buf BUF1 (N2790, N2773);
or OR3 (N2791, N2784, N2630, N526);
and AND3 (N2792, N2788, N2702, N164);
not NOT1 (N2793, N2776);
or OR3 (N2794, N2764, N763, N167);
xor XOR2 (N2795, N2790, N2396);
and AND4 (N2796, N2789, N930, N250, N2598);
or OR3 (N2797, N2796, N2538, N122);
not NOT1 (N2798, N2794);
xor XOR2 (N2799, N2793, N1667);
nand NAND3 (N2800, N2785, N791, N472);
and AND4 (N2801, N2786, N1248, N1920, N1460);
nor NOR4 (N2802, N2795, N2486, N1887, N196);
and AND2 (N2803, N2799, N1978);
xor XOR2 (N2804, N2797, N1653);
or OR2 (N2805, N2798, N407);
buf BUF1 (N2806, N2802);
or OR2 (N2807, N2792, N2756);
nor NOR3 (N2808, N2787, N543, N809);
nor NOR4 (N2809, N2807, N2441, N2700, N979);
nand NAND4 (N2810, N2808, N2455, N837, N876);
and AND4 (N2811, N2806, N1367, N2229, N2622);
buf BUF1 (N2812, N2810);
and AND3 (N2813, N2783, N923, N884);
and AND2 (N2814, N2813, N1648);
xor XOR2 (N2815, N2800, N2308);
nand NAND2 (N2816, N2803, N1099);
or OR3 (N2817, N2815, N1243, N1098);
not NOT1 (N2818, N2805);
nand NAND2 (N2819, N2811, N1697);
nor NOR4 (N2820, N2814, N875, N1877, N2444);
nand NAND2 (N2821, N2812, N1252);
not NOT1 (N2822, N2820);
or OR2 (N2823, N2801, N2765);
nor NOR3 (N2824, N2823, N840, N90);
buf BUF1 (N2825, N2819);
and AND2 (N2826, N2821, N174);
and AND3 (N2827, N2818, N654, N876);
not NOT1 (N2828, N2824);
nor NOR4 (N2829, N2822, N1320, N2061, N1542);
not NOT1 (N2830, N2809);
buf BUF1 (N2831, N2825);
xor XOR2 (N2832, N2828, N1060);
xor XOR2 (N2833, N2829, N80);
or OR2 (N2834, N2827, N1177);
buf BUF1 (N2835, N2832);
and AND3 (N2836, N2816, N2251, N1183);
xor XOR2 (N2837, N2817, N808);
or OR3 (N2838, N2834, N462, N1463);
nor NOR4 (N2839, N2804, N997, N2112, N2060);
or OR3 (N2840, N2826, N1787, N2799);
not NOT1 (N2841, N2833);
not NOT1 (N2842, N2839);
nor NOR4 (N2843, N2842, N1055, N2500, N1295);
nor NOR3 (N2844, N2843, N536, N2628);
xor XOR2 (N2845, N2791, N328);
nand NAND4 (N2846, N2840, N837, N1832, N1799);
nand NAND4 (N2847, N2841, N51, N2765, N1158);
nor NOR2 (N2848, N2847, N18);
not NOT1 (N2849, N2831);
buf BUF1 (N2850, N2837);
nand NAND2 (N2851, N2838, N2590);
nor NOR4 (N2852, N2830, N1127, N2463, N1343);
not NOT1 (N2853, N2835);
buf BUF1 (N2854, N2848);
nand NAND3 (N2855, N2852, N2186, N1724);
nand NAND4 (N2856, N2855, N527, N911, N1058);
buf BUF1 (N2857, N2851);
buf BUF1 (N2858, N2849);
and AND2 (N2859, N2857, N594);
or OR3 (N2860, N2854, N1805, N2366);
xor XOR2 (N2861, N2853, N2313);
buf BUF1 (N2862, N2846);
buf BUF1 (N2863, N2845);
buf BUF1 (N2864, N2860);
xor XOR2 (N2865, N2858, N420);
or OR3 (N2866, N2859, N1362, N1862);
nor NOR2 (N2867, N2862, N893);
xor XOR2 (N2868, N2836, N1982);
buf BUF1 (N2869, N2868);
buf BUF1 (N2870, N2856);
xor XOR2 (N2871, N2850, N2313);
and AND4 (N2872, N2844, N1080, N2647, N1595);
nand NAND2 (N2873, N2864, N828);
nor NOR4 (N2874, N2866, N299, N1664, N833);
nand NAND3 (N2875, N2861, N541, N1093);
nor NOR3 (N2876, N2872, N19, N1326);
nor NOR2 (N2877, N2870, N489);
and AND4 (N2878, N2865, N2078, N2352, N161);
or OR2 (N2879, N2874, N1697);
and AND2 (N2880, N2863, N2839);
and AND4 (N2881, N2871, N2392, N497, N993);
xor XOR2 (N2882, N2869, N375);
buf BUF1 (N2883, N2881);
and AND3 (N2884, N2882, N1956, N2203);
or OR2 (N2885, N2867, N1856);
nand NAND4 (N2886, N2878, N1407, N2884, N2567);
nand NAND3 (N2887, N375, N38, N876);
nand NAND2 (N2888, N2873, N2273);
nand NAND4 (N2889, N2879, N1816, N1063, N2791);
not NOT1 (N2890, N2887);
nor NOR2 (N2891, N2875, N1452);
not NOT1 (N2892, N2876);
and AND4 (N2893, N2890, N2489, N353, N1725);
buf BUF1 (N2894, N2888);
nor NOR4 (N2895, N2893, N337, N1717, N1095);
not NOT1 (N2896, N2894);
nand NAND3 (N2897, N2880, N1597, N1448);
nand NAND2 (N2898, N2889, N1895);
nor NOR4 (N2899, N2898, N257, N595, N1174);
nor NOR4 (N2900, N2883, N1619, N1129, N1607);
not NOT1 (N2901, N2900);
xor XOR2 (N2902, N2895, N1578);
and AND2 (N2903, N2891, N907);
xor XOR2 (N2904, N2886, N733);
not NOT1 (N2905, N2902);
or OR4 (N2906, N2892, N2438, N1976, N2637);
and AND2 (N2907, N2885, N670);
buf BUF1 (N2908, N2899);
xor XOR2 (N2909, N2897, N2455);
not NOT1 (N2910, N2896);
nand NAND3 (N2911, N2901, N573, N824);
nor NOR4 (N2912, N2903, N466, N538, N280);
not NOT1 (N2913, N2904);
and AND2 (N2914, N2910, N2014);
buf BUF1 (N2915, N2911);
nand NAND4 (N2916, N2877, N413, N809, N2833);
or OR3 (N2917, N2907, N1369, N989);
and AND3 (N2918, N2913, N2511, N1958);
not NOT1 (N2919, N2915);
nand NAND2 (N2920, N2905, N73);
nand NAND3 (N2921, N2908, N1918, N315);
xor XOR2 (N2922, N2909, N1170);
nand NAND3 (N2923, N2918, N505, N1504);
nor NOR3 (N2924, N2921, N1389, N1834);
and AND2 (N2925, N2923, N2562);
or OR2 (N2926, N2912, N2010);
or OR3 (N2927, N2906, N907, N1823);
not NOT1 (N2928, N2917);
buf BUF1 (N2929, N2924);
not NOT1 (N2930, N2920);
not NOT1 (N2931, N2929);
or OR3 (N2932, N2916, N210, N2410);
or OR3 (N2933, N2919, N213, N2931);
or OR2 (N2934, N1688, N865);
not NOT1 (N2935, N2933);
buf BUF1 (N2936, N2927);
or OR3 (N2937, N2935, N1190, N2406);
nand NAND4 (N2938, N2925, N1110, N1710, N29);
nor NOR2 (N2939, N2930, N1811);
or OR4 (N2940, N2937, N2804, N1143, N1784);
or OR3 (N2941, N2938, N2535, N1473);
and AND2 (N2942, N2941, N2936);
nand NAND3 (N2943, N1847, N2888, N376);
buf BUF1 (N2944, N2922);
nand NAND2 (N2945, N2940, N916);
not NOT1 (N2946, N2928);
nor NOR4 (N2947, N2932, N450, N194, N313);
not NOT1 (N2948, N2939);
or OR4 (N2949, N2926, N461, N217, N229);
nor NOR3 (N2950, N2946, N1727, N335);
nor NOR2 (N2951, N2943, N2391);
buf BUF1 (N2952, N2944);
or OR4 (N2953, N2945, N255, N1942, N645);
xor XOR2 (N2954, N2952, N735);
xor XOR2 (N2955, N2954, N768);
nor NOR3 (N2956, N2934, N2809, N2071);
or OR4 (N2957, N2951, N2561, N1759, N2102);
buf BUF1 (N2958, N2948);
nand NAND3 (N2959, N2942, N2287, N1405);
nand NAND3 (N2960, N2958, N2694, N2821);
nor NOR3 (N2961, N2957, N732, N1700);
buf BUF1 (N2962, N2949);
not NOT1 (N2963, N2961);
buf BUF1 (N2964, N2960);
buf BUF1 (N2965, N2947);
xor XOR2 (N2966, N2956, N526);
nand NAND3 (N2967, N2965, N509, N792);
xor XOR2 (N2968, N2962, N1114);
xor XOR2 (N2969, N2967, N2226);
nand NAND2 (N2970, N2964, N2474);
buf BUF1 (N2971, N2968);
and AND3 (N2972, N2914, N1611, N1482);
xor XOR2 (N2973, N2963, N2597);
nor NOR3 (N2974, N2972, N1549, N1685);
or OR3 (N2975, N2953, N1456, N475);
not NOT1 (N2976, N2966);
buf BUF1 (N2977, N2975);
buf BUF1 (N2978, N2970);
nor NOR2 (N2979, N2977, N804);
and AND3 (N2980, N2979, N229, N623);
nor NOR4 (N2981, N2976, N2610, N891, N1722);
nor NOR4 (N2982, N2980, N34, N871, N2202);
not NOT1 (N2983, N2978);
not NOT1 (N2984, N2971);
or OR4 (N2985, N2984, N607, N1954, N713);
nand NAND3 (N2986, N2969, N2010, N1808);
or OR3 (N2987, N2985, N2595, N221);
and AND3 (N2988, N2973, N2268, N1784);
buf BUF1 (N2989, N2959);
and AND3 (N2990, N2988, N627, N2012);
xor XOR2 (N2991, N2987, N93);
xor XOR2 (N2992, N2990, N289);
xor XOR2 (N2993, N2981, N2877);
xor XOR2 (N2994, N2993, N2253);
nor NOR2 (N2995, N2989, N1231);
not NOT1 (N2996, N2986);
not NOT1 (N2997, N2994);
nand NAND3 (N2998, N2982, N856, N1321);
xor XOR2 (N2999, N2997, N267);
or OR4 (N3000, N2998, N364, N2291, N130);
not NOT1 (N3001, N2992);
xor XOR2 (N3002, N3000, N1);
and AND2 (N3003, N3001, N2529);
and AND3 (N3004, N2955, N2150, N2499);
nor NOR3 (N3005, N2950, N517, N1159);
or OR2 (N3006, N2995, N2506);
xor XOR2 (N3007, N2991, N327);
or OR3 (N3008, N2996, N341, N509);
nand NAND4 (N3009, N3005, N159, N597, N2126);
buf BUF1 (N3010, N3006);
nor NOR4 (N3011, N3002, N1627, N684, N2915);
nand NAND4 (N3012, N2974, N2569, N1634, N517);
or OR2 (N3013, N2999, N2815);
or OR4 (N3014, N2983, N2221, N1517, N11);
nand NAND2 (N3015, N3012, N1317);
or OR4 (N3016, N3004, N2018, N91, N1150);
buf BUF1 (N3017, N3008);
nand NAND2 (N3018, N3016, N1870);
buf BUF1 (N3019, N3018);
or OR4 (N3020, N3015, N414, N333, N31);
nand NAND3 (N3021, N3020, N1209, N398);
buf BUF1 (N3022, N3009);
buf BUF1 (N3023, N3014);
and AND3 (N3024, N3013, N1810, N398);
nor NOR3 (N3025, N3024, N2578, N508);
nor NOR3 (N3026, N3017, N852, N2813);
nand NAND2 (N3027, N3025, N313);
nor NOR2 (N3028, N3011, N2948);
buf BUF1 (N3029, N3003);
buf BUF1 (N3030, N3021);
nor NOR4 (N3031, N3026, N884, N465, N2965);
not NOT1 (N3032, N3028);
nor NOR2 (N3033, N3007, N2353);
xor XOR2 (N3034, N3031, N1621);
not NOT1 (N3035, N3033);
or OR4 (N3036, N3027, N977, N819, N2983);
nand NAND2 (N3037, N3036, N204);
or OR4 (N3038, N3022, N2838, N2131, N2340);
or OR3 (N3039, N3037, N2562, N54);
xor XOR2 (N3040, N3034, N2430);
xor XOR2 (N3041, N3010, N2818);
not NOT1 (N3042, N3023);
and AND2 (N3043, N3041, N1257);
not NOT1 (N3044, N3032);
not NOT1 (N3045, N3043);
xor XOR2 (N3046, N3044, N568);
or OR3 (N3047, N3019, N699, N131);
or OR3 (N3048, N3039, N805, N1823);
nor NOR3 (N3049, N3029, N1609, N1959);
not NOT1 (N3050, N3045);
nand NAND3 (N3051, N3048, N1711, N2486);
buf BUF1 (N3052, N3051);
and AND2 (N3053, N3046, N532);
xor XOR2 (N3054, N3052, N1278);
xor XOR2 (N3055, N3038, N836);
nor NOR2 (N3056, N3047, N1917);
and AND2 (N3057, N3040, N2879);
and AND2 (N3058, N3030, N905);
and AND3 (N3059, N3056, N779, N485);
and AND4 (N3060, N3055, N1313, N2899, N2340);
xor XOR2 (N3061, N3042, N2504);
and AND3 (N3062, N3053, N96, N1437);
or OR3 (N3063, N3054, N445, N469);
or OR4 (N3064, N3049, N2994, N1044, N1078);
or OR4 (N3065, N3063, N2350, N871, N1993);
xor XOR2 (N3066, N3057, N1092);
nor NOR4 (N3067, N3065, N182, N1008, N747);
or OR3 (N3068, N3060, N2081, N2956);
and AND2 (N3069, N3062, N963);
and AND3 (N3070, N3069, N1192, N1807);
buf BUF1 (N3071, N3061);
xor XOR2 (N3072, N3071, N2742);
xor XOR2 (N3073, N3058, N758);
buf BUF1 (N3074, N3059);
nand NAND3 (N3075, N3064, N1212, N2323);
and AND3 (N3076, N3066, N504, N687);
xor XOR2 (N3077, N3067, N2800);
nor NOR3 (N3078, N3050, N566, N35);
xor XOR2 (N3079, N3074, N2686);
not NOT1 (N3080, N3076);
and AND3 (N3081, N3078, N502, N2142);
not NOT1 (N3082, N3035);
and AND2 (N3083, N3073, N705);
not NOT1 (N3084, N3072);
nand NAND2 (N3085, N3079, N2500);
or OR2 (N3086, N3084, N3021);
not NOT1 (N3087, N3075);
not NOT1 (N3088, N3081);
nand NAND4 (N3089, N3088, N2210, N741, N867);
xor XOR2 (N3090, N3087, N1033);
xor XOR2 (N3091, N3083, N1501);
nor NOR2 (N3092, N3086, N2232);
nand NAND2 (N3093, N3085, N2322);
nand NAND3 (N3094, N3080, N603, N313);
xor XOR2 (N3095, N3082, N2976);
buf BUF1 (N3096, N3092);
buf BUF1 (N3097, N3095);
nor NOR4 (N3098, N3093, N510, N1254, N2624);
or OR3 (N3099, N3090, N112, N1648);
or OR4 (N3100, N3097, N2504, N221, N283);
and AND4 (N3101, N3100, N1690, N1048, N2389);
and AND3 (N3102, N3077, N2597, N657);
nor NOR3 (N3103, N3096, N1662, N2263);
nor NOR4 (N3104, N3070, N1105, N1909, N2023);
xor XOR2 (N3105, N3094, N541);
xor XOR2 (N3106, N3101, N2836);
buf BUF1 (N3107, N3091);
nand NAND4 (N3108, N3102, N1120, N1484, N2983);
xor XOR2 (N3109, N3106, N197);
and AND4 (N3110, N3098, N2374, N647, N405);
or OR2 (N3111, N3089, N2770);
buf BUF1 (N3112, N3099);
nor NOR2 (N3113, N3105, N2645);
nand NAND3 (N3114, N3109, N511, N99);
not NOT1 (N3115, N3111);
not NOT1 (N3116, N3114);
nor NOR2 (N3117, N3115, N1045);
xor XOR2 (N3118, N3116, N1065);
xor XOR2 (N3119, N3108, N1635);
and AND4 (N3120, N3117, N2170, N449, N2707);
or OR2 (N3121, N3107, N3095);
or OR4 (N3122, N3068, N1236, N894, N969);
not NOT1 (N3123, N3112);
xor XOR2 (N3124, N3103, N2198);
nand NAND3 (N3125, N3118, N2387, N303);
nor NOR2 (N3126, N3113, N2687);
not NOT1 (N3127, N3104);
not NOT1 (N3128, N3123);
not NOT1 (N3129, N3126);
and AND2 (N3130, N3125, N1179);
nand NAND2 (N3131, N3130, N1888);
nor NOR2 (N3132, N3119, N1912);
and AND2 (N3133, N3120, N1397);
or OR2 (N3134, N3128, N459);
buf BUF1 (N3135, N3121);
xor XOR2 (N3136, N3131, N469);
not NOT1 (N3137, N3122);
and AND2 (N3138, N3132, N2375);
and AND3 (N3139, N3138, N1439, N1024);
or OR4 (N3140, N3136, N211, N1951, N1597);
buf BUF1 (N3141, N3135);
or OR4 (N3142, N3137, N1348, N2042, N707);
nor NOR4 (N3143, N3124, N2633, N356, N2369);
xor XOR2 (N3144, N3110, N2839);
xor XOR2 (N3145, N3134, N2580);
or OR2 (N3146, N3133, N1235);
nor NOR3 (N3147, N3129, N1070, N374);
nor NOR4 (N3148, N3139, N1154, N3079, N1989);
nor NOR3 (N3149, N3143, N401, N2345);
nor NOR3 (N3150, N3145, N1319, N2037);
not NOT1 (N3151, N3140);
and AND4 (N3152, N3127, N2165, N2410, N785);
xor XOR2 (N3153, N3148, N1958);
nor NOR4 (N3154, N3146, N771, N837, N279);
buf BUF1 (N3155, N3150);
or OR3 (N3156, N3144, N1771, N249);
and AND4 (N3157, N3151, N1770, N1140, N726);
nor NOR3 (N3158, N3157, N476, N1073);
buf BUF1 (N3159, N3142);
xor XOR2 (N3160, N3154, N2066);
xor XOR2 (N3161, N3156, N2649);
nand NAND3 (N3162, N3153, N1584, N2641);
or OR4 (N3163, N3161, N2573, N1111, N1021);
or OR2 (N3164, N3147, N974);
or OR2 (N3165, N3163, N578);
nand NAND4 (N3166, N3152, N774, N2352, N2464);
not NOT1 (N3167, N3141);
xor XOR2 (N3168, N3159, N1314);
and AND2 (N3169, N3166, N340);
nor NOR4 (N3170, N3169, N192, N2317, N2992);
and AND3 (N3171, N3149, N1656, N733);
and AND3 (N3172, N3167, N1015, N2754);
nor NOR2 (N3173, N3160, N3126);
xor XOR2 (N3174, N3165, N767);
xor XOR2 (N3175, N3170, N799);
buf BUF1 (N3176, N3175);
nor NOR4 (N3177, N3162, N1141, N2199, N2945);
nor NOR4 (N3178, N3155, N602, N731, N2301);
and AND3 (N3179, N3176, N1887, N2338);
buf BUF1 (N3180, N3164);
not NOT1 (N3181, N3168);
not NOT1 (N3182, N3181);
buf BUF1 (N3183, N3174);
nor NOR4 (N3184, N3183, N1633, N684, N3090);
nor NOR4 (N3185, N3173, N1337, N1754, N610);
not NOT1 (N3186, N3180);
not NOT1 (N3187, N3185);
xor XOR2 (N3188, N3158, N916);
or OR2 (N3189, N3178, N2690);
buf BUF1 (N3190, N3171);
nand NAND4 (N3191, N3182, N441, N2946, N1924);
and AND4 (N3192, N3172, N1540, N1403, N1091);
nor NOR4 (N3193, N3189, N1374, N1693, N763);
not NOT1 (N3194, N3179);
not NOT1 (N3195, N3192);
nor NOR3 (N3196, N3186, N2334, N1547);
xor XOR2 (N3197, N3194, N1678);
and AND4 (N3198, N3197, N182, N1132, N3063);
and AND2 (N3199, N3187, N1149);
and AND2 (N3200, N3184, N2039);
not NOT1 (N3201, N3196);
nor NOR3 (N3202, N3201, N863, N2978);
not NOT1 (N3203, N3198);
buf BUF1 (N3204, N3195);
nor NOR2 (N3205, N3199, N2903);
nand NAND2 (N3206, N3205, N1043);
or OR3 (N3207, N3202, N1843, N1455);
xor XOR2 (N3208, N3190, N2818);
buf BUF1 (N3209, N3191);
not NOT1 (N3210, N3188);
or OR4 (N3211, N3204, N1119, N2218, N593);
not NOT1 (N3212, N3200);
buf BUF1 (N3213, N3208);
buf BUF1 (N3214, N3177);
and AND4 (N3215, N3213, N2378, N1872, N329);
and AND4 (N3216, N3210, N1719, N3001, N456);
buf BUF1 (N3217, N3216);
buf BUF1 (N3218, N3193);
or OR4 (N3219, N3211, N1534, N1098, N1380);
and AND2 (N3220, N3215, N566);
buf BUF1 (N3221, N3219);
and AND3 (N3222, N3207, N1176, N2167);
and AND4 (N3223, N3212, N110, N988, N2200);
nand NAND2 (N3224, N3217, N398);
buf BUF1 (N3225, N3218);
or OR3 (N3226, N3221, N2624, N1894);
buf BUF1 (N3227, N3220);
not NOT1 (N3228, N3214);
and AND4 (N3229, N3226, N2669, N653, N448);
buf BUF1 (N3230, N3227);
and AND3 (N3231, N3228, N3134, N757);
not NOT1 (N3232, N3229);
nand NAND4 (N3233, N3203, N1337, N814, N2434);
or OR4 (N3234, N3206, N2756, N2218, N1449);
and AND2 (N3235, N3230, N1869);
or OR2 (N3236, N3224, N1755);
or OR4 (N3237, N3235, N2724, N2081, N828);
and AND2 (N3238, N3234, N2321);
nand NAND2 (N3239, N3237, N76);
nand NAND2 (N3240, N3231, N1861);
nor NOR4 (N3241, N3240, N920, N311, N3192);
nand NAND3 (N3242, N3236, N398, N1393);
or OR3 (N3243, N3232, N2210, N2159);
buf BUF1 (N3244, N3242);
nand NAND2 (N3245, N3239, N1743);
not NOT1 (N3246, N3241);
or OR2 (N3247, N3246, N741);
buf BUF1 (N3248, N3225);
buf BUF1 (N3249, N3247);
xor XOR2 (N3250, N3209, N1468);
not NOT1 (N3251, N3249);
nand NAND4 (N3252, N3233, N313, N325, N1456);
nand NAND3 (N3253, N3248, N1384, N390);
nor NOR4 (N3254, N3222, N2210, N1802, N1144);
xor XOR2 (N3255, N3245, N1126);
xor XOR2 (N3256, N3244, N294);
nand NAND2 (N3257, N3252, N668);
buf BUF1 (N3258, N3253);
nand NAND3 (N3259, N3258, N2595, N662);
and AND2 (N3260, N3257, N1120);
and AND4 (N3261, N3238, N2552, N1361, N1520);
nand NAND2 (N3262, N3223, N3144);
and AND3 (N3263, N3255, N3098, N428);
nand NAND3 (N3264, N3250, N2032, N2729);
or OR4 (N3265, N3260, N3221, N2855, N3121);
and AND4 (N3266, N3261, N57, N65, N1949);
nor NOR3 (N3267, N3262, N1018, N2417);
not NOT1 (N3268, N3243);
buf BUF1 (N3269, N3267);
buf BUF1 (N3270, N3265);
or OR3 (N3271, N3264, N717, N2061);
or OR2 (N3272, N3263, N1255);
and AND2 (N3273, N3256, N302);
nand NAND3 (N3274, N3266, N2825, N2850);
and AND4 (N3275, N3271, N1248, N2994, N180);
xor XOR2 (N3276, N3270, N3132);
or OR3 (N3277, N3268, N269, N2055);
not NOT1 (N3278, N3277);
and AND2 (N3279, N3276, N382);
or OR4 (N3280, N3272, N2017, N20, N1891);
nor NOR2 (N3281, N3259, N360);
nor NOR3 (N3282, N3279, N1011, N598);
or OR2 (N3283, N3278, N2556);
or OR3 (N3284, N3269, N1325, N228);
nand NAND3 (N3285, N3282, N532, N2065);
nor NOR2 (N3286, N3281, N834);
buf BUF1 (N3287, N3273);
xor XOR2 (N3288, N3251, N287);
nor NOR4 (N3289, N3280, N2501, N906, N2060);
nand NAND4 (N3290, N3289, N176, N1925, N344);
buf BUF1 (N3291, N3287);
not NOT1 (N3292, N3254);
nand NAND4 (N3293, N3288, N972, N1004, N2709);
not NOT1 (N3294, N3274);
and AND3 (N3295, N3293, N701, N3002);
not NOT1 (N3296, N3294);
nor NOR2 (N3297, N3286, N443);
nor NOR3 (N3298, N3297, N1336, N509);
nand NAND4 (N3299, N3292, N1054, N692, N2970);
nand NAND2 (N3300, N3290, N2336);
or OR3 (N3301, N3296, N399, N1824);
nor NOR3 (N3302, N3285, N1691, N2504);
xor XOR2 (N3303, N3300, N1919);
or OR2 (N3304, N3301, N1853);
nand NAND3 (N3305, N3302, N3105, N9);
not NOT1 (N3306, N3303);
or OR3 (N3307, N3291, N1458, N2522);
nand NAND3 (N3308, N3299, N2125, N3265);
or OR3 (N3309, N3295, N1667, N3224);
nand NAND3 (N3310, N3308, N550, N572);
nand NAND4 (N3311, N3307, N3305, N2483, N797);
buf BUF1 (N3312, N918);
nor NOR2 (N3313, N3284, N3060);
buf BUF1 (N3314, N3283);
nand NAND4 (N3315, N3309, N1461, N2310, N420);
not NOT1 (N3316, N3312);
not NOT1 (N3317, N3275);
and AND4 (N3318, N3317, N1223, N1850, N2465);
nor NOR4 (N3319, N3313, N1713, N409, N1959);
buf BUF1 (N3320, N3298);
nand NAND2 (N3321, N3315, N1326);
and AND4 (N3322, N3310, N237, N3293, N2342);
nor NOR3 (N3323, N3319, N2375, N2908);
nor NOR3 (N3324, N3318, N1594, N2718);
buf BUF1 (N3325, N3322);
buf BUF1 (N3326, N3323);
nand NAND3 (N3327, N3306, N2904, N2853);
nand NAND4 (N3328, N3314, N2071, N2957, N988);
buf BUF1 (N3329, N3316);
nand NAND3 (N3330, N3321, N1911, N3207);
nor NOR2 (N3331, N3325, N1924);
or OR4 (N3332, N3311, N2864, N337, N2846);
nor NOR2 (N3333, N3326, N301);
nor NOR2 (N3334, N3331, N234);
buf BUF1 (N3335, N3320);
or OR3 (N3336, N3330, N1443, N2277);
xor XOR2 (N3337, N3335, N2733);
and AND3 (N3338, N3304, N608, N546);
nand NAND3 (N3339, N3327, N2999, N518);
nor NOR2 (N3340, N3324, N938);
or OR4 (N3341, N3333, N450, N1764, N1215);
nand NAND2 (N3342, N3338, N54);
xor XOR2 (N3343, N3341, N3158);
and AND4 (N3344, N3328, N433, N1074, N2160);
or OR4 (N3345, N3329, N94, N2375, N1271);
or OR3 (N3346, N3345, N1440, N1890);
not NOT1 (N3347, N3332);
or OR2 (N3348, N3344, N1469);
and AND3 (N3349, N3346, N143, N478);
nor NOR2 (N3350, N3349, N1267);
buf BUF1 (N3351, N3348);
nand NAND4 (N3352, N3347, N920, N2445, N2507);
xor XOR2 (N3353, N3352, N140);
and AND3 (N3354, N3334, N376, N2774);
nand NAND2 (N3355, N3350, N372);
buf BUF1 (N3356, N3343);
nand NAND2 (N3357, N3354, N1925);
nor NOR3 (N3358, N3356, N2164, N2254);
not NOT1 (N3359, N3336);
nand NAND3 (N3360, N3337, N1819, N188);
not NOT1 (N3361, N3358);
not NOT1 (N3362, N3359);
nor NOR3 (N3363, N3351, N925, N339);
or OR4 (N3364, N3363, N3107, N2735, N2266);
and AND4 (N3365, N3361, N3024, N651, N1849);
and AND3 (N3366, N3342, N561, N1294);
buf BUF1 (N3367, N3360);
and AND3 (N3368, N3357, N1783, N1638);
xor XOR2 (N3369, N3340, N3044);
nand NAND4 (N3370, N3367, N451, N2785, N3066);
xor XOR2 (N3371, N3368, N1146);
nor NOR4 (N3372, N3366, N867, N2271, N1525);
nor NOR3 (N3373, N3355, N2623, N1307);
not NOT1 (N3374, N3370);
nand NAND2 (N3375, N3374, N1126);
or OR3 (N3376, N3369, N2388, N2672);
or OR3 (N3377, N3371, N175, N2664);
nor NOR3 (N3378, N3364, N2770, N1559);
not NOT1 (N3379, N3373);
and AND4 (N3380, N3378, N244, N2044, N1906);
nand NAND4 (N3381, N3375, N918, N2938, N2201);
or OR4 (N3382, N3372, N1685, N2210, N2059);
or OR2 (N3383, N3379, N148);
nand NAND2 (N3384, N3383, N28);
or OR4 (N3385, N3353, N929, N1590, N70);
nand NAND3 (N3386, N3385, N1499, N2013);
nor NOR2 (N3387, N3381, N1780);
and AND4 (N3388, N3339, N2900, N1406, N1034);
or OR2 (N3389, N3388, N3053);
not NOT1 (N3390, N3384);
nor NOR2 (N3391, N3380, N3302);
or OR2 (N3392, N3377, N2805);
or OR3 (N3393, N3392, N1538, N947);
or OR2 (N3394, N3389, N2787);
nor NOR3 (N3395, N3390, N29, N1785);
or OR3 (N3396, N3365, N3061, N451);
or OR2 (N3397, N3382, N858);
nor NOR4 (N3398, N3376, N324, N154, N1365);
or OR2 (N3399, N3386, N2093);
nand NAND4 (N3400, N3399, N3291, N3, N2824);
nand NAND2 (N3401, N3397, N516);
and AND3 (N3402, N3394, N3339, N1282);
nand NAND3 (N3403, N3398, N2419, N3282);
nor NOR3 (N3404, N3362, N3003, N3243);
buf BUF1 (N3405, N3402);
xor XOR2 (N3406, N3387, N3370);
nor NOR3 (N3407, N3395, N1655, N2803);
buf BUF1 (N3408, N3405);
nor NOR2 (N3409, N3406, N2375);
xor XOR2 (N3410, N3407, N2313);
buf BUF1 (N3411, N3396);
buf BUF1 (N3412, N3403);
or OR3 (N3413, N3393, N336, N1981);
nor NOR2 (N3414, N3409, N2466);
nor NOR2 (N3415, N3411, N1044);
buf BUF1 (N3416, N3410);
and AND3 (N3417, N3404, N100, N1811);
buf BUF1 (N3418, N3400);
or OR4 (N3419, N3408, N2830, N2555, N753);
nand NAND3 (N3420, N3418, N1560, N2315);
xor XOR2 (N3421, N3391, N1800);
not NOT1 (N3422, N3414);
and AND3 (N3423, N3412, N2469, N921);
nor NOR3 (N3424, N3417, N1718, N2366);
not NOT1 (N3425, N3420);
and AND4 (N3426, N3425, N770, N188, N895);
and AND4 (N3427, N3413, N3290, N3237, N1070);
xor XOR2 (N3428, N3421, N1826);
nand NAND3 (N3429, N3428, N120, N1350);
not NOT1 (N3430, N3416);
xor XOR2 (N3431, N3424, N2778);
not NOT1 (N3432, N3429);
or OR3 (N3433, N3432, N1271, N1294);
nor NOR4 (N3434, N3431, N139, N13, N202);
nor NOR2 (N3435, N3433, N1995);
buf BUF1 (N3436, N3435);
buf BUF1 (N3437, N3430);
not NOT1 (N3438, N3434);
xor XOR2 (N3439, N3401, N1445);
nor NOR4 (N3440, N3436, N1256, N1993, N1090);
buf BUF1 (N3441, N3437);
or OR2 (N3442, N3426, N1171);
not NOT1 (N3443, N3423);
xor XOR2 (N3444, N3439, N3421);
nand NAND2 (N3445, N3422, N14);
not NOT1 (N3446, N3438);
not NOT1 (N3447, N3440);
buf BUF1 (N3448, N3442);
nand NAND4 (N3449, N3427, N1458, N3180, N2512);
or OR3 (N3450, N3419, N869, N1936);
nor NOR4 (N3451, N3444, N2418, N3388, N1231);
not NOT1 (N3452, N3441);
xor XOR2 (N3453, N3448, N1453);
xor XOR2 (N3454, N3415, N1918);
or OR4 (N3455, N3453, N3255, N1084, N2795);
or OR3 (N3456, N3454, N2244, N810);
nand NAND2 (N3457, N3451, N276);
and AND2 (N3458, N3446, N2772);
nand NAND2 (N3459, N3449, N650);
or OR3 (N3460, N3445, N2878, N2999);
nand NAND2 (N3461, N3459, N2333);
nand NAND4 (N3462, N3447, N1716, N159, N1195);
buf BUF1 (N3463, N3452);
and AND4 (N3464, N3457, N3023, N1926, N978);
and AND4 (N3465, N3458, N1931, N3433, N2246);
not NOT1 (N3466, N3461);
and AND2 (N3467, N3466, N615);
or OR4 (N3468, N3464, N622, N1801, N2098);
nor NOR2 (N3469, N3443, N668);
nor NOR3 (N3470, N3456, N1200, N3265);
buf BUF1 (N3471, N3463);
nor NOR2 (N3472, N3462, N1284);
or OR3 (N3473, N3470, N1562, N3132);
buf BUF1 (N3474, N3473);
or OR3 (N3475, N3468, N2083, N223);
nor NOR3 (N3476, N3450, N2513, N3065);
nor NOR3 (N3477, N3455, N2695, N1560);
nor NOR4 (N3478, N3472, N1961, N2965, N2132);
not NOT1 (N3479, N3471);
or OR4 (N3480, N3475, N3047, N754, N3199);
buf BUF1 (N3481, N3460);
nor NOR2 (N3482, N3474, N2646);
not NOT1 (N3483, N3469);
nor NOR3 (N3484, N3477, N847, N2698);
buf BUF1 (N3485, N3480);
nor NOR3 (N3486, N3476, N2250, N1354);
nand NAND3 (N3487, N3465, N1414, N1019);
nand NAND2 (N3488, N3467, N208);
nor NOR2 (N3489, N3486, N1466);
buf BUF1 (N3490, N3485);
not NOT1 (N3491, N3489);
and AND3 (N3492, N3487, N2051, N1421);
or OR2 (N3493, N3482, N1833);
xor XOR2 (N3494, N3490, N774);
buf BUF1 (N3495, N3493);
nand NAND2 (N3496, N3479, N731);
not NOT1 (N3497, N3481);
or OR3 (N3498, N3478, N3263, N471);
or OR3 (N3499, N3491, N958, N3464);
or OR2 (N3500, N3497, N3224);
not NOT1 (N3501, N3500);
not NOT1 (N3502, N3488);
not NOT1 (N3503, N3484);
not NOT1 (N3504, N3483);
or OR2 (N3505, N3492, N3122);
and AND4 (N3506, N3503, N2849, N1445, N2759);
not NOT1 (N3507, N3506);
nand NAND4 (N3508, N3494, N704, N714, N1908);
not NOT1 (N3509, N3496);
xor XOR2 (N3510, N3509, N2008);
and AND4 (N3511, N3505, N1643, N131, N720);
or OR4 (N3512, N3510, N1925, N2758, N83);
nand NAND3 (N3513, N3495, N454, N2139);
xor XOR2 (N3514, N3501, N3253);
or OR4 (N3515, N3511, N534, N1111, N99);
xor XOR2 (N3516, N3515, N1189);
xor XOR2 (N3517, N3498, N2676);
and AND4 (N3518, N3508, N2487, N3344, N2154);
or OR4 (N3519, N3516, N1770, N2378, N2550);
buf BUF1 (N3520, N3513);
buf BUF1 (N3521, N3520);
buf BUF1 (N3522, N3514);
and AND4 (N3523, N3518, N197, N3077, N1140);
or OR3 (N3524, N3521, N2906, N2969);
nor NOR3 (N3525, N3523, N884, N921);
or OR4 (N3526, N3504, N2785, N571, N2819);
not NOT1 (N3527, N3512);
buf BUF1 (N3528, N3527);
not NOT1 (N3529, N3502);
and AND4 (N3530, N3529, N3388, N585, N1807);
not NOT1 (N3531, N3507);
not NOT1 (N3532, N3519);
and AND3 (N3533, N3524, N904, N2205);
not NOT1 (N3534, N3499);
xor XOR2 (N3535, N3532, N1612);
nor NOR4 (N3536, N3528, N2884, N1325, N125);
buf BUF1 (N3537, N3533);
not NOT1 (N3538, N3530);
xor XOR2 (N3539, N3534, N1609);
nand NAND2 (N3540, N3539, N2802);
or OR2 (N3541, N3531, N2557);
xor XOR2 (N3542, N3541, N2878);
xor XOR2 (N3543, N3536, N2002);
nand NAND2 (N3544, N3517, N2255);
nor NOR4 (N3545, N3542, N1464, N801, N3403);
xor XOR2 (N3546, N3538, N756);
or OR4 (N3547, N3535, N404, N614, N179);
not NOT1 (N3548, N3537);
nor NOR4 (N3549, N3544, N3042, N1820, N1089);
buf BUF1 (N3550, N3547);
nor NOR2 (N3551, N3540, N3232);
buf BUF1 (N3552, N3543);
nor NOR2 (N3553, N3550, N1320);
buf BUF1 (N3554, N3553);
buf BUF1 (N3555, N3549);
nand NAND2 (N3556, N3525, N1014);
not NOT1 (N3557, N3526);
or OR4 (N3558, N3554, N3181, N2388, N2755);
and AND4 (N3559, N3548, N2414, N1031, N1688);
nand NAND2 (N3560, N3545, N2799);
buf BUF1 (N3561, N3555);
nand NAND4 (N3562, N3560, N1871, N1816, N383);
xor XOR2 (N3563, N3561, N3008);
and AND2 (N3564, N3563, N412);
nand NAND4 (N3565, N3551, N1488, N2743, N14);
nand NAND2 (N3566, N3546, N597);
or OR2 (N3567, N3556, N3545);
or OR4 (N3568, N3566, N1328, N631, N352);
or OR2 (N3569, N3552, N660);
xor XOR2 (N3570, N3569, N1669);
buf BUF1 (N3571, N3568);
not NOT1 (N3572, N3564);
and AND3 (N3573, N3522, N636, N1592);
nand NAND3 (N3574, N3571, N2508, N2463);
xor XOR2 (N3575, N3567, N318);
not NOT1 (N3576, N3559);
or OR4 (N3577, N3570, N3011, N922, N1769);
buf BUF1 (N3578, N3576);
nand NAND2 (N3579, N3558, N1336);
not NOT1 (N3580, N3573);
nand NAND3 (N3581, N3557, N1294, N196);
buf BUF1 (N3582, N3565);
not NOT1 (N3583, N3580);
nor NOR4 (N3584, N3583, N2414, N1903, N1470);
nand NAND4 (N3585, N3577, N2405, N1955, N1482);
nand NAND4 (N3586, N3575, N1205, N2578, N1802);
or OR2 (N3587, N3584, N1518);
xor XOR2 (N3588, N3585, N3247);
xor XOR2 (N3589, N3582, N822);
not NOT1 (N3590, N3579);
xor XOR2 (N3591, N3590, N3035);
and AND4 (N3592, N3562, N1877, N121, N2379);
nand NAND2 (N3593, N3586, N3019);
not NOT1 (N3594, N3572);
not NOT1 (N3595, N3587);
nand NAND2 (N3596, N3592, N1400);
nor NOR4 (N3597, N3595, N2748, N206, N3544);
or OR4 (N3598, N3596, N2876, N495, N1629);
xor XOR2 (N3599, N3588, N779);
not NOT1 (N3600, N3589);
xor XOR2 (N3601, N3599, N3260);
xor XOR2 (N3602, N3578, N568);
nor NOR4 (N3603, N3602, N1842, N3039, N999);
nand NAND3 (N3604, N3591, N246, N2622);
xor XOR2 (N3605, N3593, N1699);
and AND3 (N3606, N3605, N2057, N3090);
xor XOR2 (N3607, N3601, N3158);
or OR3 (N3608, N3604, N2141, N389);
buf BUF1 (N3609, N3600);
nand NAND4 (N3610, N3594, N3357, N2365, N3088);
xor XOR2 (N3611, N3598, N2469);
and AND2 (N3612, N3606, N1005);
nand NAND2 (N3613, N3612, N2019);
nor NOR4 (N3614, N3574, N230, N1310, N1355);
not NOT1 (N3615, N3607);
xor XOR2 (N3616, N3597, N3171);
buf BUF1 (N3617, N3613);
not NOT1 (N3618, N3610);
buf BUF1 (N3619, N3603);
and AND2 (N3620, N3614, N2034);
nand NAND3 (N3621, N3617, N947, N1451);
xor XOR2 (N3622, N3616, N2066);
or OR3 (N3623, N3608, N2665, N2739);
buf BUF1 (N3624, N3622);
buf BUF1 (N3625, N3618);
and AND3 (N3626, N3625, N1200, N2467);
nor NOR4 (N3627, N3624, N873, N80, N3624);
xor XOR2 (N3628, N3620, N93);
and AND3 (N3629, N3609, N2773, N3244);
xor XOR2 (N3630, N3621, N2237);
nor NOR2 (N3631, N3630, N3182);
nor NOR2 (N3632, N3626, N156);
buf BUF1 (N3633, N3615);
or OR3 (N3634, N3631, N2841, N936);
xor XOR2 (N3635, N3633, N1662);
or OR3 (N3636, N3611, N2016, N1759);
and AND4 (N3637, N3581, N1550, N545, N942);
nor NOR4 (N3638, N3637, N636, N3137, N3024);
nor NOR2 (N3639, N3628, N3127);
not NOT1 (N3640, N3634);
nand NAND4 (N3641, N3627, N693, N253, N394);
and AND3 (N3642, N3623, N2721, N1181);
and AND4 (N3643, N3638, N207, N2852, N1219);
buf BUF1 (N3644, N3629);
and AND3 (N3645, N3642, N3321, N1953);
xor XOR2 (N3646, N3619, N2032);
nand NAND2 (N3647, N3645, N2017);
nor NOR3 (N3648, N3644, N601, N1094);
and AND2 (N3649, N3632, N625);
or OR4 (N3650, N3640, N2616, N577, N515);
xor XOR2 (N3651, N3641, N1412);
nand NAND2 (N3652, N3646, N879);
or OR3 (N3653, N3639, N3484, N3503);
not NOT1 (N3654, N3648);
nand NAND3 (N3655, N3653, N1783, N3596);
and AND2 (N3656, N3636, N2156);
and AND3 (N3657, N3651, N1548, N2382);
or OR3 (N3658, N3652, N1418, N3093);
nor NOR2 (N3659, N3655, N848);
nand NAND3 (N3660, N3654, N2337, N2773);
and AND4 (N3661, N3656, N831, N100, N954);
buf BUF1 (N3662, N3658);
or OR2 (N3663, N3643, N77);
and AND3 (N3664, N3661, N3176, N2655);
buf BUF1 (N3665, N3660);
and AND4 (N3666, N3664, N3586, N794, N2854);
or OR4 (N3667, N3663, N2683, N3173, N2771);
and AND2 (N3668, N3666, N1113);
not NOT1 (N3669, N3657);
xor XOR2 (N3670, N3650, N2448);
nor NOR2 (N3671, N3669, N209);
not NOT1 (N3672, N3635);
nand NAND3 (N3673, N3662, N1005, N1533);
nand NAND4 (N3674, N3668, N939, N2251, N266);
and AND2 (N3675, N3671, N3664);
xor XOR2 (N3676, N3665, N2613);
and AND2 (N3677, N3675, N981);
not NOT1 (N3678, N3673);
xor XOR2 (N3679, N3678, N1786);
nand NAND2 (N3680, N3672, N1205);
nor NOR2 (N3681, N3676, N3077);
nand NAND2 (N3682, N3677, N1242);
or OR2 (N3683, N3649, N113);
or OR2 (N3684, N3674, N1931);
or OR3 (N3685, N3684, N970, N297);
not NOT1 (N3686, N3667);
or OR4 (N3687, N3681, N2912, N6, N1147);
or OR4 (N3688, N3670, N2804, N2840, N45);
buf BUF1 (N3689, N3688);
not NOT1 (N3690, N3687);
buf BUF1 (N3691, N3686);
or OR2 (N3692, N3647, N353);
nand NAND3 (N3693, N3683, N1276, N1771);
and AND2 (N3694, N3659, N2456);
buf BUF1 (N3695, N3694);
buf BUF1 (N3696, N3693);
nor NOR4 (N3697, N3680, N905, N1750, N1838);
nand NAND3 (N3698, N3691, N398, N29);
and AND4 (N3699, N3685, N2676, N2487, N1108);
or OR4 (N3700, N3682, N3018, N3333, N2342);
and AND3 (N3701, N3698, N2571, N3350);
and AND2 (N3702, N3697, N2785);
not NOT1 (N3703, N3690);
nor NOR4 (N3704, N3703, N3213, N1333, N46);
xor XOR2 (N3705, N3702, N2281);
or OR4 (N3706, N3704, N1627, N174, N851);
not NOT1 (N3707, N3695);
nand NAND4 (N3708, N3706, N2421, N777, N1313);
nand NAND2 (N3709, N3707, N1653);
not NOT1 (N3710, N3708);
nor NOR2 (N3711, N3710, N3272);
not NOT1 (N3712, N3701);
not NOT1 (N3713, N3711);
xor XOR2 (N3714, N3696, N2170);
and AND4 (N3715, N3705, N1099, N1323, N1221);
nand NAND4 (N3716, N3679, N1795, N3109, N388);
and AND2 (N3717, N3712, N2059);
buf BUF1 (N3718, N3714);
xor XOR2 (N3719, N3716, N919);
buf BUF1 (N3720, N3715);
nor NOR4 (N3721, N3689, N2857, N210, N2781);
nor NOR3 (N3722, N3699, N2137, N89);
buf BUF1 (N3723, N3709);
not NOT1 (N3724, N3713);
nor NOR3 (N3725, N3717, N703, N1702);
or OR2 (N3726, N3700, N1875);
and AND4 (N3727, N3692, N264, N320, N2675);
buf BUF1 (N3728, N3725);
not NOT1 (N3729, N3727);
nor NOR3 (N3730, N3726, N15, N3515);
nor NOR3 (N3731, N3720, N2292, N3456);
and AND4 (N3732, N3721, N1760, N37, N3399);
not NOT1 (N3733, N3731);
buf BUF1 (N3734, N3728);
nor NOR4 (N3735, N3732, N2604, N1190, N2282);
xor XOR2 (N3736, N3730, N2807);
not NOT1 (N3737, N3729);
or OR2 (N3738, N3723, N2044);
buf BUF1 (N3739, N3738);
nor NOR2 (N3740, N3735, N1646);
buf BUF1 (N3741, N3740);
nand NAND4 (N3742, N3734, N3558, N2905, N3206);
nor NOR2 (N3743, N3742, N425);
and AND3 (N3744, N3719, N2347, N3526);
nand NAND4 (N3745, N3743, N3692, N2843, N440);
not NOT1 (N3746, N3724);
not NOT1 (N3747, N3739);
buf BUF1 (N3748, N3737);
nor NOR3 (N3749, N3744, N3569, N1529);
nand NAND2 (N3750, N3722, N486);
nand NAND3 (N3751, N3749, N2099, N3426);
nand NAND4 (N3752, N3747, N2096, N3279, N349);
nand NAND2 (N3753, N3748, N282);
nor NOR3 (N3754, N3753, N1967, N1862);
nand NAND2 (N3755, N3751, N1227);
and AND3 (N3756, N3750, N1283, N1818);
nor NOR4 (N3757, N3754, N2810, N1609, N825);
nor NOR2 (N3758, N3755, N1682);
not NOT1 (N3759, N3756);
and AND2 (N3760, N3736, N453);
or OR2 (N3761, N3745, N2545);
or OR3 (N3762, N3741, N1390, N1842);
not NOT1 (N3763, N3759);
and AND2 (N3764, N3761, N1343);
and AND2 (N3765, N3762, N2928);
buf BUF1 (N3766, N3758);
nand NAND4 (N3767, N3752, N701, N1281, N3740);
xor XOR2 (N3768, N3766, N801);
nor NOR3 (N3769, N3764, N143, N1768);
nor NOR4 (N3770, N3733, N3719, N1489, N1156);
not NOT1 (N3771, N3768);
or OR2 (N3772, N3767, N412);
nor NOR2 (N3773, N3770, N578);
not NOT1 (N3774, N3773);
not NOT1 (N3775, N3763);
not NOT1 (N3776, N3772);
not NOT1 (N3777, N3757);
buf BUF1 (N3778, N3769);
xor XOR2 (N3779, N3775, N111);
nor NOR3 (N3780, N3771, N1548, N2499);
and AND3 (N3781, N3760, N70, N539);
buf BUF1 (N3782, N3776);
nor NOR4 (N3783, N3782, N3275, N3092, N3657);
and AND4 (N3784, N3765, N3692, N2913, N2212);
not NOT1 (N3785, N3777);
and AND2 (N3786, N3718, N3362);
and AND2 (N3787, N3781, N260);
buf BUF1 (N3788, N3778);
buf BUF1 (N3789, N3783);
or OR4 (N3790, N3784, N1063, N3480, N646);
nor NOR3 (N3791, N3790, N2778, N3377);
nor NOR3 (N3792, N3789, N450, N1060);
xor XOR2 (N3793, N3786, N3155);
and AND2 (N3794, N3787, N641);
not NOT1 (N3795, N3785);
or OR3 (N3796, N3794, N966, N1960);
and AND2 (N3797, N3780, N3767);
nor NOR4 (N3798, N3796, N48, N3521, N2199);
buf BUF1 (N3799, N3791);
nand NAND3 (N3800, N3792, N3274, N807);
and AND2 (N3801, N3774, N1497);
or OR2 (N3802, N3797, N2368);
nor NOR3 (N3803, N3801, N1336, N3526);
and AND2 (N3804, N3793, N2122);
or OR3 (N3805, N3799, N2340, N899);
or OR3 (N3806, N3795, N2278, N1749);
xor XOR2 (N3807, N3746, N3744);
buf BUF1 (N3808, N3803);
nor NOR2 (N3809, N3805, N2902);
not NOT1 (N3810, N3808);
and AND4 (N3811, N3804, N2070, N2362, N678);
not NOT1 (N3812, N3811);
xor XOR2 (N3813, N3798, N3427);
or OR4 (N3814, N3806, N1381, N2393, N3369);
buf BUF1 (N3815, N3810);
buf BUF1 (N3816, N3813);
and AND4 (N3817, N3814, N3724, N583, N3169);
and AND4 (N3818, N3800, N565, N6, N3746);
or OR4 (N3819, N3802, N1979, N3257, N2994);
and AND2 (N3820, N3779, N1050);
and AND3 (N3821, N3818, N2176, N1510);
and AND4 (N3822, N3819, N50, N923, N548);
and AND4 (N3823, N3817, N3388, N1144, N3469);
and AND3 (N3824, N3816, N1198, N2198);
buf BUF1 (N3825, N3823);
nor NOR2 (N3826, N3788, N3029);
and AND4 (N3827, N3815, N2659, N3377, N1855);
buf BUF1 (N3828, N3809);
xor XOR2 (N3829, N3807, N1116);
and AND3 (N3830, N3820, N2981, N716);
and AND3 (N3831, N3826, N3674, N3830);
nand NAND4 (N3832, N1938, N2206, N1094, N3482);
nand NAND4 (N3833, N3812, N141, N1320, N1081);
or OR3 (N3834, N3821, N468, N1805);
not NOT1 (N3835, N3829);
nor NOR4 (N3836, N3834, N1626, N1925, N2301);
buf BUF1 (N3837, N3832);
nor NOR3 (N3838, N3836, N1470, N1606);
nand NAND2 (N3839, N3822, N3722);
and AND4 (N3840, N3828, N2756, N278, N1466);
not NOT1 (N3841, N3825);
xor XOR2 (N3842, N3839, N2033);
or OR3 (N3843, N3841, N1897, N2266);
xor XOR2 (N3844, N3842, N1480);
nand NAND2 (N3845, N3827, N3442);
and AND3 (N3846, N3837, N3626, N3091);
nor NOR3 (N3847, N3845, N350, N3805);
or OR2 (N3848, N3831, N1739);
or OR4 (N3849, N3843, N991, N3818, N428);
nand NAND4 (N3850, N3848, N3526, N91, N1492);
or OR2 (N3851, N3833, N2380);
or OR2 (N3852, N3840, N3556);
buf BUF1 (N3853, N3824);
and AND4 (N3854, N3850, N1840, N1955, N951);
nand NAND4 (N3855, N3854, N3575, N823, N804);
xor XOR2 (N3856, N3846, N477);
nand NAND2 (N3857, N3852, N3124);
or OR3 (N3858, N3844, N1519, N8);
xor XOR2 (N3859, N3849, N3518);
nand NAND3 (N3860, N3838, N1139, N1762);
not NOT1 (N3861, N3858);
buf BUF1 (N3862, N3835);
xor XOR2 (N3863, N3847, N2618);
buf BUF1 (N3864, N3856);
and AND3 (N3865, N3859, N3531, N1772);
buf BUF1 (N3866, N3862);
xor XOR2 (N3867, N3866, N2673);
xor XOR2 (N3868, N3853, N673);
buf BUF1 (N3869, N3868);
xor XOR2 (N3870, N3867, N2151);
and AND4 (N3871, N3851, N3845, N3357, N2115);
nor NOR4 (N3872, N3855, N3015, N3443, N3387);
or OR4 (N3873, N3872, N1475, N3541, N3177);
not NOT1 (N3874, N3870);
buf BUF1 (N3875, N3860);
buf BUF1 (N3876, N3864);
not NOT1 (N3877, N3861);
nand NAND3 (N3878, N3874, N2245, N3010);
not NOT1 (N3879, N3871);
and AND4 (N3880, N3857, N2807, N3713, N2884);
not NOT1 (N3881, N3877);
or OR4 (N3882, N3878, N1276, N2684, N2077);
nand NAND4 (N3883, N3879, N2957, N139, N343);
and AND4 (N3884, N3883, N2952, N3409, N3273);
xor XOR2 (N3885, N3884, N1204);
xor XOR2 (N3886, N3885, N2860);
xor XOR2 (N3887, N3881, N852);
or OR4 (N3888, N3887, N2650, N3146, N544);
buf BUF1 (N3889, N3886);
nor NOR4 (N3890, N3873, N1475, N2877, N910);
nand NAND3 (N3891, N3865, N2761, N2476);
or OR4 (N3892, N3891, N605, N2958, N1568);
or OR4 (N3893, N3889, N993, N2988, N2005);
nand NAND4 (N3894, N3876, N2582, N3018, N3847);
nor NOR3 (N3895, N3863, N152, N3439);
buf BUF1 (N3896, N3894);
or OR2 (N3897, N3890, N3654);
not NOT1 (N3898, N3896);
not NOT1 (N3899, N3898);
or OR3 (N3900, N3899, N1486, N2219);
buf BUF1 (N3901, N3900);
nand NAND2 (N3902, N3882, N1694);
buf BUF1 (N3903, N3902);
nand NAND3 (N3904, N3901, N693, N2898);
nand NAND2 (N3905, N3875, N698);
and AND4 (N3906, N3869, N3008, N910, N2916);
nand NAND2 (N3907, N3888, N3050);
nand NAND3 (N3908, N3904, N3781, N833);
not NOT1 (N3909, N3905);
or OR2 (N3910, N3906, N2759);
and AND2 (N3911, N3909, N1118);
nor NOR2 (N3912, N3897, N3893);
nand NAND2 (N3913, N536, N1491);
not NOT1 (N3914, N3880);
or OR4 (N3915, N3903, N1776, N2521, N1062);
buf BUF1 (N3916, N3892);
and AND4 (N3917, N3907, N3632, N883, N3688);
and AND2 (N3918, N3914, N3117);
not NOT1 (N3919, N3916);
not NOT1 (N3920, N3919);
nor NOR2 (N3921, N3913, N2028);
buf BUF1 (N3922, N3921);
nor NOR4 (N3923, N3922, N1743, N2778, N808);
nand NAND4 (N3924, N3920, N1453, N3335, N3108);
not NOT1 (N3925, N3912);
not NOT1 (N3926, N3915);
nor NOR3 (N3927, N3910, N2111, N319);
nor NOR4 (N3928, N3911, N699, N2021, N1901);
and AND3 (N3929, N3917, N591, N1042);
or OR3 (N3930, N3926, N3280, N2068);
or OR4 (N3931, N3924, N2143, N1666, N3773);
buf BUF1 (N3932, N3929);
nand NAND4 (N3933, N3895, N1046, N3539, N172);
and AND4 (N3934, N3932, N1004, N40, N417);
and AND4 (N3935, N3931, N2044, N437, N2164);
and AND2 (N3936, N3908, N1800);
nor NOR3 (N3937, N3927, N3193, N464);
xor XOR2 (N3938, N3934, N109);
not NOT1 (N3939, N3936);
buf BUF1 (N3940, N3928);
nand NAND3 (N3941, N3918, N1596, N495);
buf BUF1 (N3942, N3923);
nor NOR4 (N3943, N3937, N2317, N241, N2019);
buf BUF1 (N3944, N3939);
nand NAND4 (N3945, N3938, N2513, N2831, N3435);
buf BUF1 (N3946, N3935);
buf BUF1 (N3947, N3945);
nor NOR3 (N3948, N3942, N6, N1125);
and AND4 (N3949, N3925, N2013, N1109, N3702);
and AND3 (N3950, N3943, N2757, N137);
or OR4 (N3951, N3930, N3206, N2892, N3947);
nor NOR4 (N3952, N2931, N2117, N2385, N538);
or OR3 (N3953, N3933, N231, N1132);
nor NOR4 (N3954, N3941, N2844, N3041, N186);
not NOT1 (N3955, N3948);
nor NOR2 (N3956, N3953, N1940);
nand NAND2 (N3957, N3954, N2345);
buf BUF1 (N3958, N3956);
and AND2 (N3959, N3946, N3261);
not NOT1 (N3960, N3959);
or OR4 (N3961, N3957, N2357, N2099, N618);
and AND4 (N3962, N3950, N1850, N1368, N3328);
not NOT1 (N3963, N3961);
nor NOR3 (N3964, N3955, N840, N3230);
nor NOR2 (N3965, N3951, N390);
or OR4 (N3966, N3944, N983, N3385, N246);
or OR2 (N3967, N3940, N2317);
nand NAND3 (N3968, N3967, N1093, N1680);
xor XOR2 (N3969, N3966, N2295);
nand NAND4 (N3970, N3958, N2550, N1133, N3634);
xor XOR2 (N3971, N3960, N2131);
not NOT1 (N3972, N3971);
nor NOR2 (N3973, N3963, N2617);
or OR4 (N3974, N3969, N1079, N1134, N297);
not NOT1 (N3975, N3965);
nor NOR2 (N3976, N3975, N137);
not NOT1 (N3977, N3962);
xor XOR2 (N3978, N3949, N1837);
not NOT1 (N3979, N3974);
or OR4 (N3980, N3979, N777, N3394, N3400);
not NOT1 (N3981, N3980);
buf BUF1 (N3982, N3973);
nor NOR3 (N3983, N3976, N2699, N1082);
and AND4 (N3984, N3981, N2190, N3163, N2089);
buf BUF1 (N3985, N3952);
xor XOR2 (N3986, N3968, N2350);
nor NOR2 (N3987, N3984, N2111);
and AND4 (N3988, N3970, N2569, N1243, N1126);
xor XOR2 (N3989, N3988, N3889);
not NOT1 (N3990, N3985);
nand NAND3 (N3991, N3987, N1093, N281);
nand NAND2 (N3992, N3989, N2579);
or OR3 (N3993, N3972, N1699, N1449);
nand NAND3 (N3994, N3983, N3372, N950);
and AND4 (N3995, N3991, N1884, N2605, N3506);
not NOT1 (N3996, N3977);
nand NAND4 (N3997, N3978, N3392, N19, N1881);
xor XOR2 (N3998, N3986, N291);
nand NAND3 (N3999, N3964, N1243, N1589);
or OR4 (N4000, N3998, N1657, N381, N2729);
not NOT1 (N4001, N3996);
xor XOR2 (N4002, N3990, N754);
nor NOR3 (N4003, N3992, N2469, N865);
nor NOR2 (N4004, N3994, N265);
buf BUF1 (N4005, N3995);
nor NOR2 (N4006, N4002, N558);
buf BUF1 (N4007, N4003);
or OR3 (N4008, N4007, N2274, N2144);
or OR4 (N4009, N4000, N2699, N1259, N3262);
xor XOR2 (N4010, N3982, N3050);
nand NAND4 (N4011, N4006, N1766, N1287, N1467);
and AND2 (N4012, N3999, N3657);
xor XOR2 (N4013, N4010, N3073);
or OR4 (N4014, N4011, N1814, N1125, N3522);
not NOT1 (N4015, N4014);
not NOT1 (N4016, N4008);
xor XOR2 (N4017, N4015, N1816);
and AND4 (N4018, N4012, N80, N505, N2994);
nor NOR3 (N4019, N3993, N1487, N120);
buf BUF1 (N4020, N4013);
nand NAND4 (N4021, N4001, N2979, N3487, N938);
not NOT1 (N4022, N4018);
not NOT1 (N4023, N4016);
nand NAND3 (N4024, N4020, N3710, N2121);
xor XOR2 (N4025, N4019, N164);
buf BUF1 (N4026, N4021);
and AND2 (N4027, N4022, N1451);
nor NOR4 (N4028, N4024, N1030, N1323, N2727);
xor XOR2 (N4029, N4004, N232);
nand NAND4 (N4030, N4026, N3604, N1967, N594);
nor NOR2 (N4031, N4009, N888);
buf BUF1 (N4032, N4031);
not NOT1 (N4033, N4029);
and AND2 (N4034, N4032, N26);
buf BUF1 (N4035, N4023);
or OR3 (N4036, N4025, N699, N1279);
nand NAND4 (N4037, N4030, N1598, N3540, N2230);
nor NOR2 (N4038, N4028, N714);
nand NAND4 (N4039, N4034, N1860, N362, N2382);
buf BUF1 (N4040, N4037);
not NOT1 (N4041, N4035);
not NOT1 (N4042, N4033);
or OR4 (N4043, N4017, N2111, N3312, N1897);
or OR3 (N4044, N4042, N3860, N2251);
nand NAND4 (N4045, N4005, N3503, N3914, N1402);
xor XOR2 (N4046, N4041, N3073);
not NOT1 (N4047, N4038);
xor XOR2 (N4048, N4047, N3916);
and AND2 (N4049, N4027, N3421);
or OR3 (N4050, N4040, N3739, N4043);
xor XOR2 (N4051, N475, N1653);
or OR2 (N4052, N4046, N2874);
nor NOR2 (N4053, N4045, N3476);
and AND3 (N4054, N4036, N3616, N2128);
not NOT1 (N4055, N3997);
nand NAND3 (N4056, N4048, N3074, N1427);
buf BUF1 (N4057, N4052);
not NOT1 (N4058, N4044);
not NOT1 (N4059, N4049);
and AND2 (N4060, N4050, N2039);
nand NAND3 (N4061, N4055, N3391, N1784);
not NOT1 (N4062, N4061);
buf BUF1 (N4063, N4058);
buf BUF1 (N4064, N4039);
and AND3 (N4065, N4063, N1853, N348);
and AND3 (N4066, N4059, N853, N1364);
not NOT1 (N4067, N4060);
not NOT1 (N4068, N4065);
and AND3 (N4069, N4051, N2196, N2832);
buf BUF1 (N4070, N4057);
nor NOR3 (N4071, N4066, N3786, N3820);
xor XOR2 (N4072, N4070, N3195);
nor NOR2 (N4073, N4069, N1604);
nor NOR2 (N4074, N4067, N3415);
or OR2 (N4075, N4068, N741);
nand NAND2 (N4076, N4064, N1596);
or OR2 (N4077, N4054, N1973);
and AND3 (N4078, N4072, N1864, N1094);
and AND4 (N4079, N4056, N3425, N3328, N1064);
xor XOR2 (N4080, N4073, N2406);
not NOT1 (N4081, N4053);
not NOT1 (N4082, N4076);
xor XOR2 (N4083, N4075, N535);
xor XOR2 (N4084, N4071, N1878);
and AND3 (N4085, N4074, N2275, N3906);
not NOT1 (N4086, N4077);
nor NOR4 (N4087, N4083, N2925, N3300, N311);
nor NOR4 (N4088, N4062, N2289, N2362, N1109);
xor XOR2 (N4089, N4086, N257);
and AND4 (N4090, N4078, N3099, N2343, N1544);
buf BUF1 (N4091, N4089);
not NOT1 (N4092, N4085);
or OR2 (N4093, N4084, N3299);
not NOT1 (N4094, N4092);
buf BUF1 (N4095, N4094);
nor NOR3 (N4096, N4080, N1650, N3767);
nand NAND2 (N4097, N4093, N3211);
nor NOR2 (N4098, N4081, N3790);
or OR2 (N4099, N4097, N1737);
buf BUF1 (N4100, N4091);
nand NAND2 (N4101, N4088, N31);
and AND3 (N4102, N4099, N2703, N2065);
or OR4 (N4103, N4087, N3265, N1656, N4065);
buf BUF1 (N4104, N4100);
or OR3 (N4105, N4102, N1757, N666);
nor NOR2 (N4106, N4105, N1421);
and AND4 (N4107, N4104, N3492, N542, N2760);
nand NAND3 (N4108, N4082, N3757, N926);
nand NAND2 (N4109, N4090, N1095);
buf BUF1 (N4110, N4103);
nor NOR4 (N4111, N4096, N2395, N3051, N3912);
not NOT1 (N4112, N4106);
and AND3 (N4113, N4111, N1361, N1592);
nand NAND4 (N4114, N4107, N2339, N3085, N3263);
and AND4 (N4115, N4113, N838, N3949, N3768);
nor NOR3 (N4116, N4095, N58, N3182);
or OR2 (N4117, N4108, N1586);
not NOT1 (N4118, N4117);
xor XOR2 (N4119, N4112, N1591);
and AND3 (N4120, N4109, N2875, N891);
nor NOR3 (N4121, N4110, N1688, N2473);
not NOT1 (N4122, N4115);
not NOT1 (N4123, N4121);
nor NOR4 (N4124, N4118, N2123, N2606, N801);
not NOT1 (N4125, N4124);
nand NAND3 (N4126, N4125, N2900, N2293);
buf BUF1 (N4127, N4101);
and AND3 (N4128, N4122, N807, N387);
nand NAND4 (N4129, N4128, N321, N3791, N244);
nand NAND4 (N4130, N4126, N1246, N2768, N4118);
buf BUF1 (N4131, N4098);
or OR2 (N4132, N4120, N1356);
buf BUF1 (N4133, N4131);
buf BUF1 (N4134, N4114);
xor XOR2 (N4135, N4129, N615);
nand NAND4 (N4136, N4135, N3870, N2044, N2825);
not NOT1 (N4137, N4130);
not NOT1 (N4138, N4127);
nor NOR4 (N4139, N4138, N1588, N3714, N4023);
nor NOR3 (N4140, N4119, N3112, N3964);
xor XOR2 (N4141, N4136, N2685);
or OR4 (N4142, N4134, N1833, N1586, N1039);
buf BUF1 (N4143, N4116);
nand NAND2 (N4144, N4142, N735);
xor XOR2 (N4145, N4133, N2732);
xor XOR2 (N4146, N4123, N297);
buf BUF1 (N4147, N4141);
and AND4 (N4148, N4137, N1163, N2391, N1552);
nand NAND4 (N4149, N4139, N4023, N3434, N756);
or OR4 (N4150, N4079, N1649, N1884, N3831);
xor XOR2 (N4151, N4132, N2785);
xor XOR2 (N4152, N4143, N2386);
nor NOR2 (N4153, N4145, N1354);
and AND2 (N4154, N4144, N1463);
xor XOR2 (N4155, N4151, N1903);
not NOT1 (N4156, N4148);
nor NOR2 (N4157, N4155, N3011);
xor XOR2 (N4158, N4147, N4055);
or OR3 (N4159, N4156, N2950, N4134);
xor XOR2 (N4160, N4149, N3233);
xor XOR2 (N4161, N4157, N2251);
and AND4 (N4162, N4150, N3848, N86, N73);
and AND3 (N4163, N4158, N814, N3780);
nor NOR2 (N4164, N4161, N316);
xor XOR2 (N4165, N4146, N2924);
xor XOR2 (N4166, N4163, N978);
or OR4 (N4167, N4165, N412, N3231, N2735);
xor XOR2 (N4168, N4167, N3476);
nand NAND2 (N4169, N4153, N3405);
xor XOR2 (N4170, N4160, N542);
xor XOR2 (N4171, N4166, N2368);
nor NOR4 (N4172, N4162, N3506, N3338, N2299);
xor XOR2 (N4173, N4172, N142);
buf BUF1 (N4174, N4173);
buf BUF1 (N4175, N4164);
and AND4 (N4176, N4174, N904, N1577, N3565);
nand NAND2 (N4177, N4168, N3192);
not NOT1 (N4178, N4175);
nand NAND2 (N4179, N4169, N941);
not NOT1 (N4180, N4152);
and AND4 (N4181, N4170, N328, N1094, N3466);
not NOT1 (N4182, N4159);
and AND4 (N4183, N4182, N3535, N223, N257);
not NOT1 (N4184, N4154);
buf BUF1 (N4185, N4177);
not NOT1 (N4186, N4178);
and AND2 (N4187, N4176, N3481);
and AND3 (N4188, N4179, N2676, N1574);
and AND3 (N4189, N4180, N3082, N2526);
nor NOR4 (N4190, N4187, N2132, N645, N4102);
not NOT1 (N4191, N4184);
buf BUF1 (N4192, N4171);
nand NAND2 (N4193, N4191, N2502);
and AND4 (N4194, N4140, N491, N1267, N3766);
nor NOR3 (N4195, N4189, N1747, N2266);
and AND4 (N4196, N4193, N918, N3595, N874);
nand NAND3 (N4197, N4183, N2274, N3564);
xor XOR2 (N4198, N4181, N1737);
nor NOR3 (N4199, N4188, N230, N1566);
nand NAND4 (N4200, N4195, N1554, N3291, N102);
xor XOR2 (N4201, N4197, N3490);
nor NOR3 (N4202, N4190, N3491, N3120);
buf BUF1 (N4203, N4199);
or OR3 (N4204, N4185, N1519, N2380);
nor NOR4 (N4205, N4186, N3989, N3524, N3765);
nand NAND2 (N4206, N4204, N228);
xor XOR2 (N4207, N4198, N1479);
xor XOR2 (N4208, N4194, N176);
and AND2 (N4209, N4196, N1417);
not NOT1 (N4210, N4205);
buf BUF1 (N4211, N4208);
or OR4 (N4212, N4209, N3277, N775, N1834);
xor XOR2 (N4213, N4203, N2372);
not NOT1 (N4214, N4206);
xor XOR2 (N4215, N4200, N165);
or OR4 (N4216, N4214, N850, N2148, N3551);
buf BUF1 (N4217, N4211);
buf BUF1 (N4218, N4217);
or OR2 (N4219, N4215, N3372);
and AND4 (N4220, N4210, N2106, N628, N4147);
nand NAND2 (N4221, N4201, N373);
buf BUF1 (N4222, N4207);
buf BUF1 (N4223, N4212);
buf BUF1 (N4224, N4221);
not NOT1 (N4225, N4223);
or OR4 (N4226, N4225, N3729, N2740, N2783);
or OR3 (N4227, N4222, N2945, N1218);
or OR3 (N4228, N4226, N1738, N720);
nor NOR3 (N4229, N4202, N3627, N3403);
nor NOR4 (N4230, N4227, N1392, N975, N682);
or OR4 (N4231, N4224, N3858, N2745, N3732);
and AND2 (N4232, N4216, N4122);
nand NAND2 (N4233, N4230, N4007);
or OR3 (N4234, N4218, N73, N1033);
nor NOR3 (N4235, N4220, N4072, N1106);
buf BUF1 (N4236, N4229);
nor NOR2 (N4237, N4233, N4198);
xor XOR2 (N4238, N4231, N3720);
xor XOR2 (N4239, N4235, N615);
or OR2 (N4240, N4219, N2671);
or OR2 (N4241, N4232, N3473);
not NOT1 (N4242, N4228);
or OR2 (N4243, N4236, N1188);
and AND3 (N4244, N4237, N960, N872);
buf BUF1 (N4245, N4234);
buf BUF1 (N4246, N4239);
nor NOR3 (N4247, N4238, N4203, N331);
or OR2 (N4248, N4246, N1952);
not NOT1 (N4249, N4247);
nor NOR2 (N4250, N4242, N2802);
not NOT1 (N4251, N4250);
nor NOR2 (N4252, N4251, N2137);
or OR2 (N4253, N4249, N1007);
and AND4 (N4254, N4244, N1974, N613, N3867);
xor XOR2 (N4255, N4243, N532);
nand NAND2 (N4256, N4192, N2556);
nor NOR3 (N4257, N4240, N241, N2101);
xor XOR2 (N4258, N4248, N3789);
xor XOR2 (N4259, N4252, N2830);
nand NAND4 (N4260, N4241, N487, N1390, N328);
or OR3 (N4261, N4245, N502, N567);
nand NAND4 (N4262, N4257, N1678, N2833, N855);
nand NAND4 (N4263, N4253, N4210, N313, N1785);
nor NOR2 (N4264, N4263, N2098);
nor NOR2 (N4265, N4213, N295);
xor XOR2 (N4266, N4256, N3843);
nand NAND4 (N4267, N4255, N302, N1798, N15);
and AND2 (N4268, N4265, N8);
nor NOR2 (N4269, N4259, N3990);
and AND4 (N4270, N4266, N263, N2104, N4055);
and AND2 (N4271, N4258, N1647);
nor NOR4 (N4272, N4261, N809, N3543, N1187);
not NOT1 (N4273, N4267);
xor XOR2 (N4274, N4260, N1555);
and AND2 (N4275, N4269, N439);
xor XOR2 (N4276, N4254, N3322);
or OR3 (N4277, N4275, N2789, N1988);
nor NOR2 (N4278, N4262, N2948);
and AND3 (N4279, N4273, N405, N3992);
nand NAND2 (N4280, N4268, N1210);
nor NOR4 (N4281, N4276, N3544, N2485, N920);
buf BUF1 (N4282, N4270);
not NOT1 (N4283, N4279);
xor XOR2 (N4284, N4272, N1451);
nor NOR3 (N4285, N4264, N411, N1589);
xor XOR2 (N4286, N4277, N3158);
and AND4 (N4287, N4286, N1454, N4185, N3679);
buf BUF1 (N4288, N4285);
xor XOR2 (N4289, N4278, N3808);
xor XOR2 (N4290, N4287, N2352);
or OR3 (N4291, N4281, N3770, N2959);
nor NOR3 (N4292, N4291, N2732, N142);
not NOT1 (N4293, N4274);
or OR3 (N4294, N4293, N3941, N451);
nor NOR2 (N4295, N4289, N2303);
xor XOR2 (N4296, N4294, N2727);
nand NAND3 (N4297, N4280, N735, N508);
not NOT1 (N4298, N4296);
buf BUF1 (N4299, N4297);
buf BUF1 (N4300, N4290);
xor XOR2 (N4301, N4299, N1322);
buf BUF1 (N4302, N4301);
buf BUF1 (N4303, N4288);
buf BUF1 (N4304, N4282);
not NOT1 (N4305, N4304);
and AND3 (N4306, N4303, N2449, N3965);
or OR4 (N4307, N4271, N973, N3111, N428);
not NOT1 (N4308, N4305);
xor XOR2 (N4309, N4308, N1762);
nor NOR3 (N4310, N4309, N3263, N740);
xor XOR2 (N4311, N4307, N2172);
nand NAND2 (N4312, N4311, N1077);
nor NOR3 (N4313, N4283, N2804, N4062);
buf BUF1 (N4314, N4310);
nor NOR4 (N4315, N4298, N1764, N1839, N639);
and AND3 (N4316, N4315, N3546, N1022);
buf BUF1 (N4317, N4306);
and AND3 (N4318, N4316, N2130, N3075);
not NOT1 (N4319, N4295);
buf BUF1 (N4320, N4312);
and AND3 (N4321, N4320, N60, N2295);
nor NOR3 (N4322, N4300, N2449, N209);
xor XOR2 (N4323, N4321, N4109);
or OR4 (N4324, N4314, N4300, N1993, N4183);
xor XOR2 (N4325, N4319, N724);
and AND3 (N4326, N4324, N1320, N3947);
buf BUF1 (N4327, N4323);
or OR3 (N4328, N4318, N2735, N3550);
or OR2 (N4329, N4317, N3954);
not NOT1 (N4330, N4292);
nor NOR2 (N4331, N4326, N624);
nand NAND4 (N4332, N4330, N786, N4081, N3284);
or OR4 (N4333, N4313, N1396, N2161, N3772);
and AND4 (N4334, N4284, N1497, N3425, N1626);
xor XOR2 (N4335, N4331, N1116);
not NOT1 (N4336, N4332);
nor NOR2 (N4337, N4335, N3415);
not NOT1 (N4338, N4334);
nand NAND4 (N4339, N4333, N3863, N2784, N2154);
nor NOR2 (N4340, N4302, N2740);
and AND3 (N4341, N4329, N1552, N1582);
nor NOR3 (N4342, N4325, N1179, N1328);
nor NOR2 (N4343, N4328, N1088);
not NOT1 (N4344, N4322);
buf BUF1 (N4345, N4337);
nor NOR2 (N4346, N4338, N3377);
nand NAND2 (N4347, N4339, N3388);
and AND4 (N4348, N4340, N3844, N3903, N1469);
and AND2 (N4349, N4327, N158);
xor XOR2 (N4350, N4348, N17);
xor XOR2 (N4351, N4350, N3791);
nand NAND2 (N4352, N4343, N4262);
nor NOR4 (N4353, N4349, N582, N4034, N2480);
xor XOR2 (N4354, N4351, N517);
nor NOR2 (N4355, N4352, N2144);
nor NOR3 (N4356, N4344, N3314, N2787);
or OR4 (N4357, N4345, N253, N1966, N504);
not NOT1 (N4358, N4336);
xor XOR2 (N4359, N4353, N3417);
not NOT1 (N4360, N4354);
or OR4 (N4361, N4341, N1779, N3788, N3037);
xor XOR2 (N4362, N4346, N3829);
or OR4 (N4363, N4357, N340, N3822, N3891);
nor NOR4 (N4364, N4355, N2644, N4309, N914);
nor NOR2 (N4365, N4347, N1434);
nand NAND2 (N4366, N4356, N3572);
buf BUF1 (N4367, N4361);
nand NAND3 (N4368, N4366, N599, N812);
nand NAND2 (N4369, N4368, N4309);
nor NOR2 (N4370, N4363, N3728);
and AND4 (N4371, N4360, N3328, N1645, N543);
and AND2 (N4372, N4370, N4023);
xor XOR2 (N4373, N4359, N261);
and AND2 (N4374, N4362, N767);
and AND3 (N4375, N4367, N490, N74);
nor NOR2 (N4376, N4365, N791);
buf BUF1 (N4377, N4364);
buf BUF1 (N4378, N4373);
xor XOR2 (N4379, N4371, N4014);
nor NOR4 (N4380, N4372, N2987, N2549, N2782);
nor NOR4 (N4381, N4378, N3583, N2861, N2851);
not NOT1 (N4382, N4374);
nor NOR2 (N4383, N4381, N3572);
nor NOR4 (N4384, N4369, N475, N838, N690);
xor XOR2 (N4385, N4383, N1297);
buf BUF1 (N4386, N4379);
xor XOR2 (N4387, N4375, N882);
and AND3 (N4388, N4358, N3215, N1984);
nor NOR2 (N4389, N4387, N1642);
and AND3 (N4390, N4388, N1897, N3825);
nor NOR3 (N4391, N4386, N3262, N3570);
and AND2 (N4392, N4376, N3453);
buf BUF1 (N4393, N4380);
or OR2 (N4394, N4342, N421);
nor NOR4 (N4395, N4393, N2760, N4056, N538);
or OR3 (N4396, N4390, N1781, N935);
xor XOR2 (N4397, N4394, N2137);
nor NOR2 (N4398, N4385, N1249);
buf BUF1 (N4399, N4397);
xor XOR2 (N4400, N4384, N2510);
or OR4 (N4401, N4391, N1707, N40, N1196);
and AND4 (N4402, N4399, N912, N1456, N3149);
nand NAND4 (N4403, N4392, N445, N1214, N1393);
xor XOR2 (N4404, N4377, N2079);
buf BUF1 (N4405, N4395);
and AND3 (N4406, N4404, N4181, N1135);
buf BUF1 (N4407, N4402);
nand NAND2 (N4408, N4400, N1879);
nand NAND4 (N4409, N4407, N3969, N3845, N3956);
not NOT1 (N4410, N4408);
not NOT1 (N4411, N4389);
not NOT1 (N4412, N4410);
nor NOR4 (N4413, N4403, N173, N2574, N1048);
or OR2 (N4414, N4382, N4183);
nand NAND4 (N4415, N4406, N2186, N738, N639);
buf BUF1 (N4416, N4398);
xor XOR2 (N4417, N4411, N1781);
or OR4 (N4418, N4412, N1664, N4219, N2917);
buf BUF1 (N4419, N4405);
or OR3 (N4420, N4401, N800, N3120);
or OR4 (N4421, N4409, N1553, N1897, N93);
xor XOR2 (N4422, N4418, N1858);
buf BUF1 (N4423, N4415);
nor NOR4 (N4424, N4417, N269, N1577, N3516);
xor XOR2 (N4425, N4421, N4323);
buf BUF1 (N4426, N4420);
not NOT1 (N4427, N4413);
nor NOR2 (N4428, N4396, N3832);
not NOT1 (N4429, N4426);
and AND4 (N4430, N4427, N1945, N3579, N185);
buf BUF1 (N4431, N4429);
nor NOR3 (N4432, N4431, N3167, N1400);
nor NOR3 (N4433, N4422, N2436, N1702);
nor NOR3 (N4434, N4414, N2327, N1833);
and AND4 (N4435, N4428, N1471, N3995, N1212);
or OR4 (N4436, N4435, N2247, N3545, N321);
or OR4 (N4437, N4425, N3619, N2072, N1477);
nor NOR4 (N4438, N4436, N3422, N1810, N1146);
not NOT1 (N4439, N4423);
buf BUF1 (N4440, N4439);
not NOT1 (N4441, N4433);
not NOT1 (N4442, N4440);
buf BUF1 (N4443, N4416);
and AND3 (N4444, N4442, N2082, N1847);
and AND3 (N4445, N4424, N3647, N1639);
nand NAND3 (N4446, N4438, N1677, N1117);
buf BUF1 (N4447, N4441);
not NOT1 (N4448, N4430);
buf BUF1 (N4449, N4434);
and AND2 (N4450, N4445, N1016);
nand NAND2 (N4451, N4444, N2667);
buf BUF1 (N4452, N4451);
or OR3 (N4453, N4452, N2008, N325);
not NOT1 (N4454, N4446);
and AND2 (N4455, N4450, N214);
not NOT1 (N4456, N4437);
buf BUF1 (N4457, N4454);
and AND3 (N4458, N4448, N2705, N3425);
not NOT1 (N4459, N4457);
nor NOR4 (N4460, N4447, N576, N540, N1334);
or OR4 (N4461, N4458, N1857, N3243, N4105);
nor NOR4 (N4462, N4453, N189, N3939, N2441);
or OR3 (N4463, N4460, N4123, N1008);
nor NOR3 (N4464, N4432, N1616, N3038);
xor XOR2 (N4465, N4443, N138);
buf BUF1 (N4466, N4459);
xor XOR2 (N4467, N4461, N78);
or OR2 (N4468, N4456, N885);
not NOT1 (N4469, N4419);
not NOT1 (N4470, N4463);
nand NAND3 (N4471, N4470, N3055, N1321);
or OR3 (N4472, N4468, N1190, N3185);
nand NAND4 (N4473, N4462, N2097, N2776, N3805);
not NOT1 (N4474, N4472);
nand NAND4 (N4475, N4473, N287, N641, N4339);
or OR2 (N4476, N4475, N1942);
or OR3 (N4477, N4464, N304, N2200);
xor XOR2 (N4478, N4466, N2585);
nor NOR2 (N4479, N4476, N4287);
or OR2 (N4480, N4471, N4119);
and AND3 (N4481, N4465, N3520, N4382);
nand NAND2 (N4482, N4455, N1738);
nand NAND2 (N4483, N4477, N1156);
or OR3 (N4484, N4478, N1945, N1086);
not NOT1 (N4485, N4479);
and AND3 (N4486, N4483, N2095, N2952);
buf BUF1 (N4487, N4469);
and AND2 (N4488, N4480, N3887);
and AND3 (N4489, N4488, N506, N4458);
nand NAND4 (N4490, N4467, N900, N4149, N2194);
and AND2 (N4491, N4489, N752);
buf BUF1 (N4492, N4482);
not NOT1 (N4493, N4474);
nand NAND4 (N4494, N4493, N53, N4355, N3667);
not NOT1 (N4495, N4481);
and AND3 (N4496, N4449, N2396, N4105);
buf BUF1 (N4497, N4491);
nand NAND3 (N4498, N4484, N1240, N1043);
nand NAND2 (N4499, N4497, N3583);
and AND4 (N4500, N4499, N3356, N1517, N1366);
not NOT1 (N4501, N4498);
or OR3 (N4502, N4487, N1516, N2215);
xor XOR2 (N4503, N4501, N3992);
and AND2 (N4504, N4486, N646);
buf BUF1 (N4505, N4485);
nor NOR3 (N4506, N4503, N1407, N3075);
nand NAND2 (N4507, N4500, N1345);
or OR4 (N4508, N4495, N610, N1432, N540);
nor NOR4 (N4509, N4490, N3772, N1697, N919);
not NOT1 (N4510, N4494);
or OR2 (N4511, N4510, N743);
not NOT1 (N4512, N4505);
xor XOR2 (N4513, N4496, N928);
not NOT1 (N4514, N4509);
and AND2 (N4515, N4506, N1529);
and AND4 (N4516, N4507, N3134, N1468, N3623);
not NOT1 (N4517, N4508);
or OR3 (N4518, N4511, N2753, N3260);
not NOT1 (N4519, N4492);
buf BUF1 (N4520, N4504);
or OR3 (N4521, N4520, N3418, N3393);
not NOT1 (N4522, N4519);
or OR3 (N4523, N4515, N4429, N2288);
or OR4 (N4524, N4514, N2584, N3794, N947);
nor NOR2 (N4525, N4512, N2625);
buf BUF1 (N4526, N4517);
and AND2 (N4527, N4526, N1996);
nor NOR3 (N4528, N4521, N2766, N3006);
xor XOR2 (N4529, N4525, N3066);
xor XOR2 (N4530, N4523, N575);
nor NOR4 (N4531, N4524, N3168, N3336, N2257);
nand NAND3 (N4532, N4530, N2749, N767);
and AND3 (N4533, N4522, N87, N1042);
not NOT1 (N4534, N4516);
buf BUF1 (N4535, N4527);
and AND3 (N4536, N4531, N2161, N1677);
nor NOR2 (N4537, N4536, N192);
not NOT1 (N4538, N4537);
or OR4 (N4539, N4529, N2430, N1095, N4424);
nor NOR3 (N4540, N4539, N1472, N1953);
xor XOR2 (N4541, N4532, N2268);
xor XOR2 (N4542, N4538, N2457);
not NOT1 (N4543, N4540);
nand NAND3 (N4544, N4542, N997, N2103);
nor NOR4 (N4545, N4518, N2422, N1042, N994);
or OR2 (N4546, N4502, N467);
and AND4 (N4547, N4544, N4446, N1221, N590);
nand NAND3 (N4548, N4547, N3284, N3605);
or OR3 (N4549, N4545, N1128, N4052);
buf BUF1 (N4550, N4535);
xor XOR2 (N4551, N4543, N1369);
and AND4 (N4552, N4548, N2267, N2141, N3310);
and AND2 (N4553, N4541, N2792);
nand NAND2 (N4554, N4513, N1476);
buf BUF1 (N4555, N4546);
nor NOR3 (N4556, N4533, N1696, N1350);
xor XOR2 (N4557, N4552, N455);
or OR3 (N4558, N4551, N2923, N1602);
xor XOR2 (N4559, N4556, N2745);
or OR2 (N4560, N4557, N3857);
and AND2 (N4561, N4528, N3528);
xor XOR2 (N4562, N4559, N317);
or OR4 (N4563, N4549, N3924, N1560, N41);
and AND2 (N4564, N4558, N1923);
buf BUF1 (N4565, N4550);
or OR4 (N4566, N4534, N3610, N2258, N75);
nor NOR4 (N4567, N4562, N4006, N3891, N2557);
nor NOR4 (N4568, N4555, N3395, N1152, N3185);
xor XOR2 (N4569, N4560, N38);
nand NAND4 (N4570, N4554, N4047, N1162, N2690);
xor XOR2 (N4571, N4570, N1313);
and AND4 (N4572, N4568, N870, N2352, N4253);
not NOT1 (N4573, N4565);
and AND3 (N4574, N4566, N3202, N1924);
xor XOR2 (N4575, N4571, N3017);
nor NOR4 (N4576, N4575, N2125, N52, N368);
buf BUF1 (N4577, N4576);
nor NOR4 (N4578, N4564, N73, N47, N1583);
buf BUF1 (N4579, N4569);
nand NAND3 (N4580, N4574, N2908, N3509);
xor XOR2 (N4581, N4563, N2800);
xor XOR2 (N4582, N4573, N2715);
not NOT1 (N4583, N4581);
nand NAND3 (N4584, N4583, N3185, N2280);
and AND4 (N4585, N4584, N1760, N172, N3970);
and AND2 (N4586, N4578, N1209);
and AND3 (N4587, N4561, N2783, N2859);
or OR2 (N4588, N4567, N2060);
nor NOR4 (N4589, N4553, N3683, N3084, N4223);
buf BUF1 (N4590, N4572);
nand NAND3 (N4591, N4589, N3916, N219);
nor NOR3 (N4592, N4579, N437, N1392);
xor XOR2 (N4593, N4592, N3598);
and AND2 (N4594, N4588, N1186);
nor NOR4 (N4595, N4594, N46, N3617, N1442);
or OR3 (N4596, N4593, N101, N1472);
nor NOR2 (N4597, N4591, N58);
nand NAND3 (N4598, N4595, N1858, N1899);
not NOT1 (N4599, N4585);
xor XOR2 (N4600, N4586, N3048);
not NOT1 (N4601, N4599);
buf BUF1 (N4602, N4587);
xor XOR2 (N4603, N4602, N1486);
nand NAND3 (N4604, N4582, N2290, N2696);
not NOT1 (N4605, N4596);
nand NAND4 (N4606, N4604, N2266, N907, N1443);
nand NAND4 (N4607, N4597, N2225, N4434, N3101);
xor XOR2 (N4608, N4605, N289);
buf BUF1 (N4609, N4590);
buf BUF1 (N4610, N4607);
buf BUF1 (N4611, N4610);
or OR3 (N4612, N4598, N3283, N1549);
not NOT1 (N4613, N4601);
buf BUF1 (N4614, N4606);
nand NAND4 (N4615, N4612, N1194, N556, N3959);
or OR4 (N4616, N4600, N2563, N3600, N2427);
nor NOR2 (N4617, N4577, N1022);
buf BUF1 (N4618, N4608);
xor XOR2 (N4619, N4609, N85);
or OR2 (N4620, N4613, N640);
xor XOR2 (N4621, N4603, N1254);
nor NOR4 (N4622, N4616, N1447, N2376, N3134);
or OR3 (N4623, N4611, N3001, N2339);
and AND3 (N4624, N4614, N1058, N163);
xor XOR2 (N4625, N4622, N1513);
and AND4 (N4626, N4617, N108, N2891, N1795);
xor XOR2 (N4627, N4580, N59);
not NOT1 (N4628, N4623);
xor XOR2 (N4629, N4626, N3718);
xor XOR2 (N4630, N4615, N703);
nor NOR4 (N4631, N4621, N3149, N390, N2289);
buf BUF1 (N4632, N4627);
not NOT1 (N4633, N4628);
nand NAND4 (N4634, N4618, N3680, N3121, N4271);
or OR3 (N4635, N4624, N697, N3556);
not NOT1 (N4636, N4629);
xor XOR2 (N4637, N4619, N505);
xor XOR2 (N4638, N4632, N1096);
nand NAND2 (N4639, N4638, N3658);
not NOT1 (N4640, N4630);
or OR2 (N4641, N4637, N4198);
nand NAND2 (N4642, N4641, N646);
nor NOR4 (N4643, N4640, N3362, N2668, N2710);
not NOT1 (N4644, N4633);
nand NAND4 (N4645, N4643, N213, N3851, N169);
or OR2 (N4646, N4635, N2416);
buf BUF1 (N4647, N4639);
nor NOR4 (N4648, N4645, N2640, N476, N4005);
buf BUF1 (N4649, N4644);
nor NOR4 (N4650, N4631, N2796, N484, N3362);
nor NOR4 (N4651, N4648, N2722, N3623, N3900);
nor NOR4 (N4652, N4651, N2139, N2173, N3063);
not NOT1 (N4653, N4646);
nand NAND3 (N4654, N4652, N3327, N4120);
not NOT1 (N4655, N4636);
xor XOR2 (N4656, N4620, N994);
buf BUF1 (N4657, N4625);
nor NOR2 (N4658, N4634, N1111);
and AND3 (N4659, N4647, N1832, N2708);
nand NAND2 (N4660, N4657, N3150);
nand NAND2 (N4661, N4653, N2639);
or OR3 (N4662, N4655, N3880, N1269);
and AND2 (N4663, N4661, N142);
xor XOR2 (N4664, N4660, N1605);
buf BUF1 (N4665, N4659);
or OR2 (N4666, N4664, N3588);
xor XOR2 (N4667, N4658, N2217);
or OR4 (N4668, N4667, N27, N1909, N3921);
nand NAND2 (N4669, N4642, N1577);
xor XOR2 (N4670, N4663, N1179);
xor XOR2 (N4671, N4650, N1716);
and AND3 (N4672, N4670, N396, N1648);
nand NAND3 (N4673, N4666, N3625, N3960);
buf BUF1 (N4674, N4668);
xor XOR2 (N4675, N4665, N1444);
not NOT1 (N4676, N4662);
nand NAND3 (N4677, N4671, N3021, N351);
not NOT1 (N4678, N4675);
buf BUF1 (N4679, N4677);
nand NAND3 (N4680, N4676, N678, N604);
buf BUF1 (N4681, N4669);
nor NOR2 (N4682, N4674, N4041);
xor XOR2 (N4683, N4673, N2226);
and AND3 (N4684, N4681, N561, N4069);
and AND3 (N4685, N4680, N3736, N99);
and AND4 (N4686, N4654, N1239, N2370, N2458);
xor XOR2 (N4687, N4679, N4433);
buf BUF1 (N4688, N4683);
nand NAND3 (N4689, N4649, N2914, N3789);
and AND4 (N4690, N4687, N3147, N4065, N711);
and AND4 (N4691, N4672, N3244, N1901, N1870);
buf BUF1 (N4692, N4686);
xor XOR2 (N4693, N4684, N3632);
or OR4 (N4694, N4692, N3545, N672, N2733);
xor XOR2 (N4695, N4656, N2849);
and AND2 (N4696, N4682, N4189);
and AND4 (N4697, N4690, N777, N2384, N458);
xor XOR2 (N4698, N4694, N2325);
nor NOR3 (N4699, N4695, N2604, N1181);
nand NAND2 (N4700, N4685, N3567);
and AND4 (N4701, N4698, N1405, N2300, N4066);
buf BUF1 (N4702, N4696);
nand NAND4 (N4703, N4700, N3164, N3231, N424);
buf BUF1 (N4704, N4703);
nand NAND2 (N4705, N4688, N1259);
xor XOR2 (N4706, N4701, N2645);
xor XOR2 (N4707, N4697, N4028);
and AND2 (N4708, N4689, N4447);
buf BUF1 (N4709, N4678);
nor NOR4 (N4710, N4702, N3916, N555, N328);
or OR4 (N4711, N4691, N329, N2891, N3586);
nand NAND3 (N4712, N4699, N3626, N998);
xor XOR2 (N4713, N4705, N2615);
buf BUF1 (N4714, N4704);
nor NOR3 (N4715, N4714, N1761, N4252);
xor XOR2 (N4716, N4706, N2618);
nor NOR3 (N4717, N4707, N724, N2978);
not NOT1 (N4718, N4711);
or OR2 (N4719, N4708, N4639);
nor NOR3 (N4720, N4693, N453, N2327);
or OR3 (N4721, N4718, N1443, N3324);
nor NOR2 (N4722, N4720, N3243);
or OR4 (N4723, N4710, N1804, N352, N1200);
nor NOR2 (N4724, N4722, N4055);
xor XOR2 (N4725, N4724, N1362);
nand NAND4 (N4726, N4709, N3631, N36, N2557);
nor NOR2 (N4727, N4712, N3041);
nand NAND2 (N4728, N4723, N552);
nor NOR3 (N4729, N4715, N92, N2497);
or OR4 (N4730, N4721, N4482, N1479, N2835);
or OR2 (N4731, N4719, N196);
nor NOR2 (N4732, N4728, N1753);
nor NOR4 (N4733, N4730, N55, N1926, N2365);
or OR2 (N4734, N4733, N1836);
buf BUF1 (N4735, N4717);
nor NOR2 (N4736, N4731, N829);
nor NOR4 (N4737, N4735, N4589, N792, N2526);
xor XOR2 (N4738, N4729, N1934);
and AND2 (N4739, N4736, N3977);
or OR4 (N4740, N4713, N2188, N2474, N1955);
and AND4 (N4741, N4727, N4150, N2691, N4266);
nand NAND3 (N4742, N4732, N2778, N1256);
xor XOR2 (N4743, N4734, N734);
and AND3 (N4744, N4737, N2150, N1703);
nand NAND4 (N4745, N4716, N4284, N671, N4322);
buf BUF1 (N4746, N4745);
nor NOR2 (N4747, N4726, N2562);
nand NAND3 (N4748, N4747, N2803, N644);
not NOT1 (N4749, N4743);
not NOT1 (N4750, N4741);
nor NOR4 (N4751, N4746, N1948, N3110, N2962);
or OR2 (N4752, N4750, N4679);
buf BUF1 (N4753, N4739);
xor XOR2 (N4754, N4744, N4207);
nor NOR3 (N4755, N4748, N572, N723);
xor XOR2 (N4756, N4753, N3451);
and AND2 (N4757, N4752, N1414);
buf BUF1 (N4758, N4749);
not NOT1 (N4759, N4751);
nand NAND3 (N4760, N4756, N2513, N3341);
and AND4 (N4761, N4760, N2185, N42, N1254);
not NOT1 (N4762, N4761);
and AND2 (N4763, N4759, N1902);
or OR2 (N4764, N4762, N3839);
nand NAND3 (N4765, N4742, N3568, N3718);
nor NOR4 (N4766, N4755, N1632, N1586, N90);
buf BUF1 (N4767, N4763);
buf BUF1 (N4768, N4766);
buf BUF1 (N4769, N4738);
buf BUF1 (N4770, N4764);
and AND3 (N4771, N4767, N2646, N2873);
buf BUF1 (N4772, N4770);
nor NOR4 (N4773, N4769, N4299, N1435, N3622);
nand NAND4 (N4774, N4765, N2815, N2860, N3420);
nand NAND4 (N4775, N4768, N1077, N1619, N956);
nor NOR4 (N4776, N4740, N2062, N4374, N2205);
nand NAND4 (N4777, N4771, N933, N3666, N4519);
nand NAND2 (N4778, N4774, N2536);
not NOT1 (N4779, N4775);
nand NAND2 (N4780, N4754, N1524);
xor XOR2 (N4781, N4776, N2190);
buf BUF1 (N4782, N4781);
not NOT1 (N4783, N4773);
xor XOR2 (N4784, N4780, N3043);
nor NOR2 (N4785, N4758, N4729);
xor XOR2 (N4786, N4784, N2719);
buf BUF1 (N4787, N4786);
buf BUF1 (N4788, N4787);
or OR2 (N4789, N4785, N709);
xor XOR2 (N4790, N4725, N3834);
and AND2 (N4791, N4777, N4095);
or OR3 (N4792, N4788, N691, N2519);
and AND2 (N4793, N4772, N3423);
or OR4 (N4794, N4778, N3808, N1284, N1179);
not NOT1 (N4795, N4791);
nand NAND4 (N4796, N4792, N1625, N4123, N1968);
and AND4 (N4797, N4796, N4022, N1654, N1897);
and AND4 (N4798, N4779, N2824, N936, N4394);
buf BUF1 (N4799, N4789);
buf BUF1 (N4800, N4795);
or OR4 (N4801, N4800, N735, N1430, N610);
nor NOR2 (N4802, N4757, N2924);
not NOT1 (N4803, N4790);
nor NOR2 (N4804, N4801, N135);
or OR3 (N4805, N4803, N3324, N4655);
or OR4 (N4806, N4782, N1224, N4628, N4693);
or OR4 (N4807, N4783, N3300, N824, N4319);
buf BUF1 (N4808, N4798);
and AND4 (N4809, N4805, N2152, N2870, N3684);
nor NOR3 (N4810, N4804, N818, N1123);
nand NAND4 (N4811, N4797, N4599, N1324, N496);
nor NOR2 (N4812, N4806, N4097);
buf BUF1 (N4813, N4794);
not NOT1 (N4814, N4802);
xor XOR2 (N4815, N4810, N4497);
xor XOR2 (N4816, N4809, N2824);
and AND3 (N4817, N4793, N4089, N1605);
buf BUF1 (N4818, N4813);
nand NAND3 (N4819, N4799, N3633, N2435);
xor XOR2 (N4820, N4816, N450);
not NOT1 (N4821, N4814);
nand NAND2 (N4822, N4821, N3369);
not NOT1 (N4823, N4812);
buf BUF1 (N4824, N4823);
not NOT1 (N4825, N4818);
xor XOR2 (N4826, N4815, N3003);
or OR2 (N4827, N4808, N380);
nor NOR4 (N4828, N4817, N4706, N1297, N4603);
buf BUF1 (N4829, N4828);
not NOT1 (N4830, N4826);
buf BUF1 (N4831, N4825);
not NOT1 (N4832, N4827);
or OR2 (N4833, N4811, N4626);
not NOT1 (N4834, N4822);
not NOT1 (N4835, N4829);
and AND4 (N4836, N4831, N3295, N3540, N2511);
nor NOR4 (N4837, N4807, N2117, N2688, N2399);
not NOT1 (N4838, N4836);
nor NOR4 (N4839, N4833, N2491, N823, N3453);
xor XOR2 (N4840, N4838, N98);
and AND3 (N4841, N4837, N1175, N2506);
and AND2 (N4842, N4840, N3295);
not NOT1 (N4843, N4834);
not NOT1 (N4844, N4835);
and AND3 (N4845, N4844, N4298, N3185);
buf BUF1 (N4846, N4819);
buf BUF1 (N4847, N4820);
and AND2 (N4848, N4846, N3187);
nand NAND2 (N4849, N4845, N2081);
and AND3 (N4850, N4824, N4430, N2408);
xor XOR2 (N4851, N4842, N4363);
xor XOR2 (N4852, N4841, N3180);
buf BUF1 (N4853, N4843);
or OR3 (N4854, N4839, N2128, N4458);
buf BUF1 (N4855, N4851);
buf BUF1 (N4856, N4848);
not NOT1 (N4857, N4850);
xor XOR2 (N4858, N4852, N3749);
and AND3 (N4859, N4853, N985, N3998);
buf BUF1 (N4860, N4849);
or OR2 (N4861, N4830, N2085);
or OR4 (N4862, N4858, N3616, N3423, N3852);
nand NAND3 (N4863, N4855, N4354, N2625);
nand NAND2 (N4864, N4860, N577);
nor NOR2 (N4865, N4832, N498);
xor XOR2 (N4866, N4859, N4267);
xor XOR2 (N4867, N4861, N1764);
nand NAND3 (N4868, N4847, N2281, N672);
and AND3 (N4869, N4862, N4812, N892);
not NOT1 (N4870, N4854);
buf BUF1 (N4871, N4870);
not NOT1 (N4872, N4871);
xor XOR2 (N4873, N4865, N1440);
nor NOR4 (N4874, N4867, N1162, N1630, N1363);
xor XOR2 (N4875, N4856, N3697);
or OR2 (N4876, N4869, N3823);
or OR2 (N4877, N4876, N4077);
nand NAND2 (N4878, N4866, N3375);
not NOT1 (N4879, N4863);
not NOT1 (N4880, N4879);
buf BUF1 (N4881, N4864);
not NOT1 (N4882, N4881);
nor NOR4 (N4883, N4880, N1903, N3246, N2762);
or OR3 (N4884, N4875, N3329, N2137);
not NOT1 (N4885, N4883);
buf BUF1 (N4886, N4874);
not NOT1 (N4887, N4884);
buf BUF1 (N4888, N4885);
and AND2 (N4889, N4887, N1405);
and AND4 (N4890, N4886, N2762, N185, N2581);
and AND3 (N4891, N4878, N2357, N2518);
xor XOR2 (N4892, N4877, N3851);
xor XOR2 (N4893, N4868, N3984);
and AND3 (N4894, N4889, N2366, N3950);
buf BUF1 (N4895, N4882);
and AND2 (N4896, N4890, N2455);
or OR3 (N4897, N4872, N2805, N2158);
buf BUF1 (N4898, N4888);
buf BUF1 (N4899, N4896);
xor XOR2 (N4900, N4873, N2311);
and AND3 (N4901, N4897, N2733, N4452);
and AND3 (N4902, N4901, N1565, N428);
and AND3 (N4903, N4892, N2320, N321);
and AND3 (N4904, N4898, N1533, N2707);
or OR3 (N4905, N4893, N1097, N2629);
nor NOR4 (N4906, N4902, N3973, N1562, N983);
xor XOR2 (N4907, N4905, N971);
nand NAND4 (N4908, N4857, N2887, N793, N1478);
nand NAND4 (N4909, N4899, N212, N2985, N233);
buf BUF1 (N4910, N4895);
buf BUF1 (N4911, N4906);
xor XOR2 (N4912, N4900, N1321);
nor NOR4 (N4913, N4904, N4606, N4850, N2436);
and AND4 (N4914, N4913, N3020, N2823, N4444);
and AND2 (N4915, N4910, N2877);
buf BUF1 (N4916, N4911);
nand NAND2 (N4917, N4912, N3557);
or OR2 (N4918, N4917, N3300);
or OR4 (N4919, N4916, N111, N3096, N3845);
and AND2 (N4920, N4891, N1100);
nor NOR2 (N4921, N4915, N2163);
not NOT1 (N4922, N4918);
nor NOR4 (N4923, N4908, N3298, N4338, N3617);
buf BUF1 (N4924, N4921);
or OR2 (N4925, N4914, N3033);
and AND3 (N4926, N4920, N1321, N1648);
xor XOR2 (N4927, N4919, N2030);
buf BUF1 (N4928, N4923);
xor XOR2 (N4929, N4928, N1772);
not NOT1 (N4930, N4894);
xor XOR2 (N4931, N4930, N1508);
xor XOR2 (N4932, N4929, N4048);
and AND3 (N4933, N4932, N345, N399);
or OR4 (N4934, N4926, N2236, N4749, N2161);
nor NOR4 (N4935, N4909, N4053, N521, N1362);
nor NOR4 (N4936, N4931, N800, N3615, N1808);
buf BUF1 (N4937, N4933);
and AND2 (N4938, N4907, N3558);
xor XOR2 (N4939, N4938, N4759);
and AND2 (N4940, N4925, N871);
or OR4 (N4941, N4922, N1942, N4020, N220);
not NOT1 (N4942, N4903);
or OR3 (N4943, N4939, N1318, N4182);
xor XOR2 (N4944, N4940, N3656);
nand NAND4 (N4945, N4927, N3175, N3313, N2900);
xor XOR2 (N4946, N4924, N4561);
or OR2 (N4947, N4935, N1820);
nor NOR2 (N4948, N4943, N1137);
and AND4 (N4949, N4934, N4519, N579, N1002);
buf BUF1 (N4950, N4937);
buf BUF1 (N4951, N4944);
nand NAND4 (N4952, N4950, N2979, N2282, N4862);
nor NOR3 (N4953, N4952, N1620, N1306);
buf BUF1 (N4954, N4947);
not NOT1 (N4955, N4936);
buf BUF1 (N4956, N4941);
nor NOR4 (N4957, N4948, N2268, N1052, N1919);
and AND4 (N4958, N4954, N610, N1693, N4195);
and AND2 (N4959, N4958, N724);
or OR4 (N4960, N4959, N3248, N3396, N4104);
or OR2 (N4961, N4942, N903);
buf BUF1 (N4962, N4945);
buf BUF1 (N4963, N4951);
xor XOR2 (N4964, N4961, N3524);
and AND3 (N4965, N4956, N2568, N1684);
not NOT1 (N4966, N4949);
nand NAND4 (N4967, N4964, N4098, N35, N2632);
nor NOR3 (N4968, N4955, N716, N1036);
buf BUF1 (N4969, N4962);
or OR4 (N4970, N4967, N4235, N3914, N416);
nor NOR3 (N4971, N4960, N4864, N2598);
buf BUF1 (N4972, N4966);
not NOT1 (N4973, N4969);
or OR3 (N4974, N4970, N4575, N1016);
not NOT1 (N4975, N4963);
and AND2 (N4976, N4953, N1193);
nor NOR2 (N4977, N4974, N2687);
nand NAND3 (N4978, N4957, N154, N4819);
nand NAND3 (N4979, N4977, N3982, N4072);
or OR2 (N4980, N4972, N2903);
xor XOR2 (N4981, N4968, N1405);
not NOT1 (N4982, N4973);
and AND4 (N4983, N4978, N989, N1936, N2374);
or OR3 (N4984, N4965, N1714, N3853);
and AND4 (N4985, N4983, N2482, N1387, N968);
and AND4 (N4986, N4985, N2546, N2478, N2826);
not NOT1 (N4987, N4986);
buf BUF1 (N4988, N4975);
xor XOR2 (N4989, N4979, N871);
or OR4 (N4990, N4984, N2061, N1260, N695);
or OR3 (N4991, N4990, N1524, N4106);
and AND2 (N4992, N4982, N4916);
and AND3 (N4993, N4946, N2298, N2578);
xor XOR2 (N4994, N4988, N2738);
xor XOR2 (N4995, N4981, N3202);
or OR3 (N4996, N4976, N3803, N371);
not NOT1 (N4997, N4971);
buf BUF1 (N4998, N4995);
nand NAND4 (N4999, N4997, N656, N54, N4954);
and AND4 (N5000, N4998, N4395, N4214, N2257);
or OR4 (N5001, N4991, N624, N2723, N1317);
xor XOR2 (N5002, N4980, N2876);
nand NAND4 (N5003, N4989, N1730, N3394, N134);
buf BUF1 (N5004, N4992);
nor NOR2 (N5005, N5001, N1579);
nand NAND4 (N5006, N4993, N558, N2409, N4877);
xor XOR2 (N5007, N4999, N2445);
and AND2 (N5008, N5002, N1642);
nor NOR3 (N5009, N5005, N1321, N883);
nand NAND2 (N5010, N5009, N4874);
xor XOR2 (N5011, N4987, N2982);
nand NAND3 (N5012, N5003, N4858, N1076);
and AND3 (N5013, N5007, N525, N4067);
xor XOR2 (N5014, N4996, N3995);
xor XOR2 (N5015, N5014, N1437);
buf BUF1 (N5016, N4994);
or OR4 (N5017, N5000, N4165, N879, N4625);
and AND3 (N5018, N5006, N1331, N970);
nand NAND3 (N5019, N5017, N258, N4323);
nor NOR3 (N5020, N5004, N1325, N2415);
and AND4 (N5021, N5016, N1823, N500, N1441);
and AND3 (N5022, N5011, N588, N910);
and AND4 (N5023, N5020, N2099, N2112, N1940);
buf BUF1 (N5024, N5023);
buf BUF1 (N5025, N5024);
xor XOR2 (N5026, N5019, N546);
not NOT1 (N5027, N5022);
nand NAND2 (N5028, N5018, N4838);
not NOT1 (N5029, N5026);
and AND3 (N5030, N5028, N2714, N4335);
nand NAND4 (N5031, N5008, N956, N3002, N489);
or OR4 (N5032, N5027, N1434, N1159, N4114);
or OR4 (N5033, N5013, N2006, N659, N2629);
xor XOR2 (N5034, N5010, N2243);
nor NOR3 (N5035, N5025, N3955, N102);
nand NAND4 (N5036, N5012, N2217, N2774, N4740);
and AND4 (N5037, N5031, N4901, N297, N2987);
xor XOR2 (N5038, N5034, N102);
or OR4 (N5039, N5036, N3908, N4340, N2222);
nor NOR4 (N5040, N5032, N3257, N667, N521);
nand NAND2 (N5041, N5035, N1146);
nand NAND2 (N5042, N5033, N409);
and AND4 (N5043, N5042, N3795, N470, N1378);
nand NAND2 (N5044, N5015, N4323);
or OR2 (N5045, N5039, N2539);
and AND2 (N5046, N5030, N4407);
xor XOR2 (N5047, N5021, N421);
not NOT1 (N5048, N5046);
buf BUF1 (N5049, N5047);
buf BUF1 (N5050, N5029);
not NOT1 (N5051, N5048);
nor NOR4 (N5052, N5045, N4096, N543, N1600);
and AND3 (N5053, N5043, N937, N448);
and AND2 (N5054, N5038, N217);
and AND3 (N5055, N5040, N4448, N3873);
or OR4 (N5056, N5041, N1380, N2000, N2673);
xor XOR2 (N5057, N5051, N4880);
or OR3 (N5058, N5052, N4175, N5045);
or OR3 (N5059, N5055, N149, N1391);
nand NAND2 (N5060, N5056, N4403);
nor NOR3 (N5061, N5044, N609, N4443);
not NOT1 (N5062, N5050);
nor NOR4 (N5063, N5062, N294, N3018, N3063);
nor NOR3 (N5064, N5058, N4021, N541);
nor NOR2 (N5065, N5059, N3604);
buf BUF1 (N5066, N5060);
buf BUF1 (N5067, N5049);
not NOT1 (N5068, N5061);
nor NOR4 (N5069, N5057, N3324, N4231, N1598);
buf BUF1 (N5070, N5069);
xor XOR2 (N5071, N5054, N122);
and AND3 (N5072, N5065, N1848, N4864);
xor XOR2 (N5073, N5067, N588);
nor NOR3 (N5074, N5063, N3907, N2087);
nor NOR2 (N5075, N5068, N1335);
not NOT1 (N5076, N5072);
or OR4 (N5077, N5075, N2481, N680, N2813);
and AND4 (N5078, N5077, N5045, N311, N5046);
not NOT1 (N5079, N5053);
nor NOR3 (N5080, N5071, N2556, N757);
buf BUF1 (N5081, N5074);
and AND4 (N5082, N5064, N4603, N1197, N4134);
buf BUF1 (N5083, N5076);
nor NOR2 (N5084, N5073, N2656);
buf BUF1 (N5085, N5084);
and AND4 (N5086, N5079, N1894, N29, N1400);
and AND4 (N5087, N5078, N3312, N3912, N4087);
and AND3 (N5088, N5086, N4811, N4871);
or OR3 (N5089, N5087, N2354, N1185);
buf BUF1 (N5090, N5070);
not NOT1 (N5091, N5081);
xor XOR2 (N5092, N5082, N4710);
nand NAND3 (N5093, N5037, N3139, N1635);
not NOT1 (N5094, N5088);
nor NOR4 (N5095, N5080, N4169, N1459, N4422);
xor XOR2 (N5096, N5095, N2665);
and AND3 (N5097, N5092, N4247, N1962);
xor XOR2 (N5098, N5066, N2304);
xor XOR2 (N5099, N5093, N2055);
xor XOR2 (N5100, N5098, N2640);
and AND4 (N5101, N5089, N4847, N4960, N1951);
or OR3 (N5102, N5101, N935, N1472);
buf BUF1 (N5103, N5085);
nand NAND4 (N5104, N5099, N1106, N2996, N2714);
xor XOR2 (N5105, N5100, N3848);
not NOT1 (N5106, N5102);
nor NOR4 (N5107, N5096, N4977, N4696, N501);
or OR2 (N5108, N5091, N4360);
nor NOR2 (N5109, N5090, N1974);
nor NOR4 (N5110, N5104, N2261, N944, N2142);
and AND3 (N5111, N5105, N1507, N1894);
or OR2 (N5112, N5108, N768);
nand NAND3 (N5113, N5083, N4865, N3268);
xor XOR2 (N5114, N5112, N4186);
or OR2 (N5115, N5097, N1247);
nor NOR4 (N5116, N5109, N2554, N2516, N2288);
nand NAND3 (N5117, N5107, N1740, N4598);
nor NOR2 (N5118, N5117, N3210);
not NOT1 (N5119, N5118);
or OR3 (N5120, N5114, N1620, N2858);
nor NOR4 (N5121, N5106, N4091, N870, N4198);
nand NAND4 (N5122, N5120, N4295, N741, N779);
buf BUF1 (N5123, N5111);
buf BUF1 (N5124, N5113);
nand NAND2 (N5125, N5123, N4304);
not NOT1 (N5126, N5094);
or OR4 (N5127, N5110, N1678, N2307, N1153);
not NOT1 (N5128, N5103);
buf BUF1 (N5129, N5116);
buf BUF1 (N5130, N5115);
or OR3 (N5131, N5129, N2490, N2196);
nor NOR3 (N5132, N5121, N3294, N3991);
and AND3 (N5133, N5127, N4423, N2167);
and AND4 (N5134, N5132, N4689, N3651, N454);
nor NOR3 (N5135, N5130, N4337, N3905);
buf BUF1 (N5136, N5125);
nor NOR3 (N5137, N5131, N2235, N2131);
and AND4 (N5138, N5122, N1415, N5128, N103);
not NOT1 (N5139, N618);
not NOT1 (N5140, N5136);
nor NOR3 (N5141, N5137, N4646, N1159);
nor NOR3 (N5142, N5134, N4547, N2806);
nand NAND4 (N5143, N5126, N1697, N924, N1223);
nand NAND2 (N5144, N5142, N1942);
or OR4 (N5145, N5133, N4851, N1355, N1203);
xor XOR2 (N5146, N5141, N1023);
buf BUF1 (N5147, N5119);
or OR2 (N5148, N5143, N1503);
and AND3 (N5149, N5138, N4339, N4580);
xor XOR2 (N5150, N5147, N3707);
xor XOR2 (N5151, N5145, N795);
nand NAND2 (N5152, N5150, N2709);
nand NAND4 (N5153, N5139, N916, N4779, N1061);
xor XOR2 (N5154, N5149, N4737);
and AND4 (N5155, N5144, N3243, N3717, N4124);
not NOT1 (N5156, N5135);
buf BUF1 (N5157, N5152);
buf BUF1 (N5158, N5157);
nand NAND2 (N5159, N5154, N3642);
nand NAND2 (N5160, N5124, N5079);
or OR2 (N5161, N5140, N663);
nor NOR4 (N5162, N5156, N5130, N2293, N669);
nor NOR4 (N5163, N5153, N4351, N4923, N3091);
and AND2 (N5164, N5151, N4);
buf BUF1 (N5165, N5164);
not NOT1 (N5166, N5158);
nand NAND2 (N5167, N5148, N1407);
nand NAND3 (N5168, N5163, N2740, N623);
buf BUF1 (N5169, N5165);
xor XOR2 (N5170, N5161, N3890);
nor NOR3 (N5171, N5155, N2535, N5128);
not NOT1 (N5172, N5167);
not NOT1 (N5173, N5168);
buf BUF1 (N5174, N5169);
not NOT1 (N5175, N5172);
buf BUF1 (N5176, N5160);
nor NOR2 (N5177, N5162, N2577);
buf BUF1 (N5178, N5159);
nor NOR3 (N5179, N5174, N2833, N4406);
or OR3 (N5180, N5175, N2543, N2579);
not NOT1 (N5181, N5170);
or OR3 (N5182, N5178, N2386, N3902);
nand NAND4 (N5183, N5180, N2631, N537, N1005);
nor NOR2 (N5184, N5182, N4966);
or OR2 (N5185, N5183, N485);
nor NOR2 (N5186, N5166, N4590);
buf BUF1 (N5187, N5184);
not NOT1 (N5188, N5177);
nand NAND4 (N5189, N5181, N4822, N1322, N2443);
and AND4 (N5190, N5187, N3083, N3301, N3678);
nor NOR3 (N5191, N5189, N4054, N3805);
nor NOR2 (N5192, N5186, N3551);
or OR4 (N5193, N5173, N573, N3514, N4486);
buf BUF1 (N5194, N5146);
nand NAND3 (N5195, N5193, N4604, N1621);
nand NAND3 (N5196, N5171, N2787, N4587);
xor XOR2 (N5197, N5192, N686);
xor XOR2 (N5198, N5185, N1767);
nor NOR2 (N5199, N5176, N4224);
buf BUF1 (N5200, N5196);
nor NOR3 (N5201, N5200, N3179, N2555);
or OR4 (N5202, N5179, N855, N2591, N5070);
and AND3 (N5203, N5195, N3430, N1212);
nor NOR3 (N5204, N5194, N2180, N4736);
nor NOR3 (N5205, N5201, N2678, N2332);
nor NOR2 (N5206, N5199, N180);
and AND3 (N5207, N5205, N989, N2749);
buf BUF1 (N5208, N5207);
not NOT1 (N5209, N5190);
and AND2 (N5210, N5198, N4519);
not NOT1 (N5211, N5197);
or OR2 (N5212, N5191, N2739);
not NOT1 (N5213, N5206);
nand NAND2 (N5214, N5212, N2739);
nand NAND3 (N5215, N5203, N3360, N3645);
nor NOR2 (N5216, N5208, N3176);
buf BUF1 (N5217, N5211);
or OR2 (N5218, N5213, N1074);
nor NOR2 (N5219, N5214, N2242);
or OR3 (N5220, N5210, N357, N1433);
and AND3 (N5221, N5219, N3321, N887);
or OR4 (N5222, N5217, N34, N3276, N4138);
nand NAND3 (N5223, N5222, N715, N3024);
or OR2 (N5224, N5204, N2481);
and AND2 (N5225, N5218, N1985);
xor XOR2 (N5226, N5209, N2070);
or OR3 (N5227, N5188, N1786, N4174);
nand NAND2 (N5228, N5226, N2149);
xor XOR2 (N5229, N5216, N3310);
nor NOR4 (N5230, N5220, N1429, N6, N2857);
buf BUF1 (N5231, N5215);
nand NAND4 (N5232, N5202, N3168, N1856, N2020);
xor XOR2 (N5233, N5230, N3960);
and AND4 (N5234, N5225, N3397, N10, N4464);
and AND3 (N5235, N5234, N464, N4932);
nor NOR2 (N5236, N5221, N1867);
and AND4 (N5237, N5223, N372, N1217, N1713);
xor XOR2 (N5238, N5228, N2546);
buf BUF1 (N5239, N5227);
and AND2 (N5240, N5235, N1610);
xor XOR2 (N5241, N5224, N1393);
nand NAND4 (N5242, N5241, N1271, N3649, N4262);
xor XOR2 (N5243, N5239, N4098);
xor XOR2 (N5244, N5236, N1708);
nor NOR4 (N5245, N5229, N3968, N1992, N914);
nand NAND4 (N5246, N5237, N4533, N340, N3449);
nand NAND3 (N5247, N5233, N551, N3598);
and AND4 (N5248, N5243, N2651, N2242, N3081);
not NOT1 (N5249, N5238);
nand NAND4 (N5250, N5242, N957, N5075, N2729);
nor NOR2 (N5251, N5240, N197);
nor NOR2 (N5252, N5246, N5180);
nor NOR2 (N5253, N5245, N2637);
not NOT1 (N5254, N5250);
not NOT1 (N5255, N5231);
or OR4 (N5256, N5252, N2936, N3116, N867);
xor XOR2 (N5257, N5251, N4444);
nor NOR3 (N5258, N5248, N3882, N5014);
buf BUF1 (N5259, N5249);
and AND3 (N5260, N5258, N2739, N2530);
not NOT1 (N5261, N5232);
buf BUF1 (N5262, N5256);
or OR4 (N5263, N5247, N2100, N4035, N2136);
xor XOR2 (N5264, N5257, N4620);
buf BUF1 (N5265, N5264);
nor NOR3 (N5266, N5265, N2703, N1531);
buf BUF1 (N5267, N5260);
nand NAND2 (N5268, N5244, N4106);
and AND3 (N5269, N5261, N927, N3007);
not NOT1 (N5270, N5269);
buf BUF1 (N5271, N5259);
or OR4 (N5272, N5255, N4532, N2649, N1573);
buf BUF1 (N5273, N5262);
or OR4 (N5274, N5271, N4808, N1789, N708);
buf BUF1 (N5275, N5267);
xor XOR2 (N5276, N5270, N2265);
nand NAND2 (N5277, N5272, N4386);
xor XOR2 (N5278, N5275, N3301);
nand NAND3 (N5279, N5277, N1131, N3185);
or OR4 (N5280, N5263, N2413, N3549, N978);
nor NOR4 (N5281, N5280, N752, N2253, N2973);
xor XOR2 (N5282, N5253, N4310);
buf BUF1 (N5283, N5254);
xor XOR2 (N5284, N5283, N3063);
nand NAND2 (N5285, N5266, N2689);
nand NAND4 (N5286, N5274, N3780, N3488, N2573);
or OR2 (N5287, N5282, N2829);
and AND4 (N5288, N5279, N751, N5086, N382);
buf BUF1 (N5289, N5288);
and AND2 (N5290, N5289, N2626);
xor XOR2 (N5291, N5268, N2003);
or OR4 (N5292, N5281, N1915, N4452, N3267);
or OR2 (N5293, N5291, N4864);
or OR4 (N5294, N5278, N3523, N3243, N4247);
nor NOR4 (N5295, N5286, N2596, N3979, N3890);
xor XOR2 (N5296, N5290, N2774);
or OR3 (N5297, N5292, N2440, N4681);
xor XOR2 (N5298, N5284, N154);
and AND4 (N5299, N5293, N3151, N4597, N548);
nor NOR4 (N5300, N5294, N2336, N1398, N4719);
or OR2 (N5301, N5298, N5168);
buf BUF1 (N5302, N5297);
buf BUF1 (N5303, N5287);
xor XOR2 (N5304, N5302, N918);
not NOT1 (N5305, N5295);
xor XOR2 (N5306, N5276, N3869);
nand NAND3 (N5307, N5305, N3968, N4872);
nor NOR4 (N5308, N5273, N1685, N3815, N5135);
xor XOR2 (N5309, N5303, N4668);
xor XOR2 (N5310, N5300, N2142);
nor NOR4 (N5311, N5309, N5083, N2797, N4116);
nand NAND3 (N5312, N5311, N3222, N3792);
xor XOR2 (N5313, N5310, N725);
nor NOR4 (N5314, N5299, N706, N835, N4458);
or OR4 (N5315, N5301, N310, N3896, N1150);
nand NAND4 (N5316, N5314, N5287, N2728, N3799);
nand NAND2 (N5317, N5315, N3305);
or OR2 (N5318, N5296, N3583);
nor NOR4 (N5319, N5308, N1786, N1672, N1550);
and AND3 (N5320, N5307, N2960, N1091);
not NOT1 (N5321, N5320);
nor NOR2 (N5322, N5318, N4359);
xor XOR2 (N5323, N5312, N1114);
or OR2 (N5324, N5306, N4772);
nand NAND3 (N5325, N5304, N3033, N1667);
nor NOR4 (N5326, N5325, N2334, N2015, N216);
and AND2 (N5327, N5326, N4449);
buf BUF1 (N5328, N5322);
or OR2 (N5329, N5316, N4872);
xor XOR2 (N5330, N5321, N388);
not NOT1 (N5331, N5328);
or OR4 (N5332, N5285, N4134, N4451, N2699);
xor XOR2 (N5333, N5327, N1258);
nand NAND3 (N5334, N5329, N3285, N5054);
nand NAND3 (N5335, N5313, N4523, N918);
nand NAND2 (N5336, N5319, N4613);
or OR2 (N5337, N5331, N3980);
xor XOR2 (N5338, N5323, N1908);
xor XOR2 (N5339, N5333, N4978);
nand NAND2 (N5340, N5332, N1692);
nor NOR2 (N5341, N5330, N5090);
buf BUF1 (N5342, N5335);
not NOT1 (N5343, N5337);
and AND4 (N5344, N5343, N3556, N4240, N1904);
buf BUF1 (N5345, N5338);
nor NOR4 (N5346, N5342, N1394, N4082, N3775);
and AND4 (N5347, N5341, N4616, N5109, N2831);
nand NAND3 (N5348, N5346, N5058, N2192);
buf BUF1 (N5349, N5317);
xor XOR2 (N5350, N5349, N61);
xor XOR2 (N5351, N5350, N4673);
and AND3 (N5352, N5334, N1725, N29);
buf BUF1 (N5353, N5339);
nor NOR4 (N5354, N5336, N5021, N4682, N1560);
and AND4 (N5355, N5344, N592, N4480, N4327);
nor NOR2 (N5356, N5351, N2588);
buf BUF1 (N5357, N5355);
xor XOR2 (N5358, N5357, N2365);
nor NOR3 (N5359, N5352, N4287, N4963);
not NOT1 (N5360, N5345);
xor XOR2 (N5361, N5360, N5006);
or OR3 (N5362, N5324, N1521, N2614);
and AND2 (N5363, N5354, N3634);
buf BUF1 (N5364, N5348);
nand NAND2 (N5365, N5353, N4901);
nor NOR2 (N5366, N5362, N918);
xor XOR2 (N5367, N5365, N766);
nor NOR2 (N5368, N5347, N3912);
xor XOR2 (N5369, N5359, N3075);
xor XOR2 (N5370, N5363, N5288);
nand NAND4 (N5371, N5368, N5272, N3351, N1984);
nand NAND4 (N5372, N5371, N1571, N718, N2136);
buf BUF1 (N5373, N5367);
buf BUF1 (N5374, N5358);
buf BUF1 (N5375, N5374);
nor NOR2 (N5376, N5370, N4475);
and AND4 (N5377, N5340, N1929, N3676, N3071);
xor XOR2 (N5378, N5376, N798);
or OR4 (N5379, N5361, N2677, N825, N1850);
nand NAND4 (N5380, N5369, N332, N4401, N5235);
not NOT1 (N5381, N5375);
and AND4 (N5382, N5373, N2351, N5033, N1319);
and AND2 (N5383, N5356, N3444);
and AND4 (N5384, N5382, N966, N3318, N4531);
not NOT1 (N5385, N5380);
nand NAND3 (N5386, N5372, N1429, N1140);
and AND4 (N5387, N5366, N643, N4356, N4863);
buf BUF1 (N5388, N5386);
buf BUF1 (N5389, N5388);
nand NAND3 (N5390, N5384, N3465, N714);
nor NOR3 (N5391, N5364, N1368, N4474);
xor XOR2 (N5392, N5377, N5093);
not NOT1 (N5393, N5379);
nor NOR3 (N5394, N5391, N4982, N3073);
nor NOR4 (N5395, N5394, N2510, N1774, N3462);
not NOT1 (N5396, N5393);
xor XOR2 (N5397, N5396, N522);
or OR2 (N5398, N5392, N3333);
nor NOR2 (N5399, N5398, N3767);
nor NOR4 (N5400, N5397, N1851, N3240, N4574);
nor NOR4 (N5401, N5381, N3486, N5213, N3334);
buf BUF1 (N5402, N5395);
and AND2 (N5403, N5401, N1452);
or OR4 (N5404, N5400, N5396, N4185, N5183);
nor NOR2 (N5405, N5390, N1418);
not NOT1 (N5406, N5385);
xor XOR2 (N5407, N5403, N4281);
and AND2 (N5408, N5383, N1686);
or OR3 (N5409, N5387, N2452, N4720);
nor NOR4 (N5410, N5405, N4129, N3426, N550);
nor NOR3 (N5411, N5404, N4919, N2639);
and AND2 (N5412, N5378, N1654);
buf BUF1 (N5413, N5402);
or OR3 (N5414, N5408, N3320, N1644);
or OR3 (N5415, N5406, N4836, N3344);
or OR3 (N5416, N5389, N3355, N2683);
xor XOR2 (N5417, N5411, N2088);
nor NOR4 (N5418, N5409, N467, N1644, N4622);
nor NOR4 (N5419, N5415, N529, N3383, N2947);
xor XOR2 (N5420, N5418, N2081);
and AND2 (N5421, N5399, N5215);
not NOT1 (N5422, N5421);
buf BUF1 (N5423, N5407);
not NOT1 (N5424, N5416);
nor NOR2 (N5425, N5422, N1334);
buf BUF1 (N5426, N5413);
nand NAND4 (N5427, N5423, N2671, N4577, N1724);
or OR4 (N5428, N5426, N2564, N2063, N2696);
or OR3 (N5429, N5428, N3162, N5410);
and AND3 (N5430, N2784, N4857, N89);
buf BUF1 (N5431, N5424);
and AND2 (N5432, N5414, N120);
not NOT1 (N5433, N5425);
xor XOR2 (N5434, N5432, N313);
and AND4 (N5435, N5430, N1663, N1860, N4211);
nor NOR3 (N5436, N5433, N3467, N3274);
xor XOR2 (N5437, N5434, N571);
nand NAND3 (N5438, N5420, N3135, N1488);
and AND4 (N5439, N5412, N4759, N3120, N4454);
xor XOR2 (N5440, N5436, N4157);
buf BUF1 (N5441, N5427);
nand NAND4 (N5442, N5417, N2022, N5303, N911);
or OR3 (N5443, N5419, N3083, N542);
nor NOR2 (N5444, N5438, N590);
buf BUF1 (N5445, N5440);
xor XOR2 (N5446, N5445, N1884);
nand NAND3 (N5447, N5429, N2360, N865);
or OR2 (N5448, N5444, N558);
and AND4 (N5449, N5439, N1899, N3272, N4961);
nor NOR2 (N5450, N5443, N2726);
or OR4 (N5451, N5442, N1599, N2828, N1437);
not NOT1 (N5452, N5447);
and AND3 (N5453, N5431, N4749, N3391);
nand NAND4 (N5454, N5435, N2860, N2167, N240);
nand NAND3 (N5455, N5452, N1504, N407);
nor NOR2 (N5456, N5449, N3439);
xor XOR2 (N5457, N5454, N5298);
nand NAND4 (N5458, N5450, N1186, N15, N2476);
buf BUF1 (N5459, N5455);
nand NAND3 (N5460, N5453, N2507, N1393);
or OR2 (N5461, N5451, N3111);
nand NAND2 (N5462, N5458, N5153);
and AND2 (N5463, N5446, N4653);
nor NOR3 (N5464, N5463, N4633, N445);
and AND4 (N5465, N5457, N2671, N3839, N1700);
or OR3 (N5466, N5465, N1390, N508);
nor NOR2 (N5467, N5462, N3289);
not NOT1 (N5468, N5437);
and AND3 (N5469, N5466, N2761, N3105);
nand NAND4 (N5470, N5441, N3046, N1285, N532);
buf BUF1 (N5471, N5459);
nand NAND3 (N5472, N5469, N4915, N3847);
and AND3 (N5473, N5461, N290, N2814);
nor NOR4 (N5474, N5470, N2781, N2970, N3833);
not NOT1 (N5475, N5474);
not NOT1 (N5476, N5471);
not NOT1 (N5477, N5468);
nor NOR4 (N5478, N5464, N1872, N3660, N2002);
or OR2 (N5479, N5472, N4902);
not NOT1 (N5480, N5448);
and AND3 (N5481, N5460, N3078, N4741);
or OR2 (N5482, N5481, N1656);
and AND2 (N5483, N5482, N3777);
or OR2 (N5484, N5473, N5353);
nor NOR2 (N5485, N5478, N1231);
or OR2 (N5486, N5485, N2727);
and AND2 (N5487, N5479, N2451);
xor XOR2 (N5488, N5456, N1406);
xor XOR2 (N5489, N5477, N4494);
buf BUF1 (N5490, N5486);
not NOT1 (N5491, N5483);
nand NAND4 (N5492, N5488, N3806, N3388, N2304);
buf BUF1 (N5493, N5484);
not NOT1 (N5494, N5487);
buf BUF1 (N5495, N5492);
nor NOR2 (N5496, N5491, N126);
xor XOR2 (N5497, N5475, N5110);
and AND3 (N5498, N5494, N2570, N3039);
nand NAND4 (N5499, N5476, N1365, N1387, N3005);
xor XOR2 (N5500, N5489, N3610);
nor NOR2 (N5501, N5467, N1096);
nand NAND2 (N5502, N5500, N1360);
buf BUF1 (N5503, N5493);
not NOT1 (N5504, N5497);
and AND3 (N5505, N5490, N3644, N2569);
nor NOR3 (N5506, N5504, N1832, N1652);
buf BUF1 (N5507, N5499);
nand NAND3 (N5508, N5503, N3096, N1570);
not NOT1 (N5509, N5508);
nand NAND3 (N5510, N5498, N3902, N2634);
buf BUF1 (N5511, N5501);
and AND3 (N5512, N5511, N2981, N3630);
and AND3 (N5513, N5509, N3778, N2274);
nand NAND4 (N5514, N5495, N74, N3578, N1320);
and AND4 (N5515, N5510, N563, N862, N3336);
not NOT1 (N5516, N5513);
and AND4 (N5517, N5506, N879, N3162, N3892);
buf BUF1 (N5518, N5517);
nand NAND2 (N5519, N5507, N4147);
nor NOR3 (N5520, N5496, N4749, N4930);
nand NAND3 (N5521, N5514, N1702, N4181);
xor XOR2 (N5522, N5505, N4173);
buf BUF1 (N5523, N5502);
nand NAND4 (N5524, N5522, N3085, N3982, N1608);
not NOT1 (N5525, N5519);
nor NOR2 (N5526, N5518, N3092);
nand NAND3 (N5527, N5480, N2133, N3326);
nor NOR4 (N5528, N5521, N3393, N326, N3271);
and AND3 (N5529, N5515, N2224, N5230);
xor XOR2 (N5530, N5529, N4790);
and AND4 (N5531, N5526, N3277, N3894, N5126);
not NOT1 (N5532, N5516);
or OR2 (N5533, N5520, N4434);
or OR2 (N5534, N5532, N5401);
not NOT1 (N5535, N5524);
or OR4 (N5536, N5530, N3350, N952, N3421);
xor XOR2 (N5537, N5535, N2649);
xor XOR2 (N5538, N5536, N4394);
and AND2 (N5539, N5534, N2954);
nand NAND3 (N5540, N5512, N2261, N1883);
or OR2 (N5541, N5527, N3370);
xor XOR2 (N5542, N5541, N3843);
or OR4 (N5543, N5538, N1983, N3532, N5149);
buf BUF1 (N5544, N5528);
xor XOR2 (N5545, N5540, N5335);
not NOT1 (N5546, N5542);
nor NOR2 (N5547, N5545, N4522);
and AND2 (N5548, N5537, N1854);
not NOT1 (N5549, N5539);
or OR3 (N5550, N5523, N3946, N5125);
and AND3 (N5551, N5525, N3095, N2665);
and AND3 (N5552, N5547, N1079, N1173);
nand NAND3 (N5553, N5544, N1547, N3281);
not NOT1 (N5554, N5548);
and AND3 (N5555, N5553, N171, N240);
buf BUF1 (N5556, N5555);
buf BUF1 (N5557, N5546);
xor XOR2 (N5558, N5543, N644);
xor XOR2 (N5559, N5552, N3760);
buf BUF1 (N5560, N5557);
buf BUF1 (N5561, N5558);
xor XOR2 (N5562, N5556, N2558);
nor NOR3 (N5563, N5549, N124, N4378);
buf BUF1 (N5564, N5550);
and AND3 (N5565, N5533, N2066, N3984);
nor NOR3 (N5566, N5561, N3042, N1860);
nand NAND3 (N5567, N5566, N3554, N4800);
nand NAND3 (N5568, N5562, N1596, N2343);
xor XOR2 (N5569, N5563, N871);
buf BUF1 (N5570, N5568);
not NOT1 (N5571, N5567);
not NOT1 (N5572, N5559);
not NOT1 (N5573, N5572);
or OR4 (N5574, N5560, N1560, N4813, N3729);
and AND2 (N5575, N5574, N1633);
not NOT1 (N5576, N5571);
nand NAND4 (N5577, N5570, N2566, N4172, N898);
and AND4 (N5578, N5551, N5559, N4571, N3452);
nand NAND3 (N5579, N5565, N2240, N2171);
not NOT1 (N5580, N5569);
not NOT1 (N5581, N5573);
nor NOR3 (N5582, N5575, N4354, N5267);
nand NAND2 (N5583, N5582, N5379);
not NOT1 (N5584, N5564);
xor XOR2 (N5585, N5579, N2230);
not NOT1 (N5586, N5576);
nor NOR3 (N5587, N5578, N3436, N1801);
buf BUF1 (N5588, N5587);
not NOT1 (N5589, N5581);
and AND3 (N5590, N5583, N5536, N4463);
nor NOR4 (N5591, N5588, N1448, N4428, N1859);
buf BUF1 (N5592, N5577);
nor NOR3 (N5593, N5589, N5397, N2503);
nand NAND2 (N5594, N5531, N4497);
buf BUF1 (N5595, N5585);
or OR4 (N5596, N5584, N2635, N542, N4121);
nand NAND2 (N5597, N5593, N4300);
nor NOR4 (N5598, N5590, N3313, N1776, N2484);
not NOT1 (N5599, N5586);
buf BUF1 (N5600, N5598);
not NOT1 (N5601, N5580);
or OR2 (N5602, N5600, N896);
buf BUF1 (N5603, N5595);
or OR4 (N5604, N5602, N3868, N1261, N46);
and AND4 (N5605, N5603, N427, N4885, N5549);
buf BUF1 (N5606, N5601);
not NOT1 (N5607, N5599);
not NOT1 (N5608, N5594);
or OR4 (N5609, N5596, N3545, N2826, N2814);
nand NAND4 (N5610, N5605, N1936, N3376, N3701);
or OR2 (N5611, N5609, N4003);
xor XOR2 (N5612, N5604, N5004);
or OR4 (N5613, N5554, N2581, N3181, N2014);
or OR3 (N5614, N5608, N1960, N1130);
not NOT1 (N5615, N5597);
nand NAND4 (N5616, N5606, N411, N1804, N2978);
nor NOR4 (N5617, N5614, N4604, N3749, N1712);
nand NAND3 (N5618, N5611, N2285, N532);
not NOT1 (N5619, N5607);
or OR3 (N5620, N5613, N3101, N3517);
or OR2 (N5621, N5619, N3539);
nor NOR3 (N5622, N5616, N1579, N5440);
buf BUF1 (N5623, N5592);
nand NAND3 (N5624, N5615, N3243, N3808);
not NOT1 (N5625, N5624);
nor NOR4 (N5626, N5612, N1906, N4176, N1599);
buf BUF1 (N5627, N5622);
or OR2 (N5628, N5623, N693);
not NOT1 (N5629, N5628);
or OR2 (N5630, N5618, N1737);
and AND2 (N5631, N5610, N3795);
or OR4 (N5632, N5620, N4421, N5611, N5412);
buf BUF1 (N5633, N5621);
and AND3 (N5634, N5591, N89, N4513);
not NOT1 (N5635, N5632);
or OR3 (N5636, N5625, N4347, N1187);
or OR2 (N5637, N5626, N2188);
and AND4 (N5638, N5629, N5404, N716, N3583);
buf BUF1 (N5639, N5630);
and AND4 (N5640, N5639, N5572, N4344, N3968);
not NOT1 (N5641, N5617);
and AND4 (N5642, N5638, N3234, N3046, N3689);
not NOT1 (N5643, N5635);
not NOT1 (N5644, N5637);
nor NOR2 (N5645, N5640, N1719);
xor XOR2 (N5646, N5634, N1585);
xor XOR2 (N5647, N5643, N4217);
nor NOR4 (N5648, N5627, N208, N3567, N468);
buf BUF1 (N5649, N5642);
xor XOR2 (N5650, N5647, N1762);
and AND2 (N5651, N5650, N2564);
buf BUF1 (N5652, N5648);
or OR4 (N5653, N5651, N3682, N4594, N5457);
nor NOR3 (N5654, N5649, N1018, N439);
xor XOR2 (N5655, N5646, N4651);
and AND4 (N5656, N5644, N3027, N8, N3097);
and AND4 (N5657, N5641, N1922, N2984, N4851);
nor NOR3 (N5658, N5652, N5132, N2611);
buf BUF1 (N5659, N5633);
nand NAND4 (N5660, N5659, N4366, N4696, N4832);
nor NOR4 (N5661, N5653, N2118, N32, N4445);
and AND4 (N5662, N5636, N5650, N3941, N1530);
not NOT1 (N5663, N5661);
buf BUF1 (N5664, N5656);
or OR4 (N5665, N5658, N4793, N2181, N5370);
not NOT1 (N5666, N5654);
nand NAND2 (N5667, N5662, N1859);
not NOT1 (N5668, N5660);
and AND4 (N5669, N5666, N1871, N3637, N933);
nand NAND3 (N5670, N5655, N4053, N2289);
or OR3 (N5671, N5664, N3053, N3187);
nand NAND3 (N5672, N5670, N4244, N4954);
nor NOR4 (N5673, N5667, N2903, N2122, N2926);
not NOT1 (N5674, N5672);
not NOT1 (N5675, N5668);
nand NAND3 (N5676, N5665, N3150, N1303);
buf BUF1 (N5677, N5673);
buf BUF1 (N5678, N5674);
not NOT1 (N5679, N5645);
or OR3 (N5680, N5669, N5622, N3714);
nand NAND2 (N5681, N5657, N436);
or OR2 (N5682, N5663, N4214);
xor XOR2 (N5683, N5682, N1754);
nand NAND2 (N5684, N5680, N4239);
buf BUF1 (N5685, N5683);
or OR3 (N5686, N5681, N482, N114);
nand NAND4 (N5687, N5686, N1672, N467, N608);
or OR4 (N5688, N5685, N2516, N4984, N541);
and AND3 (N5689, N5687, N675, N2064);
xor XOR2 (N5690, N5631, N1824);
nand NAND4 (N5691, N5690, N4031, N3902, N3430);
buf BUF1 (N5692, N5679);
or OR3 (N5693, N5676, N3120, N5103);
not NOT1 (N5694, N5693);
buf BUF1 (N5695, N5677);
buf BUF1 (N5696, N5695);
not NOT1 (N5697, N5684);
xor XOR2 (N5698, N5675, N1601);
buf BUF1 (N5699, N5688);
nor NOR3 (N5700, N5671, N4184, N266);
or OR3 (N5701, N5698, N4240, N1685);
nor NOR2 (N5702, N5700, N5600);
xor XOR2 (N5703, N5689, N4577);
or OR2 (N5704, N5696, N4745);
or OR4 (N5705, N5699, N1427, N5242, N4491);
not NOT1 (N5706, N5692);
nand NAND3 (N5707, N5701, N3105, N2671);
or OR3 (N5708, N5697, N869, N5307);
buf BUF1 (N5709, N5694);
xor XOR2 (N5710, N5704, N2720);
or OR3 (N5711, N5705, N3733, N496);
nand NAND4 (N5712, N5709, N2942, N3870, N1155);
not NOT1 (N5713, N5712);
nand NAND4 (N5714, N5711, N621, N3700, N2077);
or OR3 (N5715, N5708, N473, N1278);
buf BUF1 (N5716, N5702);
nand NAND4 (N5717, N5678, N2876, N3277, N4722);
and AND2 (N5718, N5706, N324);
nor NOR4 (N5719, N5710, N4944, N4716, N2749);
nand NAND3 (N5720, N5703, N2346, N3146);
or OR3 (N5721, N5719, N695, N1301);
not NOT1 (N5722, N5721);
nand NAND3 (N5723, N5691, N4854, N5097);
and AND4 (N5724, N5715, N5328, N5588, N100);
xor XOR2 (N5725, N5724, N4746);
or OR4 (N5726, N5707, N4502, N5048, N1624);
nor NOR2 (N5727, N5722, N1383);
xor XOR2 (N5728, N5723, N1421);
not NOT1 (N5729, N5718);
nand NAND3 (N5730, N5713, N2761, N2612);
or OR3 (N5731, N5727, N2239, N3712);
nand NAND4 (N5732, N5731, N4208, N5336, N3268);
buf BUF1 (N5733, N5729);
not NOT1 (N5734, N5720);
xor XOR2 (N5735, N5725, N5648);
buf BUF1 (N5736, N5730);
or OR3 (N5737, N5716, N384, N2537);
and AND2 (N5738, N5728, N793);
nand NAND4 (N5739, N5734, N4152, N2921, N36);
or OR3 (N5740, N5736, N5500, N4889);
xor XOR2 (N5741, N5740, N99);
or OR2 (N5742, N5714, N4647);
and AND4 (N5743, N5733, N3163, N916, N1987);
or OR3 (N5744, N5742, N887, N4462);
and AND4 (N5745, N5732, N3171, N3038, N3229);
or OR4 (N5746, N5737, N5457, N3246, N1779);
xor XOR2 (N5747, N5745, N1695);
not NOT1 (N5748, N5739);
and AND3 (N5749, N5743, N1041, N413);
xor XOR2 (N5750, N5738, N4484);
xor XOR2 (N5751, N5717, N2724);
nand NAND3 (N5752, N5748, N5291, N2195);
or OR2 (N5753, N5749, N3937);
nor NOR3 (N5754, N5753, N2653, N5421);
not NOT1 (N5755, N5744);
nand NAND2 (N5756, N5750, N1428);
xor XOR2 (N5757, N5752, N1119);
or OR3 (N5758, N5726, N1198, N2011);
not NOT1 (N5759, N5746);
nor NOR4 (N5760, N5735, N1437, N3582, N1509);
nor NOR2 (N5761, N5758, N5586);
not NOT1 (N5762, N5741);
or OR2 (N5763, N5759, N5728);
not NOT1 (N5764, N5755);
xor XOR2 (N5765, N5754, N553);
buf BUF1 (N5766, N5747);
nand NAND4 (N5767, N5763, N406, N2523, N450);
buf BUF1 (N5768, N5751);
xor XOR2 (N5769, N5764, N4194);
xor XOR2 (N5770, N5757, N2966);
nand NAND4 (N5771, N5766, N5440, N780, N3020);
buf BUF1 (N5772, N5765);
not NOT1 (N5773, N5767);
not NOT1 (N5774, N5772);
nand NAND3 (N5775, N5769, N1288, N1958);
or OR4 (N5776, N5760, N1774, N32, N4167);
or OR3 (N5777, N5762, N5745, N3819);
nor NOR4 (N5778, N5771, N4517, N3986, N1204);
and AND3 (N5779, N5756, N3136, N221);
not NOT1 (N5780, N5777);
not NOT1 (N5781, N5780);
xor XOR2 (N5782, N5768, N5672);
nor NOR4 (N5783, N5776, N264, N4176, N4698);
or OR2 (N5784, N5779, N586);
not NOT1 (N5785, N5783);
not NOT1 (N5786, N5778);
xor XOR2 (N5787, N5775, N4246);
buf BUF1 (N5788, N5784);
or OR4 (N5789, N5787, N4771, N4101, N3625);
nand NAND3 (N5790, N5789, N1035, N5354);
not NOT1 (N5791, N5781);
nand NAND4 (N5792, N5773, N4087, N2280, N2102);
buf BUF1 (N5793, N5774);
and AND2 (N5794, N5792, N2506);
not NOT1 (N5795, N5785);
not NOT1 (N5796, N5790);
not NOT1 (N5797, N5793);
and AND2 (N5798, N5796, N1483);
or OR3 (N5799, N5786, N2873, N883);
or OR3 (N5800, N5788, N3531, N232);
buf BUF1 (N5801, N5761);
buf BUF1 (N5802, N5801);
nor NOR4 (N5803, N5799, N2519, N615, N1575);
not NOT1 (N5804, N5782);
and AND2 (N5805, N5795, N4032);
xor XOR2 (N5806, N5794, N906);
nand NAND3 (N5807, N5800, N4714, N1098);
nor NOR4 (N5808, N5805, N218, N2524, N1076);
nand NAND2 (N5809, N5804, N805);
nand NAND3 (N5810, N5808, N2817, N2467);
buf BUF1 (N5811, N5803);
and AND2 (N5812, N5811, N5138);
nor NOR2 (N5813, N5806, N1455);
or OR3 (N5814, N5798, N4132, N1276);
xor XOR2 (N5815, N5791, N2186);
or OR2 (N5816, N5802, N5715);
not NOT1 (N5817, N5809);
or OR2 (N5818, N5797, N648);
nor NOR2 (N5819, N5816, N394);
xor XOR2 (N5820, N5810, N1128);
and AND3 (N5821, N5820, N3163, N296);
buf BUF1 (N5822, N5813);
and AND3 (N5823, N5814, N1732, N5581);
nor NOR3 (N5824, N5822, N5543, N4569);
not NOT1 (N5825, N5823);
or OR3 (N5826, N5817, N2614, N1105);
and AND2 (N5827, N5819, N3693);
buf BUF1 (N5828, N5825);
not NOT1 (N5829, N5807);
nand NAND3 (N5830, N5829, N872, N3058);
and AND3 (N5831, N5818, N5164, N967);
nand NAND2 (N5832, N5826, N1648);
xor XOR2 (N5833, N5815, N3940);
and AND3 (N5834, N5821, N4723, N1984);
or OR3 (N5835, N5770, N4224, N5108);
not NOT1 (N5836, N5830);
or OR3 (N5837, N5833, N4905, N1859);
and AND2 (N5838, N5827, N4537);
not NOT1 (N5839, N5812);
not NOT1 (N5840, N5837);
xor XOR2 (N5841, N5828, N1243);
nand NAND2 (N5842, N5831, N5305);
buf BUF1 (N5843, N5840);
not NOT1 (N5844, N5843);
and AND4 (N5845, N5836, N1140, N1406, N23);
nor NOR4 (N5846, N5835, N237, N3213, N803);
xor XOR2 (N5847, N5824, N4214);
xor XOR2 (N5848, N5838, N4056);
nand NAND4 (N5849, N5842, N3528, N3448, N2957);
and AND3 (N5850, N5845, N5519, N5045);
or OR4 (N5851, N5850, N5298, N5654, N5634);
not NOT1 (N5852, N5832);
nand NAND4 (N5853, N5851, N2661, N534, N1658);
nor NOR4 (N5854, N5853, N1974, N5852, N5714);
nor NOR4 (N5855, N3947, N4665, N2651, N1205);
or OR2 (N5856, N5841, N4571);
nor NOR3 (N5857, N5849, N4667, N4480);
nor NOR2 (N5858, N5834, N354);
and AND3 (N5859, N5858, N415, N4184);
xor XOR2 (N5860, N5848, N5619);
not NOT1 (N5861, N5855);
xor XOR2 (N5862, N5839, N2436);
not NOT1 (N5863, N5847);
xor XOR2 (N5864, N5844, N538);
nor NOR4 (N5865, N5860, N5316, N1944, N249);
buf BUF1 (N5866, N5863);
nand NAND2 (N5867, N5862, N1683);
or OR2 (N5868, N5867, N4109);
xor XOR2 (N5869, N5861, N5489);
nand NAND4 (N5870, N5866, N1109, N2666, N736);
not NOT1 (N5871, N5865);
nand NAND3 (N5872, N5859, N161, N1175);
nand NAND3 (N5873, N5871, N3907, N4766);
xor XOR2 (N5874, N5869, N3824);
nand NAND4 (N5875, N5864, N1670, N51, N4747);
nor NOR3 (N5876, N5846, N3202, N3487);
buf BUF1 (N5877, N5874);
not NOT1 (N5878, N5875);
xor XOR2 (N5879, N5873, N3684);
xor XOR2 (N5880, N5870, N2809);
not NOT1 (N5881, N5877);
xor XOR2 (N5882, N5872, N4492);
not NOT1 (N5883, N5856);
not NOT1 (N5884, N5881);
nand NAND2 (N5885, N5854, N4561);
and AND2 (N5886, N5885, N2568);
and AND2 (N5887, N5883, N5066);
xor XOR2 (N5888, N5876, N2823);
or OR2 (N5889, N5868, N1493);
not NOT1 (N5890, N5882);
xor XOR2 (N5891, N5888, N5297);
nor NOR2 (N5892, N5857, N1034);
and AND3 (N5893, N5880, N444, N4255);
xor XOR2 (N5894, N5879, N2792);
not NOT1 (N5895, N5884);
buf BUF1 (N5896, N5887);
or OR2 (N5897, N5893, N4558);
nand NAND3 (N5898, N5890, N1242, N113);
buf BUF1 (N5899, N5894);
buf BUF1 (N5900, N5896);
not NOT1 (N5901, N5886);
or OR4 (N5902, N5895, N78, N286, N3479);
buf BUF1 (N5903, N5889);
buf BUF1 (N5904, N5903);
nand NAND3 (N5905, N5902, N4676, N2650);
nor NOR3 (N5906, N5899, N1023, N1121);
nand NAND2 (N5907, N5901, N3999);
nand NAND4 (N5908, N5906, N2914, N1069, N755);
xor XOR2 (N5909, N5891, N1292);
or OR4 (N5910, N5905, N1608, N2250, N5717);
nor NOR3 (N5911, N5909, N2683, N3837);
and AND2 (N5912, N5900, N3307);
nor NOR3 (N5913, N5878, N4384, N3988);
and AND3 (N5914, N5913, N229, N359);
not NOT1 (N5915, N5908);
nor NOR3 (N5916, N5910, N619, N4405);
buf BUF1 (N5917, N5898);
nand NAND3 (N5918, N5911, N629, N2362);
nand NAND4 (N5919, N5897, N3895, N4651, N2759);
or OR2 (N5920, N5916, N4841);
not NOT1 (N5921, N5915);
or OR3 (N5922, N5919, N1324, N2344);
xor XOR2 (N5923, N5920, N3266);
nand NAND3 (N5924, N5907, N4876, N4917);
nor NOR4 (N5925, N5923, N4161, N2481, N3888);
nand NAND4 (N5926, N5892, N4657, N805, N3965);
buf BUF1 (N5927, N5904);
and AND3 (N5928, N5926, N4920, N974);
nor NOR4 (N5929, N5917, N2638, N970, N779);
nand NAND4 (N5930, N5918, N877, N1308, N4686);
nor NOR3 (N5931, N5927, N3836, N2938);
not NOT1 (N5932, N5931);
nand NAND2 (N5933, N5929, N3070);
or OR4 (N5934, N5930, N2681, N462, N5721);
nor NOR4 (N5935, N5922, N3589, N3575, N685);
or OR4 (N5936, N5914, N61, N4204, N2320);
and AND4 (N5937, N5935, N2195, N5844, N2555);
not NOT1 (N5938, N5936);
not NOT1 (N5939, N5938);
nor NOR2 (N5940, N5939, N5858);
nor NOR3 (N5941, N5940, N1863, N1740);
not NOT1 (N5942, N5912);
or OR4 (N5943, N5925, N2070, N4911, N4210);
nand NAND3 (N5944, N5921, N4363, N5841);
not NOT1 (N5945, N5943);
nand NAND3 (N5946, N5942, N2466, N5296);
xor XOR2 (N5947, N5934, N4743);
not NOT1 (N5948, N5933);
or OR4 (N5949, N5924, N5377, N4423, N2330);
not NOT1 (N5950, N5944);
and AND3 (N5951, N5949, N4628, N2050);
or OR3 (N5952, N5945, N3236, N3005);
buf BUF1 (N5953, N5951);
nand NAND2 (N5954, N5947, N880);
xor XOR2 (N5955, N5946, N519);
nand NAND2 (N5956, N5937, N4356);
not NOT1 (N5957, N5956);
not NOT1 (N5958, N5950);
xor XOR2 (N5959, N5941, N5693);
nor NOR3 (N5960, N5958, N4335, N1107);
nor NOR4 (N5961, N5948, N3352, N5427, N2845);
nor NOR3 (N5962, N5960, N549, N2445);
and AND4 (N5963, N5932, N3668, N2164, N1172);
not NOT1 (N5964, N5928);
nand NAND2 (N5965, N5963, N2308);
not NOT1 (N5966, N5957);
buf BUF1 (N5967, N5965);
and AND2 (N5968, N5962, N5309);
and AND2 (N5969, N5955, N3092);
buf BUF1 (N5970, N5952);
nor NOR3 (N5971, N5953, N56, N5576);
nand NAND2 (N5972, N5968, N4610);
xor XOR2 (N5973, N5969, N1125);
nor NOR3 (N5974, N5973, N263, N1487);
nor NOR4 (N5975, N5974, N3881, N683, N3270);
not NOT1 (N5976, N5972);
nand NAND3 (N5977, N5966, N4013, N2926);
xor XOR2 (N5978, N5959, N5642);
not NOT1 (N5979, N5970);
and AND4 (N5980, N5954, N211, N5500, N1781);
xor XOR2 (N5981, N5964, N1434);
nand NAND2 (N5982, N5977, N221);
nand NAND2 (N5983, N5967, N3186);
and AND3 (N5984, N5983, N1771, N862);
and AND2 (N5985, N5978, N129);
nand NAND3 (N5986, N5985, N2955, N5953);
and AND3 (N5987, N5980, N2721, N2044);
nor NOR2 (N5988, N5982, N2869);
nor NOR2 (N5989, N5971, N4769);
nor NOR2 (N5990, N5984, N1421);
and AND3 (N5991, N5988, N43, N2970);
nand NAND4 (N5992, N5987, N5215, N4850, N4989);
buf BUF1 (N5993, N5991);
xor XOR2 (N5994, N5986, N1771);
nor NOR3 (N5995, N5990, N2132, N5122);
buf BUF1 (N5996, N5976);
nand NAND3 (N5997, N5975, N5330, N3079);
nor NOR4 (N5998, N5994, N4315, N2726, N182);
not NOT1 (N5999, N5998);
and AND3 (N6000, N5979, N66, N5483);
and AND3 (N6001, N5992, N4507, N4289);
buf BUF1 (N6002, N5996);
buf BUF1 (N6003, N5961);
buf BUF1 (N6004, N5995);
or OR2 (N6005, N5999, N2960);
xor XOR2 (N6006, N6005, N2458);
xor XOR2 (N6007, N5997, N869);
buf BUF1 (N6008, N5989);
and AND4 (N6009, N6003, N1668, N416, N4456);
nand NAND4 (N6010, N6008, N1186, N1314, N1253);
buf BUF1 (N6011, N6001);
and AND2 (N6012, N6007, N4257);
buf BUF1 (N6013, N6006);
or OR3 (N6014, N6013, N5197, N1558);
nor NOR2 (N6015, N6014, N3411);
nor NOR3 (N6016, N6011, N2175, N4197);
nor NOR2 (N6017, N6000, N4059);
nand NAND4 (N6018, N6004, N3709, N2011, N664);
nand NAND4 (N6019, N6017, N4572, N335, N3225);
buf BUF1 (N6020, N5981);
buf BUF1 (N6021, N6016);
nor NOR4 (N6022, N6002, N1714, N3928, N679);
buf BUF1 (N6023, N6019);
buf BUF1 (N6024, N6015);
buf BUF1 (N6025, N6023);
buf BUF1 (N6026, N5993);
or OR4 (N6027, N6022, N169, N1327, N3711);
nand NAND4 (N6028, N6027, N2236, N2699, N1737);
buf BUF1 (N6029, N6025);
or OR4 (N6030, N6020, N4909, N2818, N2207);
buf BUF1 (N6031, N6029);
and AND4 (N6032, N6026, N3440, N235, N2742);
xor XOR2 (N6033, N6012, N917);
or OR3 (N6034, N6031, N515, N1572);
not NOT1 (N6035, N6024);
and AND3 (N6036, N6032, N857, N2680);
nor NOR3 (N6037, N6009, N5428, N918);
and AND4 (N6038, N6018, N5376, N5882, N1145);
nor NOR3 (N6039, N6021, N4308, N5044);
nand NAND4 (N6040, N6034, N5044, N2821, N1599);
not NOT1 (N6041, N6037);
nor NOR2 (N6042, N6030, N5328);
and AND4 (N6043, N6039, N5882, N1209, N4687);
and AND4 (N6044, N6036, N863, N5591, N687);
and AND3 (N6045, N6040, N5163, N3847);
or OR4 (N6046, N6045, N3061, N5379, N3811);
not NOT1 (N6047, N6044);
and AND3 (N6048, N6046, N5314, N4591);
nand NAND3 (N6049, N6035, N1671, N3696);
or OR3 (N6050, N6048, N4582, N3826);
not NOT1 (N6051, N6043);
buf BUF1 (N6052, N6047);
not NOT1 (N6053, N6052);
not NOT1 (N6054, N6053);
buf BUF1 (N6055, N6010);
or OR3 (N6056, N6050, N885, N4475);
buf BUF1 (N6057, N6033);
not NOT1 (N6058, N6038);
xor XOR2 (N6059, N6042, N4370);
or OR2 (N6060, N6055, N4150);
nand NAND4 (N6061, N6056, N3470, N4915, N4305);
buf BUF1 (N6062, N6057);
not NOT1 (N6063, N6059);
xor XOR2 (N6064, N6058, N3061);
nand NAND3 (N6065, N6061, N5858, N2249);
and AND3 (N6066, N6065, N6008, N49);
nor NOR2 (N6067, N6063, N5679);
or OR3 (N6068, N6066, N3087, N2409);
xor XOR2 (N6069, N6064, N5204);
nor NOR4 (N6070, N6028, N1457, N4612, N1565);
nor NOR2 (N6071, N6068, N4682);
or OR4 (N6072, N6049, N3839, N1912, N5013);
not NOT1 (N6073, N6069);
nand NAND4 (N6074, N6041, N2671, N2396, N4994);
buf BUF1 (N6075, N6051);
or OR2 (N6076, N6072, N5153);
not NOT1 (N6077, N6075);
xor XOR2 (N6078, N6074, N661);
nor NOR4 (N6079, N6070, N5824, N2969, N4813);
or OR3 (N6080, N6060, N3130, N178);
or OR4 (N6081, N6078, N5817, N5930, N2170);
buf BUF1 (N6082, N6079);
buf BUF1 (N6083, N6071);
xor XOR2 (N6084, N6080, N4252);
nor NOR2 (N6085, N6073, N3926);
not NOT1 (N6086, N6081);
xor XOR2 (N6087, N6054, N3071);
nor NOR2 (N6088, N6085, N5501);
nand NAND3 (N6089, N6086, N3331, N4671);
nand NAND3 (N6090, N6089, N2591, N3799);
nand NAND2 (N6091, N6082, N3779);
and AND2 (N6092, N6090, N5368);
xor XOR2 (N6093, N6077, N1455);
xor XOR2 (N6094, N6087, N5934);
xor XOR2 (N6095, N6083, N5138);
and AND4 (N6096, N6094, N478, N1719, N4922);
or OR4 (N6097, N6076, N5473, N1814, N4509);
and AND4 (N6098, N6096, N3187, N162, N3319);
nand NAND3 (N6099, N6084, N2760, N653);
or OR4 (N6100, N6095, N2035, N4453, N5539);
or OR4 (N6101, N6092, N1153, N1360, N3808);
xor XOR2 (N6102, N6098, N4876);
xor XOR2 (N6103, N6099, N4005);
or OR4 (N6104, N6091, N1317, N3218, N3755);
or OR4 (N6105, N6101, N3445, N4449, N4387);
xor XOR2 (N6106, N6088, N2672);
xor XOR2 (N6107, N6097, N2559);
not NOT1 (N6108, N6103);
and AND3 (N6109, N6108, N3037, N5288);
buf BUF1 (N6110, N6093);
nand NAND4 (N6111, N6067, N3692, N477, N5766);
nand NAND4 (N6112, N6110, N4014, N1047, N5595);
xor XOR2 (N6113, N6107, N871);
and AND2 (N6114, N6105, N1459);
nor NOR4 (N6115, N6106, N4734, N1340, N2486);
nor NOR2 (N6116, N6115, N885);
and AND3 (N6117, N6113, N3329, N1403);
nand NAND3 (N6118, N6116, N1053, N2122);
not NOT1 (N6119, N6117);
nor NOR4 (N6120, N6114, N2496, N985, N2582);
xor XOR2 (N6121, N6102, N543);
xor XOR2 (N6122, N6119, N492);
and AND3 (N6123, N6104, N3426, N4647);
nand NAND3 (N6124, N6122, N5825, N2751);
and AND2 (N6125, N6062, N3876);
or OR2 (N6126, N6118, N180);
or OR4 (N6127, N6112, N1518, N3016, N3317);
xor XOR2 (N6128, N6126, N4235);
nand NAND2 (N6129, N6123, N303);
nand NAND3 (N6130, N6129, N4053, N4526);
buf BUF1 (N6131, N6121);
buf BUF1 (N6132, N6100);
not NOT1 (N6133, N6111);
xor XOR2 (N6134, N6128, N1769);
or OR4 (N6135, N6125, N3953, N7, N3436);
and AND2 (N6136, N6130, N4470);
nor NOR4 (N6137, N6109, N726, N5583, N5424);
not NOT1 (N6138, N6134);
and AND4 (N6139, N6127, N2818, N2401, N4325);
xor XOR2 (N6140, N6120, N917);
and AND4 (N6141, N6139, N966, N3846, N1141);
buf BUF1 (N6142, N6137);
not NOT1 (N6143, N6132);
buf BUF1 (N6144, N6133);
or OR2 (N6145, N6144, N4921);
not NOT1 (N6146, N6135);
nor NOR4 (N6147, N6138, N6133, N2465, N3079);
not NOT1 (N6148, N6124);
nor NOR3 (N6149, N6131, N2329, N493);
buf BUF1 (N6150, N6148);
and AND4 (N6151, N6142, N5864, N3765, N2040);
not NOT1 (N6152, N6141);
nand NAND4 (N6153, N6152, N685, N1306, N6026);
not NOT1 (N6154, N6147);
or OR3 (N6155, N6149, N4792, N2139);
nand NAND4 (N6156, N6154, N2038, N78, N248);
or OR2 (N6157, N6156, N2112);
not NOT1 (N6158, N6150);
buf BUF1 (N6159, N6145);
or OR3 (N6160, N6159, N4454, N37);
xor XOR2 (N6161, N6155, N3495);
and AND4 (N6162, N6136, N2203, N87, N5941);
and AND4 (N6163, N6153, N1689, N1752, N490);
buf BUF1 (N6164, N6140);
and AND3 (N6165, N6157, N4990, N742);
buf BUF1 (N6166, N6162);
xor XOR2 (N6167, N6160, N1992);
and AND2 (N6168, N6151, N1077);
not NOT1 (N6169, N6165);
not NOT1 (N6170, N6158);
not NOT1 (N6171, N6169);
buf BUF1 (N6172, N6146);
buf BUF1 (N6173, N6161);
not NOT1 (N6174, N6143);
nor NOR3 (N6175, N6163, N5386, N3640);
and AND4 (N6176, N6166, N2439, N6056, N5768);
and AND4 (N6177, N6173, N2095, N6139, N5680);
buf BUF1 (N6178, N6164);
or OR2 (N6179, N6170, N205);
nand NAND2 (N6180, N6176, N4758);
and AND3 (N6181, N6180, N5608, N772);
nand NAND3 (N6182, N6175, N868, N81);
buf BUF1 (N6183, N6168);
or OR4 (N6184, N6182, N2371, N1880, N3608);
or OR2 (N6185, N6177, N3382);
buf BUF1 (N6186, N6181);
or OR2 (N6187, N6184, N258);
not NOT1 (N6188, N6178);
or OR2 (N6189, N6185, N3384);
nor NOR3 (N6190, N6174, N1148, N1435);
nor NOR3 (N6191, N6167, N951, N5800);
not NOT1 (N6192, N6183);
xor XOR2 (N6193, N6186, N5252);
xor XOR2 (N6194, N6187, N5246);
nor NOR3 (N6195, N6192, N3486, N5190);
buf BUF1 (N6196, N6189);
not NOT1 (N6197, N6196);
not NOT1 (N6198, N6190);
or OR4 (N6199, N6171, N4313, N4362, N3161);
or OR3 (N6200, N6195, N5759, N3706);
xor XOR2 (N6201, N6188, N1542);
and AND2 (N6202, N6194, N2969);
and AND3 (N6203, N6193, N1955, N1903);
or OR2 (N6204, N6200, N222);
and AND2 (N6205, N6179, N3982);
or OR3 (N6206, N6197, N3093, N5756);
xor XOR2 (N6207, N6199, N5435);
xor XOR2 (N6208, N6201, N3759);
xor XOR2 (N6209, N6204, N4411);
buf BUF1 (N6210, N6191);
buf BUF1 (N6211, N6207);
not NOT1 (N6212, N6209);
nor NOR3 (N6213, N6172, N3298, N4882);
not NOT1 (N6214, N6210);
buf BUF1 (N6215, N6213);
or OR4 (N6216, N6208, N1024, N1432, N2207);
buf BUF1 (N6217, N6211);
or OR3 (N6218, N6205, N3984, N398);
xor XOR2 (N6219, N6212, N51);
and AND2 (N6220, N6214, N1164);
buf BUF1 (N6221, N6206);
nor NOR4 (N6222, N6218, N2274, N1241, N5853);
or OR4 (N6223, N6202, N1371, N774, N2441);
and AND4 (N6224, N6222, N1536, N4190, N4820);
nor NOR4 (N6225, N6223, N4223, N4303, N1222);
buf BUF1 (N6226, N6225);
nor NOR3 (N6227, N6221, N516, N3297);
nand NAND4 (N6228, N6198, N2334, N1182, N4412);
nand NAND3 (N6229, N6219, N6043, N850);
buf BUF1 (N6230, N6217);
nor NOR4 (N6231, N6224, N2925, N2202, N5890);
and AND4 (N6232, N6227, N1074, N2840, N2955);
buf BUF1 (N6233, N6203);
buf BUF1 (N6234, N6232);
or OR2 (N6235, N6228, N5355);
or OR3 (N6236, N6234, N2100, N5482);
nand NAND4 (N6237, N6215, N2791, N5333, N2667);
not NOT1 (N6238, N6216);
nor NOR3 (N6239, N6238, N1438, N4230);
nor NOR4 (N6240, N6237, N188, N2845, N5777);
or OR2 (N6241, N6229, N1045);
and AND2 (N6242, N6233, N343);
buf BUF1 (N6243, N6231);
nor NOR4 (N6244, N6239, N1009, N1542, N5208);
not NOT1 (N6245, N6226);
nand NAND4 (N6246, N6235, N1939, N5420, N5383);
and AND4 (N6247, N6220, N1366, N6145, N3276);
buf BUF1 (N6248, N6236);
buf BUF1 (N6249, N6230);
and AND3 (N6250, N6249, N5510, N2744);
nor NOR3 (N6251, N6241, N5109, N2351);
buf BUF1 (N6252, N6245);
nand NAND4 (N6253, N6242, N840, N4647, N2040);
nor NOR2 (N6254, N6248, N3180);
nor NOR3 (N6255, N6254, N5876, N2682);
buf BUF1 (N6256, N6253);
and AND2 (N6257, N6256, N2547);
not NOT1 (N6258, N6246);
nand NAND3 (N6259, N6250, N3858, N4047);
buf BUF1 (N6260, N6259);
or OR3 (N6261, N6257, N2762, N6003);
and AND4 (N6262, N6244, N842, N919, N570);
and AND2 (N6263, N6255, N5699);
not NOT1 (N6264, N6243);
not NOT1 (N6265, N6262);
buf BUF1 (N6266, N6260);
buf BUF1 (N6267, N6258);
xor XOR2 (N6268, N6251, N2654);
nand NAND3 (N6269, N6252, N1549, N777);
nand NAND4 (N6270, N6269, N4000, N4057, N1179);
not NOT1 (N6271, N6247);
nor NOR3 (N6272, N6270, N5251, N2108);
not NOT1 (N6273, N6266);
or OR3 (N6274, N6267, N5059, N489);
or OR4 (N6275, N6265, N1360, N6254, N3801);
buf BUF1 (N6276, N6275);
and AND4 (N6277, N6271, N3434, N2640, N5346);
xor XOR2 (N6278, N6263, N5028);
nand NAND4 (N6279, N6278, N1103, N5524, N4887);
nor NOR3 (N6280, N6273, N631, N1989);
xor XOR2 (N6281, N6277, N5897);
not NOT1 (N6282, N6279);
or OR4 (N6283, N6282, N5096, N4894, N3403);
nor NOR3 (N6284, N6268, N1821, N321);
nand NAND2 (N6285, N6261, N1370);
not NOT1 (N6286, N6283);
and AND3 (N6287, N6276, N4289, N811);
buf BUF1 (N6288, N6272);
nor NOR2 (N6289, N6274, N960);
or OR2 (N6290, N6289, N740);
nand NAND4 (N6291, N6287, N5422, N484, N1015);
and AND2 (N6292, N6291, N612);
or OR2 (N6293, N6240, N975);
nor NOR4 (N6294, N6292, N2668, N1163, N517);
not NOT1 (N6295, N6290);
or OR3 (N6296, N6284, N1335, N2878);
nand NAND2 (N6297, N6296, N4547);
nand NAND4 (N6298, N6286, N5287, N4883, N493);
or OR2 (N6299, N6280, N999);
nor NOR4 (N6300, N6293, N3927, N298, N4792);
nor NOR2 (N6301, N6297, N493);
not NOT1 (N6302, N6301);
not NOT1 (N6303, N6299);
or OR2 (N6304, N6295, N5810);
not NOT1 (N6305, N6294);
and AND2 (N6306, N6305, N5899);
xor XOR2 (N6307, N6285, N2660);
nor NOR2 (N6308, N6302, N6105);
xor XOR2 (N6309, N6298, N1817);
not NOT1 (N6310, N6307);
buf BUF1 (N6311, N6303);
nor NOR3 (N6312, N6281, N5038, N4695);
xor XOR2 (N6313, N6308, N3275);
buf BUF1 (N6314, N6264);
xor XOR2 (N6315, N6310, N1008);
or OR4 (N6316, N6314, N573, N4320, N636);
xor XOR2 (N6317, N6306, N3206);
nand NAND4 (N6318, N6315, N3202, N3087, N1177);
and AND3 (N6319, N6313, N2514, N2374);
nor NOR3 (N6320, N6319, N1987, N1976);
nand NAND3 (N6321, N6318, N250, N917);
or OR4 (N6322, N6316, N6265, N4258, N5239);
or OR3 (N6323, N6309, N3310, N6214);
not NOT1 (N6324, N6321);
and AND2 (N6325, N6322, N5814);
nand NAND4 (N6326, N6323, N5932, N5344, N869);
not NOT1 (N6327, N6304);
not NOT1 (N6328, N6317);
not NOT1 (N6329, N6312);
or OR4 (N6330, N6328, N4745, N4153, N88);
not NOT1 (N6331, N6320);
not NOT1 (N6332, N6300);
buf BUF1 (N6333, N6331);
nor NOR2 (N6334, N6326, N4836);
nand NAND2 (N6335, N6324, N1672);
nand NAND4 (N6336, N6288, N3757, N1392, N898);
and AND2 (N6337, N6330, N2005);
nand NAND2 (N6338, N6333, N925);
or OR4 (N6339, N6338, N2027, N352, N1512);
nor NOR2 (N6340, N6334, N2856);
or OR3 (N6341, N6337, N204, N4043);
and AND2 (N6342, N6340, N4450);
nor NOR2 (N6343, N6327, N2381);
nand NAND2 (N6344, N6341, N3672);
nor NOR4 (N6345, N6339, N3627, N288, N4648);
nand NAND2 (N6346, N6335, N5175);
nand NAND2 (N6347, N6343, N588);
nand NAND4 (N6348, N6344, N4274, N4510, N1323);
xor XOR2 (N6349, N6346, N690);
not NOT1 (N6350, N6311);
nand NAND3 (N6351, N6342, N2125, N3082);
xor XOR2 (N6352, N6332, N463);
not NOT1 (N6353, N6347);
xor XOR2 (N6354, N6351, N5060);
xor XOR2 (N6355, N6329, N4873);
nor NOR4 (N6356, N6349, N4098, N5178, N2623);
buf BUF1 (N6357, N6356);
or OR4 (N6358, N6348, N2275, N5089, N1075);
xor XOR2 (N6359, N6354, N2766);
and AND2 (N6360, N6359, N2572);
buf BUF1 (N6361, N6345);
nor NOR2 (N6362, N6350, N1325);
nor NOR3 (N6363, N6358, N5177, N1678);
xor XOR2 (N6364, N6357, N6048);
and AND2 (N6365, N6355, N3415);
nand NAND4 (N6366, N6363, N4328, N2209, N2453);
xor XOR2 (N6367, N6353, N4166);
buf BUF1 (N6368, N6336);
and AND2 (N6369, N6325, N5687);
and AND3 (N6370, N6369, N4242, N998);
nor NOR3 (N6371, N6360, N5832, N1074);
or OR2 (N6372, N6370, N5014);
and AND2 (N6373, N6364, N2065);
buf BUF1 (N6374, N6371);
nor NOR3 (N6375, N6372, N40, N1867);
and AND4 (N6376, N6373, N1795, N4534, N3181);
xor XOR2 (N6377, N6375, N5218);
nor NOR2 (N6378, N6361, N4364);
xor XOR2 (N6379, N6352, N4309);
buf BUF1 (N6380, N6377);
not NOT1 (N6381, N6362);
xor XOR2 (N6382, N6374, N3875);
buf BUF1 (N6383, N6382);
nor NOR4 (N6384, N6383, N5413, N2756, N845);
nor NOR3 (N6385, N6366, N3735, N895);
or OR4 (N6386, N6384, N3999, N6122, N1051);
and AND4 (N6387, N6365, N2864, N6382, N3102);
nor NOR4 (N6388, N6379, N3214, N3527, N3228);
and AND4 (N6389, N6388, N1325, N2227, N2180);
buf BUF1 (N6390, N6367);
not NOT1 (N6391, N6389);
and AND2 (N6392, N6376, N1321);
nor NOR3 (N6393, N6380, N4941, N2879);
buf BUF1 (N6394, N6391);
xor XOR2 (N6395, N6387, N4670);
nor NOR2 (N6396, N6385, N5988);
or OR4 (N6397, N6381, N2108, N3987, N5936);
nand NAND2 (N6398, N6378, N4215);
buf BUF1 (N6399, N6397);
nor NOR3 (N6400, N6395, N72, N2362);
and AND4 (N6401, N6399, N2526, N1053, N2885);
nand NAND2 (N6402, N6392, N5119);
not NOT1 (N6403, N6393);
or OR4 (N6404, N6402, N4401, N2989, N3764);
and AND3 (N6405, N6400, N710, N814);
nor NOR3 (N6406, N6396, N4581, N3873);
xor XOR2 (N6407, N6404, N49);
or OR3 (N6408, N6386, N2741, N4315);
xor XOR2 (N6409, N6407, N5348);
xor XOR2 (N6410, N6403, N4044);
nor NOR4 (N6411, N6408, N85, N920, N94);
and AND3 (N6412, N6411, N6145, N4713);
or OR3 (N6413, N6409, N4220, N4518);
xor XOR2 (N6414, N6413, N704);
and AND2 (N6415, N6390, N613);
not NOT1 (N6416, N6368);
or OR3 (N6417, N6401, N216, N4483);
nand NAND2 (N6418, N6417, N4389);
nand NAND4 (N6419, N6418, N764, N5198, N6316);
or OR3 (N6420, N6394, N965, N2946);
buf BUF1 (N6421, N6406);
not NOT1 (N6422, N6414);
or OR4 (N6423, N6398, N2927, N5519, N4646);
or OR2 (N6424, N6405, N4974);
not NOT1 (N6425, N6421);
or OR3 (N6426, N6424, N5842, N276);
xor XOR2 (N6427, N6426, N3178);
buf BUF1 (N6428, N6423);
buf BUF1 (N6429, N6425);
nor NOR4 (N6430, N6422, N4562, N4130, N4676);
xor XOR2 (N6431, N6428, N55);
not NOT1 (N6432, N6420);
xor XOR2 (N6433, N6415, N1429);
nand NAND2 (N6434, N6416, N3891);
xor XOR2 (N6435, N6427, N1618);
nand NAND2 (N6436, N6410, N2998);
not NOT1 (N6437, N6431);
nand NAND2 (N6438, N6436, N4379);
and AND2 (N6439, N6430, N1922);
xor XOR2 (N6440, N6438, N690);
nor NOR2 (N6441, N6433, N4541);
xor XOR2 (N6442, N6441, N4049);
xor XOR2 (N6443, N6432, N6331);
and AND4 (N6444, N6429, N4583, N5576, N235);
and AND4 (N6445, N6444, N1457, N2270, N47);
and AND3 (N6446, N6445, N6279, N1487);
nand NAND3 (N6447, N6412, N475, N4248);
or OR4 (N6448, N6439, N3097, N1923, N1975);
nor NOR3 (N6449, N6447, N6156, N2539);
nand NAND4 (N6450, N6437, N5686, N828, N5103);
and AND2 (N6451, N6450, N5594);
and AND2 (N6452, N6443, N4701);
buf BUF1 (N6453, N6448);
not NOT1 (N6454, N6451);
or OR2 (N6455, N6453, N4988);
or OR3 (N6456, N6454, N44, N1233);
xor XOR2 (N6457, N6449, N261);
and AND4 (N6458, N6446, N4999, N483, N5595);
nor NOR2 (N6459, N6452, N5151);
buf BUF1 (N6460, N6455);
nand NAND3 (N6461, N6458, N1102, N5394);
xor XOR2 (N6462, N6435, N5132);
buf BUF1 (N6463, N6460);
xor XOR2 (N6464, N6442, N5916);
buf BUF1 (N6465, N6462);
not NOT1 (N6466, N6440);
nand NAND3 (N6467, N6434, N4995, N4875);
or OR4 (N6468, N6419, N6196, N697, N4541);
nor NOR2 (N6469, N6465, N4562);
buf BUF1 (N6470, N6457);
xor XOR2 (N6471, N6456, N342);
xor XOR2 (N6472, N6467, N4065);
nand NAND3 (N6473, N6463, N3686, N5107);
not NOT1 (N6474, N6461);
buf BUF1 (N6475, N6468);
or OR3 (N6476, N6459, N2031, N4903);
and AND2 (N6477, N6471, N2266);
xor XOR2 (N6478, N6476, N833);
nor NOR3 (N6479, N6478, N5234, N3818);
and AND3 (N6480, N6466, N6430, N1684);
buf BUF1 (N6481, N6473);
or OR3 (N6482, N6477, N1451, N8);
nand NAND4 (N6483, N6470, N5502, N10, N948);
not NOT1 (N6484, N6483);
or OR3 (N6485, N6482, N1615, N1771);
nand NAND2 (N6486, N6481, N2634);
buf BUF1 (N6487, N6474);
nor NOR4 (N6488, N6475, N4538, N4325, N4913);
nor NOR3 (N6489, N6485, N3439, N4072);
nand NAND4 (N6490, N6489, N6286, N4686, N2414);
buf BUF1 (N6491, N6480);
buf BUF1 (N6492, N6490);
nand NAND2 (N6493, N6472, N367);
buf BUF1 (N6494, N6492);
not NOT1 (N6495, N6469);
and AND3 (N6496, N6487, N5398, N5980);
nor NOR2 (N6497, N6464, N1392);
nor NOR4 (N6498, N6491, N4927, N4374, N6154);
nand NAND4 (N6499, N6486, N1552, N5022, N1183);
not NOT1 (N6500, N6484);
not NOT1 (N6501, N6499);
or OR3 (N6502, N6488, N6461, N3664);
and AND4 (N6503, N6500, N4363, N3084, N3439);
not NOT1 (N6504, N6495);
nor NOR3 (N6505, N6494, N3002, N3814);
nor NOR3 (N6506, N6501, N2206, N4216);
or OR4 (N6507, N6493, N3726, N6207, N1705);
not NOT1 (N6508, N6498);
buf BUF1 (N6509, N6505);
or OR2 (N6510, N6502, N6128);
nor NOR4 (N6511, N6506, N27, N4373, N1438);
nand NAND4 (N6512, N6496, N5101, N4467, N4497);
xor XOR2 (N6513, N6508, N1999);
or OR4 (N6514, N6512, N290, N3054, N3097);
nor NOR2 (N6515, N6503, N3064);
nor NOR4 (N6516, N6514, N3000, N351, N3823);
nand NAND3 (N6517, N6504, N3063, N5702);
xor XOR2 (N6518, N6479, N802);
buf BUF1 (N6519, N6513);
not NOT1 (N6520, N6507);
buf BUF1 (N6521, N6519);
not NOT1 (N6522, N6509);
nor NOR4 (N6523, N6516, N1363, N5914, N682);
not NOT1 (N6524, N6523);
or OR2 (N6525, N6515, N4765);
not NOT1 (N6526, N6522);
or OR3 (N6527, N6525, N337, N5079);
xor XOR2 (N6528, N6521, N5152);
nor NOR2 (N6529, N6526, N4260);
nand NAND2 (N6530, N6517, N5109);
xor XOR2 (N6531, N6511, N1301);
or OR2 (N6532, N6518, N4308);
not NOT1 (N6533, N6531);
nand NAND2 (N6534, N6532, N5773);
or OR2 (N6535, N6530, N3070);
nand NAND2 (N6536, N6533, N1333);
and AND3 (N6537, N6527, N3853, N3933);
not NOT1 (N6538, N6524);
nand NAND2 (N6539, N6535, N2548);
xor XOR2 (N6540, N6537, N2868);
or OR3 (N6541, N6534, N1273, N1054);
nand NAND2 (N6542, N6497, N3307);
xor XOR2 (N6543, N6510, N2704);
nor NOR4 (N6544, N6541, N2315, N4294, N1555);
and AND2 (N6545, N6544, N1313);
nor NOR2 (N6546, N6542, N4924);
xor XOR2 (N6547, N6540, N2658);
not NOT1 (N6548, N6543);
nand NAND4 (N6549, N6536, N371, N5233, N3288);
and AND3 (N6550, N6528, N3730, N6484);
or OR3 (N6551, N6538, N2745, N4794);
not NOT1 (N6552, N6548);
xor XOR2 (N6553, N6520, N1891);
nor NOR2 (N6554, N6539, N4393);
not NOT1 (N6555, N6546);
xor XOR2 (N6556, N6547, N4353);
not NOT1 (N6557, N6554);
or OR4 (N6558, N6549, N2686, N730, N6544);
and AND4 (N6559, N6553, N4398, N2294, N2569);
or OR4 (N6560, N6557, N2035, N2418, N425);
nor NOR4 (N6561, N6529, N448, N2432, N1692);
buf BUF1 (N6562, N6556);
and AND2 (N6563, N6562, N3559);
xor XOR2 (N6564, N6550, N2168);
or OR4 (N6565, N6558, N6139, N1881, N104);
nor NOR2 (N6566, N6563, N3691);
not NOT1 (N6567, N6560);
xor XOR2 (N6568, N6555, N761);
not NOT1 (N6569, N6559);
not NOT1 (N6570, N6552);
buf BUF1 (N6571, N6567);
nand NAND3 (N6572, N6564, N508, N2641);
xor XOR2 (N6573, N6566, N2647);
nand NAND3 (N6574, N6570, N3869, N500);
nor NOR4 (N6575, N6572, N1808, N882, N6162);
and AND2 (N6576, N6575, N4811);
xor XOR2 (N6577, N6561, N3753);
buf BUF1 (N6578, N6574);
xor XOR2 (N6579, N6578, N3113);
buf BUF1 (N6580, N6565);
not NOT1 (N6581, N6577);
xor XOR2 (N6582, N6579, N6316);
nor NOR3 (N6583, N6582, N6100, N1300);
buf BUF1 (N6584, N6569);
not NOT1 (N6585, N6545);
nor NOR3 (N6586, N6571, N302, N295);
nor NOR2 (N6587, N6573, N4471);
buf BUF1 (N6588, N6580);
nand NAND2 (N6589, N6576, N574);
xor XOR2 (N6590, N6583, N1861);
nor NOR3 (N6591, N6590, N3201, N1795);
or OR3 (N6592, N6586, N174, N2679);
buf BUF1 (N6593, N6592);
nor NOR2 (N6594, N6587, N3215);
nand NAND3 (N6595, N6585, N1123, N5420);
buf BUF1 (N6596, N6595);
nand NAND3 (N6597, N6593, N3359, N5069);
buf BUF1 (N6598, N6596);
buf BUF1 (N6599, N6589);
xor XOR2 (N6600, N6551, N4662);
or OR3 (N6601, N6591, N2216, N3721);
nand NAND4 (N6602, N6599, N1540, N1897, N4508);
or OR4 (N6603, N6600, N4083, N2786, N690);
xor XOR2 (N6604, N6598, N5370);
nand NAND4 (N6605, N6601, N2772, N5134, N708);
nand NAND2 (N6606, N6604, N4613);
nor NOR2 (N6607, N6588, N686);
nand NAND3 (N6608, N6568, N2070, N2451);
or OR4 (N6609, N6606, N2439, N3513, N5796);
xor XOR2 (N6610, N6609, N2881);
and AND2 (N6611, N6602, N3534);
xor XOR2 (N6612, N6608, N4637);
or OR2 (N6613, N6581, N3822);
nor NOR3 (N6614, N6611, N3564, N5287);
nor NOR3 (N6615, N6610, N242, N2936);
buf BUF1 (N6616, N6603);
nor NOR3 (N6617, N6605, N5602, N4498);
buf BUF1 (N6618, N6607);
or OR2 (N6619, N6597, N6004);
and AND2 (N6620, N6584, N2874);
and AND4 (N6621, N6613, N2205, N6123, N1500);
and AND3 (N6622, N6594, N4764, N5705);
xor XOR2 (N6623, N6612, N216);
xor XOR2 (N6624, N6620, N110);
or OR4 (N6625, N6622, N3491, N3571, N5176);
nor NOR2 (N6626, N6623, N5482);
and AND2 (N6627, N6621, N5694);
buf BUF1 (N6628, N6615);
and AND2 (N6629, N6624, N1816);
not NOT1 (N6630, N6618);
and AND2 (N6631, N6629, N3812);
nor NOR2 (N6632, N6616, N2162);
not NOT1 (N6633, N6625);
buf BUF1 (N6634, N6628);
nand NAND4 (N6635, N6631, N1087, N4522, N4220);
nor NOR4 (N6636, N6634, N1564, N2878, N2253);
buf BUF1 (N6637, N6632);
or OR2 (N6638, N6636, N5877);
nand NAND4 (N6639, N6630, N2453, N4060, N5162);
not NOT1 (N6640, N6626);
not NOT1 (N6641, N6627);
nand NAND2 (N6642, N6638, N4174);
buf BUF1 (N6643, N6635);
buf BUF1 (N6644, N6641);
and AND3 (N6645, N6643, N5886, N5295);
not NOT1 (N6646, N6614);
not NOT1 (N6647, N6642);
not NOT1 (N6648, N6646);
nand NAND2 (N6649, N6617, N449);
nor NOR2 (N6650, N6619, N5230);
or OR2 (N6651, N6650, N2097);
xor XOR2 (N6652, N6633, N2634);
not NOT1 (N6653, N6645);
not NOT1 (N6654, N6653);
buf BUF1 (N6655, N6648);
buf BUF1 (N6656, N6647);
xor XOR2 (N6657, N6654, N1455);
nand NAND3 (N6658, N6651, N5093, N2109);
buf BUF1 (N6659, N6649);
or OR2 (N6660, N6639, N2500);
and AND4 (N6661, N6652, N871, N6422, N3819);
or OR2 (N6662, N6658, N3993);
buf BUF1 (N6663, N6655);
nand NAND4 (N6664, N6661, N5699, N3856, N3209);
nand NAND4 (N6665, N6637, N6529, N2972, N4041);
not NOT1 (N6666, N6660);
and AND2 (N6667, N6657, N5324);
nand NAND3 (N6668, N6664, N3929, N2286);
nor NOR2 (N6669, N6656, N4101);
or OR3 (N6670, N6662, N2243, N3898);
and AND2 (N6671, N6668, N3719);
buf BUF1 (N6672, N6671);
xor XOR2 (N6673, N6666, N1463);
and AND4 (N6674, N6672, N886, N1194, N2726);
xor XOR2 (N6675, N6673, N4705);
xor XOR2 (N6676, N6644, N1476);
not NOT1 (N6677, N6663);
buf BUF1 (N6678, N6675);
nor NOR2 (N6679, N6659, N404);
xor XOR2 (N6680, N6679, N2284);
nor NOR4 (N6681, N6677, N4133, N1312, N906);
nor NOR4 (N6682, N6670, N4377, N1671, N1371);
buf BUF1 (N6683, N6674);
nor NOR3 (N6684, N6681, N6298, N5810);
and AND3 (N6685, N6678, N6676, N5432);
nand NAND3 (N6686, N4600, N3307, N4921);
or OR2 (N6687, N6640, N2803);
nor NOR2 (N6688, N6665, N1372);
xor XOR2 (N6689, N6669, N1786);
buf BUF1 (N6690, N6686);
nor NOR4 (N6691, N6680, N4740, N4334, N3385);
and AND3 (N6692, N6682, N2815, N5325);
not NOT1 (N6693, N6691);
buf BUF1 (N6694, N6683);
or OR4 (N6695, N6667, N4927, N4602, N839);
xor XOR2 (N6696, N6694, N2999);
not NOT1 (N6697, N6688);
nor NOR3 (N6698, N6695, N6579, N1743);
and AND4 (N6699, N6696, N2810, N2011, N927);
and AND2 (N6700, N6693, N5506);
nor NOR3 (N6701, N6689, N6404, N2830);
xor XOR2 (N6702, N6700, N6529);
buf BUF1 (N6703, N6701);
nand NAND3 (N6704, N6698, N5665, N2955);
and AND2 (N6705, N6704, N4826);
nor NOR3 (N6706, N6705, N1602, N887);
nand NAND4 (N6707, N6697, N2686, N6440, N2132);
or OR2 (N6708, N6707, N48);
xor XOR2 (N6709, N6702, N1191);
nor NOR3 (N6710, N6687, N129, N5965);
xor XOR2 (N6711, N6708, N770);
nor NOR3 (N6712, N6711, N4084, N5066);
or OR4 (N6713, N6685, N1133, N3059, N5369);
buf BUF1 (N6714, N6706);
not NOT1 (N6715, N6703);
nor NOR2 (N6716, N6710, N1890);
not NOT1 (N6717, N6692);
nand NAND3 (N6718, N6715, N6246, N5913);
nor NOR4 (N6719, N6714, N6469, N5101, N4976);
and AND4 (N6720, N6719, N1180, N702, N1958);
and AND3 (N6721, N6718, N6017, N5228);
or OR3 (N6722, N6721, N3723, N5691);
nand NAND3 (N6723, N6684, N3741, N5219);
and AND4 (N6724, N6722, N4614, N3883, N1232);
and AND4 (N6725, N6690, N2372, N39, N3819);
nor NOR3 (N6726, N6699, N37, N3325);
and AND3 (N6727, N6717, N110, N6158);
xor XOR2 (N6728, N6727, N3141);
and AND2 (N6729, N6724, N6169);
nand NAND3 (N6730, N6712, N4635, N1893);
nor NOR4 (N6731, N6725, N5090, N90, N358);
and AND4 (N6732, N6713, N948, N6143, N2805);
not NOT1 (N6733, N6729);
not NOT1 (N6734, N6728);
not NOT1 (N6735, N6733);
nand NAND3 (N6736, N6720, N4643, N541);
nand NAND3 (N6737, N6726, N4962, N4259);
nand NAND3 (N6738, N6716, N1494, N2443);
xor XOR2 (N6739, N6735, N1391);
buf BUF1 (N6740, N6737);
nor NOR2 (N6741, N6723, N1404);
nand NAND2 (N6742, N6731, N3486);
xor XOR2 (N6743, N6736, N4658);
nand NAND4 (N6744, N6732, N4509, N511, N1362);
buf BUF1 (N6745, N6734);
nor NOR3 (N6746, N6740, N6528, N5523);
not NOT1 (N6747, N6743);
or OR2 (N6748, N6741, N6431);
nor NOR2 (N6749, N6730, N2725);
buf BUF1 (N6750, N6745);
nor NOR2 (N6751, N6746, N5689);
or OR2 (N6752, N6747, N4819);
not NOT1 (N6753, N6709);
nand NAND2 (N6754, N6749, N4915);
or OR3 (N6755, N6752, N1137, N833);
not NOT1 (N6756, N6738);
not NOT1 (N6757, N6748);
buf BUF1 (N6758, N6751);
nand NAND3 (N6759, N6754, N2048, N5088);
or OR2 (N6760, N6739, N2154);
nand NAND4 (N6761, N6760, N5232, N2123, N3916);
nand NAND4 (N6762, N6757, N3308, N747, N4412);
nand NAND3 (N6763, N6762, N6737, N1631);
or OR4 (N6764, N6763, N1576, N673, N2496);
nor NOR2 (N6765, N6758, N6615);
nand NAND3 (N6766, N6753, N2903, N727);
nand NAND2 (N6767, N6759, N6424);
xor XOR2 (N6768, N6767, N5265);
not NOT1 (N6769, N6756);
not NOT1 (N6770, N6742);
xor XOR2 (N6771, N6765, N5734);
xor XOR2 (N6772, N6761, N3889);
nand NAND3 (N6773, N6750, N4155, N1737);
not NOT1 (N6774, N6771);
nand NAND2 (N6775, N6770, N380);
or OR3 (N6776, N6768, N2622, N1552);
nor NOR2 (N6777, N6766, N2348);
nand NAND3 (N6778, N6776, N1317, N4651);
xor XOR2 (N6779, N6774, N208);
xor XOR2 (N6780, N6778, N1872);
not NOT1 (N6781, N6780);
not NOT1 (N6782, N6773);
nor NOR3 (N6783, N6779, N3479, N6112);
not NOT1 (N6784, N6755);
xor XOR2 (N6785, N6782, N5647);
or OR2 (N6786, N6744, N2971);
or OR3 (N6787, N6785, N5828, N281);
and AND4 (N6788, N6784, N1597, N2764, N3047);
and AND3 (N6789, N6783, N1268, N6668);
buf BUF1 (N6790, N6789);
xor XOR2 (N6791, N6786, N4552);
not NOT1 (N6792, N6791);
not NOT1 (N6793, N6792);
nor NOR2 (N6794, N6793, N1081);
nand NAND3 (N6795, N6787, N2438, N5976);
buf BUF1 (N6796, N6775);
xor XOR2 (N6797, N6777, N3629);
not NOT1 (N6798, N6796);
nand NAND2 (N6799, N6772, N5025);
buf BUF1 (N6800, N6788);
xor XOR2 (N6801, N6795, N2224);
not NOT1 (N6802, N6769);
not NOT1 (N6803, N6800);
xor XOR2 (N6804, N6797, N1024);
or OR3 (N6805, N6794, N5266, N3731);
xor XOR2 (N6806, N6802, N1800);
not NOT1 (N6807, N6801);
nor NOR2 (N6808, N6764, N1086);
and AND4 (N6809, N6808, N4368, N4128, N2388);
nand NAND2 (N6810, N6805, N3440);
nand NAND2 (N6811, N6807, N4601);
and AND4 (N6812, N6811, N1228, N5544, N563);
nand NAND2 (N6813, N6806, N4367);
xor XOR2 (N6814, N6809, N4267);
nor NOR3 (N6815, N6799, N6737, N1914);
buf BUF1 (N6816, N6798);
not NOT1 (N6817, N6814);
nand NAND4 (N6818, N6812, N6040, N3180, N1942);
not NOT1 (N6819, N6813);
xor XOR2 (N6820, N6804, N4463);
and AND2 (N6821, N6816, N5287);
buf BUF1 (N6822, N6781);
or OR4 (N6823, N6817, N988, N3359, N3606);
buf BUF1 (N6824, N6818);
nand NAND2 (N6825, N6824, N2926);
and AND3 (N6826, N6825, N621, N1692);
or OR4 (N6827, N6790, N3858, N890, N1700);
nand NAND2 (N6828, N6820, N1659);
nor NOR3 (N6829, N6810, N5063, N211);
and AND4 (N6830, N6819, N1225, N2751, N3041);
nand NAND4 (N6831, N6815, N3087, N4690, N1731);
buf BUF1 (N6832, N6803);
and AND4 (N6833, N6821, N4296, N1785, N2659);
nand NAND4 (N6834, N6827, N5557, N6069, N6171);
nor NOR4 (N6835, N6831, N5543, N1262, N3391);
or OR4 (N6836, N6822, N5942, N838, N6035);
nand NAND4 (N6837, N6826, N6807, N5356, N6703);
xor XOR2 (N6838, N6836, N663);
not NOT1 (N6839, N6829);
xor XOR2 (N6840, N6835, N6207);
nand NAND4 (N6841, N6830, N1396, N6743, N5637);
not NOT1 (N6842, N6828);
not NOT1 (N6843, N6839);
nand NAND3 (N6844, N6833, N4803, N1420);
nand NAND4 (N6845, N6840, N745, N372, N2303);
nand NAND2 (N6846, N6823, N796);
buf BUF1 (N6847, N6841);
xor XOR2 (N6848, N6834, N5160);
nand NAND4 (N6849, N6832, N4312, N3480, N6035);
not NOT1 (N6850, N6838);
xor XOR2 (N6851, N6843, N5549);
nor NOR3 (N6852, N6837, N3430, N2003);
xor XOR2 (N6853, N6847, N6170);
and AND2 (N6854, N6853, N159);
xor XOR2 (N6855, N6844, N4136);
not NOT1 (N6856, N6846);
nor NOR2 (N6857, N6848, N305);
and AND2 (N6858, N6850, N6035);
or OR4 (N6859, N6851, N5970, N3637, N5502);
nor NOR4 (N6860, N6856, N2311, N2061, N4902);
nand NAND4 (N6861, N6854, N1842, N1987, N5066);
and AND4 (N6862, N6842, N3452, N3420, N1702);
or OR2 (N6863, N6861, N5118);
not NOT1 (N6864, N6860);
not NOT1 (N6865, N6857);
or OR3 (N6866, N6865, N4704, N6579);
not NOT1 (N6867, N6864);
and AND4 (N6868, N6862, N3604, N2178, N5717);
or OR4 (N6869, N6855, N5648, N4639, N75);
buf BUF1 (N6870, N6852);
nor NOR2 (N6871, N6866, N2746);
xor XOR2 (N6872, N6870, N918);
nand NAND2 (N6873, N6867, N6319);
xor XOR2 (N6874, N6845, N3494);
nor NOR4 (N6875, N6868, N4196, N6355, N4144);
and AND3 (N6876, N6863, N5389, N3956);
not NOT1 (N6877, N6875);
nand NAND3 (N6878, N6877, N3865, N2232);
buf BUF1 (N6879, N6873);
nor NOR2 (N6880, N6876, N3472);
nand NAND2 (N6881, N6872, N6690);
or OR2 (N6882, N6878, N5141);
nor NOR4 (N6883, N6869, N3140, N3115, N5311);
and AND3 (N6884, N6879, N4716, N4457);
xor XOR2 (N6885, N6881, N4333);
or OR4 (N6886, N6884, N5657, N3637, N5151);
nand NAND3 (N6887, N6882, N6255, N1424);
nand NAND3 (N6888, N6883, N3342, N3144);
xor XOR2 (N6889, N6874, N1585);
not NOT1 (N6890, N6871);
xor XOR2 (N6891, N6858, N2425);
or OR3 (N6892, N6891, N522, N686);
buf BUF1 (N6893, N6886);
nor NOR2 (N6894, N6880, N3254);
not NOT1 (N6895, N6885);
xor XOR2 (N6896, N6895, N3116);
or OR3 (N6897, N6892, N3778, N2780);
nand NAND4 (N6898, N6897, N2934, N1825, N3678);
and AND4 (N6899, N6898, N1058, N546, N1858);
or OR2 (N6900, N6849, N6632);
xor XOR2 (N6901, N6894, N5294);
xor XOR2 (N6902, N6888, N4607);
xor XOR2 (N6903, N6859, N963);
and AND2 (N6904, N6896, N4952);
and AND3 (N6905, N6887, N2407, N3563);
nand NAND2 (N6906, N6902, N2994);
not NOT1 (N6907, N6890);
or OR2 (N6908, N6904, N4928);
buf BUF1 (N6909, N6906);
and AND3 (N6910, N6901, N3399, N2390);
nor NOR4 (N6911, N6903, N5353, N4508, N5148);
not NOT1 (N6912, N6900);
not NOT1 (N6913, N6908);
not NOT1 (N6914, N6910);
not NOT1 (N6915, N6907);
buf BUF1 (N6916, N6913);
nand NAND4 (N6917, N6915, N3626, N5383, N2385);
nor NOR4 (N6918, N6905, N5270, N6906, N6915);
and AND3 (N6919, N6917, N5747, N2529);
not NOT1 (N6920, N6919);
nand NAND3 (N6921, N6899, N1629, N5482);
nor NOR3 (N6922, N6889, N4841, N546);
and AND2 (N6923, N6918, N1085);
not NOT1 (N6924, N6916);
not NOT1 (N6925, N6912);
buf BUF1 (N6926, N6922);
or OR2 (N6927, N6920, N6453);
nor NOR3 (N6928, N6909, N4168, N5647);
nor NOR4 (N6929, N6914, N5954, N144, N6843);
xor XOR2 (N6930, N6893, N2781);
or OR3 (N6931, N6921, N458, N2660);
buf BUF1 (N6932, N6911);
or OR3 (N6933, N6931, N4037, N6657);
xor XOR2 (N6934, N6933, N4874);
or OR2 (N6935, N6928, N5334);
or OR2 (N6936, N6934, N3425);
buf BUF1 (N6937, N6926);
nand NAND3 (N6938, N6935, N5562, N6678);
xor XOR2 (N6939, N6927, N5784);
buf BUF1 (N6940, N6923);
and AND3 (N6941, N6929, N1394, N2105);
xor XOR2 (N6942, N6930, N3723);
and AND2 (N6943, N6924, N4392);
buf BUF1 (N6944, N6937);
xor XOR2 (N6945, N6938, N6062);
xor XOR2 (N6946, N6940, N955);
not NOT1 (N6947, N6942);
not NOT1 (N6948, N6939);
nand NAND3 (N6949, N6944, N4230, N3131);
nor NOR3 (N6950, N6941, N294, N4956);
not NOT1 (N6951, N6945);
and AND2 (N6952, N6947, N1233);
buf BUF1 (N6953, N6951);
and AND2 (N6954, N6946, N3135);
and AND4 (N6955, N6932, N3218, N2307, N6657);
buf BUF1 (N6956, N6952);
nand NAND4 (N6957, N6943, N5048, N6627, N4944);
and AND3 (N6958, N6936, N575, N1482);
buf BUF1 (N6959, N6954);
nand NAND4 (N6960, N6955, N967, N4235, N1402);
xor XOR2 (N6961, N6950, N5634);
or OR3 (N6962, N6953, N3854, N4878);
xor XOR2 (N6963, N6956, N990);
not NOT1 (N6964, N6925);
not NOT1 (N6965, N6960);
buf BUF1 (N6966, N6962);
nor NOR4 (N6967, N6958, N5155, N2157, N2791);
nand NAND2 (N6968, N6957, N229);
nor NOR2 (N6969, N6959, N3623);
nand NAND3 (N6970, N6968, N6411, N2744);
xor XOR2 (N6971, N6969, N4525);
buf BUF1 (N6972, N6964);
xor XOR2 (N6973, N6961, N998);
not NOT1 (N6974, N6971);
xor XOR2 (N6975, N6972, N3397);
nor NOR4 (N6976, N6966, N6147, N6045, N653);
and AND4 (N6977, N6973, N1754, N5926, N5221);
buf BUF1 (N6978, N6948);
nand NAND2 (N6979, N6976, N3593);
not NOT1 (N6980, N6949);
not NOT1 (N6981, N6975);
xor XOR2 (N6982, N6978, N6616);
nand NAND2 (N6983, N6981, N2521);
and AND2 (N6984, N6979, N1021);
not NOT1 (N6985, N6977);
or OR4 (N6986, N6984, N3026, N4809, N5084);
xor XOR2 (N6987, N6985, N3909);
and AND4 (N6988, N6983, N3143, N4869, N1088);
xor XOR2 (N6989, N6967, N6154);
nand NAND3 (N6990, N6987, N546, N1415);
not NOT1 (N6991, N6974);
and AND3 (N6992, N6990, N349, N95);
not NOT1 (N6993, N6965);
nor NOR3 (N6994, N6988, N2115, N3109);
nor NOR4 (N6995, N6994, N4647, N2659, N4529);
or OR4 (N6996, N6963, N6878, N6794, N2351);
nor NOR2 (N6997, N6992, N6946);
nor NOR4 (N6998, N6995, N5395, N8, N2346);
not NOT1 (N6999, N6980);
nand NAND2 (N7000, N6997, N5132);
nand NAND3 (N7001, N6999, N5900, N801);
or OR3 (N7002, N7000, N2779, N3361);
nand NAND2 (N7003, N6989, N2148);
and AND2 (N7004, N7002, N2176);
nand NAND3 (N7005, N6996, N6274, N6623);
nand NAND3 (N7006, N6986, N4481, N5089);
or OR2 (N7007, N6991, N5178);
and AND3 (N7008, N6993, N3131, N6713);
and AND4 (N7009, N7007, N4823, N4616, N5265);
and AND2 (N7010, N6998, N494);
and AND2 (N7011, N7008, N2591);
and AND3 (N7012, N7003, N2005, N3780);
or OR2 (N7013, N7010, N4166);
nor NOR3 (N7014, N7004, N6243, N5795);
nand NAND4 (N7015, N7013, N18, N3322, N5762);
buf BUF1 (N7016, N7001);
or OR4 (N7017, N7011, N5362, N1933, N3654);
buf BUF1 (N7018, N7005);
not NOT1 (N7019, N7018);
not NOT1 (N7020, N7012);
not NOT1 (N7021, N6982);
buf BUF1 (N7022, N7006);
buf BUF1 (N7023, N7020);
or OR3 (N7024, N7015, N5967, N2048);
nand NAND2 (N7025, N7014, N705);
not NOT1 (N7026, N7019);
and AND3 (N7027, N7024, N2727, N2686);
or OR2 (N7028, N7027, N3649);
nand NAND3 (N7029, N7017, N6152, N1444);
and AND4 (N7030, N7022, N2424, N727, N63);
nor NOR4 (N7031, N7025, N3323, N3797, N4647);
xor XOR2 (N7032, N7009, N1327);
and AND3 (N7033, N7030, N3224, N1553);
and AND3 (N7034, N7026, N3557, N6968);
and AND2 (N7035, N7028, N6325);
nand NAND2 (N7036, N7033, N2192);
buf BUF1 (N7037, N6970);
nand NAND3 (N7038, N7036, N2319, N1036);
not NOT1 (N7039, N7021);
xor XOR2 (N7040, N7023, N109);
not NOT1 (N7041, N7034);
not NOT1 (N7042, N7040);
not NOT1 (N7043, N7042);
nand NAND4 (N7044, N7039, N4882, N1903, N296);
buf BUF1 (N7045, N7041);
or OR2 (N7046, N7043, N1897);
nor NOR3 (N7047, N7031, N4815, N717);
nand NAND3 (N7048, N7032, N3042, N2803);
nand NAND2 (N7049, N7044, N2237);
and AND4 (N7050, N7047, N4103, N6328, N1586);
or OR3 (N7051, N7016, N2980, N3146);
nand NAND3 (N7052, N7050, N3178, N6920);
xor XOR2 (N7053, N7029, N4697);
buf BUF1 (N7054, N7053);
and AND2 (N7055, N7037, N1010);
nor NOR2 (N7056, N7048, N1922);
nand NAND3 (N7057, N7035, N3767, N4279);
nor NOR2 (N7058, N7049, N5502);
not NOT1 (N7059, N7038);
nor NOR2 (N7060, N7058, N6546);
or OR3 (N7061, N7059, N3665, N3322);
not NOT1 (N7062, N7051);
nand NAND3 (N7063, N7060, N4601, N2539);
not NOT1 (N7064, N7063);
or OR2 (N7065, N7057, N903);
not NOT1 (N7066, N7045);
buf BUF1 (N7067, N7055);
or OR4 (N7068, N7066, N1246, N4221, N6794);
not NOT1 (N7069, N7068);
nand NAND2 (N7070, N7054, N1110);
buf BUF1 (N7071, N7056);
or OR3 (N7072, N7070, N2894, N4856);
or OR3 (N7073, N7072, N1979, N3163);
nand NAND4 (N7074, N7073, N5694, N2646, N1026);
xor XOR2 (N7075, N7074, N2548);
or OR3 (N7076, N7062, N4191, N4285);
xor XOR2 (N7077, N7069, N7048);
nand NAND4 (N7078, N7065, N5113, N6124, N4580);
and AND2 (N7079, N7076, N5068);
and AND2 (N7080, N7079, N4564);
buf BUF1 (N7081, N7075);
or OR4 (N7082, N7061, N5798, N622, N3466);
buf BUF1 (N7083, N7052);
and AND3 (N7084, N7064, N4568, N2305);
not NOT1 (N7085, N7067);
and AND2 (N7086, N7078, N673);
or OR2 (N7087, N7071, N4923);
or OR4 (N7088, N7080, N4409, N5367, N4752);
or OR3 (N7089, N7084, N7082, N4399);
xor XOR2 (N7090, N4988, N5048);
buf BUF1 (N7091, N7087);
xor XOR2 (N7092, N7089, N389);
or OR2 (N7093, N7083, N1100);
or OR2 (N7094, N7092, N1786);
and AND4 (N7095, N7086, N2448, N621, N5768);
and AND2 (N7096, N7091, N4072);
nand NAND2 (N7097, N7046, N6892);
nor NOR3 (N7098, N7088, N2205, N3953);
not NOT1 (N7099, N7077);
and AND2 (N7100, N7090, N545);
or OR2 (N7101, N7096, N5478);
and AND3 (N7102, N7095, N3489, N854);
buf BUF1 (N7103, N7094);
and AND4 (N7104, N7085, N6031, N3082, N818);
and AND4 (N7105, N7098, N513, N777, N1297);
buf BUF1 (N7106, N7097);
or OR3 (N7107, N7106, N1543, N2765);
xor XOR2 (N7108, N7093, N6713);
and AND3 (N7109, N7102, N6399, N6059);
nand NAND4 (N7110, N7099, N6277, N4849, N3706);
or OR2 (N7111, N7104, N4301);
nor NOR3 (N7112, N7103, N396, N2217);
not NOT1 (N7113, N7108);
not NOT1 (N7114, N7081);
nand NAND4 (N7115, N7112, N4195, N514, N4252);
not NOT1 (N7116, N7105);
xor XOR2 (N7117, N7107, N5961);
or OR4 (N7118, N7113, N4562, N45, N521);
buf BUF1 (N7119, N7116);
or OR4 (N7120, N7111, N874, N1716, N5824);
not NOT1 (N7121, N7118);
xor XOR2 (N7122, N7115, N537);
xor XOR2 (N7123, N7110, N5060);
nand NAND2 (N7124, N7121, N1381);
and AND2 (N7125, N7120, N4605);
and AND4 (N7126, N7100, N4171, N3344, N3051);
nor NOR2 (N7127, N7124, N4278);
not NOT1 (N7128, N7101);
or OR2 (N7129, N7123, N953);
not NOT1 (N7130, N7117);
and AND3 (N7131, N7125, N2492, N6448);
xor XOR2 (N7132, N7131, N418);
nor NOR4 (N7133, N7114, N3668, N6839, N6572);
not NOT1 (N7134, N7127);
buf BUF1 (N7135, N7134);
not NOT1 (N7136, N7135);
buf BUF1 (N7137, N7129);
and AND4 (N7138, N7137, N6180, N1490, N167);
and AND3 (N7139, N7130, N167, N2365);
nand NAND3 (N7140, N7138, N5625, N3783);
xor XOR2 (N7141, N7119, N1537);
nand NAND3 (N7142, N7141, N4284, N2948);
and AND4 (N7143, N7122, N794, N3807, N5165);
xor XOR2 (N7144, N7133, N6197);
and AND4 (N7145, N7136, N5432, N2154, N2705);
nor NOR4 (N7146, N7128, N6591, N723, N678);
or OR2 (N7147, N7146, N6308);
or OR3 (N7148, N7144, N4032, N6167);
xor XOR2 (N7149, N7142, N4534);
and AND2 (N7150, N7148, N6136);
xor XOR2 (N7151, N7143, N1887);
or OR4 (N7152, N7140, N4272, N3287, N5413);
xor XOR2 (N7153, N7145, N5471);
nor NOR3 (N7154, N7152, N4955, N4941);
xor XOR2 (N7155, N7132, N2686);
nor NOR4 (N7156, N7155, N2966, N3127, N4662);
xor XOR2 (N7157, N7156, N3207);
xor XOR2 (N7158, N7109, N4102);
nor NOR3 (N7159, N7153, N5469, N260);
nor NOR4 (N7160, N7150, N6202, N1587, N199);
and AND4 (N7161, N7126, N3008, N4061, N18);
nand NAND2 (N7162, N7158, N3745);
buf BUF1 (N7163, N7160);
and AND4 (N7164, N7154, N884, N3115, N5524);
nand NAND3 (N7165, N7151, N4601, N6805);
buf BUF1 (N7166, N7163);
buf BUF1 (N7167, N7149);
xor XOR2 (N7168, N7165, N5182);
and AND3 (N7169, N7139, N6830, N5405);
not NOT1 (N7170, N7157);
nand NAND3 (N7171, N7162, N1524, N6563);
xor XOR2 (N7172, N7171, N6121);
not NOT1 (N7173, N7172);
buf BUF1 (N7174, N7169);
or OR4 (N7175, N7174, N1604, N588, N5626);
nand NAND4 (N7176, N7175, N4242, N2153, N1298);
nand NAND4 (N7177, N7166, N945, N3302, N3192);
not NOT1 (N7178, N7170);
buf BUF1 (N7179, N7159);
nor NOR4 (N7180, N7176, N4311, N3599, N975);
or OR2 (N7181, N7173, N3763);
or OR2 (N7182, N7178, N3125);
and AND4 (N7183, N7164, N4411, N367, N4758);
buf BUF1 (N7184, N7180);
xor XOR2 (N7185, N7182, N841);
xor XOR2 (N7186, N7167, N6772);
nor NOR4 (N7187, N7181, N2274, N1874, N4602);
not NOT1 (N7188, N7184);
xor XOR2 (N7189, N7186, N4562);
nand NAND4 (N7190, N7179, N1987, N2747, N4840);
nor NOR4 (N7191, N7147, N4347, N4895, N4225);
nor NOR4 (N7192, N7161, N2656, N3805, N591);
xor XOR2 (N7193, N7189, N2662);
nand NAND4 (N7194, N7188, N4341, N82, N6868);
or OR3 (N7195, N7183, N53, N800);
nor NOR4 (N7196, N7191, N6986, N2132, N6430);
xor XOR2 (N7197, N7187, N1854);
nand NAND2 (N7198, N7177, N3753);
nand NAND2 (N7199, N7185, N1400);
nand NAND3 (N7200, N7199, N7093, N1261);
nor NOR2 (N7201, N7200, N6560);
or OR2 (N7202, N7193, N2649);
nand NAND3 (N7203, N7202, N4164, N2713);
nor NOR2 (N7204, N7203, N6321);
not NOT1 (N7205, N7196);
nor NOR2 (N7206, N7204, N3794);
nand NAND3 (N7207, N7198, N7192, N4660);
nor NOR4 (N7208, N3871, N4552, N5543, N5092);
or OR4 (N7209, N7168, N4834, N175, N5010);
nor NOR2 (N7210, N7201, N6401);
xor XOR2 (N7211, N7190, N5368);
xor XOR2 (N7212, N7208, N3228);
xor XOR2 (N7213, N7205, N3282);
nand NAND3 (N7214, N7197, N3585, N1560);
nand NAND2 (N7215, N7206, N2832);
not NOT1 (N7216, N7215);
buf BUF1 (N7217, N7207);
and AND4 (N7218, N7194, N6635, N1156, N6507);
nor NOR4 (N7219, N7214, N5175, N4446, N4969);
not NOT1 (N7220, N7216);
xor XOR2 (N7221, N7195, N774);
nand NAND4 (N7222, N7213, N57, N593, N528);
buf BUF1 (N7223, N7222);
buf BUF1 (N7224, N7210);
buf BUF1 (N7225, N7220);
buf BUF1 (N7226, N7221);
nor NOR2 (N7227, N7224, N2915);
buf BUF1 (N7228, N7218);
nor NOR3 (N7229, N7211, N6333, N3133);
xor XOR2 (N7230, N7226, N3803);
or OR4 (N7231, N7230, N6626, N4807, N427);
xor XOR2 (N7232, N7212, N3114);
or OR2 (N7233, N7231, N4477);
or OR2 (N7234, N7209, N294);
buf BUF1 (N7235, N7232);
nor NOR3 (N7236, N7223, N5674, N2195);
or OR4 (N7237, N7228, N6129, N1688, N6754);
nor NOR4 (N7238, N7225, N3569, N4486, N4626);
xor XOR2 (N7239, N7227, N856);
xor XOR2 (N7240, N7239, N3180);
buf BUF1 (N7241, N7238);
not NOT1 (N7242, N7233);
not NOT1 (N7243, N7235);
not NOT1 (N7244, N7240);
or OR3 (N7245, N7217, N2148, N6513);
not NOT1 (N7246, N7244);
not NOT1 (N7247, N7234);
nand NAND3 (N7248, N7219, N2248, N2304);
nor NOR3 (N7249, N7229, N5000, N6203);
buf BUF1 (N7250, N7247);
nor NOR2 (N7251, N7242, N5446);
nand NAND2 (N7252, N7246, N2376);
xor XOR2 (N7253, N7249, N2305);
not NOT1 (N7254, N7245);
and AND2 (N7255, N7252, N4395);
buf BUF1 (N7256, N7248);
nand NAND3 (N7257, N7241, N1280, N6440);
xor XOR2 (N7258, N7256, N1602);
or OR2 (N7259, N7237, N4494);
and AND2 (N7260, N7255, N6313);
nand NAND2 (N7261, N7251, N1592);
nand NAND3 (N7262, N7253, N727, N6910);
nor NOR3 (N7263, N7257, N6771, N5353);
or OR3 (N7264, N7259, N642, N1239);
and AND2 (N7265, N7254, N7046);
and AND3 (N7266, N7260, N6078, N3097);
or OR2 (N7267, N7262, N5061);
nor NOR3 (N7268, N7265, N4429, N3680);
or OR3 (N7269, N7267, N5123, N1776);
or OR3 (N7270, N7258, N3716, N4148);
nor NOR2 (N7271, N7268, N1988);
or OR4 (N7272, N7271, N4646, N3436, N359);
and AND4 (N7273, N7236, N5645, N1990, N3702);
and AND4 (N7274, N7261, N477, N3539, N6375);
and AND4 (N7275, N7270, N6411, N2936, N1226);
nand NAND2 (N7276, N7266, N4563);
and AND4 (N7277, N7273, N6134, N7004, N6268);
or OR3 (N7278, N7269, N4897, N2041);
nor NOR3 (N7279, N7264, N5170, N4237);
buf BUF1 (N7280, N7274);
nor NOR2 (N7281, N7263, N2492);
xor XOR2 (N7282, N7250, N2346);
buf BUF1 (N7283, N7275);
not NOT1 (N7284, N7283);
nand NAND4 (N7285, N7280, N5172, N375, N6753);
nor NOR4 (N7286, N7281, N6013, N3913, N2370);
nor NOR3 (N7287, N7243, N1057, N1546);
buf BUF1 (N7288, N7278);
nor NOR2 (N7289, N7279, N5530);
buf BUF1 (N7290, N7272);
nand NAND2 (N7291, N7282, N7198);
and AND3 (N7292, N7276, N5455, N5524);
not NOT1 (N7293, N7291);
not NOT1 (N7294, N7290);
not NOT1 (N7295, N7286);
and AND3 (N7296, N7295, N4160, N3443);
nand NAND2 (N7297, N7277, N1935);
nand NAND2 (N7298, N7294, N310);
xor XOR2 (N7299, N7293, N1645);
buf BUF1 (N7300, N7289);
and AND4 (N7301, N7298, N3005, N2577, N4842);
and AND2 (N7302, N7299, N6663);
buf BUF1 (N7303, N7300);
nor NOR3 (N7304, N7284, N2724, N1820);
not NOT1 (N7305, N7303);
xor XOR2 (N7306, N7305, N4472);
not NOT1 (N7307, N7301);
not NOT1 (N7308, N7287);
and AND4 (N7309, N7302, N7121, N620, N1896);
xor XOR2 (N7310, N7292, N2406);
or OR2 (N7311, N7310, N6470);
nand NAND4 (N7312, N7297, N5572, N3424, N5705);
buf BUF1 (N7313, N7312);
not NOT1 (N7314, N7296);
nand NAND4 (N7315, N7307, N2230, N656, N1626);
xor XOR2 (N7316, N7315, N80);
xor XOR2 (N7317, N7316, N739);
or OR2 (N7318, N7311, N2092);
nor NOR4 (N7319, N7304, N4742, N167, N2650);
and AND2 (N7320, N7314, N773);
and AND2 (N7321, N7318, N3420);
and AND2 (N7322, N7317, N4090);
or OR2 (N7323, N7321, N1715);
or OR3 (N7324, N7319, N7314, N7254);
nand NAND3 (N7325, N7285, N3762, N2402);
not NOT1 (N7326, N7324);
not NOT1 (N7327, N7309);
xor XOR2 (N7328, N7323, N6573);
or OR4 (N7329, N7313, N3347, N680, N3934);
nor NOR3 (N7330, N7306, N2049, N4943);
buf BUF1 (N7331, N7329);
and AND4 (N7332, N7327, N4609, N6779, N5817);
nor NOR4 (N7333, N7325, N4015, N1262, N5587);
xor XOR2 (N7334, N7332, N5284);
nor NOR2 (N7335, N7308, N6100);
or OR2 (N7336, N7331, N1572);
or OR3 (N7337, N7335, N7265, N6383);
or OR4 (N7338, N7330, N3254, N6529, N6111);
xor XOR2 (N7339, N7338, N5794);
and AND4 (N7340, N7326, N1131, N5881, N6418);
not NOT1 (N7341, N7322);
buf BUF1 (N7342, N7336);
nor NOR4 (N7343, N7320, N1270, N3971, N124);
xor XOR2 (N7344, N7328, N2938);
or OR3 (N7345, N7333, N167, N2271);
xor XOR2 (N7346, N7345, N5369);
nand NAND4 (N7347, N7346, N4153, N7229, N4441);
or OR3 (N7348, N7341, N1108, N5016);
not NOT1 (N7349, N7347);
nand NAND4 (N7350, N7348, N6558, N5853, N3757);
not NOT1 (N7351, N7340);
and AND2 (N7352, N7342, N420);
and AND2 (N7353, N7351, N7064);
or OR4 (N7354, N7337, N5462, N6372, N1586);
or OR2 (N7355, N7334, N1699);
and AND2 (N7356, N7343, N6716);
nor NOR4 (N7357, N7352, N4267, N746, N6088);
not NOT1 (N7358, N7344);
nor NOR2 (N7359, N7353, N7104);
xor XOR2 (N7360, N7288, N4953);
nor NOR2 (N7361, N7357, N4998);
or OR3 (N7362, N7354, N1773, N810);
and AND4 (N7363, N7339, N5417, N613, N5953);
xor XOR2 (N7364, N7363, N499);
xor XOR2 (N7365, N7349, N1003);
nand NAND4 (N7366, N7350, N6881, N1082, N5923);
not NOT1 (N7367, N7361);
nor NOR4 (N7368, N7366, N2611, N200, N5388);
nor NOR2 (N7369, N7358, N3751);
not NOT1 (N7370, N7364);
not NOT1 (N7371, N7359);
not NOT1 (N7372, N7369);
not NOT1 (N7373, N7370);
xor XOR2 (N7374, N7365, N3439);
nor NOR4 (N7375, N7372, N6998, N7068, N709);
buf BUF1 (N7376, N7367);
nor NOR2 (N7377, N7360, N6271);
nor NOR2 (N7378, N7362, N1459);
not NOT1 (N7379, N7356);
nor NOR3 (N7380, N7379, N6410, N2336);
xor XOR2 (N7381, N7376, N5233);
or OR2 (N7382, N7377, N6142);
nor NOR2 (N7383, N7371, N4685);
nor NOR4 (N7384, N7382, N7102, N2665, N456);
buf BUF1 (N7385, N7381);
nor NOR4 (N7386, N7383, N1658, N6207, N7368);
nor NOR3 (N7387, N4596, N5563, N4235);
and AND4 (N7388, N7380, N1780, N2270, N4670);
or OR2 (N7389, N7388, N6077);
or OR4 (N7390, N7387, N1994, N219, N1150);
not NOT1 (N7391, N7355);
or OR2 (N7392, N7386, N2284);
nand NAND4 (N7393, N7373, N6727, N71, N5976);
and AND4 (N7394, N7390, N1804, N909, N2651);
xor XOR2 (N7395, N7389, N4438);
nand NAND2 (N7396, N7393, N4970);
nor NOR2 (N7397, N7378, N2331);
xor XOR2 (N7398, N7395, N4043);
nor NOR3 (N7399, N7397, N391, N6719);
and AND2 (N7400, N7392, N3723);
or OR2 (N7401, N7374, N3200);
and AND3 (N7402, N7396, N6499, N1520);
not NOT1 (N7403, N7375);
buf BUF1 (N7404, N7384);
and AND2 (N7405, N7403, N3844);
buf BUF1 (N7406, N7400);
or OR2 (N7407, N7405, N1712);
nand NAND4 (N7408, N7385, N5390, N4961, N4303);
nand NAND4 (N7409, N7408, N4653, N2482, N1005);
nor NOR3 (N7410, N7406, N4182, N3404);
nor NOR2 (N7411, N7407, N5506);
buf BUF1 (N7412, N7409);
nand NAND4 (N7413, N7411, N4379, N4740, N3016);
nor NOR4 (N7414, N7402, N1467, N2253, N3519);
nand NAND3 (N7415, N7401, N5210, N5843);
nand NAND4 (N7416, N7391, N173, N7356, N1798);
nor NOR4 (N7417, N7404, N4839, N6972, N3788);
nand NAND4 (N7418, N7412, N5918, N1149, N6590);
not NOT1 (N7419, N7418);
nand NAND2 (N7420, N7394, N368);
buf BUF1 (N7421, N7415);
xor XOR2 (N7422, N7413, N5248);
nor NOR3 (N7423, N7416, N2845, N5396);
nand NAND4 (N7424, N7414, N6285, N6140, N1279);
or OR3 (N7425, N7419, N5609, N1112);
nor NOR2 (N7426, N7420, N3434);
not NOT1 (N7427, N7417);
xor XOR2 (N7428, N7398, N1985);
and AND2 (N7429, N7410, N3235);
not NOT1 (N7430, N7423);
xor XOR2 (N7431, N7426, N1751);
buf BUF1 (N7432, N7425);
nand NAND2 (N7433, N7427, N2596);
nor NOR2 (N7434, N7430, N1854);
nand NAND3 (N7435, N7429, N4346, N1150);
buf BUF1 (N7436, N7399);
not NOT1 (N7437, N7428);
buf BUF1 (N7438, N7433);
or OR2 (N7439, N7435, N6804);
buf BUF1 (N7440, N7439);
not NOT1 (N7441, N7422);
not NOT1 (N7442, N7434);
or OR2 (N7443, N7436, N4986);
and AND4 (N7444, N7440, N1843, N2183, N2921);
xor XOR2 (N7445, N7432, N1354);
not NOT1 (N7446, N7444);
xor XOR2 (N7447, N7442, N3820);
buf BUF1 (N7448, N7438);
or OR2 (N7449, N7447, N7065);
and AND3 (N7450, N7431, N5954, N2051);
and AND4 (N7451, N7446, N2957, N1340, N3736);
and AND4 (N7452, N7443, N6305, N7400, N7320);
and AND4 (N7453, N7437, N6647, N1924, N5301);
xor XOR2 (N7454, N7441, N1025);
xor XOR2 (N7455, N7449, N1413);
not NOT1 (N7456, N7455);
or OR2 (N7457, N7450, N9);
or OR3 (N7458, N7456, N4843, N4418);
or OR3 (N7459, N7457, N7405, N6722);
nor NOR4 (N7460, N7448, N2835, N1649, N3588);
nor NOR3 (N7461, N7452, N2517, N5158);
not NOT1 (N7462, N7461);
buf BUF1 (N7463, N7424);
nand NAND3 (N7464, N7459, N3052, N5677);
buf BUF1 (N7465, N7445);
not NOT1 (N7466, N7458);
nor NOR2 (N7467, N7463, N6068);
and AND4 (N7468, N7464, N3015, N1766, N327);
not NOT1 (N7469, N7454);
xor XOR2 (N7470, N7460, N1222);
nor NOR4 (N7471, N7466, N5890, N4117, N1829);
or OR4 (N7472, N7470, N887, N3022, N869);
nand NAND3 (N7473, N7467, N1039, N4319);
buf BUF1 (N7474, N7462);
nand NAND3 (N7475, N7472, N5179, N3405);
nor NOR4 (N7476, N7465, N6328, N1603, N6120);
xor XOR2 (N7477, N7475, N5160);
buf BUF1 (N7478, N7476);
nand NAND2 (N7479, N7474, N2967);
or OR2 (N7480, N7479, N3705);
nor NOR3 (N7481, N7469, N7176, N7427);
nor NOR4 (N7482, N7477, N5850, N3512, N3965);
and AND2 (N7483, N7468, N158);
xor XOR2 (N7484, N7478, N726);
nor NOR2 (N7485, N7480, N715);
and AND2 (N7486, N7471, N3894);
and AND4 (N7487, N7485, N4633, N6033, N5448);
nor NOR2 (N7488, N7453, N2546);
nor NOR4 (N7489, N7483, N4823, N2571, N3126);
not NOT1 (N7490, N7484);
nor NOR3 (N7491, N7486, N803, N559);
nand NAND2 (N7492, N7451, N770);
and AND2 (N7493, N7482, N2499);
not NOT1 (N7494, N7473);
xor XOR2 (N7495, N7492, N4820);
not NOT1 (N7496, N7490);
nand NAND3 (N7497, N7491, N7120, N5770);
xor XOR2 (N7498, N7496, N5346);
buf BUF1 (N7499, N7494);
nor NOR3 (N7500, N7498, N4746, N6921);
or OR4 (N7501, N7493, N6899, N5585, N6428);
or OR4 (N7502, N7489, N3304, N3715, N3381);
and AND3 (N7503, N7497, N6425, N4498);
nand NAND4 (N7504, N7495, N4633, N462, N6500);
not NOT1 (N7505, N7499);
or OR3 (N7506, N7504, N7375, N2397);
not NOT1 (N7507, N7505);
nand NAND2 (N7508, N7500, N2394);
or OR3 (N7509, N7503, N1742, N5926);
buf BUF1 (N7510, N7501);
or OR2 (N7511, N7488, N6135);
and AND3 (N7512, N7509, N6199, N3156);
or OR4 (N7513, N7487, N6659, N5422, N3745);
not NOT1 (N7514, N7511);
not NOT1 (N7515, N7508);
nand NAND2 (N7516, N7513, N2910);
nand NAND2 (N7517, N7510, N1020);
or OR3 (N7518, N7517, N1292, N5552);
nor NOR2 (N7519, N7515, N4049);
nor NOR4 (N7520, N7507, N4742, N4627, N6346);
and AND4 (N7521, N7502, N4792, N3305, N3305);
not NOT1 (N7522, N7519);
buf BUF1 (N7523, N7521);
nor NOR4 (N7524, N7512, N4937, N4788, N1361);
buf BUF1 (N7525, N7522);
nand NAND2 (N7526, N7514, N6521);
and AND4 (N7527, N7526, N875, N980, N99);
nor NOR2 (N7528, N7516, N5870);
nand NAND2 (N7529, N7518, N3521);
and AND2 (N7530, N7523, N6241);
nor NOR4 (N7531, N7530, N631, N5595, N4347);
not NOT1 (N7532, N7525);
or OR3 (N7533, N7421, N6481, N5432);
or OR4 (N7534, N7520, N5682, N3759, N4342);
nand NAND4 (N7535, N7529, N5250, N3872, N6106);
nand NAND2 (N7536, N7533, N4467);
nor NOR4 (N7537, N7528, N6110, N4727, N4942);
or OR2 (N7538, N7481, N1022);
or OR2 (N7539, N7538, N3023);
buf BUF1 (N7540, N7534);
not NOT1 (N7541, N7531);
nor NOR2 (N7542, N7524, N1070);
not NOT1 (N7543, N7506);
nand NAND2 (N7544, N7541, N5027);
nand NAND4 (N7545, N7532, N5600, N1889, N2589);
xor XOR2 (N7546, N7543, N3120);
xor XOR2 (N7547, N7536, N2277);
buf BUF1 (N7548, N7545);
xor XOR2 (N7549, N7527, N6049);
not NOT1 (N7550, N7546);
not NOT1 (N7551, N7549);
and AND2 (N7552, N7535, N737);
xor XOR2 (N7553, N7544, N2114);
xor XOR2 (N7554, N7540, N5562);
and AND4 (N7555, N7553, N6251, N5182, N4674);
and AND2 (N7556, N7551, N4710);
and AND3 (N7557, N7547, N5115, N4150);
or OR3 (N7558, N7554, N4215, N2787);
not NOT1 (N7559, N7557);
or OR2 (N7560, N7548, N6960);
nand NAND3 (N7561, N7539, N7031, N6381);
buf BUF1 (N7562, N7542);
or OR4 (N7563, N7556, N6118, N5719, N6699);
or OR2 (N7564, N7559, N7535);
nor NOR2 (N7565, N7562, N6987);
and AND2 (N7566, N7537, N5505);
not NOT1 (N7567, N7558);
buf BUF1 (N7568, N7563);
and AND2 (N7569, N7555, N3357);
or OR3 (N7570, N7568, N6453, N883);
and AND2 (N7571, N7570, N2506);
nand NAND2 (N7572, N7560, N3849);
xor XOR2 (N7573, N7550, N5297);
not NOT1 (N7574, N7573);
nor NOR4 (N7575, N7574, N4246, N6382, N2184);
nor NOR2 (N7576, N7569, N7550);
buf BUF1 (N7577, N7571);
buf BUF1 (N7578, N7564);
buf BUF1 (N7579, N7561);
and AND3 (N7580, N7576, N6876, N415);
and AND4 (N7581, N7565, N1166, N3689, N487);
or OR3 (N7582, N7566, N6977, N4193);
xor XOR2 (N7583, N7582, N4733);
nor NOR3 (N7584, N7579, N2523, N6292);
and AND4 (N7585, N7552, N3854, N742, N6294);
xor XOR2 (N7586, N7585, N3606);
nand NAND4 (N7587, N7580, N4262, N6735, N4090);
nor NOR4 (N7588, N7578, N7418, N2474, N3267);
and AND4 (N7589, N7587, N6585, N3272, N6024);
nand NAND4 (N7590, N7586, N1926, N7521, N2798);
not NOT1 (N7591, N7584);
or OR2 (N7592, N7575, N757);
and AND3 (N7593, N7583, N3152, N3270);
and AND2 (N7594, N7572, N7123);
and AND4 (N7595, N7589, N6778, N2969, N1553);
or OR4 (N7596, N7593, N1010, N7384, N122);
not NOT1 (N7597, N7592);
or OR4 (N7598, N7567, N724, N7085, N5248);
buf BUF1 (N7599, N7598);
and AND2 (N7600, N7581, N6630);
buf BUF1 (N7601, N7596);
nand NAND2 (N7602, N7600, N5131);
buf BUF1 (N7603, N7601);
nor NOR4 (N7604, N7590, N6520, N7464, N3103);
nor NOR4 (N7605, N7591, N5288, N4226, N4427);
xor XOR2 (N7606, N7594, N6114);
buf BUF1 (N7607, N7603);
not NOT1 (N7608, N7605);
nor NOR2 (N7609, N7595, N1988);
xor XOR2 (N7610, N7599, N531);
not NOT1 (N7611, N7610);
buf BUF1 (N7612, N7577);
nor NOR4 (N7613, N7606, N560, N7302, N3382);
buf BUF1 (N7614, N7613);
nor NOR3 (N7615, N7607, N359, N1905);
not NOT1 (N7616, N7614);
nand NAND4 (N7617, N7612, N1303, N5641, N123);
or OR3 (N7618, N7588, N3170, N7245);
nor NOR3 (N7619, N7604, N4157, N1710);
not NOT1 (N7620, N7616);
nand NAND3 (N7621, N7609, N3944, N442);
and AND2 (N7622, N7608, N950);
not NOT1 (N7623, N7619);
xor XOR2 (N7624, N7611, N5129);
and AND3 (N7625, N7615, N2397, N3890);
nor NOR4 (N7626, N7624, N7236, N3201, N2667);
xor XOR2 (N7627, N7602, N6501);
and AND4 (N7628, N7597, N7104, N2594, N6768);
and AND4 (N7629, N7620, N240, N563, N6294);
and AND2 (N7630, N7618, N4509);
not NOT1 (N7631, N7628);
xor XOR2 (N7632, N7629, N5306);
buf BUF1 (N7633, N7625);
nand NAND4 (N7634, N7623, N2652, N3607, N1467);
nand NAND3 (N7635, N7632, N3925, N7058);
buf BUF1 (N7636, N7630);
buf BUF1 (N7637, N7634);
nand NAND4 (N7638, N7636, N4149, N1096, N2302);
or OR4 (N7639, N7617, N5480, N6732, N1492);
xor XOR2 (N7640, N7622, N3778);
or OR3 (N7641, N7638, N5594, N1669);
and AND4 (N7642, N7631, N6480, N3851, N7630);
nand NAND2 (N7643, N7637, N2579);
not NOT1 (N7644, N7643);
xor XOR2 (N7645, N7621, N2130);
and AND4 (N7646, N7635, N4331, N891, N2187);
not NOT1 (N7647, N7645);
nor NOR2 (N7648, N7627, N6842);
not NOT1 (N7649, N7633);
nor NOR2 (N7650, N7646, N2364);
xor XOR2 (N7651, N7642, N4562);
buf BUF1 (N7652, N7651);
buf BUF1 (N7653, N7644);
and AND2 (N7654, N7639, N850);
or OR3 (N7655, N7626, N4119, N3781);
not NOT1 (N7656, N7652);
not NOT1 (N7657, N7654);
and AND3 (N7658, N7650, N1427, N2402);
nand NAND4 (N7659, N7657, N3772, N6738, N6859);
or OR3 (N7660, N7653, N2298, N5007);
not NOT1 (N7661, N7648);
or OR2 (N7662, N7656, N3099);
xor XOR2 (N7663, N7649, N6062);
not NOT1 (N7664, N7658);
or OR4 (N7665, N7660, N6205, N5043, N2904);
xor XOR2 (N7666, N7647, N883);
nand NAND4 (N7667, N7664, N6208, N2460, N3585);
not NOT1 (N7668, N7661);
nand NAND2 (N7669, N7662, N1726);
buf BUF1 (N7670, N7663);
nand NAND2 (N7671, N7655, N1030);
or OR4 (N7672, N7665, N4268, N7582, N3804);
nand NAND3 (N7673, N7659, N4173, N5562);
xor XOR2 (N7674, N7641, N1806);
or OR2 (N7675, N7668, N6028);
or OR2 (N7676, N7673, N424);
buf BUF1 (N7677, N7669);
nor NOR4 (N7678, N7667, N4786, N7189, N2764);
or OR3 (N7679, N7675, N7219, N6783);
buf BUF1 (N7680, N7679);
buf BUF1 (N7681, N7666);
and AND2 (N7682, N7674, N829);
and AND2 (N7683, N7680, N4499);
nand NAND3 (N7684, N7683, N949, N1797);
and AND4 (N7685, N7677, N6583, N2561, N89);
and AND2 (N7686, N7681, N4744);
not NOT1 (N7687, N7678);
not NOT1 (N7688, N7686);
xor XOR2 (N7689, N7676, N6602);
or OR2 (N7690, N7688, N7345);
nand NAND4 (N7691, N7640, N4668, N977, N6894);
or OR4 (N7692, N7691, N3717, N3555, N3239);
and AND4 (N7693, N7687, N7280, N2139, N3635);
xor XOR2 (N7694, N7684, N1232);
xor XOR2 (N7695, N7671, N6411);
xor XOR2 (N7696, N7689, N3378);
not NOT1 (N7697, N7694);
buf BUF1 (N7698, N7696);
and AND4 (N7699, N7695, N567, N4711, N4697);
xor XOR2 (N7700, N7672, N6489);
not NOT1 (N7701, N7690);
or OR4 (N7702, N7697, N419, N1909, N934);
xor XOR2 (N7703, N7682, N6109);
nand NAND4 (N7704, N7699, N2556, N4552, N2787);
or OR4 (N7705, N7700, N2960, N3531, N982);
nand NAND2 (N7706, N7685, N3366);
buf BUF1 (N7707, N7670);
not NOT1 (N7708, N7703);
not NOT1 (N7709, N7706);
or OR2 (N7710, N7698, N5037);
nor NOR2 (N7711, N7710, N1531);
nor NOR2 (N7712, N7701, N3392);
nor NOR3 (N7713, N7692, N256, N7650);
and AND3 (N7714, N7713, N4945, N5691);
not NOT1 (N7715, N7705);
buf BUF1 (N7716, N7709);
and AND3 (N7717, N7716, N2765, N2945);
not NOT1 (N7718, N7715);
nor NOR3 (N7719, N7717, N1871, N2633);
xor XOR2 (N7720, N7702, N2916);
not NOT1 (N7721, N7707);
nor NOR4 (N7722, N7693, N3622, N7193, N2112);
xor XOR2 (N7723, N7721, N7679);
nor NOR3 (N7724, N7719, N5439, N6459);
not NOT1 (N7725, N7704);
buf BUF1 (N7726, N7724);
xor XOR2 (N7727, N7718, N4971);
nand NAND3 (N7728, N7725, N221, N3421);
or OR4 (N7729, N7727, N5836, N2557, N4099);
not NOT1 (N7730, N7720);
and AND4 (N7731, N7726, N5914, N4397, N741);
or OR4 (N7732, N7714, N2306, N4748, N2320);
nand NAND3 (N7733, N7708, N3972, N3989);
nor NOR3 (N7734, N7712, N2872, N4469);
and AND2 (N7735, N7730, N3732);
buf BUF1 (N7736, N7735);
or OR2 (N7737, N7711, N5408);
nor NOR2 (N7738, N7722, N4419);
buf BUF1 (N7739, N7734);
nand NAND3 (N7740, N7733, N5839, N4340);
or OR3 (N7741, N7738, N572, N4975);
buf BUF1 (N7742, N7729);
nor NOR2 (N7743, N7728, N1757);
nand NAND3 (N7744, N7732, N2447, N3839);
buf BUF1 (N7745, N7723);
xor XOR2 (N7746, N7739, N2445);
xor XOR2 (N7747, N7745, N3376);
xor XOR2 (N7748, N7736, N1377);
or OR3 (N7749, N7741, N4191, N6606);
nand NAND4 (N7750, N7740, N954, N2174, N1922);
and AND4 (N7751, N7731, N323, N7178, N3631);
and AND4 (N7752, N7737, N5273, N3630, N420);
or OR2 (N7753, N7746, N5869);
nand NAND2 (N7754, N7748, N1139);
xor XOR2 (N7755, N7742, N6803);
xor XOR2 (N7756, N7743, N2017);
buf BUF1 (N7757, N7752);
or OR4 (N7758, N7749, N5357, N855, N1236);
and AND4 (N7759, N7754, N801, N5590, N3671);
not NOT1 (N7760, N7758);
not NOT1 (N7761, N7744);
and AND4 (N7762, N7756, N7602, N13, N4432);
buf BUF1 (N7763, N7747);
or OR2 (N7764, N7762, N2984);
buf BUF1 (N7765, N7755);
and AND3 (N7766, N7761, N2466, N6514);
or OR2 (N7767, N7765, N90);
and AND2 (N7768, N7750, N1604);
not NOT1 (N7769, N7766);
xor XOR2 (N7770, N7757, N193);
nor NOR3 (N7771, N7760, N585, N4363);
xor XOR2 (N7772, N7770, N2436);
buf BUF1 (N7773, N7753);
and AND2 (N7774, N7767, N5324);
or OR4 (N7775, N7773, N6397, N2010, N1880);
xor XOR2 (N7776, N7763, N2837);
and AND2 (N7777, N7751, N5050);
buf BUF1 (N7778, N7776);
xor XOR2 (N7779, N7778, N3410);
or OR3 (N7780, N7772, N1599, N6052);
nor NOR3 (N7781, N7779, N659, N2797);
or OR2 (N7782, N7764, N2593);
not NOT1 (N7783, N7781);
nor NOR2 (N7784, N7774, N6624);
buf BUF1 (N7785, N7769);
not NOT1 (N7786, N7777);
nor NOR2 (N7787, N7780, N7698);
not NOT1 (N7788, N7771);
or OR3 (N7789, N7784, N3811, N3772);
and AND4 (N7790, N7786, N2336, N5775, N4751);
or OR3 (N7791, N7787, N7123, N4078);
not NOT1 (N7792, N7789);
or OR3 (N7793, N7791, N5637, N986);
buf BUF1 (N7794, N7790);
nand NAND2 (N7795, N7783, N2724);
not NOT1 (N7796, N7794);
not NOT1 (N7797, N7792);
xor XOR2 (N7798, N7759, N1933);
nand NAND3 (N7799, N7788, N5973, N4506);
nand NAND2 (N7800, N7798, N7648);
buf BUF1 (N7801, N7795);
nor NOR3 (N7802, N7801, N6443, N1762);
or OR2 (N7803, N7793, N4320);
not NOT1 (N7804, N7768);
buf BUF1 (N7805, N7797);
or OR4 (N7806, N7785, N4829, N6383, N1468);
not NOT1 (N7807, N7802);
xor XOR2 (N7808, N7807, N2);
not NOT1 (N7809, N7803);
and AND3 (N7810, N7809, N2432, N858);
or OR4 (N7811, N7782, N2459, N75, N5316);
nand NAND4 (N7812, N7805, N6064, N6468, N2172);
buf BUF1 (N7813, N7775);
buf BUF1 (N7814, N7808);
nor NOR2 (N7815, N7796, N2032);
xor XOR2 (N7816, N7799, N7684);
or OR2 (N7817, N7813, N4350);
nor NOR4 (N7818, N7811, N2184, N2649, N6396);
xor XOR2 (N7819, N7817, N6636);
buf BUF1 (N7820, N7806);
xor XOR2 (N7821, N7814, N1442);
and AND2 (N7822, N7800, N1978);
nor NOR4 (N7823, N7812, N692, N5774, N3760);
xor XOR2 (N7824, N7819, N1364);
and AND4 (N7825, N7822, N6691, N4543, N6342);
nand NAND3 (N7826, N7825, N4474, N4041);
not NOT1 (N7827, N7826);
or OR4 (N7828, N7804, N4986, N4152, N4484);
nand NAND4 (N7829, N7823, N5562, N4050, N2079);
not NOT1 (N7830, N7816);
not NOT1 (N7831, N7828);
not NOT1 (N7832, N7831);
xor XOR2 (N7833, N7832, N1403);
buf BUF1 (N7834, N7824);
or OR3 (N7835, N7827, N5295, N3952);
buf BUF1 (N7836, N7818);
nor NOR2 (N7837, N7830, N4091);
not NOT1 (N7838, N7834);
buf BUF1 (N7839, N7829);
and AND3 (N7840, N7837, N6430, N2599);
nor NOR4 (N7841, N7839, N2090, N7000, N2897);
or OR2 (N7842, N7836, N7130);
not NOT1 (N7843, N7810);
or OR4 (N7844, N7821, N5861, N6027, N321);
or OR3 (N7845, N7841, N3917, N5368);
or OR4 (N7846, N7840, N577, N3627, N538);
nor NOR2 (N7847, N7820, N4641);
buf BUF1 (N7848, N7842);
buf BUF1 (N7849, N7835);
or OR4 (N7850, N7848, N6518, N4988, N2921);
nand NAND2 (N7851, N7844, N5988);
nor NOR2 (N7852, N7833, N7250);
not NOT1 (N7853, N7850);
nand NAND2 (N7854, N7847, N7160);
nand NAND4 (N7855, N7845, N4926, N4046, N6875);
and AND3 (N7856, N7853, N6621, N816);
and AND2 (N7857, N7849, N7849);
and AND3 (N7858, N7855, N5474, N7608);
nand NAND3 (N7859, N7852, N631, N7003);
buf BUF1 (N7860, N7857);
or OR3 (N7861, N7859, N4234, N5332);
nor NOR2 (N7862, N7856, N6954);
buf BUF1 (N7863, N7815);
buf BUF1 (N7864, N7846);
nor NOR4 (N7865, N7854, N6292, N3057, N3993);
nor NOR4 (N7866, N7865, N1116, N2733, N2956);
buf BUF1 (N7867, N7851);
not NOT1 (N7868, N7861);
xor XOR2 (N7869, N7863, N5065);
xor XOR2 (N7870, N7868, N2767);
xor XOR2 (N7871, N7838, N3238);
and AND4 (N7872, N7860, N6940, N2570, N2555);
nor NOR2 (N7873, N7867, N2966);
xor XOR2 (N7874, N7870, N5612);
and AND2 (N7875, N7864, N2097);
not NOT1 (N7876, N7873);
nand NAND3 (N7877, N7876, N5142, N7748);
buf BUF1 (N7878, N7862);
not NOT1 (N7879, N7874);
xor XOR2 (N7880, N7872, N2441);
xor XOR2 (N7881, N7871, N6156);
nand NAND3 (N7882, N7869, N559, N6721);
nor NOR3 (N7883, N7882, N2082, N6731);
buf BUF1 (N7884, N7879);
and AND4 (N7885, N7858, N203, N1173, N2099);
or OR2 (N7886, N7880, N5492);
not NOT1 (N7887, N7878);
nor NOR4 (N7888, N7887, N603, N6764, N2340);
nand NAND4 (N7889, N7883, N7391, N2112, N5229);
or OR2 (N7890, N7888, N1584);
nand NAND2 (N7891, N7875, N5637);
not NOT1 (N7892, N7884);
or OR4 (N7893, N7843, N2672, N5759, N940);
nor NOR3 (N7894, N7886, N7547, N5541);
xor XOR2 (N7895, N7866, N364);
nand NAND4 (N7896, N7877, N4656, N604, N5406);
nand NAND3 (N7897, N7896, N3952, N2470);
not NOT1 (N7898, N7889);
not NOT1 (N7899, N7885);
nor NOR4 (N7900, N7894, N5774, N4071, N3150);
nand NAND3 (N7901, N7881, N1074, N6861);
nor NOR4 (N7902, N7892, N262, N1812, N7331);
xor XOR2 (N7903, N7902, N6644);
nand NAND4 (N7904, N7903, N675, N5285, N4402);
nand NAND2 (N7905, N7904, N1948);
or OR2 (N7906, N7901, N4688);
nor NOR3 (N7907, N7905, N1801, N3304);
or OR3 (N7908, N7900, N4741, N3273);
nor NOR4 (N7909, N7907, N6534, N554, N4976);
nand NAND4 (N7910, N7909, N5159, N2513, N5930);
xor XOR2 (N7911, N7895, N48);
buf BUF1 (N7912, N7911);
or OR4 (N7913, N7910, N5525, N6262, N7900);
xor XOR2 (N7914, N7913, N3974);
buf BUF1 (N7915, N7912);
and AND4 (N7916, N7890, N3005, N869, N1924);
nor NOR2 (N7917, N7916, N3788);
xor XOR2 (N7918, N7899, N5578);
or OR2 (N7919, N7915, N3024);
nor NOR2 (N7920, N7918, N3919);
not NOT1 (N7921, N7893);
xor XOR2 (N7922, N7897, N4656);
not NOT1 (N7923, N7908);
nor NOR3 (N7924, N7919, N4530, N4284);
buf BUF1 (N7925, N7898);
nor NOR3 (N7926, N7914, N2944, N1491);
xor XOR2 (N7927, N7922, N7306);
buf BUF1 (N7928, N7923);
buf BUF1 (N7929, N7926);
xor XOR2 (N7930, N7891, N4615);
not NOT1 (N7931, N7917);
not NOT1 (N7932, N7924);
and AND3 (N7933, N7932, N7579, N6554);
nand NAND2 (N7934, N7929, N370);
nor NOR2 (N7935, N7928, N1789);
buf BUF1 (N7936, N7931);
not NOT1 (N7937, N7930);
xor XOR2 (N7938, N7933, N362);
or OR4 (N7939, N7925, N1205, N239, N5347);
or OR2 (N7940, N7936, N7361);
nand NAND4 (N7941, N7937, N4080, N7630, N4307);
buf BUF1 (N7942, N7921);
or OR2 (N7943, N7941, N710);
nand NAND2 (N7944, N7935, N4012);
not NOT1 (N7945, N7920);
not NOT1 (N7946, N7927);
xor XOR2 (N7947, N7940, N7118);
buf BUF1 (N7948, N7939);
xor XOR2 (N7949, N7947, N7760);
not NOT1 (N7950, N7949);
not NOT1 (N7951, N7943);
buf BUF1 (N7952, N7944);
or OR4 (N7953, N7945, N5791, N7273, N2281);
nand NAND2 (N7954, N7951, N4888);
buf BUF1 (N7955, N7906);
not NOT1 (N7956, N7938);
or OR3 (N7957, N7955, N2328, N5564);
not NOT1 (N7958, N7934);
and AND4 (N7959, N7946, N138, N7586, N82);
nand NAND3 (N7960, N7948, N4656, N1101);
and AND3 (N7961, N7942, N6515, N1502);
buf BUF1 (N7962, N7950);
xor XOR2 (N7963, N7959, N4819);
buf BUF1 (N7964, N7960);
or OR2 (N7965, N7954, N2287);
or OR2 (N7966, N7965, N3591);
or OR3 (N7967, N7961, N1308, N6908);
and AND4 (N7968, N7956, N1776, N7090, N7552);
nand NAND4 (N7969, N7964, N1417, N5270, N5680);
or OR3 (N7970, N7958, N5237, N4600);
nand NAND4 (N7971, N7967, N2720, N727, N1942);
buf BUF1 (N7972, N7971);
xor XOR2 (N7973, N7968, N1146);
nand NAND4 (N7974, N7957, N3243, N989, N3267);
buf BUF1 (N7975, N7972);
or OR2 (N7976, N7966, N7648);
nor NOR4 (N7977, N7953, N884, N6047, N6481);
nand NAND2 (N7978, N7977, N5776);
or OR4 (N7979, N7952, N600, N4730, N2904);
xor XOR2 (N7980, N7970, N3523);
or OR2 (N7981, N7963, N2643);
nor NOR3 (N7982, N7980, N4041, N6750);
or OR4 (N7983, N7974, N2263, N3158, N1643);
nor NOR4 (N7984, N7978, N1008, N5599, N747);
nor NOR2 (N7985, N7975, N1571);
not NOT1 (N7986, N7981);
nor NOR4 (N7987, N7985, N6666, N133, N3614);
not NOT1 (N7988, N7982);
and AND2 (N7989, N7986, N195);
and AND4 (N7990, N7987, N4632, N5381, N6168);
and AND2 (N7991, N7973, N4722);
buf BUF1 (N7992, N7984);
buf BUF1 (N7993, N7991);
and AND3 (N7994, N7969, N6752, N7456);
and AND2 (N7995, N7988, N4094);
buf BUF1 (N7996, N7983);
not NOT1 (N7997, N7992);
xor XOR2 (N7998, N7994, N5389);
buf BUF1 (N7999, N7979);
not NOT1 (N8000, N7996);
xor XOR2 (N8001, N7990, N2667);
or OR4 (N8002, N7976, N5826, N4017, N5015);
xor XOR2 (N8003, N7993, N5177);
or OR2 (N8004, N7962, N4784);
buf BUF1 (N8005, N7997);
not NOT1 (N8006, N8005);
buf BUF1 (N8007, N7998);
xor XOR2 (N8008, N8003, N3122);
nor NOR4 (N8009, N8008, N1538, N4701, N2011);
and AND4 (N8010, N8001, N2772, N6832, N4191);
xor XOR2 (N8011, N8000, N444);
and AND2 (N8012, N7999, N371);
not NOT1 (N8013, N7989);
buf BUF1 (N8014, N8006);
nand NAND4 (N8015, N8014, N2825, N640, N7230);
and AND2 (N8016, N8010, N4531);
nor NOR4 (N8017, N8009, N3127, N3009, N685);
or OR2 (N8018, N8011, N1715);
xor XOR2 (N8019, N8004, N5083);
buf BUF1 (N8020, N7995);
nor NOR4 (N8021, N8015, N6098, N7762, N1378);
not NOT1 (N8022, N8002);
nand NAND4 (N8023, N8022, N426, N462, N1381);
xor XOR2 (N8024, N8020, N2413);
nor NOR2 (N8025, N8024, N1173);
not NOT1 (N8026, N8017);
buf BUF1 (N8027, N8019);
xor XOR2 (N8028, N8021, N3034);
nand NAND3 (N8029, N8025, N6423, N2256);
not NOT1 (N8030, N8007);
and AND3 (N8031, N8012, N3825, N5990);
or OR4 (N8032, N8018, N2955, N7581, N4637);
nor NOR3 (N8033, N8027, N5369, N805);
and AND4 (N8034, N8031, N4499, N4955, N4056);
buf BUF1 (N8035, N8032);
nor NOR2 (N8036, N8034, N808);
not NOT1 (N8037, N8028);
not NOT1 (N8038, N8026);
not NOT1 (N8039, N8029);
and AND3 (N8040, N8037, N4789, N5644);
nand NAND4 (N8041, N8036, N3996, N7364, N1848);
and AND3 (N8042, N8033, N2264, N5300);
nand NAND3 (N8043, N8030, N3538, N3930);
or OR3 (N8044, N8040, N7749, N1325);
nand NAND2 (N8045, N8044, N6343);
buf BUF1 (N8046, N8039);
and AND2 (N8047, N8042, N4310);
or OR2 (N8048, N8013, N1000);
and AND4 (N8049, N8045, N4541, N5038, N2241);
not NOT1 (N8050, N8038);
xor XOR2 (N8051, N8023, N3075);
nand NAND4 (N8052, N8046, N1113, N7183, N6765);
and AND3 (N8053, N8016, N5856, N2046);
xor XOR2 (N8054, N8050, N7384);
and AND4 (N8055, N8051, N1511, N57, N62);
or OR4 (N8056, N8049, N2330, N5939, N827);
not NOT1 (N8057, N8048);
buf BUF1 (N8058, N8043);
xor XOR2 (N8059, N8054, N4031);
nand NAND3 (N8060, N8058, N1465, N4817);
not NOT1 (N8061, N8059);
nand NAND4 (N8062, N8041, N451, N6170, N6745);
not NOT1 (N8063, N8035);
or OR2 (N8064, N8055, N4936);
buf BUF1 (N8065, N8063);
and AND4 (N8066, N8062, N404, N3246, N3273);
or OR3 (N8067, N8066, N4074, N6637);
not NOT1 (N8068, N8064);
or OR2 (N8069, N8056, N6509);
not NOT1 (N8070, N8057);
xor XOR2 (N8071, N8065, N2585);
nor NOR4 (N8072, N8047, N5000, N7697, N3352);
xor XOR2 (N8073, N8069, N7144);
nand NAND2 (N8074, N8072, N1779);
buf BUF1 (N8075, N8053);
and AND3 (N8076, N8052, N3856, N3069);
and AND3 (N8077, N8074, N3881, N3748);
nor NOR4 (N8078, N8076, N7470, N2330, N4235);
buf BUF1 (N8079, N8075);
and AND4 (N8080, N8067, N4465, N4854, N5925);
xor XOR2 (N8081, N8080, N1812);
buf BUF1 (N8082, N8078);
buf BUF1 (N8083, N8068);
nor NOR2 (N8084, N8071, N4411);
buf BUF1 (N8085, N8079);
not NOT1 (N8086, N8077);
nand NAND4 (N8087, N8084, N46, N4818, N7104);
xor XOR2 (N8088, N8060, N3157);
or OR3 (N8089, N8061, N3784, N3582);
or OR2 (N8090, N8073, N575);
not NOT1 (N8091, N8089);
or OR4 (N8092, N8090, N3160, N1869, N1865);
xor XOR2 (N8093, N8082, N4617);
nand NAND4 (N8094, N8093, N4769, N2453, N2902);
and AND2 (N8095, N8087, N4277);
or OR4 (N8096, N8083, N6988, N3668, N3452);
nand NAND2 (N8097, N8094, N3767);
buf BUF1 (N8098, N8097);
nor NOR4 (N8099, N8088, N7811, N1185, N8000);
not NOT1 (N8100, N8070);
and AND2 (N8101, N8095, N2874);
nand NAND4 (N8102, N8099, N1586, N1809, N579);
and AND4 (N8103, N8102, N5126, N3973, N3436);
not NOT1 (N8104, N8091);
and AND3 (N8105, N8081, N4539, N6824);
not NOT1 (N8106, N8100);
or OR4 (N8107, N8092, N2788, N5046, N5593);
nand NAND4 (N8108, N8098, N4566, N4932, N4272);
nand NAND2 (N8109, N8085, N149);
buf BUF1 (N8110, N8107);
not NOT1 (N8111, N8101);
not NOT1 (N8112, N8086);
and AND4 (N8113, N8105, N5389, N4077, N5187);
nand NAND4 (N8114, N8108, N1990, N1236, N7046);
or OR3 (N8115, N8104, N4739, N1455);
and AND3 (N8116, N8112, N7508, N5728);
or OR3 (N8117, N8116, N6006, N505);
nand NAND2 (N8118, N8114, N7461);
and AND3 (N8119, N8096, N4806, N4754);
nor NOR3 (N8120, N8106, N1491, N3945);
buf BUF1 (N8121, N8110);
nand NAND4 (N8122, N8109, N1686, N664, N6830);
not NOT1 (N8123, N8115);
buf BUF1 (N8124, N8113);
not NOT1 (N8125, N8122);
buf BUF1 (N8126, N8119);
or OR3 (N8127, N8126, N322, N6713);
nand NAND2 (N8128, N8124, N8074);
nor NOR3 (N8129, N8123, N2828, N2897);
buf BUF1 (N8130, N8117);
not NOT1 (N8131, N8118);
and AND2 (N8132, N8128, N604);
xor XOR2 (N8133, N8120, N5359);
xor XOR2 (N8134, N8131, N5984);
not NOT1 (N8135, N8103);
buf BUF1 (N8136, N8130);
buf BUF1 (N8137, N8133);
and AND4 (N8138, N8135, N3418, N6537, N1121);
or OR4 (N8139, N8134, N4610, N470, N2801);
nor NOR3 (N8140, N8136, N301, N4531);
nand NAND4 (N8141, N8139, N4009, N4401, N4656);
buf BUF1 (N8142, N8138);
not NOT1 (N8143, N8141);
and AND2 (N8144, N8125, N7686);
nor NOR2 (N8145, N8140, N5875);
not NOT1 (N8146, N8143);
or OR2 (N8147, N8142, N6406);
nor NOR2 (N8148, N8144, N603);
or OR3 (N8149, N8147, N3726, N6766);
buf BUF1 (N8150, N8145);
and AND2 (N8151, N8111, N1015);
nor NOR4 (N8152, N8148, N7539, N1445, N7563);
nor NOR4 (N8153, N8149, N1173, N7012, N1234);
buf BUF1 (N8154, N8121);
nor NOR4 (N8155, N8127, N1147, N2364, N4960);
or OR4 (N8156, N8146, N1403, N7082, N3538);
not NOT1 (N8157, N8151);
and AND4 (N8158, N8132, N7933, N6464, N1011);
not NOT1 (N8159, N8156);
xor XOR2 (N8160, N8159, N424);
buf BUF1 (N8161, N8150);
not NOT1 (N8162, N8160);
not NOT1 (N8163, N8158);
or OR4 (N8164, N8163, N897, N3707, N4261);
nand NAND4 (N8165, N8161, N6285, N5275, N2635);
nand NAND2 (N8166, N8162, N5671);
or OR2 (N8167, N8164, N7046);
nand NAND3 (N8168, N8166, N4307, N6154);
or OR2 (N8169, N8152, N1110);
not NOT1 (N8170, N8155);
or OR3 (N8171, N8153, N1904, N2098);
nand NAND3 (N8172, N8169, N5832, N878);
nor NOR4 (N8173, N8157, N3821, N314, N164);
nand NAND3 (N8174, N8171, N7571, N616);
nand NAND4 (N8175, N8172, N5374, N5618, N6622);
nor NOR3 (N8176, N8168, N6712, N7168);
and AND4 (N8177, N8154, N2355, N4533, N4831);
not NOT1 (N8178, N8173);
not NOT1 (N8179, N8177);
xor XOR2 (N8180, N8175, N3269);
not NOT1 (N8181, N8165);
xor XOR2 (N8182, N8178, N6624);
xor XOR2 (N8183, N8170, N2912);
nor NOR3 (N8184, N8180, N7488, N780);
xor XOR2 (N8185, N8137, N1531);
nor NOR2 (N8186, N8129, N6612);
xor XOR2 (N8187, N8186, N7896);
nor NOR2 (N8188, N8185, N4482);
and AND4 (N8189, N8187, N861, N3787, N366);
and AND4 (N8190, N8188, N4876, N213, N1998);
nor NOR2 (N8191, N8182, N1685);
nand NAND3 (N8192, N8167, N667, N5001);
xor XOR2 (N8193, N8181, N4113);
nand NAND2 (N8194, N8192, N3609);
not NOT1 (N8195, N8189);
nor NOR3 (N8196, N8191, N658, N2107);
and AND2 (N8197, N8176, N372);
buf BUF1 (N8198, N8196);
xor XOR2 (N8199, N8179, N6806);
not NOT1 (N8200, N8193);
or OR3 (N8201, N8183, N6898, N4678);
nor NOR2 (N8202, N8199, N2269);
nor NOR2 (N8203, N8197, N1246);
xor XOR2 (N8204, N8200, N2741);
nand NAND2 (N8205, N8202, N1725);
not NOT1 (N8206, N8190);
not NOT1 (N8207, N8195);
buf BUF1 (N8208, N8198);
nor NOR3 (N8209, N8194, N7527, N5524);
or OR2 (N8210, N8203, N5617);
nor NOR4 (N8211, N8207, N5304, N8039, N1718);
nor NOR2 (N8212, N8211, N3234);
not NOT1 (N8213, N8201);
not NOT1 (N8214, N8210);
or OR4 (N8215, N8213, N4877, N3777, N3894);
and AND2 (N8216, N8212, N4619);
xor XOR2 (N8217, N8214, N126);
and AND2 (N8218, N8206, N2492);
or OR3 (N8219, N8215, N7601, N3013);
not NOT1 (N8220, N8205);
or OR2 (N8221, N8174, N3341);
nand NAND4 (N8222, N8217, N5293, N4848, N5341);
xor XOR2 (N8223, N8216, N5037);
xor XOR2 (N8224, N8223, N4248);
buf BUF1 (N8225, N8219);
not NOT1 (N8226, N8218);
xor XOR2 (N8227, N8204, N130);
and AND2 (N8228, N8184, N187);
xor XOR2 (N8229, N8209, N6788);
or OR4 (N8230, N8229, N5, N7490, N7392);
xor XOR2 (N8231, N8208, N595);
or OR3 (N8232, N8222, N1928, N277);
or OR4 (N8233, N8225, N5162, N4087, N1534);
nor NOR4 (N8234, N8233, N2144, N2160, N4003);
xor XOR2 (N8235, N8220, N608);
nor NOR4 (N8236, N8221, N3095, N691, N6083);
nand NAND2 (N8237, N8231, N6244);
xor XOR2 (N8238, N8234, N7261);
nand NAND4 (N8239, N8230, N6825, N6963, N6128);
not NOT1 (N8240, N8238);
or OR4 (N8241, N8236, N3633, N5297, N1582);
buf BUF1 (N8242, N8224);
not NOT1 (N8243, N8235);
not NOT1 (N8244, N8227);
not NOT1 (N8245, N8239);
or OR3 (N8246, N8240, N275, N5834);
buf BUF1 (N8247, N8237);
nand NAND4 (N8248, N8247, N6077, N578, N919);
nor NOR4 (N8249, N8248, N6607, N510, N432);
nand NAND4 (N8250, N8241, N4161, N2871, N2556);
buf BUF1 (N8251, N8244);
nand NAND3 (N8252, N8245, N4439, N7544);
nand NAND3 (N8253, N8246, N2978, N4696);
nor NOR4 (N8254, N8251, N6280, N1625, N5054);
or OR2 (N8255, N8242, N4325);
nand NAND4 (N8256, N8226, N5168, N5686, N8018);
nand NAND3 (N8257, N8256, N6469, N7871);
or OR3 (N8258, N8255, N1158, N3402);
and AND4 (N8259, N8250, N6302, N228, N5680);
nand NAND4 (N8260, N8254, N2978, N3127, N749);
and AND4 (N8261, N8232, N3258, N2721, N1000);
or OR2 (N8262, N8228, N2329);
not NOT1 (N8263, N8249);
xor XOR2 (N8264, N8253, N7279);
buf BUF1 (N8265, N8264);
not NOT1 (N8266, N8262);
buf BUF1 (N8267, N8261);
or OR4 (N8268, N8257, N905, N4835, N8244);
not NOT1 (N8269, N8259);
nor NOR3 (N8270, N8267, N3272, N6962);
nor NOR4 (N8271, N8252, N5779, N2570, N6122);
xor XOR2 (N8272, N8260, N3637);
or OR4 (N8273, N8268, N371, N6101, N5824);
buf BUF1 (N8274, N8258);
and AND4 (N8275, N8265, N2297, N185, N8011);
buf BUF1 (N8276, N8271);
not NOT1 (N8277, N8272);
xor XOR2 (N8278, N8274, N4893);
buf BUF1 (N8279, N8276);
xor XOR2 (N8280, N8273, N5543);
xor XOR2 (N8281, N8277, N2970);
nand NAND4 (N8282, N8279, N3836, N5697, N5581);
nand NAND2 (N8283, N8269, N7657);
not NOT1 (N8284, N8266);
buf BUF1 (N8285, N8281);
buf BUF1 (N8286, N8283);
or OR4 (N8287, N8282, N6536, N5905, N2843);
nor NOR2 (N8288, N8270, N6244);
or OR2 (N8289, N8280, N3933);
xor XOR2 (N8290, N8286, N3219);
nor NOR2 (N8291, N8243, N1873);
or OR2 (N8292, N8275, N6012);
xor XOR2 (N8293, N8289, N3880);
or OR3 (N8294, N8292, N233, N2241);
nor NOR3 (N8295, N8285, N4061, N1757);
not NOT1 (N8296, N8295);
not NOT1 (N8297, N8294);
nor NOR2 (N8298, N8297, N3330);
nor NOR3 (N8299, N8278, N1599, N6010);
xor XOR2 (N8300, N8288, N4203);
nand NAND2 (N8301, N8298, N4107);
nand NAND3 (N8302, N8293, N6657, N3996);
not NOT1 (N8303, N8291);
not NOT1 (N8304, N8302);
nand NAND4 (N8305, N8301, N3416, N7513, N962);
xor XOR2 (N8306, N8303, N6029);
xor XOR2 (N8307, N8287, N6922);
buf BUF1 (N8308, N8284);
and AND2 (N8309, N8290, N4128);
nand NAND3 (N8310, N8305, N1957, N6787);
or OR2 (N8311, N8308, N1638);
nor NOR4 (N8312, N8304, N5143, N240, N3910);
and AND2 (N8313, N8311, N5265);
not NOT1 (N8314, N8263);
nor NOR2 (N8315, N8314, N5036);
not NOT1 (N8316, N8296);
buf BUF1 (N8317, N8312);
or OR3 (N8318, N8299, N1419, N3132);
nand NAND2 (N8319, N8313, N8049);
xor XOR2 (N8320, N8300, N7492);
nand NAND3 (N8321, N8319, N6523, N7342);
and AND2 (N8322, N8320, N2223);
or OR3 (N8323, N8315, N2157, N3477);
nand NAND3 (N8324, N8322, N1602, N2011);
nor NOR2 (N8325, N8317, N573);
nor NOR4 (N8326, N8325, N6810, N5154, N4790);
xor XOR2 (N8327, N8321, N3358);
nand NAND3 (N8328, N8309, N194, N4739);
nor NOR4 (N8329, N8324, N6401, N6080, N8155);
buf BUF1 (N8330, N8329);
nand NAND4 (N8331, N8323, N7227, N6032, N1628);
or OR2 (N8332, N8328, N2696);
buf BUF1 (N8333, N8310);
buf BUF1 (N8334, N8316);
not NOT1 (N8335, N8326);
and AND2 (N8336, N8333, N375);
or OR3 (N8337, N8335, N7964, N2572);
nor NOR4 (N8338, N8331, N8206, N8196, N888);
xor XOR2 (N8339, N8330, N6998);
xor XOR2 (N8340, N8338, N3466);
nor NOR4 (N8341, N8306, N6959, N1478, N7354);
or OR3 (N8342, N8337, N5772, N4796);
xor XOR2 (N8343, N8318, N5050);
xor XOR2 (N8344, N8327, N7696);
buf BUF1 (N8345, N8344);
not NOT1 (N8346, N8340);
buf BUF1 (N8347, N8341);
nor NOR3 (N8348, N8342, N4238, N324);
buf BUF1 (N8349, N8348);
nor NOR4 (N8350, N8334, N1021, N7392, N1407);
xor XOR2 (N8351, N8345, N1382);
and AND2 (N8352, N8339, N4466);
buf BUF1 (N8353, N8336);
and AND3 (N8354, N8343, N7358, N2503);
nor NOR2 (N8355, N8353, N3746);
or OR3 (N8356, N8332, N7660, N3470);
buf BUF1 (N8357, N8350);
and AND4 (N8358, N8349, N2685, N5157, N238);
nor NOR3 (N8359, N8358, N3030, N2033);
xor XOR2 (N8360, N8352, N7651);
or OR3 (N8361, N8360, N5109, N4999);
or OR3 (N8362, N8361, N443, N3613);
buf BUF1 (N8363, N8346);
buf BUF1 (N8364, N8359);
xor XOR2 (N8365, N8351, N1230);
not NOT1 (N8366, N8307);
nor NOR4 (N8367, N8357, N6379, N7891, N1769);
nand NAND4 (N8368, N8347, N2868, N3109, N2525);
nand NAND3 (N8369, N8365, N3055, N7979);
buf BUF1 (N8370, N8367);
nand NAND2 (N8371, N8368, N5359);
buf BUF1 (N8372, N8370);
buf BUF1 (N8373, N8354);
or OR2 (N8374, N8363, N826);
or OR3 (N8375, N8366, N3936, N2610);
xor XOR2 (N8376, N8364, N5476);
or OR3 (N8377, N8369, N1868, N7023);
xor XOR2 (N8378, N8375, N74);
and AND4 (N8379, N8378, N4409, N4037, N2457);
and AND2 (N8380, N8376, N6537);
and AND4 (N8381, N8373, N4853, N7902, N606);
not NOT1 (N8382, N8380);
or OR3 (N8383, N8379, N4881, N248);
nand NAND3 (N8384, N8362, N4308, N5542);
nand NAND4 (N8385, N8377, N4638, N2550, N8172);
or OR2 (N8386, N8372, N7270);
xor XOR2 (N8387, N8355, N7260);
not NOT1 (N8388, N8387);
buf BUF1 (N8389, N8385);
xor XOR2 (N8390, N8382, N5955);
or OR3 (N8391, N8381, N2463, N1190);
nor NOR3 (N8392, N8374, N1189, N8258);
not NOT1 (N8393, N8383);
nor NOR3 (N8394, N8356, N531, N244);
xor XOR2 (N8395, N8393, N7415);
or OR3 (N8396, N8389, N4959, N721);
and AND3 (N8397, N8394, N7620, N5377);
buf BUF1 (N8398, N8396);
and AND3 (N8399, N8388, N6224, N7361);
not NOT1 (N8400, N8390);
nand NAND4 (N8401, N8386, N469, N4387, N1832);
xor XOR2 (N8402, N8397, N6846);
not NOT1 (N8403, N8395);
and AND3 (N8404, N8399, N5207, N2334);
xor XOR2 (N8405, N8398, N4580);
nand NAND2 (N8406, N8402, N6130);
or OR2 (N8407, N8384, N5668);
or OR2 (N8408, N8404, N1512);
or OR2 (N8409, N8391, N2150);
not NOT1 (N8410, N8400);
buf BUF1 (N8411, N8408);
buf BUF1 (N8412, N8392);
or OR2 (N8413, N8411, N2867);
or OR2 (N8414, N8405, N1379);
not NOT1 (N8415, N8412);
or OR4 (N8416, N8406, N3470, N7513, N7711);
xor XOR2 (N8417, N8371, N3060);
and AND4 (N8418, N8407, N6893, N7553, N6161);
buf BUF1 (N8419, N8409);
nor NOR4 (N8420, N8415, N5236, N3771, N6013);
xor XOR2 (N8421, N8403, N7071);
buf BUF1 (N8422, N8418);
xor XOR2 (N8423, N8422, N5845);
xor XOR2 (N8424, N8401, N1998);
xor XOR2 (N8425, N8414, N3393);
buf BUF1 (N8426, N8421);
or OR2 (N8427, N8424, N6323);
nand NAND2 (N8428, N8423, N594);
buf BUF1 (N8429, N8417);
and AND3 (N8430, N8426, N4740, N3369);
buf BUF1 (N8431, N8419);
nor NOR2 (N8432, N8425, N5374);
not NOT1 (N8433, N8431);
buf BUF1 (N8434, N8413);
nor NOR4 (N8435, N8428, N6546, N7928, N7750);
nor NOR3 (N8436, N8420, N4300, N5786);
nor NOR3 (N8437, N8436, N7290, N1824);
not NOT1 (N8438, N8429);
and AND4 (N8439, N8432, N6287, N7156, N5996);
and AND2 (N8440, N8438, N3800);
nand NAND2 (N8441, N8427, N5220);
xor XOR2 (N8442, N8410, N1152);
xor XOR2 (N8443, N8416, N3150);
nand NAND2 (N8444, N8443, N5007);
nor NOR4 (N8445, N8441, N496, N7965, N5757);
and AND3 (N8446, N8442, N2301, N7592);
not NOT1 (N8447, N8440);
xor XOR2 (N8448, N8434, N282);
not NOT1 (N8449, N8439);
nor NOR3 (N8450, N8437, N3283, N8314);
xor XOR2 (N8451, N8449, N6814);
xor XOR2 (N8452, N8447, N2200);
and AND2 (N8453, N8450, N127);
or OR4 (N8454, N8451, N297, N7741, N6376);
nor NOR4 (N8455, N8448, N3070, N512, N7540);
nor NOR2 (N8456, N8444, N1684);
not NOT1 (N8457, N8445);
nand NAND2 (N8458, N8430, N284);
nor NOR2 (N8459, N8457, N3135);
or OR2 (N8460, N8455, N3609);
buf BUF1 (N8461, N8433);
buf BUF1 (N8462, N8453);
nor NOR3 (N8463, N8454, N5709, N3463);
and AND2 (N8464, N8452, N6258);
nor NOR3 (N8465, N8459, N4572, N3354);
nor NOR3 (N8466, N8464, N5615, N2053);
nor NOR3 (N8467, N8456, N3939, N4686);
xor XOR2 (N8468, N8463, N5853);
and AND4 (N8469, N8458, N6361, N1151, N4474);
xor XOR2 (N8470, N8446, N6131);
buf BUF1 (N8471, N8469);
xor XOR2 (N8472, N8471, N7099);
nand NAND2 (N8473, N8465, N1994);
buf BUF1 (N8474, N8467);
buf BUF1 (N8475, N8466);
and AND3 (N8476, N8475, N5684, N241);
not NOT1 (N8477, N8474);
or OR3 (N8478, N8477, N4024, N4707);
or OR4 (N8479, N8468, N5013, N6601, N3124);
xor XOR2 (N8480, N8461, N4457);
nor NOR3 (N8481, N8435, N4267, N740);
and AND4 (N8482, N8479, N7198, N8459, N1249);
and AND4 (N8483, N8462, N1749, N7558, N6800);
not NOT1 (N8484, N8478);
and AND4 (N8485, N8482, N1217, N5859, N3622);
and AND2 (N8486, N8470, N23);
xor XOR2 (N8487, N8472, N1489);
xor XOR2 (N8488, N8476, N2752);
and AND4 (N8489, N8481, N3403, N3561, N4782);
nor NOR4 (N8490, N8485, N4834, N6356, N7798);
nand NAND4 (N8491, N8490, N6124, N1948, N1873);
nand NAND3 (N8492, N8484, N7693, N701);
buf BUF1 (N8493, N8489);
or OR2 (N8494, N8480, N3742);
or OR2 (N8495, N8473, N2203);
nor NOR3 (N8496, N8494, N1092, N2249);
xor XOR2 (N8497, N8483, N1114);
not NOT1 (N8498, N8488);
nand NAND2 (N8499, N8491, N4405);
nand NAND3 (N8500, N8497, N411, N3024);
and AND4 (N8501, N8487, N5538, N3913, N2105);
buf BUF1 (N8502, N8493);
not NOT1 (N8503, N8498);
buf BUF1 (N8504, N8495);
or OR4 (N8505, N8492, N3106, N1475, N6939);
nand NAND3 (N8506, N8502, N1118, N307);
nand NAND4 (N8507, N8500, N239, N514, N3237);
buf BUF1 (N8508, N8499);
or OR2 (N8509, N8504, N6826);
or OR4 (N8510, N8506, N6826, N2090, N4458);
or OR2 (N8511, N8503, N7926);
nor NOR2 (N8512, N8508, N671);
not NOT1 (N8513, N8486);
nor NOR4 (N8514, N8496, N2873, N6035, N4451);
and AND4 (N8515, N8512, N280, N1284, N3855);
xor XOR2 (N8516, N8514, N1073);
not NOT1 (N8517, N8460);
and AND3 (N8518, N8515, N6687, N5147);
and AND2 (N8519, N8501, N4067);
buf BUF1 (N8520, N8519);
buf BUF1 (N8521, N8510);
and AND3 (N8522, N8505, N6137, N2843);
and AND3 (N8523, N8521, N4581, N3805);
nor NOR3 (N8524, N8511, N1700, N7353);
nor NOR3 (N8525, N8516, N3403, N106);
nor NOR4 (N8526, N8522, N1868, N7934, N5151);
and AND3 (N8527, N8526, N2113, N3951);
or OR4 (N8528, N8518, N3038, N3697, N5713);
xor XOR2 (N8529, N8509, N993);
xor XOR2 (N8530, N8517, N5800);
nor NOR3 (N8531, N8525, N3658, N2612);
xor XOR2 (N8532, N8507, N6018);
xor XOR2 (N8533, N8524, N5928);
buf BUF1 (N8534, N8513);
not NOT1 (N8535, N8529);
and AND2 (N8536, N8531, N7601);
xor XOR2 (N8537, N8534, N8092);
buf BUF1 (N8538, N8530);
buf BUF1 (N8539, N8520);
not NOT1 (N8540, N8532);
nand NAND2 (N8541, N8523, N4576);
xor XOR2 (N8542, N8538, N5031);
xor XOR2 (N8543, N8541, N4456);
nor NOR2 (N8544, N8536, N8254);
nand NAND2 (N8545, N8543, N5329);
nand NAND2 (N8546, N8539, N4998);
or OR4 (N8547, N8537, N521, N8076, N6396);
buf BUF1 (N8548, N8540);
xor XOR2 (N8549, N8542, N5987);
or OR3 (N8550, N8533, N7914, N6430);
or OR2 (N8551, N8528, N7694);
nand NAND3 (N8552, N8547, N6233, N4196);
buf BUF1 (N8553, N8546);
or OR2 (N8554, N8552, N6575);
and AND4 (N8555, N8554, N825, N3217, N7514);
and AND2 (N8556, N8549, N5254);
or OR2 (N8557, N8555, N3811);
or OR2 (N8558, N8545, N1161);
not NOT1 (N8559, N8553);
and AND3 (N8560, N8548, N95, N8149);
nor NOR3 (N8561, N8527, N7561, N3496);
or OR4 (N8562, N8556, N5722, N4450, N1954);
xor XOR2 (N8563, N8560, N7260);
or OR4 (N8564, N8550, N2263, N4950, N4253);
buf BUF1 (N8565, N8535);
and AND3 (N8566, N8558, N745, N6879);
buf BUF1 (N8567, N8566);
nor NOR4 (N8568, N8563, N6727, N1640, N6309);
xor XOR2 (N8569, N8561, N2791);
xor XOR2 (N8570, N8557, N4343);
nand NAND4 (N8571, N8564, N873, N6130, N3045);
and AND3 (N8572, N8544, N8051, N7439);
xor XOR2 (N8573, N8559, N8194);
nor NOR2 (N8574, N8570, N4291);
or OR2 (N8575, N8574, N2396);
or OR2 (N8576, N8567, N347);
xor XOR2 (N8577, N8569, N2810);
and AND2 (N8578, N8575, N3346);
nor NOR2 (N8579, N8562, N6965);
not NOT1 (N8580, N8565);
xor XOR2 (N8581, N8579, N871);
xor XOR2 (N8582, N8580, N7390);
nand NAND2 (N8583, N8581, N2825);
and AND3 (N8584, N8573, N2686, N6789);
nand NAND3 (N8585, N8576, N8377, N1693);
xor XOR2 (N8586, N8578, N247);
xor XOR2 (N8587, N8572, N3796);
or OR2 (N8588, N8583, N3334);
nor NOR3 (N8589, N8582, N440, N5871);
xor XOR2 (N8590, N8551, N7452);
nor NOR4 (N8591, N8590, N3469, N7196, N286);
or OR2 (N8592, N8571, N5798);
nor NOR4 (N8593, N8589, N2398, N345, N6576);
xor XOR2 (N8594, N8568, N3953);
nor NOR3 (N8595, N8588, N4008, N3948);
nor NOR4 (N8596, N8593, N4981, N1393, N1825);
nor NOR2 (N8597, N8595, N1513);
nand NAND4 (N8598, N8586, N1055, N3662, N5768);
not NOT1 (N8599, N8598);
buf BUF1 (N8600, N8599);
and AND2 (N8601, N8594, N7270);
xor XOR2 (N8602, N8577, N52);
buf BUF1 (N8603, N8587);
xor XOR2 (N8604, N8601, N742);
xor XOR2 (N8605, N8591, N873);
and AND3 (N8606, N8596, N737, N4599);
buf BUF1 (N8607, N8592);
buf BUF1 (N8608, N8606);
and AND3 (N8609, N8603, N732, N1889);
buf BUF1 (N8610, N8608);
nand NAND3 (N8611, N8584, N5909, N1750);
buf BUF1 (N8612, N8602);
and AND4 (N8613, N8607, N4002, N4073, N5843);
or OR4 (N8614, N8613, N1444, N261, N5009);
and AND3 (N8615, N8600, N7193, N6826);
nand NAND3 (N8616, N8597, N3636, N1878);
and AND3 (N8617, N8604, N347, N1611);
or OR4 (N8618, N8612, N4113, N3938, N7238);
nand NAND4 (N8619, N8618, N2526, N5045, N2421);
buf BUF1 (N8620, N8609);
or OR2 (N8621, N8620, N5969);
nor NOR2 (N8622, N8621, N722);
or OR2 (N8623, N8615, N485);
xor XOR2 (N8624, N8614, N493);
or OR3 (N8625, N8623, N1707, N192);
or OR2 (N8626, N8625, N3867);
and AND3 (N8627, N8626, N6793, N7798);
nor NOR2 (N8628, N8610, N5235);
xor XOR2 (N8629, N8624, N3014);
nand NAND3 (N8630, N8627, N3684, N5055);
nor NOR2 (N8631, N8617, N2951);
xor XOR2 (N8632, N8611, N4985);
nor NOR2 (N8633, N8605, N2912);
and AND3 (N8634, N8619, N8446, N1016);
or OR3 (N8635, N8628, N7103, N4708);
buf BUF1 (N8636, N8622);
not NOT1 (N8637, N8585);
nand NAND2 (N8638, N8636, N4208);
or OR3 (N8639, N8629, N6485, N4024);
and AND2 (N8640, N8637, N1575);
nand NAND3 (N8641, N8640, N5127, N2682);
buf BUF1 (N8642, N8630);
or OR2 (N8643, N8631, N587);
or OR4 (N8644, N8641, N4578, N4605, N5472);
buf BUF1 (N8645, N8639);
nand NAND4 (N8646, N8633, N829, N2999, N5304);
buf BUF1 (N8647, N8632);
buf BUF1 (N8648, N8638);
xor XOR2 (N8649, N8644, N4941);
and AND3 (N8650, N8647, N2638, N2047);
nor NOR4 (N8651, N8643, N319, N7724, N2761);
buf BUF1 (N8652, N8650);
buf BUF1 (N8653, N8648);
xor XOR2 (N8654, N8652, N1710);
nand NAND3 (N8655, N8642, N3318, N6485);
or OR4 (N8656, N8649, N7178, N3545, N7096);
and AND2 (N8657, N8646, N3612);
not NOT1 (N8658, N8656);
or OR2 (N8659, N8655, N1813);
and AND2 (N8660, N8616, N681);
buf BUF1 (N8661, N8659);
nand NAND3 (N8662, N8651, N8447, N4314);
xor XOR2 (N8663, N8654, N7966);
not NOT1 (N8664, N8660);
and AND3 (N8665, N8657, N1533, N6282);
not NOT1 (N8666, N8645);
buf BUF1 (N8667, N8662);
nand NAND2 (N8668, N8664, N1279);
xor XOR2 (N8669, N8663, N5307);
nand NAND2 (N8670, N8635, N234);
xor XOR2 (N8671, N8665, N8249);
or OR4 (N8672, N8658, N107, N7441, N5101);
or OR3 (N8673, N8668, N5476, N7445);
xor XOR2 (N8674, N8669, N1782);
buf BUF1 (N8675, N8670);
nand NAND3 (N8676, N8675, N434, N5907);
nor NOR3 (N8677, N8673, N6705, N2397);
xor XOR2 (N8678, N8667, N2404);
nor NOR4 (N8679, N8678, N1742, N8241, N4944);
nor NOR2 (N8680, N8666, N4);
xor XOR2 (N8681, N8653, N8144);
nor NOR3 (N8682, N8679, N7400, N6775);
and AND2 (N8683, N8672, N4805);
and AND2 (N8684, N8683, N4255);
not NOT1 (N8685, N8676);
xor XOR2 (N8686, N8677, N6007);
xor XOR2 (N8687, N8671, N6575);
or OR4 (N8688, N8681, N1, N4536, N1028);
not NOT1 (N8689, N8634);
or OR2 (N8690, N8687, N3575);
xor XOR2 (N8691, N8688, N6744);
or OR4 (N8692, N8686, N4676, N8175, N4159);
xor XOR2 (N8693, N8691, N6279);
nand NAND3 (N8694, N8692, N4999, N616);
nand NAND4 (N8695, N8694, N1186, N8228, N3933);
buf BUF1 (N8696, N8680);
and AND4 (N8697, N8695, N7217, N3362, N3446);
or OR3 (N8698, N8697, N2125, N3271);
xor XOR2 (N8699, N8685, N5364);
xor XOR2 (N8700, N8684, N2604);
or OR2 (N8701, N8661, N1176);
xor XOR2 (N8702, N8696, N2013);
buf BUF1 (N8703, N8700);
nand NAND4 (N8704, N8690, N6080, N4499, N1070);
and AND2 (N8705, N8702, N8702);
and AND4 (N8706, N8693, N2470, N7750, N4925);
nand NAND3 (N8707, N8704, N4854, N8465);
buf BUF1 (N8708, N8682);
and AND3 (N8709, N8708, N460, N8020);
buf BUF1 (N8710, N8705);
xor XOR2 (N8711, N8707, N7570);
xor XOR2 (N8712, N8701, N6803);
xor XOR2 (N8713, N8699, N2500);
xor XOR2 (N8714, N8713, N916);
and AND3 (N8715, N8689, N8114, N7280);
not NOT1 (N8716, N8710);
xor XOR2 (N8717, N8674, N3472);
nand NAND4 (N8718, N8703, N3899, N1718, N5260);
or OR3 (N8719, N8715, N8674, N2222);
not NOT1 (N8720, N8717);
buf BUF1 (N8721, N8706);
xor XOR2 (N8722, N8721, N1802);
xor XOR2 (N8723, N8722, N6104);
or OR4 (N8724, N8698, N2916, N7297, N6454);
not NOT1 (N8725, N8724);
nor NOR4 (N8726, N8720, N1037, N7512, N5885);
or OR4 (N8727, N8726, N8655, N2249, N4992);
buf BUF1 (N8728, N8712);
nand NAND3 (N8729, N8723, N6481, N6008);
xor XOR2 (N8730, N8711, N1376);
buf BUF1 (N8731, N8728);
or OR3 (N8732, N8714, N987, N7819);
nand NAND4 (N8733, N8732, N4117, N790, N5864);
xor XOR2 (N8734, N8733, N3058);
xor XOR2 (N8735, N8716, N5017);
buf BUF1 (N8736, N8735);
not NOT1 (N8737, N8727);
xor XOR2 (N8738, N8729, N8581);
nor NOR3 (N8739, N8737, N4157, N2866);
or OR4 (N8740, N8731, N3731, N4452, N5550);
not NOT1 (N8741, N8739);
buf BUF1 (N8742, N8736);
xor XOR2 (N8743, N8730, N6887);
and AND4 (N8744, N8743, N808, N642, N7236);
nor NOR2 (N8745, N8738, N929);
nor NOR4 (N8746, N8719, N2066, N7447, N6945);
or OR2 (N8747, N8742, N7866);
buf BUF1 (N8748, N8718);
nor NOR2 (N8749, N8746, N1735);
buf BUF1 (N8750, N8725);
xor XOR2 (N8751, N8734, N5803);
buf BUF1 (N8752, N8741);
and AND4 (N8753, N8752, N801, N7912, N3787);
not NOT1 (N8754, N8753);
not NOT1 (N8755, N8740);
nor NOR2 (N8756, N8754, N2246);
or OR2 (N8757, N8747, N6515);
not NOT1 (N8758, N8744);
nor NOR3 (N8759, N8749, N3869, N607);
nand NAND3 (N8760, N8751, N816, N5182);
nor NOR3 (N8761, N8750, N4151, N6173);
xor XOR2 (N8762, N8758, N3592);
not NOT1 (N8763, N8761);
buf BUF1 (N8764, N8755);
xor XOR2 (N8765, N8756, N7462);
nor NOR2 (N8766, N8762, N3888);
nand NAND2 (N8767, N8763, N56);
not NOT1 (N8768, N8766);
and AND4 (N8769, N8757, N1586, N7000, N3520);
not NOT1 (N8770, N8769);
and AND3 (N8771, N8748, N2769, N6144);
nand NAND3 (N8772, N8759, N5445, N7165);
not NOT1 (N8773, N8709);
nand NAND4 (N8774, N8765, N5052, N3513, N7236);
xor XOR2 (N8775, N8772, N5087);
not NOT1 (N8776, N8775);
not NOT1 (N8777, N8774);
and AND2 (N8778, N8760, N567);
buf BUF1 (N8779, N8776);
nand NAND3 (N8780, N8777, N4990, N1602);
nand NAND2 (N8781, N8780, N2083);
buf BUF1 (N8782, N8773);
nor NOR4 (N8783, N8778, N3761, N5111, N444);
or OR3 (N8784, N8783, N4865, N4329);
or OR2 (N8785, N8767, N8084);
nand NAND2 (N8786, N8785, N7332);
nor NOR2 (N8787, N8779, N991);
or OR4 (N8788, N8782, N3018, N1969, N8728);
nand NAND4 (N8789, N8787, N7256, N3020, N530);
nand NAND3 (N8790, N8764, N6241, N3465);
xor XOR2 (N8791, N8745, N3678);
nor NOR4 (N8792, N8790, N2514, N3554, N1658);
or OR2 (N8793, N8786, N347);
not NOT1 (N8794, N8788);
not NOT1 (N8795, N8794);
nand NAND3 (N8796, N8771, N3252, N552);
xor XOR2 (N8797, N8792, N5464);
nor NOR4 (N8798, N8793, N5781, N6797, N973);
xor XOR2 (N8799, N8791, N5227);
nand NAND4 (N8800, N8797, N2081, N638, N2608);
buf BUF1 (N8801, N8768);
nor NOR3 (N8802, N8799, N8381, N2531);
not NOT1 (N8803, N8784);
and AND2 (N8804, N8800, N3733);
nor NOR3 (N8805, N8796, N5384, N8636);
buf BUF1 (N8806, N8770);
and AND2 (N8807, N8806, N8566);
nor NOR2 (N8808, N8802, N3228);
xor XOR2 (N8809, N8795, N1640);
not NOT1 (N8810, N8789);
nand NAND2 (N8811, N8808, N6544);
not NOT1 (N8812, N8781);
or OR4 (N8813, N8810, N8665, N8023, N5882);
and AND3 (N8814, N8811, N4893, N950);
buf BUF1 (N8815, N8812);
buf BUF1 (N8816, N8809);
nand NAND2 (N8817, N8807, N8429);
nand NAND2 (N8818, N8813, N5013);
xor XOR2 (N8819, N8817, N7181);
xor XOR2 (N8820, N8798, N3852);
not NOT1 (N8821, N8801);
nor NOR2 (N8822, N8818, N4071);
nor NOR3 (N8823, N8815, N6386, N4096);
buf BUF1 (N8824, N8805);
buf BUF1 (N8825, N8823);
nor NOR2 (N8826, N8819, N3417);
and AND2 (N8827, N8820, N6075);
buf BUF1 (N8828, N8804);
or OR2 (N8829, N8827, N6861);
nor NOR3 (N8830, N8829, N5483, N7400);
and AND4 (N8831, N8803, N3551, N6721, N2827);
buf BUF1 (N8832, N8816);
buf BUF1 (N8833, N8830);
buf BUF1 (N8834, N8828);
or OR4 (N8835, N8821, N4708, N7576, N4401);
buf BUF1 (N8836, N8834);
buf BUF1 (N8837, N8835);
buf BUF1 (N8838, N8837);
xor XOR2 (N8839, N8825, N4354);
and AND2 (N8840, N8836, N2131);
and AND4 (N8841, N8833, N359, N4691, N6451);
buf BUF1 (N8842, N8814);
and AND2 (N8843, N8842, N7368);
nor NOR4 (N8844, N8839, N6928, N880, N2673);
xor XOR2 (N8845, N8824, N194);
nor NOR4 (N8846, N8844, N1068, N3222, N6863);
nand NAND4 (N8847, N8846, N2646, N7050, N8324);
xor XOR2 (N8848, N8845, N449);
nor NOR3 (N8849, N8831, N2220, N8051);
not NOT1 (N8850, N8841);
xor XOR2 (N8851, N8822, N4196);
not NOT1 (N8852, N8849);
not NOT1 (N8853, N8848);
not NOT1 (N8854, N8847);
buf BUF1 (N8855, N8838);
nand NAND3 (N8856, N8853, N140, N4153);
xor XOR2 (N8857, N8843, N6594);
and AND4 (N8858, N8826, N4250, N3544, N7475);
nand NAND4 (N8859, N8856, N123, N2631, N4508);
nor NOR2 (N8860, N8855, N8608);
nor NOR2 (N8861, N8858, N6181);
not NOT1 (N8862, N8840);
xor XOR2 (N8863, N8861, N6677);
and AND3 (N8864, N8832, N6276, N7780);
and AND3 (N8865, N8859, N7256, N473);
nor NOR2 (N8866, N8864, N7482);
xor XOR2 (N8867, N8866, N6144);
xor XOR2 (N8868, N8851, N600);
and AND2 (N8869, N8860, N8233);
nor NOR3 (N8870, N8850, N1885, N2909);
nand NAND3 (N8871, N8852, N4129, N1197);
nand NAND4 (N8872, N8870, N3872, N7325, N5306);
nand NAND4 (N8873, N8868, N7598, N8487, N395);
or OR3 (N8874, N8871, N8394, N5303);
nand NAND2 (N8875, N8872, N1822);
and AND3 (N8876, N8874, N549, N8751);
xor XOR2 (N8877, N8863, N7874);
nor NOR4 (N8878, N8875, N8846, N2110, N8111);
nand NAND3 (N8879, N8862, N6620, N2856);
nand NAND4 (N8880, N8877, N4767, N3370, N563);
buf BUF1 (N8881, N8880);
buf BUF1 (N8882, N8869);
nand NAND4 (N8883, N8881, N1975, N8433, N8766);
or OR2 (N8884, N8882, N6959);
xor XOR2 (N8885, N8867, N4601);
nand NAND3 (N8886, N8876, N1427, N7827);
or OR3 (N8887, N8873, N1863, N3445);
xor XOR2 (N8888, N8886, N6269);
not NOT1 (N8889, N8857);
not NOT1 (N8890, N8879);
buf BUF1 (N8891, N8854);
nand NAND2 (N8892, N8885, N6658);
nand NAND4 (N8893, N8888, N1828, N5033, N4328);
or OR2 (N8894, N8892, N8829);
nand NAND3 (N8895, N8865, N4086, N91);
nor NOR4 (N8896, N8887, N4311, N5778, N6828);
or OR4 (N8897, N8891, N4655, N4656, N7600);
or OR2 (N8898, N8889, N172);
not NOT1 (N8899, N8897);
not NOT1 (N8900, N8898);
or OR4 (N8901, N8895, N1364, N140, N4498);
not NOT1 (N8902, N8884);
buf BUF1 (N8903, N8902);
not NOT1 (N8904, N8903);
nand NAND3 (N8905, N8894, N7097, N681);
nand NAND3 (N8906, N8901, N1213, N4943);
or OR2 (N8907, N8883, N558);
not NOT1 (N8908, N8893);
not NOT1 (N8909, N8907);
buf BUF1 (N8910, N8896);
not NOT1 (N8911, N8906);
xor XOR2 (N8912, N8899, N5890);
buf BUF1 (N8913, N8912);
or OR3 (N8914, N8909, N5707, N7457);
nor NOR3 (N8915, N8913, N203, N7149);
nor NOR2 (N8916, N8911, N8135);
buf BUF1 (N8917, N8905);
and AND3 (N8918, N8915, N4333, N7485);
and AND2 (N8919, N8914, N3131);
xor XOR2 (N8920, N8904, N3467);
nand NAND4 (N8921, N8920, N5163, N4508, N1566);
and AND4 (N8922, N8900, N4018, N4028, N5982);
not NOT1 (N8923, N8918);
xor XOR2 (N8924, N8878, N5139);
xor XOR2 (N8925, N8922, N4284);
nor NOR4 (N8926, N8921, N1073, N3225, N6530);
nor NOR2 (N8927, N8908, N7477);
or OR3 (N8928, N8925, N8861, N8365);
nor NOR4 (N8929, N8919, N4439, N7916, N3947);
buf BUF1 (N8930, N8928);
nand NAND3 (N8931, N8923, N5204, N1592);
buf BUF1 (N8932, N8890);
not NOT1 (N8933, N8917);
not NOT1 (N8934, N8930);
and AND4 (N8935, N8910, N3818, N3372, N2800);
nand NAND3 (N8936, N8916, N106, N1338);
or OR2 (N8937, N8924, N869);
not NOT1 (N8938, N8929);
nand NAND3 (N8939, N8926, N1655, N4397);
nand NAND2 (N8940, N8935, N2206);
buf BUF1 (N8941, N8934);
buf BUF1 (N8942, N8931);
nor NOR2 (N8943, N8937, N6699);
not NOT1 (N8944, N8940);
buf BUF1 (N8945, N8933);
or OR3 (N8946, N8927, N6277, N135);
not NOT1 (N8947, N8932);
nand NAND4 (N8948, N8938, N7105, N8939, N3610);
nand NAND3 (N8949, N4149, N6015, N5978);
and AND4 (N8950, N8949, N7532, N5664, N6100);
nor NOR3 (N8951, N8942, N2400, N5093);
nor NOR4 (N8952, N8944, N8313, N6394, N1475);
buf BUF1 (N8953, N8947);
nand NAND4 (N8954, N8951, N3495, N4647, N2936);
buf BUF1 (N8955, N8950);
nor NOR2 (N8956, N8946, N440);
buf BUF1 (N8957, N8941);
or OR2 (N8958, N8954, N1372);
nand NAND4 (N8959, N8955, N7580, N8264, N1800);
xor XOR2 (N8960, N8952, N1834);
not NOT1 (N8961, N8960);
or OR4 (N8962, N8943, N1614, N6097, N6783);
not NOT1 (N8963, N8962);
nor NOR3 (N8964, N8956, N6883, N5218);
not NOT1 (N8965, N8953);
buf BUF1 (N8966, N8948);
and AND2 (N8967, N8957, N7448);
not NOT1 (N8968, N8945);
xor XOR2 (N8969, N8968, N4403);
buf BUF1 (N8970, N8969);
or OR4 (N8971, N8966, N1793, N3108, N5693);
xor XOR2 (N8972, N8936, N2591);
and AND3 (N8973, N8972, N4330, N8104);
buf BUF1 (N8974, N8965);
nor NOR4 (N8975, N8973, N2395, N290, N340);
xor XOR2 (N8976, N8971, N8138);
and AND3 (N8977, N8970, N8097, N6299);
not NOT1 (N8978, N8964);
and AND3 (N8979, N8975, N3415, N5296);
buf BUF1 (N8980, N8967);
buf BUF1 (N8981, N8963);
xor XOR2 (N8982, N8979, N7570);
buf BUF1 (N8983, N8959);
not NOT1 (N8984, N8983);
not NOT1 (N8985, N8980);
and AND4 (N8986, N8974, N6262, N261, N6690);
not NOT1 (N8987, N8961);
and AND4 (N8988, N8976, N5074, N6660, N8839);
not NOT1 (N8989, N8984);
and AND2 (N8990, N8978, N5289);
or OR4 (N8991, N8985, N7155, N8701, N6370);
nor NOR4 (N8992, N8977, N4787, N8661, N4038);
nor NOR2 (N8993, N8989, N5520);
nor NOR3 (N8994, N8987, N2058, N4286);
xor XOR2 (N8995, N8981, N1461);
nor NOR4 (N8996, N8982, N4004, N7558, N1391);
and AND3 (N8997, N8988, N1992, N2222);
buf BUF1 (N8998, N8990);
or OR3 (N8999, N8997, N4000, N8010);
and AND4 (N9000, N8995, N7263, N7069, N5634);
not NOT1 (N9001, N8986);
or OR4 (N9002, N8999, N5607, N2592, N3035);
and AND3 (N9003, N8996, N5129, N7640);
and AND3 (N9004, N8958, N3728, N7574);
not NOT1 (N9005, N8993);
or OR3 (N9006, N9004, N2194, N2814);
or OR4 (N9007, N9002, N8406, N5856, N949);
nand NAND3 (N9008, N8992, N8438, N6737);
buf BUF1 (N9009, N9008);
not NOT1 (N9010, N9001);
or OR4 (N9011, N8994, N190, N4403, N3531);
xor XOR2 (N9012, N9000, N4772);
nand NAND3 (N9013, N9012, N620, N6166);
nor NOR4 (N9014, N9003, N6661, N2126, N2071);
nor NOR4 (N9015, N9013, N8742, N7242, N1199);
xor XOR2 (N9016, N9014, N2730);
or OR3 (N9017, N9009, N8983, N2519);
and AND3 (N9018, N9017, N3279, N2938);
nand NAND4 (N9019, N9016, N4969, N6892, N8451);
buf BUF1 (N9020, N9007);
or OR3 (N9021, N9020, N1548, N7590);
buf BUF1 (N9022, N9011);
nand NAND4 (N9023, N9021, N7462, N91, N5972);
buf BUF1 (N9024, N9015);
or OR3 (N9025, N9018, N954, N8608);
nand NAND4 (N9026, N8991, N7905, N4985, N8909);
not NOT1 (N9027, N9025);
nand NAND2 (N9028, N9022, N7953);
buf BUF1 (N9029, N9027);
not NOT1 (N9030, N9028);
not NOT1 (N9031, N9019);
buf BUF1 (N9032, N9024);
buf BUF1 (N9033, N9032);
xor XOR2 (N9034, N9026, N6387);
or OR3 (N9035, N9034, N5399, N6308);
buf BUF1 (N9036, N9033);
and AND3 (N9037, N9036, N4108, N752);
buf BUF1 (N9038, N9031);
xor XOR2 (N9039, N9030, N3927);
buf BUF1 (N9040, N9010);
nand NAND2 (N9041, N9037, N814);
not NOT1 (N9042, N9038);
buf BUF1 (N9043, N9039);
nor NOR2 (N9044, N9029, N5844);
buf BUF1 (N9045, N9040);
not NOT1 (N9046, N9035);
or OR2 (N9047, N9045, N6743);
and AND3 (N9048, N9005, N6523, N3111);
nand NAND4 (N9049, N9047, N5656, N6869, N2082);
not NOT1 (N9050, N8998);
not NOT1 (N9051, N9044);
or OR2 (N9052, N9006, N7952);
nor NOR2 (N9053, N9050, N4922);
xor XOR2 (N9054, N9046, N8795);
and AND4 (N9055, N9054, N4232, N8510, N2568);
nor NOR3 (N9056, N9053, N1740, N5494);
nand NAND2 (N9057, N9052, N4786);
not NOT1 (N9058, N9049);
xor XOR2 (N9059, N9058, N2018);
not NOT1 (N9060, N9055);
and AND4 (N9061, N9051, N8010, N3823, N4316);
xor XOR2 (N9062, N9056, N8782);
xor XOR2 (N9063, N9023, N6936);
or OR4 (N9064, N9062, N7050, N406, N4551);
and AND2 (N9065, N9060, N57);
and AND4 (N9066, N9061, N5805, N3340, N2866);
nor NOR3 (N9067, N9066, N1824, N3704);
xor XOR2 (N9068, N9067, N6110);
or OR2 (N9069, N9064, N1660);
xor XOR2 (N9070, N9069, N3944);
nand NAND2 (N9071, N9048, N163);
and AND2 (N9072, N9065, N8205);
or OR3 (N9073, N9071, N3969, N4392);
and AND3 (N9074, N9073, N3369, N3244);
and AND2 (N9075, N9072, N2462);
not NOT1 (N9076, N9075);
or OR2 (N9077, N9042, N1923);
or OR4 (N9078, N9076, N81, N5526, N2956);
not NOT1 (N9079, N9043);
nand NAND4 (N9080, N9059, N1421, N6328, N8288);
and AND2 (N9081, N9041, N2813);
nand NAND3 (N9082, N9057, N8540, N6604);
xor XOR2 (N9083, N9081, N1616);
nand NAND3 (N9084, N9080, N3067, N685);
buf BUF1 (N9085, N9078);
nand NAND3 (N9086, N9084, N6812, N6054);
buf BUF1 (N9087, N9074);
nor NOR2 (N9088, N9085, N3678);
buf BUF1 (N9089, N9079);
buf BUF1 (N9090, N9068);
xor XOR2 (N9091, N9086, N6755);
and AND3 (N9092, N9077, N2486, N2880);
nor NOR2 (N9093, N9090, N8415);
nor NOR2 (N9094, N9092, N1116);
or OR4 (N9095, N9070, N4683, N6251, N3442);
not NOT1 (N9096, N9094);
buf BUF1 (N9097, N9091);
nand NAND2 (N9098, N9096, N2031);
nor NOR4 (N9099, N9087, N3173, N3924, N4043);
xor XOR2 (N9100, N9088, N4492);
nand NAND4 (N9101, N9100, N906, N6180, N1516);
nor NOR3 (N9102, N9099, N687, N8396);
nand NAND4 (N9103, N9095, N6242, N1836, N649);
and AND4 (N9104, N9102, N5979, N7576, N1614);
not NOT1 (N9105, N9097);
nand NAND3 (N9106, N9089, N3142, N4728);
buf BUF1 (N9107, N9101);
buf BUF1 (N9108, N9063);
nor NOR4 (N9109, N9082, N7073, N1659, N8308);
buf BUF1 (N9110, N9104);
or OR3 (N9111, N9105, N5430, N3699);
buf BUF1 (N9112, N9107);
or OR3 (N9113, N9098, N5042, N221);
not NOT1 (N9114, N9106);
and AND4 (N9115, N9108, N2539, N6058, N5511);
and AND4 (N9116, N9110, N8377, N7778, N6539);
or OR3 (N9117, N9114, N5159, N3976);
nand NAND2 (N9118, N9116, N8543);
or OR2 (N9119, N9109, N1016);
buf BUF1 (N9120, N9117);
nor NOR4 (N9121, N9083, N4256, N3213, N6326);
xor XOR2 (N9122, N9119, N7472);
and AND2 (N9123, N9103, N4635);
nand NAND3 (N9124, N9111, N10, N5145);
and AND2 (N9125, N9115, N8112);
nor NOR3 (N9126, N9112, N7890, N746);
buf BUF1 (N9127, N9126);
or OR2 (N9128, N9118, N8870);
not NOT1 (N9129, N9124);
and AND4 (N9130, N9122, N1098, N8805, N7330);
buf BUF1 (N9131, N9127);
nand NAND2 (N9132, N9125, N5217);
not NOT1 (N9133, N9113);
nor NOR3 (N9134, N9132, N5640, N5395);
nand NAND2 (N9135, N9123, N2932);
and AND3 (N9136, N9131, N8108, N7162);
and AND2 (N9137, N9129, N4760);
not NOT1 (N9138, N9135);
not NOT1 (N9139, N9093);
nor NOR4 (N9140, N9136, N1747, N4586, N8458);
not NOT1 (N9141, N9121);
and AND2 (N9142, N9141, N9039);
and AND3 (N9143, N9128, N7543, N5169);
and AND2 (N9144, N9138, N6557);
buf BUF1 (N9145, N9143);
not NOT1 (N9146, N9139);
and AND2 (N9147, N9145, N7641);
buf BUF1 (N9148, N9120);
xor XOR2 (N9149, N9147, N3685);
and AND2 (N9150, N9130, N6080);
and AND2 (N9151, N9149, N3139);
nor NOR4 (N9152, N9137, N4732, N6470, N2316);
buf BUF1 (N9153, N9146);
and AND3 (N9154, N9140, N2701, N2289);
xor XOR2 (N9155, N9144, N1367);
xor XOR2 (N9156, N9154, N3793);
not NOT1 (N9157, N9134);
not NOT1 (N9158, N9153);
not NOT1 (N9159, N9157);
xor XOR2 (N9160, N9156, N4463);
buf BUF1 (N9161, N9142);
buf BUF1 (N9162, N9161);
or OR4 (N9163, N9162, N6057, N1250, N4062);
nand NAND4 (N9164, N9160, N7738, N3011, N9112);
or OR4 (N9165, N9152, N1422, N3636, N4123);
nor NOR3 (N9166, N9158, N1195, N8345);
or OR2 (N9167, N9166, N718);
and AND4 (N9168, N9159, N6161, N4815, N5067);
or OR2 (N9169, N9150, N3825);
not NOT1 (N9170, N9167);
or OR2 (N9171, N9151, N5379);
nor NOR4 (N9172, N9168, N2556, N7089, N2912);
xor XOR2 (N9173, N9172, N5540);
or OR2 (N9174, N9133, N8248);
buf BUF1 (N9175, N9155);
and AND2 (N9176, N9169, N5029);
or OR2 (N9177, N9171, N3682);
not NOT1 (N9178, N9165);
xor XOR2 (N9179, N9173, N8937);
buf BUF1 (N9180, N9163);
nand NAND3 (N9181, N9170, N104, N6809);
and AND4 (N9182, N9179, N4338, N1468, N8052);
and AND2 (N9183, N9180, N4088);
or OR2 (N9184, N9177, N5674);
nand NAND3 (N9185, N9148, N8155, N6515);
nor NOR2 (N9186, N9175, N1525);
buf BUF1 (N9187, N9182);
nand NAND4 (N9188, N9181, N2497, N4169, N8764);
xor XOR2 (N9189, N9184, N4294);
and AND2 (N9190, N9188, N8993);
nand NAND2 (N9191, N9187, N2351);
not NOT1 (N9192, N9174);
and AND3 (N9193, N9185, N144, N2851);
buf BUF1 (N9194, N9193);
nand NAND2 (N9195, N9183, N1735);
and AND2 (N9196, N9186, N3676);
xor XOR2 (N9197, N9178, N6581);
nor NOR2 (N9198, N9194, N198);
buf BUF1 (N9199, N9191);
buf BUF1 (N9200, N9196);
and AND4 (N9201, N9164, N5961, N7496, N2049);
not NOT1 (N9202, N9190);
nand NAND4 (N9203, N9176, N4429, N5782, N5399);
not NOT1 (N9204, N9203);
or OR4 (N9205, N9204, N8983, N4245, N8048);
nand NAND4 (N9206, N9201, N6135, N8942, N454);
xor XOR2 (N9207, N9199, N5100);
or OR4 (N9208, N9206, N8000, N9050, N6192);
buf BUF1 (N9209, N9200);
nand NAND2 (N9210, N9198, N4039);
not NOT1 (N9211, N9195);
nand NAND4 (N9212, N9211, N6753, N4846, N915);
and AND4 (N9213, N9212, N6759, N9157, N4050);
nand NAND4 (N9214, N9205, N7813, N3359, N4939);
nor NOR4 (N9215, N9209, N6205, N5766, N2964);
or OR3 (N9216, N9189, N1200, N4033);
buf BUF1 (N9217, N9207);
and AND2 (N9218, N9202, N392);
xor XOR2 (N9219, N9218, N3641);
not NOT1 (N9220, N9215);
buf BUF1 (N9221, N9217);
nand NAND2 (N9222, N9208, N5576);
xor XOR2 (N9223, N9210, N1050);
xor XOR2 (N9224, N9214, N9169);
xor XOR2 (N9225, N9197, N3398);
nand NAND4 (N9226, N9213, N6212, N8074, N8197);
xor XOR2 (N9227, N9225, N3024);
or OR4 (N9228, N9220, N2612, N7961, N6280);
not NOT1 (N9229, N9226);
buf BUF1 (N9230, N9224);
nor NOR3 (N9231, N9228, N1864, N3630);
and AND2 (N9232, N9219, N7414);
nand NAND3 (N9233, N9192, N7984, N2721);
xor XOR2 (N9234, N9231, N1341);
nor NOR3 (N9235, N9223, N547, N2226);
xor XOR2 (N9236, N9221, N723);
or OR4 (N9237, N9232, N8476, N3555, N4133);
nand NAND3 (N9238, N9235, N6589, N8645);
nor NOR3 (N9239, N9237, N3900, N2237);
buf BUF1 (N9240, N9234);
nand NAND4 (N9241, N9227, N905, N1230, N2950);
buf BUF1 (N9242, N9239);
and AND2 (N9243, N9230, N7939);
buf BUF1 (N9244, N9242);
not NOT1 (N9245, N9244);
not NOT1 (N9246, N9229);
and AND2 (N9247, N9240, N1312);
or OR2 (N9248, N9247, N5186);
or OR2 (N9249, N9236, N485);
nor NOR3 (N9250, N9238, N3704, N8384);
buf BUF1 (N9251, N9248);
buf BUF1 (N9252, N9246);
nor NOR4 (N9253, N9250, N7428, N4751, N5324);
or OR3 (N9254, N9216, N6747, N5146);
and AND2 (N9255, N9233, N707);
xor XOR2 (N9256, N9243, N5971);
nor NOR3 (N9257, N9251, N32, N6647);
or OR3 (N9258, N9254, N5818, N197);
buf BUF1 (N9259, N9256);
xor XOR2 (N9260, N9259, N8485);
not NOT1 (N9261, N9241);
buf BUF1 (N9262, N9249);
or OR3 (N9263, N9252, N6946, N2627);
nand NAND3 (N9264, N9260, N7005, N7846);
nand NAND4 (N9265, N9261, N8038, N7593, N4550);
not NOT1 (N9266, N9264);
xor XOR2 (N9267, N9266, N7777);
xor XOR2 (N9268, N9253, N549);
or OR3 (N9269, N9267, N172, N1416);
and AND2 (N9270, N9255, N3101);
not NOT1 (N9271, N9262);
nand NAND3 (N9272, N9270, N8922, N9123);
nand NAND4 (N9273, N9263, N711, N5026, N2780);
nor NOR3 (N9274, N9271, N7769, N8079);
nor NOR4 (N9275, N9272, N4283, N8366, N7960);
nand NAND3 (N9276, N9274, N5760, N6414);
buf BUF1 (N9277, N9268);
not NOT1 (N9278, N9276);
or OR2 (N9279, N9257, N7177);
nand NAND4 (N9280, N9273, N7824, N7633, N9263);
and AND4 (N9281, N9278, N2888, N6058, N2917);
or OR3 (N9282, N9265, N8445, N8197);
nand NAND3 (N9283, N9279, N2676, N4950);
buf BUF1 (N9284, N9277);
xor XOR2 (N9285, N9269, N2704);
xor XOR2 (N9286, N9258, N5696);
xor XOR2 (N9287, N9245, N7295);
nand NAND2 (N9288, N9222, N8583);
or OR3 (N9289, N9281, N1156, N8069);
xor XOR2 (N9290, N9289, N1836);
or OR3 (N9291, N9285, N3611, N5316);
xor XOR2 (N9292, N9286, N2855);
buf BUF1 (N9293, N9287);
or OR2 (N9294, N9290, N6485);
nor NOR2 (N9295, N9280, N7828);
and AND2 (N9296, N9295, N3471);
nor NOR2 (N9297, N9296, N4582);
nand NAND2 (N9298, N9293, N3391);
and AND2 (N9299, N9297, N2884);
not NOT1 (N9300, N9298);
xor XOR2 (N9301, N9288, N4632);
and AND4 (N9302, N9300, N6045, N2094, N782);
and AND2 (N9303, N9291, N3042);
or OR3 (N9304, N9284, N1342, N5284);
nor NOR4 (N9305, N9294, N49, N5602, N5277);
nand NAND3 (N9306, N9305, N9066, N5463);
buf BUF1 (N9307, N9303);
buf BUF1 (N9308, N9283);
xor XOR2 (N9309, N9275, N457);
xor XOR2 (N9310, N9308, N6757);
or OR4 (N9311, N9306, N4471, N4101, N3275);
xor XOR2 (N9312, N9299, N9174);
buf BUF1 (N9313, N9301);
not NOT1 (N9314, N9282);
buf BUF1 (N9315, N9314);
and AND4 (N9316, N9302, N505, N6582, N5453);
nor NOR3 (N9317, N9313, N4152, N2839);
not NOT1 (N9318, N9292);
buf BUF1 (N9319, N9315);
or OR2 (N9320, N9309, N2415);
xor XOR2 (N9321, N9311, N1360);
nor NOR2 (N9322, N9320, N7010);
not NOT1 (N9323, N9316);
or OR4 (N9324, N9318, N3348, N9121, N999);
xor XOR2 (N9325, N9324, N7876);
xor XOR2 (N9326, N9325, N2066);
buf BUF1 (N9327, N9326);
nand NAND4 (N9328, N9327, N1848, N6531, N7856);
xor XOR2 (N9329, N9312, N6679);
nor NOR4 (N9330, N9328, N7809, N986, N7671);
not NOT1 (N9331, N9323);
not NOT1 (N9332, N9310);
and AND2 (N9333, N9331, N7171);
xor XOR2 (N9334, N9319, N3013);
xor XOR2 (N9335, N9330, N1129);
xor XOR2 (N9336, N9304, N2338);
nand NAND3 (N9337, N9333, N6106, N1963);
buf BUF1 (N9338, N9337);
or OR4 (N9339, N9329, N7783, N4933, N4567);
nand NAND3 (N9340, N9332, N5412, N2942);
nand NAND2 (N9341, N9338, N6510);
and AND2 (N9342, N9334, N5596);
not NOT1 (N9343, N9335);
not NOT1 (N9344, N9340);
nand NAND2 (N9345, N9344, N5576);
not NOT1 (N9346, N9317);
buf BUF1 (N9347, N9322);
nand NAND2 (N9348, N9321, N4842);
or OR2 (N9349, N9341, N7425);
nor NOR3 (N9350, N9349, N1525, N7739);
not NOT1 (N9351, N9345);
and AND2 (N9352, N9307, N8643);
xor XOR2 (N9353, N9352, N4767);
nor NOR2 (N9354, N9351, N3330);
nor NOR2 (N9355, N9347, N8940);
and AND2 (N9356, N9350, N1834);
not NOT1 (N9357, N9353);
nor NOR4 (N9358, N9336, N684, N5554, N8055);
not NOT1 (N9359, N9354);
nand NAND4 (N9360, N9359, N7788, N6421, N2595);
nand NAND4 (N9361, N9339, N5676, N2804, N5334);
xor XOR2 (N9362, N9346, N439);
and AND2 (N9363, N9358, N4011);
or OR2 (N9364, N9357, N4966);
xor XOR2 (N9365, N9363, N9084);
nand NAND4 (N9366, N9348, N8635, N7660, N5936);
nor NOR3 (N9367, N9355, N27, N5278);
not NOT1 (N9368, N9361);
nand NAND4 (N9369, N9367, N3573, N844, N3721);
and AND3 (N9370, N9369, N5458, N4061);
nand NAND4 (N9371, N9368, N8256, N8630, N2425);
xor XOR2 (N9372, N9342, N3352);
buf BUF1 (N9373, N9364);
xor XOR2 (N9374, N9370, N7232);
xor XOR2 (N9375, N9365, N334);
buf BUF1 (N9376, N9366);
buf BUF1 (N9377, N9343);
and AND3 (N9378, N9356, N66, N2568);
or OR2 (N9379, N9371, N2186);
xor XOR2 (N9380, N9376, N8468);
and AND2 (N9381, N9379, N8629);
not NOT1 (N9382, N9372);
xor XOR2 (N9383, N9377, N5942);
not NOT1 (N9384, N9381);
nand NAND2 (N9385, N9383, N351);
not NOT1 (N9386, N9374);
and AND3 (N9387, N9360, N2970, N4108);
or OR4 (N9388, N9384, N3382, N3365, N2922);
buf BUF1 (N9389, N9387);
and AND4 (N9390, N9373, N5316, N3503, N2747);
xor XOR2 (N9391, N9385, N8103);
nand NAND4 (N9392, N9380, N1035, N5891, N7624);
nor NOR4 (N9393, N9392, N6783, N7946, N8063);
not NOT1 (N9394, N9388);
nor NOR3 (N9395, N9389, N5948, N8876);
nor NOR2 (N9396, N9362, N846);
buf BUF1 (N9397, N9393);
and AND4 (N9398, N9386, N1003, N1790, N7969);
and AND4 (N9399, N9390, N5259, N8680, N6683);
or OR3 (N9400, N9399, N7971, N2216);
nor NOR4 (N9401, N9375, N8376, N4046, N6080);
nand NAND4 (N9402, N9391, N7701, N2468, N3784);
buf BUF1 (N9403, N9378);
nand NAND2 (N9404, N9382, N52);
nand NAND2 (N9405, N9400, N1128);
nand NAND4 (N9406, N9398, N132, N3786, N6669);
nor NOR3 (N9407, N9394, N2658, N3873);
buf BUF1 (N9408, N9396);
nand NAND3 (N9409, N9408, N8390, N8053);
buf BUF1 (N9410, N9395);
nor NOR4 (N9411, N9401, N4878, N1566, N3767);
buf BUF1 (N9412, N9410);
and AND4 (N9413, N9403, N8728, N6472, N7299);
buf BUF1 (N9414, N9411);
not NOT1 (N9415, N9402);
xor XOR2 (N9416, N9397, N3415);
not NOT1 (N9417, N9405);
or OR4 (N9418, N9416, N3032, N2282, N700);
nor NOR2 (N9419, N9415, N1071);
nand NAND3 (N9420, N9414, N6914, N917);
and AND4 (N9421, N9418, N7119, N8356, N5462);
nor NOR4 (N9422, N9417, N6608, N4505, N2267);
buf BUF1 (N9423, N9419);
nor NOR2 (N9424, N9413, N2065);
or OR4 (N9425, N9404, N6347, N8574, N1249);
buf BUF1 (N9426, N9423);
not NOT1 (N9427, N9426);
or OR2 (N9428, N9421, N4997);
xor XOR2 (N9429, N9412, N8716);
buf BUF1 (N9430, N9409);
nand NAND2 (N9431, N9430, N5595);
nor NOR4 (N9432, N9424, N1156, N791, N7159);
and AND4 (N9433, N9432, N8590, N7851, N2992);
xor XOR2 (N9434, N9428, N2472);
nand NAND3 (N9435, N9434, N3732, N4794);
not NOT1 (N9436, N9429);
not NOT1 (N9437, N9433);
nand NAND2 (N9438, N9420, N8675);
xor XOR2 (N9439, N9438, N6342);
xor XOR2 (N9440, N9407, N3761);
nor NOR2 (N9441, N9435, N1412);
nor NOR2 (N9442, N9439, N9258);
nand NAND3 (N9443, N9406, N575, N3216);
xor XOR2 (N9444, N9431, N4075);
and AND2 (N9445, N9443, N2805);
not NOT1 (N9446, N9442);
nand NAND2 (N9447, N9422, N4899);
buf BUF1 (N9448, N9436);
nor NOR3 (N9449, N9446, N6624, N1705);
buf BUF1 (N9450, N9425);
buf BUF1 (N9451, N9427);
nand NAND3 (N9452, N9449, N1542, N162);
nand NAND3 (N9453, N9450, N8335, N2247);
buf BUF1 (N9454, N9441);
not NOT1 (N9455, N9448);
buf BUF1 (N9456, N9437);
nor NOR4 (N9457, N9455, N1528, N8975, N6580);
or OR2 (N9458, N9445, N5365);
buf BUF1 (N9459, N9457);
or OR3 (N9460, N9447, N8868, N1637);
buf BUF1 (N9461, N9456);
or OR3 (N9462, N9461, N6090, N1496);
or OR3 (N9463, N9458, N3388, N579);
or OR2 (N9464, N9460, N4905);
and AND3 (N9465, N9452, N3581, N204);
not NOT1 (N9466, N9440);
buf BUF1 (N9467, N9465);
nand NAND4 (N9468, N9454, N807, N938, N8347);
buf BUF1 (N9469, N9464);
not NOT1 (N9470, N9444);
nand NAND2 (N9471, N9467, N6686);
buf BUF1 (N9472, N9468);
or OR3 (N9473, N9462, N1338, N1602);
or OR2 (N9474, N9453, N4996);
not NOT1 (N9475, N9463);
not NOT1 (N9476, N9471);
or OR3 (N9477, N9476, N2476, N4183);
nor NOR3 (N9478, N9474, N217, N7374);
and AND2 (N9479, N9472, N2404);
and AND4 (N9480, N9475, N3365, N3382, N8094);
or OR3 (N9481, N9480, N6188, N8150);
buf BUF1 (N9482, N9473);
nand NAND2 (N9483, N9478, N27);
not NOT1 (N9484, N9469);
not NOT1 (N9485, N9484);
nand NAND4 (N9486, N9482, N6385, N1292, N5719);
nand NAND2 (N9487, N9459, N3156);
xor XOR2 (N9488, N9451, N3291);
not NOT1 (N9489, N9477);
buf BUF1 (N9490, N9483);
xor XOR2 (N9491, N9490, N3610);
and AND3 (N9492, N9488, N2561, N6808);
or OR4 (N9493, N9489, N3560, N8435, N4919);
xor XOR2 (N9494, N9493, N4343);
buf BUF1 (N9495, N9466);
and AND3 (N9496, N9487, N4668, N7141);
xor XOR2 (N9497, N9485, N8419);
or OR4 (N9498, N9494, N3443, N6929, N314);
not NOT1 (N9499, N9470);
xor XOR2 (N9500, N9486, N9208);
buf BUF1 (N9501, N9479);
buf BUF1 (N9502, N9491);
nor NOR2 (N9503, N9501, N1810);
nor NOR3 (N9504, N9502, N5348, N4479);
nor NOR4 (N9505, N9481, N7098, N8017, N4048);
or OR4 (N9506, N9495, N8573, N401, N4018);
nand NAND2 (N9507, N9496, N5472);
nor NOR2 (N9508, N9500, N5392);
nand NAND2 (N9509, N9506, N4050);
buf BUF1 (N9510, N9503);
nand NAND3 (N9511, N9507, N1202, N5500);
nor NOR4 (N9512, N9511, N4145, N9118, N1421);
or OR4 (N9513, N9505, N1587, N1523, N6731);
xor XOR2 (N9514, N9510, N5576);
nor NOR3 (N9515, N9504, N8965, N4325);
xor XOR2 (N9516, N9514, N2302);
nand NAND4 (N9517, N9516, N8631, N8145, N1389);
or OR4 (N9518, N9513, N2696, N6865, N5711);
not NOT1 (N9519, N9509);
nand NAND4 (N9520, N9492, N8326, N9112, N1228);
and AND2 (N9521, N9512, N5446);
buf BUF1 (N9522, N9498);
buf BUF1 (N9523, N9522);
nor NOR4 (N9524, N9497, N6501, N4632, N7507);
xor XOR2 (N9525, N9517, N7560);
nand NAND2 (N9526, N9519, N4205);
not NOT1 (N9527, N9526);
or OR4 (N9528, N9521, N3373, N3777, N9263);
xor XOR2 (N9529, N9518, N6713);
or OR2 (N9530, N9524, N3541);
not NOT1 (N9531, N9528);
nor NOR4 (N9532, N9520, N2632, N444, N4518);
nand NAND3 (N9533, N9532, N5595, N7032);
xor XOR2 (N9534, N9530, N9253);
buf BUF1 (N9535, N9499);
and AND4 (N9536, N9533, N7367, N7139, N2045);
not NOT1 (N9537, N9536);
nor NOR3 (N9538, N9508, N243, N5722);
nand NAND3 (N9539, N9538, N5276, N9507);
or OR3 (N9540, N9539, N6025, N61);
and AND3 (N9541, N9537, N2008, N322);
xor XOR2 (N9542, N9523, N6597);
nand NAND2 (N9543, N9525, N7366);
nor NOR2 (N9544, N9531, N4545);
nor NOR3 (N9545, N9541, N6912, N7055);
xor XOR2 (N9546, N9544, N3826);
xor XOR2 (N9547, N9542, N8100);
buf BUF1 (N9548, N9515);
and AND3 (N9549, N9540, N8888, N2718);
or OR4 (N9550, N9549, N6219, N4649, N9120);
and AND3 (N9551, N9527, N7245, N8602);
or OR4 (N9552, N9543, N3248, N436, N3142);
or OR2 (N9553, N9548, N1840);
and AND3 (N9554, N9545, N2534, N7871);
xor XOR2 (N9555, N9554, N7730);
not NOT1 (N9556, N9534);
nand NAND3 (N9557, N9529, N5905, N6976);
or OR2 (N9558, N9551, N1533);
and AND2 (N9559, N9557, N8942);
buf BUF1 (N9560, N9552);
xor XOR2 (N9561, N9560, N8523);
or OR2 (N9562, N9559, N7880);
and AND2 (N9563, N9553, N6669);
or OR2 (N9564, N9550, N3204);
and AND4 (N9565, N9555, N5877, N114, N6561);
nand NAND2 (N9566, N9563, N5320);
nand NAND4 (N9567, N9561, N346, N4957, N1463);
nand NAND4 (N9568, N9558, N8245, N9390, N5450);
or OR3 (N9569, N9568, N1496, N9133);
xor XOR2 (N9570, N9567, N6068);
or OR3 (N9571, N9569, N8347, N2465);
nand NAND3 (N9572, N9562, N1944, N1492);
xor XOR2 (N9573, N9571, N7878);
and AND3 (N9574, N9573, N4581, N1947);
not NOT1 (N9575, N9566);
nor NOR4 (N9576, N9565, N12, N233, N6902);
nor NOR4 (N9577, N9547, N3036, N6960, N8163);
and AND2 (N9578, N9572, N9432);
not NOT1 (N9579, N9577);
xor XOR2 (N9580, N9535, N3845);
xor XOR2 (N9581, N9576, N9422);
nor NOR3 (N9582, N9578, N3523, N966);
nand NAND2 (N9583, N9570, N2767);
or OR4 (N9584, N9574, N2221, N914, N5159);
or OR4 (N9585, N9584, N6505, N4610, N4058);
nor NOR2 (N9586, N9579, N266);
or OR3 (N9587, N9586, N554, N1974);
nor NOR4 (N9588, N9575, N612, N9572, N177);
buf BUF1 (N9589, N9582);
or OR2 (N9590, N9564, N1201);
or OR2 (N9591, N9583, N3311);
buf BUF1 (N9592, N9585);
xor XOR2 (N9593, N9591, N2770);
nand NAND3 (N9594, N9592, N132, N2597);
or OR3 (N9595, N9588, N2644, N1987);
nor NOR3 (N9596, N9556, N715, N6587);
or OR3 (N9597, N9580, N4451, N3414);
buf BUF1 (N9598, N9589);
not NOT1 (N9599, N9594);
nor NOR3 (N9600, N9546, N4783, N8806);
nand NAND4 (N9601, N9581, N3448, N3812, N6613);
and AND4 (N9602, N9587, N4699, N6417, N936);
not NOT1 (N9603, N9600);
xor XOR2 (N9604, N9599, N7365);
buf BUF1 (N9605, N9602);
buf BUF1 (N9606, N9601);
nor NOR4 (N9607, N9595, N111, N9430, N4045);
and AND4 (N9608, N9597, N3851, N8552, N5073);
and AND4 (N9609, N9604, N2733, N7131, N8347);
xor XOR2 (N9610, N9606, N5922);
nand NAND2 (N9611, N9596, N5895);
not NOT1 (N9612, N9603);
nor NOR3 (N9613, N9612, N2462, N62);
nor NOR2 (N9614, N9609, N4442);
nand NAND3 (N9615, N9605, N1383, N1438);
buf BUF1 (N9616, N9611);
nor NOR3 (N9617, N9614, N5849, N9073);
nand NAND3 (N9618, N9607, N6707, N6959);
nor NOR2 (N9619, N9590, N617);
nor NOR4 (N9620, N9619, N8283, N2933, N935);
or OR2 (N9621, N9610, N1249);
or OR3 (N9622, N9615, N7765, N6642);
nor NOR4 (N9623, N9622, N5614, N6090, N1160);
buf BUF1 (N9624, N9618);
nor NOR4 (N9625, N9624, N1386, N3223, N3705);
or OR3 (N9626, N9623, N3075, N1171);
and AND2 (N9627, N9620, N5505);
nor NOR4 (N9628, N9616, N7941, N5139, N4204);
buf BUF1 (N9629, N9625);
buf BUF1 (N9630, N9617);
buf BUF1 (N9631, N9629);
and AND3 (N9632, N9593, N8939, N4275);
or OR3 (N9633, N9613, N361, N3238);
not NOT1 (N9634, N9631);
and AND3 (N9635, N9621, N2027, N1037);
or OR3 (N9636, N9626, N4400, N8223);
nand NAND2 (N9637, N9598, N1187);
nor NOR4 (N9638, N9633, N3665, N7498, N9523);
or OR3 (N9639, N9630, N4464, N8663);
nand NAND4 (N9640, N9635, N2097, N4587, N2449);
buf BUF1 (N9641, N9608);
not NOT1 (N9642, N9636);
xor XOR2 (N9643, N9627, N4520);
nor NOR2 (N9644, N9640, N672);
buf BUF1 (N9645, N9639);
buf BUF1 (N9646, N9628);
nand NAND3 (N9647, N9638, N7549, N3736);
nand NAND3 (N9648, N9646, N7176, N8402);
or OR2 (N9649, N9648, N8234);
not NOT1 (N9650, N9641);
nor NOR4 (N9651, N9644, N8423, N6942, N8233);
xor XOR2 (N9652, N9634, N8871);
nand NAND3 (N9653, N9643, N7937, N8340);
nor NOR3 (N9654, N9649, N6316, N2821);
and AND4 (N9655, N9651, N2648, N937, N4498);
or OR3 (N9656, N9642, N7159, N7799);
nand NAND3 (N9657, N9653, N7815, N1174);
not NOT1 (N9658, N9657);
or OR2 (N9659, N9658, N1087);
xor XOR2 (N9660, N9659, N7740);
nor NOR3 (N9661, N9654, N5649, N113);
nand NAND3 (N9662, N9647, N4114, N5169);
nand NAND2 (N9663, N9650, N4937);
nor NOR4 (N9664, N9655, N6810, N8363, N6190);
nand NAND3 (N9665, N9652, N6363, N6615);
and AND3 (N9666, N9661, N9174, N8854);
not NOT1 (N9667, N9662);
not NOT1 (N9668, N9656);
buf BUF1 (N9669, N9663);
not NOT1 (N9670, N9668);
and AND2 (N9671, N9670, N1695);
nor NOR2 (N9672, N9665, N9057);
xor XOR2 (N9673, N9645, N6239);
nand NAND2 (N9674, N9660, N3635);
nor NOR3 (N9675, N9666, N1564, N9435);
buf BUF1 (N9676, N9667);
and AND2 (N9677, N9672, N5918);
nor NOR4 (N9678, N9632, N527, N8587, N8919);
or OR4 (N9679, N9671, N5953, N4640, N4845);
or OR4 (N9680, N9669, N2065, N6176, N5164);
nand NAND4 (N9681, N9675, N693, N5778, N4618);
not NOT1 (N9682, N9673);
nand NAND4 (N9683, N9680, N1585, N1681, N9193);
nor NOR4 (N9684, N9682, N2913, N1291, N1652);
nor NOR3 (N9685, N9681, N8810, N8123);
buf BUF1 (N9686, N9664);
buf BUF1 (N9687, N9678);
nor NOR3 (N9688, N9676, N5018, N9470);
or OR4 (N9689, N9686, N5771, N1279, N3196);
xor XOR2 (N9690, N9689, N5199);
buf BUF1 (N9691, N9688);
xor XOR2 (N9692, N9677, N717);
and AND2 (N9693, N9685, N2277);
nand NAND2 (N9694, N9690, N6686);
nand NAND3 (N9695, N9637, N6755, N2267);
not NOT1 (N9696, N9695);
or OR2 (N9697, N9694, N2991);
not NOT1 (N9698, N9696);
buf BUF1 (N9699, N9684);
xor XOR2 (N9700, N9699, N8930);
or OR4 (N9701, N9692, N2884, N9007, N6512);
or OR2 (N9702, N9697, N3609);
nand NAND2 (N9703, N9700, N3239);
xor XOR2 (N9704, N9691, N2733);
nand NAND4 (N9705, N9704, N5109, N632, N4050);
nor NOR4 (N9706, N9698, N5733, N9498, N1003);
buf BUF1 (N9707, N9687);
xor XOR2 (N9708, N9701, N4373);
nand NAND3 (N9709, N9708, N4947, N6789);
nand NAND2 (N9710, N9707, N736);
and AND2 (N9711, N9709, N1430);
and AND4 (N9712, N9711, N2839, N1357, N8510);
xor XOR2 (N9713, N9710, N1957);
nor NOR4 (N9714, N9674, N8855, N6004, N8529);
and AND4 (N9715, N9679, N5243, N790, N5842);
and AND3 (N9716, N9715, N5824, N1387);
not NOT1 (N9717, N9705);
nor NOR2 (N9718, N9717, N9486);
and AND4 (N9719, N9714, N8738, N4873, N1249);
and AND4 (N9720, N9713, N6761, N8198, N9056);
nand NAND2 (N9721, N9702, N9288);
nand NAND4 (N9722, N9712, N1655, N3178, N4099);
nand NAND3 (N9723, N9706, N6960, N1266);
xor XOR2 (N9724, N9683, N8248);
and AND2 (N9725, N9716, N4564);
not NOT1 (N9726, N9720);
xor XOR2 (N9727, N9724, N9225);
and AND2 (N9728, N9725, N3842);
not NOT1 (N9729, N9721);
and AND3 (N9730, N9727, N3976, N329);
xor XOR2 (N9731, N9693, N4172);
buf BUF1 (N9732, N9731);
nand NAND4 (N9733, N9726, N343, N3987, N6830);
not NOT1 (N9734, N9723);
not NOT1 (N9735, N9729);
or OR4 (N9736, N9732, N8685, N9330, N7191);
buf BUF1 (N9737, N9733);
nand NAND4 (N9738, N9719, N9622, N8803, N3438);
nor NOR2 (N9739, N9730, N2355);
buf BUF1 (N9740, N9737);
nor NOR2 (N9741, N9734, N6329);
not NOT1 (N9742, N9728);
and AND2 (N9743, N9739, N6496);
buf BUF1 (N9744, N9736);
or OR2 (N9745, N9703, N8849);
xor XOR2 (N9746, N9722, N2055);
nor NOR3 (N9747, N9746, N9632, N3116);
xor XOR2 (N9748, N9742, N7114);
nand NAND2 (N9749, N9748, N4198);
nand NAND3 (N9750, N9738, N5559, N4476);
nor NOR2 (N9751, N9718, N7118);
nor NOR2 (N9752, N9743, N8694);
and AND4 (N9753, N9749, N9290, N9314, N3690);
or OR3 (N9754, N9735, N5659, N3807);
xor XOR2 (N9755, N9750, N657);
and AND3 (N9756, N9744, N9399, N219);
buf BUF1 (N9757, N9752);
xor XOR2 (N9758, N9745, N3070);
and AND2 (N9759, N9751, N8887);
buf BUF1 (N9760, N9755);
and AND2 (N9761, N9753, N2428);
nor NOR3 (N9762, N9759, N8878, N9420);
and AND3 (N9763, N9740, N6069, N6656);
not NOT1 (N9764, N9760);
and AND3 (N9765, N9762, N1655, N3593);
xor XOR2 (N9766, N9765, N8486);
nor NOR2 (N9767, N9766, N3493);
nand NAND3 (N9768, N9757, N4721, N3069);
nor NOR4 (N9769, N9754, N6195, N3593, N6214);
xor XOR2 (N9770, N9768, N6496);
buf BUF1 (N9771, N9741);
nor NOR4 (N9772, N9769, N1035, N8245, N580);
or OR2 (N9773, N9756, N6852);
or OR2 (N9774, N9758, N5174);
or OR2 (N9775, N9773, N3813);
not NOT1 (N9776, N9763);
nor NOR2 (N9777, N9775, N9751);
and AND2 (N9778, N9747, N1202);
xor XOR2 (N9779, N9774, N83);
nor NOR4 (N9780, N9778, N646, N904, N1284);
not NOT1 (N9781, N9770);
xor XOR2 (N9782, N9776, N8125);
xor XOR2 (N9783, N9777, N542);
or OR3 (N9784, N9780, N3425, N2009);
and AND4 (N9785, N9784, N6587, N6960, N5075);
or OR4 (N9786, N9771, N6699, N7840, N5845);
nand NAND4 (N9787, N9783, N5351, N8801, N4096);
xor XOR2 (N9788, N9764, N9546);
nand NAND4 (N9789, N9785, N2647, N8254, N195);
and AND2 (N9790, N9761, N6230);
buf BUF1 (N9791, N9788);
nor NOR4 (N9792, N9787, N4227, N802, N3702);
xor XOR2 (N9793, N9779, N7337);
xor XOR2 (N9794, N9792, N4914);
xor XOR2 (N9795, N9790, N3477);
nand NAND4 (N9796, N9781, N7468, N9235, N9081);
nor NOR2 (N9797, N9786, N879);
nand NAND3 (N9798, N9789, N7869, N2953);
and AND4 (N9799, N9796, N1458, N273, N6239);
nand NAND2 (N9800, N9795, N4423);
not NOT1 (N9801, N9782);
nor NOR2 (N9802, N9793, N9270);
buf BUF1 (N9803, N9799);
or OR4 (N9804, N9794, N1638, N3733, N4185);
nor NOR3 (N9805, N9798, N3460, N7083);
and AND2 (N9806, N9802, N834);
not NOT1 (N9807, N9767);
nor NOR3 (N9808, N9807, N7377, N5697);
and AND2 (N9809, N9791, N7719);
buf BUF1 (N9810, N9801);
nor NOR2 (N9811, N9808, N5417);
nor NOR2 (N9812, N9803, N2983);
or OR2 (N9813, N9797, N7694);
nand NAND4 (N9814, N9772, N6039, N8280, N3434);
not NOT1 (N9815, N9804);
nor NOR4 (N9816, N9806, N4493, N5158, N3626);
not NOT1 (N9817, N9811);
nand NAND2 (N9818, N9800, N7548);
and AND3 (N9819, N9814, N7749, N5503);
not NOT1 (N9820, N9818);
xor XOR2 (N9821, N9805, N7611);
or OR2 (N9822, N9815, N3896);
not NOT1 (N9823, N9821);
and AND3 (N9824, N9816, N3441, N1017);
not NOT1 (N9825, N9822);
and AND3 (N9826, N9819, N2553, N4341);
xor XOR2 (N9827, N9817, N5890);
and AND2 (N9828, N9809, N2027);
xor XOR2 (N9829, N9827, N7354);
or OR2 (N9830, N9825, N2348);
nand NAND4 (N9831, N9830, N7139, N2301, N5840);
not NOT1 (N9832, N9820);
nor NOR2 (N9833, N9824, N4692);
nor NOR3 (N9834, N9810, N7449, N2596);
buf BUF1 (N9835, N9833);
buf BUF1 (N9836, N9823);
or OR4 (N9837, N9828, N6925, N1965, N3821);
not NOT1 (N9838, N9832);
xor XOR2 (N9839, N9836, N3395);
buf BUF1 (N9840, N9831);
nor NOR4 (N9841, N9834, N6010, N2006, N563);
xor XOR2 (N9842, N9837, N3411);
or OR3 (N9843, N9812, N925, N9368);
or OR4 (N9844, N9839, N9781, N6259, N9450);
xor XOR2 (N9845, N9841, N5018);
nor NOR2 (N9846, N9840, N7673);
and AND2 (N9847, N9826, N721);
not NOT1 (N9848, N9843);
nor NOR3 (N9849, N9844, N5300, N9800);
or OR4 (N9850, N9813, N6206, N4507, N9123);
nand NAND2 (N9851, N9835, N2336);
buf BUF1 (N9852, N9848);
xor XOR2 (N9853, N9849, N2797);
or OR3 (N9854, N9842, N457, N2910);
and AND3 (N9855, N9847, N8709, N112);
and AND3 (N9856, N9850, N7145, N5461);
and AND4 (N9857, N9852, N3704, N7125, N6706);
nand NAND4 (N9858, N9854, N5679, N8663, N9443);
buf BUF1 (N9859, N9829);
nand NAND3 (N9860, N9838, N2036, N4303);
not NOT1 (N9861, N9846);
nand NAND2 (N9862, N9859, N1824);
nor NOR3 (N9863, N9855, N3749, N7299);
xor XOR2 (N9864, N9845, N4704);
xor XOR2 (N9865, N9863, N7665);
buf BUF1 (N9866, N9853);
or OR2 (N9867, N9866, N3103);
nand NAND2 (N9868, N9860, N4078);
buf BUF1 (N9869, N9856);
buf BUF1 (N9870, N9858);
nor NOR3 (N9871, N9870, N2795, N5800);
buf BUF1 (N9872, N9864);
or OR2 (N9873, N9865, N3453);
nor NOR4 (N9874, N9872, N332, N4647, N1099);
nor NOR2 (N9875, N9868, N2203);
nor NOR3 (N9876, N9857, N3055, N3828);
not NOT1 (N9877, N9861);
xor XOR2 (N9878, N9851, N7716);
nor NOR2 (N9879, N9875, N9286);
nand NAND3 (N9880, N9862, N5871, N4811);
and AND2 (N9881, N9878, N6105);
not NOT1 (N9882, N9873);
or OR4 (N9883, N9874, N9480, N8060, N1298);
buf BUF1 (N9884, N9871);
not NOT1 (N9885, N9883);
nand NAND4 (N9886, N9882, N3938, N6468, N3398);
or OR4 (N9887, N9884, N4315, N4073, N3374);
or OR2 (N9888, N9867, N3969);
buf BUF1 (N9889, N9886);
and AND3 (N9890, N9885, N5733, N1925);
xor XOR2 (N9891, N9877, N3496);
xor XOR2 (N9892, N9891, N5090);
xor XOR2 (N9893, N9869, N921);
not NOT1 (N9894, N9879);
not NOT1 (N9895, N9890);
nor NOR2 (N9896, N9880, N7041);
or OR3 (N9897, N9888, N5169, N4566);
buf BUF1 (N9898, N9896);
and AND2 (N9899, N9881, N6519);
nor NOR3 (N9900, N9898, N6241, N2854);
nor NOR2 (N9901, N9895, N4449);
nor NOR3 (N9902, N9876, N1235, N7256);
nand NAND2 (N9903, N9889, N2006);
and AND3 (N9904, N9902, N7652, N9033);
nor NOR3 (N9905, N9894, N170, N8961);
and AND3 (N9906, N9905, N4903, N5524);
xor XOR2 (N9907, N9904, N3401);
nor NOR3 (N9908, N9897, N3445, N5605);
or OR2 (N9909, N9907, N4299);
or OR3 (N9910, N9892, N8160, N2710);
nand NAND3 (N9911, N9887, N1107, N4004);
nand NAND3 (N9912, N9908, N5464, N2947);
and AND3 (N9913, N9910, N8322, N3783);
nand NAND2 (N9914, N9906, N4872);
and AND2 (N9915, N9912, N4926);
and AND4 (N9916, N9900, N5355, N3122, N1903);
buf BUF1 (N9917, N9899);
or OR3 (N9918, N9917, N9244, N283);
buf BUF1 (N9919, N9901);
not NOT1 (N9920, N9913);
nor NOR2 (N9921, N9914, N678);
not NOT1 (N9922, N9893);
xor XOR2 (N9923, N9921, N3576);
and AND4 (N9924, N9920, N3940, N593, N301);
buf BUF1 (N9925, N9915);
not NOT1 (N9926, N9918);
nand NAND2 (N9927, N9903, N5512);
nor NOR2 (N9928, N9926, N874);
not NOT1 (N9929, N9923);
buf BUF1 (N9930, N9909);
and AND3 (N9931, N9930, N9295, N192);
nand NAND4 (N9932, N9927, N8808, N8763, N9422);
or OR4 (N9933, N9931, N4118, N2033, N177);
nand NAND3 (N9934, N9932, N8055, N1065);
nand NAND2 (N9935, N9933, N2011);
nor NOR2 (N9936, N9916, N6334);
buf BUF1 (N9937, N9922);
xor XOR2 (N9938, N9919, N8017);
nor NOR3 (N9939, N9911, N4490, N1426);
and AND3 (N9940, N9935, N4122, N1107);
or OR3 (N9941, N9937, N4859, N5067);
nor NOR4 (N9942, N9939, N254, N4358, N1648);
nor NOR3 (N9943, N9941, N1992, N4317);
buf BUF1 (N9944, N9934);
nand NAND4 (N9945, N9943, N7308, N1901, N1527);
or OR4 (N9946, N9925, N6033, N6561, N2837);
or OR2 (N9947, N9946, N1659);
xor XOR2 (N9948, N9944, N3562);
not NOT1 (N9949, N9928);
not NOT1 (N9950, N9940);
nor NOR4 (N9951, N9949, N5189, N3007, N1007);
nand NAND2 (N9952, N9929, N1430);
or OR2 (N9953, N9950, N7855);
buf BUF1 (N9954, N9938);
buf BUF1 (N9955, N9952);
xor XOR2 (N9956, N9955, N9606);
nand NAND3 (N9957, N9951, N8426, N7127);
and AND4 (N9958, N9942, N9114, N6995, N2779);
buf BUF1 (N9959, N9948);
or OR3 (N9960, N9953, N9149, N8470);
nand NAND2 (N9961, N9924, N8322);
nor NOR2 (N9962, N9961, N2474);
xor XOR2 (N9963, N9960, N9786);
not NOT1 (N9964, N9957);
buf BUF1 (N9965, N9958);
or OR2 (N9966, N9962, N8400);
buf BUF1 (N9967, N9965);
not NOT1 (N9968, N9964);
buf BUF1 (N9969, N9967);
not NOT1 (N9970, N9966);
nor NOR4 (N9971, N9947, N7524, N5157, N6167);
nand NAND4 (N9972, N9956, N7212, N2900, N6656);
nand NAND3 (N9973, N9954, N4259, N2437);
nand NAND3 (N9974, N9969, N7111, N3899);
nor NOR4 (N9975, N9959, N3724, N9950, N5811);
nor NOR3 (N9976, N9963, N5742, N8221);
buf BUF1 (N9977, N9976);
nor NOR2 (N9978, N9973, N4435);
not NOT1 (N9979, N9977);
nand NAND4 (N9980, N9974, N7049, N7228, N5019);
or OR3 (N9981, N9970, N4539, N1280);
nand NAND4 (N9982, N9945, N8191, N3530, N7812);
xor XOR2 (N9983, N9978, N5852);
and AND2 (N9984, N9980, N669);
buf BUF1 (N9985, N9968);
xor XOR2 (N9986, N9979, N428);
xor XOR2 (N9987, N9986, N1774);
and AND3 (N9988, N9936, N2407, N6666);
nand NAND2 (N9989, N9983, N8282);
buf BUF1 (N9990, N9981);
nor NOR4 (N9991, N9975, N5892, N7637, N634);
buf BUF1 (N9992, N9987);
not NOT1 (N9993, N9992);
nand NAND2 (N9994, N9982, N7057);
and AND2 (N9995, N9972, N2717);
buf BUF1 (N9996, N9995);
buf BUF1 (N9997, N9989);
buf BUF1 (N9998, N9997);
or OR3 (N9999, N9984, N2091, N7184);
xor XOR2 (N10000, N9998, N5859);
and AND3 (N10001, N10000, N5520, N9823);
nand NAND4 (N10002, N9971, N6594, N3136, N3329);
nor NOR2 (N10003, N9999, N403);
and AND4 (N10004, N9996, N3323, N8222, N4793);
nor NOR2 (N10005, N9994, N3486);
and AND3 (N10006, N9985, N6481, N5576);
nand NAND4 (N10007, N10003, N5897, N7520, N4851);
and AND4 (N10008, N9988, N5726, N5346, N3969);
xor XOR2 (N10009, N9990, N3407);
buf BUF1 (N10010, N10009);
not NOT1 (N10011, N10005);
buf BUF1 (N10012, N10004);
buf BUF1 (N10013, N9993);
nand NAND3 (N10014, N10011, N1529, N1617);
nand NAND4 (N10015, N10010, N3317, N4824, N7179);
buf BUF1 (N10016, N10015);
not NOT1 (N10017, N10014);
nand NAND2 (N10018, N9991, N7062);
and AND3 (N10019, N10018, N7443, N8587);
xor XOR2 (N10020, N10006, N2582);
and AND4 (N10021, N10008, N5169, N162, N6821);
nor NOR4 (N10022, N10017, N1391, N9296, N7760);
buf BUF1 (N10023, N10022);
xor XOR2 (N10024, N10007, N8777);
buf BUF1 (N10025, N10012);
nand NAND4 (N10026, N10025, N9973, N3421, N5943);
xor XOR2 (N10027, N10021, N2049);
nand NAND2 (N10028, N10013, N7682);
not NOT1 (N10029, N10019);
buf BUF1 (N10030, N10027);
xor XOR2 (N10031, N10028, N9703);
nor NOR2 (N10032, N10016, N7811);
nand NAND3 (N10033, N10031, N1269, N1092);
not NOT1 (N10034, N10026);
xor XOR2 (N10035, N10029, N11);
xor XOR2 (N10036, N10001, N3426);
nand NAND3 (N10037, N10024, N6876, N1229);
and AND3 (N10038, N10030, N3807, N9462);
or OR4 (N10039, N10034, N2847, N6803, N2596);
and AND4 (N10040, N10002, N9208, N8718, N9668);
or OR2 (N10041, N10023, N528);
not NOT1 (N10042, N10035);
nand NAND3 (N10043, N10036, N8438, N4469);
not NOT1 (N10044, N10038);
or OR2 (N10045, N10032, N1899);
not NOT1 (N10046, N10043);
and AND4 (N10047, N10033, N6634, N2692, N4653);
buf BUF1 (N10048, N10044);
and AND4 (N10049, N10020, N8465, N9765, N5593);
xor XOR2 (N10050, N10049, N1491);
and AND2 (N10051, N10047, N4364);
xor XOR2 (N10052, N10050, N4559);
not NOT1 (N10053, N10041);
nand NAND2 (N10054, N10053, N852);
buf BUF1 (N10055, N10037);
xor XOR2 (N10056, N10054, N9805);
and AND3 (N10057, N10048, N5626, N9002);
xor XOR2 (N10058, N10039, N6913);
and AND3 (N10059, N10040, N6617, N4005);
buf BUF1 (N10060, N10045);
and AND2 (N10061, N10046, N5619);
buf BUF1 (N10062, N10055);
or OR3 (N10063, N10059, N3476, N480);
nor NOR4 (N10064, N10051, N1910, N1732, N647);
or OR3 (N10065, N10057, N6420, N9980);
nand NAND3 (N10066, N10065, N6468, N10045);
not NOT1 (N10067, N10064);
nand NAND2 (N10068, N10052, N4346);
or OR4 (N10069, N10068, N2338, N6471, N990);
buf BUF1 (N10070, N10042);
xor XOR2 (N10071, N10058, N2912);
not NOT1 (N10072, N10066);
nor NOR4 (N10073, N10067, N1417, N6883, N8858);
nand NAND2 (N10074, N10070, N1677);
nand NAND2 (N10075, N10061, N2550);
nor NOR2 (N10076, N10062, N4249);
and AND2 (N10077, N10069, N6542);
or OR2 (N10078, N10056, N1849);
buf BUF1 (N10079, N10078);
xor XOR2 (N10080, N10060, N5916);
nor NOR4 (N10081, N10077, N2133, N4822, N5810);
or OR3 (N10082, N10072, N7128, N4384);
xor XOR2 (N10083, N10080, N612);
and AND3 (N10084, N10081, N3448, N788);
and AND2 (N10085, N10076, N3015);
or OR4 (N10086, N10071, N3531, N2554, N1008);
or OR2 (N10087, N10083, N4889);
or OR4 (N10088, N10085, N8621, N139, N8679);
nand NAND2 (N10089, N10087, N4367);
xor XOR2 (N10090, N10075, N8896);
or OR3 (N10091, N10088, N6049, N9136);
nor NOR2 (N10092, N10090, N1601);
xor XOR2 (N10093, N10063, N5031);
xor XOR2 (N10094, N10092, N865);
or OR3 (N10095, N10074, N3276, N2078);
and AND4 (N10096, N10091, N9915, N7283, N8554);
buf BUF1 (N10097, N10082);
or OR4 (N10098, N10093, N9555, N1933, N9164);
xor XOR2 (N10099, N10096, N6861);
buf BUF1 (N10100, N10089);
buf BUF1 (N10101, N10095);
or OR4 (N10102, N10094, N9817, N8975, N9756);
xor XOR2 (N10103, N10086, N2348);
and AND2 (N10104, N10101, N2510);
and AND2 (N10105, N10100, N1661);
nor NOR4 (N10106, N10073, N5011, N5265, N8125);
xor XOR2 (N10107, N10102, N6886);
xor XOR2 (N10108, N10107, N781);
or OR4 (N10109, N10098, N1333, N820, N383);
buf BUF1 (N10110, N10099);
nand NAND4 (N10111, N10079, N4144, N1002, N5161);
and AND3 (N10112, N10103, N438, N256);
buf BUF1 (N10113, N10112);
xor XOR2 (N10114, N10111, N4348);
nor NOR3 (N10115, N10106, N3818, N4343);
not NOT1 (N10116, N10115);
and AND2 (N10117, N10097, N2979);
or OR2 (N10118, N10109, N2958);
nand NAND2 (N10119, N10105, N2187);
or OR2 (N10120, N10104, N5444);
buf BUF1 (N10121, N10108);
nand NAND4 (N10122, N10121, N1506, N8296, N9682);
and AND3 (N10123, N10118, N4774, N4274);
nor NOR4 (N10124, N10113, N10002, N7783, N5775);
buf BUF1 (N10125, N10119);
nor NOR4 (N10126, N10114, N9654, N8105, N7080);
nor NOR4 (N10127, N10124, N8614, N9845, N8918);
or OR2 (N10128, N10110, N1351);
or OR2 (N10129, N10084, N5831);
or OR2 (N10130, N10116, N2385);
and AND4 (N10131, N10122, N9868, N7722, N5235);
nor NOR3 (N10132, N10130, N9187, N4595);
nand NAND4 (N10133, N10131, N10114, N116, N7828);
not NOT1 (N10134, N10117);
and AND4 (N10135, N10132, N1880, N5192, N969);
or OR3 (N10136, N10126, N176, N4074);
and AND4 (N10137, N10128, N6100, N5453, N9170);
not NOT1 (N10138, N10123);
nand NAND2 (N10139, N10129, N3740);
nor NOR2 (N10140, N10133, N10080);
nand NAND4 (N10141, N10127, N6913, N1727, N1423);
and AND2 (N10142, N10137, N3820);
not NOT1 (N10143, N10134);
nand NAND4 (N10144, N10139, N5844, N6561, N2674);
nor NOR3 (N10145, N10143, N3122, N3935);
xor XOR2 (N10146, N10142, N146);
buf BUF1 (N10147, N10145);
or OR4 (N10148, N10144, N5552, N4726, N6496);
xor XOR2 (N10149, N10140, N1402);
nor NOR2 (N10150, N10148, N8040);
and AND4 (N10151, N10136, N2163, N7480, N3284);
nand NAND4 (N10152, N10150, N2828, N8965, N9196);
or OR2 (N10153, N10149, N3072);
xor XOR2 (N10154, N10138, N6002);
and AND2 (N10155, N10135, N9731);
xor XOR2 (N10156, N10153, N4693);
nand NAND3 (N10157, N10152, N5859, N4492);
xor XOR2 (N10158, N10156, N626);
xor XOR2 (N10159, N10158, N1813);
not NOT1 (N10160, N10151);
buf BUF1 (N10161, N10154);
or OR3 (N10162, N10146, N8070, N4031);
or OR3 (N10163, N10160, N7020, N9260);
nand NAND2 (N10164, N10163, N10140);
buf BUF1 (N10165, N10161);
xor XOR2 (N10166, N10120, N4099);
xor XOR2 (N10167, N10125, N4656);
and AND2 (N10168, N10141, N3907);
not NOT1 (N10169, N10159);
nand NAND2 (N10170, N10164, N634);
buf BUF1 (N10171, N10167);
nor NOR3 (N10172, N10169, N3282, N7473);
xor XOR2 (N10173, N10172, N2441);
nand NAND4 (N10174, N10168, N2889, N767, N1452);
not NOT1 (N10175, N10165);
xor XOR2 (N10176, N10170, N8426);
not NOT1 (N10177, N10166);
and AND3 (N10178, N10157, N3640, N4150);
nor NOR4 (N10179, N10171, N4572, N8701, N989);
xor XOR2 (N10180, N10174, N1048);
and AND3 (N10181, N10155, N9233, N1718);
and AND3 (N10182, N10179, N7674, N733);
xor XOR2 (N10183, N10176, N5249);
not NOT1 (N10184, N10162);
nor NOR4 (N10185, N10173, N5603, N541, N7430);
buf BUF1 (N10186, N10181);
not NOT1 (N10187, N10177);
buf BUF1 (N10188, N10182);
buf BUF1 (N10189, N10147);
nand NAND4 (N10190, N10185, N1448, N1201, N1144);
xor XOR2 (N10191, N10186, N2378);
nand NAND2 (N10192, N10183, N3162);
nor NOR4 (N10193, N10191, N2188, N303, N4151);
xor XOR2 (N10194, N10190, N6315);
and AND3 (N10195, N10184, N7397, N1825);
not NOT1 (N10196, N10193);
not NOT1 (N10197, N10175);
and AND2 (N10198, N10189, N3724);
nand NAND4 (N10199, N10180, N9273, N3114, N8581);
or OR3 (N10200, N10196, N1078, N510);
nand NAND2 (N10201, N10195, N4105);
not NOT1 (N10202, N10194);
nand NAND2 (N10203, N10197, N8173);
or OR2 (N10204, N10202, N7824);
nor NOR3 (N10205, N10198, N3734, N1221);
not NOT1 (N10206, N10204);
nand NAND4 (N10207, N10205, N8554, N2501, N4062);
nand NAND4 (N10208, N10188, N2211, N3651, N6308);
buf BUF1 (N10209, N10208);
not NOT1 (N10210, N10201);
or OR2 (N10211, N10192, N8112);
nand NAND4 (N10212, N10187, N3161, N1232, N8360);
xor XOR2 (N10213, N10209, N8027);
and AND2 (N10214, N10203, N5501);
xor XOR2 (N10215, N10210, N3506);
not NOT1 (N10216, N10178);
or OR2 (N10217, N10213, N5465);
not NOT1 (N10218, N10215);
nand NAND2 (N10219, N10217, N3170);
or OR2 (N10220, N10211, N2113);
or OR2 (N10221, N10218, N2407);
buf BUF1 (N10222, N10221);
or OR2 (N10223, N10220, N9530);
and AND4 (N10224, N10212, N3620, N2167, N3543);
not NOT1 (N10225, N10199);
and AND2 (N10226, N10207, N7909);
xor XOR2 (N10227, N10223, N4109);
xor XOR2 (N10228, N10219, N1759);
nand NAND3 (N10229, N10216, N8766, N5976);
xor XOR2 (N10230, N10228, N3275);
and AND4 (N10231, N10226, N4100, N8046, N10223);
nor NOR3 (N10232, N10230, N2097, N200);
and AND2 (N10233, N10214, N8873);
xor XOR2 (N10234, N10229, N3334);
nor NOR3 (N10235, N10233, N6422, N4705);
nor NOR4 (N10236, N10224, N73, N278, N4973);
or OR4 (N10237, N10206, N8018, N10204, N8594);
nand NAND3 (N10238, N10235, N8476, N10203);
xor XOR2 (N10239, N10236, N7174);
or OR2 (N10240, N10231, N2579);
and AND2 (N10241, N10232, N7770);
not NOT1 (N10242, N10227);
or OR4 (N10243, N10241, N681, N9409, N1886);
not NOT1 (N10244, N10240);
or OR3 (N10245, N10238, N342, N1669);
xor XOR2 (N10246, N10242, N5729);
and AND2 (N10247, N10200, N806);
or OR4 (N10248, N10246, N2112, N8493, N6454);
not NOT1 (N10249, N10237);
not NOT1 (N10250, N10248);
and AND4 (N10251, N10239, N9268, N7403, N628);
not NOT1 (N10252, N10243);
xor XOR2 (N10253, N10245, N5150);
and AND3 (N10254, N10250, N391, N6696);
and AND3 (N10255, N10252, N3911, N7863);
nand NAND2 (N10256, N10249, N6263);
not NOT1 (N10257, N10234);
or OR3 (N10258, N10255, N6842, N4008);
not NOT1 (N10259, N10254);
nor NOR4 (N10260, N10258, N665, N2743, N8499);
or OR3 (N10261, N10257, N7180, N1260);
buf BUF1 (N10262, N10244);
nor NOR3 (N10263, N10259, N3647, N734);
not NOT1 (N10264, N10253);
nor NOR2 (N10265, N10247, N1266);
nand NAND3 (N10266, N10261, N1800, N3543);
nand NAND3 (N10267, N10264, N7317, N3193);
xor XOR2 (N10268, N10267, N3043);
not NOT1 (N10269, N10225);
buf BUF1 (N10270, N10265);
buf BUF1 (N10271, N10268);
or OR2 (N10272, N10222, N2724);
not NOT1 (N10273, N10256);
nand NAND2 (N10274, N10266, N2529);
nor NOR3 (N10275, N10269, N504, N5357);
or OR3 (N10276, N10272, N2945, N3464);
or OR2 (N10277, N10262, N4903);
or OR4 (N10278, N10275, N4918, N8431, N5673);
and AND4 (N10279, N10274, N10237, N7653, N983);
buf BUF1 (N10280, N10270);
and AND3 (N10281, N10251, N9473, N1049);
nand NAND3 (N10282, N10263, N6710, N9523);
nor NOR4 (N10283, N10260, N6653, N5158, N6466);
nor NOR2 (N10284, N10273, N8593);
and AND2 (N10285, N10271, N8820);
or OR2 (N10286, N10281, N3589);
not NOT1 (N10287, N10278);
and AND2 (N10288, N10280, N5596);
xor XOR2 (N10289, N10286, N9315);
buf BUF1 (N10290, N10282);
buf BUF1 (N10291, N10284);
buf BUF1 (N10292, N10289);
xor XOR2 (N10293, N10288, N3918);
xor XOR2 (N10294, N10290, N2042);
not NOT1 (N10295, N10292);
not NOT1 (N10296, N10295);
nand NAND3 (N10297, N10279, N1804, N4980);
nor NOR2 (N10298, N10291, N3496);
buf BUF1 (N10299, N10298);
or OR4 (N10300, N10296, N7097, N9377, N8237);
nor NOR3 (N10301, N10283, N3795, N2153);
xor XOR2 (N10302, N10297, N9000);
nand NAND4 (N10303, N10299, N2145, N8728, N5979);
or OR4 (N10304, N10301, N2826, N8349, N855);
or OR4 (N10305, N10287, N6593, N1101, N1197);
not NOT1 (N10306, N10277);
xor XOR2 (N10307, N10300, N7026);
nand NAND3 (N10308, N10304, N5411, N8056);
nor NOR4 (N10309, N10285, N8193, N987, N6578);
not NOT1 (N10310, N10307);
buf BUF1 (N10311, N10308);
nor NOR4 (N10312, N10302, N822, N3599, N4213);
nand NAND4 (N10313, N10311, N291, N2817, N8928);
and AND2 (N10314, N10294, N4094);
xor XOR2 (N10315, N10313, N6848);
xor XOR2 (N10316, N10293, N6502);
nand NAND2 (N10317, N10316, N1798);
or OR3 (N10318, N10312, N3795, N1015);
or OR2 (N10319, N10318, N4598);
xor XOR2 (N10320, N10306, N867);
xor XOR2 (N10321, N10314, N7324);
buf BUF1 (N10322, N10321);
xor XOR2 (N10323, N10309, N2879);
xor XOR2 (N10324, N10319, N2561);
xor XOR2 (N10325, N10322, N7813);
nor NOR2 (N10326, N10303, N9134);
xor XOR2 (N10327, N10317, N4711);
and AND3 (N10328, N10323, N2985, N6218);
nand NAND3 (N10329, N10315, N1504, N2686);
buf BUF1 (N10330, N10325);
xor XOR2 (N10331, N10276, N1921);
buf BUF1 (N10332, N10330);
xor XOR2 (N10333, N10310, N2866);
buf BUF1 (N10334, N10326);
nor NOR3 (N10335, N10320, N4286, N6296);
or OR2 (N10336, N10333, N258);
or OR3 (N10337, N10331, N9861, N9346);
buf BUF1 (N10338, N10334);
nor NOR3 (N10339, N10324, N5696, N4115);
or OR4 (N10340, N10335, N8048, N4413, N780);
and AND4 (N10341, N10339, N1635, N4433, N3692);
and AND3 (N10342, N10338, N649, N565);
xor XOR2 (N10343, N10336, N497);
buf BUF1 (N10344, N10305);
nand NAND4 (N10345, N10340, N6612, N7334, N60);
buf BUF1 (N10346, N10344);
nand NAND2 (N10347, N10346, N3991);
xor XOR2 (N10348, N10328, N11);
not NOT1 (N10349, N10347);
buf BUF1 (N10350, N10332);
buf BUF1 (N10351, N10343);
xor XOR2 (N10352, N10351, N6212);
buf BUF1 (N10353, N10342);
buf BUF1 (N10354, N10350);
nor NOR3 (N10355, N10329, N6214, N2873);
or OR2 (N10356, N10337, N8449);
or OR3 (N10357, N10327, N2188, N4263);
and AND4 (N10358, N10348, N5633, N6614, N1412);
nor NOR2 (N10359, N10349, N2621);
or OR4 (N10360, N10345, N4274, N2529, N1634);
nand NAND3 (N10361, N10356, N10247, N8690);
xor XOR2 (N10362, N10359, N7698);
nor NOR4 (N10363, N10354, N2382, N2902, N3387);
and AND2 (N10364, N10355, N2105);
not NOT1 (N10365, N10363);
nor NOR4 (N10366, N10353, N8429, N3057, N1326);
or OR3 (N10367, N10357, N6766, N10321);
xor XOR2 (N10368, N10358, N5414);
not NOT1 (N10369, N10360);
or OR2 (N10370, N10365, N4155);
not NOT1 (N10371, N10361);
nor NOR2 (N10372, N10341, N1023);
nor NOR2 (N10373, N10372, N7743);
nor NOR2 (N10374, N10352, N7120);
buf BUF1 (N10375, N10370);
xor XOR2 (N10376, N10375, N5339);
and AND3 (N10377, N10364, N5955, N6317);
buf BUF1 (N10378, N10368);
and AND2 (N10379, N10371, N63);
not NOT1 (N10380, N10379);
not NOT1 (N10381, N10380);
not NOT1 (N10382, N10381);
nand NAND4 (N10383, N10367, N802, N150, N6224);
not NOT1 (N10384, N10369);
not NOT1 (N10385, N10378);
or OR4 (N10386, N10382, N970, N9076, N4674);
xor XOR2 (N10387, N10386, N6577);
buf BUF1 (N10388, N10385);
not NOT1 (N10389, N10388);
not NOT1 (N10390, N10389);
xor XOR2 (N10391, N10383, N9867);
not NOT1 (N10392, N10390);
nor NOR4 (N10393, N10384, N43, N1926, N449);
or OR2 (N10394, N10393, N8306);
xor XOR2 (N10395, N10391, N748);
xor XOR2 (N10396, N10394, N3382);
buf BUF1 (N10397, N10366);
nor NOR4 (N10398, N10362, N53, N4153, N1958);
nand NAND2 (N10399, N10392, N8598);
xor XOR2 (N10400, N10376, N845);
and AND4 (N10401, N10373, N3512, N6280, N3743);
buf BUF1 (N10402, N10377);
or OR3 (N10403, N10374, N6774, N389);
buf BUF1 (N10404, N10398);
or OR2 (N10405, N10387, N9542);
or OR2 (N10406, N10405, N4826);
nor NOR4 (N10407, N10401, N5605, N8492, N10004);
nand NAND4 (N10408, N10402, N1732, N7840, N8588);
and AND3 (N10409, N10407, N9274, N2662);
xor XOR2 (N10410, N10409, N3548);
xor XOR2 (N10411, N10396, N2230);
buf BUF1 (N10412, N10408);
nor NOR4 (N10413, N10403, N8060, N702, N340);
and AND4 (N10414, N10400, N9340, N8387, N2105);
and AND4 (N10415, N10397, N7620, N9629, N5287);
not NOT1 (N10416, N10412);
and AND3 (N10417, N10411, N2003, N3415);
nor NOR3 (N10418, N10416, N3598, N9243);
not NOT1 (N10419, N10413);
nor NOR2 (N10420, N10406, N8296);
buf BUF1 (N10421, N10404);
buf BUF1 (N10422, N10419);
xor XOR2 (N10423, N10418, N9525);
not NOT1 (N10424, N10420);
nand NAND4 (N10425, N10417, N3410, N479, N1954);
nor NOR2 (N10426, N10414, N9316);
nand NAND2 (N10427, N10423, N2022);
not NOT1 (N10428, N10415);
nand NAND4 (N10429, N10399, N9480, N3316, N5030);
or OR4 (N10430, N10425, N9654, N8222, N787);
nand NAND2 (N10431, N10429, N423);
and AND2 (N10432, N10424, N2708);
not NOT1 (N10433, N10395);
nand NAND4 (N10434, N10430, N645, N2780, N3018);
and AND2 (N10435, N10427, N541);
buf BUF1 (N10436, N10432);
and AND4 (N10437, N10434, N1912, N1543, N3287);
xor XOR2 (N10438, N10435, N1809);
or OR2 (N10439, N10421, N729);
xor XOR2 (N10440, N10438, N4078);
nand NAND4 (N10441, N10422, N3838, N46, N5669);
or OR4 (N10442, N10436, N5957, N3516, N5636);
nand NAND3 (N10443, N10442, N8697, N2027);
or OR4 (N10444, N10431, N377, N9603, N8539);
nor NOR2 (N10445, N10440, N3628);
and AND3 (N10446, N10410, N6787, N2031);
xor XOR2 (N10447, N10428, N893);
and AND2 (N10448, N10437, N2620);
or OR4 (N10449, N10433, N5238, N5240, N8751);
nand NAND2 (N10450, N10439, N7463);
xor XOR2 (N10451, N10441, N4384);
buf BUF1 (N10452, N10449);
nand NAND3 (N10453, N10426, N2288, N4686);
nand NAND4 (N10454, N10445, N7035, N4518, N8966);
nor NOR3 (N10455, N10450, N10080, N6687);
buf BUF1 (N10456, N10455);
not NOT1 (N10457, N10453);
and AND4 (N10458, N10447, N3060, N9915, N5699);
and AND3 (N10459, N10458, N9253, N10319);
and AND2 (N10460, N10457, N4405);
xor XOR2 (N10461, N10448, N5806);
buf BUF1 (N10462, N10460);
nor NOR4 (N10463, N10462, N5672, N8798, N9562);
and AND4 (N10464, N10456, N9108, N497, N6677);
nor NOR4 (N10465, N10451, N4080, N5834, N6744);
not NOT1 (N10466, N10464);
nand NAND3 (N10467, N10463, N9747, N7715);
nor NOR2 (N10468, N10454, N4882);
or OR2 (N10469, N10459, N8197);
or OR3 (N10470, N10443, N1359, N6570);
buf BUF1 (N10471, N10452);
nand NAND4 (N10472, N10471, N5637, N2127, N4440);
or OR4 (N10473, N10465, N5422, N7226, N2859);
nor NOR3 (N10474, N10446, N4358, N6553);
nand NAND2 (N10475, N10473, N4820);
nor NOR4 (N10476, N10466, N8983, N8577, N7480);
buf BUF1 (N10477, N10467);
buf BUF1 (N10478, N10475);
xor XOR2 (N10479, N10444, N3184);
not NOT1 (N10480, N10469);
and AND3 (N10481, N10477, N8570, N2982);
buf BUF1 (N10482, N10478);
nand NAND4 (N10483, N10461, N5597, N8226, N704);
buf BUF1 (N10484, N10480);
not NOT1 (N10485, N10468);
nand NAND2 (N10486, N10470, N10394);
not NOT1 (N10487, N10472);
nor NOR2 (N10488, N10487, N1235);
and AND3 (N10489, N10481, N9248, N3718);
nand NAND2 (N10490, N10485, N4832);
nor NOR4 (N10491, N10482, N3503, N10034, N9342);
nand NAND4 (N10492, N10483, N1838, N6820, N10243);
buf BUF1 (N10493, N10490);
nand NAND3 (N10494, N10491, N3599, N7769);
or OR4 (N10495, N10493, N4284, N6646, N1496);
buf BUF1 (N10496, N10479);
or OR3 (N10497, N10489, N1965, N8460);
nand NAND3 (N10498, N10488, N8563, N4239);
not NOT1 (N10499, N10498);
not NOT1 (N10500, N10497);
xor XOR2 (N10501, N10496, N8383);
nor NOR4 (N10502, N10474, N4842, N8785, N4400);
buf BUF1 (N10503, N10476);
and AND3 (N10504, N10484, N1671, N1732);
nor NOR3 (N10505, N10502, N8151, N2776);
not NOT1 (N10506, N10504);
or OR3 (N10507, N10506, N4517, N9293);
nand NAND4 (N10508, N10501, N2660, N10165, N1140);
or OR2 (N10509, N10505, N1420);
xor XOR2 (N10510, N10509, N499);
xor XOR2 (N10511, N10495, N5053);
nor NOR4 (N10512, N10510, N8383, N3711, N1047);
and AND2 (N10513, N10511, N9613);
not NOT1 (N10514, N10486);
nor NOR3 (N10515, N10492, N4097, N5201);
xor XOR2 (N10516, N10514, N7823);
nor NOR3 (N10517, N10516, N5710, N184);
not NOT1 (N10518, N10503);
xor XOR2 (N10519, N10518, N5450);
buf BUF1 (N10520, N10494);
or OR3 (N10521, N10508, N2531, N3243);
and AND3 (N10522, N10513, N3940, N8554);
or OR4 (N10523, N10522, N6044, N616, N4369);
buf BUF1 (N10524, N10517);
buf BUF1 (N10525, N10515);
buf BUF1 (N10526, N10512);
nand NAND2 (N10527, N10507, N4983);
and AND2 (N10528, N10519, N5887);
xor XOR2 (N10529, N10525, N4657);
and AND3 (N10530, N10526, N1448, N500);
buf BUF1 (N10531, N10520);
xor XOR2 (N10532, N10528, N9068);
or OR4 (N10533, N10523, N7681, N83, N7598);
xor XOR2 (N10534, N10524, N6149);
or OR4 (N10535, N10521, N2534, N3087, N5390);
nor NOR2 (N10536, N10529, N2111);
not NOT1 (N10537, N10531);
xor XOR2 (N10538, N10537, N6921);
not NOT1 (N10539, N10527);
xor XOR2 (N10540, N10536, N36);
not NOT1 (N10541, N10538);
buf BUF1 (N10542, N10500);
nor NOR2 (N10543, N10541, N1617);
and AND3 (N10544, N10542, N8454, N7735);
or OR2 (N10545, N10539, N5423);
xor XOR2 (N10546, N10544, N9442);
or OR4 (N10547, N10532, N9451, N1646, N7294);
nand NAND2 (N10548, N10533, N1712);
nor NOR3 (N10549, N10540, N5300, N9381);
and AND2 (N10550, N10535, N446);
nand NAND4 (N10551, N10548, N6346, N8255, N3138);
and AND2 (N10552, N10545, N748);
and AND2 (N10553, N10546, N3319);
xor XOR2 (N10554, N10530, N6718);
buf BUF1 (N10555, N10543);
not NOT1 (N10556, N10551);
nor NOR3 (N10557, N10547, N8163, N3479);
and AND4 (N10558, N10549, N8103, N3066, N8159);
and AND3 (N10559, N10552, N1988, N8904);
buf BUF1 (N10560, N10555);
nor NOR3 (N10561, N10534, N1909, N589);
nor NOR4 (N10562, N10554, N7287, N5401, N399);
and AND4 (N10563, N10553, N6211, N1583, N9739);
nor NOR4 (N10564, N10561, N9582, N462, N10121);
or OR4 (N10565, N10558, N3892, N5916, N995);
not NOT1 (N10566, N10560);
or OR4 (N10567, N10550, N4240, N3516, N4759);
nand NAND3 (N10568, N10564, N7801, N6381);
or OR3 (N10569, N10565, N8306, N4988);
xor XOR2 (N10570, N10556, N7475);
xor XOR2 (N10571, N10559, N10520);
buf BUF1 (N10572, N10562);
xor XOR2 (N10573, N10571, N9113);
and AND2 (N10574, N10563, N3524);
xor XOR2 (N10575, N10574, N2193);
nor NOR3 (N10576, N10570, N4031, N2246);
not NOT1 (N10577, N10499);
and AND4 (N10578, N10567, N9798, N6514, N9814);
or OR4 (N10579, N10578, N8712, N2235, N4048);
and AND2 (N10580, N10575, N6772);
xor XOR2 (N10581, N10569, N3520);
or OR2 (N10582, N10572, N1613);
and AND4 (N10583, N10568, N2352, N9607, N271);
nand NAND4 (N10584, N10579, N4036, N8901, N4513);
nor NOR2 (N10585, N10581, N5944);
buf BUF1 (N10586, N10573);
buf BUF1 (N10587, N10584);
or OR2 (N10588, N10557, N8714);
xor XOR2 (N10589, N10586, N10404);
buf BUF1 (N10590, N10588);
not NOT1 (N10591, N10577);
not NOT1 (N10592, N10580);
nand NAND3 (N10593, N10576, N9954, N7385);
xor XOR2 (N10594, N10592, N8856);
xor XOR2 (N10595, N10587, N9632);
nor NOR4 (N10596, N10594, N529, N8526, N9155);
or OR4 (N10597, N10596, N1143, N5791, N9285);
buf BUF1 (N10598, N10566);
xor XOR2 (N10599, N10595, N281);
xor XOR2 (N10600, N10590, N4519);
and AND4 (N10601, N10593, N10019, N8948, N5881);
nand NAND4 (N10602, N10597, N7943, N2753, N1822);
nor NOR3 (N10603, N10585, N10058, N7341);
nor NOR4 (N10604, N10591, N1991, N4581, N7404);
or OR3 (N10605, N10598, N3579, N5459);
not NOT1 (N10606, N10605);
nor NOR4 (N10607, N10599, N9078, N511, N7197);
nand NAND3 (N10608, N10603, N8279, N8563);
and AND4 (N10609, N10607, N9838, N3418, N6617);
not NOT1 (N10610, N10608);
nand NAND2 (N10611, N10610, N6727);
and AND2 (N10612, N10582, N2678);
xor XOR2 (N10613, N10604, N8696);
and AND3 (N10614, N10589, N4972, N293);
nand NAND2 (N10615, N10614, N3606);
nand NAND3 (N10616, N10613, N1841, N3882);
xor XOR2 (N10617, N10601, N9404);
and AND4 (N10618, N10616, N7643, N8283, N1494);
nor NOR3 (N10619, N10617, N970, N1010);
nor NOR4 (N10620, N10609, N9277, N6291, N7328);
xor XOR2 (N10621, N10612, N3639);
not NOT1 (N10622, N10620);
or OR3 (N10623, N10622, N3147, N1176);
not NOT1 (N10624, N10611);
buf BUF1 (N10625, N10623);
and AND3 (N10626, N10625, N2363, N4799);
or OR2 (N10627, N10600, N2761);
not NOT1 (N10628, N10619);
not NOT1 (N10629, N10624);
nor NOR4 (N10630, N10583, N2054, N6703, N6122);
nand NAND3 (N10631, N10602, N5786, N3095);
nor NOR2 (N10632, N10615, N8078);
and AND2 (N10633, N10626, N3669);
buf BUF1 (N10634, N10627);
or OR3 (N10635, N10633, N9290, N4111);
nor NOR3 (N10636, N10618, N990, N3948);
buf BUF1 (N10637, N10635);
not NOT1 (N10638, N10634);
xor XOR2 (N10639, N10621, N6887);
nor NOR2 (N10640, N10632, N4719);
and AND4 (N10641, N10628, N5010, N627, N5034);
or OR2 (N10642, N10630, N7480);
or OR4 (N10643, N10638, N2328, N8506, N3865);
not NOT1 (N10644, N10642);
xor XOR2 (N10645, N10636, N6924);
nand NAND2 (N10646, N10637, N3045);
xor XOR2 (N10647, N10606, N10161);
nor NOR2 (N10648, N10640, N5145);
and AND2 (N10649, N10631, N425);
not NOT1 (N10650, N10639);
xor XOR2 (N10651, N10648, N3392);
not NOT1 (N10652, N10647);
or OR2 (N10653, N10646, N5493);
nor NOR3 (N10654, N10653, N10571, N5649);
and AND4 (N10655, N10643, N5882, N6248, N1546);
and AND4 (N10656, N10652, N7216, N3968, N578);
xor XOR2 (N10657, N10655, N4939);
nand NAND2 (N10658, N10650, N730);
nand NAND2 (N10659, N10658, N7470);
or OR3 (N10660, N10656, N5907, N7434);
buf BUF1 (N10661, N10654);
or OR2 (N10662, N10629, N1311);
and AND3 (N10663, N10641, N4, N10404);
nand NAND4 (N10664, N10660, N9279, N4198, N10239);
not NOT1 (N10665, N10657);
buf BUF1 (N10666, N10662);
and AND4 (N10667, N10651, N3998, N1549, N5537);
and AND3 (N10668, N10645, N7110, N2464);
or OR2 (N10669, N10644, N8937);
xor XOR2 (N10670, N10668, N2252);
and AND3 (N10671, N10669, N1264, N8323);
or OR2 (N10672, N10663, N4973);
not NOT1 (N10673, N10670);
or OR3 (N10674, N10659, N9014, N7729);
or OR2 (N10675, N10664, N5607);
and AND3 (N10676, N10675, N3406, N2152);
not NOT1 (N10677, N10673);
buf BUF1 (N10678, N10666);
xor XOR2 (N10679, N10677, N1906);
or OR3 (N10680, N10674, N593, N4041);
nor NOR4 (N10681, N10679, N2549, N8850, N10199);
buf BUF1 (N10682, N10681);
buf BUF1 (N10683, N10661);
nand NAND4 (N10684, N10676, N7789, N4604, N9204);
buf BUF1 (N10685, N10665);
or OR2 (N10686, N10672, N8927);
and AND3 (N10687, N10671, N3564, N9417);
nand NAND2 (N10688, N10682, N9165);
or OR4 (N10689, N10687, N2129, N2958, N2424);
not NOT1 (N10690, N10649);
xor XOR2 (N10691, N10667, N8377);
xor XOR2 (N10692, N10689, N5212);
not NOT1 (N10693, N10678);
xor XOR2 (N10694, N10692, N4279);
and AND3 (N10695, N10694, N7631, N6322);
or OR3 (N10696, N10690, N203, N7731);
nor NOR2 (N10697, N10686, N9364);
and AND3 (N10698, N10693, N4518, N5418);
not NOT1 (N10699, N10691);
buf BUF1 (N10700, N10696);
buf BUF1 (N10701, N10685);
nor NOR3 (N10702, N10688, N7987, N807);
buf BUF1 (N10703, N10680);
not NOT1 (N10704, N10695);
not NOT1 (N10705, N10698);
and AND3 (N10706, N10702, N5469, N9537);
and AND4 (N10707, N10704, N6334, N7715, N1326);
xor XOR2 (N10708, N10701, N10607);
and AND4 (N10709, N10683, N4958, N8709, N2057);
or OR4 (N10710, N10700, N6258, N3375, N4510);
buf BUF1 (N10711, N10697);
nand NAND2 (N10712, N10703, N2587);
buf BUF1 (N10713, N10705);
or OR4 (N10714, N10712, N4205, N6895, N8225);
not NOT1 (N10715, N10707);
not NOT1 (N10716, N10708);
buf BUF1 (N10717, N10714);
not NOT1 (N10718, N10711);
nand NAND3 (N10719, N10715, N5554, N5207);
xor XOR2 (N10720, N10684, N6513);
nor NOR3 (N10721, N10709, N7793, N612);
not NOT1 (N10722, N10719);
buf BUF1 (N10723, N10720);
xor XOR2 (N10724, N10706, N10043);
and AND4 (N10725, N10724, N10455, N409, N6587);
or OR2 (N10726, N10713, N281);
or OR3 (N10727, N10722, N7777, N1031);
and AND2 (N10728, N10723, N7716);
or OR2 (N10729, N10727, N8942);
xor XOR2 (N10730, N10728, N10568);
or OR3 (N10731, N10726, N1129, N1275);
nand NAND2 (N10732, N10729, N3477);
buf BUF1 (N10733, N10716);
not NOT1 (N10734, N10733);
nand NAND2 (N10735, N10699, N4057);
and AND4 (N10736, N10717, N9894, N4620, N10604);
xor XOR2 (N10737, N10710, N8780);
nand NAND3 (N10738, N10734, N1766, N4497);
not NOT1 (N10739, N10738);
nor NOR2 (N10740, N10737, N739);
xor XOR2 (N10741, N10721, N2102);
xor XOR2 (N10742, N10740, N6563);
xor XOR2 (N10743, N10736, N7206);
and AND3 (N10744, N10743, N7252, N10020);
or OR3 (N10745, N10730, N7360, N1383);
nand NAND3 (N10746, N10735, N9477, N4275);
not NOT1 (N10747, N10741);
and AND2 (N10748, N10725, N1123);
and AND2 (N10749, N10718, N9846);
and AND4 (N10750, N10739, N6943, N1662, N3278);
nand NAND3 (N10751, N10750, N6782, N1533);
nand NAND3 (N10752, N10742, N5965, N934);
buf BUF1 (N10753, N10731);
buf BUF1 (N10754, N10746);
not NOT1 (N10755, N10753);
nor NOR4 (N10756, N10752, N912, N8004, N2231);
buf BUF1 (N10757, N10744);
nand NAND2 (N10758, N10747, N489);
nor NOR4 (N10759, N10748, N7855, N10416, N9608);
nor NOR4 (N10760, N10745, N3907, N7083, N6026);
xor XOR2 (N10761, N10732, N833);
nor NOR4 (N10762, N10756, N6856, N1780, N7097);
buf BUF1 (N10763, N10759);
or OR3 (N10764, N10751, N8112, N5911);
nor NOR2 (N10765, N10755, N8998);
xor XOR2 (N10766, N10762, N7255);
buf BUF1 (N10767, N10757);
or OR2 (N10768, N10763, N1044);
xor XOR2 (N10769, N10767, N6219);
xor XOR2 (N10770, N10760, N1027);
xor XOR2 (N10771, N10766, N5116);
nor NOR2 (N10772, N10749, N7913);
not NOT1 (N10773, N10761);
and AND3 (N10774, N10764, N6692, N3055);
nor NOR2 (N10775, N10772, N8278);
nor NOR3 (N10776, N10765, N1444, N1725);
nand NAND4 (N10777, N10768, N7555, N10024, N2146);
and AND3 (N10778, N10758, N5704, N10734);
nor NOR2 (N10779, N10771, N7687);
and AND3 (N10780, N10769, N787, N1269);
nor NOR3 (N10781, N10779, N2028, N10199);
xor XOR2 (N10782, N10775, N7450);
buf BUF1 (N10783, N10776);
nor NOR4 (N10784, N10781, N6665, N8679, N1939);
and AND2 (N10785, N10773, N3278);
not NOT1 (N10786, N10785);
and AND2 (N10787, N10784, N1129);
nand NAND3 (N10788, N10774, N6802, N1070);
nand NAND2 (N10789, N10778, N2922);
and AND2 (N10790, N10782, N2416);
or OR2 (N10791, N10788, N8229);
nor NOR4 (N10792, N10783, N4618, N2433, N541);
buf BUF1 (N10793, N10787);
buf BUF1 (N10794, N10792);
and AND4 (N10795, N10780, N331, N295, N3072);
nor NOR4 (N10796, N10770, N5108, N8037, N3600);
nor NOR4 (N10797, N10791, N4327, N5791, N3547);
xor XOR2 (N10798, N10794, N1968);
nand NAND2 (N10799, N10786, N3061);
buf BUF1 (N10800, N10754);
buf BUF1 (N10801, N10793);
not NOT1 (N10802, N10789);
not NOT1 (N10803, N10802);
nor NOR2 (N10804, N10790, N2131);
and AND4 (N10805, N10797, N7973, N230, N1977);
or OR3 (N10806, N10798, N5865, N4312);
buf BUF1 (N10807, N10801);
or OR3 (N10808, N10807, N4823, N8534);
and AND3 (N10809, N10777, N4766, N1012);
not NOT1 (N10810, N10796);
nand NAND4 (N10811, N10799, N10539, N2448, N2574);
buf BUF1 (N10812, N10809);
buf BUF1 (N10813, N10808);
and AND2 (N10814, N10811, N5010);
nand NAND4 (N10815, N10800, N10427, N4052, N3436);
nand NAND2 (N10816, N10806, N6251);
not NOT1 (N10817, N10804);
nand NAND2 (N10818, N10810, N4712);
or OR3 (N10819, N10805, N10124, N4297);
or OR2 (N10820, N10816, N1095);
buf BUF1 (N10821, N10803);
xor XOR2 (N10822, N10817, N1762);
nand NAND2 (N10823, N10818, N4761);
nor NOR2 (N10824, N10820, N10038);
buf BUF1 (N10825, N10821);
nand NAND4 (N10826, N10815, N9129, N3271, N1144);
buf BUF1 (N10827, N10822);
not NOT1 (N10828, N10814);
and AND2 (N10829, N10813, N9491);
not NOT1 (N10830, N10828);
and AND3 (N10831, N10825, N8238, N3999);
xor XOR2 (N10832, N10831, N4786);
nand NAND2 (N10833, N10829, N8860);
buf BUF1 (N10834, N10830);
buf BUF1 (N10835, N10832);
and AND4 (N10836, N10795, N2140, N4549, N8424);
and AND3 (N10837, N10823, N7313, N214);
nand NAND4 (N10838, N10824, N9593, N332, N2174);
nand NAND4 (N10839, N10833, N4256, N4641, N7609);
nor NOR2 (N10840, N10838, N5655);
or OR2 (N10841, N10835, N3949);
nand NAND3 (N10842, N10826, N8401, N3287);
not NOT1 (N10843, N10837);
or OR4 (N10844, N10827, N3446, N2980, N7257);
nor NOR4 (N10845, N10844, N814, N8415, N1791);
or OR4 (N10846, N10841, N2144, N2785, N2899);
xor XOR2 (N10847, N10812, N2368);
or OR4 (N10848, N10836, N1554, N5678, N6529);
nor NOR3 (N10849, N10847, N4508, N2820);
nor NOR3 (N10850, N10842, N7119, N1082);
xor XOR2 (N10851, N10845, N6876);
or OR4 (N10852, N10846, N10005, N1099, N8397);
xor XOR2 (N10853, N10840, N2419);
not NOT1 (N10854, N10834);
nand NAND4 (N10855, N10848, N7331, N912, N10125);
or OR2 (N10856, N10852, N9340);
buf BUF1 (N10857, N10849);
or OR2 (N10858, N10853, N3411);
buf BUF1 (N10859, N10850);
nand NAND2 (N10860, N10843, N6186);
or OR2 (N10861, N10860, N10439);
and AND3 (N10862, N10861, N6544, N4463);
and AND3 (N10863, N10856, N5845, N5896);
buf BUF1 (N10864, N10839);
nand NAND2 (N10865, N10862, N6244);
xor XOR2 (N10866, N10864, N6555);
nor NOR3 (N10867, N10854, N9670, N7462);
nor NOR2 (N10868, N10863, N3990);
and AND3 (N10869, N10851, N2948, N6523);
not NOT1 (N10870, N10868);
or OR4 (N10871, N10855, N6542, N2246, N9251);
nand NAND2 (N10872, N10871, N6090);
xor XOR2 (N10873, N10858, N3987);
not NOT1 (N10874, N10866);
or OR3 (N10875, N10869, N9631, N9857);
xor XOR2 (N10876, N10819, N3057);
nand NAND3 (N10877, N10867, N1712, N10291);
nand NAND2 (N10878, N10865, N10517);
xor XOR2 (N10879, N10878, N3974);
buf BUF1 (N10880, N10875);
buf BUF1 (N10881, N10857);
or OR2 (N10882, N10881, N1474);
and AND2 (N10883, N10882, N1795);
buf BUF1 (N10884, N10874);
nor NOR2 (N10885, N10877, N1304);
nor NOR3 (N10886, N10870, N1248, N1558);
not NOT1 (N10887, N10859);
buf BUF1 (N10888, N10887);
xor XOR2 (N10889, N10880, N5229);
nor NOR4 (N10890, N10885, N135, N1342, N5660);
nor NOR3 (N10891, N10872, N5823, N2801);
nor NOR2 (N10892, N10888, N8515);
xor XOR2 (N10893, N10873, N2705);
not NOT1 (N10894, N10883);
and AND2 (N10895, N10893, N6081);
xor XOR2 (N10896, N10891, N2148);
not NOT1 (N10897, N10889);
not NOT1 (N10898, N10897);
xor XOR2 (N10899, N10886, N6263);
nor NOR3 (N10900, N10895, N7501, N7024);
or OR3 (N10901, N10884, N5719, N5792);
and AND3 (N10902, N10896, N10451, N8699);
buf BUF1 (N10903, N10898);
nand NAND3 (N10904, N10890, N8325, N5671);
xor XOR2 (N10905, N10879, N5356);
xor XOR2 (N10906, N10900, N4767);
nor NOR4 (N10907, N10906, N4234, N8964, N1602);
nand NAND2 (N10908, N10907, N8178);
and AND3 (N10909, N10905, N6751, N8324);
xor XOR2 (N10910, N10899, N7384);
nand NAND4 (N10911, N10902, N4871, N6563, N9390);
and AND2 (N10912, N10910, N5870);
or OR4 (N10913, N10911, N179, N2671, N559);
or OR3 (N10914, N10892, N5824, N10337);
nand NAND2 (N10915, N10908, N135);
nor NOR3 (N10916, N10915, N839, N274);
or OR3 (N10917, N10913, N1830, N534);
or OR2 (N10918, N10909, N6622);
or OR3 (N10919, N10903, N8568, N1392);
nor NOR4 (N10920, N10904, N2879, N8132, N8941);
nor NOR4 (N10921, N10894, N9098, N10874, N4049);
or OR4 (N10922, N10920, N203, N10713, N2752);
and AND3 (N10923, N10912, N5123, N9196);
or OR2 (N10924, N10919, N3852);
nand NAND2 (N10925, N10917, N9233);
xor XOR2 (N10926, N10923, N10494);
buf BUF1 (N10927, N10918);
and AND2 (N10928, N10926, N2541);
and AND4 (N10929, N10927, N8741, N358, N6491);
nor NOR3 (N10930, N10876, N10602, N6717);
nor NOR3 (N10931, N10914, N9324, N10912);
not NOT1 (N10932, N10931);
nand NAND3 (N10933, N10901, N7943, N4061);
and AND2 (N10934, N10929, N6233);
nor NOR3 (N10935, N10933, N1042, N6320);
or OR3 (N10936, N10916, N5043, N986);
not NOT1 (N10937, N10921);
nand NAND3 (N10938, N10934, N4912, N9250);
buf BUF1 (N10939, N10922);
or OR2 (N10940, N10925, N10778);
and AND2 (N10941, N10939, N4263);
buf BUF1 (N10942, N10937);
nor NOR3 (N10943, N10938, N4787, N1458);
and AND3 (N10944, N10928, N7153, N5473);
xor XOR2 (N10945, N10936, N2065);
or OR4 (N10946, N10924, N253, N3453, N1729);
xor XOR2 (N10947, N10940, N3279);
buf BUF1 (N10948, N10941);
nor NOR3 (N10949, N10944, N9442, N1517);
nor NOR3 (N10950, N10945, N300, N10872);
nor NOR4 (N10951, N10935, N9998, N5450, N5020);
nor NOR2 (N10952, N10948, N6986);
not NOT1 (N10953, N10952);
buf BUF1 (N10954, N10951);
not NOT1 (N10955, N10932);
or OR3 (N10956, N10942, N1214, N6946);
nor NOR3 (N10957, N10947, N8318, N7152);
buf BUF1 (N10958, N10955);
or OR4 (N10959, N10953, N4269, N10565, N2856);
and AND2 (N10960, N10957, N1955);
and AND4 (N10961, N10959, N5649, N7322, N4639);
buf BUF1 (N10962, N10960);
or OR2 (N10963, N10950, N9298);
or OR3 (N10964, N10949, N7391, N10168);
nand NAND4 (N10965, N10964, N6309, N5925, N2820);
buf BUF1 (N10966, N10965);
xor XOR2 (N10967, N10930, N227);
nor NOR2 (N10968, N10962, N8178);
nor NOR2 (N10969, N10956, N4568);
buf BUF1 (N10970, N10966);
or OR3 (N10971, N10954, N2457, N4375);
xor XOR2 (N10972, N10967, N2271);
and AND4 (N10973, N10970, N3488, N6860, N1636);
or OR4 (N10974, N10963, N1539, N10590, N5510);
or OR2 (N10975, N10943, N9138);
buf BUF1 (N10976, N10946);
xor XOR2 (N10977, N10975, N7132);
nor NOR4 (N10978, N10977, N5314, N6717, N8291);
and AND2 (N10979, N10972, N7633);
not NOT1 (N10980, N10961);
buf BUF1 (N10981, N10958);
nand NAND4 (N10982, N10971, N9612, N1301, N9025);
and AND2 (N10983, N10969, N9095);
xor XOR2 (N10984, N10973, N8251);
xor XOR2 (N10985, N10974, N1471);
nor NOR4 (N10986, N10983, N6907, N1499, N1364);
xor XOR2 (N10987, N10968, N361);
not NOT1 (N10988, N10987);
buf BUF1 (N10989, N10988);
nand NAND4 (N10990, N10989, N3748, N10698, N2767);
or OR2 (N10991, N10976, N581);
buf BUF1 (N10992, N10991);
buf BUF1 (N10993, N10978);
nand NAND2 (N10994, N10982, N8314);
not NOT1 (N10995, N10990);
or OR3 (N10996, N10985, N6449, N10407);
nor NOR2 (N10997, N10996, N7035);
buf BUF1 (N10998, N10979);
not NOT1 (N10999, N10994);
not NOT1 (N11000, N10998);
or OR2 (N11001, N10980, N9192);
or OR4 (N11002, N10995, N3851, N210, N2977);
buf BUF1 (N11003, N10984);
xor XOR2 (N11004, N11003, N8272);
nand NAND4 (N11005, N11000, N9649, N3291, N8981);
nor NOR3 (N11006, N10997, N1367, N5778);
xor XOR2 (N11007, N10999, N7818);
nor NOR4 (N11008, N10986, N7175, N4896, N8142);
xor XOR2 (N11009, N11008, N9876);
nand NAND4 (N11010, N10981, N10941, N3188, N3247);
or OR2 (N11011, N11005, N4338);
and AND3 (N11012, N11004, N7897, N3445);
xor XOR2 (N11013, N11012, N4700);
or OR2 (N11014, N10992, N1469);
buf BUF1 (N11015, N11009);
nor NOR2 (N11016, N11006, N2035);
xor XOR2 (N11017, N11011, N10526);
xor XOR2 (N11018, N11015, N724);
or OR3 (N11019, N11002, N6620, N747);
nor NOR2 (N11020, N11018, N9394);
and AND2 (N11021, N11020, N5250);
xor XOR2 (N11022, N11001, N6894);
nor NOR4 (N11023, N11010, N4544, N10789, N9514);
xor XOR2 (N11024, N11023, N1324);
not NOT1 (N11025, N11007);
buf BUF1 (N11026, N11016);
and AND4 (N11027, N11019, N7979, N4962, N1492);
and AND2 (N11028, N11024, N3792);
xor XOR2 (N11029, N11021, N5321);
nor NOR3 (N11030, N11026, N8229, N3223);
not NOT1 (N11031, N11022);
or OR3 (N11032, N11017, N2976, N2285);
not NOT1 (N11033, N11029);
buf BUF1 (N11034, N11033);
not NOT1 (N11035, N11028);
not NOT1 (N11036, N11032);
and AND3 (N11037, N11036, N406, N4599);
buf BUF1 (N11038, N11025);
not NOT1 (N11039, N11035);
nor NOR3 (N11040, N11031, N3972, N8706);
nor NOR2 (N11041, N10993, N2957);
not NOT1 (N11042, N11014);
buf BUF1 (N11043, N11038);
or OR4 (N11044, N11043, N10230, N1618, N7408);
and AND4 (N11045, N11039, N9269, N9662, N7875);
not NOT1 (N11046, N11044);
xor XOR2 (N11047, N11045, N3384);
nand NAND2 (N11048, N11041, N9426);
nor NOR3 (N11049, N11046, N1079, N4934);
and AND3 (N11050, N11034, N4014, N42);
xor XOR2 (N11051, N11027, N6076);
xor XOR2 (N11052, N11037, N8910);
and AND3 (N11053, N11047, N9559, N7942);
and AND2 (N11054, N11049, N5257);
or OR2 (N11055, N11053, N1458);
buf BUF1 (N11056, N11040);
xor XOR2 (N11057, N11042, N3691);
xor XOR2 (N11058, N11056, N7643);
or OR3 (N11059, N11057, N10006, N5424);
nor NOR3 (N11060, N11048, N7869, N789);
and AND3 (N11061, N11060, N4706, N5527);
buf BUF1 (N11062, N11030);
not NOT1 (N11063, N11062);
nor NOR4 (N11064, N11054, N3717, N10178, N6835);
and AND3 (N11065, N11063, N4445, N10565);
nor NOR3 (N11066, N11055, N4421, N6328);
xor XOR2 (N11067, N11065, N1664);
buf BUF1 (N11068, N11050);
xor XOR2 (N11069, N11066, N10728);
nand NAND4 (N11070, N11064, N6946, N2522, N875);
nor NOR2 (N11071, N11067, N10385);
buf BUF1 (N11072, N11068);
xor XOR2 (N11073, N11058, N1013);
buf BUF1 (N11074, N11013);
not NOT1 (N11075, N11059);
nand NAND2 (N11076, N11072, N3871);
xor XOR2 (N11077, N11051, N1923);
nand NAND4 (N11078, N11070, N1185, N9064, N4094);
or OR3 (N11079, N11052, N8398, N3490);
not NOT1 (N11080, N11079);
or OR3 (N11081, N11076, N10264, N245);
buf BUF1 (N11082, N11078);
nor NOR4 (N11083, N11080, N4536, N4980, N8556);
or OR3 (N11084, N11082, N1605, N4710);
nand NAND2 (N11085, N11061, N1361);
and AND4 (N11086, N11071, N4185, N3213, N9840);
buf BUF1 (N11087, N11075);
xor XOR2 (N11088, N11074, N7152);
not NOT1 (N11089, N11087);
or OR2 (N11090, N11081, N7029);
and AND2 (N11091, N11090, N3663);
xor XOR2 (N11092, N11077, N5318);
nand NAND4 (N11093, N11092, N7004, N2993, N7883);
or OR4 (N11094, N11073, N3654, N5613, N3610);
nand NAND3 (N11095, N11085, N1403, N5026);
nand NAND2 (N11096, N11069, N3160);
buf BUF1 (N11097, N11095);
nor NOR2 (N11098, N11094, N6700);
nor NOR4 (N11099, N11098, N74, N6593, N5389);
not NOT1 (N11100, N11091);
not NOT1 (N11101, N11097);
nor NOR4 (N11102, N11100, N7300, N9199, N9837);
buf BUF1 (N11103, N11101);
buf BUF1 (N11104, N11102);
buf BUF1 (N11105, N11083);
nor NOR3 (N11106, N11084, N1645, N5921);
nand NAND4 (N11107, N11099, N5259, N5857, N4432);
and AND3 (N11108, N11106, N5178, N5863);
and AND3 (N11109, N11103, N8151, N10884);
buf BUF1 (N11110, N11086);
or OR2 (N11111, N11089, N10578);
nand NAND2 (N11112, N11108, N5878);
and AND3 (N11113, N11105, N240, N10981);
not NOT1 (N11114, N11113);
or OR4 (N11115, N11114, N5609, N9281, N1796);
nand NAND3 (N11116, N11111, N3487, N4215);
and AND3 (N11117, N11107, N7950, N6439);
and AND3 (N11118, N11110, N480, N9206);
xor XOR2 (N11119, N11117, N5075);
or OR3 (N11120, N11109, N4459, N6334);
and AND4 (N11121, N11118, N5281, N5905, N6318);
nand NAND4 (N11122, N11104, N6503, N7733, N8730);
nor NOR3 (N11123, N11119, N7102, N2129);
not NOT1 (N11124, N11116);
buf BUF1 (N11125, N11124);
xor XOR2 (N11126, N11120, N9617);
and AND4 (N11127, N11125, N616, N8048, N6522);
nand NAND2 (N11128, N11112, N3045);
nand NAND2 (N11129, N11123, N8482);
xor XOR2 (N11130, N11122, N10908);
buf BUF1 (N11131, N11126);
xor XOR2 (N11132, N11088, N7378);
nor NOR3 (N11133, N11115, N1760, N7992);
not NOT1 (N11134, N11130);
not NOT1 (N11135, N11096);
nand NAND4 (N11136, N11134, N8906, N10312, N9911);
nor NOR4 (N11137, N11135, N8211, N5786, N8145);
xor XOR2 (N11138, N11127, N6491);
not NOT1 (N11139, N11121);
nor NOR2 (N11140, N11131, N2311);
nor NOR3 (N11141, N11128, N5111, N10737);
xor XOR2 (N11142, N11133, N5013);
not NOT1 (N11143, N11138);
xor XOR2 (N11144, N11093, N6539);
buf BUF1 (N11145, N11142);
not NOT1 (N11146, N11136);
buf BUF1 (N11147, N11143);
nor NOR2 (N11148, N11146, N498);
nand NAND3 (N11149, N11129, N693, N2348);
not NOT1 (N11150, N11147);
or OR2 (N11151, N11145, N8738);
and AND4 (N11152, N11140, N5263, N5436, N4102);
nor NOR3 (N11153, N11150, N547, N1933);
nand NAND4 (N11154, N11144, N4745, N4558, N2336);
buf BUF1 (N11155, N11132);
nor NOR3 (N11156, N11155, N6648, N10546);
buf BUF1 (N11157, N11139);
nor NOR2 (N11158, N11149, N4385);
or OR3 (N11159, N11157, N10408, N4289);
buf BUF1 (N11160, N11156);
nand NAND3 (N11161, N11154, N6608, N11072);
nand NAND4 (N11162, N11153, N8571, N7591, N11012);
or OR3 (N11163, N11151, N705, N5807);
buf BUF1 (N11164, N11161);
not NOT1 (N11165, N11164);
or OR4 (N11166, N11148, N7826, N3121, N1234);
not NOT1 (N11167, N11160);
nand NAND4 (N11168, N11163, N5493, N10216, N11044);
nand NAND3 (N11169, N11159, N4285, N2456);
xor XOR2 (N11170, N11168, N5158);
xor XOR2 (N11171, N11137, N4923);
or OR2 (N11172, N11171, N6480);
or OR4 (N11173, N11166, N1637, N10955, N4436);
not NOT1 (N11174, N11167);
buf BUF1 (N11175, N11141);
nor NOR3 (N11176, N11169, N4658, N5593);
nand NAND2 (N11177, N11162, N3180);
buf BUF1 (N11178, N11172);
and AND4 (N11179, N11175, N8195, N9179, N10394);
buf BUF1 (N11180, N11152);
or OR3 (N11181, N11180, N7855, N544);
not NOT1 (N11182, N11165);
and AND3 (N11183, N11174, N5206, N909);
not NOT1 (N11184, N11170);
or OR4 (N11185, N11158, N4663, N3, N1708);
xor XOR2 (N11186, N11185, N643);
nand NAND2 (N11187, N11179, N8743);
xor XOR2 (N11188, N11181, N8716);
nor NOR4 (N11189, N11188, N3595, N4968, N6175);
nor NOR4 (N11190, N11176, N5069, N10995, N10037);
and AND4 (N11191, N11184, N4325, N6339, N10733);
xor XOR2 (N11192, N11178, N130);
xor XOR2 (N11193, N11183, N8796);
buf BUF1 (N11194, N11193);
nand NAND4 (N11195, N11187, N2819, N6334, N4715);
not NOT1 (N11196, N11189);
nor NOR4 (N11197, N11191, N6201, N1042, N6553);
buf BUF1 (N11198, N11192);
or OR2 (N11199, N11198, N11139);
or OR4 (N11200, N11199, N10019, N4135, N4533);
and AND3 (N11201, N11195, N9669, N5853);
and AND2 (N11202, N11200, N9107);
not NOT1 (N11203, N11182);
xor XOR2 (N11204, N11177, N8928);
or OR4 (N11205, N11201, N6455, N1481, N9507);
and AND4 (N11206, N11196, N4161, N1428, N4233);
or OR2 (N11207, N11186, N6453);
xor XOR2 (N11208, N11190, N7868);
xor XOR2 (N11209, N11207, N9028);
and AND2 (N11210, N11173, N1630);
and AND2 (N11211, N11203, N5242);
and AND2 (N11212, N11209, N5977);
nand NAND2 (N11213, N11206, N273);
xor XOR2 (N11214, N11211, N1022);
buf BUF1 (N11215, N11194);
not NOT1 (N11216, N11202);
xor XOR2 (N11217, N11216, N8060);
buf BUF1 (N11218, N11208);
nor NOR2 (N11219, N11205, N4051);
and AND3 (N11220, N11213, N4541, N7856);
and AND4 (N11221, N11220, N9372, N5632, N10300);
nor NOR2 (N11222, N11214, N3556);
nand NAND2 (N11223, N11218, N10039);
nor NOR3 (N11224, N11222, N2827, N2260);
nor NOR2 (N11225, N11223, N5115);
not NOT1 (N11226, N11212);
xor XOR2 (N11227, N11217, N5483);
and AND4 (N11228, N11204, N7640, N5606, N413);
nor NOR2 (N11229, N11210, N9684);
nand NAND4 (N11230, N11225, N4814, N9242, N4423);
or OR2 (N11231, N11227, N10506);
or OR3 (N11232, N11226, N3188, N3809);
not NOT1 (N11233, N11224);
not NOT1 (N11234, N11230);
xor XOR2 (N11235, N11229, N3015);
nand NAND2 (N11236, N11197, N5233);
xor XOR2 (N11237, N11215, N4921);
and AND4 (N11238, N11232, N7622, N3056, N6141);
xor XOR2 (N11239, N11234, N7698);
nor NOR4 (N11240, N11239, N10910, N3550, N6072);
buf BUF1 (N11241, N11238);
nor NOR3 (N11242, N11233, N7684, N1671);
buf BUF1 (N11243, N11240);
xor XOR2 (N11244, N11219, N292);
buf BUF1 (N11245, N11221);
and AND4 (N11246, N11231, N2373, N9673, N232);
nor NOR2 (N11247, N11236, N10269);
not NOT1 (N11248, N11246);
buf BUF1 (N11249, N11243);
nor NOR4 (N11250, N11235, N4787, N10421, N4541);
buf BUF1 (N11251, N11248);
not NOT1 (N11252, N11249);
buf BUF1 (N11253, N11252);
nor NOR3 (N11254, N11245, N8647, N788);
not NOT1 (N11255, N11254);
not NOT1 (N11256, N11253);
nor NOR4 (N11257, N11242, N7701, N10566, N1029);
xor XOR2 (N11258, N11244, N8278);
nor NOR3 (N11259, N11257, N643, N5349);
xor XOR2 (N11260, N11247, N1497);
not NOT1 (N11261, N11250);
or OR3 (N11262, N11258, N2889, N319);
and AND2 (N11263, N11251, N6121);
nand NAND2 (N11264, N11237, N956);
or OR4 (N11265, N11255, N9963, N6568, N3841);
and AND3 (N11266, N11263, N555, N5706);
nor NOR4 (N11267, N11264, N1445, N6717, N5769);
nor NOR4 (N11268, N11266, N1532, N7266, N1519);
xor XOR2 (N11269, N11265, N6649);
buf BUF1 (N11270, N11269);
nor NOR4 (N11271, N11228, N141, N3172, N5573);
nor NOR3 (N11272, N11259, N10489, N10506);
not NOT1 (N11273, N11260);
xor XOR2 (N11274, N11262, N7474);
not NOT1 (N11275, N11271);
nor NOR4 (N11276, N11275, N2285, N4280, N8839);
buf BUF1 (N11277, N11256);
xor XOR2 (N11278, N11267, N9359);
nand NAND4 (N11279, N11272, N389, N4398, N2324);
or OR4 (N11280, N11273, N9691, N698, N7009);
or OR2 (N11281, N11280, N1876);
nor NOR3 (N11282, N11261, N2902, N8780);
nand NAND2 (N11283, N11270, N8536);
not NOT1 (N11284, N11241);
and AND3 (N11285, N11268, N6589, N147);
xor XOR2 (N11286, N11274, N2456);
nor NOR2 (N11287, N11279, N416);
buf BUF1 (N11288, N11281);
nor NOR3 (N11289, N11286, N4899, N10775);
nand NAND3 (N11290, N11277, N8755, N9927);
and AND3 (N11291, N11283, N6098, N5527);
buf BUF1 (N11292, N11278);
nor NOR3 (N11293, N11292, N3400, N9234);
xor XOR2 (N11294, N11287, N1348);
nor NOR4 (N11295, N11288, N7469, N6513, N3962);
and AND2 (N11296, N11289, N3774);
xor XOR2 (N11297, N11284, N4917);
or OR2 (N11298, N11290, N8026);
and AND2 (N11299, N11295, N9383);
buf BUF1 (N11300, N11297);
xor XOR2 (N11301, N11298, N851);
and AND2 (N11302, N11300, N5875);
buf BUF1 (N11303, N11301);
not NOT1 (N11304, N11299);
nand NAND4 (N11305, N11304, N10091, N4844, N9371);
not NOT1 (N11306, N11302);
xor XOR2 (N11307, N11276, N9670);
or OR4 (N11308, N11305, N430, N10583, N10158);
not NOT1 (N11309, N11307);
nand NAND4 (N11310, N11282, N6670, N8168, N972);
xor XOR2 (N11311, N11309, N5129);
or OR4 (N11312, N11294, N4806, N1443, N3105);
or OR4 (N11313, N11311, N6889, N1900, N9047);
not NOT1 (N11314, N11296);
nor NOR2 (N11315, N11285, N10643);
not NOT1 (N11316, N11313);
buf BUF1 (N11317, N11303);
and AND2 (N11318, N11314, N4666);
nor NOR2 (N11319, N11291, N7221);
xor XOR2 (N11320, N11317, N8501);
buf BUF1 (N11321, N11315);
or OR2 (N11322, N11316, N1776);
xor XOR2 (N11323, N11312, N11054);
nand NAND3 (N11324, N11319, N5469, N7472);
not NOT1 (N11325, N11306);
not NOT1 (N11326, N11325);
xor XOR2 (N11327, N11318, N711);
nand NAND4 (N11328, N11321, N484, N5751, N3806);
xor XOR2 (N11329, N11320, N1120);
nand NAND4 (N11330, N11322, N2072, N8679, N9732);
or OR2 (N11331, N11329, N9791);
nand NAND2 (N11332, N11310, N2963);
nor NOR2 (N11333, N11323, N89);
nor NOR2 (N11334, N11330, N5760);
buf BUF1 (N11335, N11331);
and AND4 (N11336, N11308, N6453, N4180, N10026);
not NOT1 (N11337, N11336);
not NOT1 (N11338, N11334);
nor NOR4 (N11339, N11333, N3712, N11046, N2954);
or OR2 (N11340, N11328, N3169);
xor XOR2 (N11341, N11327, N6414);
buf BUF1 (N11342, N11337);
or OR2 (N11343, N11340, N2303);
or OR2 (N11344, N11335, N8245);
nor NOR2 (N11345, N11324, N1061);
or OR4 (N11346, N11344, N829, N4910, N4122);
and AND3 (N11347, N11332, N8898, N123);
or OR2 (N11348, N11343, N5086);
nand NAND3 (N11349, N11341, N8769, N9169);
or OR4 (N11350, N11339, N6300, N4076, N3797);
nor NOR3 (N11351, N11342, N6104, N6041);
buf BUF1 (N11352, N11349);
or OR4 (N11353, N11338, N607, N8112, N1104);
not NOT1 (N11354, N11353);
and AND2 (N11355, N11346, N7215);
and AND3 (N11356, N11354, N5987, N878);
or OR2 (N11357, N11355, N6268);
or OR2 (N11358, N11293, N9090);
or OR4 (N11359, N11358, N5315, N1373, N1427);
nand NAND4 (N11360, N11359, N4717, N4608, N2275);
nor NOR2 (N11361, N11351, N9289);
xor XOR2 (N11362, N11326, N6184);
buf BUF1 (N11363, N11352);
xor XOR2 (N11364, N11350, N5792);
xor XOR2 (N11365, N11362, N730);
xor XOR2 (N11366, N11364, N6488);
and AND2 (N11367, N11347, N7556);
not NOT1 (N11368, N11356);
or OR2 (N11369, N11345, N4533);
buf BUF1 (N11370, N11369);
and AND3 (N11371, N11361, N3607, N6715);
and AND3 (N11372, N11365, N3832, N1854);
nand NAND3 (N11373, N11363, N3226, N35);
nand NAND3 (N11374, N11373, N9732, N10487);
or OR4 (N11375, N11371, N7483, N6570, N4507);
nor NOR3 (N11376, N11372, N4311, N7941);
nand NAND3 (N11377, N11366, N10501, N8938);
nand NAND3 (N11378, N11376, N11276, N7052);
nor NOR3 (N11379, N11367, N1370, N2209);
nor NOR2 (N11380, N11377, N502);
not NOT1 (N11381, N11357);
nor NOR4 (N11382, N11379, N1165, N4058, N4551);
buf BUF1 (N11383, N11375);
xor XOR2 (N11384, N11381, N10958);
or OR2 (N11385, N11370, N4147);
xor XOR2 (N11386, N11385, N5702);
or OR2 (N11387, N11380, N6935);
and AND3 (N11388, N11348, N8716, N5674);
buf BUF1 (N11389, N11368);
nand NAND3 (N11390, N11382, N2449, N7001);
xor XOR2 (N11391, N11389, N4486);
buf BUF1 (N11392, N11386);
buf BUF1 (N11393, N11390);
nor NOR2 (N11394, N11378, N2520);
nand NAND3 (N11395, N11392, N287, N7012);
or OR4 (N11396, N11387, N9147, N731, N9745);
and AND2 (N11397, N11395, N339);
buf BUF1 (N11398, N11397);
and AND3 (N11399, N11360, N9278, N9579);
xor XOR2 (N11400, N11384, N9462);
buf BUF1 (N11401, N11396);
xor XOR2 (N11402, N11399, N1952);
and AND2 (N11403, N11398, N9984);
buf BUF1 (N11404, N11374);
xor XOR2 (N11405, N11391, N925);
nand NAND2 (N11406, N11400, N10498);
not NOT1 (N11407, N11388);
nand NAND4 (N11408, N11402, N2842, N382, N1548);
buf BUF1 (N11409, N11408);
buf BUF1 (N11410, N11404);
or OR4 (N11411, N11393, N8442, N11096, N223);
and AND2 (N11412, N11401, N11285);
buf BUF1 (N11413, N11412);
xor XOR2 (N11414, N11413, N462);
xor XOR2 (N11415, N11403, N5024);
not NOT1 (N11416, N11414);
nor NOR3 (N11417, N11383, N7843, N9527);
not NOT1 (N11418, N11415);
nor NOR3 (N11419, N11394, N5798, N4485);
nor NOR3 (N11420, N11410, N71, N5168);
not NOT1 (N11421, N11409);
nor NOR4 (N11422, N11421, N5808, N10347, N3504);
xor XOR2 (N11423, N11406, N7743);
or OR4 (N11424, N11423, N5978, N8986, N706);
nor NOR4 (N11425, N11420, N7730, N2025, N1126);
and AND3 (N11426, N11419, N9990, N2111);
nand NAND2 (N11427, N11416, N2233);
nand NAND3 (N11428, N11422, N2517, N9761);
or OR4 (N11429, N11424, N4932, N4368, N1454);
xor XOR2 (N11430, N11426, N10529);
not NOT1 (N11431, N11425);
buf BUF1 (N11432, N11417);
nand NAND2 (N11433, N11429, N6953);
not NOT1 (N11434, N11411);
nor NOR4 (N11435, N11431, N3572, N5747, N11303);
or OR3 (N11436, N11405, N1225, N2334);
nor NOR2 (N11437, N11433, N5832);
not NOT1 (N11438, N11430);
not NOT1 (N11439, N11427);
xor XOR2 (N11440, N11435, N5685);
buf BUF1 (N11441, N11432);
or OR4 (N11442, N11436, N9899, N7443, N2936);
xor XOR2 (N11443, N11441, N4846);
and AND4 (N11444, N11438, N112, N10221, N10109);
buf BUF1 (N11445, N11439);
or OR2 (N11446, N11418, N5256);
and AND3 (N11447, N11434, N6632, N5388);
nor NOR3 (N11448, N11445, N4648, N646);
or OR4 (N11449, N11428, N2209, N6083, N5024);
nor NOR3 (N11450, N11407, N7016, N3970);
nand NAND2 (N11451, N11449, N3390);
not NOT1 (N11452, N11448);
nor NOR2 (N11453, N11447, N8101);
nor NOR4 (N11454, N11451, N5148, N1254, N4140);
nor NOR2 (N11455, N11446, N6323);
nand NAND2 (N11456, N11454, N7104);
nand NAND3 (N11457, N11452, N2838, N545);
xor XOR2 (N11458, N11440, N10595);
nor NOR4 (N11459, N11437, N9261, N5120, N2358);
nor NOR4 (N11460, N11444, N8487, N538, N2344);
buf BUF1 (N11461, N11455);
and AND3 (N11462, N11458, N10777, N4919);
not NOT1 (N11463, N11457);
nor NOR4 (N11464, N11456, N10188, N3018, N10604);
nor NOR2 (N11465, N11462, N162);
not NOT1 (N11466, N11463);
and AND4 (N11467, N11442, N8514, N4581, N983);
nand NAND4 (N11468, N11459, N5340, N4667, N4269);
buf BUF1 (N11469, N11465);
and AND3 (N11470, N11453, N1729, N9510);
xor XOR2 (N11471, N11443, N5117);
xor XOR2 (N11472, N11468, N4552);
and AND4 (N11473, N11461, N1556, N9009, N10961);
nand NAND4 (N11474, N11467, N4614, N134, N10624);
xor XOR2 (N11475, N11471, N4364);
nor NOR3 (N11476, N11460, N393, N6516);
and AND4 (N11477, N11450, N11004, N7428, N10432);
buf BUF1 (N11478, N11470);
nor NOR3 (N11479, N11477, N1798, N4691);
nand NAND2 (N11480, N11473, N4547);
xor XOR2 (N11481, N11475, N10108);
or OR4 (N11482, N11464, N8605, N5527, N8312);
buf BUF1 (N11483, N11481);
buf BUF1 (N11484, N11478);
nand NAND3 (N11485, N11483, N9390, N805);
and AND3 (N11486, N11474, N1631, N356);
buf BUF1 (N11487, N11466);
or OR3 (N11488, N11480, N6000, N9673);
not NOT1 (N11489, N11487);
nor NOR3 (N11490, N11489, N1552, N770);
nand NAND4 (N11491, N11485, N11307, N6514, N8902);
xor XOR2 (N11492, N11482, N1075);
nor NOR2 (N11493, N11476, N3808);
xor XOR2 (N11494, N11488, N6906);
nand NAND4 (N11495, N11494, N7795, N2370, N8667);
and AND4 (N11496, N11486, N5151, N3054, N9534);
and AND3 (N11497, N11484, N8939, N8797);
xor XOR2 (N11498, N11469, N7586);
xor XOR2 (N11499, N11479, N2431);
nand NAND3 (N11500, N11498, N6091, N5555);
and AND3 (N11501, N11499, N1278, N6662);
or OR3 (N11502, N11492, N10426, N4392);
xor XOR2 (N11503, N11497, N8758);
buf BUF1 (N11504, N11495);
xor XOR2 (N11505, N11496, N1190);
nand NAND2 (N11506, N11472, N2847);
nor NOR2 (N11507, N11493, N2040);
buf BUF1 (N11508, N11500);
or OR2 (N11509, N11503, N10463);
nor NOR3 (N11510, N11491, N9659, N8608);
nand NAND2 (N11511, N11509, N2871);
nor NOR4 (N11512, N11490, N6425, N8277, N8548);
nor NOR2 (N11513, N11505, N6305);
xor XOR2 (N11514, N11504, N1890);
nor NOR4 (N11515, N11513, N7949, N28, N8594);
xor XOR2 (N11516, N11515, N8943);
nand NAND4 (N11517, N11507, N4880, N2608, N7431);
or OR4 (N11518, N11511, N2941, N4711, N714);
nand NAND3 (N11519, N11501, N10791, N10661);
and AND2 (N11520, N11518, N2650);
or OR2 (N11521, N11514, N3856);
buf BUF1 (N11522, N11502);
nand NAND2 (N11523, N11516, N5473);
buf BUF1 (N11524, N11519);
or OR3 (N11525, N11524, N9819, N8793);
nor NOR2 (N11526, N11508, N4774);
not NOT1 (N11527, N11526);
not NOT1 (N11528, N11521);
and AND4 (N11529, N11517, N4417, N9112, N11004);
or OR4 (N11530, N11528, N9409, N10170, N7473);
nand NAND4 (N11531, N11510, N7818, N8879, N5866);
buf BUF1 (N11532, N11527);
nand NAND3 (N11533, N11532, N7626, N8453);
not NOT1 (N11534, N11506);
xor XOR2 (N11535, N11533, N7565);
nand NAND3 (N11536, N11522, N5780, N4729);
and AND3 (N11537, N11534, N6028, N1714);
xor XOR2 (N11538, N11535, N235);
xor XOR2 (N11539, N11512, N8375);
not NOT1 (N11540, N11529);
or OR2 (N11541, N11539, N7265);
buf BUF1 (N11542, N11538);
nor NOR4 (N11543, N11541, N11108, N3272, N8330);
or OR4 (N11544, N11540, N846, N11521, N1626);
or OR3 (N11545, N11531, N10495, N9662);
xor XOR2 (N11546, N11545, N2607);
nor NOR2 (N11547, N11525, N1242);
nand NAND3 (N11548, N11542, N4973, N8671);
not NOT1 (N11549, N11546);
nand NAND3 (N11550, N11530, N6797, N11075);
nand NAND3 (N11551, N11549, N4794, N8924);
not NOT1 (N11552, N11536);
xor XOR2 (N11553, N11543, N1913);
and AND4 (N11554, N11552, N8980, N189, N11443);
not NOT1 (N11555, N11554);
not NOT1 (N11556, N11520);
buf BUF1 (N11557, N11544);
nor NOR3 (N11558, N11556, N366, N3255);
or OR4 (N11559, N11551, N393, N3068, N2736);
and AND4 (N11560, N11523, N4458, N11106, N8097);
not NOT1 (N11561, N11537);
buf BUF1 (N11562, N11550);
nand NAND4 (N11563, N11558, N5443, N7086, N5300);
buf BUF1 (N11564, N11561);
or OR2 (N11565, N11555, N2652);
buf BUF1 (N11566, N11565);
not NOT1 (N11567, N11560);
nand NAND4 (N11568, N11563, N6421, N7088, N861);
or OR2 (N11569, N11559, N3796);
and AND2 (N11570, N11568, N4934);
and AND4 (N11571, N11569, N1521, N10092, N3956);
nand NAND4 (N11572, N11564, N8830, N6725, N73);
or OR3 (N11573, N11562, N938, N8723);
or OR3 (N11574, N11571, N802, N7003);
xor XOR2 (N11575, N11566, N640);
or OR3 (N11576, N11553, N9094, N5797);
xor XOR2 (N11577, N11576, N618);
and AND4 (N11578, N11574, N2857, N2806, N9884);
nor NOR3 (N11579, N11578, N2966, N4293);
and AND3 (N11580, N11548, N11328, N9383);
or OR4 (N11581, N11547, N6932, N3397, N8121);
buf BUF1 (N11582, N11579);
nor NOR3 (N11583, N11580, N3951, N859);
nand NAND4 (N11584, N11572, N10352, N8475, N8325);
not NOT1 (N11585, N11570);
not NOT1 (N11586, N11585);
nor NOR3 (N11587, N11583, N717, N4621);
buf BUF1 (N11588, N11575);
not NOT1 (N11589, N11557);
not NOT1 (N11590, N11573);
xor XOR2 (N11591, N11577, N5499);
or OR2 (N11592, N11581, N1323);
and AND2 (N11593, N11591, N8645);
and AND4 (N11594, N11589, N2303, N2283, N266);
not NOT1 (N11595, N11582);
nor NOR3 (N11596, N11595, N7927, N3462);
nand NAND3 (N11597, N11596, N7819, N9821);
nor NOR3 (N11598, N11586, N8756, N6056);
not NOT1 (N11599, N11594);
xor XOR2 (N11600, N11593, N8368);
not NOT1 (N11601, N11598);
and AND4 (N11602, N11590, N8249, N6313, N3237);
buf BUF1 (N11603, N11584);
or OR4 (N11604, N11600, N178, N3369, N9075);
xor XOR2 (N11605, N11588, N401);
buf BUF1 (N11606, N11599);
and AND4 (N11607, N11604, N9199, N8087, N9932);
or OR3 (N11608, N11597, N6404, N11277);
xor XOR2 (N11609, N11587, N4860);
and AND4 (N11610, N11592, N3240, N9324, N4523);
not NOT1 (N11611, N11601);
nor NOR4 (N11612, N11567, N1212, N5278, N9655);
nand NAND3 (N11613, N11603, N1587, N5230);
nand NAND4 (N11614, N11613, N3516, N4641, N1406);
and AND2 (N11615, N11606, N457);
and AND3 (N11616, N11612, N8141, N6774);
xor XOR2 (N11617, N11610, N3436);
buf BUF1 (N11618, N11607);
and AND4 (N11619, N11611, N3449, N8214, N8299);
xor XOR2 (N11620, N11617, N5866);
nor NOR4 (N11621, N11605, N1041, N5463, N7051);
and AND2 (N11622, N11618, N1543);
buf BUF1 (N11623, N11619);
nand NAND3 (N11624, N11608, N10823, N2960);
xor XOR2 (N11625, N11615, N1525);
nor NOR4 (N11626, N11621, N9652, N9031, N2822);
nor NOR4 (N11627, N11602, N2470, N2062, N227);
xor XOR2 (N11628, N11616, N1102);
not NOT1 (N11629, N11624);
xor XOR2 (N11630, N11629, N7002);
xor XOR2 (N11631, N11614, N781);
or OR4 (N11632, N11609, N722, N11050, N5073);
or OR4 (N11633, N11626, N5503, N3362, N3474);
buf BUF1 (N11634, N11628);
xor XOR2 (N11635, N11632, N7602);
and AND2 (N11636, N11627, N4954);
and AND2 (N11637, N11625, N6607);
nand NAND3 (N11638, N11637, N8494, N3379);
or OR3 (N11639, N11635, N9309, N694);
xor XOR2 (N11640, N11639, N9280);
nand NAND4 (N11641, N11623, N900, N8291, N6348);
not NOT1 (N11642, N11634);
and AND2 (N11643, N11641, N9145);
and AND4 (N11644, N11633, N396, N5384, N5460);
or OR4 (N11645, N11642, N6962, N2506, N8428);
xor XOR2 (N11646, N11622, N8043);
buf BUF1 (N11647, N11631);
xor XOR2 (N11648, N11646, N5212);
nand NAND2 (N11649, N11643, N3097);
and AND3 (N11650, N11640, N9002, N22);
buf BUF1 (N11651, N11647);
xor XOR2 (N11652, N11649, N2639);
or OR4 (N11653, N11644, N7964, N5338, N8232);
xor XOR2 (N11654, N11653, N10324);
or OR3 (N11655, N11630, N8280, N4040);
nand NAND2 (N11656, N11638, N5703);
not NOT1 (N11657, N11655);
buf BUF1 (N11658, N11652);
or OR3 (N11659, N11657, N7584, N851);
and AND3 (N11660, N11654, N4014, N9114);
and AND2 (N11661, N11648, N4875);
not NOT1 (N11662, N11636);
xor XOR2 (N11663, N11661, N581);
nor NOR4 (N11664, N11620, N1788, N6894, N1806);
and AND4 (N11665, N11651, N10860, N6019, N912);
not NOT1 (N11666, N11664);
nor NOR2 (N11667, N11650, N11138);
xor XOR2 (N11668, N11666, N6819);
not NOT1 (N11669, N11663);
nand NAND2 (N11670, N11645, N9285);
not NOT1 (N11671, N11670);
or OR4 (N11672, N11656, N8364, N10399, N1275);
and AND4 (N11673, N11669, N771, N6707, N786);
not NOT1 (N11674, N11665);
nand NAND2 (N11675, N11667, N8758);
or OR3 (N11676, N11673, N2349, N1279);
and AND2 (N11677, N11658, N491);
nand NAND3 (N11678, N11659, N4710, N4933);
not NOT1 (N11679, N11662);
not NOT1 (N11680, N11674);
and AND3 (N11681, N11679, N2434, N6289);
and AND4 (N11682, N11681, N11036, N1419, N4673);
or OR2 (N11683, N11680, N5696);
or OR3 (N11684, N11660, N7903, N7221);
nor NOR3 (N11685, N11672, N1037, N516);
nor NOR2 (N11686, N11685, N886);
xor XOR2 (N11687, N11682, N3919);
and AND3 (N11688, N11676, N5029, N6406);
buf BUF1 (N11689, N11688);
not NOT1 (N11690, N11689);
nor NOR3 (N11691, N11686, N2617, N10458);
not NOT1 (N11692, N11677);
xor XOR2 (N11693, N11684, N4547);
buf BUF1 (N11694, N11671);
xor XOR2 (N11695, N11668, N1102);
nor NOR2 (N11696, N11693, N7463);
buf BUF1 (N11697, N11695);
buf BUF1 (N11698, N11697);
and AND3 (N11699, N11694, N2387, N5095);
xor XOR2 (N11700, N11675, N2576);
nand NAND3 (N11701, N11698, N577, N2005);
and AND4 (N11702, N11701, N4037, N5761, N1536);
nor NOR4 (N11703, N11700, N4568, N2981, N2988);
nor NOR4 (N11704, N11696, N330, N9716, N1984);
and AND4 (N11705, N11702, N3655, N1592, N1276);
or OR2 (N11706, N11691, N3308);
or OR4 (N11707, N11678, N245, N5548, N7004);
not NOT1 (N11708, N11707);
not NOT1 (N11709, N11690);
xor XOR2 (N11710, N11706, N3120);
nand NAND4 (N11711, N11683, N1774, N11411, N5904);
nor NOR2 (N11712, N11703, N8971);
or OR2 (N11713, N11709, N9574);
xor XOR2 (N11714, N11712, N10158);
nor NOR3 (N11715, N11687, N1435, N5113);
and AND3 (N11716, N11710, N10925, N8868);
not NOT1 (N11717, N11714);
buf BUF1 (N11718, N11704);
buf BUF1 (N11719, N11716);
nand NAND2 (N11720, N11715, N7186);
nand NAND3 (N11721, N11705, N10910, N3009);
or OR3 (N11722, N11692, N7436, N7295);
and AND3 (N11723, N11721, N182, N5316);
or OR4 (N11724, N11719, N4696, N708, N6258);
nor NOR3 (N11725, N11713, N244, N5295);
nand NAND4 (N11726, N11718, N7696, N4793, N874);
and AND2 (N11727, N11708, N11671);
nand NAND2 (N11728, N11717, N8608);
not NOT1 (N11729, N11727);
nand NAND4 (N11730, N11723, N10972, N6184, N2494);
nor NOR3 (N11731, N11699, N348, N4239);
nor NOR3 (N11732, N11725, N9586, N4813);
or OR3 (N11733, N11728, N4263, N9360);
nor NOR3 (N11734, N11724, N4342, N10220);
nor NOR4 (N11735, N11731, N11569, N5424, N3775);
buf BUF1 (N11736, N11711);
nor NOR4 (N11737, N11736, N9064, N2727, N2654);
not NOT1 (N11738, N11722);
not NOT1 (N11739, N11730);
not NOT1 (N11740, N11729);
not NOT1 (N11741, N11733);
not NOT1 (N11742, N11720);
nand NAND4 (N11743, N11741, N869, N10818, N1482);
and AND3 (N11744, N11739, N4479, N2093);
buf BUF1 (N11745, N11742);
nor NOR4 (N11746, N11745, N8449, N3881, N2250);
nor NOR2 (N11747, N11726, N9596);
nand NAND4 (N11748, N11734, N9815, N6042, N1362);
xor XOR2 (N11749, N11746, N6167);
nand NAND2 (N11750, N11732, N9135);
buf BUF1 (N11751, N11744);
nand NAND3 (N11752, N11751, N7919, N3078);
or OR4 (N11753, N11738, N1275, N3601, N9945);
or OR2 (N11754, N11740, N3020);
buf BUF1 (N11755, N11752);
nor NOR3 (N11756, N11735, N7360, N4450);
not NOT1 (N11757, N11755);
buf BUF1 (N11758, N11747);
xor XOR2 (N11759, N11758, N1490);
nor NOR2 (N11760, N11737, N7740);
and AND4 (N11761, N11748, N6989, N4399, N9519);
or OR4 (N11762, N11743, N4169, N10190, N4061);
nor NOR4 (N11763, N11757, N11309, N3954, N4105);
or OR4 (N11764, N11760, N4883, N9274, N3108);
not NOT1 (N11765, N11762);
not NOT1 (N11766, N11765);
xor XOR2 (N11767, N11753, N5557);
buf BUF1 (N11768, N11754);
or OR3 (N11769, N11756, N10557, N7748);
xor XOR2 (N11770, N11766, N8084);
not NOT1 (N11771, N11749);
nand NAND4 (N11772, N11759, N7785, N1390, N7833);
buf BUF1 (N11773, N11750);
and AND3 (N11774, N11772, N4984, N2947);
xor XOR2 (N11775, N11767, N3679);
xor XOR2 (N11776, N11775, N3848);
nand NAND4 (N11777, N11774, N2511, N3722, N7600);
and AND3 (N11778, N11776, N593, N4617);
xor XOR2 (N11779, N11770, N5589);
nand NAND2 (N11780, N11771, N11221);
buf BUF1 (N11781, N11780);
buf BUF1 (N11782, N11773);
not NOT1 (N11783, N11768);
not NOT1 (N11784, N11761);
or OR3 (N11785, N11778, N9755, N11703);
nand NAND4 (N11786, N11781, N962, N10287, N5521);
nor NOR2 (N11787, N11784, N2344);
or OR2 (N11788, N11783, N5133);
not NOT1 (N11789, N11764);
xor XOR2 (N11790, N11769, N30);
buf BUF1 (N11791, N11782);
or OR4 (N11792, N11787, N9524, N6444, N7789);
xor XOR2 (N11793, N11785, N4416);
not NOT1 (N11794, N11779);
not NOT1 (N11795, N11789);
not NOT1 (N11796, N11791);
not NOT1 (N11797, N11777);
or OR2 (N11798, N11794, N4639);
buf BUF1 (N11799, N11795);
or OR4 (N11800, N11799, N2822, N2791, N7763);
nand NAND2 (N11801, N11796, N5119);
and AND4 (N11802, N11788, N10063, N11375, N11244);
nand NAND2 (N11803, N11763, N9679);
xor XOR2 (N11804, N11801, N8784);
xor XOR2 (N11805, N11803, N7205);
buf BUF1 (N11806, N11800);
nor NOR2 (N11807, N11786, N202);
nor NOR4 (N11808, N11805, N11738, N5692, N4340);
or OR3 (N11809, N11806, N11447, N561);
and AND3 (N11810, N11798, N5837, N6216);
nand NAND3 (N11811, N11809, N8746, N724);
buf BUF1 (N11812, N11792);
and AND4 (N11813, N11793, N3639, N158, N2975);
or OR4 (N11814, N11804, N8390, N9456, N9015);
not NOT1 (N11815, N11813);
or OR2 (N11816, N11808, N10183);
nor NOR2 (N11817, N11802, N7254);
xor XOR2 (N11818, N11812, N7691);
nand NAND3 (N11819, N11797, N1387, N11363);
xor XOR2 (N11820, N11811, N1021);
and AND4 (N11821, N11817, N538, N1214, N9145);
nand NAND2 (N11822, N11821, N9741);
or OR2 (N11823, N11814, N136);
buf BUF1 (N11824, N11816);
nor NOR4 (N11825, N11818, N2476, N9937, N10005);
or OR2 (N11826, N11820, N4452);
not NOT1 (N11827, N11815);
buf BUF1 (N11828, N11827);
and AND4 (N11829, N11824, N8078, N11358, N4198);
buf BUF1 (N11830, N11810);
buf BUF1 (N11831, N11830);
or OR2 (N11832, N11825, N10452);
nor NOR2 (N11833, N11790, N10727);
xor XOR2 (N11834, N11826, N3170);
and AND3 (N11835, N11822, N8066, N5223);
xor XOR2 (N11836, N11832, N4548);
and AND4 (N11837, N11807, N10875, N10777, N4240);
or OR3 (N11838, N11831, N5050, N7610);
not NOT1 (N11839, N11834);
xor XOR2 (N11840, N11819, N10641);
buf BUF1 (N11841, N11823);
or OR2 (N11842, N11835, N2455);
nor NOR2 (N11843, N11836, N5403);
nor NOR3 (N11844, N11842, N555, N10629);
or OR2 (N11845, N11840, N9101);
not NOT1 (N11846, N11829);
buf BUF1 (N11847, N11837);
buf BUF1 (N11848, N11839);
and AND4 (N11849, N11841, N11563, N3162, N11543);
xor XOR2 (N11850, N11848, N5653);
nor NOR4 (N11851, N11849, N8210, N2133, N8041);
not NOT1 (N11852, N11844);
nor NOR2 (N11853, N11846, N3544);
or OR3 (N11854, N11852, N3771, N610);
xor XOR2 (N11855, N11853, N1642);
not NOT1 (N11856, N11833);
or OR4 (N11857, N11845, N9073, N10280, N530);
buf BUF1 (N11858, N11855);
or OR4 (N11859, N11854, N8090, N8170, N3543);
and AND2 (N11860, N11843, N6397);
or OR2 (N11861, N11847, N423);
and AND4 (N11862, N11851, N4651, N6731, N6358);
and AND4 (N11863, N11860, N4638, N1805, N8752);
not NOT1 (N11864, N11858);
nor NOR4 (N11865, N11828, N78, N5051, N5885);
xor XOR2 (N11866, N11861, N2105);
xor XOR2 (N11867, N11850, N2276);
xor XOR2 (N11868, N11859, N9049);
and AND3 (N11869, N11838, N9826, N4338);
and AND4 (N11870, N11863, N2088, N7798, N2042);
or OR2 (N11871, N11868, N5671);
xor XOR2 (N11872, N11869, N430);
nor NOR2 (N11873, N11870, N3632);
nand NAND3 (N11874, N11866, N10296, N10916);
nor NOR3 (N11875, N11856, N847, N9476);
not NOT1 (N11876, N11872);
nor NOR3 (N11877, N11873, N2437, N1114);
nor NOR4 (N11878, N11862, N1099, N2048, N6701);
buf BUF1 (N11879, N11875);
or OR2 (N11880, N11877, N1672);
nand NAND2 (N11881, N11878, N5323);
and AND3 (N11882, N11857, N852, N4583);
and AND3 (N11883, N11879, N4207, N11669);
xor XOR2 (N11884, N11867, N10166);
and AND4 (N11885, N11874, N4849, N255, N819);
not NOT1 (N11886, N11881);
nand NAND3 (N11887, N11883, N5822, N5275);
buf BUF1 (N11888, N11882);
nand NAND2 (N11889, N11864, N9335);
xor XOR2 (N11890, N11865, N428);
not NOT1 (N11891, N11884);
nor NOR2 (N11892, N11888, N3974);
nand NAND3 (N11893, N11876, N1527, N8121);
buf BUF1 (N11894, N11893);
nor NOR2 (N11895, N11871, N7815);
buf BUF1 (N11896, N11885);
xor XOR2 (N11897, N11891, N3058);
nand NAND4 (N11898, N11890, N201, N5652, N7963);
not NOT1 (N11899, N11880);
nand NAND4 (N11900, N11896, N631, N10667, N10166);
and AND2 (N11901, N11900, N9013);
nand NAND4 (N11902, N11899, N5028, N3503, N877);
or OR3 (N11903, N11898, N4513, N10940);
not NOT1 (N11904, N11902);
xor XOR2 (N11905, N11904, N3596);
nand NAND3 (N11906, N11895, N7911, N723);
not NOT1 (N11907, N11906);
buf BUF1 (N11908, N11897);
nand NAND3 (N11909, N11889, N259, N3578);
not NOT1 (N11910, N11903);
or OR3 (N11911, N11892, N2652, N8645);
nand NAND2 (N11912, N11909, N7994);
and AND3 (N11913, N11905, N3779, N1377);
not NOT1 (N11914, N11886);
buf BUF1 (N11915, N11901);
nand NAND3 (N11916, N11907, N11063, N232);
or OR4 (N11917, N11911, N2651, N7938, N4842);
not NOT1 (N11918, N11916);
nand NAND4 (N11919, N11912, N8914, N1277, N7141);
and AND4 (N11920, N11918, N8785, N7317, N6575);
nand NAND4 (N11921, N11920, N10074, N2285, N4331);
or OR2 (N11922, N11921, N3285);
nand NAND2 (N11923, N11887, N8908);
nor NOR2 (N11924, N11908, N4390);
and AND4 (N11925, N11917, N11701, N770, N3124);
or OR4 (N11926, N11915, N11779, N4398, N2054);
and AND3 (N11927, N11923, N11590, N6637);
xor XOR2 (N11928, N11894, N6085);
xor XOR2 (N11929, N11924, N8155);
xor XOR2 (N11930, N11919, N5817);
and AND3 (N11931, N11922, N901, N10370);
xor XOR2 (N11932, N11930, N1883);
nor NOR4 (N11933, N11927, N492, N2146, N6156);
not NOT1 (N11934, N11910);
not NOT1 (N11935, N11928);
or OR4 (N11936, N11934, N4960, N2836, N902);
nor NOR4 (N11937, N11914, N7011, N1817, N9106);
nand NAND4 (N11938, N11925, N9727, N1191, N119);
or OR3 (N11939, N11937, N9445, N10131);
nor NOR3 (N11940, N11931, N3313, N1138);
nand NAND3 (N11941, N11913, N654, N2315);
nand NAND3 (N11942, N11941, N1151, N9173);
and AND2 (N11943, N11939, N10881);
nor NOR3 (N11944, N11933, N10295, N7028);
nor NOR4 (N11945, N11936, N6719, N8187, N9977);
and AND2 (N11946, N11932, N403);
or OR2 (N11947, N11945, N8563);
or OR3 (N11948, N11942, N8116, N5339);
nand NAND4 (N11949, N11926, N2455, N5451, N9791);
nor NOR3 (N11950, N11943, N5959, N8716);
nand NAND2 (N11951, N11948, N11068);
xor XOR2 (N11952, N11950, N7921);
nor NOR2 (N11953, N11935, N11320);
nor NOR3 (N11954, N11940, N1422, N10723);
or OR3 (N11955, N11954, N9232, N4208);
nor NOR3 (N11956, N11951, N11153, N6118);
buf BUF1 (N11957, N11953);
or OR2 (N11958, N11946, N3072);
buf BUF1 (N11959, N11938);
and AND4 (N11960, N11929, N8480, N10460, N9090);
or OR2 (N11961, N11958, N8119);
xor XOR2 (N11962, N11944, N2485);
or OR2 (N11963, N11949, N7543);
nor NOR3 (N11964, N11962, N1207, N1153);
buf BUF1 (N11965, N11959);
and AND2 (N11966, N11965, N2396);
and AND3 (N11967, N11961, N11685, N4636);
nand NAND3 (N11968, N11947, N9081, N3912);
nor NOR3 (N11969, N11968, N11372, N5990);
nand NAND3 (N11970, N11967, N5593, N7115);
xor XOR2 (N11971, N11955, N10475);
and AND3 (N11972, N11960, N2611, N8885);
and AND3 (N11973, N11956, N7750, N10306);
or OR2 (N11974, N11969, N1602);
not NOT1 (N11975, N11966);
nand NAND2 (N11976, N11971, N1250);
xor XOR2 (N11977, N11957, N3206);
or OR4 (N11978, N11964, N8163, N1248, N8791);
buf BUF1 (N11979, N11978);
nor NOR4 (N11980, N11975, N10442, N6018, N9427);
and AND2 (N11981, N11963, N11616);
nor NOR3 (N11982, N11979, N264, N3611);
nand NAND4 (N11983, N11980, N4122, N824, N8248);
and AND2 (N11984, N11972, N8156);
nand NAND2 (N11985, N11970, N7203);
buf BUF1 (N11986, N11982);
buf BUF1 (N11987, N11977);
or OR2 (N11988, N11983, N2721);
buf BUF1 (N11989, N11986);
or OR3 (N11990, N11985, N1816, N4147);
not NOT1 (N11991, N11987);
and AND3 (N11992, N11991, N9579, N11782);
nor NOR3 (N11993, N11976, N5287, N7927);
not NOT1 (N11994, N11990);
not NOT1 (N11995, N11981);
nor NOR2 (N11996, N11995, N3265);
or OR2 (N11997, N11992, N5756);
nand NAND2 (N11998, N11993, N10451);
nand NAND2 (N11999, N11984, N8041);
or OR2 (N12000, N11996, N8106);
nor NOR3 (N12001, N12000, N11489, N8097);
nor NOR2 (N12002, N11989, N117);
and AND2 (N12003, N11988, N6864);
xor XOR2 (N12004, N11998, N2186);
and AND2 (N12005, N11973, N431);
or OR4 (N12006, N11994, N3950, N8390, N5777);
buf BUF1 (N12007, N12002);
and AND2 (N12008, N12001, N490);
xor XOR2 (N12009, N11997, N7071);
nor NOR4 (N12010, N12006, N2698, N2670, N1379);
and AND3 (N12011, N11952, N6309, N6177);
and AND3 (N12012, N12003, N756, N9099);
and AND2 (N12013, N11974, N11886);
buf BUF1 (N12014, N12012);
or OR4 (N12015, N12008, N7691, N8153, N11121);
not NOT1 (N12016, N11999);
and AND3 (N12017, N12005, N2378, N5709);
xor XOR2 (N12018, N12017, N3679);
buf BUF1 (N12019, N12009);
or OR3 (N12020, N12014, N3455, N1556);
not NOT1 (N12021, N12020);
nor NOR3 (N12022, N12007, N11958, N6353);
or OR3 (N12023, N12018, N7218, N936);
buf BUF1 (N12024, N12022);
buf BUF1 (N12025, N12015);
nand NAND3 (N12026, N12023, N2604, N11962);
or OR2 (N12027, N12019, N5401);
not NOT1 (N12028, N12013);
nor NOR4 (N12029, N12026, N11934, N7775, N266);
not NOT1 (N12030, N12010);
buf BUF1 (N12031, N12030);
nor NOR3 (N12032, N12004, N3800, N1787);
buf BUF1 (N12033, N12028);
buf BUF1 (N12034, N12011);
not NOT1 (N12035, N12027);
buf BUF1 (N12036, N12021);
not NOT1 (N12037, N12016);
xor XOR2 (N12038, N12034, N7418);
or OR2 (N12039, N12024, N1974);
and AND4 (N12040, N12032, N1449, N9343, N11127);
nor NOR2 (N12041, N12035, N3354);
nand NAND4 (N12042, N12038, N10999, N45, N2206);
buf BUF1 (N12043, N12025);
nand NAND3 (N12044, N12037, N10015, N10648);
buf BUF1 (N12045, N12041);
nand NAND2 (N12046, N12029, N1232);
nor NOR3 (N12047, N12039, N7911, N10456);
or OR4 (N12048, N12042, N5369, N10464, N8728);
not NOT1 (N12049, N12033);
nand NAND3 (N12050, N12040, N8161, N9805);
buf BUF1 (N12051, N12043);
or OR3 (N12052, N12047, N11678, N2283);
or OR4 (N12053, N12045, N10235, N8419, N113);
nor NOR2 (N12054, N12052, N10944);
and AND4 (N12055, N12046, N5053, N9134, N9974);
or OR3 (N12056, N12054, N951, N4173);
nand NAND4 (N12057, N12049, N9937, N2911, N2595);
nor NOR2 (N12058, N12053, N504);
buf BUF1 (N12059, N12050);
buf BUF1 (N12060, N12057);
or OR3 (N12061, N12036, N10325, N837);
or OR2 (N12062, N12060, N4005);
nand NAND4 (N12063, N12051, N678, N3843, N10025);
and AND2 (N12064, N12062, N8496);
buf BUF1 (N12065, N12048);
not NOT1 (N12066, N12059);
or OR4 (N12067, N12031, N3785, N6105, N455);
and AND4 (N12068, N12063, N2619, N86, N7807);
and AND2 (N12069, N12061, N3775);
buf BUF1 (N12070, N12068);
not NOT1 (N12071, N12056);
not NOT1 (N12072, N12071);
not NOT1 (N12073, N12070);
not NOT1 (N12074, N12066);
nor NOR3 (N12075, N12067, N777, N3884);
nor NOR3 (N12076, N12073, N3189, N3798);
xor XOR2 (N12077, N12075, N1251);
nand NAND2 (N12078, N12055, N5325);
or OR4 (N12079, N12065, N9295, N9249, N10171);
buf BUF1 (N12080, N12069);
nor NOR3 (N12081, N12079, N6588, N3896);
nor NOR4 (N12082, N12078, N3528, N6606, N8808);
xor XOR2 (N12083, N12072, N191);
nor NOR4 (N12084, N12077, N11767, N11245, N4405);
buf BUF1 (N12085, N12081);
xor XOR2 (N12086, N12082, N3008);
and AND2 (N12087, N12044, N6621);
buf BUF1 (N12088, N12083);
and AND3 (N12089, N12074, N4964, N4589);
not NOT1 (N12090, N12080);
and AND2 (N12091, N12076, N930);
not NOT1 (N12092, N12084);
nand NAND3 (N12093, N12085, N8569, N10138);
or OR3 (N12094, N12058, N3777, N4124);
and AND2 (N12095, N12086, N3370);
buf BUF1 (N12096, N12091);
nand NAND2 (N12097, N12092, N11197);
nor NOR3 (N12098, N12064, N4998, N3933);
nand NAND2 (N12099, N12098, N8242);
and AND4 (N12100, N12089, N10001, N3163, N5644);
and AND4 (N12101, N12097, N1061, N8248, N5227);
buf BUF1 (N12102, N12096);
nand NAND3 (N12103, N12100, N6385, N1547);
not NOT1 (N12104, N12099);
not NOT1 (N12105, N12090);
or OR3 (N12106, N12087, N8568, N7142);
or OR4 (N12107, N12105, N2572, N2799, N6978);
nor NOR3 (N12108, N12101, N3005, N6899);
or OR2 (N12109, N12088, N3060);
or OR2 (N12110, N12094, N6823);
nand NAND3 (N12111, N12102, N11195, N6435);
and AND4 (N12112, N12106, N9616, N5615, N2857);
not NOT1 (N12113, N12108);
not NOT1 (N12114, N12093);
and AND4 (N12115, N12107, N5266, N8452, N8908);
and AND2 (N12116, N12111, N857);
or OR2 (N12117, N12116, N10769);
nor NOR2 (N12118, N12112, N9474);
or OR3 (N12119, N12109, N12076, N815);
nand NAND3 (N12120, N12115, N2917, N405);
buf BUF1 (N12121, N12117);
and AND4 (N12122, N12118, N8145, N2422, N8050);
nand NAND2 (N12123, N12113, N7283);
xor XOR2 (N12124, N12123, N3269);
xor XOR2 (N12125, N12121, N6465);
xor XOR2 (N12126, N12104, N5713);
and AND3 (N12127, N12120, N9578, N10338);
and AND4 (N12128, N12103, N6865, N9060, N5695);
buf BUF1 (N12129, N12114);
and AND4 (N12130, N12125, N9244, N4144, N9321);
xor XOR2 (N12131, N12122, N2581);
and AND4 (N12132, N12128, N957, N4343, N4403);
and AND4 (N12133, N12126, N3972, N1075, N11457);
xor XOR2 (N12134, N12129, N10871);
buf BUF1 (N12135, N12127);
nand NAND2 (N12136, N12131, N10485);
nand NAND3 (N12137, N12124, N4355, N3632);
not NOT1 (N12138, N12137);
buf BUF1 (N12139, N12119);
or OR4 (N12140, N12139, N349, N8811, N2527);
and AND2 (N12141, N12133, N6633);
xor XOR2 (N12142, N12095, N7179);
and AND2 (N12143, N12132, N10285);
not NOT1 (N12144, N12143);
xor XOR2 (N12145, N12144, N3019);
not NOT1 (N12146, N12138);
not NOT1 (N12147, N12145);
nor NOR2 (N12148, N12141, N11378);
xor XOR2 (N12149, N12110, N3110);
and AND3 (N12150, N12140, N8949, N7602);
xor XOR2 (N12151, N12150, N4496);
buf BUF1 (N12152, N12135);
buf BUF1 (N12153, N12136);
not NOT1 (N12154, N12153);
buf BUF1 (N12155, N12146);
xor XOR2 (N12156, N12148, N9546);
nor NOR2 (N12157, N12151, N8623);
not NOT1 (N12158, N12154);
nor NOR2 (N12159, N12156, N6557);
not NOT1 (N12160, N12149);
or OR3 (N12161, N12147, N1101, N7452);
not NOT1 (N12162, N12134);
nor NOR4 (N12163, N12159, N4234, N8525, N8594);
or OR2 (N12164, N12162, N6946);
buf BUF1 (N12165, N12155);
nor NOR2 (N12166, N12142, N3092);
nor NOR3 (N12167, N12160, N9448, N7701);
not NOT1 (N12168, N12163);
xor XOR2 (N12169, N12164, N5623);
nor NOR3 (N12170, N12161, N6775, N1970);
nand NAND2 (N12171, N12130, N4840);
nor NOR3 (N12172, N12167, N1008, N2925);
and AND2 (N12173, N12152, N3358);
not NOT1 (N12174, N12173);
not NOT1 (N12175, N12166);
nor NOR3 (N12176, N12169, N7643, N11648);
or OR3 (N12177, N12172, N7179, N2799);
xor XOR2 (N12178, N12165, N8967);
buf BUF1 (N12179, N12168);
not NOT1 (N12180, N12170);
xor XOR2 (N12181, N12174, N3432);
nor NOR3 (N12182, N12158, N5656, N430);
nand NAND3 (N12183, N12176, N11700, N2613);
not NOT1 (N12184, N12171);
and AND4 (N12185, N12183, N9586, N6068, N2084);
nand NAND3 (N12186, N12184, N2304, N6805);
buf BUF1 (N12187, N12179);
or OR2 (N12188, N12186, N2324);
and AND2 (N12189, N12178, N7806);
xor XOR2 (N12190, N12177, N8827);
and AND3 (N12191, N12190, N7844, N8655);
and AND3 (N12192, N12187, N833, N1316);
nor NOR4 (N12193, N12180, N2946, N4810, N10760);
xor XOR2 (N12194, N12192, N348);
buf BUF1 (N12195, N12157);
buf BUF1 (N12196, N12195);
and AND4 (N12197, N12188, N6902, N7603, N5753);
or OR2 (N12198, N12194, N10968);
or OR2 (N12199, N12182, N104);
not NOT1 (N12200, N12181);
xor XOR2 (N12201, N12197, N8810);
nand NAND4 (N12202, N12201, N2742, N6539, N11648);
buf BUF1 (N12203, N12202);
or OR4 (N12204, N12199, N12166, N3067, N4735);
xor XOR2 (N12205, N12185, N1120);
and AND4 (N12206, N12204, N11585, N6912, N42);
nand NAND3 (N12207, N12206, N10926, N1384);
and AND4 (N12208, N12203, N962, N4361, N5403);
buf BUF1 (N12209, N12208);
xor XOR2 (N12210, N12175, N7545);
buf BUF1 (N12211, N12196);
nor NOR3 (N12212, N12189, N2443, N2811);
xor XOR2 (N12213, N12198, N10919);
xor XOR2 (N12214, N12213, N4896);
xor XOR2 (N12215, N12191, N5244);
xor XOR2 (N12216, N12200, N616);
nand NAND2 (N12217, N12209, N10209);
buf BUF1 (N12218, N12216);
xor XOR2 (N12219, N12211, N1025);
nor NOR4 (N12220, N12215, N5529, N8492, N6410);
or OR4 (N12221, N12210, N4034, N7515, N3428);
buf BUF1 (N12222, N12214);
buf BUF1 (N12223, N12220);
and AND2 (N12224, N12193, N9069);
nor NOR4 (N12225, N12222, N8850, N5225, N10451);
or OR4 (N12226, N12224, N1644, N12114, N6819);
and AND4 (N12227, N12221, N8554, N5574, N11402);
nand NAND3 (N12228, N12223, N5119, N3338);
buf BUF1 (N12229, N12228);
buf BUF1 (N12230, N12217);
and AND4 (N12231, N12230, N3671, N2563, N9903);
not NOT1 (N12232, N12207);
not NOT1 (N12233, N12232);
not NOT1 (N12234, N12225);
nor NOR4 (N12235, N12218, N11925, N908, N7953);
or OR2 (N12236, N12226, N4174);
xor XOR2 (N12237, N12212, N8594);
nor NOR4 (N12238, N12231, N6617, N11378, N10578);
buf BUF1 (N12239, N12205);
and AND3 (N12240, N12227, N7116, N2285);
and AND4 (N12241, N12236, N1697, N551, N9646);
xor XOR2 (N12242, N12240, N1419);
not NOT1 (N12243, N12234);
and AND4 (N12244, N12241, N2490, N11061, N2950);
or OR2 (N12245, N12219, N6495);
buf BUF1 (N12246, N12244);
xor XOR2 (N12247, N12243, N8839);
buf BUF1 (N12248, N12247);
buf BUF1 (N12249, N12246);
or OR4 (N12250, N12238, N7363, N4736, N10953);
not NOT1 (N12251, N12245);
nor NOR4 (N12252, N12239, N86, N1234, N7631);
nand NAND2 (N12253, N12252, N9663);
or OR2 (N12254, N12235, N11428);
buf BUF1 (N12255, N12249);
xor XOR2 (N12256, N12250, N3335);
or OR2 (N12257, N12251, N2035);
and AND3 (N12258, N12257, N3928, N11990);
nor NOR3 (N12259, N12253, N808, N3614);
nor NOR4 (N12260, N12258, N3905, N6647, N4347);
and AND3 (N12261, N12248, N7316, N2814);
or OR2 (N12262, N12237, N2871);
nor NOR2 (N12263, N12229, N10216);
or OR3 (N12264, N12255, N7673, N566);
nor NOR2 (N12265, N12233, N10976);
buf BUF1 (N12266, N12259);
and AND3 (N12267, N12242, N1342, N3758);
buf BUF1 (N12268, N12264);
not NOT1 (N12269, N12256);
xor XOR2 (N12270, N12269, N4655);
or OR2 (N12271, N12265, N485);
xor XOR2 (N12272, N12266, N1576);
nand NAND3 (N12273, N12263, N5949, N7570);
nor NOR2 (N12274, N12273, N9432);
xor XOR2 (N12275, N12274, N729);
buf BUF1 (N12276, N12268);
not NOT1 (N12277, N12270);
buf BUF1 (N12278, N12260);
xor XOR2 (N12279, N12278, N2004);
nand NAND3 (N12280, N12275, N7677, N894);
and AND3 (N12281, N12279, N2420, N8890);
not NOT1 (N12282, N12281);
not NOT1 (N12283, N12271);
or OR4 (N12284, N12267, N9978, N10120, N2393);
not NOT1 (N12285, N12277);
xor XOR2 (N12286, N12284, N3591);
buf BUF1 (N12287, N12272);
and AND4 (N12288, N12262, N3631, N11031, N2238);
buf BUF1 (N12289, N12287);
nor NOR3 (N12290, N12276, N4622, N7959);
nor NOR3 (N12291, N12254, N3489, N8936);
nand NAND3 (N12292, N12291, N6050, N11430);
or OR3 (N12293, N12283, N809, N12006);
not NOT1 (N12294, N12292);
and AND4 (N12295, N12285, N11461, N11701, N2248);
and AND4 (N12296, N12289, N6965, N642, N11988);
and AND2 (N12297, N12288, N2060);
nor NOR4 (N12298, N12296, N2754, N10317, N2493);
and AND2 (N12299, N12290, N10206);
nand NAND3 (N12300, N12299, N8796, N3943);
and AND2 (N12301, N12286, N5175);
xor XOR2 (N12302, N12294, N8196);
xor XOR2 (N12303, N12302, N1040);
nand NAND2 (N12304, N12298, N281);
and AND4 (N12305, N12261, N4630, N11521, N3740);
buf BUF1 (N12306, N12295);
xor XOR2 (N12307, N12300, N4191);
buf BUF1 (N12308, N12306);
or OR4 (N12309, N12305, N915, N3613, N9084);
buf BUF1 (N12310, N12280);
nor NOR4 (N12311, N12307, N3826, N7738, N5182);
nand NAND4 (N12312, N12310, N5213, N2651, N1644);
or OR3 (N12313, N12303, N11701, N2910);
nand NAND4 (N12314, N12301, N9661, N319, N10108);
buf BUF1 (N12315, N12297);
nor NOR2 (N12316, N12308, N7423);
and AND2 (N12317, N12315, N259);
buf BUF1 (N12318, N12282);
and AND2 (N12319, N12311, N2673);
or OR3 (N12320, N12314, N4586, N7466);
and AND4 (N12321, N12318, N7122, N6067, N7128);
nand NAND4 (N12322, N12313, N6548, N6129, N10075);
and AND3 (N12323, N12322, N4159, N10594);
or OR4 (N12324, N12317, N1916, N10634, N2384);
nand NAND3 (N12325, N12293, N4542, N2379);
nor NOR2 (N12326, N12325, N892);
not NOT1 (N12327, N12309);
buf BUF1 (N12328, N12319);
xor XOR2 (N12329, N12328, N27);
buf BUF1 (N12330, N12321);
or OR3 (N12331, N12329, N6229, N3188);
xor XOR2 (N12332, N12331, N1669);
buf BUF1 (N12333, N12323);
and AND4 (N12334, N12333, N3910, N3104, N11828);
and AND4 (N12335, N12320, N8845, N11350, N2851);
nor NOR3 (N12336, N12312, N10207, N960);
xor XOR2 (N12337, N12327, N9627);
and AND4 (N12338, N12334, N3983, N11277, N10566);
or OR4 (N12339, N12337, N9498, N52, N7783);
or OR2 (N12340, N12336, N944);
nor NOR4 (N12341, N12335, N5624, N11808, N1963);
or OR2 (N12342, N12339, N2058);
not NOT1 (N12343, N12338);
nor NOR3 (N12344, N12316, N9885, N2870);
buf BUF1 (N12345, N12340);
xor XOR2 (N12346, N12344, N4064);
and AND4 (N12347, N12341, N10291, N838, N1790);
nand NAND4 (N12348, N12346, N6816, N6901, N1802);
nor NOR4 (N12349, N12326, N8008, N7943, N7625);
nand NAND3 (N12350, N12348, N11778, N6626);
nor NOR3 (N12351, N12345, N12009, N7667);
nor NOR4 (N12352, N12304, N2152, N4508, N6719);
not NOT1 (N12353, N12332);
not NOT1 (N12354, N12342);
and AND3 (N12355, N12352, N7734, N1207);
nor NOR2 (N12356, N12347, N9617);
nand NAND2 (N12357, N12351, N6259);
xor XOR2 (N12358, N12343, N1693);
not NOT1 (N12359, N12353);
not NOT1 (N12360, N12359);
nand NAND4 (N12361, N12356, N5774, N461, N7959);
nand NAND3 (N12362, N12324, N11576, N544);
nor NOR3 (N12363, N12358, N12089, N10151);
and AND4 (N12364, N12360, N5077, N6847, N10499);
or OR4 (N12365, N12354, N1388, N6976, N7789);
or OR3 (N12366, N12364, N10093, N4856);
buf BUF1 (N12367, N12355);
nor NOR3 (N12368, N12366, N5656, N9034);
and AND2 (N12369, N12363, N8461);
and AND3 (N12370, N12350, N9087, N4841);
not NOT1 (N12371, N12349);
nand NAND4 (N12372, N12357, N10489, N2224, N7614);
or OR3 (N12373, N12371, N10182, N1760);
xor XOR2 (N12374, N12370, N3323);
nor NOR3 (N12375, N12369, N2207, N323);
xor XOR2 (N12376, N12367, N10622);
and AND2 (N12377, N12361, N504);
xor XOR2 (N12378, N12372, N5950);
nand NAND2 (N12379, N12373, N7042);
not NOT1 (N12380, N12330);
not NOT1 (N12381, N12374);
and AND3 (N12382, N12368, N8583, N3908);
and AND2 (N12383, N12378, N8446);
buf BUF1 (N12384, N12365);
buf BUF1 (N12385, N12381);
and AND3 (N12386, N12377, N1040, N5695);
and AND2 (N12387, N12375, N2484);
or OR2 (N12388, N12383, N10729);
nor NOR4 (N12389, N12362, N8448, N8873, N6952);
nand NAND4 (N12390, N12376, N7610, N7462, N1002);
xor XOR2 (N12391, N12382, N6136);
xor XOR2 (N12392, N12391, N4158);
not NOT1 (N12393, N12389);
nand NAND4 (N12394, N12385, N983, N5699, N7491);
nand NAND4 (N12395, N12386, N850, N10715, N5623);
xor XOR2 (N12396, N12387, N6966);
nor NOR4 (N12397, N12390, N11750, N11739, N2193);
xor XOR2 (N12398, N12392, N1589);
xor XOR2 (N12399, N12397, N10726);
nor NOR4 (N12400, N12384, N11194, N1469, N734);
not NOT1 (N12401, N12380);
buf BUF1 (N12402, N12388);
and AND3 (N12403, N12401, N5972, N10680);
or OR2 (N12404, N12398, N10795);
not NOT1 (N12405, N12404);
xor XOR2 (N12406, N12379, N6218);
or OR2 (N12407, N12400, N10891);
nor NOR3 (N12408, N12394, N1990, N8950);
and AND2 (N12409, N12405, N3660);
nor NOR4 (N12410, N12403, N1385, N5196, N2914);
nand NAND2 (N12411, N12395, N8369);
nor NOR3 (N12412, N12407, N5843, N11069);
buf BUF1 (N12413, N12396);
xor XOR2 (N12414, N12408, N5872);
xor XOR2 (N12415, N12413, N6816);
nor NOR4 (N12416, N12410, N6074, N6645, N6347);
or OR3 (N12417, N12402, N8859, N351);
and AND2 (N12418, N12406, N2870);
or OR2 (N12419, N12409, N6789);
nand NAND2 (N12420, N12393, N10501);
nor NOR3 (N12421, N12416, N4546, N575);
or OR2 (N12422, N12414, N12400);
xor XOR2 (N12423, N12419, N5458);
not NOT1 (N12424, N12411);
and AND2 (N12425, N12415, N8662);
nand NAND2 (N12426, N12425, N8904);
xor XOR2 (N12427, N12424, N2046);
xor XOR2 (N12428, N12427, N12259);
or OR2 (N12429, N12423, N10507);
xor XOR2 (N12430, N12422, N9073);
nor NOR2 (N12431, N12420, N1340);
xor XOR2 (N12432, N12430, N6035);
buf BUF1 (N12433, N12417);
and AND4 (N12434, N12428, N1529, N8252, N3818);
or OR4 (N12435, N12418, N10893, N1454, N3646);
nand NAND2 (N12436, N12432, N4180);
xor XOR2 (N12437, N12435, N6253);
not NOT1 (N12438, N12437);
buf BUF1 (N12439, N12399);
nand NAND2 (N12440, N12436, N11082);
nand NAND3 (N12441, N12434, N6953, N7210);
nor NOR3 (N12442, N12440, N8014, N4618);
buf BUF1 (N12443, N12433);
or OR4 (N12444, N12438, N5589, N2179, N2583);
and AND4 (N12445, N12443, N8806, N2106, N6389);
xor XOR2 (N12446, N12439, N11352);
not NOT1 (N12447, N12412);
nand NAND2 (N12448, N12441, N3217);
xor XOR2 (N12449, N12446, N9653);
buf BUF1 (N12450, N12447);
nand NAND3 (N12451, N12448, N4703, N4288);
not NOT1 (N12452, N12445);
nor NOR4 (N12453, N12450, N11536, N1849, N12137);
buf BUF1 (N12454, N12444);
xor XOR2 (N12455, N12429, N11075);
not NOT1 (N12456, N12452);
not NOT1 (N12457, N12453);
not NOT1 (N12458, N12451);
xor XOR2 (N12459, N12458, N11054);
or OR3 (N12460, N12421, N5919, N7089);
nand NAND4 (N12461, N12426, N11467, N3873, N10775);
buf BUF1 (N12462, N12459);
not NOT1 (N12463, N12462);
not NOT1 (N12464, N12457);
not NOT1 (N12465, N12460);
nor NOR2 (N12466, N12463, N131);
or OR2 (N12467, N12454, N5833);
or OR4 (N12468, N12442, N9791, N7898, N3907);
not NOT1 (N12469, N12468);
or OR2 (N12470, N12455, N7882);
not NOT1 (N12471, N12464);
and AND2 (N12472, N12470, N9277);
buf BUF1 (N12473, N12472);
nor NOR3 (N12474, N12465, N4871, N187);
nand NAND4 (N12475, N12471, N2306, N9811, N4877);
nor NOR3 (N12476, N12474, N10787, N4299);
or OR4 (N12477, N12473, N2186, N5887, N6130);
xor XOR2 (N12478, N12467, N7656);
or OR2 (N12479, N12469, N10693);
and AND2 (N12480, N12461, N3550);
xor XOR2 (N12481, N12466, N1642);
xor XOR2 (N12482, N12478, N8470);
or OR3 (N12483, N12456, N8499, N4429);
and AND4 (N12484, N12475, N4888, N4535, N10465);
buf BUF1 (N12485, N12484);
nor NOR4 (N12486, N12479, N3448, N8133, N984);
buf BUF1 (N12487, N12485);
nand NAND3 (N12488, N12477, N610, N10993);
buf BUF1 (N12489, N12481);
nand NAND2 (N12490, N12449, N93);
and AND4 (N12491, N12486, N10715, N7888, N9125);
xor XOR2 (N12492, N12491, N6548);
nor NOR2 (N12493, N12489, N779);
xor XOR2 (N12494, N12483, N495);
not NOT1 (N12495, N12493);
xor XOR2 (N12496, N12495, N6324);
or OR3 (N12497, N12494, N11332, N7102);
and AND2 (N12498, N12476, N10877);
nand NAND4 (N12499, N12492, N11373, N3384, N11194);
buf BUF1 (N12500, N12496);
nor NOR4 (N12501, N12488, N8812, N9993, N5476);
buf BUF1 (N12502, N12490);
and AND4 (N12503, N12502, N6521, N4747, N8411);
nand NAND2 (N12504, N12487, N827);
buf BUF1 (N12505, N12499);
nor NOR2 (N12506, N12497, N5278);
not NOT1 (N12507, N12504);
nor NOR3 (N12508, N12506, N6559, N5003);
buf BUF1 (N12509, N12500);
nor NOR4 (N12510, N12508, N8823, N864, N11375);
not NOT1 (N12511, N12503);
nor NOR4 (N12512, N12482, N8899, N858, N10068);
nor NOR3 (N12513, N12510, N7435, N590);
nand NAND2 (N12514, N12509, N3922);
nor NOR3 (N12515, N12513, N8820, N2412);
or OR2 (N12516, N12480, N3575);
nand NAND4 (N12517, N12498, N4506, N6383, N875);
nor NOR4 (N12518, N12501, N9647, N7659, N1818);
and AND3 (N12519, N12517, N8151, N3283);
nand NAND2 (N12520, N12515, N3266);
and AND3 (N12521, N12516, N1322, N11742);
and AND2 (N12522, N12505, N6323);
not NOT1 (N12523, N12519);
xor XOR2 (N12524, N12521, N10230);
not NOT1 (N12525, N12518);
nor NOR2 (N12526, N12507, N7427);
and AND4 (N12527, N12522, N7113, N933, N4210);
and AND2 (N12528, N12527, N2035);
or OR2 (N12529, N12524, N647);
nand NAND4 (N12530, N12511, N1898, N6929, N9233);
nor NOR3 (N12531, N12514, N6064, N3386);
and AND3 (N12532, N12431, N1020, N7010);
not NOT1 (N12533, N12526);
and AND2 (N12534, N12530, N5242);
or OR3 (N12535, N12529, N10101, N4590);
nand NAND3 (N12536, N12523, N4258, N2041);
or OR4 (N12537, N12533, N7664, N9164, N5780);
and AND4 (N12538, N12536, N11562, N2995, N7075);
nand NAND3 (N12539, N12537, N8046, N1199);
and AND2 (N12540, N12534, N6347);
nand NAND2 (N12541, N12539, N5721);
and AND2 (N12542, N12532, N4204);
or OR3 (N12543, N12531, N4194, N5992);
nand NAND4 (N12544, N12538, N1423, N4673, N5993);
and AND2 (N12545, N12544, N8675);
not NOT1 (N12546, N12540);
or OR4 (N12547, N12528, N9871, N6843, N11065);
buf BUF1 (N12548, N12547);
nand NAND3 (N12549, N12520, N10839, N7669);
or OR3 (N12550, N12549, N1422, N2439);
or OR4 (N12551, N12541, N5223, N4227, N5989);
and AND3 (N12552, N12512, N7317, N5505);
or OR4 (N12553, N12548, N6387, N3433, N6697);
or OR3 (N12554, N12543, N8195, N9645);
or OR3 (N12555, N12551, N2085, N571);
xor XOR2 (N12556, N12525, N573);
or OR4 (N12557, N12556, N2387, N11297, N8305);
nor NOR4 (N12558, N12535, N8624, N1669, N1344);
nor NOR4 (N12559, N12552, N11841, N9600, N2875);
not NOT1 (N12560, N12554);
not NOT1 (N12561, N12560);
or OR4 (N12562, N12546, N1341, N3042, N2857);
xor XOR2 (N12563, N12561, N850);
nand NAND3 (N12564, N12553, N11880, N476);
or OR3 (N12565, N12557, N3408, N10617);
nand NAND2 (N12566, N12564, N5259);
or OR2 (N12567, N12555, N1731);
nor NOR4 (N12568, N12566, N7533, N1285, N3134);
nor NOR4 (N12569, N12562, N11357, N10175, N7459);
xor XOR2 (N12570, N12565, N8518);
nor NOR4 (N12571, N12550, N9661, N1822, N4580);
nor NOR3 (N12572, N12571, N7953, N529);
nand NAND4 (N12573, N12558, N1933, N7334, N7842);
xor XOR2 (N12574, N12559, N10287);
nand NAND2 (N12575, N12545, N1327);
nor NOR3 (N12576, N12575, N6538, N12515);
nor NOR3 (N12577, N12569, N1560, N5843);
xor XOR2 (N12578, N12574, N522);
nor NOR2 (N12579, N12578, N602);
not NOT1 (N12580, N12563);
or OR2 (N12581, N12572, N5977);
nor NOR4 (N12582, N12580, N7893, N37, N5694);
nand NAND3 (N12583, N12542, N8258, N5931);
not NOT1 (N12584, N12577);
or OR4 (N12585, N12581, N6491, N11647, N5748);
nand NAND3 (N12586, N12583, N10731, N6155);
xor XOR2 (N12587, N12570, N2359);
or OR3 (N12588, N12576, N5658, N4356);
nor NOR4 (N12589, N12579, N12442, N10562, N6909);
or OR3 (N12590, N12584, N62, N8408);
nand NAND2 (N12591, N12568, N8146);
buf BUF1 (N12592, N12586);
buf BUF1 (N12593, N12587);
xor XOR2 (N12594, N12588, N11349);
xor XOR2 (N12595, N12591, N11477);
nand NAND2 (N12596, N12594, N9551);
or OR2 (N12597, N12592, N1442);
and AND2 (N12598, N12573, N8957);
or OR2 (N12599, N12597, N7694);
nor NOR4 (N12600, N12599, N1172, N778, N5405);
or OR2 (N12601, N12593, N7356);
and AND3 (N12602, N12582, N722, N4840);
buf BUF1 (N12603, N12567);
buf BUF1 (N12604, N12596);
buf BUF1 (N12605, N12602);
and AND4 (N12606, N12590, N7913, N11928, N6909);
and AND3 (N12607, N12605, N4741, N3954);
nand NAND3 (N12608, N12603, N11577, N3680);
buf BUF1 (N12609, N12608);
and AND4 (N12610, N12589, N2425, N12520, N8647);
nor NOR2 (N12611, N12606, N5611);
xor XOR2 (N12612, N12611, N8823);
and AND2 (N12613, N12601, N10313);
buf BUF1 (N12614, N12609);
and AND2 (N12615, N12598, N9529);
nand NAND3 (N12616, N12610, N4145, N1586);
nor NOR4 (N12617, N12616, N5315, N11427, N11510);
or OR4 (N12618, N12614, N8095, N9688, N3344);
nand NAND4 (N12619, N12595, N5098, N10693, N6547);
not NOT1 (N12620, N12612);
buf BUF1 (N12621, N12620);
not NOT1 (N12622, N12615);
nor NOR2 (N12623, N12585, N818);
not NOT1 (N12624, N12617);
buf BUF1 (N12625, N12624);
buf BUF1 (N12626, N12618);
nand NAND3 (N12627, N12607, N7233, N2497);
and AND3 (N12628, N12626, N3045, N7899);
or OR4 (N12629, N12613, N3843, N8601, N990);
or OR4 (N12630, N12621, N2778, N6424, N11331);
nor NOR4 (N12631, N12630, N10507, N7131, N5);
and AND4 (N12632, N12600, N10889, N516, N2372);
and AND3 (N12633, N12622, N9946, N715);
nand NAND4 (N12634, N12631, N2224, N4916, N4085);
or OR2 (N12635, N12633, N6750);
nand NAND3 (N12636, N12635, N10273, N12344);
buf BUF1 (N12637, N12619);
buf BUF1 (N12638, N12632);
nand NAND4 (N12639, N12623, N12549, N7754, N4142);
buf BUF1 (N12640, N12625);
not NOT1 (N12641, N12640);
buf BUF1 (N12642, N12637);
xor XOR2 (N12643, N12641, N9009);
and AND3 (N12644, N12629, N2273, N5185);
buf BUF1 (N12645, N12627);
or OR3 (N12646, N12645, N768, N8061);
or OR3 (N12647, N12604, N8432, N11843);
xor XOR2 (N12648, N12643, N6452);
and AND4 (N12649, N12628, N3523, N1517, N12399);
nor NOR4 (N12650, N12649, N9938, N4961, N12054);
xor XOR2 (N12651, N12634, N9821);
xor XOR2 (N12652, N12646, N7915);
not NOT1 (N12653, N12652);
nor NOR4 (N12654, N12650, N4286, N7061, N7870);
or OR2 (N12655, N12653, N578);
nor NOR2 (N12656, N12642, N4393);
not NOT1 (N12657, N12654);
nand NAND3 (N12658, N12638, N11499, N442);
buf BUF1 (N12659, N12655);
xor XOR2 (N12660, N12644, N8164);
nand NAND3 (N12661, N12636, N7431, N11947);
and AND4 (N12662, N12659, N6131, N8507, N3227);
xor XOR2 (N12663, N12658, N5467);
xor XOR2 (N12664, N12663, N9488);
nand NAND4 (N12665, N12660, N2995, N6717, N2088);
nand NAND4 (N12666, N12648, N9449, N5554, N2284);
or OR4 (N12667, N12664, N5881, N10279, N6334);
nand NAND3 (N12668, N12639, N743, N1048);
xor XOR2 (N12669, N12662, N10510);
or OR3 (N12670, N12656, N4530, N4307);
not NOT1 (N12671, N12669);
xor XOR2 (N12672, N12665, N5211);
xor XOR2 (N12673, N12670, N10079);
not NOT1 (N12674, N12666);
not NOT1 (N12675, N12672);
xor XOR2 (N12676, N12661, N8702);
not NOT1 (N12677, N12651);
or OR4 (N12678, N12675, N3911, N8859, N1865);
xor XOR2 (N12679, N12677, N9187);
nor NOR2 (N12680, N12673, N11504);
and AND4 (N12681, N12674, N429, N1661, N8117);
xor XOR2 (N12682, N12647, N1817);
buf BUF1 (N12683, N12671);
and AND2 (N12684, N12680, N9457);
nor NOR4 (N12685, N12679, N6662, N8866, N6781);
nor NOR4 (N12686, N12684, N5302, N11986, N8184);
and AND2 (N12687, N12676, N4288);
or OR3 (N12688, N12685, N9856, N1927);
nand NAND3 (N12689, N12688, N5983, N2423);
nand NAND4 (N12690, N12686, N3097, N4471, N7660);
nand NAND4 (N12691, N12683, N6425, N7227, N363);
buf BUF1 (N12692, N12691);
and AND4 (N12693, N12690, N4072, N9210, N10514);
not NOT1 (N12694, N12667);
nor NOR2 (N12695, N12657, N8929);
or OR2 (N12696, N12668, N6716);
and AND2 (N12697, N12682, N2309);
xor XOR2 (N12698, N12687, N4310);
xor XOR2 (N12699, N12695, N3586);
buf BUF1 (N12700, N12698);
xor XOR2 (N12701, N12693, N7193);
nand NAND2 (N12702, N12678, N795);
nand NAND4 (N12703, N12701, N9637, N9798, N8822);
buf BUF1 (N12704, N12700);
and AND2 (N12705, N12697, N10175);
nand NAND3 (N12706, N12699, N2667, N10083);
xor XOR2 (N12707, N12705, N9114);
not NOT1 (N12708, N12689);
or OR4 (N12709, N12694, N10341, N1370, N10509);
or OR4 (N12710, N12681, N5825, N10041, N11870);
buf BUF1 (N12711, N12696);
buf BUF1 (N12712, N12709);
nor NOR4 (N12713, N12712, N10824, N4379, N8528);
not NOT1 (N12714, N12692);
and AND3 (N12715, N12704, N2462, N10198);
not NOT1 (N12716, N12714);
and AND3 (N12717, N12702, N11602, N7742);
not NOT1 (N12718, N12717);
buf BUF1 (N12719, N12715);
nor NOR3 (N12720, N12718, N10274, N9248);
buf BUF1 (N12721, N12720);
xor XOR2 (N12722, N12716, N7665);
xor XOR2 (N12723, N12708, N5145);
xor XOR2 (N12724, N12710, N5211);
nand NAND2 (N12725, N12703, N3805);
nand NAND4 (N12726, N12719, N9146, N5860, N9693);
nor NOR2 (N12727, N12726, N2650);
or OR4 (N12728, N12725, N4363, N10314, N1820);
buf BUF1 (N12729, N12722);
and AND3 (N12730, N12706, N242, N10028);
or OR2 (N12731, N12713, N8517);
nand NAND3 (N12732, N12721, N1336, N6967);
not NOT1 (N12733, N12724);
buf BUF1 (N12734, N12729);
xor XOR2 (N12735, N12733, N3672);
nor NOR2 (N12736, N12728, N5555);
nand NAND2 (N12737, N12707, N10888);
and AND2 (N12738, N12727, N5649);
or OR2 (N12739, N12735, N8252);
or OR4 (N12740, N12738, N1756, N12585, N197);
xor XOR2 (N12741, N12740, N7826);
nor NOR3 (N12742, N12723, N4493, N3702);
nor NOR3 (N12743, N12731, N1117, N9005);
nor NOR3 (N12744, N12743, N2037, N7665);
or OR4 (N12745, N12739, N7559, N482, N5315);
buf BUF1 (N12746, N12711);
nor NOR4 (N12747, N12746, N2724, N960, N4979);
nand NAND4 (N12748, N12737, N9250, N1277, N6999);
and AND4 (N12749, N12736, N10622, N8560, N7261);
nand NAND3 (N12750, N12748, N8219, N4962);
or OR4 (N12751, N12747, N3312, N248, N5848);
nand NAND2 (N12752, N12730, N8257);
xor XOR2 (N12753, N12745, N9912);
or OR4 (N12754, N12749, N12128, N4395, N11785);
and AND4 (N12755, N12750, N2241, N6724, N6732);
not NOT1 (N12756, N12732);
nor NOR4 (N12757, N12751, N8120, N10309, N5910);
not NOT1 (N12758, N12752);
and AND2 (N12759, N12758, N12634);
buf BUF1 (N12760, N12756);
xor XOR2 (N12761, N12754, N10573);
buf BUF1 (N12762, N12755);
nor NOR3 (N12763, N12741, N1982, N11346);
and AND4 (N12764, N12753, N7195, N2976, N8083);
xor XOR2 (N12765, N12759, N1200);
not NOT1 (N12766, N12761);
buf BUF1 (N12767, N12762);
or OR2 (N12768, N12744, N5473);
and AND4 (N12769, N12767, N12436, N9609, N11118);
buf BUF1 (N12770, N12768);
nor NOR2 (N12771, N12757, N5761);
nor NOR3 (N12772, N12766, N3491, N4702);
xor XOR2 (N12773, N12771, N6709);
and AND3 (N12774, N12773, N6973, N12623);
buf BUF1 (N12775, N12764);
buf BUF1 (N12776, N12769);
xor XOR2 (N12777, N12775, N8624);
xor XOR2 (N12778, N12763, N6605);
xor XOR2 (N12779, N12774, N12235);
or OR2 (N12780, N12765, N3013);
xor XOR2 (N12781, N12772, N7541);
and AND4 (N12782, N12780, N3640, N8660, N12758);
not NOT1 (N12783, N12778);
or OR3 (N12784, N12781, N751, N2557);
nand NAND2 (N12785, N12742, N6560);
and AND2 (N12786, N12779, N9116);
xor XOR2 (N12787, N12776, N7175);
or OR2 (N12788, N12787, N6851);
and AND2 (N12789, N12734, N12587);
and AND2 (N12790, N12785, N5067);
buf BUF1 (N12791, N12784);
not NOT1 (N12792, N12790);
buf BUF1 (N12793, N12786);
not NOT1 (N12794, N12792);
and AND3 (N12795, N12783, N4632, N2339);
nand NAND3 (N12796, N12793, N4603, N2079);
nand NAND2 (N12797, N12782, N3043);
nand NAND2 (N12798, N12777, N1205);
buf BUF1 (N12799, N12796);
nand NAND2 (N12800, N12788, N11158);
buf BUF1 (N12801, N12791);
buf BUF1 (N12802, N12798);
nand NAND3 (N12803, N12795, N4476, N6500);
and AND3 (N12804, N12799, N11686, N5961);
nor NOR3 (N12805, N12797, N4440, N6572);
xor XOR2 (N12806, N12801, N12431);
not NOT1 (N12807, N12760);
and AND3 (N12808, N12802, N11616, N5333);
nor NOR2 (N12809, N12794, N447);
nor NOR3 (N12810, N12770, N10692, N7021);
and AND4 (N12811, N12809, N3300, N4798, N7181);
or OR2 (N12812, N12807, N10178);
and AND3 (N12813, N12806, N12197, N10008);
buf BUF1 (N12814, N12804);
xor XOR2 (N12815, N12789, N2598);
and AND4 (N12816, N12810, N4763, N664, N11400);
or OR3 (N12817, N12800, N1158, N7866);
and AND4 (N12818, N12808, N198, N12504, N11239);
nand NAND4 (N12819, N12818, N2615, N6494, N4516);
buf BUF1 (N12820, N12814);
and AND2 (N12821, N12813, N1474);
not NOT1 (N12822, N12820);
buf BUF1 (N12823, N12812);
buf BUF1 (N12824, N12815);
and AND4 (N12825, N12811, N4805, N5260, N10348);
nor NOR4 (N12826, N12805, N5650, N4390, N5417);
and AND2 (N12827, N12825, N3884);
buf BUF1 (N12828, N12816);
nor NOR4 (N12829, N12822, N3960, N6602, N11064);
buf BUF1 (N12830, N12829);
nor NOR4 (N12831, N12826, N5815, N5176, N12356);
nor NOR4 (N12832, N12803, N1177, N7303, N3048);
not NOT1 (N12833, N12830);
not NOT1 (N12834, N12832);
not NOT1 (N12835, N12827);
buf BUF1 (N12836, N12828);
not NOT1 (N12837, N12823);
or OR2 (N12838, N12819, N2999);
or OR2 (N12839, N12824, N6018);
and AND3 (N12840, N12833, N7243, N7239);
nand NAND4 (N12841, N12836, N9230, N1908, N10894);
buf BUF1 (N12842, N12831);
xor XOR2 (N12843, N12834, N99);
nor NOR4 (N12844, N12817, N7034, N7142, N7598);
buf BUF1 (N12845, N12837);
nor NOR4 (N12846, N12821, N12005, N618, N3381);
or OR3 (N12847, N12838, N130, N3409);
or OR4 (N12848, N12835, N12822, N675, N4813);
or OR4 (N12849, N12847, N9667, N4716, N6017);
buf BUF1 (N12850, N12840);
xor XOR2 (N12851, N12849, N10314);
nor NOR4 (N12852, N12842, N1132, N12517, N9594);
or OR4 (N12853, N12839, N11204, N6355, N548);
buf BUF1 (N12854, N12844);
buf BUF1 (N12855, N12851);
nor NOR3 (N12856, N12850, N10624, N10494);
xor XOR2 (N12857, N12845, N9092);
and AND2 (N12858, N12853, N2366);
nor NOR4 (N12859, N12846, N4319, N5957, N3213);
nand NAND3 (N12860, N12848, N665, N12283);
buf BUF1 (N12861, N12858);
nand NAND3 (N12862, N12857, N12671, N8787);
nor NOR4 (N12863, N12860, N6221, N11363, N12568);
or OR3 (N12864, N12862, N7638, N10610);
xor XOR2 (N12865, N12861, N4886);
nand NAND2 (N12866, N12852, N6036);
xor XOR2 (N12867, N12865, N9616);
not NOT1 (N12868, N12859);
not NOT1 (N12869, N12856);
xor XOR2 (N12870, N12841, N3583);
and AND4 (N12871, N12867, N7705, N7153, N6800);
xor XOR2 (N12872, N12854, N9667);
or OR3 (N12873, N12871, N8346, N3069);
xor XOR2 (N12874, N12866, N10118);
buf BUF1 (N12875, N12870);
nor NOR2 (N12876, N12864, N9650);
not NOT1 (N12877, N12876);
not NOT1 (N12878, N12872);
buf BUF1 (N12879, N12863);
buf BUF1 (N12880, N12875);
or OR2 (N12881, N12877, N4332);
not NOT1 (N12882, N12873);
and AND3 (N12883, N12881, N1786, N4895);
and AND4 (N12884, N12843, N1112, N4854, N9768);
not NOT1 (N12885, N12878);
or OR2 (N12886, N12874, N131);
or OR3 (N12887, N12883, N8780, N11321);
buf BUF1 (N12888, N12879);
xor XOR2 (N12889, N12880, N10066);
and AND4 (N12890, N12869, N4134, N11958, N4603);
or OR4 (N12891, N12886, N5982, N2099, N11581);
nor NOR3 (N12892, N12890, N5932, N3615);
and AND2 (N12893, N12884, N1856);
nor NOR2 (N12894, N12855, N10768);
and AND2 (N12895, N12894, N8643);
nor NOR3 (N12896, N12885, N7095, N6794);
xor XOR2 (N12897, N12896, N2352);
buf BUF1 (N12898, N12895);
nor NOR2 (N12899, N12887, N4561);
and AND4 (N12900, N12899, N5345, N5012, N10406);
xor XOR2 (N12901, N12897, N617);
xor XOR2 (N12902, N12901, N5512);
nor NOR3 (N12903, N12893, N4777, N6321);
xor XOR2 (N12904, N12882, N5585);
xor XOR2 (N12905, N12888, N10751);
xor XOR2 (N12906, N12905, N2828);
xor XOR2 (N12907, N12902, N7749);
and AND3 (N12908, N12906, N4416, N1554);
buf BUF1 (N12909, N12891);
nor NOR2 (N12910, N12907, N2037);
nand NAND3 (N12911, N12889, N12306, N3348);
or OR2 (N12912, N12892, N113);
buf BUF1 (N12913, N12909);
nand NAND2 (N12914, N12913, N2778);
buf BUF1 (N12915, N12904);
buf BUF1 (N12916, N12911);
or OR3 (N12917, N12915, N10403, N1241);
and AND2 (N12918, N12900, N8741);
nor NOR4 (N12919, N12916, N701, N9622, N6764);
buf BUF1 (N12920, N12903);
buf BUF1 (N12921, N12919);
xor XOR2 (N12922, N12898, N2844);
not NOT1 (N12923, N12920);
nand NAND2 (N12924, N12918, N12240);
xor XOR2 (N12925, N12922, N12461);
buf BUF1 (N12926, N12924);
nor NOR2 (N12927, N12923, N1953);
and AND2 (N12928, N12912, N4044);
buf BUF1 (N12929, N12926);
nor NOR4 (N12930, N12925, N12424, N5105, N5253);
and AND3 (N12931, N12910, N8348, N1297);
not NOT1 (N12932, N12929);
buf BUF1 (N12933, N12917);
nor NOR3 (N12934, N12930, N7730, N6096);
nand NAND4 (N12935, N12928, N10952, N8922, N5375);
and AND2 (N12936, N12914, N3096);
or OR3 (N12937, N12931, N10972, N10738);
nand NAND4 (N12938, N12935, N10472, N6885, N9024);
xor XOR2 (N12939, N12933, N3012);
and AND2 (N12940, N12934, N743);
or OR4 (N12941, N12932, N6114, N7130, N6982);
nor NOR2 (N12942, N12927, N11083);
buf BUF1 (N12943, N12939);
xor XOR2 (N12944, N12936, N9170);
not NOT1 (N12945, N12938);
not NOT1 (N12946, N12940);
xor XOR2 (N12947, N12868, N3930);
xor XOR2 (N12948, N12945, N7892);
not NOT1 (N12949, N12947);
nand NAND4 (N12950, N12943, N12438, N10633, N9968);
buf BUF1 (N12951, N12921);
nand NAND3 (N12952, N12941, N9027, N5650);
nor NOR2 (N12953, N12948, N11826);
buf BUF1 (N12954, N12908);
not NOT1 (N12955, N12953);
xor XOR2 (N12956, N12955, N4995);
nor NOR3 (N12957, N12951, N3729, N9536);
nand NAND4 (N12958, N12944, N126, N7219, N9912);
buf BUF1 (N12959, N12958);
and AND4 (N12960, N12937, N7140, N3538, N8467);
nor NOR4 (N12961, N12946, N189, N12672, N1579);
xor XOR2 (N12962, N12942, N7085);
buf BUF1 (N12963, N12950);
not NOT1 (N12964, N12949);
xor XOR2 (N12965, N12959, N7410);
buf BUF1 (N12966, N12952);
not NOT1 (N12967, N12964);
xor XOR2 (N12968, N12967, N8602);
not NOT1 (N12969, N12957);
buf BUF1 (N12970, N12966);
buf BUF1 (N12971, N12963);
xor XOR2 (N12972, N12960, N4028);
nor NOR3 (N12973, N12968, N11993, N11145);
nor NOR2 (N12974, N12971, N8507);
and AND4 (N12975, N12961, N12735, N3645, N11251);
nor NOR2 (N12976, N12975, N2881);
not NOT1 (N12977, N12976);
and AND2 (N12978, N12972, N4293);
buf BUF1 (N12979, N12954);
buf BUF1 (N12980, N12979);
or OR4 (N12981, N12973, N6728, N10038, N9716);
not NOT1 (N12982, N12956);
or OR2 (N12983, N12962, N4086);
xor XOR2 (N12984, N12974, N6276);
nor NOR3 (N12985, N12970, N8313, N1667);
and AND2 (N12986, N12985, N232);
nand NAND3 (N12987, N12981, N3694, N6817);
nor NOR3 (N12988, N12980, N12577, N5639);
not NOT1 (N12989, N12983);
buf BUF1 (N12990, N12987);
or OR3 (N12991, N12989, N245, N4550);
buf BUF1 (N12992, N12969);
and AND3 (N12993, N12992, N6268, N6533);
or OR3 (N12994, N12982, N5340, N719);
xor XOR2 (N12995, N12984, N8787);
xor XOR2 (N12996, N12993, N6624);
or OR4 (N12997, N12994, N12844, N12394, N9783);
nand NAND2 (N12998, N12986, N7308);
and AND2 (N12999, N12991, N1925);
nand NAND2 (N13000, N12999, N8069);
nor NOR2 (N13001, N12996, N1730);
not NOT1 (N13002, N12997);
and AND4 (N13003, N13002, N7978, N8627, N6274);
xor XOR2 (N13004, N12965, N6267);
or OR3 (N13005, N13000, N2767, N4685);
not NOT1 (N13006, N13003);
xor XOR2 (N13007, N12988, N6887);
buf BUF1 (N13008, N12995);
or OR2 (N13009, N13006, N1148);
nand NAND2 (N13010, N12998, N6948);
or OR4 (N13011, N13005, N10405, N2202, N8225);
nand NAND2 (N13012, N13008, N12804);
nand NAND4 (N13013, N13011, N12815, N8775, N9995);
and AND3 (N13014, N13001, N12633, N7717);
nand NAND2 (N13015, N12977, N636);
nand NAND3 (N13016, N13014, N2940, N7586);
nor NOR4 (N13017, N13015, N10369, N3794, N3405);
xor XOR2 (N13018, N13009, N4618);
nand NAND3 (N13019, N13004, N10276, N6732);
or OR3 (N13020, N13017, N10447, N2859);
buf BUF1 (N13021, N12990);
and AND2 (N13022, N13020, N11551);
or OR4 (N13023, N13013, N1310, N9125, N12446);
buf BUF1 (N13024, N13021);
and AND3 (N13025, N13018, N8516, N11547);
nand NAND2 (N13026, N12978, N6659);
buf BUF1 (N13027, N13010);
and AND3 (N13028, N13022, N4277, N6035);
xor XOR2 (N13029, N13025, N6535);
xor XOR2 (N13030, N13019, N10153);
buf BUF1 (N13031, N13028);
nand NAND3 (N13032, N13029, N9372, N5751);
buf BUF1 (N13033, N13007);
buf BUF1 (N13034, N13031);
nand NAND4 (N13035, N13033, N7216, N11917, N8974);
and AND3 (N13036, N13023, N4684, N4131);
xor XOR2 (N13037, N13016, N11183);
and AND2 (N13038, N13030, N2404);
or OR4 (N13039, N13034, N6728, N12948, N4163);
or OR2 (N13040, N13012, N12472);
not NOT1 (N13041, N13040);
xor XOR2 (N13042, N13027, N12749);
nor NOR3 (N13043, N13024, N6648, N6322);
nor NOR2 (N13044, N13042, N1494);
buf BUF1 (N13045, N13035);
xor XOR2 (N13046, N13043, N11623);
not NOT1 (N13047, N13037);
xor XOR2 (N13048, N13046, N4585);
xor XOR2 (N13049, N13038, N5169);
nand NAND3 (N13050, N13047, N9828, N8698);
buf BUF1 (N13051, N13032);
buf BUF1 (N13052, N13050);
nor NOR2 (N13053, N13045, N11432);
nor NOR4 (N13054, N13052, N6498, N3619, N1491);
nand NAND4 (N13055, N13051, N5081, N5631, N9611);
nor NOR4 (N13056, N13039, N2524, N6474, N12649);
or OR4 (N13057, N13026, N1593, N6960, N11821);
xor XOR2 (N13058, N13057, N3102);
or OR2 (N13059, N13044, N8287);
and AND4 (N13060, N13055, N6138, N11458, N996);
nor NOR3 (N13061, N13054, N3698, N206);
or OR3 (N13062, N13060, N4470, N10671);
or OR3 (N13063, N13059, N11497, N10949);
xor XOR2 (N13064, N13061, N319);
xor XOR2 (N13065, N13041, N11451);
xor XOR2 (N13066, N13049, N1647);
nand NAND3 (N13067, N13063, N1630, N11999);
nand NAND3 (N13068, N13036, N6878, N11910);
or OR4 (N13069, N13056, N776, N2596, N2205);
xor XOR2 (N13070, N13048, N12490);
and AND4 (N13071, N13053, N12945, N3509, N2787);
nor NOR4 (N13072, N13066, N13071, N6407, N1427);
and AND2 (N13073, N7173, N9478);
not NOT1 (N13074, N13072);
or OR4 (N13075, N13067, N8307, N8203, N7568);
not NOT1 (N13076, N13073);
nand NAND2 (N13077, N13076, N8212);
buf BUF1 (N13078, N13064);
or OR4 (N13079, N13077, N9065, N95, N2624);
and AND2 (N13080, N13065, N6630);
nand NAND3 (N13081, N13062, N1800, N4205);
not NOT1 (N13082, N13069);
nand NAND3 (N13083, N13081, N12995, N2605);
xor XOR2 (N13084, N13083, N4200);
or OR3 (N13085, N13058, N106, N6253);
buf BUF1 (N13086, N13074);
xor XOR2 (N13087, N13068, N10040);
not NOT1 (N13088, N13087);
xor XOR2 (N13089, N13088, N1823);
nand NAND3 (N13090, N13086, N6127, N12292);
xor XOR2 (N13091, N13075, N11713);
xor XOR2 (N13092, N13091, N12937);
and AND4 (N13093, N13085, N8909, N9434, N12544);
nand NAND3 (N13094, N13093, N1371, N2301);
or OR3 (N13095, N13070, N8835, N1047);
xor XOR2 (N13096, N13079, N5731);
nor NOR3 (N13097, N13090, N12583, N5890);
and AND3 (N13098, N13092, N7236, N11438);
and AND2 (N13099, N13095, N5167);
nor NOR4 (N13100, N13084, N10180, N10955, N6383);
nand NAND2 (N13101, N13089, N4977);
not NOT1 (N13102, N13098);
xor XOR2 (N13103, N13102, N5818);
nor NOR4 (N13104, N13096, N670, N7640, N11475);
nor NOR4 (N13105, N13097, N11424, N5126, N6799);
xor XOR2 (N13106, N13094, N11369);
xor XOR2 (N13107, N13103, N4492);
buf BUF1 (N13108, N13107);
nor NOR4 (N13109, N13101, N5652, N998, N2139);
xor XOR2 (N13110, N13109, N3702);
and AND3 (N13111, N13105, N5163, N1916);
xor XOR2 (N13112, N13099, N12042);
or OR2 (N13113, N13110, N1930);
not NOT1 (N13114, N13106);
xor XOR2 (N13115, N13113, N323);
not NOT1 (N13116, N13111);
not NOT1 (N13117, N13115);
nand NAND2 (N13118, N13078, N11493);
not NOT1 (N13119, N13116);
buf BUF1 (N13120, N13104);
and AND2 (N13121, N13118, N11460);
buf BUF1 (N13122, N13119);
and AND3 (N13123, N13080, N1412, N3501);
not NOT1 (N13124, N13122);
xor XOR2 (N13125, N13121, N3046);
xor XOR2 (N13126, N13114, N6147);
nand NAND4 (N13127, N13112, N8747, N6649, N9845);
buf BUF1 (N13128, N13127);
or OR4 (N13129, N13108, N8860, N10603, N8824);
or OR3 (N13130, N13082, N2131, N9776);
buf BUF1 (N13131, N13130);
or OR4 (N13132, N13123, N6654, N8931, N2549);
not NOT1 (N13133, N13132);
nand NAND2 (N13134, N13117, N561);
buf BUF1 (N13135, N13126);
nor NOR2 (N13136, N13100, N4035);
not NOT1 (N13137, N13125);
xor XOR2 (N13138, N13129, N6676);
nor NOR4 (N13139, N13120, N11509, N10421, N11525);
and AND4 (N13140, N13137, N3174, N3709, N251);
nand NAND2 (N13141, N13134, N6398);
or OR4 (N13142, N13133, N1011, N1416, N2519);
or OR2 (N13143, N13138, N11471);
nand NAND3 (N13144, N13143, N3689, N11998);
xor XOR2 (N13145, N13131, N2193);
not NOT1 (N13146, N13144);
and AND4 (N13147, N13140, N1916, N12808, N5378);
buf BUF1 (N13148, N13124);
not NOT1 (N13149, N13142);
or OR3 (N13150, N13148, N7487, N605);
and AND4 (N13151, N13128, N8553, N10095, N3102);
buf BUF1 (N13152, N13136);
or OR3 (N13153, N13147, N9681, N317);
not NOT1 (N13154, N13149);
nand NAND3 (N13155, N13154, N9121, N8672);
nand NAND2 (N13156, N13139, N12628);
not NOT1 (N13157, N13151);
not NOT1 (N13158, N13155);
or OR3 (N13159, N13156, N7473, N13082);
nor NOR4 (N13160, N13158, N5443, N4541, N3130);
not NOT1 (N13161, N13153);
and AND3 (N13162, N13146, N5273, N8598);
and AND3 (N13163, N13152, N13152, N6474);
xor XOR2 (N13164, N13159, N3623);
nor NOR2 (N13165, N13141, N4258);
nand NAND3 (N13166, N13135, N1871, N3396);
buf BUF1 (N13167, N13150);
nor NOR3 (N13168, N13160, N9040, N10922);
buf BUF1 (N13169, N13165);
or OR3 (N13170, N13169, N13067, N3832);
buf BUF1 (N13171, N13170);
not NOT1 (N13172, N13164);
or OR4 (N13173, N13167, N5402, N10494, N2661);
buf BUF1 (N13174, N13172);
xor XOR2 (N13175, N13161, N3286);
nor NOR4 (N13176, N13173, N11888, N120, N6742);
or OR2 (N13177, N13166, N4320);
nor NOR3 (N13178, N13145, N11965, N12200);
nand NAND4 (N13179, N13178, N6528, N9883, N10379);
buf BUF1 (N13180, N13171);
nand NAND4 (N13181, N13157, N9817, N645, N7278);
or OR2 (N13182, N13176, N2047);
nor NOR4 (N13183, N13182, N5886, N1623, N6326);
and AND3 (N13184, N13168, N5993, N4261);
nor NOR4 (N13185, N13184, N391, N12721, N1609);
not NOT1 (N13186, N13177);
buf BUF1 (N13187, N13180);
and AND2 (N13188, N13183, N10927);
and AND3 (N13189, N13188, N4114, N11317);
buf BUF1 (N13190, N13189);
buf BUF1 (N13191, N13179);
not NOT1 (N13192, N13174);
not NOT1 (N13193, N13163);
or OR3 (N13194, N13193, N3062, N13101);
and AND4 (N13195, N13187, N11249, N4951, N232);
and AND2 (N13196, N13191, N3447);
xor XOR2 (N13197, N13185, N11924);
xor XOR2 (N13198, N13181, N3780);
nor NOR4 (N13199, N13190, N9175, N11620, N4251);
not NOT1 (N13200, N13175);
xor XOR2 (N13201, N13200, N3551);
nand NAND4 (N13202, N13194, N1479, N787, N290);
nand NAND3 (N13203, N13192, N9440, N11120);
or OR2 (N13204, N13198, N1414);
nand NAND4 (N13205, N13203, N11040, N11361, N393);
and AND3 (N13206, N13162, N2318, N6295);
xor XOR2 (N13207, N13195, N129);
or OR2 (N13208, N13205, N10516);
not NOT1 (N13209, N13199);
or OR2 (N13210, N13209, N8305);
nand NAND3 (N13211, N13207, N12802, N12174);
buf BUF1 (N13212, N13196);
xor XOR2 (N13213, N13202, N5108);
not NOT1 (N13214, N13211);
nor NOR3 (N13215, N13208, N12234, N9055);
xor XOR2 (N13216, N13201, N1696);
not NOT1 (N13217, N13204);
nand NAND3 (N13218, N13212, N12676, N9103);
nand NAND3 (N13219, N13197, N3410, N1030);
nand NAND2 (N13220, N13219, N11603);
or OR3 (N13221, N13213, N6419, N12301);
and AND2 (N13222, N13220, N2923);
not NOT1 (N13223, N13210);
nand NAND4 (N13224, N13223, N9710, N6705, N10910);
buf BUF1 (N13225, N13222);
nor NOR3 (N13226, N13215, N9260, N6821);
not NOT1 (N13227, N13225);
or OR4 (N13228, N13186, N4986, N11767, N9108);
xor XOR2 (N13229, N13226, N5549);
nand NAND2 (N13230, N13206, N2009);
nand NAND4 (N13231, N13224, N10548, N10819, N1106);
not NOT1 (N13232, N13217);
and AND4 (N13233, N13231, N453, N3519, N9747);
not NOT1 (N13234, N13227);
not NOT1 (N13235, N13230);
buf BUF1 (N13236, N13229);
or OR2 (N13237, N13235, N3276);
nand NAND2 (N13238, N13221, N10123);
nand NAND3 (N13239, N13216, N9991, N11879);
and AND3 (N13240, N13214, N8779, N5628);
or OR2 (N13241, N13239, N260);
or OR3 (N13242, N13240, N10631, N10059);
and AND3 (N13243, N13232, N9670, N2303);
nand NAND4 (N13244, N13237, N1739, N2512, N6208);
and AND3 (N13245, N13236, N5218, N4348);
nand NAND2 (N13246, N13218, N4399);
or OR3 (N13247, N13238, N4703, N9442);
nand NAND4 (N13248, N13234, N7413, N5036, N7188);
and AND2 (N13249, N13242, N1380);
and AND4 (N13250, N13246, N2904, N4190, N11462);
buf BUF1 (N13251, N13245);
or OR2 (N13252, N13241, N3764);
or OR4 (N13253, N13250, N12770, N3822, N11511);
xor XOR2 (N13254, N13251, N7282);
buf BUF1 (N13255, N13249);
nor NOR4 (N13256, N13255, N12254, N2415, N13217);
nor NOR2 (N13257, N13228, N3948);
xor XOR2 (N13258, N13256, N7434);
or OR3 (N13259, N13243, N10824, N9881);
buf BUF1 (N13260, N13233);
buf BUF1 (N13261, N13248);
or OR2 (N13262, N13254, N12749);
not NOT1 (N13263, N13247);
and AND3 (N13264, N13262, N6621, N2200);
or OR4 (N13265, N13261, N11140, N10402, N13160);
buf BUF1 (N13266, N13257);
nor NOR2 (N13267, N13253, N4943);
and AND4 (N13268, N13259, N2090, N2325, N6369);
not NOT1 (N13269, N13267);
nor NOR2 (N13270, N13266, N3214);
nor NOR4 (N13271, N13264, N474, N5730, N2566);
or OR3 (N13272, N13268, N10619, N707);
not NOT1 (N13273, N13272);
or OR2 (N13274, N13258, N2358);
xor XOR2 (N13275, N13263, N5739);
xor XOR2 (N13276, N13260, N3805);
buf BUF1 (N13277, N13269);
xor XOR2 (N13278, N13274, N7987);
nand NAND3 (N13279, N13271, N5921, N6282);
not NOT1 (N13280, N13277);
not NOT1 (N13281, N13276);
or OR3 (N13282, N13278, N4336, N6896);
and AND4 (N13283, N13282, N2430, N1710, N5991);
buf BUF1 (N13284, N13265);
and AND4 (N13285, N13281, N7099, N11804, N12509);
or OR4 (N13286, N13283, N11111, N9527, N10945);
nor NOR3 (N13287, N13286, N13206, N12131);
xor XOR2 (N13288, N13287, N794);
not NOT1 (N13289, N13244);
or OR4 (N13290, N13289, N7964, N10074, N1736);
or OR3 (N13291, N13285, N3255, N6800);
nor NOR3 (N13292, N13280, N7959, N2307);
nand NAND2 (N13293, N13279, N9396);
or OR3 (N13294, N13284, N3949, N2345);
nor NOR4 (N13295, N13275, N4243, N4254, N160);
nor NOR3 (N13296, N13273, N164, N6331);
buf BUF1 (N13297, N13294);
not NOT1 (N13298, N13296);
xor XOR2 (N13299, N13297, N8180);
nand NAND2 (N13300, N13290, N11525);
xor XOR2 (N13301, N13288, N10466);
or OR4 (N13302, N13295, N9753, N3629, N7163);
nand NAND2 (N13303, N13252, N2294);
or OR2 (N13304, N13301, N5747);
xor XOR2 (N13305, N13292, N5525);
and AND4 (N13306, N13298, N8692, N5396, N7724);
xor XOR2 (N13307, N13299, N8402);
or OR3 (N13308, N13305, N10388, N69);
buf BUF1 (N13309, N13307);
nand NAND4 (N13310, N13306, N9405, N11160, N11382);
and AND4 (N13311, N13293, N12510, N7098, N9845);
xor XOR2 (N13312, N13311, N9392);
buf BUF1 (N13313, N13270);
buf BUF1 (N13314, N13313);
buf BUF1 (N13315, N13303);
xor XOR2 (N13316, N13314, N6612);
not NOT1 (N13317, N13291);
nand NAND2 (N13318, N13317, N7379);
and AND2 (N13319, N13310, N13038);
xor XOR2 (N13320, N13302, N7638);
or OR4 (N13321, N13315, N10232, N5750, N10386);
buf BUF1 (N13322, N13320);
or OR2 (N13323, N13300, N432);
nand NAND3 (N13324, N13322, N9420, N10736);
nand NAND3 (N13325, N13318, N5839, N7249);
not NOT1 (N13326, N13304);
and AND4 (N13327, N13325, N5472, N7376, N10018);
and AND3 (N13328, N13324, N10796, N9689);
nor NOR2 (N13329, N13321, N4245);
not NOT1 (N13330, N13328);
nor NOR4 (N13331, N13309, N1348, N1397, N7497);
nand NAND2 (N13332, N13319, N989);
buf BUF1 (N13333, N13326);
buf BUF1 (N13334, N13312);
not NOT1 (N13335, N13331);
and AND3 (N13336, N13333, N4577, N1093);
not NOT1 (N13337, N13332);
xor XOR2 (N13338, N13334, N11220);
not NOT1 (N13339, N13337);
xor XOR2 (N13340, N13327, N7466);
nand NAND3 (N13341, N13340, N12351, N5655);
xor XOR2 (N13342, N13338, N7871);
nor NOR4 (N13343, N13341, N10972, N12403, N2308);
or OR3 (N13344, N13330, N8453, N2048);
xor XOR2 (N13345, N13323, N3271);
or OR4 (N13346, N13336, N8209, N5251, N10733);
not NOT1 (N13347, N13344);
buf BUF1 (N13348, N13308);
and AND2 (N13349, N13329, N3799);
or OR2 (N13350, N13347, N3901);
not NOT1 (N13351, N13335);
not NOT1 (N13352, N13345);
buf BUF1 (N13353, N13350);
xor XOR2 (N13354, N13348, N720);
buf BUF1 (N13355, N13342);
xor XOR2 (N13356, N13355, N3344);
or OR4 (N13357, N13346, N12462, N10279, N5110);
and AND3 (N13358, N13356, N6442, N140);
not NOT1 (N13359, N13349);
and AND2 (N13360, N13358, N3018);
nor NOR4 (N13361, N13360, N13174, N10428, N1810);
nand NAND3 (N13362, N13351, N12334, N3822);
and AND2 (N13363, N13361, N1020);
xor XOR2 (N13364, N13343, N12685);
and AND3 (N13365, N13339, N2883, N2161);
not NOT1 (N13366, N13354);
and AND2 (N13367, N13363, N8097);
xor XOR2 (N13368, N13362, N5406);
buf BUF1 (N13369, N13352);
not NOT1 (N13370, N13367);
and AND3 (N13371, N13353, N10802, N8510);
buf BUF1 (N13372, N13359);
or OR4 (N13373, N13316, N6346, N11888, N10438);
nand NAND4 (N13374, N13371, N5334, N195, N2331);
xor XOR2 (N13375, N13368, N61);
buf BUF1 (N13376, N13373);
buf BUF1 (N13377, N13365);
xor XOR2 (N13378, N13370, N12716);
nor NOR4 (N13379, N13364, N6586, N12507, N7507);
or OR3 (N13380, N13366, N1808, N12654);
nor NOR3 (N13381, N13378, N9708, N2434);
buf BUF1 (N13382, N13380);
nand NAND3 (N13383, N13375, N1219, N3203);
nor NOR2 (N13384, N13382, N1803);
buf BUF1 (N13385, N13381);
xor XOR2 (N13386, N13357, N9613);
or OR3 (N13387, N13379, N10184, N9907);
or OR3 (N13388, N13384, N12950, N5144);
not NOT1 (N13389, N13388);
and AND4 (N13390, N13383, N10977, N3545, N4447);
nand NAND2 (N13391, N13374, N6098);
and AND2 (N13392, N13387, N5420);
and AND2 (N13393, N13372, N5054);
and AND2 (N13394, N13369, N6279);
xor XOR2 (N13395, N13376, N12613);
and AND3 (N13396, N13385, N10009, N8592);
nor NOR3 (N13397, N13394, N9641, N4950);
not NOT1 (N13398, N13386);
not NOT1 (N13399, N13392);
xor XOR2 (N13400, N13390, N8874);
nand NAND3 (N13401, N13399, N1426, N3889);
not NOT1 (N13402, N13377);
nand NAND4 (N13403, N13395, N10413, N11918, N4074);
and AND4 (N13404, N13402, N9534, N8626, N11196);
nor NOR4 (N13405, N13401, N11327, N7030, N6828);
not NOT1 (N13406, N13398);
buf BUF1 (N13407, N13397);
nand NAND4 (N13408, N13400, N2352, N4464, N7335);
nand NAND4 (N13409, N13396, N9165, N4549, N2984);
nor NOR4 (N13410, N13391, N1572, N1873, N6566);
xor XOR2 (N13411, N13404, N642);
not NOT1 (N13412, N13393);
xor XOR2 (N13413, N13412, N4888);
xor XOR2 (N13414, N13408, N4737);
buf BUF1 (N13415, N13405);
buf BUF1 (N13416, N13403);
nand NAND3 (N13417, N13407, N2750, N2364);
nand NAND2 (N13418, N13406, N7678);
or OR3 (N13419, N13409, N2572, N13108);
not NOT1 (N13420, N13416);
nor NOR3 (N13421, N13389, N11845, N989);
xor XOR2 (N13422, N13421, N11997);
xor XOR2 (N13423, N13418, N9045);
xor XOR2 (N13424, N13420, N10095);
or OR2 (N13425, N13415, N2287);
xor XOR2 (N13426, N13417, N12755);
buf BUF1 (N13427, N13413);
or OR3 (N13428, N13414, N11749, N3360);
nand NAND4 (N13429, N13425, N7022, N8181, N11948);
or OR2 (N13430, N13419, N2911);
nand NAND2 (N13431, N13422, N8690);
xor XOR2 (N13432, N13431, N1799);
xor XOR2 (N13433, N13432, N8339);
nand NAND2 (N13434, N13428, N4634);
nand NAND4 (N13435, N13423, N3675, N424, N3428);
and AND3 (N13436, N13433, N10701, N10521);
not NOT1 (N13437, N13426);
buf BUF1 (N13438, N13436);
nand NAND3 (N13439, N13430, N4468, N5689);
or OR4 (N13440, N13437, N2935, N2894, N1734);
buf BUF1 (N13441, N13440);
and AND2 (N13442, N13410, N6145);
nor NOR3 (N13443, N13439, N5107, N11482);
nand NAND3 (N13444, N13434, N8467, N2355);
nand NAND3 (N13445, N13435, N3377, N10784);
nor NOR2 (N13446, N13443, N11029);
xor XOR2 (N13447, N13441, N7306);
and AND4 (N13448, N13442, N13394, N825, N7466);
nand NAND3 (N13449, N13445, N6311, N11338);
xor XOR2 (N13450, N13448, N12968);
nand NAND4 (N13451, N13450, N2469, N3591, N1711);
and AND4 (N13452, N13427, N12948, N4916, N7324);
not NOT1 (N13453, N13451);
and AND4 (N13454, N13411, N6491, N11030, N6135);
buf BUF1 (N13455, N13454);
xor XOR2 (N13456, N13444, N10589);
nand NAND2 (N13457, N13449, N6374);
nor NOR3 (N13458, N13424, N2206, N13141);
nand NAND3 (N13459, N13456, N5493, N10589);
nor NOR4 (N13460, N13457, N4159, N7164, N2774);
buf BUF1 (N13461, N13447);
not NOT1 (N13462, N13461);
nor NOR3 (N13463, N13462, N10735, N9159);
nor NOR2 (N13464, N13460, N10233);
nand NAND3 (N13465, N13459, N5229, N12350);
buf BUF1 (N13466, N13453);
and AND2 (N13467, N13452, N1504);
nand NAND4 (N13468, N13446, N12313, N2947, N3300);
xor XOR2 (N13469, N13438, N12116);
not NOT1 (N13470, N13458);
buf BUF1 (N13471, N13429);
or OR3 (N13472, N13466, N1743, N8178);
nand NAND2 (N13473, N13463, N5913);
and AND3 (N13474, N13473, N9756, N12428);
not NOT1 (N13475, N13472);
xor XOR2 (N13476, N13455, N9002);
or OR3 (N13477, N13475, N6769, N13138);
nand NAND4 (N13478, N13464, N1655, N10465, N9325);
buf BUF1 (N13479, N13476);
nand NAND2 (N13480, N13471, N7389);
nand NAND2 (N13481, N13468, N1449);
nor NOR4 (N13482, N13478, N3774, N5337, N10401);
nand NAND2 (N13483, N13479, N5323);
or OR2 (N13484, N13482, N3520);
not NOT1 (N13485, N13465);
buf BUF1 (N13486, N13481);
nand NAND4 (N13487, N13467, N7488, N1769, N615);
nor NOR3 (N13488, N13484, N11738, N5054);
or OR4 (N13489, N13470, N5703, N9054, N11167);
nand NAND4 (N13490, N13483, N11634, N13051, N5096);
or OR4 (N13491, N13474, N3487, N11493, N7017);
not NOT1 (N13492, N13485);
buf BUF1 (N13493, N13492);
xor XOR2 (N13494, N13469, N13154);
not NOT1 (N13495, N13488);
xor XOR2 (N13496, N13494, N1298);
buf BUF1 (N13497, N13477);
not NOT1 (N13498, N13493);
nand NAND2 (N13499, N13497, N3862);
and AND3 (N13500, N13489, N2465, N12296);
nand NAND3 (N13501, N13499, N3141, N12589);
nand NAND2 (N13502, N13500, N2340);
and AND2 (N13503, N13496, N3447);
not NOT1 (N13504, N13495);
nand NAND2 (N13505, N13498, N5963);
buf BUF1 (N13506, N13487);
and AND3 (N13507, N13504, N6461, N8362);
xor XOR2 (N13508, N13480, N2574);
xor XOR2 (N13509, N13506, N2793);
not NOT1 (N13510, N13501);
buf BUF1 (N13511, N13509);
nand NAND3 (N13512, N13490, N4877, N2796);
not NOT1 (N13513, N13510);
not NOT1 (N13514, N13486);
and AND4 (N13515, N13507, N1011, N12292, N8702);
nor NOR3 (N13516, N13514, N10055, N13074);
or OR3 (N13517, N13513, N265, N17);
nand NAND4 (N13518, N13503, N13308, N2369, N384);
not NOT1 (N13519, N13512);
nor NOR4 (N13520, N13518, N9910, N13487, N13273);
nor NOR2 (N13521, N13508, N669);
buf BUF1 (N13522, N13491);
nand NAND4 (N13523, N13520, N2322, N8410, N12693);
xor XOR2 (N13524, N13511, N12970);
and AND3 (N13525, N13524, N4894, N8466);
xor XOR2 (N13526, N13502, N8895);
and AND4 (N13527, N13523, N2122, N2894, N8601);
not NOT1 (N13528, N13521);
nor NOR3 (N13529, N13522, N4714, N9002);
not NOT1 (N13530, N13528);
nor NOR3 (N13531, N13519, N3060, N3247);
not NOT1 (N13532, N13505);
nand NAND3 (N13533, N13526, N4045, N11951);
or OR3 (N13534, N13533, N360, N6206);
not NOT1 (N13535, N13532);
and AND4 (N13536, N13530, N3568, N5037, N5040);
and AND3 (N13537, N13531, N3361, N12989);
buf BUF1 (N13538, N13527);
not NOT1 (N13539, N13529);
or OR2 (N13540, N13539, N1468);
not NOT1 (N13541, N13535);
not NOT1 (N13542, N13536);
or OR3 (N13543, N13525, N6988, N9446);
buf BUF1 (N13544, N13515);
nor NOR3 (N13545, N13516, N7269, N1192);
not NOT1 (N13546, N13541);
nand NAND4 (N13547, N13534, N8888, N7582, N11122);
nand NAND3 (N13548, N13544, N2148, N362);
or OR4 (N13549, N13538, N1899, N2738, N4607);
buf BUF1 (N13550, N13546);
and AND4 (N13551, N13549, N8962, N5251, N10348);
nor NOR4 (N13552, N13542, N6973, N7713, N9626);
not NOT1 (N13553, N13548);
and AND4 (N13554, N13543, N808, N1858, N162);
xor XOR2 (N13555, N13552, N4952);
not NOT1 (N13556, N13555);
nand NAND3 (N13557, N13554, N1280, N3766);
or OR3 (N13558, N13550, N7972, N2388);
not NOT1 (N13559, N13558);
not NOT1 (N13560, N13557);
buf BUF1 (N13561, N13553);
buf BUF1 (N13562, N13537);
or OR4 (N13563, N13551, N10037, N2662, N12715);
nor NOR2 (N13564, N13560, N5200);
buf BUF1 (N13565, N13517);
buf BUF1 (N13566, N13561);
xor XOR2 (N13567, N13556, N12134);
or OR3 (N13568, N13565, N6673, N9112);
nand NAND3 (N13569, N13547, N13074, N4393);
xor XOR2 (N13570, N13545, N2118);
nand NAND3 (N13571, N13563, N10084, N5520);
or OR4 (N13572, N13567, N3002, N7536, N11918);
or OR2 (N13573, N13562, N10408);
and AND2 (N13574, N13564, N3836);
xor XOR2 (N13575, N13570, N9523);
buf BUF1 (N13576, N13540);
and AND2 (N13577, N13575, N12477);
xor XOR2 (N13578, N13576, N12817);
buf BUF1 (N13579, N13578);
xor XOR2 (N13580, N13559, N8196);
and AND3 (N13581, N13569, N5227, N606);
and AND2 (N13582, N13574, N2018);
not NOT1 (N13583, N13573);
or OR2 (N13584, N13568, N11826);
buf BUF1 (N13585, N13577);
xor XOR2 (N13586, N13580, N11168);
xor XOR2 (N13587, N13572, N10130);
nor NOR3 (N13588, N13587, N6639, N8563);
nand NAND2 (N13589, N13579, N113);
or OR4 (N13590, N13582, N2846, N1169, N1671);
or OR4 (N13591, N13586, N2290, N10641, N4753);
not NOT1 (N13592, N13584);
xor XOR2 (N13593, N13588, N11099);
nand NAND3 (N13594, N13591, N1809, N5413);
nand NAND2 (N13595, N13592, N3502);
and AND2 (N13596, N13571, N11140);
xor XOR2 (N13597, N13595, N296);
and AND2 (N13598, N13583, N3912);
nor NOR4 (N13599, N13589, N11545, N6783, N8137);
buf BUF1 (N13600, N13566);
buf BUF1 (N13601, N13596);
buf BUF1 (N13602, N13598);
buf BUF1 (N13603, N13602);
not NOT1 (N13604, N13594);
nand NAND4 (N13605, N13603, N10504, N1063, N2315);
nor NOR4 (N13606, N13590, N11961, N6367, N10548);
xor XOR2 (N13607, N13593, N11170);
xor XOR2 (N13608, N13585, N9115);
nand NAND4 (N13609, N13607, N3778, N10657, N8531);
nand NAND3 (N13610, N13581, N3251, N7099);
not NOT1 (N13611, N13600);
xor XOR2 (N13612, N13605, N10982);
buf BUF1 (N13613, N13606);
and AND2 (N13614, N13610, N8899);
not NOT1 (N13615, N13612);
xor XOR2 (N13616, N13609, N2616);
not NOT1 (N13617, N13616);
buf BUF1 (N13618, N13617);
buf BUF1 (N13619, N13608);
buf BUF1 (N13620, N13611);
and AND4 (N13621, N13599, N11026, N6267, N13076);
and AND3 (N13622, N13620, N13127, N3334);
or OR3 (N13623, N13615, N7177, N3226);
nor NOR2 (N13624, N13601, N7293);
xor XOR2 (N13625, N13614, N8249);
xor XOR2 (N13626, N13604, N3571);
nand NAND4 (N13627, N13623, N4961, N13081, N7478);
buf BUF1 (N13628, N13622);
and AND3 (N13629, N13621, N7405, N5779);
not NOT1 (N13630, N13628);
nor NOR3 (N13631, N13597, N8382, N1063);
buf BUF1 (N13632, N13624);
and AND3 (N13633, N13619, N9352, N8385);
nor NOR2 (N13634, N13632, N13338);
nand NAND3 (N13635, N13627, N103, N9992);
xor XOR2 (N13636, N13630, N13304);
or OR2 (N13637, N13629, N9350);
not NOT1 (N13638, N13633);
not NOT1 (N13639, N13635);
nand NAND3 (N13640, N13638, N2866, N2380);
nand NAND4 (N13641, N13639, N8805, N5110, N1439);
nand NAND3 (N13642, N13636, N2465, N6097);
xor XOR2 (N13643, N13625, N3878);
nor NOR3 (N13644, N13618, N6508, N5911);
and AND4 (N13645, N13644, N205, N8713, N458);
nor NOR3 (N13646, N13637, N8187, N5823);
and AND2 (N13647, N13642, N9086);
xor XOR2 (N13648, N13643, N4645);
not NOT1 (N13649, N13641);
or OR4 (N13650, N13649, N1498, N10321, N11421);
not NOT1 (N13651, N13634);
and AND3 (N13652, N13631, N11624, N3810);
and AND4 (N13653, N13651, N6372, N6386, N10501);
xor XOR2 (N13654, N13648, N2838);
nand NAND4 (N13655, N13613, N4666, N5488, N6942);
buf BUF1 (N13656, N13647);
nand NAND4 (N13657, N13656, N12701, N5585, N3817);
or OR2 (N13658, N13640, N6758);
nand NAND2 (N13659, N13645, N4724);
and AND3 (N13660, N13655, N2152, N9009);
and AND2 (N13661, N13654, N145);
buf BUF1 (N13662, N13653);
nand NAND3 (N13663, N13650, N6402, N7499);
xor XOR2 (N13664, N13657, N3711);
and AND4 (N13665, N13659, N12409, N3183, N7472);
buf BUF1 (N13666, N13658);
nor NOR4 (N13667, N13660, N4577, N7016, N6190);
or OR3 (N13668, N13646, N12671, N310);
and AND3 (N13669, N13668, N469, N3380);
or OR3 (N13670, N13665, N5069, N8201);
and AND2 (N13671, N13667, N13540);
nand NAND2 (N13672, N13670, N1545);
and AND4 (N13673, N13671, N11723, N13553, N9787);
or OR4 (N13674, N13663, N59, N13096, N5367);
not NOT1 (N13675, N13626);
or OR2 (N13676, N13674, N1892);
nor NOR2 (N13677, N13662, N11214);
nand NAND2 (N13678, N13652, N11955);
and AND2 (N13679, N13678, N7355);
or OR2 (N13680, N13673, N5185);
not NOT1 (N13681, N13679);
not NOT1 (N13682, N13664);
nand NAND3 (N13683, N13666, N9854, N5158);
and AND3 (N13684, N13669, N6579, N1430);
nor NOR3 (N13685, N13684, N12901, N10713);
and AND4 (N13686, N13677, N2894, N8, N6118);
nand NAND2 (N13687, N13683, N12915);
xor XOR2 (N13688, N13672, N3893);
xor XOR2 (N13689, N13676, N6641);
xor XOR2 (N13690, N13682, N10121);
or OR2 (N13691, N13689, N5721);
and AND4 (N13692, N13686, N3362, N7592, N2316);
nor NOR3 (N13693, N13692, N11824, N3615);
xor XOR2 (N13694, N13675, N11942);
buf BUF1 (N13695, N13687);
buf BUF1 (N13696, N13693);
not NOT1 (N13697, N13694);
xor XOR2 (N13698, N13688, N1233);
and AND3 (N13699, N13681, N3168, N3476);
nand NAND2 (N13700, N13696, N3250);
nor NOR3 (N13701, N13690, N7486, N951);
xor XOR2 (N13702, N13661, N5463);
xor XOR2 (N13703, N13702, N5765);
buf BUF1 (N13704, N13697);
buf BUF1 (N13705, N13685);
nand NAND2 (N13706, N13680, N9793);
nand NAND2 (N13707, N13703, N11262);
and AND2 (N13708, N13691, N5576);
and AND3 (N13709, N13699, N28, N9609);
and AND3 (N13710, N13700, N2183, N1427);
and AND3 (N13711, N13710, N6167, N10005);
and AND3 (N13712, N13698, N8633, N2603);
xor XOR2 (N13713, N13701, N5764);
nand NAND3 (N13714, N13708, N2236, N2613);
nand NAND4 (N13715, N13706, N10489, N1839, N8958);
buf BUF1 (N13716, N13715);
not NOT1 (N13717, N13712);
buf BUF1 (N13718, N13717);
buf BUF1 (N13719, N13716);
not NOT1 (N13720, N13707);
and AND2 (N13721, N13718, N11063);
not NOT1 (N13722, N13719);
nand NAND4 (N13723, N13713, N7706, N1271, N3843);
buf BUF1 (N13724, N13720);
not NOT1 (N13725, N13721);
or OR4 (N13726, N13724, N8624, N4187, N13581);
nor NOR3 (N13727, N13722, N13486, N5526);
xor XOR2 (N13728, N13714, N1472);
or OR3 (N13729, N13695, N7414, N13338);
xor XOR2 (N13730, N13729, N9831);
nor NOR3 (N13731, N13726, N2580, N7982);
nor NOR4 (N13732, N13730, N5258, N265, N4368);
and AND2 (N13733, N13711, N10302);
and AND2 (N13734, N13709, N12232);
nor NOR2 (N13735, N13723, N10107);
nor NOR2 (N13736, N13735, N3261);
and AND2 (N13737, N13736, N8448);
or OR4 (N13738, N13728, N6797, N1454, N11617);
not NOT1 (N13739, N13731);
and AND4 (N13740, N13725, N4212, N670, N8872);
nand NAND3 (N13741, N13734, N11592, N1372);
nor NOR3 (N13742, N13733, N6588, N4298);
nor NOR3 (N13743, N13742, N11540, N4219);
nand NAND2 (N13744, N13741, N7292);
or OR2 (N13745, N13744, N5131);
not NOT1 (N13746, N13745);
or OR4 (N13747, N13743, N1320, N5255, N4341);
buf BUF1 (N13748, N13732);
buf BUF1 (N13749, N13704);
and AND2 (N13750, N13749, N9332);
nor NOR4 (N13751, N13740, N9263, N6252, N7927);
nor NOR4 (N13752, N13705, N4355, N286, N2942);
nand NAND3 (N13753, N13748, N3264, N828);
not NOT1 (N13754, N13750);
buf BUF1 (N13755, N13746);
nand NAND2 (N13756, N13738, N9223);
nand NAND4 (N13757, N13752, N6165, N1963, N5655);
buf BUF1 (N13758, N13737);
buf BUF1 (N13759, N13757);
or OR2 (N13760, N13754, N6907);
buf BUF1 (N13761, N13753);
buf BUF1 (N13762, N13758);
or OR4 (N13763, N13755, N2755, N11658, N10336);
and AND3 (N13764, N13756, N12346, N12740);
buf BUF1 (N13765, N13762);
not NOT1 (N13766, N13764);
nor NOR2 (N13767, N13727, N11419);
nor NOR4 (N13768, N13747, N3552, N6889, N46);
nand NAND4 (N13769, N13763, N3772, N3721, N11324);
buf BUF1 (N13770, N13760);
xor XOR2 (N13771, N13769, N1023);
or OR4 (N13772, N13771, N8292, N1983, N4311);
and AND3 (N13773, N13751, N12334, N2613);
and AND4 (N13774, N13766, N309, N12314, N2727);
not NOT1 (N13775, N13761);
nor NOR3 (N13776, N13770, N1894, N3302);
or OR3 (N13777, N13775, N1390, N8283);
nand NAND3 (N13778, N13773, N10502, N4354);
nor NOR4 (N13779, N13777, N13093, N11890, N12205);
or OR2 (N13780, N13779, N12463);
nand NAND4 (N13781, N13774, N3375, N11876, N2702);
and AND2 (N13782, N13778, N999);
and AND4 (N13783, N13776, N8111, N5921, N5162);
nand NAND2 (N13784, N13768, N7532);
nor NOR3 (N13785, N13739, N6712, N76);
or OR3 (N13786, N13767, N7262, N2634);
buf BUF1 (N13787, N13759);
nand NAND3 (N13788, N13785, N10621, N8503);
nor NOR2 (N13789, N13788, N6933);
or OR3 (N13790, N13787, N4229, N7770);
xor XOR2 (N13791, N13765, N1360);
nand NAND4 (N13792, N13791, N2162, N11254, N9451);
not NOT1 (N13793, N13783);
xor XOR2 (N13794, N13793, N8854);
nand NAND2 (N13795, N13794, N13524);
nand NAND3 (N13796, N13790, N1508, N7059);
nor NOR3 (N13797, N13796, N8203, N995);
nand NAND2 (N13798, N13784, N1193);
or OR2 (N13799, N13780, N10426);
nor NOR4 (N13800, N13789, N13157, N10356, N5885);
xor XOR2 (N13801, N13772, N8926);
nor NOR2 (N13802, N13795, N3605);
xor XOR2 (N13803, N13799, N11714);
not NOT1 (N13804, N13786);
xor XOR2 (N13805, N13797, N3558);
and AND2 (N13806, N13781, N10495);
nor NOR3 (N13807, N13805, N8148, N225);
xor XOR2 (N13808, N13804, N5448);
nand NAND3 (N13809, N13801, N9101, N4971);
not NOT1 (N13810, N13807);
nor NOR2 (N13811, N13809, N6838);
xor XOR2 (N13812, N13803, N11215);
nor NOR3 (N13813, N13782, N12694, N4604);
or OR2 (N13814, N13798, N6008);
or OR4 (N13815, N13808, N1536, N7235, N8086);
nand NAND3 (N13816, N13813, N12260, N9110);
or OR3 (N13817, N13812, N5037, N12852);
not NOT1 (N13818, N13800);
nand NAND4 (N13819, N13817, N8108, N3004, N9787);
not NOT1 (N13820, N13792);
not NOT1 (N13821, N13819);
and AND2 (N13822, N13814, N1333);
nand NAND4 (N13823, N13811, N2719, N5578, N7823);
nor NOR2 (N13824, N13818, N6327);
not NOT1 (N13825, N13823);
xor XOR2 (N13826, N13806, N13103);
nor NOR2 (N13827, N13826, N8809);
xor XOR2 (N13828, N13824, N4676);
and AND2 (N13829, N13822, N11166);
and AND2 (N13830, N13810, N3579);
nand NAND4 (N13831, N13828, N3093, N1568, N7195);
or OR4 (N13832, N13827, N8838, N9892, N11902);
buf BUF1 (N13833, N13816);
and AND2 (N13834, N13820, N11424);
not NOT1 (N13835, N13829);
buf BUF1 (N13836, N13825);
not NOT1 (N13837, N13830);
not NOT1 (N13838, N13832);
nor NOR2 (N13839, N13802, N1575);
not NOT1 (N13840, N13837);
nor NOR4 (N13841, N13838, N4521, N8072, N13189);
buf BUF1 (N13842, N13834);
buf BUF1 (N13843, N13831);
xor XOR2 (N13844, N13839, N7962);
nor NOR2 (N13845, N13840, N6479);
and AND3 (N13846, N13843, N4880, N987);
or OR4 (N13847, N13821, N729, N3663, N4464);
and AND2 (N13848, N13815, N3308);
and AND4 (N13849, N13844, N7347, N8638, N12953);
nor NOR4 (N13850, N13842, N9390, N4517, N5218);
or OR3 (N13851, N13845, N10604, N1727);
xor XOR2 (N13852, N13841, N2414);
not NOT1 (N13853, N13836);
xor XOR2 (N13854, N13853, N2973);
nor NOR4 (N13855, N13849, N6868, N140, N6880);
not NOT1 (N13856, N13851);
nor NOR2 (N13857, N13833, N10867);
not NOT1 (N13858, N13855);
and AND4 (N13859, N13846, N6885, N826, N6950);
or OR4 (N13860, N13850, N5374, N961, N4163);
buf BUF1 (N13861, N13860);
and AND4 (N13862, N13861, N12592, N9996, N10628);
buf BUF1 (N13863, N13858);
xor XOR2 (N13864, N13859, N4055);
buf BUF1 (N13865, N13863);
xor XOR2 (N13866, N13862, N5150);
nor NOR3 (N13867, N13847, N11564, N10434);
buf BUF1 (N13868, N13852);
or OR2 (N13869, N13854, N6591);
buf BUF1 (N13870, N13868);
nand NAND2 (N13871, N13867, N13446);
nor NOR2 (N13872, N13857, N10806);
or OR2 (N13873, N13866, N1228);
buf BUF1 (N13874, N13869);
nand NAND4 (N13875, N13864, N722, N3150, N6941);
or OR2 (N13876, N13865, N3000);
and AND2 (N13877, N13876, N7684);
and AND4 (N13878, N13856, N4976, N11528, N12392);
or OR2 (N13879, N13870, N6140);
or OR3 (N13880, N13878, N12485, N5628);
or OR4 (N13881, N13873, N5419, N2327, N4260);
nor NOR4 (N13882, N13880, N7599, N2950, N4142);
buf BUF1 (N13883, N13879);
xor XOR2 (N13884, N13882, N3517);
nor NOR4 (N13885, N13884, N5838, N7517, N4760);
or OR4 (N13886, N13875, N4195, N9743, N7415);
nor NOR4 (N13887, N13877, N4263, N12784, N1792);
xor XOR2 (N13888, N13885, N10852);
nor NOR4 (N13889, N13872, N8208, N10412, N8987);
xor XOR2 (N13890, N13871, N8352);
not NOT1 (N13891, N13890);
nor NOR4 (N13892, N13888, N10743, N8783, N10512);
not NOT1 (N13893, N13886);
nand NAND4 (N13894, N13881, N6331, N813, N5651);
xor XOR2 (N13895, N13892, N10309);
nand NAND2 (N13896, N13848, N5563);
or OR2 (N13897, N13887, N754);
nand NAND2 (N13898, N13894, N12685);
xor XOR2 (N13899, N13895, N9152);
xor XOR2 (N13900, N13893, N1205);
nor NOR3 (N13901, N13899, N1803, N13175);
and AND3 (N13902, N13889, N8726, N6724);
or OR4 (N13903, N13902, N9008, N3300, N7841);
nand NAND2 (N13904, N13883, N12602);
and AND2 (N13905, N13897, N9224);
or OR3 (N13906, N13835, N866, N10476);
nand NAND3 (N13907, N13891, N6353, N13839);
nand NAND2 (N13908, N13896, N11278);
buf BUF1 (N13909, N13905);
nand NAND3 (N13910, N13898, N6569, N4084);
and AND3 (N13911, N13907, N12773, N11417);
or OR2 (N13912, N13901, N3567);
and AND3 (N13913, N13874, N11049, N8654);
not NOT1 (N13914, N13900);
and AND4 (N13915, N13904, N151, N2881, N11604);
not NOT1 (N13916, N13909);
nor NOR2 (N13917, N13913, N1390);
not NOT1 (N13918, N13916);
nand NAND2 (N13919, N13910, N5962);
and AND3 (N13920, N13919, N10435, N4278);
xor XOR2 (N13921, N13903, N4377);
or OR4 (N13922, N13918, N9802, N3830, N11452);
nand NAND2 (N13923, N13920, N6405);
or OR3 (N13924, N13923, N6522, N12987);
buf BUF1 (N13925, N13906);
or OR2 (N13926, N13924, N2353);
xor XOR2 (N13927, N13922, N12718);
and AND2 (N13928, N13925, N8949);
nor NOR2 (N13929, N13927, N6462);
and AND2 (N13930, N13908, N9028);
buf BUF1 (N13931, N13930);
xor XOR2 (N13932, N13912, N11858);
xor XOR2 (N13933, N13926, N3605);
and AND2 (N13934, N13915, N3191);
buf BUF1 (N13935, N13932);
xor XOR2 (N13936, N13928, N3874);
not NOT1 (N13937, N13931);
and AND4 (N13938, N13917, N10964, N13232, N13023);
and AND4 (N13939, N13934, N12140, N12897, N9693);
not NOT1 (N13940, N13914);
nand NAND4 (N13941, N13940, N6502, N7074, N10194);
or OR2 (N13942, N13936, N2483);
buf BUF1 (N13943, N13935);
nor NOR3 (N13944, N13911, N3760, N11646);
or OR3 (N13945, N13944, N5661, N13496);
or OR2 (N13946, N13945, N5555);
xor XOR2 (N13947, N13942, N1388);
and AND4 (N13948, N13939, N9513, N9902, N6496);
and AND3 (N13949, N13929, N984, N7328);
buf BUF1 (N13950, N13943);
or OR2 (N13951, N13947, N4823);
not NOT1 (N13952, N13921);
nand NAND4 (N13953, N13949, N4984, N8900, N4039);
nand NAND4 (N13954, N13946, N4506, N3849, N5783);
and AND3 (N13955, N13937, N2926, N10972);
or OR3 (N13956, N13941, N10163, N7152);
not NOT1 (N13957, N13950);
and AND3 (N13958, N13938, N12811, N7485);
xor XOR2 (N13959, N13933, N8900);
or OR3 (N13960, N13958, N8922, N2346);
or OR3 (N13961, N13954, N4654, N2991);
nand NAND4 (N13962, N13951, N1673, N10675, N2554);
or OR2 (N13963, N13962, N10985);
nor NOR2 (N13964, N13961, N4834);
buf BUF1 (N13965, N13948);
buf BUF1 (N13966, N13957);
nor NOR4 (N13967, N13956, N13902, N2945, N5929);
or OR2 (N13968, N13963, N5284);
or OR3 (N13969, N13955, N10857, N2616);
xor XOR2 (N13970, N13968, N4216);
buf BUF1 (N13971, N13965);
nand NAND2 (N13972, N13959, N4982);
nand NAND4 (N13973, N13964, N2695, N5575, N350);
and AND3 (N13974, N13970, N1516, N2572);
xor XOR2 (N13975, N13952, N11779);
xor XOR2 (N13976, N13953, N1056);
nand NAND4 (N13977, N13967, N11876, N5226, N285);
nor NOR2 (N13978, N13969, N598);
nand NAND4 (N13979, N13976, N7837, N12751, N9334);
not NOT1 (N13980, N13978);
buf BUF1 (N13981, N13973);
not NOT1 (N13982, N13971);
nand NAND4 (N13983, N13979, N906, N60, N12239);
xor XOR2 (N13984, N13972, N162);
or OR3 (N13985, N13974, N10900, N6850);
buf BUF1 (N13986, N13984);
not NOT1 (N13987, N13981);
nor NOR2 (N13988, N13983, N11447);
not NOT1 (N13989, N13960);
xor XOR2 (N13990, N13989, N3727);
nor NOR3 (N13991, N13980, N8255, N4280);
and AND3 (N13992, N13991, N14, N6655);
buf BUF1 (N13993, N13982);
nor NOR3 (N13994, N13985, N9015, N5175);
and AND4 (N13995, N13977, N8472, N9252, N12985);
or OR3 (N13996, N13990, N8415, N5522);
nand NAND3 (N13997, N13992, N691, N13596);
and AND4 (N13998, N13993, N9850, N7077, N9747);
or OR2 (N13999, N13966, N972);
and AND3 (N14000, N13986, N10199, N9302);
buf BUF1 (N14001, N13988);
nand NAND2 (N14002, N13975, N5469);
and AND4 (N14003, N13994, N6286, N12947, N12789);
nand NAND2 (N14004, N13997, N8670);
xor XOR2 (N14005, N13999, N4153);
xor XOR2 (N14006, N13987, N2387);
and AND4 (N14007, N14002, N6301, N2295, N12294);
buf BUF1 (N14008, N14005);
buf BUF1 (N14009, N14008);
buf BUF1 (N14010, N14004);
nor NOR4 (N14011, N13998, N11217, N2087, N5957);
nand NAND3 (N14012, N14007, N9900, N571);
xor XOR2 (N14013, N14009, N3176);
or OR4 (N14014, N14012, N3767, N1703, N8211);
nand NAND4 (N14015, N14011, N2806, N7148, N11446);
or OR2 (N14016, N14001, N11238);
buf BUF1 (N14017, N14006);
and AND4 (N14018, N14003, N9590, N1897, N2095);
or OR2 (N14019, N14000, N11523);
nand NAND3 (N14020, N13996, N5591, N7577);
xor XOR2 (N14021, N14019, N12162);
or OR3 (N14022, N14018, N3164, N12544);
buf BUF1 (N14023, N14017);
not NOT1 (N14024, N14010);
nand NAND4 (N14025, N14021, N2703, N877, N5376);
xor XOR2 (N14026, N14013, N10943);
buf BUF1 (N14027, N14014);
nor NOR4 (N14028, N14020, N6072, N13978, N8504);
nand NAND4 (N14029, N14022, N12729, N4694, N6386);
or OR2 (N14030, N13995, N2818);
and AND4 (N14031, N14026, N7095, N10639, N4665);
xor XOR2 (N14032, N14015, N8290);
or OR2 (N14033, N14027, N8795);
buf BUF1 (N14034, N14030);
nand NAND2 (N14035, N14031, N3954);
buf BUF1 (N14036, N14016);
and AND3 (N14037, N14036, N11876, N550);
nor NOR4 (N14038, N14029, N631, N11922, N1499);
not NOT1 (N14039, N14028);
buf BUF1 (N14040, N14035);
nor NOR4 (N14041, N14025, N326, N4703, N4453);
buf BUF1 (N14042, N14037);
or OR2 (N14043, N14041, N6077);
buf BUF1 (N14044, N14042);
buf BUF1 (N14045, N14033);
xor XOR2 (N14046, N14024, N8756);
buf BUF1 (N14047, N14034);
and AND4 (N14048, N14043, N1867, N1559, N12850);
or OR4 (N14049, N14045, N5751, N9575, N1318);
not NOT1 (N14050, N14048);
not NOT1 (N14051, N14044);
or OR3 (N14052, N14049, N920, N121);
xor XOR2 (N14053, N14040, N2488);
and AND2 (N14054, N14032, N6853);
nand NAND3 (N14055, N14039, N1508, N10622);
nor NOR2 (N14056, N14046, N2236);
and AND4 (N14057, N14047, N3318, N7218, N12034);
nor NOR2 (N14058, N14050, N7380);
xor XOR2 (N14059, N14038, N6845);
and AND3 (N14060, N14056, N9783, N13280);
nor NOR4 (N14061, N14051, N3540, N8655, N7201);
nor NOR2 (N14062, N14060, N3776);
nor NOR4 (N14063, N14055, N6390, N4059, N8926);
xor XOR2 (N14064, N14061, N3235);
xor XOR2 (N14065, N14058, N3594);
nand NAND3 (N14066, N14057, N13715, N5493);
and AND4 (N14067, N14062, N3099, N3217, N5366);
nor NOR4 (N14068, N14065, N747, N9071, N6560);
xor XOR2 (N14069, N14059, N9414);
nor NOR3 (N14070, N14067, N3364, N10227);
nand NAND3 (N14071, N14053, N10646, N9947);
or OR3 (N14072, N14069, N10309, N4799);
xor XOR2 (N14073, N14064, N2581);
buf BUF1 (N14074, N14071);
nand NAND3 (N14075, N14072, N3002, N13579);
buf BUF1 (N14076, N14052);
nand NAND3 (N14077, N14070, N6967, N8992);
nand NAND4 (N14078, N14068, N596, N2831, N3322);
not NOT1 (N14079, N14077);
nor NOR3 (N14080, N14073, N5755, N3365);
and AND4 (N14081, N14066, N10894, N11815, N11247);
not NOT1 (N14082, N14079);
not NOT1 (N14083, N14063);
not NOT1 (N14084, N14078);
or OR2 (N14085, N14054, N11280);
nor NOR3 (N14086, N14080, N11866, N11182);
or OR4 (N14087, N14085, N312, N12626, N8434);
nand NAND4 (N14088, N14087, N5739, N360, N13186);
or OR2 (N14089, N14084, N6981);
not NOT1 (N14090, N14082);
nand NAND4 (N14091, N14088, N938, N2357, N11836);
xor XOR2 (N14092, N14075, N4502);
and AND3 (N14093, N14081, N8964, N5063);
xor XOR2 (N14094, N14093, N2647);
xor XOR2 (N14095, N14094, N8803);
xor XOR2 (N14096, N14095, N106);
buf BUF1 (N14097, N14096);
nor NOR3 (N14098, N14023, N9763, N13933);
or OR3 (N14099, N14091, N8269, N8954);
nand NAND4 (N14100, N14074, N823, N2521, N5935);
nand NAND4 (N14101, N14097, N12752, N4594, N174);
or OR4 (N14102, N14100, N9635, N4625, N12968);
nand NAND4 (N14103, N14076, N10310, N4177, N639);
nand NAND3 (N14104, N14099, N11960, N1567);
buf BUF1 (N14105, N14104);
or OR4 (N14106, N14083, N4845, N10548, N914);
or OR3 (N14107, N14090, N12283, N591);
nor NOR3 (N14108, N14089, N3930, N6129);
nor NOR4 (N14109, N14108, N13103, N3443, N13061);
buf BUF1 (N14110, N14103);
xor XOR2 (N14111, N14098, N741);
and AND3 (N14112, N14110, N10327, N6065);
nand NAND3 (N14113, N14109, N2635, N9742);
not NOT1 (N14114, N14107);
not NOT1 (N14115, N14112);
not NOT1 (N14116, N14086);
or OR3 (N14117, N14116, N9741, N14087);
not NOT1 (N14118, N14115);
not NOT1 (N14119, N14111);
buf BUF1 (N14120, N14106);
not NOT1 (N14121, N14102);
buf BUF1 (N14122, N14092);
nand NAND2 (N14123, N14117, N5108);
not NOT1 (N14124, N14114);
or OR4 (N14125, N14105, N9910, N5032, N1835);
nand NAND3 (N14126, N14122, N969, N6548);
not NOT1 (N14127, N14118);
or OR3 (N14128, N14123, N4657, N11903);
nor NOR4 (N14129, N14120, N11484, N9152, N8361);
not NOT1 (N14130, N14121);
or OR4 (N14131, N14113, N8532, N6889, N9528);
buf BUF1 (N14132, N14119);
or OR4 (N14133, N14125, N4695, N6264, N2451);
xor XOR2 (N14134, N14127, N1896);
buf BUF1 (N14135, N14130);
and AND3 (N14136, N14129, N3201, N4104);
nor NOR3 (N14137, N14135, N806, N6991);
or OR2 (N14138, N14128, N11733);
nor NOR3 (N14139, N14124, N11777, N1264);
not NOT1 (N14140, N14138);
not NOT1 (N14141, N14140);
xor XOR2 (N14142, N14133, N10035);
buf BUF1 (N14143, N14126);
xor XOR2 (N14144, N14101, N10017);
xor XOR2 (N14145, N14134, N328);
not NOT1 (N14146, N14145);
and AND4 (N14147, N14146, N12065, N5721, N7399);
xor XOR2 (N14148, N14139, N3012);
nor NOR2 (N14149, N14142, N7700);
not NOT1 (N14150, N14149);
xor XOR2 (N14151, N14132, N9852);
nor NOR2 (N14152, N14143, N8357);
buf BUF1 (N14153, N14144);
or OR3 (N14154, N14137, N6740, N7490);
and AND3 (N14155, N14147, N12942, N11662);
nor NOR2 (N14156, N14141, N10917);
nor NOR4 (N14157, N14153, N12688, N2887, N6562);
or OR2 (N14158, N14136, N13914);
nor NOR2 (N14159, N14156, N10020);
nand NAND4 (N14160, N14150, N7896, N8659, N1418);
nor NOR2 (N14161, N14152, N4525);
not NOT1 (N14162, N14161);
nand NAND3 (N14163, N14151, N1523, N5189);
xor XOR2 (N14164, N14160, N6228);
nor NOR3 (N14165, N14157, N11888, N2826);
xor XOR2 (N14166, N14163, N1598);
or OR2 (N14167, N14131, N4656);
nor NOR3 (N14168, N14154, N10673, N1695);
and AND2 (N14169, N14168, N3554);
buf BUF1 (N14170, N14148);
buf BUF1 (N14171, N14169);
or OR4 (N14172, N14171, N709, N697, N243);
buf BUF1 (N14173, N14164);
nand NAND3 (N14174, N14166, N8622, N11864);
and AND2 (N14175, N14165, N9152);
buf BUF1 (N14176, N14174);
xor XOR2 (N14177, N14172, N13467);
buf BUF1 (N14178, N14167);
or OR2 (N14179, N14158, N10499);
nor NOR2 (N14180, N14177, N8437);
nor NOR2 (N14181, N14178, N14136);
buf BUF1 (N14182, N14176);
or OR3 (N14183, N14162, N3559, N4784);
or OR4 (N14184, N14181, N1788, N4012, N11965);
buf BUF1 (N14185, N14184);
nor NOR4 (N14186, N14173, N10497, N12359, N1963);
and AND2 (N14187, N14183, N898);
buf BUF1 (N14188, N14186);
or OR2 (N14189, N14179, N3610);
xor XOR2 (N14190, N14189, N10877);
or OR4 (N14191, N14190, N13983, N10033, N2676);
or OR3 (N14192, N14188, N8903, N4505);
xor XOR2 (N14193, N14187, N3620);
not NOT1 (N14194, N14155);
not NOT1 (N14195, N14194);
buf BUF1 (N14196, N14195);
xor XOR2 (N14197, N14182, N5622);
nor NOR4 (N14198, N14191, N9875, N11022, N9371);
or OR4 (N14199, N14170, N4151, N1188, N9593);
xor XOR2 (N14200, N14159, N11277);
nand NAND2 (N14201, N14180, N13906);
and AND4 (N14202, N14199, N13453, N4770, N10277);
or OR4 (N14203, N14193, N466, N8090, N13599);
xor XOR2 (N14204, N14197, N11407);
and AND3 (N14205, N14198, N9336, N5774);
not NOT1 (N14206, N14203);
not NOT1 (N14207, N14175);
nor NOR2 (N14208, N14196, N590);
and AND3 (N14209, N14207, N5733, N4444);
xor XOR2 (N14210, N14209, N261);
not NOT1 (N14211, N14185);
and AND2 (N14212, N14205, N9125);
not NOT1 (N14213, N14211);
and AND4 (N14214, N14210, N4849, N6709, N8499);
xor XOR2 (N14215, N14201, N6136);
buf BUF1 (N14216, N14208);
buf BUF1 (N14217, N14200);
xor XOR2 (N14218, N14204, N1890);
nor NOR4 (N14219, N14216, N10432, N2473, N7847);
nand NAND4 (N14220, N14202, N13518, N9818, N13613);
nand NAND2 (N14221, N14218, N6550);
nor NOR4 (N14222, N14215, N5838, N2024, N693);
or OR4 (N14223, N14213, N9968, N4433, N7848);
or OR2 (N14224, N14206, N2098);
xor XOR2 (N14225, N14219, N5135);
or OR2 (N14226, N14221, N9671);
xor XOR2 (N14227, N14226, N10883);
nor NOR3 (N14228, N14227, N6324, N3890);
or OR4 (N14229, N14214, N9623, N4799, N5425);
buf BUF1 (N14230, N14222);
not NOT1 (N14231, N14228);
nor NOR3 (N14232, N14229, N2237, N1060);
nor NOR4 (N14233, N14192, N7031, N9350, N13379);
or OR4 (N14234, N14224, N12557, N12746, N5291);
or OR2 (N14235, N14217, N6071);
and AND4 (N14236, N14212, N10917, N5094, N12684);
buf BUF1 (N14237, N14230);
or OR4 (N14238, N14232, N14183, N3461, N694);
buf BUF1 (N14239, N14238);
not NOT1 (N14240, N14220);
not NOT1 (N14241, N14225);
nand NAND2 (N14242, N14233, N119);
nand NAND2 (N14243, N14242, N2693);
and AND4 (N14244, N14240, N2209, N14153, N10228);
nand NAND2 (N14245, N14241, N4628);
and AND2 (N14246, N14243, N11517);
buf BUF1 (N14247, N14231);
buf BUF1 (N14248, N14244);
and AND3 (N14249, N14237, N5255, N1765);
xor XOR2 (N14250, N14234, N14244);
xor XOR2 (N14251, N14249, N1335);
nand NAND4 (N14252, N14250, N13596, N2804, N4968);
buf BUF1 (N14253, N14235);
xor XOR2 (N14254, N14223, N7504);
nand NAND4 (N14255, N14239, N1585, N9662, N5532);
buf BUF1 (N14256, N14246);
buf BUF1 (N14257, N14254);
and AND2 (N14258, N14248, N8477);
buf BUF1 (N14259, N14251);
or OR2 (N14260, N14258, N1628);
nor NOR4 (N14261, N14253, N10003, N6360, N11046);
and AND3 (N14262, N14255, N10086, N1968);
buf BUF1 (N14263, N14262);
xor XOR2 (N14264, N14252, N8380);
not NOT1 (N14265, N14259);
buf BUF1 (N14266, N14265);
not NOT1 (N14267, N14245);
not NOT1 (N14268, N14261);
nor NOR4 (N14269, N14236, N9155, N7816, N13145);
or OR3 (N14270, N14268, N1346, N14264);
and AND3 (N14271, N13597, N12179, N1813);
nand NAND2 (N14272, N14257, N9731);
buf BUF1 (N14273, N14272);
buf BUF1 (N14274, N14260);
and AND4 (N14275, N14271, N9136, N302, N4034);
nand NAND2 (N14276, N14275, N11317);
and AND4 (N14277, N14256, N9026, N12946, N11329);
or OR4 (N14278, N14276, N1691, N2135, N2296);
nand NAND2 (N14279, N14277, N6211);
buf BUF1 (N14280, N14270);
xor XOR2 (N14281, N14247, N9693);
not NOT1 (N14282, N14266);
nand NAND3 (N14283, N14281, N13417, N6269);
nor NOR2 (N14284, N14283, N10901);
not NOT1 (N14285, N14278);
buf BUF1 (N14286, N14263);
xor XOR2 (N14287, N14274, N5842);
nor NOR3 (N14288, N14285, N1034, N2285);
xor XOR2 (N14289, N14288, N14150);
buf BUF1 (N14290, N14269);
buf BUF1 (N14291, N14290);
nor NOR4 (N14292, N14273, N8740, N3868, N3300);
xor XOR2 (N14293, N14292, N11259);
nand NAND4 (N14294, N14291, N3526, N11841, N2872);
not NOT1 (N14295, N14280);
not NOT1 (N14296, N14295);
nand NAND3 (N14297, N14267, N753, N10788);
or OR3 (N14298, N14287, N3256, N6727);
buf BUF1 (N14299, N14284);
xor XOR2 (N14300, N14298, N7135);
nor NOR4 (N14301, N14289, N11643, N7946, N942);
buf BUF1 (N14302, N14294);
nand NAND2 (N14303, N14299, N618);
not NOT1 (N14304, N14303);
and AND3 (N14305, N14304, N7480, N2875);
not NOT1 (N14306, N14301);
and AND2 (N14307, N14286, N13935);
xor XOR2 (N14308, N14305, N4873);
nand NAND2 (N14309, N14282, N10295);
xor XOR2 (N14310, N14308, N9601);
nand NAND4 (N14311, N14309, N9906, N11438, N9276);
nor NOR2 (N14312, N14307, N8610);
nand NAND4 (N14313, N14297, N1155, N4893, N2417);
xor XOR2 (N14314, N14310, N13779);
nand NAND2 (N14315, N14293, N10608);
and AND3 (N14316, N14296, N3798, N5442);
or OR2 (N14317, N14302, N3502);
nand NAND3 (N14318, N14316, N1226, N4594);
nand NAND2 (N14319, N14318, N13368);
not NOT1 (N14320, N14279);
not NOT1 (N14321, N14312);
or OR2 (N14322, N14300, N9879);
xor XOR2 (N14323, N14311, N32);
or OR3 (N14324, N14322, N4101, N13641);
buf BUF1 (N14325, N14315);
xor XOR2 (N14326, N14313, N1092);
not NOT1 (N14327, N14317);
and AND4 (N14328, N14325, N11342, N1738, N8077);
and AND2 (N14329, N14314, N4979);
not NOT1 (N14330, N14321);
buf BUF1 (N14331, N14306);
nor NOR3 (N14332, N14326, N5035, N2891);
nand NAND2 (N14333, N14330, N5171);
nand NAND3 (N14334, N14327, N14229, N7176);
or OR2 (N14335, N14329, N4619);
nand NAND2 (N14336, N14332, N10725);
and AND3 (N14337, N14331, N7860, N4682);
nor NOR4 (N14338, N14319, N4219, N10887, N10169);
nor NOR4 (N14339, N14324, N4750, N7383, N1726);
not NOT1 (N14340, N14323);
or OR3 (N14341, N14338, N1978, N4574);
and AND4 (N14342, N14320, N5597, N9791, N12498);
or OR3 (N14343, N14341, N4758, N8071);
buf BUF1 (N14344, N14328);
or OR2 (N14345, N14342, N2805);
or OR4 (N14346, N14334, N12930, N8162, N10063);
buf BUF1 (N14347, N14340);
xor XOR2 (N14348, N14346, N14235);
or OR3 (N14349, N14347, N11410, N2344);
nand NAND2 (N14350, N14348, N4511);
xor XOR2 (N14351, N14337, N11039);
nor NOR2 (N14352, N14351, N8498);
or OR2 (N14353, N14339, N868);
nor NOR2 (N14354, N14349, N1575);
and AND2 (N14355, N14336, N5787);
xor XOR2 (N14356, N14335, N4247);
buf BUF1 (N14357, N14333);
not NOT1 (N14358, N14344);
not NOT1 (N14359, N14356);
xor XOR2 (N14360, N14357, N5469);
buf BUF1 (N14361, N14353);
not NOT1 (N14362, N14359);
or OR2 (N14363, N14362, N11077);
buf BUF1 (N14364, N14350);
and AND2 (N14365, N14363, N2932);
and AND4 (N14366, N14361, N7305, N2077, N9020);
and AND3 (N14367, N14366, N13803, N8614);
nand NAND2 (N14368, N14352, N11614);
and AND3 (N14369, N14355, N4877, N7920);
nand NAND2 (N14370, N14369, N13699);
nand NAND4 (N14371, N14365, N9726, N12619, N7777);
nand NAND2 (N14372, N14367, N13291);
nor NOR4 (N14373, N14372, N13621, N13360, N13545);
not NOT1 (N14374, N14345);
xor XOR2 (N14375, N14358, N3172);
not NOT1 (N14376, N14375);
nand NAND3 (N14377, N14368, N3607, N5150);
nor NOR3 (N14378, N14354, N4439, N3301);
nor NOR3 (N14379, N14373, N12212, N5020);
buf BUF1 (N14380, N14377);
nand NAND2 (N14381, N14379, N1984);
not NOT1 (N14382, N14370);
nand NAND3 (N14383, N14381, N9264, N4549);
nand NAND2 (N14384, N14364, N12230);
or OR3 (N14385, N14374, N7418, N1624);
buf BUF1 (N14386, N14383);
and AND4 (N14387, N14380, N599, N2736, N6606);
nand NAND4 (N14388, N14385, N13589, N623, N8397);
or OR2 (N14389, N14388, N13871);
nand NAND2 (N14390, N14343, N1779);
and AND4 (N14391, N14387, N1240, N9451, N3420);
nand NAND3 (N14392, N14384, N9052, N3764);
nand NAND3 (N14393, N14376, N7186, N12681);
not NOT1 (N14394, N14393);
nor NOR3 (N14395, N14390, N13424, N12042);
not NOT1 (N14396, N14392);
and AND3 (N14397, N14386, N3812, N11991);
nor NOR4 (N14398, N14397, N14093, N12768, N14294);
buf BUF1 (N14399, N14378);
nand NAND3 (N14400, N14382, N7038, N1009);
nand NAND3 (N14401, N14400, N3758, N6195);
or OR4 (N14402, N14371, N12309, N9045, N6436);
and AND2 (N14403, N14398, N10967);
xor XOR2 (N14404, N14391, N12227);
not NOT1 (N14405, N14395);
nand NAND2 (N14406, N14401, N5169);
and AND3 (N14407, N14360, N3863, N6658);
and AND3 (N14408, N14406, N1255, N9151);
nand NAND4 (N14409, N14404, N2889, N3163, N1819);
buf BUF1 (N14410, N14389);
not NOT1 (N14411, N14399);
and AND4 (N14412, N14396, N11245, N13921, N2946);
xor XOR2 (N14413, N14402, N12789);
or OR3 (N14414, N14394, N10671, N9985);
not NOT1 (N14415, N14413);
buf BUF1 (N14416, N14411);
buf BUF1 (N14417, N14416);
or OR4 (N14418, N14407, N7145, N7852, N11681);
xor XOR2 (N14419, N14409, N1039);
not NOT1 (N14420, N14417);
nor NOR3 (N14421, N14408, N13544, N4193);
nand NAND2 (N14422, N14419, N5182);
and AND3 (N14423, N14414, N11021, N12774);
and AND2 (N14424, N14422, N13165);
nor NOR3 (N14425, N14423, N13447, N2337);
and AND4 (N14426, N14403, N4256, N9656, N11172);
or OR2 (N14427, N14421, N7020);
nor NOR3 (N14428, N14424, N5633, N211);
nor NOR3 (N14429, N14415, N9680, N2558);
xor XOR2 (N14430, N14420, N9694);
xor XOR2 (N14431, N14430, N6247);
not NOT1 (N14432, N14427);
buf BUF1 (N14433, N14410);
xor XOR2 (N14434, N14429, N9228);
and AND2 (N14435, N14418, N10734);
buf BUF1 (N14436, N14435);
nand NAND3 (N14437, N14432, N9402, N3085);
nor NOR3 (N14438, N14436, N556, N2119);
buf BUF1 (N14439, N14428);
not NOT1 (N14440, N14431);
xor XOR2 (N14441, N14412, N12994);
buf BUF1 (N14442, N14405);
nor NOR4 (N14443, N14440, N5796, N11241, N6527);
buf BUF1 (N14444, N14434);
not NOT1 (N14445, N14425);
nand NAND3 (N14446, N14445, N7801, N7991);
nor NOR4 (N14447, N14426, N2354, N14104, N11492);
xor XOR2 (N14448, N14433, N2154);
not NOT1 (N14449, N14446);
nor NOR4 (N14450, N14441, N8872, N12092, N13162);
nand NAND2 (N14451, N14450, N12124);
xor XOR2 (N14452, N14447, N13264);
nand NAND4 (N14453, N14444, N11533, N2265, N9186);
nand NAND3 (N14454, N14439, N13932, N10719);
and AND2 (N14455, N14442, N13857);
xor XOR2 (N14456, N14451, N13641);
not NOT1 (N14457, N14438);
nor NOR4 (N14458, N14452, N2825, N6764, N12922);
buf BUF1 (N14459, N14449);
nor NOR2 (N14460, N14443, N8869);
nand NAND3 (N14461, N14460, N2700, N13109);
or OR3 (N14462, N14457, N2925, N3794);
nor NOR4 (N14463, N14456, N3343, N1600, N11131);
buf BUF1 (N14464, N14453);
not NOT1 (N14465, N14463);
or OR2 (N14466, N14461, N10631);
and AND2 (N14467, N14455, N1129);
nor NOR2 (N14468, N14464, N6186);
nand NAND2 (N14469, N14437, N3278);
xor XOR2 (N14470, N14468, N12175);
or OR3 (N14471, N14467, N13325, N9458);
or OR4 (N14472, N14448, N10780, N11966, N3494);
and AND2 (N14473, N14459, N1780);
or OR4 (N14474, N14470, N7640, N7131, N10446);
not NOT1 (N14475, N14472);
xor XOR2 (N14476, N14466, N3497);
not NOT1 (N14477, N14474);
and AND3 (N14478, N14454, N12686, N12206);
xor XOR2 (N14479, N14458, N8174);
not NOT1 (N14480, N14476);
nand NAND2 (N14481, N14465, N2169);
nor NOR3 (N14482, N14473, N10909, N2724);
nand NAND3 (N14483, N14475, N5735, N11765);
not NOT1 (N14484, N14477);
and AND3 (N14485, N14484, N6931, N9635);
nor NOR2 (N14486, N14469, N12170);
or OR4 (N14487, N14481, N12532, N4517, N13361);
or OR2 (N14488, N14487, N4078);
nand NAND4 (N14489, N14485, N12328, N10746, N871);
and AND3 (N14490, N14489, N3820, N11282);
or OR3 (N14491, N14479, N11422, N554);
nand NAND2 (N14492, N14483, N11823);
not NOT1 (N14493, N14490);
nor NOR2 (N14494, N14488, N5957);
not NOT1 (N14495, N14492);
and AND2 (N14496, N14493, N12939);
and AND4 (N14497, N14482, N13348, N6024, N2759);
nand NAND4 (N14498, N14496, N10467, N12421, N1928);
nor NOR2 (N14499, N14480, N10518);
nand NAND3 (N14500, N14462, N2685, N6815);
or OR2 (N14501, N14500, N13914);
xor XOR2 (N14502, N14486, N12161);
or OR4 (N14503, N14471, N8031, N1752, N11671);
nand NAND2 (N14504, N14503, N11823);
nand NAND2 (N14505, N14499, N12066);
buf BUF1 (N14506, N14501);
nor NOR3 (N14507, N14491, N4814, N8300);
not NOT1 (N14508, N14502);
and AND4 (N14509, N14504, N6443, N1509, N7199);
xor XOR2 (N14510, N14505, N10588);
nand NAND2 (N14511, N14478, N1333);
or OR3 (N14512, N14497, N4998, N5664);
and AND3 (N14513, N14509, N7733, N4036);
and AND4 (N14514, N14511, N4138, N12902, N6863);
and AND3 (N14515, N14508, N11344, N3233);
not NOT1 (N14516, N14513);
buf BUF1 (N14517, N14506);
or OR3 (N14518, N14495, N548, N11981);
buf BUF1 (N14519, N14516);
or OR3 (N14520, N14519, N8129, N12031);
nor NOR3 (N14521, N14510, N8288, N9043);
not NOT1 (N14522, N14494);
buf BUF1 (N14523, N14498);
nand NAND2 (N14524, N14520, N5268);
and AND4 (N14525, N14522, N1699, N6823, N2716);
not NOT1 (N14526, N14518);
buf BUF1 (N14527, N14507);
not NOT1 (N14528, N14515);
not NOT1 (N14529, N14514);
xor XOR2 (N14530, N14527, N13340);
nor NOR4 (N14531, N14523, N2126, N8149, N8235);
or OR2 (N14532, N14528, N9616);
not NOT1 (N14533, N14521);
xor XOR2 (N14534, N14530, N7196);
and AND3 (N14535, N14512, N4287, N8617);
nor NOR3 (N14536, N14517, N12925, N4349);
and AND3 (N14537, N14526, N10957, N14362);
xor XOR2 (N14538, N14537, N1254);
and AND4 (N14539, N14538, N10930, N10617, N6326);
buf BUF1 (N14540, N14531);
and AND3 (N14541, N14535, N4583, N12135);
not NOT1 (N14542, N14532);
or OR3 (N14543, N14533, N1025, N13994);
xor XOR2 (N14544, N14541, N7413);
xor XOR2 (N14545, N14534, N9250);
buf BUF1 (N14546, N14542);
nor NOR2 (N14547, N14536, N13306);
not NOT1 (N14548, N14547);
buf BUF1 (N14549, N14544);
nor NOR2 (N14550, N14546, N11982);
and AND2 (N14551, N14540, N5889);
not NOT1 (N14552, N14524);
and AND2 (N14553, N14550, N10720);
xor XOR2 (N14554, N14539, N6439);
buf BUF1 (N14555, N14548);
nand NAND3 (N14556, N14549, N4227, N7570);
xor XOR2 (N14557, N14529, N14188);
not NOT1 (N14558, N14557);
and AND3 (N14559, N14543, N12416, N9588);
or OR2 (N14560, N14555, N3522);
nand NAND2 (N14561, N14553, N4540);
nor NOR3 (N14562, N14556, N2911, N12863);
nand NAND3 (N14563, N14562, N8213, N11349);
xor XOR2 (N14564, N14558, N5945);
or OR4 (N14565, N14559, N9846, N4292, N1522);
nand NAND2 (N14566, N14552, N12028);
buf BUF1 (N14567, N14564);
buf BUF1 (N14568, N14554);
nor NOR3 (N14569, N14566, N4675, N12898);
xor XOR2 (N14570, N14560, N755);
nand NAND2 (N14571, N14569, N12560);
not NOT1 (N14572, N14525);
xor XOR2 (N14573, N14561, N3339);
not NOT1 (N14574, N14565);
or OR4 (N14575, N14573, N1222, N3558, N642);
not NOT1 (N14576, N14575);
buf BUF1 (N14577, N14571);
not NOT1 (N14578, N14551);
xor XOR2 (N14579, N14577, N14508);
buf BUF1 (N14580, N14578);
buf BUF1 (N14581, N14576);
nor NOR3 (N14582, N14563, N13390, N171);
xor XOR2 (N14583, N14568, N11511);
and AND4 (N14584, N14570, N3384, N10299, N953);
nor NOR4 (N14585, N14581, N3046, N11109, N14317);
buf BUF1 (N14586, N14580);
nor NOR4 (N14587, N14585, N12267, N3204, N2839);
xor XOR2 (N14588, N14545, N8219);
and AND3 (N14589, N14574, N1728, N2311);
or OR3 (N14590, N14579, N7799, N14459);
and AND4 (N14591, N14583, N5082, N10533, N8392);
nand NAND3 (N14592, N14567, N14361, N3192);
buf BUF1 (N14593, N14587);
or OR3 (N14594, N14589, N7739, N1884);
not NOT1 (N14595, N14594);
not NOT1 (N14596, N14584);
buf BUF1 (N14597, N14590);
not NOT1 (N14598, N14593);
not NOT1 (N14599, N14596);
nor NOR3 (N14600, N14586, N2500, N4560);
or OR3 (N14601, N14582, N11268, N14038);
nor NOR4 (N14602, N14599, N7303, N13020, N8233);
nand NAND4 (N14603, N14588, N11684, N3584, N14016);
or OR2 (N14604, N14572, N13573);
and AND3 (N14605, N14602, N11721, N1523);
and AND3 (N14606, N14603, N4914, N2250);
and AND4 (N14607, N14598, N3240, N13691, N12796);
or OR3 (N14608, N14606, N9189, N4321);
nor NOR3 (N14609, N14608, N1062, N3593);
nor NOR2 (N14610, N14605, N11793);
and AND4 (N14611, N14600, N8280, N11352, N14117);
xor XOR2 (N14612, N14607, N3905);
and AND2 (N14613, N14610, N7421);
buf BUF1 (N14614, N14591);
nand NAND4 (N14615, N14611, N12254, N7837, N6588);
buf BUF1 (N14616, N14612);
not NOT1 (N14617, N14609);
buf BUF1 (N14618, N14595);
buf BUF1 (N14619, N14617);
or OR3 (N14620, N14604, N3537, N10009);
xor XOR2 (N14621, N14597, N9843);
and AND2 (N14622, N14618, N6627);
buf BUF1 (N14623, N14614);
and AND2 (N14624, N14613, N8359);
or OR3 (N14625, N14615, N1318, N11503);
and AND4 (N14626, N14624, N9719, N12473, N6813);
not NOT1 (N14627, N14616);
xor XOR2 (N14628, N14619, N1442);
nor NOR4 (N14629, N14620, N4514, N8436, N1527);
not NOT1 (N14630, N14601);
buf BUF1 (N14631, N14592);
or OR3 (N14632, N14630, N14423, N10774);
nand NAND4 (N14633, N14623, N6659, N7454, N11116);
nand NAND2 (N14634, N14622, N3718);
xor XOR2 (N14635, N14632, N9974);
or OR4 (N14636, N14633, N3060, N10950, N5132);
xor XOR2 (N14637, N14631, N10104);
or OR4 (N14638, N14634, N4977, N8871, N2034);
and AND2 (N14639, N14628, N4058);
and AND2 (N14640, N14637, N6183);
or OR2 (N14641, N14625, N13336);
nand NAND4 (N14642, N14626, N3612, N11619, N14251);
nand NAND3 (N14643, N14621, N10676, N11503);
xor XOR2 (N14644, N14635, N12020);
and AND3 (N14645, N14644, N14013, N4290);
not NOT1 (N14646, N14638);
nor NOR2 (N14647, N14646, N3563);
nor NOR3 (N14648, N14639, N1014, N7248);
nand NAND2 (N14649, N14645, N5824);
nor NOR4 (N14650, N14636, N13755, N6679, N13633);
xor XOR2 (N14651, N14629, N3444);
xor XOR2 (N14652, N14643, N1764);
nand NAND2 (N14653, N14642, N13362);
xor XOR2 (N14654, N14650, N7904);
buf BUF1 (N14655, N14651);
xor XOR2 (N14656, N14655, N9400);
nand NAND4 (N14657, N14640, N14187, N7255, N13785);
nor NOR3 (N14658, N14648, N4633, N13264);
xor XOR2 (N14659, N14641, N11206);
nor NOR2 (N14660, N14652, N3201);
buf BUF1 (N14661, N14659);
and AND2 (N14662, N14627, N11342);
and AND4 (N14663, N14649, N3578, N11088, N12076);
nand NAND3 (N14664, N14657, N3792, N11631);
not NOT1 (N14665, N14660);
xor XOR2 (N14666, N14665, N10070);
nand NAND2 (N14667, N14653, N14313);
and AND4 (N14668, N14664, N2136, N10060, N11551);
nand NAND3 (N14669, N14668, N6115, N1025);
nor NOR3 (N14670, N14669, N783, N8722);
nand NAND3 (N14671, N14666, N6719, N2545);
not NOT1 (N14672, N14663);
and AND3 (N14673, N14658, N6844, N8832);
nor NOR2 (N14674, N14672, N12094);
and AND3 (N14675, N14670, N12915, N2536);
and AND2 (N14676, N14673, N4139);
or OR3 (N14677, N14675, N1266, N6222);
nand NAND2 (N14678, N14654, N3503);
xor XOR2 (N14679, N14671, N1460);
xor XOR2 (N14680, N14679, N13707);
nand NAND3 (N14681, N14647, N6881, N4300);
or OR4 (N14682, N14661, N14597, N13337, N10957);
not NOT1 (N14683, N14667);
not NOT1 (N14684, N14683);
buf BUF1 (N14685, N14656);
nor NOR3 (N14686, N14682, N1100, N14681);
buf BUF1 (N14687, N3343);
or OR2 (N14688, N14685, N3515);
and AND3 (N14689, N14686, N8842, N4540);
or OR3 (N14690, N14688, N12139, N11344);
buf BUF1 (N14691, N14680);
xor XOR2 (N14692, N14674, N3539);
buf BUF1 (N14693, N14676);
nor NOR2 (N14694, N14677, N7095);
nand NAND2 (N14695, N14693, N13799);
xor XOR2 (N14696, N14687, N948);
not NOT1 (N14697, N14678);
nor NOR3 (N14698, N14696, N2718, N476);
nand NAND2 (N14699, N14662, N14146);
nor NOR2 (N14700, N14684, N13650);
or OR4 (N14701, N14691, N3481, N5964, N1772);
nor NOR3 (N14702, N14701, N8286, N820);
buf BUF1 (N14703, N14700);
not NOT1 (N14704, N14695);
or OR3 (N14705, N14697, N9096, N6193);
buf BUF1 (N14706, N14689);
buf BUF1 (N14707, N14694);
and AND3 (N14708, N14706, N947, N12446);
nor NOR2 (N14709, N14705, N11879);
or OR4 (N14710, N14709, N7961, N2668, N4816);
or OR2 (N14711, N14707, N5693);
buf BUF1 (N14712, N14698);
nand NAND2 (N14713, N14710, N10693);
buf BUF1 (N14714, N14690);
or OR3 (N14715, N14708, N7927, N5348);
or OR4 (N14716, N14703, N2005, N8895, N1578);
not NOT1 (N14717, N14714);
xor XOR2 (N14718, N14704, N13373);
buf BUF1 (N14719, N14702);
and AND4 (N14720, N14713, N9537, N6074, N1697);
buf BUF1 (N14721, N14692);
buf BUF1 (N14722, N14716);
xor XOR2 (N14723, N14718, N10670);
or OR4 (N14724, N14722, N7294, N11437, N9416);
xor XOR2 (N14725, N14699, N12169);
or OR4 (N14726, N14715, N14543, N1845, N8900);
buf BUF1 (N14727, N14717);
or OR3 (N14728, N14727, N7220, N492);
or OR3 (N14729, N14719, N6538, N2273);
nand NAND4 (N14730, N14712, N947, N7359, N7180);
and AND4 (N14731, N14724, N8601, N6611, N1575);
or OR2 (N14732, N14723, N5737);
or OR2 (N14733, N14728, N4270);
buf BUF1 (N14734, N14730);
buf BUF1 (N14735, N14725);
nand NAND2 (N14736, N14733, N11053);
buf BUF1 (N14737, N14736);
and AND3 (N14738, N14729, N13553, N4361);
and AND2 (N14739, N14738, N2768);
nor NOR4 (N14740, N14731, N7648, N5794, N11390);
or OR3 (N14741, N14739, N3599, N14433);
nand NAND4 (N14742, N14737, N7843, N3286, N11633);
and AND4 (N14743, N14735, N10373, N13419, N1711);
and AND3 (N14744, N14732, N12938, N9121);
buf BUF1 (N14745, N14711);
nor NOR4 (N14746, N14744, N5194, N1568, N4802);
xor XOR2 (N14747, N14745, N10884);
or OR4 (N14748, N14743, N8529, N898, N5684);
not NOT1 (N14749, N14741);
not NOT1 (N14750, N14740);
buf BUF1 (N14751, N14721);
or OR2 (N14752, N14742, N12437);
and AND2 (N14753, N14749, N3321);
or OR3 (N14754, N14720, N14071, N4599);
nand NAND2 (N14755, N14726, N4172);
and AND3 (N14756, N14755, N5830, N9986);
nand NAND3 (N14757, N14747, N11340, N9809);
and AND3 (N14758, N14752, N5434, N9852);
nor NOR3 (N14759, N14748, N1854, N5943);
xor XOR2 (N14760, N14734, N2218);
nand NAND2 (N14761, N14754, N6361);
not NOT1 (N14762, N14750);
not NOT1 (N14763, N14758);
nand NAND3 (N14764, N14756, N8975, N8525);
not NOT1 (N14765, N14763);
or OR3 (N14766, N14765, N13310, N7051);
nand NAND4 (N14767, N14746, N1997, N8611, N14437);
and AND3 (N14768, N14764, N1708, N5474);
buf BUF1 (N14769, N14761);
and AND3 (N14770, N14757, N1367, N8513);
buf BUF1 (N14771, N14760);
nor NOR3 (N14772, N14770, N9273, N2585);
nand NAND3 (N14773, N14753, N5084, N14624);
nand NAND3 (N14774, N14769, N838, N7941);
or OR3 (N14775, N14774, N401, N5757);
nor NOR4 (N14776, N14773, N13518, N2192, N10528);
and AND2 (N14777, N14776, N8004);
not NOT1 (N14778, N14777);
buf BUF1 (N14779, N14768);
not NOT1 (N14780, N14771);
xor XOR2 (N14781, N14759, N13302);
not NOT1 (N14782, N14775);
xor XOR2 (N14783, N14778, N8965);
nor NOR2 (N14784, N14779, N9916);
nand NAND2 (N14785, N14766, N924);
not NOT1 (N14786, N14780);
xor XOR2 (N14787, N14784, N3398);
or OR2 (N14788, N14785, N12227);
or OR3 (N14789, N14751, N8863, N9096);
and AND2 (N14790, N14772, N6064);
not NOT1 (N14791, N14782);
xor XOR2 (N14792, N14789, N11190);
not NOT1 (N14793, N14787);
not NOT1 (N14794, N14783);
not NOT1 (N14795, N14767);
nand NAND2 (N14796, N14781, N12167);
not NOT1 (N14797, N14796);
not NOT1 (N14798, N14762);
xor XOR2 (N14799, N14792, N13843);
nor NOR2 (N14800, N14786, N6758);
or OR4 (N14801, N14798, N10486, N8103, N11083);
nand NAND4 (N14802, N14797, N12205, N12657, N7788);
or OR2 (N14803, N14793, N13170);
not NOT1 (N14804, N14794);
buf BUF1 (N14805, N14802);
not NOT1 (N14806, N14795);
xor XOR2 (N14807, N14791, N11326);
not NOT1 (N14808, N14801);
buf BUF1 (N14809, N14806);
not NOT1 (N14810, N14808);
and AND3 (N14811, N14810, N4554, N2411);
and AND3 (N14812, N14805, N11941, N3280);
nor NOR2 (N14813, N14800, N3511);
xor XOR2 (N14814, N14807, N3702);
not NOT1 (N14815, N14799);
buf BUF1 (N14816, N14811);
or OR2 (N14817, N14803, N10172);
nand NAND4 (N14818, N14812, N7181, N9267, N8910);
nor NOR3 (N14819, N14814, N8056, N14062);
or OR3 (N14820, N14818, N7358, N13391);
nor NOR2 (N14821, N14804, N3866);
and AND4 (N14822, N14815, N8121, N12484, N10025);
xor XOR2 (N14823, N14817, N8129);
or OR2 (N14824, N14813, N72);
and AND3 (N14825, N14821, N10804, N1192);
nor NOR4 (N14826, N14823, N8252, N10381, N7714);
buf BUF1 (N14827, N14820);
and AND3 (N14828, N14826, N2306, N5191);
not NOT1 (N14829, N14809);
nand NAND3 (N14830, N14829, N4620, N3465);
and AND4 (N14831, N14825, N1022, N13634, N5442);
nor NOR3 (N14832, N14827, N5344, N5327);
buf BUF1 (N14833, N14819);
or OR2 (N14834, N14831, N5037);
buf BUF1 (N14835, N14824);
nand NAND2 (N14836, N14822, N4594);
nor NOR2 (N14837, N14830, N1720);
nor NOR4 (N14838, N14790, N12814, N4927, N6693);
xor XOR2 (N14839, N14834, N10287);
and AND3 (N14840, N14833, N14470, N10689);
xor XOR2 (N14841, N14839, N7573);
buf BUF1 (N14842, N14838);
xor XOR2 (N14843, N14837, N725);
nor NOR2 (N14844, N14840, N5258);
nand NAND3 (N14845, N14841, N5093, N2962);
nand NAND3 (N14846, N14845, N2222, N6468);
or OR2 (N14847, N14842, N1185);
xor XOR2 (N14848, N14843, N14701);
nor NOR2 (N14849, N14828, N483);
nand NAND3 (N14850, N14848, N11826, N13123);
xor XOR2 (N14851, N14849, N8291);
nor NOR2 (N14852, N14846, N1509);
nor NOR4 (N14853, N14836, N9433, N11352, N10972);
and AND3 (N14854, N14835, N12366, N4657);
nor NOR3 (N14855, N14852, N7672, N13979);
nor NOR4 (N14856, N14855, N1068, N1337, N11730);
and AND3 (N14857, N14853, N6940, N9321);
or OR2 (N14858, N14847, N14281);
nand NAND4 (N14859, N14854, N234, N1997, N403);
and AND4 (N14860, N14832, N10068, N747, N11547);
or OR4 (N14861, N14788, N1134, N3890, N10893);
or OR2 (N14862, N14816, N10084);
nor NOR3 (N14863, N14862, N8947, N4052);
buf BUF1 (N14864, N14850);
and AND3 (N14865, N14851, N191, N14494);
xor XOR2 (N14866, N14865, N8324);
or OR2 (N14867, N14856, N5905);
buf BUF1 (N14868, N14866);
buf BUF1 (N14869, N14863);
buf BUF1 (N14870, N14869);
nor NOR3 (N14871, N14867, N2459, N13632);
xor XOR2 (N14872, N14857, N11799);
and AND4 (N14873, N14870, N4182, N1349, N10536);
not NOT1 (N14874, N14858);
xor XOR2 (N14875, N14874, N749);
not NOT1 (N14876, N14864);
not NOT1 (N14877, N14876);
nand NAND3 (N14878, N14871, N4577, N12018);
buf BUF1 (N14879, N14872);
xor XOR2 (N14880, N14875, N7909);
nor NOR2 (N14881, N14880, N901);
nor NOR2 (N14882, N14860, N8744);
nand NAND2 (N14883, N14844, N13392);
and AND3 (N14884, N14877, N8498, N11934);
not NOT1 (N14885, N14868);
not NOT1 (N14886, N14861);
buf BUF1 (N14887, N14859);
nand NAND4 (N14888, N14873, N6642, N994, N9004);
buf BUF1 (N14889, N14878);
and AND4 (N14890, N14886, N13687, N11779, N8593);
buf BUF1 (N14891, N14884);
nor NOR3 (N14892, N14890, N5444, N14609);
buf BUF1 (N14893, N14889);
or OR3 (N14894, N14893, N1415, N408);
buf BUF1 (N14895, N14887);
nor NOR2 (N14896, N14892, N6165);
or OR2 (N14897, N14895, N8136);
nor NOR2 (N14898, N14879, N12672);
nand NAND3 (N14899, N14888, N1824, N11525);
nor NOR2 (N14900, N14894, N2606);
nor NOR2 (N14901, N14897, N1039);
buf BUF1 (N14902, N14881);
nor NOR2 (N14903, N14896, N10218);
nand NAND3 (N14904, N14901, N4981, N6789);
nor NOR3 (N14905, N14891, N4727, N5503);
nand NAND3 (N14906, N14903, N10210, N9550);
buf BUF1 (N14907, N14906);
and AND3 (N14908, N14907, N8101, N13420);
or OR3 (N14909, N14904, N7979, N14821);
not NOT1 (N14910, N14899);
buf BUF1 (N14911, N14900);
xor XOR2 (N14912, N14898, N10535);
nor NOR2 (N14913, N14902, N4443);
nor NOR2 (N14914, N14883, N12117);
and AND3 (N14915, N14910, N7393, N828);
nand NAND4 (N14916, N14913, N12985, N7826, N10953);
nor NOR4 (N14917, N14909, N14257, N4279, N6875);
xor XOR2 (N14918, N14916, N5972);
or OR2 (N14919, N14885, N13000);
not NOT1 (N14920, N14911);
or OR3 (N14921, N14908, N11256, N10649);
xor XOR2 (N14922, N14915, N1966);
and AND2 (N14923, N14920, N2189);
xor XOR2 (N14924, N14923, N14569);
buf BUF1 (N14925, N14918);
buf BUF1 (N14926, N14914);
xor XOR2 (N14927, N14917, N10563);
nand NAND4 (N14928, N14921, N3548, N2294, N14253);
and AND3 (N14929, N14922, N7959, N11789);
or OR2 (N14930, N14912, N10616);
buf BUF1 (N14931, N14927);
and AND4 (N14932, N14919, N5557, N3967, N683);
and AND3 (N14933, N14905, N12103, N4039);
not NOT1 (N14934, N14933);
nand NAND3 (N14935, N14931, N14034, N1122);
buf BUF1 (N14936, N14929);
not NOT1 (N14937, N14926);
or OR3 (N14938, N14936, N13668, N3817);
not NOT1 (N14939, N14934);
buf BUF1 (N14940, N14939);
nand NAND2 (N14941, N14940, N3508);
not NOT1 (N14942, N14928);
and AND3 (N14943, N14942, N6425, N6129);
buf BUF1 (N14944, N14935);
buf BUF1 (N14945, N14925);
nor NOR2 (N14946, N14941, N5695);
and AND3 (N14947, N14944, N43, N4202);
nor NOR2 (N14948, N14938, N2211);
and AND3 (N14949, N14946, N7738, N119);
or OR3 (N14950, N14930, N13265, N9805);
nand NAND2 (N14951, N14949, N4276);
and AND4 (N14952, N14943, N3625, N6975, N9389);
not NOT1 (N14953, N14952);
not NOT1 (N14954, N14948);
nand NAND4 (N14955, N14945, N4030, N9078, N9487);
and AND4 (N14956, N14954, N986, N12925, N12487);
and AND4 (N14957, N14882, N7139, N9348, N6103);
or OR3 (N14958, N14950, N5572, N782);
and AND4 (N14959, N14924, N8674, N1451, N8919);
not NOT1 (N14960, N14932);
and AND4 (N14961, N14947, N14839, N653, N3200);
or OR2 (N14962, N14959, N12423);
nor NOR4 (N14963, N14951, N5554, N3124, N3673);
and AND2 (N14964, N14955, N13437);
nand NAND2 (N14965, N14937, N13225);
xor XOR2 (N14966, N14965, N13341);
buf BUF1 (N14967, N14956);
or OR3 (N14968, N14967, N8715, N3672);
nor NOR4 (N14969, N14968, N14668, N9397, N10041);
buf BUF1 (N14970, N14969);
nand NAND2 (N14971, N14961, N1289);
xor XOR2 (N14972, N14971, N13083);
nand NAND4 (N14973, N14963, N4027, N7770, N6501);
or OR2 (N14974, N14953, N7440);
xor XOR2 (N14975, N14962, N14311);
not NOT1 (N14976, N14975);
or OR2 (N14977, N14964, N3199);
nand NAND2 (N14978, N14972, N8291);
not NOT1 (N14979, N14958);
and AND2 (N14980, N14957, N9522);
not NOT1 (N14981, N14976);
and AND3 (N14982, N14970, N2510, N12972);
nor NOR4 (N14983, N14973, N8682, N5158, N5138);
buf BUF1 (N14984, N14982);
or OR2 (N14985, N14960, N11523);
xor XOR2 (N14986, N14984, N1651);
buf BUF1 (N14987, N14974);
nand NAND2 (N14988, N14979, N389);
xor XOR2 (N14989, N14988, N6112);
not NOT1 (N14990, N14980);
buf BUF1 (N14991, N14990);
or OR3 (N14992, N14989, N4670, N12750);
nand NAND2 (N14993, N14985, N97);
not NOT1 (N14994, N14977);
xor XOR2 (N14995, N14981, N13638);
and AND2 (N14996, N14978, N6295);
buf BUF1 (N14997, N14983);
or OR3 (N14998, N14996, N6843, N11042);
or OR4 (N14999, N14992, N6173, N4142, N13958);
not NOT1 (N15000, N14986);
or OR4 (N15001, N14987, N10803, N8493, N8763);
and AND4 (N15002, N14966, N5168, N7866, N7332);
nor NOR3 (N15003, N14991, N11645, N1372);
nand NAND4 (N15004, N14997, N4792, N13078, N8960);
not NOT1 (N15005, N15003);
xor XOR2 (N15006, N15004, N3250);
nor NOR3 (N15007, N14998, N1672, N1951);
nand NAND3 (N15008, N14995, N2380, N7798);
not NOT1 (N15009, N15007);
or OR2 (N15010, N14994, N1702);
and AND3 (N15011, N15002, N14147, N14218);
not NOT1 (N15012, N14993);
nand NAND4 (N15013, N15005, N12851, N1885, N4116);
nor NOR2 (N15014, N15010, N9922);
xor XOR2 (N15015, N15011, N6109);
buf BUF1 (N15016, N15014);
nand NAND2 (N15017, N15015, N5414);
or OR2 (N15018, N15016, N52);
xor XOR2 (N15019, N15017, N6335);
or OR2 (N15020, N15012, N9966);
or OR3 (N15021, N15019, N6863, N1458);
not NOT1 (N15022, N14999);
buf BUF1 (N15023, N15001);
nor NOR2 (N15024, N15008, N11029);
and AND2 (N15025, N15023, N3065);
or OR2 (N15026, N15025, N8990);
xor XOR2 (N15027, N15013, N11677);
nor NOR2 (N15028, N15006, N11184);
or OR4 (N15029, N15026, N3272, N3493, N446);
xor XOR2 (N15030, N15018, N3444);
or OR4 (N15031, N15030, N4620, N7369, N3453);
nand NAND4 (N15032, N15021, N5757, N5441, N14915);
buf BUF1 (N15033, N15022);
and AND2 (N15034, N15024, N3192);
xor XOR2 (N15035, N15020, N7475);
or OR2 (N15036, N15009, N9583);
nor NOR4 (N15037, N15029, N12028, N785, N4468);
nor NOR3 (N15038, N15031, N2040, N9565);
nand NAND3 (N15039, N15034, N5630, N2210);
or OR3 (N15040, N15036, N8358, N2191);
or OR2 (N15041, N15038, N14740);
nand NAND2 (N15042, N15037, N7495);
not NOT1 (N15043, N15028);
nand NAND2 (N15044, N15041, N9662);
and AND4 (N15045, N15043, N9821, N1870, N3639);
nor NOR3 (N15046, N15042, N10233, N13433);
and AND3 (N15047, N15040, N1967, N14961);
and AND4 (N15048, N15035, N4495, N12906, N13820);
nor NOR3 (N15049, N15039, N12804, N5368);
nor NOR3 (N15050, N15046, N11879, N10160);
buf BUF1 (N15051, N15000);
not NOT1 (N15052, N15033);
xor XOR2 (N15053, N15032, N6527);
buf BUF1 (N15054, N15051);
and AND2 (N15055, N15045, N87);
xor XOR2 (N15056, N15052, N6605);
or OR2 (N15057, N15055, N13802);
nand NAND3 (N15058, N15047, N12056, N10902);
not NOT1 (N15059, N15057);
or OR4 (N15060, N15058, N7610, N4896, N1169);
not NOT1 (N15061, N15050);
not NOT1 (N15062, N15054);
and AND4 (N15063, N15062, N2349, N3303, N11304);
not NOT1 (N15064, N15049);
buf BUF1 (N15065, N15048);
xor XOR2 (N15066, N15064, N7316);
buf BUF1 (N15067, N15027);
or OR2 (N15068, N15059, N14073);
and AND4 (N15069, N15067, N4356, N1716, N9423);
xor XOR2 (N15070, N15069, N13032);
buf BUF1 (N15071, N15056);
nand NAND2 (N15072, N15068, N12606);
xor XOR2 (N15073, N15071, N3113);
and AND4 (N15074, N15063, N11980, N10995, N6102);
and AND4 (N15075, N15061, N11507, N1863, N3674);
nor NOR2 (N15076, N15065, N9235);
nand NAND4 (N15077, N15072, N11234, N5077, N546);
or OR3 (N15078, N15070, N7019, N4218);
not NOT1 (N15079, N15073);
or OR2 (N15080, N15077, N4891);
and AND3 (N15081, N15060, N12545, N7939);
and AND4 (N15082, N15076, N5553, N12701, N8066);
and AND2 (N15083, N15082, N13968);
nor NOR4 (N15084, N15079, N6016, N8564, N4036);
nand NAND4 (N15085, N15084, N3910, N3379, N7782);
or OR4 (N15086, N15078, N13114, N9552, N14603);
and AND4 (N15087, N15066, N6161, N5830, N583);
nand NAND4 (N15088, N15087, N2189, N2176, N4686);
and AND3 (N15089, N15081, N2155, N14666);
nand NAND2 (N15090, N15085, N6278);
or OR2 (N15091, N15075, N6239);
and AND4 (N15092, N15088, N7346, N6441, N4491);
xor XOR2 (N15093, N15083, N5821);
or OR3 (N15094, N15089, N11019, N3164);
xor XOR2 (N15095, N15090, N9848);
buf BUF1 (N15096, N15044);
nand NAND4 (N15097, N15086, N11817, N3963, N9196);
buf BUF1 (N15098, N15094);
or OR2 (N15099, N15074, N14734);
buf BUF1 (N15100, N15095);
and AND3 (N15101, N15098, N1773, N6565);
nand NAND2 (N15102, N15100, N2686);
not NOT1 (N15103, N15096);
not NOT1 (N15104, N15091);
and AND4 (N15105, N15103, N1368, N2087, N12890);
buf BUF1 (N15106, N15105);
or OR2 (N15107, N15097, N12261);
or OR3 (N15108, N15092, N11610, N8952);
nand NAND4 (N15109, N15106, N6799, N231, N7893);
xor XOR2 (N15110, N15107, N4078);
xor XOR2 (N15111, N15108, N9438);
buf BUF1 (N15112, N15109);
nor NOR2 (N15113, N15053, N8229);
nor NOR2 (N15114, N15110, N14988);
or OR3 (N15115, N15080, N6419, N7909);
and AND2 (N15116, N15101, N7484);
nand NAND2 (N15117, N15112, N11937);
buf BUF1 (N15118, N15099);
and AND4 (N15119, N15111, N14076, N49, N2438);
xor XOR2 (N15120, N15118, N11410);
and AND3 (N15121, N15120, N11423, N3635);
nand NAND3 (N15122, N15115, N9182, N11131);
nand NAND4 (N15123, N15121, N14996, N6378, N8937);
nand NAND2 (N15124, N15114, N1549);
nor NOR4 (N15125, N15116, N8913, N14755, N14824);
buf BUF1 (N15126, N15102);
nor NOR2 (N15127, N15122, N1192);
xor XOR2 (N15128, N15113, N13195);
and AND2 (N15129, N15128, N5602);
and AND3 (N15130, N15119, N9541, N2731);
nand NAND3 (N15131, N15127, N9969, N10438);
xor XOR2 (N15132, N15130, N183);
nor NOR3 (N15133, N15131, N8916, N12728);
or OR3 (N15134, N15117, N2884, N4743);
nor NOR2 (N15135, N15132, N10331);
buf BUF1 (N15136, N15134);
nor NOR4 (N15137, N15125, N13456, N8521, N1161);
and AND4 (N15138, N15135, N4860, N1928, N14857);
buf BUF1 (N15139, N15104);
or OR4 (N15140, N15093, N5060, N4289, N13838);
or OR4 (N15141, N15126, N7579, N4245, N5584);
not NOT1 (N15142, N15137);
and AND2 (N15143, N15124, N14074);
xor XOR2 (N15144, N15136, N2560);
nor NOR4 (N15145, N15140, N1365, N7364, N12611);
buf BUF1 (N15146, N15139);
nor NOR4 (N15147, N15146, N14333, N5335, N8907);
and AND2 (N15148, N15129, N3740);
nand NAND2 (N15149, N15147, N12662);
and AND2 (N15150, N15141, N13682);
buf BUF1 (N15151, N15123);
nor NOR2 (N15152, N15145, N128);
buf BUF1 (N15153, N15151);
nand NAND3 (N15154, N15143, N9102, N4422);
xor XOR2 (N15155, N15142, N7843);
xor XOR2 (N15156, N15149, N5550);
buf BUF1 (N15157, N15152);
xor XOR2 (N15158, N15133, N1059);
xor XOR2 (N15159, N15157, N7156);
and AND3 (N15160, N15155, N11355, N9192);
or OR2 (N15161, N15148, N11171);
not NOT1 (N15162, N15161);
not NOT1 (N15163, N15144);
nand NAND3 (N15164, N15138, N10749, N14292);
or OR4 (N15165, N15164, N12812, N4886, N766);
and AND2 (N15166, N15156, N12131);
nor NOR3 (N15167, N15165, N5573, N11519);
buf BUF1 (N15168, N15166);
nand NAND2 (N15169, N15160, N1942);
xor XOR2 (N15170, N15154, N4335);
and AND2 (N15171, N15170, N3309);
and AND4 (N15172, N15163, N5443, N11589, N9099);
not NOT1 (N15173, N15162);
not NOT1 (N15174, N15171);
nand NAND3 (N15175, N15168, N9435, N14583);
nor NOR3 (N15176, N15150, N8149, N5533);
and AND2 (N15177, N15176, N10473);
buf BUF1 (N15178, N15177);
and AND2 (N15179, N15159, N3087);
nand NAND2 (N15180, N15179, N4471);
and AND2 (N15181, N15169, N14214);
or OR2 (N15182, N15174, N8030);
buf BUF1 (N15183, N15178);
and AND3 (N15184, N15153, N2083, N11303);
xor XOR2 (N15185, N15184, N4066);
and AND4 (N15186, N15158, N12476, N5390, N4916);
nor NOR4 (N15187, N15180, N4058, N2054, N11589);
xor XOR2 (N15188, N15173, N12996);
and AND2 (N15189, N15185, N13062);
and AND2 (N15190, N15187, N10506);
and AND2 (N15191, N15181, N1860);
nand NAND3 (N15192, N15182, N7492, N5595);
nand NAND2 (N15193, N15189, N14536);
not NOT1 (N15194, N15193);
buf BUF1 (N15195, N15188);
not NOT1 (N15196, N15190);
or OR4 (N15197, N15191, N7822, N14054, N8306);
xor XOR2 (N15198, N15192, N6390);
nand NAND4 (N15199, N15196, N1584, N8144, N5576);
not NOT1 (N15200, N15198);
nor NOR2 (N15201, N15200, N12551);
xor XOR2 (N15202, N15167, N1512);
nand NAND2 (N15203, N15186, N197);
nor NOR2 (N15204, N15203, N8583);
not NOT1 (N15205, N15201);
buf BUF1 (N15206, N15175);
and AND3 (N15207, N15197, N14578, N3130);
xor XOR2 (N15208, N15202, N7794);
and AND2 (N15209, N15194, N4703);
nor NOR2 (N15210, N15183, N6417);
and AND4 (N15211, N15208, N1609, N9101, N13765);
and AND2 (N15212, N15207, N5186);
nor NOR3 (N15213, N15172, N2394, N14292);
or OR4 (N15214, N15213, N4650, N2082, N7927);
not NOT1 (N15215, N15211);
and AND4 (N15216, N15212, N1091, N11964, N9014);
buf BUF1 (N15217, N15214);
buf BUF1 (N15218, N15195);
nand NAND3 (N15219, N15204, N7974, N14694);
and AND2 (N15220, N15219, N8176);
and AND2 (N15221, N15209, N14286);
nand NAND4 (N15222, N15199, N902, N2138, N6743);
nand NAND4 (N15223, N15221, N3805, N10186, N11784);
nor NOR3 (N15224, N15215, N6783, N13152);
and AND2 (N15225, N15223, N7081);
and AND4 (N15226, N15218, N6072, N5895, N11048);
and AND2 (N15227, N15216, N425);
nor NOR3 (N15228, N15220, N7271, N13288);
nand NAND4 (N15229, N15228, N2830, N9813, N2206);
not NOT1 (N15230, N15224);
not NOT1 (N15231, N15217);
xor XOR2 (N15232, N15229, N3179);
buf BUF1 (N15233, N15226);
not NOT1 (N15234, N15225);
nor NOR3 (N15235, N15205, N9205, N7092);
or OR3 (N15236, N15210, N1513, N14722);
buf BUF1 (N15237, N15230);
or OR4 (N15238, N15233, N6516, N1098, N3271);
nand NAND4 (N15239, N15231, N6343, N5167, N6949);
nor NOR4 (N15240, N15234, N12116, N11487, N7534);
buf BUF1 (N15241, N15238);
or OR4 (N15242, N15241, N11367, N3772, N4163);
nor NOR2 (N15243, N15232, N3454);
xor XOR2 (N15244, N15206, N12682);
xor XOR2 (N15245, N15244, N6347);
nor NOR4 (N15246, N15239, N1752, N12819, N5738);
nor NOR2 (N15247, N15235, N9008);
xor XOR2 (N15248, N15222, N9075);
not NOT1 (N15249, N15247);
xor XOR2 (N15250, N15248, N9912);
nor NOR2 (N15251, N15240, N4567);
xor XOR2 (N15252, N15237, N6659);
nand NAND2 (N15253, N15246, N647);
buf BUF1 (N15254, N15253);
nor NOR3 (N15255, N15249, N10668, N1122);
nand NAND3 (N15256, N15243, N13363, N8462);
xor XOR2 (N15257, N15242, N8431);
and AND3 (N15258, N15250, N4105, N6457);
nand NAND2 (N15259, N15252, N4212);
buf BUF1 (N15260, N15256);
xor XOR2 (N15261, N15251, N12894);
xor XOR2 (N15262, N15236, N4571);
xor XOR2 (N15263, N15262, N13490);
buf BUF1 (N15264, N15263);
and AND3 (N15265, N15257, N5913, N13526);
nand NAND4 (N15266, N15265, N14214, N3323, N11079);
not NOT1 (N15267, N15255);
nand NAND2 (N15268, N15227, N12092);
or OR2 (N15269, N15267, N1381);
not NOT1 (N15270, N15266);
buf BUF1 (N15271, N15258);
and AND4 (N15272, N15271, N8223, N10716, N2685);
nand NAND4 (N15273, N15259, N3320, N10443, N13589);
nor NOR4 (N15274, N15270, N1851, N201, N2864);
and AND2 (N15275, N15264, N531);
nand NAND2 (N15276, N15268, N13045);
buf BUF1 (N15277, N15276);
xor XOR2 (N15278, N15260, N11210);
xor XOR2 (N15279, N15261, N14360);
or OR3 (N15280, N15269, N13220, N7571);
not NOT1 (N15281, N15279);
and AND3 (N15282, N15274, N203, N8615);
nor NOR2 (N15283, N15273, N12799);
or OR4 (N15284, N15280, N117, N7087, N414);
buf BUF1 (N15285, N15282);
nor NOR4 (N15286, N15278, N7831, N6055, N3051);
not NOT1 (N15287, N15275);
nand NAND4 (N15288, N15287, N4036, N3381, N11383);
nor NOR2 (N15289, N15288, N9941);
xor XOR2 (N15290, N15285, N12399);
not NOT1 (N15291, N15245);
buf BUF1 (N15292, N15283);
or OR2 (N15293, N15281, N2324);
or OR4 (N15294, N15293, N7848, N13097, N2413);
buf BUF1 (N15295, N15254);
or OR2 (N15296, N15289, N4411);
buf BUF1 (N15297, N15291);
not NOT1 (N15298, N15296);
xor XOR2 (N15299, N15286, N4503);
and AND4 (N15300, N15294, N8066, N5168, N14320);
xor XOR2 (N15301, N15284, N2524);
xor XOR2 (N15302, N15292, N14884);
nand NAND2 (N15303, N15272, N9222);
buf BUF1 (N15304, N15277);
or OR4 (N15305, N15304, N5593, N14343, N2015);
and AND2 (N15306, N15300, N11972);
and AND3 (N15307, N15302, N1758, N2321);
and AND3 (N15308, N15298, N9651, N6934);
and AND3 (N15309, N15308, N12849, N14480);
buf BUF1 (N15310, N15307);
nand NAND3 (N15311, N15299, N3736, N4939);
nor NOR3 (N15312, N15301, N8409, N10074);
not NOT1 (N15313, N15290);
and AND4 (N15314, N15303, N7847, N14893, N3354);
xor XOR2 (N15315, N15305, N8800);
not NOT1 (N15316, N15310);
buf BUF1 (N15317, N15312);
not NOT1 (N15318, N15314);
buf BUF1 (N15319, N15318);
xor XOR2 (N15320, N15315, N9189);
not NOT1 (N15321, N15311);
nor NOR2 (N15322, N15295, N7599);
buf BUF1 (N15323, N15316);
nand NAND2 (N15324, N15317, N11405);
buf BUF1 (N15325, N15306);
not NOT1 (N15326, N15321);
xor XOR2 (N15327, N15322, N13681);
nor NOR3 (N15328, N15327, N7542, N6623);
and AND2 (N15329, N15309, N7685);
nor NOR4 (N15330, N15319, N12404, N6341, N12268);
xor XOR2 (N15331, N15329, N1369);
nor NOR3 (N15332, N15313, N9594, N2630);
not NOT1 (N15333, N15324);
not NOT1 (N15334, N15323);
not NOT1 (N15335, N15333);
buf BUF1 (N15336, N15320);
buf BUF1 (N15337, N15335);
not NOT1 (N15338, N15297);
nand NAND3 (N15339, N15330, N5642, N11417);
or OR4 (N15340, N15338, N13420, N13824, N8036);
or OR4 (N15341, N15326, N10276, N7597, N1116);
buf BUF1 (N15342, N15337);
not NOT1 (N15343, N15331);
buf BUF1 (N15344, N15328);
not NOT1 (N15345, N15341);
nor NOR4 (N15346, N15340, N7033, N3931, N11962);
buf BUF1 (N15347, N15345);
buf BUF1 (N15348, N15325);
or OR2 (N15349, N15332, N13576);
xor XOR2 (N15350, N15344, N4823);
not NOT1 (N15351, N15343);
not NOT1 (N15352, N15334);
buf BUF1 (N15353, N15349);
buf BUF1 (N15354, N15352);
not NOT1 (N15355, N15348);
buf BUF1 (N15356, N15350);
not NOT1 (N15357, N15356);
and AND2 (N15358, N15342, N8294);
nor NOR3 (N15359, N15354, N9230, N5377);
buf BUF1 (N15360, N15346);
not NOT1 (N15361, N15351);
nand NAND3 (N15362, N15360, N9838, N11479);
or OR4 (N15363, N15361, N15169, N4232, N44);
xor XOR2 (N15364, N15336, N9840);
or OR4 (N15365, N15364, N12914, N744, N11890);
buf BUF1 (N15366, N15355);
nand NAND3 (N15367, N15363, N1513, N3948);
xor XOR2 (N15368, N15347, N14225);
and AND4 (N15369, N15367, N14190, N839, N2047);
or OR4 (N15370, N15368, N9468, N7974, N15015);
nand NAND3 (N15371, N15339, N9896, N11607);
or OR3 (N15372, N15362, N7333, N3804);
not NOT1 (N15373, N15359);
buf BUF1 (N15374, N15372);
nand NAND3 (N15375, N15366, N14429, N12258);
or OR2 (N15376, N15374, N3065);
not NOT1 (N15377, N15370);
not NOT1 (N15378, N15377);
xor XOR2 (N15379, N15365, N9562);
or OR2 (N15380, N15379, N183);
nor NOR4 (N15381, N15380, N3069, N12150, N5068);
nand NAND3 (N15382, N15358, N12211, N8855);
xor XOR2 (N15383, N15382, N3619);
and AND3 (N15384, N15383, N5703, N8308);
buf BUF1 (N15385, N15371);
xor XOR2 (N15386, N15378, N6644);
xor XOR2 (N15387, N15357, N1072);
and AND4 (N15388, N15381, N6827, N2142, N13316);
xor XOR2 (N15389, N15353, N8992);
nor NOR4 (N15390, N15386, N12427, N7916, N13019);
nor NOR3 (N15391, N15389, N15308, N7723);
and AND3 (N15392, N15385, N13942, N2693);
not NOT1 (N15393, N15373);
nand NAND3 (N15394, N15375, N6321, N14916);
buf BUF1 (N15395, N15393);
and AND3 (N15396, N15384, N4845, N8824);
and AND4 (N15397, N15369, N15158, N8695, N13239);
xor XOR2 (N15398, N15391, N9246);
not NOT1 (N15399, N15394);
nor NOR4 (N15400, N15388, N12687, N13701, N2449);
xor XOR2 (N15401, N15395, N8006);
xor XOR2 (N15402, N15401, N14439);
nand NAND3 (N15403, N15376, N14671, N5838);
not NOT1 (N15404, N15399);
nand NAND2 (N15405, N15402, N11603);
or OR3 (N15406, N15390, N6550, N12112);
nor NOR4 (N15407, N15405, N203, N3621, N9625);
or OR2 (N15408, N15398, N15106);
buf BUF1 (N15409, N15397);
buf BUF1 (N15410, N15392);
buf BUF1 (N15411, N15406);
and AND2 (N15412, N15403, N8073);
nor NOR4 (N15413, N15412, N8170, N9112, N6784);
or OR2 (N15414, N15407, N9586);
nand NAND2 (N15415, N15414, N14891);
and AND3 (N15416, N15413, N3785, N8942);
nor NOR2 (N15417, N15387, N9987);
nand NAND3 (N15418, N15408, N1946, N12214);
and AND3 (N15419, N15410, N8813, N1748);
nor NOR2 (N15420, N15400, N2085);
and AND4 (N15421, N15404, N12156, N4903, N9904);
buf BUF1 (N15422, N15416);
xor XOR2 (N15423, N15396, N13294);
buf BUF1 (N15424, N15423);
nand NAND3 (N15425, N15415, N14933, N5728);
buf BUF1 (N15426, N15420);
or OR4 (N15427, N15425, N9141, N2714, N1742);
nor NOR3 (N15428, N15417, N266, N6705);
nor NOR3 (N15429, N15411, N13510, N431);
buf BUF1 (N15430, N15409);
xor XOR2 (N15431, N15430, N8978);
nand NAND4 (N15432, N15418, N12125, N5776, N10991);
not NOT1 (N15433, N15429);
nand NAND4 (N15434, N15422, N224, N14685, N10176);
xor XOR2 (N15435, N15419, N10595);
not NOT1 (N15436, N15431);
buf BUF1 (N15437, N15432);
not NOT1 (N15438, N15437);
and AND3 (N15439, N15434, N9179, N544);
buf BUF1 (N15440, N15439);
and AND4 (N15441, N15428, N12100, N12371, N221);
or OR2 (N15442, N15436, N8285);
or OR4 (N15443, N15427, N13772, N12297, N3232);
or OR4 (N15444, N15438, N8632, N9571, N9874);
nand NAND3 (N15445, N15433, N7863, N7491);
or OR4 (N15446, N15442, N13446, N12852, N13348);
and AND2 (N15447, N15440, N9085);
not NOT1 (N15448, N15446);
not NOT1 (N15449, N15426);
and AND4 (N15450, N15449, N10222, N7427, N11719);
not NOT1 (N15451, N15441);
nor NOR2 (N15452, N15444, N10174);
or OR4 (N15453, N15448, N12026, N2961, N5064);
nor NOR2 (N15454, N15435, N14149);
not NOT1 (N15455, N15452);
nand NAND3 (N15456, N15443, N6110, N5237);
buf BUF1 (N15457, N15447);
or OR3 (N15458, N15453, N13496, N7678);
nor NOR3 (N15459, N15457, N8744, N13814);
not NOT1 (N15460, N15450);
and AND2 (N15461, N15459, N10612);
or OR4 (N15462, N15421, N280, N14823, N11516);
buf BUF1 (N15463, N15455);
and AND2 (N15464, N15458, N9135);
or OR4 (N15465, N15464, N10205, N4496, N5069);
not NOT1 (N15466, N15463);
and AND4 (N15467, N15466, N13532, N9729, N6348);
xor XOR2 (N15468, N15424, N6755);
and AND3 (N15469, N15465, N12781, N13180);
xor XOR2 (N15470, N15456, N8934);
and AND3 (N15471, N15461, N9506, N7573);
not NOT1 (N15472, N15462);
not NOT1 (N15473, N15472);
or OR3 (N15474, N15471, N10095, N2455);
not NOT1 (N15475, N15470);
xor XOR2 (N15476, N15454, N2910);
nor NOR3 (N15477, N15468, N14379, N306);
not NOT1 (N15478, N15473);
not NOT1 (N15479, N15460);
nand NAND4 (N15480, N15479, N14123, N7232, N3229);
not NOT1 (N15481, N15451);
nor NOR3 (N15482, N15475, N7948, N7521);
xor XOR2 (N15483, N15467, N5064);
or OR3 (N15484, N15481, N15048, N6437);
nand NAND2 (N15485, N15477, N1475);
nor NOR4 (N15486, N15445, N11386, N2733, N15029);
or OR4 (N15487, N15480, N12611, N1083, N1230);
buf BUF1 (N15488, N15482);
not NOT1 (N15489, N15486);
buf BUF1 (N15490, N15487);
nor NOR3 (N15491, N15485, N12523, N88);
not NOT1 (N15492, N15483);
or OR4 (N15493, N15484, N12840, N11389, N7936);
and AND2 (N15494, N15469, N7859);
xor XOR2 (N15495, N15492, N796);
not NOT1 (N15496, N15490);
nand NAND3 (N15497, N15478, N7428, N11681);
not NOT1 (N15498, N15489);
not NOT1 (N15499, N15495);
and AND4 (N15500, N15491, N10108, N12495, N11);
nor NOR4 (N15501, N15488, N950, N12786, N6304);
or OR2 (N15502, N15501, N13411);
buf BUF1 (N15503, N15493);
or OR3 (N15504, N15476, N4000, N10977);
nor NOR4 (N15505, N15494, N14664, N8137, N1804);
nand NAND3 (N15506, N15496, N13435, N11636);
or OR4 (N15507, N15503, N1210, N13734, N9782);
and AND2 (N15508, N15474, N3002);
nand NAND2 (N15509, N15504, N9985);
xor XOR2 (N15510, N15507, N1789);
nand NAND3 (N15511, N15502, N11635, N8671);
buf BUF1 (N15512, N15500);
and AND2 (N15513, N15512, N10340);
nand NAND4 (N15514, N15509, N7570, N10539, N5824);
and AND3 (N15515, N15506, N15459, N7333);
buf BUF1 (N15516, N15511);
buf BUF1 (N15517, N15510);
not NOT1 (N15518, N15513);
not NOT1 (N15519, N15498);
nand NAND4 (N15520, N15515, N5271, N4438, N5388);
xor XOR2 (N15521, N15505, N9489);
not NOT1 (N15522, N15499);
nand NAND4 (N15523, N15521, N8727, N8521, N11715);
not NOT1 (N15524, N15517);
buf BUF1 (N15525, N15508);
buf BUF1 (N15526, N15497);
not NOT1 (N15527, N15523);
or OR3 (N15528, N15525, N7031, N12265);
nor NOR2 (N15529, N15527, N14949);
xor XOR2 (N15530, N15528, N562);
nor NOR2 (N15531, N15518, N8530);
and AND3 (N15532, N15526, N3363, N10120);
nor NOR3 (N15533, N15520, N3234, N5559);
not NOT1 (N15534, N15514);
xor XOR2 (N15535, N15516, N7078);
not NOT1 (N15536, N15532);
xor XOR2 (N15537, N15522, N7344);
nand NAND3 (N15538, N15535, N9689, N13577);
and AND4 (N15539, N15530, N9084, N11405, N7330);
nor NOR3 (N15540, N15529, N12, N13130);
xor XOR2 (N15541, N15519, N7914);
and AND2 (N15542, N15537, N2477);
nor NOR3 (N15543, N15539, N1937, N1543);
or OR2 (N15544, N15531, N3461);
and AND2 (N15545, N15533, N2000);
and AND2 (N15546, N15534, N10649);
not NOT1 (N15547, N15536);
nand NAND2 (N15548, N15545, N12717);
buf BUF1 (N15549, N15543);
or OR4 (N15550, N15544, N7524, N3057, N1924);
and AND3 (N15551, N15541, N15381, N1853);
not NOT1 (N15552, N15538);
nand NAND2 (N15553, N15548, N13900);
buf BUF1 (N15554, N15553);
xor XOR2 (N15555, N15551, N11911);
and AND2 (N15556, N15554, N3519);
nand NAND4 (N15557, N15540, N5300, N14357, N3066);
buf BUF1 (N15558, N15547);
buf BUF1 (N15559, N15552);
buf BUF1 (N15560, N15559);
or OR3 (N15561, N15560, N1142, N14245);
nand NAND4 (N15562, N15556, N8246, N10626, N7031);
not NOT1 (N15563, N15546);
xor XOR2 (N15564, N15563, N4842);
xor XOR2 (N15565, N15542, N8091);
not NOT1 (N15566, N15558);
buf BUF1 (N15567, N15564);
not NOT1 (N15568, N15566);
nor NOR4 (N15569, N15550, N3273, N1643, N11813);
or OR3 (N15570, N15524, N8207, N6569);
nor NOR4 (N15571, N15555, N1385, N8097, N7535);
or OR3 (N15572, N15569, N3128, N8916);
xor XOR2 (N15573, N15562, N15015);
buf BUF1 (N15574, N15572);
xor XOR2 (N15575, N15573, N13911);
and AND3 (N15576, N15568, N3134, N3025);
nor NOR2 (N15577, N15576, N1154);
or OR4 (N15578, N15549, N2008, N11852, N1032);
buf BUF1 (N15579, N15570);
and AND3 (N15580, N15574, N6612, N6809);
nor NOR3 (N15581, N15561, N8124, N1782);
nor NOR3 (N15582, N15567, N9360, N11513);
or OR2 (N15583, N15565, N7887);
buf BUF1 (N15584, N15578);
xor XOR2 (N15585, N15582, N11664);
and AND4 (N15586, N15577, N9780, N1760, N6255);
and AND2 (N15587, N15580, N11673);
and AND4 (N15588, N15587, N961, N15551, N3407);
or OR3 (N15589, N15586, N10477, N8226);
xor XOR2 (N15590, N15589, N3585);
and AND2 (N15591, N15585, N12515);
or OR2 (N15592, N15583, N11891);
and AND3 (N15593, N15575, N11868, N2348);
or OR4 (N15594, N15590, N10721, N6139, N13056);
and AND4 (N15595, N15594, N11457, N11915, N2460);
or OR3 (N15596, N15592, N4279, N12666);
nor NOR4 (N15597, N15591, N11088, N7070, N9483);
nand NAND3 (N15598, N15593, N4497, N10835);
xor XOR2 (N15599, N15557, N13255);
or OR2 (N15600, N15596, N8628);
not NOT1 (N15601, N15581);
and AND3 (N15602, N15588, N7211, N7543);
nor NOR3 (N15603, N15579, N9583, N4721);
and AND4 (N15604, N15600, N8702, N7907, N12660);
xor XOR2 (N15605, N15598, N4010);
and AND2 (N15606, N15571, N13466);
not NOT1 (N15607, N15584);
nand NAND4 (N15608, N15601, N6408, N659, N6766);
xor XOR2 (N15609, N15603, N13199);
nor NOR4 (N15610, N15595, N3633, N253, N3568);
xor XOR2 (N15611, N15599, N14809);
nor NOR2 (N15612, N15609, N5042);
and AND4 (N15613, N15606, N12533, N12507, N314);
buf BUF1 (N15614, N15611);
nor NOR3 (N15615, N15612, N4666, N12015);
and AND2 (N15616, N15602, N6673);
not NOT1 (N15617, N15597);
or OR4 (N15618, N15614, N1566, N11031, N1060);
and AND4 (N15619, N15605, N12423, N11697, N6682);
xor XOR2 (N15620, N15616, N15038);
not NOT1 (N15621, N15613);
nand NAND4 (N15622, N15617, N2373, N6765, N6760);
and AND3 (N15623, N15620, N14829, N1926);
and AND3 (N15624, N15618, N5525, N13713);
nand NAND2 (N15625, N15615, N1319);
and AND3 (N15626, N15607, N13278, N12211);
buf BUF1 (N15627, N15604);
nand NAND3 (N15628, N15627, N6418, N13348);
not NOT1 (N15629, N15626);
nand NAND3 (N15630, N15628, N14168, N4118);
nor NOR4 (N15631, N15625, N10941, N14529, N2584);
not NOT1 (N15632, N15608);
nor NOR3 (N15633, N15619, N10819, N3271);
not NOT1 (N15634, N15624);
nand NAND4 (N15635, N15610, N7128, N8771, N12683);
nor NOR4 (N15636, N15633, N12365, N13417, N6770);
or OR2 (N15637, N15621, N11896);
nor NOR3 (N15638, N15632, N316, N7629);
xor XOR2 (N15639, N15623, N9155);
xor XOR2 (N15640, N15638, N4535);
xor XOR2 (N15641, N15634, N14047);
nor NOR3 (N15642, N15636, N3388, N2430);
nor NOR4 (N15643, N15642, N8041, N4600, N9658);
and AND2 (N15644, N15641, N10459);
buf BUF1 (N15645, N15631);
nor NOR3 (N15646, N15635, N6929, N10167);
and AND2 (N15647, N15643, N2551);
nor NOR4 (N15648, N15622, N11194, N11832, N13467);
not NOT1 (N15649, N15646);
or OR2 (N15650, N15649, N15091);
buf BUF1 (N15651, N15650);
xor XOR2 (N15652, N15644, N14744);
and AND3 (N15653, N15637, N13668, N12217);
nor NOR3 (N15654, N15639, N12, N2014);
buf BUF1 (N15655, N15654);
not NOT1 (N15656, N15648);
or OR4 (N15657, N15652, N7551, N891, N768);
and AND2 (N15658, N15651, N14470);
not NOT1 (N15659, N15655);
nand NAND4 (N15660, N15658, N461, N5883, N9750);
nand NAND4 (N15661, N15657, N6662, N6994, N14950);
and AND2 (N15662, N15660, N6533);
not NOT1 (N15663, N15656);
not NOT1 (N15664, N15647);
xor XOR2 (N15665, N15629, N12529);
buf BUF1 (N15666, N15640);
not NOT1 (N15667, N15645);
not NOT1 (N15668, N15661);
nor NOR4 (N15669, N15664, N1586, N2601, N6243);
buf BUF1 (N15670, N15663);
or OR2 (N15671, N15653, N749);
not NOT1 (N15672, N15630);
not NOT1 (N15673, N15662);
xor XOR2 (N15674, N15665, N8863);
xor XOR2 (N15675, N15666, N11904);
not NOT1 (N15676, N15671);
nor NOR4 (N15677, N15674, N9787, N10859, N4484);
buf BUF1 (N15678, N15669);
nand NAND3 (N15679, N15675, N8249, N12124);
buf BUF1 (N15680, N15659);
not NOT1 (N15681, N15677);
not NOT1 (N15682, N15680);
xor XOR2 (N15683, N15681, N8412);
xor XOR2 (N15684, N15668, N983);
not NOT1 (N15685, N15679);
not NOT1 (N15686, N15684);
or OR2 (N15687, N15667, N12535);
or OR2 (N15688, N15686, N5964);
or OR3 (N15689, N15676, N10632, N657);
xor XOR2 (N15690, N15670, N13308);
and AND4 (N15691, N15687, N15159, N4161, N11833);
nor NOR4 (N15692, N15689, N5562, N3325, N8399);
buf BUF1 (N15693, N15692);
nand NAND4 (N15694, N15688, N2354, N166, N8625);
not NOT1 (N15695, N15678);
xor XOR2 (N15696, N15691, N10764);
nand NAND4 (N15697, N15695, N14464, N2765, N4815);
buf BUF1 (N15698, N15683);
and AND2 (N15699, N15696, N8155);
nand NAND2 (N15700, N15694, N6254);
and AND4 (N15701, N15697, N13395, N8544, N3809);
nor NOR3 (N15702, N15673, N7019, N5286);
not NOT1 (N15703, N15693);
not NOT1 (N15704, N15701);
xor XOR2 (N15705, N15690, N10537);
and AND2 (N15706, N15682, N9438);
or OR3 (N15707, N15706, N1, N1687);
xor XOR2 (N15708, N15705, N15097);
nand NAND2 (N15709, N15708, N8354);
buf BUF1 (N15710, N15700);
not NOT1 (N15711, N15710);
nor NOR2 (N15712, N15711, N2080);
and AND4 (N15713, N15709, N4721, N8046, N6768);
or OR2 (N15714, N15698, N10781);
nor NOR4 (N15715, N15704, N12049, N6622, N15140);
not NOT1 (N15716, N15714);
and AND2 (N15717, N15699, N5951);
not NOT1 (N15718, N15703);
or OR3 (N15719, N15718, N8112, N6282);
buf BUF1 (N15720, N15712);
buf BUF1 (N15721, N15685);
or OR4 (N15722, N15672, N7084, N15678, N9757);
nor NOR4 (N15723, N15721, N4012, N11021, N11110);
buf BUF1 (N15724, N15715);
nand NAND3 (N15725, N15707, N6110, N11870);
and AND4 (N15726, N15716, N11501, N7460, N288);
nor NOR4 (N15727, N15722, N7469, N14234, N11167);
not NOT1 (N15728, N15726);
or OR3 (N15729, N15717, N5483, N6652);
nor NOR2 (N15730, N15713, N1887);
or OR3 (N15731, N15724, N2288, N11373);
nor NOR2 (N15732, N15731, N3142);
or OR4 (N15733, N15732, N3496, N15502, N14534);
not NOT1 (N15734, N15727);
nor NOR3 (N15735, N15719, N9804, N6260);
not NOT1 (N15736, N15729);
nand NAND2 (N15737, N15734, N10249);
or OR2 (N15738, N15735, N4088);
nor NOR3 (N15739, N15728, N10510, N12067);
or OR4 (N15740, N15738, N5124, N15572, N11651);
buf BUF1 (N15741, N15736);
not NOT1 (N15742, N15730);
or OR3 (N15743, N15723, N5279, N11570);
nor NOR3 (N15744, N15737, N9795, N11091);
xor XOR2 (N15745, N15739, N4333);
buf BUF1 (N15746, N15743);
nor NOR2 (N15747, N15741, N1189);
nor NOR4 (N15748, N15746, N1930, N14435, N6888);
not NOT1 (N15749, N15742);
buf BUF1 (N15750, N15702);
or OR4 (N15751, N15740, N10355, N2779, N13797);
nand NAND2 (N15752, N15720, N4491);
xor XOR2 (N15753, N15748, N6312);
or OR3 (N15754, N15745, N2390, N13143);
buf BUF1 (N15755, N15733);
buf BUF1 (N15756, N15754);
buf BUF1 (N15757, N15751);
nand NAND3 (N15758, N15752, N405, N14178);
nand NAND2 (N15759, N15758, N7984);
buf BUF1 (N15760, N15744);
not NOT1 (N15761, N15749);
nor NOR4 (N15762, N15760, N5692, N4871, N15704);
nand NAND2 (N15763, N15756, N2527);
xor XOR2 (N15764, N15759, N10448);
buf BUF1 (N15765, N15757);
not NOT1 (N15766, N15761);
buf BUF1 (N15767, N15766);
nand NAND2 (N15768, N15725, N6099);
xor XOR2 (N15769, N15753, N5530);
buf BUF1 (N15770, N15769);
nand NAND2 (N15771, N15750, N13053);
and AND2 (N15772, N15765, N12988);
buf BUF1 (N15773, N15771);
buf BUF1 (N15774, N15755);
or OR4 (N15775, N15763, N4911, N2860, N13046);
or OR4 (N15776, N15772, N10232, N1013, N13301);
not NOT1 (N15777, N15773);
not NOT1 (N15778, N15762);
xor XOR2 (N15779, N15747, N1859);
or OR4 (N15780, N15770, N12942, N3209, N10365);
nor NOR4 (N15781, N15768, N7662, N7838, N6222);
and AND2 (N15782, N15775, N6673);
nor NOR4 (N15783, N15778, N373, N5696, N8171);
not NOT1 (N15784, N15776);
buf BUF1 (N15785, N15783);
or OR2 (N15786, N15774, N4380);
nand NAND2 (N15787, N15780, N2257);
nand NAND2 (N15788, N15784, N2589);
nor NOR2 (N15789, N15785, N13600);
not NOT1 (N15790, N15789);
or OR3 (N15791, N15767, N5965, N2563);
nand NAND4 (N15792, N15787, N1633, N10124, N5881);
nand NAND4 (N15793, N15790, N15214, N5412, N5358);
nor NOR2 (N15794, N15779, N5767);
or OR4 (N15795, N15791, N4662, N4363, N15674);
buf BUF1 (N15796, N15786);
and AND3 (N15797, N15795, N13217, N1674);
or OR3 (N15798, N15781, N15602, N4173);
nand NAND3 (N15799, N15796, N14899, N15368);
not NOT1 (N15800, N15798);
nand NAND2 (N15801, N15792, N11717);
xor XOR2 (N15802, N15777, N12723);
or OR4 (N15803, N15788, N8472, N13096, N12917);
or OR2 (N15804, N15800, N9080);
not NOT1 (N15805, N15793);
or OR3 (N15806, N15803, N5653, N7399);
nand NAND4 (N15807, N15802, N8976, N1337, N15535);
nand NAND4 (N15808, N15799, N957, N2731, N13918);
buf BUF1 (N15809, N15807);
nand NAND2 (N15810, N15805, N3442);
not NOT1 (N15811, N15809);
and AND2 (N15812, N15801, N2141);
or OR2 (N15813, N15782, N9705);
nor NOR3 (N15814, N15764, N7538, N15222);
nor NOR4 (N15815, N15811, N9647, N2317, N1802);
and AND2 (N15816, N15814, N5277);
nand NAND3 (N15817, N15812, N8044, N13247);
buf BUF1 (N15818, N15816);
and AND2 (N15819, N15815, N15149);
or OR2 (N15820, N15808, N2023);
or OR3 (N15821, N15813, N9181, N2493);
buf BUF1 (N15822, N15821);
buf BUF1 (N15823, N15794);
buf BUF1 (N15824, N15818);
or OR3 (N15825, N15822, N5467, N7284);
and AND4 (N15826, N15797, N10115, N13731, N15011);
nor NOR2 (N15827, N15817, N6065);
buf BUF1 (N15828, N15806);
nand NAND2 (N15829, N15823, N12608);
or OR2 (N15830, N15826, N15228);
nor NOR4 (N15831, N15830, N11461, N1601, N4976);
buf BUF1 (N15832, N15810);
buf BUF1 (N15833, N15827);
buf BUF1 (N15834, N15825);
xor XOR2 (N15835, N15829, N2416);
not NOT1 (N15836, N15804);
buf BUF1 (N15837, N15832);
nand NAND3 (N15838, N15831, N7458, N6502);
buf BUF1 (N15839, N15833);
or OR2 (N15840, N15820, N13059);
not NOT1 (N15841, N15836);
or OR2 (N15842, N15840, N8847);
not NOT1 (N15843, N15839);
buf BUF1 (N15844, N15819);
or OR2 (N15845, N15837, N14661);
xor XOR2 (N15846, N15835, N7720);
and AND2 (N15847, N15838, N879);
xor XOR2 (N15848, N15843, N2925);
and AND3 (N15849, N15841, N5162, N9122);
nand NAND2 (N15850, N15849, N5108);
xor XOR2 (N15851, N15844, N13460);
nor NOR2 (N15852, N15846, N9354);
and AND4 (N15853, N15824, N11346, N4164, N8634);
nand NAND4 (N15854, N15845, N5964, N9142, N6107);
nor NOR3 (N15855, N15852, N3946, N1019);
nand NAND4 (N15856, N15842, N10841, N3377, N7329);
nand NAND3 (N15857, N15847, N7316, N6365);
and AND2 (N15858, N15853, N6400);
xor XOR2 (N15859, N15858, N1303);
buf BUF1 (N15860, N15855);
buf BUF1 (N15861, N15834);
or OR4 (N15862, N15857, N1019, N4451, N14282);
nand NAND4 (N15863, N15862, N4522, N15406, N10444);
buf BUF1 (N15864, N15850);
nor NOR2 (N15865, N15861, N4360);
nor NOR4 (N15866, N15865, N12014, N13963, N3640);
and AND4 (N15867, N15864, N9580, N14706, N15322);
not NOT1 (N15868, N15828);
not NOT1 (N15869, N15856);
nand NAND3 (N15870, N15867, N11318, N3167);
not NOT1 (N15871, N15868);
xor XOR2 (N15872, N15866, N6699);
nand NAND3 (N15873, N15870, N8473, N14047);
and AND4 (N15874, N15873, N7898, N1313, N6727);
or OR4 (N15875, N15859, N1057, N6585, N14573);
xor XOR2 (N15876, N15875, N12015);
not NOT1 (N15877, N15860);
buf BUF1 (N15878, N15863);
nor NOR3 (N15879, N15874, N6150, N1432);
buf BUF1 (N15880, N15854);
not NOT1 (N15881, N15872);
nand NAND2 (N15882, N15881, N4076);
not NOT1 (N15883, N15882);
xor XOR2 (N15884, N15878, N13072);
or OR4 (N15885, N15869, N5311, N7274, N4997);
and AND4 (N15886, N15851, N13170, N1116, N6034);
nand NAND4 (N15887, N15885, N4153, N1074, N14774);
nor NOR3 (N15888, N15871, N11713, N9029);
nand NAND3 (N15889, N15887, N2293, N3367);
buf BUF1 (N15890, N15884);
not NOT1 (N15891, N15888);
or OR4 (N15892, N15879, N11748, N11369, N897);
or OR3 (N15893, N15880, N13070, N5276);
nor NOR3 (N15894, N15891, N4919, N5829);
xor XOR2 (N15895, N15877, N5369);
buf BUF1 (N15896, N15883);
not NOT1 (N15897, N15896);
xor XOR2 (N15898, N15895, N9322);
nor NOR3 (N15899, N15848, N4677, N6217);
not NOT1 (N15900, N15897);
and AND4 (N15901, N15899, N11682, N3152, N6732);
nand NAND4 (N15902, N15893, N7933, N13963, N6847);
xor XOR2 (N15903, N15890, N4509);
nand NAND4 (N15904, N15902, N748, N6830, N12275);
not NOT1 (N15905, N15898);
nor NOR4 (N15906, N15892, N15104, N14572, N14282);
xor XOR2 (N15907, N15886, N13881);
or OR4 (N15908, N15904, N6572, N5305, N14574);
buf BUF1 (N15909, N15906);
and AND3 (N15910, N15900, N5400, N114);
xor XOR2 (N15911, N15905, N14078);
nand NAND4 (N15912, N15907, N11811, N11531, N11210);
and AND4 (N15913, N15894, N1809, N8941, N13706);
and AND4 (N15914, N15901, N6577, N4826, N15470);
not NOT1 (N15915, N15908);
nor NOR2 (N15916, N15909, N6512);
not NOT1 (N15917, N15876);
or OR3 (N15918, N15914, N9099, N2963);
nor NOR2 (N15919, N15918, N11116);
or OR2 (N15920, N15912, N7868);
nand NAND4 (N15921, N15917, N8021, N12733, N12816);
xor XOR2 (N15922, N15889, N1519);
xor XOR2 (N15923, N15919, N3582);
not NOT1 (N15924, N15922);
nand NAND4 (N15925, N15923, N15417, N9650, N11364);
or OR4 (N15926, N15916, N5482, N13919, N7568);
nor NOR2 (N15927, N15921, N8865);
buf BUF1 (N15928, N15903);
nand NAND4 (N15929, N15915, N2089, N8890, N14672);
or OR4 (N15930, N15927, N8349, N9625, N5123);
or OR3 (N15931, N15920, N6282, N11236);
buf BUF1 (N15932, N15911);
not NOT1 (N15933, N15929);
not NOT1 (N15934, N15910);
buf BUF1 (N15935, N15924);
nor NOR4 (N15936, N15913, N14717, N13858, N11064);
xor XOR2 (N15937, N15931, N8210);
or OR4 (N15938, N15934, N10172, N196, N14694);
nand NAND4 (N15939, N15933, N840, N14212, N5949);
buf BUF1 (N15940, N15935);
and AND4 (N15941, N15928, N9819, N8997, N12904);
nor NOR4 (N15942, N15936, N11753, N15562, N10891);
nand NAND2 (N15943, N15939, N781);
nand NAND3 (N15944, N15926, N8129, N1223);
or OR2 (N15945, N15932, N1259);
buf BUF1 (N15946, N15937);
buf BUF1 (N15947, N15925);
or OR4 (N15948, N15938, N7796, N9016, N5314);
nand NAND4 (N15949, N15942, N3554, N3836, N6137);
nor NOR4 (N15950, N15949, N8860, N6625, N2077);
buf BUF1 (N15951, N15950);
or OR2 (N15952, N15946, N5942);
xor XOR2 (N15953, N15945, N12495);
nor NOR3 (N15954, N15944, N8506, N11667);
xor XOR2 (N15955, N15953, N8367);
nand NAND2 (N15956, N15955, N5840);
not NOT1 (N15957, N15943);
and AND3 (N15958, N15951, N12277, N14152);
xor XOR2 (N15959, N15957, N6754);
xor XOR2 (N15960, N15959, N14612);
buf BUF1 (N15961, N15947);
nor NOR2 (N15962, N15941, N15079);
or OR2 (N15963, N15956, N6487);
nand NAND2 (N15964, N15960, N4462);
and AND4 (N15965, N15930, N2426, N15548, N15956);
not NOT1 (N15966, N15958);
buf BUF1 (N15967, N15962);
nand NAND2 (N15968, N15965, N10424);
or OR2 (N15969, N15967, N4835);
nand NAND4 (N15970, N15969, N9557, N9575, N9193);
nor NOR3 (N15971, N15966, N12612, N5262);
not NOT1 (N15972, N15968);
or OR2 (N15973, N15964, N4590);
nor NOR2 (N15974, N15973, N813);
not NOT1 (N15975, N15971);
buf BUF1 (N15976, N15948);
or OR4 (N15977, N15976, N706, N14783, N4854);
not NOT1 (N15978, N15940);
nor NOR3 (N15979, N15975, N12050, N3161);
nand NAND3 (N15980, N15977, N13027, N7251);
xor XOR2 (N15981, N15980, N8541);
buf BUF1 (N15982, N15961);
nor NOR2 (N15983, N15979, N3143);
xor XOR2 (N15984, N15972, N6608);
nand NAND3 (N15985, N15984, N3990, N11476);
xor XOR2 (N15986, N15974, N3249);
and AND4 (N15987, N15981, N10083, N8887, N3485);
nor NOR4 (N15988, N15987, N1819, N2191, N5851);
xor XOR2 (N15989, N15986, N3445);
nor NOR2 (N15990, N15970, N7516);
nand NAND4 (N15991, N15963, N426, N6484, N9553);
or OR2 (N15992, N15982, N6148);
xor XOR2 (N15993, N15992, N5831);
xor XOR2 (N15994, N15983, N15984);
xor XOR2 (N15995, N15954, N4881);
xor XOR2 (N15996, N15995, N1143);
nand NAND4 (N15997, N15985, N12990, N13559, N10097);
nor NOR2 (N15998, N15988, N5172);
or OR2 (N15999, N15993, N3817);
or OR4 (N16000, N15996, N6299, N14635, N5627);
and AND2 (N16001, N15991, N8611);
nor NOR2 (N16002, N15952, N15820);
or OR4 (N16003, N15990, N14217, N1889, N1451);
nor NOR3 (N16004, N16002, N345, N10761);
buf BUF1 (N16005, N15998);
and AND3 (N16006, N16005, N10103, N15516);
xor XOR2 (N16007, N15978, N6950);
or OR2 (N16008, N16007, N9278);
buf BUF1 (N16009, N15997);
nand NAND4 (N16010, N16004, N3965, N5591, N1798);
nor NOR2 (N16011, N16000, N6052);
xor XOR2 (N16012, N16009, N6609);
not NOT1 (N16013, N15999);
nand NAND3 (N16014, N16010, N12882, N11105);
not NOT1 (N16015, N16001);
and AND3 (N16016, N16003, N15900, N12987);
or OR4 (N16017, N16006, N6144, N4246, N11806);
and AND4 (N16018, N16013, N11367, N11129, N1409);
buf BUF1 (N16019, N16008);
or OR4 (N16020, N16014, N2803, N7172, N9938);
not NOT1 (N16021, N16018);
xor XOR2 (N16022, N16015, N6128);
endmodule