// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22;

output N1508,N1516,N1489,N1517,N1518,N1515,N1521,N1488,N1520,N1522;

buf BUF1 (N23, N5);
or OR4 (N24, N8, N3, N6, N7);
nand NAND3 (N25, N7, N8, N15);
buf BUF1 (N26, N22);
and AND4 (N27, N5, N10, N23, N21);
or OR4 (N28, N27, N1, N11, N27);
nor NOR4 (N29, N8, N14, N23, N5);
or OR2 (N30, N11, N17);
and AND2 (N31, N16, N11);
xor XOR2 (N32, N11, N29);
buf BUF1 (N33, N9);
not NOT1 (N34, N21);
buf BUF1 (N35, N34);
nand NAND4 (N36, N34, N22, N14, N26);
or OR2 (N37, N21, N11);
or OR2 (N38, N32, N1);
nand NAND2 (N39, N35, N21);
or OR2 (N40, N28, N18);
and AND4 (N41, N31, N38, N16, N24);
nor NOR3 (N42, N25, N8, N21);
nand NAND2 (N43, N19, N1);
not NOT1 (N44, N26);
or OR2 (N45, N42, N1);
xor XOR2 (N46, N36, N2);
nand NAND4 (N47, N43, N1, N37, N2);
buf BUF1 (N48, N38);
not NOT1 (N49, N41);
buf BUF1 (N50, N49);
or OR2 (N51, N48, N26);
nand NAND4 (N52, N47, N16, N25, N12);
not NOT1 (N53, N50);
buf BUF1 (N54, N46);
or OR2 (N55, N44, N8);
or OR2 (N56, N55, N24);
not NOT1 (N57, N52);
buf BUF1 (N58, N51);
buf BUF1 (N59, N45);
buf BUF1 (N60, N57);
or OR2 (N61, N30, N51);
not NOT1 (N62, N59);
xor XOR2 (N63, N62, N15);
not NOT1 (N64, N60);
or OR3 (N65, N56, N51, N7);
and AND4 (N66, N65, N47, N17, N18);
buf BUF1 (N67, N54);
nor NOR2 (N68, N66, N19);
nor NOR3 (N69, N58, N16, N22);
and AND3 (N70, N33, N56, N32);
xor XOR2 (N71, N64, N70);
or OR2 (N72, N56, N70);
not NOT1 (N73, N63);
nand NAND3 (N74, N69, N52, N41);
buf BUF1 (N75, N72);
xor XOR2 (N76, N67, N43);
xor XOR2 (N77, N75, N60);
not NOT1 (N78, N77);
not NOT1 (N79, N40);
and AND2 (N80, N74, N46);
or OR2 (N81, N68, N26);
not NOT1 (N82, N78);
or OR4 (N83, N79, N70, N61, N18);
nor NOR2 (N84, N36, N13);
and AND2 (N85, N83, N79);
not NOT1 (N86, N85);
nand NAND3 (N87, N84, N23, N4);
xor XOR2 (N88, N86, N46);
or OR4 (N89, N71, N44, N36, N58);
xor XOR2 (N90, N89, N88);
and AND2 (N91, N29, N8);
and AND2 (N92, N39, N45);
buf BUF1 (N93, N73);
and AND2 (N94, N91, N83);
buf BUF1 (N95, N80);
not NOT1 (N96, N90);
or OR4 (N97, N95, N45, N38, N66);
nand NAND3 (N98, N93, N36, N69);
and AND4 (N99, N81, N60, N18, N39);
and AND3 (N100, N96, N14, N9);
or OR2 (N101, N97, N55);
or OR2 (N102, N92, N87);
xor XOR2 (N103, N54, N58);
or OR4 (N104, N82, N32, N36, N29);
buf BUF1 (N105, N76);
not NOT1 (N106, N104);
or OR2 (N107, N103, N29);
not NOT1 (N108, N107);
not NOT1 (N109, N101);
not NOT1 (N110, N100);
xor XOR2 (N111, N94, N83);
not NOT1 (N112, N110);
nor NOR2 (N113, N109, N27);
xor XOR2 (N114, N106, N7);
nor NOR2 (N115, N99, N18);
not NOT1 (N116, N112);
xor XOR2 (N117, N53, N30);
not NOT1 (N118, N115);
nor NOR3 (N119, N118, N110, N63);
xor XOR2 (N120, N108, N81);
nor NOR2 (N121, N105, N10);
nor NOR2 (N122, N111, N65);
not NOT1 (N123, N113);
or OR4 (N124, N98, N25, N120, N4);
and AND3 (N125, N82, N109, N88);
buf BUF1 (N126, N117);
buf BUF1 (N127, N116);
not NOT1 (N128, N124);
and AND2 (N129, N125, N95);
nor NOR2 (N130, N119, N63);
xor XOR2 (N131, N128, N88);
nand NAND3 (N132, N127, N71, N84);
xor XOR2 (N133, N129, N78);
buf BUF1 (N134, N126);
nor NOR4 (N135, N114, N107, N31, N98);
nand NAND2 (N136, N135, N92);
nor NOR4 (N137, N102, N35, N128, N25);
buf BUF1 (N138, N131);
not NOT1 (N139, N130);
xor XOR2 (N140, N137, N74);
nor NOR3 (N141, N140, N67, N46);
buf BUF1 (N142, N139);
nand NAND4 (N143, N122, N48, N51, N38);
xor XOR2 (N144, N132, N114);
not NOT1 (N145, N142);
and AND3 (N146, N138, N67, N87);
or OR3 (N147, N144, N10, N95);
or OR4 (N148, N123, N56, N21, N87);
or OR2 (N149, N141, N109);
and AND4 (N150, N134, N20, N93, N117);
and AND4 (N151, N146, N6, N88, N128);
nor NOR2 (N152, N136, N126);
or OR4 (N153, N152, N17, N124, N57);
or OR4 (N154, N151, N3, N50, N149);
and AND3 (N155, N124, N113, N143);
and AND4 (N156, N35, N114, N62, N143);
or OR2 (N157, N150, N144);
not NOT1 (N158, N121);
buf BUF1 (N159, N158);
not NOT1 (N160, N157);
not NOT1 (N161, N159);
xor XOR2 (N162, N133, N52);
or OR4 (N163, N161, N31, N134, N3);
nor NOR2 (N164, N160, N153);
not NOT1 (N165, N111);
xor XOR2 (N166, N154, N69);
not NOT1 (N167, N148);
buf BUF1 (N168, N165);
not NOT1 (N169, N167);
or OR3 (N170, N145, N126, N8);
nor NOR4 (N171, N156, N117, N53, N79);
buf BUF1 (N172, N155);
not NOT1 (N173, N166);
nor NOR3 (N174, N173, N86, N116);
nand NAND2 (N175, N169, N100);
xor XOR2 (N176, N164, N94);
or OR3 (N177, N176, N72, N39);
and AND2 (N178, N171, N26);
xor XOR2 (N179, N172, N49);
buf BUF1 (N180, N177);
buf BUF1 (N181, N180);
nand NAND2 (N182, N163, N158);
or OR4 (N183, N178, N179, N32, N39);
buf BUF1 (N184, N106);
not NOT1 (N185, N162);
not NOT1 (N186, N168);
and AND3 (N187, N183, N60, N179);
nor NOR2 (N188, N184, N37);
xor XOR2 (N189, N187, N124);
not NOT1 (N190, N188);
xor XOR2 (N191, N189, N103);
or OR2 (N192, N175, N73);
buf BUF1 (N193, N191);
buf BUF1 (N194, N174);
and AND2 (N195, N185, N163);
nand NAND2 (N196, N192, N117);
xor XOR2 (N197, N170, N52);
nor NOR4 (N198, N181, N106, N109, N81);
or OR3 (N199, N195, N9, N111);
not NOT1 (N200, N186);
not NOT1 (N201, N200);
xor XOR2 (N202, N147, N165);
not NOT1 (N203, N201);
not NOT1 (N204, N194);
nor NOR3 (N205, N204, N10, N115);
buf BUF1 (N206, N203);
not NOT1 (N207, N198);
nor NOR2 (N208, N205, N34);
xor XOR2 (N209, N202, N123);
nor NOR4 (N210, N197, N30, N206, N177);
buf BUF1 (N211, N170);
nor NOR3 (N212, N190, N27, N52);
or OR2 (N213, N209, N9);
xor XOR2 (N214, N182, N12);
and AND3 (N215, N212, N148, N124);
and AND3 (N216, N207, N211, N207);
nor NOR2 (N217, N84, N150);
and AND2 (N218, N214, N1);
or OR4 (N219, N218, N111, N115, N139);
xor XOR2 (N220, N210, N81);
or OR2 (N221, N219, N164);
nor NOR4 (N222, N217, N93, N21, N71);
nor NOR2 (N223, N208, N208);
nand NAND2 (N224, N216, N169);
nor NOR3 (N225, N220, N127, N175);
nand NAND2 (N226, N222, N154);
buf BUF1 (N227, N193);
nand NAND3 (N228, N215, N120, N29);
and AND3 (N229, N223, N39, N160);
or OR2 (N230, N196, N11);
nor NOR3 (N231, N199, N31, N207);
nor NOR4 (N232, N225, N117, N101, N101);
and AND2 (N233, N213, N51);
and AND2 (N234, N228, N221);
nor NOR4 (N235, N78, N171, N41, N232);
and AND2 (N236, N31, N54);
or OR3 (N237, N234, N131, N34);
or OR2 (N238, N229, N142);
not NOT1 (N239, N227);
buf BUF1 (N240, N237);
buf BUF1 (N241, N235);
not NOT1 (N242, N241);
not NOT1 (N243, N242);
or OR4 (N244, N230, N137, N75, N52);
or OR3 (N245, N236, N234, N202);
nand NAND3 (N246, N233, N216, N57);
buf BUF1 (N247, N238);
or OR3 (N248, N247, N114, N1);
buf BUF1 (N249, N226);
xor XOR2 (N250, N240, N203);
nand NAND4 (N251, N249, N189, N55, N37);
nor NOR4 (N252, N239, N220, N155, N232);
and AND4 (N253, N252, N56, N58, N144);
buf BUF1 (N254, N248);
not NOT1 (N255, N254);
buf BUF1 (N256, N244);
buf BUF1 (N257, N243);
or OR3 (N258, N251, N129, N107);
or OR3 (N259, N245, N229, N26);
and AND2 (N260, N255, N65);
buf BUF1 (N261, N253);
buf BUF1 (N262, N257);
not NOT1 (N263, N224);
xor XOR2 (N264, N246, N67);
buf BUF1 (N265, N261);
buf BUF1 (N266, N264);
nor NOR2 (N267, N231, N103);
nor NOR3 (N268, N263, N196, N88);
not NOT1 (N269, N250);
or OR3 (N270, N256, N138, N153);
buf BUF1 (N271, N266);
buf BUF1 (N272, N267);
or OR4 (N273, N258, N133, N148, N177);
not NOT1 (N274, N268);
buf BUF1 (N275, N262);
and AND2 (N276, N275, N207);
nor NOR2 (N277, N259, N158);
buf BUF1 (N278, N277);
xor XOR2 (N279, N273, N158);
not NOT1 (N280, N272);
nand NAND2 (N281, N270, N15);
nand NAND4 (N282, N274, N228, N194, N224);
and AND2 (N283, N280, N242);
nor NOR3 (N284, N281, N87, N39);
and AND3 (N285, N265, N157, N114);
not NOT1 (N286, N285);
buf BUF1 (N287, N260);
and AND2 (N288, N276, N214);
or OR2 (N289, N269, N193);
buf BUF1 (N290, N283);
xor XOR2 (N291, N287, N42);
nand NAND4 (N292, N288, N36, N186, N287);
or OR3 (N293, N290, N205, N24);
nand NAND2 (N294, N278, N241);
xor XOR2 (N295, N291, N153);
buf BUF1 (N296, N289);
and AND2 (N297, N284, N91);
and AND3 (N298, N293, N48, N261);
xor XOR2 (N299, N282, N70);
not NOT1 (N300, N286);
nor NOR2 (N301, N294, N261);
nor NOR3 (N302, N297, N275, N243);
nor NOR2 (N303, N302, N170);
xor XOR2 (N304, N303, N109);
buf BUF1 (N305, N296);
or OR2 (N306, N305, N182);
and AND4 (N307, N295, N254, N32, N73);
not NOT1 (N308, N299);
not NOT1 (N309, N292);
not NOT1 (N310, N300);
nor NOR3 (N311, N310, N192, N295);
nor NOR3 (N312, N309, N220, N10);
buf BUF1 (N313, N279);
not NOT1 (N314, N301);
buf BUF1 (N315, N311);
nand NAND2 (N316, N298, N300);
nand NAND4 (N317, N304, N81, N26, N213);
nor NOR4 (N318, N271, N33, N242, N135);
or OR3 (N319, N312, N174, N85);
nor NOR4 (N320, N307, N98, N98, N159);
not NOT1 (N321, N308);
or OR4 (N322, N316, N125, N191, N8);
not NOT1 (N323, N317);
nand NAND2 (N324, N323, N91);
and AND4 (N325, N324, N164, N313, N323);
not NOT1 (N326, N247);
nand NAND2 (N327, N321, N215);
nor NOR2 (N328, N322, N147);
nand NAND2 (N329, N320, N293);
or OR3 (N330, N306, N127, N317);
nor NOR4 (N331, N328, N174, N293, N170);
nand NAND3 (N332, N329, N216, N102);
nand NAND3 (N333, N319, N182, N201);
nand NAND2 (N334, N327, N231);
not NOT1 (N335, N326);
not NOT1 (N336, N330);
nand NAND3 (N337, N333, N120, N3);
or OR4 (N338, N318, N199, N224, N183);
xor XOR2 (N339, N338, N139);
nand NAND4 (N340, N331, N318, N186, N106);
buf BUF1 (N341, N340);
nor NOR3 (N342, N341, N212, N341);
nand NAND2 (N343, N342, N75);
or OR4 (N344, N334, N171, N322, N124);
buf BUF1 (N345, N339);
not NOT1 (N346, N325);
and AND3 (N347, N343, N257, N20);
and AND2 (N348, N347, N162);
xor XOR2 (N349, N314, N243);
not NOT1 (N350, N346);
nor NOR2 (N351, N336, N84);
buf BUF1 (N352, N332);
or OR2 (N353, N345, N263);
xor XOR2 (N354, N348, N195);
or OR3 (N355, N352, N122, N126);
not NOT1 (N356, N349);
or OR2 (N357, N337, N113);
nor NOR4 (N358, N357, N197, N5, N214);
buf BUF1 (N359, N353);
and AND4 (N360, N358, N254, N145, N249);
nor NOR4 (N361, N350, N37, N75, N338);
and AND3 (N362, N344, N334, N75);
nand NAND3 (N363, N351, N3, N165);
buf BUF1 (N364, N363);
not NOT1 (N365, N360);
nor NOR3 (N366, N356, N175, N161);
or OR3 (N367, N315, N82, N151);
not NOT1 (N368, N355);
xor XOR2 (N369, N335, N255);
xor XOR2 (N370, N365, N294);
buf BUF1 (N371, N368);
and AND4 (N372, N361, N22, N267, N69);
buf BUF1 (N373, N371);
not NOT1 (N374, N369);
and AND2 (N375, N359, N61);
buf BUF1 (N376, N366);
xor XOR2 (N377, N372, N372);
nand NAND3 (N378, N364, N151, N12);
nand NAND2 (N379, N375, N365);
or OR4 (N380, N370, N145, N215, N30);
nor NOR4 (N381, N374, N181, N346, N23);
and AND3 (N382, N376, N276, N294);
or OR3 (N383, N362, N370, N374);
xor XOR2 (N384, N367, N6);
buf BUF1 (N385, N381);
nand NAND2 (N386, N383, N151);
nand NAND2 (N387, N384, N248);
and AND2 (N388, N387, N216);
nand NAND2 (N389, N382, N250);
buf BUF1 (N390, N389);
buf BUF1 (N391, N354);
nand NAND4 (N392, N388, N115, N257, N226);
and AND4 (N393, N385, N242, N311, N109);
nand NAND3 (N394, N390, N257, N44);
nand NAND4 (N395, N386, N103, N89, N394);
or OR3 (N396, N149, N220, N57);
nor NOR3 (N397, N396, N109, N231);
and AND2 (N398, N397, N283);
and AND3 (N399, N377, N176, N119);
and AND4 (N400, N380, N122, N364, N169);
not NOT1 (N401, N391);
or OR2 (N402, N400, N242);
and AND3 (N403, N392, N15, N166);
and AND4 (N404, N403, N101, N34, N375);
and AND4 (N405, N402, N41, N344, N140);
xor XOR2 (N406, N379, N401);
buf BUF1 (N407, N325);
or OR3 (N408, N404, N376, N43);
not NOT1 (N409, N395);
not NOT1 (N410, N373);
and AND4 (N411, N378, N237, N399, N355);
and AND3 (N412, N146, N225, N316);
nor NOR3 (N413, N409, N212, N328);
and AND2 (N414, N408, N203);
buf BUF1 (N415, N412);
and AND2 (N416, N406, N77);
or OR2 (N417, N393, N44);
nor NOR2 (N418, N416, N125);
nand NAND4 (N419, N415, N198, N212, N285);
or OR4 (N420, N410, N132, N136, N87);
not NOT1 (N421, N407);
and AND4 (N422, N411, N61, N17, N26);
or OR2 (N423, N420, N154);
buf BUF1 (N424, N423);
nor NOR2 (N425, N418, N169);
nand NAND2 (N426, N421, N305);
nand NAND3 (N427, N398, N404, N8);
buf BUF1 (N428, N413);
nor NOR3 (N429, N425, N190, N200);
or OR3 (N430, N426, N141, N10);
xor XOR2 (N431, N430, N208);
not NOT1 (N432, N417);
and AND3 (N433, N414, N79, N380);
buf BUF1 (N434, N422);
and AND2 (N435, N431, N408);
buf BUF1 (N436, N434);
xor XOR2 (N437, N405, N143);
and AND4 (N438, N419, N294, N68, N263);
nor NOR2 (N439, N427, N275);
and AND3 (N440, N436, N249, N276);
nand NAND4 (N441, N428, N146, N243, N299);
xor XOR2 (N442, N424, N136);
buf BUF1 (N443, N441);
or OR4 (N444, N438, N124, N376, N181);
or OR4 (N445, N429, N2, N406, N350);
nand NAND3 (N446, N443, N268, N299);
and AND2 (N447, N445, N270);
buf BUF1 (N448, N442);
nor NOR4 (N449, N439, N31, N110, N322);
or OR3 (N450, N432, N321, N421);
or OR3 (N451, N449, N48, N133);
buf BUF1 (N452, N440);
nor NOR2 (N453, N433, N75);
nand NAND3 (N454, N451, N202, N384);
nor NOR2 (N455, N453, N289);
nor NOR3 (N456, N452, N41, N266);
or OR2 (N457, N435, N330);
buf BUF1 (N458, N448);
not NOT1 (N459, N454);
or OR2 (N460, N456, N127);
xor XOR2 (N461, N437, N160);
nand NAND2 (N462, N457, N21);
and AND2 (N463, N460, N269);
nand NAND4 (N464, N444, N215, N453, N222);
xor XOR2 (N465, N464, N359);
or OR2 (N466, N458, N216);
not NOT1 (N467, N466);
and AND2 (N468, N465, N92);
not NOT1 (N469, N467);
nand NAND3 (N470, N455, N432, N233);
nand NAND2 (N471, N446, N223);
xor XOR2 (N472, N470, N189);
buf BUF1 (N473, N459);
xor XOR2 (N474, N461, N289);
and AND2 (N475, N447, N55);
buf BUF1 (N476, N450);
buf BUF1 (N477, N476);
nor NOR3 (N478, N462, N103, N285);
nand NAND2 (N479, N473, N278);
nand NAND3 (N480, N469, N238, N115);
not NOT1 (N481, N471);
xor XOR2 (N482, N478, N422);
buf BUF1 (N483, N481);
or OR2 (N484, N477, N148);
nand NAND3 (N485, N480, N245, N305);
or OR3 (N486, N482, N334, N282);
or OR4 (N487, N486, N410, N138, N134);
xor XOR2 (N488, N475, N162);
nand NAND2 (N489, N479, N2);
buf BUF1 (N490, N468);
xor XOR2 (N491, N488, N345);
nor NOR3 (N492, N490, N297, N412);
not NOT1 (N493, N491);
xor XOR2 (N494, N487, N255);
buf BUF1 (N495, N489);
and AND4 (N496, N483, N136, N2, N270);
xor XOR2 (N497, N495, N490);
nand NAND3 (N498, N493, N33, N103);
nand NAND4 (N499, N485, N221, N340, N51);
buf BUF1 (N500, N497);
nand NAND3 (N501, N498, N488, N437);
nor NOR2 (N502, N492, N35);
nor NOR3 (N503, N501, N115, N61);
buf BUF1 (N504, N494);
nor NOR2 (N505, N474, N412);
xor XOR2 (N506, N500, N21);
buf BUF1 (N507, N505);
nor NOR4 (N508, N504, N2, N56, N235);
and AND3 (N509, N508, N395, N445);
xor XOR2 (N510, N484, N106);
and AND3 (N511, N496, N278, N345);
nand NAND4 (N512, N509, N95, N165, N24);
and AND2 (N513, N472, N428);
and AND2 (N514, N513, N441);
and AND2 (N515, N499, N227);
xor XOR2 (N516, N507, N493);
xor XOR2 (N517, N503, N202);
xor XOR2 (N518, N463, N420);
nand NAND4 (N519, N502, N378, N303, N399);
not NOT1 (N520, N515);
nand NAND4 (N521, N520, N186, N128, N414);
buf BUF1 (N522, N521);
and AND4 (N523, N510, N188, N111, N125);
buf BUF1 (N524, N516);
nand NAND4 (N525, N506, N266, N148, N412);
or OR4 (N526, N514, N430, N479, N14);
and AND4 (N527, N524, N80, N56, N139);
nor NOR4 (N528, N527, N216, N76, N410);
not NOT1 (N529, N525);
nand NAND2 (N530, N522, N160);
or OR2 (N531, N526, N62);
buf BUF1 (N532, N529);
and AND2 (N533, N517, N520);
not NOT1 (N534, N530);
not NOT1 (N535, N518);
not NOT1 (N536, N533);
not NOT1 (N537, N519);
buf BUF1 (N538, N534);
nor NOR2 (N539, N535, N245);
xor XOR2 (N540, N511, N439);
or OR2 (N541, N540, N183);
or OR4 (N542, N512, N407, N143, N367);
and AND3 (N543, N541, N386, N211);
nand NAND4 (N544, N542, N148, N10, N516);
not NOT1 (N545, N536);
xor XOR2 (N546, N538, N177);
nand NAND2 (N547, N523, N105);
nand NAND4 (N548, N537, N383, N282, N301);
nand NAND3 (N549, N547, N68, N330);
xor XOR2 (N550, N549, N125);
and AND4 (N551, N546, N163, N54, N72);
buf BUF1 (N552, N550);
and AND3 (N553, N539, N295, N232);
and AND4 (N554, N531, N147, N487, N76);
or OR4 (N555, N553, N539, N198, N473);
nand NAND4 (N556, N545, N409, N509, N247);
nor NOR4 (N557, N554, N171, N351, N462);
or OR4 (N558, N532, N493, N159, N538);
not NOT1 (N559, N556);
nand NAND2 (N560, N551, N240);
buf BUF1 (N561, N543);
and AND2 (N562, N559, N241);
not NOT1 (N563, N562);
and AND3 (N564, N528, N39, N82);
nor NOR3 (N565, N548, N113, N534);
not NOT1 (N566, N555);
buf BUF1 (N567, N564);
buf BUF1 (N568, N561);
nand NAND3 (N569, N563, N455, N415);
nor NOR3 (N570, N557, N456, N285);
or OR3 (N571, N570, N213, N436);
nand NAND2 (N572, N544, N243);
or OR4 (N573, N567, N235, N402, N139);
and AND2 (N574, N573, N75);
nor NOR4 (N575, N566, N330, N78, N551);
buf BUF1 (N576, N572);
xor XOR2 (N577, N574, N40);
nand NAND2 (N578, N569, N548);
xor XOR2 (N579, N560, N363);
buf BUF1 (N580, N565);
not NOT1 (N581, N552);
or OR2 (N582, N577, N338);
and AND2 (N583, N578, N533);
nand NAND4 (N584, N575, N503, N497, N231);
xor XOR2 (N585, N584, N4);
nand NAND3 (N586, N580, N573, N96);
buf BUF1 (N587, N581);
nand NAND2 (N588, N568, N476);
nor NOR3 (N589, N582, N121, N418);
nand NAND4 (N590, N571, N157, N207, N495);
and AND4 (N591, N587, N95, N469, N450);
buf BUF1 (N592, N585);
nand NAND2 (N593, N558, N565);
or OR4 (N594, N592, N114, N379, N40);
and AND2 (N595, N579, N319);
nand NAND2 (N596, N595, N257);
nor NOR2 (N597, N589, N236);
or OR2 (N598, N583, N554);
not NOT1 (N599, N593);
nand NAND3 (N600, N591, N194, N515);
or OR4 (N601, N590, N538, N363, N247);
nand NAND4 (N602, N600, N224, N429, N434);
nand NAND4 (N603, N586, N291, N326, N137);
or OR4 (N604, N596, N232, N297, N16);
and AND4 (N605, N588, N245, N214, N240);
buf BUF1 (N606, N602);
nand NAND2 (N607, N604, N566);
xor XOR2 (N608, N598, N6);
buf BUF1 (N609, N603);
nand NAND3 (N610, N594, N601, N298);
xor XOR2 (N611, N351, N254);
nor NOR3 (N612, N609, N88, N207);
nor NOR2 (N613, N612, N536);
not NOT1 (N614, N608);
xor XOR2 (N615, N611, N130);
xor XOR2 (N616, N605, N290);
not NOT1 (N617, N614);
nand NAND2 (N618, N615, N384);
or OR4 (N619, N610, N318, N60, N487);
and AND2 (N620, N606, N64);
or OR2 (N621, N613, N372);
not NOT1 (N622, N576);
buf BUF1 (N623, N620);
not NOT1 (N624, N618);
not NOT1 (N625, N599);
or OR3 (N626, N619, N292, N164);
buf BUF1 (N627, N617);
or OR2 (N628, N626, N402);
and AND3 (N629, N621, N331, N362);
not NOT1 (N630, N628);
nand NAND2 (N631, N597, N392);
and AND2 (N632, N631, N64);
not NOT1 (N633, N627);
buf BUF1 (N634, N623);
not NOT1 (N635, N629);
not NOT1 (N636, N633);
and AND3 (N637, N624, N134, N181);
and AND2 (N638, N622, N193);
not NOT1 (N639, N638);
buf BUF1 (N640, N630);
and AND2 (N641, N640, N297);
not NOT1 (N642, N636);
and AND4 (N643, N641, N24, N137, N364);
buf BUF1 (N644, N625);
xor XOR2 (N645, N635, N481);
not NOT1 (N646, N643);
nand NAND3 (N647, N642, N536, N56);
xor XOR2 (N648, N645, N213);
xor XOR2 (N649, N644, N195);
not NOT1 (N650, N646);
not NOT1 (N651, N616);
nor NOR4 (N652, N634, N217, N635, N129);
not NOT1 (N653, N632);
or OR4 (N654, N650, N507, N538, N493);
or OR2 (N655, N652, N206);
nor NOR2 (N656, N649, N123);
and AND2 (N657, N653, N527);
buf BUF1 (N658, N657);
and AND3 (N659, N639, N185, N559);
and AND3 (N660, N607, N584, N58);
buf BUF1 (N661, N656);
buf BUF1 (N662, N660);
and AND2 (N663, N637, N326);
xor XOR2 (N664, N651, N310);
xor XOR2 (N665, N662, N93);
xor XOR2 (N666, N647, N3);
buf BUF1 (N667, N661);
xor XOR2 (N668, N666, N444);
xor XOR2 (N669, N654, N20);
buf BUF1 (N670, N663);
nor NOR4 (N671, N655, N238, N8, N321);
xor XOR2 (N672, N659, N180);
not NOT1 (N673, N667);
and AND3 (N674, N664, N347, N524);
nand NAND4 (N675, N648, N490, N138, N576);
not NOT1 (N676, N669);
nand NAND4 (N677, N675, N433, N388, N615);
and AND3 (N678, N670, N99, N93);
and AND3 (N679, N658, N519, N455);
xor XOR2 (N680, N671, N163);
not NOT1 (N681, N665);
nor NOR2 (N682, N679, N2);
xor XOR2 (N683, N668, N337);
or OR4 (N684, N681, N228, N262, N239);
xor XOR2 (N685, N682, N32);
not NOT1 (N686, N684);
and AND4 (N687, N678, N623, N474, N124);
or OR2 (N688, N683, N103);
not NOT1 (N689, N673);
not NOT1 (N690, N680);
or OR3 (N691, N676, N359, N147);
xor XOR2 (N692, N690, N318);
not NOT1 (N693, N685);
nor NOR3 (N694, N672, N439, N568);
not NOT1 (N695, N694);
nand NAND4 (N696, N687, N629, N289, N225);
nor NOR4 (N697, N691, N38, N212, N434);
and AND2 (N698, N688, N198);
and AND3 (N699, N674, N232, N188);
and AND4 (N700, N686, N616, N619, N601);
xor XOR2 (N701, N695, N611);
xor XOR2 (N702, N699, N60);
and AND4 (N703, N696, N308, N311, N319);
buf BUF1 (N704, N693);
nor NOR2 (N705, N702, N291);
and AND2 (N706, N700, N506);
nor NOR2 (N707, N706, N155);
nand NAND4 (N708, N704, N330, N62, N258);
not NOT1 (N709, N705);
and AND3 (N710, N692, N271, N405);
and AND2 (N711, N709, N633);
nor NOR4 (N712, N698, N61, N219, N708);
buf BUF1 (N713, N151);
nor NOR2 (N714, N701, N162);
nand NAND2 (N715, N712, N667);
or OR3 (N716, N713, N475, N201);
buf BUF1 (N717, N707);
or OR4 (N718, N716, N445, N274, N176);
nand NAND2 (N719, N718, N481);
or OR2 (N720, N703, N643);
and AND4 (N721, N719, N97, N674, N153);
or OR2 (N722, N710, N281);
xor XOR2 (N723, N711, N406);
buf BUF1 (N724, N720);
nand NAND4 (N725, N715, N328, N231, N363);
or OR2 (N726, N722, N586);
not NOT1 (N727, N677);
xor XOR2 (N728, N726, N370);
nor NOR4 (N729, N717, N140, N123, N334);
nor NOR3 (N730, N714, N463, N247);
or OR4 (N731, N725, N324, N535, N681);
buf BUF1 (N732, N728);
or OR3 (N733, N730, N670, N326);
or OR3 (N734, N697, N670, N657);
or OR2 (N735, N721, N186);
not NOT1 (N736, N735);
not NOT1 (N737, N732);
nor NOR2 (N738, N731, N492);
xor XOR2 (N739, N738, N712);
nor NOR3 (N740, N727, N164, N200);
buf BUF1 (N741, N724);
nor NOR3 (N742, N736, N426, N39);
not NOT1 (N743, N742);
xor XOR2 (N744, N737, N225);
or OR4 (N745, N743, N237, N502, N690);
buf BUF1 (N746, N723);
and AND2 (N747, N689, N720);
nand NAND2 (N748, N740, N445);
xor XOR2 (N749, N748, N221);
and AND2 (N750, N734, N97);
and AND2 (N751, N739, N658);
not NOT1 (N752, N744);
and AND4 (N753, N733, N141, N586, N255);
xor XOR2 (N754, N746, N468);
nor NOR4 (N755, N754, N345, N143, N225);
nor NOR4 (N756, N752, N446, N452, N422);
and AND2 (N757, N741, N139);
xor XOR2 (N758, N747, N524);
or OR4 (N759, N729, N355, N492, N731);
nand NAND2 (N760, N759, N243);
xor XOR2 (N761, N750, N418);
xor XOR2 (N762, N749, N518);
not NOT1 (N763, N745);
nand NAND3 (N764, N756, N202, N123);
xor XOR2 (N765, N751, N575);
xor XOR2 (N766, N758, N261);
not NOT1 (N767, N766);
xor XOR2 (N768, N753, N277);
and AND4 (N769, N755, N636, N98, N550);
xor XOR2 (N770, N767, N282);
nand NAND4 (N771, N761, N7, N630, N674);
and AND2 (N772, N764, N207);
nand NAND4 (N773, N769, N164, N99, N409);
buf BUF1 (N774, N773);
buf BUF1 (N775, N770);
nor NOR4 (N776, N757, N115, N189, N180);
buf BUF1 (N777, N771);
nor NOR4 (N778, N774, N192, N483, N490);
nor NOR3 (N779, N776, N706, N74);
buf BUF1 (N780, N772);
xor XOR2 (N781, N768, N213);
nor NOR3 (N782, N780, N434, N671);
or OR2 (N783, N763, N17);
nor NOR3 (N784, N778, N347, N242);
or OR2 (N785, N784, N712);
and AND4 (N786, N775, N352, N513, N563);
xor XOR2 (N787, N760, N769);
nor NOR4 (N788, N787, N546, N423, N243);
nor NOR2 (N789, N788, N456);
or OR4 (N790, N789, N429, N772, N135);
nand NAND3 (N791, N782, N342, N178);
buf BUF1 (N792, N762);
not NOT1 (N793, N790);
nor NOR4 (N794, N791, N170, N507, N659);
not NOT1 (N795, N779);
or OR3 (N796, N793, N725, N520);
nor NOR4 (N797, N786, N796, N476, N732);
nor NOR4 (N798, N573, N141, N232, N165);
xor XOR2 (N799, N785, N542);
and AND2 (N800, N797, N400);
nor NOR3 (N801, N777, N253, N660);
buf BUF1 (N802, N795);
nor NOR2 (N803, N798, N123);
nand NAND3 (N804, N803, N50, N540);
or OR2 (N805, N783, N672);
not NOT1 (N806, N804);
nor NOR3 (N807, N765, N423, N468);
or OR2 (N808, N805, N322);
nand NAND2 (N809, N806, N120);
buf BUF1 (N810, N792);
nand NAND4 (N811, N800, N632, N435, N585);
not NOT1 (N812, N794);
xor XOR2 (N813, N799, N224);
or OR2 (N814, N808, N219);
not NOT1 (N815, N813);
and AND3 (N816, N811, N57, N617);
nand NAND4 (N817, N807, N636, N427, N692);
buf BUF1 (N818, N815);
xor XOR2 (N819, N812, N518);
xor XOR2 (N820, N819, N230);
nand NAND4 (N821, N810, N102, N45, N129);
and AND4 (N822, N814, N205, N779, N789);
nor NOR2 (N823, N809, N300);
nor NOR4 (N824, N801, N441, N474, N332);
not NOT1 (N825, N816);
and AND4 (N826, N825, N518, N517, N650);
or OR3 (N827, N823, N197, N181);
nand NAND2 (N828, N817, N371);
not NOT1 (N829, N824);
nor NOR4 (N830, N828, N141, N326, N447);
or OR4 (N831, N827, N548, N211, N22);
nor NOR2 (N832, N829, N822);
and AND2 (N833, N795, N777);
nor NOR4 (N834, N826, N157, N357, N84);
nand NAND3 (N835, N781, N331, N137);
xor XOR2 (N836, N835, N701);
nor NOR2 (N837, N818, N265);
or OR3 (N838, N832, N154, N562);
not NOT1 (N839, N830);
and AND3 (N840, N820, N575, N444);
not NOT1 (N841, N834);
buf BUF1 (N842, N821);
not NOT1 (N843, N840);
xor XOR2 (N844, N802, N54);
or OR4 (N845, N839, N489, N460, N403);
not NOT1 (N846, N838);
xor XOR2 (N847, N833, N525);
buf BUF1 (N848, N847);
xor XOR2 (N849, N831, N465);
not NOT1 (N850, N842);
nor NOR3 (N851, N845, N409, N727);
or OR4 (N852, N849, N333, N457, N328);
nand NAND3 (N853, N841, N256, N494);
xor XOR2 (N854, N850, N650);
nand NAND2 (N855, N853, N133);
not NOT1 (N856, N844);
nand NAND3 (N857, N837, N517, N373);
nand NAND3 (N858, N836, N726, N590);
not NOT1 (N859, N855);
or OR4 (N860, N848, N807, N438, N698);
and AND2 (N861, N854, N699);
or OR3 (N862, N843, N725, N846);
or OR4 (N863, N160, N231, N461, N660);
nand NAND3 (N864, N857, N130, N487);
or OR2 (N865, N860, N451);
nand NAND3 (N866, N863, N626, N744);
or OR3 (N867, N861, N643, N390);
and AND4 (N868, N862, N717, N371, N648);
buf BUF1 (N869, N868);
xor XOR2 (N870, N867, N242);
xor XOR2 (N871, N851, N342);
xor XOR2 (N872, N866, N739);
nand NAND3 (N873, N865, N21, N826);
buf BUF1 (N874, N869);
nor NOR4 (N875, N871, N646, N627, N111);
nand NAND2 (N876, N864, N327);
and AND2 (N877, N873, N528);
and AND2 (N878, N859, N535);
not NOT1 (N879, N878);
nor NOR4 (N880, N852, N244, N541, N409);
or OR2 (N881, N875, N215);
xor XOR2 (N882, N880, N738);
or OR4 (N883, N856, N347, N171, N664);
xor XOR2 (N884, N870, N627);
or OR4 (N885, N879, N819, N785, N140);
and AND2 (N886, N881, N59);
xor XOR2 (N887, N882, N573);
nor NOR2 (N888, N884, N842);
nand NAND3 (N889, N874, N589, N399);
not NOT1 (N890, N876);
buf BUF1 (N891, N883);
nand NAND3 (N892, N887, N689, N591);
and AND3 (N893, N891, N568, N766);
nand NAND3 (N894, N888, N611, N878);
xor XOR2 (N895, N894, N275);
not NOT1 (N896, N885);
or OR4 (N897, N896, N36, N596, N76);
not NOT1 (N898, N858);
nand NAND3 (N899, N877, N72, N261);
nor NOR3 (N900, N899, N761, N878);
nor NOR2 (N901, N872, N615);
and AND4 (N902, N893, N88, N84, N39);
nand NAND4 (N903, N902, N555, N363, N630);
not NOT1 (N904, N900);
or OR3 (N905, N904, N141, N758);
nand NAND3 (N906, N886, N417, N270);
nand NAND2 (N907, N895, N190);
not NOT1 (N908, N897);
xor XOR2 (N909, N903, N321);
xor XOR2 (N910, N907, N662);
or OR4 (N911, N898, N193, N273, N538);
and AND2 (N912, N911, N358);
xor XOR2 (N913, N908, N535);
and AND3 (N914, N913, N823, N604);
and AND4 (N915, N901, N318, N50, N245);
not NOT1 (N916, N905);
xor XOR2 (N917, N914, N212);
nand NAND2 (N918, N892, N38);
not NOT1 (N919, N910);
nor NOR4 (N920, N890, N79, N903, N276);
buf BUF1 (N921, N920);
buf BUF1 (N922, N921);
xor XOR2 (N923, N915, N372);
nand NAND3 (N924, N916, N819, N197);
nand NAND2 (N925, N906, N708);
not NOT1 (N926, N918);
nand NAND2 (N927, N923, N641);
nor NOR4 (N928, N917, N581, N163, N364);
not NOT1 (N929, N925);
nand NAND3 (N930, N928, N542, N52);
xor XOR2 (N931, N924, N123);
nand NAND2 (N932, N922, N573);
and AND3 (N933, N929, N381, N576);
or OR2 (N934, N912, N3);
and AND3 (N935, N932, N856, N213);
buf BUF1 (N936, N927);
and AND3 (N937, N936, N663, N627);
nor NOR2 (N938, N937, N15);
nor NOR2 (N939, N919, N521);
nor NOR4 (N940, N935, N603, N753, N434);
nand NAND3 (N941, N889, N241, N473);
nor NOR2 (N942, N931, N504);
not NOT1 (N943, N909);
xor XOR2 (N944, N938, N205);
nor NOR2 (N945, N934, N274);
and AND4 (N946, N940, N852, N926, N437);
xor XOR2 (N947, N472, N669);
buf BUF1 (N948, N944);
nand NAND2 (N949, N930, N440);
xor XOR2 (N950, N942, N272);
and AND2 (N951, N943, N605);
or OR3 (N952, N945, N410, N208);
and AND2 (N953, N933, N482);
or OR3 (N954, N952, N594, N255);
nor NOR3 (N955, N939, N269, N932);
nand NAND4 (N956, N951, N757, N48, N543);
and AND4 (N957, N956, N261, N705, N247);
xor XOR2 (N958, N941, N55);
not NOT1 (N959, N958);
nand NAND4 (N960, N948, N567, N482, N869);
or OR3 (N961, N947, N583, N209);
not NOT1 (N962, N959);
nor NOR3 (N963, N960, N350, N938);
buf BUF1 (N964, N957);
xor XOR2 (N965, N964, N292);
nand NAND3 (N966, N953, N232, N81);
or OR2 (N967, N966, N941);
nor NOR2 (N968, N950, N962);
buf BUF1 (N969, N375);
or OR3 (N970, N946, N492, N964);
and AND4 (N971, N967, N337, N101, N661);
nand NAND2 (N972, N969, N848);
nand NAND4 (N973, N949, N82, N588, N723);
nand NAND4 (N974, N968, N291, N637, N784);
or OR3 (N975, N961, N939, N697);
or OR2 (N976, N972, N703);
xor XOR2 (N977, N963, N298);
nand NAND4 (N978, N973, N608, N374, N215);
buf BUF1 (N979, N970);
buf BUF1 (N980, N976);
nand NAND3 (N981, N980, N633, N412);
buf BUF1 (N982, N977);
not NOT1 (N983, N954);
nor NOR3 (N984, N978, N770, N255);
nand NAND2 (N985, N955, N601);
nor NOR3 (N986, N971, N642, N566);
xor XOR2 (N987, N986, N416);
xor XOR2 (N988, N983, N279);
xor XOR2 (N989, N982, N342);
nand NAND4 (N990, N987, N802, N432, N378);
xor XOR2 (N991, N975, N784);
and AND4 (N992, N988, N591, N590, N669);
buf BUF1 (N993, N965);
nor NOR3 (N994, N993, N495, N252);
and AND2 (N995, N991, N10);
buf BUF1 (N996, N994);
and AND4 (N997, N990, N485, N48, N36);
or OR4 (N998, N989, N9, N880, N804);
or OR4 (N999, N997, N72, N258, N608);
buf BUF1 (N1000, N999);
and AND4 (N1001, N974, N91, N186, N91);
or OR2 (N1002, N996, N645);
not NOT1 (N1003, N979);
not NOT1 (N1004, N1002);
and AND3 (N1005, N1003, N931, N304);
xor XOR2 (N1006, N1005, N404);
buf BUF1 (N1007, N1006);
not NOT1 (N1008, N1007);
and AND3 (N1009, N981, N548, N171);
xor XOR2 (N1010, N998, N484);
buf BUF1 (N1011, N1008);
nor NOR3 (N1012, N1001, N100, N145);
buf BUF1 (N1013, N1012);
buf BUF1 (N1014, N985);
nor NOR3 (N1015, N1009, N576, N390);
or OR4 (N1016, N984, N104, N644, N216);
nand NAND4 (N1017, N1013, N472, N293, N825);
not NOT1 (N1018, N1011);
not NOT1 (N1019, N992);
nand NAND2 (N1020, N1019, N670);
and AND2 (N1021, N1018, N428);
nor NOR4 (N1022, N1000, N749, N85, N685);
or OR4 (N1023, N1020, N729, N794, N739);
buf BUF1 (N1024, N1016);
or OR2 (N1025, N1017, N535);
not NOT1 (N1026, N1022);
nand NAND4 (N1027, N995, N30, N111, N380);
xor XOR2 (N1028, N1014, N833);
or OR3 (N1029, N1021, N851, N839);
not NOT1 (N1030, N1026);
nand NAND3 (N1031, N1030, N566, N928);
not NOT1 (N1032, N1023);
or OR4 (N1033, N1015, N485, N961, N490);
or OR3 (N1034, N1027, N584, N787);
xor XOR2 (N1035, N1025, N456);
or OR3 (N1036, N1004, N1021, N179);
or OR4 (N1037, N1031, N199, N202, N254);
or OR4 (N1038, N1010, N537, N609, N237);
nand NAND3 (N1039, N1033, N431, N567);
and AND4 (N1040, N1036, N158, N997, N194);
and AND3 (N1041, N1028, N644, N1007);
and AND2 (N1042, N1035, N845);
nand NAND3 (N1043, N1037, N173, N315);
nand NAND3 (N1044, N1038, N919, N485);
and AND2 (N1045, N1042, N363);
nand NAND2 (N1046, N1044, N1027);
and AND4 (N1047, N1034, N189, N509, N721);
nor NOR4 (N1048, N1024, N334, N583, N422);
nor NOR4 (N1049, N1046, N482, N850, N892);
xor XOR2 (N1050, N1029, N773);
xor XOR2 (N1051, N1045, N1009);
and AND3 (N1052, N1041, N508, N153);
xor XOR2 (N1053, N1048, N339);
or OR2 (N1054, N1032, N45);
nand NAND2 (N1055, N1047, N60);
nor NOR4 (N1056, N1040, N614, N321, N122);
not NOT1 (N1057, N1053);
and AND4 (N1058, N1052, N897, N908, N500);
nand NAND2 (N1059, N1057, N61);
buf BUF1 (N1060, N1058);
xor XOR2 (N1061, N1055, N1057);
nor NOR2 (N1062, N1056, N426);
and AND2 (N1063, N1039, N207);
and AND2 (N1064, N1063, N558);
buf BUF1 (N1065, N1060);
buf BUF1 (N1066, N1061);
and AND2 (N1067, N1064, N956);
nand NAND4 (N1068, N1049, N820, N647, N592);
buf BUF1 (N1069, N1043);
not NOT1 (N1070, N1068);
or OR2 (N1071, N1070, N242);
not NOT1 (N1072, N1050);
and AND2 (N1073, N1051, N448);
or OR4 (N1074, N1072, N74, N456, N646);
buf BUF1 (N1075, N1062);
buf BUF1 (N1076, N1059);
buf BUF1 (N1077, N1067);
not NOT1 (N1078, N1054);
nand NAND2 (N1079, N1076, N738);
or OR2 (N1080, N1065, N323);
buf BUF1 (N1081, N1066);
not NOT1 (N1082, N1075);
xor XOR2 (N1083, N1077, N722);
or OR3 (N1084, N1083, N400, N551);
or OR4 (N1085, N1079, N651, N412, N431);
or OR4 (N1086, N1071, N382, N915, N589);
buf BUF1 (N1087, N1074);
not NOT1 (N1088, N1085);
not NOT1 (N1089, N1082);
nand NAND4 (N1090, N1084, N945, N409, N918);
and AND3 (N1091, N1088, N1004, N1054);
nand NAND2 (N1092, N1069, N43);
buf BUF1 (N1093, N1091);
not NOT1 (N1094, N1089);
and AND4 (N1095, N1073, N948, N125, N898);
not NOT1 (N1096, N1086);
nand NAND2 (N1097, N1080, N541);
and AND3 (N1098, N1092, N546, N180);
buf BUF1 (N1099, N1090);
and AND2 (N1100, N1093, N98);
and AND2 (N1101, N1098, N623);
nand NAND4 (N1102, N1081, N527, N243, N1000);
not NOT1 (N1103, N1087);
or OR4 (N1104, N1096, N860, N758, N758);
buf BUF1 (N1105, N1101);
nor NOR3 (N1106, N1102, N1062, N193);
not NOT1 (N1107, N1099);
nand NAND3 (N1108, N1105, N431, N703);
buf BUF1 (N1109, N1106);
nand NAND2 (N1110, N1107, N165);
and AND3 (N1111, N1110, N974, N257);
not NOT1 (N1112, N1104);
or OR3 (N1113, N1112, N838, N793);
nor NOR4 (N1114, N1108, N900, N435, N400);
nor NOR2 (N1115, N1113, N101);
buf BUF1 (N1116, N1103);
not NOT1 (N1117, N1078);
and AND2 (N1118, N1095, N545);
nor NOR4 (N1119, N1114, N611, N522, N605);
buf BUF1 (N1120, N1118);
xor XOR2 (N1121, N1120, N136);
or OR3 (N1122, N1117, N167, N104);
not NOT1 (N1123, N1115);
xor XOR2 (N1124, N1109, N656);
xor XOR2 (N1125, N1116, N837);
not NOT1 (N1126, N1111);
nand NAND4 (N1127, N1122, N236, N780, N362);
nand NAND4 (N1128, N1097, N754, N997, N485);
buf BUF1 (N1129, N1123);
xor XOR2 (N1130, N1100, N737);
not NOT1 (N1131, N1129);
nor NOR4 (N1132, N1130, N119, N41, N53);
or OR3 (N1133, N1132, N53, N711);
nor NOR3 (N1134, N1131, N582, N360);
nor NOR3 (N1135, N1126, N634, N931);
or OR2 (N1136, N1127, N1033);
buf BUF1 (N1137, N1128);
xor XOR2 (N1138, N1137, N42);
or OR4 (N1139, N1125, N183, N1124, N548);
xor XOR2 (N1140, N425, N67);
xor XOR2 (N1141, N1135, N1096);
buf BUF1 (N1142, N1134);
not NOT1 (N1143, N1119);
and AND4 (N1144, N1142, N841, N950, N398);
or OR4 (N1145, N1138, N180, N488, N319);
nand NAND3 (N1146, N1145, N688, N574);
or OR4 (N1147, N1144, N831, N40, N683);
nand NAND4 (N1148, N1141, N756, N934, N551);
xor XOR2 (N1149, N1146, N270);
or OR4 (N1150, N1140, N475, N581, N620);
and AND2 (N1151, N1121, N229);
nor NOR3 (N1152, N1150, N264, N335);
nand NAND2 (N1153, N1133, N425);
nor NOR4 (N1154, N1139, N1010, N990, N208);
xor XOR2 (N1155, N1152, N456);
xor XOR2 (N1156, N1153, N850);
nor NOR4 (N1157, N1143, N306, N732, N219);
not NOT1 (N1158, N1094);
xor XOR2 (N1159, N1154, N1139);
buf BUF1 (N1160, N1151);
buf BUF1 (N1161, N1156);
not NOT1 (N1162, N1147);
nor NOR3 (N1163, N1160, N20, N256);
nor NOR2 (N1164, N1157, N354);
nand NAND2 (N1165, N1158, N275);
nand NAND2 (N1166, N1136, N517);
or OR3 (N1167, N1155, N4, N601);
or OR3 (N1168, N1166, N204, N663);
or OR4 (N1169, N1167, N155, N398, N408);
buf BUF1 (N1170, N1169);
nor NOR4 (N1171, N1148, N706, N725, N223);
nand NAND3 (N1172, N1162, N23, N279);
not NOT1 (N1173, N1168);
xor XOR2 (N1174, N1149, N371);
nor NOR4 (N1175, N1174, N216, N237, N63);
not NOT1 (N1176, N1172);
and AND4 (N1177, N1159, N240, N677, N930);
or OR3 (N1178, N1170, N129, N451);
nor NOR4 (N1179, N1176, N276, N1153, N1058);
and AND4 (N1180, N1161, N795, N952, N568);
buf BUF1 (N1181, N1163);
nand NAND3 (N1182, N1171, N1036, N990);
nand NAND2 (N1183, N1177, N608);
nor NOR4 (N1184, N1181, N86, N1085, N501);
buf BUF1 (N1185, N1183);
nand NAND2 (N1186, N1173, N772);
xor XOR2 (N1187, N1165, N907);
and AND2 (N1188, N1185, N13);
nor NOR4 (N1189, N1164, N715, N186, N747);
not NOT1 (N1190, N1186);
nor NOR2 (N1191, N1178, N190);
and AND2 (N1192, N1188, N1178);
and AND4 (N1193, N1184, N1092, N30, N1183);
or OR4 (N1194, N1189, N419, N832, N927);
nor NOR2 (N1195, N1190, N1019);
buf BUF1 (N1196, N1192);
nor NOR3 (N1197, N1196, N495, N196);
or OR2 (N1198, N1182, N387);
nand NAND3 (N1199, N1180, N895, N481);
nand NAND2 (N1200, N1193, N864);
or OR2 (N1201, N1200, N492);
and AND4 (N1202, N1195, N1032, N769, N422);
nand NAND2 (N1203, N1179, N93);
nand NAND2 (N1204, N1191, N31);
and AND3 (N1205, N1204, N185, N885);
not NOT1 (N1206, N1203);
buf BUF1 (N1207, N1199);
and AND3 (N1208, N1175, N1112, N935);
buf BUF1 (N1209, N1187);
nand NAND3 (N1210, N1207, N998, N124);
nand NAND3 (N1211, N1205, N417, N194);
not NOT1 (N1212, N1198);
nor NOR3 (N1213, N1211, N819, N238);
or OR3 (N1214, N1210, N658, N618);
nor NOR3 (N1215, N1197, N257, N986);
nand NAND3 (N1216, N1209, N814, N480);
or OR3 (N1217, N1213, N1029, N14);
nor NOR2 (N1218, N1216, N440);
buf BUF1 (N1219, N1206);
xor XOR2 (N1220, N1208, N437);
or OR3 (N1221, N1218, N353, N294);
buf BUF1 (N1222, N1221);
nor NOR3 (N1223, N1215, N116, N110);
and AND3 (N1224, N1220, N181, N498);
nor NOR2 (N1225, N1202, N146);
nand NAND4 (N1226, N1224, N629, N486, N768);
xor XOR2 (N1227, N1225, N808);
buf BUF1 (N1228, N1194);
or OR2 (N1229, N1217, N800);
or OR4 (N1230, N1222, N610, N1060, N327);
nand NAND2 (N1231, N1219, N734);
and AND4 (N1232, N1229, N176, N35, N164);
not NOT1 (N1233, N1214);
or OR3 (N1234, N1231, N673, N193);
and AND3 (N1235, N1230, N932, N751);
buf BUF1 (N1236, N1227);
buf BUF1 (N1237, N1232);
or OR4 (N1238, N1236, N808, N487, N128);
and AND3 (N1239, N1212, N752, N448);
not NOT1 (N1240, N1235);
and AND3 (N1241, N1233, N329, N391);
nand NAND4 (N1242, N1237, N1165, N1231, N922);
not NOT1 (N1243, N1239);
nand NAND3 (N1244, N1240, N806, N972);
nand NAND4 (N1245, N1241, N1202, N574, N128);
xor XOR2 (N1246, N1201, N849);
not NOT1 (N1247, N1238);
not NOT1 (N1248, N1247);
buf BUF1 (N1249, N1245);
or OR2 (N1250, N1228, N204);
nor NOR3 (N1251, N1248, N109, N430);
nand NAND3 (N1252, N1234, N594, N603);
buf BUF1 (N1253, N1244);
buf BUF1 (N1254, N1250);
or OR3 (N1255, N1249, N1151, N179);
nand NAND2 (N1256, N1253, N476);
nand NAND3 (N1257, N1242, N837, N930);
nand NAND4 (N1258, N1254, N1180, N1015, N976);
and AND3 (N1259, N1258, N135, N398);
nand NAND3 (N1260, N1252, N290, N483);
buf BUF1 (N1261, N1243);
buf BUF1 (N1262, N1259);
buf BUF1 (N1263, N1260);
not NOT1 (N1264, N1256);
and AND3 (N1265, N1261, N114, N578);
buf BUF1 (N1266, N1251);
buf BUF1 (N1267, N1255);
buf BUF1 (N1268, N1264);
buf BUF1 (N1269, N1267);
nand NAND4 (N1270, N1266, N324, N600, N496);
and AND2 (N1271, N1226, N405);
buf BUF1 (N1272, N1265);
or OR3 (N1273, N1270, N430, N1124);
or OR2 (N1274, N1257, N721);
or OR2 (N1275, N1273, N596);
xor XOR2 (N1276, N1269, N1196);
not NOT1 (N1277, N1263);
xor XOR2 (N1278, N1223, N324);
xor XOR2 (N1279, N1246, N1007);
or OR2 (N1280, N1279, N686);
nand NAND2 (N1281, N1275, N111);
not NOT1 (N1282, N1281);
and AND2 (N1283, N1271, N241);
buf BUF1 (N1284, N1278);
xor XOR2 (N1285, N1262, N139);
and AND4 (N1286, N1272, N247, N879, N1247);
nor NOR2 (N1287, N1268, N315);
or OR4 (N1288, N1274, N1007, N657, N814);
buf BUF1 (N1289, N1286);
buf BUF1 (N1290, N1287);
nor NOR2 (N1291, N1283, N400);
not NOT1 (N1292, N1289);
nor NOR4 (N1293, N1291, N594, N47, N622);
nor NOR2 (N1294, N1277, N181);
buf BUF1 (N1295, N1290);
xor XOR2 (N1296, N1292, N1094);
nor NOR4 (N1297, N1280, N317, N618, N1013);
and AND3 (N1298, N1295, N160, N628);
or OR3 (N1299, N1284, N694, N1006);
xor XOR2 (N1300, N1293, N741);
and AND3 (N1301, N1297, N264, N301);
nand NAND2 (N1302, N1301, N641);
or OR4 (N1303, N1285, N581, N914, N242);
and AND3 (N1304, N1298, N586, N799);
buf BUF1 (N1305, N1300);
or OR4 (N1306, N1276, N508, N636, N120);
nor NOR2 (N1307, N1288, N984);
xor XOR2 (N1308, N1303, N940);
not NOT1 (N1309, N1305);
not NOT1 (N1310, N1294);
xor XOR2 (N1311, N1282, N944);
and AND3 (N1312, N1308, N857, N93);
nand NAND4 (N1313, N1302, N475, N702, N496);
or OR4 (N1314, N1296, N867, N266, N246);
and AND3 (N1315, N1313, N890, N969);
and AND3 (N1316, N1311, N645, N1072);
not NOT1 (N1317, N1310);
xor XOR2 (N1318, N1307, N721);
nand NAND3 (N1319, N1312, N694, N329);
xor XOR2 (N1320, N1299, N575);
xor XOR2 (N1321, N1315, N594);
and AND2 (N1322, N1316, N1109);
xor XOR2 (N1323, N1306, N136);
not NOT1 (N1324, N1323);
nor NOR4 (N1325, N1304, N896, N1153, N509);
nand NAND2 (N1326, N1321, N756);
and AND3 (N1327, N1319, N209, N749);
or OR4 (N1328, N1318, N386, N1124, N628);
not NOT1 (N1329, N1322);
nand NAND3 (N1330, N1309, N724, N1055);
buf BUF1 (N1331, N1325);
or OR3 (N1332, N1328, N674, N1085);
not NOT1 (N1333, N1330);
and AND2 (N1334, N1326, N463);
nor NOR4 (N1335, N1324, N493, N221, N401);
not NOT1 (N1336, N1335);
nor NOR3 (N1337, N1333, N284, N873);
nand NAND3 (N1338, N1332, N122, N714);
and AND3 (N1339, N1320, N763, N890);
nand NAND3 (N1340, N1327, N1229, N1062);
and AND3 (N1341, N1314, N66, N293);
buf BUF1 (N1342, N1331);
and AND2 (N1343, N1329, N64);
xor XOR2 (N1344, N1339, N559);
nand NAND3 (N1345, N1336, N841, N1034);
buf BUF1 (N1346, N1342);
buf BUF1 (N1347, N1346);
and AND2 (N1348, N1345, N941);
xor XOR2 (N1349, N1340, N1086);
or OR2 (N1350, N1349, N1193);
not NOT1 (N1351, N1350);
nor NOR4 (N1352, N1338, N265, N600, N1137);
and AND2 (N1353, N1351, N34);
buf BUF1 (N1354, N1337);
buf BUF1 (N1355, N1353);
buf BUF1 (N1356, N1352);
nor NOR4 (N1357, N1317, N937, N971, N927);
and AND4 (N1358, N1347, N171, N263, N863);
not NOT1 (N1359, N1348);
and AND2 (N1360, N1334, N461);
not NOT1 (N1361, N1359);
buf BUF1 (N1362, N1358);
buf BUF1 (N1363, N1362);
or OR3 (N1364, N1356, N97, N1130);
buf BUF1 (N1365, N1355);
nor NOR2 (N1366, N1363, N347);
and AND2 (N1367, N1366, N1065);
buf BUF1 (N1368, N1367);
buf BUF1 (N1369, N1357);
not NOT1 (N1370, N1343);
nor NOR2 (N1371, N1360, N198);
nand NAND4 (N1372, N1364, N1078, N462, N337);
not NOT1 (N1373, N1341);
and AND3 (N1374, N1370, N364, N392);
nand NAND2 (N1375, N1354, N94);
and AND4 (N1376, N1365, N1023, N661, N124);
and AND3 (N1377, N1375, N1043, N62);
and AND3 (N1378, N1374, N784, N211);
nand NAND3 (N1379, N1361, N1100, N1228);
not NOT1 (N1380, N1344);
xor XOR2 (N1381, N1380, N1290);
and AND2 (N1382, N1373, N993);
or OR3 (N1383, N1376, N869, N1171);
or OR4 (N1384, N1379, N1343, N1115, N1045);
buf BUF1 (N1385, N1384);
nor NOR4 (N1386, N1371, N1156, N902, N474);
nor NOR4 (N1387, N1383, N545, N734, N1089);
and AND2 (N1388, N1377, N798);
nor NOR4 (N1389, N1382, N1387, N1153, N1245);
buf BUF1 (N1390, N759);
xor XOR2 (N1391, N1389, N232);
nor NOR2 (N1392, N1368, N150);
and AND2 (N1393, N1391, N151);
nand NAND3 (N1394, N1372, N16, N582);
buf BUF1 (N1395, N1394);
and AND2 (N1396, N1393, N979);
and AND3 (N1397, N1386, N1200, N605);
buf BUF1 (N1398, N1369);
not NOT1 (N1399, N1396);
nor NOR3 (N1400, N1378, N745, N402);
or OR3 (N1401, N1398, N452, N983);
not NOT1 (N1402, N1392);
not NOT1 (N1403, N1401);
buf BUF1 (N1404, N1395);
xor XOR2 (N1405, N1397, N642);
xor XOR2 (N1406, N1385, N354);
not NOT1 (N1407, N1402);
buf BUF1 (N1408, N1400);
or OR2 (N1409, N1408, N1270);
xor XOR2 (N1410, N1405, N327);
and AND4 (N1411, N1407, N1127, N76, N862);
nor NOR2 (N1412, N1403, N150);
and AND4 (N1413, N1406, N793, N415, N1023);
or OR2 (N1414, N1399, N776);
buf BUF1 (N1415, N1411);
xor XOR2 (N1416, N1413, N1274);
not NOT1 (N1417, N1404);
xor XOR2 (N1418, N1414, N1292);
and AND2 (N1419, N1409, N1137);
and AND2 (N1420, N1390, N1107);
buf BUF1 (N1421, N1388);
buf BUF1 (N1422, N1381);
or OR4 (N1423, N1422, N897, N936, N212);
nand NAND3 (N1424, N1412, N517, N575);
nor NOR2 (N1425, N1417, N83);
nor NOR2 (N1426, N1410, N481);
and AND3 (N1427, N1415, N1399, N281);
and AND2 (N1428, N1427, N1393);
xor XOR2 (N1429, N1420, N1353);
nand NAND2 (N1430, N1426, N567);
buf BUF1 (N1431, N1421);
nor NOR3 (N1432, N1428, N690, N1110);
xor XOR2 (N1433, N1429, N826);
nand NAND4 (N1434, N1432, N930, N1396, N127);
and AND3 (N1435, N1423, N701, N857);
buf BUF1 (N1436, N1435);
not NOT1 (N1437, N1425);
xor XOR2 (N1438, N1416, N1095);
not NOT1 (N1439, N1437);
and AND4 (N1440, N1436, N914, N838, N309);
or OR3 (N1441, N1418, N798, N463);
and AND3 (N1442, N1441, N1209, N907);
buf BUF1 (N1443, N1430);
nand NAND2 (N1444, N1419, N1436);
not NOT1 (N1445, N1434);
and AND2 (N1446, N1438, N462);
not NOT1 (N1447, N1442);
nor NOR3 (N1448, N1424, N816, N425);
buf BUF1 (N1449, N1446);
xor XOR2 (N1450, N1443, N472);
not NOT1 (N1451, N1445);
buf BUF1 (N1452, N1433);
not NOT1 (N1453, N1448);
xor XOR2 (N1454, N1440, N1070);
xor XOR2 (N1455, N1439, N1247);
nor NOR4 (N1456, N1452, N17, N1271, N642);
or OR4 (N1457, N1453, N541, N449, N1022);
or OR3 (N1458, N1449, N843, N688);
nand NAND2 (N1459, N1444, N88);
xor XOR2 (N1460, N1454, N1202);
or OR2 (N1461, N1431, N842);
or OR2 (N1462, N1459, N1132);
and AND2 (N1463, N1455, N540);
not NOT1 (N1464, N1462);
xor XOR2 (N1465, N1464, N466);
and AND4 (N1466, N1458, N820, N601, N1339);
not NOT1 (N1467, N1466);
or OR3 (N1468, N1447, N132, N27);
nand NAND4 (N1469, N1460, N1062, N1071, N506);
or OR4 (N1470, N1467, N292, N867, N928);
not NOT1 (N1471, N1465);
and AND3 (N1472, N1470, N481, N979);
not NOT1 (N1473, N1463);
or OR2 (N1474, N1451, N1075);
and AND4 (N1475, N1469, N821, N1152, N1391);
xor XOR2 (N1476, N1471, N867);
buf BUF1 (N1477, N1472);
xor XOR2 (N1478, N1450, N1315);
nand NAND2 (N1479, N1477, N1211);
and AND2 (N1480, N1474, N1223);
and AND4 (N1481, N1457, N1299, N1344, N830);
nor NOR3 (N1482, N1468, N1191, N425);
buf BUF1 (N1483, N1475);
nand NAND2 (N1484, N1481, N739);
nor NOR2 (N1485, N1478, N567);
buf BUF1 (N1486, N1461);
nor NOR4 (N1487, N1473, N613, N902, N598);
nand NAND4 (N1488, N1484, N1415, N181, N984);
not NOT1 (N1489, N1487);
buf BUF1 (N1490, N1482);
not NOT1 (N1491, N1483);
xor XOR2 (N1492, N1480, N1259);
nor NOR2 (N1493, N1476, N1280);
buf BUF1 (N1494, N1492);
buf BUF1 (N1495, N1485);
or OR2 (N1496, N1494, N715);
nor NOR2 (N1497, N1456, N1155);
nand NAND2 (N1498, N1479, N447);
and AND2 (N1499, N1497, N740);
or OR3 (N1500, N1495, N1227, N507);
or OR2 (N1501, N1491, N1028);
buf BUF1 (N1502, N1496);
buf BUF1 (N1503, N1490);
or OR2 (N1504, N1501, N791);
xor XOR2 (N1505, N1486, N907);
or OR2 (N1506, N1500, N1130);
nand NAND3 (N1507, N1502, N1113, N905);
and AND4 (N1508, N1499, N443, N955, N345);
buf BUF1 (N1509, N1504);
or OR3 (N1510, N1503, N1365, N1296);
nor NOR4 (N1511, N1509, N389, N226, N1485);
or OR2 (N1512, N1507, N1051);
or OR4 (N1513, N1505, N1267, N1079, N1256);
buf BUF1 (N1514, N1513);
or OR3 (N1515, N1514, N330, N414);
not NOT1 (N1516, N1510);
buf BUF1 (N1517, N1512);
not NOT1 (N1518, N1511);
not NOT1 (N1519, N1493);
nor NOR2 (N1520, N1506, N674);
xor XOR2 (N1521, N1498, N1130);
and AND3 (N1522, N1519, N13, N1024);
endmodule