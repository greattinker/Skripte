// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11;

output N2003,N2007,N2010,N2000,N2005,N1998,N1999,N2009,N2006,N2011;

or OR3 (N12, N9, N6, N6);
xor XOR2 (N13, N5, N4);
or OR2 (N14, N1, N4);
not NOT1 (N15, N11);
nor NOR4 (N16, N8, N15, N13, N8);
and AND3 (N17, N5, N9, N3);
and AND4 (N18, N14, N2, N3, N2);
or OR2 (N19, N13, N7);
and AND4 (N20, N13, N17, N16, N19);
or OR4 (N21, N10, N16, N2, N10);
xor XOR2 (N22, N3, N16);
nand NAND2 (N23, N8, N2);
nor NOR2 (N24, N12, N17);
nor NOR2 (N25, N10, N5);
buf BUF1 (N26, N15);
buf BUF1 (N27, N15);
nor NOR3 (N28, N2, N14, N3);
buf BUF1 (N29, N25);
buf BUF1 (N30, N21);
and AND3 (N31, N18, N22, N2);
nor NOR3 (N32, N4, N18, N18);
buf BUF1 (N33, N24);
or OR2 (N34, N30, N12);
or OR4 (N35, N20, N22, N26, N1);
and AND3 (N36, N30, N20, N8);
or OR4 (N37, N23, N2, N16, N3);
nor NOR3 (N38, N36, N10, N31);
not NOT1 (N39, N22);
nor NOR3 (N40, N34, N28, N23);
not NOT1 (N41, N4);
nor NOR3 (N42, N27, N16, N26);
and AND4 (N43, N35, N8, N6, N36);
nand NAND4 (N44, N38, N17, N4, N24);
or OR2 (N45, N43, N1);
nor NOR3 (N46, N40, N28, N36);
and AND4 (N47, N46, N10, N37, N36);
xor XOR2 (N48, N38, N45);
and AND3 (N49, N23, N21, N35);
or OR3 (N50, N48, N25, N8);
nor NOR2 (N51, N47, N20);
nand NAND3 (N52, N41, N16, N43);
not NOT1 (N53, N52);
xor XOR2 (N54, N32, N39);
nor NOR3 (N55, N49, N11, N40);
nand NAND3 (N56, N52, N47, N43);
buf BUF1 (N57, N33);
not NOT1 (N58, N56);
nor NOR3 (N59, N50, N18, N35);
xor XOR2 (N60, N54, N2);
nor NOR4 (N61, N58, N28, N33, N46);
not NOT1 (N62, N59);
xor XOR2 (N63, N42, N7);
and AND3 (N64, N29, N50, N39);
or OR2 (N65, N44, N25);
nor NOR2 (N66, N53, N58);
buf BUF1 (N67, N63);
nor NOR4 (N68, N60, N12, N65, N55);
nand NAND2 (N69, N5, N20);
or OR2 (N70, N69, N19);
not NOT1 (N71, N32);
buf BUF1 (N72, N71);
not NOT1 (N73, N62);
and AND2 (N74, N51, N48);
nand NAND3 (N75, N74, N26, N68);
nand NAND4 (N76, N61, N69, N33, N14);
xor XOR2 (N77, N21, N2);
nor NOR3 (N78, N75, N1, N67);
buf BUF1 (N79, N29);
buf BUF1 (N80, N70);
and AND4 (N81, N77, N2, N14, N9);
or OR3 (N82, N66, N50, N35);
buf BUF1 (N83, N64);
and AND2 (N84, N82, N67);
nand NAND3 (N85, N80, N46, N71);
xor XOR2 (N86, N57, N78);
or OR3 (N87, N20, N57, N50);
buf BUF1 (N88, N87);
buf BUF1 (N89, N79);
xor XOR2 (N90, N83, N23);
and AND3 (N91, N72, N77, N80);
buf BUF1 (N92, N81);
nor NOR4 (N93, N85, N39, N38, N90);
and AND3 (N94, N25, N86, N32);
nand NAND2 (N95, N62, N52);
and AND3 (N96, N91, N79, N86);
not NOT1 (N97, N76);
or OR2 (N98, N89, N2);
nand NAND4 (N99, N94, N26, N34, N82);
nor NOR3 (N100, N95, N10, N11);
or OR2 (N101, N84, N83);
or OR3 (N102, N92, N14, N89);
buf BUF1 (N103, N101);
xor XOR2 (N104, N73, N93);
nand NAND4 (N105, N17, N57, N60, N61);
xor XOR2 (N106, N100, N47);
nor NOR2 (N107, N98, N100);
nor NOR4 (N108, N102, N7, N34, N67);
buf BUF1 (N109, N96);
buf BUF1 (N110, N88);
nand NAND4 (N111, N99, N15, N100, N69);
nor NOR4 (N112, N97, N90, N45, N70);
nand NAND2 (N113, N110, N111);
not NOT1 (N114, N17);
nor NOR4 (N115, N103, N91, N46, N86);
nor NOR2 (N116, N104, N99);
nor NOR3 (N117, N113, N66, N19);
nand NAND4 (N118, N117, N43, N28, N90);
not NOT1 (N119, N114);
nor NOR4 (N120, N118, N45, N20, N55);
and AND2 (N121, N119, N31);
nand NAND3 (N122, N106, N26, N67);
nand NAND4 (N123, N112, N35, N121, N2);
or OR4 (N124, N87, N117, N71, N54);
not NOT1 (N125, N108);
nor NOR3 (N126, N120, N51, N87);
or OR3 (N127, N126, N19, N1);
buf BUF1 (N128, N122);
xor XOR2 (N129, N125, N71);
buf BUF1 (N130, N124);
nor NOR3 (N131, N105, N86, N59);
xor XOR2 (N132, N129, N92);
buf BUF1 (N133, N130);
and AND2 (N134, N133, N46);
and AND3 (N135, N132, N63, N48);
nor NOR2 (N136, N109, N74);
xor XOR2 (N137, N134, N70);
xor XOR2 (N138, N135, N107);
not NOT1 (N139, N29);
or OR4 (N140, N123, N21, N93, N104);
nand NAND3 (N141, N127, N84, N54);
nand NAND2 (N142, N131, N135);
nand NAND3 (N143, N128, N66, N85);
and AND4 (N144, N142, N31, N67, N53);
nor NOR3 (N145, N138, N16, N73);
nand NAND2 (N146, N136, N79);
xor XOR2 (N147, N141, N57);
xor XOR2 (N148, N139, N88);
not NOT1 (N149, N116);
and AND3 (N150, N146, N100, N148);
nand NAND3 (N151, N133, N26, N59);
nand NAND4 (N152, N143, N135, N27, N60);
nand NAND3 (N153, N140, N144, N103);
not NOT1 (N154, N99);
or OR3 (N155, N151, N128, N55);
xor XOR2 (N156, N153, N50);
xor XOR2 (N157, N115, N14);
buf BUF1 (N158, N150);
xor XOR2 (N159, N145, N56);
xor XOR2 (N160, N155, N106);
xor XOR2 (N161, N154, N19);
nand NAND4 (N162, N137, N97, N149, N119);
or OR2 (N163, N131, N70);
not NOT1 (N164, N160);
nand NAND3 (N165, N157, N162, N59);
buf BUF1 (N166, N135);
buf BUF1 (N167, N163);
not NOT1 (N168, N156);
buf BUF1 (N169, N158);
nand NAND2 (N170, N166, N55);
nand NAND2 (N171, N164, N109);
buf BUF1 (N172, N167);
nand NAND3 (N173, N159, N101, N47);
nand NAND3 (N174, N152, N112, N159);
nand NAND2 (N175, N165, N28);
not NOT1 (N176, N174);
nand NAND3 (N177, N175, N135, N106);
and AND3 (N178, N168, N19, N153);
nor NOR4 (N179, N176, N11, N127, N93);
buf BUF1 (N180, N170);
xor XOR2 (N181, N172, N152);
nor NOR3 (N182, N171, N84, N52);
nor NOR3 (N183, N181, N100, N61);
not NOT1 (N184, N173);
buf BUF1 (N185, N179);
xor XOR2 (N186, N184, N178);
buf BUF1 (N187, N28);
not NOT1 (N188, N187);
buf BUF1 (N189, N180);
not NOT1 (N190, N186);
or OR4 (N191, N188, N37, N114, N129);
nand NAND4 (N192, N191, N100, N161, N29);
xor XOR2 (N193, N91, N115);
xor XOR2 (N194, N193, N186);
buf BUF1 (N195, N183);
nand NAND4 (N196, N177, N163, N7, N176);
buf BUF1 (N197, N189);
nand NAND4 (N198, N194, N27, N58, N102);
and AND3 (N199, N196, N89, N178);
and AND3 (N200, N185, N30, N52);
not NOT1 (N201, N190);
not NOT1 (N202, N192);
buf BUF1 (N203, N199);
and AND2 (N204, N200, N192);
or OR2 (N205, N201, N169);
nand NAND3 (N206, N40, N50, N78);
nor NOR4 (N207, N198, N30, N96, N85);
or OR4 (N208, N206, N15, N177, N81);
and AND3 (N209, N195, N111, N39);
buf BUF1 (N210, N208);
xor XOR2 (N211, N147, N164);
and AND3 (N212, N211, N154, N128);
nand NAND2 (N213, N204, N116);
nor NOR4 (N214, N182, N56, N177, N70);
not NOT1 (N215, N210);
buf BUF1 (N216, N202);
and AND2 (N217, N216, N137);
buf BUF1 (N218, N203);
or OR4 (N219, N218, N199, N153, N125);
nand NAND2 (N220, N212, N198);
xor XOR2 (N221, N215, N183);
nor NOR4 (N222, N214, N159, N201, N122);
buf BUF1 (N223, N217);
and AND2 (N224, N207, N73);
nand NAND3 (N225, N205, N187, N57);
nor NOR2 (N226, N220, N6);
buf BUF1 (N227, N197);
buf BUF1 (N228, N227);
nor NOR3 (N229, N223, N11, N153);
nand NAND2 (N230, N228, N137);
or OR2 (N231, N213, N66);
or OR3 (N232, N209, N51, N9);
nand NAND3 (N233, N226, N213, N107);
nor NOR4 (N234, N230, N114, N197, N66);
and AND3 (N235, N231, N89, N221);
not NOT1 (N236, N62);
nor NOR2 (N237, N224, N101);
buf BUF1 (N238, N235);
not NOT1 (N239, N219);
nand NAND4 (N240, N238, N198, N129, N44);
nor NOR4 (N241, N229, N24, N190, N79);
nand NAND3 (N242, N222, N54, N88);
not NOT1 (N243, N242);
xor XOR2 (N244, N236, N192);
xor XOR2 (N245, N239, N163);
and AND2 (N246, N243, N145);
or OR3 (N247, N232, N118, N178);
nor NOR2 (N248, N234, N113);
nand NAND3 (N249, N237, N110, N168);
not NOT1 (N250, N225);
and AND2 (N251, N244, N65);
nand NAND2 (N252, N241, N151);
nand NAND4 (N253, N240, N96, N36, N142);
nand NAND4 (N254, N248, N186, N41, N120);
buf BUF1 (N255, N254);
xor XOR2 (N256, N246, N102);
or OR2 (N257, N247, N117);
not NOT1 (N258, N251);
and AND4 (N259, N255, N237, N57, N120);
not NOT1 (N260, N257);
or OR3 (N261, N258, N54, N106);
buf BUF1 (N262, N261);
xor XOR2 (N263, N256, N184);
and AND3 (N264, N250, N245, N6);
nor NOR3 (N265, N22, N83, N26);
not NOT1 (N266, N253);
or OR4 (N267, N265, N185, N34, N39);
xor XOR2 (N268, N233, N87);
nand NAND3 (N269, N260, N22, N65);
xor XOR2 (N270, N267, N139);
nor NOR4 (N271, N270, N240, N55, N170);
xor XOR2 (N272, N262, N74);
and AND4 (N273, N259, N85, N192, N144);
and AND2 (N274, N268, N116);
or OR2 (N275, N266, N70);
buf BUF1 (N276, N271);
and AND3 (N277, N252, N187, N193);
not NOT1 (N278, N264);
nand NAND2 (N279, N263, N73);
and AND2 (N280, N276, N168);
or OR4 (N281, N277, N103, N202, N161);
xor XOR2 (N282, N273, N22);
buf BUF1 (N283, N274);
not NOT1 (N284, N278);
nand NAND2 (N285, N279, N77);
nor NOR2 (N286, N249, N196);
nand NAND2 (N287, N284, N132);
nand NAND4 (N288, N282, N66, N30, N79);
xor XOR2 (N289, N275, N148);
buf BUF1 (N290, N287);
nand NAND3 (N291, N288, N238, N216);
nand NAND2 (N292, N281, N111);
or OR4 (N293, N272, N225, N286, N87);
and AND3 (N294, N124, N255, N193);
buf BUF1 (N295, N292);
nand NAND2 (N296, N289, N128);
and AND4 (N297, N295, N270, N288, N62);
or OR4 (N298, N285, N255, N185, N213);
or OR2 (N299, N290, N239);
not NOT1 (N300, N298);
or OR2 (N301, N300, N278);
or OR2 (N302, N293, N162);
or OR3 (N303, N296, N169, N235);
buf BUF1 (N304, N269);
nand NAND4 (N305, N294, N127, N83, N204);
nor NOR4 (N306, N283, N223, N242, N177);
not NOT1 (N307, N302);
or OR4 (N308, N304, N203, N65, N38);
not NOT1 (N309, N305);
or OR4 (N310, N308, N192, N228, N115);
nand NAND4 (N311, N291, N6, N142, N32);
buf BUF1 (N312, N310);
or OR3 (N313, N301, N297, N133);
nor NOR3 (N314, N280, N213, N29);
buf BUF1 (N315, N271);
nand NAND2 (N316, N309, N41);
nor NOR3 (N317, N303, N124, N24);
or OR3 (N318, N315, N117, N164);
not NOT1 (N319, N317);
or OR2 (N320, N306, N208);
and AND3 (N321, N312, N84, N185);
xor XOR2 (N322, N311, N13);
xor XOR2 (N323, N322, N104);
nor NOR4 (N324, N307, N72, N299, N7);
nor NOR4 (N325, N315, N154, N252, N288);
and AND3 (N326, N319, N59, N287);
or OR3 (N327, N314, N94, N193);
or OR3 (N328, N326, N72, N283);
xor XOR2 (N329, N316, N73);
xor XOR2 (N330, N327, N218);
xor XOR2 (N331, N325, N141);
nand NAND3 (N332, N328, N60, N218);
xor XOR2 (N333, N321, N29);
or OR3 (N334, N323, N61, N331);
and AND3 (N335, N270, N185, N309);
buf BUF1 (N336, N320);
buf BUF1 (N337, N333);
or OR3 (N338, N334, N281, N45);
or OR2 (N339, N329, N64);
nand NAND3 (N340, N336, N323, N270);
xor XOR2 (N341, N332, N279);
buf BUF1 (N342, N337);
or OR2 (N343, N335, N114);
or OR3 (N344, N324, N334, N158);
and AND4 (N345, N338, N206, N60, N173);
not NOT1 (N346, N342);
nand NAND3 (N347, N318, N331, N123);
nor NOR2 (N348, N313, N87);
not NOT1 (N349, N341);
xor XOR2 (N350, N339, N317);
not NOT1 (N351, N343);
not NOT1 (N352, N340);
nor NOR4 (N353, N347, N181, N73, N93);
nand NAND3 (N354, N348, N67, N265);
not NOT1 (N355, N349);
or OR3 (N356, N353, N184, N178);
and AND3 (N357, N344, N313, N234);
and AND2 (N358, N357, N114);
nand NAND4 (N359, N351, N305, N245, N276);
and AND3 (N360, N356, N124, N84);
and AND3 (N361, N355, N4, N261);
or OR4 (N362, N350, N318, N146, N54);
and AND3 (N363, N354, N120, N178);
nor NOR2 (N364, N352, N273);
and AND3 (N365, N360, N233, N348);
and AND4 (N366, N362, N83, N52, N219);
buf BUF1 (N367, N365);
nand NAND4 (N368, N366, N98, N142, N219);
nand NAND2 (N369, N368, N241);
xor XOR2 (N370, N346, N189);
xor XOR2 (N371, N359, N106);
not NOT1 (N372, N370);
nor NOR3 (N373, N345, N342, N111);
buf BUF1 (N374, N367);
or OR4 (N375, N364, N73, N39, N99);
not NOT1 (N376, N371);
xor XOR2 (N377, N375, N108);
nand NAND3 (N378, N377, N218, N147);
xor XOR2 (N379, N358, N113);
xor XOR2 (N380, N373, N159);
nor NOR3 (N381, N379, N103, N313);
nand NAND4 (N382, N374, N128, N274, N90);
and AND3 (N383, N382, N41, N244);
xor XOR2 (N384, N383, N82);
or OR4 (N385, N363, N135, N366, N283);
xor XOR2 (N386, N385, N82);
nor NOR3 (N387, N361, N64, N143);
and AND3 (N388, N387, N355, N273);
or OR3 (N389, N376, N87, N9);
or OR2 (N390, N380, N170);
and AND4 (N391, N330, N32, N386, N6);
and AND3 (N392, N381, N295, N296);
nor NOR3 (N393, N220, N174, N379);
or OR3 (N394, N391, N278, N138);
and AND2 (N395, N372, N195);
buf BUF1 (N396, N395);
and AND4 (N397, N392, N222, N207, N69);
or OR2 (N398, N393, N333);
nor NOR3 (N399, N384, N255, N388);
xor XOR2 (N400, N138, N138);
buf BUF1 (N401, N396);
buf BUF1 (N402, N401);
and AND3 (N403, N402, N22, N161);
buf BUF1 (N404, N378);
not NOT1 (N405, N404);
nand NAND2 (N406, N369, N136);
not NOT1 (N407, N398);
not NOT1 (N408, N397);
or OR3 (N409, N389, N56, N314);
and AND3 (N410, N399, N51, N22);
buf BUF1 (N411, N408);
nand NAND4 (N412, N406, N14, N150, N404);
xor XOR2 (N413, N407, N171);
not NOT1 (N414, N413);
or OR4 (N415, N403, N376, N113, N184);
and AND2 (N416, N409, N82);
buf BUF1 (N417, N394);
nand NAND2 (N418, N412, N93);
buf BUF1 (N419, N410);
buf BUF1 (N420, N418);
not NOT1 (N421, N414);
nor NOR4 (N422, N421, N298, N297, N94);
and AND2 (N423, N415, N230);
nand NAND2 (N424, N390, N42);
nor NOR3 (N425, N417, N417, N270);
xor XOR2 (N426, N424, N256);
not NOT1 (N427, N423);
buf BUF1 (N428, N426);
or OR2 (N429, N422, N358);
nand NAND2 (N430, N416, N350);
and AND4 (N431, N425, N196, N309, N22);
buf BUF1 (N432, N405);
not NOT1 (N433, N411);
not NOT1 (N434, N429);
nor NOR2 (N435, N400, N41);
xor XOR2 (N436, N420, N358);
nor NOR4 (N437, N435, N164, N116, N436);
or OR2 (N438, N223, N427);
buf BUF1 (N439, N266);
nor NOR4 (N440, N428, N176, N31, N140);
not NOT1 (N441, N434);
or OR2 (N442, N432, N233);
nor NOR3 (N443, N433, N442, N390);
xor XOR2 (N444, N414, N312);
buf BUF1 (N445, N430);
nor NOR4 (N446, N437, N20, N314, N368);
nand NAND2 (N447, N445, N364);
nor NOR3 (N448, N446, N35, N56);
not NOT1 (N449, N431);
buf BUF1 (N450, N443);
or OR3 (N451, N448, N176, N167);
not NOT1 (N452, N419);
xor XOR2 (N453, N440, N409);
xor XOR2 (N454, N439, N372);
xor XOR2 (N455, N438, N58);
and AND3 (N456, N441, N437, N331);
and AND3 (N457, N454, N157, N27);
or OR3 (N458, N455, N78, N435);
not NOT1 (N459, N444);
buf BUF1 (N460, N459);
nand NAND4 (N461, N453, N77, N347, N79);
and AND2 (N462, N452, N122);
xor XOR2 (N463, N461, N89);
buf BUF1 (N464, N450);
nor NOR3 (N465, N462, N154, N402);
nand NAND4 (N466, N460, N159, N172, N262);
xor XOR2 (N467, N458, N384);
and AND4 (N468, N456, N288, N302, N405);
or OR2 (N469, N451, N112);
nor NOR3 (N470, N464, N189, N278);
xor XOR2 (N471, N457, N446);
or OR3 (N472, N469, N206, N157);
or OR4 (N473, N472, N11, N296, N120);
nor NOR3 (N474, N473, N194, N39);
or OR4 (N475, N470, N48, N449, N164);
nor NOR2 (N476, N335, N130);
xor XOR2 (N477, N465, N323);
or OR4 (N478, N477, N362, N31, N348);
or OR3 (N479, N476, N247, N245);
nor NOR4 (N480, N471, N376, N409, N416);
nand NAND4 (N481, N478, N226, N351, N329);
xor XOR2 (N482, N479, N156);
nand NAND2 (N483, N468, N19);
nand NAND3 (N484, N483, N56, N399);
and AND4 (N485, N467, N426, N351, N235);
and AND3 (N486, N447, N100, N264);
nor NOR2 (N487, N463, N158);
and AND3 (N488, N482, N366, N265);
xor XOR2 (N489, N480, N69);
not NOT1 (N490, N487);
and AND2 (N491, N474, N40);
not NOT1 (N492, N490);
or OR4 (N493, N466, N87, N382, N248);
buf BUF1 (N494, N493);
and AND3 (N495, N494, N22, N29);
xor XOR2 (N496, N484, N152);
xor XOR2 (N497, N485, N70);
or OR4 (N498, N496, N444, N341, N425);
not NOT1 (N499, N491);
buf BUF1 (N500, N497);
and AND4 (N501, N498, N439, N121, N19);
nor NOR4 (N502, N475, N46, N85, N20);
or OR3 (N503, N486, N450, N406);
xor XOR2 (N504, N500, N326);
nand NAND4 (N505, N501, N364, N352, N302);
buf BUF1 (N506, N499);
or OR4 (N507, N503, N316, N169, N411);
nor NOR3 (N508, N492, N455, N91);
and AND3 (N509, N495, N278, N42);
and AND2 (N510, N509, N39);
buf BUF1 (N511, N510);
nor NOR2 (N512, N506, N30);
xor XOR2 (N513, N489, N274);
and AND2 (N514, N512, N271);
buf BUF1 (N515, N504);
buf BUF1 (N516, N511);
and AND3 (N517, N513, N131, N422);
buf BUF1 (N518, N515);
xor XOR2 (N519, N502, N349);
xor XOR2 (N520, N518, N346);
and AND2 (N521, N516, N307);
not NOT1 (N522, N481);
xor XOR2 (N523, N488, N446);
or OR4 (N524, N507, N85, N211, N278);
and AND4 (N525, N524, N351, N31, N445);
not NOT1 (N526, N514);
or OR2 (N527, N505, N247);
and AND3 (N528, N508, N206, N368);
xor XOR2 (N529, N521, N371);
buf BUF1 (N530, N527);
and AND3 (N531, N519, N107, N342);
nor NOR3 (N532, N530, N185, N48);
nand NAND3 (N533, N517, N125, N78);
or OR4 (N534, N531, N134, N25, N521);
or OR3 (N535, N534, N458, N494);
and AND3 (N536, N532, N510, N102);
and AND4 (N537, N526, N474, N15, N111);
or OR2 (N538, N522, N115);
nand NAND4 (N539, N538, N17, N327, N440);
xor XOR2 (N540, N535, N53);
nand NAND4 (N541, N540, N403, N125, N271);
nor NOR2 (N542, N537, N219);
buf BUF1 (N543, N529);
not NOT1 (N544, N543);
not NOT1 (N545, N528);
nor NOR4 (N546, N544, N445, N114, N214);
buf BUF1 (N547, N533);
and AND4 (N548, N539, N141, N54, N108);
nand NAND3 (N549, N546, N326, N349);
nand NAND2 (N550, N520, N440);
or OR4 (N551, N547, N30, N221, N35);
xor XOR2 (N552, N541, N23);
nor NOR4 (N553, N536, N466, N530, N29);
and AND2 (N554, N523, N69);
buf BUF1 (N555, N554);
nor NOR3 (N556, N549, N352, N48);
not NOT1 (N557, N551);
and AND4 (N558, N553, N84, N156, N213);
nor NOR4 (N559, N545, N501, N154, N544);
and AND3 (N560, N550, N379, N5);
nand NAND4 (N561, N558, N117, N8, N10);
xor XOR2 (N562, N542, N279);
not NOT1 (N563, N525);
nor NOR2 (N564, N562, N514);
nor NOR4 (N565, N552, N292, N539, N69);
nor NOR3 (N566, N561, N353, N251);
and AND4 (N567, N563, N440, N343, N515);
nor NOR2 (N568, N556, N21);
or OR2 (N569, N565, N353);
nand NAND4 (N570, N548, N149, N40, N75);
buf BUF1 (N571, N567);
xor XOR2 (N572, N571, N68);
not NOT1 (N573, N568);
or OR3 (N574, N566, N376, N104);
or OR3 (N575, N555, N419, N416);
not NOT1 (N576, N557);
xor XOR2 (N577, N576, N250);
not NOT1 (N578, N570);
nand NAND2 (N579, N559, N57);
and AND2 (N580, N577, N442);
or OR2 (N581, N569, N409);
or OR2 (N582, N572, N111);
not NOT1 (N583, N574);
xor XOR2 (N584, N564, N463);
and AND4 (N585, N581, N373, N362, N584);
and AND2 (N586, N512, N304);
and AND3 (N587, N582, N544, N115);
buf BUF1 (N588, N586);
and AND3 (N589, N583, N18, N96);
and AND4 (N590, N573, N556, N323, N492);
xor XOR2 (N591, N590, N378);
buf BUF1 (N592, N575);
nand NAND2 (N593, N585, N250);
or OR3 (N594, N593, N381, N548);
or OR3 (N595, N592, N180, N233);
xor XOR2 (N596, N580, N405);
xor XOR2 (N597, N587, N349);
xor XOR2 (N598, N595, N340);
and AND2 (N599, N589, N3);
nand NAND3 (N600, N598, N216, N121);
buf BUF1 (N601, N599);
not NOT1 (N602, N601);
xor XOR2 (N603, N591, N169);
buf BUF1 (N604, N597);
buf BUF1 (N605, N604);
not NOT1 (N606, N605);
nand NAND3 (N607, N594, N226, N384);
not NOT1 (N608, N600);
or OR3 (N609, N596, N577, N242);
not NOT1 (N610, N608);
or OR2 (N611, N578, N69);
buf BUF1 (N612, N607);
or OR3 (N613, N606, N131, N365);
buf BUF1 (N614, N612);
and AND4 (N615, N602, N345, N94, N527);
or OR2 (N616, N603, N160);
nor NOR2 (N617, N613, N244);
buf BUF1 (N618, N579);
nand NAND3 (N619, N616, N24, N165);
xor XOR2 (N620, N618, N117);
nor NOR4 (N621, N609, N547, N167, N350);
not NOT1 (N622, N610);
nor NOR3 (N623, N622, N197, N319);
or OR3 (N624, N619, N608, N612);
buf BUF1 (N625, N624);
or OR3 (N626, N588, N249, N566);
and AND3 (N627, N621, N256, N366);
or OR4 (N628, N614, N47, N449, N355);
buf BUF1 (N629, N625);
xor XOR2 (N630, N620, N605);
not NOT1 (N631, N627);
xor XOR2 (N632, N623, N447);
nand NAND4 (N633, N629, N277, N627, N41);
and AND4 (N634, N632, N460, N14, N50);
buf BUF1 (N635, N628);
not NOT1 (N636, N635);
nand NAND3 (N637, N615, N48, N153);
nor NOR3 (N638, N636, N535, N95);
or OR4 (N639, N638, N384, N253, N231);
nor NOR4 (N640, N630, N469, N349, N537);
nand NAND3 (N641, N633, N621, N448);
and AND2 (N642, N617, N591);
xor XOR2 (N643, N626, N89);
xor XOR2 (N644, N631, N138);
xor XOR2 (N645, N642, N246);
nand NAND2 (N646, N644, N91);
and AND4 (N647, N637, N437, N95, N474);
nand NAND4 (N648, N611, N224, N605, N265);
buf BUF1 (N649, N641);
or OR4 (N650, N639, N68, N102, N364);
xor XOR2 (N651, N647, N228);
nand NAND3 (N652, N640, N501, N494);
not NOT1 (N653, N649);
nor NOR3 (N654, N650, N84, N236);
xor XOR2 (N655, N648, N167);
nand NAND3 (N656, N634, N310, N59);
nand NAND2 (N657, N655, N229);
buf BUF1 (N658, N657);
nor NOR2 (N659, N645, N285);
or OR2 (N660, N652, N296);
nand NAND4 (N661, N643, N136, N637, N250);
and AND4 (N662, N656, N652, N450, N62);
xor XOR2 (N663, N646, N52);
or OR2 (N664, N653, N217);
not NOT1 (N665, N658);
xor XOR2 (N666, N560, N178);
or OR4 (N667, N654, N135, N425, N15);
or OR3 (N668, N664, N459, N239);
nand NAND4 (N669, N668, N20, N608, N627);
buf BUF1 (N670, N660);
or OR3 (N671, N663, N284, N54);
not NOT1 (N672, N659);
buf BUF1 (N673, N661);
or OR3 (N674, N672, N162, N503);
or OR3 (N675, N673, N69, N254);
nor NOR4 (N676, N669, N628, N369, N634);
buf BUF1 (N677, N667);
buf BUF1 (N678, N670);
nand NAND2 (N679, N675, N521);
nor NOR4 (N680, N676, N32, N196, N60);
and AND4 (N681, N666, N415, N137, N363);
buf BUF1 (N682, N671);
nor NOR4 (N683, N677, N582, N527, N197);
not NOT1 (N684, N651);
nor NOR4 (N685, N680, N46, N117, N515);
not NOT1 (N686, N685);
buf BUF1 (N687, N686);
not NOT1 (N688, N674);
xor XOR2 (N689, N687, N128);
not NOT1 (N690, N688);
nand NAND4 (N691, N662, N375, N337, N222);
and AND4 (N692, N679, N118, N476, N261);
and AND2 (N693, N681, N46);
buf BUF1 (N694, N693);
not NOT1 (N695, N692);
buf BUF1 (N696, N695);
not NOT1 (N697, N691);
not NOT1 (N698, N682);
nor NOR4 (N699, N683, N647, N643, N396);
nand NAND4 (N700, N698, N525, N637, N68);
buf BUF1 (N701, N700);
nor NOR3 (N702, N678, N524, N74);
nor NOR3 (N703, N684, N463, N656);
nand NAND3 (N704, N699, N609, N72);
nand NAND4 (N705, N697, N617, N121, N229);
nand NAND4 (N706, N704, N442, N652, N462);
xor XOR2 (N707, N690, N24);
nand NAND3 (N708, N696, N612, N400);
or OR2 (N709, N707, N360);
buf BUF1 (N710, N689);
nor NOR3 (N711, N665, N142, N57);
nand NAND2 (N712, N694, N325);
and AND3 (N713, N712, N172, N611);
nand NAND4 (N714, N709, N340, N117, N471);
not NOT1 (N715, N713);
buf BUF1 (N716, N715);
nor NOR4 (N717, N711, N611, N315, N125);
and AND2 (N718, N705, N689);
nand NAND4 (N719, N703, N609, N27, N284);
xor XOR2 (N720, N706, N59);
nand NAND4 (N721, N701, N330, N499, N19);
not NOT1 (N722, N702);
nand NAND4 (N723, N721, N396, N621, N226);
and AND2 (N724, N714, N306);
nor NOR4 (N725, N722, N453, N621, N584);
or OR2 (N726, N717, N65);
or OR2 (N727, N710, N622);
not NOT1 (N728, N724);
or OR2 (N729, N708, N275);
and AND3 (N730, N718, N138, N482);
xor XOR2 (N731, N728, N295);
nor NOR2 (N732, N730, N8);
buf BUF1 (N733, N725);
xor XOR2 (N734, N731, N373);
buf BUF1 (N735, N726);
xor XOR2 (N736, N734, N220);
nand NAND3 (N737, N732, N136, N190);
buf BUF1 (N738, N737);
or OR2 (N739, N719, N168);
and AND4 (N740, N729, N117, N497, N241);
or OR4 (N741, N739, N305, N554, N337);
nor NOR2 (N742, N736, N279);
nor NOR2 (N743, N742, N118);
or OR4 (N744, N716, N332, N628, N217);
nor NOR4 (N745, N735, N716, N467, N405);
nand NAND3 (N746, N743, N309, N15);
buf BUF1 (N747, N744);
nor NOR2 (N748, N723, N381);
xor XOR2 (N749, N741, N598);
nor NOR2 (N750, N733, N33);
xor XOR2 (N751, N745, N471);
xor XOR2 (N752, N720, N217);
not NOT1 (N753, N747);
xor XOR2 (N754, N752, N317);
and AND2 (N755, N738, N596);
nand NAND3 (N756, N749, N451, N533);
buf BUF1 (N757, N751);
xor XOR2 (N758, N727, N571);
not NOT1 (N759, N740);
not NOT1 (N760, N750);
and AND4 (N761, N757, N728, N532, N473);
nand NAND4 (N762, N754, N57, N666, N211);
buf BUF1 (N763, N756);
buf BUF1 (N764, N763);
nand NAND4 (N765, N748, N436, N622, N226);
or OR2 (N766, N764, N367);
not NOT1 (N767, N759);
and AND3 (N768, N755, N669, N82);
buf BUF1 (N769, N766);
nor NOR4 (N770, N769, N257, N670, N333);
nor NOR3 (N771, N753, N552, N214);
or OR4 (N772, N762, N164, N570, N338);
nand NAND2 (N773, N767, N577);
or OR4 (N774, N768, N208, N52, N103);
buf BUF1 (N775, N771);
nor NOR4 (N776, N770, N609, N100, N629);
buf BUF1 (N777, N773);
nand NAND2 (N778, N760, N359);
not NOT1 (N779, N778);
and AND4 (N780, N779, N201, N646, N716);
not NOT1 (N781, N746);
nand NAND2 (N782, N775, N184);
buf BUF1 (N783, N765);
buf BUF1 (N784, N774);
xor XOR2 (N785, N782, N281);
xor XOR2 (N786, N783, N188);
nand NAND2 (N787, N780, N408);
xor XOR2 (N788, N761, N33);
nor NOR4 (N789, N788, N383, N152, N725);
xor XOR2 (N790, N772, N340);
or OR3 (N791, N758, N105, N670);
and AND3 (N792, N784, N313, N122);
nand NAND4 (N793, N792, N573, N779, N600);
xor XOR2 (N794, N791, N466);
buf BUF1 (N795, N794);
not NOT1 (N796, N787);
not NOT1 (N797, N793);
not NOT1 (N798, N795);
buf BUF1 (N799, N777);
or OR3 (N800, N785, N266, N95);
buf BUF1 (N801, N799);
not NOT1 (N802, N800);
and AND2 (N803, N781, N707);
nand NAND2 (N804, N798, N53);
and AND2 (N805, N802, N570);
buf BUF1 (N806, N805);
nand NAND3 (N807, N806, N725, N56);
nor NOR3 (N808, N789, N714, N651);
xor XOR2 (N809, N796, N22);
nand NAND4 (N810, N804, N104, N394, N128);
and AND2 (N811, N803, N642);
nand NAND4 (N812, N790, N9, N131, N429);
buf BUF1 (N813, N801);
buf BUF1 (N814, N811);
and AND2 (N815, N812, N494);
nor NOR4 (N816, N797, N295, N194, N502);
and AND3 (N817, N807, N89, N781);
nand NAND3 (N818, N816, N470, N460);
xor XOR2 (N819, N813, N814);
not NOT1 (N820, N305);
not NOT1 (N821, N809);
and AND3 (N822, N818, N299, N253);
nand NAND3 (N823, N822, N821, N103);
buf BUF1 (N824, N431);
or OR3 (N825, N815, N152, N51);
nand NAND3 (N826, N825, N72, N451);
nand NAND2 (N827, N808, N317);
buf BUF1 (N828, N819);
and AND2 (N829, N823, N419);
buf BUF1 (N830, N776);
xor XOR2 (N831, N810, N555);
xor XOR2 (N832, N826, N788);
nor NOR4 (N833, N832, N360, N391, N446);
or OR3 (N834, N827, N337, N293);
not NOT1 (N835, N828);
not NOT1 (N836, N835);
buf BUF1 (N837, N834);
nand NAND2 (N838, N833, N19);
or OR3 (N839, N837, N690, N466);
xor XOR2 (N840, N839, N58);
not NOT1 (N841, N840);
nand NAND3 (N842, N824, N701, N623);
and AND2 (N843, N836, N365);
and AND4 (N844, N843, N808, N790, N487);
or OR2 (N845, N838, N340);
not NOT1 (N846, N842);
or OR2 (N847, N820, N22);
not NOT1 (N848, N841);
nor NOR3 (N849, N830, N527, N302);
not NOT1 (N850, N829);
nor NOR2 (N851, N844, N314);
and AND3 (N852, N845, N389, N114);
not NOT1 (N853, N846);
buf BUF1 (N854, N817);
and AND2 (N855, N852, N25);
nand NAND2 (N856, N847, N688);
nand NAND3 (N857, N848, N801, N685);
xor XOR2 (N858, N849, N851);
not NOT1 (N859, N304);
buf BUF1 (N860, N853);
nand NAND3 (N861, N856, N267, N165);
or OR2 (N862, N850, N166);
not NOT1 (N863, N860);
buf BUF1 (N864, N863);
buf BUF1 (N865, N786);
nand NAND3 (N866, N864, N309, N178);
and AND3 (N867, N858, N178, N396);
or OR2 (N868, N862, N28);
or OR3 (N869, N857, N492, N862);
nand NAND4 (N870, N869, N38, N79, N767);
or OR3 (N871, N854, N72, N457);
or OR4 (N872, N831, N848, N294, N769);
buf BUF1 (N873, N855);
xor XOR2 (N874, N867, N1);
or OR2 (N875, N871, N849);
xor XOR2 (N876, N859, N89);
or OR3 (N877, N874, N686, N256);
nand NAND3 (N878, N866, N311, N852);
xor XOR2 (N879, N861, N676);
buf BUF1 (N880, N865);
and AND3 (N881, N873, N371, N183);
buf BUF1 (N882, N881);
and AND4 (N883, N870, N102, N160, N661);
nor NOR3 (N884, N880, N744, N170);
nor NOR4 (N885, N875, N342, N445, N419);
buf BUF1 (N886, N878);
and AND4 (N887, N882, N196, N767, N221);
xor XOR2 (N888, N872, N306);
xor XOR2 (N889, N887, N390);
not NOT1 (N890, N877);
nand NAND4 (N891, N884, N481, N185, N835);
nand NAND3 (N892, N883, N122, N311);
or OR2 (N893, N891, N211);
buf BUF1 (N894, N868);
nor NOR4 (N895, N879, N303, N398, N213);
and AND2 (N896, N888, N588);
nand NAND2 (N897, N885, N637);
nor NOR3 (N898, N890, N396, N735);
not NOT1 (N899, N898);
nand NAND2 (N900, N896, N710);
and AND2 (N901, N895, N2);
nor NOR4 (N902, N886, N268, N399, N344);
not NOT1 (N903, N899);
nand NAND2 (N904, N889, N70);
and AND2 (N905, N903, N147);
and AND4 (N906, N900, N314, N436, N474);
nand NAND2 (N907, N892, N114);
and AND2 (N908, N893, N476);
not NOT1 (N909, N906);
xor XOR2 (N910, N902, N239);
and AND2 (N911, N908, N622);
not NOT1 (N912, N901);
not NOT1 (N913, N909);
and AND4 (N914, N907, N548, N219, N58);
nand NAND3 (N915, N910, N98, N392);
nor NOR2 (N916, N904, N335);
nand NAND4 (N917, N913, N679, N195, N262);
xor XOR2 (N918, N914, N628);
or OR3 (N919, N897, N510, N659);
nand NAND4 (N920, N919, N133, N311, N483);
buf BUF1 (N921, N918);
buf BUF1 (N922, N876);
or OR3 (N923, N922, N837, N336);
nand NAND4 (N924, N905, N131, N117, N2);
or OR4 (N925, N924, N643, N763, N511);
xor XOR2 (N926, N925, N666);
buf BUF1 (N927, N915);
xor XOR2 (N928, N927, N488);
and AND4 (N929, N894, N142, N911, N580);
or OR4 (N930, N353, N917, N66, N792);
xor XOR2 (N931, N33, N71);
not NOT1 (N932, N931);
or OR3 (N933, N921, N750, N366);
xor XOR2 (N934, N928, N689);
buf BUF1 (N935, N932);
buf BUF1 (N936, N934);
and AND4 (N937, N929, N213, N105, N461);
buf BUF1 (N938, N926);
not NOT1 (N939, N937);
xor XOR2 (N940, N939, N90);
or OR3 (N941, N916, N109, N400);
nor NOR3 (N942, N923, N294, N919);
and AND4 (N943, N933, N408, N490, N353);
buf BUF1 (N944, N940);
nor NOR3 (N945, N943, N41, N696);
nand NAND4 (N946, N942, N474, N159, N768);
and AND3 (N947, N944, N134, N396);
nand NAND2 (N948, N938, N721);
buf BUF1 (N949, N945);
buf BUF1 (N950, N930);
nand NAND4 (N951, N948, N722, N921, N453);
buf BUF1 (N952, N950);
nor NOR2 (N953, N952, N656);
or OR3 (N954, N946, N580, N938);
nor NOR4 (N955, N947, N686, N867, N70);
xor XOR2 (N956, N941, N613);
and AND3 (N957, N912, N28, N886);
or OR4 (N958, N920, N931, N626, N704);
buf BUF1 (N959, N951);
buf BUF1 (N960, N958);
nand NAND2 (N961, N959, N599);
and AND3 (N962, N954, N581, N473);
and AND3 (N963, N953, N262, N414);
nor NOR4 (N964, N936, N43, N49, N684);
nor NOR3 (N965, N960, N392, N103);
buf BUF1 (N966, N962);
nor NOR4 (N967, N963, N299, N166, N498);
xor XOR2 (N968, N965, N799);
not NOT1 (N969, N935);
nor NOR2 (N970, N957, N531);
nor NOR2 (N971, N968, N348);
buf BUF1 (N972, N966);
or OR4 (N973, N967, N208, N631, N789);
buf BUF1 (N974, N955);
nand NAND3 (N975, N974, N951, N271);
not NOT1 (N976, N973);
nor NOR3 (N977, N972, N182, N626);
not NOT1 (N978, N976);
nand NAND4 (N979, N970, N416, N842, N288);
not NOT1 (N980, N978);
and AND2 (N981, N975, N613);
and AND2 (N982, N980, N531);
not NOT1 (N983, N981);
nor NOR2 (N984, N949, N469);
nand NAND2 (N985, N979, N721);
xor XOR2 (N986, N983, N389);
and AND4 (N987, N984, N26, N958, N492);
and AND2 (N988, N985, N354);
nor NOR2 (N989, N982, N673);
and AND3 (N990, N977, N735, N358);
not NOT1 (N991, N987);
nand NAND2 (N992, N986, N320);
buf BUF1 (N993, N988);
buf BUF1 (N994, N990);
xor XOR2 (N995, N991, N698);
or OR4 (N996, N969, N423, N866, N82);
nand NAND3 (N997, N971, N432, N257);
nand NAND3 (N998, N997, N892, N395);
not NOT1 (N999, N989);
xor XOR2 (N1000, N992, N897);
not NOT1 (N1001, N956);
not NOT1 (N1002, N995);
not NOT1 (N1003, N999);
xor XOR2 (N1004, N1003, N717);
nand NAND4 (N1005, N1002, N213, N442, N644);
or OR2 (N1006, N1000, N113);
nor NOR4 (N1007, N996, N6, N676, N779);
xor XOR2 (N1008, N994, N711);
not NOT1 (N1009, N961);
and AND3 (N1010, N964, N756, N6);
nor NOR4 (N1011, N1005, N407, N413, N226);
and AND4 (N1012, N1009, N729, N800, N196);
not NOT1 (N1013, N1010);
and AND3 (N1014, N1007, N409, N156);
xor XOR2 (N1015, N993, N988);
not NOT1 (N1016, N1001);
nand NAND2 (N1017, N1014, N1006);
xor XOR2 (N1018, N886, N46);
not NOT1 (N1019, N1011);
or OR4 (N1020, N1008, N246, N669, N812);
xor XOR2 (N1021, N1020, N25);
nand NAND3 (N1022, N1017, N794, N897);
or OR4 (N1023, N1016, N958, N950, N82);
xor XOR2 (N1024, N998, N84);
nand NAND2 (N1025, N1024, N657);
xor XOR2 (N1026, N1021, N1021);
buf BUF1 (N1027, N1023);
not NOT1 (N1028, N1025);
and AND2 (N1029, N1012, N417);
buf BUF1 (N1030, N1028);
nor NOR3 (N1031, N1018, N862, N437);
and AND3 (N1032, N1027, N881, N449);
buf BUF1 (N1033, N1004);
nand NAND2 (N1034, N1013, N930);
not NOT1 (N1035, N1030);
nand NAND4 (N1036, N1032, N545, N672, N215);
and AND2 (N1037, N1034, N138);
or OR3 (N1038, N1019, N748, N904);
nor NOR4 (N1039, N1022, N823, N486, N500);
nor NOR2 (N1040, N1015, N193);
buf BUF1 (N1041, N1040);
xor XOR2 (N1042, N1029, N929);
buf BUF1 (N1043, N1033);
nand NAND2 (N1044, N1041, N251);
buf BUF1 (N1045, N1031);
or OR2 (N1046, N1044, N934);
or OR4 (N1047, N1037, N624, N669, N928);
and AND4 (N1048, N1042, N772, N87, N197);
xor XOR2 (N1049, N1036, N386);
nand NAND2 (N1050, N1038, N543);
nor NOR2 (N1051, N1048, N43);
buf BUF1 (N1052, N1049);
xor XOR2 (N1053, N1047, N639);
xor XOR2 (N1054, N1026, N719);
xor XOR2 (N1055, N1043, N728);
and AND4 (N1056, N1053, N523, N225, N67);
not NOT1 (N1057, N1051);
and AND4 (N1058, N1057, N583, N96, N174);
nand NAND2 (N1059, N1052, N873);
nor NOR2 (N1060, N1054, N477);
xor XOR2 (N1061, N1055, N335);
nand NAND2 (N1062, N1035, N536);
or OR3 (N1063, N1060, N100, N909);
buf BUF1 (N1064, N1046);
nor NOR2 (N1065, N1062, N845);
nand NAND2 (N1066, N1061, N206);
buf BUF1 (N1067, N1039);
and AND3 (N1068, N1066, N806, N865);
and AND4 (N1069, N1059, N39, N425, N361);
not NOT1 (N1070, N1045);
nor NOR2 (N1071, N1070, N411);
nand NAND2 (N1072, N1064, N788);
xor XOR2 (N1073, N1072, N542);
not NOT1 (N1074, N1050);
nor NOR2 (N1075, N1058, N586);
or OR2 (N1076, N1071, N551);
xor XOR2 (N1077, N1056, N595);
not NOT1 (N1078, N1065);
or OR4 (N1079, N1069, N504, N444, N553);
nor NOR2 (N1080, N1063, N1055);
nand NAND3 (N1081, N1068, N678, N97);
buf BUF1 (N1082, N1079);
nand NAND2 (N1083, N1077, N869);
and AND3 (N1084, N1076, N1066, N794);
nor NOR2 (N1085, N1080, N868);
nor NOR2 (N1086, N1085, N757);
nand NAND4 (N1087, N1078, N1004, N7, N1076);
buf BUF1 (N1088, N1073);
nor NOR2 (N1089, N1081, N370);
or OR4 (N1090, N1084, N87, N767, N1052);
nor NOR2 (N1091, N1089, N30);
nand NAND4 (N1092, N1067, N296, N51, N885);
not NOT1 (N1093, N1082);
or OR4 (N1094, N1087, N723, N187, N1065);
buf BUF1 (N1095, N1075);
nor NOR2 (N1096, N1086, N910);
and AND4 (N1097, N1074, N880, N248, N355);
nor NOR3 (N1098, N1094, N870, N351);
buf BUF1 (N1099, N1083);
xor XOR2 (N1100, N1090, N631);
buf BUF1 (N1101, N1096);
or OR2 (N1102, N1092, N726);
xor XOR2 (N1103, N1088, N577);
or OR3 (N1104, N1101, N242, N1007);
nor NOR3 (N1105, N1095, N537, N713);
xor XOR2 (N1106, N1105, N993);
nor NOR4 (N1107, N1103, N252, N854, N1101);
nand NAND3 (N1108, N1102, N164, N467);
or OR3 (N1109, N1097, N785, N1060);
buf BUF1 (N1110, N1091);
or OR3 (N1111, N1110, N44, N516);
nor NOR3 (N1112, N1100, N779, N897);
xor XOR2 (N1113, N1104, N188);
xor XOR2 (N1114, N1113, N963);
nor NOR3 (N1115, N1112, N683, N792);
nand NAND4 (N1116, N1093, N780, N387, N126);
nor NOR3 (N1117, N1098, N15, N779);
nand NAND4 (N1118, N1107, N341, N137, N705);
nand NAND3 (N1119, N1115, N603, N966);
not NOT1 (N1120, N1106);
xor XOR2 (N1121, N1109, N970);
nor NOR4 (N1122, N1116, N936, N818, N550);
nor NOR2 (N1123, N1108, N592);
and AND4 (N1124, N1099, N525, N607, N837);
buf BUF1 (N1125, N1121);
buf BUF1 (N1126, N1114);
or OR4 (N1127, N1122, N380, N774, N786);
nand NAND3 (N1128, N1111, N488, N1054);
xor XOR2 (N1129, N1120, N888);
buf BUF1 (N1130, N1126);
or OR3 (N1131, N1118, N863, N1037);
buf BUF1 (N1132, N1124);
xor XOR2 (N1133, N1127, N283);
and AND3 (N1134, N1130, N1015, N226);
nand NAND4 (N1135, N1119, N776, N729, N966);
or OR2 (N1136, N1131, N482);
nand NAND2 (N1137, N1125, N799);
and AND2 (N1138, N1133, N930);
nand NAND2 (N1139, N1138, N332);
xor XOR2 (N1140, N1117, N597);
or OR3 (N1141, N1129, N522, N361);
nand NAND4 (N1142, N1132, N82, N284, N180);
or OR3 (N1143, N1142, N860, N309);
or OR3 (N1144, N1123, N559, N32);
xor XOR2 (N1145, N1140, N881);
nor NOR2 (N1146, N1135, N653);
xor XOR2 (N1147, N1139, N261);
or OR4 (N1148, N1143, N913, N366, N61);
nor NOR3 (N1149, N1146, N313, N286);
buf BUF1 (N1150, N1144);
buf BUF1 (N1151, N1134);
nand NAND3 (N1152, N1148, N873, N368);
and AND4 (N1153, N1145, N780, N1116, N634);
buf BUF1 (N1154, N1147);
nor NOR4 (N1155, N1128, N152, N838, N231);
nor NOR3 (N1156, N1152, N232, N704);
or OR3 (N1157, N1151, N174, N139);
and AND3 (N1158, N1154, N478, N534);
nor NOR4 (N1159, N1156, N395, N290, N511);
nand NAND4 (N1160, N1136, N782, N679, N869);
nor NOR2 (N1161, N1137, N902);
not NOT1 (N1162, N1155);
xor XOR2 (N1163, N1158, N623);
nor NOR3 (N1164, N1141, N16, N141);
buf BUF1 (N1165, N1149);
buf BUF1 (N1166, N1160);
nand NAND4 (N1167, N1162, N532, N706, N739);
not NOT1 (N1168, N1161);
and AND4 (N1169, N1153, N882, N360, N201);
nand NAND2 (N1170, N1157, N479);
nor NOR2 (N1171, N1166, N368);
not NOT1 (N1172, N1164);
not NOT1 (N1173, N1150);
nand NAND3 (N1174, N1171, N45, N139);
and AND3 (N1175, N1173, N561, N1037);
not NOT1 (N1176, N1167);
buf BUF1 (N1177, N1169);
nand NAND4 (N1178, N1165, N39, N531, N490);
xor XOR2 (N1179, N1177, N938);
xor XOR2 (N1180, N1178, N714);
and AND2 (N1181, N1159, N942);
or OR4 (N1182, N1174, N850, N762, N468);
nand NAND2 (N1183, N1182, N757);
and AND4 (N1184, N1176, N242, N37, N916);
or OR4 (N1185, N1175, N666, N680, N330);
not NOT1 (N1186, N1179);
xor XOR2 (N1187, N1170, N949);
not NOT1 (N1188, N1163);
or OR3 (N1189, N1187, N359, N425);
buf BUF1 (N1190, N1181);
not NOT1 (N1191, N1190);
and AND3 (N1192, N1183, N765, N1039);
and AND2 (N1193, N1189, N254);
not NOT1 (N1194, N1191);
and AND3 (N1195, N1194, N1009, N1008);
or OR4 (N1196, N1193, N802, N892, N1143);
or OR4 (N1197, N1185, N733, N211, N523);
nand NAND2 (N1198, N1197, N646);
nor NOR2 (N1199, N1188, N791);
not NOT1 (N1200, N1195);
nand NAND2 (N1201, N1180, N100);
not NOT1 (N1202, N1186);
xor XOR2 (N1203, N1198, N270);
not NOT1 (N1204, N1202);
xor XOR2 (N1205, N1192, N1033);
and AND3 (N1206, N1201, N874, N642);
and AND2 (N1207, N1168, N892);
and AND2 (N1208, N1199, N92);
nand NAND3 (N1209, N1172, N475, N872);
buf BUF1 (N1210, N1196);
xor XOR2 (N1211, N1184, N988);
nand NAND4 (N1212, N1206, N723, N333, N231);
or OR2 (N1213, N1200, N222);
and AND4 (N1214, N1211, N24, N903, N779);
xor XOR2 (N1215, N1209, N173);
not NOT1 (N1216, N1212);
xor XOR2 (N1217, N1210, N810);
nand NAND4 (N1218, N1214, N468, N194, N583);
nand NAND4 (N1219, N1216, N439, N1042, N11);
not NOT1 (N1220, N1203);
xor XOR2 (N1221, N1218, N262);
nor NOR4 (N1222, N1204, N532, N633, N457);
nand NAND4 (N1223, N1217, N1165, N642, N802);
buf BUF1 (N1224, N1220);
buf BUF1 (N1225, N1213);
buf BUF1 (N1226, N1207);
xor XOR2 (N1227, N1222, N684);
nor NOR2 (N1228, N1215, N467);
and AND2 (N1229, N1228, N788);
not NOT1 (N1230, N1221);
buf BUF1 (N1231, N1223);
xor XOR2 (N1232, N1208, N1006);
not NOT1 (N1233, N1226);
and AND4 (N1234, N1219, N966, N355, N531);
nor NOR3 (N1235, N1224, N202, N1229);
buf BUF1 (N1236, N114);
not NOT1 (N1237, N1231);
not NOT1 (N1238, N1232);
not NOT1 (N1239, N1205);
not NOT1 (N1240, N1225);
or OR2 (N1241, N1238, N74);
not NOT1 (N1242, N1240);
or OR4 (N1243, N1233, N1022, N657, N447);
buf BUF1 (N1244, N1239);
or OR3 (N1245, N1234, N515, N1213);
not NOT1 (N1246, N1243);
nand NAND2 (N1247, N1245, N195);
buf BUF1 (N1248, N1227);
nor NOR4 (N1249, N1247, N981, N613, N1085);
nand NAND4 (N1250, N1236, N1115, N1014, N284);
or OR4 (N1251, N1242, N570, N249, N299);
nor NOR2 (N1252, N1230, N1006);
and AND2 (N1253, N1241, N1160);
buf BUF1 (N1254, N1235);
not NOT1 (N1255, N1237);
nor NOR2 (N1256, N1254, N572);
xor XOR2 (N1257, N1250, N196);
xor XOR2 (N1258, N1255, N707);
buf BUF1 (N1259, N1251);
and AND3 (N1260, N1256, N151, N397);
nor NOR4 (N1261, N1246, N135, N994, N477);
and AND3 (N1262, N1248, N294, N464);
not NOT1 (N1263, N1261);
xor XOR2 (N1264, N1249, N936);
or OR3 (N1265, N1259, N217, N487);
or OR3 (N1266, N1263, N652, N533);
xor XOR2 (N1267, N1264, N155);
buf BUF1 (N1268, N1258);
nor NOR4 (N1269, N1260, N354, N230, N960);
xor XOR2 (N1270, N1265, N1249);
xor XOR2 (N1271, N1268, N185);
not NOT1 (N1272, N1253);
and AND2 (N1273, N1267, N324);
and AND3 (N1274, N1252, N255, N950);
and AND4 (N1275, N1262, N822, N128, N441);
nor NOR2 (N1276, N1272, N381);
buf BUF1 (N1277, N1274);
and AND3 (N1278, N1276, N135, N527);
nor NOR2 (N1279, N1277, N480);
nand NAND4 (N1280, N1244, N1092, N416, N740);
or OR3 (N1281, N1278, N929, N977);
xor XOR2 (N1282, N1275, N906);
and AND2 (N1283, N1270, N180);
or OR3 (N1284, N1269, N1225, N657);
and AND2 (N1285, N1273, N896);
not NOT1 (N1286, N1280);
xor XOR2 (N1287, N1279, N2);
buf BUF1 (N1288, N1266);
and AND3 (N1289, N1288, N233, N651);
xor XOR2 (N1290, N1286, N744);
buf BUF1 (N1291, N1271);
and AND4 (N1292, N1285, N966, N1037, N507);
and AND3 (N1293, N1282, N261, N257);
not NOT1 (N1294, N1281);
xor XOR2 (N1295, N1292, N344);
xor XOR2 (N1296, N1283, N85);
buf BUF1 (N1297, N1289);
nor NOR4 (N1298, N1296, N1119, N74, N182);
not NOT1 (N1299, N1290);
and AND3 (N1300, N1287, N353, N813);
not NOT1 (N1301, N1297);
or OR3 (N1302, N1294, N515, N100);
or OR4 (N1303, N1293, N942, N96, N431);
buf BUF1 (N1304, N1284);
not NOT1 (N1305, N1302);
xor XOR2 (N1306, N1295, N144);
buf BUF1 (N1307, N1298);
or OR4 (N1308, N1307, N934, N148, N100);
xor XOR2 (N1309, N1304, N913);
buf BUF1 (N1310, N1309);
and AND4 (N1311, N1299, N555, N1275, N304);
xor XOR2 (N1312, N1300, N1052);
and AND3 (N1313, N1305, N989, N74);
nand NAND3 (N1314, N1257, N1202, N277);
nand NAND3 (N1315, N1308, N1266, N837);
buf BUF1 (N1316, N1310);
buf BUF1 (N1317, N1316);
and AND2 (N1318, N1311, N916);
and AND4 (N1319, N1314, N1155, N221, N27);
nand NAND2 (N1320, N1306, N1144);
nor NOR2 (N1321, N1315, N170);
nor NOR2 (N1322, N1312, N572);
not NOT1 (N1323, N1317);
buf BUF1 (N1324, N1320);
buf BUF1 (N1325, N1319);
buf BUF1 (N1326, N1291);
nor NOR2 (N1327, N1324, N163);
nand NAND3 (N1328, N1325, N1085, N192);
and AND3 (N1329, N1318, N81, N262);
nor NOR2 (N1330, N1328, N253);
and AND4 (N1331, N1322, N1270, N782, N467);
nor NOR4 (N1332, N1327, N581, N264, N473);
buf BUF1 (N1333, N1326);
nand NAND3 (N1334, N1321, N430, N122);
buf BUF1 (N1335, N1330);
xor XOR2 (N1336, N1313, N433);
or OR3 (N1337, N1303, N783, N24);
or OR4 (N1338, N1332, N353, N534, N844);
and AND2 (N1339, N1301, N251);
and AND4 (N1340, N1339, N489, N389, N711);
xor XOR2 (N1341, N1333, N293);
xor XOR2 (N1342, N1335, N40);
nor NOR3 (N1343, N1331, N54, N52);
nand NAND3 (N1344, N1329, N953, N542);
buf BUF1 (N1345, N1337);
or OR4 (N1346, N1343, N695, N90, N484);
or OR3 (N1347, N1342, N1210, N649);
buf BUF1 (N1348, N1334);
and AND2 (N1349, N1336, N1084);
xor XOR2 (N1350, N1346, N1316);
and AND2 (N1351, N1323, N1074);
not NOT1 (N1352, N1341);
and AND3 (N1353, N1338, N265, N1103);
nand NAND4 (N1354, N1350, N743, N1284, N685);
and AND2 (N1355, N1348, N1234);
and AND2 (N1356, N1352, N25);
nand NAND4 (N1357, N1356, N183, N367, N865);
buf BUF1 (N1358, N1351);
xor XOR2 (N1359, N1344, N1018);
nor NOR2 (N1360, N1353, N208);
buf BUF1 (N1361, N1355);
buf BUF1 (N1362, N1347);
and AND3 (N1363, N1360, N1050, N575);
or OR2 (N1364, N1358, N73);
nor NOR3 (N1365, N1361, N873, N546);
nor NOR2 (N1366, N1340, N1058);
nor NOR4 (N1367, N1365, N682, N1185, N281);
or OR3 (N1368, N1345, N74, N1298);
nand NAND3 (N1369, N1354, N582, N135);
and AND3 (N1370, N1369, N720, N81);
nor NOR2 (N1371, N1349, N930);
and AND4 (N1372, N1371, N230, N860, N1150);
or OR3 (N1373, N1363, N1, N120);
or OR2 (N1374, N1368, N209);
nor NOR3 (N1375, N1372, N491, N1229);
and AND4 (N1376, N1366, N1219, N598, N1251);
xor XOR2 (N1377, N1357, N1249);
xor XOR2 (N1378, N1367, N285);
and AND3 (N1379, N1377, N645, N546);
xor XOR2 (N1380, N1370, N1213);
nor NOR2 (N1381, N1376, N1274);
not NOT1 (N1382, N1378);
and AND3 (N1383, N1375, N707, N895);
nor NOR3 (N1384, N1359, N811, N59);
and AND4 (N1385, N1373, N1203, N851, N1022);
not NOT1 (N1386, N1385);
nand NAND2 (N1387, N1379, N613);
or OR3 (N1388, N1386, N109, N196);
nor NOR3 (N1389, N1388, N844, N646);
nor NOR3 (N1390, N1382, N626, N912);
and AND4 (N1391, N1364, N39, N492, N973);
not NOT1 (N1392, N1387);
xor XOR2 (N1393, N1392, N1088);
xor XOR2 (N1394, N1374, N1193);
nor NOR4 (N1395, N1380, N981, N1126, N232);
and AND2 (N1396, N1394, N795);
nand NAND3 (N1397, N1381, N730, N563);
buf BUF1 (N1398, N1391);
and AND2 (N1399, N1390, N1344);
and AND4 (N1400, N1393, N175, N1263, N1102);
and AND3 (N1401, N1399, N288, N69);
not NOT1 (N1402, N1401);
buf BUF1 (N1403, N1383);
xor XOR2 (N1404, N1397, N19);
not NOT1 (N1405, N1400);
not NOT1 (N1406, N1362);
or OR3 (N1407, N1389, N614, N1144);
nor NOR3 (N1408, N1406, N43, N490);
not NOT1 (N1409, N1396);
xor XOR2 (N1410, N1398, N251);
or OR2 (N1411, N1407, N408);
not NOT1 (N1412, N1409);
and AND4 (N1413, N1384, N922, N140, N237);
or OR4 (N1414, N1402, N920, N461, N228);
and AND4 (N1415, N1395, N78, N1087, N58);
buf BUF1 (N1416, N1413);
not NOT1 (N1417, N1415);
not NOT1 (N1418, N1404);
buf BUF1 (N1419, N1403);
not NOT1 (N1420, N1418);
nor NOR3 (N1421, N1412, N552, N252);
or OR3 (N1422, N1416, N621, N883);
and AND4 (N1423, N1414, N489, N1236, N51);
not NOT1 (N1424, N1417);
xor XOR2 (N1425, N1422, N567);
xor XOR2 (N1426, N1410, N1422);
not NOT1 (N1427, N1424);
not NOT1 (N1428, N1427);
xor XOR2 (N1429, N1425, N663);
nand NAND2 (N1430, N1420, N386);
not NOT1 (N1431, N1408);
nand NAND3 (N1432, N1431, N890, N685);
and AND4 (N1433, N1432, N59, N47, N1121);
nand NAND2 (N1434, N1423, N948);
or OR3 (N1435, N1428, N1397, N323);
nand NAND2 (N1436, N1429, N929);
not NOT1 (N1437, N1426);
xor XOR2 (N1438, N1411, N933);
nand NAND3 (N1439, N1437, N116, N793);
and AND2 (N1440, N1434, N722);
xor XOR2 (N1441, N1439, N93);
xor XOR2 (N1442, N1421, N1134);
nand NAND4 (N1443, N1433, N1342, N1317, N1216);
buf BUF1 (N1444, N1435);
nand NAND4 (N1445, N1438, N362, N46, N1432);
buf BUF1 (N1446, N1405);
and AND4 (N1447, N1443, N978, N248, N841);
and AND3 (N1448, N1445, N319, N1291);
xor XOR2 (N1449, N1441, N1126);
nor NOR4 (N1450, N1442, N443, N1404, N244);
buf BUF1 (N1451, N1430);
and AND2 (N1452, N1419, N811);
or OR3 (N1453, N1450, N606, N756);
or OR4 (N1454, N1440, N230, N604, N993);
not NOT1 (N1455, N1452);
buf BUF1 (N1456, N1453);
nor NOR2 (N1457, N1444, N481);
xor XOR2 (N1458, N1436, N561);
xor XOR2 (N1459, N1449, N547);
nor NOR3 (N1460, N1451, N674, N802);
or OR3 (N1461, N1456, N1370, N1301);
not NOT1 (N1462, N1461);
nor NOR2 (N1463, N1458, N248);
nand NAND2 (N1464, N1448, N277);
xor XOR2 (N1465, N1457, N127);
or OR3 (N1466, N1454, N69, N181);
or OR3 (N1467, N1455, N1386, N296);
buf BUF1 (N1468, N1446);
buf BUF1 (N1469, N1460);
not NOT1 (N1470, N1466);
nand NAND4 (N1471, N1467, N869, N813, N910);
nor NOR3 (N1472, N1469, N1365, N672);
nand NAND3 (N1473, N1462, N205, N221);
not NOT1 (N1474, N1473);
buf BUF1 (N1475, N1465);
not NOT1 (N1476, N1474);
xor XOR2 (N1477, N1464, N17);
and AND4 (N1478, N1459, N1312, N21, N880);
xor XOR2 (N1479, N1478, N1434);
nor NOR2 (N1480, N1476, N1054);
nor NOR2 (N1481, N1463, N928);
nor NOR3 (N1482, N1475, N992, N1416);
nand NAND3 (N1483, N1471, N862, N1386);
nand NAND2 (N1484, N1470, N495);
or OR2 (N1485, N1479, N364);
not NOT1 (N1486, N1447);
nand NAND4 (N1487, N1481, N241, N949, N1002);
nand NAND3 (N1488, N1483, N1320, N1031);
not NOT1 (N1489, N1480);
nand NAND2 (N1490, N1468, N550);
not NOT1 (N1491, N1472);
xor XOR2 (N1492, N1491, N871);
buf BUF1 (N1493, N1492);
or OR2 (N1494, N1486, N563);
or OR2 (N1495, N1485, N430);
not NOT1 (N1496, N1490);
nand NAND2 (N1497, N1496, N1198);
xor XOR2 (N1498, N1487, N697);
not NOT1 (N1499, N1489);
not NOT1 (N1500, N1477);
buf BUF1 (N1501, N1500);
or OR4 (N1502, N1501, N53, N1115, N1229);
not NOT1 (N1503, N1498);
and AND4 (N1504, N1488, N573, N502, N7);
buf BUF1 (N1505, N1493);
and AND4 (N1506, N1494, N495, N799, N21);
xor XOR2 (N1507, N1497, N1084);
nor NOR4 (N1508, N1499, N824, N1348, N183);
nor NOR3 (N1509, N1502, N1113, N816);
nor NOR3 (N1510, N1495, N792, N76);
or OR2 (N1511, N1503, N617);
xor XOR2 (N1512, N1509, N29);
and AND3 (N1513, N1508, N497, N786);
or OR2 (N1514, N1510, N363);
nand NAND4 (N1515, N1512, N1199, N870, N1247);
or OR3 (N1516, N1515, N97, N528);
buf BUF1 (N1517, N1516);
not NOT1 (N1518, N1511);
or OR3 (N1519, N1484, N563, N1430);
nand NAND4 (N1520, N1514, N576, N1514, N1399);
nand NAND4 (N1521, N1505, N1009, N572, N599);
nor NOR4 (N1522, N1521, N600, N1392, N1389);
not NOT1 (N1523, N1513);
nor NOR3 (N1524, N1482, N751, N207);
buf BUF1 (N1525, N1524);
xor XOR2 (N1526, N1522, N1369);
and AND4 (N1527, N1519, N679, N66, N609);
buf BUF1 (N1528, N1527);
buf BUF1 (N1529, N1520);
nand NAND4 (N1530, N1504, N268, N542, N86);
nand NAND2 (N1531, N1528, N478);
buf BUF1 (N1532, N1507);
and AND2 (N1533, N1529, N1025);
nor NOR3 (N1534, N1532, N1038, N420);
nand NAND2 (N1535, N1506, N457);
or OR3 (N1536, N1535, N258, N1238);
xor XOR2 (N1537, N1531, N1529);
or OR2 (N1538, N1536, N940);
nor NOR3 (N1539, N1530, N1525, N385);
xor XOR2 (N1540, N1185, N781);
buf BUF1 (N1541, N1538);
or OR4 (N1542, N1533, N1011, N1243, N733);
buf BUF1 (N1543, N1541);
and AND2 (N1544, N1543, N206);
nand NAND3 (N1545, N1526, N638, N187);
nor NOR4 (N1546, N1539, N1223, N328, N290);
not NOT1 (N1547, N1537);
or OR4 (N1548, N1517, N1293, N1508, N585);
nand NAND2 (N1549, N1548, N1484);
buf BUF1 (N1550, N1549);
buf BUF1 (N1551, N1545);
nor NOR2 (N1552, N1523, N1143);
nand NAND4 (N1553, N1550, N1502, N1281, N1190);
nor NOR3 (N1554, N1542, N1340, N461);
and AND3 (N1555, N1546, N879, N1262);
nor NOR3 (N1556, N1554, N475, N570);
not NOT1 (N1557, N1540);
nand NAND4 (N1558, N1556, N855, N1429, N1414);
or OR3 (N1559, N1558, N90, N1273);
nand NAND4 (N1560, N1534, N1323, N1302, N1041);
or OR4 (N1561, N1551, N807, N207, N667);
not NOT1 (N1562, N1552);
nor NOR4 (N1563, N1561, N366, N853, N1477);
nor NOR4 (N1564, N1557, N60, N252, N598);
buf BUF1 (N1565, N1560);
not NOT1 (N1566, N1547);
nor NOR4 (N1567, N1553, N1341, N1513, N1237);
not NOT1 (N1568, N1518);
nand NAND3 (N1569, N1566, N159, N301);
not NOT1 (N1570, N1567);
xor XOR2 (N1571, N1565, N76);
or OR2 (N1572, N1544, N100);
buf BUF1 (N1573, N1568);
xor XOR2 (N1574, N1563, N892);
nor NOR2 (N1575, N1562, N700);
nand NAND4 (N1576, N1572, N660, N1407, N1203);
and AND2 (N1577, N1574, N397);
nor NOR4 (N1578, N1564, N1182, N1520, N1134);
nor NOR3 (N1579, N1576, N53, N118);
or OR4 (N1580, N1555, N962, N199, N627);
nor NOR2 (N1581, N1580, N149);
xor XOR2 (N1582, N1575, N639);
or OR4 (N1583, N1570, N1573, N560, N308);
and AND4 (N1584, N1065, N1132, N1183, N754);
and AND4 (N1585, N1582, N367, N406, N1204);
nand NAND4 (N1586, N1578, N283, N1355, N866);
xor XOR2 (N1587, N1584, N122);
xor XOR2 (N1588, N1569, N585);
or OR3 (N1589, N1588, N634, N870);
not NOT1 (N1590, N1587);
or OR4 (N1591, N1577, N309, N1552, N746);
not NOT1 (N1592, N1579);
and AND4 (N1593, N1592, N851, N1525, N422);
not NOT1 (N1594, N1571);
and AND2 (N1595, N1590, N1335);
and AND3 (N1596, N1559, N313, N104);
and AND2 (N1597, N1589, N329);
or OR2 (N1598, N1585, N369);
nand NAND4 (N1599, N1598, N1063, N776, N888);
xor XOR2 (N1600, N1594, N689);
not NOT1 (N1601, N1596);
xor XOR2 (N1602, N1599, N1080);
nand NAND2 (N1603, N1601, N914);
nand NAND3 (N1604, N1583, N848, N595);
and AND2 (N1605, N1600, N545);
buf BUF1 (N1606, N1595);
xor XOR2 (N1607, N1597, N926);
not NOT1 (N1608, N1586);
and AND2 (N1609, N1607, N791);
and AND3 (N1610, N1605, N598, N972);
and AND3 (N1611, N1610, N947, N914);
xor XOR2 (N1612, N1609, N1404);
and AND2 (N1613, N1603, N1011);
and AND4 (N1614, N1593, N131, N1104, N470);
nand NAND4 (N1615, N1604, N602, N1103, N405);
or OR2 (N1616, N1608, N1162);
or OR4 (N1617, N1612, N996, N720, N136);
and AND4 (N1618, N1606, N602, N64, N1389);
buf BUF1 (N1619, N1602);
xor XOR2 (N1620, N1614, N684);
or OR4 (N1621, N1617, N1609, N254, N650);
nor NOR2 (N1622, N1591, N1181);
buf BUF1 (N1623, N1616);
buf BUF1 (N1624, N1623);
not NOT1 (N1625, N1618);
xor XOR2 (N1626, N1620, N599);
and AND2 (N1627, N1621, N1071);
not NOT1 (N1628, N1627);
buf BUF1 (N1629, N1581);
or OR4 (N1630, N1611, N1526, N28, N349);
buf BUF1 (N1631, N1629);
nor NOR3 (N1632, N1626, N328, N866);
not NOT1 (N1633, N1624);
nand NAND2 (N1634, N1631, N1037);
nor NOR3 (N1635, N1628, N1438, N126);
or OR2 (N1636, N1632, N591);
xor XOR2 (N1637, N1634, N1353);
or OR2 (N1638, N1625, N1041);
not NOT1 (N1639, N1633);
nand NAND4 (N1640, N1622, N743, N52, N739);
and AND4 (N1641, N1637, N472, N1541, N427);
nand NAND4 (N1642, N1630, N474, N524, N235);
buf BUF1 (N1643, N1641);
xor XOR2 (N1644, N1639, N1413);
and AND4 (N1645, N1613, N1427, N416, N1504);
buf BUF1 (N1646, N1643);
xor XOR2 (N1647, N1645, N855);
buf BUF1 (N1648, N1647);
nor NOR3 (N1649, N1615, N708, N1505);
or OR4 (N1650, N1640, N781, N1433, N501);
nor NOR4 (N1651, N1619, N471, N1456, N1504);
and AND4 (N1652, N1651, N688, N499, N1499);
or OR3 (N1653, N1642, N1383, N722);
nor NOR3 (N1654, N1650, N542, N551);
and AND2 (N1655, N1646, N590);
xor XOR2 (N1656, N1644, N324);
nor NOR4 (N1657, N1653, N1119, N1573, N992);
nand NAND2 (N1658, N1636, N1112);
and AND4 (N1659, N1635, N447, N1186, N651);
nand NAND3 (N1660, N1654, N208, N285);
buf BUF1 (N1661, N1649);
nand NAND4 (N1662, N1659, N476, N538, N486);
and AND4 (N1663, N1662, N360, N1477, N485);
nor NOR3 (N1664, N1648, N206, N59);
buf BUF1 (N1665, N1656);
buf BUF1 (N1666, N1652);
xor XOR2 (N1667, N1661, N639);
or OR3 (N1668, N1666, N294, N737);
and AND3 (N1669, N1657, N1190, N240);
nor NOR2 (N1670, N1669, N253);
or OR3 (N1671, N1664, N1661, N646);
xor XOR2 (N1672, N1668, N1149);
nor NOR2 (N1673, N1671, N412);
nand NAND4 (N1674, N1672, N106, N1141, N893);
nand NAND2 (N1675, N1674, N1058);
or OR4 (N1676, N1660, N1607, N1523, N501);
buf BUF1 (N1677, N1675);
not NOT1 (N1678, N1676);
and AND2 (N1679, N1638, N1241);
xor XOR2 (N1680, N1665, N546);
nand NAND3 (N1681, N1658, N302, N800);
nor NOR3 (N1682, N1678, N351, N877);
nor NOR2 (N1683, N1681, N546);
not NOT1 (N1684, N1667);
not NOT1 (N1685, N1673);
buf BUF1 (N1686, N1655);
xor XOR2 (N1687, N1679, N154);
not NOT1 (N1688, N1680);
or OR3 (N1689, N1686, N536, N235);
nor NOR2 (N1690, N1684, N1586);
not NOT1 (N1691, N1689);
and AND2 (N1692, N1685, N1189);
or OR4 (N1693, N1663, N546, N119, N994);
nand NAND4 (N1694, N1683, N502, N757, N1570);
or OR4 (N1695, N1670, N248, N657, N78);
nor NOR2 (N1696, N1695, N328);
nand NAND3 (N1697, N1696, N135, N713);
xor XOR2 (N1698, N1677, N1003);
xor XOR2 (N1699, N1694, N1486);
or OR2 (N1700, N1699, N221);
buf BUF1 (N1701, N1693);
buf BUF1 (N1702, N1692);
xor XOR2 (N1703, N1697, N220);
nor NOR3 (N1704, N1701, N1207, N606);
and AND4 (N1705, N1688, N1647, N730, N766);
or OR4 (N1706, N1705, N56, N430, N908);
buf BUF1 (N1707, N1687);
nand NAND3 (N1708, N1682, N1611, N537);
xor XOR2 (N1709, N1700, N1551);
and AND3 (N1710, N1708, N1301, N1495);
buf BUF1 (N1711, N1706);
not NOT1 (N1712, N1702);
or OR4 (N1713, N1712, N1361, N1527, N939);
and AND2 (N1714, N1698, N1077);
nand NAND2 (N1715, N1711, N1697);
not NOT1 (N1716, N1715);
xor XOR2 (N1717, N1716, N801);
nand NAND4 (N1718, N1704, N235, N757, N648);
and AND2 (N1719, N1703, N669);
and AND4 (N1720, N1709, N524, N164, N375);
and AND4 (N1721, N1717, N481, N1084, N372);
nor NOR4 (N1722, N1691, N370, N846, N519);
nand NAND2 (N1723, N1690, N172);
nor NOR2 (N1724, N1718, N1021);
not NOT1 (N1725, N1714);
and AND4 (N1726, N1724, N1525, N514, N954);
or OR3 (N1727, N1707, N156, N987);
xor XOR2 (N1728, N1721, N396);
and AND3 (N1729, N1722, N1220, N1434);
or OR3 (N1730, N1719, N1223, N1028);
or OR4 (N1731, N1720, N718, N343, N1060);
buf BUF1 (N1732, N1710);
not NOT1 (N1733, N1725);
nor NOR3 (N1734, N1727, N809, N314);
not NOT1 (N1735, N1734);
and AND3 (N1736, N1732, N1643, N729);
xor XOR2 (N1737, N1731, N271);
buf BUF1 (N1738, N1736);
or OR2 (N1739, N1713, N894);
nor NOR2 (N1740, N1728, N1034);
not NOT1 (N1741, N1733);
xor XOR2 (N1742, N1730, N814);
buf BUF1 (N1743, N1737);
nand NAND4 (N1744, N1742, N1308, N1164, N1584);
and AND4 (N1745, N1738, N896, N1063, N1332);
and AND3 (N1746, N1729, N1, N47);
or OR3 (N1747, N1743, N938, N1299);
xor XOR2 (N1748, N1746, N1673);
nor NOR3 (N1749, N1747, N1157, N1082);
and AND4 (N1750, N1735, N1037, N202, N1075);
buf BUF1 (N1751, N1750);
xor XOR2 (N1752, N1741, N1472);
nand NAND2 (N1753, N1748, N576);
and AND3 (N1754, N1740, N166, N1611);
or OR2 (N1755, N1754, N465);
nand NAND4 (N1756, N1744, N544, N1457, N559);
nor NOR2 (N1757, N1755, N38);
buf BUF1 (N1758, N1745);
buf BUF1 (N1759, N1753);
nor NOR4 (N1760, N1759, N1442, N878, N936);
or OR2 (N1761, N1726, N748);
nand NAND2 (N1762, N1739, N1706);
or OR3 (N1763, N1761, N1617, N836);
buf BUF1 (N1764, N1758);
or OR3 (N1765, N1760, N1376, N37);
buf BUF1 (N1766, N1757);
xor XOR2 (N1767, N1756, N1064);
xor XOR2 (N1768, N1752, N281);
or OR4 (N1769, N1751, N1315, N855, N1504);
not NOT1 (N1770, N1765);
and AND4 (N1771, N1763, N1166, N1612, N1534);
and AND2 (N1772, N1771, N58);
or OR3 (N1773, N1749, N128, N1541);
not NOT1 (N1774, N1768);
nor NOR2 (N1775, N1767, N1268);
nor NOR4 (N1776, N1769, N545, N1680, N1078);
or OR2 (N1777, N1773, N384);
not NOT1 (N1778, N1766);
and AND3 (N1779, N1723, N584, N723);
xor XOR2 (N1780, N1778, N1188);
xor XOR2 (N1781, N1770, N1039);
buf BUF1 (N1782, N1762);
nor NOR2 (N1783, N1777, N305);
and AND4 (N1784, N1783, N1296, N847, N483);
buf BUF1 (N1785, N1775);
xor XOR2 (N1786, N1776, N55);
nor NOR2 (N1787, N1781, N1568);
not NOT1 (N1788, N1764);
nor NOR2 (N1789, N1779, N815);
xor XOR2 (N1790, N1789, N106);
or OR4 (N1791, N1787, N655, N719, N191);
or OR2 (N1792, N1772, N619);
nor NOR3 (N1793, N1774, N1400, N1176);
not NOT1 (N1794, N1792);
or OR4 (N1795, N1780, N754, N1417, N1217);
buf BUF1 (N1796, N1782);
nand NAND2 (N1797, N1795, N147);
or OR3 (N1798, N1791, N316, N724);
or OR4 (N1799, N1796, N877, N365, N201);
nand NAND3 (N1800, N1797, N1428, N945);
or OR4 (N1801, N1785, N550, N854, N1576);
and AND2 (N1802, N1788, N381);
nor NOR3 (N1803, N1798, N673, N76);
not NOT1 (N1804, N1790);
xor XOR2 (N1805, N1802, N1755);
nor NOR4 (N1806, N1801, N593, N1329, N714);
xor XOR2 (N1807, N1786, N1780);
buf BUF1 (N1808, N1800);
nand NAND3 (N1809, N1793, N1495, N1779);
and AND3 (N1810, N1799, N19, N1145);
or OR4 (N1811, N1803, N1516, N1393, N1467);
nand NAND4 (N1812, N1807, N1081, N1294, N1691);
and AND2 (N1813, N1794, N411);
nor NOR4 (N1814, N1813, N506, N857, N564);
or OR2 (N1815, N1806, N210);
or OR3 (N1816, N1814, N1361, N188);
or OR3 (N1817, N1784, N743, N1260);
or OR3 (N1818, N1815, N1797, N214);
not NOT1 (N1819, N1817);
or OR2 (N1820, N1811, N17);
and AND2 (N1821, N1809, N418);
nand NAND4 (N1822, N1812, N575, N170, N410);
xor XOR2 (N1823, N1810, N530);
nor NOR3 (N1824, N1818, N1643, N1056);
buf BUF1 (N1825, N1816);
buf BUF1 (N1826, N1819);
nor NOR2 (N1827, N1805, N909);
nor NOR2 (N1828, N1808, N912);
and AND4 (N1829, N1826, N1151, N1681, N948);
and AND4 (N1830, N1820, N1324, N180, N205);
buf BUF1 (N1831, N1828);
not NOT1 (N1832, N1821);
or OR4 (N1833, N1823, N1325, N1132, N1001);
nor NOR2 (N1834, N1833, N364);
nand NAND3 (N1835, N1832, N1461, N779);
xor XOR2 (N1836, N1835, N1024);
xor XOR2 (N1837, N1829, N640);
not NOT1 (N1838, N1831);
nand NAND2 (N1839, N1837, N1474);
nand NAND4 (N1840, N1825, N857, N177, N1787);
not NOT1 (N1841, N1836);
buf BUF1 (N1842, N1830);
xor XOR2 (N1843, N1804, N183);
nand NAND4 (N1844, N1838, N140, N1146, N684);
or OR3 (N1845, N1822, N1742, N1512);
buf BUF1 (N1846, N1843);
nor NOR3 (N1847, N1824, N194, N1782);
nor NOR4 (N1848, N1840, N16, N98, N927);
and AND4 (N1849, N1842, N1133, N540, N1668);
and AND2 (N1850, N1844, N1811);
buf BUF1 (N1851, N1839);
nor NOR3 (N1852, N1841, N320, N1177);
and AND2 (N1853, N1849, N715);
or OR2 (N1854, N1846, N699);
nand NAND4 (N1855, N1852, N5, N1344, N1186);
nand NAND3 (N1856, N1847, N109, N1088);
xor XOR2 (N1857, N1851, N1625);
or OR3 (N1858, N1853, N49, N614);
nand NAND3 (N1859, N1848, N404, N1191);
buf BUF1 (N1860, N1856);
or OR4 (N1861, N1834, N190, N1012, N605);
or OR3 (N1862, N1845, N827, N1473);
nand NAND4 (N1863, N1862, N189, N781, N1412);
xor XOR2 (N1864, N1861, N842);
xor XOR2 (N1865, N1857, N1541);
nor NOR4 (N1866, N1855, N325, N803, N925);
and AND2 (N1867, N1860, N868);
nand NAND3 (N1868, N1866, N224, N86);
not NOT1 (N1869, N1850);
and AND2 (N1870, N1864, N569);
or OR3 (N1871, N1868, N1259, N256);
or OR2 (N1872, N1858, N1512);
nor NOR3 (N1873, N1867, N63, N382);
or OR4 (N1874, N1871, N374, N517, N1551);
or OR4 (N1875, N1870, N761, N1501, N373);
and AND3 (N1876, N1854, N1850, N739);
not NOT1 (N1877, N1875);
or OR2 (N1878, N1869, N981);
nand NAND3 (N1879, N1878, N311, N1824);
not NOT1 (N1880, N1859);
nand NAND3 (N1881, N1876, N429, N211);
xor XOR2 (N1882, N1879, N1615);
or OR2 (N1883, N1872, N353);
and AND2 (N1884, N1865, N1847);
or OR3 (N1885, N1881, N1792, N1324);
not NOT1 (N1886, N1873);
and AND2 (N1887, N1884, N1023);
or OR4 (N1888, N1883, N229, N223, N1500);
xor XOR2 (N1889, N1886, N691);
xor XOR2 (N1890, N1889, N1779);
xor XOR2 (N1891, N1885, N44);
not NOT1 (N1892, N1827);
not NOT1 (N1893, N1863);
nor NOR3 (N1894, N1882, N948, N609);
or OR2 (N1895, N1887, N1381);
and AND3 (N1896, N1890, N1495, N1282);
buf BUF1 (N1897, N1880);
nor NOR3 (N1898, N1897, N773, N724);
nor NOR2 (N1899, N1874, N1634);
or OR3 (N1900, N1888, N934, N114);
buf BUF1 (N1901, N1894);
or OR4 (N1902, N1898, N1532, N1545, N1443);
nand NAND2 (N1903, N1896, N438);
not NOT1 (N1904, N1877);
and AND3 (N1905, N1899, N1246, N341);
and AND3 (N1906, N1891, N1080, N840);
not NOT1 (N1907, N1892);
not NOT1 (N1908, N1902);
nand NAND3 (N1909, N1900, N698, N210);
or OR3 (N1910, N1895, N1284, N1743);
and AND3 (N1911, N1910, N967, N786);
and AND3 (N1912, N1906, N256, N414);
or OR3 (N1913, N1901, N470, N621);
nor NOR4 (N1914, N1909, N417, N214, N502);
xor XOR2 (N1915, N1914, N626);
or OR3 (N1916, N1911, N923, N1194);
and AND3 (N1917, N1908, N1148, N341);
and AND4 (N1918, N1915, N1765, N1710, N1401);
and AND3 (N1919, N1904, N506, N1258);
xor XOR2 (N1920, N1916, N271);
not NOT1 (N1921, N1893);
nand NAND4 (N1922, N1918, N864, N735, N854);
xor XOR2 (N1923, N1922, N1709);
nand NAND4 (N1924, N1913, N1183, N1516, N700);
xor XOR2 (N1925, N1920, N1617);
nand NAND4 (N1926, N1919, N996, N1766, N846);
and AND2 (N1927, N1917, N806);
xor XOR2 (N1928, N1905, N784);
or OR3 (N1929, N1927, N1464, N1710);
nand NAND2 (N1930, N1929, N126);
xor XOR2 (N1931, N1903, N163);
or OR4 (N1932, N1930, N95, N1383, N1192);
nor NOR2 (N1933, N1912, N140);
nor NOR2 (N1934, N1931, N1282);
not NOT1 (N1935, N1934);
nor NOR2 (N1936, N1924, N572);
nand NAND2 (N1937, N1935, N714);
xor XOR2 (N1938, N1936, N1205);
nor NOR4 (N1939, N1932, N591, N428, N1042);
not NOT1 (N1940, N1907);
nor NOR3 (N1941, N1925, N689, N479);
not NOT1 (N1942, N1941);
or OR4 (N1943, N1937, N1834, N1020, N1398);
not NOT1 (N1944, N1938);
xor XOR2 (N1945, N1933, N1516);
xor XOR2 (N1946, N1943, N1845);
buf BUF1 (N1947, N1944);
nand NAND3 (N1948, N1940, N945, N1748);
or OR2 (N1949, N1926, N302);
nand NAND3 (N1950, N1923, N204, N211);
nor NOR3 (N1951, N1946, N1296, N953);
not NOT1 (N1952, N1942);
not NOT1 (N1953, N1947);
and AND4 (N1954, N1945, N926, N960, N1649);
xor XOR2 (N1955, N1921, N1633);
buf BUF1 (N1956, N1950);
and AND4 (N1957, N1956, N1238, N1453, N1550);
xor XOR2 (N1958, N1955, N1505);
or OR4 (N1959, N1948, N1335, N1446, N1723);
and AND4 (N1960, N1951, N580, N68, N1290);
buf BUF1 (N1961, N1949);
not NOT1 (N1962, N1959);
not NOT1 (N1963, N1960);
or OR2 (N1964, N1939, N1504);
nor NOR2 (N1965, N1954, N1641);
nand NAND3 (N1966, N1957, N327, N1950);
or OR3 (N1967, N1958, N492, N283);
not NOT1 (N1968, N1963);
not NOT1 (N1969, N1964);
not NOT1 (N1970, N1965);
buf BUF1 (N1971, N1961);
xor XOR2 (N1972, N1967, N1237);
or OR4 (N1973, N1953, N1735, N752, N1621);
buf BUF1 (N1974, N1968);
xor XOR2 (N1975, N1928, N1);
buf BUF1 (N1976, N1974);
not NOT1 (N1977, N1971);
not NOT1 (N1978, N1975);
nand NAND4 (N1979, N1973, N729, N493, N1037);
buf BUF1 (N1980, N1976);
not NOT1 (N1981, N1962);
not NOT1 (N1982, N1978);
and AND2 (N1983, N1969, N1716);
nor NOR4 (N1984, N1966, N59, N821, N1564);
and AND3 (N1985, N1980, N321, N807);
xor XOR2 (N1986, N1952, N786);
and AND4 (N1987, N1972, N686, N1596, N1057);
buf BUF1 (N1988, N1987);
or OR4 (N1989, N1988, N1010, N1339, N658);
xor XOR2 (N1990, N1970, N117);
buf BUF1 (N1991, N1984);
nand NAND2 (N1992, N1990, N1950);
xor XOR2 (N1993, N1981, N153);
xor XOR2 (N1994, N1993, N1219);
not NOT1 (N1995, N1985);
nand NAND2 (N1996, N1992, N991);
buf BUF1 (N1997, N1989);
nand NAND2 (N1998, N1995, N1990);
buf BUF1 (N1999, N1994);
xor XOR2 (N2000, N1982, N582);
not NOT1 (N2001, N1983);
not NOT1 (N2002, N1991);
xor XOR2 (N2003, N1986, N1658);
not NOT1 (N2004, N1997);
buf BUF1 (N2005, N2001);
or OR3 (N2006, N2002, N1352, N1424);
not NOT1 (N2007, N2004);
xor XOR2 (N2008, N1977, N407);
and AND4 (N2009, N1979, N1129, N829, N1321);
not NOT1 (N2010, N2008);
not NOT1 (N2011, N1996);
endmodule