// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17;

output N1015,N981,N1014,N995,N1005,N998,N1009,N1010,N1016,N1017;

nor NOR4 (N18, N13, N1, N17, N15);
nor NOR2 (N19, N6, N1);
or OR3 (N20, N16, N14, N10);
or OR4 (N21, N11, N15, N11, N2);
nor NOR3 (N22, N7, N8, N5);
not NOT1 (N23, N14);
xor XOR2 (N24, N8, N5);
or OR4 (N25, N7, N15, N11, N8);
or OR4 (N26, N14, N18, N14, N21);
nand NAND4 (N27, N22, N10, N11, N20);
xor XOR2 (N28, N21, N18);
buf BUF1 (N29, N24);
nand NAND3 (N30, N23, N14, N5);
xor XOR2 (N31, N7, N16);
nand NAND2 (N32, N1, N24);
and AND2 (N33, N7, N20);
and AND4 (N34, N33, N25, N17, N29);
not NOT1 (N35, N21);
nand NAND4 (N36, N18, N21, N17, N32);
xor XOR2 (N37, N30, N22);
and AND4 (N38, N34, N28, N1, N35);
not NOT1 (N39, N34);
nand NAND3 (N40, N16, N25, N23);
not NOT1 (N41, N31);
or OR2 (N42, N4, N30);
or OR2 (N43, N19, N23);
or OR2 (N44, N36, N34);
or OR2 (N45, N38, N10);
and AND2 (N46, N40, N36);
buf BUF1 (N47, N45);
xor XOR2 (N48, N44, N29);
nor NOR4 (N49, N42, N37, N47, N20);
nor NOR2 (N50, N48, N7);
and AND3 (N51, N1, N49, N39);
buf BUF1 (N52, N3);
or OR3 (N53, N4, N41, N39);
not NOT1 (N54, N34);
xor XOR2 (N55, N23, N48);
and AND2 (N56, N54, N19);
and AND2 (N57, N50, N6);
nor NOR3 (N58, N56, N17, N42);
and AND4 (N59, N55, N37, N22, N11);
buf BUF1 (N60, N58);
and AND2 (N61, N43, N11);
and AND2 (N62, N57, N23);
buf BUF1 (N63, N53);
buf BUF1 (N64, N60);
or OR2 (N65, N26, N25);
xor XOR2 (N66, N27, N24);
or OR3 (N67, N66, N57, N10);
nor NOR2 (N68, N64, N1);
or OR2 (N69, N51, N39);
and AND4 (N70, N62, N39, N22, N53);
nand NAND3 (N71, N70, N27, N31);
buf BUF1 (N72, N68);
not NOT1 (N73, N46);
nand NAND3 (N74, N61, N26, N67);
nand NAND4 (N75, N63, N2, N55, N66);
xor XOR2 (N76, N36, N23);
xor XOR2 (N77, N76, N23);
or OR4 (N78, N65, N62, N52, N19);
xor XOR2 (N79, N46, N32);
not NOT1 (N80, N74);
xor XOR2 (N81, N73, N3);
nor NOR4 (N82, N79, N33, N4, N15);
buf BUF1 (N83, N82);
nor NOR2 (N84, N72, N25);
nand NAND3 (N85, N59, N55, N18);
and AND4 (N86, N78, N68, N71, N58);
buf BUF1 (N87, N45);
and AND4 (N88, N69, N62, N52, N24);
nand NAND4 (N89, N84, N48, N51, N11);
and AND4 (N90, N88, N11, N45, N5);
nand NAND2 (N91, N81, N34);
or OR4 (N92, N86, N55, N48, N69);
or OR4 (N93, N91, N51, N88, N52);
or OR4 (N94, N77, N36, N68, N89);
not NOT1 (N95, N40);
buf BUF1 (N96, N87);
buf BUF1 (N97, N94);
nand NAND2 (N98, N92, N93);
not NOT1 (N99, N12);
buf BUF1 (N100, N75);
or OR2 (N101, N80, N15);
nand NAND4 (N102, N90, N36, N28, N101);
buf BUF1 (N103, N34);
buf BUF1 (N104, N85);
xor XOR2 (N105, N99, N33);
not NOT1 (N106, N103);
nand NAND4 (N107, N105, N85, N75, N13);
buf BUF1 (N108, N100);
not NOT1 (N109, N96);
buf BUF1 (N110, N107);
buf BUF1 (N111, N95);
not NOT1 (N112, N83);
nand NAND4 (N113, N106, N38, N60, N28);
or OR3 (N114, N97, N27, N87);
buf BUF1 (N115, N113);
buf BUF1 (N116, N111);
or OR2 (N117, N102, N13);
nand NAND4 (N118, N114, N107, N38, N84);
and AND3 (N119, N118, N57, N26);
nor NOR4 (N120, N117, N119, N26, N98);
buf BUF1 (N121, N104);
buf BUF1 (N122, N108);
or OR3 (N123, N74, N20, N13);
or OR3 (N124, N25, N104, N115);
not NOT1 (N125, N58);
or OR4 (N126, N124, N92, N66, N82);
and AND4 (N127, N109, N124, N5, N21);
not NOT1 (N128, N120);
nand NAND3 (N129, N116, N39, N43);
xor XOR2 (N130, N123, N21);
nand NAND4 (N131, N110, N93, N88, N71);
or OR2 (N132, N121, N43);
or OR3 (N133, N127, N3, N81);
not NOT1 (N134, N132);
not NOT1 (N135, N122);
or OR4 (N136, N128, N52, N72, N26);
xor XOR2 (N137, N129, N39);
and AND4 (N138, N112, N1, N1, N10);
and AND2 (N139, N136, N34);
xor XOR2 (N140, N139, N67);
nand NAND2 (N141, N133, N55);
or OR3 (N142, N138, N74, N32);
or OR3 (N143, N137, N100, N1);
buf BUF1 (N144, N141);
not NOT1 (N145, N130);
not NOT1 (N146, N140);
nor NOR3 (N147, N144, N130, N105);
xor XOR2 (N148, N146, N32);
nor NOR3 (N149, N145, N54, N88);
and AND3 (N150, N149, N131, N134);
xor XOR2 (N151, N99, N124);
xor XOR2 (N152, N122, N80);
buf BUF1 (N153, N126);
and AND2 (N154, N152, N102);
not NOT1 (N155, N153);
nand NAND4 (N156, N135, N102, N61, N49);
buf BUF1 (N157, N148);
buf BUF1 (N158, N155);
not NOT1 (N159, N125);
buf BUF1 (N160, N154);
nand NAND3 (N161, N160, N126, N52);
and AND2 (N162, N156, N137);
not NOT1 (N163, N158);
buf BUF1 (N164, N142);
or OR4 (N165, N147, N88, N127, N130);
nand NAND4 (N166, N143, N52, N114, N10);
and AND2 (N167, N163, N47);
buf BUF1 (N168, N151);
buf BUF1 (N169, N166);
buf BUF1 (N170, N169);
xor XOR2 (N171, N162, N45);
nor NOR4 (N172, N157, N26, N93, N101);
buf BUF1 (N173, N172);
nand NAND2 (N174, N168, N9);
nor NOR2 (N175, N171, N14);
buf BUF1 (N176, N167);
nor NOR2 (N177, N150, N61);
nor NOR4 (N178, N175, N95, N128, N23);
and AND3 (N179, N170, N5, N144);
or OR4 (N180, N165, N54, N29, N132);
or OR4 (N181, N178, N116, N120, N127);
buf BUF1 (N182, N164);
nor NOR3 (N183, N174, N23, N46);
and AND3 (N184, N183, N111, N4);
and AND2 (N185, N161, N144);
not NOT1 (N186, N179);
xor XOR2 (N187, N159, N42);
buf BUF1 (N188, N184);
not NOT1 (N189, N182);
buf BUF1 (N190, N176);
nor NOR2 (N191, N185, N104);
nor NOR4 (N192, N180, N39, N149, N79);
buf BUF1 (N193, N177);
or OR4 (N194, N188, N10, N50, N37);
and AND3 (N195, N187, N88, N46);
nor NOR2 (N196, N193, N32);
and AND2 (N197, N192, N125);
and AND3 (N198, N173, N65, N8);
or OR3 (N199, N190, N125, N140);
buf BUF1 (N200, N194);
or OR2 (N201, N199, N152);
nor NOR3 (N202, N197, N104, N82);
xor XOR2 (N203, N189, N12);
xor XOR2 (N204, N195, N152);
buf BUF1 (N205, N181);
nor NOR3 (N206, N191, N96, N162);
not NOT1 (N207, N205);
xor XOR2 (N208, N203, N180);
and AND2 (N209, N204, N32);
and AND2 (N210, N200, N160);
and AND4 (N211, N207, N52, N188, N114);
not NOT1 (N212, N211);
buf BUF1 (N213, N186);
xor XOR2 (N214, N209, N180);
buf BUF1 (N215, N202);
xor XOR2 (N216, N212, N117);
or OR3 (N217, N198, N206, N152);
not NOT1 (N218, N149);
or OR4 (N219, N196, N33, N122, N77);
or OR4 (N220, N219, N45, N107, N116);
xor XOR2 (N221, N213, N127);
or OR4 (N222, N218, N200, N6, N198);
nor NOR3 (N223, N220, N217, N136);
and AND2 (N224, N125, N102);
and AND2 (N225, N208, N78);
nand NAND2 (N226, N224, N220);
not NOT1 (N227, N226);
and AND3 (N228, N225, N178, N2);
nand NAND2 (N229, N214, N183);
and AND4 (N230, N227, N134, N121, N135);
xor XOR2 (N231, N229, N98);
nand NAND3 (N232, N230, N202, N163);
or OR3 (N233, N215, N204, N61);
nor NOR2 (N234, N232, N230);
or OR4 (N235, N210, N109, N161, N214);
and AND2 (N236, N221, N44);
not NOT1 (N237, N201);
buf BUF1 (N238, N237);
or OR2 (N239, N228, N52);
or OR2 (N240, N222, N104);
nor NOR2 (N241, N216, N36);
or OR4 (N242, N240, N171, N167, N13);
xor XOR2 (N243, N231, N41);
nor NOR2 (N244, N236, N63);
nor NOR2 (N245, N235, N178);
buf BUF1 (N246, N242);
or OR3 (N247, N223, N224, N185);
or OR2 (N248, N234, N140);
nor NOR3 (N249, N233, N134, N115);
or OR3 (N250, N244, N47, N151);
xor XOR2 (N251, N239, N200);
xor XOR2 (N252, N249, N68);
buf BUF1 (N253, N248);
xor XOR2 (N254, N238, N213);
buf BUF1 (N255, N247);
not NOT1 (N256, N253);
not NOT1 (N257, N241);
xor XOR2 (N258, N255, N119);
nor NOR3 (N259, N250, N30, N124);
nand NAND4 (N260, N252, N144, N183, N7);
and AND2 (N261, N259, N43);
not NOT1 (N262, N254);
buf BUF1 (N263, N243);
nor NOR3 (N264, N263, N73, N182);
and AND4 (N265, N246, N87, N66, N109);
nand NAND3 (N266, N260, N230, N123);
nor NOR2 (N267, N266, N42);
nor NOR3 (N268, N261, N135, N209);
nor NOR2 (N269, N251, N32);
not NOT1 (N270, N256);
and AND2 (N271, N245, N252);
and AND2 (N272, N268, N241);
and AND2 (N273, N257, N258);
or OR4 (N274, N253, N40, N64, N124);
or OR4 (N275, N271, N9, N239, N209);
and AND3 (N276, N270, N112, N81);
nand NAND4 (N277, N269, N2, N127, N195);
nand NAND4 (N278, N277, N275, N32, N153);
nand NAND2 (N279, N134, N16);
nor NOR3 (N280, N265, N13, N143);
nand NAND3 (N281, N262, N278, N186);
nor NOR2 (N282, N53, N56);
xor XOR2 (N283, N264, N95);
and AND4 (N284, N267, N276, N213, N58);
not NOT1 (N285, N45);
xor XOR2 (N286, N274, N96);
nand NAND3 (N287, N282, N121, N12);
and AND4 (N288, N286, N137, N146, N80);
xor XOR2 (N289, N288, N103);
nand NAND2 (N290, N279, N237);
and AND2 (N291, N284, N266);
buf BUF1 (N292, N280);
xor XOR2 (N293, N292, N287);
nand NAND3 (N294, N58, N252, N34);
buf BUF1 (N295, N285);
xor XOR2 (N296, N289, N165);
nand NAND3 (N297, N293, N183, N44);
not NOT1 (N298, N281);
buf BUF1 (N299, N297);
not NOT1 (N300, N272);
and AND4 (N301, N283, N224, N273, N262);
not NOT1 (N302, N153);
buf BUF1 (N303, N296);
nand NAND2 (N304, N299, N189);
nor NOR3 (N305, N303, N123, N224);
buf BUF1 (N306, N302);
nand NAND2 (N307, N295, N272);
or OR4 (N308, N307, N42, N307, N289);
nor NOR2 (N309, N290, N156);
not NOT1 (N310, N301);
xor XOR2 (N311, N309, N262);
not NOT1 (N312, N310);
not NOT1 (N313, N308);
not NOT1 (N314, N291);
and AND3 (N315, N305, N136, N296);
buf BUF1 (N316, N315);
and AND4 (N317, N306, N232, N193, N111);
and AND4 (N318, N294, N193, N60, N207);
xor XOR2 (N319, N313, N78);
and AND4 (N320, N300, N203, N21, N79);
or OR4 (N321, N319, N289, N206, N94);
nor NOR4 (N322, N311, N15, N16, N246);
not NOT1 (N323, N320);
buf BUF1 (N324, N317);
and AND2 (N325, N324, N44);
nand NAND4 (N326, N321, N146, N14, N3);
not NOT1 (N327, N318);
and AND2 (N328, N304, N173);
and AND3 (N329, N328, N308, N228);
buf BUF1 (N330, N322);
nand NAND4 (N331, N312, N230, N262, N16);
not NOT1 (N332, N330);
nor NOR4 (N333, N323, N188, N36, N124);
xor XOR2 (N334, N333, N60);
buf BUF1 (N335, N331);
and AND2 (N336, N316, N196);
nand NAND4 (N337, N314, N71, N196, N116);
buf BUF1 (N338, N325);
not NOT1 (N339, N334);
xor XOR2 (N340, N298, N126);
and AND4 (N341, N326, N136, N338, N177);
nand NAND4 (N342, N183, N14, N266, N224);
buf BUF1 (N343, N327);
and AND3 (N344, N339, N244, N199);
nor NOR4 (N345, N332, N231, N128, N106);
buf BUF1 (N346, N341);
nor NOR2 (N347, N342, N183);
nor NOR2 (N348, N337, N115);
and AND4 (N349, N329, N186, N158, N8);
xor XOR2 (N350, N348, N77);
xor XOR2 (N351, N345, N200);
nor NOR2 (N352, N335, N324);
and AND2 (N353, N350, N81);
not NOT1 (N354, N347);
nand NAND4 (N355, N340, N48, N198, N42);
nand NAND2 (N356, N353, N36);
and AND4 (N357, N346, N21, N62, N35);
buf BUF1 (N358, N336);
or OR2 (N359, N344, N62);
xor XOR2 (N360, N359, N119);
and AND2 (N361, N355, N177);
nand NAND3 (N362, N357, N111, N36);
or OR4 (N363, N349, N290, N314, N210);
or OR3 (N364, N354, N94, N120);
not NOT1 (N365, N358);
nand NAND3 (N366, N360, N147, N60);
or OR3 (N367, N361, N222, N108);
xor XOR2 (N368, N362, N247);
or OR4 (N369, N352, N145, N244, N54);
buf BUF1 (N370, N368);
buf BUF1 (N371, N356);
and AND4 (N372, N351, N236, N225, N191);
xor XOR2 (N373, N366, N187);
nand NAND4 (N374, N373, N283, N313, N68);
and AND2 (N375, N364, N31);
nand NAND3 (N376, N365, N203, N27);
nand NAND2 (N377, N367, N220);
nor NOR2 (N378, N370, N104);
or OR3 (N379, N375, N284, N143);
and AND2 (N380, N378, N279);
or OR2 (N381, N377, N35);
or OR3 (N382, N363, N43, N11);
nand NAND2 (N383, N376, N378);
not NOT1 (N384, N383);
and AND3 (N385, N371, N189, N34);
not NOT1 (N386, N369);
and AND4 (N387, N381, N70, N3, N278);
and AND4 (N388, N385, N202, N312, N245);
xor XOR2 (N389, N387, N168);
not NOT1 (N390, N382);
nand NAND3 (N391, N343, N94, N384);
xor XOR2 (N392, N7, N314);
nand NAND3 (N393, N389, N265, N141);
not NOT1 (N394, N372);
not NOT1 (N395, N392);
buf BUF1 (N396, N391);
nor NOR4 (N397, N393, N140, N146, N395);
xor XOR2 (N398, N280, N77);
nand NAND3 (N399, N397, N89, N320);
not NOT1 (N400, N379);
or OR4 (N401, N390, N62, N152, N130);
or OR2 (N402, N374, N300);
nand NAND4 (N403, N400, N381, N180, N162);
xor XOR2 (N404, N403, N381);
buf BUF1 (N405, N398);
or OR2 (N406, N401, N123);
not NOT1 (N407, N399);
not NOT1 (N408, N402);
and AND4 (N409, N386, N99, N326, N50);
and AND4 (N410, N388, N78, N239, N66);
not NOT1 (N411, N407);
buf BUF1 (N412, N406);
nor NOR3 (N413, N412, N21, N329);
or OR3 (N414, N405, N227, N115);
not NOT1 (N415, N410);
buf BUF1 (N416, N409);
buf BUF1 (N417, N416);
buf BUF1 (N418, N417);
or OR4 (N419, N394, N326, N160, N385);
not NOT1 (N420, N414);
not NOT1 (N421, N408);
nor NOR4 (N422, N413, N50, N118, N365);
nand NAND4 (N423, N421, N341, N235, N126);
buf BUF1 (N424, N396);
nand NAND3 (N425, N424, N144, N267);
nand NAND4 (N426, N419, N112, N150, N421);
or OR2 (N427, N380, N324);
buf BUF1 (N428, N422);
xor XOR2 (N429, N423, N73);
buf BUF1 (N430, N425);
nor NOR2 (N431, N429, N9);
or OR3 (N432, N427, N198, N152);
and AND2 (N433, N426, N73);
buf BUF1 (N434, N428);
nor NOR3 (N435, N432, N91, N163);
and AND3 (N436, N418, N324, N417);
not NOT1 (N437, N436);
and AND4 (N438, N411, N236, N382, N39);
not NOT1 (N439, N437);
nand NAND3 (N440, N435, N229, N312);
and AND4 (N441, N404, N279, N305, N160);
or OR3 (N442, N415, N109, N238);
and AND3 (N443, N420, N408, N121);
buf BUF1 (N444, N443);
not NOT1 (N445, N442);
and AND2 (N446, N431, N175);
not NOT1 (N447, N433);
or OR3 (N448, N447, N180, N17);
nor NOR4 (N449, N439, N170, N254, N249);
or OR3 (N450, N449, N77, N228);
buf BUF1 (N451, N440);
not NOT1 (N452, N451);
nand NAND4 (N453, N430, N69, N18, N406);
nand NAND3 (N454, N441, N206, N309);
nor NOR2 (N455, N444, N65);
xor XOR2 (N456, N453, N420);
nand NAND2 (N457, N448, N443);
nand NAND2 (N458, N457, N358);
or OR2 (N459, N452, N129);
buf BUF1 (N460, N456);
nand NAND2 (N461, N458, N156);
or OR3 (N462, N434, N81, N347);
nand NAND2 (N463, N445, N337);
nor NOR3 (N464, N462, N12, N403);
not NOT1 (N465, N463);
buf BUF1 (N466, N454);
nor NOR4 (N467, N438, N297, N321, N385);
and AND2 (N468, N460, N210);
nand NAND3 (N469, N450, N343, N386);
nor NOR3 (N470, N464, N347, N117);
buf BUF1 (N471, N459);
and AND2 (N472, N469, N374);
nor NOR4 (N473, N461, N74, N357, N112);
not NOT1 (N474, N467);
not NOT1 (N475, N446);
xor XOR2 (N476, N470, N289);
or OR3 (N477, N465, N340, N110);
xor XOR2 (N478, N473, N42);
buf BUF1 (N479, N468);
not NOT1 (N480, N478);
xor XOR2 (N481, N476, N317);
buf BUF1 (N482, N472);
xor XOR2 (N483, N466, N282);
nor NOR4 (N484, N480, N75, N82, N370);
not NOT1 (N485, N481);
buf BUF1 (N486, N482);
xor XOR2 (N487, N484, N464);
and AND2 (N488, N475, N457);
and AND3 (N489, N479, N12, N467);
nand NAND4 (N490, N486, N300, N264, N489);
buf BUF1 (N491, N111);
or OR4 (N492, N477, N81, N285, N161);
or OR2 (N493, N471, N46);
xor XOR2 (N494, N491, N473);
xor XOR2 (N495, N493, N248);
or OR2 (N496, N494, N487);
xor XOR2 (N497, N210, N471);
and AND2 (N498, N496, N107);
xor XOR2 (N499, N488, N432);
not NOT1 (N500, N492);
and AND3 (N501, N490, N134, N325);
or OR2 (N502, N455, N282);
nor NOR2 (N503, N499, N91);
buf BUF1 (N504, N485);
nor NOR2 (N505, N500, N451);
not NOT1 (N506, N495);
nand NAND2 (N507, N505, N452);
and AND4 (N508, N501, N440, N103, N14);
and AND3 (N509, N506, N307, N438);
or OR3 (N510, N474, N354, N98);
nor NOR3 (N511, N502, N351, N67);
not NOT1 (N512, N497);
nor NOR2 (N513, N511, N5);
and AND2 (N514, N512, N453);
buf BUF1 (N515, N503);
not NOT1 (N516, N483);
nor NOR3 (N517, N509, N376, N75);
xor XOR2 (N518, N508, N252);
not NOT1 (N519, N516);
nor NOR4 (N520, N513, N405, N405, N385);
buf BUF1 (N521, N518);
and AND2 (N522, N519, N511);
and AND2 (N523, N507, N15);
nor NOR3 (N524, N514, N90, N452);
not NOT1 (N525, N504);
or OR2 (N526, N525, N317);
xor XOR2 (N527, N510, N455);
and AND3 (N528, N520, N449, N441);
and AND4 (N529, N517, N421, N196, N211);
nor NOR4 (N530, N521, N279, N506, N198);
xor XOR2 (N531, N528, N365);
not NOT1 (N532, N498);
and AND3 (N533, N515, N355, N86);
nand NAND2 (N534, N529, N419);
buf BUF1 (N535, N526);
or OR2 (N536, N533, N335);
and AND2 (N537, N524, N244);
xor XOR2 (N538, N523, N469);
or OR2 (N539, N536, N459);
not NOT1 (N540, N535);
and AND3 (N541, N539, N300, N114);
buf BUF1 (N542, N540);
nand NAND3 (N543, N534, N536, N531);
not NOT1 (N544, N222);
or OR3 (N545, N538, N308, N490);
nand NAND4 (N546, N542, N507, N102, N467);
nand NAND2 (N547, N545, N386);
not NOT1 (N548, N527);
nor NOR3 (N549, N532, N392, N403);
or OR4 (N550, N546, N493, N398, N38);
nand NAND4 (N551, N543, N343, N87, N523);
xor XOR2 (N552, N541, N324);
buf BUF1 (N553, N530);
nand NAND3 (N554, N547, N368, N454);
not NOT1 (N555, N554);
or OR4 (N556, N522, N186, N257, N410);
and AND3 (N557, N549, N210, N31);
nand NAND2 (N558, N552, N58);
buf BUF1 (N559, N558);
nor NOR3 (N560, N556, N101, N521);
nor NOR4 (N561, N551, N376, N371, N67);
not NOT1 (N562, N548);
nor NOR4 (N563, N555, N46, N464, N414);
xor XOR2 (N564, N537, N4);
and AND4 (N565, N557, N290, N449, N280);
and AND2 (N566, N550, N146);
xor XOR2 (N567, N560, N180);
or OR4 (N568, N565, N134, N80, N261);
or OR2 (N569, N559, N203);
xor XOR2 (N570, N563, N495);
and AND3 (N571, N561, N523, N188);
or OR4 (N572, N568, N458, N15, N335);
and AND2 (N573, N572, N512);
not NOT1 (N574, N562);
nand NAND2 (N575, N571, N499);
nand NAND3 (N576, N570, N52, N84);
nand NAND4 (N577, N575, N302, N459, N88);
nor NOR2 (N578, N564, N469);
nor NOR2 (N579, N567, N67);
and AND3 (N580, N579, N575, N239);
not NOT1 (N581, N576);
not NOT1 (N582, N544);
and AND2 (N583, N582, N327);
or OR2 (N584, N569, N533);
buf BUF1 (N585, N573);
not NOT1 (N586, N566);
or OR3 (N587, N583, N85, N498);
or OR3 (N588, N587, N240, N519);
nand NAND2 (N589, N577, N327);
not NOT1 (N590, N586);
not NOT1 (N591, N578);
buf BUF1 (N592, N589);
nor NOR4 (N593, N585, N364, N91, N101);
xor XOR2 (N594, N591, N4);
nor NOR3 (N595, N590, N270, N253);
nand NAND3 (N596, N593, N462, N131);
buf BUF1 (N597, N595);
and AND3 (N598, N594, N198, N112);
or OR4 (N599, N598, N248, N340, N369);
buf BUF1 (N600, N553);
buf BUF1 (N601, N584);
not NOT1 (N602, N588);
nand NAND2 (N603, N596, N528);
or OR4 (N604, N574, N274, N362, N201);
nor NOR4 (N605, N602, N74, N107, N229);
not NOT1 (N606, N599);
nor NOR3 (N607, N581, N110, N183);
nor NOR3 (N608, N607, N140, N269);
nor NOR4 (N609, N580, N379, N590, N546);
or OR2 (N610, N597, N558);
nand NAND4 (N611, N601, N189, N549, N141);
nand NAND4 (N612, N608, N600, N14, N228);
buf BUF1 (N613, N57);
xor XOR2 (N614, N592, N592);
nand NAND3 (N615, N612, N358, N259);
nand NAND2 (N616, N609, N41);
nor NOR2 (N617, N604, N419);
not NOT1 (N618, N610);
and AND2 (N619, N615, N197);
nand NAND2 (N620, N605, N131);
nor NOR2 (N621, N620, N197);
buf BUF1 (N622, N621);
and AND2 (N623, N616, N246);
and AND3 (N624, N617, N164, N24);
xor XOR2 (N625, N606, N291);
not NOT1 (N626, N619);
and AND4 (N627, N625, N245, N586, N192);
nor NOR2 (N628, N614, N145);
nor NOR4 (N629, N611, N295, N124, N469);
xor XOR2 (N630, N618, N55);
or OR3 (N631, N630, N550, N153);
nor NOR3 (N632, N623, N271, N306);
nor NOR4 (N633, N624, N339, N265, N82);
buf BUF1 (N634, N603);
xor XOR2 (N635, N627, N319);
or OR4 (N636, N613, N343, N570, N8);
xor XOR2 (N637, N634, N197);
and AND2 (N638, N628, N162);
nor NOR2 (N639, N638, N581);
xor XOR2 (N640, N639, N241);
nand NAND3 (N641, N626, N129, N445);
nor NOR3 (N642, N629, N525, N396);
nand NAND2 (N643, N622, N221);
or OR3 (N644, N642, N450, N241);
nor NOR4 (N645, N632, N117, N353, N178);
not NOT1 (N646, N637);
nand NAND3 (N647, N641, N64, N58);
nor NOR3 (N648, N645, N13, N608);
or OR2 (N649, N647, N320);
or OR3 (N650, N643, N627, N46);
xor XOR2 (N651, N635, N493);
nand NAND2 (N652, N648, N358);
and AND3 (N653, N631, N634, N533);
buf BUF1 (N654, N633);
buf BUF1 (N655, N651);
nand NAND4 (N656, N640, N236, N496, N646);
or OR2 (N657, N291, N203);
or OR3 (N658, N653, N459, N222);
nor NOR3 (N659, N650, N217, N209);
nand NAND2 (N660, N649, N271);
buf BUF1 (N661, N644);
nor NOR4 (N662, N636, N485, N367, N218);
buf BUF1 (N663, N654);
not NOT1 (N664, N656);
buf BUF1 (N665, N658);
nand NAND3 (N666, N655, N569, N626);
xor XOR2 (N667, N652, N316);
or OR4 (N668, N666, N59, N431, N144);
nand NAND4 (N669, N662, N568, N103, N514);
buf BUF1 (N670, N667);
and AND3 (N671, N663, N183, N432);
or OR3 (N672, N664, N113, N266);
and AND3 (N673, N670, N346, N26);
nor NOR4 (N674, N661, N329, N525, N228);
or OR3 (N675, N660, N582, N352);
buf BUF1 (N676, N665);
not NOT1 (N677, N674);
not NOT1 (N678, N677);
or OR4 (N679, N672, N289, N222, N311);
not NOT1 (N680, N669);
buf BUF1 (N681, N673);
nor NOR2 (N682, N678, N378);
nor NOR3 (N683, N676, N151, N513);
nor NOR4 (N684, N683, N497, N152, N365);
buf BUF1 (N685, N675);
not NOT1 (N686, N681);
nor NOR3 (N687, N686, N453, N485);
xor XOR2 (N688, N679, N301);
buf BUF1 (N689, N671);
nor NOR2 (N690, N689, N468);
xor XOR2 (N691, N657, N436);
nand NAND3 (N692, N687, N224, N560);
or OR2 (N693, N685, N640);
not NOT1 (N694, N659);
nor NOR4 (N695, N688, N632, N443, N386);
not NOT1 (N696, N668);
nor NOR4 (N697, N696, N25, N389, N480);
or OR4 (N698, N695, N396, N582, N425);
and AND2 (N699, N680, N49);
xor XOR2 (N700, N690, N640);
nor NOR3 (N701, N691, N321, N696);
nand NAND3 (N702, N694, N403, N123);
and AND4 (N703, N692, N207, N372, N188);
buf BUF1 (N704, N698);
or OR2 (N705, N699, N641);
nand NAND2 (N706, N703, N175);
xor XOR2 (N707, N697, N482);
or OR2 (N708, N693, N595);
buf BUF1 (N709, N701);
xor XOR2 (N710, N707, N418);
nor NOR4 (N711, N702, N19, N110, N274);
buf BUF1 (N712, N700);
nand NAND4 (N713, N712, N564, N571, N259);
or OR2 (N714, N704, N693);
buf BUF1 (N715, N709);
nor NOR3 (N716, N684, N457, N378);
and AND2 (N717, N715, N377);
nand NAND3 (N718, N708, N542, N708);
and AND4 (N719, N718, N71, N170, N520);
and AND3 (N720, N714, N412, N431);
nor NOR3 (N721, N716, N219, N601);
not NOT1 (N722, N710);
and AND2 (N723, N706, N687);
or OR2 (N724, N717, N652);
xor XOR2 (N725, N721, N620);
buf BUF1 (N726, N719);
or OR3 (N727, N705, N186, N214);
or OR2 (N728, N727, N270);
buf BUF1 (N729, N724);
nand NAND2 (N730, N723, N83);
or OR4 (N731, N720, N233, N79, N528);
buf BUF1 (N732, N731);
not NOT1 (N733, N732);
xor XOR2 (N734, N711, N688);
buf BUF1 (N735, N726);
buf BUF1 (N736, N734);
or OR2 (N737, N722, N90);
and AND2 (N738, N728, N374);
nand NAND3 (N739, N738, N113, N110);
xor XOR2 (N740, N730, N352);
buf BUF1 (N741, N739);
xor XOR2 (N742, N741, N384);
buf BUF1 (N743, N729);
buf BUF1 (N744, N743);
nand NAND4 (N745, N682, N668, N30, N702);
buf BUF1 (N746, N713);
or OR3 (N747, N746, N229, N394);
nand NAND4 (N748, N736, N715, N411, N582);
nand NAND2 (N749, N740, N255);
and AND3 (N750, N745, N461, N138);
nor NOR3 (N751, N748, N237, N427);
and AND2 (N752, N747, N231);
nand NAND2 (N753, N750, N559);
not NOT1 (N754, N752);
buf BUF1 (N755, N744);
nand NAND2 (N756, N735, N555);
xor XOR2 (N757, N751, N95);
nor NOR4 (N758, N757, N667, N580, N166);
buf BUF1 (N759, N737);
nand NAND2 (N760, N756, N77);
or OR2 (N761, N753, N119);
xor XOR2 (N762, N742, N356);
buf BUF1 (N763, N725);
nand NAND4 (N764, N762, N604, N731, N341);
or OR4 (N765, N764, N448, N351, N307);
nand NAND4 (N766, N761, N429, N756, N750);
not NOT1 (N767, N759);
xor XOR2 (N768, N765, N728);
nand NAND3 (N769, N749, N507, N396);
xor XOR2 (N770, N767, N297);
nand NAND2 (N771, N769, N372);
xor XOR2 (N772, N768, N364);
buf BUF1 (N773, N763);
buf BUF1 (N774, N766);
xor XOR2 (N775, N774, N758);
or OR3 (N776, N127, N440, N475);
buf BUF1 (N777, N771);
buf BUF1 (N778, N760);
and AND3 (N779, N733, N442, N598);
or OR2 (N780, N770, N407);
nor NOR2 (N781, N773, N661);
nand NAND4 (N782, N755, N596, N432, N38);
or OR3 (N783, N776, N462, N142);
nor NOR3 (N784, N779, N737, N366);
xor XOR2 (N785, N778, N105);
nor NOR3 (N786, N777, N382, N320);
xor XOR2 (N787, N754, N329);
nor NOR2 (N788, N782, N691);
nand NAND2 (N789, N787, N294);
nand NAND3 (N790, N788, N436, N559);
buf BUF1 (N791, N786);
xor XOR2 (N792, N781, N733);
or OR4 (N793, N785, N593, N656, N240);
not NOT1 (N794, N780);
buf BUF1 (N795, N783);
not NOT1 (N796, N793);
and AND3 (N797, N772, N393, N26);
nand NAND3 (N798, N795, N64, N113);
nand NAND3 (N799, N791, N328, N209);
xor XOR2 (N800, N799, N323);
xor XOR2 (N801, N789, N262);
nand NAND4 (N802, N796, N342, N496, N523);
nand NAND3 (N803, N775, N201, N694);
nand NAND4 (N804, N803, N98, N87, N445);
not NOT1 (N805, N784);
nand NAND2 (N806, N804, N652);
buf BUF1 (N807, N797);
and AND4 (N808, N805, N39, N320, N381);
or OR4 (N809, N800, N47, N129, N669);
nor NOR2 (N810, N806, N478);
nor NOR2 (N811, N792, N258);
or OR3 (N812, N798, N249, N577);
and AND2 (N813, N810, N578);
not NOT1 (N814, N802);
or OR4 (N815, N814, N313, N435, N97);
not NOT1 (N816, N812);
not NOT1 (N817, N816);
xor XOR2 (N818, N794, N404);
or OR3 (N819, N818, N784, N251);
and AND3 (N820, N809, N364, N743);
nor NOR3 (N821, N815, N373, N802);
not NOT1 (N822, N813);
buf BUF1 (N823, N801);
buf BUF1 (N824, N807);
xor XOR2 (N825, N820, N733);
nor NOR4 (N826, N808, N425, N223, N444);
buf BUF1 (N827, N790);
nor NOR4 (N828, N821, N49, N651, N785);
nor NOR3 (N829, N826, N419, N299);
or OR2 (N830, N811, N558);
and AND4 (N831, N828, N385, N84, N135);
and AND4 (N832, N819, N767, N396, N641);
or OR3 (N833, N830, N201, N103);
nor NOR3 (N834, N831, N603, N616);
nand NAND4 (N835, N834, N118, N363, N163);
and AND4 (N836, N832, N441, N581, N215);
nand NAND2 (N837, N829, N824);
nand NAND3 (N838, N809, N108, N831);
and AND3 (N839, N822, N404, N568);
buf BUF1 (N840, N825);
nand NAND3 (N841, N839, N257, N834);
nor NOR4 (N842, N833, N182, N481, N665);
and AND2 (N843, N842, N804);
and AND3 (N844, N823, N118, N718);
not NOT1 (N845, N837);
not NOT1 (N846, N838);
buf BUF1 (N847, N841);
nand NAND4 (N848, N836, N590, N427, N111);
not NOT1 (N849, N843);
and AND4 (N850, N840, N749, N492, N635);
not NOT1 (N851, N817);
or OR3 (N852, N827, N761, N328);
nor NOR2 (N853, N850, N98);
xor XOR2 (N854, N846, N93);
nand NAND4 (N855, N847, N39, N305, N553);
buf BUF1 (N856, N854);
xor XOR2 (N857, N855, N417);
nand NAND4 (N858, N852, N472, N566, N145);
nand NAND3 (N859, N845, N258, N632);
buf BUF1 (N860, N851);
nand NAND4 (N861, N857, N620, N515, N534);
and AND2 (N862, N860, N643);
nor NOR2 (N863, N848, N196);
nor NOR2 (N864, N859, N33);
nand NAND2 (N865, N853, N667);
buf BUF1 (N866, N856);
and AND2 (N867, N844, N578);
not NOT1 (N868, N863);
nor NOR3 (N869, N866, N757, N263);
and AND4 (N870, N862, N859, N835, N742);
nor NOR2 (N871, N389, N91);
or OR2 (N872, N868, N527);
xor XOR2 (N873, N867, N314);
nand NAND2 (N874, N865, N470);
not NOT1 (N875, N861);
and AND2 (N876, N858, N19);
nand NAND2 (N877, N870, N392);
nand NAND2 (N878, N877, N405);
nand NAND4 (N879, N873, N195, N435, N401);
and AND2 (N880, N869, N302);
xor XOR2 (N881, N849, N76);
and AND3 (N882, N875, N200, N421);
nor NOR3 (N883, N871, N664, N868);
not NOT1 (N884, N883);
nand NAND3 (N885, N874, N80, N591);
nand NAND4 (N886, N864, N648, N94, N508);
xor XOR2 (N887, N879, N253);
not NOT1 (N888, N885);
or OR2 (N889, N878, N53);
nand NAND3 (N890, N880, N485, N339);
and AND2 (N891, N884, N763);
nand NAND3 (N892, N881, N640, N702);
or OR2 (N893, N890, N339);
not NOT1 (N894, N876);
or OR2 (N895, N887, N173);
buf BUF1 (N896, N891);
nand NAND4 (N897, N882, N731, N375, N401);
and AND4 (N898, N889, N468, N255, N177);
nand NAND3 (N899, N892, N623, N198);
and AND3 (N900, N899, N377, N466);
nor NOR3 (N901, N872, N152, N508);
and AND2 (N902, N896, N583);
and AND4 (N903, N900, N154, N479, N132);
xor XOR2 (N904, N888, N397);
not NOT1 (N905, N886);
and AND3 (N906, N904, N652, N311);
xor XOR2 (N907, N902, N429);
nand NAND4 (N908, N907, N330, N840, N385);
nand NAND3 (N909, N893, N509, N430);
not NOT1 (N910, N906);
xor XOR2 (N911, N909, N720);
nor NOR2 (N912, N910, N895);
buf BUF1 (N913, N210);
nand NAND4 (N914, N903, N649, N42, N658);
or OR3 (N915, N897, N463, N50);
buf BUF1 (N916, N901);
buf BUF1 (N917, N908);
xor XOR2 (N918, N917, N843);
and AND4 (N919, N915, N274, N462, N451);
nor NOR4 (N920, N894, N239, N472, N874);
nand NAND2 (N921, N898, N526);
nand NAND4 (N922, N921, N723, N150, N156);
buf BUF1 (N923, N905);
not NOT1 (N924, N918);
nor NOR2 (N925, N924, N285);
not NOT1 (N926, N923);
not NOT1 (N927, N922);
buf BUF1 (N928, N920);
nand NAND4 (N929, N926, N120, N906, N705);
or OR2 (N930, N916, N860);
or OR4 (N931, N911, N340, N378, N113);
xor XOR2 (N932, N913, N619);
nor NOR4 (N933, N931, N215, N122, N369);
xor XOR2 (N934, N930, N525);
and AND4 (N935, N928, N23, N450, N518);
xor XOR2 (N936, N935, N346);
and AND3 (N937, N927, N60, N315);
nor NOR3 (N938, N925, N3, N928);
and AND4 (N939, N912, N753, N365, N806);
not NOT1 (N940, N932);
not NOT1 (N941, N933);
xor XOR2 (N942, N929, N624);
nor NOR4 (N943, N939, N809, N89, N84);
nor NOR3 (N944, N919, N704, N107);
and AND2 (N945, N937, N318);
nor NOR2 (N946, N943, N560);
or OR4 (N947, N936, N311, N99, N860);
buf BUF1 (N948, N945);
or OR4 (N949, N938, N279, N136, N524);
buf BUF1 (N950, N946);
nand NAND2 (N951, N950, N51);
not NOT1 (N952, N940);
buf BUF1 (N953, N947);
or OR2 (N954, N952, N529);
buf BUF1 (N955, N941);
nand NAND2 (N956, N951, N729);
and AND2 (N957, N955, N549);
and AND2 (N958, N948, N604);
and AND2 (N959, N953, N565);
nor NOR2 (N960, N949, N211);
nor NOR3 (N961, N934, N773, N431);
nor NOR3 (N962, N954, N334, N385);
buf BUF1 (N963, N960);
or OR2 (N964, N963, N919);
buf BUF1 (N965, N956);
nor NOR4 (N966, N958, N288, N300, N652);
and AND4 (N967, N965, N379, N84, N213);
xor XOR2 (N968, N961, N454);
and AND4 (N969, N968, N357, N565, N191);
or OR3 (N970, N967, N214, N69);
and AND3 (N971, N914, N66, N172);
buf BUF1 (N972, N966);
and AND2 (N973, N962, N167);
xor XOR2 (N974, N971, N298);
and AND3 (N975, N970, N259, N720);
or OR3 (N976, N957, N926, N449);
buf BUF1 (N977, N944);
buf BUF1 (N978, N972);
or OR2 (N979, N977, N536);
nand NAND3 (N980, N942, N819, N207);
not NOT1 (N981, N969);
nand NAND2 (N982, N973, N943);
buf BUF1 (N983, N975);
buf BUF1 (N984, N982);
buf BUF1 (N985, N984);
or OR3 (N986, N978, N536, N767);
or OR3 (N987, N976, N847, N425);
not NOT1 (N988, N983);
nand NAND3 (N989, N964, N370, N215);
or OR2 (N990, N987, N759);
buf BUF1 (N991, N974);
nand NAND2 (N992, N959, N207);
not NOT1 (N993, N986);
buf BUF1 (N994, N991);
nand NAND2 (N995, N992, N200);
not NOT1 (N996, N979);
buf BUF1 (N997, N994);
nand NAND4 (N998, N997, N62, N261, N935);
nor NOR4 (N999, N996, N371, N579, N303);
and AND2 (N1000, N990, N231);
and AND2 (N1001, N1000, N26);
nand NAND3 (N1002, N993, N409, N596);
and AND3 (N1003, N1002, N146, N986);
xor XOR2 (N1004, N989, N336);
or OR2 (N1005, N1004, N301);
buf BUF1 (N1006, N999);
not NOT1 (N1007, N1001);
or OR4 (N1008, N988, N615, N553, N13);
or OR4 (N1009, N985, N929, N858, N253);
nor NOR2 (N1010, N1008, N830);
and AND3 (N1011, N1003, N445, N866);
or OR2 (N1012, N980, N874);
buf BUF1 (N1013, N1006);
buf BUF1 (N1014, N1012);
or OR3 (N1015, N1007, N605, N525);
nor NOR3 (N1016, N1013, N976, N636);
and AND3 (N1017, N1011, N579, N850);
endmodule