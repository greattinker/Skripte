// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;

output N509,N512,N515,N511,N513,N516,N474,N517,N493,N518;

buf BUF1 (N19, N7);
nand NAND2 (N20, N7, N8);
nor NOR2 (N21, N6, N10);
nor NOR3 (N22, N11, N16, N7);
nand NAND3 (N23, N19, N6, N15);
not NOT1 (N24, N18);
or OR3 (N25, N15, N6, N6);
not NOT1 (N26, N11);
xor XOR2 (N27, N10, N8);
buf BUF1 (N28, N12);
nor NOR3 (N29, N3, N5, N15);
and AND4 (N30, N29, N14, N26, N14);
nor NOR4 (N31, N22, N29, N24, N4);
buf BUF1 (N32, N22);
xor XOR2 (N33, N18, N21);
nor NOR4 (N34, N7, N19, N29, N11);
buf BUF1 (N35, N32);
buf BUF1 (N36, N25);
and AND3 (N37, N20, N20, N22);
or OR2 (N38, N33, N31);
buf BUF1 (N39, N3);
and AND4 (N40, N36, N21, N23, N22);
or OR2 (N41, N19, N13);
not NOT1 (N42, N41);
or OR2 (N43, N30, N3);
or OR4 (N44, N42, N14, N40, N14);
and AND4 (N45, N44, N9, N25, N35);
and AND3 (N46, N37, N32, N30);
and AND2 (N47, N11, N11);
and AND2 (N48, N28, N14);
nand NAND2 (N49, N36, N4);
and AND2 (N50, N38, N14);
buf BUF1 (N51, N48);
and AND3 (N52, N49, N44, N22);
xor XOR2 (N53, N50, N20);
and AND3 (N54, N43, N43, N8);
nand NAND4 (N55, N52, N4, N7, N33);
nand NAND3 (N56, N53, N26, N30);
nand NAND4 (N57, N55, N12, N8, N47);
nor NOR3 (N58, N3, N23, N43);
xor XOR2 (N59, N57, N13);
nand NAND4 (N60, N45, N3, N16, N10);
buf BUF1 (N61, N51);
nand NAND4 (N62, N39, N40, N32, N44);
or OR3 (N63, N61, N52, N24);
xor XOR2 (N64, N34, N34);
and AND4 (N65, N46, N50, N21, N19);
and AND4 (N66, N65, N17, N35, N35);
or OR4 (N67, N62, N17, N33, N28);
xor XOR2 (N68, N67, N17);
nor NOR2 (N69, N68, N32);
nand NAND3 (N70, N64, N28, N34);
or OR4 (N71, N60, N62, N20, N4);
not NOT1 (N72, N63);
or OR2 (N73, N66, N2);
not NOT1 (N74, N56);
nand NAND3 (N75, N71, N35, N18);
nor NOR3 (N76, N58, N30, N44);
nand NAND4 (N77, N74, N71, N68, N32);
buf BUF1 (N78, N69);
not NOT1 (N79, N78);
xor XOR2 (N80, N75, N70);
buf BUF1 (N81, N17);
not NOT1 (N82, N81);
xor XOR2 (N83, N82, N1);
not NOT1 (N84, N27);
buf BUF1 (N85, N83);
buf BUF1 (N86, N79);
or OR3 (N87, N77, N1, N16);
nor NOR3 (N88, N54, N55, N49);
buf BUF1 (N89, N59);
not NOT1 (N90, N88);
and AND3 (N91, N85, N60, N55);
not NOT1 (N92, N73);
or OR4 (N93, N92, N80, N5, N13);
or OR2 (N94, N90, N22);
buf BUF1 (N95, N33);
or OR3 (N96, N93, N7, N41);
nand NAND3 (N97, N87, N89, N5);
xor XOR2 (N98, N36, N3);
not NOT1 (N99, N72);
xor XOR2 (N100, N86, N8);
nand NAND2 (N101, N97, N87);
xor XOR2 (N102, N84, N30);
nand NAND4 (N103, N99, N82, N102, N59);
nor NOR4 (N104, N100, N60, N73, N9);
nor NOR3 (N105, N82, N36, N27);
not NOT1 (N106, N98);
nand NAND3 (N107, N91, N42, N65);
xor XOR2 (N108, N76, N35);
or OR2 (N109, N94, N87);
nand NAND3 (N110, N108, N47, N105);
and AND3 (N111, N34, N27, N27);
not NOT1 (N112, N107);
nand NAND4 (N113, N112, N88, N53, N45);
or OR2 (N114, N101, N73);
and AND4 (N115, N111, N108, N73, N109);
nor NOR3 (N116, N59, N31, N88);
and AND4 (N117, N103, N2, N13, N69);
buf BUF1 (N118, N96);
xor XOR2 (N119, N115, N13);
nand NAND3 (N120, N114, N54, N96);
not NOT1 (N121, N104);
nand NAND2 (N122, N119, N67);
not NOT1 (N123, N106);
xor XOR2 (N124, N116, N108);
nand NAND2 (N125, N121, N90);
buf BUF1 (N126, N95);
nand NAND4 (N127, N117, N76, N79, N66);
nand NAND2 (N128, N118, N32);
buf BUF1 (N129, N126);
nand NAND3 (N130, N124, N113, N95);
nand NAND2 (N131, N55, N100);
or OR3 (N132, N110, N15, N50);
or OR2 (N133, N125, N112);
and AND2 (N134, N131, N7);
or OR4 (N135, N122, N124, N76, N55);
nor NOR2 (N136, N120, N124);
not NOT1 (N137, N129);
nor NOR3 (N138, N135, N69, N58);
not NOT1 (N139, N133);
buf BUF1 (N140, N138);
xor XOR2 (N141, N128, N13);
or OR3 (N142, N141, N22, N70);
and AND2 (N143, N123, N76);
nor NOR2 (N144, N137, N28);
nor NOR4 (N145, N144, N40, N34, N23);
or OR3 (N146, N136, N1, N41);
nor NOR4 (N147, N145, N80, N145, N33);
buf BUF1 (N148, N147);
not NOT1 (N149, N142);
nor NOR4 (N150, N127, N66, N131, N23);
nor NOR4 (N151, N134, N120, N111, N129);
nand NAND4 (N152, N150, N83, N61, N98);
nor NOR2 (N153, N143, N54);
nor NOR4 (N154, N151, N55, N91, N4);
not NOT1 (N155, N149);
nor NOR4 (N156, N130, N63, N101, N50);
nand NAND4 (N157, N132, N36, N146, N12);
and AND2 (N158, N153, N11);
buf BUF1 (N159, N136);
nand NAND4 (N160, N154, N80, N121, N82);
and AND3 (N161, N155, N76, N104);
not NOT1 (N162, N148);
xor XOR2 (N163, N160, N48);
buf BUF1 (N164, N158);
not NOT1 (N165, N162);
not NOT1 (N166, N164);
buf BUF1 (N167, N159);
buf BUF1 (N168, N157);
or OR3 (N169, N163, N100, N97);
nor NOR4 (N170, N169, N5, N6, N11);
nand NAND4 (N171, N166, N151, N94, N96);
xor XOR2 (N172, N152, N60);
buf BUF1 (N173, N167);
buf BUF1 (N174, N172);
nand NAND4 (N175, N161, N54, N89, N10);
not NOT1 (N176, N156);
xor XOR2 (N177, N174, N8);
not NOT1 (N178, N171);
not NOT1 (N179, N170);
buf BUF1 (N180, N139);
buf BUF1 (N181, N179);
not NOT1 (N182, N173);
and AND3 (N183, N180, N29, N103);
and AND4 (N184, N165, N145, N135, N103);
nor NOR4 (N185, N168, N133, N172, N142);
buf BUF1 (N186, N175);
or OR3 (N187, N182, N121, N20);
or OR4 (N188, N183, N139, N25, N52);
or OR3 (N189, N176, N158, N149);
nor NOR4 (N190, N181, N22, N81, N28);
xor XOR2 (N191, N186, N90);
nand NAND4 (N192, N178, N58, N182, N160);
and AND4 (N193, N185, N101, N108, N81);
nand NAND4 (N194, N189, N60, N12, N27);
nand NAND2 (N195, N188, N74);
and AND2 (N196, N184, N75);
or OR4 (N197, N191, N49, N37, N147);
buf BUF1 (N198, N140);
nand NAND3 (N199, N187, N187, N26);
and AND3 (N200, N198, N175, N21);
buf BUF1 (N201, N200);
or OR4 (N202, N199, N164, N82, N82);
nand NAND4 (N203, N196, N108, N81, N114);
xor XOR2 (N204, N195, N199);
buf BUF1 (N205, N177);
nand NAND3 (N206, N194, N69, N135);
nand NAND4 (N207, N197, N191, N122, N91);
not NOT1 (N208, N205);
and AND3 (N209, N208, N174, N116);
buf BUF1 (N210, N192);
and AND4 (N211, N203, N78, N149, N41);
nor NOR2 (N212, N209, N211);
nand NAND4 (N213, N87, N203, N165, N111);
nor NOR3 (N214, N202, N59, N123);
xor XOR2 (N215, N201, N117);
nor NOR4 (N216, N214, N5, N8, N197);
buf BUF1 (N217, N212);
xor XOR2 (N218, N210, N202);
nor NOR2 (N219, N193, N31);
not NOT1 (N220, N207);
not NOT1 (N221, N219);
nand NAND4 (N222, N218, N206, N128, N112);
xor XOR2 (N223, N92, N38);
or OR2 (N224, N204, N23);
nand NAND2 (N225, N221, N82);
and AND4 (N226, N225, N132, N186, N121);
nand NAND3 (N227, N222, N197, N169);
nand NAND4 (N228, N224, N49, N47, N48);
not NOT1 (N229, N217);
nand NAND4 (N230, N223, N173, N106, N47);
or OR4 (N231, N226, N31, N29, N221);
buf BUF1 (N232, N215);
nand NAND3 (N233, N220, N95, N8);
nand NAND4 (N234, N213, N189, N161, N221);
xor XOR2 (N235, N229, N33);
nand NAND4 (N236, N232, N147, N124, N218);
xor XOR2 (N237, N216, N35);
and AND3 (N238, N230, N11, N103);
xor XOR2 (N239, N236, N160);
buf BUF1 (N240, N227);
and AND4 (N241, N235, N85, N176, N167);
buf BUF1 (N242, N190);
nand NAND4 (N243, N241, N43, N61, N169);
and AND3 (N244, N228, N183, N138);
xor XOR2 (N245, N237, N142);
nand NAND2 (N246, N231, N210);
xor XOR2 (N247, N245, N206);
not NOT1 (N248, N243);
not NOT1 (N249, N240);
or OR4 (N250, N238, N238, N47, N150);
buf BUF1 (N251, N247);
xor XOR2 (N252, N242, N150);
buf BUF1 (N253, N249);
or OR2 (N254, N251, N100);
nand NAND3 (N255, N253, N142, N145);
or OR2 (N256, N248, N61);
not NOT1 (N257, N246);
or OR2 (N258, N256, N143);
not NOT1 (N259, N234);
nand NAND3 (N260, N255, N54, N14);
or OR2 (N261, N252, N260);
not NOT1 (N262, N123);
and AND3 (N263, N259, N172, N71);
xor XOR2 (N264, N244, N142);
xor XOR2 (N265, N239, N258);
not NOT1 (N266, N14);
xor XOR2 (N267, N257, N47);
xor XOR2 (N268, N264, N202);
not NOT1 (N269, N268);
buf BUF1 (N270, N262);
or OR4 (N271, N266, N210, N98, N82);
buf BUF1 (N272, N265);
nand NAND4 (N273, N270, N149, N128, N9);
nand NAND2 (N274, N269, N173);
xor XOR2 (N275, N274, N151);
nor NOR2 (N276, N271, N205);
not NOT1 (N277, N267);
nor NOR2 (N278, N263, N75);
nand NAND3 (N279, N250, N139, N73);
nor NOR2 (N280, N277, N24);
nand NAND3 (N281, N275, N197, N83);
nor NOR4 (N282, N233, N113, N239, N128);
xor XOR2 (N283, N254, N274);
or OR3 (N284, N273, N172, N36);
buf BUF1 (N285, N276);
nand NAND3 (N286, N279, N195, N75);
or OR4 (N287, N286, N208, N9, N73);
xor XOR2 (N288, N280, N278);
nor NOR2 (N289, N111, N148);
nand NAND2 (N290, N285, N154);
nor NOR2 (N291, N289, N26);
xor XOR2 (N292, N284, N203);
buf BUF1 (N293, N283);
nor NOR4 (N294, N261, N230, N251, N127);
nand NAND3 (N295, N290, N21, N252);
not NOT1 (N296, N282);
buf BUF1 (N297, N291);
xor XOR2 (N298, N292, N24);
not NOT1 (N299, N298);
buf BUF1 (N300, N288);
xor XOR2 (N301, N297, N197);
not NOT1 (N302, N295);
buf BUF1 (N303, N272);
nand NAND2 (N304, N301, N205);
nand NAND3 (N305, N304, N170, N110);
and AND3 (N306, N294, N146, N29);
not NOT1 (N307, N296);
xor XOR2 (N308, N293, N102);
nand NAND3 (N309, N305, N306, N249);
not NOT1 (N310, N46);
buf BUF1 (N311, N300);
xor XOR2 (N312, N307, N18);
xor XOR2 (N313, N312, N16);
nand NAND3 (N314, N310, N293, N15);
not NOT1 (N315, N281);
and AND2 (N316, N302, N120);
not NOT1 (N317, N309);
buf BUF1 (N318, N287);
nand NAND3 (N319, N308, N122, N311);
nor NOR4 (N320, N27, N235, N304, N28);
xor XOR2 (N321, N303, N305);
xor XOR2 (N322, N318, N245);
and AND2 (N323, N315, N113);
nand NAND3 (N324, N321, N206, N236);
not NOT1 (N325, N317);
nor NOR4 (N326, N320, N121, N231, N302);
and AND4 (N327, N314, N142, N307, N173);
not NOT1 (N328, N326);
nor NOR4 (N329, N316, N70, N11, N67);
not NOT1 (N330, N324);
xor XOR2 (N331, N313, N316);
not NOT1 (N332, N299);
and AND2 (N333, N328, N261);
or OR2 (N334, N330, N74);
nor NOR4 (N335, N322, N137, N201, N172);
xor XOR2 (N336, N329, N104);
not NOT1 (N337, N319);
nand NAND3 (N338, N323, N276, N35);
xor XOR2 (N339, N338, N268);
not NOT1 (N340, N327);
xor XOR2 (N341, N336, N105);
xor XOR2 (N342, N334, N7);
nand NAND4 (N343, N342, N34, N296, N17);
xor XOR2 (N344, N335, N76);
nand NAND3 (N345, N332, N215, N138);
and AND2 (N346, N331, N133);
or OR4 (N347, N325, N229, N125, N103);
buf BUF1 (N348, N340);
nand NAND3 (N349, N339, N187, N1);
and AND4 (N350, N337, N240, N61, N197);
buf BUF1 (N351, N343);
and AND4 (N352, N351, N78, N14, N224);
and AND2 (N353, N348, N219);
not NOT1 (N354, N353);
or OR3 (N355, N350, N341, N327);
nand NAND3 (N356, N301, N62, N337);
xor XOR2 (N357, N346, N133);
nor NOR3 (N358, N355, N135, N27);
buf BUF1 (N359, N349);
buf BUF1 (N360, N356);
nand NAND3 (N361, N354, N25, N270);
nand NAND2 (N362, N357, N272);
buf BUF1 (N363, N362);
nand NAND3 (N364, N363, N274, N80);
not NOT1 (N365, N361);
buf BUF1 (N366, N359);
or OR2 (N367, N358, N151);
buf BUF1 (N368, N352);
or OR2 (N369, N360, N344);
nand NAND3 (N370, N333, N203, N69);
and AND2 (N371, N210, N136);
buf BUF1 (N372, N345);
not NOT1 (N373, N347);
buf BUF1 (N374, N365);
nor NOR3 (N375, N371, N189, N75);
or OR3 (N376, N372, N263, N144);
nor NOR3 (N377, N369, N185, N125);
or OR2 (N378, N375, N217);
or OR2 (N379, N367, N106);
nand NAND2 (N380, N373, N24);
nor NOR4 (N381, N364, N193, N284, N117);
buf BUF1 (N382, N379);
nand NAND3 (N383, N370, N302, N304);
xor XOR2 (N384, N382, N159);
or OR4 (N385, N381, N277, N310, N315);
buf BUF1 (N386, N384);
nand NAND2 (N387, N378, N220);
and AND4 (N388, N366, N197, N123, N227);
and AND3 (N389, N374, N243, N90);
and AND3 (N390, N377, N197, N111);
or OR3 (N391, N386, N353, N82);
nor NOR3 (N392, N387, N23, N236);
nor NOR3 (N393, N388, N25, N138);
nand NAND2 (N394, N383, N306);
or OR2 (N395, N385, N315);
not NOT1 (N396, N368);
and AND3 (N397, N396, N278, N71);
nand NAND3 (N398, N393, N196, N112);
not NOT1 (N399, N398);
nor NOR3 (N400, N399, N306, N392);
xor XOR2 (N401, N74, N59);
or OR3 (N402, N390, N145, N122);
not NOT1 (N403, N397);
or OR4 (N404, N400, N37, N24, N138);
nor NOR2 (N405, N380, N103);
xor XOR2 (N406, N389, N181);
nor NOR4 (N407, N394, N20, N55, N117);
nand NAND4 (N408, N376, N326, N168, N156);
or OR2 (N409, N408, N49);
or OR2 (N410, N407, N158);
not NOT1 (N411, N409);
buf BUF1 (N412, N391);
nand NAND2 (N413, N404, N206);
xor XOR2 (N414, N402, N35);
and AND4 (N415, N401, N157, N400, N354);
and AND2 (N416, N403, N195);
nor NOR2 (N417, N414, N194);
nor NOR3 (N418, N416, N326, N220);
nand NAND3 (N419, N405, N369, N351);
nand NAND2 (N420, N413, N100);
nor NOR4 (N421, N415, N35, N289, N305);
or OR2 (N422, N412, N39);
not NOT1 (N423, N395);
buf BUF1 (N424, N406);
nor NOR3 (N425, N422, N388, N132);
and AND4 (N426, N419, N252, N74, N70);
not NOT1 (N427, N425);
buf BUF1 (N428, N427);
nor NOR2 (N429, N426, N331);
and AND3 (N430, N417, N323, N156);
nor NOR4 (N431, N430, N343, N21, N333);
xor XOR2 (N432, N421, N357);
nor NOR2 (N433, N418, N199);
nor NOR4 (N434, N432, N349, N156, N404);
nor NOR4 (N435, N433, N425, N426, N85);
nor NOR2 (N436, N431, N28);
and AND3 (N437, N410, N345, N339);
and AND2 (N438, N436, N325);
nand NAND3 (N439, N420, N89, N45);
not NOT1 (N440, N423);
and AND2 (N441, N428, N82);
nor NOR2 (N442, N440, N161);
nand NAND4 (N443, N441, N160, N195, N58);
not NOT1 (N444, N434);
xor XOR2 (N445, N435, N375);
nand NAND2 (N446, N429, N3);
not NOT1 (N447, N445);
and AND2 (N448, N443, N401);
buf BUF1 (N449, N439);
or OR4 (N450, N442, N261, N157, N364);
not NOT1 (N451, N437);
nand NAND2 (N452, N449, N227);
buf BUF1 (N453, N447);
buf BUF1 (N454, N452);
nor NOR2 (N455, N453, N75);
not NOT1 (N456, N454);
and AND3 (N457, N446, N423, N383);
xor XOR2 (N458, N455, N229);
and AND3 (N459, N450, N401, N275);
not NOT1 (N460, N456);
not NOT1 (N461, N438);
nand NAND2 (N462, N460, N51);
buf BUF1 (N463, N444);
xor XOR2 (N464, N411, N90);
or OR4 (N465, N451, N444, N413, N109);
nand NAND3 (N466, N464, N370, N42);
nand NAND4 (N467, N458, N417, N8, N393);
and AND4 (N468, N463, N165, N443, N60);
xor XOR2 (N469, N467, N95);
and AND3 (N470, N469, N455, N267);
or OR4 (N471, N424, N222, N110, N48);
or OR2 (N472, N470, N391);
buf BUF1 (N473, N462);
not NOT1 (N474, N466);
or OR4 (N475, N472, N199, N32, N282);
not NOT1 (N476, N465);
nand NAND4 (N477, N457, N224, N331, N173);
xor XOR2 (N478, N477, N312);
nand NAND3 (N479, N475, N255, N299);
xor XOR2 (N480, N468, N417);
xor XOR2 (N481, N480, N353);
xor XOR2 (N482, N459, N378);
not NOT1 (N483, N478);
nand NAND2 (N484, N483, N113);
not NOT1 (N485, N484);
nand NAND4 (N486, N471, N311, N182, N216);
nor NOR3 (N487, N479, N354, N239);
not NOT1 (N488, N481);
and AND4 (N489, N482, N270, N106, N453);
xor XOR2 (N490, N485, N190);
not NOT1 (N491, N461);
or OR2 (N492, N491, N381);
buf BUF1 (N493, N492);
nor NOR3 (N494, N473, N124, N390);
xor XOR2 (N495, N476, N11);
nor NOR4 (N496, N486, N55, N388, N155);
or OR2 (N497, N448, N209);
nand NAND3 (N498, N490, N418, N105);
buf BUF1 (N499, N488);
not NOT1 (N500, N494);
buf BUF1 (N501, N497);
xor XOR2 (N502, N489, N28);
not NOT1 (N503, N487);
nand NAND4 (N504, N498, N454, N285, N142);
xor XOR2 (N505, N495, N298);
and AND4 (N506, N499, N280, N412, N380);
buf BUF1 (N507, N505);
or OR2 (N508, N500, N323);
xor XOR2 (N509, N507, N79);
nand NAND3 (N510, N502, N502, N347);
and AND3 (N511, N501, N110, N465);
nor NOR3 (N512, N510, N8, N62);
buf BUF1 (N513, N503);
xor XOR2 (N514, N506, N120);
and AND2 (N515, N514, N390);
or OR2 (N516, N504, N453);
nor NOR4 (N517, N496, N100, N317, N10);
nor NOR3 (N518, N508, N115, N142);
endmodule