// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10;

output N3508,N3504,N3506,N3479,N3498,N3485,N3475,N3502,N3509,N3510;

not NOT1 (N11, N8);
and AND2 (N12, N8, N4);
or OR3 (N13, N10, N2, N2);
or OR4 (N14, N4, N3, N4, N1);
not NOT1 (N15, N6);
nand NAND3 (N16, N4, N7, N10);
xor XOR2 (N17, N11, N5);
and AND3 (N18, N15, N15, N5);
nor NOR3 (N19, N10, N14, N4);
xor XOR2 (N20, N9, N18);
nor NOR3 (N21, N2, N10, N11);
nand NAND2 (N22, N5, N1);
xor XOR2 (N23, N22, N5);
or OR3 (N24, N16, N6, N19);
nand NAND3 (N25, N24, N1, N3);
and AND4 (N26, N23, N14, N10, N23);
not NOT1 (N27, N26);
not NOT1 (N28, N3);
or OR2 (N29, N19, N1);
xor XOR2 (N30, N18, N9);
and AND2 (N31, N25, N5);
xor XOR2 (N32, N31, N23);
nand NAND4 (N33, N13, N14, N21, N11);
nand NAND2 (N34, N22, N25);
buf BUF1 (N35, N17);
or OR2 (N36, N12, N14);
buf BUF1 (N37, N32);
nor NOR2 (N38, N28, N3);
and AND4 (N39, N34, N28, N4, N4);
or OR3 (N40, N36, N27, N19);
nor NOR4 (N41, N37, N35, N4, N4);
or OR3 (N42, N24, N19, N27);
or OR4 (N43, N2, N33, N33, N25);
and AND3 (N44, N15, N30, N34);
not NOT1 (N45, N16);
nand NAND3 (N46, N29, N9, N36);
or OR2 (N47, N43, N7);
nand NAND3 (N48, N39, N15, N33);
nor NOR4 (N49, N48, N31, N38, N24);
xor XOR2 (N50, N41, N24);
nand NAND4 (N51, N38, N47, N10, N6);
nand NAND3 (N52, N42, N41, N11);
nand NAND3 (N53, N20, N19, N37);
xor XOR2 (N54, N13, N15);
or OR4 (N55, N51, N5, N34, N23);
and AND2 (N56, N40, N20);
and AND3 (N57, N50, N16, N31);
and AND3 (N58, N44, N53, N15);
nor NOR4 (N59, N41, N50, N57, N24);
and AND4 (N60, N33, N39, N33, N15);
buf BUF1 (N61, N55);
or OR2 (N62, N59, N46);
not NOT1 (N63, N31);
not NOT1 (N64, N49);
and AND4 (N65, N64, N21, N29, N23);
buf BUF1 (N66, N63);
or OR3 (N67, N56, N60, N45);
xor XOR2 (N68, N35, N40);
not NOT1 (N69, N27);
or OR2 (N70, N58, N23);
nor NOR2 (N71, N66, N32);
or OR3 (N72, N54, N23, N12);
nor NOR2 (N73, N52, N57);
nor NOR2 (N74, N68, N64);
xor XOR2 (N75, N72, N69);
and AND2 (N76, N16, N11);
nand NAND2 (N77, N62, N25);
nand NAND2 (N78, N76, N75);
or OR4 (N79, N29, N5, N28, N11);
not NOT1 (N80, N65);
buf BUF1 (N81, N71);
buf BUF1 (N82, N79);
xor XOR2 (N83, N80, N22);
xor XOR2 (N84, N70, N47);
and AND3 (N85, N84, N37, N15);
and AND3 (N86, N73, N49, N62);
nor NOR2 (N87, N77, N48);
and AND4 (N88, N78, N22, N81, N57);
not NOT1 (N89, N67);
nor NOR2 (N90, N28, N18);
and AND3 (N91, N86, N24, N83);
or OR3 (N92, N51, N50, N70);
buf BUF1 (N93, N85);
or OR2 (N94, N90, N45);
or OR2 (N95, N61, N10);
xor XOR2 (N96, N82, N13);
and AND3 (N97, N91, N62, N84);
nand NAND4 (N98, N96, N38, N91, N60);
and AND3 (N99, N95, N65, N36);
not NOT1 (N100, N93);
not NOT1 (N101, N74);
nand NAND3 (N102, N97, N75, N41);
buf BUF1 (N103, N87);
and AND3 (N104, N92, N28, N45);
nor NOR2 (N105, N104, N60);
not NOT1 (N106, N94);
not NOT1 (N107, N105);
buf BUF1 (N108, N101);
not NOT1 (N109, N88);
not NOT1 (N110, N106);
nand NAND3 (N111, N102, N61, N25);
and AND2 (N112, N100, N32);
or OR2 (N113, N107, N50);
nand NAND3 (N114, N110, N64, N69);
or OR4 (N115, N113, N10, N4, N4);
buf BUF1 (N116, N89);
not NOT1 (N117, N116);
not NOT1 (N118, N103);
nor NOR3 (N119, N114, N65, N22);
and AND3 (N120, N109, N61, N63);
not NOT1 (N121, N119);
nor NOR3 (N122, N115, N19, N33);
not NOT1 (N123, N121);
nand NAND2 (N124, N98, N98);
xor XOR2 (N125, N112, N120);
and AND4 (N126, N105, N34, N111, N103);
nand NAND2 (N127, N101, N97);
or OR3 (N128, N123, N74, N84);
and AND4 (N129, N124, N63, N26, N124);
nor NOR3 (N130, N118, N36, N9);
and AND2 (N131, N130, N64);
and AND3 (N132, N122, N91, N65);
and AND3 (N133, N126, N15, N27);
xor XOR2 (N134, N131, N128);
not NOT1 (N135, N102);
xor XOR2 (N136, N127, N100);
or OR2 (N137, N117, N121);
xor XOR2 (N138, N134, N76);
not NOT1 (N139, N138);
not NOT1 (N140, N125);
not NOT1 (N141, N140);
not NOT1 (N142, N129);
nor NOR4 (N143, N137, N97, N49, N61);
not NOT1 (N144, N141);
nand NAND2 (N145, N142, N127);
nand NAND3 (N146, N145, N60, N137);
and AND3 (N147, N133, N78, N145);
buf BUF1 (N148, N139);
not NOT1 (N149, N108);
nand NAND3 (N150, N149, N43, N113);
and AND4 (N151, N136, N89, N11, N26);
xor XOR2 (N152, N143, N104);
not NOT1 (N153, N99);
not NOT1 (N154, N153);
not NOT1 (N155, N150);
nand NAND4 (N156, N151, N37, N89, N145);
or OR2 (N157, N155, N125);
buf BUF1 (N158, N157);
nor NOR4 (N159, N132, N106, N49, N1);
and AND2 (N160, N158, N113);
nor NOR4 (N161, N144, N39, N63, N9);
buf BUF1 (N162, N156);
or OR4 (N163, N148, N116, N125, N2);
or OR3 (N164, N154, N122, N141);
nand NAND4 (N165, N147, N154, N62, N46);
xor XOR2 (N166, N165, N103);
and AND3 (N167, N146, N40, N145);
not NOT1 (N168, N160);
or OR2 (N169, N166, N57);
not NOT1 (N170, N164);
nand NAND3 (N171, N161, N18, N46);
buf BUF1 (N172, N159);
or OR3 (N173, N152, N114, N152);
and AND2 (N174, N172, N109);
xor XOR2 (N175, N167, N39);
or OR4 (N176, N174, N36, N131, N31);
buf BUF1 (N177, N135);
and AND4 (N178, N175, N126, N129, N114);
and AND2 (N179, N178, N118);
xor XOR2 (N180, N163, N59);
not NOT1 (N181, N171);
or OR3 (N182, N173, N156, N59);
not NOT1 (N183, N182);
nand NAND4 (N184, N176, N25, N18, N77);
and AND3 (N185, N183, N78, N27);
nand NAND4 (N186, N177, N39, N27, N104);
buf BUF1 (N187, N162);
xor XOR2 (N188, N181, N165);
or OR3 (N189, N179, N141, N4);
and AND2 (N190, N186, N3);
not NOT1 (N191, N168);
nand NAND4 (N192, N185, N47, N94, N117);
nand NAND3 (N193, N170, N16, N66);
and AND4 (N194, N193, N85, N159, N184);
nor NOR4 (N195, N187, N52, N155, N28);
nand NAND2 (N196, N176, N170);
and AND2 (N197, N188, N102);
not NOT1 (N198, N196);
not NOT1 (N199, N192);
nor NOR3 (N200, N197, N142, N65);
xor XOR2 (N201, N189, N152);
buf BUF1 (N202, N199);
nand NAND4 (N203, N195, N6, N55, N152);
nor NOR3 (N204, N180, N192, N183);
buf BUF1 (N205, N204);
and AND2 (N206, N202, N84);
not NOT1 (N207, N191);
not NOT1 (N208, N207);
not NOT1 (N209, N208);
nand NAND3 (N210, N205, N37, N97);
nand NAND2 (N211, N200, N129);
and AND3 (N212, N169, N137, N181);
not NOT1 (N213, N190);
not NOT1 (N214, N203);
not NOT1 (N215, N212);
buf BUF1 (N216, N213);
xor XOR2 (N217, N215, N96);
xor XOR2 (N218, N210, N117);
or OR2 (N219, N209, N86);
or OR3 (N220, N206, N198, N29);
nand NAND3 (N221, N35, N49, N51);
not NOT1 (N222, N217);
or OR4 (N223, N216, N215, N36, N106);
xor XOR2 (N224, N220, N117);
nor NOR3 (N225, N218, N34, N222);
and AND4 (N226, N150, N79, N67, N140);
xor XOR2 (N227, N221, N92);
xor XOR2 (N228, N219, N93);
and AND4 (N229, N226, N7, N211, N41);
nor NOR4 (N230, N57, N169, N225, N199);
xor XOR2 (N231, N187, N30);
xor XOR2 (N232, N230, N85);
nand NAND4 (N233, N228, N12, N152, N94);
nor NOR2 (N234, N227, N229);
nor NOR4 (N235, N134, N3, N143, N187);
nor NOR2 (N236, N201, N41);
not NOT1 (N237, N232);
or OR2 (N238, N194, N171);
xor XOR2 (N239, N233, N174);
not NOT1 (N240, N236);
not NOT1 (N241, N234);
and AND4 (N242, N239, N67, N169, N73);
nand NAND3 (N243, N242, N73, N145);
and AND4 (N244, N237, N230, N15, N225);
nand NAND4 (N245, N224, N162, N79, N185);
nand NAND4 (N246, N231, N245, N174, N54);
or OR2 (N247, N20, N90);
and AND4 (N248, N246, N139, N207, N212);
not NOT1 (N249, N247);
buf BUF1 (N250, N249);
xor XOR2 (N251, N250, N163);
xor XOR2 (N252, N240, N165);
and AND4 (N253, N251, N216, N194, N89);
or OR4 (N254, N238, N140, N199, N149);
nand NAND2 (N255, N248, N192);
nand NAND4 (N256, N255, N248, N161, N214);
nand NAND4 (N257, N22, N17, N33, N6);
and AND3 (N258, N241, N73, N58);
and AND2 (N259, N244, N56);
or OR4 (N260, N254, N185, N22, N174);
or OR4 (N261, N259, N198, N159, N88);
buf BUF1 (N262, N223);
nand NAND3 (N263, N235, N46, N218);
buf BUF1 (N264, N256);
nand NAND4 (N265, N243, N106, N68, N165);
and AND3 (N266, N257, N167, N62);
and AND3 (N267, N263, N49, N189);
and AND4 (N268, N266, N118, N102, N11);
nand NAND4 (N269, N260, N93, N248, N90);
and AND4 (N270, N253, N51, N126, N41);
xor XOR2 (N271, N269, N125);
and AND4 (N272, N262, N121, N98, N161);
or OR4 (N273, N271, N6, N220, N203);
buf BUF1 (N274, N273);
nor NOR2 (N275, N270, N166);
xor XOR2 (N276, N274, N269);
nand NAND4 (N277, N252, N122, N14, N84);
or OR3 (N278, N258, N224, N266);
not NOT1 (N279, N267);
nand NAND3 (N280, N272, N205, N8);
not NOT1 (N281, N261);
not NOT1 (N282, N278);
and AND3 (N283, N277, N72, N64);
and AND2 (N284, N281, N91);
buf BUF1 (N285, N282);
or OR2 (N286, N276, N176);
buf BUF1 (N287, N279);
nor NOR2 (N288, N280, N230);
and AND4 (N289, N285, N192, N272, N267);
not NOT1 (N290, N264);
and AND2 (N291, N286, N275);
nor NOR4 (N292, N32, N106, N156, N72);
nand NAND4 (N293, N283, N274, N103, N261);
not NOT1 (N294, N265);
nand NAND2 (N295, N268, N152);
or OR2 (N296, N289, N133);
xor XOR2 (N297, N287, N2);
nor NOR3 (N298, N296, N53, N107);
nand NAND2 (N299, N294, N90);
nor NOR2 (N300, N299, N211);
nor NOR2 (N301, N290, N80);
buf BUF1 (N302, N288);
and AND4 (N303, N298, N286, N61, N187);
xor XOR2 (N304, N301, N123);
nand NAND3 (N305, N297, N110, N115);
not NOT1 (N306, N302);
nor NOR2 (N307, N291, N139);
buf BUF1 (N308, N306);
or OR2 (N309, N308, N226);
buf BUF1 (N310, N307);
buf BUF1 (N311, N305);
nand NAND3 (N312, N311, N165, N12);
nand NAND2 (N313, N304, N184);
not NOT1 (N314, N309);
buf BUF1 (N315, N312);
buf BUF1 (N316, N300);
xor XOR2 (N317, N303, N300);
nor NOR4 (N318, N317, N221, N230, N25);
nor NOR2 (N319, N293, N292);
nor NOR2 (N320, N98, N104);
or OR3 (N321, N314, N308, N130);
or OR4 (N322, N310, N188, N228, N23);
and AND4 (N323, N320, N4, N94, N266);
xor XOR2 (N324, N295, N266);
buf BUF1 (N325, N313);
not NOT1 (N326, N316);
xor XOR2 (N327, N318, N113);
xor XOR2 (N328, N327, N269);
and AND2 (N329, N325, N280);
xor XOR2 (N330, N319, N194);
nor NOR2 (N331, N330, N32);
xor XOR2 (N332, N326, N176);
nor NOR4 (N333, N331, N234, N199, N299);
and AND2 (N334, N328, N98);
nor NOR2 (N335, N321, N42);
nand NAND3 (N336, N315, N44, N183);
buf BUF1 (N337, N332);
and AND3 (N338, N337, N27, N300);
not NOT1 (N339, N324);
not NOT1 (N340, N323);
nor NOR2 (N341, N284, N322);
nand NAND3 (N342, N91, N71, N292);
or OR2 (N343, N333, N149);
or OR3 (N344, N338, N86, N14);
nand NAND2 (N345, N340, N67);
xor XOR2 (N346, N336, N44);
nor NOR3 (N347, N329, N258, N235);
buf BUF1 (N348, N342);
nor NOR3 (N349, N341, N139, N43);
xor XOR2 (N350, N344, N216);
and AND4 (N351, N343, N24, N135, N35);
xor XOR2 (N352, N351, N157);
xor XOR2 (N353, N348, N44);
buf BUF1 (N354, N347);
buf BUF1 (N355, N335);
nand NAND4 (N356, N334, N163, N316, N67);
nand NAND3 (N357, N356, N166, N143);
nor NOR4 (N358, N353, N323, N57, N113);
xor XOR2 (N359, N350, N332);
nor NOR4 (N360, N357, N54, N195, N311);
nand NAND3 (N361, N359, N31, N268);
and AND3 (N362, N349, N11, N65);
not NOT1 (N363, N355);
not NOT1 (N364, N354);
not NOT1 (N365, N363);
buf BUF1 (N366, N364);
nand NAND2 (N367, N352, N34);
or OR4 (N368, N362, N55, N315, N366);
not NOT1 (N369, N42);
nand NAND4 (N370, N369, N168, N285, N43);
not NOT1 (N371, N339);
not NOT1 (N372, N371);
or OR3 (N373, N370, N166, N131);
xor XOR2 (N374, N368, N77);
not NOT1 (N375, N373);
or OR2 (N376, N365, N220);
buf BUF1 (N377, N367);
not NOT1 (N378, N374);
nand NAND2 (N379, N360, N283);
not NOT1 (N380, N377);
buf BUF1 (N381, N376);
xor XOR2 (N382, N345, N336);
and AND3 (N383, N361, N122, N217);
xor XOR2 (N384, N375, N311);
nor NOR2 (N385, N346, N229);
and AND3 (N386, N382, N280, N86);
not NOT1 (N387, N386);
and AND4 (N388, N372, N311, N225, N335);
xor XOR2 (N389, N384, N97);
or OR4 (N390, N380, N319, N120, N239);
not NOT1 (N391, N378);
nor NOR3 (N392, N388, N216, N359);
not NOT1 (N393, N383);
and AND4 (N394, N391, N204, N35, N202);
or OR2 (N395, N387, N52);
not NOT1 (N396, N390);
and AND4 (N397, N358, N318, N101, N373);
or OR3 (N398, N393, N364, N22);
or OR3 (N399, N392, N193, N91);
xor XOR2 (N400, N399, N230);
not NOT1 (N401, N379);
nor NOR2 (N402, N389, N38);
not NOT1 (N403, N400);
buf BUF1 (N404, N395);
not NOT1 (N405, N403);
or OR2 (N406, N398, N116);
or OR2 (N407, N394, N45);
buf BUF1 (N408, N381);
xor XOR2 (N409, N405, N3);
and AND3 (N410, N406, N365, N152);
xor XOR2 (N411, N410, N223);
buf BUF1 (N412, N407);
or OR3 (N413, N396, N355, N138);
or OR2 (N414, N409, N42);
not NOT1 (N415, N404);
buf BUF1 (N416, N402);
and AND3 (N417, N385, N264, N155);
nor NOR3 (N418, N411, N246, N307);
xor XOR2 (N419, N413, N242);
nand NAND4 (N420, N401, N14, N295, N233);
not NOT1 (N421, N420);
or OR4 (N422, N408, N26, N142, N227);
or OR2 (N423, N419, N300);
nor NOR3 (N424, N416, N200, N413);
not NOT1 (N425, N421);
or OR2 (N426, N418, N367);
buf BUF1 (N427, N425);
and AND3 (N428, N415, N228, N132);
buf BUF1 (N429, N428);
buf BUF1 (N430, N429);
and AND2 (N431, N423, N119);
not NOT1 (N432, N412);
and AND2 (N433, N431, N291);
nor NOR2 (N434, N426, N217);
or OR2 (N435, N433, N355);
or OR2 (N436, N424, N92);
or OR3 (N437, N435, N14, N339);
not NOT1 (N438, N427);
or OR3 (N439, N430, N318, N10);
not NOT1 (N440, N397);
and AND2 (N441, N438, N310);
not NOT1 (N442, N440);
nand NAND2 (N443, N437, N120);
nand NAND2 (N444, N436, N383);
nand NAND3 (N445, N442, N273, N24);
xor XOR2 (N446, N432, N50);
nand NAND4 (N447, N443, N429, N111, N325);
not NOT1 (N448, N422);
nor NOR2 (N449, N441, N25);
buf BUF1 (N450, N445);
nand NAND3 (N451, N439, N326, N89);
buf BUF1 (N452, N450);
or OR2 (N453, N434, N47);
or OR2 (N454, N452, N368);
nand NAND3 (N455, N449, N111, N252);
xor XOR2 (N456, N448, N165);
nand NAND2 (N457, N455, N393);
not NOT1 (N458, N453);
not NOT1 (N459, N458);
nor NOR3 (N460, N444, N238, N170);
or OR2 (N461, N414, N438);
not NOT1 (N462, N461);
nand NAND3 (N463, N417, N173, N10);
nand NAND2 (N464, N454, N114);
or OR2 (N465, N456, N273);
and AND3 (N466, N464, N273, N391);
nor NOR3 (N467, N459, N5, N152);
xor XOR2 (N468, N465, N218);
nor NOR2 (N469, N463, N48);
buf BUF1 (N470, N451);
xor XOR2 (N471, N447, N119);
not NOT1 (N472, N466);
nor NOR3 (N473, N467, N169, N101);
nand NAND2 (N474, N473, N61);
buf BUF1 (N475, N470);
not NOT1 (N476, N475);
nand NAND4 (N477, N474, N378, N343, N14);
xor XOR2 (N478, N457, N414);
not NOT1 (N479, N476);
nor NOR2 (N480, N471, N431);
and AND4 (N481, N469, N383, N140, N84);
nand NAND4 (N482, N481, N391, N348, N379);
nor NOR3 (N483, N472, N77, N279);
and AND3 (N484, N477, N75, N129);
not NOT1 (N485, N479);
and AND2 (N486, N482, N258);
xor XOR2 (N487, N484, N326);
not NOT1 (N488, N446);
xor XOR2 (N489, N462, N488);
nor NOR2 (N490, N486, N472);
buf BUF1 (N491, N434);
xor XOR2 (N492, N480, N273);
xor XOR2 (N493, N483, N209);
nor NOR4 (N494, N485, N205, N153, N491);
not NOT1 (N495, N278);
or OR4 (N496, N495, N331, N198, N422);
and AND2 (N497, N487, N319);
and AND2 (N498, N497, N45);
or OR3 (N499, N478, N39, N430);
not NOT1 (N500, N468);
nor NOR4 (N501, N493, N465, N266, N235);
buf BUF1 (N502, N489);
nor NOR4 (N503, N499, N480, N190, N434);
not NOT1 (N504, N496);
or OR4 (N505, N460, N89, N215, N419);
and AND2 (N506, N502, N110);
buf BUF1 (N507, N506);
or OR4 (N508, N490, N309, N127, N219);
nand NAND4 (N509, N498, N22, N159, N283);
and AND2 (N510, N501, N442);
and AND2 (N511, N503, N431);
not NOT1 (N512, N510);
nand NAND3 (N513, N492, N415, N325);
not NOT1 (N514, N494);
nor NOR3 (N515, N507, N97, N9);
not NOT1 (N516, N500);
not NOT1 (N517, N511);
or OR3 (N518, N512, N407, N263);
or OR2 (N519, N515, N102);
and AND4 (N520, N504, N337, N194, N27);
or OR3 (N521, N516, N427, N66);
xor XOR2 (N522, N514, N119);
buf BUF1 (N523, N522);
buf BUF1 (N524, N521);
nor NOR3 (N525, N523, N322, N243);
and AND4 (N526, N517, N173, N110, N81);
or OR2 (N527, N508, N523);
and AND2 (N528, N526, N417);
nor NOR2 (N529, N518, N121);
or OR4 (N530, N529, N76, N429, N327);
buf BUF1 (N531, N519);
nand NAND2 (N532, N525, N248);
and AND2 (N533, N505, N51);
nor NOR3 (N534, N530, N108, N223);
not NOT1 (N535, N513);
not NOT1 (N536, N533);
nand NAND2 (N537, N520, N511);
nand NAND3 (N538, N509, N319, N387);
or OR3 (N539, N537, N303, N1);
xor XOR2 (N540, N536, N262);
nand NAND2 (N541, N534, N537);
nand NAND2 (N542, N531, N209);
or OR2 (N543, N528, N42);
buf BUF1 (N544, N532);
nand NAND2 (N545, N540, N135);
nor NOR2 (N546, N545, N320);
and AND4 (N547, N543, N120, N260, N526);
and AND2 (N548, N544, N118);
xor XOR2 (N549, N524, N525);
nor NOR2 (N550, N527, N428);
not NOT1 (N551, N546);
and AND4 (N552, N551, N270, N89, N439);
nor NOR3 (N553, N538, N548, N450);
and AND4 (N554, N217, N113, N434, N122);
nor NOR2 (N555, N547, N336);
xor XOR2 (N556, N550, N331);
buf BUF1 (N557, N535);
buf BUF1 (N558, N554);
xor XOR2 (N559, N552, N444);
and AND3 (N560, N557, N377, N8);
buf BUF1 (N561, N542);
not NOT1 (N562, N559);
or OR3 (N563, N561, N278, N193);
and AND3 (N564, N555, N386, N277);
buf BUF1 (N565, N564);
nand NAND3 (N566, N556, N182, N541);
nand NAND4 (N567, N315, N141, N516, N486);
nor NOR2 (N568, N549, N192);
not NOT1 (N569, N553);
nand NAND4 (N570, N562, N67, N455, N77);
nand NAND4 (N571, N565, N539, N314, N125);
and AND4 (N572, N250, N484, N220, N75);
nand NAND3 (N573, N571, N193, N71);
nand NAND2 (N574, N568, N465);
or OR4 (N575, N558, N2, N225, N293);
buf BUF1 (N576, N574);
nor NOR3 (N577, N572, N304, N212);
or OR3 (N578, N575, N182, N184);
nand NAND2 (N579, N577, N362);
not NOT1 (N580, N578);
buf BUF1 (N581, N563);
xor XOR2 (N582, N576, N70);
xor XOR2 (N583, N580, N129);
nor NOR2 (N584, N583, N113);
not NOT1 (N585, N570);
and AND2 (N586, N584, N31);
not NOT1 (N587, N560);
nor NOR4 (N588, N581, N570, N232, N575);
nand NAND3 (N589, N587, N138, N511);
and AND4 (N590, N579, N58, N363, N174);
and AND3 (N591, N582, N108, N315);
and AND4 (N592, N588, N558, N144, N171);
xor XOR2 (N593, N589, N67);
xor XOR2 (N594, N590, N29);
or OR4 (N595, N593, N479, N43, N111);
xor XOR2 (N596, N566, N548);
xor XOR2 (N597, N573, N214);
not NOT1 (N598, N594);
or OR2 (N599, N592, N213);
not NOT1 (N600, N567);
buf BUF1 (N601, N596);
not NOT1 (N602, N591);
and AND3 (N603, N585, N438, N197);
xor XOR2 (N604, N600, N554);
xor XOR2 (N605, N604, N501);
and AND2 (N606, N569, N260);
and AND4 (N607, N597, N198, N164, N167);
and AND3 (N608, N599, N418, N389);
nor NOR3 (N609, N603, N521, N169);
not NOT1 (N610, N602);
nand NAND2 (N611, N598, N377);
and AND4 (N612, N609, N246, N554, N404);
or OR3 (N613, N601, N313, N585);
or OR4 (N614, N610, N91, N342, N179);
buf BUF1 (N615, N605);
and AND2 (N616, N611, N419);
nor NOR4 (N617, N614, N450, N334, N336);
or OR3 (N618, N616, N3, N596);
buf BUF1 (N619, N586);
nor NOR4 (N620, N607, N483, N227, N515);
nor NOR4 (N621, N612, N25, N432, N391);
and AND3 (N622, N618, N446, N74);
nand NAND2 (N623, N615, N9);
not NOT1 (N624, N623);
xor XOR2 (N625, N622, N485);
nor NOR4 (N626, N620, N231, N498, N63);
not NOT1 (N627, N613);
not NOT1 (N628, N595);
and AND2 (N629, N608, N193);
nor NOR2 (N630, N624, N106);
nand NAND4 (N631, N626, N111, N115, N244);
or OR4 (N632, N631, N416, N121, N169);
or OR3 (N633, N628, N540, N624);
xor XOR2 (N634, N625, N65);
nor NOR2 (N635, N617, N516);
nand NAND2 (N636, N630, N120);
buf BUF1 (N637, N619);
nand NAND3 (N638, N627, N474, N227);
nand NAND3 (N639, N629, N105, N476);
nor NOR2 (N640, N634, N256);
buf BUF1 (N641, N633);
and AND2 (N642, N621, N635);
and AND3 (N643, N430, N101, N405);
and AND2 (N644, N643, N28);
or OR2 (N645, N638, N140);
nand NAND3 (N646, N645, N17, N86);
nand NAND3 (N647, N646, N247, N410);
xor XOR2 (N648, N636, N627);
buf BUF1 (N649, N648);
or OR2 (N650, N639, N326);
not NOT1 (N651, N637);
not NOT1 (N652, N651);
and AND3 (N653, N652, N82, N590);
xor XOR2 (N654, N641, N456);
and AND4 (N655, N640, N496, N310, N127);
nor NOR4 (N656, N647, N600, N511, N498);
nand NAND4 (N657, N644, N397, N407, N348);
nor NOR3 (N658, N606, N373, N616);
or OR4 (N659, N632, N357, N314, N172);
xor XOR2 (N660, N655, N199);
buf BUF1 (N661, N649);
and AND2 (N662, N656, N298);
xor XOR2 (N663, N660, N326);
nand NAND4 (N664, N661, N176, N254, N40);
nand NAND4 (N665, N650, N62, N149, N577);
buf BUF1 (N666, N663);
nor NOR3 (N667, N642, N201, N605);
and AND2 (N668, N657, N498);
xor XOR2 (N669, N654, N497);
nor NOR3 (N670, N658, N633, N387);
buf BUF1 (N671, N666);
and AND4 (N672, N671, N167, N94, N239);
nand NAND4 (N673, N668, N109, N119, N116);
buf BUF1 (N674, N662);
or OR4 (N675, N673, N76, N161, N493);
or OR2 (N676, N669, N429);
buf BUF1 (N677, N659);
buf BUF1 (N678, N664);
buf BUF1 (N679, N674);
or OR3 (N680, N677, N255, N233);
and AND4 (N681, N675, N215, N369, N562);
or OR2 (N682, N681, N471);
nand NAND2 (N683, N670, N295);
nand NAND4 (N684, N676, N482, N136, N116);
not NOT1 (N685, N680);
and AND4 (N686, N685, N400, N571, N630);
buf BUF1 (N687, N682);
or OR2 (N688, N679, N174);
or OR2 (N689, N653, N376);
buf BUF1 (N690, N684);
not NOT1 (N691, N686);
and AND3 (N692, N691, N14, N354);
not NOT1 (N693, N692);
or OR2 (N694, N667, N544);
or OR3 (N695, N687, N624, N300);
or OR2 (N696, N695, N292);
nand NAND4 (N697, N693, N565, N339, N395);
nor NOR3 (N698, N683, N146, N437);
xor XOR2 (N699, N697, N184);
buf BUF1 (N700, N694);
not NOT1 (N701, N690);
not NOT1 (N702, N672);
not NOT1 (N703, N698);
and AND3 (N704, N699, N335, N78);
xor XOR2 (N705, N665, N539);
and AND2 (N706, N689, N589);
and AND3 (N707, N705, N545, N583);
buf BUF1 (N708, N696);
nand NAND4 (N709, N707, N376, N606, N91);
xor XOR2 (N710, N708, N268);
xor XOR2 (N711, N710, N50);
not NOT1 (N712, N678);
nor NOR3 (N713, N704, N52, N275);
buf BUF1 (N714, N701);
xor XOR2 (N715, N702, N105);
not NOT1 (N716, N715);
xor XOR2 (N717, N709, N294);
nand NAND2 (N718, N712, N242);
not NOT1 (N719, N688);
or OR2 (N720, N717, N527);
buf BUF1 (N721, N719);
nor NOR4 (N722, N718, N358, N669, N139);
not NOT1 (N723, N716);
nor NOR4 (N724, N722, N26, N407, N627);
xor XOR2 (N725, N723, N444);
and AND4 (N726, N720, N480, N582, N695);
xor XOR2 (N727, N703, N97);
nor NOR4 (N728, N726, N644, N132, N439);
nand NAND2 (N729, N727, N204);
and AND4 (N730, N721, N6, N56, N566);
or OR3 (N731, N713, N481, N482);
xor XOR2 (N732, N725, N658);
and AND4 (N733, N728, N21, N213, N401);
nand NAND4 (N734, N730, N499, N346, N58);
not NOT1 (N735, N706);
not NOT1 (N736, N735);
nor NOR3 (N737, N714, N513, N107);
xor XOR2 (N738, N731, N501);
not NOT1 (N739, N734);
or OR4 (N740, N700, N103, N492, N100);
and AND3 (N741, N736, N363, N320);
xor XOR2 (N742, N724, N222);
and AND3 (N743, N729, N614, N566);
or OR4 (N744, N733, N685, N623, N246);
buf BUF1 (N745, N743);
nand NAND2 (N746, N741, N241);
and AND3 (N747, N737, N69, N474);
or OR3 (N748, N742, N51, N195);
nor NOR3 (N749, N739, N107, N457);
nor NOR2 (N750, N748, N8);
buf BUF1 (N751, N747);
xor XOR2 (N752, N744, N290);
buf BUF1 (N753, N746);
or OR3 (N754, N749, N207, N447);
and AND3 (N755, N751, N365, N462);
or OR3 (N756, N754, N307, N339);
and AND4 (N757, N711, N187, N578, N613);
not NOT1 (N758, N745);
not NOT1 (N759, N758);
buf BUF1 (N760, N756);
or OR3 (N761, N750, N743, N339);
nand NAND4 (N762, N755, N409, N222, N30);
nor NOR2 (N763, N760, N32);
xor XOR2 (N764, N753, N45);
not NOT1 (N765, N740);
and AND4 (N766, N761, N548, N301, N353);
and AND4 (N767, N738, N623, N298, N30);
xor XOR2 (N768, N764, N215);
nand NAND3 (N769, N763, N485, N341);
xor XOR2 (N770, N765, N627);
not NOT1 (N771, N768);
buf BUF1 (N772, N762);
xor XOR2 (N773, N759, N50);
and AND4 (N774, N752, N164, N421, N221);
and AND2 (N775, N732, N671);
nand NAND2 (N776, N775, N314);
nor NOR4 (N777, N757, N682, N373, N618);
nor NOR4 (N778, N769, N71, N240, N339);
or OR3 (N779, N766, N96, N583);
not NOT1 (N780, N770);
xor XOR2 (N781, N777, N666);
xor XOR2 (N782, N778, N302);
nand NAND4 (N783, N771, N519, N651, N429);
not NOT1 (N784, N780);
xor XOR2 (N785, N781, N575);
nand NAND2 (N786, N779, N415);
xor XOR2 (N787, N783, N409);
nand NAND2 (N788, N772, N229);
xor XOR2 (N789, N784, N612);
buf BUF1 (N790, N786);
buf BUF1 (N791, N782);
or OR3 (N792, N788, N314, N686);
nand NAND4 (N793, N792, N358, N364, N657);
nor NOR2 (N794, N791, N364);
nor NOR4 (N795, N793, N543, N628, N8);
or OR3 (N796, N789, N473, N82);
not NOT1 (N797, N776);
nor NOR3 (N798, N785, N166, N219);
nor NOR3 (N799, N790, N329, N427);
not NOT1 (N800, N787);
and AND4 (N801, N797, N640, N486, N474);
and AND4 (N802, N800, N121, N547, N649);
nor NOR3 (N803, N795, N343, N579);
buf BUF1 (N804, N799);
nor NOR2 (N805, N767, N488);
xor XOR2 (N806, N802, N308);
and AND4 (N807, N801, N610, N87, N757);
buf BUF1 (N808, N806);
not NOT1 (N809, N774);
and AND2 (N810, N773, N650);
nand NAND3 (N811, N796, N386, N742);
xor XOR2 (N812, N794, N772);
xor XOR2 (N813, N811, N191);
nand NAND3 (N814, N805, N803, N632);
and AND2 (N815, N458, N765);
xor XOR2 (N816, N812, N491);
or OR3 (N817, N798, N94, N685);
not NOT1 (N818, N804);
not NOT1 (N819, N808);
xor XOR2 (N820, N815, N206);
buf BUF1 (N821, N818);
not NOT1 (N822, N810);
nor NOR4 (N823, N809, N269, N612, N611);
and AND3 (N824, N821, N180, N676);
not NOT1 (N825, N814);
xor XOR2 (N826, N820, N33);
or OR2 (N827, N822, N480);
nand NAND2 (N828, N824, N430);
not NOT1 (N829, N828);
not NOT1 (N830, N825);
and AND4 (N831, N816, N220, N513, N102);
nor NOR3 (N832, N813, N117, N729);
xor XOR2 (N833, N827, N695);
and AND2 (N834, N833, N677);
not NOT1 (N835, N817);
nand NAND3 (N836, N834, N361, N171);
not NOT1 (N837, N835);
and AND3 (N838, N829, N340, N629);
nor NOR3 (N839, N830, N814, N230);
buf BUF1 (N840, N807);
buf BUF1 (N841, N840);
not NOT1 (N842, N841);
nand NAND4 (N843, N838, N110, N336, N606);
or OR3 (N844, N819, N601, N355);
buf BUF1 (N845, N837);
xor XOR2 (N846, N836, N384);
or OR2 (N847, N842, N370);
buf BUF1 (N848, N823);
nor NOR4 (N849, N843, N61, N615, N806);
and AND3 (N850, N849, N405, N277);
and AND2 (N851, N847, N570);
xor XOR2 (N852, N839, N90);
not NOT1 (N853, N846);
nor NOR4 (N854, N845, N461, N359, N134);
and AND3 (N855, N844, N562, N679);
nor NOR3 (N856, N855, N644, N339);
and AND2 (N857, N850, N381);
or OR3 (N858, N857, N653, N210);
or OR2 (N859, N854, N189);
or OR2 (N860, N826, N267);
buf BUF1 (N861, N848);
or OR4 (N862, N831, N557, N679, N284);
not NOT1 (N863, N862);
and AND2 (N864, N856, N138);
or OR4 (N865, N832, N564, N707, N406);
buf BUF1 (N866, N858);
nand NAND3 (N867, N853, N208, N274);
nand NAND2 (N868, N852, N3);
not NOT1 (N869, N860);
buf BUF1 (N870, N867);
not NOT1 (N871, N869);
nand NAND3 (N872, N870, N404, N819);
not NOT1 (N873, N859);
buf BUF1 (N874, N864);
nand NAND2 (N875, N866, N268);
nor NOR4 (N876, N863, N600, N547, N537);
not NOT1 (N877, N874);
buf BUF1 (N878, N861);
not NOT1 (N879, N876);
nand NAND2 (N880, N873, N289);
xor XOR2 (N881, N871, N640);
not NOT1 (N882, N875);
nand NAND3 (N883, N877, N111, N214);
buf BUF1 (N884, N880);
xor XOR2 (N885, N884, N256);
and AND3 (N886, N883, N544, N246);
buf BUF1 (N887, N881);
nand NAND3 (N888, N851, N449, N676);
buf BUF1 (N889, N868);
nand NAND3 (N890, N888, N56, N338);
xor XOR2 (N891, N878, N796);
and AND3 (N892, N872, N634, N684);
nor NOR2 (N893, N879, N425);
buf BUF1 (N894, N885);
nor NOR2 (N895, N865, N252);
or OR3 (N896, N894, N228, N641);
and AND2 (N897, N889, N143);
buf BUF1 (N898, N890);
and AND3 (N899, N886, N74, N478);
buf BUF1 (N900, N895);
xor XOR2 (N901, N896, N287);
and AND4 (N902, N899, N424, N858, N469);
not NOT1 (N903, N901);
xor XOR2 (N904, N902, N350);
xor XOR2 (N905, N898, N197);
nor NOR4 (N906, N882, N681, N468, N856);
nand NAND3 (N907, N891, N134, N799);
not NOT1 (N908, N906);
nand NAND3 (N909, N897, N95, N694);
xor XOR2 (N910, N903, N739);
xor XOR2 (N911, N887, N583);
nand NAND2 (N912, N910, N238);
and AND2 (N913, N907, N772);
xor XOR2 (N914, N900, N227);
or OR4 (N915, N909, N462, N125, N695);
nand NAND2 (N916, N911, N803);
not NOT1 (N917, N916);
or OR2 (N918, N905, N662);
xor XOR2 (N919, N893, N737);
nor NOR2 (N920, N919, N811);
or OR2 (N921, N908, N282);
nor NOR4 (N922, N915, N759, N688, N300);
not NOT1 (N923, N914);
nand NAND3 (N924, N921, N899, N830);
nor NOR4 (N925, N913, N327, N92, N556);
not NOT1 (N926, N922);
or OR4 (N927, N920, N632, N510, N284);
nand NAND4 (N928, N917, N480, N86, N279);
not NOT1 (N929, N904);
buf BUF1 (N930, N924);
not NOT1 (N931, N912);
nor NOR3 (N932, N928, N681, N554);
buf BUF1 (N933, N931);
buf BUF1 (N934, N918);
xor XOR2 (N935, N892, N92);
nand NAND2 (N936, N935, N241);
nand NAND4 (N937, N936, N191, N688, N203);
xor XOR2 (N938, N925, N497);
and AND2 (N939, N929, N760);
or OR2 (N940, N932, N167);
nand NAND4 (N941, N930, N900, N502, N13);
xor XOR2 (N942, N926, N34);
not NOT1 (N943, N941);
xor XOR2 (N944, N934, N98);
or OR2 (N945, N923, N168);
buf BUF1 (N946, N943);
xor XOR2 (N947, N927, N477);
not NOT1 (N948, N947);
nor NOR4 (N949, N933, N28, N713, N25);
and AND3 (N950, N945, N103, N333);
nor NOR3 (N951, N946, N661, N110);
nand NAND4 (N952, N938, N457, N692, N563);
or OR2 (N953, N940, N482);
or OR4 (N954, N944, N620, N456, N942);
or OR2 (N955, N524, N898);
and AND3 (N956, N937, N647, N234);
nor NOR4 (N957, N949, N421, N934, N557);
not NOT1 (N958, N955);
xor XOR2 (N959, N957, N590);
or OR2 (N960, N958, N426);
nor NOR4 (N961, N939, N762, N316, N345);
buf BUF1 (N962, N954);
or OR4 (N963, N952, N556, N174, N358);
or OR2 (N964, N953, N505);
and AND3 (N965, N963, N386, N80);
nand NAND4 (N966, N951, N505, N947, N248);
nor NOR2 (N967, N959, N731);
not NOT1 (N968, N960);
nor NOR2 (N969, N962, N931);
nor NOR3 (N970, N964, N252, N621);
nor NOR4 (N971, N968, N335, N285, N368);
nor NOR4 (N972, N948, N648, N23, N29);
xor XOR2 (N973, N971, N820);
not NOT1 (N974, N966);
nand NAND4 (N975, N972, N574, N506, N48);
nand NAND2 (N976, N969, N159);
buf BUF1 (N977, N976);
or OR2 (N978, N974, N961);
or OR4 (N979, N304, N629, N296, N745);
and AND3 (N980, N967, N293, N599);
xor XOR2 (N981, N978, N970);
xor XOR2 (N982, N682, N837);
xor XOR2 (N983, N950, N567);
not NOT1 (N984, N982);
nand NAND3 (N985, N973, N626, N547);
and AND2 (N986, N984, N423);
or OR4 (N987, N985, N19, N962, N960);
or OR2 (N988, N983, N938);
nand NAND2 (N989, N977, N553);
nand NAND4 (N990, N965, N944, N237, N36);
nand NAND3 (N991, N956, N499, N171);
nor NOR2 (N992, N975, N688);
buf BUF1 (N993, N991);
xor XOR2 (N994, N980, N252);
buf BUF1 (N995, N987);
or OR4 (N996, N992, N932, N750, N672);
buf BUF1 (N997, N989);
and AND2 (N998, N993, N405);
xor XOR2 (N999, N997, N651);
nand NAND3 (N1000, N986, N496, N531);
and AND4 (N1001, N990, N421, N355, N104);
or OR2 (N1002, N999, N329);
buf BUF1 (N1003, N994);
buf BUF1 (N1004, N981);
buf BUF1 (N1005, N1002);
or OR3 (N1006, N995, N412, N46);
not NOT1 (N1007, N1001);
xor XOR2 (N1008, N996, N574);
not NOT1 (N1009, N1007);
or OR2 (N1010, N979, N361);
or OR4 (N1011, N1010, N122, N596, N388);
nor NOR2 (N1012, N998, N858);
xor XOR2 (N1013, N1000, N128);
xor XOR2 (N1014, N1009, N811);
or OR3 (N1015, N1006, N367, N742);
buf BUF1 (N1016, N1003);
or OR3 (N1017, N1004, N68, N806);
and AND2 (N1018, N1012, N963);
xor XOR2 (N1019, N1015, N483);
xor XOR2 (N1020, N1013, N1018);
nor NOR2 (N1021, N283, N418);
nor NOR4 (N1022, N1020, N155, N673, N117);
or OR2 (N1023, N1021, N589);
nand NAND2 (N1024, N1016, N11);
xor XOR2 (N1025, N1011, N571);
nor NOR4 (N1026, N1008, N576, N968, N662);
not NOT1 (N1027, N1026);
not NOT1 (N1028, N1005);
and AND4 (N1029, N1025, N467, N39, N691);
or OR3 (N1030, N1029, N129, N563);
xor XOR2 (N1031, N1028, N966);
nor NOR2 (N1032, N1022, N517);
buf BUF1 (N1033, N1017);
and AND4 (N1034, N1023, N984, N369, N406);
not NOT1 (N1035, N1014);
xor XOR2 (N1036, N1019, N977);
buf BUF1 (N1037, N1031);
buf BUF1 (N1038, N1035);
and AND2 (N1039, N1036, N917);
nand NAND3 (N1040, N1032, N380, N312);
nand NAND3 (N1041, N1040, N55, N457);
and AND4 (N1042, N988, N159, N897, N350);
buf BUF1 (N1043, N1027);
nor NOR4 (N1044, N1041, N362, N767, N983);
not NOT1 (N1045, N1030);
and AND4 (N1046, N1042, N23, N729, N519);
nor NOR4 (N1047, N1046, N63, N258, N127);
xor XOR2 (N1048, N1043, N198);
or OR2 (N1049, N1048, N112);
xor XOR2 (N1050, N1047, N741);
xor XOR2 (N1051, N1034, N152);
nand NAND2 (N1052, N1050, N648);
or OR3 (N1053, N1051, N254, N885);
and AND3 (N1054, N1038, N615, N226);
or OR2 (N1055, N1039, N364);
nand NAND3 (N1056, N1054, N200, N521);
or OR4 (N1057, N1053, N271, N625, N1035);
nand NAND3 (N1058, N1055, N951, N342);
not NOT1 (N1059, N1045);
nor NOR4 (N1060, N1058, N279, N624, N919);
nand NAND3 (N1061, N1024, N442, N955);
nand NAND4 (N1062, N1044, N589, N774, N517);
nand NAND3 (N1063, N1060, N247, N330);
nand NAND4 (N1064, N1049, N701, N302, N654);
nor NOR3 (N1065, N1063, N851, N322);
or OR3 (N1066, N1062, N669, N141);
not NOT1 (N1067, N1065);
nor NOR3 (N1068, N1037, N364, N554);
xor XOR2 (N1069, N1057, N570);
nor NOR4 (N1070, N1069, N895, N715, N736);
nor NOR2 (N1071, N1064, N203);
xor XOR2 (N1072, N1068, N266);
xor XOR2 (N1073, N1067, N355);
or OR4 (N1074, N1033, N655, N302, N886);
xor XOR2 (N1075, N1052, N282);
and AND2 (N1076, N1056, N802);
not NOT1 (N1077, N1059);
buf BUF1 (N1078, N1076);
nand NAND4 (N1079, N1070, N687, N335, N852);
buf BUF1 (N1080, N1074);
nor NOR2 (N1081, N1078, N917);
or OR3 (N1082, N1075, N953, N318);
not NOT1 (N1083, N1079);
xor XOR2 (N1084, N1082, N1081);
nor NOR4 (N1085, N909, N224, N972, N543);
nor NOR4 (N1086, N1077, N318, N401, N890);
nor NOR3 (N1087, N1085, N302, N55);
or OR3 (N1088, N1071, N916, N1037);
or OR3 (N1089, N1088, N5, N56);
buf BUF1 (N1090, N1061);
not NOT1 (N1091, N1083);
not NOT1 (N1092, N1084);
nand NAND2 (N1093, N1066, N472);
xor XOR2 (N1094, N1092, N144);
or OR2 (N1095, N1089, N924);
xor XOR2 (N1096, N1094, N508);
and AND4 (N1097, N1090, N681, N889, N860);
or OR3 (N1098, N1091, N379, N915);
or OR2 (N1099, N1072, N599);
not NOT1 (N1100, N1093);
nand NAND2 (N1101, N1080, N1085);
xor XOR2 (N1102, N1100, N397);
nand NAND4 (N1103, N1098, N949, N415, N742);
xor XOR2 (N1104, N1102, N960);
nor NOR4 (N1105, N1099, N60, N655, N389);
or OR2 (N1106, N1104, N20);
and AND2 (N1107, N1095, N454);
xor XOR2 (N1108, N1103, N53);
xor XOR2 (N1109, N1108, N471);
xor XOR2 (N1110, N1107, N62);
not NOT1 (N1111, N1110);
and AND2 (N1112, N1087, N804);
nand NAND2 (N1113, N1073, N721);
and AND4 (N1114, N1097, N470, N705, N529);
nand NAND4 (N1115, N1105, N849, N390, N234);
nand NAND2 (N1116, N1112, N446);
or OR2 (N1117, N1086, N1044);
and AND3 (N1118, N1109, N730, N620);
xor XOR2 (N1119, N1096, N1052);
xor XOR2 (N1120, N1119, N1096);
and AND3 (N1121, N1111, N875, N321);
xor XOR2 (N1122, N1121, N881);
or OR4 (N1123, N1101, N582, N589, N772);
xor XOR2 (N1124, N1115, N681);
or OR3 (N1125, N1122, N900, N927);
or OR2 (N1126, N1116, N659);
or OR3 (N1127, N1106, N267, N231);
not NOT1 (N1128, N1127);
nand NAND2 (N1129, N1120, N734);
nand NAND4 (N1130, N1125, N374, N459, N71);
nand NAND2 (N1131, N1126, N455);
not NOT1 (N1132, N1129);
nand NAND3 (N1133, N1131, N264, N999);
nor NOR3 (N1134, N1113, N511, N951);
xor XOR2 (N1135, N1123, N99);
buf BUF1 (N1136, N1128);
buf BUF1 (N1137, N1124);
buf BUF1 (N1138, N1137);
not NOT1 (N1139, N1114);
nor NOR4 (N1140, N1132, N318, N827, N57);
buf BUF1 (N1141, N1140);
nor NOR4 (N1142, N1133, N480, N792, N316);
nor NOR2 (N1143, N1118, N1142);
nor NOR2 (N1144, N23, N377);
not NOT1 (N1145, N1144);
and AND4 (N1146, N1139, N31, N21, N623);
and AND3 (N1147, N1146, N322, N1090);
buf BUF1 (N1148, N1130);
or OR3 (N1149, N1134, N116, N315);
buf BUF1 (N1150, N1117);
not NOT1 (N1151, N1141);
xor XOR2 (N1152, N1147, N348);
xor XOR2 (N1153, N1151, N361);
nand NAND2 (N1154, N1152, N922);
nand NAND2 (N1155, N1136, N108);
nand NAND4 (N1156, N1138, N501, N459, N406);
xor XOR2 (N1157, N1153, N253);
not NOT1 (N1158, N1148);
nand NAND2 (N1159, N1158, N472);
xor XOR2 (N1160, N1143, N993);
nand NAND4 (N1161, N1135, N251, N1027, N647);
nor NOR3 (N1162, N1145, N361, N583);
not NOT1 (N1163, N1156);
or OR2 (N1164, N1155, N87);
buf BUF1 (N1165, N1150);
buf BUF1 (N1166, N1164);
and AND2 (N1167, N1159, N461);
or OR2 (N1168, N1160, N763);
not NOT1 (N1169, N1165);
xor XOR2 (N1170, N1162, N197);
nor NOR2 (N1171, N1163, N631);
xor XOR2 (N1172, N1168, N281);
buf BUF1 (N1173, N1154);
buf BUF1 (N1174, N1173);
xor XOR2 (N1175, N1161, N311);
xor XOR2 (N1176, N1157, N559);
nand NAND4 (N1177, N1172, N162, N1044, N158);
nand NAND2 (N1178, N1167, N747);
buf BUF1 (N1179, N1170);
xor XOR2 (N1180, N1149, N1178);
xor XOR2 (N1181, N94, N248);
not NOT1 (N1182, N1171);
xor XOR2 (N1183, N1179, N426);
buf BUF1 (N1184, N1177);
buf BUF1 (N1185, N1182);
buf BUF1 (N1186, N1176);
nand NAND4 (N1187, N1184, N112, N436, N541);
nand NAND4 (N1188, N1185, N1012, N226, N903);
or OR4 (N1189, N1166, N1051, N791, N428);
not NOT1 (N1190, N1181);
not NOT1 (N1191, N1174);
nand NAND4 (N1192, N1190, N129, N581, N678);
not NOT1 (N1193, N1169);
xor XOR2 (N1194, N1191, N552);
nor NOR3 (N1195, N1186, N1187, N1027);
nor NOR4 (N1196, N865, N797, N76, N649);
buf BUF1 (N1197, N1196);
or OR2 (N1198, N1188, N122);
xor XOR2 (N1199, N1180, N105);
buf BUF1 (N1200, N1175);
nand NAND4 (N1201, N1192, N37, N250, N1063);
and AND2 (N1202, N1193, N57);
nor NOR4 (N1203, N1200, N776, N903, N1007);
buf BUF1 (N1204, N1197);
and AND2 (N1205, N1201, N989);
buf BUF1 (N1206, N1198);
buf BUF1 (N1207, N1189);
not NOT1 (N1208, N1205);
xor XOR2 (N1209, N1183, N507);
buf BUF1 (N1210, N1207);
nor NOR4 (N1211, N1204, N134, N1161, N679);
or OR4 (N1212, N1203, N1126, N897, N966);
nand NAND3 (N1213, N1194, N796, N341);
buf BUF1 (N1214, N1208);
or OR2 (N1215, N1202, N339);
not NOT1 (N1216, N1215);
nand NAND2 (N1217, N1212, N196);
nand NAND3 (N1218, N1216, N840, N1020);
and AND2 (N1219, N1218, N576);
or OR3 (N1220, N1206, N132, N228);
and AND4 (N1221, N1220, N768, N806, N238);
xor XOR2 (N1222, N1217, N646);
or OR2 (N1223, N1210, N44);
xor XOR2 (N1224, N1195, N398);
or OR4 (N1225, N1223, N531, N1063, N569);
not NOT1 (N1226, N1224);
buf BUF1 (N1227, N1209);
and AND4 (N1228, N1213, N752, N599, N833);
nand NAND2 (N1229, N1222, N89);
xor XOR2 (N1230, N1225, N541);
not NOT1 (N1231, N1214);
xor XOR2 (N1232, N1231, N28);
nor NOR2 (N1233, N1221, N940);
nand NAND4 (N1234, N1230, N13, N1157, N176);
not NOT1 (N1235, N1226);
nand NAND2 (N1236, N1228, N288);
or OR4 (N1237, N1232, N506, N369, N136);
xor XOR2 (N1238, N1236, N184);
and AND3 (N1239, N1219, N1126, N256);
and AND4 (N1240, N1235, N919, N805, N827);
nand NAND4 (N1241, N1237, N1128, N733, N34);
not NOT1 (N1242, N1211);
or OR4 (N1243, N1241, N939, N286, N997);
or OR4 (N1244, N1240, N1011, N698, N134);
and AND4 (N1245, N1242, N272, N418, N962);
buf BUF1 (N1246, N1227);
nand NAND3 (N1247, N1243, N922, N640);
nand NAND2 (N1248, N1233, N233);
and AND2 (N1249, N1244, N1189);
not NOT1 (N1250, N1246);
and AND4 (N1251, N1248, N745, N85, N414);
xor XOR2 (N1252, N1229, N241);
or OR2 (N1253, N1250, N826);
and AND2 (N1254, N1245, N1242);
not NOT1 (N1255, N1247);
nand NAND2 (N1256, N1239, N629);
or OR3 (N1257, N1249, N404, N194);
and AND4 (N1258, N1238, N868, N1055, N1012);
buf BUF1 (N1259, N1255);
not NOT1 (N1260, N1257);
and AND2 (N1261, N1254, N84);
and AND4 (N1262, N1251, N764, N443, N832);
not NOT1 (N1263, N1262);
not NOT1 (N1264, N1260);
nor NOR2 (N1265, N1256, N219);
nand NAND2 (N1266, N1265, N419);
buf BUF1 (N1267, N1258);
nor NOR2 (N1268, N1234, N820);
buf BUF1 (N1269, N1268);
or OR3 (N1270, N1199, N1156, N284);
or OR2 (N1271, N1269, N1059);
not NOT1 (N1272, N1266);
buf BUF1 (N1273, N1267);
xor XOR2 (N1274, N1270, N716);
xor XOR2 (N1275, N1263, N990);
and AND4 (N1276, N1273, N527, N1215, N189);
nor NOR3 (N1277, N1252, N878, N1074);
and AND2 (N1278, N1261, N215);
and AND2 (N1279, N1259, N688);
buf BUF1 (N1280, N1271);
xor XOR2 (N1281, N1264, N1232);
or OR3 (N1282, N1280, N835, N811);
not NOT1 (N1283, N1275);
or OR3 (N1284, N1279, N108, N92);
buf BUF1 (N1285, N1277);
nor NOR3 (N1286, N1272, N1119, N1059);
nor NOR3 (N1287, N1281, N831, N143);
nor NOR3 (N1288, N1276, N993, N680);
not NOT1 (N1289, N1253);
buf BUF1 (N1290, N1283);
and AND4 (N1291, N1282, N525, N637, N1184);
or OR4 (N1292, N1286, N1249, N226, N219);
or OR4 (N1293, N1292, N719, N219, N168);
or OR2 (N1294, N1293, N1111);
or OR3 (N1295, N1278, N602, N531);
xor XOR2 (N1296, N1274, N625);
nor NOR3 (N1297, N1290, N372, N1120);
xor XOR2 (N1298, N1291, N1282);
and AND2 (N1299, N1289, N740);
nand NAND4 (N1300, N1298, N1258, N1283, N62);
not NOT1 (N1301, N1285);
and AND2 (N1302, N1296, N739);
or OR2 (N1303, N1302, N312);
nor NOR4 (N1304, N1288, N617, N44, N636);
or OR3 (N1305, N1284, N924, N128);
xor XOR2 (N1306, N1305, N635);
nor NOR2 (N1307, N1303, N262);
buf BUF1 (N1308, N1307);
not NOT1 (N1309, N1299);
xor XOR2 (N1310, N1300, N146);
not NOT1 (N1311, N1287);
not NOT1 (N1312, N1306);
nor NOR3 (N1313, N1308, N185, N310);
nand NAND3 (N1314, N1295, N318, N168);
not NOT1 (N1315, N1309);
nor NOR4 (N1316, N1312, N832, N1276, N63);
xor XOR2 (N1317, N1311, N670);
nand NAND4 (N1318, N1316, N239, N282, N331);
xor XOR2 (N1319, N1318, N592);
not NOT1 (N1320, N1319);
or OR2 (N1321, N1304, N266);
nand NAND3 (N1322, N1315, N645, N956);
or OR3 (N1323, N1310, N465, N418);
nor NOR2 (N1324, N1322, N942);
nor NOR4 (N1325, N1301, N131, N360, N456);
nor NOR4 (N1326, N1313, N489, N1168, N991);
buf BUF1 (N1327, N1297);
nand NAND4 (N1328, N1323, N939, N252, N876);
nor NOR3 (N1329, N1294, N711, N209);
or OR2 (N1330, N1317, N914);
and AND2 (N1331, N1320, N928);
xor XOR2 (N1332, N1321, N945);
nor NOR2 (N1333, N1328, N658);
buf BUF1 (N1334, N1326);
not NOT1 (N1335, N1332);
xor XOR2 (N1336, N1314, N1303);
xor XOR2 (N1337, N1330, N1315);
and AND4 (N1338, N1331, N1258, N222, N315);
xor XOR2 (N1339, N1334, N949);
nand NAND3 (N1340, N1337, N1159, N1294);
not NOT1 (N1341, N1333);
xor XOR2 (N1342, N1329, N1119);
and AND3 (N1343, N1335, N297, N857);
xor XOR2 (N1344, N1343, N1218);
nor NOR3 (N1345, N1338, N363, N1069);
or OR3 (N1346, N1341, N928, N221);
nand NAND2 (N1347, N1327, N1064);
or OR2 (N1348, N1340, N1068);
nand NAND3 (N1349, N1347, N970, N814);
buf BUF1 (N1350, N1342);
not NOT1 (N1351, N1348);
nand NAND4 (N1352, N1351, N1119, N519, N906);
or OR4 (N1353, N1339, N1197, N546, N1054);
and AND3 (N1354, N1344, N313, N247);
or OR3 (N1355, N1349, N1077, N112);
nor NOR4 (N1356, N1325, N89, N1186, N156);
nor NOR2 (N1357, N1352, N782);
nor NOR2 (N1358, N1353, N436);
and AND4 (N1359, N1324, N160, N360, N229);
nor NOR4 (N1360, N1350, N511, N1023, N1011);
nor NOR3 (N1361, N1360, N59, N1265);
and AND3 (N1362, N1359, N2, N1299);
not NOT1 (N1363, N1354);
buf BUF1 (N1364, N1355);
nor NOR2 (N1365, N1357, N587);
or OR3 (N1366, N1346, N185, N1188);
xor XOR2 (N1367, N1361, N18);
not NOT1 (N1368, N1362);
and AND2 (N1369, N1363, N1167);
xor XOR2 (N1370, N1358, N980);
nand NAND4 (N1371, N1367, N1292, N587, N910);
buf BUF1 (N1372, N1356);
not NOT1 (N1373, N1365);
and AND3 (N1374, N1373, N1161, N1038);
or OR2 (N1375, N1368, N1062);
nor NOR2 (N1376, N1345, N1332);
not NOT1 (N1377, N1366);
nor NOR3 (N1378, N1374, N637, N874);
or OR3 (N1379, N1371, N1324, N429);
or OR4 (N1380, N1369, N524, N190, N32);
or OR3 (N1381, N1380, N887, N97);
not NOT1 (N1382, N1377);
and AND4 (N1383, N1370, N463, N741, N1373);
nor NOR2 (N1384, N1381, N278);
xor XOR2 (N1385, N1378, N653);
or OR3 (N1386, N1385, N568, N72);
or OR3 (N1387, N1376, N916, N1335);
buf BUF1 (N1388, N1383);
buf BUF1 (N1389, N1387);
buf BUF1 (N1390, N1386);
nor NOR2 (N1391, N1336, N1063);
not NOT1 (N1392, N1391);
and AND4 (N1393, N1372, N953, N136, N432);
not NOT1 (N1394, N1364);
and AND2 (N1395, N1384, N289);
xor XOR2 (N1396, N1375, N1215);
xor XOR2 (N1397, N1393, N1176);
not NOT1 (N1398, N1394);
buf BUF1 (N1399, N1395);
or OR3 (N1400, N1389, N837, N998);
and AND3 (N1401, N1379, N1393, N1039);
or OR3 (N1402, N1399, N335, N1310);
nor NOR4 (N1403, N1401, N166, N695, N367);
nand NAND3 (N1404, N1396, N24, N1145);
and AND2 (N1405, N1398, N1271);
or OR4 (N1406, N1382, N1113, N646, N1236);
not NOT1 (N1407, N1403);
xor XOR2 (N1408, N1407, N1303);
nand NAND4 (N1409, N1402, N1054, N1174, N471);
xor XOR2 (N1410, N1390, N400);
buf BUF1 (N1411, N1392);
not NOT1 (N1412, N1408);
buf BUF1 (N1413, N1406);
xor XOR2 (N1414, N1413, N411);
or OR3 (N1415, N1412, N1310, N770);
buf BUF1 (N1416, N1397);
nand NAND3 (N1417, N1414, N760, N676);
nor NOR3 (N1418, N1405, N469, N280);
and AND3 (N1419, N1417, N1364, N1190);
buf BUF1 (N1420, N1416);
nand NAND4 (N1421, N1420, N203, N725, N1214);
not NOT1 (N1422, N1415);
nand NAND3 (N1423, N1411, N1411, N113);
and AND3 (N1424, N1421, N54, N1153);
and AND3 (N1425, N1404, N162, N792);
xor XOR2 (N1426, N1419, N721);
nand NAND3 (N1427, N1410, N110, N293);
xor XOR2 (N1428, N1425, N511);
nand NAND2 (N1429, N1427, N28);
nor NOR2 (N1430, N1429, N1049);
and AND2 (N1431, N1423, N364);
nand NAND2 (N1432, N1426, N80);
nor NOR3 (N1433, N1388, N594, N266);
not NOT1 (N1434, N1418);
nor NOR3 (N1435, N1400, N75, N1403);
not NOT1 (N1436, N1422);
buf BUF1 (N1437, N1424);
and AND4 (N1438, N1432, N205, N657, N858);
or OR3 (N1439, N1409, N214, N150);
and AND3 (N1440, N1433, N244, N932);
nor NOR4 (N1441, N1435, N651, N1243, N389);
or OR2 (N1442, N1434, N1055);
not NOT1 (N1443, N1439);
buf BUF1 (N1444, N1441);
nor NOR2 (N1445, N1438, N1071);
not NOT1 (N1446, N1431);
or OR2 (N1447, N1428, N899);
or OR4 (N1448, N1437, N348, N1436, N1361);
or OR2 (N1449, N469, N140);
and AND2 (N1450, N1449, N75);
nor NOR2 (N1451, N1440, N102);
not NOT1 (N1452, N1447);
or OR4 (N1453, N1444, N89, N343, N1207);
xor XOR2 (N1454, N1451, N863);
or OR3 (N1455, N1448, N802, N711);
not NOT1 (N1456, N1445);
nand NAND3 (N1457, N1430, N469, N893);
or OR2 (N1458, N1454, N489);
nor NOR3 (N1459, N1458, N407, N128);
and AND4 (N1460, N1446, N326, N1230, N1459);
or OR3 (N1461, N378, N661, N911);
nand NAND2 (N1462, N1461, N564);
buf BUF1 (N1463, N1457);
or OR4 (N1464, N1460, N690, N778, N1111);
not NOT1 (N1465, N1453);
nor NOR4 (N1466, N1450, N743, N1396, N663);
not NOT1 (N1467, N1452);
buf BUF1 (N1468, N1464);
not NOT1 (N1469, N1442);
and AND4 (N1470, N1468, N1000, N138, N1267);
and AND3 (N1471, N1465, N1051, N1273);
and AND2 (N1472, N1463, N909);
xor XOR2 (N1473, N1466, N1399);
buf BUF1 (N1474, N1471);
nand NAND4 (N1475, N1455, N72, N336, N1173);
xor XOR2 (N1476, N1443, N1242);
not NOT1 (N1477, N1476);
xor XOR2 (N1478, N1477, N682);
nand NAND3 (N1479, N1474, N453, N1393);
buf BUF1 (N1480, N1470);
nor NOR4 (N1481, N1469, N1458, N73, N863);
not NOT1 (N1482, N1481);
buf BUF1 (N1483, N1478);
or OR3 (N1484, N1472, N1482, N1111);
nand NAND4 (N1485, N991, N582, N295, N1038);
nand NAND4 (N1486, N1483, N267, N1419, N199);
xor XOR2 (N1487, N1480, N350);
and AND4 (N1488, N1485, N100, N1101, N833);
buf BUF1 (N1489, N1486);
and AND4 (N1490, N1487, N1257, N1036, N990);
not NOT1 (N1491, N1467);
xor XOR2 (N1492, N1479, N528);
not NOT1 (N1493, N1488);
not NOT1 (N1494, N1484);
nand NAND4 (N1495, N1456, N506, N384, N1311);
buf BUF1 (N1496, N1495);
nand NAND3 (N1497, N1473, N561, N374);
buf BUF1 (N1498, N1475);
buf BUF1 (N1499, N1496);
not NOT1 (N1500, N1498);
nand NAND2 (N1501, N1500, N870);
xor XOR2 (N1502, N1489, N1334);
nor NOR3 (N1503, N1490, N277, N1239);
nand NAND4 (N1504, N1491, N285, N302, N457);
not NOT1 (N1505, N1492);
nor NOR4 (N1506, N1505, N1048, N467, N41);
not NOT1 (N1507, N1499);
or OR3 (N1508, N1493, N945, N323);
and AND2 (N1509, N1501, N172);
not NOT1 (N1510, N1494);
buf BUF1 (N1511, N1506);
or OR2 (N1512, N1508, N60);
nand NAND4 (N1513, N1512, N598, N577, N558);
not NOT1 (N1514, N1513);
nand NAND4 (N1515, N1514, N124, N501, N125);
nand NAND3 (N1516, N1515, N184, N650);
or OR3 (N1517, N1497, N498, N587);
or OR4 (N1518, N1517, N618, N742, N1221);
and AND2 (N1519, N1507, N503);
nand NAND3 (N1520, N1502, N838, N1267);
xor XOR2 (N1521, N1504, N124);
not NOT1 (N1522, N1503);
nand NAND3 (N1523, N1462, N939, N786);
and AND4 (N1524, N1516, N1218, N138, N97);
or OR2 (N1525, N1521, N187);
xor XOR2 (N1526, N1509, N963);
and AND4 (N1527, N1523, N701, N861, N303);
or OR3 (N1528, N1527, N478, N683);
or OR2 (N1529, N1511, N1431);
buf BUF1 (N1530, N1510);
xor XOR2 (N1531, N1519, N753);
not NOT1 (N1532, N1525);
or OR3 (N1533, N1526, N1338, N1112);
nor NOR2 (N1534, N1532, N694);
buf BUF1 (N1535, N1518);
nor NOR2 (N1536, N1533, N917);
xor XOR2 (N1537, N1534, N1507);
and AND4 (N1538, N1531, N842, N76, N818);
not NOT1 (N1539, N1520);
buf BUF1 (N1540, N1524);
or OR4 (N1541, N1528, N854, N505, N348);
and AND2 (N1542, N1537, N943);
and AND3 (N1543, N1542, N649, N689);
buf BUF1 (N1544, N1539);
and AND2 (N1545, N1544, N1362);
and AND3 (N1546, N1530, N530, N40);
not NOT1 (N1547, N1538);
xor XOR2 (N1548, N1522, N14);
and AND2 (N1549, N1547, N879);
xor XOR2 (N1550, N1545, N1531);
or OR3 (N1551, N1540, N1228, N1297);
nand NAND2 (N1552, N1546, N1440);
not NOT1 (N1553, N1550);
nand NAND4 (N1554, N1552, N1248, N685, N429);
and AND3 (N1555, N1551, N1471, N125);
xor XOR2 (N1556, N1549, N1009);
nand NAND4 (N1557, N1555, N1179, N1067, N1168);
and AND4 (N1558, N1543, N828, N119, N520);
xor XOR2 (N1559, N1554, N853);
or OR3 (N1560, N1529, N183, N476);
nand NAND4 (N1561, N1535, N1468, N412, N337);
not NOT1 (N1562, N1560);
xor XOR2 (N1563, N1561, N1121);
nand NAND4 (N1564, N1563, N550, N267, N584);
buf BUF1 (N1565, N1541);
nor NOR2 (N1566, N1558, N1074);
and AND2 (N1567, N1536, N1054);
not NOT1 (N1568, N1565);
or OR4 (N1569, N1567, N397, N335, N1182);
buf BUF1 (N1570, N1559);
xor XOR2 (N1571, N1568, N712);
not NOT1 (N1572, N1548);
xor XOR2 (N1573, N1572, N1541);
and AND3 (N1574, N1557, N518, N714);
nor NOR2 (N1575, N1553, N762);
buf BUF1 (N1576, N1562);
and AND3 (N1577, N1569, N795, N316);
buf BUF1 (N1578, N1576);
or OR2 (N1579, N1574, N543);
buf BUF1 (N1580, N1570);
or OR2 (N1581, N1571, N1381);
nand NAND3 (N1582, N1564, N1221, N62);
nor NOR4 (N1583, N1566, N55, N664, N1326);
or OR3 (N1584, N1583, N576, N784);
nand NAND4 (N1585, N1580, N1550, N938, N725);
not NOT1 (N1586, N1585);
xor XOR2 (N1587, N1581, N659);
not NOT1 (N1588, N1575);
xor XOR2 (N1589, N1588, N1224);
and AND4 (N1590, N1584, N576, N239, N1264);
or OR2 (N1591, N1587, N706);
xor XOR2 (N1592, N1590, N1006);
nand NAND3 (N1593, N1582, N336, N356);
not NOT1 (N1594, N1579);
or OR2 (N1595, N1573, N220);
not NOT1 (N1596, N1592);
not NOT1 (N1597, N1595);
buf BUF1 (N1598, N1596);
nor NOR3 (N1599, N1578, N1356, N515);
not NOT1 (N1600, N1598);
not NOT1 (N1601, N1599);
or OR2 (N1602, N1597, N1214);
buf BUF1 (N1603, N1593);
or OR3 (N1604, N1601, N1507, N567);
nand NAND2 (N1605, N1603, N656);
nor NOR4 (N1606, N1594, N1024, N1381, N1339);
buf BUF1 (N1607, N1591);
nand NAND4 (N1608, N1556, N494, N858, N1358);
nor NOR4 (N1609, N1606, N39, N849, N1420);
nor NOR4 (N1610, N1604, N1519, N277, N70);
and AND4 (N1611, N1600, N1582, N364, N49);
buf BUF1 (N1612, N1607);
not NOT1 (N1613, N1586);
and AND4 (N1614, N1589, N337, N1386, N469);
or OR2 (N1615, N1612, N790);
xor XOR2 (N1616, N1610, N1306);
not NOT1 (N1617, N1602);
not NOT1 (N1618, N1615);
or OR4 (N1619, N1611, N1232, N82, N1315);
or OR2 (N1620, N1613, N277);
nor NOR3 (N1621, N1577, N1500, N353);
buf BUF1 (N1622, N1608);
and AND3 (N1623, N1614, N584, N1588);
and AND3 (N1624, N1617, N1327, N782);
nand NAND2 (N1625, N1616, N675);
nand NAND2 (N1626, N1605, N957);
nor NOR2 (N1627, N1618, N1602);
not NOT1 (N1628, N1626);
nor NOR4 (N1629, N1625, N1137, N896, N1429);
xor XOR2 (N1630, N1627, N41);
xor XOR2 (N1631, N1623, N895);
and AND4 (N1632, N1620, N926, N327, N1297);
or OR2 (N1633, N1619, N258);
or OR4 (N1634, N1628, N1500, N566, N1582);
xor XOR2 (N1635, N1609, N520);
not NOT1 (N1636, N1633);
nor NOR3 (N1637, N1629, N658, N1617);
xor XOR2 (N1638, N1630, N376);
and AND2 (N1639, N1631, N747);
and AND2 (N1640, N1637, N918);
or OR2 (N1641, N1640, N1075);
not NOT1 (N1642, N1639);
nor NOR3 (N1643, N1634, N581, N115);
buf BUF1 (N1644, N1636);
not NOT1 (N1645, N1644);
or OR4 (N1646, N1638, N1434, N1628, N655);
nor NOR3 (N1647, N1635, N73, N244);
not NOT1 (N1648, N1632);
not NOT1 (N1649, N1647);
nor NOR2 (N1650, N1649, N1311);
buf BUF1 (N1651, N1642);
buf BUF1 (N1652, N1648);
or OR2 (N1653, N1645, N1144);
nand NAND4 (N1654, N1653, N1492, N156, N1434);
nor NOR3 (N1655, N1643, N83, N562);
or OR3 (N1656, N1652, N1070, N132);
or OR3 (N1657, N1650, N458, N1119);
or OR2 (N1658, N1624, N5);
nand NAND2 (N1659, N1651, N453);
not NOT1 (N1660, N1622);
not NOT1 (N1661, N1641);
buf BUF1 (N1662, N1655);
not NOT1 (N1663, N1656);
not NOT1 (N1664, N1654);
not NOT1 (N1665, N1661);
buf BUF1 (N1666, N1657);
nand NAND4 (N1667, N1646, N609, N448, N1311);
nand NAND3 (N1668, N1665, N1291, N1598);
xor XOR2 (N1669, N1659, N685);
nand NAND4 (N1670, N1621, N884, N1385, N321);
nor NOR4 (N1671, N1664, N936, N306, N951);
not NOT1 (N1672, N1658);
nand NAND3 (N1673, N1667, N1230, N1545);
and AND4 (N1674, N1673, N617, N748, N1449);
nor NOR3 (N1675, N1662, N358, N1037);
xor XOR2 (N1676, N1668, N1273);
nor NOR2 (N1677, N1672, N537);
and AND3 (N1678, N1669, N1479, N899);
or OR4 (N1679, N1663, N1503, N949, N880);
not NOT1 (N1680, N1677);
xor XOR2 (N1681, N1680, N450);
not NOT1 (N1682, N1660);
or OR3 (N1683, N1682, N148, N168);
buf BUF1 (N1684, N1676);
not NOT1 (N1685, N1683);
nand NAND4 (N1686, N1674, N1285, N62, N768);
and AND3 (N1687, N1679, N856, N1120);
nand NAND3 (N1688, N1681, N1353, N1125);
not NOT1 (N1689, N1688);
buf BUF1 (N1690, N1687);
buf BUF1 (N1691, N1666);
not NOT1 (N1692, N1685);
nor NOR2 (N1693, N1689, N684);
and AND3 (N1694, N1691, N1230, N1492);
nor NOR4 (N1695, N1692, N821, N1236, N1077);
nor NOR2 (N1696, N1686, N1146);
or OR4 (N1697, N1684, N78, N803, N1306);
buf BUF1 (N1698, N1696);
buf BUF1 (N1699, N1697);
or OR4 (N1700, N1670, N66, N1442, N1591);
not NOT1 (N1701, N1678);
not NOT1 (N1702, N1675);
or OR2 (N1703, N1698, N735);
nand NAND4 (N1704, N1701, N559, N1020, N932);
and AND3 (N1705, N1695, N224, N367);
and AND2 (N1706, N1694, N1548);
nor NOR2 (N1707, N1704, N1130);
xor XOR2 (N1708, N1690, N1440);
xor XOR2 (N1709, N1708, N883);
nor NOR4 (N1710, N1709, N1343, N1153, N1253);
nand NAND4 (N1711, N1699, N468, N967, N122);
nor NOR3 (N1712, N1700, N1459, N764);
buf BUF1 (N1713, N1711);
not NOT1 (N1714, N1703);
and AND2 (N1715, N1712, N335);
or OR4 (N1716, N1713, N425, N788, N1686);
not NOT1 (N1717, N1714);
buf BUF1 (N1718, N1706);
or OR2 (N1719, N1671, N18);
buf BUF1 (N1720, N1717);
buf BUF1 (N1721, N1705);
and AND4 (N1722, N1693, N1587, N1418, N1673);
nor NOR4 (N1723, N1707, N1273, N424, N1566);
nor NOR4 (N1724, N1710, N1338, N192, N1417);
nand NAND4 (N1725, N1724, N1377, N1580, N1502);
nand NAND2 (N1726, N1722, N1627);
nand NAND3 (N1727, N1721, N1365, N1602);
buf BUF1 (N1728, N1720);
or OR3 (N1729, N1719, N504, N629);
buf BUF1 (N1730, N1726);
nor NOR4 (N1731, N1715, N1242, N450, N1692);
nor NOR4 (N1732, N1723, N1673, N202, N457);
xor XOR2 (N1733, N1732, N1459);
nand NAND3 (N1734, N1730, N450, N1322);
not NOT1 (N1735, N1728);
not NOT1 (N1736, N1733);
nand NAND4 (N1737, N1736, N198, N651, N806);
or OR4 (N1738, N1727, N1414, N1259, N449);
buf BUF1 (N1739, N1716);
nor NOR2 (N1740, N1737, N25);
nor NOR3 (N1741, N1729, N903, N1506);
buf BUF1 (N1742, N1738);
nand NAND4 (N1743, N1718, N912, N1231, N756);
nand NAND4 (N1744, N1739, N1425, N33, N1016);
and AND3 (N1745, N1734, N1093, N939);
nand NAND4 (N1746, N1735, N37, N1103, N556);
nand NAND4 (N1747, N1741, N1664, N535, N429);
and AND4 (N1748, N1745, N14, N613, N940);
and AND3 (N1749, N1743, N136, N1014);
xor XOR2 (N1750, N1740, N1520);
xor XOR2 (N1751, N1750, N467);
xor XOR2 (N1752, N1746, N301);
xor XOR2 (N1753, N1742, N372);
xor XOR2 (N1754, N1748, N865);
nor NOR4 (N1755, N1752, N213, N757, N24);
buf BUF1 (N1756, N1731);
buf BUF1 (N1757, N1747);
or OR4 (N1758, N1725, N1146, N1468, N724);
nor NOR4 (N1759, N1749, N498, N641, N373);
xor XOR2 (N1760, N1754, N1444);
nand NAND3 (N1761, N1755, N1446, N1329);
not NOT1 (N1762, N1760);
or OR4 (N1763, N1744, N1119, N1092, N1597);
buf BUF1 (N1764, N1759);
xor XOR2 (N1765, N1763, N1043);
xor XOR2 (N1766, N1751, N1521);
nand NAND4 (N1767, N1758, N726, N441, N798);
not NOT1 (N1768, N1702);
nand NAND3 (N1769, N1753, N1451, N579);
nand NAND2 (N1770, N1756, N1072);
xor XOR2 (N1771, N1768, N686);
nand NAND3 (N1772, N1761, N867, N1612);
buf BUF1 (N1773, N1772);
nand NAND3 (N1774, N1762, N1276, N69);
nand NAND2 (N1775, N1767, N1070);
not NOT1 (N1776, N1757);
xor XOR2 (N1777, N1770, N1501);
buf BUF1 (N1778, N1771);
nor NOR3 (N1779, N1773, N711, N721);
or OR2 (N1780, N1778, N78);
buf BUF1 (N1781, N1766);
not NOT1 (N1782, N1777);
nor NOR2 (N1783, N1780, N267);
nand NAND4 (N1784, N1779, N768, N1137, N1396);
xor XOR2 (N1785, N1781, N647);
or OR4 (N1786, N1775, N86, N1531, N12);
buf BUF1 (N1787, N1782);
nand NAND3 (N1788, N1783, N399, N1041);
nand NAND2 (N1789, N1764, N62);
not NOT1 (N1790, N1776);
nand NAND3 (N1791, N1765, N1066, N559);
or OR2 (N1792, N1787, N385);
nor NOR2 (N1793, N1792, N396);
nor NOR2 (N1794, N1791, N245);
or OR4 (N1795, N1785, N1047, N920, N49);
not NOT1 (N1796, N1793);
xor XOR2 (N1797, N1789, N619);
or OR2 (N1798, N1796, N301);
xor XOR2 (N1799, N1794, N1490);
not NOT1 (N1800, N1786);
xor XOR2 (N1801, N1788, N802);
buf BUF1 (N1802, N1795);
nand NAND2 (N1803, N1798, N851);
not NOT1 (N1804, N1802);
nor NOR3 (N1805, N1801, N416, N904);
and AND4 (N1806, N1774, N1283, N1231, N1458);
and AND3 (N1807, N1799, N1450, N277);
nor NOR3 (N1808, N1805, N1152, N358);
or OR4 (N1809, N1769, N137, N1519, N513);
nand NAND2 (N1810, N1807, N812);
and AND3 (N1811, N1797, N1041, N966);
or OR4 (N1812, N1810, N990, N1147, N854);
buf BUF1 (N1813, N1808);
nand NAND2 (N1814, N1813, N600);
and AND2 (N1815, N1804, N812);
nor NOR3 (N1816, N1812, N180, N1482);
nand NAND3 (N1817, N1790, N972, N119);
and AND4 (N1818, N1814, N497, N241, N904);
xor XOR2 (N1819, N1806, N3);
or OR3 (N1820, N1803, N258, N1148);
or OR4 (N1821, N1818, N915, N1710, N503);
nand NAND4 (N1822, N1817, N377, N980, N444);
nand NAND3 (N1823, N1820, N1414, N1039);
buf BUF1 (N1824, N1784);
nor NOR3 (N1825, N1811, N1376, N936);
xor XOR2 (N1826, N1809, N53);
nand NAND4 (N1827, N1826, N1576, N1817, N949);
xor XOR2 (N1828, N1827, N726);
xor XOR2 (N1829, N1819, N197);
nand NAND4 (N1830, N1816, N414, N905, N841);
nand NAND2 (N1831, N1824, N1451);
and AND2 (N1832, N1829, N429);
nand NAND2 (N1833, N1800, N542);
xor XOR2 (N1834, N1830, N722);
not NOT1 (N1835, N1828);
nor NOR4 (N1836, N1833, N1079, N1049, N1210);
xor XOR2 (N1837, N1836, N591);
not NOT1 (N1838, N1832);
buf BUF1 (N1839, N1838);
and AND2 (N1840, N1823, N1582);
nand NAND3 (N1841, N1837, N135, N482);
not NOT1 (N1842, N1841);
buf BUF1 (N1843, N1839);
buf BUF1 (N1844, N1822);
not NOT1 (N1845, N1843);
or OR3 (N1846, N1834, N1694, N879);
buf BUF1 (N1847, N1835);
nor NOR3 (N1848, N1847, N171, N1658);
not NOT1 (N1849, N1831);
and AND3 (N1850, N1844, N339, N1647);
nand NAND2 (N1851, N1821, N1769);
buf BUF1 (N1852, N1842);
buf BUF1 (N1853, N1851);
nor NOR4 (N1854, N1853, N1389, N417, N1277);
or OR4 (N1855, N1850, N1666, N289, N1425);
nor NOR2 (N1856, N1815, N914);
xor XOR2 (N1857, N1855, N1588);
not NOT1 (N1858, N1825);
buf BUF1 (N1859, N1849);
not NOT1 (N1860, N1840);
not NOT1 (N1861, N1860);
buf BUF1 (N1862, N1856);
xor XOR2 (N1863, N1854, N843);
or OR4 (N1864, N1861, N170, N1691, N1687);
and AND4 (N1865, N1864, N1279, N565, N969);
buf BUF1 (N1866, N1857);
xor XOR2 (N1867, N1863, N1552);
or OR4 (N1868, N1865, N1422, N977, N291);
and AND2 (N1869, N1862, N951);
buf BUF1 (N1870, N1848);
nor NOR4 (N1871, N1868, N340, N736, N1739);
xor XOR2 (N1872, N1852, N233);
and AND3 (N1873, N1845, N1501, N1653);
not NOT1 (N1874, N1872);
buf BUF1 (N1875, N1866);
and AND4 (N1876, N1874, N1867, N1537, N84);
xor XOR2 (N1877, N1498, N1374);
buf BUF1 (N1878, N1870);
xor XOR2 (N1879, N1859, N1758);
nand NAND2 (N1880, N1876, N1181);
and AND4 (N1881, N1869, N823, N1628, N1150);
and AND4 (N1882, N1881, N148, N1382, N1467);
nand NAND2 (N1883, N1846, N1429);
and AND2 (N1884, N1882, N1640);
nor NOR4 (N1885, N1884, N1158, N460, N1496);
and AND3 (N1886, N1858, N1667, N1019);
xor XOR2 (N1887, N1871, N1743);
nand NAND4 (N1888, N1887, N1367, N1380, N1113);
not NOT1 (N1889, N1875);
not NOT1 (N1890, N1877);
or OR4 (N1891, N1889, N1102, N1326, N1878);
and AND2 (N1892, N532, N839);
or OR2 (N1893, N1886, N1750);
nor NOR2 (N1894, N1891, N1599);
xor XOR2 (N1895, N1885, N1121);
xor XOR2 (N1896, N1880, N1715);
buf BUF1 (N1897, N1896);
or OR4 (N1898, N1892, N96, N1834, N1615);
buf BUF1 (N1899, N1883);
and AND3 (N1900, N1898, N195, N1028);
nand NAND4 (N1901, N1890, N1777, N1583, N1289);
and AND2 (N1902, N1888, N105);
buf BUF1 (N1903, N1879);
xor XOR2 (N1904, N1900, N222);
buf BUF1 (N1905, N1899);
not NOT1 (N1906, N1894);
or OR3 (N1907, N1873, N186, N560);
buf BUF1 (N1908, N1895);
not NOT1 (N1909, N1904);
and AND4 (N1910, N1897, N366, N1120, N461);
or OR4 (N1911, N1893, N607, N1098, N1830);
nor NOR4 (N1912, N1906, N1904, N1643, N1106);
or OR2 (N1913, N1911, N392);
not NOT1 (N1914, N1905);
or OR3 (N1915, N1909, N1697, N1481);
buf BUF1 (N1916, N1902);
buf BUF1 (N1917, N1916);
xor XOR2 (N1918, N1913, N1745);
xor XOR2 (N1919, N1908, N629);
or OR4 (N1920, N1919, N731, N36, N1537);
or OR3 (N1921, N1910, N1154, N451);
buf BUF1 (N1922, N1918);
xor XOR2 (N1923, N1921, N940);
and AND4 (N1924, N1920, N600, N1468, N936);
nor NOR3 (N1925, N1901, N702, N731);
buf BUF1 (N1926, N1907);
and AND2 (N1927, N1926, N413);
buf BUF1 (N1928, N1922);
and AND3 (N1929, N1928, N256, N605);
or OR4 (N1930, N1915, N360, N386, N1576);
and AND3 (N1931, N1903, N1455, N190);
and AND4 (N1932, N1924, N1364, N224, N696);
not NOT1 (N1933, N1930);
xor XOR2 (N1934, N1914, N1406);
not NOT1 (N1935, N1923);
not NOT1 (N1936, N1933);
xor XOR2 (N1937, N1927, N760);
buf BUF1 (N1938, N1931);
not NOT1 (N1939, N1917);
or OR3 (N1940, N1929, N484, N86);
and AND2 (N1941, N1939, N197);
xor XOR2 (N1942, N1937, N746);
nor NOR3 (N1943, N1942, N761, N963);
not NOT1 (N1944, N1935);
nand NAND3 (N1945, N1912, N170, N1899);
nand NAND2 (N1946, N1934, N1721);
xor XOR2 (N1947, N1936, N1907);
buf BUF1 (N1948, N1938);
and AND3 (N1949, N1946, N1385, N1793);
not NOT1 (N1950, N1948);
xor XOR2 (N1951, N1947, N918);
and AND2 (N1952, N1944, N1525);
buf BUF1 (N1953, N1941);
not NOT1 (N1954, N1943);
xor XOR2 (N1955, N1932, N1491);
or OR2 (N1956, N1925, N1769);
nor NOR2 (N1957, N1949, N379);
or OR3 (N1958, N1945, N1789, N1816);
xor XOR2 (N1959, N1950, N1332);
buf BUF1 (N1960, N1953);
or OR2 (N1961, N1952, N408);
buf BUF1 (N1962, N1959);
and AND4 (N1963, N1958, N1796, N764, N118);
buf BUF1 (N1964, N1963);
or OR2 (N1965, N1954, N1409);
or OR3 (N1966, N1955, N1803, N1305);
nor NOR2 (N1967, N1966, N1620);
and AND4 (N1968, N1957, N1596, N566, N1356);
nand NAND2 (N1969, N1956, N11);
xor XOR2 (N1970, N1951, N824);
nand NAND4 (N1971, N1964, N1770, N559, N396);
or OR2 (N1972, N1960, N306);
and AND4 (N1973, N1965, N323, N1908, N606);
not NOT1 (N1974, N1970);
xor XOR2 (N1975, N1961, N197);
not NOT1 (N1976, N1972);
not NOT1 (N1977, N1971);
xor XOR2 (N1978, N1975, N1475);
xor XOR2 (N1979, N1978, N666);
nor NOR3 (N1980, N1976, N180, N664);
buf BUF1 (N1981, N1940);
nand NAND2 (N1982, N1962, N1685);
buf BUF1 (N1983, N1968);
nand NAND3 (N1984, N1974, N830, N1886);
nor NOR2 (N1985, N1977, N1279);
xor XOR2 (N1986, N1969, N616);
nor NOR4 (N1987, N1980, N1064, N745, N1825);
nor NOR2 (N1988, N1984, N1820);
not NOT1 (N1989, N1988);
buf BUF1 (N1990, N1987);
buf BUF1 (N1991, N1967);
xor XOR2 (N1992, N1983, N152);
buf BUF1 (N1993, N1979);
and AND2 (N1994, N1992, N1923);
xor XOR2 (N1995, N1985, N1654);
or OR3 (N1996, N1986, N1262, N1907);
nor NOR3 (N1997, N1993, N471, N1124);
and AND3 (N1998, N1991, N1884, N900);
nor NOR2 (N1999, N1981, N431);
and AND3 (N2000, N1990, N490, N1228);
and AND4 (N2001, N1997, N1772, N609, N1444);
or OR3 (N2002, N1998, N570, N668);
nor NOR4 (N2003, N2001, N134, N1049, N1589);
or OR3 (N2004, N2003, N804, N1829);
not NOT1 (N2005, N1999);
or OR2 (N2006, N2005, N714);
nor NOR2 (N2007, N1994, N465);
buf BUF1 (N2008, N1973);
or OR4 (N2009, N2002, N1113, N1264, N231);
nor NOR2 (N2010, N1996, N180);
nor NOR3 (N2011, N1982, N1469, N1733);
or OR2 (N2012, N2010, N1804);
xor XOR2 (N2013, N1995, N356);
not NOT1 (N2014, N2008);
xor XOR2 (N2015, N2014, N1701);
nand NAND3 (N2016, N2007, N159, N397);
buf BUF1 (N2017, N2004);
nand NAND3 (N2018, N2000, N107, N1966);
xor XOR2 (N2019, N2016, N1607);
or OR2 (N2020, N2015, N889);
not NOT1 (N2021, N2009);
nand NAND3 (N2022, N2013, N1053, N1211);
or OR2 (N2023, N2011, N1585);
not NOT1 (N2024, N2023);
and AND4 (N2025, N2024, N173, N167, N1857);
not NOT1 (N2026, N2012);
xor XOR2 (N2027, N2025, N909);
xor XOR2 (N2028, N2026, N1648);
and AND4 (N2029, N2006, N1707, N1168, N1494);
buf BUF1 (N2030, N2020);
xor XOR2 (N2031, N2028, N346);
xor XOR2 (N2032, N2021, N1499);
and AND4 (N2033, N2030, N1997, N790, N1870);
nand NAND3 (N2034, N2019, N1983, N1593);
not NOT1 (N2035, N2022);
not NOT1 (N2036, N2018);
not NOT1 (N2037, N2032);
not NOT1 (N2038, N2029);
not NOT1 (N2039, N2034);
and AND2 (N2040, N2033, N712);
not NOT1 (N2041, N2031);
or OR3 (N2042, N2037, N1394, N621);
not NOT1 (N2043, N1989);
buf BUF1 (N2044, N2040);
or OR3 (N2045, N2041, N201, N301);
xor XOR2 (N2046, N2038, N115);
xor XOR2 (N2047, N2043, N1590);
xor XOR2 (N2048, N2045, N1347);
not NOT1 (N2049, N2044);
xor XOR2 (N2050, N2046, N28);
xor XOR2 (N2051, N2050, N1895);
buf BUF1 (N2052, N2039);
and AND4 (N2053, N2047, N2043, N1888, N1364);
buf BUF1 (N2054, N2048);
and AND4 (N2055, N2054, N1665, N60, N1742);
and AND4 (N2056, N2017, N1477, N1387, N1185);
buf BUF1 (N2057, N2053);
nor NOR3 (N2058, N2057, N281, N656);
nand NAND2 (N2059, N2058, N614);
nor NOR2 (N2060, N2049, N1702);
buf BUF1 (N2061, N2055);
nor NOR3 (N2062, N2042, N557, N2033);
and AND3 (N2063, N2056, N1057, N348);
or OR2 (N2064, N2052, N1737);
or OR3 (N2065, N2063, N50, N2039);
nor NOR2 (N2066, N2051, N1893);
or OR2 (N2067, N2059, N302);
xor XOR2 (N2068, N2060, N817);
nor NOR4 (N2069, N2061, N289, N118, N1411);
xor XOR2 (N2070, N2027, N1462);
not NOT1 (N2071, N2070);
and AND2 (N2072, N2064, N999);
xor XOR2 (N2073, N2036, N390);
nor NOR4 (N2074, N2066, N101, N329, N1936);
xor XOR2 (N2075, N2072, N40);
xor XOR2 (N2076, N2035, N1905);
buf BUF1 (N2077, N2075);
and AND4 (N2078, N2073, N1250, N1246, N468);
nor NOR3 (N2079, N2062, N1707, N1255);
nor NOR3 (N2080, N2077, N478, N37);
nand NAND4 (N2081, N2080, N1033, N186, N352);
nor NOR2 (N2082, N2071, N1594);
and AND3 (N2083, N2078, N1352, N928);
nor NOR4 (N2084, N2082, N751, N1166, N1635);
not NOT1 (N2085, N2084);
and AND3 (N2086, N2065, N886, N1474);
or OR2 (N2087, N2067, N1788);
nand NAND4 (N2088, N2068, N1170, N1494, N371);
nand NAND3 (N2089, N2085, N692, N1866);
nor NOR4 (N2090, N2088, N951, N903, N73);
nor NOR4 (N2091, N2079, N117, N2081, N601);
xor XOR2 (N2092, N448, N1992);
buf BUF1 (N2093, N2090);
nor NOR4 (N2094, N2076, N1638, N619, N843);
nand NAND3 (N2095, N2074, N232, N1185);
nand NAND2 (N2096, N2089, N1649);
nand NAND3 (N2097, N2083, N1662, N769);
not NOT1 (N2098, N2093);
nor NOR2 (N2099, N2096, N1357);
not NOT1 (N2100, N2092);
nand NAND3 (N2101, N2094, N1837, N838);
and AND2 (N2102, N2098, N752);
buf BUF1 (N2103, N2069);
and AND3 (N2104, N2103, N1960, N1481);
or OR4 (N2105, N2087, N1440, N947, N505);
not NOT1 (N2106, N2100);
and AND4 (N2107, N2104, N1351, N167, N817);
and AND3 (N2108, N2099, N2064, N355);
not NOT1 (N2109, N2097);
and AND2 (N2110, N2107, N1065);
not NOT1 (N2111, N2095);
nand NAND4 (N2112, N2101, N1562, N640, N712);
or OR2 (N2113, N2091, N1663);
not NOT1 (N2114, N2111);
buf BUF1 (N2115, N2105);
not NOT1 (N2116, N2115);
nor NOR2 (N2117, N2114, N929);
not NOT1 (N2118, N2102);
not NOT1 (N2119, N2106);
and AND3 (N2120, N2113, N873, N391);
nand NAND3 (N2121, N2110, N1063, N1654);
nor NOR3 (N2122, N2121, N507, N1241);
buf BUF1 (N2123, N2122);
xor XOR2 (N2124, N2117, N1116);
not NOT1 (N2125, N2118);
or OR2 (N2126, N2108, N878);
nand NAND2 (N2127, N2112, N325);
nand NAND3 (N2128, N2123, N1132, N633);
nand NAND3 (N2129, N2125, N33, N1605);
buf BUF1 (N2130, N2129);
xor XOR2 (N2131, N2119, N1859);
nor NOR4 (N2132, N2120, N536, N266, N1210);
buf BUF1 (N2133, N2128);
nand NAND4 (N2134, N2131, N923, N584, N845);
xor XOR2 (N2135, N2086, N219);
not NOT1 (N2136, N2124);
nor NOR4 (N2137, N2126, N1848, N750, N1390);
not NOT1 (N2138, N2137);
nor NOR4 (N2139, N2134, N927, N1158, N89);
not NOT1 (N2140, N2130);
xor XOR2 (N2141, N2136, N1081);
nand NAND4 (N2142, N2132, N1259, N1515, N2109);
and AND3 (N2143, N790, N1944, N1890);
xor XOR2 (N2144, N2133, N1559);
xor XOR2 (N2145, N2140, N816);
nor NOR4 (N2146, N2143, N71, N1124, N1573);
nand NAND3 (N2147, N2145, N273, N1765);
and AND3 (N2148, N2135, N617, N115);
buf BUF1 (N2149, N2147);
nor NOR2 (N2150, N2144, N1938);
buf BUF1 (N2151, N2139);
nor NOR2 (N2152, N2148, N2058);
and AND2 (N2153, N2151, N1308);
nor NOR3 (N2154, N2152, N1586, N527);
buf BUF1 (N2155, N2127);
buf BUF1 (N2156, N2142);
not NOT1 (N2157, N2155);
or OR4 (N2158, N2153, N1291, N337, N384);
nand NAND3 (N2159, N2150, N605, N298);
or OR3 (N2160, N2116, N2142, N1718);
xor XOR2 (N2161, N2146, N754);
buf BUF1 (N2162, N2154);
nand NAND3 (N2163, N2159, N326, N1342);
not NOT1 (N2164, N2162);
or OR3 (N2165, N2164, N357, N1940);
buf BUF1 (N2166, N2165);
nor NOR3 (N2167, N2166, N2094, N2048);
and AND4 (N2168, N2141, N1830, N1809, N2001);
not NOT1 (N2169, N2161);
not NOT1 (N2170, N2167);
nor NOR4 (N2171, N2169, N106, N667, N396);
not NOT1 (N2172, N2163);
not NOT1 (N2173, N2160);
buf BUF1 (N2174, N2138);
not NOT1 (N2175, N2149);
buf BUF1 (N2176, N2175);
and AND2 (N2177, N2172, N1460);
and AND3 (N2178, N2171, N238, N431);
not NOT1 (N2179, N2177);
nand NAND3 (N2180, N2173, N692, N947);
xor XOR2 (N2181, N2157, N517);
and AND4 (N2182, N2158, N1139, N753, N1072);
and AND4 (N2183, N2178, N1739, N714, N1905);
nand NAND2 (N2184, N2170, N100);
not NOT1 (N2185, N2168);
and AND4 (N2186, N2183, N849, N101, N1523);
or OR3 (N2187, N2182, N1630, N1087);
or OR2 (N2188, N2176, N604);
or OR3 (N2189, N2188, N1418, N315);
xor XOR2 (N2190, N2185, N1321);
and AND2 (N2191, N2179, N554);
xor XOR2 (N2192, N2190, N535);
and AND3 (N2193, N2174, N2022, N1668);
not NOT1 (N2194, N2180);
xor XOR2 (N2195, N2192, N452);
or OR3 (N2196, N2191, N1329, N988);
nor NOR2 (N2197, N2184, N810);
xor XOR2 (N2198, N2156, N2082);
buf BUF1 (N2199, N2198);
nor NOR2 (N2200, N2195, N235);
nor NOR4 (N2201, N2197, N1501, N1876, N20);
and AND3 (N2202, N2193, N1587, N1564);
nand NAND2 (N2203, N2187, N1873);
xor XOR2 (N2204, N2202, N1118);
and AND4 (N2205, N2189, N745, N1170, N1104);
xor XOR2 (N2206, N2204, N1828);
and AND3 (N2207, N2186, N1959, N1543);
not NOT1 (N2208, N2196);
or OR3 (N2209, N2206, N1368, N127);
or OR2 (N2210, N2207, N1788);
not NOT1 (N2211, N2201);
not NOT1 (N2212, N2209);
not NOT1 (N2213, N2200);
xor XOR2 (N2214, N2203, N1840);
not NOT1 (N2215, N2214);
nor NOR3 (N2216, N2211, N433, N1758);
or OR4 (N2217, N2199, N677, N1403, N1568);
buf BUF1 (N2218, N2213);
buf BUF1 (N2219, N2205);
not NOT1 (N2220, N2181);
xor XOR2 (N2221, N2208, N623);
buf BUF1 (N2222, N2219);
nand NAND4 (N2223, N2218, N1047, N62, N1087);
nand NAND2 (N2224, N2194, N1677);
not NOT1 (N2225, N2216);
nor NOR3 (N2226, N2221, N1315, N294);
nand NAND3 (N2227, N2212, N2197, N303);
nor NOR2 (N2228, N2223, N1515);
xor XOR2 (N2229, N2226, N2101);
not NOT1 (N2230, N2210);
nor NOR4 (N2231, N2225, N2211, N997, N1504);
buf BUF1 (N2232, N2224);
nand NAND4 (N2233, N2215, N2101, N522, N1968);
nand NAND2 (N2234, N2228, N1793);
not NOT1 (N2235, N2231);
or OR4 (N2236, N2233, N506, N908, N2127);
nor NOR4 (N2237, N2232, N1015, N1334, N34);
nor NOR4 (N2238, N2220, N486, N1975, N1701);
nand NAND2 (N2239, N2229, N1936);
nand NAND4 (N2240, N2237, N435, N889, N197);
buf BUF1 (N2241, N2222);
and AND3 (N2242, N2227, N1322, N1176);
buf BUF1 (N2243, N2240);
and AND4 (N2244, N2234, N668, N389, N78);
nor NOR2 (N2245, N2238, N1822);
buf BUF1 (N2246, N2244);
or OR4 (N2247, N2242, N164, N1183, N341);
or OR3 (N2248, N2247, N1226, N1187);
and AND2 (N2249, N2243, N91);
and AND3 (N2250, N2235, N2165, N423);
nor NOR4 (N2251, N2241, N133, N889, N1912);
and AND3 (N2252, N2230, N1819, N2037);
not NOT1 (N2253, N2251);
not NOT1 (N2254, N2217);
and AND2 (N2255, N2236, N1345);
or OR2 (N2256, N2253, N2002);
buf BUF1 (N2257, N2252);
buf BUF1 (N2258, N2239);
nand NAND3 (N2259, N2258, N2161, N1182);
nand NAND4 (N2260, N2254, N372, N1964, N1491);
or OR3 (N2261, N2256, N192, N779);
and AND4 (N2262, N2250, N1473, N1789, N1025);
buf BUF1 (N2263, N2261);
buf BUF1 (N2264, N2262);
or OR2 (N2265, N2259, N521);
buf BUF1 (N2266, N2255);
nand NAND3 (N2267, N2249, N732, N470);
nand NAND3 (N2268, N2263, N2070, N1209);
buf BUF1 (N2269, N2260);
or OR2 (N2270, N2257, N2072);
nand NAND4 (N2271, N2270, N1130, N1311, N481);
buf BUF1 (N2272, N2264);
xor XOR2 (N2273, N2265, N1196);
nand NAND4 (N2274, N2267, N1798, N1395, N1430);
or OR2 (N2275, N2266, N396);
and AND4 (N2276, N2271, N162, N538, N1747);
nor NOR2 (N2277, N2248, N586);
xor XOR2 (N2278, N2275, N667);
xor XOR2 (N2279, N2278, N333);
or OR2 (N2280, N2269, N1102);
or OR2 (N2281, N2276, N770);
and AND3 (N2282, N2280, N1670, N672);
or OR3 (N2283, N2272, N1684, N806);
nor NOR4 (N2284, N2273, N622, N277, N1658);
nand NAND4 (N2285, N2284, N352, N2219, N60);
and AND2 (N2286, N2274, N1952);
nor NOR2 (N2287, N2282, N445);
or OR2 (N2288, N2277, N1125);
xor XOR2 (N2289, N2288, N2128);
or OR2 (N2290, N2245, N294);
nand NAND3 (N2291, N2286, N1558, N515);
buf BUF1 (N2292, N2246);
and AND4 (N2293, N2292, N1481, N1740, N2224);
not NOT1 (N2294, N2289);
nor NOR4 (N2295, N2290, N954, N49, N952);
nand NAND2 (N2296, N2294, N1990);
nand NAND4 (N2297, N2296, N1666, N2256, N1136);
buf BUF1 (N2298, N2281);
not NOT1 (N2299, N2291);
nand NAND3 (N2300, N2287, N398, N1635);
nand NAND4 (N2301, N2285, N1227, N1085, N1513);
xor XOR2 (N2302, N2283, N1605);
nand NAND2 (N2303, N2295, N817);
nor NOR4 (N2304, N2293, N1238, N1266, N1229);
not NOT1 (N2305, N2304);
nor NOR4 (N2306, N2305, N687, N1884, N347);
buf BUF1 (N2307, N2306);
buf BUF1 (N2308, N2268);
not NOT1 (N2309, N2299);
or OR3 (N2310, N2279, N2285, N2013);
xor XOR2 (N2311, N2302, N54);
buf BUF1 (N2312, N2307);
nor NOR3 (N2313, N2298, N52, N591);
and AND4 (N2314, N2308, N1280, N1067, N1941);
nand NAND4 (N2315, N2300, N1634, N380, N1889);
not NOT1 (N2316, N2311);
or OR3 (N2317, N2303, N2145, N683);
nand NAND2 (N2318, N2312, N732);
or OR3 (N2319, N2316, N1480, N598);
not NOT1 (N2320, N2319);
nor NOR4 (N2321, N2317, N1251, N485, N584);
nand NAND3 (N2322, N2313, N1626, N964);
nand NAND2 (N2323, N2321, N460);
nor NOR2 (N2324, N2323, N817);
not NOT1 (N2325, N2297);
and AND4 (N2326, N2310, N2066, N804, N1068);
buf BUF1 (N2327, N2301);
and AND2 (N2328, N2326, N1050);
or OR3 (N2329, N2314, N1249, N2137);
xor XOR2 (N2330, N2327, N189);
xor XOR2 (N2331, N2328, N2285);
xor XOR2 (N2332, N2322, N1613);
nand NAND3 (N2333, N2330, N1572, N1737);
nand NAND4 (N2334, N2332, N2125, N686, N422);
not NOT1 (N2335, N2329);
not NOT1 (N2336, N2331);
not NOT1 (N2337, N2335);
not NOT1 (N2338, N2315);
or OR3 (N2339, N2336, N1503, N1496);
and AND3 (N2340, N2309, N807, N983);
buf BUF1 (N2341, N2337);
and AND2 (N2342, N2341, N759);
xor XOR2 (N2343, N2318, N1849);
not NOT1 (N2344, N2325);
xor XOR2 (N2345, N2339, N1506);
xor XOR2 (N2346, N2343, N1960);
and AND4 (N2347, N2324, N631, N943, N440);
and AND4 (N2348, N2334, N2255, N1311, N713);
buf BUF1 (N2349, N2345);
and AND3 (N2350, N2347, N880, N1556);
xor XOR2 (N2351, N2340, N50);
and AND4 (N2352, N2320, N1861, N280, N1723);
buf BUF1 (N2353, N2344);
buf BUF1 (N2354, N2353);
nand NAND4 (N2355, N2349, N21, N2005, N1875);
or OR2 (N2356, N2348, N2291);
nand NAND2 (N2357, N2333, N1143);
nand NAND3 (N2358, N2338, N10, N1037);
nor NOR2 (N2359, N2358, N725);
and AND2 (N2360, N2359, N1156);
xor XOR2 (N2361, N2350, N2209);
xor XOR2 (N2362, N2355, N1473);
buf BUF1 (N2363, N2362);
buf BUF1 (N2364, N2360);
buf BUF1 (N2365, N2342);
not NOT1 (N2366, N2365);
xor XOR2 (N2367, N2352, N2320);
nor NOR4 (N2368, N2363, N567, N6, N1710);
not NOT1 (N2369, N2346);
buf BUF1 (N2370, N2369);
nand NAND4 (N2371, N2366, N23, N665, N1671);
nor NOR3 (N2372, N2368, N1998, N1099);
nand NAND2 (N2373, N2370, N1723);
buf BUF1 (N2374, N2354);
nor NOR4 (N2375, N2364, N1491, N1670, N1651);
nand NAND4 (N2376, N2356, N183, N2364, N1379);
buf BUF1 (N2377, N2376);
not NOT1 (N2378, N2373);
buf BUF1 (N2379, N2375);
xor XOR2 (N2380, N2351, N2320);
or OR4 (N2381, N2374, N1758, N14, N323);
nor NOR3 (N2382, N2379, N474, N245);
nand NAND4 (N2383, N2372, N2082, N2263, N41);
not NOT1 (N2384, N2382);
xor XOR2 (N2385, N2378, N515);
xor XOR2 (N2386, N2381, N1715);
and AND2 (N2387, N2367, N751);
and AND3 (N2388, N2383, N1917, N1844);
nor NOR2 (N2389, N2380, N1827);
and AND3 (N2390, N2361, N1323, N514);
xor XOR2 (N2391, N2385, N1500);
nand NAND4 (N2392, N2387, N2295, N477, N293);
or OR4 (N2393, N2377, N343, N1632, N1918);
nor NOR3 (N2394, N2384, N541, N1259);
nand NAND2 (N2395, N2386, N1894);
buf BUF1 (N2396, N2395);
nor NOR2 (N2397, N2357, N433);
or OR4 (N2398, N2391, N1308, N2269, N737);
not NOT1 (N2399, N2388);
and AND3 (N2400, N2394, N2016, N1526);
not NOT1 (N2401, N2389);
nand NAND3 (N2402, N2371, N2115, N1021);
or OR2 (N2403, N2390, N1941);
not NOT1 (N2404, N2392);
not NOT1 (N2405, N2398);
nand NAND2 (N2406, N2397, N811);
not NOT1 (N2407, N2402);
xor XOR2 (N2408, N2407, N854);
nor NOR4 (N2409, N2405, N1374, N838, N2227);
nand NAND2 (N2410, N2406, N654);
buf BUF1 (N2411, N2404);
and AND3 (N2412, N2410, N97, N800);
nor NOR3 (N2413, N2411, N2281, N1634);
nand NAND2 (N2414, N2399, N876);
xor XOR2 (N2415, N2400, N2160);
nor NOR2 (N2416, N2403, N265);
not NOT1 (N2417, N2415);
nor NOR4 (N2418, N2408, N1138, N1908, N1751);
or OR3 (N2419, N2417, N1197, N872);
and AND2 (N2420, N2396, N602);
buf BUF1 (N2421, N2409);
not NOT1 (N2422, N2421);
xor XOR2 (N2423, N2416, N1589);
and AND2 (N2424, N2418, N476);
or OR3 (N2425, N2414, N30, N663);
nor NOR4 (N2426, N2423, N121, N1231, N1862);
and AND4 (N2427, N2422, N1015, N897, N174);
xor XOR2 (N2428, N2412, N941);
buf BUF1 (N2429, N2393);
and AND4 (N2430, N2428, N2378, N562, N269);
buf BUF1 (N2431, N2401);
xor XOR2 (N2432, N2429, N1764);
not NOT1 (N2433, N2413);
xor XOR2 (N2434, N2430, N1970);
and AND3 (N2435, N2420, N72, N199);
xor XOR2 (N2436, N2434, N1546);
or OR4 (N2437, N2431, N2002, N739, N1044);
nor NOR2 (N2438, N2432, N441);
buf BUF1 (N2439, N2437);
xor XOR2 (N2440, N2438, N67);
nor NOR3 (N2441, N2427, N1153, N2134);
not NOT1 (N2442, N2441);
or OR4 (N2443, N2435, N1170, N1379, N475);
not NOT1 (N2444, N2419);
buf BUF1 (N2445, N2442);
nand NAND2 (N2446, N2433, N334);
buf BUF1 (N2447, N2425);
not NOT1 (N2448, N2436);
xor XOR2 (N2449, N2426, N72);
or OR2 (N2450, N2448, N439);
buf BUF1 (N2451, N2440);
not NOT1 (N2452, N2447);
and AND4 (N2453, N2449, N1095, N2265, N105);
buf BUF1 (N2454, N2453);
not NOT1 (N2455, N2439);
xor XOR2 (N2456, N2443, N1116);
xor XOR2 (N2457, N2454, N614);
xor XOR2 (N2458, N2456, N1613);
not NOT1 (N2459, N2455);
buf BUF1 (N2460, N2444);
buf BUF1 (N2461, N2445);
or OR4 (N2462, N2450, N2212, N1489, N2187);
not NOT1 (N2463, N2451);
not NOT1 (N2464, N2458);
nor NOR3 (N2465, N2464, N1402, N1421);
buf BUF1 (N2466, N2457);
buf BUF1 (N2467, N2462);
not NOT1 (N2468, N2461);
nor NOR3 (N2469, N2468, N452, N1439);
nor NOR2 (N2470, N2424, N1582);
not NOT1 (N2471, N2446);
or OR2 (N2472, N2467, N1150);
or OR3 (N2473, N2459, N1120, N1534);
xor XOR2 (N2474, N2465, N1286);
and AND4 (N2475, N2466, N2459, N2362, N2337);
nand NAND3 (N2476, N2474, N938, N2424);
xor XOR2 (N2477, N2471, N1348);
xor XOR2 (N2478, N2472, N1224);
nand NAND3 (N2479, N2460, N1166, N635);
or OR4 (N2480, N2470, N504, N2015, N656);
or OR2 (N2481, N2473, N1295);
xor XOR2 (N2482, N2476, N413);
or OR3 (N2483, N2479, N2339, N2229);
nand NAND4 (N2484, N2482, N1667, N972, N658);
and AND2 (N2485, N2452, N1584);
xor XOR2 (N2486, N2463, N2199);
nor NOR3 (N2487, N2486, N866, N2211);
and AND4 (N2488, N2469, N414, N473, N1482);
not NOT1 (N2489, N2481);
and AND4 (N2490, N2483, N1516, N647, N2268);
xor XOR2 (N2491, N2489, N580);
xor XOR2 (N2492, N2478, N1796);
not NOT1 (N2493, N2491);
nor NOR3 (N2494, N2475, N318, N2244);
xor XOR2 (N2495, N2492, N687);
buf BUF1 (N2496, N2494);
nand NAND2 (N2497, N2488, N1277);
buf BUF1 (N2498, N2484);
or OR2 (N2499, N2497, N1943);
xor XOR2 (N2500, N2499, N511);
buf BUF1 (N2501, N2477);
nor NOR2 (N2502, N2490, N903);
nor NOR4 (N2503, N2501, N1198, N96, N2342);
or OR2 (N2504, N2485, N1574);
xor XOR2 (N2505, N2496, N2216);
xor XOR2 (N2506, N2500, N517);
nand NAND3 (N2507, N2502, N2182, N1081);
xor XOR2 (N2508, N2503, N2231);
nor NOR2 (N2509, N2480, N464);
and AND3 (N2510, N2504, N897, N986);
or OR3 (N2511, N2505, N1366, N2386);
buf BUF1 (N2512, N2507);
nor NOR3 (N2513, N2498, N2318, N713);
and AND2 (N2514, N2495, N1157);
xor XOR2 (N2515, N2509, N1659);
xor XOR2 (N2516, N2493, N879);
or OR4 (N2517, N2515, N1440, N1448, N1462);
or OR3 (N2518, N2510, N996, N1851);
nand NAND3 (N2519, N2516, N888, N2066);
nor NOR4 (N2520, N2517, N390, N2279, N1996);
nand NAND2 (N2521, N2519, N1977);
and AND2 (N2522, N2508, N2142);
buf BUF1 (N2523, N2518);
or OR3 (N2524, N2511, N2133, N241);
and AND2 (N2525, N2514, N885);
xor XOR2 (N2526, N2523, N1857);
xor XOR2 (N2527, N2521, N722);
not NOT1 (N2528, N2513);
nand NAND4 (N2529, N2487, N326, N2325, N923);
and AND2 (N2530, N2528, N628);
or OR3 (N2531, N2526, N1123, N519);
nand NAND2 (N2532, N2529, N2130);
xor XOR2 (N2533, N2520, N593);
buf BUF1 (N2534, N2533);
and AND3 (N2535, N2512, N2172, N1004);
or OR2 (N2536, N2534, N1398);
nand NAND4 (N2537, N2530, N1489, N2531, N1717);
or OR2 (N2538, N1020, N110);
or OR2 (N2539, N2538, N2065);
or OR3 (N2540, N2532, N141, N1343);
xor XOR2 (N2541, N2525, N1320);
buf BUF1 (N2542, N2536);
or OR4 (N2543, N2541, N1171, N1408, N1521);
and AND2 (N2544, N2539, N880);
buf BUF1 (N2545, N2537);
nand NAND3 (N2546, N2535, N521, N582);
xor XOR2 (N2547, N2540, N878);
nor NOR2 (N2548, N2543, N1908);
and AND2 (N2549, N2524, N1431);
not NOT1 (N2550, N2506);
or OR2 (N2551, N2547, N2538);
nor NOR2 (N2552, N2527, N2509);
nor NOR4 (N2553, N2549, N992, N749, N648);
and AND3 (N2554, N2553, N1381, N2193);
buf BUF1 (N2555, N2551);
nor NOR4 (N2556, N2554, N1827, N468, N421);
not NOT1 (N2557, N2548);
nor NOR2 (N2558, N2550, N103);
buf BUF1 (N2559, N2555);
nor NOR4 (N2560, N2558, N338, N253, N1007);
or OR3 (N2561, N2552, N1694, N198);
xor XOR2 (N2562, N2545, N413);
nand NAND4 (N2563, N2556, N1480, N1943, N2039);
not NOT1 (N2564, N2559);
nor NOR3 (N2565, N2561, N1778, N1765);
nor NOR4 (N2566, N2563, N97, N792, N1578);
not NOT1 (N2567, N2546);
nand NAND3 (N2568, N2565, N1003, N345);
nand NAND2 (N2569, N2568, N1549);
nand NAND2 (N2570, N2542, N1793);
not NOT1 (N2571, N2570);
and AND2 (N2572, N2571, N2389);
not NOT1 (N2573, N2557);
nand NAND4 (N2574, N2564, N702, N126, N1245);
xor XOR2 (N2575, N2566, N163);
nor NOR4 (N2576, N2560, N833, N2330, N61);
or OR3 (N2577, N2567, N1386, N111);
or OR3 (N2578, N2572, N301, N32);
nand NAND2 (N2579, N2578, N2083);
buf BUF1 (N2580, N2544);
nand NAND4 (N2581, N2522, N1345, N2314, N1304);
and AND2 (N2582, N2576, N2249);
or OR2 (N2583, N2569, N2200);
buf BUF1 (N2584, N2574);
xor XOR2 (N2585, N2573, N2263);
xor XOR2 (N2586, N2584, N1531);
buf BUF1 (N2587, N2575);
nor NOR4 (N2588, N2587, N1997, N1770, N1687);
buf BUF1 (N2589, N2583);
or OR2 (N2590, N2585, N508);
and AND4 (N2591, N2589, N437, N284, N1851);
xor XOR2 (N2592, N2591, N907);
or OR3 (N2593, N2588, N23, N406);
nand NAND2 (N2594, N2590, N768);
and AND2 (N2595, N2594, N1573);
not NOT1 (N2596, N2579);
xor XOR2 (N2597, N2580, N507);
and AND3 (N2598, N2592, N1131, N1141);
nor NOR4 (N2599, N2593, N1384, N958, N626);
nand NAND3 (N2600, N2581, N1578, N2046);
nand NAND3 (N2601, N2582, N1627, N168);
buf BUF1 (N2602, N2577);
nor NOR3 (N2603, N2599, N1016, N527);
not NOT1 (N2604, N2586);
xor XOR2 (N2605, N2597, N557);
nor NOR2 (N2606, N2595, N1932);
nand NAND3 (N2607, N2603, N784, N171);
nor NOR3 (N2608, N2600, N2014, N376);
or OR2 (N2609, N2608, N2425);
xor XOR2 (N2610, N2601, N274);
nor NOR2 (N2611, N2610, N1056);
nor NOR3 (N2612, N2602, N1467, N278);
buf BUF1 (N2613, N2605);
or OR3 (N2614, N2607, N1922, N30);
or OR2 (N2615, N2613, N1907);
nand NAND3 (N2616, N2611, N931, N670);
nand NAND3 (N2617, N2596, N862, N292);
xor XOR2 (N2618, N2612, N2179);
not NOT1 (N2619, N2598);
xor XOR2 (N2620, N2609, N237);
nor NOR4 (N2621, N2616, N279, N1286, N2081);
and AND3 (N2622, N2614, N365, N955);
not NOT1 (N2623, N2621);
and AND4 (N2624, N2622, N1671, N1495, N86);
xor XOR2 (N2625, N2619, N443);
nand NAND2 (N2626, N2617, N633);
nor NOR2 (N2627, N2623, N719);
xor XOR2 (N2628, N2627, N2063);
and AND2 (N2629, N2625, N1169);
not NOT1 (N2630, N2620);
not NOT1 (N2631, N2618);
not NOT1 (N2632, N2631);
or OR2 (N2633, N2630, N100);
nor NOR4 (N2634, N2604, N1508, N2529, N1812);
buf BUF1 (N2635, N2633);
nor NOR3 (N2636, N2606, N71, N946);
not NOT1 (N2637, N2562);
buf BUF1 (N2638, N2634);
nand NAND3 (N2639, N2629, N994, N1942);
nand NAND3 (N2640, N2626, N1229, N1523);
not NOT1 (N2641, N2635);
not NOT1 (N2642, N2615);
xor XOR2 (N2643, N2636, N911);
buf BUF1 (N2644, N2641);
not NOT1 (N2645, N2643);
not NOT1 (N2646, N2638);
and AND4 (N2647, N2642, N1560, N30, N1961);
not NOT1 (N2648, N2644);
xor XOR2 (N2649, N2640, N2001);
buf BUF1 (N2650, N2639);
not NOT1 (N2651, N2624);
buf BUF1 (N2652, N2628);
buf BUF1 (N2653, N2651);
xor XOR2 (N2654, N2652, N376);
not NOT1 (N2655, N2645);
or OR4 (N2656, N2655, N470, N1984, N332);
xor XOR2 (N2657, N2632, N2324);
nand NAND3 (N2658, N2653, N2331, N137);
nor NOR4 (N2659, N2648, N1708, N2489, N1365);
not NOT1 (N2660, N2654);
or OR2 (N2661, N2637, N2434);
or OR2 (N2662, N2660, N2253);
nor NOR4 (N2663, N2658, N2569, N2034, N2384);
or OR4 (N2664, N2649, N1250, N2548, N1324);
not NOT1 (N2665, N2646);
buf BUF1 (N2666, N2659);
xor XOR2 (N2667, N2666, N755);
nor NOR4 (N2668, N2665, N1762, N2054, N549);
nand NAND3 (N2669, N2657, N1605, N2616);
nand NAND3 (N2670, N2650, N2247, N1290);
or OR4 (N2671, N2647, N2635, N1598, N492);
and AND2 (N2672, N2663, N2293);
nand NAND4 (N2673, N2672, N2244, N338, N2331);
xor XOR2 (N2674, N2664, N2169);
not NOT1 (N2675, N2668);
nand NAND3 (N2676, N2673, N274, N2441);
buf BUF1 (N2677, N2656);
and AND3 (N2678, N2667, N1615, N2456);
xor XOR2 (N2679, N2669, N1174);
or OR3 (N2680, N2677, N2028, N2172);
nand NAND2 (N2681, N2675, N702);
xor XOR2 (N2682, N2679, N2581);
and AND3 (N2683, N2680, N2173, N847);
not NOT1 (N2684, N2683);
buf BUF1 (N2685, N2681);
not NOT1 (N2686, N2671);
and AND4 (N2687, N2676, N322, N141, N1026);
and AND2 (N2688, N2685, N2456);
buf BUF1 (N2689, N2688);
or OR2 (N2690, N2662, N467);
or OR3 (N2691, N2690, N120, N2402);
not NOT1 (N2692, N2670);
buf BUF1 (N2693, N2691);
buf BUF1 (N2694, N2689);
xor XOR2 (N2695, N2692, N1294);
and AND2 (N2696, N2674, N1411);
buf BUF1 (N2697, N2684);
nor NOR4 (N2698, N2686, N1554, N2066, N1151);
nor NOR2 (N2699, N2678, N388);
nand NAND4 (N2700, N2682, N238, N2078, N1705);
not NOT1 (N2701, N2700);
nor NOR3 (N2702, N2699, N204, N2494);
not NOT1 (N2703, N2702);
nand NAND3 (N2704, N2687, N2404, N219);
or OR4 (N2705, N2693, N2242, N866, N662);
buf BUF1 (N2706, N2695);
or OR4 (N2707, N2698, N510, N298, N771);
buf BUF1 (N2708, N2704);
nor NOR3 (N2709, N2705, N2372, N1789);
nor NOR4 (N2710, N2697, N934, N207, N2109);
or OR2 (N2711, N2694, N1125);
or OR2 (N2712, N2696, N2580);
and AND2 (N2713, N2709, N2698);
nand NAND4 (N2714, N2701, N899, N1064, N1400);
nor NOR3 (N2715, N2714, N980, N1909);
or OR2 (N2716, N2707, N86);
or OR3 (N2717, N2712, N2142, N2213);
nand NAND2 (N2718, N2703, N1663);
nor NOR2 (N2719, N2716, N706);
nand NAND4 (N2720, N2719, N1384, N1767, N895);
nor NOR2 (N2721, N2717, N1620);
nor NOR3 (N2722, N2715, N567, N1457);
or OR2 (N2723, N2710, N1872);
and AND4 (N2724, N2722, N1523, N887, N1202);
and AND4 (N2725, N2713, N1500, N449, N1458);
nor NOR3 (N2726, N2708, N2060, N1500);
or OR4 (N2727, N2724, N1846, N310, N1270);
nand NAND2 (N2728, N2720, N17);
nor NOR2 (N2729, N2711, N2359);
nand NAND4 (N2730, N2729, N532, N2078, N795);
xor XOR2 (N2731, N2727, N1382);
or OR4 (N2732, N2725, N2699, N210, N1603);
and AND3 (N2733, N2723, N1416, N984);
xor XOR2 (N2734, N2718, N319);
xor XOR2 (N2735, N2726, N402);
buf BUF1 (N2736, N2730);
not NOT1 (N2737, N2721);
xor XOR2 (N2738, N2734, N1000);
nand NAND4 (N2739, N2736, N1664, N1844, N127);
nand NAND4 (N2740, N2737, N1347, N2345, N498);
buf BUF1 (N2741, N2731);
not NOT1 (N2742, N2661);
xor XOR2 (N2743, N2728, N475);
not NOT1 (N2744, N2738);
buf BUF1 (N2745, N2740);
xor XOR2 (N2746, N2741, N146);
not NOT1 (N2747, N2746);
buf BUF1 (N2748, N2742);
and AND3 (N2749, N2733, N2577, N1444);
or OR4 (N2750, N2749, N1410, N1883, N1932);
nor NOR3 (N2751, N2706, N919, N2177);
and AND3 (N2752, N2732, N642, N2622);
xor XOR2 (N2753, N2750, N342);
buf BUF1 (N2754, N2735);
nand NAND4 (N2755, N2747, N2320, N2561, N1730);
or OR2 (N2756, N2755, N1548);
or OR4 (N2757, N2754, N1105, N172, N817);
and AND4 (N2758, N2739, N1081, N2168, N175);
or OR2 (N2759, N2748, N2540);
nand NAND4 (N2760, N2743, N101, N258, N1100);
buf BUF1 (N2761, N2753);
or OR4 (N2762, N2756, N688, N1182, N433);
nor NOR4 (N2763, N2762, N1787, N841, N945);
or OR3 (N2764, N2760, N2668, N1495);
buf BUF1 (N2765, N2763);
xor XOR2 (N2766, N2757, N150);
buf BUF1 (N2767, N2752);
buf BUF1 (N2768, N2767);
nor NOR3 (N2769, N2745, N2654, N2426);
xor XOR2 (N2770, N2761, N531);
nand NAND4 (N2771, N2758, N2292, N2441, N1431);
nor NOR2 (N2772, N2764, N487);
and AND4 (N2773, N2768, N471, N883, N963);
or OR4 (N2774, N2772, N91, N673, N2080);
buf BUF1 (N2775, N2771);
nor NOR2 (N2776, N2775, N1947);
xor XOR2 (N2777, N2766, N1529);
and AND2 (N2778, N2777, N394);
and AND2 (N2779, N2744, N2299);
nor NOR2 (N2780, N2769, N308);
or OR3 (N2781, N2759, N966, N627);
nand NAND2 (N2782, N2779, N1565);
not NOT1 (N2783, N2765);
nor NOR4 (N2784, N2773, N2624, N1733, N153);
buf BUF1 (N2785, N2782);
buf BUF1 (N2786, N2774);
xor XOR2 (N2787, N2770, N876);
nand NAND2 (N2788, N2776, N2476);
nor NOR3 (N2789, N2787, N2101, N449);
nor NOR4 (N2790, N2789, N2461, N2017, N362);
and AND4 (N2791, N2790, N2670, N799, N1198);
nor NOR3 (N2792, N2785, N2760, N944);
and AND4 (N2793, N2751, N2119, N461, N2350);
not NOT1 (N2794, N2786);
or OR4 (N2795, N2778, N2709, N1266, N1607);
buf BUF1 (N2796, N2781);
nand NAND4 (N2797, N2793, N2546, N1244, N597);
nor NOR3 (N2798, N2795, N503, N422);
or OR3 (N2799, N2792, N1646, N2644);
buf BUF1 (N2800, N2780);
and AND4 (N2801, N2797, N114, N486, N1173);
not NOT1 (N2802, N2800);
buf BUF1 (N2803, N2791);
or OR3 (N2804, N2794, N78, N817);
not NOT1 (N2805, N2803);
nor NOR3 (N2806, N2788, N2619, N5);
nor NOR4 (N2807, N2796, N590, N2464, N765);
buf BUF1 (N2808, N2799);
nand NAND2 (N2809, N2806, N1968);
nor NOR4 (N2810, N2807, N1620, N2249, N2287);
and AND3 (N2811, N2798, N2254, N2082);
buf BUF1 (N2812, N2809);
xor XOR2 (N2813, N2784, N378);
nor NOR4 (N2814, N2805, N2283, N2652, N113);
and AND4 (N2815, N2801, N2092, N299, N2453);
and AND3 (N2816, N2813, N1179, N1928);
or OR3 (N2817, N2815, N1566, N980);
nand NAND2 (N2818, N2812, N1883);
and AND3 (N2819, N2814, N391, N150);
xor XOR2 (N2820, N2819, N124);
nor NOR3 (N2821, N2820, N513, N2481);
xor XOR2 (N2822, N2821, N121);
buf BUF1 (N2823, N2816);
nand NAND3 (N2824, N2783, N639, N1369);
nand NAND2 (N2825, N2818, N292);
not NOT1 (N2826, N2824);
nand NAND2 (N2827, N2822, N249);
nor NOR2 (N2828, N2810, N2233);
nor NOR2 (N2829, N2804, N2462);
xor XOR2 (N2830, N2823, N2714);
xor XOR2 (N2831, N2825, N1419);
nand NAND4 (N2832, N2829, N2760, N937, N1141);
not NOT1 (N2833, N2811);
nor NOR2 (N2834, N2831, N1748);
xor XOR2 (N2835, N2833, N2067);
not NOT1 (N2836, N2802);
and AND3 (N2837, N2828, N749, N1956);
not NOT1 (N2838, N2830);
buf BUF1 (N2839, N2836);
buf BUF1 (N2840, N2839);
buf BUF1 (N2841, N2838);
buf BUF1 (N2842, N2826);
or OR2 (N2843, N2832, N1525);
buf BUF1 (N2844, N2841);
buf BUF1 (N2845, N2842);
and AND2 (N2846, N2808, N122);
nor NOR3 (N2847, N2827, N664, N2725);
or OR3 (N2848, N2837, N1723, N2273);
nand NAND4 (N2849, N2843, N1373, N2690, N1486);
nor NOR4 (N2850, N2840, N1916, N306, N2334);
nand NAND4 (N2851, N2845, N1184, N875, N296);
or OR2 (N2852, N2835, N221);
nand NAND2 (N2853, N2851, N1843);
buf BUF1 (N2854, N2853);
not NOT1 (N2855, N2848);
xor XOR2 (N2856, N2834, N2728);
buf BUF1 (N2857, N2850);
and AND4 (N2858, N2857, N897, N1538, N1085);
not NOT1 (N2859, N2852);
nor NOR2 (N2860, N2859, N1445);
and AND3 (N2861, N2844, N727, N1490);
not NOT1 (N2862, N2847);
buf BUF1 (N2863, N2854);
buf BUF1 (N2864, N2860);
buf BUF1 (N2865, N2863);
nand NAND4 (N2866, N2861, N2847, N1481, N1913);
not NOT1 (N2867, N2866);
nor NOR2 (N2868, N2856, N313);
buf BUF1 (N2869, N2864);
nor NOR3 (N2870, N2862, N1425, N1278);
nand NAND2 (N2871, N2817, N1744);
buf BUF1 (N2872, N2870);
nor NOR2 (N2873, N2868, N853);
not NOT1 (N2874, N2869);
xor XOR2 (N2875, N2858, N1784);
not NOT1 (N2876, N2871);
and AND4 (N2877, N2867, N2305, N1037, N2394);
and AND2 (N2878, N2873, N1739);
and AND2 (N2879, N2874, N1578);
not NOT1 (N2880, N2875);
buf BUF1 (N2881, N2849);
xor XOR2 (N2882, N2876, N1877);
nand NAND4 (N2883, N2865, N422, N1549, N2029);
xor XOR2 (N2884, N2879, N157);
or OR3 (N2885, N2878, N692, N19);
buf BUF1 (N2886, N2881);
not NOT1 (N2887, N2872);
nand NAND3 (N2888, N2883, N895, N2480);
xor XOR2 (N2889, N2846, N1279);
nand NAND4 (N2890, N2886, N2781, N927, N1200);
xor XOR2 (N2891, N2884, N2101);
buf BUF1 (N2892, N2887);
not NOT1 (N2893, N2877);
nor NOR2 (N2894, N2888, N1022);
nand NAND4 (N2895, N2880, N2554, N1535, N2028);
or OR2 (N2896, N2885, N1073);
nor NOR4 (N2897, N2896, N1916, N2341, N1338);
or OR4 (N2898, N2890, N1060, N1660, N29);
buf BUF1 (N2899, N2897);
not NOT1 (N2900, N2892);
xor XOR2 (N2901, N2898, N603);
not NOT1 (N2902, N2889);
xor XOR2 (N2903, N2901, N277);
nor NOR2 (N2904, N2894, N1935);
and AND4 (N2905, N2895, N2559, N1158, N2031);
not NOT1 (N2906, N2905);
not NOT1 (N2907, N2904);
and AND3 (N2908, N2900, N1431, N170);
buf BUF1 (N2909, N2906);
buf BUF1 (N2910, N2908);
not NOT1 (N2911, N2882);
or OR4 (N2912, N2893, N2664, N1077, N2709);
nand NAND3 (N2913, N2911, N1384, N2507);
and AND3 (N2914, N2891, N2544, N1115);
or OR2 (N2915, N2913, N2182);
and AND3 (N2916, N2902, N399, N425);
and AND4 (N2917, N2912, N691, N2340, N2913);
nand NAND2 (N2918, N2910, N2809);
nor NOR3 (N2919, N2915, N1124, N1250);
buf BUF1 (N2920, N2855);
or OR4 (N2921, N2916, N1899, N1394, N262);
xor XOR2 (N2922, N2918, N1412);
xor XOR2 (N2923, N2907, N178);
not NOT1 (N2924, N2922);
not NOT1 (N2925, N2921);
nor NOR2 (N2926, N2925, N2193);
or OR3 (N2927, N2923, N835, N2096);
not NOT1 (N2928, N2926);
buf BUF1 (N2929, N2924);
nor NOR4 (N2930, N2909, N2127, N2819, N216);
or OR2 (N2931, N2927, N2756);
and AND3 (N2932, N2903, N624, N2438);
nor NOR4 (N2933, N2932, N2051, N570, N1973);
nand NAND4 (N2934, N2919, N2314, N2580, N1920);
nor NOR3 (N2935, N2929, N582, N1998);
buf BUF1 (N2936, N2934);
xor XOR2 (N2937, N2917, N1984);
and AND3 (N2938, N2920, N176, N2181);
not NOT1 (N2939, N2936);
not NOT1 (N2940, N2935);
or OR4 (N2941, N2933, N334, N833, N2212);
nand NAND2 (N2942, N2939, N1285);
buf BUF1 (N2943, N2899);
xor XOR2 (N2944, N2937, N2818);
or OR3 (N2945, N2943, N1043, N85);
or OR3 (N2946, N2942, N541, N1915);
not NOT1 (N2947, N2928);
xor XOR2 (N2948, N2945, N2406);
nor NOR2 (N2949, N2940, N963);
nor NOR4 (N2950, N2947, N1992, N954, N1794);
and AND3 (N2951, N2914, N1579, N2581);
nor NOR3 (N2952, N2938, N2899, N2231);
nor NOR4 (N2953, N2931, N1516, N361, N1617);
not NOT1 (N2954, N2944);
nor NOR3 (N2955, N2949, N2569, N1955);
not NOT1 (N2956, N2951);
or OR3 (N2957, N2930, N617, N876);
xor XOR2 (N2958, N2946, N2592);
nor NOR3 (N2959, N2941, N2539, N882);
buf BUF1 (N2960, N2953);
not NOT1 (N2961, N2948);
nor NOR4 (N2962, N2960, N879, N1284, N955);
or OR2 (N2963, N2959, N930);
not NOT1 (N2964, N2957);
buf BUF1 (N2965, N2950);
or OR2 (N2966, N2952, N135);
or OR2 (N2967, N2954, N2687);
nor NOR3 (N2968, N2958, N1140, N844);
nor NOR2 (N2969, N2966, N2088);
xor XOR2 (N2970, N2964, N1643);
xor XOR2 (N2971, N2968, N452);
and AND2 (N2972, N2962, N2502);
and AND4 (N2973, N2971, N792, N87, N265);
xor XOR2 (N2974, N2963, N1234);
buf BUF1 (N2975, N2972);
xor XOR2 (N2976, N2955, N1868);
nor NOR3 (N2977, N2969, N1647, N2114);
nor NOR3 (N2978, N2965, N415, N2453);
nand NAND2 (N2979, N2967, N1732);
nor NOR2 (N2980, N2975, N2391);
nand NAND2 (N2981, N2970, N2761);
buf BUF1 (N2982, N2961);
nand NAND2 (N2983, N2979, N2065);
nor NOR3 (N2984, N2978, N2047, N683);
not NOT1 (N2985, N2983);
xor XOR2 (N2986, N2980, N33);
not NOT1 (N2987, N2977);
or OR2 (N2988, N2981, N318);
buf BUF1 (N2989, N2988);
nor NOR2 (N2990, N2985, N2742);
buf BUF1 (N2991, N2986);
not NOT1 (N2992, N2984);
nand NAND2 (N2993, N2990, N1557);
or OR4 (N2994, N2973, N1987, N142, N2536);
nand NAND3 (N2995, N2992, N2911, N1640);
or OR3 (N2996, N2982, N1159, N1992);
nor NOR4 (N2997, N2991, N1634, N490, N556);
or OR2 (N2998, N2994, N2314);
buf BUF1 (N2999, N2996);
nor NOR3 (N3000, N2976, N2841, N1990);
nor NOR2 (N3001, N2974, N1856);
nand NAND4 (N3002, N2998, N1383, N2386, N2416);
nand NAND3 (N3003, N2997, N1636, N50);
not NOT1 (N3004, N2987);
buf BUF1 (N3005, N2993);
and AND4 (N3006, N3005, N2881, N60, N2020);
nand NAND3 (N3007, N3006, N1963, N2255);
buf BUF1 (N3008, N2956);
or OR3 (N3009, N3000, N1384, N16);
or OR3 (N3010, N3004, N1712, N1236);
and AND2 (N3011, N3009, N750);
and AND3 (N3012, N3007, N2301, N2036);
buf BUF1 (N3013, N3010);
buf BUF1 (N3014, N3003);
xor XOR2 (N3015, N2995, N419);
and AND3 (N3016, N3013, N374, N1826);
not NOT1 (N3017, N3001);
xor XOR2 (N3018, N3008, N2103);
xor XOR2 (N3019, N3002, N1761);
nor NOR4 (N3020, N3015, N1745, N228, N1224);
xor XOR2 (N3021, N2999, N1851);
nand NAND2 (N3022, N3012, N1225);
nor NOR2 (N3023, N2989, N59);
nor NOR3 (N3024, N3021, N2589, N2560);
xor XOR2 (N3025, N3018, N2207);
not NOT1 (N3026, N3011);
nand NAND3 (N3027, N3014, N100, N2443);
nand NAND2 (N3028, N3016, N1966);
nand NAND2 (N3029, N3024, N1719);
nand NAND2 (N3030, N3022, N2628);
not NOT1 (N3031, N3025);
nor NOR4 (N3032, N3028, N2129, N1025, N2320);
nand NAND3 (N3033, N3031, N195, N1458);
not NOT1 (N3034, N3029);
nand NAND4 (N3035, N3023, N1618, N1170, N2459);
and AND3 (N3036, N3020, N526, N442);
and AND3 (N3037, N3030, N362, N1750);
nor NOR4 (N3038, N3026, N1522, N1406, N717);
xor XOR2 (N3039, N3019, N1908);
nor NOR2 (N3040, N3017, N2018);
buf BUF1 (N3041, N3027);
nor NOR3 (N3042, N3037, N1857, N1507);
nand NAND2 (N3043, N3035, N2578);
nor NOR2 (N3044, N3042, N38);
or OR2 (N3045, N3032, N2375);
xor XOR2 (N3046, N3033, N1981);
buf BUF1 (N3047, N3034);
xor XOR2 (N3048, N3046, N2839);
nor NOR2 (N3049, N3044, N456);
buf BUF1 (N3050, N3049);
buf BUF1 (N3051, N3050);
xor XOR2 (N3052, N3036, N1798);
or OR4 (N3053, N3039, N2275, N2674, N2804);
xor XOR2 (N3054, N3043, N1580);
nor NOR3 (N3055, N3054, N740, N1081);
nand NAND2 (N3056, N3041, N2065);
nand NAND3 (N3057, N3051, N1520, N1638);
and AND4 (N3058, N3057, N1872, N2914, N2467);
nor NOR4 (N3059, N3053, N3056, N1771, N1773);
xor XOR2 (N3060, N1755, N1128);
nor NOR4 (N3061, N3060, N1296, N2345, N1614);
xor XOR2 (N3062, N3058, N757);
xor XOR2 (N3063, N3061, N2690);
not NOT1 (N3064, N3055);
buf BUF1 (N3065, N3047);
or OR2 (N3066, N3059, N1156);
buf BUF1 (N3067, N3064);
nor NOR3 (N3068, N3066, N2747, N175);
xor XOR2 (N3069, N3052, N1108);
and AND2 (N3070, N3062, N2144);
and AND2 (N3071, N3048, N2820);
or OR4 (N3072, N3068, N2988, N36, N899);
nand NAND2 (N3073, N3065, N1464);
xor XOR2 (N3074, N3040, N2064);
nor NOR2 (N3075, N3069, N603);
nand NAND3 (N3076, N3038, N1992, N725);
xor XOR2 (N3077, N3074, N2399);
or OR4 (N3078, N3072, N1861, N1187, N249);
not NOT1 (N3079, N3077);
nand NAND3 (N3080, N3045, N1904, N1141);
xor XOR2 (N3081, N3070, N2610);
xor XOR2 (N3082, N3080, N2141);
buf BUF1 (N3083, N3075);
not NOT1 (N3084, N3083);
and AND4 (N3085, N3079, N2728, N1260, N1516);
and AND2 (N3086, N3063, N2736);
buf BUF1 (N3087, N3067);
xor XOR2 (N3088, N3084, N1673);
not NOT1 (N3089, N3085);
xor XOR2 (N3090, N3089, N1501);
and AND2 (N3091, N3082, N2675);
buf BUF1 (N3092, N3090);
nand NAND4 (N3093, N3076, N114, N1317, N1928);
nand NAND2 (N3094, N3071, N298);
and AND3 (N3095, N3073, N599, N926);
and AND2 (N3096, N3094, N2586);
nand NAND2 (N3097, N3081, N2128);
or OR4 (N3098, N3093, N1335, N993, N551);
not NOT1 (N3099, N3088);
buf BUF1 (N3100, N3087);
buf BUF1 (N3101, N3078);
or OR2 (N3102, N3091, N1222);
not NOT1 (N3103, N3095);
and AND2 (N3104, N3102, N2645);
nor NOR4 (N3105, N3099, N59, N519, N2500);
or OR3 (N3106, N3105, N2260, N1546);
not NOT1 (N3107, N3100);
or OR3 (N3108, N3098, N2823, N1466);
or OR3 (N3109, N3107, N2600, N411);
nand NAND3 (N3110, N3092, N2735, N1477);
not NOT1 (N3111, N3104);
or OR2 (N3112, N3108, N2840);
xor XOR2 (N3113, N3101, N181);
or OR4 (N3114, N3109, N2293, N2978, N692);
or OR4 (N3115, N3106, N572, N1499, N2830);
buf BUF1 (N3116, N3096);
xor XOR2 (N3117, N3112, N1382);
not NOT1 (N3118, N3111);
nand NAND4 (N3119, N3103, N1358, N1836, N2621);
xor XOR2 (N3120, N3116, N2935);
and AND2 (N3121, N3117, N1504);
and AND3 (N3122, N3121, N733, N3093);
not NOT1 (N3123, N3097);
xor XOR2 (N3124, N3119, N2565);
and AND2 (N3125, N3113, N2258);
buf BUF1 (N3126, N3086);
or OR3 (N3127, N3114, N1791, N622);
nor NOR2 (N3128, N3110, N2434);
nor NOR4 (N3129, N3128, N1776, N822, N1064);
nor NOR2 (N3130, N3120, N1656);
nand NAND2 (N3131, N3127, N1148);
not NOT1 (N3132, N3126);
nand NAND4 (N3133, N3115, N2849, N2862, N2697);
xor XOR2 (N3134, N3129, N1638);
buf BUF1 (N3135, N3118);
or OR2 (N3136, N3135, N608);
xor XOR2 (N3137, N3122, N2641);
nor NOR2 (N3138, N3137, N370);
not NOT1 (N3139, N3132);
not NOT1 (N3140, N3125);
buf BUF1 (N3141, N3139);
nor NOR3 (N3142, N3123, N3011, N3064);
nor NOR4 (N3143, N3136, N1117, N2745, N935);
and AND4 (N3144, N3131, N1409, N377, N228);
or OR4 (N3145, N3141, N1068, N128, N318);
xor XOR2 (N3146, N3130, N1579);
or OR4 (N3147, N3142, N1421, N2509, N648);
xor XOR2 (N3148, N3133, N492);
or OR4 (N3149, N3134, N1314, N2176, N1042);
not NOT1 (N3150, N3145);
nor NOR4 (N3151, N3138, N316, N474, N700);
or OR2 (N3152, N3144, N1613);
not NOT1 (N3153, N3146);
not NOT1 (N3154, N3124);
or OR3 (N3155, N3140, N1201, N1427);
not NOT1 (N3156, N3147);
buf BUF1 (N3157, N3151);
nand NAND2 (N3158, N3156, N92);
xor XOR2 (N3159, N3149, N479);
or OR2 (N3160, N3157, N1252);
nand NAND2 (N3161, N3152, N2911);
xor XOR2 (N3162, N3143, N1937);
or OR4 (N3163, N3162, N269, N2961, N3070);
and AND3 (N3164, N3159, N3141, N2529);
and AND2 (N3165, N3164, N899);
or OR3 (N3166, N3161, N1436, N1345);
xor XOR2 (N3167, N3153, N2560);
nand NAND2 (N3168, N3167, N1138);
nand NAND3 (N3169, N3168, N2259, N80);
not NOT1 (N3170, N3155);
not NOT1 (N3171, N3169);
nand NAND4 (N3172, N3154, N3016, N1259, N2359);
nor NOR3 (N3173, N3171, N623, N1313);
xor XOR2 (N3174, N3172, N1514);
nor NOR2 (N3175, N3173, N1776);
nor NOR3 (N3176, N3165, N1543, N2154);
and AND2 (N3177, N3174, N1148);
not NOT1 (N3178, N3170);
buf BUF1 (N3179, N3166);
or OR4 (N3180, N3177, N2129, N157, N1027);
or OR3 (N3181, N3175, N195, N1618);
xor XOR2 (N3182, N3181, N1043);
and AND2 (N3183, N3150, N1959);
xor XOR2 (N3184, N3158, N2590);
xor XOR2 (N3185, N3176, N2558);
not NOT1 (N3186, N3184);
not NOT1 (N3187, N3178);
nand NAND3 (N3188, N3186, N2685, N3141);
buf BUF1 (N3189, N3160);
buf BUF1 (N3190, N3180);
nand NAND4 (N3191, N3188, N3016, N2355, N332);
nand NAND2 (N3192, N3189, N1953);
or OR3 (N3193, N3191, N2332, N1128);
and AND4 (N3194, N3179, N791, N1916, N2926);
nand NAND4 (N3195, N3183, N2524, N2369, N2384);
xor XOR2 (N3196, N3190, N1298);
or OR4 (N3197, N3193, N2326, N2115, N2076);
and AND3 (N3198, N3197, N1249, N1071);
buf BUF1 (N3199, N3194);
not NOT1 (N3200, N3192);
not NOT1 (N3201, N3196);
nor NOR4 (N3202, N3182, N2008, N2030, N1648);
not NOT1 (N3203, N3198);
nand NAND2 (N3204, N3195, N1282);
nand NAND2 (N3205, N3163, N373);
nor NOR4 (N3206, N3201, N1603, N968, N797);
buf BUF1 (N3207, N3148);
nand NAND2 (N3208, N3199, N2476);
nor NOR3 (N3209, N3203, N1919, N902);
xor XOR2 (N3210, N3205, N1936);
nand NAND4 (N3211, N3208, N312, N1369, N828);
buf BUF1 (N3212, N3206);
buf BUF1 (N3213, N3185);
or OR4 (N3214, N3209, N949, N3045, N2429);
or OR2 (N3215, N3214, N1829);
or OR2 (N3216, N3200, N2582);
nand NAND4 (N3217, N3204, N675, N2034, N1593);
not NOT1 (N3218, N3207);
buf BUF1 (N3219, N3211);
nor NOR4 (N3220, N3216, N389, N537, N1773);
nand NAND4 (N3221, N3217, N3064, N1761, N2658);
and AND2 (N3222, N3221, N214);
or OR3 (N3223, N3219, N1265, N2753);
and AND3 (N3224, N3223, N348, N900);
or OR3 (N3225, N3210, N1112, N2618);
not NOT1 (N3226, N3187);
and AND3 (N3227, N3224, N1361, N1066);
or OR2 (N3228, N3225, N1156);
buf BUF1 (N3229, N3222);
or OR2 (N3230, N3202, N243);
nor NOR2 (N3231, N3218, N2544);
nand NAND3 (N3232, N3226, N2209, N2309);
or OR2 (N3233, N3232, N36);
buf BUF1 (N3234, N3229);
and AND3 (N3235, N3234, N2162, N11);
or OR3 (N3236, N3228, N1835, N242);
or OR2 (N3237, N3231, N2490);
buf BUF1 (N3238, N3220);
not NOT1 (N3239, N3215);
and AND2 (N3240, N3236, N123);
xor XOR2 (N3241, N3238, N482);
or OR3 (N3242, N3233, N1070, N1404);
buf BUF1 (N3243, N3237);
nor NOR4 (N3244, N3243, N2286, N1577, N746);
nand NAND2 (N3245, N3235, N868);
buf BUF1 (N3246, N3227);
not NOT1 (N3247, N3213);
and AND2 (N3248, N3239, N2414);
nand NAND4 (N3249, N3245, N772, N421, N813);
nor NOR4 (N3250, N3212, N1220, N3131, N2569);
xor XOR2 (N3251, N3244, N1982);
buf BUF1 (N3252, N3240);
xor XOR2 (N3253, N3246, N1794);
xor XOR2 (N3254, N3249, N1491);
nor NOR2 (N3255, N3252, N529);
buf BUF1 (N3256, N3241);
not NOT1 (N3257, N3230);
xor XOR2 (N3258, N3242, N371);
not NOT1 (N3259, N3251);
and AND4 (N3260, N3257, N28, N507, N1958);
not NOT1 (N3261, N3248);
nor NOR2 (N3262, N3259, N319);
xor XOR2 (N3263, N3247, N71);
or OR3 (N3264, N3250, N3131, N2396);
nand NAND2 (N3265, N3260, N977);
not NOT1 (N3266, N3265);
nand NAND2 (N3267, N3261, N1368);
buf BUF1 (N3268, N3256);
nor NOR2 (N3269, N3255, N895);
xor XOR2 (N3270, N3263, N1157);
nand NAND2 (N3271, N3269, N448);
not NOT1 (N3272, N3267);
buf BUF1 (N3273, N3266);
or OR3 (N3274, N3254, N2039, N1992);
and AND4 (N3275, N3258, N1722, N1675, N2033);
xor XOR2 (N3276, N3272, N3050);
nor NOR3 (N3277, N3270, N1755, N885);
not NOT1 (N3278, N3264);
xor XOR2 (N3279, N3262, N321);
nor NOR3 (N3280, N3268, N1301, N1842);
buf BUF1 (N3281, N3277);
xor XOR2 (N3282, N3274, N1313);
nor NOR3 (N3283, N3281, N908, N2180);
nand NAND3 (N3284, N3276, N1509, N3178);
not NOT1 (N3285, N3282);
xor XOR2 (N3286, N3285, N2906);
buf BUF1 (N3287, N3275);
xor XOR2 (N3288, N3271, N6);
buf BUF1 (N3289, N3288);
buf BUF1 (N3290, N3278);
xor XOR2 (N3291, N3283, N2523);
or OR3 (N3292, N3279, N1186, N1985);
xor XOR2 (N3293, N3292, N2080);
and AND4 (N3294, N3253, N2327, N2513, N2211);
not NOT1 (N3295, N3293);
buf BUF1 (N3296, N3290);
buf BUF1 (N3297, N3286);
xor XOR2 (N3298, N3295, N489);
and AND4 (N3299, N3284, N915, N1625, N678);
not NOT1 (N3300, N3273);
nand NAND4 (N3301, N3298, N3099, N1094, N1021);
buf BUF1 (N3302, N3300);
and AND2 (N3303, N3297, N2920);
nand NAND3 (N3304, N3303, N62, N143);
not NOT1 (N3305, N3302);
and AND2 (N3306, N3291, N2782);
nor NOR2 (N3307, N3299, N157);
nor NOR3 (N3308, N3289, N631, N2229);
or OR2 (N3309, N3306, N1005);
or OR3 (N3310, N3309, N838, N2298);
and AND3 (N3311, N3304, N1080, N1418);
not NOT1 (N3312, N3305);
xor XOR2 (N3313, N3280, N80);
xor XOR2 (N3314, N3287, N2771);
nor NOR3 (N3315, N3311, N1074, N2829);
and AND3 (N3316, N3301, N1077, N146);
and AND3 (N3317, N3315, N1893, N2252);
buf BUF1 (N3318, N3294);
not NOT1 (N3319, N3314);
nor NOR2 (N3320, N3310, N2899);
nor NOR3 (N3321, N3320, N323, N1138);
and AND2 (N3322, N3308, N1384);
nor NOR3 (N3323, N3322, N2637, N1055);
nand NAND4 (N3324, N3316, N1344, N2362, N1771);
not NOT1 (N3325, N3296);
and AND2 (N3326, N3319, N3032);
xor XOR2 (N3327, N3317, N1464);
nor NOR4 (N3328, N3323, N3263, N2614, N1497);
nor NOR4 (N3329, N3324, N71, N1714, N1939);
or OR4 (N3330, N3321, N1130, N503, N1020);
and AND2 (N3331, N3325, N1717);
xor XOR2 (N3332, N3318, N2732);
nor NOR4 (N3333, N3332, N645, N2016, N2732);
buf BUF1 (N3334, N3312);
nand NAND2 (N3335, N3330, N303);
nand NAND4 (N3336, N3307, N2599, N1086, N2417);
nor NOR4 (N3337, N3326, N858, N1140, N932);
not NOT1 (N3338, N3329);
or OR2 (N3339, N3313, N2204);
not NOT1 (N3340, N3339);
xor XOR2 (N3341, N3327, N725);
not NOT1 (N3342, N3328);
xor XOR2 (N3343, N3341, N2612);
xor XOR2 (N3344, N3338, N2231);
nand NAND2 (N3345, N3336, N2859);
not NOT1 (N3346, N3333);
buf BUF1 (N3347, N3337);
nand NAND3 (N3348, N3334, N870, N2926);
nor NOR3 (N3349, N3331, N1138, N869);
xor XOR2 (N3350, N3348, N2233);
nor NOR3 (N3351, N3342, N282, N138);
nor NOR2 (N3352, N3343, N1285);
xor XOR2 (N3353, N3335, N2471);
or OR3 (N3354, N3346, N629, N874);
not NOT1 (N3355, N3354);
or OR4 (N3356, N3352, N90, N1878, N1269);
xor XOR2 (N3357, N3350, N253);
not NOT1 (N3358, N3347);
and AND4 (N3359, N3357, N45, N1062, N1936);
xor XOR2 (N3360, N3356, N791);
and AND2 (N3361, N3351, N2935);
and AND4 (N3362, N3355, N1093, N1285, N1413);
and AND2 (N3363, N3344, N1521);
nand NAND3 (N3364, N3362, N2324, N1700);
buf BUF1 (N3365, N3345);
nand NAND3 (N3366, N3340, N493, N2862);
nor NOR4 (N3367, N3349, N2597, N723, N3308);
xor XOR2 (N3368, N3364, N3264);
or OR2 (N3369, N3367, N1289);
buf BUF1 (N3370, N3358);
buf BUF1 (N3371, N3359);
nor NOR4 (N3372, N3360, N499, N3063, N451);
or OR4 (N3373, N3361, N934, N3236, N382);
buf BUF1 (N3374, N3369);
or OR2 (N3375, N3363, N282);
xor XOR2 (N3376, N3353, N1805);
and AND3 (N3377, N3370, N1795, N1659);
buf BUF1 (N3378, N3377);
not NOT1 (N3379, N3368);
or OR2 (N3380, N3374, N2709);
xor XOR2 (N3381, N3376, N1865);
xor XOR2 (N3382, N3372, N903);
nor NOR2 (N3383, N3382, N3367);
or OR2 (N3384, N3378, N788);
and AND2 (N3385, N3384, N3282);
xor XOR2 (N3386, N3375, N691);
nand NAND4 (N3387, N3373, N3232, N2857, N3166);
and AND4 (N3388, N3371, N1983, N1782, N891);
and AND4 (N3389, N3365, N2647, N2128, N1872);
not NOT1 (N3390, N3389);
buf BUF1 (N3391, N3385);
or OR4 (N3392, N3383, N214, N2899, N1633);
not NOT1 (N3393, N3366);
xor XOR2 (N3394, N3391, N3108);
xor XOR2 (N3395, N3387, N39);
and AND4 (N3396, N3388, N1297, N2150, N446);
buf BUF1 (N3397, N3390);
and AND2 (N3398, N3380, N2908);
not NOT1 (N3399, N3398);
not NOT1 (N3400, N3399);
and AND4 (N3401, N3394, N1939, N780, N1520);
nand NAND3 (N3402, N3392, N2301, N1510);
and AND4 (N3403, N3397, N2559, N2486, N2378);
nand NAND4 (N3404, N3395, N2396, N35, N968);
nor NOR3 (N3405, N3396, N481, N547);
and AND3 (N3406, N3404, N2702, N977);
nand NAND3 (N3407, N3400, N85, N1261);
xor XOR2 (N3408, N3407, N2379);
not NOT1 (N3409, N3393);
nand NAND3 (N3410, N3402, N458, N1314);
and AND2 (N3411, N3379, N3010);
not NOT1 (N3412, N3405);
and AND4 (N3413, N3406, N3138, N911, N250);
nand NAND4 (N3414, N3409, N225, N1385, N2651);
buf BUF1 (N3415, N3414);
and AND2 (N3416, N3386, N1916);
not NOT1 (N3417, N3401);
buf BUF1 (N3418, N3411);
xor XOR2 (N3419, N3403, N2438);
nor NOR2 (N3420, N3412, N1883);
xor XOR2 (N3421, N3419, N1988);
nand NAND3 (N3422, N3410, N1562, N2345);
xor XOR2 (N3423, N3416, N1670);
or OR2 (N3424, N3418, N3042);
xor XOR2 (N3425, N3381, N2300);
nor NOR4 (N3426, N3422, N1429, N969, N1985);
xor XOR2 (N3427, N3415, N240);
xor XOR2 (N3428, N3423, N1325);
xor XOR2 (N3429, N3424, N1384);
and AND4 (N3430, N3420, N2509, N3389, N1455);
not NOT1 (N3431, N3421);
not NOT1 (N3432, N3426);
not NOT1 (N3433, N3417);
nand NAND4 (N3434, N3408, N927, N2078, N1403);
not NOT1 (N3435, N3427);
nor NOR4 (N3436, N3432, N2180, N2147, N2120);
xor XOR2 (N3437, N3430, N486);
or OR2 (N3438, N3437, N2401);
buf BUF1 (N3439, N3438);
and AND2 (N3440, N3436, N199);
xor XOR2 (N3441, N3425, N738);
or OR2 (N3442, N3439, N1309);
not NOT1 (N3443, N3441);
buf BUF1 (N3444, N3429);
and AND2 (N3445, N3444, N1816);
or OR4 (N3446, N3435, N2296, N1138, N3237);
or OR2 (N3447, N3433, N789);
nand NAND2 (N3448, N3442, N965);
xor XOR2 (N3449, N3413, N529);
nor NOR2 (N3450, N3428, N2787);
nor NOR2 (N3451, N3446, N1043);
buf BUF1 (N3452, N3450);
and AND4 (N3453, N3447, N584, N617, N1800);
nand NAND2 (N3454, N3445, N1307);
nor NOR4 (N3455, N3451, N3068, N75, N2461);
xor XOR2 (N3456, N3452, N1427);
and AND4 (N3457, N3454, N3196, N2571, N2737);
not NOT1 (N3458, N3443);
or OR3 (N3459, N3440, N716, N2532);
or OR2 (N3460, N3449, N2049);
nand NAND3 (N3461, N3431, N2539, N430);
nand NAND3 (N3462, N3455, N1595, N2922);
xor XOR2 (N3463, N3458, N1201);
nor NOR2 (N3464, N3459, N2960);
nand NAND2 (N3465, N3463, N2935);
and AND2 (N3466, N3456, N2177);
nor NOR2 (N3467, N3466, N1361);
or OR3 (N3468, N3460, N667, N1687);
nand NAND2 (N3469, N3464, N3138);
and AND4 (N3470, N3467, N1981, N1180, N555);
and AND4 (N3471, N3453, N719, N3265, N684);
and AND2 (N3472, N3457, N3356);
and AND3 (N3473, N3461, N676, N3217);
buf BUF1 (N3474, N3469);
not NOT1 (N3475, N3465);
buf BUF1 (N3476, N3470);
not NOT1 (N3477, N3473);
buf BUF1 (N3478, N3448);
xor XOR2 (N3479, N3472, N2512);
or OR2 (N3480, N3434, N2688);
not NOT1 (N3481, N3476);
xor XOR2 (N3482, N3462, N1215);
nor NOR4 (N3483, N3471, N894, N2912, N29);
and AND4 (N3484, N3477, N1554, N779, N614);
not NOT1 (N3485, N3480);
or OR2 (N3486, N3481, N567);
buf BUF1 (N3487, N3468);
or OR3 (N3488, N3486, N2228, N2193);
nor NOR3 (N3489, N3474, N992, N403);
buf BUF1 (N3490, N3483);
nand NAND3 (N3491, N3478, N790, N2006);
or OR2 (N3492, N3484, N3249);
not NOT1 (N3493, N3492);
xor XOR2 (N3494, N3490, N2059);
buf BUF1 (N3495, N3494);
nand NAND2 (N3496, N3491, N1896);
buf BUF1 (N3497, N3487);
buf BUF1 (N3498, N3495);
nor NOR2 (N3499, N3488, N1000);
or OR4 (N3500, N3482, N1127, N2073, N616);
buf BUF1 (N3501, N3489);
or OR2 (N3502, N3501, N3138);
and AND4 (N3503, N3493, N1336, N2351, N2274);
xor XOR2 (N3504, N3497, N1205);
buf BUF1 (N3505, N3496);
and AND3 (N3506, N3500, N2882, N207);
and AND3 (N3507, N3505, N1949, N2723);
xor XOR2 (N3508, N3507, N177);
not NOT1 (N3509, N3499);
buf BUF1 (N3510, N3503);
endmodule