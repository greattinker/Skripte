// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;

output N3018,N3023,N3014,N3020,N3009,N3015,N3021,N3019,N3016,N3024;

or OR4 (N25, N7, N12, N5, N22);
xor XOR2 (N26, N17, N20);
and AND3 (N27, N8, N9, N26);
nand NAND2 (N28, N5, N6);
xor XOR2 (N29, N28, N28);
nor NOR4 (N30, N13, N8, N22, N19);
buf BUF1 (N31, N19);
or OR3 (N32, N10, N31, N2);
nor NOR4 (N33, N25, N14, N25, N25);
not NOT1 (N34, N18);
not NOT1 (N35, N20);
or OR4 (N36, N20, N17, N28, N19);
nand NAND3 (N37, N5, N25, N5);
nor NOR3 (N38, N1, N25, N22);
buf BUF1 (N39, N33);
buf BUF1 (N40, N29);
xor XOR2 (N41, N40, N9);
nor NOR2 (N42, N38, N10);
buf BUF1 (N43, N39);
buf BUF1 (N44, N30);
not NOT1 (N45, N36);
not NOT1 (N46, N44);
not NOT1 (N47, N35);
xor XOR2 (N48, N45, N30);
not NOT1 (N49, N46);
not NOT1 (N50, N34);
nor NOR3 (N51, N32, N49, N30);
or OR4 (N52, N17, N50, N16, N20);
and AND2 (N53, N35, N41);
or OR3 (N54, N48, N2, N28);
not NOT1 (N55, N25);
nand NAND2 (N56, N42, N47);
nor NOR3 (N57, N2, N1, N15);
nor NOR2 (N58, N37, N52);
nor NOR4 (N59, N38, N4, N9, N15);
or OR2 (N60, N59, N14);
buf BUF1 (N61, N51);
or OR2 (N62, N60, N48);
xor XOR2 (N63, N58, N53);
xor XOR2 (N64, N17, N36);
or OR2 (N65, N63, N17);
nand NAND2 (N66, N43, N25);
nor NOR3 (N67, N64, N64, N34);
not NOT1 (N68, N66);
or OR3 (N69, N54, N37, N47);
or OR2 (N70, N62, N24);
and AND4 (N71, N55, N34, N7, N12);
nor NOR2 (N72, N57, N9);
and AND4 (N73, N67, N41, N20, N7);
not NOT1 (N74, N68);
or OR3 (N75, N61, N53, N32);
buf BUF1 (N76, N56);
nor NOR3 (N77, N70, N75, N16);
nand NAND3 (N78, N48, N76, N46);
nand NAND3 (N79, N10, N18, N67);
and AND4 (N80, N78, N21, N5, N55);
and AND2 (N81, N65, N52);
buf BUF1 (N82, N74);
xor XOR2 (N83, N77, N23);
not NOT1 (N84, N71);
and AND2 (N85, N82, N7);
xor XOR2 (N86, N79, N37);
xor XOR2 (N87, N81, N61);
xor XOR2 (N88, N87, N13);
nor NOR4 (N89, N88, N18, N22, N47);
xor XOR2 (N90, N69, N70);
not NOT1 (N91, N80);
and AND3 (N92, N91, N44, N35);
not NOT1 (N93, N85);
xor XOR2 (N94, N84, N42);
nand NAND3 (N95, N94, N14, N32);
and AND2 (N96, N73, N70);
or OR3 (N97, N86, N41, N24);
xor XOR2 (N98, N83, N64);
buf BUF1 (N99, N98);
or OR4 (N100, N96, N17, N2, N60);
not NOT1 (N101, N99);
buf BUF1 (N102, N72);
buf BUF1 (N103, N92);
not NOT1 (N104, N90);
nor NOR2 (N105, N104, N25);
nor NOR2 (N106, N100, N59);
not NOT1 (N107, N89);
not NOT1 (N108, N101);
not NOT1 (N109, N106);
nand NAND3 (N110, N105, N82, N77);
xor XOR2 (N111, N103, N52);
buf BUF1 (N112, N97);
nand NAND2 (N113, N110, N10);
not NOT1 (N114, N108);
not NOT1 (N115, N109);
and AND2 (N116, N113, N55);
xor XOR2 (N117, N27, N114);
xor XOR2 (N118, N15, N44);
buf BUF1 (N119, N111);
nand NAND3 (N120, N93, N63, N30);
not NOT1 (N121, N120);
or OR3 (N122, N95, N2, N75);
buf BUF1 (N123, N119);
nor NOR3 (N124, N102, N4, N56);
or OR2 (N125, N122, N56);
buf BUF1 (N126, N117);
or OR2 (N127, N112, N71);
or OR2 (N128, N121, N19);
xor XOR2 (N129, N124, N45);
nand NAND4 (N130, N123, N82, N2, N75);
buf BUF1 (N131, N130);
nand NAND3 (N132, N115, N84, N36);
xor XOR2 (N133, N107, N102);
or OR2 (N134, N118, N87);
not NOT1 (N135, N125);
xor XOR2 (N136, N129, N95);
buf BUF1 (N137, N116);
and AND3 (N138, N131, N21, N8);
or OR3 (N139, N135, N82, N92);
xor XOR2 (N140, N134, N134);
xor XOR2 (N141, N126, N126);
not NOT1 (N142, N128);
xor XOR2 (N143, N142, N108);
and AND2 (N144, N127, N89);
not NOT1 (N145, N143);
or OR3 (N146, N136, N108, N51);
nand NAND4 (N147, N132, N63, N53, N144);
nor NOR2 (N148, N68, N85);
and AND4 (N149, N141, N103, N136, N138);
nor NOR4 (N150, N122, N148, N102, N86);
nor NOR2 (N151, N13, N115);
and AND4 (N152, N151, N68, N70, N15);
buf BUF1 (N153, N137);
xor XOR2 (N154, N145, N133);
and AND4 (N155, N126, N111, N63, N9);
buf BUF1 (N156, N154);
buf BUF1 (N157, N153);
nor NOR3 (N158, N156, N50, N69);
nand NAND4 (N159, N157, N113, N70, N9);
and AND2 (N160, N155, N26);
nand NAND2 (N161, N158, N83);
not NOT1 (N162, N147);
xor XOR2 (N163, N149, N112);
buf BUF1 (N164, N140);
not NOT1 (N165, N163);
not NOT1 (N166, N162);
not NOT1 (N167, N161);
buf BUF1 (N168, N159);
nor NOR3 (N169, N146, N135, N42);
or OR3 (N170, N166, N18, N163);
nand NAND3 (N171, N160, N133, N89);
nor NOR2 (N172, N164, N88);
buf BUF1 (N173, N172);
nor NOR4 (N174, N165, N112, N58, N147);
xor XOR2 (N175, N168, N116);
not NOT1 (N176, N152);
xor XOR2 (N177, N174, N28);
not NOT1 (N178, N169);
buf BUF1 (N179, N170);
nand NAND3 (N180, N167, N22, N140);
nand NAND4 (N181, N139, N102, N114, N171);
or OR2 (N182, N134, N48);
or OR3 (N183, N176, N131, N129);
buf BUF1 (N184, N178);
and AND4 (N185, N182, N96, N9, N175);
nand NAND2 (N186, N134, N8);
nor NOR4 (N187, N177, N95, N52, N185);
not NOT1 (N188, N86);
nand NAND2 (N189, N150, N3);
xor XOR2 (N190, N180, N88);
or OR4 (N191, N179, N171, N14, N180);
nor NOR3 (N192, N173, N167, N151);
nor NOR2 (N193, N187, N84);
nand NAND3 (N194, N189, N91, N110);
not NOT1 (N195, N186);
or OR2 (N196, N184, N49);
not NOT1 (N197, N194);
not NOT1 (N198, N196);
xor XOR2 (N199, N195, N133);
buf BUF1 (N200, N198);
nor NOR2 (N201, N200, N177);
not NOT1 (N202, N197);
and AND3 (N203, N188, N27, N152);
not NOT1 (N204, N202);
not NOT1 (N205, N204);
xor XOR2 (N206, N205, N145);
or OR2 (N207, N190, N14);
xor XOR2 (N208, N207, N41);
nor NOR2 (N209, N206, N115);
buf BUF1 (N210, N203);
nor NOR4 (N211, N193, N177, N167, N142);
nand NAND4 (N212, N208, N47, N42, N141);
and AND4 (N213, N210, N42, N164, N35);
xor XOR2 (N214, N183, N82);
or OR3 (N215, N181, N104, N133);
buf BUF1 (N216, N214);
and AND3 (N217, N213, N180, N130);
and AND3 (N218, N216, N98, N85);
buf BUF1 (N219, N212);
and AND3 (N220, N209, N171, N76);
not NOT1 (N221, N211);
or OR3 (N222, N219, N187, N111);
not NOT1 (N223, N222);
xor XOR2 (N224, N218, N222);
buf BUF1 (N225, N191);
and AND2 (N226, N223, N208);
buf BUF1 (N227, N224);
not NOT1 (N228, N226);
and AND2 (N229, N192, N165);
nor NOR4 (N230, N201, N27, N172, N68);
not NOT1 (N231, N225);
xor XOR2 (N232, N227, N93);
and AND4 (N233, N229, N179, N73, N222);
nor NOR4 (N234, N228, N195, N176, N30);
not NOT1 (N235, N217);
nand NAND4 (N236, N234, N119, N219, N61);
xor XOR2 (N237, N236, N172);
not NOT1 (N238, N221);
not NOT1 (N239, N235);
or OR3 (N240, N220, N230, N101);
buf BUF1 (N241, N61);
buf BUF1 (N242, N239);
nand NAND3 (N243, N240, N74, N169);
and AND2 (N244, N215, N217);
or OR4 (N245, N237, N42, N34, N129);
or OR2 (N246, N238, N193);
buf BUF1 (N247, N233);
nor NOR4 (N248, N232, N220, N12, N42);
buf BUF1 (N249, N243);
not NOT1 (N250, N244);
and AND2 (N251, N249, N10);
nand NAND2 (N252, N250, N117);
not NOT1 (N253, N242);
nand NAND3 (N254, N252, N231, N95);
nor NOR3 (N255, N37, N101, N188);
not NOT1 (N256, N246);
or OR3 (N257, N253, N141, N232);
nand NAND3 (N258, N247, N230, N181);
nand NAND3 (N259, N257, N7, N181);
xor XOR2 (N260, N241, N204);
buf BUF1 (N261, N254);
xor XOR2 (N262, N248, N80);
nand NAND2 (N263, N255, N201);
and AND3 (N264, N199, N11, N223);
not NOT1 (N265, N256);
or OR2 (N266, N245, N177);
buf BUF1 (N267, N266);
and AND4 (N268, N264, N78, N51, N240);
xor XOR2 (N269, N261, N15);
and AND3 (N270, N263, N257, N111);
nand NAND2 (N271, N251, N174);
xor XOR2 (N272, N267, N127);
nor NOR4 (N273, N260, N260, N208, N50);
nand NAND3 (N274, N265, N148, N193);
xor XOR2 (N275, N268, N108);
buf BUF1 (N276, N259);
xor XOR2 (N277, N273, N14);
xor XOR2 (N278, N272, N241);
xor XOR2 (N279, N275, N87);
not NOT1 (N280, N269);
nor NOR4 (N281, N258, N156, N265, N6);
nand NAND3 (N282, N274, N190, N219);
buf BUF1 (N283, N276);
not NOT1 (N284, N282);
xor XOR2 (N285, N271, N226);
nand NAND3 (N286, N278, N85, N250);
nand NAND4 (N287, N277, N175, N222, N191);
xor XOR2 (N288, N280, N256);
or OR4 (N289, N283, N271, N215, N35);
nor NOR3 (N290, N286, N121, N16);
and AND2 (N291, N289, N198);
not NOT1 (N292, N262);
buf BUF1 (N293, N290);
buf BUF1 (N294, N287);
or OR3 (N295, N270, N231, N49);
xor XOR2 (N296, N294, N232);
and AND4 (N297, N293, N91, N138, N71);
xor XOR2 (N298, N281, N295);
buf BUF1 (N299, N111);
buf BUF1 (N300, N297);
or OR3 (N301, N300, N111, N68);
xor XOR2 (N302, N296, N70);
nor NOR2 (N303, N292, N269);
nand NAND2 (N304, N284, N298);
nand NAND3 (N305, N159, N207, N144);
and AND3 (N306, N303, N28, N200);
buf BUF1 (N307, N301);
buf BUF1 (N308, N279);
and AND3 (N309, N305, N139, N305);
xor XOR2 (N310, N309, N18);
xor XOR2 (N311, N306, N82);
nor NOR4 (N312, N304, N50, N23, N237);
xor XOR2 (N313, N308, N303);
or OR4 (N314, N299, N36, N42, N233);
not NOT1 (N315, N291);
nor NOR4 (N316, N313, N23, N283, N200);
nor NOR3 (N317, N315, N230, N84);
nor NOR3 (N318, N316, N226, N93);
xor XOR2 (N319, N318, N48);
nand NAND2 (N320, N317, N109);
nand NAND4 (N321, N285, N319, N166, N193);
or OR2 (N322, N209, N6);
nand NAND2 (N323, N322, N63);
or OR4 (N324, N320, N182, N274, N119);
xor XOR2 (N325, N302, N236);
and AND3 (N326, N321, N279, N166);
and AND2 (N327, N310, N273);
nor NOR2 (N328, N288, N284);
and AND2 (N329, N312, N260);
nand NAND4 (N330, N324, N311, N208, N221);
buf BUF1 (N331, N26);
or OR2 (N332, N323, N238);
nor NOR2 (N333, N328, N2);
nor NOR3 (N334, N325, N155, N106);
nand NAND3 (N335, N327, N206, N96);
buf BUF1 (N336, N335);
nor NOR2 (N337, N336, N198);
and AND3 (N338, N333, N49, N26);
buf BUF1 (N339, N334);
or OR4 (N340, N332, N59, N268, N46);
buf BUF1 (N341, N329);
nand NAND4 (N342, N338, N278, N216, N68);
nand NAND3 (N343, N341, N34, N128);
buf BUF1 (N344, N340);
xor XOR2 (N345, N326, N64);
and AND2 (N346, N344, N147);
nor NOR4 (N347, N330, N198, N327, N215);
and AND3 (N348, N314, N287, N233);
buf BUF1 (N349, N347);
xor XOR2 (N350, N337, N136);
and AND3 (N351, N307, N349, N200);
not NOT1 (N352, N55);
or OR2 (N353, N346, N237);
and AND2 (N354, N351, N123);
nor NOR2 (N355, N343, N26);
buf BUF1 (N356, N342);
xor XOR2 (N357, N339, N304);
not NOT1 (N358, N352);
nand NAND2 (N359, N358, N85);
nand NAND4 (N360, N345, N42, N324, N219);
buf BUF1 (N361, N355);
buf BUF1 (N362, N360);
and AND2 (N363, N353, N340);
and AND3 (N364, N331, N187, N229);
buf BUF1 (N365, N363);
not NOT1 (N366, N365);
buf BUF1 (N367, N359);
and AND4 (N368, N348, N136, N42, N47);
or OR2 (N369, N368, N73);
and AND3 (N370, N362, N259, N86);
nand NAND2 (N371, N354, N220);
or OR4 (N372, N371, N54, N294, N82);
not NOT1 (N373, N366);
or OR2 (N374, N361, N358);
nor NOR2 (N375, N374, N9);
and AND2 (N376, N370, N239);
and AND3 (N377, N369, N164, N238);
nand NAND3 (N378, N373, N2, N38);
xor XOR2 (N379, N356, N134);
not NOT1 (N380, N367);
nand NAND2 (N381, N380, N120);
xor XOR2 (N382, N376, N240);
nand NAND2 (N383, N381, N36);
xor XOR2 (N384, N383, N272);
or OR3 (N385, N382, N155, N362);
not NOT1 (N386, N364);
or OR2 (N387, N375, N36);
buf BUF1 (N388, N377);
nor NOR3 (N389, N387, N378, N284);
not NOT1 (N390, N189);
or OR4 (N391, N385, N117, N118, N165);
xor XOR2 (N392, N386, N105);
nor NOR4 (N393, N388, N110, N76, N348);
xor XOR2 (N394, N389, N63);
nand NAND3 (N395, N391, N218, N197);
and AND2 (N396, N357, N187);
nor NOR2 (N397, N379, N195);
not NOT1 (N398, N390);
and AND2 (N399, N372, N341);
and AND2 (N400, N396, N115);
or OR4 (N401, N350, N168, N115, N217);
buf BUF1 (N402, N394);
nand NAND2 (N403, N400, N161);
not NOT1 (N404, N401);
buf BUF1 (N405, N397);
nor NOR2 (N406, N398, N157);
or OR4 (N407, N395, N5, N214, N181);
or OR3 (N408, N384, N117, N225);
or OR4 (N409, N393, N103, N259, N162);
and AND3 (N410, N399, N287, N85);
xor XOR2 (N411, N408, N358);
xor XOR2 (N412, N407, N325);
nand NAND2 (N413, N404, N170);
buf BUF1 (N414, N413);
nand NAND4 (N415, N409, N407, N308, N362);
buf BUF1 (N416, N411);
nor NOR3 (N417, N412, N356, N205);
xor XOR2 (N418, N416, N189);
buf BUF1 (N419, N392);
xor XOR2 (N420, N419, N377);
buf BUF1 (N421, N415);
xor XOR2 (N422, N410, N415);
xor XOR2 (N423, N414, N20);
and AND2 (N424, N420, N366);
nand NAND4 (N425, N402, N101, N197, N77);
and AND2 (N426, N403, N321);
nor NOR4 (N427, N426, N190, N278, N20);
xor XOR2 (N428, N417, N232);
nand NAND4 (N429, N418, N252, N227, N7);
nand NAND3 (N430, N427, N375, N237);
buf BUF1 (N431, N428);
or OR4 (N432, N430, N75, N19, N126);
or OR4 (N433, N432, N319, N133, N24);
buf BUF1 (N434, N425);
or OR2 (N435, N423, N344);
buf BUF1 (N436, N434);
xor XOR2 (N437, N405, N80);
nor NOR2 (N438, N422, N2);
and AND4 (N439, N421, N12, N133, N148);
or OR2 (N440, N436, N152);
buf BUF1 (N441, N439);
nor NOR3 (N442, N435, N129, N313);
buf BUF1 (N443, N429);
buf BUF1 (N444, N424);
or OR4 (N445, N442, N308, N24, N440);
and AND3 (N446, N115, N39, N388);
xor XOR2 (N447, N437, N309);
or OR2 (N448, N447, N394);
and AND4 (N449, N406, N343, N215, N86);
or OR4 (N450, N444, N348, N333, N420);
xor XOR2 (N451, N450, N61);
and AND4 (N452, N448, N16, N84, N39);
and AND3 (N453, N438, N219, N407);
and AND3 (N454, N445, N405, N161);
xor XOR2 (N455, N433, N236);
nor NOR4 (N456, N452, N351, N130, N83);
nor NOR2 (N457, N454, N334);
or OR4 (N458, N431, N206, N162, N435);
or OR3 (N459, N455, N456, N228);
not NOT1 (N460, N430);
nand NAND3 (N461, N441, N293, N111);
nor NOR3 (N462, N446, N310, N157);
not NOT1 (N463, N451);
buf BUF1 (N464, N461);
or OR4 (N465, N459, N417, N13, N448);
buf BUF1 (N466, N460);
nand NAND3 (N467, N443, N308, N232);
xor XOR2 (N468, N463, N226);
not NOT1 (N469, N466);
buf BUF1 (N470, N464);
xor XOR2 (N471, N470, N22);
nor NOR4 (N472, N457, N360, N242, N25);
and AND3 (N473, N467, N38, N293);
nand NAND4 (N474, N449, N84, N175, N71);
nor NOR3 (N475, N471, N159, N372);
buf BUF1 (N476, N458);
and AND4 (N477, N475, N472, N175, N153);
not NOT1 (N478, N334);
and AND4 (N479, N453, N101, N89, N406);
and AND4 (N480, N468, N268, N100, N467);
nand NAND2 (N481, N479, N312);
and AND2 (N482, N465, N278);
buf BUF1 (N483, N469);
nand NAND3 (N484, N477, N348, N89);
nand NAND3 (N485, N478, N422, N88);
nor NOR4 (N486, N483, N188, N233, N453);
xor XOR2 (N487, N481, N289);
not NOT1 (N488, N487);
not NOT1 (N489, N484);
buf BUF1 (N490, N473);
nor NOR3 (N491, N482, N392, N158);
and AND4 (N492, N485, N201, N181, N461);
not NOT1 (N493, N476);
xor XOR2 (N494, N493, N458);
nor NOR3 (N495, N494, N438, N462);
nand NAND2 (N496, N156, N154);
xor XOR2 (N497, N495, N116);
buf BUF1 (N498, N491);
xor XOR2 (N499, N496, N392);
and AND2 (N500, N499, N6);
nand NAND3 (N501, N474, N137, N2);
buf BUF1 (N502, N492);
nor NOR2 (N503, N502, N269);
xor XOR2 (N504, N497, N373);
xor XOR2 (N505, N490, N397);
xor XOR2 (N506, N480, N66);
not NOT1 (N507, N488);
and AND4 (N508, N503, N162, N113, N43);
or OR4 (N509, N506, N140, N28, N72);
and AND3 (N510, N500, N312, N346);
not NOT1 (N511, N489);
nand NAND2 (N512, N486, N159);
nand NAND2 (N513, N511, N14);
buf BUF1 (N514, N501);
or OR3 (N515, N509, N165, N179);
and AND2 (N516, N510, N491);
not NOT1 (N517, N515);
not NOT1 (N518, N512);
not NOT1 (N519, N507);
xor XOR2 (N520, N508, N193);
or OR3 (N521, N498, N394, N194);
not NOT1 (N522, N516);
nor NOR3 (N523, N518, N430, N290);
xor XOR2 (N524, N522, N205);
or OR2 (N525, N513, N46);
or OR3 (N526, N523, N289, N468);
buf BUF1 (N527, N524);
nor NOR4 (N528, N519, N21, N344, N461);
not NOT1 (N529, N517);
not NOT1 (N530, N514);
nor NOR2 (N531, N527, N239);
and AND2 (N532, N529, N518);
nand NAND2 (N533, N530, N104);
nor NOR3 (N534, N525, N52, N443);
buf BUF1 (N535, N531);
xor XOR2 (N536, N532, N153);
and AND2 (N537, N526, N453);
nand NAND3 (N538, N505, N149, N301);
or OR2 (N539, N528, N13);
nor NOR2 (N540, N521, N88);
not NOT1 (N541, N534);
or OR2 (N542, N535, N236);
buf BUF1 (N543, N520);
or OR2 (N544, N541, N134);
nor NOR3 (N545, N539, N418, N97);
nand NAND3 (N546, N536, N447, N79);
nor NOR2 (N547, N504, N341);
nor NOR4 (N548, N547, N457, N30, N248);
nor NOR2 (N549, N538, N57);
nor NOR3 (N550, N548, N333, N247);
or OR2 (N551, N545, N402);
and AND3 (N552, N542, N246, N222);
nand NAND3 (N553, N537, N549, N99);
nor NOR3 (N554, N151, N522, N382);
buf BUF1 (N555, N533);
buf BUF1 (N556, N543);
and AND4 (N557, N550, N349, N131, N279);
nand NAND4 (N558, N544, N187, N142, N2);
buf BUF1 (N559, N558);
buf BUF1 (N560, N557);
buf BUF1 (N561, N553);
nor NOR4 (N562, N559, N530, N495, N212);
and AND4 (N563, N561, N89, N238, N447);
and AND3 (N564, N556, N271, N289);
or OR3 (N565, N546, N165, N402);
not NOT1 (N566, N554);
or OR2 (N567, N565, N433);
xor XOR2 (N568, N563, N13);
buf BUF1 (N569, N555);
nand NAND2 (N570, N540, N369);
xor XOR2 (N571, N569, N163);
or OR3 (N572, N570, N142, N314);
not NOT1 (N573, N552);
not NOT1 (N574, N572);
buf BUF1 (N575, N566);
nand NAND3 (N576, N562, N149, N39);
nand NAND3 (N577, N571, N203, N552);
xor XOR2 (N578, N575, N14);
nand NAND4 (N579, N578, N267, N141, N29);
and AND3 (N580, N577, N424, N404);
not NOT1 (N581, N564);
xor XOR2 (N582, N567, N26);
nor NOR4 (N583, N581, N166, N229, N497);
or OR4 (N584, N573, N100, N473, N171);
nor NOR2 (N585, N576, N316);
or OR3 (N586, N568, N517, N565);
nand NAND3 (N587, N586, N359, N543);
buf BUF1 (N588, N587);
buf BUF1 (N589, N583);
nand NAND2 (N590, N560, N397);
not NOT1 (N591, N590);
or OR3 (N592, N591, N463, N418);
buf BUF1 (N593, N580);
xor XOR2 (N594, N574, N470);
and AND2 (N595, N582, N582);
xor XOR2 (N596, N589, N138);
nor NOR4 (N597, N595, N349, N391, N146);
not NOT1 (N598, N594);
nor NOR2 (N599, N588, N392);
nor NOR3 (N600, N585, N431, N387);
and AND4 (N601, N584, N133, N578, N428);
buf BUF1 (N602, N598);
nor NOR4 (N603, N601, N106, N478, N337);
nand NAND3 (N604, N551, N444, N29);
not NOT1 (N605, N604);
and AND4 (N606, N593, N434, N569, N604);
not NOT1 (N607, N596);
nor NOR3 (N608, N597, N243, N309);
not NOT1 (N609, N603);
nand NAND4 (N610, N599, N299, N120, N229);
nand NAND2 (N611, N608, N110);
buf BUF1 (N612, N600);
nand NAND3 (N613, N607, N248, N119);
buf BUF1 (N614, N579);
xor XOR2 (N615, N611, N570);
or OR4 (N616, N610, N447, N580, N592);
and AND3 (N617, N205, N88, N614);
xor XOR2 (N618, N259, N32);
and AND3 (N619, N612, N153, N515);
nand NAND2 (N620, N615, N118);
and AND2 (N621, N602, N41);
or OR4 (N622, N621, N189, N472, N435);
nor NOR4 (N623, N617, N3, N583, N279);
nor NOR4 (N624, N618, N350, N281, N16);
buf BUF1 (N625, N605);
not NOT1 (N626, N609);
buf BUF1 (N627, N619);
buf BUF1 (N628, N625);
nor NOR2 (N629, N616, N93);
buf BUF1 (N630, N626);
nor NOR4 (N631, N629, N561, N123, N8);
nor NOR4 (N632, N613, N160, N2, N388);
xor XOR2 (N633, N630, N609);
xor XOR2 (N634, N622, N211);
nor NOR4 (N635, N606, N558, N217, N595);
nand NAND4 (N636, N633, N364, N509, N526);
xor XOR2 (N637, N627, N464);
and AND2 (N638, N620, N526);
nand NAND2 (N639, N628, N83);
nand NAND4 (N640, N638, N401, N494, N182);
not NOT1 (N641, N637);
xor XOR2 (N642, N632, N293);
and AND3 (N643, N634, N224, N265);
or OR4 (N644, N624, N122, N504, N241);
buf BUF1 (N645, N641);
or OR3 (N646, N636, N435, N577);
xor XOR2 (N647, N642, N49);
nand NAND4 (N648, N646, N294, N346, N511);
buf BUF1 (N649, N644);
and AND2 (N650, N623, N425);
xor XOR2 (N651, N647, N466);
and AND2 (N652, N648, N562);
buf BUF1 (N653, N650);
xor XOR2 (N654, N631, N12);
nand NAND4 (N655, N643, N394, N580, N313);
buf BUF1 (N656, N654);
and AND4 (N657, N639, N335, N92, N568);
and AND3 (N658, N640, N524, N154);
buf BUF1 (N659, N655);
and AND3 (N660, N653, N646, N158);
nor NOR3 (N661, N652, N61, N621);
xor XOR2 (N662, N660, N70);
and AND4 (N663, N658, N552, N385, N478);
nor NOR2 (N664, N645, N156);
xor XOR2 (N665, N651, N558);
xor XOR2 (N666, N661, N228);
nor NOR2 (N667, N666, N603);
xor XOR2 (N668, N663, N577);
not NOT1 (N669, N635);
nand NAND4 (N670, N668, N465, N207, N205);
xor XOR2 (N671, N665, N62);
buf BUF1 (N672, N649);
and AND2 (N673, N672, N485);
nand NAND3 (N674, N670, N314, N333);
buf BUF1 (N675, N657);
nand NAND2 (N676, N659, N216);
nand NAND2 (N677, N669, N188);
buf BUF1 (N678, N673);
nor NOR3 (N679, N656, N252, N311);
xor XOR2 (N680, N675, N379);
nand NAND4 (N681, N676, N152, N620, N551);
nand NAND3 (N682, N681, N149, N577);
or OR2 (N683, N667, N419);
nand NAND3 (N684, N664, N441, N5);
nor NOR3 (N685, N682, N385, N656);
or OR4 (N686, N678, N252, N636, N25);
buf BUF1 (N687, N677);
or OR2 (N688, N674, N645);
buf BUF1 (N689, N687);
xor XOR2 (N690, N686, N136);
nand NAND4 (N691, N662, N673, N494, N640);
xor XOR2 (N692, N688, N74);
buf BUF1 (N693, N690);
xor XOR2 (N694, N679, N232);
nand NAND4 (N695, N692, N36, N402, N36);
nand NAND2 (N696, N684, N82);
nand NAND3 (N697, N696, N299, N450);
nor NOR2 (N698, N671, N396);
or OR3 (N699, N698, N638, N386);
buf BUF1 (N700, N699);
xor XOR2 (N701, N693, N79);
nand NAND3 (N702, N694, N526, N311);
or OR3 (N703, N691, N144, N459);
not NOT1 (N704, N697);
nand NAND4 (N705, N701, N265, N489, N505);
nor NOR3 (N706, N683, N509, N231);
nor NOR4 (N707, N706, N550, N547, N306);
and AND3 (N708, N703, N58, N674);
not NOT1 (N709, N705);
nor NOR3 (N710, N708, N204, N522);
nand NAND4 (N711, N707, N631, N553, N89);
nand NAND2 (N712, N685, N323);
nor NOR2 (N713, N711, N340);
nor NOR2 (N714, N710, N579);
xor XOR2 (N715, N702, N121);
nand NAND3 (N716, N700, N507, N534);
nand NAND2 (N717, N689, N446);
xor XOR2 (N718, N695, N186);
and AND3 (N719, N715, N703, N236);
xor XOR2 (N720, N714, N559);
not NOT1 (N721, N680);
or OR4 (N722, N717, N22, N498, N504);
nor NOR4 (N723, N713, N294, N377, N704);
or OR2 (N724, N517, N683);
or OR2 (N725, N721, N334);
xor XOR2 (N726, N722, N354);
or OR4 (N727, N726, N350, N317, N419);
and AND3 (N728, N718, N253, N723);
or OR4 (N729, N512, N477, N181, N123);
or OR3 (N730, N720, N654, N599);
and AND2 (N731, N730, N526);
xor XOR2 (N732, N719, N510);
and AND4 (N733, N725, N596, N289, N145);
and AND3 (N734, N712, N279, N328);
buf BUF1 (N735, N727);
buf BUF1 (N736, N728);
not NOT1 (N737, N736);
or OR3 (N738, N716, N730, N89);
nand NAND2 (N739, N737, N28);
xor XOR2 (N740, N724, N22);
nor NOR4 (N741, N729, N256, N18, N344);
and AND4 (N742, N733, N406, N23, N11);
buf BUF1 (N743, N734);
nor NOR2 (N744, N735, N616);
xor XOR2 (N745, N740, N604);
and AND3 (N746, N745, N635, N127);
nor NOR4 (N747, N739, N319, N640, N206);
xor XOR2 (N748, N738, N95);
buf BUF1 (N749, N746);
nand NAND4 (N750, N748, N700, N45, N710);
or OR4 (N751, N731, N447, N687, N360);
or OR2 (N752, N742, N333);
xor XOR2 (N753, N732, N520);
xor XOR2 (N754, N744, N245);
or OR4 (N755, N751, N313, N714, N419);
nor NOR4 (N756, N752, N568, N473, N529);
or OR2 (N757, N747, N308);
and AND3 (N758, N749, N305, N214);
xor XOR2 (N759, N741, N526);
buf BUF1 (N760, N754);
xor XOR2 (N761, N755, N39);
nor NOR4 (N762, N753, N156, N422, N66);
and AND4 (N763, N759, N650, N475, N738);
nand NAND2 (N764, N758, N320);
or OR4 (N765, N763, N462, N175, N394);
not NOT1 (N766, N764);
nand NAND4 (N767, N756, N300, N604, N687);
not NOT1 (N768, N765);
buf BUF1 (N769, N750);
xor XOR2 (N770, N767, N115);
nand NAND2 (N771, N757, N74);
buf BUF1 (N772, N770);
nand NAND2 (N773, N771, N708);
or OR2 (N774, N768, N510);
not NOT1 (N775, N774);
or OR2 (N776, N775, N241);
or OR4 (N777, N776, N133, N600, N478);
or OR2 (N778, N709, N682);
or OR3 (N779, N778, N453, N279);
or OR2 (N780, N760, N214);
buf BUF1 (N781, N772);
and AND3 (N782, N780, N738, N179);
nand NAND4 (N783, N761, N84, N410, N537);
nand NAND4 (N784, N773, N34, N391, N248);
or OR4 (N785, N762, N734, N411, N585);
and AND4 (N786, N779, N479, N513, N326);
and AND2 (N787, N782, N265);
or OR3 (N788, N783, N442, N736);
xor XOR2 (N789, N787, N497);
xor XOR2 (N790, N788, N538);
and AND4 (N791, N789, N494, N459, N196);
xor XOR2 (N792, N785, N410);
and AND3 (N793, N791, N367, N743);
nand NAND3 (N794, N692, N530, N392);
not NOT1 (N795, N766);
and AND3 (N796, N781, N393, N441);
xor XOR2 (N797, N796, N207);
buf BUF1 (N798, N786);
buf BUF1 (N799, N794);
and AND4 (N800, N798, N584, N145, N165);
and AND4 (N801, N795, N796, N603, N105);
nor NOR2 (N802, N801, N155);
not NOT1 (N803, N784);
xor XOR2 (N804, N792, N549);
and AND4 (N805, N803, N14, N244, N790);
not NOT1 (N806, N297);
buf BUF1 (N807, N806);
xor XOR2 (N808, N769, N543);
nor NOR3 (N809, N802, N691, N210);
not NOT1 (N810, N809);
nor NOR2 (N811, N797, N385);
not NOT1 (N812, N799);
and AND3 (N813, N807, N620, N682);
and AND3 (N814, N811, N665, N522);
nand NAND2 (N815, N808, N257);
not NOT1 (N816, N813);
and AND4 (N817, N816, N782, N727, N345);
nand NAND3 (N818, N817, N118, N212);
xor XOR2 (N819, N777, N725);
buf BUF1 (N820, N814);
xor XOR2 (N821, N815, N468);
buf BUF1 (N822, N804);
nor NOR2 (N823, N810, N711);
nand NAND4 (N824, N819, N680, N819, N167);
not NOT1 (N825, N805);
xor XOR2 (N826, N818, N744);
nor NOR2 (N827, N826, N798);
xor XOR2 (N828, N820, N460);
xor XOR2 (N829, N825, N653);
xor XOR2 (N830, N793, N755);
or OR4 (N831, N828, N376, N796, N665);
or OR3 (N832, N812, N711, N729);
buf BUF1 (N833, N823);
nand NAND2 (N834, N821, N119);
nor NOR4 (N835, N829, N614, N665, N253);
or OR2 (N836, N832, N164);
buf BUF1 (N837, N831);
nor NOR4 (N838, N836, N360, N814, N449);
xor XOR2 (N839, N824, N443);
and AND2 (N840, N830, N287);
not NOT1 (N841, N827);
not NOT1 (N842, N840);
and AND3 (N843, N839, N310, N104);
and AND2 (N844, N835, N402);
and AND2 (N845, N841, N800);
not NOT1 (N846, N366);
buf BUF1 (N847, N833);
or OR4 (N848, N838, N803, N460, N417);
not NOT1 (N849, N848);
buf BUF1 (N850, N842);
nor NOR2 (N851, N822, N814);
and AND4 (N852, N850, N501, N237, N836);
and AND4 (N853, N852, N409, N744, N668);
xor XOR2 (N854, N847, N484);
xor XOR2 (N855, N849, N777);
buf BUF1 (N856, N844);
nand NAND4 (N857, N845, N400, N830, N154);
xor XOR2 (N858, N843, N627);
not NOT1 (N859, N837);
nor NOR3 (N860, N856, N242, N846);
nor NOR2 (N861, N17, N661);
xor XOR2 (N862, N858, N371);
xor XOR2 (N863, N857, N243);
and AND2 (N864, N851, N133);
nand NAND3 (N865, N834, N855, N368);
xor XOR2 (N866, N842, N467);
not NOT1 (N867, N863);
not NOT1 (N868, N867);
nor NOR2 (N869, N866, N850);
nor NOR2 (N870, N869, N684);
nor NOR3 (N871, N868, N298, N521);
and AND4 (N872, N859, N240, N33, N785);
nand NAND3 (N873, N860, N707, N107);
not NOT1 (N874, N853);
nand NAND3 (N875, N874, N824, N862);
nor NOR3 (N876, N321, N162, N794);
nand NAND2 (N877, N875, N768);
buf BUF1 (N878, N854);
nand NAND3 (N879, N878, N508, N108);
nor NOR2 (N880, N861, N223);
nor NOR3 (N881, N877, N283, N730);
buf BUF1 (N882, N873);
xor XOR2 (N883, N880, N37);
buf BUF1 (N884, N864);
xor XOR2 (N885, N883, N611);
not NOT1 (N886, N870);
xor XOR2 (N887, N876, N456);
xor XOR2 (N888, N886, N136);
nand NAND3 (N889, N872, N38, N365);
and AND4 (N890, N882, N387, N174, N860);
buf BUF1 (N891, N889);
not NOT1 (N892, N885);
and AND4 (N893, N881, N625, N553, N278);
nand NAND3 (N894, N879, N696, N170);
not NOT1 (N895, N891);
not NOT1 (N896, N884);
nand NAND3 (N897, N895, N678, N327);
or OR3 (N898, N897, N172, N504);
nand NAND3 (N899, N871, N660, N388);
or OR3 (N900, N894, N846, N787);
and AND2 (N901, N888, N336);
nor NOR3 (N902, N899, N339, N683);
nor NOR3 (N903, N890, N253, N851);
buf BUF1 (N904, N903);
nor NOR3 (N905, N900, N70, N542);
buf BUF1 (N906, N887);
not NOT1 (N907, N898);
and AND3 (N908, N865, N311, N797);
and AND4 (N909, N902, N308, N570, N669);
nand NAND2 (N910, N901, N480);
nor NOR2 (N911, N908, N357);
and AND2 (N912, N896, N350);
and AND3 (N913, N906, N716, N510);
not NOT1 (N914, N911);
nor NOR4 (N915, N904, N371, N261, N526);
buf BUF1 (N916, N914);
nand NAND3 (N917, N893, N555, N161);
nor NOR2 (N918, N915, N284);
or OR4 (N919, N910, N602, N603, N653);
and AND3 (N920, N918, N604, N149);
or OR4 (N921, N916, N500, N555, N236);
or OR3 (N922, N913, N653, N658);
nand NAND3 (N923, N905, N449, N922);
nor NOR2 (N924, N644, N16);
not NOT1 (N925, N920);
xor XOR2 (N926, N923, N153);
buf BUF1 (N927, N917);
nor NOR3 (N928, N924, N722, N663);
not NOT1 (N929, N928);
or OR4 (N930, N929, N882, N910, N724);
or OR4 (N931, N927, N705, N316, N79);
buf BUF1 (N932, N925);
and AND4 (N933, N921, N552, N45, N462);
and AND4 (N934, N931, N70, N550, N320);
buf BUF1 (N935, N919);
xor XOR2 (N936, N926, N144);
buf BUF1 (N937, N934);
nand NAND2 (N938, N892, N788);
or OR3 (N939, N937, N89, N365);
nand NAND3 (N940, N935, N798, N790);
nand NAND4 (N941, N933, N90, N758, N244);
or OR3 (N942, N941, N81, N703);
buf BUF1 (N943, N942);
nand NAND3 (N944, N930, N254, N474);
not NOT1 (N945, N936);
buf BUF1 (N946, N932);
nor NOR4 (N947, N909, N916, N49, N388);
not NOT1 (N948, N907);
nor NOR2 (N949, N939, N108);
not NOT1 (N950, N945);
not NOT1 (N951, N949);
buf BUF1 (N952, N940);
not NOT1 (N953, N938);
nor NOR3 (N954, N947, N857, N337);
buf BUF1 (N955, N951);
or OR3 (N956, N946, N773, N327);
nor NOR3 (N957, N953, N75, N193);
nor NOR3 (N958, N912, N802, N283);
nand NAND3 (N959, N944, N611, N609);
nand NAND3 (N960, N958, N625, N81);
xor XOR2 (N961, N952, N721);
nand NAND2 (N962, N956, N571);
nor NOR3 (N963, N960, N708, N318);
nor NOR4 (N964, N955, N925, N511, N254);
buf BUF1 (N965, N963);
xor XOR2 (N966, N961, N108);
nor NOR2 (N967, N959, N774);
nand NAND4 (N968, N943, N133, N421, N927);
buf BUF1 (N969, N950);
not NOT1 (N970, N969);
and AND2 (N971, N962, N8);
buf BUF1 (N972, N957);
nand NAND2 (N973, N970, N664);
not NOT1 (N974, N948);
nand NAND2 (N975, N972, N279);
not NOT1 (N976, N964);
and AND2 (N977, N976, N582);
buf BUF1 (N978, N971);
not NOT1 (N979, N967);
nand NAND2 (N980, N965, N774);
nand NAND4 (N981, N977, N548, N484, N498);
and AND2 (N982, N979, N940);
xor XOR2 (N983, N980, N617);
and AND2 (N984, N973, N687);
and AND4 (N985, N981, N758, N159, N562);
buf BUF1 (N986, N985);
nor NOR3 (N987, N982, N683, N591);
nand NAND4 (N988, N974, N60, N203, N908);
buf BUF1 (N989, N987);
not NOT1 (N990, N989);
nand NAND3 (N991, N984, N323, N823);
and AND3 (N992, N968, N445, N205);
nor NOR3 (N993, N966, N276, N467);
xor XOR2 (N994, N986, N838);
buf BUF1 (N995, N978);
nor NOR2 (N996, N988, N169);
buf BUF1 (N997, N975);
buf BUF1 (N998, N997);
and AND3 (N999, N992, N469, N392);
xor XOR2 (N1000, N954, N769);
nor NOR4 (N1001, N991, N322, N282, N189);
xor XOR2 (N1002, N994, N848);
buf BUF1 (N1003, N998);
buf BUF1 (N1004, N1000);
nor NOR3 (N1005, N999, N823, N729);
and AND3 (N1006, N1004, N681, N209);
xor XOR2 (N1007, N990, N921);
nand NAND2 (N1008, N1005, N679);
nor NOR3 (N1009, N993, N595, N159);
buf BUF1 (N1010, N1003);
and AND3 (N1011, N1010, N627, N513);
or OR2 (N1012, N983, N582);
or OR2 (N1013, N1007, N564);
or OR4 (N1014, N1011, N395, N672, N569);
nand NAND4 (N1015, N1009, N173, N548, N707);
not NOT1 (N1016, N1013);
xor XOR2 (N1017, N1014, N934);
buf BUF1 (N1018, N995);
not NOT1 (N1019, N1012);
xor XOR2 (N1020, N1016, N967);
buf BUF1 (N1021, N1002);
and AND3 (N1022, N1019, N710, N1000);
nand NAND3 (N1023, N1008, N715, N1008);
buf BUF1 (N1024, N1020);
and AND2 (N1025, N1023, N146);
not NOT1 (N1026, N1017);
nor NOR3 (N1027, N996, N847, N464);
not NOT1 (N1028, N1022);
or OR2 (N1029, N1021, N506);
and AND4 (N1030, N1015, N729, N903, N276);
nand NAND2 (N1031, N1001, N317);
and AND2 (N1032, N1025, N986);
buf BUF1 (N1033, N1006);
not NOT1 (N1034, N1030);
nand NAND2 (N1035, N1031, N962);
nor NOR2 (N1036, N1018, N214);
and AND2 (N1037, N1034, N620);
or OR3 (N1038, N1029, N843, N1031);
nor NOR3 (N1039, N1033, N611, N759);
or OR2 (N1040, N1026, N351);
not NOT1 (N1041, N1040);
and AND3 (N1042, N1037, N77, N625);
nand NAND4 (N1043, N1024, N55, N631, N465);
xor XOR2 (N1044, N1027, N584);
nand NAND4 (N1045, N1044, N210, N289, N37);
or OR4 (N1046, N1036, N284, N635, N407);
buf BUF1 (N1047, N1046);
xor XOR2 (N1048, N1045, N260);
nor NOR2 (N1049, N1042, N880);
buf BUF1 (N1050, N1039);
nand NAND2 (N1051, N1028, N216);
or OR4 (N1052, N1038, N73, N836, N483);
or OR2 (N1053, N1041, N341);
or OR2 (N1054, N1051, N618);
and AND4 (N1055, N1054, N442, N564, N847);
nand NAND2 (N1056, N1032, N1032);
not NOT1 (N1057, N1049);
xor XOR2 (N1058, N1055, N185);
not NOT1 (N1059, N1057);
nor NOR3 (N1060, N1052, N336, N802);
or OR4 (N1061, N1056, N630, N365, N143);
xor XOR2 (N1062, N1060, N333);
and AND2 (N1063, N1059, N341);
nand NAND2 (N1064, N1035, N597);
not NOT1 (N1065, N1063);
buf BUF1 (N1066, N1062);
nor NOR2 (N1067, N1064, N426);
and AND2 (N1068, N1048, N47);
nor NOR3 (N1069, N1066, N261, N255);
nand NAND3 (N1070, N1043, N249, N832);
xor XOR2 (N1071, N1058, N661);
not NOT1 (N1072, N1070);
not NOT1 (N1073, N1053);
not NOT1 (N1074, N1068);
nand NAND3 (N1075, N1074, N853, N445);
not NOT1 (N1076, N1069);
buf BUF1 (N1077, N1065);
xor XOR2 (N1078, N1061, N803);
or OR3 (N1079, N1078, N510, N1058);
buf BUF1 (N1080, N1075);
buf BUF1 (N1081, N1073);
nand NAND4 (N1082, N1072, N150, N397, N60);
nand NAND3 (N1083, N1067, N833, N50);
xor XOR2 (N1084, N1077, N36);
and AND3 (N1085, N1081, N778, N576);
nor NOR4 (N1086, N1084, N492, N763, N830);
nor NOR3 (N1087, N1083, N1073, N84);
not NOT1 (N1088, N1080);
or OR4 (N1089, N1079, N289, N130, N258);
nand NAND2 (N1090, N1071, N133);
not NOT1 (N1091, N1082);
buf BUF1 (N1092, N1088);
not NOT1 (N1093, N1047);
nor NOR3 (N1094, N1089, N420, N956);
nor NOR2 (N1095, N1091, N990);
xor XOR2 (N1096, N1092, N150);
xor XOR2 (N1097, N1094, N803);
and AND2 (N1098, N1097, N784);
or OR2 (N1099, N1086, N1002);
or OR4 (N1100, N1098, N313, N1071, N382);
or OR3 (N1101, N1087, N175, N423);
not NOT1 (N1102, N1085);
nor NOR2 (N1103, N1102, N461);
not NOT1 (N1104, N1099);
not NOT1 (N1105, N1093);
and AND4 (N1106, N1095, N484, N261, N896);
xor XOR2 (N1107, N1106, N417);
or OR4 (N1108, N1096, N254, N713, N1050);
buf BUF1 (N1109, N701);
or OR3 (N1110, N1103, N556, N142);
not NOT1 (N1111, N1108);
nor NOR2 (N1112, N1100, N288);
not NOT1 (N1113, N1112);
not NOT1 (N1114, N1110);
nand NAND3 (N1115, N1090, N520, N405);
nor NOR3 (N1116, N1113, N66, N958);
and AND4 (N1117, N1109, N618, N897, N692);
and AND4 (N1118, N1116, N665, N187, N356);
and AND4 (N1119, N1101, N926, N693, N752);
buf BUF1 (N1120, N1107);
buf BUF1 (N1121, N1119);
not NOT1 (N1122, N1120);
or OR4 (N1123, N1105, N837, N8, N838);
nand NAND4 (N1124, N1076, N942, N259, N750);
nor NOR3 (N1125, N1121, N802, N436);
and AND3 (N1126, N1115, N342, N1076);
buf BUF1 (N1127, N1118);
nor NOR3 (N1128, N1125, N660, N41);
nand NAND2 (N1129, N1124, N831);
buf BUF1 (N1130, N1128);
and AND3 (N1131, N1130, N229, N451);
xor XOR2 (N1132, N1123, N300);
or OR3 (N1133, N1127, N759, N637);
nor NOR3 (N1134, N1133, N286, N810);
and AND3 (N1135, N1104, N254, N319);
or OR4 (N1136, N1117, N935, N643, N733);
buf BUF1 (N1137, N1136);
not NOT1 (N1138, N1129);
and AND3 (N1139, N1134, N537, N424);
not NOT1 (N1140, N1137);
or OR3 (N1141, N1126, N1136, N870);
not NOT1 (N1142, N1122);
or OR3 (N1143, N1142, N1061, N474);
nor NOR4 (N1144, N1143, N49, N239, N404);
not NOT1 (N1145, N1135);
not NOT1 (N1146, N1139);
nor NOR3 (N1147, N1132, N1060, N374);
xor XOR2 (N1148, N1146, N1116);
xor XOR2 (N1149, N1141, N519);
xor XOR2 (N1150, N1140, N207);
nand NAND4 (N1151, N1149, N635, N1119, N45);
xor XOR2 (N1152, N1145, N99);
xor XOR2 (N1153, N1138, N97);
and AND3 (N1154, N1131, N1015, N585);
nor NOR3 (N1155, N1154, N711, N1125);
or OR4 (N1156, N1150, N261, N900, N966);
or OR4 (N1157, N1151, N905, N478, N166);
buf BUF1 (N1158, N1144);
nor NOR2 (N1159, N1152, N488);
or OR2 (N1160, N1148, N803);
nor NOR4 (N1161, N1114, N1006, N174, N938);
xor XOR2 (N1162, N1161, N580);
and AND4 (N1163, N1153, N1057, N720, N426);
not NOT1 (N1164, N1162);
nor NOR2 (N1165, N1155, N1078);
and AND2 (N1166, N1156, N239);
not NOT1 (N1167, N1159);
or OR2 (N1168, N1164, N383);
and AND3 (N1169, N1168, N646, N23);
or OR3 (N1170, N1111, N1144, N1045);
buf BUF1 (N1171, N1147);
nand NAND4 (N1172, N1167, N1103, N640, N953);
or OR4 (N1173, N1171, N1020, N559, N533);
nor NOR3 (N1174, N1163, N410, N55);
nand NAND4 (N1175, N1166, N922, N528, N596);
buf BUF1 (N1176, N1160);
buf BUF1 (N1177, N1172);
xor XOR2 (N1178, N1170, N489);
nand NAND3 (N1179, N1169, N264, N923);
or OR4 (N1180, N1176, N375, N16, N996);
xor XOR2 (N1181, N1177, N397);
nor NOR4 (N1182, N1173, N114, N1072, N822);
not NOT1 (N1183, N1158);
and AND2 (N1184, N1181, N792);
and AND3 (N1185, N1184, N79, N674);
or OR3 (N1186, N1179, N189, N90);
nor NOR2 (N1187, N1183, N503);
xor XOR2 (N1188, N1186, N619);
or OR4 (N1189, N1178, N538, N440, N800);
buf BUF1 (N1190, N1188);
nand NAND4 (N1191, N1175, N63, N91, N1016);
or OR2 (N1192, N1190, N404);
xor XOR2 (N1193, N1180, N906);
nand NAND2 (N1194, N1174, N154);
buf BUF1 (N1195, N1187);
nor NOR2 (N1196, N1185, N444);
buf BUF1 (N1197, N1157);
buf BUF1 (N1198, N1195);
and AND3 (N1199, N1193, N205, N219);
nand NAND3 (N1200, N1182, N141, N197);
buf BUF1 (N1201, N1197);
or OR4 (N1202, N1198, N756, N725, N128);
nand NAND3 (N1203, N1191, N725, N456);
nor NOR3 (N1204, N1199, N606, N1046);
or OR2 (N1205, N1201, N454);
not NOT1 (N1206, N1202);
nand NAND3 (N1207, N1189, N145, N208);
buf BUF1 (N1208, N1165);
nand NAND4 (N1209, N1208, N141, N719, N1125);
not NOT1 (N1210, N1205);
xor XOR2 (N1211, N1209, N678);
xor XOR2 (N1212, N1210, N372);
nand NAND2 (N1213, N1204, N340);
and AND2 (N1214, N1211, N520);
not NOT1 (N1215, N1200);
nand NAND2 (N1216, N1214, N343);
nand NAND3 (N1217, N1216, N577, N299);
and AND4 (N1218, N1217, N446, N1042, N580);
and AND2 (N1219, N1203, N245);
nor NOR3 (N1220, N1215, N23, N992);
buf BUF1 (N1221, N1218);
nor NOR4 (N1222, N1196, N338, N1071, N184);
or OR4 (N1223, N1221, N50, N767, N102);
or OR2 (N1224, N1219, N901);
nand NAND2 (N1225, N1223, N613);
not NOT1 (N1226, N1206);
nor NOR2 (N1227, N1194, N755);
or OR2 (N1228, N1224, N540);
and AND3 (N1229, N1226, N751, N81);
nor NOR3 (N1230, N1222, N94, N773);
not NOT1 (N1231, N1220);
buf BUF1 (N1232, N1229);
buf BUF1 (N1233, N1227);
nand NAND3 (N1234, N1231, N568, N1082);
not NOT1 (N1235, N1192);
nand NAND2 (N1236, N1213, N1135);
nand NAND2 (N1237, N1233, N571);
or OR4 (N1238, N1230, N982, N1041, N999);
buf BUF1 (N1239, N1234);
nand NAND3 (N1240, N1232, N1042, N668);
nand NAND2 (N1241, N1235, N1059);
xor XOR2 (N1242, N1237, N1200);
buf BUF1 (N1243, N1241);
xor XOR2 (N1244, N1239, N265);
and AND2 (N1245, N1236, N439);
buf BUF1 (N1246, N1228);
xor XOR2 (N1247, N1246, N1063);
buf BUF1 (N1248, N1247);
xor XOR2 (N1249, N1248, N560);
not NOT1 (N1250, N1242);
nand NAND4 (N1251, N1212, N67, N860, N192);
xor XOR2 (N1252, N1251, N707);
xor XOR2 (N1253, N1245, N710);
or OR4 (N1254, N1243, N773, N1071, N60);
or OR3 (N1255, N1252, N409, N424);
not NOT1 (N1256, N1254);
nor NOR3 (N1257, N1250, N1088, N981);
or OR4 (N1258, N1256, N945, N747, N1142);
and AND4 (N1259, N1257, N24, N527, N1070);
nand NAND3 (N1260, N1253, N481, N634);
and AND2 (N1261, N1240, N455);
not NOT1 (N1262, N1258);
not NOT1 (N1263, N1262);
or OR3 (N1264, N1225, N515, N718);
and AND3 (N1265, N1260, N716, N778);
nor NOR2 (N1266, N1244, N586);
buf BUF1 (N1267, N1265);
and AND2 (N1268, N1255, N378);
and AND4 (N1269, N1266, N855, N1009, N449);
or OR4 (N1270, N1269, N1007, N21, N810);
or OR2 (N1271, N1263, N1226);
buf BUF1 (N1272, N1259);
nor NOR2 (N1273, N1264, N813);
not NOT1 (N1274, N1249);
nor NOR2 (N1275, N1268, N172);
not NOT1 (N1276, N1267);
nor NOR3 (N1277, N1271, N25, N956);
xor XOR2 (N1278, N1207, N199);
nand NAND4 (N1279, N1276, N1021, N1128, N133);
nand NAND4 (N1280, N1272, N1254, N749, N16);
xor XOR2 (N1281, N1270, N7);
buf BUF1 (N1282, N1275);
buf BUF1 (N1283, N1277);
or OR3 (N1284, N1282, N614, N239);
nor NOR4 (N1285, N1274, N638, N928, N751);
nand NAND2 (N1286, N1285, N386);
nand NAND3 (N1287, N1283, N168, N69);
and AND3 (N1288, N1281, N156, N151);
buf BUF1 (N1289, N1288);
and AND3 (N1290, N1278, N59, N473);
nand NAND3 (N1291, N1287, N293, N470);
nand NAND3 (N1292, N1284, N30, N280);
and AND2 (N1293, N1291, N745);
and AND3 (N1294, N1238, N26, N1100);
nor NOR2 (N1295, N1280, N310);
or OR4 (N1296, N1286, N149, N1260, N1129);
nor NOR2 (N1297, N1261, N43);
nand NAND3 (N1298, N1289, N1279, N704);
buf BUF1 (N1299, N1025);
nor NOR2 (N1300, N1273, N1096);
buf BUF1 (N1301, N1290);
buf BUF1 (N1302, N1301);
nor NOR4 (N1303, N1293, N1032, N126, N959);
or OR2 (N1304, N1302, N566);
xor XOR2 (N1305, N1295, N293);
nand NAND2 (N1306, N1304, N352);
xor XOR2 (N1307, N1292, N1195);
nand NAND4 (N1308, N1299, N280, N344, N82);
nor NOR3 (N1309, N1294, N1052, N916);
not NOT1 (N1310, N1300);
xor XOR2 (N1311, N1303, N993);
or OR2 (N1312, N1298, N414);
nand NAND3 (N1313, N1305, N1155, N1220);
buf BUF1 (N1314, N1309);
xor XOR2 (N1315, N1307, N270);
nor NOR4 (N1316, N1312, N900, N1101, N929);
nand NAND2 (N1317, N1311, N764);
buf BUF1 (N1318, N1315);
xor XOR2 (N1319, N1313, N499);
and AND4 (N1320, N1319, N495, N659, N1317);
not NOT1 (N1321, N688);
or OR4 (N1322, N1318, N285, N1151, N79);
nand NAND2 (N1323, N1306, N598);
buf BUF1 (N1324, N1323);
nor NOR4 (N1325, N1316, N577, N46, N909);
not NOT1 (N1326, N1310);
or OR3 (N1327, N1308, N427, N136);
or OR3 (N1328, N1297, N373, N340);
nor NOR3 (N1329, N1296, N174, N501);
nand NAND2 (N1330, N1321, N113);
xor XOR2 (N1331, N1328, N111);
nor NOR4 (N1332, N1327, N973, N991, N803);
or OR4 (N1333, N1325, N509, N657, N689);
xor XOR2 (N1334, N1322, N325);
buf BUF1 (N1335, N1329);
nor NOR2 (N1336, N1334, N1331);
nor NOR4 (N1337, N237, N126, N1029, N137);
and AND3 (N1338, N1332, N754, N393);
not NOT1 (N1339, N1314);
not NOT1 (N1340, N1324);
xor XOR2 (N1341, N1330, N1044);
and AND3 (N1342, N1339, N1245, N853);
nor NOR4 (N1343, N1336, N526, N1191, N506);
not NOT1 (N1344, N1333);
nor NOR2 (N1345, N1341, N557);
nand NAND3 (N1346, N1335, N763, N518);
xor XOR2 (N1347, N1320, N958);
not NOT1 (N1348, N1337);
and AND3 (N1349, N1340, N255, N262);
buf BUF1 (N1350, N1342);
xor XOR2 (N1351, N1348, N36);
buf BUF1 (N1352, N1346);
nand NAND4 (N1353, N1344, N724, N560, N1130);
xor XOR2 (N1354, N1349, N1254);
xor XOR2 (N1355, N1354, N319);
or OR2 (N1356, N1353, N572);
and AND3 (N1357, N1343, N452, N95);
or OR2 (N1358, N1356, N1212);
xor XOR2 (N1359, N1352, N1194);
and AND2 (N1360, N1350, N966);
and AND4 (N1361, N1355, N284, N1028, N1261);
nand NAND4 (N1362, N1359, N664, N220, N822);
nor NOR3 (N1363, N1338, N632, N317);
and AND4 (N1364, N1362, N1143, N1161, N899);
or OR3 (N1365, N1363, N682, N449);
or OR2 (N1366, N1361, N1066);
and AND4 (N1367, N1326, N1243, N1331, N983);
not NOT1 (N1368, N1365);
xor XOR2 (N1369, N1345, N265);
buf BUF1 (N1370, N1357);
nor NOR3 (N1371, N1370, N750, N1039);
nand NAND2 (N1372, N1360, N116);
nor NOR3 (N1373, N1368, N356, N1170);
nand NAND4 (N1374, N1351, N477, N680, N761);
xor XOR2 (N1375, N1366, N1045);
or OR4 (N1376, N1374, N1340, N1095, N1262);
xor XOR2 (N1377, N1369, N783);
nor NOR3 (N1378, N1376, N408, N247);
nand NAND3 (N1379, N1367, N243, N11);
buf BUF1 (N1380, N1347);
xor XOR2 (N1381, N1372, N1114);
or OR4 (N1382, N1375, N54, N761, N893);
buf BUF1 (N1383, N1364);
or OR2 (N1384, N1381, N445);
and AND3 (N1385, N1373, N771, N883);
and AND3 (N1386, N1377, N1260, N1128);
buf BUF1 (N1387, N1380);
and AND2 (N1388, N1385, N1235);
nor NOR2 (N1389, N1387, N1215);
buf BUF1 (N1390, N1384);
buf BUF1 (N1391, N1358);
xor XOR2 (N1392, N1388, N365);
or OR2 (N1393, N1382, N636);
or OR2 (N1394, N1386, N128);
and AND3 (N1395, N1371, N57, N1040);
xor XOR2 (N1396, N1383, N269);
not NOT1 (N1397, N1379);
or OR3 (N1398, N1394, N1003, N397);
buf BUF1 (N1399, N1391);
nor NOR3 (N1400, N1396, N224, N289);
nand NAND4 (N1401, N1392, N167, N980, N105);
and AND4 (N1402, N1399, N400, N262, N891);
nand NAND4 (N1403, N1401, N818, N511, N405);
buf BUF1 (N1404, N1378);
buf BUF1 (N1405, N1402);
nor NOR4 (N1406, N1404, N1060, N1348, N1133);
nand NAND2 (N1407, N1390, N480);
and AND2 (N1408, N1398, N354);
buf BUF1 (N1409, N1389);
buf BUF1 (N1410, N1393);
xor XOR2 (N1411, N1408, N463);
nand NAND4 (N1412, N1407, N536, N1174, N275);
xor XOR2 (N1413, N1395, N404);
xor XOR2 (N1414, N1400, N439);
nand NAND3 (N1415, N1412, N241, N292);
nor NOR2 (N1416, N1403, N582);
nor NOR3 (N1417, N1415, N444, N525);
or OR3 (N1418, N1411, N748, N1348);
buf BUF1 (N1419, N1413);
nor NOR4 (N1420, N1417, N1051, N586, N702);
or OR4 (N1421, N1410, N514, N34, N864);
xor XOR2 (N1422, N1418, N1211);
buf BUF1 (N1423, N1409);
or OR2 (N1424, N1420, N560);
nand NAND2 (N1425, N1416, N537);
nor NOR2 (N1426, N1414, N820);
xor XOR2 (N1427, N1423, N844);
not NOT1 (N1428, N1422);
xor XOR2 (N1429, N1421, N1398);
not NOT1 (N1430, N1425);
and AND3 (N1431, N1430, N1253, N498);
xor XOR2 (N1432, N1424, N948);
xor XOR2 (N1433, N1432, N1376);
nor NOR2 (N1434, N1433, N833);
and AND3 (N1435, N1426, N342, N1390);
xor XOR2 (N1436, N1406, N259);
nor NOR4 (N1437, N1405, N1072, N1204, N452);
xor XOR2 (N1438, N1437, N997);
and AND2 (N1439, N1431, N376);
nand NAND2 (N1440, N1435, N1168);
nand NAND3 (N1441, N1439, N422, N109);
xor XOR2 (N1442, N1440, N77);
and AND4 (N1443, N1436, N1377, N636, N807);
not NOT1 (N1444, N1434);
xor XOR2 (N1445, N1419, N999);
xor XOR2 (N1446, N1443, N726);
and AND2 (N1447, N1442, N1069);
not NOT1 (N1448, N1444);
nor NOR4 (N1449, N1397, N169, N614, N1310);
and AND4 (N1450, N1441, N677, N11, N676);
or OR2 (N1451, N1427, N537);
not NOT1 (N1452, N1428);
not NOT1 (N1453, N1445);
buf BUF1 (N1454, N1453);
and AND2 (N1455, N1450, N292);
buf BUF1 (N1456, N1451);
or OR3 (N1457, N1447, N1330, N1156);
not NOT1 (N1458, N1452);
not NOT1 (N1459, N1455);
or OR2 (N1460, N1429, N911);
nand NAND3 (N1461, N1454, N1355, N484);
or OR3 (N1462, N1449, N1347, N672);
buf BUF1 (N1463, N1457);
nor NOR3 (N1464, N1460, N199, N669);
nand NAND2 (N1465, N1456, N17);
xor XOR2 (N1466, N1438, N435);
buf BUF1 (N1467, N1463);
buf BUF1 (N1468, N1466);
nor NOR4 (N1469, N1448, N1297, N430, N191);
or OR3 (N1470, N1467, N1256, N787);
not NOT1 (N1471, N1458);
buf BUF1 (N1472, N1469);
nor NOR2 (N1473, N1472, N1006);
and AND2 (N1474, N1465, N305);
xor XOR2 (N1475, N1461, N289);
buf BUF1 (N1476, N1464);
not NOT1 (N1477, N1475);
nor NOR3 (N1478, N1468, N1367, N68);
not NOT1 (N1479, N1478);
and AND3 (N1480, N1479, N260, N1126);
nand NAND3 (N1481, N1462, N15, N987);
and AND2 (N1482, N1476, N1407);
buf BUF1 (N1483, N1471);
xor XOR2 (N1484, N1446, N557);
nand NAND4 (N1485, N1480, N217, N1383, N915);
not NOT1 (N1486, N1481);
nor NOR3 (N1487, N1484, N1270, N811);
or OR3 (N1488, N1485, N149, N1111);
nor NOR2 (N1489, N1488, N1138);
not NOT1 (N1490, N1470);
nor NOR4 (N1491, N1486, N1243, N1124, N805);
and AND4 (N1492, N1489, N249, N753, N444);
or OR2 (N1493, N1487, N596);
not NOT1 (N1494, N1459);
not NOT1 (N1495, N1494);
xor XOR2 (N1496, N1473, N1094);
not NOT1 (N1497, N1477);
and AND2 (N1498, N1497, N748);
nand NAND2 (N1499, N1491, N202);
nor NOR2 (N1500, N1490, N453);
nor NOR4 (N1501, N1495, N68, N401, N293);
xor XOR2 (N1502, N1498, N429);
and AND4 (N1503, N1474, N224, N1148, N406);
buf BUF1 (N1504, N1482);
and AND2 (N1505, N1503, N576);
and AND3 (N1506, N1501, N1249, N154);
and AND4 (N1507, N1492, N809, N637, N1152);
not NOT1 (N1508, N1483);
and AND2 (N1509, N1493, N964);
and AND2 (N1510, N1509, N1450);
nor NOR2 (N1511, N1502, N1085);
nand NAND4 (N1512, N1508, N1311, N543, N1144);
not NOT1 (N1513, N1510);
not NOT1 (N1514, N1512);
or OR4 (N1515, N1511, N643, N1492, N640);
or OR3 (N1516, N1515, N659, N1006);
nand NAND2 (N1517, N1513, N1071);
or OR2 (N1518, N1499, N1010);
buf BUF1 (N1519, N1505);
or OR2 (N1520, N1516, N1248);
not NOT1 (N1521, N1500);
buf BUF1 (N1522, N1504);
nand NAND2 (N1523, N1520, N466);
nand NAND4 (N1524, N1521, N1353, N1201, N241);
nor NOR4 (N1525, N1523, N955, N1421, N141);
xor XOR2 (N1526, N1519, N1408);
and AND4 (N1527, N1526, N1092, N452, N1146);
and AND4 (N1528, N1506, N793, N1181, N1292);
or OR3 (N1529, N1514, N1434, N1304);
nand NAND4 (N1530, N1529, N923, N1191, N522);
nor NOR3 (N1531, N1524, N544, N526);
and AND3 (N1532, N1496, N735, N592);
nor NOR4 (N1533, N1517, N1407, N1392, N1234);
and AND3 (N1534, N1507, N1469, N913);
xor XOR2 (N1535, N1522, N212);
xor XOR2 (N1536, N1518, N650);
nand NAND4 (N1537, N1525, N617, N90, N123);
xor XOR2 (N1538, N1527, N1529);
nor NOR2 (N1539, N1535, N1349);
or OR2 (N1540, N1536, N25);
buf BUF1 (N1541, N1538);
and AND3 (N1542, N1530, N1533, N79);
nor NOR2 (N1543, N1063, N516);
nand NAND4 (N1544, N1532, N556, N824, N964);
nand NAND2 (N1545, N1528, N1535);
and AND3 (N1546, N1531, N1129, N1082);
not NOT1 (N1547, N1540);
xor XOR2 (N1548, N1543, N1128);
and AND4 (N1549, N1548, N568, N1506, N1207);
and AND3 (N1550, N1542, N717, N701);
not NOT1 (N1551, N1534);
or OR2 (N1552, N1549, N1274);
xor XOR2 (N1553, N1545, N693);
and AND4 (N1554, N1553, N550, N1065, N1486);
buf BUF1 (N1555, N1552);
and AND3 (N1556, N1555, N994, N1002);
and AND4 (N1557, N1537, N522, N1070, N588);
nor NOR4 (N1558, N1544, N87, N254, N482);
and AND4 (N1559, N1554, N302, N1147, N309);
nand NAND4 (N1560, N1559, N1527, N1294, N1342);
buf BUF1 (N1561, N1560);
or OR4 (N1562, N1547, N292, N351, N1346);
nand NAND4 (N1563, N1539, N377, N735, N1081);
or OR4 (N1564, N1546, N912, N538, N694);
nand NAND3 (N1565, N1551, N941, N888);
or OR4 (N1566, N1564, N866, N1384, N1462);
nand NAND3 (N1567, N1563, N17, N43);
nor NOR2 (N1568, N1541, N1501);
nor NOR3 (N1569, N1566, N1447, N801);
and AND3 (N1570, N1561, N1461, N39);
not NOT1 (N1571, N1569);
buf BUF1 (N1572, N1562);
or OR4 (N1573, N1550, N367, N496, N188);
nor NOR2 (N1574, N1556, N1097);
and AND3 (N1575, N1571, N173, N1485);
buf BUF1 (N1576, N1573);
nor NOR2 (N1577, N1575, N152);
not NOT1 (N1578, N1557);
xor XOR2 (N1579, N1577, N892);
and AND3 (N1580, N1558, N1546, N910);
not NOT1 (N1581, N1578);
and AND3 (N1582, N1567, N1506, N1227);
not NOT1 (N1583, N1582);
nand NAND2 (N1584, N1568, N911);
or OR4 (N1585, N1565, N125, N1564, N689);
xor XOR2 (N1586, N1570, N894);
xor XOR2 (N1587, N1586, N341);
nor NOR3 (N1588, N1585, N1004, N292);
or OR2 (N1589, N1579, N1508);
not NOT1 (N1590, N1587);
or OR2 (N1591, N1589, N1328);
not NOT1 (N1592, N1591);
and AND4 (N1593, N1590, N413, N934, N624);
not NOT1 (N1594, N1576);
buf BUF1 (N1595, N1574);
not NOT1 (N1596, N1594);
nand NAND3 (N1597, N1588, N805, N704);
and AND2 (N1598, N1593, N178);
and AND3 (N1599, N1592, N1206, N159);
nand NAND4 (N1600, N1572, N669, N93, N1495);
xor XOR2 (N1601, N1597, N434);
xor XOR2 (N1602, N1600, N1104);
and AND2 (N1603, N1581, N1168);
not NOT1 (N1604, N1599);
or OR4 (N1605, N1595, N1480, N895, N1343);
nand NAND4 (N1606, N1584, N1038, N202, N586);
nor NOR3 (N1607, N1603, N1468, N18);
xor XOR2 (N1608, N1605, N531);
nor NOR2 (N1609, N1580, N196);
xor XOR2 (N1610, N1604, N1433);
xor XOR2 (N1611, N1596, N1109);
xor XOR2 (N1612, N1607, N387);
and AND4 (N1613, N1610, N712, N53, N1044);
nor NOR3 (N1614, N1608, N812, N923);
or OR2 (N1615, N1606, N1143);
buf BUF1 (N1616, N1611);
buf BUF1 (N1617, N1602);
and AND2 (N1618, N1598, N1590);
xor XOR2 (N1619, N1583, N1130);
not NOT1 (N1620, N1609);
or OR4 (N1621, N1615, N706, N420, N1275);
buf BUF1 (N1622, N1612);
buf BUF1 (N1623, N1622);
not NOT1 (N1624, N1621);
and AND3 (N1625, N1614, N385, N1197);
and AND2 (N1626, N1620, N1461);
and AND3 (N1627, N1617, N269, N1545);
xor XOR2 (N1628, N1626, N1180);
or OR4 (N1629, N1619, N1607, N248, N676);
or OR4 (N1630, N1616, N597, N762, N236);
or OR3 (N1631, N1618, N1617, N1420);
nand NAND2 (N1632, N1625, N296);
nor NOR2 (N1633, N1601, N1103);
not NOT1 (N1634, N1632);
or OR2 (N1635, N1624, N1138);
and AND2 (N1636, N1628, N27);
and AND4 (N1637, N1630, N353, N114, N1323);
nand NAND2 (N1638, N1623, N586);
and AND4 (N1639, N1633, N1153, N174, N1271);
nand NAND2 (N1640, N1631, N1241);
nor NOR2 (N1641, N1639, N822);
nor NOR4 (N1642, N1627, N368, N433, N704);
and AND3 (N1643, N1638, N248, N7);
buf BUF1 (N1644, N1642);
nand NAND2 (N1645, N1635, N542);
and AND3 (N1646, N1636, N1394, N245);
nor NOR3 (N1647, N1613, N1619, N1084);
nand NAND3 (N1648, N1644, N1500, N106);
nor NOR3 (N1649, N1629, N184, N937);
nor NOR4 (N1650, N1649, N876, N698, N219);
not NOT1 (N1651, N1641);
not NOT1 (N1652, N1640);
nor NOR2 (N1653, N1646, N1013);
nand NAND2 (N1654, N1645, N1509);
xor XOR2 (N1655, N1634, N566);
not NOT1 (N1656, N1643);
nand NAND3 (N1657, N1647, N1219, N902);
not NOT1 (N1658, N1653);
and AND3 (N1659, N1655, N95, N1602);
xor XOR2 (N1660, N1654, N361);
not NOT1 (N1661, N1657);
not NOT1 (N1662, N1648);
nand NAND3 (N1663, N1651, N578, N983);
nand NAND4 (N1664, N1661, N917, N919, N1129);
nor NOR4 (N1665, N1637, N85, N1143, N1113);
and AND2 (N1666, N1662, N408);
buf BUF1 (N1667, N1650);
buf BUF1 (N1668, N1658);
nand NAND4 (N1669, N1667, N457, N444, N1271);
buf BUF1 (N1670, N1668);
or OR3 (N1671, N1670, N516, N1039);
nand NAND4 (N1672, N1663, N161, N1213, N64);
nand NAND2 (N1673, N1671, N153);
and AND3 (N1674, N1673, N198, N1243);
nand NAND4 (N1675, N1672, N689, N1493, N163);
buf BUF1 (N1676, N1660);
xor XOR2 (N1677, N1665, N1222);
not NOT1 (N1678, N1669);
nor NOR2 (N1679, N1678, N980);
not NOT1 (N1680, N1674);
not NOT1 (N1681, N1666);
not NOT1 (N1682, N1664);
buf BUF1 (N1683, N1675);
not NOT1 (N1684, N1683);
xor XOR2 (N1685, N1681, N615);
nand NAND3 (N1686, N1685, N877, N55);
nor NOR4 (N1687, N1684, N1068, N437, N285);
nand NAND3 (N1688, N1680, N474, N1252);
nor NOR4 (N1689, N1686, N1072, N837, N101);
not NOT1 (N1690, N1656);
and AND3 (N1691, N1652, N1404, N317);
not NOT1 (N1692, N1688);
or OR2 (N1693, N1691, N692);
xor XOR2 (N1694, N1687, N1328);
or OR3 (N1695, N1676, N813, N1689);
not NOT1 (N1696, N1554);
xor XOR2 (N1697, N1659, N937);
not NOT1 (N1698, N1690);
not NOT1 (N1699, N1693);
or OR4 (N1700, N1697, N495, N265, N1614);
or OR3 (N1701, N1696, N1004, N883);
xor XOR2 (N1702, N1701, N41);
or OR4 (N1703, N1679, N1433, N1173, N102);
buf BUF1 (N1704, N1698);
nand NAND4 (N1705, N1682, N1548, N457, N552);
nor NOR4 (N1706, N1694, N1444, N1130, N1579);
and AND3 (N1707, N1692, N1232, N1686);
nand NAND3 (N1708, N1706, N167, N533);
buf BUF1 (N1709, N1699);
or OR4 (N1710, N1709, N332, N529, N1347);
nand NAND2 (N1711, N1677, N481);
nor NOR3 (N1712, N1707, N1376, N52);
not NOT1 (N1713, N1704);
buf BUF1 (N1714, N1712);
xor XOR2 (N1715, N1710, N1696);
or OR3 (N1716, N1702, N1652, N1260);
not NOT1 (N1717, N1703);
not NOT1 (N1718, N1714);
and AND2 (N1719, N1713, N1596);
nand NAND4 (N1720, N1719, N49, N114, N1645);
nor NOR3 (N1721, N1700, N1424, N1031);
and AND3 (N1722, N1711, N411, N1396);
xor XOR2 (N1723, N1717, N79);
and AND3 (N1724, N1715, N1263, N920);
buf BUF1 (N1725, N1695);
not NOT1 (N1726, N1708);
xor XOR2 (N1727, N1723, N897);
buf BUF1 (N1728, N1716);
or OR3 (N1729, N1727, N562, N766);
nand NAND3 (N1730, N1726, N1177, N6);
not NOT1 (N1731, N1722);
xor XOR2 (N1732, N1721, N742);
and AND3 (N1733, N1731, N1384, N1348);
buf BUF1 (N1734, N1733);
nand NAND4 (N1735, N1729, N834, N91, N1665);
or OR3 (N1736, N1705, N432, N1564);
nand NAND2 (N1737, N1724, N1503);
xor XOR2 (N1738, N1730, N917);
buf BUF1 (N1739, N1728);
or OR3 (N1740, N1739, N1394, N1354);
buf BUF1 (N1741, N1735);
buf BUF1 (N1742, N1718);
buf BUF1 (N1743, N1741);
xor XOR2 (N1744, N1737, N1348);
nand NAND3 (N1745, N1743, N575, N3);
xor XOR2 (N1746, N1745, N913);
nand NAND2 (N1747, N1742, N660);
nor NOR4 (N1748, N1725, N531, N991, N154);
nor NOR3 (N1749, N1734, N1701, N692);
nand NAND2 (N1750, N1748, N534);
or OR2 (N1751, N1744, N840);
nor NOR3 (N1752, N1750, N534, N710);
or OR3 (N1753, N1740, N1009, N131);
nor NOR4 (N1754, N1747, N456, N786, N62);
not NOT1 (N1755, N1754);
nand NAND4 (N1756, N1753, N1015, N1586, N1057);
nor NOR4 (N1757, N1720, N937, N90, N501);
and AND3 (N1758, N1757, N1319, N99);
not NOT1 (N1759, N1758);
xor XOR2 (N1760, N1759, N1264);
not NOT1 (N1761, N1732);
and AND3 (N1762, N1736, N862, N655);
nand NAND3 (N1763, N1749, N1114, N298);
not NOT1 (N1764, N1755);
not NOT1 (N1765, N1738);
buf BUF1 (N1766, N1752);
or OR3 (N1767, N1765, N375, N953);
or OR4 (N1768, N1761, N1234, N858, N190);
xor XOR2 (N1769, N1763, N1627);
or OR4 (N1770, N1760, N1512, N903, N513);
or OR3 (N1771, N1766, N1295, N854);
or OR2 (N1772, N1751, N716);
nor NOR3 (N1773, N1767, N874, N129);
or OR4 (N1774, N1762, N1754, N1539, N105);
nand NAND4 (N1775, N1764, N1425, N1610, N1);
nand NAND2 (N1776, N1774, N1565);
nor NOR4 (N1777, N1746, N1678, N723, N187);
and AND4 (N1778, N1773, N1701, N1380, N1212);
nand NAND2 (N1779, N1776, N749);
nor NOR4 (N1780, N1778, N520, N328, N195);
buf BUF1 (N1781, N1768);
nand NAND2 (N1782, N1777, N1442);
not NOT1 (N1783, N1779);
buf BUF1 (N1784, N1756);
or OR4 (N1785, N1782, N1692, N61, N1450);
not NOT1 (N1786, N1783);
or OR3 (N1787, N1786, N938, N1410);
not NOT1 (N1788, N1775);
not NOT1 (N1789, N1788);
nor NOR4 (N1790, N1784, N889, N109, N526);
buf BUF1 (N1791, N1781);
nor NOR4 (N1792, N1789, N705, N1342, N36);
nor NOR3 (N1793, N1771, N1268, N608);
nor NOR2 (N1794, N1791, N434);
nor NOR4 (N1795, N1772, N732, N1696, N799);
or OR2 (N1796, N1795, N814);
nor NOR2 (N1797, N1793, N1296);
not NOT1 (N1798, N1797);
or OR3 (N1799, N1790, N1400, N1129);
not NOT1 (N1800, N1792);
xor XOR2 (N1801, N1794, N339);
or OR2 (N1802, N1785, N972);
nand NAND4 (N1803, N1798, N907, N211, N85);
nand NAND3 (N1804, N1803, N49, N278);
or OR2 (N1805, N1804, N874);
or OR3 (N1806, N1800, N119, N161);
not NOT1 (N1807, N1770);
or OR3 (N1808, N1799, N1002, N1768);
or OR2 (N1809, N1780, N986);
not NOT1 (N1810, N1808);
nand NAND2 (N1811, N1805, N1186);
not NOT1 (N1812, N1802);
and AND4 (N1813, N1801, N1531, N1188, N722);
or OR3 (N1814, N1809, N89, N495);
xor XOR2 (N1815, N1787, N336);
or OR2 (N1816, N1813, N1780);
buf BUF1 (N1817, N1812);
buf BUF1 (N1818, N1807);
xor XOR2 (N1819, N1816, N469);
and AND2 (N1820, N1819, N1559);
not NOT1 (N1821, N1810);
not NOT1 (N1822, N1811);
or OR3 (N1823, N1821, N1465, N725);
nor NOR2 (N1824, N1823, N120);
xor XOR2 (N1825, N1814, N1327);
and AND2 (N1826, N1822, N1126);
buf BUF1 (N1827, N1769);
or OR2 (N1828, N1820, N926);
or OR4 (N1829, N1826, N159, N677, N344);
buf BUF1 (N1830, N1824);
and AND2 (N1831, N1806, N351);
nor NOR2 (N1832, N1827, N1040);
nor NOR2 (N1833, N1818, N1628);
or OR3 (N1834, N1817, N880, N1586);
and AND2 (N1835, N1825, N1663);
not NOT1 (N1836, N1830);
xor XOR2 (N1837, N1834, N1137);
xor XOR2 (N1838, N1836, N1184);
xor XOR2 (N1839, N1796, N618);
or OR3 (N1840, N1828, N585, N665);
and AND3 (N1841, N1837, N40, N404);
nor NOR4 (N1842, N1832, N1397, N975, N1318);
and AND2 (N1843, N1842, N908);
nor NOR2 (N1844, N1831, N1654);
nor NOR3 (N1845, N1840, N162, N576);
xor XOR2 (N1846, N1839, N905);
xor XOR2 (N1847, N1845, N1204);
nand NAND4 (N1848, N1841, N1196, N622, N825);
not NOT1 (N1849, N1838);
not NOT1 (N1850, N1835);
nand NAND4 (N1851, N1844, N747, N456, N46);
xor XOR2 (N1852, N1829, N83);
or OR4 (N1853, N1848, N469, N139, N205);
nor NOR2 (N1854, N1852, N611);
nand NAND2 (N1855, N1853, N1582);
nand NAND3 (N1856, N1855, N1386, N929);
and AND2 (N1857, N1849, N994);
or OR2 (N1858, N1854, N802);
buf BUF1 (N1859, N1856);
and AND2 (N1860, N1851, N73);
and AND4 (N1861, N1858, N446, N391, N664);
nand NAND3 (N1862, N1860, N592, N1395);
buf BUF1 (N1863, N1861);
buf BUF1 (N1864, N1815);
buf BUF1 (N1865, N1857);
xor XOR2 (N1866, N1864, N1034);
xor XOR2 (N1867, N1862, N959);
and AND3 (N1868, N1865, N1411, N282);
xor XOR2 (N1869, N1846, N1126);
xor XOR2 (N1870, N1863, N949);
xor XOR2 (N1871, N1867, N1692);
or OR4 (N1872, N1833, N1536, N1551, N681);
not NOT1 (N1873, N1859);
xor XOR2 (N1874, N1850, N32);
nor NOR2 (N1875, N1872, N952);
buf BUF1 (N1876, N1874);
nor NOR2 (N1877, N1876, N409);
xor XOR2 (N1878, N1866, N995);
or OR4 (N1879, N1871, N732, N1427, N910);
nor NOR2 (N1880, N1879, N718);
or OR3 (N1881, N1875, N795, N1795);
xor XOR2 (N1882, N1843, N1207);
or OR2 (N1883, N1873, N165);
or OR2 (N1884, N1868, N1157);
nand NAND2 (N1885, N1878, N216);
xor XOR2 (N1886, N1885, N1445);
or OR4 (N1887, N1877, N1291, N882, N1518);
and AND4 (N1888, N1881, N1436, N715, N263);
and AND2 (N1889, N1882, N361);
not NOT1 (N1890, N1869);
xor XOR2 (N1891, N1883, N540);
or OR2 (N1892, N1889, N50);
not NOT1 (N1893, N1884);
not NOT1 (N1894, N1880);
or OR3 (N1895, N1891, N1680, N317);
or OR4 (N1896, N1893, N1656, N511, N765);
nor NOR4 (N1897, N1888, N1524, N835, N1399);
and AND4 (N1898, N1870, N46, N1160, N795);
xor XOR2 (N1899, N1886, N424);
or OR4 (N1900, N1896, N308, N1037, N1064);
nor NOR4 (N1901, N1890, N985, N748, N1537);
and AND2 (N1902, N1901, N1161);
and AND2 (N1903, N1902, N1570);
nand NAND2 (N1904, N1895, N1360);
nand NAND3 (N1905, N1898, N1428, N709);
xor XOR2 (N1906, N1905, N31);
buf BUF1 (N1907, N1899);
xor XOR2 (N1908, N1894, N852);
not NOT1 (N1909, N1907);
nand NAND3 (N1910, N1909, N1880, N623);
not NOT1 (N1911, N1904);
nor NOR2 (N1912, N1906, N201);
not NOT1 (N1913, N1900);
xor XOR2 (N1914, N1892, N769);
and AND2 (N1915, N1911, N1293);
buf BUF1 (N1916, N1912);
nor NOR3 (N1917, N1910, N262, N1065);
buf BUF1 (N1918, N1897);
xor XOR2 (N1919, N1918, N835);
or OR3 (N1920, N1919, N1510, N1802);
nor NOR4 (N1921, N1913, N49, N1389, N1780);
or OR2 (N1922, N1916, N1587);
nand NAND2 (N1923, N1921, N419);
and AND3 (N1924, N1920, N1369, N1548);
nor NOR4 (N1925, N1924, N1321, N417, N51);
not NOT1 (N1926, N1923);
buf BUF1 (N1927, N1926);
nor NOR3 (N1928, N1922, N1099, N764);
or OR4 (N1929, N1925, N669, N941, N1310);
not NOT1 (N1930, N1928);
or OR4 (N1931, N1914, N405, N167, N1244);
and AND3 (N1932, N1908, N836, N1439);
buf BUF1 (N1933, N1903);
nor NOR2 (N1934, N1931, N344);
nand NAND2 (N1935, N1929, N1305);
and AND2 (N1936, N1930, N960);
nor NOR4 (N1937, N1936, N487, N1829, N144);
and AND3 (N1938, N1932, N874, N286);
buf BUF1 (N1939, N1933);
xor XOR2 (N1940, N1939, N1123);
nand NAND2 (N1941, N1940, N300);
and AND4 (N1942, N1915, N1204, N4, N1059);
nand NAND2 (N1943, N1937, N799);
not NOT1 (N1944, N1935);
xor XOR2 (N1945, N1934, N1077);
and AND3 (N1946, N1917, N262, N1088);
or OR4 (N1947, N1944, N231, N98, N49);
nor NOR3 (N1948, N1887, N1325, N1375);
buf BUF1 (N1949, N1942);
buf BUF1 (N1950, N1847);
xor XOR2 (N1951, N1941, N1754);
buf BUF1 (N1952, N1927);
and AND4 (N1953, N1950, N1264, N1282, N1281);
xor XOR2 (N1954, N1947, N747);
not NOT1 (N1955, N1945);
nor NOR4 (N1956, N1949, N1190, N1792, N1470);
nand NAND4 (N1957, N1938, N304, N241, N28);
not NOT1 (N1958, N1948);
nand NAND4 (N1959, N1952, N1213, N311, N1545);
and AND3 (N1960, N1956, N178, N1925);
buf BUF1 (N1961, N1954);
not NOT1 (N1962, N1946);
not NOT1 (N1963, N1957);
and AND3 (N1964, N1951, N85, N1893);
not NOT1 (N1965, N1960);
not NOT1 (N1966, N1965);
nand NAND2 (N1967, N1955, N802);
and AND3 (N1968, N1958, N721, N452);
not NOT1 (N1969, N1968);
nand NAND2 (N1970, N1963, N1658);
and AND2 (N1971, N1970, N1382);
or OR4 (N1972, N1943, N535, N71, N68);
buf BUF1 (N1973, N1964);
and AND2 (N1974, N1972, N251);
not NOT1 (N1975, N1961);
buf BUF1 (N1976, N1971);
not NOT1 (N1977, N1967);
xor XOR2 (N1978, N1974, N1714);
nor NOR2 (N1979, N1969, N454);
nor NOR3 (N1980, N1977, N1067, N899);
or OR4 (N1981, N1980, N319, N1379, N725);
and AND2 (N1982, N1959, N190);
nand NAND3 (N1983, N1966, N1780, N634);
xor XOR2 (N1984, N1953, N1294);
not NOT1 (N1985, N1973);
xor XOR2 (N1986, N1979, N1608);
nor NOR3 (N1987, N1976, N1149, N45);
buf BUF1 (N1988, N1984);
and AND3 (N1989, N1985, N972, N1132);
nand NAND3 (N1990, N1978, N10, N1967);
not NOT1 (N1991, N1962);
nand NAND2 (N1992, N1989, N936);
nand NAND2 (N1993, N1981, N338);
nand NAND4 (N1994, N1983, N1721, N1514, N522);
buf BUF1 (N1995, N1982);
nor NOR3 (N1996, N1987, N1542, N1851);
not NOT1 (N1997, N1991);
nand NAND4 (N1998, N1986, N1765, N588, N1869);
nand NAND3 (N1999, N1975, N664, N1660);
nand NAND4 (N2000, N1994, N1166, N1719, N948);
nor NOR4 (N2001, N1988, N735, N940, N1430);
nor NOR3 (N2002, N1995, N608, N1818);
buf BUF1 (N2003, N1997);
nand NAND4 (N2004, N1999, N1586, N147, N609);
buf BUF1 (N2005, N2004);
nand NAND2 (N2006, N1993, N468);
not NOT1 (N2007, N1992);
and AND4 (N2008, N2003, N507, N803, N541);
nor NOR3 (N2009, N2007, N803, N226);
buf BUF1 (N2010, N1998);
nand NAND4 (N2011, N1996, N193, N1005, N1210);
or OR3 (N2012, N1990, N355, N312);
xor XOR2 (N2013, N2011, N397);
and AND3 (N2014, N2012, N82, N1717);
buf BUF1 (N2015, N2006);
and AND4 (N2016, N2008, N397, N55, N1748);
or OR2 (N2017, N2009, N770);
nand NAND4 (N2018, N2005, N2004, N174, N1307);
and AND2 (N2019, N2014, N1772);
or OR3 (N2020, N2017, N1431, N1489);
and AND3 (N2021, N2013, N452, N580);
nand NAND3 (N2022, N2010, N1276, N218);
and AND4 (N2023, N2020, N659, N775, N758);
not NOT1 (N2024, N2016);
nor NOR3 (N2025, N2001, N1294, N970);
nand NAND2 (N2026, N2000, N214);
not NOT1 (N2027, N2002);
nand NAND4 (N2028, N2024, N745, N1727, N1080);
buf BUF1 (N2029, N2019);
nand NAND3 (N2030, N2028, N1016, N1038);
not NOT1 (N2031, N2030);
and AND3 (N2032, N2027, N1279, N1785);
and AND3 (N2033, N2026, N1008, N1773);
xor XOR2 (N2034, N2032, N440);
nand NAND4 (N2035, N2029, N483, N365, N1687);
or OR2 (N2036, N2034, N460);
not NOT1 (N2037, N2022);
or OR4 (N2038, N2023, N1743, N229, N1838);
xor XOR2 (N2039, N2036, N743);
or OR4 (N2040, N2031, N709, N1310, N201);
and AND4 (N2041, N2025, N1959, N966, N1185);
or OR2 (N2042, N2035, N295);
not NOT1 (N2043, N2015);
or OR3 (N2044, N2040, N1226, N408);
nand NAND4 (N2045, N2041, N944, N1311, N1017);
or OR2 (N2046, N2042, N1867);
not NOT1 (N2047, N2043);
nand NAND2 (N2048, N2044, N384);
and AND4 (N2049, N2046, N1627, N1955, N220);
buf BUF1 (N2050, N2038);
not NOT1 (N2051, N2047);
xor XOR2 (N2052, N2048, N1507);
nor NOR4 (N2053, N2050, N1714, N456, N1404);
and AND4 (N2054, N2045, N1674, N343, N51);
or OR3 (N2055, N2018, N186, N430);
not NOT1 (N2056, N2054);
buf BUF1 (N2057, N2055);
nand NAND3 (N2058, N2037, N1084, N2014);
nand NAND4 (N2059, N2049, N1096, N1950, N1860);
not NOT1 (N2060, N2052);
nand NAND3 (N2061, N2039, N506, N516);
nor NOR2 (N2062, N2061, N1511);
not NOT1 (N2063, N2056);
or OR2 (N2064, N2021, N2003);
nor NOR3 (N2065, N2033, N268, N107);
not NOT1 (N2066, N2059);
buf BUF1 (N2067, N2063);
or OR2 (N2068, N2066, N1040);
nor NOR4 (N2069, N2053, N1628, N1124, N1927);
not NOT1 (N2070, N2058);
nand NAND2 (N2071, N2057, N1133);
xor XOR2 (N2072, N2067, N1336);
xor XOR2 (N2073, N2065, N1646);
nand NAND4 (N2074, N2062, N95, N1889, N795);
not NOT1 (N2075, N2070);
nor NOR3 (N2076, N2075, N906, N1367);
or OR4 (N2077, N2068, N127, N1435, N505);
xor XOR2 (N2078, N2072, N1649);
not NOT1 (N2079, N2078);
nand NAND3 (N2080, N2077, N178, N50);
buf BUF1 (N2081, N2080);
not NOT1 (N2082, N2081);
nand NAND2 (N2083, N2071, N1770);
buf BUF1 (N2084, N2076);
and AND3 (N2085, N2083, N1396, N1743);
or OR3 (N2086, N2064, N223, N1334);
not NOT1 (N2087, N2073);
nor NOR2 (N2088, N2085, N1105);
nand NAND2 (N2089, N2086, N522);
nor NOR4 (N2090, N2079, N559, N2066, N1019);
not NOT1 (N2091, N2060);
buf BUF1 (N2092, N2051);
xor XOR2 (N2093, N2084, N278);
and AND4 (N2094, N2069, N1095, N982, N2030);
buf BUF1 (N2095, N2090);
nor NOR4 (N2096, N2091, N1361, N273, N681);
and AND3 (N2097, N2082, N1852, N1707);
and AND4 (N2098, N2097, N2016, N1587, N721);
buf BUF1 (N2099, N2092);
or OR4 (N2100, N2095, N206, N1360, N164);
nor NOR2 (N2101, N2074, N1758);
not NOT1 (N2102, N2089);
nand NAND3 (N2103, N2096, N1815, N97);
not NOT1 (N2104, N2098);
nor NOR2 (N2105, N2093, N443);
nand NAND4 (N2106, N2087, N1524, N678, N4);
or OR3 (N2107, N2094, N49, N850);
xor XOR2 (N2108, N2102, N322);
or OR2 (N2109, N2103, N500);
xor XOR2 (N2110, N2088, N496);
not NOT1 (N2111, N2105);
nor NOR2 (N2112, N2107, N2024);
xor XOR2 (N2113, N2108, N495);
and AND4 (N2114, N2106, N1488, N1753, N1010);
not NOT1 (N2115, N2112);
xor XOR2 (N2116, N2099, N430);
and AND4 (N2117, N2115, N740, N1077, N2060);
not NOT1 (N2118, N2100);
xor XOR2 (N2119, N2118, N846);
xor XOR2 (N2120, N2114, N1252);
and AND4 (N2121, N2109, N886, N1236, N1659);
xor XOR2 (N2122, N2121, N931);
or OR3 (N2123, N2111, N148, N1409);
nor NOR2 (N2124, N2122, N1996);
buf BUF1 (N2125, N2113);
xor XOR2 (N2126, N2101, N476);
nor NOR2 (N2127, N2126, N1214);
xor XOR2 (N2128, N2120, N1021);
buf BUF1 (N2129, N2117);
nor NOR3 (N2130, N2104, N852, N1743);
and AND3 (N2131, N2125, N34, N454);
and AND4 (N2132, N2116, N909, N1724, N1772);
nor NOR4 (N2133, N2129, N468, N1770, N405);
not NOT1 (N2134, N2130);
or OR3 (N2135, N2123, N1699, N732);
nand NAND3 (N2136, N2127, N507, N382);
not NOT1 (N2137, N2136);
not NOT1 (N2138, N2124);
nand NAND4 (N2139, N2133, N2029, N1324, N616);
nand NAND4 (N2140, N2134, N844, N340, N1271);
not NOT1 (N2141, N2131);
nor NOR2 (N2142, N2137, N1775);
xor XOR2 (N2143, N2142, N1284);
xor XOR2 (N2144, N2139, N501);
nor NOR3 (N2145, N2135, N1536, N1802);
and AND2 (N2146, N2132, N117);
nand NAND4 (N2147, N2146, N278, N100, N1845);
buf BUF1 (N2148, N2141);
nand NAND2 (N2149, N2148, N565);
or OR4 (N2150, N2149, N372, N483, N538);
or OR3 (N2151, N2128, N371, N570);
xor XOR2 (N2152, N2138, N1328);
not NOT1 (N2153, N2110);
or OR4 (N2154, N2153, N1511, N547, N349);
xor XOR2 (N2155, N2151, N1595);
not NOT1 (N2156, N2155);
not NOT1 (N2157, N2140);
nor NOR4 (N2158, N2156, N2103, N1568, N1769);
or OR2 (N2159, N2147, N649);
and AND3 (N2160, N2145, N1237, N118);
or OR4 (N2161, N2154, N760, N1673, N1863);
and AND4 (N2162, N2143, N1271, N1657, N811);
buf BUF1 (N2163, N2150);
nand NAND3 (N2164, N2157, N1541, N1320);
or OR4 (N2165, N2162, N5, N389, N807);
buf BUF1 (N2166, N2119);
or OR4 (N2167, N2144, N1558, N1769, N458);
not NOT1 (N2168, N2160);
or OR4 (N2169, N2165, N427, N309, N1391);
not NOT1 (N2170, N2167);
nand NAND4 (N2171, N2152, N57, N1820, N1830);
xor XOR2 (N2172, N2158, N278);
not NOT1 (N2173, N2171);
buf BUF1 (N2174, N2173);
buf BUF1 (N2175, N2166);
not NOT1 (N2176, N2172);
buf BUF1 (N2177, N2168);
nor NOR3 (N2178, N2159, N1360, N2119);
nor NOR3 (N2179, N2178, N426, N1345);
nor NOR2 (N2180, N2164, N2153);
not NOT1 (N2181, N2174);
xor XOR2 (N2182, N2179, N1926);
not NOT1 (N2183, N2161);
or OR4 (N2184, N2176, N2086, N705, N1865);
xor XOR2 (N2185, N2184, N482);
not NOT1 (N2186, N2181);
or OR2 (N2187, N2163, N1746);
nor NOR4 (N2188, N2180, N1089, N2018, N1669);
and AND4 (N2189, N2175, N1213, N1905, N1168);
nand NAND4 (N2190, N2187, N554, N1790, N1299);
xor XOR2 (N2191, N2170, N1864);
and AND2 (N2192, N2188, N1801);
and AND2 (N2193, N2189, N1581);
not NOT1 (N2194, N2186);
buf BUF1 (N2195, N2169);
nand NAND2 (N2196, N2185, N1413);
nor NOR2 (N2197, N2195, N701);
not NOT1 (N2198, N2192);
xor XOR2 (N2199, N2197, N1436);
or OR2 (N2200, N2177, N936);
xor XOR2 (N2201, N2190, N1119);
xor XOR2 (N2202, N2196, N666);
nand NAND4 (N2203, N2201, N152, N15, N1157);
xor XOR2 (N2204, N2194, N310);
not NOT1 (N2205, N2191);
xor XOR2 (N2206, N2205, N1180);
nor NOR4 (N2207, N2204, N747, N1428, N521);
nor NOR3 (N2208, N2183, N1487, N1874);
nor NOR3 (N2209, N2208, N1266, N165);
and AND2 (N2210, N2198, N733);
or OR4 (N2211, N2203, N738, N157, N204);
nor NOR2 (N2212, N2206, N924);
not NOT1 (N2213, N2202);
xor XOR2 (N2214, N2212, N910);
buf BUF1 (N2215, N2193);
nor NOR4 (N2216, N2210, N491, N1041, N76);
not NOT1 (N2217, N2214);
and AND2 (N2218, N2199, N1425);
and AND3 (N2219, N2218, N632, N527);
nor NOR3 (N2220, N2211, N185, N1553);
not NOT1 (N2221, N2219);
buf BUF1 (N2222, N2213);
buf BUF1 (N2223, N2222);
not NOT1 (N2224, N2220);
buf BUF1 (N2225, N2223);
nor NOR4 (N2226, N2207, N41, N591, N1216);
buf BUF1 (N2227, N2226);
buf BUF1 (N2228, N2182);
not NOT1 (N2229, N2216);
nor NOR2 (N2230, N2228, N1813);
buf BUF1 (N2231, N2215);
or OR4 (N2232, N2230, N698, N1566, N345);
buf BUF1 (N2233, N2229);
xor XOR2 (N2234, N2200, N1236);
not NOT1 (N2235, N2234);
nor NOR2 (N2236, N2224, N2113);
and AND4 (N2237, N2225, N1020, N1950, N2097);
or OR3 (N2238, N2233, N742, N885);
buf BUF1 (N2239, N2235);
or OR2 (N2240, N2239, N773);
nand NAND3 (N2241, N2209, N1419, N875);
buf BUF1 (N2242, N2237);
xor XOR2 (N2243, N2238, N40);
buf BUF1 (N2244, N2221);
or OR2 (N2245, N2241, N689);
buf BUF1 (N2246, N2242);
buf BUF1 (N2247, N2246);
xor XOR2 (N2248, N2243, N1844);
nand NAND3 (N2249, N2240, N60, N1709);
not NOT1 (N2250, N2227);
nor NOR4 (N2251, N2247, N2084, N68, N240);
or OR2 (N2252, N2249, N1451);
and AND2 (N2253, N2231, N152);
xor XOR2 (N2254, N2244, N2030);
not NOT1 (N2255, N2232);
buf BUF1 (N2256, N2251);
or OR3 (N2257, N2236, N597, N519);
buf BUF1 (N2258, N2250);
and AND4 (N2259, N2254, N301, N849, N2033);
and AND3 (N2260, N2245, N1836, N2175);
nand NAND3 (N2261, N2258, N1474, N1469);
nand NAND3 (N2262, N2257, N1898, N1557);
buf BUF1 (N2263, N2262);
nor NOR3 (N2264, N2253, N69, N202);
nor NOR3 (N2265, N2263, N831, N930);
nor NOR3 (N2266, N2264, N1165, N740);
xor XOR2 (N2267, N2265, N1112);
buf BUF1 (N2268, N2255);
buf BUF1 (N2269, N2217);
xor XOR2 (N2270, N2267, N1488);
not NOT1 (N2271, N2256);
xor XOR2 (N2272, N2260, N950);
buf BUF1 (N2273, N2261);
nand NAND2 (N2274, N2266, N2084);
not NOT1 (N2275, N2274);
or OR3 (N2276, N2272, N1050, N584);
buf BUF1 (N2277, N2275);
not NOT1 (N2278, N2268);
not NOT1 (N2279, N2259);
or OR4 (N2280, N2269, N674, N615, N1678);
or OR3 (N2281, N2277, N1915, N1526);
buf BUF1 (N2282, N2276);
nor NOR4 (N2283, N2278, N1577, N274, N1628);
not NOT1 (N2284, N2248);
nand NAND4 (N2285, N2283, N1885, N499, N905);
nor NOR4 (N2286, N2284, N1446, N846, N201);
nor NOR4 (N2287, N2282, N1852, N720, N2067);
and AND3 (N2288, N2273, N723, N1010);
nand NAND3 (N2289, N2280, N351, N1805);
nand NAND4 (N2290, N2286, N19, N774, N83);
xor XOR2 (N2291, N2290, N2173);
and AND3 (N2292, N2279, N223, N2056);
or OR3 (N2293, N2281, N1694, N1432);
buf BUF1 (N2294, N2289);
nand NAND3 (N2295, N2287, N2040, N1428);
and AND4 (N2296, N2295, N660, N2003, N1867);
not NOT1 (N2297, N2271);
nor NOR4 (N2298, N2252, N543, N1555, N1560);
and AND4 (N2299, N2293, N123, N453, N319);
buf BUF1 (N2300, N2285);
and AND2 (N2301, N2300, N2154);
not NOT1 (N2302, N2296);
buf BUF1 (N2303, N2292);
nor NOR4 (N2304, N2288, N2296, N548, N1211);
or OR2 (N2305, N2299, N1750);
nand NAND2 (N2306, N2303, N1847);
or OR4 (N2307, N2270, N1376, N737, N137);
or OR4 (N2308, N2302, N78, N72, N1361);
buf BUF1 (N2309, N2305);
nand NAND2 (N2310, N2304, N1621);
nor NOR3 (N2311, N2301, N596, N1185);
nand NAND3 (N2312, N2291, N1241, N2161);
nor NOR2 (N2313, N2307, N96);
buf BUF1 (N2314, N2310);
xor XOR2 (N2315, N2313, N1013);
and AND3 (N2316, N2312, N131, N321);
nand NAND3 (N2317, N2294, N302, N521);
xor XOR2 (N2318, N2308, N160);
nor NOR3 (N2319, N2314, N1198, N359);
nor NOR4 (N2320, N2306, N1519, N1600, N795);
xor XOR2 (N2321, N2318, N284);
not NOT1 (N2322, N2311);
or OR2 (N2323, N2315, N642);
buf BUF1 (N2324, N2316);
nand NAND2 (N2325, N2309, N1252);
and AND4 (N2326, N2322, N1871, N801, N483);
not NOT1 (N2327, N2317);
or OR3 (N2328, N2321, N1216, N1625);
and AND2 (N2329, N2324, N1523);
buf BUF1 (N2330, N2320);
xor XOR2 (N2331, N2323, N38);
buf BUF1 (N2332, N2319);
and AND2 (N2333, N2330, N1837);
nor NOR3 (N2334, N2297, N2286, N2244);
not NOT1 (N2335, N2298);
nor NOR4 (N2336, N2331, N1550, N1833, N71);
xor XOR2 (N2337, N2327, N990);
buf BUF1 (N2338, N2335);
buf BUF1 (N2339, N2325);
buf BUF1 (N2340, N2328);
or OR3 (N2341, N2326, N1025, N2004);
nor NOR3 (N2342, N2341, N1570, N2142);
xor XOR2 (N2343, N2339, N685);
and AND4 (N2344, N2338, N156, N923, N1606);
or OR4 (N2345, N2342, N1310, N1609, N1689);
nand NAND3 (N2346, N2343, N1281, N1079);
buf BUF1 (N2347, N2336);
nand NAND3 (N2348, N2334, N1174, N1745);
nand NAND2 (N2349, N2346, N2297);
not NOT1 (N2350, N2344);
or OR3 (N2351, N2340, N2183, N283);
buf BUF1 (N2352, N2329);
nand NAND3 (N2353, N2348, N609, N1129);
and AND3 (N2354, N2345, N618, N1646);
or OR2 (N2355, N2349, N9);
nor NOR4 (N2356, N2333, N4, N898, N791);
and AND4 (N2357, N2356, N1557, N478, N52);
and AND3 (N2358, N2351, N454, N931);
buf BUF1 (N2359, N2350);
or OR3 (N2360, N2337, N1068, N310);
and AND2 (N2361, N2352, N312);
or OR3 (N2362, N2359, N603, N869);
or OR2 (N2363, N2361, N691);
nand NAND2 (N2364, N2332, N2016);
nand NAND3 (N2365, N2354, N1522, N198);
not NOT1 (N2366, N2355);
nor NOR3 (N2367, N2365, N1403, N1811);
or OR3 (N2368, N2364, N1612, N1371);
nor NOR2 (N2369, N2347, N515);
xor XOR2 (N2370, N2366, N385);
nor NOR3 (N2371, N2358, N1070, N2033);
or OR4 (N2372, N2369, N448, N760, N1744);
xor XOR2 (N2373, N2353, N957);
and AND2 (N2374, N2372, N2168);
or OR2 (N2375, N2374, N1802);
or OR3 (N2376, N2375, N1352, N712);
not NOT1 (N2377, N2373);
xor XOR2 (N2378, N2376, N1450);
or OR3 (N2379, N2367, N1130, N1884);
buf BUF1 (N2380, N2371);
and AND2 (N2381, N2379, N1910);
buf BUF1 (N2382, N2363);
and AND2 (N2383, N2377, N368);
xor XOR2 (N2384, N2381, N1125);
nor NOR3 (N2385, N2382, N2188, N2275);
nand NAND4 (N2386, N2380, N1987, N1309, N471);
not NOT1 (N2387, N2383);
not NOT1 (N2388, N2385);
not NOT1 (N2389, N2388);
nor NOR4 (N2390, N2387, N356, N263, N1731);
buf BUF1 (N2391, N2368);
nand NAND3 (N2392, N2386, N2168, N783);
and AND3 (N2393, N2389, N637, N1580);
not NOT1 (N2394, N2362);
nand NAND2 (N2395, N2394, N285);
xor XOR2 (N2396, N2392, N1838);
nand NAND4 (N2397, N2384, N1743, N1015, N1476);
and AND3 (N2398, N2357, N2100, N2112);
and AND3 (N2399, N2397, N1956, N1945);
buf BUF1 (N2400, N2393);
buf BUF1 (N2401, N2390);
or OR3 (N2402, N2400, N287, N900);
and AND2 (N2403, N2395, N1450);
nor NOR2 (N2404, N2378, N1601);
xor XOR2 (N2405, N2402, N607);
nor NOR2 (N2406, N2360, N370);
not NOT1 (N2407, N2399);
buf BUF1 (N2408, N2391);
xor XOR2 (N2409, N2398, N68);
xor XOR2 (N2410, N2406, N1477);
and AND3 (N2411, N2396, N1343, N2084);
nand NAND2 (N2412, N2410, N741);
xor XOR2 (N2413, N2411, N1666);
or OR4 (N2414, N2401, N281, N2310, N2114);
and AND2 (N2415, N2403, N1582);
not NOT1 (N2416, N2415);
xor XOR2 (N2417, N2412, N119);
and AND3 (N2418, N2409, N1947, N2098);
nand NAND3 (N2419, N2417, N1596, N1100);
nor NOR4 (N2420, N2407, N1685, N847, N446);
nand NAND2 (N2421, N2419, N780);
not NOT1 (N2422, N2370);
buf BUF1 (N2423, N2413);
buf BUF1 (N2424, N2416);
or OR4 (N2425, N2424, N1604, N96, N1501);
buf BUF1 (N2426, N2405);
xor XOR2 (N2427, N2422, N447);
nand NAND4 (N2428, N2423, N73, N1739, N213);
or OR4 (N2429, N2404, N386, N52, N528);
buf BUF1 (N2430, N2418);
nand NAND3 (N2431, N2428, N1616, N1803);
nand NAND2 (N2432, N2431, N347);
or OR2 (N2433, N2421, N2189);
nand NAND3 (N2434, N2433, N1527, N1926);
and AND4 (N2435, N2434, N1573, N1698, N586);
not NOT1 (N2436, N2426);
buf BUF1 (N2437, N2420);
buf BUF1 (N2438, N2408);
xor XOR2 (N2439, N2427, N2386);
buf BUF1 (N2440, N2436);
or OR2 (N2441, N2438, N1069);
or OR2 (N2442, N2425, N2390);
not NOT1 (N2443, N2441);
and AND2 (N2444, N2443, N678);
xor XOR2 (N2445, N2429, N1677);
xor XOR2 (N2446, N2430, N1164);
nand NAND3 (N2447, N2432, N236, N435);
not NOT1 (N2448, N2437);
nand NAND3 (N2449, N2445, N225, N2408);
xor XOR2 (N2450, N2439, N468);
buf BUF1 (N2451, N2447);
or OR3 (N2452, N2440, N1533, N440);
and AND2 (N2453, N2452, N13);
or OR4 (N2454, N2446, N942, N308, N1808);
and AND3 (N2455, N2453, N1558, N938);
xor XOR2 (N2456, N2455, N11);
nor NOR3 (N2457, N2454, N713, N847);
buf BUF1 (N2458, N2450);
and AND3 (N2459, N2414, N365, N1252);
or OR4 (N2460, N2448, N1031, N2082, N827);
nand NAND3 (N2461, N2451, N1648, N1425);
nor NOR4 (N2462, N2458, N1457, N663, N1092);
or OR4 (N2463, N2460, N1967, N1373, N2317);
nand NAND3 (N2464, N2444, N1514, N1520);
xor XOR2 (N2465, N2449, N2078);
not NOT1 (N2466, N2459);
or OR4 (N2467, N2435, N1298, N2458, N2280);
nor NOR2 (N2468, N2461, N196);
not NOT1 (N2469, N2456);
and AND3 (N2470, N2463, N1440, N843);
not NOT1 (N2471, N2442);
and AND2 (N2472, N2467, N549);
nor NOR3 (N2473, N2466, N2227, N1432);
xor XOR2 (N2474, N2469, N2372);
or OR2 (N2475, N2470, N1137);
and AND3 (N2476, N2474, N559, N91);
nand NAND2 (N2477, N2471, N1897);
and AND3 (N2478, N2477, N1173, N849);
and AND4 (N2479, N2462, N565, N1031, N461);
nor NOR2 (N2480, N2479, N892);
nor NOR3 (N2481, N2476, N1457, N1493);
and AND3 (N2482, N2464, N278, N2182);
and AND4 (N2483, N2481, N859, N2431, N2434);
nand NAND3 (N2484, N2472, N355, N1558);
not NOT1 (N2485, N2475);
or OR3 (N2486, N2457, N983, N2129);
nand NAND2 (N2487, N2468, N1552);
or OR4 (N2488, N2482, N1777, N1291, N2003);
nand NAND4 (N2489, N2480, N2279, N32, N665);
xor XOR2 (N2490, N2488, N1460);
or OR4 (N2491, N2484, N727, N397, N1226);
not NOT1 (N2492, N2489);
nand NAND4 (N2493, N2465, N826, N830, N2214);
not NOT1 (N2494, N2483);
xor XOR2 (N2495, N2487, N2186);
xor XOR2 (N2496, N2494, N2443);
xor XOR2 (N2497, N2493, N1508);
nand NAND3 (N2498, N2478, N1132, N2393);
not NOT1 (N2499, N2497);
or OR3 (N2500, N2491, N746, N2235);
nand NAND4 (N2501, N2492, N1686, N2106, N1747);
or OR2 (N2502, N2498, N1041);
xor XOR2 (N2503, N2486, N1063);
or OR3 (N2504, N2485, N2102, N343);
xor XOR2 (N2505, N2503, N1037);
nor NOR3 (N2506, N2496, N1796, N501);
xor XOR2 (N2507, N2505, N1540);
buf BUF1 (N2508, N2501);
xor XOR2 (N2509, N2508, N705);
and AND3 (N2510, N2504, N252, N842);
nor NOR4 (N2511, N2500, N146, N1579, N1205);
and AND2 (N2512, N2507, N1281);
not NOT1 (N2513, N2509);
nand NAND2 (N2514, N2511, N1652);
or OR4 (N2515, N2510, N1771, N2115, N202);
not NOT1 (N2516, N2512);
nand NAND2 (N2517, N2514, N2434);
nor NOR4 (N2518, N2513, N104, N798, N480);
nand NAND2 (N2519, N2516, N32);
or OR4 (N2520, N2502, N1989, N863, N601);
nand NAND3 (N2521, N2517, N512, N2049);
not NOT1 (N2522, N2521);
nand NAND3 (N2523, N2499, N1936, N21);
nand NAND3 (N2524, N2490, N2322, N1924);
buf BUF1 (N2525, N2520);
and AND3 (N2526, N2515, N2252, N1950);
xor XOR2 (N2527, N2506, N1784);
nand NAND2 (N2528, N2519, N562);
nor NOR2 (N2529, N2473, N2266);
or OR2 (N2530, N2527, N2179);
buf BUF1 (N2531, N2495);
not NOT1 (N2532, N2525);
nor NOR4 (N2533, N2518, N737, N1126, N83);
or OR2 (N2534, N2529, N1670);
not NOT1 (N2535, N2526);
buf BUF1 (N2536, N2524);
nand NAND2 (N2537, N2528, N54);
or OR3 (N2538, N2535, N2166, N458);
nand NAND3 (N2539, N2532, N632, N2533);
not NOT1 (N2540, N2317);
xor XOR2 (N2541, N2523, N493);
buf BUF1 (N2542, N2536);
and AND3 (N2543, N2540, N1252, N116);
nand NAND2 (N2544, N2534, N536);
nand NAND4 (N2545, N2541, N1787, N568, N2400);
nor NOR3 (N2546, N2537, N1063, N565);
not NOT1 (N2547, N2531);
or OR4 (N2548, N2546, N29, N1085, N1343);
or OR3 (N2549, N2542, N918, N1435);
nor NOR4 (N2550, N2548, N70, N1846, N1199);
or OR2 (N2551, N2538, N2296);
nor NOR3 (N2552, N2545, N735, N1793);
buf BUF1 (N2553, N2522);
xor XOR2 (N2554, N2550, N1412);
nor NOR3 (N2555, N2549, N1297, N663);
nand NAND4 (N2556, N2530, N1844, N1142, N2282);
or OR2 (N2557, N2555, N2007);
nor NOR2 (N2558, N2557, N2530);
nand NAND4 (N2559, N2551, N1900, N346, N975);
and AND2 (N2560, N2554, N2216);
nor NOR4 (N2561, N2552, N328, N849, N267);
or OR4 (N2562, N2561, N1837, N1993, N61);
nor NOR4 (N2563, N2547, N2416, N607, N2241);
not NOT1 (N2564, N2559);
not NOT1 (N2565, N2563);
not NOT1 (N2566, N2564);
xor XOR2 (N2567, N2566, N1231);
buf BUF1 (N2568, N2553);
or OR2 (N2569, N2543, N2214);
and AND4 (N2570, N2569, N884, N296, N1250);
not NOT1 (N2571, N2562);
nand NAND4 (N2572, N2544, N2125, N1745, N2425);
not NOT1 (N2573, N2568);
buf BUF1 (N2574, N2571);
or OR2 (N2575, N2558, N51);
xor XOR2 (N2576, N2573, N1335);
not NOT1 (N2577, N2570);
xor XOR2 (N2578, N2565, N1930);
nor NOR2 (N2579, N2572, N715);
xor XOR2 (N2580, N2576, N1887);
xor XOR2 (N2581, N2560, N2027);
nand NAND4 (N2582, N2575, N2337, N1819, N1430);
not NOT1 (N2583, N2577);
not NOT1 (N2584, N2556);
not NOT1 (N2585, N2578);
nor NOR2 (N2586, N2580, N66);
nand NAND4 (N2587, N2579, N1646, N1117, N90);
xor XOR2 (N2588, N2583, N2159);
xor XOR2 (N2589, N2539, N821);
or OR3 (N2590, N2582, N1998, N1576);
xor XOR2 (N2591, N2584, N2052);
not NOT1 (N2592, N2574);
and AND4 (N2593, N2581, N279, N2407, N991);
nor NOR2 (N2594, N2586, N1817);
and AND4 (N2595, N2591, N832, N1865, N2184);
buf BUF1 (N2596, N2567);
xor XOR2 (N2597, N2585, N1535);
not NOT1 (N2598, N2588);
not NOT1 (N2599, N2598);
buf BUF1 (N2600, N2589);
not NOT1 (N2601, N2592);
nor NOR4 (N2602, N2599, N218, N2203, N1377);
xor XOR2 (N2603, N2596, N2037);
buf BUF1 (N2604, N2601);
and AND2 (N2605, N2603, N1820);
nor NOR4 (N2606, N2597, N428, N920, N1092);
and AND2 (N2607, N2604, N2136);
not NOT1 (N2608, N2605);
nand NAND4 (N2609, N2600, N1740, N2595, N725);
nor NOR4 (N2610, N68, N594, N837, N934);
nand NAND2 (N2611, N2606, N379);
buf BUF1 (N2612, N2593);
nor NOR4 (N2613, N2607, N65, N2550, N619);
not NOT1 (N2614, N2608);
nor NOR4 (N2615, N2594, N1451, N502, N1273);
buf BUF1 (N2616, N2614);
and AND2 (N2617, N2587, N1719);
xor XOR2 (N2618, N2602, N1212);
buf BUF1 (N2619, N2610);
buf BUF1 (N2620, N2590);
nor NOR3 (N2621, N2613, N1167, N1667);
nand NAND3 (N2622, N2616, N1461, N312);
buf BUF1 (N2623, N2617);
and AND3 (N2624, N2619, N2141, N2504);
not NOT1 (N2625, N2623);
nand NAND2 (N2626, N2622, N2187);
and AND4 (N2627, N2624, N1909, N47, N766);
not NOT1 (N2628, N2618);
nor NOR4 (N2629, N2620, N316, N1760, N1983);
not NOT1 (N2630, N2609);
buf BUF1 (N2631, N2629);
nand NAND4 (N2632, N2615, N11, N2493, N360);
nor NOR3 (N2633, N2627, N1647, N259);
nand NAND3 (N2634, N2612, N118, N888);
xor XOR2 (N2635, N2628, N897);
or OR2 (N2636, N2626, N1374);
nor NOR4 (N2637, N2635, N312, N2493, N1529);
not NOT1 (N2638, N2631);
nor NOR2 (N2639, N2634, N1459);
nand NAND3 (N2640, N2638, N521, N1239);
xor XOR2 (N2641, N2636, N79);
not NOT1 (N2642, N2630);
and AND4 (N2643, N2639, N1716, N204, N593);
xor XOR2 (N2644, N2637, N544);
xor XOR2 (N2645, N2644, N2288);
buf BUF1 (N2646, N2640);
nor NOR4 (N2647, N2643, N2564, N62, N370);
buf BUF1 (N2648, N2642);
and AND2 (N2649, N2648, N2019);
not NOT1 (N2650, N2649);
or OR4 (N2651, N2625, N66, N523, N2415);
and AND4 (N2652, N2633, N519, N364, N393);
or OR3 (N2653, N2652, N14, N126);
buf BUF1 (N2654, N2650);
or OR2 (N2655, N2647, N1899);
xor XOR2 (N2656, N2655, N2302);
or OR3 (N2657, N2646, N1704, N997);
not NOT1 (N2658, N2621);
or OR4 (N2659, N2641, N213, N380, N1503);
buf BUF1 (N2660, N2656);
nor NOR2 (N2661, N2611, N2366);
nand NAND4 (N2662, N2651, N1241, N1394, N6);
or OR4 (N2663, N2654, N170, N2581, N379);
buf BUF1 (N2664, N2657);
and AND4 (N2665, N2661, N2513, N1760, N1282);
nand NAND3 (N2666, N2658, N1555, N2251);
nor NOR2 (N2667, N2662, N495);
buf BUF1 (N2668, N2666);
xor XOR2 (N2669, N2663, N1888);
nand NAND4 (N2670, N2659, N1101, N2520, N631);
and AND2 (N2671, N2668, N1318);
xor XOR2 (N2672, N2669, N1837);
not NOT1 (N2673, N2665);
nand NAND3 (N2674, N2672, N532, N606);
nand NAND4 (N2675, N2670, N1420, N809, N2225);
nor NOR4 (N2676, N2671, N220, N409, N2439);
and AND3 (N2677, N2675, N1645, N2447);
xor XOR2 (N2678, N2664, N1417);
or OR3 (N2679, N2660, N237, N2570);
not NOT1 (N2680, N2653);
nor NOR3 (N2681, N2674, N303, N1447);
nor NOR4 (N2682, N2676, N2464, N1473, N2024);
not NOT1 (N2683, N2677);
xor XOR2 (N2684, N2682, N866);
not NOT1 (N2685, N2632);
or OR2 (N2686, N2681, N558);
or OR3 (N2687, N2680, N2076, N1970);
nor NOR3 (N2688, N2678, N387, N1164);
and AND2 (N2689, N2684, N36);
and AND2 (N2690, N2687, N2430);
nand NAND2 (N2691, N2679, N2228);
and AND2 (N2692, N2686, N2287);
and AND3 (N2693, N2688, N1085, N2555);
not NOT1 (N2694, N2691);
and AND3 (N2695, N2690, N1071, N2052);
nor NOR2 (N2696, N2693, N1543);
nand NAND3 (N2697, N2692, N1776, N2168);
or OR2 (N2698, N2645, N1654);
nand NAND3 (N2699, N2689, N2053, N1290);
not NOT1 (N2700, N2695);
nor NOR3 (N2701, N2667, N1865, N607);
and AND3 (N2702, N2700, N1151, N457);
xor XOR2 (N2703, N2673, N2219);
nand NAND2 (N2704, N2696, N2498);
nor NOR4 (N2705, N2704, N2533, N6, N298);
xor XOR2 (N2706, N2699, N2561);
buf BUF1 (N2707, N2694);
nand NAND3 (N2708, N2703, N1542, N1596);
and AND2 (N2709, N2685, N2246);
buf BUF1 (N2710, N2702);
nor NOR2 (N2711, N2707, N2624);
not NOT1 (N2712, N2705);
nand NAND3 (N2713, N2711, N1829, N978);
buf BUF1 (N2714, N2683);
nand NAND2 (N2715, N2708, N1163);
or OR2 (N2716, N2701, N1883);
nor NOR3 (N2717, N2713, N305, N1362);
not NOT1 (N2718, N2716);
nor NOR3 (N2719, N2714, N2545, N1497);
and AND2 (N2720, N2698, N164);
and AND3 (N2721, N2706, N1340, N235);
xor XOR2 (N2722, N2718, N528);
or OR3 (N2723, N2719, N765, N996);
and AND4 (N2724, N2723, N2289, N1989, N2464);
not NOT1 (N2725, N2721);
buf BUF1 (N2726, N2725);
buf BUF1 (N2727, N2720);
nor NOR3 (N2728, N2724, N683, N293);
and AND4 (N2729, N2710, N1655, N2636, N1166);
buf BUF1 (N2730, N2697);
or OR4 (N2731, N2728, N607, N2018, N682);
not NOT1 (N2732, N2722);
nor NOR3 (N2733, N2709, N1432, N670);
nor NOR2 (N2734, N2726, N740);
and AND2 (N2735, N2730, N2278);
and AND2 (N2736, N2729, N958);
xor XOR2 (N2737, N2734, N267);
xor XOR2 (N2738, N2733, N455);
xor XOR2 (N2739, N2738, N2125);
nor NOR4 (N2740, N2732, N469, N243, N1058);
xor XOR2 (N2741, N2712, N1532);
not NOT1 (N2742, N2727);
buf BUF1 (N2743, N2731);
nor NOR2 (N2744, N2715, N1641);
nor NOR3 (N2745, N2737, N1251, N569);
xor XOR2 (N2746, N2717, N1876);
or OR3 (N2747, N2743, N1027, N1713);
or OR3 (N2748, N2736, N2454, N598);
or OR3 (N2749, N2748, N2694, N2591);
and AND2 (N2750, N2739, N2233);
nor NOR3 (N2751, N2744, N191, N1705);
not NOT1 (N2752, N2746);
nand NAND2 (N2753, N2745, N919);
nor NOR4 (N2754, N2747, N360, N289, N113);
nand NAND3 (N2755, N2751, N1722, N552);
nand NAND3 (N2756, N2740, N1350, N1318);
not NOT1 (N2757, N2753);
nor NOR3 (N2758, N2735, N1646, N2524);
nand NAND4 (N2759, N2757, N273, N202, N2586);
buf BUF1 (N2760, N2759);
nand NAND4 (N2761, N2758, N2539, N1012, N2268);
xor XOR2 (N2762, N2749, N1625);
nor NOR4 (N2763, N2760, N751, N1741, N2326);
buf BUF1 (N2764, N2761);
buf BUF1 (N2765, N2750);
nand NAND3 (N2766, N2762, N831, N1184);
or OR4 (N2767, N2756, N1577, N328, N1650);
or OR3 (N2768, N2742, N1067, N734);
or OR4 (N2769, N2754, N476, N1481, N2448);
nand NAND3 (N2770, N2769, N2352, N1747);
or OR3 (N2771, N2755, N1071, N415);
not NOT1 (N2772, N2771);
and AND2 (N2773, N2772, N631);
nor NOR3 (N2774, N2763, N504, N78);
and AND3 (N2775, N2774, N1507, N861);
not NOT1 (N2776, N2768);
not NOT1 (N2777, N2775);
buf BUF1 (N2778, N2767);
not NOT1 (N2779, N2777);
nand NAND3 (N2780, N2741, N472, N885);
nor NOR4 (N2781, N2752, N1235, N2129, N1395);
xor XOR2 (N2782, N2779, N533);
buf BUF1 (N2783, N2770);
nand NAND2 (N2784, N2773, N374);
or OR4 (N2785, N2778, N1208, N732, N2064);
and AND3 (N2786, N2766, N2178, N511);
and AND3 (N2787, N2785, N726, N411);
nand NAND2 (N2788, N2765, N917);
not NOT1 (N2789, N2776);
nand NAND3 (N2790, N2789, N772, N2318);
xor XOR2 (N2791, N2764, N368);
or OR3 (N2792, N2782, N2138, N1614);
not NOT1 (N2793, N2780);
nor NOR2 (N2794, N2792, N502);
and AND3 (N2795, N2787, N1331, N922);
nand NAND3 (N2796, N2786, N1493, N1736);
nor NOR3 (N2797, N2784, N1447, N2713);
or OR3 (N2798, N2796, N1981, N2445);
and AND3 (N2799, N2798, N255, N1822);
not NOT1 (N2800, N2793);
nand NAND2 (N2801, N2795, N754);
xor XOR2 (N2802, N2783, N167);
buf BUF1 (N2803, N2800);
xor XOR2 (N2804, N2801, N1013);
nand NAND2 (N2805, N2791, N2390);
nand NAND3 (N2806, N2803, N158, N2051);
xor XOR2 (N2807, N2781, N1344);
nand NAND4 (N2808, N2794, N2405, N1903, N1965);
and AND3 (N2809, N2790, N2591, N1852);
not NOT1 (N2810, N2797);
nor NOR4 (N2811, N2807, N1571, N1766, N2466);
nor NOR3 (N2812, N2788, N51, N254);
nor NOR2 (N2813, N2811, N840);
xor XOR2 (N2814, N2799, N1786);
nand NAND2 (N2815, N2802, N64);
or OR4 (N2816, N2813, N1680, N59, N889);
nand NAND2 (N2817, N2815, N2422);
not NOT1 (N2818, N2808);
and AND3 (N2819, N2814, N633, N2545);
xor XOR2 (N2820, N2812, N240);
nand NAND4 (N2821, N2819, N2731, N1017, N1763);
and AND3 (N2822, N2821, N2226, N227);
or OR4 (N2823, N2817, N1362, N2807, N884);
xor XOR2 (N2824, N2806, N2084);
xor XOR2 (N2825, N2809, N1307);
buf BUF1 (N2826, N2820);
nand NAND3 (N2827, N2823, N1945, N1146);
nor NOR4 (N2828, N2824, N2307, N1569, N2381);
nor NOR3 (N2829, N2804, N1066, N2374);
nor NOR4 (N2830, N2827, N2440, N1820, N1323);
not NOT1 (N2831, N2826);
or OR2 (N2832, N2822, N92);
nand NAND4 (N2833, N2810, N2502, N2009, N1801);
or OR3 (N2834, N2825, N1675, N1882);
nand NAND3 (N2835, N2830, N563, N347);
nor NOR3 (N2836, N2816, N2041, N2513);
and AND4 (N2837, N2828, N149, N568, N1767);
buf BUF1 (N2838, N2837);
or OR3 (N2839, N2818, N516, N195);
and AND3 (N2840, N2836, N630, N2513);
or OR4 (N2841, N2805, N1348, N2751, N974);
nand NAND2 (N2842, N2833, N1742);
nand NAND4 (N2843, N2829, N2499, N1233, N2743);
nand NAND3 (N2844, N2839, N641, N52);
buf BUF1 (N2845, N2844);
xor XOR2 (N2846, N2842, N2665);
nand NAND2 (N2847, N2843, N949);
and AND3 (N2848, N2840, N1698, N489);
and AND3 (N2849, N2845, N2779, N608);
xor XOR2 (N2850, N2834, N803);
and AND2 (N2851, N2832, N721);
or OR4 (N2852, N2848, N414, N896, N863);
xor XOR2 (N2853, N2852, N1603);
xor XOR2 (N2854, N2846, N2407);
or OR2 (N2855, N2831, N1561);
or OR4 (N2856, N2854, N2722, N887, N1755);
nand NAND4 (N2857, N2850, N839, N1523, N2358);
buf BUF1 (N2858, N2855);
or OR3 (N2859, N2838, N425, N700);
buf BUF1 (N2860, N2849);
or OR2 (N2861, N2851, N278);
and AND3 (N2862, N2841, N7, N1069);
and AND3 (N2863, N2835, N296, N715);
nor NOR2 (N2864, N2860, N1338);
xor XOR2 (N2865, N2856, N2507);
and AND3 (N2866, N2857, N2602, N2803);
or OR4 (N2867, N2847, N827, N2617, N1521);
nor NOR3 (N2868, N2858, N1664, N128);
not NOT1 (N2869, N2853);
nor NOR4 (N2870, N2866, N2028, N2356, N1160);
not NOT1 (N2871, N2864);
and AND3 (N2872, N2859, N1865, N298);
nor NOR4 (N2873, N2868, N2734, N1836, N521);
nor NOR3 (N2874, N2865, N2025, N2520);
nand NAND4 (N2875, N2874, N1375, N1687, N2236);
buf BUF1 (N2876, N2870);
nor NOR3 (N2877, N2861, N116, N1280);
and AND3 (N2878, N2872, N1736, N1633);
buf BUF1 (N2879, N2876);
buf BUF1 (N2880, N2871);
nor NOR4 (N2881, N2880, N2776, N147, N285);
nand NAND4 (N2882, N2881, N1877, N253, N1530);
and AND2 (N2883, N2862, N1089);
xor XOR2 (N2884, N2883, N2721);
or OR2 (N2885, N2877, N1834);
xor XOR2 (N2886, N2878, N808);
nand NAND3 (N2887, N2886, N540, N780);
or OR2 (N2888, N2875, N1083);
nor NOR4 (N2889, N2869, N2393, N2066, N2211);
buf BUF1 (N2890, N2887);
not NOT1 (N2891, N2884);
or OR3 (N2892, N2867, N1753, N316);
xor XOR2 (N2893, N2882, N2148);
not NOT1 (N2894, N2892);
not NOT1 (N2895, N2890);
xor XOR2 (N2896, N2893, N266);
xor XOR2 (N2897, N2873, N1198);
nand NAND2 (N2898, N2894, N2360);
nor NOR2 (N2899, N2896, N410);
not NOT1 (N2900, N2863);
buf BUF1 (N2901, N2889);
xor XOR2 (N2902, N2885, N677);
and AND2 (N2903, N2897, N464);
not NOT1 (N2904, N2895);
xor XOR2 (N2905, N2901, N856);
not NOT1 (N2906, N2905);
or OR4 (N2907, N2906, N2115, N2306, N1293);
buf BUF1 (N2908, N2891);
nor NOR4 (N2909, N2902, N866, N2465, N554);
or OR2 (N2910, N2909, N2652);
and AND4 (N2911, N2900, N2396, N288, N1056);
nor NOR4 (N2912, N2907, N2124, N1095, N2735);
xor XOR2 (N2913, N2899, N2452);
and AND2 (N2914, N2912, N1638);
and AND4 (N2915, N2911, N52, N1781, N663);
buf BUF1 (N2916, N2913);
xor XOR2 (N2917, N2908, N1239);
nor NOR2 (N2918, N2914, N332);
not NOT1 (N2919, N2917);
nor NOR4 (N2920, N2898, N782, N466, N1480);
nand NAND2 (N2921, N2888, N2375);
nor NOR4 (N2922, N2916, N2334, N1158, N1831);
and AND4 (N2923, N2904, N1997, N837, N1186);
nand NAND3 (N2924, N2920, N1108, N1249);
xor XOR2 (N2925, N2903, N414);
nor NOR4 (N2926, N2879, N742, N809, N2628);
buf BUF1 (N2927, N2922);
not NOT1 (N2928, N2924);
buf BUF1 (N2929, N2915);
nand NAND2 (N2930, N2919, N153);
buf BUF1 (N2931, N2923);
nor NOR3 (N2932, N2929, N700, N2559);
and AND4 (N2933, N2931, N2586, N1321, N1308);
or OR3 (N2934, N2927, N990, N417);
nand NAND3 (N2935, N2933, N799, N101);
and AND2 (N2936, N2918, N2209);
nor NOR4 (N2937, N2910, N2690, N222, N1863);
nor NOR3 (N2938, N2928, N2341, N1790);
xor XOR2 (N2939, N2935, N1714);
and AND3 (N2940, N2936, N1470, N1114);
xor XOR2 (N2941, N2932, N1663);
buf BUF1 (N2942, N2926);
nor NOR3 (N2943, N2937, N472, N2680);
and AND4 (N2944, N2930, N2011, N1214, N1676);
buf BUF1 (N2945, N2942);
nor NOR3 (N2946, N2943, N1163, N1058);
and AND4 (N2947, N2938, N1854, N460, N1232);
nor NOR3 (N2948, N2940, N2700, N1759);
buf BUF1 (N2949, N2939);
buf BUF1 (N2950, N2944);
or OR3 (N2951, N2949, N2004, N1545);
or OR3 (N2952, N2950, N213, N1161);
buf BUF1 (N2953, N2934);
buf BUF1 (N2954, N2941);
not NOT1 (N2955, N2925);
or OR3 (N2956, N2952, N2541, N189);
and AND3 (N2957, N2948, N2781, N2472);
xor XOR2 (N2958, N2953, N1271);
xor XOR2 (N2959, N2921, N1124);
xor XOR2 (N2960, N2958, N77);
xor XOR2 (N2961, N2945, N2157);
xor XOR2 (N2962, N2947, N508);
not NOT1 (N2963, N2951);
xor XOR2 (N2964, N2955, N255);
buf BUF1 (N2965, N2959);
nor NOR2 (N2966, N2956, N203);
nand NAND3 (N2967, N2965, N1300, N2592);
or OR3 (N2968, N2964, N311, N640);
not NOT1 (N2969, N2967);
nor NOR3 (N2970, N2946, N1921, N836);
not NOT1 (N2971, N2963);
nand NAND3 (N2972, N2954, N1284, N960);
xor XOR2 (N2973, N2972, N2926);
buf BUF1 (N2974, N2969);
xor XOR2 (N2975, N2971, N1598);
buf BUF1 (N2976, N2962);
xor XOR2 (N2977, N2970, N2909);
nor NOR4 (N2978, N2974, N1144, N1951, N1758);
or OR2 (N2979, N2976, N68);
nor NOR2 (N2980, N2979, N2668);
nand NAND3 (N2981, N2957, N744, N1345);
and AND3 (N2982, N2966, N751, N617);
nand NAND4 (N2983, N2981, N932, N2848, N2077);
nand NAND4 (N2984, N2975, N2159, N75, N446);
nor NOR2 (N2985, N2978, N2964);
and AND3 (N2986, N2960, N555, N1665);
buf BUF1 (N2987, N2982);
or OR2 (N2988, N2973, N1287);
buf BUF1 (N2989, N2980);
not NOT1 (N2990, N2988);
buf BUF1 (N2991, N2987);
or OR2 (N2992, N2961, N2932);
xor XOR2 (N2993, N2989, N2337);
nor NOR2 (N2994, N2968, N1853);
nor NOR3 (N2995, N2984, N2960, N1830);
not NOT1 (N2996, N2991);
xor XOR2 (N2997, N2983, N1000);
and AND2 (N2998, N2997, N2244);
nor NOR3 (N2999, N2993, N2419, N522);
nand NAND3 (N3000, N2998, N331, N1213);
nand NAND2 (N3001, N2977, N1838);
not NOT1 (N3002, N2994);
or OR2 (N3003, N3001, N1863);
or OR3 (N3004, N2995, N818, N2900);
buf BUF1 (N3005, N2996);
or OR2 (N3006, N2992, N1980);
and AND4 (N3007, N3000, N256, N2504, N2027);
or OR2 (N3008, N3004, N1970);
buf BUF1 (N3009, N3008);
nand NAND2 (N3010, N3002, N1807);
xor XOR2 (N3011, N2985, N2437);
and AND4 (N3012, N2999, N399, N1265, N2212);
buf BUF1 (N3013, N3005);
buf BUF1 (N3014, N2986);
not NOT1 (N3015, N3003);
xor XOR2 (N3016, N3012, N2893);
and AND2 (N3017, N3006, N611);
nand NAND3 (N3018, N3010, N1056, N1222);
not NOT1 (N3019, N3017);
xor XOR2 (N3020, N3013, N1552);
and AND3 (N3021, N3011, N2875, N2091);
not NOT1 (N3022, N3007);
not NOT1 (N3023, N3022);
buf BUF1 (N3024, N2990);
endmodule