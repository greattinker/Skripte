// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16;

output N1993,N2015,N1998,N2013,N1985,N2006,N2012,N2014,N2011,N2016;

not NOT1 (N17, N7);
buf BUF1 (N18, N7);
nand NAND2 (N19, N15, N9);
and AND3 (N20, N6, N7, N1);
xor XOR2 (N21, N5, N7);
not NOT1 (N22, N15);
nor NOR3 (N23, N11, N21, N14);
or OR4 (N24, N23, N1, N20, N23);
nor NOR4 (N25, N20, N7, N18, N4);
xor XOR2 (N26, N13, N23);
and AND3 (N27, N4, N24, N14);
nor NOR2 (N28, N4, N17);
buf BUF1 (N29, N26);
buf BUF1 (N30, N2);
not NOT1 (N31, N11);
xor XOR2 (N32, N12, N20);
or OR2 (N33, N2, N10);
not NOT1 (N34, N29);
buf BUF1 (N35, N34);
or OR4 (N36, N35, N20, N2, N13);
xor XOR2 (N37, N19, N19);
nor NOR4 (N38, N25, N9, N15, N34);
not NOT1 (N39, N37);
buf BUF1 (N40, N28);
xor XOR2 (N41, N32, N19);
buf BUF1 (N42, N40);
nand NAND3 (N43, N38, N23, N1);
xor XOR2 (N44, N31, N2);
xor XOR2 (N45, N39, N12);
or OR2 (N46, N44, N33);
nand NAND3 (N47, N4, N16, N46);
xor XOR2 (N48, N4, N26);
nor NOR4 (N49, N36, N1, N19, N31);
xor XOR2 (N50, N27, N20);
xor XOR2 (N51, N47, N5);
not NOT1 (N52, N45);
not NOT1 (N53, N50);
not NOT1 (N54, N53);
xor XOR2 (N55, N51, N20);
or OR3 (N56, N42, N17, N44);
nor NOR3 (N57, N52, N42, N21);
nor NOR2 (N58, N22, N13);
buf BUF1 (N59, N49);
buf BUF1 (N60, N54);
and AND4 (N61, N30, N38, N38, N19);
nand NAND3 (N62, N61, N45, N24);
nand NAND3 (N63, N57, N8, N16);
not NOT1 (N64, N48);
buf BUF1 (N65, N60);
nor NOR3 (N66, N65, N30, N5);
not NOT1 (N67, N64);
nor NOR2 (N68, N59, N37);
or OR3 (N69, N43, N67, N15);
nand NAND2 (N70, N38, N63);
not NOT1 (N71, N15);
or OR3 (N72, N55, N1, N59);
xor XOR2 (N73, N62, N32);
and AND3 (N74, N58, N38, N2);
and AND4 (N75, N72, N40, N12, N61);
or OR3 (N76, N75, N54, N29);
nor NOR4 (N77, N68, N62, N48, N53);
not NOT1 (N78, N76);
xor XOR2 (N79, N41, N1);
nor NOR2 (N80, N79, N55);
and AND2 (N81, N74, N73);
not NOT1 (N82, N41);
xor XOR2 (N83, N81, N18);
nor NOR3 (N84, N78, N20, N18);
or OR2 (N85, N84, N38);
xor XOR2 (N86, N70, N6);
or OR4 (N87, N69, N71, N24, N50);
and AND4 (N88, N61, N25, N84, N50);
or OR3 (N89, N83, N11, N74);
and AND4 (N90, N86, N36, N29, N15);
or OR4 (N91, N88, N85, N43, N22);
xor XOR2 (N92, N3, N83);
and AND2 (N93, N77, N7);
xor XOR2 (N94, N90, N1);
nor NOR2 (N95, N56, N83);
or OR4 (N96, N80, N87, N16, N31);
nand NAND2 (N97, N22, N1);
or OR3 (N98, N95, N23, N86);
buf BUF1 (N99, N89);
or OR2 (N100, N66, N14);
nand NAND3 (N101, N100, N72, N88);
xor XOR2 (N102, N93, N18);
not NOT1 (N103, N97);
nor NOR2 (N104, N96, N43);
and AND3 (N105, N101, N103, N60);
nor NOR3 (N106, N46, N10, N41);
not NOT1 (N107, N99);
buf BUF1 (N108, N106);
buf BUF1 (N109, N107);
and AND4 (N110, N102, N26, N48, N53);
not NOT1 (N111, N91);
not NOT1 (N112, N105);
not NOT1 (N113, N104);
xor XOR2 (N114, N98, N95);
nand NAND4 (N115, N94, N49, N13, N108);
nand NAND2 (N116, N114, N47);
and AND4 (N117, N33, N41, N56, N13);
xor XOR2 (N118, N115, N12);
xor XOR2 (N119, N109, N5);
and AND3 (N120, N113, N40, N22);
or OR4 (N121, N110, N56, N86, N38);
nor NOR3 (N122, N121, N25, N61);
nand NAND3 (N123, N117, N54, N25);
nor NOR3 (N124, N122, N40, N66);
xor XOR2 (N125, N118, N121);
nor NOR2 (N126, N123, N122);
and AND2 (N127, N111, N115);
xor XOR2 (N128, N82, N84);
nor NOR3 (N129, N127, N67, N60);
nand NAND3 (N130, N119, N20, N74);
buf BUF1 (N131, N92);
and AND3 (N132, N129, N46, N114);
or OR4 (N133, N120, N96, N103, N24);
nor NOR4 (N134, N133, N78, N67, N58);
and AND2 (N135, N128, N117);
or OR2 (N136, N134, N76);
nand NAND2 (N137, N126, N7);
or OR2 (N138, N112, N16);
and AND3 (N139, N136, N44, N58);
and AND4 (N140, N137, N70, N82, N14);
or OR3 (N141, N125, N36, N47);
nand NAND2 (N142, N138, N136);
or OR2 (N143, N135, N114);
not NOT1 (N144, N130);
buf BUF1 (N145, N139);
nor NOR2 (N146, N142, N2);
not NOT1 (N147, N116);
or OR2 (N148, N146, N92);
nor NOR2 (N149, N148, N58);
xor XOR2 (N150, N143, N49);
nor NOR2 (N151, N145, N65);
not NOT1 (N152, N131);
xor XOR2 (N153, N151, N19);
and AND2 (N154, N152, N62);
nand NAND4 (N155, N154, N39, N22, N55);
not NOT1 (N156, N132);
not NOT1 (N157, N141);
or OR4 (N158, N140, N98, N64, N95);
and AND3 (N159, N157, N139, N12);
or OR4 (N160, N156, N88, N5, N146);
nand NAND4 (N161, N124, N76, N79, N13);
buf BUF1 (N162, N158);
or OR4 (N163, N149, N118, N58, N42);
nand NAND3 (N164, N150, N25, N155);
and AND2 (N165, N70, N146);
nand NAND4 (N166, N144, N110, N1, N36);
and AND3 (N167, N164, N113, N1);
nor NOR3 (N168, N162, N39, N70);
buf BUF1 (N169, N147);
nor NOR2 (N170, N153, N154);
not NOT1 (N171, N163);
and AND4 (N172, N169, N151, N148, N64);
xor XOR2 (N173, N161, N49);
nor NOR4 (N174, N159, N65, N148, N12);
xor XOR2 (N175, N168, N80);
nor NOR2 (N176, N171, N167);
xor XOR2 (N177, N88, N139);
and AND4 (N178, N173, N103, N122, N89);
or OR2 (N179, N172, N81);
buf BUF1 (N180, N165);
buf BUF1 (N181, N166);
nor NOR3 (N182, N181, N32, N159);
buf BUF1 (N183, N180);
or OR4 (N184, N178, N126, N48, N116);
and AND2 (N185, N179, N169);
nand NAND4 (N186, N175, N183, N119, N172);
buf BUF1 (N187, N121);
buf BUF1 (N188, N182);
and AND4 (N189, N176, N95, N158, N92);
xor XOR2 (N190, N187, N86);
xor XOR2 (N191, N188, N94);
not NOT1 (N192, N170);
nor NOR2 (N193, N189, N11);
xor XOR2 (N194, N186, N63);
xor XOR2 (N195, N192, N44);
nand NAND4 (N196, N190, N54, N28, N171);
nor NOR2 (N197, N185, N124);
xor XOR2 (N198, N174, N103);
and AND4 (N199, N198, N87, N155, N27);
or OR2 (N200, N196, N25);
or OR2 (N201, N191, N149);
not NOT1 (N202, N199);
or OR3 (N203, N200, N111, N81);
xor XOR2 (N204, N193, N61);
buf BUF1 (N205, N203);
xor XOR2 (N206, N205, N24);
buf BUF1 (N207, N202);
xor XOR2 (N208, N177, N52);
nor NOR2 (N209, N208, N139);
not NOT1 (N210, N206);
nand NAND2 (N211, N207, N127);
nand NAND2 (N212, N201, N48);
or OR3 (N213, N209, N125, N6);
not NOT1 (N214, N160);
and AND3 (N215, N184, N64, N144);
buf BUF1 (N216, N212);
not NOT1 (N217, N204);
buf BUF1 (N218, N210);
and AND3 (N219, N211, N216, N130);
or OR4 (N220, N38, N99, N36, N156);
buf BUF1 (N221, N214);
nand NAND3 (N222, N217, N84, N169);
or OR3 (N223, N194, N181, N111);
nand NAND2 (N224, N197, N81);
buf BUF1 (N225, N224);
not NOT1 (N226, N220);
or OR4 (N227, N215, N190, N115, N152);
nand NAND3 (N228, N227, N15, N86);
buf BUF1 (N229, N225);
nand NAND4 (N230, N222, N140, N97, N60);
and AND4 (N231, N228, N168, N192, N111);
and AND4 (N232, N218, N173, N25, N129);
buf BUF1 (N233, N226);
not NOT1 (N234, N221);
not NOT1 (N235, N195);
nor NOR4 (N236, N235, N222, N129, N197);
or OR2 (N237, N230, N139);
and AND2 (N238, N231, N207);
nand NAND4 (N239, N213, N171, N192, N8);
nor NOR4 (N240, N229, N217, N222, N38);
buf BUF1 (N241, N232);
nor NOR2 (N242, N219, N49);
and AND3 (N243, N238, N79, N198);
nor NOR2 (N244, N233, N70);
or OR2 (N245, N241, N37);
or OR2 (N246, N239, N143);
buf BUF1 (N247, N244);
not NOT1 (N248, N246);
or OR3 (N249, N237, N69, N16);
not NOT1 (N250, N236);
nand NAND3 (N251, N250, N229, N117);
or OR4 (N252, N234, N149, N231, N204);
or OR4 (N253, N252, N68, N230, N162);
nor NOR2 (N254, N249, N232);
or OR4 (N255, N242, N248, N1, N236);
or OR3 (N256, N130, N75, N17);
nand NAND3 (N257, N223, N78, N183);
or OR2 (N258, N245, N74);
or OR2 (N259, N254, N143);
xor XOR2 (N260, N253, N61);
and AND3 (N261, N258, N124, N96);
nand NAND2 (N262, N257, N89);
nor NOR3 (N263, N260, N61, N179);
buf BUF1 (N264, N261);
nor NOR3 (N265, N262, N262, N182);
buf BUF1 (N266, N251);
buf BUF1 (N267, N259);
and AND2 (N268, N255, N182);
or OR4 (N269, N266, N248, N152, N202);
xor XOR2 (N270, N256, N260);
buf BUF1 (N271, N265);
xor XOR2 (N272, N264, N206);
not NOT1 (N273, N272);
xor XOR2 (N274, N273, N269);
not NOT1 (N275, N138);
nor NOR3 (N276, N267, N218, N189);
buf BUF1 (N277, N247);
xor XOR2 (N278, N270, N189);
or OR3 (N279, N243, N18, N208);
not NOT1 (N280, N274);
buf BUF1 (N281, N275);
not NOT1 (N282, N281);
and AND3 (N283, N280, N107, N12);
or OR2 (N284, N279, N233);
buf BUF1 (N285, N278);
buf BUF1 (N286, N268);
and AND3 (N287, N263, N172, N194);
nand NAND4 (N288, N285, N23, N56, N272);
nor NOR2 (N289, N283, N112);
nor NOR3 (N290, N277, N265, N252);
nor NOR2 (N291, N284, N121);
buf BUF1 (N292, N290);
or OR3 (N293, N287, N220, N53);
nand NAND2 (N294, N286, N147);
not NOT1 (N295, N276);
nor NOR3 (N296, N294, N220, N225);
buf BUF1 (N297, N291);
xor XOR2 (N298, N271, N158);
and AND4 (N299, N297, N150, N169, N157);
xor XOR2 (N300, N240, N116);
nor NOR2 (N301, N296, N77);
and AND2 (N302, N289, N19);
not NOT1 (N303, N300);
not NOT1 (N304, N301);
nand NAND3 (N305, N302, N74, N293);
nand NAND2 (N306, N160, N273);
nor NOR4 (N307, N306, N177, N248, N69);
buf BUF1 (N308, N305);
nand NAND2 (N309, N308, N249);
buf BUF1 (N310, N309);
buf BUF1 (N311, N310);
nand NAND3 (N312, N303, N207, N242);
not NOT1 (N313, N292);
nor NOR3 (N314, N295, N122, N18);
xor XOR2 (N315, N298, N58);
not NOT1 (N316, N307);
or OR2 (N317, N282, N160);
not NOT1 (N318, N313);
not NOT1 (N319, N312);
nor NOR2 (N320, N288, N86);
buf BUF1 (N321, N311);
xor XOR2 (N322, N321, N73);
or OR3 (N323, N320, N27, N271);
or OR3 (N324, N319, N196, N82);
nand NAND4 (N325, N315, N290, N109, N107);
nand NAND3 (N326, N317, N254, N238);
nand NAND2 (N327, N299, N29);
nand NAND3 (N328, N316, N33, N259);
nand NAND3 (N329, N325, N199, N261);
not NOT1 (N330, N323);
and AND2 (N331, N318, N321);
and AND2 (N332, N331, N207);
xor XOR2 (N333, N332, N222);
xor XOR2 (N334, N326, N208);
buf BUF1 (N335, N328);
buf BUF1 (N336, N335);
not NOT1 (N337, N324);
xor XOR2 (N338, N322, N129);
nand NAND4 (N339, N327, N83, N292, N219);
not NOT1 (N340, N339);
nor NOR4 (N341, N336, N146, N204, N18);
nor NOR2 (N342, N330, N289);
or OR3 (N343, N338, N6, N289);
nand NAND3 (N344, N341, N106, N333);
xor XOR2 (N345, N263, N193);
nor NOR3 (N346, N304, N233, N208);
or OR4 (N347, N314, N212, N100, N207);
not NOT1 (N348, N345);
buf BUF1 (N349, N340);
buf BUF1 (N350, N329);
buf BUF1 (N351, N337);
or OR2 (N352, N351, N243);
nor NOR2 (N353, N347, N28);
nand NAND3 (N354, N350, N130, N134);
and AND4 (N355, N354, N218, N317, N285);
nand NAND3 (N356, N343, N342, N242);
and AND3 (N357, N276, N127, N264);
and AND4 (N358, N349, N307, N325, N297);
nand NAND3 (N359, N357, N184, N138);
buf BUF1 (N360, N356);
buf BUF1 (N361, N355);
and AND4 (N362, N348, N187, N303, N156);
not NOT1 (N363, N334);
nor NOR2 (N364, N353, N142);
and AND4 (N365, N358, N120, N37, N129);
and AND3 (N366, N363, N106, N197);
xor XOR2 (N367, N366, N234);
buf BUF1 (N368, N362);
not NOT1 (N369, N346);
nand NAND3 (N370, N367, N133, N345);
and AND3 (N371, N360, N278, N15);
buf BUF1 (N372, N361);
xor XOR2 (N373, N371, N316);
or OR2 (N374, N370, N332);
and AND3 (N375, N365, N102, N31);
nand NAND2 (N376, N352, N338);
nand NAND4 (N377, N364, N127, N324, N351);
nor NOR2 (N378, N344, N5);
or OR2 (N379, N368, N159);
nand NAND2 (N380, N374, N95);
nor NOR4 (N381, N372, N277, N12, N120);
and AND4 (N382, N378, N41, N71, N30);
and AND2 (N383, N380, N14);
nor NOR2 (N384, N369, N249);
and AND3 (N385, N381, N119, N273);
not NOT1 (N386, N379);
nand NAND3 (N387, N375, N295, N50);
buf BUF1 (N388, N382);
or OR3 (N389, N377, N82, N225);
or OR3 (N390, N383, N221, N160);
not NOT1 (N391, N388);
buf BUF1 (N392, N384);
and AND2 (N393, N390, N75);
and AND4 (N394, N386, N217, N291, N339);
nor NOR3 (N395, N373, N393, N102);
buf BUF1 (N396, N376);
not NOT1 (N397, N89);
not NOT1 (N398, N394);
buf BUF1 (N399, N387);
buf BUF1 (N400, N396);
and AND4 (N401, N389, N252, N203, N323);
buf BUF1 (N402, N395);
xor XOR2 (N403, N398, N40);
xor XOR2 (N404, N397, N118);
or OR2 (N405, N403, N385);
not NOT1 (N406, N320);
and AND4 (N407, N392, N323, N136, N310);
xor XOR2 (N408, N359, N294);
not NOT1 (N409, N399);
buf BUF1 (N410, N407);
not NOT1 (N411, N408);
buf BUF1 (N412, N402);
buf BUF1 (N413, N391);
nor NOR3 (N414, N413, N310, N266);
xor XOR2 (N415, N414, N162);
nand NAND4 (N416, N401, N220, N121, N164);
or OR4 (N417, N411, N20, N82, N66);
xor XOR2 (N418, N416, N239);
nor NOR4 (N419, N409, N261, N286, N326);
or OR2 (N420, N406, N158);
and AND4 (N421, N405, N57, N51, N247);
and AND2 (N422, N418, N12);
nand NAND4 (N423, N410, N221, N218, N180);
or OR3 (N424, N420, N226, N82);
xor XOR2 (N425, N422, N291);
buf BUF1 (N426, N423);
nand NAND3 (N427, N426, N362, N155);
buf BUF1 (N428, N427);
or OR4 (N429, N421, N334, N189, N290);
xor XOR2 (N430, N428, N406);
and AND4 (N431, N419, N5, N35, N69);
buf BUF1 (N432, N417);
nand NAND4 (N433, N431, N28, N343, N417);
xor XOR2 (N434, N429, N256);
not NOT1 (N435, N424);
or OR3 (N436, N412, N104, N252);
nand NAND2 (N437, N434, N436);
xor XOR2 (N438, N204, N310);
nor NOR3 (N439, N433, N10, N12);
not NOT1 (N440, N430);
buf BUF1 (N441, N404);
and AND2 (N442, N432, N242);
nor NOR4 (N443, N440, N288, N35, N441);
and AND3 (N444, N131, N303, N65);
nand NAND2 (N445, N438, N336);
and AND2 (N446, N400, N402);
and AND2 (N447, N444, N40);
xor XOR2 (N448, N443, N432);
nand NAND4 (N449, N442, N242, N296, N402);
or OR2 (N450, N446, N126);
nor NOR2 (N451, N449, N39);
or OR3 (N452, N448, N146, N333);
xor XOR2 (N453, N425, N53);
xor XOR2 (N454, N415, N253);
nor NOR3 (N455, N447, N213, N241);
nand NAND4 (N456, N439, N71, N115, N235);
buf BUF1 (N457, N453);
and AND4 (N458, N452, N133, N366, N349);
nor NOR4 (N459, N445, N346, N395, N164);
buf BUF1 (N460, N437);
xor XOR2 (N461, N457, N457);
not NOT1 (N462, N459);
not NOT1 (N463, N460);
buf BUF1 (N464, N454);
or OR2 (N465, N458, N66);
nor NOR2 (N466, N461, N19);
xor XOR2 (N467, N466, N259);
nor NOR3 (N468, N455, N280, N234);
buf BUF1 (N469, N451);
nor NOR4 (N470, N462, N77, N455, N215);
xor XOR2 (N471, N467, N395);
or OR4 (N472, N456, N378, N185, N120);
not NOT1 (N473, N471);
buf BUF1 (N474, N472);
xor XOR2 (N475, N463, N91);
nor NOR3 (N476, N468, N175, N77);
nand NAND4 (N477, N435, N275, N228, N225);
xor XOR2 (N478, N474, N254);
buf BUF1 (N479, N450);
buf BUF1 (N480, N478);
nand NAND2 (N481, N477, N87);
buf BUF1 (N482, N464);
not NOT1 (N483, N480);
nor NOR3 (N484, N465, N388, N393);
and AND4 (N485, N476, N81, N169, N336);
buf BUF1 (N486, N479);
nand NAND4 (N487, N475, N107, N44, N262);
buf BUF1 (N488, N481);
nand NAND3 (N489, N485, N18, N365);
or OR2 (N490, N489, N462);
buf BUF1 (N491, N490);
nor NOR2 (N492, N488, N198);
or OR4 (N493, N470, N271, N192, N61);
nand NAND4 (N494, N482, N471, N239, N409);
buf BUF1 (N495, N492);
not NOT1 (N496, N494);
xor XOR2 (N497, N486, N475);
not NOT1 (N498, N483);
or OR2 (N499, N493, N86);
or OR4 (N500, N469, N241, N400, N93);
nand NAND4 (N501, N473, N485, N204, N183);
and AND2 (N502, N487, N479);
and AND4 (N503, N495, N348, N251, N190);
and AND4 (N504, N496, N194, N110, N65);
and AND4 (N505, N502, N233, N449, N147);
buf BUF1 (N506, N501);
nand NAND2 (N507, N497, N155);
and AND2 (N508, N498, N468);
not NOT1 (N509, N503);
nor NOR2 (N510, N499, N411);
nand NAND4 (N511, N508, N469, N94, N365);
or OR2 (N512, N491, N64);
or OR3 (N513, N510, N162, N475);
or OR4 (N514, N507, N226, N316, N268);
buf BUF1 (N515, N500);
buf BUF1 (N516, N512);
not NOT1 (N517, N511);
buf BUF1 (N518, N516);
nor NOR2 (N519, N518, N245);
and AND2 (N520, N513, N372);
xor XOR2 (N521, N484, N349);
nand NAND4 (N522, N517, N204, N464, N71);
not NOT1 (N523, N504);
xor XOR2 (N524, N520, N364);
not NOT1 (N525, N524);
and AND3 (N526, N525, N326, N503);
not NOT1 (N527, N505);
xor XOR2 (N528, N527, N510);
and AND2 (N529, N514, N298);
and AND2 (N530, N528, N284);
not NOT1 (N531, N522);
xor XOR2 (N532, N515, N148);
xor XOR2 (N533, N521, N19);
nor NOR4 (N534, N531, N280, N174, N362);
or OR2 (N535, N526, N101);
nand NAND4 (N536, N519, N153, N387, N240);
nand NAND3 (N537, N533, N223, N335);
nor NOR4 (N538, N509, N398, N515, N86);
buf BUF1 (N539, N538);
nand NAND4 (N540, N523, N76, N459, N343);
nor NOR2 (N541, N530, N22);
nand NAND2 (N542, N506, N71);
or OR3 (N543, N534, N369, N425);
nand NAND4 (N544, N540, N257, N338, N251);
xor XOR2 (N545, N536, N206);
nor NOR4 (N546, N542, N265, N191, N251);
nor NOR2 (N547, N546, N406);
nor NOR4 (N548, N537, N233, N47, N384);
nor NOR4 (N549, N545, N170, N55, N353);
nor NOR3 (N550, N529, N262, N78);
nand NAND4 (N551, N532, N261, N167, N97);
nor NOR2 (N552, N547, N501);
or OR4 (N553, N541, N288, N326, N5);
and AND4 (N554, N544, N170, N516, N283);
or OR2 (N555, N543, N307);
nand NAND3 (N556, N552, N246, N528);
or OR2 (N557, N539, N516);
xor XOR2 (N558, N557, N380);
xor XOR2 (N559, N553, N388);
buf BUF1 (N560, N551);
nor NOR3 (N561, N558, N226, N41);
or OR4 (N562, N556, N300, N234, N289);
buf BUF1 (N563, N561);
and AND3 (N564, N560, N246, N168);
buf BUF1 (N565, N555);
nor NOR3 (N566, N535, N39, N5);
nor NOR2 (N567, N559, N129);
xor XOR2 (N568, N565, N474);
xor XOR2 (N569, N562, N180);
or OR2 (N570, N549, N354);
or OR3 (N571, N569, N510, N250);
nor NOR3 (N572, N568, N567, N354);
xor XOR2 (N573, N265, N327);
not NOT1 (N574, N548);
nand NAND2 (N575, N564, N427);
and AND4 (N576, N554, N478, N505, N455);
nor NOR4 (N577, N574, N318, N281, N91);
and AND3 (N578, N566, N399, N545);
nand NAND4 (N579, N550, N248, N465, N343);
or OR4 (N580, N570, N177, N69, N293);
and AND2 (N581, N579, N147);
nand NAND2 (N582, N577, N432);
xor XOR2 (N583, N582, N223);
and AND2 (N584, N573, N319);
buf BUF1 (N585, N576);
or OR2 (N586, N583, N325);
not NOT1 (N587, N584);
and AND3 (N588, N575, N122, N358);
and AND3 (N589, N588, N236, N373);
not NOT1 (N590, N580);
nor NOR4 (N591, N563, N511, N291, N557);
not NOT1 (N592, N591);
nor NOR3 (N593, N581, N537, N586);
nor NOR4 (N594, N4, N249, N433, N520);
buf BUF1 (N595, N585);
buf BUF1 (N596, N587);
not NOT1 (N597, N578);
nor NOR2 (N598, N589, N74);
nand NAND3 (N599, N593, N560, N457);
buf BUF1 (N600, N599);
or OR3 (N601, N598, N266, N230);
or OR4 (N602, N600, N471, N387, N541);
and AND2 (N603, N596, N166);
buf BUF1 (N604, N590);
and AND3 (N605, N601, N37, N330);
nand NAND3 (N606, N603, N498, N372);
xor XOR2 (N607, N604, N31);
nand NAND2 (N608, N597, N79);
xor XOR2 (N609, N594, N71);
nor NOR2 (N610, N572, N377);
buf BUF1 (N611, N571);
and AND4 (N612, N610, N6, N174, N206);
buf BUF1 (N613, N605);
or OR4 (N614, N592, N107, N291, N253);
buf BUF1 (N615, N612);
xor XOR2 (N616, N615, N308);
or OR3 (N617, N611, N210, N180);
nand NAND2 (N618, N614, N261);
and AND2 (N619, N609, N94);
xor XOR2 (N620, N606, N83);
buf BUF1 (N621, N620);
nor NOR4 (N622, N617, N209, N46, N560);
xor XOR2 (N623, N613, N177);
xor XOR2 (N624, N622, N415);
buf BUF1 (N625, N616);
nand NAND3 (N626, N602, N316, N141);
not NOT1 (N627, N624);
or OR2 (N628, N595, N553);
nor NOR4 (N629, N618, N182, N242, N363);
buf BUF1 (N630, N621);
buf BUF1 (N631, N608);
buf BUF1 (N632, N630);
xor XOR2 (N633, N631, N421);
xor XOR2 (N634, N628, N173);
buf BUF1 (N635, N629);
buf BUF1 (N636, N634);
xor XOR2 (N637, N636, N299);
not NOT1 (N638, N632);
nand NAND2 (N639, N619, N21);
and AND3 (N640, N633, N282, N189);
xor XOR2 (N641, N639, N415);
not NOT1 (N642, N625);
buf BUF1 (N643, N627);
nor NOR3 (N644, N640, N324, N176);
nor NOR4 (N645, N643, N226, N168, N256);
not NOT1 (N646, N635);
not NOT1 (N647, N607);
nand NAND3 (N648, N623, N517, N393);
and AND2 (N649, N644, N196);
nand NAND4 (N650, N638, N322, N324, N517);
buf BUF1 (N651, N645);
nand NAND2 (N652, N641, N337);
not NOT1 (N653, N642);
buf BUF1 (N654, N651);
nor NOR2 (N655, N646, N49);
or OR3 (N656, N649, N484, N470);
not NOT1 (N657, N637);
xor XOR2 (N658, N656, N460);
and AND2 (N659, N657, N15);
and AND3 (N660, N648, N549, N538);
buf BUF1 (N661, N660);
xor XOR2 (N662, N650, N526);
not NOT1 (N663, N655);
and AND4 (N664, N661, N573, N347, N300);
not NOT1 (N665, N653);
nand NAND3 (N666, N658, N257, N368);
not NOT1 (N667, N626);
nand NAND4 (N668, N664, N123, N509, N467);
not NOT1 (N669, N663);
nor NOR3 (N670, N666, N65, N526);
nor NOR2 (N671, N652, N132);
buf BUF1 (N672, N654);
xor XOR2 (N673, N647, N339);
or OR2 (N674, N673, N631);
or OR2 (N675, N671, N338);
nor NOR4 (N676, N659, N286, N29, N619);
not NOT1 (N677, N672);
and AND4 (N678, N677, N187, N548, N302);
nor NOR4 (N679, N665, N229, N325, N157);
buf BUF1 (N680, N675);
nand NAND3 (N681, N680, N350, N150);
nor NOR2 (N682, N668, N554);
xor XOR2 (N683, N682, N71);
nor NOR3 (N684, N662, N415, N55);
xor XOR2 (N685, N667, N573);
nand NAND2 (N686, N684, N168);
xor XOR2 (N687, N686, N611);
and AND3 (N688, N681, N226, N58);
not NOT1 (N689, N685);
nand NAND3 (N690, N688, N152, N595);
nor NOR3 (N691, N674, N464, N492);
and AND3 (N692, N669, N527, N455);
or OR3 (N693, N691, N65, N178);
and AND3 (N694, N683, N197, N601);
not NOT1 (N695, N676);
nand NAND2 (N696, N679, N76);
buf BUF1 (N697, N678);
not NOT1 (N698, N689);
not NOT1 (N699, N692);
nor NOR3 (N700, N696, N356, N199);
nand NAND2 (N701, N700, N572);
and AND4 (N702, N697, N460, N464, N210);
and AND2 (N703, N687, N442);
nand NAND2 (N704, N694, N184);
buf BUF1 (N705, N703);
buf BUF1 (N706, N670);
nand NAND2 (N707, N706, N170);
buf BUF1 (N708, N690);
not NOT1 (N709, N705);
xor XOR2 (N710, N704, N323);
buf BUF1 (N711, N707);
and AND4 (N712, N709, N411, N120, N123);
not NOT1 (N713, N711);
not NOT1 (N714, N712);
or OR4 (N715, N710, N378, N153, N421);
xor XOR2 (N716, N701, N31);
and AND4 (N717, N708, N506, N258, N57);
not NOT1 (N718, N693);
and AND3 (N719, N695, N60, N497);
buf BUF1 (N720, N713);
and AND4 (N721, N719, N408, N471, N486);
nand NAND2 (N722, N721, N507);
and AND3 (N723, N699, N346, N678);
or OR2 (N724, N722, N506);
nor NOR4 (N725, N720, N236, N368, N443);
or OR3 (N726, N718, N586, N395);
not NOT1 (N727, N724);
buf BUF1 (N728, N727);
nor NOR2 (N729, N725, N206);
and AND2 (N730, N698, N30);
nand NAND4 (N731, N728, N475, N703, N525);
not NOT1 (N732, N715);
nand NAND3 (N733, N732, N35, N631);
xor XOR2 (N734, N702, N22);
or OR2 (N735, N729, N648);
not NOT1 (N736, N716);
and AND3 (N737, N717, N257, N173);
not NOT1 (N738, N733);
nand NAND3 (N739, N737, N161, N371);
xor XOR2 (N740, N734, N310);
nor NOR4 (N741, N714, N431, N449, N454);
buf BUF1 (N742, N726);
not NOT1 (N743, N738);
nor NOR4 (N744, N739, N518, N152, N735);
or OR4 (N745, N109, N211, N717, N712);
and AND4 (N746, N745, N554, N571, N394);
nand NAND4 (N747, N742, N230, N269, N378);
nand NAND3 (N748, N741, N389, N550);
xor XOR2 (N749, N743, N509);
nor NOR2 (N750, N723, N347);
nand NAND4 (N751, N731, N185, N695, N544);
and AND2 (N752, N744, N227);
nand NAND2 (N753, N748, N141);
buf BUF1 (N754, N736);
buf BUF1 (N755, N750);
xor XOR2 (N756, N746, N248);
not NOT1 (N757, N751);
xor XOR2 (N758, N756, N164);
xor XOR2 (N759, N755, N713);
or OR3 (N760, N747, N581, N192);
nand NAND2 (N761, N758, N326);
and AND4 (N762, N753, N743, N593, N729);
not NOT1 (N763, N752);
and AND4 (N764, N730, N731, N503, N353);
xor XOR2 (N765, N757, N597);
and AND2 (N766, N759, N627);
and AND4 (N767, N749, N34, N727, N501);
nor NOR3 (N768, N761, N264, N254);
or OR3 (N769, N766, N542, N469);
nor NOR3 (N770, N765, N307, N522);
xor XOR2 (N771, N769, N189);
and AND2 (N772, N767, N629);
buf BUF1 (N773, N772);
not NOT1 (N774, N740);
xor XOR2 (N775, N773, N507);
buf BUF1 (N776, N763);
or OR2 (N777, N754, N244);
xor XOR2 (N778, N768, N146);
xor XOR2 (N779, N776, N355);
and AND3 (N780, N774, N701, N119);
or OR4 (N781, N779, N599, N167, N585);
not NOT1 (N782, N771);
nand NAND4 (N783, N777, N458, N83, N556);
not NOT1 (N784, N782);
and AND2 (N785, N780, N492);
buf BUF1 (N786, N785);
xor XOR2 (N787, N786, N93);
and AND4 (N788, N778, N58, N217, N431);
or OR2 (N789, N784, N574);
nand NAND2 (N790, N760, N473);
buf BUF1 (N791, N787);
or OR3 (N792, N791, N81, N385);
nand NAND2 (N793, N781, N141);
xor XOR2 (N794, N775, N658);
buf BUF1 (N795, N790);
and AND4 (N796, N789, N308, N432, N261);
or OR4 (N797, N794, N733, N316, N242);
buf BUF1 (N798, N762);
not NOT1 (N799, N783);
nor NOR4 (N800, N793, N769, N758, N758);
xor XOR2 (N801, N788, N70);
buf BUF1 (N802, N770);
xor XOR2 (N803, N798, N26);
and AND4 (N804, N799, N374, N338, N730);
and AND3 (N805, N804, N436, N101);
buf BUF1 (N806, N792);
buf BUF1 (N807, N795);
buf BUF1 (N808, N764);
xor XOR2 (N809, N796, N657);
not NOT1 (N810, N802);
not NOT1 (N811, N810);
nor NOR4 (N812, N809, N213, N371, N430);
or OR2 (N813, N800, N627);
buf BUF1 (N814, N812);
xor XOR2 (N815, N808, N723);
nand NAND3 (N816, N807, N228, N343);
nand NAND4 (N817, N816, N443, N63, N811);
xor XOR2 (N818, N200, N753);
or OR3 (N819, N817, N368, N771);
nor NOR2 (N820, N797, N647);
nand NAND4 (N821, N814, N280, N378, N453);
nand NAND2 (N822, N820, N743);
or OR2 (N823, N819, N392);
not NOT1 (N824, N818);
nor NOR2 (N825, N823, N655);
nor NOR3 (N826, N805, N454, N479);
buf BUF1 (N827, N822);
or OR2 (N828, N806, N451);
nor NOR4 (N829, N821, N395, N752, N515);
xor XOR2 (N830, N825, N725);
not NOT1 (N831, N827);
buf BUF1 (N832, N813);
or OR2 (N833, N803, N269);
or OR3 (N834, N828, N794, N230);
xor XOR2 (N835, N826, N236);
and AND3 (N836, N834, N783, N688);
buf BUF1 (N837, N801);
nor NOR3 (N838, N815, N271, N625);
or OR4 (N839, N832, N116, N283, N813);
not NOT1 (N840, N830);
not NOT1 (N841, N829);
and AND3 (N842, N831, N572, N84);
or OR2 (N843, N836, N620);
xor XOR2 (N844, N838, N556);
buf BUF1 (N845, N841);
buf BUF1 (N846, N833);
not NOT1 (N847, N846);
nand NAND2 (N848, N844, N194);
buf BUF1 (N849, N835);
xor XOR2 (N850, N837, N211);
nand NAND2 (N851, N843, N124);
or OR4 (N852, N848, N138, N616, N444);
and AND4 (N853, N852, N552, N404, N802);
and AND4 (N854, N849, N464, N357, N71);
xor XOR2 (N855, N840, N609);
nand NAND4 (N856, N853, N838, N591, N335);
and AND2 (N857, N856, N361);
or OR3 (N858, N839, N815, N539);
nand NAND4 (N859, N824, N195, N454, N166);
or OR3 (N860, N855, N235, N240);
nand NAND3 (N861, N857, N446, N159);
buf BUF1 (N862, N850);
nor NOR2 (N863, N860, N101);
or OR2 (N864, N842, N165);
not NOT1 (N865, N858);
and AND3 (N866, N854, N192, N70);
or OR3 (N867, N845, N655, N595);
buf BUF1 (N868, N867);
and AND4 (N869, N847, N15, N25, N137);
buf BUF1 (N870, N869);
nor NOR2 (N871, N865, N96);
or OR4 (N872, N870, N314, N777, N486);
buf BUF1 (N873, N866);
xor XOR2 (N874, N873, N200);
nand NAND3 (N875, N861, N269, N511);
and AND4 (N876, N864, N193, N419, N148);
nand NAND3 (N877, N862, N820, N425);
not NOT1 (N878, N851);
or OR2 (N879, N876, N449);
not NOT1 (N880, N875);
nor NOR4 (N881, N874, N28, N567, N855);
xor XOR2 (N882, N878, N56);
and AND3 (N883, N880, N712, N755);
nand NAND4 (N884, N879, N688, N5, N337);
not NOT1 (N885, N881);
nor NOR2 (N886, N885, N432);
nand NAND4 (N887, N871, N170, N296, N104);
xor XOR2 (N888, N884, N760);
buf BUF1 (N889, N868);
xor XOR2 (N890, N859, N458);
nand NAND4 (N891, N882, N610, N390, N422);
nand NAND4 (N892, N887, N339, N3, N719);
nand NAND2 (N893, N890, N225);
not NOT1 (N894, N889);
buf BUF1 (N895, N894);
buf BUF1 (N896, N892);
and AND2 (N897, N895, N699);
buf BUF1 (N898, N863);
nor NOR3 (N899, N897, N162, N387);
nor NOR2 (N900, N886, N31);
xor XOR2 (N901, N900, N107);
buf BUF1 (N902, N898);
nor NOR2 (N903, N899, N708);
and AND2 (N904, N888, N708);
or OR2 (N905, N872, N68);
nand NAND4 (N906, N905, N274, N499, N785);
buf BUF1 (N907, N903);
xor XOR2 (N908, N901, N805);
and AND2 (N909, N906, N573);
and AND2 (N910, N883, N680);
xor XOR2 (N911, N908, N402);
xor XOR2 (N912, N910, N155);
nand NAND2 (N913, N911, N248);
and AND3 (N914, N896, N705, N95);
or OR4 (N915, N913, N122, N95, N844);
buf BUF1 (N916, N902);
not NOT1 (N917, N914);
and AND2 (N918, N877, N347);
xor XOR2 (N919, N916, N40);
not NOT1 (N920, N893);
or OR2 (N921, N918, N436);
or OR2 (N922, N912, N620);
buf BUF1 (N923, N915);
or OR2 (N924, N920, N902);
and AND4 (N925, N907, N514, N479, N101);
buf BUF1 (N926, N909);
xor XOR2 (N927, N922, N263);
xor XOR2 (N928, N926, N458);
not NOT1 (N929, N921);
buf BUF1 (N930, N923);
buf BUF1 (N931, N924);
or OR4 (N932, N904, N724, N201, N685);
or OR4 (N933, N930, N381, N671, N717);
nor NOR2 (N934, N932, N83);
buf BUF1 (N935, N927);
nand NAND2 (N936, N891, N517);
not NOT1 (N937, N925);
not NOT1 (N938, N933);
and AND3 (N939, N928, N723, N785);
nand NAND3 (N940, N936, N4, N461);
buf BUF1 (N941, N937);
nor NOR4 (N942, N917, N738, N545, N125);
nand NAND4 (N943, N929, N668, N835, N877);
buf BUF1 (N944, N935);
and AND4 (N945, N919, N179, N864, N769);
nand NAND3 (N946, N944, N48, N305);
and AND4 (N947, N940, N352, N530, N312);
buf BUF1 (N948, N945);
nand NAND3 (N949, N931, N38, N614);
and AND3 (N950, N938, N224, N314);
nor NOR4 (N951, N941, N81, N869, N227);
xor XOR2 (N952, N950, N941);
buf BUF1 (N953, N942);
nor NOR2 (N954, N952, N743);
buf BUF1 (N955, N946);
not NOT1 (N956, N955);
not NOT1 (N957, N951);
and AND2 (N958, N934, N954);
nand NAND4 (N959, N161, N520, N53, N806);
nand NAND2 (N960, N949, N648);
nand NAND4 (N961, N960, N940, N426, N386);
buf BUF1 (N962, N961);
nor NOR2 (N963, N959, N313);
xor XOR2 (N964, N953, N746);
nand NAND2 (N965, N964, N620);
xor XOR2 (N966, N958, N280);
and AND4 (N967, N963, N773, N414, N591);
or OR2 (N968, N967, N368);
nand NAND3 (N969, N966, N721, N847);
buf BUF1 (N970, N947);
buf BUF1 (N971, N970);
nor NOR2 (N972, N939, N9);
nor NOR3 (N973, N968, N792, N648);
buf BUF1 (N974, N971);
and AND2 (N975, N965, N174);
and AND4 (N976, N969, N934, N382, N190);
not NOT1 (N977, N957);
nor NOR4 (N978, N948, N974, N791, N317);
nand NAND2 (N979, N37, N102);
xor XOR2 (N980, N973, N685);
buf BUF1 (N981, N956);
not NOT1 (N982, N962);
not NOT1 (N983, N981);
xor XOR2 (N984, N980, N678);
and AND4 (N985, N972, N844, N273, N246);
xor XOR2 (N986, N985, N341);
not NOT1 (N987, N976);
or OR4 (N988, N979, N509, N312, N986);
not NOT1 (N989, N186);
nand NAND2 (N990, N987, N298);
not NOT1 (N991, N990);
or OR3 (N992, N984, N1, N16);
or OR3 (N993, N988, N720, N394);
nand NAND4 (N994, N977, N766, N898, N418);
not NOT1 (N995, N982);
nor NOR2 (N996, N991, N831);
buf BUF1 (N997, N989);
not NOT1 (N998, N995);
nand NAND2 (N999, N983, N282);
buf BUF1 (N1000, N997);
xor XOR2 (N1001, N975, N265);
not NOT1 (N1002, N1000);
nor NOR4 (N1003, N1002, N652, N788, N787);
not NOT1 (N1004, N1001);
buf BUF1 (N1005, N996);
buf BUF1 (N1006, N998);
not NOT1 (N1007, N992);
and AND2 (N1008, N999, N26);
buf BUF1 (N1009, N978);
not NOT1 (N1010, N1005);
buf BUF1 (N1011, N1009);
and AND3 (N1012, N943, N602, N103);
xor XOR2 (N1013, N1012, N933);
buf BUF1 (N1014, N1008);
buf BUF1 (N1015, N1011);
not NOT1 (N1016, N1003);
nor NOR4 (N1017, N1013, N468, N921, N990);
xor XOR2 (N1018, N993, N210);
buf BUF1 (N1019, N1017);
and AND2 (N1020, N1010, N249);
nor NOR4 (N1021, N1015, N927, N817, N145);
buf BUF1 (N1022, N1004);
not NOT1 (N1023, N1021);
buf BUF1 (N1024, N1023);
or OR4 (N1025, N1014, N1024, N433, N555);
or OR3 (N1026, N441, N299, N106);
and AND2 (N1027, N1019, N29);
and AND3 (N1028, N1027, N921, N802);
not NOT1 (N1029, N1006);
buf BUF1 (N1030, N1016);
nand NAND3 (N1031, N1030, N344, N1025);
nand NAND4 (N1032, N457, N706, N113, N825);
not NOT1 (N1033, N994);
nand NAND2 (N1034, N1007, N779);
xor XOR2 (N1035, N1028, N800);
or OR2 (N1036, N1029, N969);
nand NAND4 (N1037, N1032, N812, N358, N449);
nor NOR4 (N1038, N1018, N295, N427, N825);
buf BUF1 (N1039, N1034);
nand NAND4 (N1040, N1031, N625, N4, N1023);
buf BUF1 (N1041, N1040);
or OR3 (N1042, N1035, N608, N511);
xor XOR2 (N1043, N1038, N334);
nor NOR4 (N1044, N1022, N395, N590, N601);
xor XOR2 (N1045, N1042, N874);
not NOT1 (N1046, N1039);
and AND2 (N1047, N1033, N167);
or OR2 (N1048, N1045, N224);
not NOT1 (N1049, N1036);
xor XOR2 (N1050, N1044, N785);
not NOT1 (N1051, N1037);
not NOT1 (N1052, N1047);
or OR3 (N1053, N1041, N61, N342);
nand NAND4 (N1054, N1046, N347, N609, N253);
nand NAND3 (N1055, N1053, N502, N173);
buf BUF1 (N1056, N1020);
nor NOR2 (N1057, N1052, N773);
buf BUF1 (N1058, N1057);
buf BUF1 (N1059, N1049);
buf BUF1 (N1060, N1051);
xor XOR2 (N1061, N1048, N34);
xor XOR2 (N1062, N1059, N217);
nor NOR2 (N1063, N1058, N1037);
not NOT1 (N1064, N1055);
xor XOR2 (N1065, N1063, N721);
not NOT1 (N1066, N1060);
nand NAND3 (N1067, N1050, N55, N823);
nor NOR3 (N1068, N1066, N392, N398);
nor NOR3 (N1069, N1064, N524, N27);
not NOT1 (N1070, N1069);
buf BUF1 (N1071, N1062);
not NOT1 (N1072, N1067);
not NOT1 (N1073, N1071);
buf BUF1 (N1074, N1073);
or OR4 (N1075, N1072, N505, N870, N889);
buf BUF1 (N1076, N1075);
nor NOR2 (N1077, N1054, N937);
or OR4 (N1078, N1056, N531, N737, N686);
xor XOR2 (N1079, N1077, N152);
buf BUF1 (N1080, N1070);
and AND3 (N1081, N1074, N16, N956);
not NOT1 (N1082, N1076);
not NOT1 (N1083, N1068);
xor XOR2 (N1084, N1080, N548);
xor XOR2 (N1085, N1084, N47);
nand NAND3 (N1086, N1061, N225, N250);
not NOT1 (N1087, N1086);
nand NAND3 (N1088, N1085, N448, N454);
nand NAND2 (N1089, N1078, N1031);
nand NAND3 (N1090, N1088, N260, N287);
not NOT1 (N1091, N1090);
nor NOR4 (N1092, N1081, N1000, N142, N857);
nor NOR4 (N1093, N1091, N700, N942, N703);
nor NOR3 (N1094, N1093, N155, N230);
not NOT1 (N1095, N1082);
not NOT1 (N1096, N1065);
xor XOR2 (N1097, N1095, N1083);
nor NOR3 (N1098, N607, N838, N787);
xor XOR2 (N1099, N1098, N1044);
xor XOR2 (N1100, N1089, N449);
not NOT1 (N1101, N1092);
buf BUF1 (N1102, N1079);
or OR4 (N1103, N1094, N50, N860, N101);
xor XOR2 (N1104, N1087, N712);
nand NAND3 (N1105, N1102, N360, N298);
not NOT1 (N1106, N1026);
not NOT1 (N1107, N1104);
or OR3 (N1108, N1099, N1083, N25);
or OR4 (N1109, N1108, N575, N869, N546);
and AND2 (N1110, N1107, N1069);
or OR3 (N1111, N1109, N528, N381);
nand NAND2 (N1112, N1101, N455);
nand NAND4 (N1113, N1096, N569, N993, N430);
or OR4 (N1114, N1111, N323, N930, N1029);
nor NOR4 (N1115, N1100, N415, N341, N240);
buf BUF1 (N1116, N1097);
nand NAND3 (N1117, N1103, N842, N398);
and AND3 (N1118, N1116, N147, N837);
nor NOR3 (N1119, N1043, N30, N284);
or OR3 (N1120, N1105, N324, N227);
buf BUF1 (N1121, N1118);
buf BUF1 (N1122, N1112);
not NOT1 (N1123, N1106);
not NOT1 (N1124, N1115);
not NOT1 (N1125, N1122);
buf BUF1 (N1126, N1113);
nor NOR3 (N1127, N1123, N713, N1008);
and AND4 (N1128, N1127, N962, N166, N128);
xor XOR2 (N1129, N1120, N428);
xor XOR2 (N1130, N1119, N726);
not NOT1 (N1131, N1129);
xor XOR2 (N1132, N1121, N162);
buf BUF1 (N1133, N1124);
nor NOR2 (N1134, N1130, N381);
xor XOR2 (N1135, N1114, N945);
nor NOR3 (N1136, N1125, N240, N983);
buf BUF1 (N1137, N1126);
buf BUF1 (N1138, N1128);
not NOT1 (N1139, N1136);
or OR4 (N1140, N1135, N469, N1090, N911);
nor NOR4 (N1141, N1117, N749, N153, N617);
and AND3 (N1142, N1131, N1047, N132);
buf BUF1 (N1143, N1132);
or OR3 (N1144, N1133, N1137, N457);
xor XOR2 (N1145, N1067, N1121);
nand NAND4 (N1146, N1110, N1121, N278, N93);
or OR3 (N1147, N1138, N557, N84);
nor NOR3 (N1148, N1143, N366, N944);
xor XOR2 (N1149, N1144, N1070);
xor XOR2 (N1150, N1134, N800);
or OR4 (N1151, N1147, N150, N644, N235);
nor NOR4 (N1152, N1150, N819, N319, N63);
buf BUF1 (N1153, N1142);
or OR3 (N1154, N1146, N101, N447);
xor XOR2 (N1155, N1141, N529);
xor XOR2 (N1156, N1145, N342);
and AND4 (N1157, N1151, N1053, N221, N228);
and AND3 (N1158, N1153, N92, N10);
or OR4 (N1159, N1154, N11, N1017, N172);
nor NOR3 (N1160, N1158, N193, N828);
or OR2 (N1161, N1140, N1127);
nor NOR3 (N1162, N1148, N1118, N430);
buf BUF1 (N1163, N1152);
or OR4 (N1164, N1139, N465, N1150, N358);
xor XOR2 (N1165, N1161, N852);
nor NOR3 (N1166, N1165, N296, N1090);
nand NAND2 (N1167, N1157, N117);
nand NAND3 (N1168, N1160, N982, N177);
buf BUF1 (N1169, N1164);
nand NAND2 (N1170, N1166, N260);
and AND3 (N1171, N1162, N564, N552);
xor XOR2 (N1172, N1155, N274);
buf BUF1 (N1173, N1149);
not NOT1 (N1174, N1173);
xor XOR2 (N1175, N1174, N573);
and AND2 (N1176, N1163, N594);
xor XOR2 (N1177, N1170, N629);
and AND2 (N1178, N1172, N632);
nand NAND2 (N1179, N1171, N1177);
not NOT1 (N1180, N427);
nand NAND4 (N1181, N1178, N732, N1089, N1164);
buf BUF1 (N1182, N1181);
buf BUF1 (N1183, N1179);
or OR3 (N1184, N1169, N924, N833);
nand NAND2 (N1185, N1159, N517);
not NOT1 (N1186, N1180);
or OR2 (N1187, N1185, N612);
nand NAND2 (N1188, N1186, N834);
and AND2 (N1189, N1183, N263);
not NOT1 (N1190, N1188);
buf BUF1 (N1191, N1176);
nor NOR3 (N1192, N1182, N1047, N236);
nor NOR2 (N1193, N1189, N49);
not NOT1 (N1194, N1167);
buf BUF1 (N1195, N1168);
nand NAND4 (N1196, N1156, N139, N568, N946);
buf BUF1 (N1197, N1190);
nor NOR2 (N1198, N1195, N584);
nand NAND2 (N1199, N1184, N1170);
not NOT1 (N1200, N1196);
buf BUF1 (N1201, N1197);
or OR3 (N1202, N1193, N366, N306);
or OR3 (N1203, N1201, N1079, N989);
and AND4 (N1204, N1203, N198, N506, N1139);
and AND3 (N1205, N1200, N822, N1174);
nand NAND4 (N1206, N1192, N912, N626, N13);
and AND2 (N1207, N1204, N195);
and AND3 (N1208, N1207, N200, N337);
xor XOR2 (N1209, N1191, N845);
buf BUF1 (N1210, N1198);
not NOT1 (N1211, N1202);
nor NOR3 (N1212, N1208, N24, N1168);
and AND4 (N1213, N1187, N943, N926, N944);
not NOT1 (N1214, N1175);
not NOT1 (N1215, N1209);
xor XOR2 (N1216, N1212, N97);
not NOT1 (N1217, N1215);
nand NAND4 (N1218, N1199, N1185, N847, N913);
nand NAND2 (N1219, N1213, N483);
nor NOR3 (N1220, N1216, N806, N365);
not NOT1 (N1221, N1194);
not NOT1 (N1222, N1219);
nand NAND4 (N1223, N1206, N1016, N167, N867);
not NOT1 (N1224, N1218);
xor XOR2 (N1225, N1224, N1106);
not NOT1 (N1226, N1214);
and AND2 (N1227, N1217, N857);
xor XOR2 (N1228, N1227, N273);
nand NAND3 (N1229, N1222, N225, N290);
not NOT1 (N1230, N1226);
buf BUF1 (N1231, N1210);
buf BUF1 (N1232, N1229);
nor NOR4 (N1233, N1232, N1166, N1086, N1001);
and AND2 (N1234, N1205, N1016);
nand NAND3 (N1235, N1231, N465, N904);
nand NAND4 (N1236, N1211, N1126, N309, N797);
xor XOR2 (N1237, N1233, N1044);
xor XOR2 (N1238, N1220, N280);
and AND2 (N1239, N1221, N357);
or OR3 (N1240, N1230, N689, N918);
xor XOR2 (N1241, N1237, N1147);
xor XOR2 (N1242, N1223, N119);
buf BUF1 (N1243, N1242);
nor NOR3 (N1244, N1228, N487, N763);
nor NOR4 (N1245, N1236, N64, N8, N891);
not NOT1 (N1246, N1244);
xor XOR2 (N1247, N1235, N510);
and AND3 (N1248, N1225, N1022, N462);
nand NAND2 (N1249, N1240, N330);
or OR2 (N1250, N1241, N25);
and AND2 (N1251, N1234, N790);
or OR3 (N1252, N1249, N485, N763);
xor XOR2 (N1253, N1239, N123);
buf BUF1 (N1254, N1248);
and AND4 (N1255, N1243, N940, N154, N880);
buf BUF1 (N1256, N1255);
or OR2 (N1257, N1247, N1032);
xor XOR2 (N1258, N1238, N443);
nand NAND2 (N1259, N1246, N150);
nand NAND3 (N1260, N1256, N116, N353);
nor NOR2 (N1261, N1254, N546);
and AND3 (N1262, N1261, N110, N1082);
xor XOR2 (N1263, N1259, N1006);
xor XOR2 (N1264, N1258, N142);
or OR3 (N1265, N1257, N657, N1046);
not NOT1 (N1266, N1263);
nand NAND2 (N1267, N1262, N839);
or OR3 (N1268, N1250, N1018, N1115);
or OR2 (N1269, N1267, N672);
buf BUF1 (N1270, N1251);
and AND3 (N1271, N1269, N763, N1162);
not NOT1 (N1272, N1271);
not NOT1 (N1273, N1266);
xor XOR2 (N1274, N1253, N221);
nand NAND4 (N1275, N1264, N176, N1099, N228);
nand NAND3 (N1276, N1272, N692, N71);
nand NAND2 (N1277, N1273, N1272);
or OR2 (N1278, N1277, N130);
not NOT1 (N1279, N1260);
and AND2 (N1280, N1274, N643);
nor NOR2 (N1281, N1245, N982);
nand NAND3 (N1282, N1270, N98, N875);
xor XOR2 (N1283, N1252, N526);
not NOT1 (N1284, N1275);
or OR3 (N1285, N1268, N603, N656);
not NOT1 (N1286, N1281);
nand NAND4 (N1287, N1283, N446, N765, N849);
nor NOR4 (N1288, N1285, N190, N74, N953);
or OR3 (N1289, N1265, N1258, N942);
buf BUF1 (N1290, N1284);
or OR4 (N1291, N1286, N560, N824, N264);
nor NOR3 (N1292, N1291, N247, N94);
buf BUF1 (N1293, N1290);
xor XOR2 (N1294, N1279, N88);
buf BUF1 (N1295, N1287);
buf BUF1 (N1296, N1295);
and AND3 (N1297, N1278, N1223, N180);
or OR3 (N1298, N1282, N477, N1096);
buf BUF1 (N1299, N1292);
or OR3 (N1300, N1294, N775, N1200);
not NOT1 (N1301, N1298);
xor XOR2 (N1302, N1301, N586);
buf BUF1 (N1303, N1293);
nor NOR2 (N1304, N1297, N1014);
nand NAND4 (N1305, N1300, N1119, N1139, N1009);
buf BUF1 (N1306, N1276);
or OR2 (N1307, N1299, N165);
not NOT1 (N1308, N1305);
not NOT1 (N1309, N1306);
nor NOR4 (N1310, N1308, N666, N814, N223);
buf BUF1 (N1311, N1307);
and AND2 (N1312, N1288, N812);
buf BUF1 (N1313, N1310);
nor NOR4 (N1314, N1311, N788, N720, N411);
not NOT1 (N1315, N1313);
and AND3 (N1316, N1302, N350, N374);
and AND3 (N1317, N1280, N261, N602);
nand NAND2 (N1318, N1314, N422);
buf BUF1 (N1319, N1304);
not NOT1 (N1320, N1309);
not NOT1 (N1321, N1316);
xor XOR2 (N1322, N1312, N1239);
nand NAND4 (N1323, N1315, N455, N903, N675);
nand NAND2 (N1324, N1320, N1093);
not NOT1 (N1325, N1324);
and AND3 (N1326, N1296, N423, N1290);
nand NAND4 (N1327, N1303, N380, N661, N970);
xor XOR2 (N1328, N1319, N685);
and AND3 (N1329, N1317, N908, N249);
or OR2 (N1330, N1325, N435);
buf BUF1 (N1331, N1323);
and AND3 (N1332, N1331, N926, N887);
and AND2 (N1333, N1328, N1012);
buf BUF1 (N1334, N1322);
nand NAND4 (N1335, N1330, N670, N1277, N930);
nand NAND2 (N1336, N1334, N1178);
buf BUF1 (N1337, N1321);
xor XOR2 (N1338, N1329, N52);
nand NAND2 (N1339, N1338, N221);
and AND2 (N1340, N1335, N1175);
nand NAND2 (N1341, N1340, N179);
and AND3 (N1342, N1289, N27, N92);
buf BUF1 (N1343, N1327);
nand NAND2 (N1344, N1333, N138);
not NOT1 (N1345, N1343);
buf BUF1 (N1346, N1344);
xor XOR2 (N1347, N1336, N128);
not NOT1 (N1348, N1332);
nand NAND3 (N1349, N1326, N789, N1068);
or OR3 (N1350, N1341, N253, N335);
or OR3 (N1351, N1346, N1296, N197);
not NOT1 (N1352, N1345);
and AND2 (N1353, N1352, N248);
not NOT1 (N1354, N1318);
buf BUF1 (N1355, N1342);
xor XOR2 (N1356, N1348, N357);
or OR2 (N1357, N1337, N1093);
not NOT1 (N1358, N1349);
xor XOR2 (N1359, N1354, N436);
nor NOR3 (N1360, N1339, N77, N833);
or OR2 (N1361, N1357, N622);
nand NAND4 (N1362, N1351, N1122, N1117, N554);
or OR3 (N1363, N1350, N817, N1042);
nand NAND4 (N1364, N1353, N465, N34, N609);
nor NOR2 (N1365, N1355, N141);
not NOT1 (N1366, N1365);
nand NAND3 (N1367, N1366, N316, N1042);
not NOT1 (N1368, N1359);
or OR4 (N1369, N1367, N809, N825, N172);
nor NOR4 (N1370, N1362, N487, N941, N919);
buf BUF1 (N1371, N1368);
buf BUF1 (N1372, N1371);
and AND2 (N1373, N1360, N1241);
not NOT1 (N1374, N1373);
xor XOR2 (N1375, N1363, N202);
buf BUF1 (N1376, N1361);
and AND3 (N1377, N1358, N975, N1223);
nor NOR3 (N1378, N1347, N819, N532);
nor NOR2 (N1379, N1374, N1061);
buf BUF1 (N1380, N1372);
xor XOR2 (N1381, N1378, N912);
and AND2 (N1382, N1364, N245);
nand NAND2 (N1383, N1370, N417);
xor XOR2 (N1384, N1383, N981);
nand NAND2 (N1385, N1379, N391);
nand NAND4 (N1386, N1375, N504, N1121, N1372);
xor XOR2 (N1387, N1380, N998);
nand NAND4 (N1388, N1386, N672, N528, N1369);
nor NOR3 (N1389, N265, N259, N312);
not NOT1 (N1390, N1377);
xor XOR2 (N1391, N1376, N1145);
nor NOR2 (N1392, N1388, N837);
buf BUF1 (N1393, N1391);
nor NOR2 (N1394, N1392, N404);
buf BUF1 (N1395, N1356);
or OR3 (N1396, N1384, N78, N804);
or OR2 (N1397, N1395, N247);
and AND2 (N1398, N1393, N1336);
or OR3 (N1399, N1389, N965, N404);
nor NOR4 (N1400, N1390, N97, N1212, N938);
buf BUF1 (N1401, N1397);
not NOT1 (N1402, N1400);
nand NAND2 (N1403, N1398, N349);
not NOT1 (N1404, N1396);
or OR4 (N1405, N1387, N562, N604, N411);
or OR2 (N1406, N1382, N400);
not NOT1 (N1407, N1403);
nor NOR3 (N1408, N1405, N603, N1389);
and AND3 (N1409, N1399, N413, N1381);
buf BUF1 (N1410, N475);
or OR2 (N1411, N1394, N1132);
buf BUF1 (N1412, N1409);
xor XOR2 (N1413, N1401, N911);
nor NOR4 (N1414, N1408, N238, N997, N491);
xor XOR2 (N1415, N1407, N30);
nor NOR4 (N1416, N1415, N682, N341, N1244);
nor NOR3 (N1417, N1416, N191, N1051);
nor NOR4 (N1418, N1414, N1004, N588, N1152);
buf BUF1 (N1419, N1411);
xor XOR2 (N1420, N1410, N316);
nand NAND4 (N1421, N1417, N61, N1152, N130);
or OR2 (N1422, N1413, N945);
buf BUF1 (N1423, N1385);
nor NOR4 (N1424, N1422, N15, N1304, N32);
and AND3 (N1425, N1420, N582, N689);
or OR3 (N1426, N1425, N792, N951);
nand NAND2 (N1427, N1412, N893);
or OR2 (N1428, N1402, N119);
xor XOR2 (N1429, N1419, N1129);
and AND2 (N1430, N1428, N1133);
buf BUF1 (N1431, N1427);
not NOT1 (N1432, N1418);
not NOT1 (N1433, N1424);
not NOT1 (N1434, N1430);
nor NOR3 (N1435, N1406, N1360, N57);
nor NOR4 (N1436, N1432, N1193, N770, N108);
or OR2 (N1437, N1429, N555);
or OR2 (N1438, N1423, N198);
not NOT1 (N1439, N1435);
xor XOR2 (N1440, N1438, N1357);
nand NAND3 (N1441, N1436, N266, N285);
nor NOR4 (N1442, N1437, N969, N371, N326);
or OR3 (N1443, N1440, N709, N1136);
nor NOR3 (N1444, N1431, N538, N305);
and AND4 (N1445, N1439, N1285, N917, N1422);
nand NAND4 (N1446, N1404, N11, N310, N406);
or OR4 (N1447, N1442, N386, N725, N1344);
xor XOR2 (N1448, N1434, N685);
or OR4 (N1449, N1444, N1237, N250, N1178);
nor NOR4 (N1450, N1441, N1108, N1063, N197);
nor NOR4 (N1451, N1426, N1142, N378, N535);
not NOT1 (N1452, N1433);
xor XOR2 (N1453, N1452, N364);
nor NOR2 (N1454, N1446, N786);
nor NOR2 (N1455, N1447, N341);
xor XOR2 (N1456, N1451, N272);
nor NOR2 (N1457, N1449, N877);
nand NAND2 (N1458, N1443, N340);
or OR3 (N1459, N1421, N481, N835);
and AND3 (N1460, N1457, N574, N79);
not NOT1 (N1461, N1454);
and AND3 (N1462, N1461, N261, N1040);
and AND4 (N1463, N1456, N623, N1162, N627);
nand NAND4 (N1464, N1460, N1415, N1341, N549);
or OR4 (N1465, N1445, N464, N1452, N929);
not NOT1 (N1466, N1463);
or OR2 (N1467, N1466, N491);
xor XOR2 (N1468, N1450, N1208);
nor NOR4 (N1469, N1464, N255, N1374, N1380);
xor XOR2 (N1470, N1458, N697);
and AND4 (N1471, N1468, N957, N161, N357);
xor XOR2 (N1472, N1459, N100);
or OR4 (N1473, N1465, N138, N1156, N1265);
and AND4 (N1474, N1469, N1102, N110, N695);
buf BUF1 (N1475, N1472);
nor NOR3 (N1476, N1474, N1390, N1213);
and AND2 (N1477, N1475, N1343);
not NOT1 (N1478, N1448);
not NOT1 (N1479, N1471);
xor XOR2 (N1480, N1453, N1243);
nor NOR3 (N1481, N1480, N330, N527);
not NOT1 (N1482, N1481);
or OR3 (N1483, N1479, N322, N157);
nor NOR3 (N1484, N1473, N79, N577);
and AND4 (N1485, N1462, N777, N824, N893);
and AND3 (N1486, N1485, N277, N264);
xor XOR2 (N1487, N1486, N1103);
nor NOR4 (N1488, N1478, N1009, N1060, N1410);
xor XOR2 (N1489, N1467, N236);
nor NOR3 (N1490, N1489, N701, N36);
xor XOR2 (N1491, N1484, N66);
or OR2 (N1492, N1482, N1173);
xor XOR2 (N1493, N1492, N461);
and AND3 (N1494, N1493, N922, N1395);
or OR4 (N1495, N1490, N1033, N932, N261);
or OR2 (N1496, N1477, N1332);
not NOT1 (N1497, N1487);
or OR3 (N1498, N1494, N1020, N249);
nand NAND2 (N1499, N1498, N1298);
buf BUF1 (N1500, N1476);
nor NOR4 (N1501, N1455, N507, N1362, N865);
xor XOR2 (N1502, N1491, N327);
buf BUF1 (N1503, N1500);
or OR4 (N1504, N1502, N59, N876, N1210);
and AND2 (N1505, N1504, N676);
not NOT1 (N1506, N1501);
and AND2 (N1507, N1506, N615);
xor XOR2 (N1508, N1496, N301);
nand NAND2 (N1509, N1470, N1382);
or OR4 (N1510, N1505, N1243, N1474, N817);
nor NOR4 (N1511, N1509, N1155, N442, N161);
not NOT1 (N1512, N1510);
and AND4 (N1513, N1503, N1067, N115, N1377);
nor NOR2 (N1514, N1497, N1259);
and AND2 (N1515, N1507, N449);
nand NAND3 (N1516, N1512, N830, N1438);
and AND4 (N1517, N1516, N657, N562, N1045);
not NOT1 (N1518, N1508);
not NOT1 (N1519, N1483);
or OR3 (N1520, N1518, N110, N1156);
nand NAND4 (N1521, N1495, N650, N803, N81);
and AND2 (N1522, N1488, N248);
or OR4 (N1523, N1521, N1359, N360, N1256);
xor XOR2 (N1524, N1513, N1158);
xor XOR2 (N1525, N1499, N963);
nand NAND4 (N1526, N1524, N1481, N1125, N236);
nor NOR3 (N1527, N1522, N1211, N280);
or OR3 (N1528, N1515, N839, N439);
and AND3 (N1529, N1517, N756, N890);
xor XOR2 (N1530, N1519, N505);
nand NAND3 (N1531, N1528, N127, N286);
nor NOR3 (N1532, N1527, N1458, N1219);
and AND3 (N1533, N1530, N1460, N718);
or OR4 (N1534, N1533, N100, N714, N1022);
not NOT1 (N1535, N1534);
xor XOR2 (N1536, N1526, N572);
nor NOR3 (N1537, N1514, N975, N177);
or OR3 (N1538, N1532, N58, N468);
nand NAND2 (N1539, N1523, N1330);
or OR2 (N1540, N1536, N225);
nand NAND3 (N1541, N1529, N1111, N1074);
or OR2 (N1542, N1531, N997);
buf BUF1 (N1543, N1525);
nor NOR3 (N1544, N1537, N322, N1326);
or OR4 (N1545, N1541, N675, N1125, N452);
or OR4 (N1546, N1535, N429, N1327, N1209);
and AND2 (N1547, N1542, N920);
and AND3 (N1548, N1544, N385, N798);
or OR2 (N1549, N1547, N768);
xor XOR2 (N1550, N1540, N919);
xor XOR2 (N1551, N1538, N867);
nand NAND3 (N1552, N1543, N662, N1345);
and AND3 (N1553, N1549, N1243, N223);
and AND4 (N1554, N1520, N70, N1141, N1467);
xor XOR2 (N1555, N1553, N1425);
buf BUF1 (N1556, N1552);
nor NOR3 (N1557, N1556, N1138, N1125);
nand NAND3 (N1558, N1545, N818, N491);
or OR4 (N1559, N1550, N181, N491, N258);
not NOT1 (N1560, N1551);
or OR2 (N1561, N1546, N1432);
nor NOR3 (N1562, N1561, N1324, N621);
and AND3 (N1563, N1539, N1171, N583);
nor NOR2 (N1564, N1558, N409);
and AND4 (N1565, N1564, N92, N1138, N37);
nor NOR4 (N1566, N1511, N568, N1327, N1022);
nand NAND4 (N1567, N1566, N1362, N749, N1072);
nand NAND2 (N1568, N1548, N1139);
buf BUF1 (N1569, N1568);
xor XOR2 (N1570, N1569, N400);
not NOT1 (N1571, N1554);
or OR4 (N1572, N1571, N1074, N1435, N1034);
not NOT1 (N1573, N1565);
or OR3 (N1574, N1567, N1364, N755);
nor NOR3 (N1575, N1573, N885, N533);
or OR3 (N1576, N1574, N824, N319);
not NOT1 (N1577, N1559);
and AND2 (N1578, N1563, N21);
and AND3 (N1579, N1557, N1554, N348);
not NOT1 (N1580, N1578);
not NOT1 (N1581, N1580);
or OR3 (N1582, N1562, N401, N1029);
xor XOR2 (N1583, N1555, N658);
nor NOR3 (N1584, N1583, N1201, N363);
nor NOR2 (N1585, N1577, N943);
not NOT1 (N1586, N1584);
not NOT1 (N1587, N1570);
nand NAND3 (N1588, N1585, N1430, N1177);
or OR4 (N1589, N1576, N544, N312, N1116);
nor NOR3 (N1590, N1588, N1119, N578);
or OR4 (N1591, N1572, N251, N1386, N600);
buf BUF1 (N1592, N1582);
xor XOR2 (N1593, N1586, N996);
not NOT1 (N1594, N1592);
or OR2 (N1595, N1581, N406);
not NOT1 (N1596, N1590);
or OR3 (N1597, N1596, N270, N80);
nor NOR3 (N1598, N1579, N726, N742);
nor NOR3 (N1599, N1598, N723, N512);
nor NOR4 (N1600, N1591, N1174, N164, N1351);
not NOT1 (N1601, N1600);
xor XOR2 (N1602, N1587, N574);
and AND4 (N1603, N1593, N1155, N249, N543);
or OR3 (N1604, N1589, N58, N1424);
xor XOR2 (N1605, N1603, N1429);
not NOT1 (N1606, N1597);
nor NOR3 (N1607, N1595, N1285, N823);
nand NAND4 (N1608, N1606, N337, N1066, N507);
xor XOR2 (N1609, N1575, N397);
not NOT1 (N1610, N1609);
not NOT1 (N1611, N1601);
or OR2 (N1612, N1605, N933);
nand NAND4 (N1613, N1599, N1324, N429, N1478);
and AND2 (N1614, N1602, N495);
not NOT1 (N1615, N1594);
xor XOR2 (N1616, N1614, N1556);
or OR2 (N1617, N1608, N1491);
xor XOR2 (N1618, N1612, N1059);
xor XOR2 (N1619, N1618, N679);
and AND3 (N1620, N1610, N33, N184);
nand NAND3 (N1621, N1615, N1508, N728);
nand NAND2 (N1622, N1560, N1360);
and AND4 (N1623, N1620, N1066, N165, N984);
and AND2 (N1624, N1613, N431);
xor XOR2 (N1625, N1607, N1012);
and AND4 (N1626, N1621, N512, N1065, N1333);
xor XOR2 (N1627, N1604, N336);
nor NOR3 (N1628, N1623, N1192, N1139);
nor NOR2 (N1629, N1628, N1429);
buf BUF1 (N1630, N1619);
not NOT1 (N1631, N1617);
not NOT1 (N1632, N1622);
or OR3 (N1633, N1625, N800, N48);
not NOT1 (N1634, N1624);
buf BUF1 (N1635, N1616);
or OR2 (N1636, N1630, N483);
nor NOR2 (N1637, N1635, N848);
or OR4 (N1638, N1633, N238, N14, N41);
xor XOR2 (N1639, N1627, N776);
nand NAND4 (N1640, N1631, N1234, N1502, N1488);
xor XOR2 (N1641, N1640, N191);
nor NOR4 (N1642, N1629, N1100, N154, N1262);
buf BUF1 (N1643, N1636);
or OR2 (N1644, N1638, N817);
buf BUF1 (N1645, N1632);
buf BUF1 (N1646, N1634);
xor XOR2 (N1647, N1643, N535);
nor NOR2 (N1648, N1639, N1432);
nand NAND4 (N1649, N1626, N1384, N1375, N1227);
buf BUF1 (N1650, N1644);
or OR2 (N1651, N1647, N1535);
xor XOR2 (N1652, N1637, N649);
nand NAND3 (N1653, N1645, N565, N1523);
not NOT1 (N1654, N1652);
or OR2 (N1655, N1653, N1077);
xor XOR2 (N1656, N1651, N1193);
xor XOR2 (N1657, N1656, N1274);
nor NOR2 (N1658, N1611, N582);
and AND4 (N1659, N1642, N1467, N1287, N161);
buf BUF1 (N1660, N1648);
and AND3 (N1661, N1659, N664, N1121);
xor XOR2 (N1662, N1655, N371);
not NOT1 (N1663, N1658);
and AND2 (N1664, N1657, N1222);
xor XOR2 (N1665, N1662, N915);
buf BUF1 (N1666, N1663);
or OR2 (N1667, N1665, N1240);
nor NOR3 (N1668, N1664, N1603, N1485);
or OR4 (N1669, N1650, N1061, N1066, N495);
nand NAND2 (N1670, N1649, N1644);
or OR3 (N1671, N1667, N1086, N244);
buf BUF1 (N1672, N1661);
xor XOR2 (N1673, N1668, N541);
and AND4 (N1674, N1673, N1315, N371, N596);
buf BUF1 (N1675, N1660);
not NOT1 (N1676, N1669);
not NOT1 (N1677, N1676);
not NOT1 (N1678, N1654);
xor XOR2 (N1679, N1641, N1160);
buf BUF1 (N1680, N1672);
buf BUF1 (N1681, N1666);
and AND3 (N1682, N1670, N459, N1340);
nand NAND4 (N1683, N1675, N899, N1325, N151);
xor XOR2 (N1684, N1680, N483);
nor NOR2 (N1685, N1678, N565);
nor NOR2 (N1686, N1681, N87);
xor XOR2 (N1687, N1685, N63);
not NOT1 (N1688, N1683);
nand NAND4 (N1689, N1682, N414, N1375, N906);
xor XOR2 (N1690, N1671, N690);
nor NOR4 (N1691, N1677, N941, N1547, N1451);
xor XOR2 (N1692, N1688, N1436);
nand NAND4 (N1693, N1686, N1175, N846, N1313);
and AND4 (N1694, N1691, N761, N1652, N61);
buf BUF1 (N1695, N1693);
and AND3 (N1696, N1692, N944, N1442);
or OR2 (N1697, N1684, N655);
or OR3 (N1698, N1694, N469, N105);
and AND3 (N1699, N1690, N1694, N450);
and AND3 (N1700, N1646, N1324, N340);
and AND2 (N1701, N1679, N740);
nor NOR4 (N1702, N1674, N742, N447, N582);
or OR4 (N1703, N1702, N1443, N879, N171);
xor XOR2 (N1704, N1695, N431);
nand NAND3 (N1705, N1701, N661, N1393);
buf BUF1 (N1706, N1696);
nand NAND3 (N1707, N1697, N1148, N253);
nand NAND2 (N1708, N1705, N377);
nor NOR2 (N1709, N1698, N534);
nand NAND4 (N1710, N1708, N1147, N87, N532);
not NOT1 (N1711, N1703);
nand NAND2 (N1712, N1706, N1423);
not NOT1 (N1713, N1709);
or OR4 (N1714, N1713, N1393, N570, N445);
or OR2 (N1715, N1710, N355);
xor XOR2 (N1716, N1700, N802);
nor NOR3 (N1717, N1711, N1531, N927);
nand NAND4 (N1718, N1704, N1213, N1561, N18);
and AND4 (N1719, N1716, N1597, N1337, N1183);
and AND4 (N1720, N1712, N1474, N363, N1524);
xor XOR2 (N1721, N1689, N281);
xor XOR2 (N1722, N1714, N578);
or OR4 (N1723, N1707, N152, N141, N1059);
and AND4 (N1724, N1687, N1464, N1604, N36);
or OR4 (N1725, N1719, N1579, N1549, N1303);
nand NAND4 (N1726, N1722, N384, N580, N1015);
nor NOR2 (N1727, N1721, N508);
or OR2 (N1728, N1724, N503);
xor XOR2 (N1729, N1726, N1170);
and AND3 (N1730, N1717, N1520, N802);
nor NOR2 (N1731, N1718, N1542);
nand NAND4 (N1732, N1729, N1219, N1420, N462);
not NOT1 (N1733, N1727);
xor XOR2 (N1734, N1730, N855);
xor XOR2 (N1735, N1715, N411);
and AND3 (N1736, N1720, N1602, N957);
or OR4 (N1737, N1723, N510, N1718, N1643);
and AND4 (N1738, N1735, N529, N252, N40);
and AND3 (N1739, N1734, N1673, N373);
not NOT1 (N1740, N1731);
or OR2 (N1741, N1738, N526);
nand NAND4 (N1742, N1740, N1535, N143, N1458);
nor NOR2 (N1743, N1732, N1502);
buf BUF1 (N1744, N1743);
or OR2 (N1745, N1744, N409);
or OR4 (N1746, N1742, N1107, N364, N449);
nor NOR3 (N1747, N1745, N340, N1273);
nor NOR3 (N1748, N1725, N753, N1381);
xor XOR2 (N1749, N1746, N896);
nand NAND2 (N1750, N1728, N1038);
buf BUF1 (N1751, N1699);
or OR3 (N1752, N1733, N1332, N1654);
nand NAND2 (N1753, N1747, N642);
buf BUF1 (N1754, N1752);
nor NOR3 (N1755, N1754, N1114, N102);
buf BUF1 (N1756, N1749);
buf BUF1 (N1757, N1739);
nor NOR3 (N1758, N1756, N332, N1382);
not NOT1 (N1759, N1757);
buf BUF1 (N1760, N1741);
buf BUF1 (N1761, N1759);
or OR2 (N1762, N1760, N1613);
xor XOR2 (N1763, N1758, N1437);
and AND4 (N1764, N1762, N1287, N1658, N1024);
nor NOR3 (N1765, N1750, N1012, N1653);
nand NAND2 (N1766, N1748, N1042);
buf BUF1 (N1767, N1751);
nand NAND3 (N1768, N1764, N672, N1153);
or OR4 (N1769, N1763, N1416, N1732, N1531);
not NOT1 (N1770, N1761);
xor XOR2 (N1771, N1736, N1544);
and AND2 (N1772, N1766, N46);
nand NAND3 (N1773, N1771, N1219, N287);
buf BUF1 (N1774, N1753);
nand NAND2 (N1775, N1769, N650);
not NOT1 (N1776, N1767);
not NOT1 (N1777, N1774);
xor XOR2 (N1778, N1776, N617);
or OR4 (N1779, N1765, N251, N1644, N924);
not NOT1 (N1780, N1737);
xor XOR2 (N1781, N1777, N1169);
nor NOR3 (N1782, N1778, N1558, N49);
not NOT1 (N1783, N1770);
xor XOR2 (N1784, N1780, N1573);
nor NOR3 (N1785, N1783, N469, N813);
not NOT1 (N1786, N1785);
or OR4 (N1787, N1755, N1166, N1424, N63);
or OR2 (N1788, N1779, N675);
buf BUF1 (N1789, N1782);
nand NAND3 (N1790, N1773, N1606, N169);
xor XOR2 (N1791, N1775, N1705);
xor XOR2 (N1792, N1788, N1005);
buf BUF1 (N1793, N1792);
nor NOR2 (N1794, N1790, N177);
nor NOR3 (N1795, N1789, N344, N331);
nor NOR4 (N1796, N1786, N449, N1064, N1237);
nor NOR2 (N1797, N1772, N1193);
nand NAND3 (N1798, N1793, N617, N1428);
buf BUF1 (N1799, N1795);
nand NAND4 (N1800, N1768, N404, N885, N356);
nor NOR2 (N1801, N1800, N1210);
buf BUF1 (N1802, N1797);
nand NAND4 (N1803, N1801, N1104, N222, N872);
and AND3 (N1804, N1787, N1414, N1275);
buf BUF1 (N1805, N1794);
nor NOR3 (N1806, N1802, N1529, N1556);
or OR4 (N1807, N1804, N55, N1170, N1222);
not NOT1 (N1808, N1791);
and AND4 (N1809, N1803, N532, N1134, N1308);
not NOT1 (N1810, N1784);
nand NAND2 (N1811, N1807, N595);
xor XOR2 (N1812, N1805, N795);
xor XOR2 (N1813, N1809, N992);
not NOT1 (N1814, N1798);
buf BUF1 (N1815, N1813);
and AND3 (N1816, N1799, N1340, N691);
nor NOR3 (N1817, N1816, N1293, N396);
and AND4 (N1818, N1815, N475, N126, N271);
and AND3 (N1819, N1810, N418, N1639);
buf BUF1 (N1820, N1811);
xor XOR2 (N1821, N1796, N1342);
or OR3 (N1822, N1820, N732, N617);
xor XOR2 (N1823, N1812, N961);
nor NOR4 (N1824, N1817, N400, N1723, N1285);
nor NOR2 (N1825, N1814, N1458);
or OR2 (N1826, N1781, N1304);
or OR4 (N1827, N1808, N1731, N938, N179);
buf BUF1 (N1828, N1818);
and AND3 (N1829, N1824, N985, N907);
or OR2 (N1830, N1821, N450);
not NOT1 (N1831, N1827);
and AND4 (N1832, N1823, N602, N435, N216);
or OR2 (N1833, N1806, N1097);
and AND4 (N1834, N1819, N1493, N1825, N1354);
and AND2 (N1835, N133, N1731);
not NOT1 (N1836, N1826);
not NOT1 (N1837, N1831);
xor XOR2 (N1838, N1828, N1556);
xor XOR2 (N1839, N1830, N127);
not NOT1 (N1840, N1836);
xor XOR2 (N1841, N1839, N1068);
and AND4 (N1842, N1837, N1760, N896, N874);
xor XOR2 (N1843, N1842, N1456);
not NOT1 (N1844, N1835);
nand NAND2 (N1845, N1833, N702);
not NOT1 (N1846, N1840);
nand NAND2 (N1847, N1832, N1109);
xor XOR2 (N1848, N1847, N1361);
not NOT1 (N1849, N1841);
nor NOR2 (N1850, N1846, N205);
nor NOR2 (N1851, N1829, N904);
nand NAND4 (N1852, N1848, N511, N1093, N1677);
nand NAND4 (N1853, N1845, N158, N1462, N498);
buf BUF1 (N1854, N1822);
and AND3 (N1855, N1853, N1360, N716);
xor XOR2 (N1856, N1838, N1272);
not NOT1 (N1857, N1834);
and AND2 (N1858, N1849, N409);
or OR3 (N1859, N1851, N1683, N831);
buf BUF1 (N1860, N1850);
and AND3 (N1861, N1844, N934, N169);
buf BUF1 (N1862, N1852);
buf BUF1 (N1863, N1856);
not NOT1 (N1864, N1861);
and AND2 (N1865, N1855, N581);
and AND4 (N1866, N1864, N1037, N1461, N1363);
nand NAND2 (N1867, N1854, N1211);
nor NOR3 (N1868, N1863, N412, N104);
or OR3 (N1869, N1866, N1187, N1011);
nand NAND2 (N1870, N1857, N323);
nor NOR2 (N1871, N1859, N1435);
or OR3 (N1872, N1860, N872, N652);
and AND2 (N1873, N1858, N1520);
nand NAND4 (N1874, N1869, N255, N237, N818);
and AND2 (N1875, N1870, N745);
buf BUF1 (N1876, N1843);
nand NAND3 (N1877, N1868, N693, N1822);
not NOT1 (N1878, N1877);
buf BUF1 (N1879, N1867);
or OR2 (N1880, N1862, N687);
buf BUF1 (N1881, N1871);
or OR4 (N1882, N1873, N1070, N65, N394);
not NOT1 (N1883, N1875);
not NOT1 (N1884, N1872);
buf BUF1 (N1885, N1879);
nor NOR4 (N1886, N1876, N1885, N1363, N405);
or OR3 (N1887, N1086, N127, N674);
buf BUF1 (N1888, N1884);
buf BUF1 (N1889, N1882);
or OR2 (N1890, N1878, N769);
xor XOR2 (N1891, N1890, N947);
nand NAND2 (N1892, N1881, N1451);
or OR3 (N1893, N1880, N594, N1510);
or OR2 (N1894, N1888, N598);
not NOT1 (N1895, N1886);
not NOT1 (N1896, N1895);
or OR4 (N1897, N1865, N1207, N1254, N883);
xor XOR2 (N1898, N1892, N1690);
or OR3 (N1899, N1889, N1403, N945);
nor NOR2 (N1900, N1898, N101);
or OR3 (N1901, N1893, N504, N1533);
xor XOR2 (N1902, N1883, N1436);
and AND4 (N1903, N1901, N891, N314, N1433);
or OR3 (N1904, N1894, N753, N90);
nand NAND2 (N1905, N1900, N744);
xor XOR2 (N1906, N1902, N1738);
and AND3 (N1907, N1891, N1902, N766);
not NOT1 (N1908, N1897);
buf BUF1 (N1909, N1896);
nand NAND2 (N1910, N1909, N343);
nor NOR2 (N1911, N1904, N1317);
and AND3 (N1912, N1908, N1678, N967);
not NOT1 (N1913, N1887);
or OR4 (N1914, N1913, N595, N1803, N1146);
xor XOR2 (N1915, N1906, N1069);
nand NAND2 (N1916, N1914, N909);
not NOT1 (N1917, N1874);
or OR4 (N1918, N1915, N399, N1751, N912);
xor XOR2 (N1919, N1910, N1521);
xor XOR2 (N1920, N1905, N459);
not NOT1 (N1921, N1917);
nand NAND2 (N1922, N1912, N65);
or OR4 (N1923, N1916, N393, N701, N1201);
buf BUF1 (N1924, N1922);
and AND3 (N1925, N1899, N293, N1523);
not NOT1 (N1926, N1924);
buf BUF1 (N1927, N1921);
or OR4 (N1928, N1918, N681, N1195, N1211);
not NOT1 (N1929, N1926);
xor XOR2 (N1930, N1925, N418);
nor NOR3 (N1931, N1920, N137, N1507);
xor XOR2 (N1932, N1911, N862);
or OR2 (N1933, N1928, N127);
or OR4 (N1934, N1930, N907, N414, N212);
not NOT1 (N1935, N1929);
not NOT1 (N1936, N1934);
xor XOR2 (N1937, N1931, N1220);
nor NOR2 (N1938, N1936, N1167);
nor NOR3 (N1939, N1927, N948, N56);
buf BUF1 (N1940, N1903);
not NOT1 (N1941, N1935);
not NOT1 (N1942, N1923);
nor NOR3 (N1943, N1932, N1638, N858);
nor NOR4 (N1944, N1938, N1238, N1218, N1244);
xor XOR2 (N1945, N1907, N1200);
and AND4 (N1946, N1941, N1897, N1735, N1411);
xor XOR2 (N1947, N1933, N1249);
nand NAND3 (N1948, N1919, N1628, N1299);
buf BUF1 (N1949, N1947);
and AND2 (N1950, N1943, N961);
or OR2 (N1951, N1937, N739);
nor NOR3 (N1952, N1944, N177, N1039);
or OR3 (N1953, N1950, N1695, N990);
nand NAND4 (N1954, N1949, N340, N1357, N693);
xor XOR2 (N1955, N1948, N37);
nand NAND4 (N1956, N1945, N669, N1495, N1634);
buf BUF1 (N1957, N1946);
nand NAND4 (N1958, N1952, N48, N1908, N526);
nand NAND4 (N1959, N1939, N1678, N787, N1490);
nor NOR3 (N1960, N1953, N1957, N926);
not NOT1 (N1961, N404);
buf BUF1 (N1962, N1960);
nand NAND3 (N1963, N1961, N426, N1472);
xor XOR2 (N1964, N1940, N71);
nor NOR4 (N1965, N1951, N742, N509, N1099);
and AND2 (N1966, N1963, N1532);
and AND3 (N1967, N1965, N1506, N958);
nor NOR4 (N1968, N1964, N751, N1612, N1121);
buf BUF1 (N1969, N1968);
buf BUF1 (N1970, N1966);
xor XOR2 (N1971, N1956, N526);
nor NOR2 (N1972, N1959, N712);
not NOT1 (N1973, N1954);
xor XOR2 (N1974, N1955, N790);
nand NAND3 (N1975, N1971, N177, N204);
buf BUF1 (N1976, N1962);
buf BUF1 (N1977, N1942);
buf BUF1 (N1978, N1969);
buf BUF1 (N1979, N1975);
nor NOR4 (N1980, N1972, N1398, N1641, N1820);
or OR2 (N1981, N1977, N1713);
xor XOR2 (N1982, N1978, N705);
not NOT1 (N1983, N1967);
and AND4 (N1984, N1970, N880, N81, N857);
nand NAND2 (N1985, N1976, N1055);
not NOT1 (N1986, N1981);
nor NOR3 (N1987, N1983, N1676, N855);
and AND3 (N1988, N1980, N1200, N271);
nand NAND4 (N1989, N1958, N1891, N215, N1468);
or OR2 (N1990, N1984, N1956);
and AND2 (N1991, N1982, N1816);
or OR2 (N1992, N1986, N1284);
or OR3 (N1993, N1988, N1457, N678);
buf BUF1 (N1994, N1992);
and AND3 (N1995, N1987, N405, N1953);
nor NOR2 (N1996, N1994, N75);
xor XOR2 (N1997, N1974, N136);
and AND4 (N1998, N1991, N913, N1475, N1796);
or OR2 (N1999, N1979, N59);
not NOT1 (N2000, N1996);
nand NAND3 (N2001, N1997, N352, N857);
nor NOR4 (N2002, N1999, N174, N1255, N634);
buf BUF1 (N2003, N2001);
or OR2 (N2004, N1973, N1830);
xor XOR2 (N2005, N1989, N1603);
nor NOR4 (N2006, N1995, N1038, N790, N1345);
or OR2 (N2007, N2002, N1423);
nand NAND4 (N2008, N2004, N1561, N692, N439);
xor XOR2 (N2009, N2007, N1967);
and AND4 (N2010, N2003, N1315, N1410, N1454);
nor NOR3 (N2011, N2000, N502, N769);
nand NAND4 (N2012, N1990, N1465, N474, N1660);
or OR2 (N2013, N2009, N286);
xor XOR2 (N2014, N2005, N1656);
or OR4 (N2015, N2010, N1550, N1690, N668);
buf BUF1 (N2016, N2008);
endmodule