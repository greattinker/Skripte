// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;

output N1615,N1618,N1620,N1612,N1621,N1619,N1597,N1623,N1622,N1624;

xor XOR2 (N25, N13, N20);
and AND4 (N26, N22, N3, N9, N17);
or OR2 (N27, N2, N14);
xor XOR2 (N28, N6, N27);
not NOT1 (N29, N11);
nor NOR3 (N30, N22, N15, N18);
nor NOR2 (N31, N23, N17);
not NOT1 (N32, N12);
or OR3 (N33, N29, N4, N14);
xor XOR2 (N34, N17, N20);
and AND4 (N35, N1, N12, N19, N25);
and AND3 (N36, N29, N32, N18);
and AND4 (N37, N28, N13, N31, N25);
nand NAND2 (N38, N28, N6);
and AND4 (N39, N14, N16, N4, N19);
xor XOR2 (N40, N16, N20);
or OR4 (N41, N33, N7, N18, N40);
xor XOR2 (N42, N17, N7);
nor NOR4 (N43, N36, N20, N21, N19);
nor NOR2 (N44, N34, N18);
buf BUF1 (N45, N43);
xor XOR2 (N46, N39, N38);
buf BUF1 (N47, N7);
nand NAND2 (N48, N47, N16);
and AND2 (N49, N42, N19);
and AND4 (N50, N35, N48, N2, N27);
not NOT1 (N51, N34);
xor XOR2 (N52, N44, N31);
nand NAND3 (N53, N46, N52, N39);
buf BUF1 (N54, N34);
and AND4 (N55, N45, N47, N17, N41);
not NOT1 (N56, N14);
nor NOR2 (N57, N54, N38);
or OR3 (N58, N56, N33, N3);
not NOT1 (N59, N51);
buf BUF1 (N60, N53);
nand NAND2 (N61, N55, N34);
or OR4 (N62, N26, N35, N36, N19);
not NOT1 (N63, N60);
and AND2 (N64, N62, N1);
and AND3 (N65, N30, N24, N41);
and AND3 (N66, N58, N37, N51);
and AND3 (N67, N23, N9, N35);
xor XOR2 (N68, N67, N36);
xor XOR2 (N69, N50, N9);
xor XOR2 (N70, N65, N9);
not NOT1 (N71, N68);
xor XOR2 (N72, N70, N22);
and AND3 (N73, N64, N23, N61);
nand NAND3 (N74, N8, N47, N17);
not NOT1 (N75, N49);
and AND3 (N76, N74, N61, N54);
nand NAND3 (N77, N66, N49, N71);
nor NOR2 (N78, N1, N13);
nand NAND3 (N79, N76, N71, N60);
not NOT1 (N80, N72);
and AND2 (N81, N69, N59);
nor NOR4 (N82, N36, N81, N79, N76);
nor NOR2 (N83, N17, N48);
xor XOR2 (N84, N73, N27);
buf BUF1 (N85, N54);
or OR2 (N86, N63, N4);
nand NAND3 (N87, N86, N78, N59);
not NOT1 (N88, N66);
buf BUF1 (N89, N84);
nand NAND3 (N90, N88, N89, N23);
and AND4 (N91, N23, N28, N51, N42);
xor XOR2 (N92, N90, N12);
and AND2 (N93, N92, N41);
xor XOR2 (N94, N91, N34);
xor XOR2 (N95, N85, N76);
buf BUF1 (N96, N83);
not NOT1 (N97, N93);
buf BUF1 (N98, N95);
or OR2 (N99, N57, N35);
or OR2 (N100, N94, N60);
not NOT1 (N101, N98);
xor XOR2 (N102, N80, N75);
buf BUF1 (N103, N13);
or OR3 (N104, N87, N82, N46);
buf BUF1 (N105, N75);
xor XOR2 (N106, N104, N52);
xor XOR2 (N107, N101, N46);
nor NOR2 (N108, N96, N74);
nand NAND2 (N109, N100, N87);
not NOT1 (N110, N107);
nand NAND4 (N111, N97, N6, N91, N101);
nor NOR4 (N112, N111, N81, N77, N73);
or OR4 (N113, N45, N79, N32, N89);
xor XOR2 (N114, N105, N3);
nor NOR4 (N115, N110, N2, N41, N111);
nor NOR3 (N116, N113, N41, N104);
not NOT1 (N117, N112);
or OR3 (N118, N116, N108, N80);
or OR4 (N119, N44, N5, N113, N2);
nand NAND3 (N120, N117, N14, N1);
not NOT1 (N121, N115);
not NOT1 (N122, N102);
buf BUF1 (N123, N119);
buf BUF1 (N124, N109);
or OR4 (N125, N123, N6, N58, N47);
not NOT1 (N126, N106);
nand NAND2 (N127, N125, N25);
nand NAND2 (N128, N126, N3);
xor XOR2 (N129, N127, N80);
not NOT1 (N130, N124);
or OR4 (N131, N130, N120, N76, N76);
nor NOR3 (N132, N125, N98, N96);
not NOT1 (N133, N114);
and AND2 (N134, N121, N59);
or OR4 (N135, N131, N36, N59, N91);
and AND3 (N136, N132, N12, N65);
nand NAND4 (N137, N118, N80, N111, N10);
nand NAND2 (N138, N103, N72);
nor NOR4 (N139, N122, N138, N42, N120);
nor NOR4 (N140, N135, N98, N8, N44);
nand NAND2 (N141, N6, N63);
and AND3 (N142, N141, N15, N81);
or OR3 (N143, N142, N22, N111);
nor NOR4 (N144, N134, N139, N55, N101);
nand NAND2 (N145, N82, N84);
not NOT1 (N146, N144);
nor NOR4 (N147, N128, N131, N136, N24);
buf BUF1 (N148, N124);
or OR4 (N149, N145, N33, N71, N80);
nor NOR3 (N150, N137, N78, N78);
not NOT1 (N151, N148);
and AND3 (N152, N151, N44, N131);
xor XOR2 (N153, N143, N115);
and AND4 (N154, N150, N57, N84, N64);
and AND2 (N155, N152, N3);
buf BUF1 (N156, N149);
nand NAND4 (N157, N146, N92, N132, N57);
xor XOR2 (N158, N133, N41);
or OR4 (N159, N155, N29, N5, N24);
xor XOR2 (N160, N158, N53);
or OR2 (N161, N154, N20);
or OR2 (N162, N99, N109);
nand NAND3 (N163, N140, N30, N122);
nand NAND2 (N164, N161, N76);
xor XOR2 (N165, N147, N5);
nand NAND4 (N166, N129, N56, N141, N9);
xor XOR2 (N167, N165, N105);
nor NOR2 (N168, N159, N61);
not NOT1 (N169, N164);
buf BUF1 (N170, N153);
nor NOR2 (N171, N166, N105);
nand NAND3 (N172, N171, N17, N45);
or OR4 (N173, N160, N30, N135, N28);
nand NAND4 (N174, N168, N169, N39, N59);
and AND3 (N175, N46, N159, N105);
nand NAND2 (N176, N167, N172);
or OR4 (N177, N175, N117, N71, N158);
buf BUF1 (N178, N171);
nor NOR3 (N179, N163, N107, N90);
or OR2 (N180, N179, N142);
not NOT1 (N181, N156);
nand NAND3 (N182, N177, N9, N59);
and AND3 (N183, N173, N9, N84);
nand NAND4 (N184, N170, N47, N78, N172);
xor XOR2 (N185, N184, N60);
or OR2 (N186, N183, N61);
and AND3 (N187, N182, N96, N97);
or OR4 (N188, N162, N156, N106, N12);
not NOT1 (N189, N174);
and AND2 (N190, N185, N135);
not NOT1 (N191, N187);
and AND2 (N192, N186, N36);
or OR3 (N193, N180, N130, N148);
xor XOR2 (N194, N181, N17);
not NOT1 (N195, N157);
not NOT1 (N196, N178);
buf BUF1 (N197, N190);
nor NOR2 (N198, N189, N194);
and AND4 (N199, N77, N65, N63, N128);
xor XOR2 (N200, N198, N84);
nand NAND3 (N201, N188, N6, N80);
xor XOR2 (N202, N176, N107);
xor XOR2 (N203, N193, N184);
or OR3 (N204, N199, N119, N87);
nand NAND4 (N205, N200, N171, N1, N48);
xor XOR2 (N206, N201, N61);
nor NOR4 (N207, N203, N58, N136, N108);
xor XOR2 (N208, N204, N54);
nand NAND3 (N209, N192, N16, N40);
nand NAND4 (N210, N191, N11, N168, N77);
nand NAND4 (N211, N206, N55, N190, N20);
xor XOR2 (N212, N195, N30);
and AND3 (N213, N196, N153, N108);
and AND2 (N214, N207, N132);
or OR3 (N215, N197, N99, N79);
not NOT1 (N216, N202);
and AND3 (N217, N208, N160, N85);
not NOT1 (N218, N205);
not NOT1 (N219, N214);
and AND3 (N220, N213, N95, N166);
buf BUF1 (N221, N211);
not NOT1 (N222, N210);
nor NOR3 (N223, N209, N100, N209);
buf BUF1 (N224, N219);
or OR3 (N225, N221, N203, N95);
nor NOR3 (N226, N217, N153, N125);
and AND2 (N227, N218, N192);
buf BUF1 (N228, N215);
buf BUF1 (N229, N216);
xor XOR2 (N230, N223, N170);
or OR2 (N231, N212, N16);
xor XOR2 (N232, N222, N103);
xor XOR2 (N233, N229, N202);
nand NAND4 (N234, N227, N106, N36, N155);
xor XOR2 (N235, N226, N118);
or OR4 (N236, N235, N29, N14, N163);
xor XOR2 (N237, N231, N78);
xor XOR2 (N238, N232, N21);
xor XOR2 (N239, N224, N39);
not NOT1 (N240, N230);
xor XOR2 (N241, N234, N83);
nor NOR4 (N242, N233, N30, N202, N181);
and AND3 (N243, N220, N36, N242);
nor NOR3 (N244, N223, N20, N232);
buf BUF1 (N245, N241);
nand NAND2 (N246, N240, N99);
not NOT1 (N247, N237);
xor XOR2 (N248, N246, N35);
or OR4 (N249, N245, N52, N206, N234);
xor XOR2 (N250, N225, N61);
xor XOR2 (N251, N247, N208);
not NOT1 (N252, N236);
not NOT1 (N253, N248);
and AND3 (N254, N250, N228, N100);
xor XOR2 (N255, N190, N82);
buf BUF1 (N256, N254);
nand NAND2 (N257, N249, N24);
not NOT1 (N258, N239);
not NOT1 (N259, N238);
or OR2 (N260, N256, N150);
nand NAND2 (N261, N257, N142);
nand NAND2 (N262, N255, N108);
buf BUF1 (N263, N244);
nand NAND2 (N264, N243, N20);
buf BUF1 (N265, N263);
buf BUF1 (N266, N264);
nand NAND3 (N267, N258, N260, N194);
or OR4 (N268, N122, N45, N130, N161);
or OR4 (N269, N262, N31, N250, N160);
buf BUF1 (N270, N261);
xor XOR2 (N271, N267, N140);
or OR3 (N272, N251, N29, N38);
xor XOR2 (N273, N268, N160);
buf BUF1 (N274, N259);
and AND3 (N275, N265, N57, N274);
or OR3 (N276, N235, N87, N105);
and AND3 (N277, N270, N249, N221);
not NOT1 (N278, N277);
buf BUF1 (N279, N269);
or OR2 (N280, N271, N31);
nand NAND4 (N281, N280, N54, N141, N117);
xor XOR2 (N282, N279, N91);
or OR2 (N283, N273, N99);
buf BUF1 (N284, N272);
not NOT1 (N285, N282);
buf BUF1 (N286, N266);
or OR2 (N287, N286, N81);
not NOT1 (N288, N283);
buf BUF1 (N289, N252);
buf BUF1 (N290, N276);
buf BUF1 (N291, N253);
nand NAND3 (N292, N287, N85, N35);
xor XOR2 (N293, N278, N123);
nand NAND3 (N294, N290, N219, N132);
or OR2 (N295, N291, N123);
nor NOR3 (N296, N284, N2, N55);
nor NOR3 (N297, N275, N115, N220);
and AND3 (N298, N297, N55, N282);
buf BUF1 (N299, N281);
buf BUF1 (N300, N292);
nor NOR4 (N301, N296, N262, N192, N62);
buf BUF1 (N302, N294);
or OR3 (N303, N300, N139, N133);
nor NOR2 (N304, N295, N85);
nor NOR3 (N305, N285, N62, N114);
and AND4 (N306, N304, N57, N223, N156);
not NOT1 (N307, N298);
nand NAND4 (N308, N288, N257, N260, N33);
and AND3 (N309, N306, N132, N169);
nor NOR4 (N310, N302, N286, N134, N121);
not NOT1 (N311, N308);
xor XOR2 (N312, N307, N182);
nand NAND3 (N313, N299, N84, N132);
xor XOR2 (N314, N305, N134);
xor XOR2 (N315, N312, N34);
buf BUF1 (N316, N309);
and AND3 (N317, N314, N146, N33);
buf BUF1 (N318, N315);
nor NOR3 (N319, N317, N257, N269);
buf BUF1 (N320, N310);
buf BUF1 (N321, N313);
not NOT1 (N322, N311);
or OR2 (N323, N318, N147);
and AND2 (N324, N293, N153);
xor XOR2 (N325, N322, N7);
not NOT1 (N326, N316);
nand NAND3 (N327, N301, N176, N265);
nand NAND4 (N328, N319, N127, N229, N244);
nand NAND2 (N329, N328, N139);
and AND4 (N330, N320, N194, N4, N290);
nor NOR4 (N331, N324, N151, N232, N9);
nand NAND4 (N332, N289, N169, N62, N55);
or OR4 (N333, N321, N65, N203, N170);
not NOT1 (N334, N329);
not NOT1 (N335, N334);
and AND4 (N336, N330, N23, N194, N41);
or OR2 (N337, N331, N41);
or OR4 (N338, N303, N126, N223, N68);
buf BUF1 (N339, N332);
or OR2 (N340, N336, N276);
nor NOR2 (N341, N326, N26);
not NOT1 (N342, N333);
or OR3 (N343, N341, N144, N225);
and AND4 (N344, N338, N43, N26, N261);
nand NAND3 (N345, N342, N343, N309);
xor XOR2 (N346, N265, N341);
and AND2 (N347, N339, N276);
nand NAND2 (N348, N346, N139);
or OR2 (N349, N327, N184);
not NOT1 (N350, N345);
or OR3 (N351, N323, N331, N4);
nor NOR4 (N352, N344, N103, N3, N304);
buf BUF1 (N353, N352);
nor NOR3 (N354, N340, N185, N146);
and AND3 (N355, N337, N2, N86);
and AND3 (N356, N350, N254, N235);
nand NAND4 (N357, N349, N313, N349, N293);
nor NOR3 (N358, N351, N104, N196);
or OR2 (N359, N358, N93);
or OR2 (N360, N347, N32);
nand NAND2 (N361, N325, N279);
buf BUF1 (N362, N360);
or OR4 (N363, N335, N233, N264, N95);
nand NAND3 (N364, N363, N188, N98);
and AND3 (N365, N357, N1, N256);
nor NOR2 (N366, N365, N54);
not NOT1 (N367, N359);
and AND4 (N368, N367, N96, N344, N334);
and AND4 (N369, N364, N343, N208, N345);
xor XOR2 (N370, N362, N209);
nor NOR2 (N371, N355, N326);
and AND4 (N372, N371, N9, N258, N20);
and AND3 (N373, N353, N70, N359);
and AND2 (N374, N354, N251);
not NOT1 (N375, N374);
xor XOR2 (N376, N372, N11);
xor XOR2 (N377, N376, N42);
nand NAND3 (N378, N369, N227, N22);
nor NOR2 (N379, N377, N36);
not NOT1 (N380, N348);
nand NAND3 (N381, N370, N162, N120);
nand NAND3 (N382, N379, N152, N217);
nand NAND2 (N383, N381, N1);
or OR3 (N384, N373, N104, N100);
buf BUF1 (N385, N366);
nand NAND3 (N386, N378, N40, N254);
nor NOR2 (N387, N361, N299);
buf BUF1 (N388, N356);
buf BUF1 (N389, N384);
and AND4 (N390, N383, N57, N249, N374);
not NOT1 (N391, N388);
xor XOR2 (N392, N382, N88);
nor NOR4 (N393, N389, N194, N75, N237);
or OR4 (N394, N380, N179, N120, N352);
xor XOR2 (N395, N391, N388);
not NOT1 (N396, N393);
buf BUF1 (N397, N375);
nor NOR4 (N398, N387, N96, N56, N214);
or OR3 (N399, N386, N15, N132);
or OR4 (N400, N390, N91, N250, N240);
and AND2 (N401, N398, N358);
or OR4 (N402, N395, N203, N35, N27);
nor NOR2 (N403, N401, N139);
or OR2 (N404, N399, N162);
nand NAND4 (N405, N397, N351, N107, N339);
and AND3 (N406, N403, N335, N238);
not NOT1 (N407, N400);
nand NAND3 (N408, N407, N1, N172);
buf BUF1 (N409, N404);
or OR3 (N410, N368, N65, N66);
and AND3 (N411, N392, N23, N206);
not NOT1 (N412, N405);
nor NOR2 (N413, N409, N103);
buf BUF1 (N414, N402);
xor XOR2 (N415, N413, N185);
nand NAND4 (N416, N406, N369, N338, N201);
nor NOR3 (N417, N416, N274, N166);
xor XOR2 (N418, N414, N413);
not NOT1 (N419, N408);
not NOT1 (N420, N411);
or OR4 (N421, N417, N147, N301, N203);
nor NOR3 (N422, N421, N258, N183);
and AND4 (N423, N385, N118, N67, N296);
not NOT1 (N424, N412);
nor NOR4 (N425, N419, N75, N134, N361);
xor XOR2 (N426, N415, N45);
buf BUF1 (N427, N396);
and AND2 (N428, N420, N391);
buf BUF1 (N429, N426);
not NOT1 (N430, N422);
nor NOR4 (N431, N427, N169, N304, N229);
and AND3 (N432, N418, N279, N198);
and AND3 (N433, N410, N23, N215);
nand NAND4 (N434, N423, N312, N134, N236);
and AND2 (N435, N394, N196);
not NOT1 (N436, N434);
nand NAND2 (N437, N436, N220);
buf BUF1 (N438, N435);
or OR4 (N439, N437, N342, N121, N43);
and AND3 (N440, N424, N161, N353);
and AND4 (N441, N438, N65, N396, N341);
not NOT1 (N442, N430);
nor NOR4 (N443, N431, N49, N332, N144);
nor NOR3 (N444, N425, N410, N260);
xor XOR2 (N445, N439, N227);
nand NAND2 (N446, N428, N250);
xor XOR2 (N447, N445, N90);
or OR3 (N448, N444, N366, N352);
not NOT1 (N449, N448);
not NOT1 (N450, N440);
and AND3 (N451, N433, N282, N201);
nor NOR2 (N452, N449, N260);
nor NOR2 (N453, N442, N103);
nand NAND4 (N454, N452, N286, N368, N188);
xor XOR2 (N455, N454, N242);
and AND4 (N456, N446, N390, N38, N77);
not NOT1 (N457, N450);
xor XOR2 (N458, N456, N49);
nand NAND3 (N459, N455, N348, N254);
nor NOR3 (N460, N459, N235, N288);
not NOT1 (N461, N429);
buf BUF1 (N462, N443);
xor XOR2 (N463, N458, N12);
nand NAND2 (N464, N453, N143);
not NOT1 (N465, N464);
not NOT1 (N466, N441);
nor NOR2 (N467, N466, N4);
xor XOR2 (N468, N447, N264);
or OR4 (N469, N457, N269, N64, N269);
or OR3 (N470, N468, N398, N100);
or OR4 (N471, N470, N87, N387, N365);
xor XOR2 (N472, N467, N443);
and AND3 (N473, N463, N102, N224);
or OR2 (N474, N462, N374);
xor XOR2 (N475, N461, N70);
buf BUF1 (N476, N469);
buf BUF1 (N477, N472);
nor NOR3 (N478, N475, N251, N255);
and AND3 (N479, N478, N137, N456);
xor XOR2 (N480, N460, N70);
and AND2 (N481, N473, N257);
nand NAND4 (N482, N476, N384, N102, N432);
xor XOR2 (N483, N70, N237);
or OR3 (N484, N451, N88, N449);
and AND2 (N485, N482, N125);
xor XOR2 (N486, N480, N36);
and AND3 (N487, N477, N53, N460);
and AND2 (N488, N465, N318);
or OR4 (N489, N486, N456, N221, N29);
and AND4 (N490, N483, N317, N166, N257);
or OR3 (N491, N479, N193, N357);
xor XOR2 (N492, N474, N227);
and AND4 (N493, N490, N113, N230, N322);
and AND2 (N494, N485, N239);
and AND4 (N495, N484, N248, N432, N271);
buf BUF1 (N496, N492);
buf BUF1 (N497, N494);
not NOT1 (N498, N481);
or OR2 (N499, N488, N288);
xor XOR2 (N500, N487, N431);
or OR3 (N501, N489, N449, N100);
nand NAND3 (N502, N501, N202, N315);
not NOT1 (N503, N498);
nand NAND3 (N504, N496, N312, N144);
and AND4 (N505, N502, N481, N37, N154);
and AND3 (N506, N499, N217, N353);
not NOT1 (N507, N491);
not NOT1 (N508, N495);
buf BUF1 (N509, N497);
xor XOR2 (N510, N505, N392);
not NOT1 (N511, N510);
nand NAND4 (N512, N471, N19, N501, N211);
nand NAND4 (N513, N512, N433, N166, N444);
or OR4 (N514, N513, N69, N119, N453);
and AND4 (N515, N511, N478, N310, N210);
or OR4 (N516, N508, N454, N432, N61);
and AND2 (N517, N506, N166);
nor NOR2 (N518, N509, N78);
xor XOR2 (N519, N516, N283);
buf BUF1 (N520, N518);
buf BUF1 (N521, N515);
xor XOR2 (N522, N520, N509);
or OR4 (N523, N519, N500, N306, N1);
buf BUF1 (N524, N391);
not NOT1 (N525, N524);
not NOT1 (N526, N507);
not NOT1 (N527, N517);
not NOT1 (N528, N493);
nand NAND4 (N529, N514, N171, N208, N49);
buf BUF1 (N530, N523);
or OR4 (N531, N503, N30, N368, N101);
and AND3 (N532, N531, N115, N351);
xor XOR2 (N533, N521, N183);
or OR3 (N534, N526, N1, N342);
buf BUF1 (N535, N534);
buf BUF1 (N536, N535);
nand NAND3 (N537, N532, N150, N266);
xor XOR2 (N538, N527, N220);
buf BUF1 (N539, N528);
or OR4 (N540, N530, N100, N287, N391);
or OR3 (N541, N539, N526, N347);
and AND2 (N542, N525, N320);
nor NOR4 (N543, N542, N297, N46, N58);
and AND2 (N544, N537, N263);
nor NOR2 (N545, N544, N485);
nand NAND4 (N546, N541, N124, N148, N478);
and AND4 (N547, N546, N473, N316, N114);
nor NOR2 (N548, N533, N285);
xor XOR2 (N549, N536, N46);
buf BUF1 (N550, N540);
not NOT1 (N551, N547);
buf BUF1 (N552, N551);
buf BUF1 (N553, N538);
or OR4 (N554, N552, N485, N95, N192);
xor XOR2 (N555, N554, N154);
not NOT1 (N556, N543);
not NOT1 (N557, N504);
not NOT1 (N558, N550);
and AND4 (N559, N557, N288, N341, N338);
nor NOR2 (N560, N558, N548);
or OR2 (N561, N143, N363);
nand NAND3 (N562, N545, N403, N303);
buf BUF1 (N563, N561);
not NOT1 (N564, N549);
nand NAND2 (N565, N529, N111);
buf BUF1 (N566, N562);
buf BUF1 (N567, N556);
buf BUF1 (N568, N565);
xor XOR2 (N569, N553, N568);
or OR4 (N570, N232, N250, N164, N158);
xor XOR2 (N571, N563, N336);
buf BUF1 (N572, N559);
buf BUF1 (N573, N566);
xor XOR2 (N574, N555, N142);
nor NOR2 (N575, N569, N437);
nor NOR2 (N576, N575, N344);
or OR4 (N577, N573, N61, N271, N542);
or OR3 (N578, N577, N15, N345);
nor NOR3 (N579, N567, N433, N176);
not NOT1 (N580, N578);
or OR3 (N581, N579, N26, N361);
or OR4 (N582, N570, N473, N290, N80);
nand NAND3 (N583, N522, N569, N133);
nand NAND4 (N584, N574, N291, N218, N506);
xor XOR2 (N585, N571, N96);
nand NAND2 (N586, N576, N133);
nor NOR3 (N587, N580, N428, N517);
buf BUF1 (N588, N586);
or OR4 (N589, N588, N363, N289, N384);
not NOT1 (N590, N589);
and AND2 (N591, N581, N73);
nor NOR4 (N592, N572, N236, N260, N111);
nand NAND3 (N593, N591, N121, N482);
buf BUF1 (N594, N564);
nor NOR2 (N595, N593, N184);
and AND3 (N596, N587, N84, N363);
and AND2 (N597, N594, N536);
nand NAND2 (N598, N590, N49);
buf BUF1 (N599, N560);
or OR3 (N600, N598, N276, N508);
xor XOR2 (N601, N583, N479);
or OR2 (N602, N596, N387);
nand NAND2 (N603, N599, N464);
and AND4 (N604, N585, N535, N420, N63);
buf BUF1 (N605, N592);
nor NOR3 (N606, N595, N138, N516);
nor NOR3 (N607, N605, N239, N551);
xor XOR2 (N608, N600, N58);
nor NOR3 (N609, N597, N134, N134);
nor NOR3 (N610, N604, N528, N499);
buf BUF1 (N611, N584);
and AND3 (N612, N611, N389, N118);
buf BUF1 (N613, N608);
or OR4 (N614, N601, N319, N494, N260);
and AND4 (N615, N609, N529, N70, N530);
xor XOR2 (N616, N615, N571);
buf BUF1 (N617, N614);
nand NAND4 (N618, N603, N367, N143, N543);
xor XOR2 (N619, N618, N106);
buf BUF1 (N620, N606);
nand NAND2 (N621, N610, N89);
not NOT1 (N622, N607);
not NOT1 (N623, N622);
buf BUF1 (N624, N619);
not NOT1 (N625, N602);
and AND4 (N626, N623, N9, N241, N486);
xor XOR2 (N627, N612, N320);
nand NAND4 (N628, N620, N344, N423, N227);
buf BUF1 (N629, N625);
buf BUF1 (N630, N582);
xor XOR2 (N631, N621, N44);
not NOT1 (N632, N624);
not NOT1 (N633, N616);
or OR3 (N634, N626, N555, N356);
xor XOR2 (N635, N627, N445);
not NOT1 (N636, N617);
buf BUF1 (N637, N632);
buf BUF1 (N638, N613);
nand NAND2 (N639, N635, N34);
buf BUF1 (N640, N629);
nor NOR2 (N641, N628, N28);
or OR3 (N642, N634, N17, N636);
not NOT1 (N643, N398);
xor XOR2 (N644, N641, N394);
xor XOR2 (N645, N640, N471);
buf BUF1 (N646, N644);
not NOT1 (N647, N643);
and AND2 (N648, N647, N213);
xor XOR2 (N649, N633, N175);
nand NAND2 (N650, N638, N347);
nor NOR2 (N651, N631, N646);
nor NOR4 (N652, N464, N617, N571, N288);
nor NOR2 (N653, N637, N362);
not NOT1 (N654, N630);
nand NAND3 (N655, N648, N429, N117);
and AND4 (N656, N642, N630, N246, N165);
not NOT1 (N657, N654);
nand NAND2 (N658, N652, N252);
or OR4 (N659, N657, N141, N478, N512);
and AND3 (N660, N651, N373, N396);
xor XOR2 (N661, N658, N508);
not NOT1 (N662, N639);
and AND2 (N663, N656, N233);
or OR4 (N664, N650, N146, N276, N486);
nand NAND3 (N665, N663, N596, N118);
xor XOR2 (N666, N655, N146);
buf BUF1 (N667, N664);
and AND4 (N668, N653, N13, N186, N282);
not NOT1 (N669, N661);
buf BUF1 (N670, N659);
and AND2 (N671, N649, N83);
buf BUF1 (N672, N667);
xor XOR2 (N673, N668, N18);
nand NAND3 (N674, N660, N654, N221);
not NOT1 (N675, N666);
not NOT1 (N676, N662);
xor XOR2 (N677, N675, N429);
nor NOR3 (N678, N669, N212, N367);
and AND2 (N679, N670, N482);
nor NOR3 (N680, N671, N616, N154);
nand NAND2 (N681, N677, N647);
or OR4 (N682, N673, N116, N180, N465);
and AND3 (N683, N679, N29, N590);
not NOT1 (N684, N676);
xor XOR2 (N685, N682, N546);
nand NAND4 (N686, N645, N243, N579, N211);
not NOT1 (N687, N678);
and AND2 (N688, N672, N598);
buf BUF1 (N689, N683);
xor XOR2 (N690, N680, N91);
and AND4 (N691, N684, N603, N474, N652);
nand NAND2 (N692, N689, N483);
nor NOR4 (N693, N690, N633, N76, N229);
not NOT1 (N694, N665);
nor NOR2 (N695, N687, N221);
or OR2 (N696, N694, N298);
or OR3 (N697, N688, N361, N576);
not NOT1 (N698, N674);
or OR2 (N699, N698, N171);
or OR2 (N700, N685, N513);
xor XOR2 (N701, N700, N601);
and AND4 (N702, N686, N472, N690, N128);
nand NAND4 (N703, N695, N672, N693, N450);
and AND3 (N704, N133, N509, N685);
nand NAND4 (N705, N681, N632, N283, N509);
xor XOR2 (N706, N701, N252);
and AND2 (N707, N692, N512);
nor NOR4 (N708, N703, N538, N140, N72);
not NOT1 (N709, N699);
xor XOR2 (N710, N705, N571);
nor NOR2 (N711, N706, N308);
not NOT1 (N712, N708);
or OR4 (N713, N711, N99, N472, N487);
nand NAND4 (N714, N704, N638, N607, N472);
nor NOR3 (N715, N713, N303, N633);
nand NAND2 (N716, N697, N567);
not NOT1 (N717, N709);
not NOT1 (N718, N715);
or OR4 (N719, N702, N96, N403, N251);
nand NAND2 (N720, N718, N114);
not NOT1 (N721, N707);
xor XOR2 (N722, N712, N623);
nand NAND2 (N723, N691, N591);
buf BUF1 (N724, N716);
and AND4 (N725, N696, N686, N39, N163);
buf BUF1 (N726, N722);
nor NOR3 (N727, N724, N579, N545);
not NOT1 (N728, N720);
or OR4 (N729, N714, N96, N340, N444);
nor NOR4 (N730, N717, N6, N250, N350);
and AND3 (N731, N726, N608, N425);
and AND4 (N732, N731, N447, N526, N48);
xor XOR2 (N733, N710, N446);
or OR2 (N734, N733, N28);
nand NAND4 (N735, N728, N632, N445, N128);
and AND2 (N736, N721, N359);
or OR4 (N737, N732, N198, N567, N656);
xor XOR2 (N738, N729, N643);
buf BUF1 (N739, N730);
or OR2 (N740, N723, N525);
or OR3 (N741, N738, N69, N431);
or OR2 (N742, N739, N672);
nand NAND3 (N743, N741, N529, N318);
nor NOR4 (N744, N742, N50, N261, N297);
or OR4 (N745, N735, N103, N710, N430);
not NOT1 (N746, N719);
or OR2 (N747, N745, N380);
not NOT1 (N748, N746);
xor XOR2 (N749, N737, N172);
not NOT1 (N750, N740);
and AND3 (N751, N736, N617, N98);
and AND4 (N752, N725, N652, N434, N500);
nor NOR4 (N753, N744, N332, N569, N357);
nand NAND3 (N754, N734, N68, N184);
nor NOR4 (N755, N752, N561, N108, N514);
xor XOR2 (N756, N754, N715);
nand NAND4 (N757, N750, N735, N20, N274);
nor NOR4 (N758, N743, N45, N681, N485);
nor NOR2 (N759, N751, N421);
buf BUF1 (N760, N749);
or OR3 (N761, N755, N7, N505);
or OR3 (N762, N761, N237, N115);
not NOT1 (N763, N748);
not NOT1 (N764, N727);
nand NAND2 (N765, N759, N15);
nor NOR4 (N766, N764, N36, N741, N457);
nand NAND3 (N767, N747, N320, N6);
nand NAND3 (N768, N762, N710, N505);
buf BUF1 (N769, N763);
or OR4 (N770, N757, N310, N715, N746);
and AND2 (N771, N766, N205);
nand NAND3 (N772, N760, N662, N653);
nand NAND3 (N773, N769, N156, N324);
nor NOR4 (N774, N758, N581, N715, N81);
not NOT1 (N775, N770);
buf BUF1 (N776, N756);
not NOT1 (N777, N776);
xor XOR2 (N778, N768, N497);
or OR2 (N779, N773, N356);
nor NOR2 (N780, N753, N429);
not NOT1 (N781, N774);
not NOT1 (N782, N779);
not NOT1 (N783, N781);
buf BUF1 (N784, N778);
nor NOR4 (N785, N775, N520, N366, N75);
not NOT1 (N786, N777);
buf BUF1 (N787, N783);
nor NOR2 (N788, N771, N87);
nor NOR4 (N789, N780, N132, N596, N569);
and AND2 (N790, N767, N673);
nand NAND2 (N791, N788, N398);
nor NOR4 (N792, N785, N694, N790, N739);
buf BUF1 (N793, N527);
nand NAND2 (N794, N792, N792);
and AND3 (N795, N791, N239, N557);
buf BUF1 (N796, N765);
and AND2 (N797, N782, N538);
nand NAND2 (N798, N795, N56);
nand NAND3 (N799, N786, N39, N145);
nand NAND4 (N800, N789, N136, N408, N514);
and AND2 (N801, N796, N642);
nand NAND3 (N802, N798, N229, N712);
or OR2 (N803, N793, N207);
xor XOR2 (N804, N787, N574);
nand NAND4 (N805, N797, N265, N87, N84);
nand NAND2 (N806, N803, N266);
xor XOR2 (N807, N802, N227);
nand NAND3 (N808, N804, N609, N767);
xor XOR2 (N809, N808, N202);
nor NOR2 (N810, N807, N455);
nor NOR2 (N811, N806, N73);
buf BUF1 (N812, N784);
or OR2 (N813, N811, N58);
buf BUF1 (N814, N813);
or OR3 (N815, N812, N193, N219);
and AND2 (N816, N799, N766);
buf BUF1 (N817, N794);
or OR3 (N818, N815, N67, N293);
nand NAND3 (N819, N800, N749, N599);
nand NAND3 (N820, N810, N259, N277);
nor NOR2 (N821, N816, N305);
and AND2 (N822, N818, N694);
xor XOR2 (N823, N805, N304);
and AND4 (N824, N823, N360, N241, N192);
nand NAND4 (N825, N817, N101, N576, N24);
nor NOR2 (N826, N821, N305);
nand NAND3 (N827, N809, N563, N506);
nor NOR4 (N828, N827, N142, N352, N270);
not NOT1 (N829, N828);
not NOT1 (N830, N772);
nor NOR2 (N831, N830, N789);
buf BUF1 (N832, N822);
not NOT1 (N833, N820);
buf BUF1 (N834, N801);
xor XOR2 (N835, N826, N676);
or OR2 (N836, N829, N299);
buf BUF1 (N837, N819);
nand NAND4 (N838, N837, N91, N363, N496);
nand NAND2 (N839, N814, N220);
nor NOR3 (N840, N832, N90, N809);
nand NAND4 (N841, N836, N664, N638, N497);
nand NAND3 (N842, N838, N542, N345);
not NOT1 (N843, N839);
and AND2 (N844, N825, N555);
nand NAND4 (N845, N835, N407, N769, N695);
and AND4 (N846, N840, N807, N279, N600);
nand NAND4 (N847, N833, N651, N380, N702);
nor NOR2 (N848, N842, N329);
not NOT1 (N849, N824);
nand NAND3 (N850, N845, N822, N812);
or OR3 (N851, N849, N412, N554);
nor NOR3 (N852, N850, N692, N167);
and AND4 (N853, N843, N457, N747, N262);
nand NAND2 (N854, N841, N19);
xor XOR2 (N855, N848, N571);
xor XOR2 (N856, N851, N515);
or OR3 (N857, N831, N533, N386);
not NOT1 (N858, N844);
xor XOR2 (N859, N852, N837);
buf BUF1 (N860, N859);
nor NOR4 (N861, N855, N23, N526, N378);
buf BUF1 (N862, N856);
and AND2 (N863, N860, N459);
or OR2 (N864, N861, N115);
buf BUF1 (N865, N863);
and AND2 (N866, N862, N116);
nor NOR3 (N867, N834, N383, N404);
nor NOR4 (N868, N865, N480, N242, N518);
nand NAND2 (N869, N854, N734);
xor XOR2 (N870, N868, N519);
not NOT1 (N871, N870);
buf BUF1 (N872, N858);
nand NAND2 (N873, N866, N412);
xor XOR2 (N874, N847, N608);
buf BUF1 (N875, N864);
or OR3 (N876, N867, N739, N542);
not NOT1 (N877, N875);
xor XOR2 (N878, N874, N365);
xor XOR2 (N879, N857, N398);
and AND2 (N880, N876, N752);
and AND2 (N881, N877, N349);
nor NOR3 (N882, N871, N29, N543);
and AND3 (N883, N879, N7, N400);
nor NOR3 (N884, N880, N384, N66);
or OR2 (N885, N883, N776);
or OR2 (N886, N869, N148);
nor NOR2 (N887, N885, N748);
and AND2 (N888, N881, N877);
not NOT1 (N889, N884);
or OR3 (N890, N872, N453, N540);
nor NOR2 (N891, N889, N55);
nand NAND2 (N892, N853, N66);
and AND3 (N893, N886, N117, N659);
or OR3 (N894, N887, N119, N267);
nor NOR4 (N895, N882, N19, N263, N815);
or OR2 (N896, N846, N294);
buf BUF1 (N897, N873);
and AND2 (N898, N893, N74);
and AND2 (N899, N895, N441);
and AND2 (N900, N888, N521);
not NOT1 (N901, N897);
nor NOR4 (N902, N901, N836, N376, N286);
or OR4 (N903, N894, N686, N389, N35);
and AND4 (N904, N890, N28, N748, N207);
not NOT1 (N905, N898);
or OR2 (N906, N902, N879);
or OR4 (N907, N896, N810, N763, N568);
nor NOR4 (N908, N899, N219, N537, N194);
and AND2 (N909, N891, N607);
nand NAND2 (N910, N878, N84);
xor XOR2 (N911, N907, N460);
nand NAND4 (N912, N909, N227, N150, N853);
not NOT1 (N913, N905);
not NOT1 (N914, N912);
not NOT1 (N915, N892);
not NOT1 (N916, N913);
xor XOR2 (N917, N904, N371);
or OR3 (N918, N900, N38, N559);
and AND2 (N919, N911, N854);
not NOT1 (N920, N915);
nor NOR2 (N921, N914, N740);
or OR3 (N922, N921, N4, N240);
xor XOR2 (N923, N906, N162);
and AND4 (N924, N908, N455, N134, N168);
nor NOR2 (N925, N918, N670);
nor NOR3 (N926, N923, N599, N642);
nor NOR4 (N927, N916, N776, N536, N163);
buf BUF1 (N928, N917);
xor XOR2 (N929, N903, N791);
nor NOR2 (N930, N928, N282);
and AND2 (N931, N926, N466);
nor NOR4 (N932, N922, N111, N408, N627);
and AND3 (N933, N910, N313, N446);
not NOT1 (N934, N932);
not NOT1 (N935, N929);
nor NOR3 (N936, N930, N288, N553);
xor XOR2 (N937, N934, N815);
buf BUF1 (N938, N937);
not NOT1 (N939, N927);
not NOT1 (N940, N924);
not NOT1 (N941, N931);
xor XOR2 (N942, N940, N938);
nor NOR3 (N943, N22, N720, N915);
xor XOR2 (N944, N941, N684);
buf BUF1 (N945, N925);
buf BUF1 (N946, N945);
and AND4 (N947, N939, N480, N209, N107);
buf BUF1 (N948, N944);
nor NOR4 (N949, N946, N948, N831, N561);
xor XOR2 (N950, N563, N100);
nor NOR4 (N951, N936, N699, N656, N337);
nand NAND2 (N952, N920, N365);
or OR4 (N953, N942, N102, N296, N841);
xor XOR2 (N954, N951, N562);
and AND3 (N955, N947, N236, N369);
nor NOR2 (N956, N949, N737);
nor NOR2 (N957, N950, N30);
or OR4 (N958, N955, N383, N391, N304);
not NOT1 (N959, N956);
nor NOR4 (N960, N943, N449, N275, N848);
and AND4 (N961, N919, N835, N671, N617);
xor XOR2 (N962, N960, N199);
buf BUF1 (N963, N962);
xor XOR2 (N964, N963, N268);
not NOT1 (N965, N953);
and AND3 (N966, N933, N902, N161);
and AND4 (N967, N961, N706, N643, N470);
or OR4 (N968, N952, N467, N538, N621);
or OR4 (N969, N958, N640, N949, N878);
nor NOR3 (N970, N967, N475, N201);
not NOT1 (N971, N959);
buf BUF1 (N972, N971);
nand NAND3 (N973, N966, N836, N571);
not NOT1 (N974, N964);
xor XOR2 (N975, N973, N416);
xor XOR2 (N976, N974, N373);
buf BUF1 (N977, N935);
nand NAND4 (N978, N975, N505, N826, N8);
xor XOR2 (N979, N954, N368);
not NOT1 (N980, N965);
xor XOR2 (N981, N968, N545);
xor XOR2 (N982, N976, N252);
nand NAND4 (N983, N972, N594, N301, N272);
or OR4 (N984, N969, N291, N56, N324);
xor XOR2 (N985, N957, N983);
not NOT1 (N986, N796);
xor XOR2 (N987, N970, N314);
not NOT1 (N988, N978);
xor XOR2 (N989, N987, N230);
buf BUF1 (N990, N977);
or OR2 (N991, N988, N657);
buf BUF1 (N992, N989);
xor XOR2 (N993, N981, N200);
or OR3 (N994, N992, N207, N481);
not NOT1 (N995, N990);
and AND4 (N996, N995, N283, N668, N937);
nand NAND3 (N997, N996, N240, N993);
xor XOR2 (N998, N548, N615);
nand NAND4 (N999, N982, N633, N411, N265);
or OR2 (N1000, N998, N381);
buf BUF1 (N1001, N979);
nand NAND2 (N1002, N1001, N741);
or OR2 (N1003, N994, N621);
buf BUF1 (N1004, N991);
buf BUF1 (N1005, N984);
buf BUF1 (N1006, N1002);
and AND3 (N1007, N1003, N77, N709);
xor XOR2 (N1008, N1005, N695);
nand NAND2 (N1009, N1006, N115);
nor NOR2 (N1010, N1007, N622);
not NOT1 (N1011, N999);
xor XOR2 (N1012, N980, N730);
nor NOR4 (N1013, N1010, N711, N532, N701);
nand NAND2 (N1014, N1008, N315);
and AND3 (N1015, N1012, N625, N16);
or OR3 (N1016, N985, N69, N425);
and AND3 (N1017, N1014, N491, N211);
not NOT1 (N1018, N1000);
nand NAND3 (N1019, N986, N542, N771);
xor XOR2 (N1020, N997, N167);
or OR2 (N1021, N1018, N442);
nor NOR3 (N1022, N1017, N862, N859);
buf BUF1 (N1023, N1015);
and AND4 (N1024, N1016, N471, N820, N53);
and AND2 (N1025, N1020, N291);
buf BUF1 (N1026, N1022);
nor NOR3 (N1027, N1026, N505, N969);
or OR2 (N1028, N1025, N959);
and AND4 (N1029, N1028, N956, N631, N579);
xor XOR2 (N1030, N1029, N819);
nor NOR3 (N1031, N1019, N784, N116);
nand NAND2 (N1032, N1031, N926);
xor XOR2 (N1033, N1021, N667);
not NOT1 (N1034, N1013);
nand NAND3 (N1035, N1009, N694, N467);
xor XOR2 (N1036, N1032, N803);
or OR2 (N1037, N1034, N697);
and AND4 (N1038, N1033, N839, N849, N562);
and AND2 (N1039, N1027, N416);
buf BUF1 (N1040, N1037);
or OR3 (N1041, N1030, N827, N266);
buf BUF1 (N1042, N1038);
buf BUF1 (N1043, N1023);
nor NOR3 (N1044, N1039, N927, N110);
nor NOR4 (N1045, N1040, N778, N309, N902);
buf BUF1 (N1046, N1024);
not NOT1 (N1047, N1004);
or OR2 (N1048, N1035, N1016);
and AND2 (N1049, N1048, N889);
not NOT1 (N1050, N1043);
or OR2 (N1051, N1036, N792);
buf BUF1 (N1052, N1049);
xor XOR2 (N1053, N1047, N581);
nor NOR3 (N1054, N1053, N450, N994);
or OR2 (N1055, N1052, N981);
buf BUF1 (N1056, N1050);
not NOT1 (N1057, N1046);
nand NAND4 (N1058, N1044, N1024, N322, N303);
xor XOR2 (N1059, N1058, N509);
xor XOR2 (N1060, N1056, N460);
or OR4 (N1061, N1055, N455, N189, N337);
or OR3 (N1062, N1011, N410, N323);
xor XOR2 (N1063, N1059, N820);
buf BUF1 (N1064, N1051);
not NOT1 (N1065, N1045);
not NOT1 (N1066, N1042);
and AND4 (N1067, N1054, N1003, N67, N6);
or OR3 (N1068, N1062, N745, N829);
buf BUF1 (N1069, N1067);
xor XOR2 (N1070, N1069, N872);
not NOT1 (N1071, N1066);
buf BUF1 (N1072, N1061);
and AND4 (N1073, N1072, N378, N381, N652);
nand NAND3 (N1074, N1063, N600, N302);
or OR3 (N1075, N1064, N410, N61);
not NOT1 (N1076, N1070);
or OR3 (N1077, N1068, N288, N737);
and AND3 (N1078, N1073, N777, N456);
buf BUF1 (N1079, N1076);
nor NOR4 (N1080, N1075, N351, N965, N209);
xor XOR2 (N1081, N1057, N519);
and AND4 (N1082, N1077, N603, N580, N453);
xor XOR2 (N1083, N1074, N819);
xor XOR2 (N1084, N1071, N23);
xor XOR2 (N1085, N1081, N128);
and AND4 (N1086, N1083, N192, N777, N89);
xor XOR2 (N1087, N1078, N206);
nand NAND3 (N1088, N1065, N90, N468);
xor XOR2 (N1089, N1080, N316);
not NOT1 (N1090, N1089);
buf BUF1 (N1091, N1090);
not NOT1 (N1092, N1087);
buf BUF1 (N1093, N1085);
nand NAND3 (N1094, N1092, N679, N347);
and AND2 (N1095, N1079, N816);
not NOT1 (N1096, N1095);
or OR3 (N1097, N1041, N55, N20);
not NOT1 (N1098, N1094);
and AND2 (N1099, N1097, N370);
and AND4 (N1100, N1093, N318, N974, N166);
buf BUF1 (N1101, N1060);
not NOT1 (N1102, N1099);
and AND4 (N1103, N1086, N1031, N43, N119);
buf BUF1 (N1104, N1084);
nor NOR4 (N1105, N1103, N637, N535, N278);
xor XOR2 (N1106, N1104, N831);
xor XOR2 (N1107, N1102, N879);
nand NAND2 (N1108, N1107, N274);
and AND2 (N1109, N1100, N1077);
xor XOR2 (N1110, N1108, N4);
not NOT1 (N1111, N1105);
and AND3 (N1112, N1101, N668, N500);
nand NAND3 (N1113, N1109, N501, N695);
xor XOR2 (N1114, N1112, N1017);
nor NOR3 (N1115, N1091, N805, N987);
nand NAND2 (N1116, N1088, N174);
or OR4 (N1117, N1116, N601, N82, N765);
or OR4 (N1118, N1098, N753, N924, N856);
or OR2 (N1119, N1118, N988);
buf BUF1 (N1120, N1082);
and AND3 (N1121, N1113, N978, N1116);
xor XOR2 (N1122, N1106, N487);
not NOT1 (N1123, N1096);
and AND4 (N1124, N1114, N581, N1025, N205);
nand NAND4 (N1125, N1122, N224, N1052, N817);
buf BUF1 (N1126, N1124);
and AND2 (N1127, N1111, N945);
xor XOR2 (N1128, N1125, N505);
and AND3 (N1129, N1115, N597, N1061);
and AND2 (N1130, N1119, N257);
nor NOR2 (N1131, N1120, N793);
nand NAND2 (N1132, N1117, N183);
nor NOR4 (N1133, N1132, N1055, N436, N375);
nor NOR3 (N1134, N1126, N612, N94);
xor XOR2 (N1135, N1110, N62);
buf BUF1 (N1136, N1127);
or OR2 (N1137, N1131, N45);
buf BUF1 (N1138, N1129);
nand NAND4 (N1139, N1134, N288, N427, N252);
nor NOR4 (N1140, N1138, N776, N548, N43);
nand NAND2 (N1141, N1139, N658);
xor XOR2 (N1142, N1137, N37);
nor NOR2 (N1143, N1135, N987);
nand NAND3 (N1144, N1128, N1060, N306);
xor XOR2 (N1145, N1123, N493);
xor XOR2 (N1146, N1141, N52);
and AND3 (N1147, N1121, N903, N670);
nand NAND3 (N1148, N1146, N502, N106);
and AND2 (N1149, N1130, N461);
buf BUF1 (N1150, N1133);
nand NAND3 (N1151, N1145, N1099, N1013);
nand NAND4 (N1152, N1136, N175, N336, N933);
or OR2 (N1153, N1143, N138);
nor NOR2 (N1154, N1140, N378);
and AND4 (N1155, N1147, N1017, N645, N24);
or OR4 (N1156, N1155, N1148, N1142, N247);
or OR4 (N1157, N404, N1020, N273, N926);
and AND3 (N1158, N587, N122, N340);
nand NAND4 (N1159, N1156, N238, N792, N338);
xor XOR2 (N1160, N1149, N1000);
and AND3 (N1161, N1157, N859, N185);
xor XOR2 (N1162, N1144, N172);
not NOT1 (N1163, N1151);
buf BUF1 (N1164, N1158);
and AND3 (N1165, N1161, N621, N450);
nand NAND4 (N1166, N1160, N919, N872, N496);
nor NOR2 (N1167, N1164, N352);
nor NOR2 (N1168, N1165, N352);
not NOT1 (N1169, N1162);
xor XOR2 (N1170, N1168, N786);
buf BUF1 (N1171, N1163);
buf BUF1 (N1172, N1154);
buf BUF1 (N1173, N1170);
and AND2 (N1174, N1171, N305);
xor XOR2 (N1175, N1167, N1113);
xor XOR2 (N1176, N1172, N493);
nor NOR4 (N1177, N1174, N94, N776, N301);
not NOT1 (N1178, N1150);
not NOT1 (N1179, N1176);
not NOT1 (N1180, N1169);
or OR4 (N1181, N1179, N463, N502, N219);
and AND2 (N1182, N1175, N5);
and AND4 (N1183, N1152, N863, N670, N1024);
nand NAND3 (N1184, N1178, N791, N997);
xor XOR2 (N1185, N1166, N61);
not NOT1 (N1186, N1183);
not NOT1 (N1187, N1182);
xor XOR2 (N1188, N1187, N220);
xor XOR2 (N1189, N1181, N945);
not NOT1 (N1190, N1185);
or OR3 (N1191, N1186, N1185, N593);
nor NOR2 (N1192, N1177, N399);
or OR2 (N1193, N1189, N332);
and AND2 (N1194, N1192, N860);
nand NAND2 (N1195, N1188, N926);
xor XOR2 (N1196, N1195, N1098);
nand NAND2 (N1197, N1180, N163);
and AND3 (N1198, N1159, N536, N926);
not NOT1 (N1199, N1190);
nand NAND3 (N1200, N1153, N225, N780);
or OR2 (N1201, N1198, N831);
xor XOR2 (N1202, N1191, N123);
not NOT1 (N1203, N1173);
not NOT1 (N1204, N1193);
and AND4 (N1205, N1199, N666, N735, N1090);
or OR3 (N1206, N1184, N363, N381);
not NOT1 (N1207, N1201);
nor NOR3 (N1208, N1205, N496, N1107);
nand NAND3 (N1209, N1206, N1104, N811);
or OR2 (N1210, N1203, N915);
xor XOR2 (N1211, N1204, N45);
or OR3 (N1212, N1200, N1094, N711);
nor NOR4 (N1213, N1194, N692, N581, N193);
or OR3 (N1214, N1197, N170, N209);
nand NAND2 (N1215, N1207, N795);
xor XOR2 (N1216, N1202, N782);
and AND3 (N1217, N1215, N628, N316);
nand NAND3 (N1218, N1217, N662, N704);
or OR2 (N1219, N1211, N286);
not NOT1 (N1220, N1196);
buf BUF1 (N1221, N1218);
or OR2 (N1222, N1221, N172);
nor NOR2 (N1223, N1210, N1066);
nand NAND2 (N1224, N1213, N464);
and AND3 (N1225, N1208, N468, N871);
nor NOR4 (N1226, N1222, N263, N345, N578);
nor NOR4 (N1227, N1214, N220, N1186, N1006);
nor NOR4 (N1228, N1224, N830, N525, N829);
nor NOR2 (N1229, N1223, N395);
nand NAND3 (N1230, N1216, N936, N791);
nor NOR4 (N1231, N1220, N1230, N396, N744);
xor XOR2 (N1232, N596, N1028);
nor NOR3 (N1233, N1225, N256, N825);
not NOT1 (N1234, N1219);
not NOT1 (N1235, N1227);
xor XOR2 (N1236, N1231, N1111);
nor NOR3 (N1237, N1236, N628, N120);
xor XOR2 (N1238, N1209, N458);
or OR2 (N1239, N1229, N1128);
nand NAND2 (N1240, N1237, N331);
and AND3 (N1241, N1234, N774, N216);
or OR3 (N1242, N1238, N245, N623);
xor XOR2 (N1243, N1228, N859);
nor NOR2 (N1244, N1243, N584);
buf BUF1 (N1245, N1232);
and AND4 (N1246, N1241, N38, N111, N5);
not NOT1 (N1247, N1245);
nor NOR4 (N1248, N1246, N149, N471, N879);
nor NOR4 (N1249, N1244, N51, N848, N292);
xor XOR2 (N1250, N1240, N790);
nand NAND3 (N1251, N1212, N888, N103);
or OR3 (N1252, N1247, N510, N1248);
not NOT1 (N1253, N741);
xor XOR2 (N1254, N1226, N1211);
nor NOR2 (N1255, N1249, N519);
not NOT1 (N1256, N1254);
not NOT1 (N1257, N1255);
xor XOR2 (N1258, N1242, N935);
and AND4 (N1259, N1256, N948, N578, N700);
nor NOR2 (N1260, N1253, N920);
nand NAND2 (N1261, N1258, N637);
and AND4 (N1262, N1261, N651, N1154, N801);
or OR3 (N1263, N1233, N612, N223);
nand NAND4 (N1264, N1262, N1098, N1171, N273);
buf BUF1 (N1265, N1239);
xor XOR2 (N1266, N1252, N158);
or OR3 (N1267, N1250, N172, N603);
not NOT1 (N1268, N1263);
nand NAND2 (N1269, N1235, N406);
and AND4 (N1270, N1268, N223, N1235, N426);
nand NAND4 (N1271, N1269, N1241, N715, N676);
nor NOR3 (N1272, N1270, N1009, N750);
xor XOR2 (N1273, N1260, N1053);
xor XOR2 (N1274, N1267, N407);
nor NOR4 (N1275, N1273, N186, N838, N63);
nand NAND3 (N1276, N1275, N954, N687);
nand NAND3 (N1277, N1259, N170, N1198);
nand NAND3 (N1278, N1251, N1132, N1178);
xor XOR2 (N1279, N1264, N674);
buf BUF1 (N1280, N1276);
not NOT1 (N1281, N1274);
not NOT1 (N1282, N1271);
or OR3 (N1283, N1278, N462, N950);
not NOT1 (N1284, N1272);
nor NOR3 (N1285, N1283, N134, N1057);
and AND2 (N1286, N1281, N172);
nand NAND4 (N1287, N1265, N319, N821, N716);
or OR2 (N1288, N1257, N274);
xor XOR2 (N1289, N1280, N305);
and AND2 (N1290, N1284, N128);
xor XOR2 (N1291, N1288, N635);
nor NOR4 (N1292, N1291, N91, N302, N1267);
nor NOR3 (N1293, N1287, N1116, N833);
nand NAND2 (N1294, N1266, N1121);
nor NOR4 (N1295, N1289, N229, N949, N188);
buf BUF1 (N1296, N1286);
not NOT1 (N1297, N1293);
and AND4 (N1298, N1296, N496, N469, N1261);
xor XOR2 (N1299, N1298, N1165);
nand NAND4 (N1300, N1277, N559, N823, N288);
nand NAND3 (N1301, N1290, N988, N462);
not NOT1 (N1302, N1295);
nand NAND4 (N1303, N1279, N581, N1285, N787);
nand NAND4 (N1304, N1173, N976, N424, N1188);
buf BUF1 (N1305, N1300);
xor XOR2 (N1306, N1304, N662);
buf BUF1 (N1307, N1282);
not NOT1 (N1308, N1299);
not NOT1 (N1309, N1292);
nand NAND3 (N1310, N1306, N478, N1148);
buf BUF1 (N1311, N1310);
not NOT1 (N1312, N1311);
or OR4 (N1313, N1308, N796, N1106, N256);
not NOT1 (N1314, N1309);
nor NOR4 (N1315, N1303, N933, N597, N641);
and AND4 (N1316, N1313, N1186, N1037, N871);
and AND4 (N1317, N1315, N333, N1274, N184);
xor XOR2 (N1318, N1314, N416);
and AND2 (N1319, N1301, N357);
xor XOR2 (N1320, N1317, N1075);
not NOT1 (N1321, N1316);
nand NAND2 (N1322, N1312, N936);
or OR4 (N1323, N1302, N998, N401, N268);
buf BUF1 (N1324, N1297);
xor XOR2 (N1325, N1324, N698);
and AND2 (N1326, N1322, N367);
xor XOR2 (N1327, N1325, N94);
not NOT1 (N1328, N1319);
xor XOR2 (N1329, N1307, N257);
xor XOR2 (N1330, N1320, N104);
xor XOR2 (N1331, N1328, N224);
nand NAND3 (N1332, N1294, N425, N1266);
xor XOR2 (N1333, N1331, N896);
and AND2 (N1334, N1330, N1302);
nor NOR4 (N1335, N1318, N134, N80, N152);
nor NOR4 (N1336, N1333, N23, N835, N313);
nand NAND4 (N1337, N1336, N737, N662, N739);
and AND4 (N1338, N1335, N1284, N51, N353);
and AND4 (N1339, N1326, N913, N1033, N1217);
xor XOR2 (N1340, N1329, N1204);
buf BUF1 (N1341, N1323);
xor XOR2 (N1342, N1341, N1100);
nand NAND4 (N1343, N1321, N257, N151, N1166);
buf BUF1 (N1344, N1342);
or OR3 (N1345, N1327, N1306, N278);
nand NAND4 (N1346, N1340, N504, N604, N33);
xor XOR2 (N1347, N1332, N1285);
xor XOR2 (N1348, N1345, N211);
nand NAND4 (N1349, N1344, N1291, N661, N23);
nand NAND4 (N1350, N1343, N313, N731, N28);
buf BUF1 (N1351, N1350);
and AND2 (N1352, N1305, N987);
xor XOR2 (N1353, N1347, N977);
or OR4 (N1354, N1346, N66, N1207, N470);
nand NAND3 (N1355, N1348, N1075, N515);
and AND3 (N1356, N1338, N1045, N771);
xor XOR2 (N1357, N1337, N365);
nor NOR2 (N1358, N1353, N967);
xor XOR2 (N1359, N1356, N635);
buf BUF1 (N1360, N1354);
or OR3 (N1361, N1360, N426, N691);
not NOT1 (N1362, N1349);
nand NAND4 (N1363, N1359, N777, N1021, N142);
or OR2 (N1364, N1334, N918);
or OR3 (N1365, N1339, N100, N1098);
nand NAND3 (N1366, N1365, N1158, N1265);
xor XOR2 (N1367, N1362, N121);
xor XOR2 (N1368, N1366, N470);
not NOT1 (N1369, N1364);
not NOT1 (N1370, N1352);
xor XOR2 (N1371, N1361, N1061);
nor NOR2 (N1372, N1357, N144);
xor XOR2 (N1373, N1368, N813);
xor XOR2 (N1374, N1370, N1064);
nand NAND2 (N1375, N1358, N209);
xor XOR2 (N1376, N1367, N1272);
and AND3 (N1377, N1369, N1095, N645);
and AND4 (N1378, N1373, N1368, N573, N1221);
not NOT1 (N1379, N1378);
not NOT1 (N1380, N1355);
nor NOR4 (N1381, N1376, N129, N888, N401);
nor NOR3 (N1382, N1381, N746, N46);
not NOT1 (N1383, N1372);
or OR2 (N1384, N1380, N422);
or OR3 (N1385, N1377, N913, N602);
and AND2 (N1386, N1385, N339);
nand NAND4 (N1387, N1371, N168, N1059, N397);
nand NAND4 (N1388, N1383, N681, N833, N116);
or OR3 (N1389, N1363, N611, N680);
or OR4 (N1390, N1386, N176, N154, N252);
xor XOR2 (N1391, N1389, N362);
xor XOR2 (N1392, N1390, N642);
or OR3 (N1393, N1391, N547, N844);
and AND3 (N1394, N1375, N858, N522);
nand NAND3 (N1395, N1374, N298, N1316);
not NOT1 (N1396, N1395);
xor XOR2 (N1397, N1394, N19);
not NOT1 (N1398, N1387);
xor XOR2 (N1399, N1379, N320);
nand NAND4 (N1400, N1398, N338, N1006, N638);
buf BUF1 (N1401, N1393);
not NOT1 (N1402, N1400);
nand NAND4 (N1403, N1399, N559, N898, N47);
and AND2 (N1404, N1384, N205);
nand NAND4 (N1405, N1401, N1019, N517, N978);
xor XOR2 (N1406, N1405, N377);
or OR4 (N1407, N1382, N1221, N151, N797);
nand NAND4 (N1408, N1407, N214, N1221, N1169);
nor NOR2 (N1409, N1388, N445);
or OR2 (N1410, N1402, N1273);
buf BUF1 (N1411, N1409);
or OR4 (N1412, N1392, N1008, N1316, N59);
not NOT1 (N1413, N1404);
not NOT1 (N1414, N1412);
and AND3 (N1415, N1414, N1333, N1132);
buf BUF1 (N1416, N1415);
xor XOR2 (N1417, N1413, N782);
not NOT1 (N1418, N1416);
nor NOR4 (N1419, N1351, N800, N1383, N963);
and AND3 (N1420, N1406, N221, N1101);
buf BUF1 (N1421, N1396);
and AND2 (N1422, N1403, N949);
buf BUF1 (N1423, N1419);
nand NAND4 (N1424, N1420, N640, N291, N797);
nor NOR3 (N1425, N1411, N82, N791);
buf BUF1 (N1426, N1397);
xor XOR2 (N1427, N1423, N766);
or OR4 (N1428, N1421, N805, N924, N661);
not NOT1 (N1429, N1422);
buf BUF1 (N1430, N1425);
not NOT1 (N1431, N1418);
nand NAND3 (N1432, N1431, N733, N1274);
buf BUF1 (N1433, N1432);
nand NAND3 (N1434, N1424, N883, N749);
nor NOR4 (N1435, N1417, N1333, N645, N1227);
buf BUF1 (N1436, N1429);
buf BUF1 (N1437, N1427);
xor XOR2 (N1438, N1410, N19);
nor NOR4 (N1439, N1430, N1052, N1248, N1196);
or OR3 (N1440, N1436, N1162, N194);
nor NOR3 (N1441, N1437, N220, N726);
and AND4 (N1442, N1441, N530, N1229, N723);
nor NOR2 (N1443, N1435, N55);
xor XOR2 (N1444, N1442, N996);
nor NOR2 (N1445, N1438, N1259);
xor XOR2 (N1446, N1408, N1170);
buf BUF1 (N1447, N1440);
xor XOR2 (N1448, N1434, N310);
nor NOR2 (N1449, N1426, N1039);
nor NOR3 (N1450, N1439, N751, N507);
nand NAND4 (N1451, N1444, N248, N648, N21);
nor NOR4 (N1452, N1447, N540, N1048, N1168);
buf BUF1 (N1453, N1448);
nor NOR3 (N1454, N1433, N304, N1023);
not NOT1 (N1455, N1445);
and AND2 (N1456, N1428, N271);
or OR3 (N1457, N1455, N26, N276);
and AND3 (N1458, N1446, N5, N536);
nor NOR4 (N1459, N1458, N61, N831, N1042);
not NOT1 (N1460, N1456);
buf BUF1 (N1461, N1459);
buf BUF1 (N1462, N1452);
nand NAND4 (N1463, N1443, N1374, N822, N103);
buf BUF1 (N1464, N1453);
nor NOR4 (N1465, N1460, N417, N810, N1144);
or OR2 (N1466, N1449, N368);
nor NOR4 (N1467, N1466, N83, N1148, N639);
and AND4 (N1468, N1461, N1117, N256, N1303);
buf BUF1 (N1469, N1463);
not NOT1 (N1470, N1467);
not NOT1 (N1471, N1464);
nor NOR4 (N1472, N1470, N1322, N10, N880);
nor NOR4 (N1473, N1454, N326, N363, N356);
nand NAND3 (N1474, N1471, N1120, N752);
and AND3 (N1475, N1457, N514, N235);
or OR2 (N1476, N1465, N893);
and AND4 (N1477, N1468, N417, N236, N1018);
not NOT1 (N1478, N1477);
nand NAND2 (N1479, N1478, N566);
xor XOR2 (N1480, N1469, N651);
or OR3 (N1481, N1480, N127, N1419);
buf BUF1 (N1482, N1472);
nor NOR3 (N1483, N1462, N482, N1351);
nand NAND2 (N1484, N1481, N365);
and AND4 (N1485, N1474, N256, N965, N1356);
or OR2 (N1486, N1475, N8);
nor NOR2 (N1487, N1451, N769);
nor NOR4 (N1488, N1482, N682, N46, N1110);
nand NAND3 (N1489, N1479, N206, N769);
xor XOR2 (N1490, N1483, N979);
nor NOR2 (N1491, N1476, N703);
xor XOR2 (N1492, N1487, N955);
not NOT1 (N1493, N1485);
nand NAND4 (N1494, N1492, N651, N1116, N1293);
xor XOR2 (N1495, N1489, N1166);
or OR3 (N1496, N1491, N1452, N1003);
xor XOR2 (N1497, N1473, N864);
nor NOR4 (N1498, N1490, N996, N34, N2);
nor NOR2 (N1499, N1496, N1414);
nand NAND2 (N1500, N1493, N1224);
or OR2 (N1501, N1499, N1374);
nor NOR2 (N1502, N1495, N1464);
not NOT1 (N1503, N1497);
nor NOR2 (N1504, N1501, N1416);
xor XOR2 (N1505, N1488, N1128);
not NOT1 (N1506, N1450);
nand NAND3 (N1507, N1498, N257, N1337);
nor NOR3 (N1508, N1486, N1037, N703);
and AND3 (N1509, N1502, N1390, N225);
buf BUF1 (N1510, N1484);
not NOT1 (N1511, N1507);
xor XOR2 (N1512, N1500, N562);
xor XOR2 (N1513, N1505, N405);
buf BUF1 (N1514, N1511);
and AND2 (N1515, N1509, N1002);
and AND3 (N1516, N1510, N373, N320);
buf BUF1 (N1517, N1512);
nand NAND3 (N1518, N1504, N455, N1483);
nand NAND3 (N1519, N1517, N1197, N1372);
or OR2 (N1520, N1494, N1191);
xor XOR2 (N1521, N1519, N919);
nand NAND3 (N1522, N1506, N119, N1040);
nor NOR3 (N1523, N1514, N747, N1219);
and AND2 (N1524, N1522, N980);
and AND2 (N1525, N1516, N470);
not NOT1 (N1526, N1525);
and AND3 (N1527, N1503, N1421, N1341);
buf BUF1 (N1528, N1524);
not NOT1 (N1529, N1518);
xor XOR2 (N1530, N1508, N188);
nand NAND2 (N1531, N1530, N191);
buf BUF1 (N1532, N1520);
nand NAND4 (N1533, N1529, N446, N870, N582);
nor NOR3 (N1534, N1532, N559, N1250);
or OR4 (N1535, N1513, N709, N573, N287);
nand NAND3 (N1536, N1523, N376, N1208);
nand NAND2 (N1537, N1526, N682);
or OR2 (N1538, N1536, N1230);
not NOT1 (N1539, N1535);
nor NOR4 (N1540, N1537, N326, N187, N436);
buf BUF1 (N1541, N1533);
xor XOR2 (N1542, N1531, N1007);
not NOT1 (N1543, N1528);
not NOT1 (N1544, N1542);
nand NAND3 (N1545, N1540, N1221, N1359);
nor NOR4 (N1546, N1545, N626, N1400, N1172);
xor XOR2 (N1547, N1543, N656);
or OR4 (N1548, N1546, N462, N1084, N794);
and AND4 (N1549, N1521, N479, N1174, N950);
not NOT1 (N1550, N1527);
or OR3 (N1551, N1534, N566, N233);
and AND3 (N1552, N1541, N1008, N559);
or OR4 (N1553, N1552, N1389, N282, N134);
and AND2 (N1554, N1538, N1213);
buf BUF1 (N1555, N1549);
buf BUF1 (N1556, N1553);
or OR2 (N1557, N1556, N1012);
or OR2 (N1558, N1548, N795);
buf BUF1 (N1559, N1555);
or OR3 (N1560, N1515, N55, N664);
or OR3 (N1561, N1557, N839, N1340);
and AND2 (N1562, N1558, N307);
nand NAND2 (N1563, N1561, N125);
nor NOR4 (N1564, N1539, N346, N998, N201);
nand NAND2 (N1565, N1550, N928);
or OR4 (N1566, N1565, N1103, N962, N1552);
xor XOR2 (N1567, N1560, N1363);
buf BUF1 (N1568, N1554);
or OR4 (N1569, N1568, N1562, N256, N913);
nand NAND2 (N1570, N1085, N809);
xor XOR2 (N1571, N1570, N744);
and AND3 (N1572, N1569, N1473, N1332);
xor XOR2 (N1573, N1559, N273);
or OR2 (N1574, N1564, N151);
buf BUF1 (N1575, N1573);
nand NAND2 (N1576, N1551, N1088);
and AND4 (N1577, N1571, N973, N453, N129);
buf BUF1 (N1578, N1577);
and AND4 (N1579, N1563, N109, N143, N882);
not NOT1 (N1580, N1574);
nor NOR2 (N1581, N1580, N379);
nor NOR4 (N1582, N1572, N1326, N1096, N1279);
not NOT1 (N1583, N1576);
xor XOR2 (N1584, N1582, N1353);
nor NOR4 (N1585, N1566, N43, N1520, N987);
not NOT1 (N1586, N1584);
or OR4 (N1587, N1583, N28, N1440, N273);
xor XOR2 (N1588, N1547, N785);
buf BUF1 (N1589, N1575);
nor NOR4 (N1590, N1544, N1354, N312, N538);
nand NAND3 (N1591, N1588, N1455, N1366);
xor XOR2 (N1592, N1585, N683);
or OR2 (N1593, N1579, N28);
xor XOR2 (N1594, N1581, N1497);
nand NAND4 (N1595, N1590, N1112, N281, N1114);
and AND4 (N1596, N1587, N163, N228, N672);
and AND3 (N1597, N1592, N670, N1021);
and AND4 (N1598, N1586, N1500, N1574, N500);
nand NAND3 (N1599, N1567, N855, N623);
not NOT1 (N1600, N1595);
xor XOR2 (N1601, N1596, N726);
xor XOR2 (N1602, N1601, N436);
nand NAND3 (N1603, N1602, N663, N1389);
buf BUF1 (N1604, N1598);
not NOT1 (N1605, N1604);
not NOT1 (N1606, N1599);
not NOT1 (N1607, N1589);
or OR3 (N1608, N1603, N194, N26);
nand NAND3 (N1609, N1578, N379, N1441);
buf BUF1 (N1610, N1591);
or OR2 (N1611, N1606, N508);
nand NAND2 (N1612, N1607, N82);
nor NOR4 (N1613, N1605, N433, N527, N1303);
nor NOR3 (N1614, N1608, N1065, N393);
xor XOR2 (N1615, N1611, N556);
nor NOR3 (N1616, N1614, N18, N535);
xor XOR2 (N1617, N1613, N1101);
or OR3 (N1618, N1600, N1539, N703);
or OR3 (N1619, N1616, N117, N203);
buf BUF1 (N1620, N1594);
or OR3 (N1621, N1593, N1286, N1275);
nand NAND4 (N1622, N1617, N1051, N1267, N568);
or OR4 (N1623, N1610, N649, N1423, N1605);
and AND4 (N1624, N1609, N99, N342, N1409);
endmodule