// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17;

output N1604,N1594,N1603,N1616,N1606,N1614,N1607,N1612,N1608,N1617;

and AND2 (N18, N1, N12);
buf BUF1 (N19, N6);
or OR4 (N20, N13, N7, N17, N19);
not NOT1 (N21, N2);
nor NOR3 (N22, N6, N6, N2);
xor XOR2 (N23, N3, N5);
not NOT1 (N24, N9);
nor NOR4 (N25, N7, N4, N1, N19);
nand NAND2 (N26, N23, N12);
nor NOR3 (N27, N2, N21, N2);
xor XOR2 (N28, N22, N15);
buf BUF1 (N29, N12);
buf BUF1 (N30, N13);
xor XOR2 (N31, N2, N20);
or OR3 (N32, N10, N18, N16);
or OR3 (N33, N11, N15, N23);
not NOT1 (N34, N28);
and AND3 (N35, N32, N18, N3);
xor XOR2 (N36, N27, N20);
nor NOR4 (N37, N24, N19, N10, N32);
and AND4 (N38, N30, N3, N7, N24);
nor NOR2 (N39, N25, N13);
or OR3 (N40, N37, N32, N2);
nor NOR2 (N41, N31, N39);
not NOT1 (N42, N29);
buf BUF1 (N43, N18);
and AND3 (N44, N38, N20, N18);
or OR2 (N45, N36, N10);
nand NAND4 (N46, N43, N40, N45, N20);
or OR2 (N47, N21, N35);
xor XOR2 (N48, N28, N39);
and AND2 (N49, N4, N21);
nand NAND4 (N50, N42, N20, N45, N39);
and AND2 (N51, N44, N25);
and AND4 (N52, N34, N39, N24, N46);
xor XOR2 (N53, N14, N47);
and AND3 (N54, N12, N22, N37);
and AND3 (N55, N54, N24, N46);
nand NAND4 (N56, N33, N54, N50, N34);
nor NOR4 (N57, N44, N46, N18, N55);
and AND2 (N58, N34, N29);
and AND3 (N59, N26, N33, N19);
nand NAND4 (N60, N56, N19, N59, N12);
and AND2 (N61, N57, N5);
or OR3 (N62, N9, N30, N10);
nor NOR3 (N63, N61, N4, N23);
nand NAND2 (N64, N51, N38);
or OR3 (N65, N63, N1, N16);
nand NAND2 (N66, N52, N35);
or OR4 (N67, N53, N55, N55, N34);
not NOT1 (N68, N64);
nand NAND3 (N69, N49, N53, N38);
buf BUF1 (N70, N60);
nand NAND2 (N71, N65, N57);
and AND4 (N72, N69, N60, N32, N31);
nor NOR3 (N73, N48, N35, N70);
xor XOR2 (N74, N45, N23);
buf BUF1 (N75, N58);
buf BUF1 (N76, N67);
nor NOR3 (N77, N71, N74, N30);
xor XOR2 (N78, N61, N7);
nand NAND3 (N79, N75, N38, N35);
nand NAND2 (N80, N62, N75);
xor XOR2 (N81, N79, N34);
xor XOR2 (N82, N72, N59);
or OR3 (N83, N76, N77, N42);
buf BUF1 (N84, N12);
nand NAND4 (N85, N81, N29, N59, N43);
nand NAND4 (N86, N80, N43, N76, N85);
or OR3 (N87, N26, N19, N13);
or OR4 (N88, N87, N62, N4, N37);
nor NOR4 (N89, N86, N3, N63, N30);
nand NAND3 (N90, N82, N42, N79);
and AND4 (N91, N89, N46, N54, N34);
nand NAND2 (N92, N78, N54);
nand NAND3 (N93, N68, N89, N49);
buf BUF1 (N94, N66);
xor XOR2 (N95, N41, N43);
and AND4 (N96, N91, N55, N16, N35);
xor XOR2 (N97, N90, N8);
xor XOR2 (N98, N93, N5);
nand NAND2 (N99, N83, N54);
buf BUF1 (N100, N95);
nand NAND3 (N101, N97, N46, N26);
xor XOR2 (N102, N99, N69);
and AND2 (N103, N96, N69);
buf BUF1 (N104, N92);
buf BUF1 (N105, N84);
nand NAND4 (N106, N88, N28, N26, N36);
xor XOR2 (N107, N98, N54);
nor NOR2 (N108, N105, N66);
nor NOR3 (N109, N103, N33, N9);
nand NAND2 (N110, N106, N14);
not NOT1 (N111, N104);
nand NAND3 (N112, N109, N15, N83);
or OR2 (N113, N111, N47);
and AND4 (N114, N112, N44, N113, N93);
not NOT1 (N115, N92);
not NOT1 (N116, N114);
or OR3 (N117, N116, N89, N43);
nand NAND4 (N118, N110, N50, N27, N44);
nand NAND2 (N119, N107, N40);
xor XOR2 (N120, N94, N38);
nand NAND2 (N121, N101, N11);
nand NAND3 (N122, N100, N76, N100);
not NOT1 (N123, N115);
nand NAND3 (N124, N117, N1, N101);
nor NOR4 (N125, N120, N12, N98, N97);
buf BUF1 (N126, N73);
not NOT1 (N127, N102);
and AND4 (N128, N119, N66, N37, N121);
nor NOR2 (N129, N70, N13);
and AND2 (N130, N118, N24);
buf BUF1 (N131, N130);
xor XOR2 (N132, N127, N65);
buf BUF1 (N133, N124);
nor NOR4 (N134, N132, N4, N131, N131);
buf BUF1 (N135, N129);
xor XOR2 (N136, N24, N29);
and AND4 (N137, N123, N109, N112, N126);
nor NOR3 (N138, N72, N133, N28);
or OR2 (N139, N20, N82);
nor NOR3 (N140, N135, N53, N124);
or OR3 (N141, N108, N78, N3);
nor NOR2 (N142, N125, N27);
or OR3 (N143, N137, N69, N133);
xor XOR2 (N144, N138, N122);
buf BUF1 (N145, N27);
and AND3 (N146, N134, N53, N122);
nor NOR3 (N147, N143, N21, N110);
nand NAND2 (N148, N128, N93);
or OR4 (N149, N145, N3, N77, N124);
or OR2 (N150, N149, N58);
buf BUF1 (N151, N144);
nor NOR4 (N152, N146, N81, N5, N147);
xor XOR2 (N153, N124, N16);
nor NOR4 (N154, N151, N109, N72, N39);
buf BUF1 (N155, N141);
or OR4 (N156, N155, N144, N6, N75);
nor NOR2 (N157, N136, N147);
nand NAND3 (N158, N139, N136, N14);
nand NAND4 (N159, N152, N147, N88, N4);
or OR3 (N160, N156, N150, N8);
nor NOR4 (N161, N14, N57, N119, N83);
buf BUF1 (N162, N154);
not NOT1 (N163, N159);
or OR3 (N164, N163, N37, N20);
or OR4 (N165, N153, N49, N102, N81);
nand NAND4 (N166, N140, N12, N112, N133);
or OR3 (N167, N164, N111, N154);
nor NOR3 (N168, N158, N116, N96);
and AND2 (N169, N142, N91);
buf BUF1 (N170, N160);
not NOT1 (N171, N148);
xor XOR2 (N172, N168, N159);
or OR3 (N173, N157, N13, N137);
buf BUF1 (N174, N165);
nand NAND4 (N175, N162, N96, N144, N164);
not NOT1 (N176, N161);
nand NAND4 (N177, N172, N109, N97, N83);
buf BUF1 (N178, N173);
or OR4 (N179, N170, N111, N29, N120);
and AND4 (N180, N175, N86, N62, N96);
buf BUF1 (N181, N176);
nand NAND4 (N182, N180, N10, N80, N167);
nand NAND3 (N183, N83, N105, N63);
or OR2 (N184, N174, N176);
not NOT1 (N185, N171);
nor NOR3 (N186, N182, N31, N23);
buf BUF1 (N187, N181);
xor XOR2 (N188, N166, N85);
nand NAND4 (N189, N183, N121, N163, N135);
nand NAND4 (N190, N186, N44, N53, N4);
and AND3 (N191, N169, N31, N117);
nand NAND4 (N192, N185, N54, N134, N133);
xor XOR2 (N193, N184, N60);
buf BUF1 (N194, N188);
nor NOR3 (N195, N192, N178, N127);
or OR3 (N196, N51, N127, N145);
buf BUF1 (N197, N190);
xor XOR2 (N198, N187, N164);
or OR2 (N199, N177, N122);
xor XOR2 (N200, N193, N104);
nor NOR2 (N201, N197, N61);
xor XOR2 (N202, N189, N23);
buf BUF1 (N203, N196);
or OR3 (N204, N195, N123, N130);
and AND3 (N205, N204, N133, N96);
or OR2 (N206, N194, N62);
or OR2 (N207, N191, N19);
nor NOR2 (N208, N203, N37);
nor NOR2 (N209, N202, N75);
nand NAND3 (N210, N205, N152, N182);
nand NAND2 (N211, N206, N53);
nand NAND2 (N212, N179, N93);
not NOT1 (N213, N209);
buf BUF1 (N214, N212);
not NOT1 (N215, N199);
buf BUF1 (N216, N211);
not NOT1 (N217, N208);
and AND2 (N218, N200, N152);
xor XOR2 (N219, N214, N46);
and AND4 (N220, N198, N146, N216, N101);
or OR4 (N221, N114, N86, N75, N219);
xor XOR2 (N222, N93, N166);
nand NAND4 (N223, N217, N25, N99, N178);
buf BUF1 (N224, N213);
or OR2 (N225, N220, N215);
buf BUF1 (N226, N21);
nor NOR3 (N227, N210, N74, N11);
nand NAND2 (N228, N226, N67);
not NOT1 (N229, N225);
nand NAND2 (N230, N229, N30);
or OR3 (N231, N221, N6, N55);
nand NAND4 (N232, N228, N25, N158, N211);
nand NAND4 (N233, N231, N72, N218, N145);
xor XOR2 (N234, N221, N146);
nand NAND3 (N235, N230, N222, N9);
or OR3 (N236, N110, N67, N220);
nor NOR4 (N237, N234, N230, N164, N18);
and AND3 (N238, N233, N95, N118);
xor XOR2 (N239, N224, N74);
buf BUF1 (N240, N239);
nand NAND2 (N241, N238, N233);
buf BUF1 (N242, N235);
xor XOR2 (N243, N223, N35);
buf BUF1 (N244, N207);
and AND2 (N245, N241, N200);
buf BUF1 (N246, N236);
buf BUF1 (N247, N246);
xor XOR2 (N248, N243, N189);
nor NOR2 (N249, N240, N216);
nor NOR4 (N250, N249, N31, N214, N67);
and AND3 (N251, N232, N145, N8);
xor XOR2 (N252, N201, N88);
or OR2 (N253, N252, N134);
or OR3 (N254, N251, N117, N183);
nand NAND3 (N255, N242, N19, N34);
buf BUF1 (N256, N247);
nand NAND4 (N257, N244, N33, N183, N103);
nand NAND4 (N258, N256, N45, N199, N184);
nand NAND4 (N259, N250, N149, N107, N184);
nor NOR3 (N260, N254, N127, N191);
buf BUF1 (N261, N248);
buf BUF1 (N262, N261);
and AND3 (N263, N245, N79, N255);
nand NAND2 (N264, N183, N55);
nor NOR2 (N265, N264, N168);
or OR2 (N266, N258, N134);
not NOT1 (N267, N262);
nand NAND2 (N268, N265, N130);
nand NAND4 (N269, N237, N154, N175, N66);
and AND3 (N270, N260, N5, N3);
and AND4 (N271, N266, N153, N230, N265);
not NOT1 (N272, N227);
nand NAND2 (N273, N257, N209);
nor NOR2 (N274, N271, N207);
buf BUF1 (N275, N274);
or OR4 (N276, N269, N181, N21, N52);
buf BUF1 (N277, N273);
nor NOR2 (N278, N268, N102);
and AND3 (N279, N259, N179, N197);
buf BUF1 (N280, N272);
or OR3 (N281, N267, N76, N127);
nand NAND3 (N282, N278, N63, N56);
nand NAND4 (N283, N253, N248, N143, N273);
or OR2 (N284, N283, N188);
nand NAND4 (N285, N275, N99, N178, N140);
buf BUF1 (N286, N282);
nand NAND2 (N287, N263, N247);
xor XOR2 (N288, N277, N42);
xor XOR2 (N289, N284, N260);
buf BUF1 (N290, N279);
nor NOR2 (N291, N285, N83);
or OR3 (N292, N281, N139, N7);
nand NAND3 (N293, N276, N41, N63);
or OR3 (N294, N280, N250, N35);
and AND3 (N295, N286, N260, N30);
buf BUF1 (N296, N292);
or OR3 (N297, N295, N121, N67);
buf BUF1 (N298, N294);
not NOT1 (N299, N296);
and AND3 (N300, N297, N249, N136);
xor XOR2 (N301, N290, N256);
xor XOR2 (N302, N288, N289);
buf BUF1 (N303, N125);
buf BUF1 (N304, N291);
nor NOR3 (N305, N302, N195, N233);
xor XOR2 (N306, N304, N84);
nand NAND2 (N307, N305, N22);
and AND3 (N308, N307, N21, N174);
not NOT1 (N309, N308);
and AND3 (N310, N299, N289, N157);
buf BUF1 (N311, N301);
or OR4 (N312, N306, N205, N259, N101);
or OR4 (N313, N287, N248, N269, N194);
buf BUF1 (N314, N312);
and AND3 (N315, N298, N140, N127);
buf BUF1 (N316, N313);
xor XOR2 (N317, N303, N210);
buf BUF1 (N318, N270);
or OR2 (N319, N314, N192);
and AND3 (N320, N316, N197, N25);
nand NAND3 (N321, N315, N135, N66);
xor XOR2 (N322, N311, N156);
xor XOR2 (N323, N319, N292);
and AND4 (N324, N309, N211, N136, N144);
xor XOR2 (N325, N321, N29);
xor XOR2 (N326, N310, N137);
xor XOR2 (N327, N325, N93);
not NOT1 (N328, N317);
not NOT1 (N329, N300);
not NOT1 (N330, N328);
or OR2 (N331, N293, N9);
nor NOR3 (N332, N320, N223, N108);
not NOT1 (N333, N327);
xor XOR2 (N334, N333, N42);
xor XOR2 (N335, N318, N323);
xor XOR2 (N336, N127, N197);
xor XOR2 (N337, N330, N84);
nor NOR4 (N338, N336, N84, N260, N45);
nor NOR3 (N339, N331, N260, N4);
nand NAND4 (N340, N322, N87, N317, N64);
xor XOR2 (N341, N332, N266);
buf BUF1 (N342, N329);
or OR2 (N343, N324, N270);
buf BUF1 (N344, N334);
not NOT1 (N345, N343);
nor NOR3 (N346, N345, N75, N107);
buf BUF1 (N347, N337);
buf BUF1 (N348, N339);
nor NOR4 (N349, N344, N164, N77, N66);
not NOT1 (N350, N347);
buf BUF1 (N351, N346);
nand NAND2 (N352, N351, N52);
xor XOR2 (N353, N348, N13);
and AND3 (N354, N350, N309, N25);
nor NOR4 (N355, N341, N235, N5, N101);
nand NAND4 (N356, N338, N117, N166, N307);
not NOT1 (N357, N354);
not NOT1 (N358, N326);
not NOT1 (N359, N355);
nand NAND2 (N360, N342, N291);
buf BUF1 (N361, N340);
not NOT1 (N362, N356);
nand NAND2 (N363, N353, N42);
nand NAND3 (N364, N361, N195, N363);
and AND2 (N365, N91, N58);
or OR3 (N366, N335, N310, N290);
xor XOR2 (N367, N366, N11);
not NOT1 (N368, N360);
xor XOR2 (N369, N368, N60);
not NOT1 (N370, N358);
nand NAND4 (N371, N352, N296, N250, N40);
and AND4 (N372, N362, N109, N127, N247);
buf BUF1 (N373, N349);
nand NAND3 (N374, N359, N156, N124);
or OR2 (N375, N357, N306);
xor XOR2 (N376, N369, N259);
xor XOR2 (N377, N365, N317);
not NOT1 (N378, N372);
and AND2 (N379, N364, N356);
nand NAND3 (N380, N373, N32, N3);
nand NAND4 (N381, N376, N141, N368, N132);
or OR3 (N382, N370, N157, N204);
or OR4 (N383, N379, N80, N253, N368);
buf BUF1 (N384, N378);
xor XOR2 (N385, N375, N231);
buf BUF1 (N386, N374);
not NOT1 (N387, N386);
and AND3 (N388, N387, N322, N60);
not NOT1 (N389, N384);
nand NAND2 (N390, N382, N171);
and AND4 (N391, N383, N19, N42, N84);
not NOT1 (N392, N381);
nand NAND2 (N393, N380, N146);
or OR4 (N394, N389, N322, N333, N17);
nand NAND4 (N395, N394, N232, N269, N222);
not NOT1 (N396, N391);
buf BUF1 (N397, N371);
or OR4 (N398, N385, N264, N23, N132);
not NOT1 (N399, N393);
xor XOR2 (N400, N395, N268);
xor XOR2 (N401, N388, N215);
or OR4 (N402, N401, N302, N383, N303);
nor NOR3 (N403, N377, N367, N357);
nand NAND2 (N404, N2, N286);
buf BUF1 (N405, N397);
nor NOR2 (N406, N402, N401);
and AND4 (N407, N399, N396, N361, N392);
xor XOR2 (N408, N249, N300);
not NOT1 (N409, N245);
not NOT1 (N410, N390);
and AND3 (N411, N405, N279, N199);
or OR2 (N412, N408, N357);
or OR2 (N413, N404, N29);
xor XOR2 (N414, N413, N413);
nor NOR4 (N415, N406, N350, N381, N380);
not NOT1 (N416, N400);
xor XOR2 (N417, N398, N363);
or OR2 (N418, N417, N247);
not NOT1 (N419, N412);
nand NAND3 (N420, N416, N232, N354);
nand NAND3 (N421, N403, N247, N346);
and AND3 (N422, N418, N112, N409);
buf BUF1 (N423, N327);
xor XOR2 (N424, N422, N257);
xor XOR2 (N425, N415, N263);
nor NOR4 (N426, N423, N248, N110, N104);
buf BUF1 (N427, N411);
and AND3 (N428, N410, N170, N383);
buf BUF1 (N429, N424);
and AND4 (N430, N421, N69, N327, N176);
xor XOR2 (N431, N420, N144);
nand NAND3 (N432, N426, N210, N185);
nand NAND2 (N433, N427, N296);
nor NOR3 (N434, N425, N120, N286);
buf BUF1 (N435, N432);
not NOT1 (N436, N419);
nand NAND3 (N437, N435, N158, N220);
nand NAND3 (N438, N437, N364, N118);
nor NOR3 (N439, N434, N138, N326);
or OR4 (N440, N431, N15, N111, N86);
and AND3 (N441, N439, N266, N156);
not NOT1 (N442, N407);
nand NAND3 (N443, N441, N159, N89);
nand NAND2 (N444, N433, N220);
not NOT1 (N445, N428);
buf BUF1 (N446, N443);
nor NOR2 (N447, N414, N416);
or OR2 (N448, N447, N109);
nor NOR3 (N449, N448, N20, N347);
not NOT1 (N450, N449);
and AND4 (N451, N450, N49, N441, N127);
and AND2 (N452, N445, N406);
xor XOR2 (N453, N446, N138);
and AND2 (N454, N442, N184);
and AND3 (N455, N454, N111, N47);
not NOT1 (N456, N453);
buf BUF1 (N457, N430);
xor XOR2 (N458, N456, N211);
or OR2 (N459, N452, N85);
nor NOR3 (N460, N459, N63, N382);
xor XOR2 (N461, N451, N419);
xor XOR2 (N462, N444, N359);
buf BUF1 (N463, N458);
nand NAND4 (N464, N463, N230, N391, N178);
xor XOR2 (N465, N461, N122);
xor XOR2 (N466, N438, N337);
or OR2 (N467, N429, N399);
xor XOR2 (N468, N460, N355);
and AND3 (N469, N455, N378, N45);
or OR4 (N470, N468, N22, N419, N126);
or OR4 (N471, N466, N235, N66, N96);
buf BUF1 (N472, N470);
buf BUF1 (N473, N467);
nand NAND3 (N474, N465, N230, N57);
or OR3 (N475, N471, N148, N389);
or OR2 (N476, N474, N413);
not NOT1 (N477, N469);
nor NOR2 (N478, N440, N429);
nand NAND3 (N479, N476, N354, N109);
nand NAND2 (N480, N473, N410);
nor NOR4 (N481, N478, N189, N480, N256);
and AND4 (N482, N391, N193, N481, N268);
not NOT1 (N483, N381);
or OR4 (N484, N475, N349, N385, N73);
not NOT1 (N485, N482);
not NOT1 (N486, N436);
nor NOR2 (N487, N472, N119);
and AND3 (N488, N457, N7, N403);
or OR2 (N489, N488, N64);
not NOT1 (N490, N487);
nor NOR2 (N491, N490, N124);
or OR4 (N492, N485, N238, N392, N236);
nand NAND2 (N493, N492, N312);
nor NOR4 (N494, N462, N49, N222, N115);
not NOT1 (N495, N477);
buf BUF1 (N496, N484);
not NOT1 (N497, N489);
not NOT1 (N498, N496);
nor NOR2 (N499, N479, N122);
buf BUF1 (N500, N483);
xor XOR2 (N501, N464, N443);
and AND3 (N502, N501, N223, N333);
xor XOR2 (N503, N486, N375);
nand NAND2 (N504, N497, N174);
nor NOR4 (N505, N495, N192, N16, N77);
nand NAND3 (N506, N500, N109, N343);
or OR3 (N507, N502, N478, N445);
buf BUF1 (N508, N491);
buf BUF1 (N509, N508);
nand NAND2 (N510, N499, N112);
or OR2 (N511, N505, N140);
nand NAND4 (N512, N511, N466, N261, N43);
buf BUF1 (N513, N509);
xor XOR2 (N514, N512, N483);
or OR3 (N515, N514, N510, N181);
not NOT1 (N516, N355);
nor NOR2 (N517, N498, N65);
buf BUF1 (N518, N515);
xor XOR2 (N519, N516, N182);
nor NOR3 (N520, N504, N138, N178);
xor XOR2 (N521, N517, N383);
not NOT1 (N522, N506);
not NOT1 (N523, N507);
nor NOR3 (N524, N494, N92, N355);
or OR3 (N525, N521, N106, N224);
or OR2 (N526, N519, N290);
nand NAND3 (N527, N525, N217, N197);
xor XOR2 (N528, N523, N72);
and AND3 (N529, N518, N512, N226);
nand NAND2 (N530, N524, N459);
or OR3 (N531, N522, N213, N197);
and AND2 (N532, N528, N65);
xor XOR2 (N533, N527, N465);
xor XOR2 (N534, N526, N121);
nor NOR3 (N535, N531, N457, N346);
not NOT1 (N536, N529);
xor XOR2 (N537, N536, N318);
xor XOR2 (N538, N520, N434);
not NOT1 (N539, N513);
nor NOR4 (N540, N532, N510, N405, N140);
buf BUF1 (N541, N530);
and AND3 (N542, N533, N294, N213);
nor NOR4 (N543, N539, N106, N50, N326);
buf BUF1 (N544, N493);
and AND4 (N545, N540, N141, N522, N141);
nand NAND4 (N546, N543, N469, N317, N441);
nor NOR2 (N547, N542, N49);
and AND4 (N548, N541, N336, N267, N277);
or OR2 (N549, N535, N104);
or OR4 (N550, N538, N244, N159, N392);
and AND3 (N551, N547, N86, N158);
nand NAND3 (N552, N534, N94, N441);
not NOT1 (N553, N549);
and AND3 (N554, N537, N377, N418);
not NOT1 (N555, N552);
or OR3 (N556, N548, N223, N536);
nand NAND3 (N557, N556, N289, N149);
buf BUF1 (N558, N503);
and AND4 (N559, N554, N235, N122, N167);
xor XOR2 (N560, N550, N220);
buf BUF1 (N561, N557);
xor XOR2 (N562, N546, N24);
nor NOR4 (N563, N562, N364, N282, N200);
nand NAND4 (N564, N560, N130, N360, N433);
and AND3 (N565, N544, N133, N188);
not NOT1 (N566, N564);
nor NOR4 (N567, N563, N401, N458, N285);
xor XOR2 (N568, N551, N288);
xor XOR2 (N569, N553, N389);
nor NOR3 (N570, N559, N76, N22);
buf BUF1 (N571, N570);
nor NOR3 (N572, N561, N422, N458);
and AND3 (N573, N545, N99, N131);
buf BUF1 (N574, N568);
buf BUF1 (N575, N571);
nor NOR2 (N576, N567, N226);
and AND3 (N577, N565, N117, N279);
nor NOR4 (N578, N576, N449, N182, N349);
not NOT1 (N579, N566);
xor XOR2 (N580, N572, N500);
and AND2 (N581, N578, N565);
xor XOR2 (N582, N555, N114);
buf BUF1 (N583, N575);
xor XOR2 (N584, N573, N388);
xor XOR2 (N585, N577, N134);
not NOT1 (N586, N574);
nand NAND2 (N587, N558, N95);
nand NAND2 (N588, N586, N329);
nor NOR3 (N589, N585, N116, N536);
not NOT1 (N590, N589);
nand NAND2 (N591, N590, N153);
buf BUF1 (N592, N583);
xor XOR2 (N593, N582, N333);
and AND3 (N594, N592, N469, N447);
or OR4 (N595, N588, N142, N325, N125);
buf BUF1 (N596, N579);
or OR4 (N597, N596, N441, N300, N591);
nand NAND3 (N598, N375, N402, N260);
nand NAND3 (N599, N595, N216, N559);
nand NAND4 (N600, N584, N540, N229, N488);
or OR2 (N601, N597, N175);
nor NOR2 (N602, N600, N542);
and AND4 (N603, N598, N451, N333, N336);
not NOT1 (N604, N581);
nor NOR4 (N605, N587, N293, N279, N20);
nand NAND4 (N606, N569, N488, N501, N324);
and AND4 (N607, N604, N507, N592, N134);
xor XOR2 (N608, N601, N131);
not NOT1 (N609, N594);
xor XOR2 (N610, N599, N491);
xor XOR2 (N611, N609, N228);
not NOT1 (N612, N602);
not NOT1 (N613, N603);
or OR4 (N614, N608, N237, N596, N158);
buf BUF1 (N615, N606);
xor XOR2 (N616, N614, N21);
not NOT1 (N617, N615);
nor NOR3 (N618, N605, N359, N312);
or OR4 (N619, N612, N485, N306, N413);
not NOT1 (N620, N619);
and AND3 (N621, N620, N351, N512);
xor XOR2 (N622, N611, N404);
not NOT1 (N623, N613);
nand NAND2 (N624, N580, N106);
nor NOR2 (N625, N610, N493);
nor NOR2 (N626, N593, N319);
buf BUF1 (N627, N618);
and AND4 (N628, N616, N507, N41, N469);
xor XOR2 (N629, N623, N205);
and AND3 (N630, N628, N376, N296);
xor XOR2 (N631, N621, N252);
xor XOR2 (N632, N626, N131);
and AND2 (N633, N617, N484);
nor NOR3 (N634, N607, N483, N184);
nor NOR2 (N635, N622, N102);
and AND4 (N636, N632, N275, N332, N398);
nor NOR2 (N637, N624, N304);
not NOT1 (N638, N637);
buf BUF1 (N639, N629);
and AND3 (N640, N635, N58, N270);
xor XOR2 (N641, N639, N155);
or OR2 (N642, N636, N83);
buf BUF1 (N643, N634);
buf BUF1 (N644, N631);
or OR3 (N645, N627, N389, N308);
nor NOR2 (N646, N638, N235);
and AND2 (N647, N642, N352);
nor NOR3 (N648, N646, N453, N235);
not NOT1 (N649, N633);
and AND2 (N650, N630, N384);
xor XOR2 (N651, N625, N413);
and AND3 (N652, N651, N87, N244);
nand NAND3 (N653, N649, N433, N110);
buf BUF1 (N654, N653);
buf BUF1 (N655, N643);
xor XOR2 (N656, N641, N139);
and AND4 (N657, N652, N450, N280, N624);
or OR4 (N658, N657, N519, N91, N173);
or OR3 (N659, N658, N476, N482);
not NOT1 (N660, N644);
xor XOR2 (N661, N656, N490);
or OR3 (N662, N645, N353, N598);
not NOT1 (N663, N662);
or OR2 (N664, N647, N548);
xor XOR2 (N665, N659, N344);
buf BUF1 (N666, N660);
nand NAND2 (N667, N650, N427);
or OR3 (N668, N648, N395, N79);
nor NOR3 (N669, N655, N441, N55);
nor NOR4 (N670, N640, N356, N210, N639);
nor NOR3 (N671, N667, N403, N135);
nand NAND2 (N672, N661, N548);
nand NAND3 (N673, N664, N170, N557);
xor XOR2 (N674, N663, N663);
or OR2 (N675, N665, N330);
buf BUF1 (N676, N675);
buf BUF1 (N677, N668);
and AND4 (N678, N670, N209, N531, N14);
not NOT1 (N679, N678);
and AND4 (N680, N672, N350, N179, N586);
xor XOR2 (N681, N673, N362);
nand NAND2 (N682, N681, N298);
buf BUF1 (N683, N674);
nor NOR3 (N684, N679, N280, N337);
nand NAND4 (N685, N671, N515, N119, N354);
not NOT1 (N686, N676);
and AND4 (N687, N686, N654, N201, N537);
nand NAND3 (N688, N57, N686, N173);
not NOT1 (N689, N685);
not NOT1 (N690, N689);
or OR2 (N691, N666, N685);
nor NOR2 (N692, N682, N31);
xor XOR2 (N693, N669, N227);
buf BUF1 (N694, N684);
nor NOR4 (N695, N688, N215, N624, N188);
nand NAND4 (N696, N677, N538, N327, N584);
not NOT1 (N697, N691);
nor NOR4 (N698, N697, N275, N361, N555);
nand NAND3 (N699, N698, N79, N594);
and AND4 (N700, N690, N594, N305, N612);
and AND2 (N701, N680, N424);
or OR2 (N702, N699, N167);
or OR2 (N703, N687, N139);
not NOT1 (N704, N701);
nand NAND2 (N705, N693, N507);
or OR4 (N706, N700, N534, N90, N78);
or OR3 (N707, N692, N262, N115);
nor NOR3 (N708, N703, N389, N242);
and AND2 (N709, N683, N57);
not NOT1 (N710, N705);
buf BUF1 (N711, N696);
not NOT1 (N712, N694);
xor XOR2 (N713, N707, N550);
not NOT1 (N714, N709);
nor NOR3 (N715, N704, N322, N473);
nand NAND3 (N716, N695, N584, N112);
nor NOR3 (N717, N713, N10, N516);
nand NAND3 (N718, N715, N341, N598);
nand NAND4 (N719, N711, N448, N625, N322);
nor NOR3 (N720, N717, N632, N573);
nor NOR3 (N721, N718, N625, N706);
nor NOR2 (N722, N345, N493);
nand NAND4 (N723, N708, N513, N600, N240);
not NOT1 (N724, N710);
xor XOR2 (N725, N712, N653);
buf BUF1 (N726, N719);
nor NOR3 (N727, N720, N1, N566);
and AND2 (N728, N716, N203);
xor XOR2 (N729, N722, N642);
xor XOR2 (N730, N729, N303);
nand NAND4 (N731, N725, N320, N516, N637);
and AND2 (N732, N728, N68);
buf BUF1 (N733, N714);
and AND2 (N734, N726, N368);
or OR4 (N735, N702, N501, N217, N352);
buf BUF1 (N736, N724);
and AND3 (N737, N735, N591, N420);
buf BUF1 (N738, N721);
not NOT1 (N739, N732);
nand NAND3 (N740, N727, N568, N695);
not NOT1 (N741, N734);
xor XOR2 (N742, N738, N314);
xor XOR2 (N743, N737, N426);
not NOT1 (N744, N741);
xor XOR2 (N745, N744, N574);
buf BUF1 (N746, N723);
and AND2 (N747, N745, N725);
or OR3 (N748, N742, N462, N547);
buf BUF1 (N749, N731);
xor XOR2 (N750, N739, N579);
xor XOR2 (N751, N736, N736);
or OR4 (N752, N746, N193, N407, N598);
and AND4 (N753, N740, N737, N399, N90);
xor XOR2 (N754, N747, N527);
and AND2 (N755, N730, N749);
xor XOR2 (N756, N20, N131);
or OR2 (N757, N750, N128);
and AND2 (N758, N757, N684);
nor NOR2 (N759, N752, N614);
nor NOR2 (N760, N743, N410);
and AND3 (N761, N756, N114, N247);
buf BUF1 (N762, N748);
xor XOR2 (N763, N755, N390);
nand NAND4 (N764, N759, N394, N271, N92);
not NOT1 (N765, N760);
nand NAND3 (N766, N765, N710, N594);
not NOT1 (N767, N762);
or OR4 (N768, N763, N152, N104, N392);
nand NAND3 (N769, N767, N618, N659);
nor NOR2 (N770, N754, N209);
xor XOR2 (N771, N769, N768);
nand NAND3 (N772, N216, N461, N139);
xor XOR2 (N773, N771, N238);
or OR3 (N774, N733, N436, N628);
and AND4 (N775, N772, N70, N48, N245);
nand NAND4 (N776, N775, N539, N37, N261);
not NOT1 (N777, N753);
buf BUF1 (N778, N758);
xor XOR2 (N779, N766, N235);
nor NOR3 (N780, N774, N460, N367);
nand NAND3 (N781, N764, N669, N282);
or OR4 (N782, N770, N640, N9, N267);
nand NAND3 (N783, N773, N687, N207);
buf BUF1 (N784, N782);
and AND2 (N785, N779, N320);
nand NAND4 (N786, N780, N600, N296, N312);
not NOT1 (N787, N751);
nor NOR2 (N788, N787, N30);
and AND2 (N789, N784, N579);
nor NOR4 (N790, N789, N142, N456, N311);
nor NOR3 (N791, N785, N188, N464);
or OR3 (N792, N761, N381, N382);
nand NAND2 (N793, N777, N784);
xor XOR2 (N794, N781, N778);
and AND2 (N795, N37, N301);
not NOT1 (N796, N788);
nor NOR4 (N797, N786, N436, N51, N35);
buf BUF1 (N798, N791);
nand NAND3 (N799, N798, N204, N729);
nand NAND2 (N800, N783, N147);
or OR2 (N801, N800, N735);
buf BUF1 (N802, N776);
nand NAND4 (N803, N799, N563, N207, N681);
or OR2 (N804, N790, N320);
not NOT1 (N805, N796);
not NOT1 (N806, N805);
not NOT1 (N807, N803);
buf BUF1 (N808, N794);
xor XOR2 (N809, N807, N295);
nor NOR2 (N810, N797, N550);
buf BUF1 (N811, N801);
or OR3 (N812, N795, N459, N604);
and AND3 (N813, N811, N780, N214);
xor XOR2 (N814, N808, N241);
not NOT1 (N815, N792);
xor XOR2 (N816, N793, N586);
nor NOR3 (N817, N813, N266, N612);
buf BUF1 (N818, N815);
buf BUF1 (N819, N817);
not NOT1 (N820, N812);
or OR4 (N821, N819, N663, N50, N541);
nor NOR2 (N822, N816, N12);
or OR2 (N823, N810, N520);
and AND2 (N824, N804, N375);
nand NAND4 (N825, N823, N550, N493, N718);
and AND4 (N826, N814, N153, N674, N229);
and AND2 (N827, N822, N434);
not NOT1 (N828, N821);
not NOT1 (N829, N826);
nor NOR3 (N830, N818, N798, N40);
not NOT1 (N831, N802);
not NOT1 (N832, N828);
nor NOR4 (N833, N809, N319, N648, N714);
nand NAND3 (N834, N832, N190, N104);
not NOT1 (N835, N830);
buf BUF1 (N836, N834);
and AND4 (N837, N824, N60, N423, N68);
nor NOR2 (N838, N820, N738);
xor XOR2 (N839, N825, N511);
nor NOR3 (N840, N838, N784, N58);
or OR3 (N841, N836, N722, N171);
not NOT1 (N842, N806);
buf BUF1 (N843, N839);
xor XOR2 (N844, N831, N792);
not NOT1 (N845, N841);
or OR2 (N846, N833, N113);
buf BUF1 (N847, N835);
nand NAND3 (N848, N846, N843, N390);
nor NOR2 (N849, N624, N249);
nand NAND3 (N850, N849, N830, N221);
nor NOR4 (N851, N827, N534, N102, N444);
and AND4 (N852, N851, N484, N685, N376);
not NOT1 (N853, N837);
and AND4 (N854, N847, N336, N264, N474);
buf BUF1 (N855, N852);
xor XOR2 (N856, N845, N501);
xor XOR2 (N857, N856, N589);
not NOT1 (N858, N844);
xor XOR2 (N859, N854, N615);
nor NOR3 (N860, N840, N724, N842);
or OR2 (N861, N843, N182);
or OR4 (N862, N853, N204, N421, N2);
nor NOR4 (N863, N861, N268, N640, N200);
or OR4 (N864, N857, N414, N407, N540);
not NOT1 (N865, N860);
or OR4 (N866, N863, N365, N89, N444);
or OR2 (N867, N829, N506);
nand NAND3 (N868, N864, N116, N677);
and AND3 (N869, N859, N782, N747);
or OR3 (N870, N858, N383, N106);
not NOT1 (N871, N869);
nand NAND4 (N872, N850, N508, N603, N825);
xor XOR2 (N873, N871, N783);
not NOT1 (N874, N867);
nand NAND3 (N875, N862, N586, N357);
not NOT1 (N876, N874);
and AND4 (N877, N855, N202, N194, N468);
not NOT1 (N878, N865);
nor NOR2 (N879, N868, N844);
not NOT1 (N880, N878);
and AND2 (N881, N876, N640);
buf BUF1 (N882, N872);
xor XOR2 (N883, N870, N356);
buf BUF1 (N884, N877);
not NOT1 (N885, N848);
xor XOR2 (N886, N879, N833);
buf BUF1 (N887, N886);
buf BUF1 (N888, N883);
not NOT1 (N889, N887);
xor XOR2 (N890, N881, N243);
nand NAND3 (N891, N873, N465, N49);
xor XOR2 (N892, N888, N190);
nor NOR2 (N893, N866, N254);
or OR4 (N894, N875, N306, N299, N430);
xor XOR2 (N895, N894, N552);
xor XOR2 (N896, N891, N387);
or OR2 (N897, N896, N126);
buf BUF1 (N898, N880);
nor NOR4 (N899, N885, N680, N508, N843);
nor NOR2 (N900, N899, N607);
not NOT1 (N901, N882);
and AND4 (N902, N895, N236, N351, N676);
buf BUF1 (N903, N900);
nand NAND3 (N904, N884, N203, N500);
nand NAND3 (N905, N893, N852, N351);
or OR4 (N906, N901, N818, N86, N737);
nor NOR3 (N907, N890, N642, N332);
buf BUF1 (N908, N905);
nor NOR2 (N909, N906, N862);
nand NAND3 (N910, N898, N180, N482);
or OR4 (N911, N910, N228, N682, N594);
buf BUF1 (N912, N908);
not NOT1 (N913, N909);
xor XOR2 (N914, N892, N17);
xor XOR2 (N915, N897, N27);
and AND4 (N916, N889, N40, N442, N601);
xor XOR2 (N917, N904, N764);
xor XOR2 (N918, N911, N711);
buf BUF1 (N919, N913);
nor NOR2 (N920, N917, N443);
xor XOR2 (N921, N903, N346);
nand NAND3 (N922, N921, N385, N612);
or OR4 (N923, N920, N788, N458, N813);
and AND4 (N924, N919, N76, N371, N555);
not NOT1 (N925, N914);
buf BUF1 (N926, N907);
or OR3 (N927, N924, N493, N238);
not NOT1 (N928, N927);
nor NOR3 (N929, N915, N1, N578);
buf BUF1 (N930, N923);
xor XOR2 (N931, N902, N50);
nor NOR4 (N932, N928, N79, N590, N245);
buf BUF1 (N933, N929);
xor XOR2 (N934, N925, N159);
and AND2 (N935, N916, N611);
nand NAND4 (N936, N932, N298, N920, N506);
not NOT1 (N937, N930);
not NOT1 (N938, N935);
nor NOR4 (N939, N936, N165, N353, N548);
nand NAND2 (N940, N926, N389);
xor XOR2 (N941, N940, N442);
buf BUF1 (N942, N941);
xor XOR2 (N943, N918, N809);
and AND3 (N944, N937, N323, N785);
buf BUF1 (N945, N934);
nand NAND2 (N946, N912, N176);
or OR4 (N947, N938, N895, N828, N461);
nand NAND2 (N948, N939, N590);
nor NOR2 (N949, N931, N869);
or OR4 (N950, N922, N459, N349, N628);
nor NOR2 (N951, N942, N552);
xor XOR2 (N952, N944, N384);
nor NOR4 (N953, N948, N224, N548, N276);
and AND3 (N954, N943, N50, N161);
buf BUF1 (N955, N946);
and AND3 (N956, N945, N299, N2);
nor NOR2 (N957, N951, N188);
buf BUF1 (N958, N950);
and AND4 (N959, N956, N441, N641, N317);
not NOT1 (N960, N947);
and AND3 (N961, N959, N342, N173);
buf BUF1 (N962, N953);
not NOT1 (N963, N962);
or OR4 (N964, N955, N829, N493, N699);
xor XOR2 (N965, N961, N46);
xor XOR2 (N966, N965, N939);
and AND4 (N967, N966, N487, N454, N518);
or OR4 (N968, N960, N62, N13, N157);
nand NAND3 (N969, N952, N967, N762);
nor NOR2 (N970, N134, N361);
xor XOR2 (N971, N968, N636);
xor XOR2 (N972, N949, N277);
buf BUF1 (N973, N963);
nand NAND3 (N974, N973, N358, N324);
xor XOR2 (N975, N972, N262);
nor NOR4 (N976, N954, N465, N788, N101);
or OR2 (N977, N933, N764);
and AND2 (N978, N977, N699);
or OR2 (N979, N964, N627);
not NOT1 (N980, N958);
xor XOR2 (N981, N970, N83);
or OR2 (N982, N978, N590);
not NOT1 (N983, N974);
nor NOR2 (N984, N976, N28);
and AND2 (N985, N957, N840);
nand NAND3 (N986, N971, N58, N625);
nor NOR3 (N987, N979, N15, N596);
buf BUF1 (N988, N983);
nand NAND2 (N989, N987, N694);
nor NOR2 (N990, N975, N131);
xor XOR2 (N991, N982, N243);
and AND2 (N992, N990, N81);
or OR4 (N993, N991, N174, N486, N818);
or OR2 (N994, N969, N313);
xor XOR2 (N995, N993, N362);
buf BUF1 (N996, N984);
nor NOR3 (N997, N989, N298, N617);
and AND2 (N998, N985, N972);
nor NOR3 (N999, N980, N499, N222);
buf BUF1 (N1000, N992);
and AND4 (N1001, N986, N487, N667, N583);
nor NOR2 (N1002, N994, N845);
or OR4 (N1003, N999, N202, N725, N170);
nor NOR3 (N1004, N998, N191, N609);
buf BUF1 (N1005, N1004);
buf BUF1 (N1006, N1002);
or OR3 (N1007, N1001, N197, N566);
nor NOR3 (N1008, N1003, N310, N989);
not NOT1 (N1009, N1005);
buf BUF1 (N1010, N997);
nor NOR3 (N1011, N1006, N305, N534);
not NOT1 (N1012, N995);
or OR4 (N1013, N1008, N696, N742, N99);
xor XOR2 (N1014, N1010, N159);
xor XOR2 (N1015, N988, N662);
not NOT1 (N1016, N1013);
or OR4 (N1017, N1009, N484, N837, N785);
nand NAND3 (N1018, N1000, N584, N332);
and AND4 (N1019, N1018, N608, N322, N920);
or OR3 (N1020, N1014, N197, N288);
nor NOR2 (N1021, N981, N650);
nor NOR4 (N1022, N1019, N826, N390, N198);
xor XOR2 (N1023, N1022, N563);
not NOT1 (N1024, N1023);
buf BUF1 (N1025, N1015);
and AND3 (N1026, N1020, N157, N412);
not NOT1 (N1027, N1026);
not NOT1 (N1028, N1025);
nand NAND3 (N1029, N1012, N246, N374);
xor XOR2 (N1030, N1029, N994);
buf BUF1 (N1031, N1027);
nor NOR2 (N1032, N1031, N742);
xor XOR2 (N1033, N1007, N304);
nand NAND3 (N1034, N1030, N556, N602);
not NOT1 (N1035, N1011);
nor NOR4 (N1036, N1035, N25, N770, N857);
buf BUF1 (N1037, N1016);
and AND3 (N1038, N1032, N127, N915);
or OR4 (N1039, N1024, N470, N541, N224);
xor XOR2 (N1040, N1021, N549);
nand NAND3 (N1041, N1039, N92, N374);
nand NAND2 (N1042, N1038, N15);
nor NOR2 (N1043, N1028, N537);
and AND4 (N1044, N1017, N997, N666, N531);
nand NAND4 (N1045, N1040, N725, N578, N834);
nand NAND4 (N1046, N1033, N579, N144, N570);
xor XOR2 (N1047, N1044, N338);
not NOT1 (N1048, N1045);
xor XOR2 (N1049, N1034, N787);
and AND3 (N1050, N1043, N265, N508);
nand NAND2 (N1051, N1041, N621);
buf BUF1 (N1052, N996);
not NOT1 (N1053, N1051);
buf BUF1 (N1054, N1047);
buf BUF1 (N1055, N1042);
nand NAND3 (N1056, N1048, N52, N342);
nand NAND2 (N1057, N1052, N617);
nor NOR3 (N1058, N1049, N254, N263);
xor XOR2 (N1059, N1054, N211);
nand NAND2 (N1060, N1058, N225);
buf BUF1 (N1061, N1036);
nand NAND3 (N1062, N1056, N319, N687);
nand NAND3 (N1063, N1053, N876, N249);
or OR4 (N1064, N1063, N902, N981, N150);
buf BUF1 (N1065, N1055);
or OR3 (N1066, N1062, N864, N867);
nand NAND3 (N1067, N1050, N72, N1016);
xor XOR2 (N1068, N1059, N67);
nor NOR4 (N1069, N1037, N806, N822, N466);
or OR4 (N1070, N1068, N170, N1030, N305);
and AND2 (N1071, N1065, N810);
xor XOR2 (N1072, N1060, N699);
or OR3 (N1073, N1071, N351, N19);
not NOT1 (N1074, N1061);
nor NOR3 (N1075, N1070, N990, N127);
nand NAND2 (N1076, N1057, N84);
buf BUF1 (N1077, N1069);
buf BUF1 (N1078, N1073);
and AND4 (N1079, N1078, N1024, N1045, N861);
nor NOR3 (N1080, N1046, N546, N451);
nand NAND2 (N1081, N1080, N71);
xor XOR2 (N1082, N1066, N460);
buf BUF1 (N1083, N1072);
nand NAND2 (N1084, N1079, N317);
nor NOR4 (N1085, N1084, N228, N177, N509);
and AND3 (N1086, N1077, N341, N72);
nand NAND2 (N1087, N1075, N690);
nand NAND3 (N1088, N1074, N491, N1076);
and AND2 (N1089, N743, N544);
nand NAND3 (N1090, N1082, N578, N391);
buf BUF1 (N1091, N1087);
nor NOR4 (N1092, N1083, N802, N323, N983);
not NOT1 (N1093, N1090);
xor XOR2 (N1094, N1088, N705);
and AND3 (N1095, N1086, N722, N675);
xor XOR2 (N1096, N1095, N202);
and AND3 (N1097, N1091, N940, N545);
or OR3 (N1098, N1097, N462, N370);
buf BUF1 (N1099, N1067);
xor XOR2 (N1100, N1094, N355);
xor XOR2 (N1101, N1092, N897);
nor NOR4 (N1102, N1100, N624, N340, N267);
buf BUF1 (N1103, N1096);
nand NAND4 (N1104, N1085, N295, N1025, N947);
or OR3 (N1105, N1093, N707, N873);
and AND2 (N1106, N1098, N924);
nor NOR2 (N1107, N1104, N1074);
not NOT1 (N1108, N1105);
not NOT1 (N1109, N1106);
not NOT1 (N1110, N1108);
nor NOR4 (N1111, N1107, N118, N171, N1090);
or OR2 (N1112, N1109, N561);
nand NAND3 (N1113, N1081, N744, N580);
nor NOR4 (N1114, N1064, N1070, N631, N28);
nand NAND3 (N1115, N1099, N134, N895);
buf BUF1 (N1116, N1089);
xor XOR2 (N1117, N1112, N659);
nor NOR2 (N1118, N1115, N541);
nand NAND4 (N1119, N1118, N473, N431, N1068);
not NOT1 (N1120, N1114);
nor NOR2 (N1121, N1103, N728);
nor NOR2 (N1122, N1116, N943);
nor NOR4 (N1123, N1121, N871, N772, N124);
and AND4 (N1124, N1110, N939, N268, N963);
nor NOR4 (N1125, N1113, N245, N1091, N169);
buf BUF1 (N1126, N1125);
buf BUF1 (N1127, N1111);
xor XOR2 (N1128, N1122, N800);
or OR3 (N1129, N1124, N194, N801);
and AND2 (N1130, N1126, N909);
not NOT1 (N1131, N1128);
or OR3 (N1132, N1102, N828, N389);
nand NAND3 (N1133, N1127, N913, N942);
or OR4 (N1134, N1132, N510, N197, N757);
nor NOR2 (N1135, N1101, N60);
nand NAND2 (N1136, N1120, N380);
xor XOR2 (N1137, N1136, N816);
and AND3 (N1138, N1134, N897, N122);
xor XOR2 (N1139, N1131, N1095);
or OR3 (N1140, N1138, N117, N323);
not NOT1 (N1141, N1130);
buf BUF1 (N1142, N1133);
nand NAND2 (N1143, N1129, N817);
or OR2 (N1144, N1117, N507);
xor XOR2 (N1145, N1119, N1120);
not NOT1 (N1146, N1141);
nor NOR2 (N1147, N1135, N352);
or OR4 (N1148, N1139, N540, N826, N442);
or OR4 (N1149, N1143, N407, N827, N559);
buf BUF1 (N1150, N1148);
or OR2 (N1151, N1150, N768);
not NOT1 (N1152, N1137);
and AND4 (N1153, N1146, N117, N974, N546);
buf BUF1 (N1154, N1147);
not NOT1 (N1155, N1145);
xor XOR2 (N1156, N1123, N742);
nor NOR3 (N1157, N1155, N115, N1094);
and AND4 (N1158, N1144, N1074, N1017, N395);
nor NOR4 (N1159, N1153, N1071, N1020, N596);
and AND2 (N1160, N1152, N279);
xor XOR2 (N1161, N1151, N915);
nor NOR3 (N1162, N1140, N409, N494);
nand NAND2 (N1163, N1158, N865);
nor NOR3 (N1164, N1160, N777, N245);
and AND3 (N1165, N1142, N93, N25);
xor XOR2 (N1166, N1154, N554);
or OR4 (N1167, N1159, N77, N442, N82);
not NOT1 (N1168, N1161);
nor NOR3 (N1169, N1166, N913, N626);
nand NAND2 (N1170, N1169, N888);
nand NAND2 (N1171, N1164, N40);
nor NOR4 (N1172, N1170, N505, N465, N158);
nand NAND3 (N1173, N1163, N53, N362);
not NOT1 (N1174, N1173);
buf BUF1 (N1175, N1157);
and AND2 (N1176, N1171, N686);
buf BUF1 (N1177, N1174);
not NOT1 (N1178, N1165);
nor NOR4 (N1179, N1162, N479, N468, N774);
not NOT1 (N1180, N1176);
buf BUF1 (N1181, N1172);
and AND4 (N1182, N1149, N1114, N1149, N1007);
or OR4 (N1183, N1177, N153, N587, N913);
and AND2 (N1184, N1156, N179);
nor NOR2 (N1185, N1181, N111);
nor NOR2 (N1186, N1180, N562);
not NOT1 (N1187, N1175);
buf BUF1 (N1188, N1187);
and AND4 (N1189, N1188, N13, N278, N768);
nand NAND3 (N1190, N1183, N676, N185);
xor XOR2 (N1191, N1178, N378);
not NOT1 (N1192, N1167);
and AND4 (N1193, N1189, N465, N901, N983);
or OR4 (N1194, N1179, N1078, N11, N797);
and AND3 (N1195, N1168, N721, N388);
not NOT1 (N1196, N1190);
buf BUF1 (N1197, N1196);
and AND3 (N1198, N1193, N15, N454);
buf BUF1 (N1199, N1192);
nand NAND3 (N1200, N1182, N992, N177);
xor XOR2 (N1201, N1197, N1081);
buf BUF1 (N1202, N1185);
not NOT1 (N1203, N1184);
xor XOR2 (N1204, N1194, N751);
and AND2 (N1205, N1203, N1058);
xor XOR2 (N1206, N1198, N338);
nand NAND3 (N1207, N1195, N1175, N1000);
nor NOR2 (N1208, N1199, N729);
or OR3 (N1209, N1207, N1144, N301);
buf BUF1 (N1210, N1209);
nor NOR2 (N1211, N1191, N592);
nand NAND2 (N1212, N1202, N65);
and AND3 (N1213, N1201, N807, N471);
nor NOR3 (N1214, N1205, N429, N337);
not NOT1 (N1215, N1214);
not NOT1 (N1216, N1211);
xor XOR2 (N1217, N1204, N332);
buf BUF1 (N1218, N1213);
and AND2 (N1219, N1208, N816);
buf BUF1 (N1220, N1186);
or OR2 (N1221, N1215, N832);
nor NOR3 (N1222, N1217, N829, N8);
nand NAND4 (N1223, N1220, N1044, N832, N713);
xor XOR2 (N1224, N1210, N124);
or OR3 (N1225, N1206, N459, N561);
or OR2 (N1226, N1223, N134);
xor XOR2 (N1227, N1200, N524);
nor NOR2 (N1228, N1226, N33);
nor NOR3 (N1229, N1227, N1091, N997);
or OR4 (N1230, N1221, N1043, N330, N23);
nor NOR3 (N1231, N1218, N1068, N596);
xor XOR2 (N1232, N1231, N240);
nor NOR2 (N1233, N1229, N54);
nand NAND4 (N1234, N1230, N683, N41, N333);
not NOT1 (N1235, N1219);
xor XOR2 (N1236, N1235, N148);
not NOT1 (N1237, N1233);
nor NOR3 (N1238, N1224, N248, N524);
buf BUF1 (N1239, N1234);
not NOT1 (N1240, N1239);
nand NAND4 (N1241, N1238, N663, N822, N1196);
or OR4 (N1242, N1222, N1026, N775, N1092);
xor XOR2 (N1243, N1241, N603);
xor XOR2 (N1244, N1232, N1194);
not NOT1 (N1245, N1225);
buf BUF1 (N1246, N1216);
xor XOR2 (N1247, N1236, N691);
nor NOR2 (N1248, N1212, N705);
xor XOR2 (N1249, N1243, N603);
nor NOR3 (N1250, N1240, N386, N712);
or OR4 (N1251, N1246, N755, N1093, N907);
not NOT1 (N1252, N1247);
and AND3 (N1253, N1237, N1244, N49);
nor NOR2 (N1254, N589, N483);
nand NAND2 (N1255, N1228, N389);
or OR3 (N1256, N1248, N403, N36);
not NOT1 (N1257, N1251);
xor XOR2 (N1258, N1257, N246);
not NOT1 (N1259, N1258);
or OR4 (N1260, N1259, N826, N421, N1251);
or OR3 (N1261, N1245, N361, N508);
nor NOR2 (N1262, N1256, N498);
nor NOR4 (N1263, N1254, N588, N1209, N1253);
nand NAND2 (N1264, N633, N671);
not NOT1 (N1265, N1260);
or OR4 (N1266, N1242, N307, N737, N834);
nor NOR3 (N1267, N1249, N116, N9);
or OR2 (N1268, N1250, N1);
or OR4 (N1269, N1263, N276, N514, N728);
xor XOR2 (N1270, N1266, N731);
and AND2 (N1271, N1261, N1111);
nand NAND4 (N1272, N1267, N859, N1172, N400);
not NOT1 (N1273, N1262);
xor XOR2 (N1274, N1273, N369);
or OR2 (N1275, N1265, N503);
xor XOR2 (N1276, N1252, N556);
not NOT1 (N1277, N1274);
buf BUF1 (N1278, N1269);
or OR3 (N1279, N1272, N1008, N685);
nor NOR2 (N1280, N1268, N1017);
not NOT1 (N1281, N1255);
or OR2 (N1282, N1278, N558);
nor NOR3 (N1283, N1270, N979, N429);
nand NAND4 (N1284, N1264, N720, N195, N57);
nor NOR4 (N1285, N1279, N213, N260, N64);
or OR4 (N1286, N1280, N429, N788, N315);
xor XOR2 (N1287, N1277, N333);
or OR4 (N1288, N1286, N193, N698, N310);
xor XOR2 (N1289, N1276, N1174);
buf BUF1 (N1290, N1281);
and AND2 (N1291, N1288, N1045);
and AND3 (N1292, N1271, N421, N75);
not NOT1 (N1293, N1292);
and AND3 (N1294, N1283, N10, N1251);
not NOT1 (N1295, N1284);
nand NAND3 (N1296, N1290, N992, N1194);
nor NOR2 (N1297, N1285, N575);
xor XOR2 (N1298, N1296, N44);
xor XOR2 (N1299, N1289, N361);
nor NOR2 (N1300, N1275, N268);
nand NAND4 (N1301, N1294, N669, N255, N1033);
buf BUF1 (N1302, N1301);
nand NAND2 (N1303, N1282, N265);
buf BUF1 (N1304, N1299);
nand NAND2 (N1305, N1300, N1291);
or OR4 (N1306, N923, N1104, N645, N413);
or OR3 (N1307, N1297, N31, N1058);
xor XOR2 (N1308, N1305, N207);
buf BUF1 (N1309, N1306);
xor XOR2 (N1310, N1298, N243);
nand NAND3 (N1311, N1310, N117, N421);
xor XOR2 (N1312, N1293, N1281);
nand NAND2 (N1313, N1307, N930);
xor XOR2 (N1314, N1311, N557);
nand NAND2 (N1315, N1303, N843);
nand NAND4 (N1316, N1314, N415, N372, N146);
not NOT1 (N1317, N1313);
nor NOR4 (N1318, N1317, N999, N399, N1198);
nor NOR2 (N1319, N1304, N1108);
and AND2 (N1320, N1302, N973);
nand NAND2 (N1321, N1287, N545);
xor XOR2 (N1322, N1316, N1310);
nand NAND3 (N1323, N1322, N1148, N933);
and AND2 (N1324, N1308, N1102);
nand NAND4 (N1325, N1312, N1313, N691, N189);
nor NOR3 (N1326, N1321, N713, N201);
not NOT1 (N1327, N1319);
nand NAND3 (N1328, N1325, N421, N179);
buf BUF1 (N1329, N1324);
not NOT1 (N1330, N1327);
or OR3 (N1331, N1326, N303, N287);
buf BUF1 (N1332, N1309);
xor XOR2 (N1333, N1323, N726);
nand NAND3 (N1334, N1331, N975, N1261);
buf BUF1 (N1335, N1332);
xor XOR2 (N1336, N1320, N416);
xor XOR2 (N1337, N1329, N24);
buf BUF1 (N1338, N1333);
buf BUF1 (N1339, N1335);
not NOT1 (N1340, N1330);
nor NOR3 (N1341, N1318, N1038, N673);
nand NAND3 (N1342, N1336, N231, N407);
nor NOR3 (N1343, N1315, N243, N825);
nor NOR2 (N1344, N1334, N329);
nand NAND3 (N1345, N1342, N1070, N720);
and AND4 (N1346, N1341, N1078, N820, N1117);
buf BUF1 (N1347, N1345);
nand NAND2 (N1348, N1328, N518);
nand NAND2 (N1349, N1340, N408);
nand NAND3 (N1350, N1339, N1247, N1073);
and AND2 (N1351, N1295, N72);
xor XOR2 (N1352, N1349, N167);
not NOT1 (N1353, N1352);
not NOT1 (N1354, N1338);
xor XOR2 (N1355, N1344, N958);
not NOT1 (N1356, N1348);
xor XOR2 (N1357, N1337, N849);
xor XOR2 (N1358, N1350, N339);
nand NAND4 (N1359, N1354, N726, N677, N887);
and AND4 (N1360, N1357, N290, N386, N581);
or OR3 (N1361, N1356, N539, N358);
xor XOR2 (N1362, N1358, N645);
nor NOR2 (N1363, N1360, N327);
xor XOR2 (N1364, N1362, N1222);
or OR4 (N1365, N1359, N216, N1339, N1215);
or OR3 (N1366, N1353, N1213, N814);
nand NAND3 (N1367, N1343, N741, N451);
not NOT1 (N1368, N1366);
xor XOR2 (N1369, N1365, N1072);
nor NOR2 (N1370, N1347, N1127);
and AND3 (N1371, N1351, N879, N1251);
or OR4 (N1372, N1371, N149, N871, N445);
buf BUF1 (N1373, N1372);
or OR3 (N1374, N1361, N597, N1316);
nand NAND2 (N1375, N1368, N682);
nand NAND4 (N1376, N1369, N440, N308, N1174);
buf BUF1 (N1377, N1373);
xor XOR2 (N1378, N1364, N676);
and AND3 (N1379, N1374, N1112, N1372);
or OR3 (N1380, N1379, N1025, N693);
buf BUF1 (N1381, N1346);
nor NOR2 (N1382, N1381, N357);
nor NOR2 (N1383, N1380, N1328);
xor XOR2 (N1384, N1367, N68);
or OR2 (N1385, N1370, N1192);
buf BUF1 (N1386, N1383);
not NOT1 (N1387, N1355);
buf BUF1 (N1388, N1378);
xor XOR2 (N1389, N1376, N987);
buf BUF1 (N1390, N1382);
and AND3 (N1391, N1388, N544, N54);
nand NAND4 (N1392, N1390, N752, N931, N1103);
and AND4 (N1393, N1389, N685, N685, N397);
not NOT1 (N1394, N1384);
nand NAND2 (N1395, N1392, N800);
buf BUF1 (N1396, N1387);
nand NAND2 (N1397, N1363, N522);
xor XOR2 (N1398, N1393, N709);
buf BUF1 (N1399, N1375);
nand NAND3 (N1400, N1391, N457, N470);
nor NOR3 (N1401, N1398, N148, N474);
nor NOR4 (N1402, N1377, N849, N58, N1004);
not NOT1 (N1403, N1399);
xor XOR2 (N1404, N1403, N1174);
not NOT1 (N1405, N1401);
not NOT1 (N1406, N1385);
xor XOR2 (N1407, N1397, N852);
and AND4 (N1408, N1394, N858, N1392, N1064);
xor XOR2 (N1409, N1400, N788);
and AND3 (N1410, N1407, N1136, N187);
and AND4 (N1411, N1386, N683, N243, N584);
or OR2 (N1412, N1410, N1389);
not NOT1 (N1413, N1402);
xor XOR2 (N1414, N1395, N390);
xor XOR2 (N1415, N1396, N1263);
not NOT1 (N1416, N1411);
or OR3 (N1417, N1406, N1045, N169);
nor NOR4 (N1418, N1413, N583, N360, N700);
not NOT1 (N1419, N1409);
and AND4 (N1420, N1412, N482, N309, N31);
and AND2 (N1421, N1416, N1220);
or OR2 (N1422, N1415, N808);
or OR4 (N1423, N1421, N598, N338, N1289);
nor NOR3 (N1424, N1417, N547, N1046);
not NOT1 (N1425, N1418);
nor NOR4 (N1426, N1405, N689, N321, N724);
or OR2 (N1427, N1422, N673);
xor XOR2 (N1428, N1426, N837);
not NOT1 (N1429, N1414);
nand NAND3 (N1430, N1428, N775, N393);
not NOT1 (N1431, N1408);
not NOT1 (N1432, N1425);
and AND4 (N1433, N1423, N1109, N162, N766);
nor NOR4 (N1434, N1424, N115, N339, N34);
nand NAND3 (N1435, N1419, N26, N1078);
nand NAND4 (N1436, N1434, N983, N277, N748);
xor XOR2 (N1437, N1436, N1064);
xor XOR2 (N1438, N1427, N335);
and AND2 (N1439, N1438, N717);
xor XOR2 (N1440, N1432, N256);
not NOT1 (N1441, N1430);
nand NAND4 (N1442, N1441, N795, N314, N1235);
buf BUF1 (N1443, N1429);
not NOT1 (N1444, N1420);
xor XOR2 (N1445, N1437, N787);
or OR2 (N1446, N1444, N1032);
or OR4 (N1447, N1433, N556, N585, N1266);
nand NAND3 (N1448, N1431, N1131, N1223);
and AND4 (N1449, N1439, N438, N259, N912);
or OR2 (N1450, N1435, N677);
xor XOR2 (N1451, N1449, N291);
or OR3 (N1452, N1442, N954, N1284);
buf BUF1 (N1453, N1447);
not NOT1 (N1454, N1445);
xor XOR2 (N1455, N1440, N161);
nand NAND4 (N1456, N1454, N915, N1267, N1370);
nand NAND2 (N1457, N1455, N575);
buf BUF1 (N1458, N1443);
nor NOR4 (N1459, N1456, N889, N1076, N175);
buf BUF1 (N1460, N1404);
xor XOR2 (N1461, N1453, N265);
buf BUF1 (N1462, N1458);
and AND3 (N1463, N1452, N932, N334);
not NOT1 (N1464, N1450);
xor XOR2 (N1465, N1462, N1179);
xor XOR2 (N1466, N1457, N1200);
xor XOR2 (N1467, N1464, N1332);
buf BUF1 (N1468, N1463);
not NOT1 (N1469, N1459);
xor XOR2 (N1470, N1460, N892);
buf BUF1 (N1471, N1465);
or OR2 (N1472, N1467, N1249);
or OR3 (N1473, N1470, N1347, N1358);
and AND3 (N1474, N1448, N1179, N107);
and AND2 (N1475, N1446, N1299);
and AND4 (N1476, N1466, N394, N260, N1093);
nor NOR3 (N1477, N1475, N376, N1396);
nand NAND3 (N1478, N1468, N1442, N395);
and AND3 (N1479, N1474, N718, N505);
nand NAND2 (N1480, N1471, N461);
or OR2 (N1481, N1476, N585);
buf BUF1 (N1482, N1473);
buf BUF1 (N1483, N1480);
xor XOR2 (N1484, N1478, N537);
or OR2 (N1485, N1481, N17);
or OR2 (N1486, N1451, N1304);
buf BUF1 (N1487, N1485);
xor XOR2 (N1488, N1469, N213);
nand NAND4 (N1489, N1461, N15, N1176, N183);
not NOT1 (N1490, N1472);
buf BUF1 (N1491, N1483);
nand NAND2 (N1492, N1479, N163);
nand NAND2 (N1493, N1491, N262);
buf BUF1 (N1494, N1484);
not NOT1 (N1495, N1493);
or OR3 (N1496, N1477, N562, N243);
not NOT1 (N1497, N1488);
and AND3 (N1498, N1494, N649, N715);
and AND2 (N1499, N1487, N20);
not NOT1 (N1500, N1499);
xor XOR2 (N1501, N1496, N973);
xor XOR2 (N1502, N1486, N107);
nor NOR4 (N1503, N1495, N1120, N1479, N1440);
nor NOR2 (N1504, N1503, N822);
not NOT1 (N1505, N1502);
buf BUF1 (N1506, N1498);
not NOT1 (N1507, N1482);
nor NOR3 (N1508, N1490, N949, N166);
xor XOR2 (N1509, N1506, N1146);
not NOT1 (N1510, N1489);
xor XOR2 (N1511, N1500, N468);
or OR3 (N1512, N1504, N919, N1273);
and AND4 (N1513, N1508, N799, N1463, N415);
nand NAND4 (N1514, N1510, N17, N958, N1182);
nand NAND3 (N1515, N1509, N625, N1176);
nor NOR4 (N1516, N1497, N1105, N125, N1329);
xor XOR2 (N1517, N1515, N1086);
buf BUF1 (N1518, N1514);
xor XOR2 (N1519, N1511, N68);
xor XOR2 (N1520, N1517, N1327);
nor NOR2 (N1521, N1507, N1198);
nor NOR4 (N1522, N1512, N1024, N950, N250);
or OR2 (N1523, N1520, N750);
or OR3 (N1524, N1519, N486, N1158);
and AND3 (N1525, N1513, N1286, N1270);
nand NAND2 (N1526, N1505, N1434);
and AND4 (N1527, N1523, N181, N987, N778);
or OR3 (N1528, N1518, N295, N1447);
or OR2 (N1529, N1526, N701);
nand NAND4 (N1530, N1521, N541, N1009, N1411);
buf BUF1 (N1531, N1528);
nor NOR2 (N1532, N1531, N1264);
xor XOR2 (N1533, N1516, N1152);
nor NOR3 (N1534, N1492, N1242, N700);
buf BUF1 (N1535, N1522);
nand NAND2 (N1536, N1527, N114);
buf BUF1 (N1537, N1525);
buf BUF1 (N1538, N1532);
xor XOR2 (N1539, N1537, N808);
and AND4 (N1540, N1535, N880, N862, N1530);
buf BUF1 (N1541, N844);
or OR4 (N1542, N1529, N6, N183, N977);
buf BUF1 (N1543, N1542);
buf BUF1 (N1544, N1538);
and AND3 (N1545, N1539, N689, N516);
xor XOR2 (N1546, N1540, N241);
nor NOR3 (N1547, N1545, N1250, N633);
nand NAND3 (N1548, N1547, N433, N828);
xor XOR2 (N1549, N1534, N570);
or OR4 (N1550, N1543, N816, N1131, N1306);
and AND2 (N1551, N1548, N994);
and AND2 (N1552, N1524, N956);
not NOT1 (N1553, N1533);
buf BUF1 (N1554, N1501);
or OR4 (N1555, N1550, N141, N314, N1415);
buf BUF1 (N1556, N1536);
nor NOR3 (N1557, N1556, N1451, N179);
xor XOR2 (N1558, N1555, N646);
not NOT1 (N1559, N1552);
or OR2 (N1560, N1559, N555);
nor NOR2 (N1561, N1549, N1038);
xor XOR2 (N1562, N1541, N378);
nand NAND4 (N1563, N1561, N556, N1540, N334);
nand NAND4 (N1564, N1553, N923, N154, N200);
nand NAND3 (N1565, N1558, N1181, N1477);
or OR3 (N1566, N1551, N750, N1314);
not NOT1 (N1567, N1562);
xor XOR2 (N1568, N1567, N1370);
buf BUF1 (N1569, N1557);
buf BUF1 (N1570, N1554);
and AND4 (N1571, N1564, N958, N1260, N942);
not NOT1 (N1572, N1544);
and AND4 (N1573, N1546, N427, N1285, N451);
nor NOR3 (N1574, N1565, N208, N840);
nor NOR4 (N1575, N1574, N971, N530, N574);
and AND3 (N1576, N1569, N1157, N561);
xor XOR2 (N1577, N1570, N691);
and AND3 (N1578, N1576, N784, N1230);
nand NAND3 (N1579, N1575, N1323, N913);
and AND2 (N1580, N1579, N519);
xor XOR2 (N1581, N1571, N855);
xor XOR2 (N1582, N1560, N1308);
buf BUF1 (N1583, N1573);
not NOT1 (N1584, N1582);
and AND4 (N1585, N1580, N1322, N1446, N90);
and AND2 (N1586, N1568, N772);
buf BUF1 (N1587, N1585);
nor NOR2 (N1588, N1578, N285);
nor NOR4 (N1589, N1588, N1061, N1288, N1105);
buf BUF1 (N1590, N1589);
not NOT1 (N1591, N1586);
buf BUF1 (N1592, N1584);
nand NAND4 (N1593, N1583, N905, N18, N567);
nor NOR4 (N1594, N1590, N1394, N826, N907);
nor NOR2 (N1595, N1566, N293);
and AND2 (N1596, N1595, N701);
or OR4 (N1597, N1563, N403, N321, N709);
xor XOR2 (N1598, N1591, N1353);
or OR4 (N1599, N1598, N78, N1346, N243);
xor XOR2 (N1600, N1577, N1213);
and AND4 (N1601, N1587, N1505, N807, N263);
nor NOR4 (N1602, N1599, N131, N438, N1248);
buf BUF1 (N1603, N1597);
buf BUF1 (N1604, N1593);
or OR2 (N1605, N1592, N1521);
or OR2 (N1606, N1605, N1065);
xor XOR2 (N1607, N1581, N96);
xor XOR2 (N1608, N1602, N1290);
nor NOR2 (N1609, N1572, N318);
xor XOR2 (N1610, N1609, N583);
buf BUF1 (N1611, N1610);
and AND4 (N1612, N1611, N392, N1115, N1098);
buf BUF1 (N1613, N1596);
nand NAND4 (N1614, N1601, N993, N1453, N1114);
nand NAND2 (N1615, N1600, N782);
xor XOR2 (N1616, N1613, N593);
and AND3 (N1617, N1615, N864, N88);
endmodule