// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14;

output N3993,N4006,N4008,N4010,N4003,N4009,N4013,N4011,N4012,N4014;

xor XOR2 (N15, N10, N12);
xor XOR2 (N16, N10, N3);
not NOT1 (N17, N5);
not NOT1 (N18, N1);
or OR3 (N19, N14, N18, N17);
xor XOR2 (N20, N19, N3);
or OR4 (N21, N10, N19, N6, N17);
buf BUF1 (N22, N5);
buf BUF1 (N23, N22);
nor NOR3 (N24, N1, N17, N19);
xor XOR2 (N25, N17, N11);
and AND4 (N26, N19, N8, N24, N16);
nand NAND2 (N27, N6, N15);
and AND3 (N28, N14, N14, N7);
buf BUF1 (N29, N14);
xor XOR2 (N30, N21, N13);
and AND2 (N31, N5, N23);
buf BUF1 (N32, N23);
buf BUF1 (N33, N18);
nand NAND2 (N34, N31, N30);
nor NOR4 (N35, N23, N5, N20, N1);
or OR2 (N36, N18, N15);
or OR3 (N37, N28, N17, N6);
buf BUF1 (N38, N26);
nor NOR2 (N39, N36, N24);
and AND2 (N40, N34, N20);
nand NAND4 (N41, N37, N35, N3, N9);
and AND2 (N42, N18, N34);
not NOT1 (N43, N27);
nand NAND2 (N44, N40, N12);
xor XOR2 (N45, N44, N11);
nand NAND2 (N46, N33, N39);
not NOT1 (N47, N37);
or OR3 (N48, N43, N4, N35);
not NOT1 (N49, N32);
nor NOR2 (N50, N49, N18);
xor XOR2 (N51, N25, N2);
and AND4 (N52, N47, N30, N29, N17);
nor NOR3 (N53, N11, N46, N40);
or OR4 (N54, N23, N46, N25, N14);
and AND2 (N55, N41, N11);
nand NAND4 (N56, N52, N15, N37, N55);
not NOT1 (N57, N16);
and AND3 (N58, N45, N8, N6);
and AND2 (N59, N51, N10);
and AND3 (N60, N59, N53, N8);
buf BUF1 (N61, N36);
buf BUF1 (N62, N54);
not NOT1 (N63, N58);
or OR4 (N64, N50, N33, N35, N21);
xor XOR2 (N65, N57, N53);
and AND2 (N66, N38, N36);
and AND2 (N67, N62, N38);
not NOT1 (N68, N56);
or OR3 (N69, N63, N39, N26);
or OR3 (N70, N42, N30, N6);
or OR2 (N71, N48, N27);
nand NAND2 (N72, N60, N5);
buf BUF1 (N73, N64);
xor XOR2 (N74, N72, N3);
nand NAND4 (N75, N61, N43, N35, N58);
or OR2 (N76, N65, N34);
buf BUF1 (N77, N73);
not NOT1 (N78, N75);
or OR3 (N79, N70, N19, N64);
buf BUF1 (N80, N77);
not NOT1 (N81, N67);
not NOT1 (N82, N79);
not NOT1 (N83, N66);
and AND4 (N84, N76, N8, N12, N65);
buf BUF1 (N85, N71);
not NOT1 (N86, N81);
nand NAND2 (N87, N84, N37);
buf BUF1 (N88, N78);
or OR3 (N89, N87, N72, N39);
and AND3 (N90, N80, N21, N52);
nor NOR2 (N91, N82, N47);
or OR3 (N92, N69, N85, N49);
xor XOR2 (N93, N82, N63);
and AND3 (N94, N92, N36, N2);
or OR2 (N95, N93, N32);
not NOT1 (N96, N95);
nor NOR4 (N97, N90, N87, N23, N9);
nand NAND4 (N98, N83, N42, N95, N46);
nor NOR3 (N99, N74, N29, N98);
nor NOR4 (N100, N36, N59, N44, N50);
or OR2 (N101, N91, N14);
xor XOR2 (N102, N86, N35);
buf BUF1 (N103, N100);
and AND3 (N104, N102, N27, N19);
nor NOR3 (N105, N103, N91, N83);
buf BUF1 (N106, N97);
xor XOR2 (N107, N89, N49);
xor XOR2 (N108, N101, N11);
not NOT1 (N109, N107);
xor XOR2 (N110, N68, N106);
buf BUF1 (N111, N45);
nand NAND3 (N112, N94, N33, N72);
buf BUF1 (N113, N105);
xor XOR2 (N114, N113, N16);
nor NOR3 (N115, N110, N24, N78);
xor XOR2 (N116, N99, N72);
nand NAND2 (N117, N112, N28);
or OR4 (N118, N116, N79, N93, N93);
not NOT1 (N119, N88);
nor NOR4 (N120, N117, N54, N7, N19);
buf BUF1 (N121, N108);
nor NOR4 (N122, N111, N30, N72, N95);
and AND2 (N123, N121, N95);
or OR2 (N124, N109, N36);
nand NAND3 (N125, N118, N24, N123);
nand NAND3 (N126, N7, N44, N46);
or OR4 (N127, N122, N31, N19, N58);
not NOT1 (N128, N119);
and AND4 (N129, N114, N65, N31, N33);
and AND2 (N130, N125, N63);
buf BUF1 (N131, N128);
nand NAND4 (N132, N124, N37, N111, N103);
buf BUF1 (N133, N120);
nor NOR4 (N134, N104, N24, N103, N99);
and AND4 (N135, N115, N45, N41, N49);
or OR4 (N136, N130, N20, N70, N21);
and AND3 (N137, N126, N113, N2);
nand NAND2 (N138, N135, N64);
nand NAND4 (N139, N127, N10, N136, N130);
nor NOR3 (N140, N30, N111, N136);
xor XOR2 (N141, N138, N120);
not NOT1 (N142, N132);
or OR4 (N143, N142, N51, N102, N100);
or OR2 (N144, N134, N104);
xor XOR2 (N145, N137, N113);
nand NAND3 (N146, N139, N70, N111);
xor XOR2 (N147, N146, N33);
nand NAND2 (N148, N96, N108);
xor XOR2 (N149, N144, N30);
or OR4 (N150, N145, N26, N80, N119);
or OR3 (N151, N129, N26, N106);
buf BUF1 (N152, N149);
xor XOR2 (N153, N141, N123);
nand NAND2 (N154, N153, N121);
nor NOR4 (N155, N131, N68, N104, N104);
nor NOR4 (N156, N150, N71, N17, N65);
xor XOR2 (N157, N143, N77);
nor NOR2 (N158, N140, N76);
xor XOR2 (N159, N155, N35);
and AND3 (N160, N152, N153, N107);
or OR2 (N161, N158, N143);
xor XOR2 (N162, N151, N45);
and AND3 (N163, N133, N100, N99);
not NOT1 (N164, N147);
not NOT1 (N165, N157);
and AND3 (N166, N165, N122, N114);
nor NOR2 (N167, N163, N52);
buf BUF1 (N168, N154);
not NOT1 (N169, N166);
xor XOR2 (N170, N160, N63);
and AND2 (N171, N161, N80);
xor XOR2 (N172, N171, N5);
or OR2 (N173, N159, N153);
nand NAND3 (N174, N172, N85, N139);
not NOT1 (N175, N156);
or OR4 (N176, N173, N175, N52, N131);
buf BUF1 (N177, N7);
or OR3 (N178, N164, N58, N128);
or OR2 (N179, N169, N167);
or OR3 (N180, N19, N62, N8);
nor NOR3 (N181, N180, N126, N96);
nand NAND4 (N182, N178, N62, N173, N174);
or OR3 (N183, N125, N134, N97);
buf BUF1 (N184, N162);
nor NOR4 (N185, N179, N126, N8, N168);
xor XOR2 (N186, N113, N17);
nor NOR3 (N187, N182, N44, N73);
and AND3 (N188, N183, N26, N70);
xor XOR2 (N189, N181, N11);
or OR2 (N190, N189, N108);
nor NOR2 (N191, N188, N61);
nor NOR3 (N192, N187, N167, N181);
not NOT1 (N193, N191);
nor NOR2 (N194, N186, N143);
xor XOR2 (N195, N177, N55);
or OR3 (N196, N170, N10, N168);
or OR3 (N197, N184, N160, N1);
nor NOR2 (N198, N176, N12);
or OR3 (N199, N193, N129, N94);
nor NOR3 (N200, N197, N124, N70);
nor NOR3 (N201, N185, N191, N47);
or OR2 (N202, N194, N91);
xor XOR2 (N203, N148, N152);
not NOT1 (N204, N198);
and AND2 (N205, N201, N13);
not NOT1 (N206, N200);
and AND4 (N207, N192, N119, N134, N97);
or OR4 (N208, N207, N103, N151, N106);
xor XOR2 (N209, N203, N11);
not NOT1 (N210, N195);
nand NAND2 (N211, N190, N182);
or OR3 (N212, N209, N34, N169);
nor NOR3 (N213, N211, N15, N139);
and AND2 (N214, N205, N131);
and AND2 (N215, N213, N64);
not NOT1 (N216, N196);
buf BUF1 (N217, N210);
not NOT1 (N218, N202);
xor XOR2 (N219, N204, N96);
and AND2 (N220, N199, N82);
and AND2 (N221, N220, N174);
buf BUF1 (N222, N219);
nor NOR2 (N223, N217, N166);
buf BUF1 (N224, N212);
xor XOR2 (N225, N224, N46);
and AND2 (N226, N225, N20);
not NOT1 (N227, N216);
xor XOR2 (N228, N215, N148);
nor NOR3 (N229, N208, N152, N140);
and AND2 (N230, N221, N106);
or OR3 (N231, N218, N20, N114);
buf BUF1 (N232, N223);
and AND2 (N233, N228, N200);
xor XOR2 (N234, N231, N233);
buf BUF1 (N235, N37);
and AND3 (N236, N214, N27, N22);
not NOT1 (N237, N234);
xor XOR2 (N238, N222, N57);
nor NOR4 (N239, N235, N24, N48, N210);
buf BUF1 (N240, N226);
buf BUF1 (N241, N227);
xor XOR2 (N242, N206, N142);
or OR4 (N243, N238, N98, N146, N186);
nor NOR4 (N244, N242, N147, N11, N190);
nand NAND4 (N245, N243, N216, N118, N76);
not NOT1 (N246, N236);
or OR4 (N247, N240, N185, N170, N160);
not NOT1 (N248, N229);
not NOT1 (N249, N237);
xor XOR2 (N250, N249, N119);
and AND3 (N251, N230, N41, N174);
nand NAND3 (N252, N245, N53, N111);
not NOT1 (N253, N244);
not NOT1 (N254, N247);
buf BUF1 (N255, N253);
or OR3 (N256, N246, N103, N199);
nand NAND3 (N257, N241, N117, N121);
buf BUF1 (N258, N257);
nor NOR2 (N259, N255, N10);
or OR2 (N260, N258, N254);
buf BUF1 (N261, N217);
xor XOR2 (N262, N251, N114);
nor NOR3 (N263, N248, N71, N88);
nand NAND4 (N264, N239, N102, N92, N204);
xor XOR2 (N265, N252, N127);
xor XOR2 (N266, N264, N126);
or OR4 (N267, N263, N175, N28, N52);
buf BUF1 (N268, N256);
and AND4 (N269, N265, N245, N80, N21);
and AND2 (N270, N262, N213);
nor NOR3 (N271, N269, N26, N201);
xor XOR2 (N272, N250, N102);
not NOT1 (N273, N266);
nand NAND4 (N274, N270, N213, N96, N250);
and AND2 (N275, N261, N18);
buf BUF1 (N276, N273);
nand NAND3 (N277, N232, N205, N141);
xor XOR2 (N278, N274, N144);
not NOT1 (N279, N267);
xor XOR2 (N280, N259, N255);
nor NOR3 (N281, N278, N200, N186);
nor NOR2 (N282, N272, N53);
or OR2 (N283, N277, N24);
buf BUF1 (N284, N280);
and AND4 (N285, N283, N162, N84, N93);
nor NOR3 (N286, N285, N246, N105);
not NOT1 (N287, N281);
xor XOR2 (N288, N275, N186);
and AND4 (N289, N284, N211, N42, N124);
not NOT1 (N290, N260);
not NOT1 (N291, N290);
buf BUF1 (N292, N291);
and AND2 (N293, N282, N238);
nor NOR2 (N294, N287, N16);
not NOT1 (N295, N293);
nand NAND4 (N296, N276, N179, N99, N250);
not NOT1 (N297, N268);
nand NAND4 (N298, N297, N73, N80, N236);
and AND2 (N299, N289, N82);
or OR3 (N300, N299, N49, N121);
and AND3 (N301, N271, N103, N72);
nand NAND2 (N302, N288, N66);
nand NAND2 (N303, N292, N87);
nor NOR2 (N304, N294, N4);
and AND3 (N305, N279, N38, N298);
xor XOR2 (N306, N54, N120);
buf BUF1 (N307, N286);
nand NAND4 (N308, N304, N122, N205, N182);
nor NOR2 (N309, N301, N266);
or OR2 (N310, N305, N93);
nor NOR4 (N311, N306, N37, N8, N54);
and AND3 (N312, N310, N212, N152);
or OR4 (N313, N303, N227, N295, N124);
buf BUF1 (N314, N242);
and AND3 (N315, N296, N240, N257);
and AND3 (N316, N307, N91, N61);
nand NAND3 (N317, N311, N30, N13);
or OR3 (N318, N308, N102, N27);
xor XOR2 (N319, N318, N281);
and AND2 (N320, N302, N43);
buf BUF1 (N321, N312);
nand NAND2 (N322, N300, N208);
nand NAND3 (N323, N322, N44, N152);
not NOT1 (N324, N315);
buf BUF1 (N325, N320);
buf BUF1 (N326, N316);
and AND2 (N327, N326, N291);
or OR4 (N328, N314, N169, N320, N180);
or OR2 (N329, N309, N119);
not NOT1 (N330, N328);
nand NAND4 (N331, N313, N54, N290, N316);
xor XOR2 (N332, N330, N24);
buf BUF1 (N333, N331);
not NOT1 (N334, N317);
or OR4 (N335, N329, N294, N135, N105);
nand NAND3 (N336, N335, N128, N285);
or OR3 (N337, N319, N250, N30);
nor NOR3 (N338, N321, N125, N251);
or OR4 (N339, N325, N86, N106, N61);
nand NAND4 (N340, N338, N290, N229, N294);
nand NAND3 (N341, N340, N66, N246);
nor NOR3 (N342, N333, N159, N208);
nor NOR2 (N343, N327, N101);
and AND2 (N344, N341, N228);
not NOT1 (N345, N332);
or OR4 (N346, N344, N124, N62, N237);
nand NAND2 (N347, N346, N170);
buf BUF1 (N348, N336);
or OR4 (N349, N323, N333, N193, N310);
and AND2 (N350, N347, N302);
nand NAND4 (N351, N342, N273, N309, N219);
and AND3 (N352, N349, N232, N86);
nand NAND2 (N353, N334, N168);
and AND2 (N354, N339, N35);
and AND2 (N355, N353, N157);
xor XOR2 (N356, N354, N278);
nor NOR3 (N357, N343, N243, N158);
xor XOR2 (N358, N345, N197);
nor NOR2 (N359, N357, N212);
nand NAND3 (N360, N358, N60, N220);
or OR2 (N361, N337, N112);
or OR4 (N362, N355, N225, N213, N290);
not NOT1 (N363, N360);
and AND2 (N364, N361, N12);
buf BUF1 (N365, N348);
xor XOR2 (N366, N362, N24);
not NOT1 (N367, N364);
nor NOR3 (N368, N356, N334, N148);
nor NOR4 (N369, N366, N112, N245, N28);
and AND4 (N370, N350, N154, N228, N313);
nand NAND4 (N371, N368, N49, N146, N318);
buf BUF1 (N372, N363);
not NOT1 (N373, N370);
buf BUF1 (N374, N371);
or OR4 (N375, N324, N9, N168, N167);
not NOT1 (N376, N365);
nor NOR4 (N377, N375, N208, N284, N300);
and AND2 (N378, N372, N136);
buf BUF1 (N379, N369);
xor XOR2 (N380, N351, N114);
and AND2 (N381, N379, N314);
nand NAND2 (N382, N381, N230);
or OR4 (N383, N374, N266, N97, N382);
nand NAND2 (N384, N271, N195);
and AND3 (N385, N359, N338, N160);
buf BUF1 (N386, N373);
nand NAND3 (N387, N383, N333, N331);
xor XOR2 (N388, N378, N210);
nand NAND2 (N389, N386, N55);
nor NOR4 (N390, N380, N299, N192, N124);
not NOT1 (N391, N377);
not NOT1 (N392, N367);
not NOT1 (N393, N390);
xor XOR2 (N394, N384, N229);
nand NAND4 (N395, N391, N249, N309, N46);
nand NAND4 (N396, N392, N293, N258, N300);
and AND3 (N397, N376, N350, N106);
and AND4 (N398, N352, N173, N73, N253);
and AND3 (N399, N389, N307, N344);
xor XOR2 (N400, N399, N334);
buf BUF1 (N401, N387);
nor NOR4 (N402, N401, N118, N28, N343);
buf BUF1 (N403, N388);
not NOT1 (N404, N403);
nor NOR2 (N405, N393, N228);
and AND2 (N406, N395, N333);
or OR2 (N407, N400, N338);
buf BUF1 (N408, N405);
xor XOR2 (N409, N398, N359);
and AND3 (N410, N402, N239, N20);
buf BUF1 (N411, N404);
not NOT1 (N412, N411);
nor NOR4 (N413, N385, N183, N84, N398);
not NOT1 (N414, N396);
nor NOR2 (N415, N413, N217);
buf BUF1 (N416, N409);
nand NAND2 (N417, N410, N59);
or OR4 (N418, N415, N115, N248, N251);
and AND2 (N419, N414, N278);
nor NOR4 (N420, N397, N116, N294, N159);
buf BUF1 (N421, N394);
and AND3 (N422, N408, N296, N36);
or OR3 (N423, N412, N303, N330);
xor XOR2 (N424, N421, N171);
nand NAND2 (N425, N423, N80);
buf BUF1 (N426, N406);
or OR3 (N427, N419, N201, N417);
and AND4 (N428, N163, N57, N216, N386);
nor NOR3 (N429, N416, N101, N144);
and AND3 (N430, N422, N255, N44);
not NOT1 (N431, N428);
not NOT1 (N432, N420);
xor XOR2 (N433, N424, N29);
nand NAND4 (N434, N426, N40, N220, N375);
or OR2 (N435, N434, N63);
and AND2 (N436, N407, N422);
and AND2 (N437, N436, N307);
buf BUF1 (N438, N418);
xor XOR2 (N439, N435, N285);
or OR4 (N440, N425, N151, N292, N63);
and AND3 (N441, N437, N41, N229);
xor XOR2 (N442, N430, N429);
not NOT1 (N443, N192);
nor NOR2 (N444, N433, N212);
buf BUF1 (N445, N441);
buf BUF1 (N446, N439);
or OR2 (N447, N446, N392);
and AND4 (N448, N432, N436, N309, N32);
or OR4 (N449, N447, N447, N70, N275);
and AND3 (N450, N444, N162, N37);
buf BUF1 (N451, N443);
or OR4 (N452, N450, N186, N25, N325);
not NOT1 (N453, N451);
nor NOR4 (N454, N438, N383, N267, N450);
buf BUF1 (N455, N453);
not NOT1 (N456, N445);
buf BUF1 (N457, N455);
and AND4 (N458, N448, N173, N282, N317);
nor NOR3 (N459, N457, N67, N145);
nand NAND2 (N460, N442, N209);
not NOT1 (N461, N427);
nand NAND2 (N462, N460, N34);
nor NOR4 (N463, N449, N222, N325, N168);
nor NOR2 (N464, N461, N388);
nand NAND2 (N465, N454, N323);
nand NAND2 (N466, N459, N207);
xor XOR2 (N467, N452, N73);
nor NOR3 (N468, N456, N80, N395);
xor XOR2 (N469, N467, N194);
buf BUF1 (N470, N458);
nand NAND4 (N471, N465, N441, N111, N189);
not NOT1 (N472, N431);
nor NOR2 (N473, N466, N359);
buf BUF1 (N474, N463);
or OR4 (N475, N473, N225, N107, N419);
or OR2 (N476, N472, N453);
not NOT1 (N477, N469);
buf BUF1 (N478, N470);
nand NAND3 (N479, N475, N397, N208);
buf BUF1 (N480, N464);
buf BUF1 (N481, N440);
or OR3 (N482, N462, N309, N65);
and AND2 (N483, N478, N227);
not NOT1 (N484, N483);
not NOT1 (N485, N471);
xor XOR2 (N486, N484, N425);
or OR3 (N487, N468, N379, N221);
and AND3 (N488, N486, N82, N219);
xor XOR2 (N489, N477, N374);
or OR2 (N490, N480, N61);
not NOT1 (N491, N481);
buf BUF1 (N492, N488);
nor NOR4 (N493, N489, N140, N465, N143);
buf BUF1 (N494, N482);
xor XOR2 (N495, N487, N303);
or OR2 (N496, N476, N303);
not NOT1 (N497, N485);
buf BUF1 (N498, N495);
and AND3 (N499, N498, N240, N163);
nor NOR2 (N500, N491, N12);
or OR3 (N501, N490, N94, N5);
or OR3 (N502, N500, N58, N44);
nand NAND4 (N503, N497, N424, N12, N66);
not NOT1 (N504, N501);
or OR2 (N505, N504, N436);
and AND4 (N506, N502, N379, N424, N54);
and AND3 (N507, N506, N118, N365);
buf BUF1 (N508, N479);
nand NAND2 (N509, N496, N389);
or OR4 (N510, N493, N274, N267, N414);
or OR4 (N511, N494, N205, N6, N48);
nand NAND3 (N512, N499, N79, N250);
nand NAND2 (N513, N511, N346);
not NOT1 (N514, N512);
or OR4 (N515, N510, N18, N398, N65);
xor XOR2 (N516, N513, N140);
and AND4 (N517, N514, N450, N261, N400);
or OR3 (N518, N505, N310, N56);
xor XOR2 (N519, N517, N420);
xor XOR2 (N520, N507, N404);
or OR3 (N521, N509, N108, N334);
or OR2 (N522, N508, N307);
or OR2 (N523, N521, N304);
nor NOR4 (N524, N492, N277, N73, N290);
nand NAND4 (N525, N523, N281, N174, N18);
buf BUF1 (N526, N518);
nor NOR2 (N527, N522, N410);
not NOT1 (N528, N527);
nand NAND3 (N529, N528, N249, N189);
buf BUF1 (N530, N520);
buf BUF1 (N531, N516);
or OR4 (N532, N515, N240, N33, N209);
not NOT1 (N533, N529);
or OR4 (N534, N474, N340, N216, N384);
and AND4 (N535, N533, N388, N393, N135);
buf BUF1 (N536, N531);
buf BUF1 (N537, N536);
and AND3 (N538, N530, N429, N93);
nor NOR2 (N539, N535, N3);
or OR2 (N540, N526, N358);
and AND4 (N541, N525, N430, N203, N336);
nand NAND4 (N542, N539, N381, N533, N338);
xor XOR2 (N543, N541, N446);
nor NOR3 (N544, N503, N374, N37);
not NOT1 (N545, N544);
buf BUF1 (N546, N543);
nor NOR4 (N547, N546, N308, N449, N408);
buf BUF1 (N548, N545);
xor XOR2 (N549, N532, N355);
not NOT1 (N550, N537);
not NOT1 (N551, N549);
nor NOR4 (N552, N524, N346, N234, N59);
and AND2 (N553, N519, N74);
xor XOR2 (N554, N552, N371);
not NOT1 (N555, N551);
buf BUF1 (N556, N538);
xor XOR2 (N557, N548, N228);
not NOT1 (N558, N553);
xor XOR2 (N559, N547, N135);
or OR4 (N560, N557, N442, N222, N34);
buf BUF1 (N561, N555);
xor XOR2 (N562, N540, N48);
or OR4 (N563, N562, N399, N201, N24);
buf BUF1 (N564, N558);
and AND2 (N565, N563, N345);
buf BUF1 (N566, N542);
not NOT1 (N567, N550);
and AND4 (N568, N560, N9, N393, N521);
or OR2 (N569, N566, N138);
and AND3 (N570, N568, N98, N373);
or OR4 (N571, N569, N147, N566, N320);
not NOT1 (N572, N564);
not NOT1 (N573, N572);
nand NAND4 (N574, N567, N139, N182, N291);
nor NOR4 (N575, N570, N155, N500, N73);
buf BUF1 (N576, N554);
and AND4 (N577, N565, N514, N519, N151);
or OR2 (N578, N575, N30);
and AND2 (N579, N571, N67);
xor XOR2 (N580, N576, N294);
not NOT1 (N581, N578);
nor NOR4 (N582, N581, N191, N394, N321);
not NOT1 (N583, N580);
not NOT1 (N584, N556);
buf BUF1 (N585, N574);
nor NOR4 (N586, N583, N447, N383, N435);
buf BUF1 (N587, N577);
nor NOR4 (N588, N534, N183, N464, N350);
and AND2 (N589, N588, N423);
xor XOR2 (N590, N586, N161);
buf BUF1 (N591, N590);
not NOT1 (N592, N559);
nor NOR2 (N593, N584, N96);
and AND4 (N594, N561, N532, N43, N180);
buf BUF1 (N595, N587);
or OR2 (N596, N591, N396);
nand NAND4 (N597, N585, N255, N148, N167);
buf BUF1 (N598, N582);
nor NOR4 (N599, N593, N86, N234, N326);
buf BUF1 (N600, N592);
buf BUF1 (N601, N594);
nand NAND2 (N602, N573, N75);
not NOT1 (N603, N598);
buf BUF1 (N604, N597);
xor XOR2 (N605, N579, N413);
not NOT1 (N606, N599);
xor XOR2 (N607, N602, N148);
not NOT1 (N608, N600);
and AND4 (N609, N606, N446, N437, N350);
and AND3 (N610, N604, N386, N477);
buf BUF1 (N611, N595);
xor XOR2 (N612, N601, N373);
buf BUF1 (N613, N612);
buf BUF1 (N614, N607);
and AND4 (N615, N610, N579, N240, N591);
not NOT1 (N616, N603);
buf BUF1 (N617, N596);
nor NOR4 (N618, N589, N547, N236, N358);
and AND3 (N619, N613, N469, N128);
and AND4 (N620, N615, N151, N408, N536);
and AND4 (N621, N617, N23, N210, N502);
nor NOR3 (N622, N620, N407, N513);
or OR3 (N623, N605, N337, N341);
or OR3 (N624, N609, N105, N90);
not NOT1 (N625, N623);
nor NOR2 (N626, N619, N558);
or OR2 (N627, N626, N223);
nor NOR4 (N628, N625, N621, N276, N415);
nand NAND3 (N629, N575, N92, N379);
xor XOR2 (N630, N624, N175);
buf BUF1 (N631, N629);
xor XOR2 (N632, N630, N247);
not NOT1 (N633, N631);
and AND2 (N634, N618, N576);
or OR2 (N635, N608, N416);
and AND2 (N636, N633, N49);
or OR4 (N637, N635, N461, N588, N403);
or OR3 (N638, N614, N128, N398);
and AND4 (N639, N638, N275, N593, N429);
nor NOR4 (N640, N628, N638, N559, N246);
nor NOR4 (N641, N634, N617, N495, N432);
nor NOR4 (N642, N637, N233, N467, N545);
nand NAND4 (N643, N636, N514, N577, N55);
and AND4 (N644, N611, N611, N150, N110);
nand NAND2 (N645, N641, N14);
buf BUF1 (N646, N632);
nand NAND4 (N647, N639, N185, N216, N280);
not NOT1 (N648, N622);
and AND2 (N649, N640, N63);
and AND2 (N650, N642, N343);
and AND3 (N651, N627, N313, N365);
and AND4 (N652, N649, N40, N334, N202);
buf BUF1 (N653, N646);
buf BUF1 (N654, N651);
xor XOR2 (N655, N653, N522);
buf BUF1 (N656, N650);
not NOT1 (N657, N644);
buf BUF1 (N658, N655);
xor XOR2 (N659, N657, N252);
nand NAND3 (N660, N658, N121, N55);
nand NAND4 (N661, N643, N433, N585, N219);
nor NOR2 (N662, N647, N284);
nor NOR3 (N663, N654, N29, N552);
nand NAND3 (N664, N662, N423, N235);
not NOT1 (N665, N652);
not NOT1 (N666, N659);
buf BUF1 (N667, N660);
not NOT1 (N668, N645);
not NOT1 (N669, N668);
nor NOR3 (N670, N616, N170, N296);
and AND2 (N671, N648, N210);
nor NOR2 (N672, N666, N593);
nor NOR3 (N673, N667, N2, N581);
or OR3 (N674, N656, N649, N135);
or OR2 (N675, N672, N328);
and AND3 (N676, N675, N73, N228);
buf BUF1 (N677, N671);
not NOT1 (N678, N663);
nand NAND2 (N679, N673, N284);
nand NAND4 (N680, N669, N526, N436, N561);
and AND3 (N681, N670, N661, N378);
and AND4 (N682, N335, N393, N311, N139);
or OR2 (N683, N677, N235);
or OR3 (N684, N676, N618, N213);
buf BUF1 (N685, N684);
and AND2 (N686, N679, N17);
nand NAND4 (N687, N664, N29, N424, N352);
nand NAND2 (N688, N682, N620);
buf BUF1 (N689, N680);
and AND4 (N690, N681, N499, N265, N587);
nand NAND3 (N691, N690, N225, N426);
nand NAND4 (N692, N689, N475, N292, N423);
buf BUF1 (N693, N686);
or OR2 (N694, N678, N117);
and AND4 (N695, N674, N126, N572, N593);
not NOT1 (N696, N665);
nor NOR3 (N697, N692, N684, N142);
and AND2 (N698, N688, N173);
and AND3 (N699, N695, N80, N676);
nand NAND4 (N700, N697, N593, N326, N590);
nor NOR4 (N701, N685, N249, N37, N434);
not NOT1 (N702, N698);
xor XOR2 (N703, N694, N183);
and AND2 (N704, N687, N242);
or OR4 (N705, N704, N123, N303, N314);
not NOT1 (N706, N700);
nand NAND2 (N707, N702, N557);
and AND3 (N708, N701, N222, N327);
xor XOR2 (N709, N696, N444);
nand NAND4 (N710, N683, N189, N139, N493);
xor XOR2 (N711, N706, N646);
nor NOR3 (N712, N703, N61, N582);
nand NAND3 (N713, N691, N242, N706);
not NOT1 (N714, N707);
xor XOR2 (N715, N708, N51);
buf BUF1 (N716, N715);
not NOT1 (N717, N693);
xor XOR2 (N718, N705, N211);
buf BUF1 (N719, N711);
not NOT1 (N720, N719);
xor XOR2 (N721, N709, N323);
or OR4 (N722, N710, N241, N173, N195);
xor XOR2 (N723, N722, N20);
nand NAND4 (N724, N699, N118, N465, N246);
and AND4 (N725, N712, N53, N266, N155);
xor XOR2 (N726, N714, N725);
and AND2 (N727, N203, N219);
nand NAND3 (N728, N718, N291, N527);
buf BUF1 (N729, N728);
buf BUF1 (N730, N727);
and AND4 (N731, N717, N35, N147, N690);
and AND3 (N732, N721, N570, N281);
not NOT1 (N733, N731);
xor XOR2 (N734, N726, N207);
and AND4 (N735, N732, N108, N164, N600);
nor NOR4 (N736, N724, N214, N414, N618);
nand NAND4 (N737, N729, N406, N7, N333);
buf BUF1 (N738, N716);
nor NOR2 (N739, N738, N694);
nand NAND4 (N740, N737, N595, N35, N205);
xor XOR2 (N741, N720, N416);
nor NOR2 (N742, N733, N70);
nand NAND3 (N743, N742, N163, N548);
and AND2 (N744, N713, N208);
and AND4 (N745, N740, N499, N16, N676);
nand NAND3 (N746, N736, N5, N150);
buf BUF1 (N747, N730);
xor XOR2 (N748, N723, N237);
and AND4 (N749, N741, N352, N407, N177);
buf BUF1 (N750, N743);
xor XOR2 (N751, N734, N298);
buf BUF1 (N752, N739);
or OR4 (N753, N746, N509, N712, N593);
nor NOR3 (N754, N735, N606, N717);
or OR3 (N755, N754, N81, N473);
nor NOR2 (N756, N751, N560);
not NOT1 (N757, N752);
and AND4 (N758, N748, N502, N541, N141);
nor NOR2 (N759, N749, N166);
xor XOR2 (N760, N756, N535);
nand NAND4 (N761, N744, N689, N28, N486);
buf BUF1 (N762, N760);
not NOT1 (N763, N759);
nor NOR3 (N764, N758, N353, N581);
xor XOR2 (N765, N753, N549);
not NOT1 (N766, N763);
nand NAND3 (N767, N762, N390, N650);
nor NOR4 (N768, N747, N401, N134, N745);
buf BUF1 (N769, N617);
nand NAND4 (N770, N766, N621, N369, N54);
nand NAND4 (N771, N767, N92, N706, N438);
and AND3 (N772, N764, N723, N640);
nand NAND3 (N773, N757, N635, N270);
and AND4 (N774, N772, N58, N556, N19);
nand NAND3 (N775, N750, N256, N446);
xor XOR2 (N776, N768, N247);
nor NOR3 (N777, N775, N375, N78);
or OR4 (N778, N771, N654, N586, N219);
nor NOR3 (N779, N777, N163, N88);
nand NAND4 (N780, N779, N662, N385, N152);
nor NOR2 (N781, N776, N476);
nor NOR3 (N782, N755, N639, N189);
nand NAND3 (N783, N769, N119, N1);
nand NAND3 (N784, N782, N154, N562);
and AND3 (N785, N770, N699, N445);
not NOT1 (N786, N781);
nor NOR3 (N787, N765, N555, N621);
buf BUF1 (N788, N761);
buf BUF1 (N789, N785);
buf BUF1 (N790, N789);
buf BUF1 (N791, N783);
nand NAND2 (N792, N791, N313);
buf BUF1 (N793, N774);
or OR3 (N794, N788, N108, N81);
buf BUF1 (N795, N794);
xor XOR2 (N796, N778, N205);
xor XOR2 (N797, N787, N176);
buf BUF1 (N798, N795);
nor NOR3 (N799, N784, N234, N478);
buf BUF1 (N800, N780);
not NOT1 (N801, N773);
and AND4 (N802, N799, N783, N224, N90);
buf BUF1 (N803, N796);
not NOT1 (N804, N803);
not NOT1 (N805, N797);
not NOT1 (N806, N800);
nand NAND3 (N807, N806, N258, N323);
nand NAND4 (N808, N805, N355, N391, N664);
buf BUF1 (N809, N790);
not NOT1 (N810, N792);
nand NAND4 (N811, N808, N556, N656, N89);
nor NOR2 (N812, N811, N390);
buf BUF1 (N813, N804);
not NOT1 (N814, N810);
nand NAND3 (N815, N801, N213, N11);
xor XOR2 (N816, N798, N400);
or OR2 (N817, N812, N416);
and AND3 (N818, N815, N613, N790);
nor NOR3 (N819, N814, N523, N736);
nand NAND3 (N820, N807, N629, N798);
and AND4 (N821, N820, N808, N152, N489);
or OR3 (N822, N793, N270, N695);
nor NOR4 (N823, N816, N81, N332, N458);
and AND3 (N824, N809, N89, N149);
buf BUF1 (N825, N813);
nor NOR4 (N826, N818, N211, N655, N531);
not NOT1 (N827, N821);
buf BUF1 (N828, N826);
or OR2 (N829, N824, N54);
buf BUF1 (N830, N825);
or OR3 (N831, N786, N115, N332);
buf BUF1 (N832, N829);
nand NAND3 (N833, N831, N41, N634);
nand NAND3 (N834, N832, N620, N48);
or OR3 (N835, N822, N723, N715);
nor NOR3 (N836, N823, N699, N53);
xor XOR2 (N837, N833, N833);
xor XOR2 (N838, N802, N337);
xor XOR2 (N839, N827, N619);
buf BUF1 (N840, N828);
xor XOR2 (N841, N839, N744);
and AND4 (N842, N837, N305, N706, N709);
and AND4 (N843, N817, N149, N519, N326);
nand NAND2 (N844, N830, N581);
nor NOR3 (N845, N843, N21, N763);
and AND2 (N846, N841, N309);
or OR4 (N847, N835, N494, N732, N284);
nor NOR2 (N848, N842, N706);
nand NAND2 (N849, N844, N492);
or OR3 (N850, N849, N69, N165);
xor XOR2 (N851, N848, N814);
not NOT1 (N852, N851);
nor NOR4 (N853, N845, N846, N836, N687);
buf BUF1 (N854, N429);
and AND4 (N855, N51, N674, N79, N848);
xor XOR2 (N856, N855, N729);
buf BUF1 (N857, N847);
and AND4 (N858, N857, N271, N508, N319);
nor NOR4 (N859, N854, N234, N489, N367);
not NOT1 (N860, N859);
xor XOR2 (N861, N838, N204);
or OR3 (N862, N850, N75, N769);
and AND3 (N863, N834, N52, N458);
nor NOR2 (N864, N819, N107);
or OR3 (N865, N860, N347, N388);
buf BUF1 (N866, N840);
and AND4 (N867, N864, N477, N574, N529);
or OR4 (N868, N856, N449, N633, N746);
and AND4 (N869, N865, N69, N223, N68);
xor XOR2 (N870, N866, N379);
buf BUF1 (N871, N861);
buf BUF1 (N872, N853);
or OR3 (N873, N867, N476, N471);
buf BUF1 (N874, N868);
nand NAND3 (N875, N869, N46, N602);
or OR2 (N876, N862, N52);
buf BUF1 (N877, N863);
nand NAND2 (N878, N873, N724);
and AND4 (N879, N852, N679, N623, N813);
or OR4 (N880, N871, N704, N204, N457);
or OR4 (N881, N877, N861, N329, N127);
or OR2 (N882, N858, N562);
nand NAND2 (N883, N870, N585);
buf BUF1 (N884, N876);
xor XOR2 (N885, N880, N433);
buf BUF1 (N886, N879);
nor NOR3 (N887, N885, N782, N60);
or OR3 (N888, N874, N195, N4);
buf BUF1 (N889, N884);
nand NAND2 (N890, N882, N819);
and AND2 (N891, N875, N309);
and AND3 (N892, N872, N847, N253);
xor XOR2 (N893, N883, N614);
and AND4 (N894, N881, N75, N869, N836);
xor XOR2 (N895, N894, N727);
buf BUF1 (N896, N892);
nor NOR3 (N897, N893, N216, N390);
buf BUF1 (N898, N886);
xor XOR2 (N899, N891, N846);
nand NAND4 (N900, N895, N511, N520, N186);
nor NOR4 (N901, N896, N549, N878, N51);
xor XOR2 (N902, N45, N465);
and AND4 (N903, N889, N144, N122, N275);
and AND2 (N904, N903, N620);
or OR3 (N905, N899, N564, N356);
not NOT1 (N906, N887);
buf BUF1 (N907, N902);
and AND2 (N908, N897, N491);
and AND2 (N909, N906, N413);
nor NOR4 (N910, N904, N195, N674, N272);
nand NAND3 (N911, N909, N157, N844);
or OR2 (N912, N898, N723);
nand NAND3 (N913, N908, N661, N786);
and AND3 (N914, N912, N675, N153);
or OR4 (N915, N900, N333, N285, N801);
and AND2 (N916, N888, N54);
buf BUF1 (N917, N911);
and AND3 (N918, N915, N717, N703);
or OR3 (N919, N901, N171, N519);
not NOT1 (N920, N919);
or OR2 (N921, N913, N50);
nand NAND2 (N922, N905, N406);
nor NOR3 (N923, N920, N478, N223);
nor NOR3 (N924, N923, N516, N139);
and AND4 (N925, N914, N494, N267, N388);
nor NOR4 (N926, N916, N483, N888, N907);
or OR4 (N927, N595, N173, N568, N570);
not NOT1 (N928, N926);
and AND4 (N929, N924, N516, N171, N404);
and AND3 (N930, N910, N845, N152);
and AND3 (N931, N928, N526, N559);
or OR3 (N932, N929, N261, N786);
and AND2 (N933, N918, N109);
nor NOR4 (N934, N930, N103, N725, N108);
or OR4 (N935, N927, N541, N934, N762);
nor NOR2 (N936, N261, N22);
nor NOR3 (N937, N917, N229, N531);
or OR3 (N938, N937, N56, N583);
nand NAND2 (N939, N921, N502);
nor NOR3 (N940, N932, N639, N204);
and AND2 (N941, N890, N786);
or OR4 (N942, N933, N633, N928, N698);
or OR4 (N943, N931, N97, N286, N451);
xor XOR2 (N944, N925, N675);
nand NAND4 (N945, N922, N348, N674, N268);
nand NAND2 (N946, N942, N686);
nand NAND2 (N947, N938, N767);
or OR2 (N948, N936, N187);
and AND4 (N949, N940, N632, N244, N550);
not NOT1 (N950, N948);
or OR3 (N951, N944, N764, N288);
or OR2 (N952, N949, N228);
or OR2 (N953, N946, N394);
nand NAND3 (N954, N939, N649, N815);
xor XOR2 (N955, N953, N658);
buf BUF1 (N956, N951);
nor NOR2 (N957, N941, N464);
buf BUF1 (N958, N947);
nand NAND2 (N959, N943, N488);
buf BUF1 (N960, N935);
or OR2 (N961, N950, N701);
nor NOR4 (N962, N957, N907, N406, N702);
nand NAND2 (N963, N955, N180);
or OR3 (N964, N956, N453, N287);
buf BUF1 (N965, N961);
nor NOR2 (N966, N945, N488);
not NOT1 (N967, N954);
or OR4 (N968, N965, N515, N923, N494);
nor NOR3 (N969, N967, N556, N657);
or OR3 (N970, N966, N191, N139);
xor XOR2 (N971, N960, N42);
xor XOR2 (N972, N963, N684);
and AND4 (N973, N968, N940, N523, N420);
nor NOR4 (N974, N971, N681, N239, N511);
nor NOR2 (N975, N964, N638);
and AND2 (N976, N952, N328);
buf BUF1 (N977, N970);
or OR3 (N978, N976, N192, N956);
xor XOR2 (N979, N973, N486);
and AND3 (N980, N969, N34, N696);
nor NOR2 (N981, N978, N464);
and AND2 (N982, N980, N103);
nor NOR3 (N983, N977, N571, N382);
nand NAND3 (N984, N979, N40, N713);
xor XOR2 (N985, N962, N145);
nor NOR2 (N986, N975, N11);
or OR3 (N987, N983, N369, N850);
and AND2 (N988, N974, N288);
or OR4 (N989, N985, N441, N564, N93);
and AND2 (N990, N982, N701);
xor XOR2 (N991, N989, N990);
nand NAND3 (N992, N916, N262, N919);
not NOT1 (N993, N986);
nor NOR4 (N994, N988, N149, N613, N482);
nor NOR3 (N995, N994, N61, N806);
buf BUF1 (N996, N992);
nor NOR4 (N997, N991, N767, N833, N458);
not NOT1 (N998, N993);
xor XOR2 (N999, N959, N721);
or OR3 (N1000, N984, N299, N89);
buf BUF1 (N1001, N998);
xor XOR2 (N1002, N987, N432);
and AND4 (N1003, N999, N751, N251, N127);
or OR4 (N1004, N1001, N378, N957, N570);
buf BUF1 (N1005, N1000);
nand NAND3 (N1006, N981, N360, N674);
nand NAND2 (N1007, N1003, N342);
nand NAND4 (N1008, N1002, N945, N152, N678);
and AND4 (N1009, N1007, N625, N179, N572);
buf BUF1 (N1010, N1006);
xor XOR2 (N1011, N995, N658);
buf BUF1 (N1012, N958);
nor NOR4 (N1013, N1004, N806, N565, N385);
not NOT1 (N1014, N1008);
not NOT1 (N1015, N1005);
xor XOR2 (N1016, N1015, N167);
or OR4 (N1017, N1011, N17, N770, N910);
or OR3 (N1018, N1017, N511, N780);
nand NAND3 (N1019, N1010, N322, N965);
not NOT1 (N1020, N1013);
not NOT1 (N1021, N1016);
nand NAND3 (N1022, N1009, N304, N299);
nor NOR2 (N1023, N1019, N419);
xor XOR2 (N1024, N997, N815);
buf BUF1 (N1025, N1024);
xor XOR2 (N1026, N1012, N45);
not NOT1 (N1027, N1021);
and AND3 (N1028, N1023, N556, N880);
or OR3 (N1029, N1020, N41, N551);
xor XOR2 (N1030, N1026, N635);
buf BUF1 (N1031, N1030);
nor NOR2 (N1032, N1027, N392);
not NOT1 (N1033, N1025);
nor NOR3 (N1034, N1029, N687, N561);
nand NAND4 (N1035, N1034, N924, N391, N886);
or OR2 (N1036, N1032, N808);
nor NOR4 (N1037, N996, N270, N410, N471);
buf BUF1 (N1038, N1018);
xor XOR2 (N1039, N1033, N43);
and AND2 (N1040, N1014, N838);
xor XOR2 (N1041, N1031, N602);
xor XOR2 (N1042, N1040, N265);
nor NOR2 (N1043, N1038, N916);
nor NOR4 (N1044, N1041, N783, N780, N257);
not NOT1 (N1045, N1042);
nand NAND4 (N1046, N1022, N35, N210, N702);
nor NOR4 (N1047, N1043, N449, N535, N910);
or OR2 (N1048, N1047, N958);
and AND3 (N1049, N1037, N662, N731);
xor XOR2 (N1050, N1028, N372);
nor NOR2 (N1051, N1049, N670);
xor XOR2 (N1052, N1051, N268);
and AND2 (N1053, N1045, N645);
nand NAND2 (N1054, N1039, N610);
not NOT1 (N1055, N1052);
not NOT1 (N1056, N1044);
nand NAND2 (N1057, N1056, N173);
nand NAND3 (N1058, N1050, N249, N264);
or OR3 (N1059, N1048, N893, N145);
and AND4 (N1060, N1035, N634, N895, N637);
or OR2 (N1061, N1036, N68);
not NOT1 (N1062, N1061);
nor NOR3 (N1063, N1058, N873, N607);
not NOT1 (N1064, N1057);
buf BUF1 (N1065, N1046);
nand NAND2 (N1066, N1064, N813);
nand NAND4 (N1067, N1053, N822, N52, N756);
nand NAND3 (N1068, N1062, N432, N814);
buf BUF1 (N1069, N1054);
and AND4 (N1070, N1069, N997, N926, N245);
xor XOR2 (N1071, N1055, N937);
not NOT1 (N1072, N1071);
or OR3 (N1073, N1068, N157, N852);
buf BUF1 (N1074, N972);
and AND2 (N1075, N1060, N983);
and AND3 (N1076, N1059, N147, N460);
nand NAND3 (N1077, N1075, N502, N357);
not NOT1 (N1078, N1070);
not NOT1 (N1079, N1065);
not NOT1 (N1080, N1079);
nand NAND2 (N1081, N1066, N113);
or OR3 (N1082, N1074, N935, N173);
xor XOR2 (N1083, N1080, N534);
or OR3 (N1084, N1072, N629, N51);
nand NAND3 (N1085, N1082, N484, N437);
not NOT1 (N1086, N1085);
not NOT1 (N1087, N1081);
nand NAND2 (N1088, N1086, N921);
and AND4 (N1089, N1073, N834, N874, N718);
and AND4 (N1090, N1067, N329, N751, N856);
and AND2 (N1091, N1090, N863);
and AND4 (N1092, N1087, N838, N595, N344);
not NOT1 (N1093, N1063);
xor XOR2 (N1094, N1076, N1016);
and AND3 (N1095, N1077, N354, N307);
buf BUF1 (N1096, N1089);
buf BUF1 (N1097, N1091);
nand NAND4 (N1098, N1093, N1078, N765, N835);
or OR2 (N1099, N846, N156);
nand NAND2 (N1100, N1084, N988);
or OR2 (N1101, N1099, N994);
and AND2 (N1102, N1083, N420);
not NOT1 (N1103, N1098);
xor XOR2 (N1104, N1100, N878);
nand NAND2 (N1105, N1103, N782);
not NOT1 (N1106, N1096);
not NOT1 (N1107, N1102);
buf BUF1 (N1108, N1094);
nor NOR2 (N1109, N1108, N826);
xor XOR2 (N1110, N1106, N304);
nand NAND2 (N1111, N1097, N1041);
xor XOR2 (N1112, N1092, N444);
nor NOR4 (N1113, N1110, N465, N558, N674);
not NOT1 (N1114, N1113);
xor XOR2 (N1115, N1114, N945);
xor XOR2 (N1116, N1104, N823);
or OR2 (N1117, N1116, N223);
nand NAND4 (N1118, N1107, N31, N379, N492);
or OR3 (N1119, N1115, N1105, N864);
nor NOR2 (N1120, N324, N115);
xor XOR2 (N1121, N1101, N65);
nand NAND3 (N1122, N1118, N1036, N869);
buf BUF1 (N1123, N1117);
nor NOR3 (N1124, N1120, N135, N27);
not NOT1 (N1125, N1088);
nor NOR4 (N1126, N1121, N795, N490, N364);
or OR2 (N1127, N1109, N544);
nor NOR2 (N1128, N1095, N911);
not NOT1 (N1129, N1123);
nand NAND3 (N1130, N1126, N792, N901);
and AND3 (N1131, N1130, N429, N787);
nor NOR2 (N1132, N1129, N1013);
xor XOR2 (N1133, N1131, N959);
buf BUF1 (N1134, N1125);
not NOT1 (N1135, N1119);
nand NAND2 (N1136, N1122, N228);
buf BUF1 (N1137, N1133);
nand NAND2 (N1138, N1134, N565);
and AND2 (N1139, N1135, N206);
nand NAND3 (N1140, N1139, N558, N573);
buf BUF1 (N1141, N1127);
buf BUF1 (N1142, N1140);
buf BUF1 (N1143, N1136);
or OR3 (N1144, N1124, N1013, N261);
buf BUF1 (N1145, N1144);
not NOT1 (N1146, N1138);
xor XOR2 (N1147, N1128, N1118);
or OR2 (N1148, N1141, N849);
nor NOR2 (N1149, N1148, N831);
nand NAND4 (N1150, N1145, N396, N1050, N495);
buf BUF1 (N1151, N1112);
or OR3 (N1152, N1147, N773, N430);
buf BUF1 (N1153, N1111);
xor XOR2 (N1154, N1142, N18);
or OR4 (N1155, N1150, N814, N823, N895);
nor NOR4 (N1156, N1152, N864, N1088, N757);
buf BUF1 (N1157, N1149);
not NOT1 (N1158, N1155);
xor XOR2 (N1159, N1146, N736);
xor XOR2 (N1160, N1153, N731);
xor XOR2 (N1161, N1137, N870);
and AND3 (N1162, N1161, N334, N1012);
or OR3 (N1163, N1160, N568, N870);
xor XOR2 (N1164, N1159, N1038);
or OR2 (N1165, N1151, N404);
not NOT1 (N1166, N1132);
buf BUF1 (N1167, N1165);
buf BUF1 (N1168, N1163);
nor NOR2 (N1169, N1156, N877);
nor NOR2 (N1170, N1164, N599);
nor NOR3 (N1171, N1158, N216, N1051);
nand NAND3 (N1172, N1157, N1002, N206);
and AND2 (N1173, N1167, N791);
buf BUF1 (N1174, N1154);
and AND4 (N1175, N1143, N55, N565, N1017);
and AND3 (N1176, N1175, N1134, N57);
nor NOR3 (N1177, N1162, N499, N760);
or OR4 (N1178, N1177, N402, N870, N724);
nor NOR3 (N1179, N1174, N802, N505);
not NOT1 (N1180, N1170);
xor XOR2 (N1181, N1171, N948);
xor XOR2 (N1182, N1176, N129);
not NOT1 (N1183, N1182);
and AND4 (N1184, N1183, N863, N73, N860);
buf BUF1 (N1185, N1178);
xor XOR2 (N1186, N1166, N129);
nand NAND4 (N1187, N1179, N226, N563, N668);
or OR3 (N1188, N1184, N560, N801);
not NOT1 (N1189, N1181);
xor XOR2 (N1190, N1187, N1123);
nand NAND2 (N1191, N1188, N531);
nand NAND2 (N1192, N1185, N588);
buf BUF1 (N1193, N1186);
not NOT1 (N1194, N1189);
nand NAND4 (N1195, N1172, N486, N685, N9);
not NOT1 (N1196, N1190);
nand NAND4 (N1197, N1173, N983, N120, N739);
buf BUF1 (N1198, N1191);
not NOT1 (N1199, N1169);
buf BUF1 (N1200, N1199);
buf BUF1 (N1201, N1195);
and AND4 (N1202, N1197, N868, N950, N864);
buf BUF1 (N1203, N1200);
nand NAND4 (N1204, N1198, N793, N693, N596);
or OR4 (N1205, N1180, N323, N1107, N1161);
buf BUF1 (N1206, N1196);
xor XOR2 (N1207, N1205, N761);
nand NAND3 (N1208, N1201, N510, N1126);
xor XOR2 (N1209, N1203, N22);
or OR3 (N1210, N1168, N528, N1032);
and AND2 (N1211, N1207, N988);
or OR3 (N1212, N1206, N851, N313);
nor NOR4 (N1213, N1212, N656, N856, N898);
xor XOR2 (N1214, N1192, N426);
nand NAND2 (N1215, N1211, N917);
or OR3 (N1216, N1202, N728, N240);
not NOT1 (N1217, N1213);
and AND2 (N1218, N1204, N52);
xor XOR2 (N1219, N1210, N831);
nor NOR2 (N1220, N1217, N277);
nor NOR4 (N1221, N1216, N429, N142, N547);
or OR3 (N1222, N1221, N997, N560);
buf BUF1 (N1223, N1209);
buf BUF1 (N1224, N1220);
not NOT1 (N1225, N1218);
not NOT1 (N1226, N1219);
or OR3 (N1227, N1193, N177, N1200);
not NOT1 (N1228, N1215);
xor XOR2 (N1229, N1222, N491);
nand NAND3 (N1230, N1223, N478, N239);
nand NAND2 (N1231, N1226, N417);
nor NOR2 (N1232, N1231, N49);
not NOT1 (N1233, N1227);
or OR4 (N1234, N1214, N185, N939, N625);
not NOT1 (N1235, N1225);
nand NAND4 (N1236, N1230, N1, N739, N151);
and AND4 (N1237, N1208, N890, N745, N563);
or OR2 (N1238, N1233, N1089);
and AND3 (N1239, N1234, N847, N310);
nand NAND2 (N1240, N1235, N403);
buf BUF1 (N1241, N1232);
xor XOR2 (N1242, N1194, N806);
xor XOR2 (N1243, N1224, N149);
not NOT1 (N1244, N1229);
nor NOR3 (N1245, N1243, N292, N809);
and AND3 (N1246, N1244, N465, N134);
and AND3 (N1247, N1228, N681, N19);
nand NAND4 (N1248, N1246, N661, N762, N1071);
and AND4 (N1249, N1241, N437, N18, N1085);
buf BUF1 (N1250, N1237);
nor NOR4 (N1251, N1242, N217, N1084, N344);
not NOT1 (N1252, N1249);
not NOT1 (N1253, N1236);
nand NAND3 (N1254, N1252, N610, N224);
nand NAND4 (N1255, N1239, N66, N877, N653);
nor NOR3 (N1256, N1245, N777, N1120);
nor NOR3 (N1257, N1256, N874, N440);
not NOT1 (N1258, N1250);
and AND3 (N1259, N1248, N212, N932);
xor XOR2 (N1260, N1258, N112);
xor XOR2 (N1261, N1257, N1);
nand NAND3 (N1262, N1240, N397, N936);
or OR3 (N1263, N1238, N612, N1257);
buf BUF1 (N1264, N1255);
xor XOR2 (N1265, N1262, N410);
buf BUF1 (N1266, N1251);
buf BUF1 (N1267, N1263);
not NOT1 (N1268, N1264);
buf BUF1 (N1269, N1268);
nor NOR2 (N1270, N1265, N551);
xor XOR2 (N1271, N1270, N444);
not NOT1 (N1272, N1253);
buf BUF1 (N1273, N1247);
not NOT1 (N1274, N1272);
nor NOR2 (N1275, N1271, N997);
and AND2 (N1276, N1259, N828);
xor XOR2 (N1277, N1261, N776);
nand NAND4 (N1278, N1260, N331, N838, N714);
not NOT1 (N1279, N1254);
or OR2 (N1280, N1274, N856);
or OR2 (N1281, N1273, N868);
and AND2 (N1282, N1279, N936);
xor XOR2 (N1283, N1282, N767);
xor XOR2 (N1284, N1283, N671);
nand NAND4 (N1285, N1266, N587, N233, N1232);
and AND2 (N1286, N1280, N156);
not NOT1 (N1287, N1284);
not NOT1 (N1288, N1267);
and AND4 (N1289, N1286, N704, N729, N453);
or OR2 (N1290, N1281, N1014);
nand NAND3 (N1291, N1287, N796, N175);
buf BUF1 (N1292, N1290);
xor XOR2 (N1293, N1292, N287);
nor NOR3 (N1294, N1277, N267, N68);
or OR2 (N1295, N1285, N1059);
and AND3 (N1296, N1291, N474, N330);
xor XOR2 (N1297, N1289, N741);
nor NOR3 (N1298, N1293, N972, N136);
buf BUF1 (N1299, N1295);
nand NAND4 (N1300, N1275, N268, N1088, N576);
or OR2 (N1301, N1298, N1288);
nand NAND2 (N1302, N822, N972);
buf BUF1 (N1303, N1269);
not NOT1 (N1304, N1294);
or OR4 (N1305, N1300, N210, N1202, N1005);
not NOT1 (N1306, N1303);
nand NAND2 (N1307, N1305, N621);
not NOT1 (N1308, N1301);
not NOT1 (N1309, N1296);
nor NOR4 (N1310, N1306, N275, N10, N1267);
or OR3 (N1311, N1299, N153, N239);
and AND3 (N1312, N1302, N823, N656);
nor NOR4 (N1313, N1297, N785, N374, N948);
buf BUF1 (N1314, N1278);
not NOT1 (N1315, N1311);
or OR4 (N1316, N1304, N515, N1307, N318);
xor XOR2 (N1317, N851, N124);
nand NAND2 (N1318, N1317, N839);
or OR3 (N1319, N1276, N835, N833);
nand NAND4 (N1320, N1309, N1156, N1301, N921);
nor NOR3 (N1321, N1314, N41, N1052);
xor XOR2 (N1322, N1320, N992);
xor XOR2 (N1323, N1319, N649);
xor XOR2 (N1324, N1312, N586);
and AND3 (N1325, N1310, N1213, N703);
xor XOR2 (N1326, N1323, N1209);
and AND3 (N1327, N1315, N816, N1022);
nor NOR3 (N1328, N1327, N120, N467);
nor NOR4 (N1329, N1322, N1225, N975, N1269);
and AND2 (N1330, N1313, N1135);
xor XOR2 (N1331, N1330, N361);
not NOT1 (N1332, N1329);
xor XOR2 (N1333, N1308, N252);
and AND2 (N1334, N1331, N80);
xor XOR2 (N1335, N1321, N1193);
xor XOR2 (N1336, N1328, N770);
and AND2 (N1337, N1316, N635);
xor XOR2 (N1338, N1335, N724);
nand NAND3 (N1339, N1338, N330, N657);
or OR4 (N1340, N1326, N300, N487, N54);
and AND4 (N1341, N1318, N1276, N1120, N845);
not NOT1 (N1342, N1332);
xor XOR2 (N1343, N1342, N1117);
buf BUF1 (N1344, N1339);
nor NOR4 (N1345, N1343, N525, N1188, N783);
nand NAND2 (N1346, N1333, N950);
nand NAND4 (N1347, N1346, N713, N754, N182);
xor XOR2 (N1348, N1324, N193);
nand NAND4 (N1349, N1337, N1053, N612, N1159);
xor XOR2 (N1350, N1348, N289);
or OR2 (N1351, N1341, N42);
and AND3 (N1352, N1350, N201, N1280);
not NOT1 (N1353, N1347);
or OR3 (N1354, N1340, N892, N1249);
buf BUF1 (N1355, N1344);
nor NOR2 (N1356, N1349, N375);
xor XOR2 (N1357, N1345, N670);
buf BUF1 (N1358, N1357);
or OR3 (N1359, N1355, N981, N828);
buf BUF1 (N1360, N1359);
nor NOR3 (N1361, N1352, N270, N764);
nor NOR4 (N1362, N1334, N988, N900, N323);
nor NOR2 (N1363, N1354, N1073);
not NOT1 (N1364, N1351);
buf BUF1 (N1365, N1325);
nor NOR2 (N1366, N1336, N905);
not NOT1 (N1367, N1356);
nor NOR4 (N1368, N1366, N482, N616, N1092);
xor XOR2 (N1369, N1361, N1073);
xor XOR2 (N1370, N1369, N735);
nor NOR3 (N1371, N1368, N1315, N1153);
nand NAND2 (N1372, N1360, N1276);
xor XOR2 (N1373, N1362, N961);
or OR3 (N1374, N1363, N780, N716);
or OR4 (N1375, N1371, N127, N216, N149);
xor XOR2 (N1376, N1370, N437);
and AND3 (N1377, N1374, N1213, N527);
xor XOR2 (N1378, N1358, N1311);
and AND3 (N1379, N1377, N301, N23);
and AND3 (N1380, N1365, N995, N1234);
nor NOR2 (N1381, N1375, N282);
or OR3 (N1382, N1381, N966, N237);
not NOT1 (N1383, N1353);
not NOT1 (N1384, N1383);
xor XOR2 (N1385, N1364, N638);
nand NAND2 (N1386, N1378, N1208);
nor NOR4 (N1387, N1386, N518, N246, N1216);
and AND4 (N1388, N1379, N548, N650, N639);
nand NAND4 (N1389, N1380, N1242, N1016, N487);
and AND2 (N1390, N1387, N236);
nand NAND2 (N1391, N1390, N437);
buf BUF1 (N1392, N1376);
nand NAND3 (N1393, N1389, N926, N275);
or OR4 (N1394, N1372, N1373, N588, N1314);
nor NOR2 (N1395, N1071, N1274);
xor XOR2 (N1396, N1391, N473);
buf BUF1 (N1397, N1382);
and AND3 (N1398, N1384, N1227, N840);
nand NAND3 (N1399, N1388, N706, N937);
not NOT1 (N1400, N1367);
and AND3 (N1401, N1400, N634, N965);
buf BUF1 (N1402, N1394);
and AND2 (N1403, N1402, N1271);
nand NAND3 (N1404, N1395, N630, N1395);
and AND3 (N1405, N1397, N219, N527);
xor XOR2 (N1406, N1385, N116);
and AND2 (N1407, N1393, N1238);
or OR2 (N1408, N1398, N481);
nor NOR2 (N1409, N1408, N153);
not NOT1 (N1410, N1403);
or OR4 (N1411, N1396, N1102, N1062, N196);
buf BUF1 (N1412, N1407);
nor NOR3 (N1413, N1411, N188, N174);
xor XOR2 (N1414, N1401, N442);
buf BUF1 (N1415, N1409);
or OR4 (N1416, N1413, N287, N308, N1128);
nand NAND4 (N1417, N1404, N467, N763, N205);
not NOT1 (N1418, N1412);
nand NAND4 (N1419, N1410, N183, N1372, N1310);
xor XOR2 (N1420, N1406, N760);
xor XOR2 (N1421, N1418, N290);
xor XOR2 (N1422, N1392, N388);
buf BUF1 (N1423, N1405);
or OR3 (N1424, N1414, N1405, N344);
xor XOR2 (N1425, N1422, N1067);
nor NOR3 (N1426, N1424, N895, N447);
buf BUF1 (N1427, N1420);
xor XOR2 (N1428, N1426, N81);
and AND2 (N1429, N1421, N1085);
nor NOR2 (N1430, N1427, N556);
xor XOR2 (N1431, N1415, N1070);
or OR2 (N1432, N1417, N592);
xor XOR2 (N1433, N1416, N1287);
xor XOR2 (N1434, N1399, N536);
and AND3 (N1435, N1425, N1008, N386);
buf BUF1 (N1436, N1435);
and AND3 (N1437, N1423, N100, N39);
not NOT1 (N1438, N1437);
nand NAND2 (N1439, N1438, N1069);
buf BUF1 (N1440, N1432);
or OR2 (N1441, N1434, N827);
not NOT1 (N1442, N1436);
nor NOR2 (N1443, N1428, N376);
nand NAND3 (N1444, N1443, N618, N149);
xor XOR2 (N1445, N1429, N562);
buf BUF1 (N1446, N1442);
not NOT1 (N1447, N1433);
and AND3 (N1448, N1431, N597, N229);
xor XOR2 (N1449, N1419, N1439);
nand NAND2 (N1450, N1266, N664);
nand NAND2 (N1451, N1450, N1405);
not NOT1 (N1452, N1444);
buf BUF1 (N1453, N1446);
buf BUF1 (N1454, N1430);
not NOT1 (N1455, N1448);
nor NOR2 (N1456, N1441, N720);
nor NOR2 (N1457, N1452, N1230);
nand NAND4 (N1458, N1449, N443, N1225, N666);
nand NAND3 (N1459, N1453, N614, N1271);
nor NOR3 (N1460, N1455, N1335, N682);
nor NOR4 (N1461, N1457, N185, N1324, N125);
nand NAND2 (N1462, N1454, N105);
nor NOR4 (N1463, N1460, N1060, N844, N904);
xor XOR2 (N1464, N1461, N875);
buf BUF1 (N1465, N1463);
nor NOR4 (N1466, N1445, N126, N1117, N526);
buf BUF1 (N1467, N1464);
and AND3 (N1468, N1451, N381, N500);
or OR4 (N1469, N1465, N714, N1285, N1003);
and AND2 (N1470, N1456, N190);
not NOT1 (N1471, N1459);
nand NAND4 (N1472, N1470, N1182, N384, N331);
not NOT1 (N1473, N1462);
not NOT1 (N1474, N1471);
nor NOR3 (N1475, N1469, N1160, N1123);
not NOT1 (N1476, N1472);
or OR3 (N1477, N1473, N417, N433);
and AND4 (N1478, N1440, N824, N1362, N457);
and AND2 (N1479, N1475, N647);
nor NOR3 (N1480, N1466, N954, N475);
not NOT1 (N1481, N1477);
nand NAND3 (N1482, N1468, N519, N1175);
nand NAND4 (N1483, N1481, N560, N792, N926);
nand NAND4 (N1484, N1480, N966, N304, N296);
buf BUF1 (N1485, N1476);
nand NAND2 (N1486, N1479, N851);
not NOT1 (N1487, N1447);
and AND4 (N1488, N1485, N1120, N935, N804);
not NOT1 (N1489, N1482);
buf BUF1 (N1490, N1478);
nor NOR2 (N1491, N1467, N677);
or OR4 (N1492, N1488, N788, N18, N667);
xor XOR2 (N1493, N1483, N545);
nor NOR4 (N1494, N1458, N794, N1241, N233);
xor XOR2 (N1495, N1489, N1014);
xor XOR2 (N1496, N1490, N819);
or OR4 (N1497, N1491, N1132, N918, N99);
nand NAND3 (N1498, N1493, N493, N836);
nor NOR2 (N1499, N1474, N1163);
or OR4 (N1500, N1484, N1316, N1467, N1105);
or OR3 (N1501, N1496, N151, N318);
nor NOR2 (N1502, N1499, N253);
or OR3 (N1503, N1501, N280, N606);
xor XOR2 (N1504, N1495, N1131);
buf BUF1 (N1505, N1502);
or OR3 (N1506, N1494, N1128, N258);
xor XOR2 (N1507, N1487, N687);
and AND3 (N1508, N1497, N901, N298);
not NOT1 (N1509, N1504);
nand NAND3 (N1510, N1509, N1488, N309);
xor XOR2 (N1511, N1486, N259);
and AND4 (N1512, N1508, N464, N611, N475);
or OR3 (N1513, N1505, N733, N324);
xor XOR2 (N1514, N1507, N1181);
buf BUF1 (N1515, N1498);
nor NOR3 (N1516, N1515, N236, N669);
xor XOR2 (N1517, N1500, N233);
not NOT1 (N1518, N1492);
nand NAND4 (N1519, N1513, N664, N289, N833);
xor XOR2 (N1520, N1519, N820);
xor XOR2 (N1521, N1503, N1064);
xor XOR2 (N1522, N1511, N1166);
xor XOR2 (N1523, N1516, N1095);
not NOT1 (N1524, N1521);
xor XOR2 (N1525, N1523, N869);
buf BUF1 (N1526, N1510);
xor XOR2 (N1527, N1506, N143);
or OR3 (N1528, N1514, N504, N135);
nor NOR2 (N1529, N1520, N146);
nand NAND4 (N1530, N1522, N929, N1400, N735);
xor XOR2 (N1531, N1530, N54);
or OR4 (N1532, N1529, N100, N236, N804);
and AND3 (N1533, N1526, N637, N1305);
or OR4 (N1534, N1533, N862, N82, N135);
not NOT1 (N1535, N1525);
not NOT1 (N1536, N1518);
and AND4 (N1537, N1512, N1301, N936, N997);
and AND2 (N1538, N1528, N1261);
not NOT1 (N1539, N1536);
and AND2 (N1540, N1537, N951);
not NOT1 (N1541, N1532);
not NOT1 (N1542, N1531);
nor NOR3 (N1543, N1517, N736, N590);
or OR3 (N1544, N1535, N1487, N405);
buf BUF1 (N1545, N1540);
not NOT1 (N1546, N1539);
nor NOR3 (N1547, N1542, N52, N1416);
nand NAND2 (N1548, N1546, N481);
or OR4 (N1549, N1545, N1276, N331, N849);
not NOT1 (N1550, N1538);
xor XOR2 (N1551, N1547, N406);
or OR2 (N1552, N1541, N236);
and AND3 (N1553, N1544, N904, N821);
xor XOR2 (N1554, N1534, N400);
xor XOR2 (N1555, N1548, N1394);
nand NAND3 (N1556, N1554, N1536, N1402);
or OR3 (N1557, N1551, N300, N1500);
nand NAND4 (N1558, N1527, N97, N1111, N694);
and AND4 (N1559, N1556, N227, N536, N1435);
buf BUF1 (N1560, N1559);
nand NAND2 (N1561, N1560, N740);
buf BUF1 (N1562, N1550);
and AND3 (N1563, N1555, N769, N674);
not NOT1 (N1564, N1563);
or OR2 (N1565, N1562, N960);
nand NAND2 (N1566, N1565, N813);
nand NAND3 (N1567, N1549, N1385, N1296);
not NOT1 (N1568, N1543);
xor XOR2 (N1569, N1557, N1126);
or OR3 (N1570, N1564, N1133, N1142);
buf BUF1 (N1571, N1552);
nand NAND2 (N1572, N1524, N57);
not NOT1 (N1573, N1571);
nand NAND3 (N1574, N1568, N1066, N713);
not NOT1 (N1575, N1572);
and AND3 (N1576, N1566, N356, N766);
and AND2 (N1577, N1576, N1181);
nand NAND3 (N1578, N1558, N1536, N911);
buf BUF1 (N1579, N1570);
or OR4 (N1580, N1567, N521, N1446, N1327);
or OR3 (N1581, N1569, N116, N1197);
or OR4 (N1582, N1581, N1147, N168, N146);
buf BUF1 (N1583, N1574);
not NOT1 (N1584, N1561);
not NOT1 (N1585, N1580);
buf BUF1 (N1586, N1585);
nor NOR3 (N1587, N1582, N1106, N757);
xor XOR2 (N1588, N1578, N1523);
xor XOR2 (N1589, N1587, N450);
or OR2 (N1590, N1579, N766);
not NOT1 (N1591, N1589);
xor XOR2 (N1592, N1575, N1495);
and AND2 (N1593, N1584, N728);
nor NOR4 (N1594, N1583, N1073, N623, N1208);
and AND2 (N1595, N1553, N1576);
not NOT1 (N1596, N1591);
nand NAND4 (N1597, N1596, N910, N1016, N586);
and AND2 (N1598, N1588, N1343);
buf BUF1 (N1599, N1597);
nor NOR3 (N1600, N1590, N1305, N64);
xor XOR2 (N1601, N1598, N425);
nand NAND2 (N1602, N1573, N68);
nand NAND4 (N1603, N1600, N878, N720, N1433);
xor XOR2 (N1604, N1577, N994);
buf BUF1 (N1605, N1586);
and AND3 (N1606, N1592, N1322, N884);
and AND2 (N1607, N1603, N120);
or OR4 (N1608, N1606, N1514, N226, N844);
xor XOR2 (N1609, N1601, N1056);
and AND4 (N1610, N1605, N474, N1490, N1571);
xor XOR2 (N1611, N1593, N463);
buf BUF1 (N1612, N1607);
and AND3 (N1613, N1594, N754, N881);
nor NOR4 (N1614, N1604, N724, N1415, N1021);
nand NAND4 (N1615, N1595, N690, N248, N867);
buf BUF1 (N1616, N1614);
or OR4 (N1617, N1599, N263, N1479, N464);
xor XOR2 (N1618, N1616, N1407);
and AND4 (N1619, N1602, N13, N1334, N431);
and AND3 (N1620, N1608, N1135, N18);
not NOT1 (N1621, N1609);
buf BUF1 (N1622, N1612);
nor NOR3 (N1623, N1619, N1511, N1236);
not NOT1 (N1624, N1613);
not NOT1 (N1625, N1617);
not NOT1 (N1626, N1615);
and AND3 (N1627, N1624, N832, N1214);
nand NAND4 (N1628, N1623, N1233, N1470, N836);
and AND4 (N1629, N1627, N1458, N496, N565);
buf BUF1 (N1630, N1621);
nand NAND3 (N1631, N1628, N799, N571);
buf BUF1 (N1632, N1629);
and AND2 (N1633, N1632, N346);
xor XOR2 (N1634, N1622, N896);
or OR2 (N1635, N1625, N60);
xor XOR2 (N1636, N1631, N1562);
or OR4 (N1637, N1618, N1143, N288, N618);
or OR4 (N1638, N1637, N779, N701, N1026);
or OR4 (N1639, N1611, N1392, N326, N357);
xor XOR2 (N1640, N1630, N643);
xor XOR2 (N1641, N1610, N118);
and AND4 (N1642, N1620, N1305, N1633, N822);
and AND2 (N1643, N1084, N87);
xor XOR2 (N1644, N1626, N166);
nor NOR4 (N1645, N1639, N1350, N1431, N654);
nand NAND4 (N1646, N1645, N1273, N510, N579);
nor NOR2 (N1647, N1635, N642);
buf BUF1 (N1648, N1641);
and AND3 (N1649, N1644, N1639, N1441);
not NOT1 (N1650, N1648);
not NOT1 (N1651, N1646);
nand NAND4 (N1652, N1651, N1171, N1027, N551);
and AND4 (N1653, N1638, N1111, N1175, N1283);
not NOT1 (N1654, N1643);
nor NOR2 (N1655, N1652, N1590);
nor NOR2 (N1656, N1634, N19);
nand NAND4 (N1657, N1656, N1364, N992, N1513);
or OR2 (N1658, N1650, N1099);
xor XOR2 (N1659, N1647, N1648);
buf BUF1 (N1660, N1642);
nand NAND2 (N1661, N1653, N180);
nand NAND3 (N1662, N1660, N246, N1317);
or OR3 (N1663, N1662, N1551, N1077);
or OR3 (N1664, N1655, N1444, N1225);
and AND4 (N1665, N1663, N875, N1119, N489);
nor NOR4 (N1666, N1665, N881, N1564, N592);
buf BUF1 (N1667, N1636);
buf BUF1 (N1668, N1661);
or OR3 (N1669, N1658, N1379, N1066);
nand NAND4 (N1670, N1640, N1476, N1634, N720);
nand NAND4 (N1671, N1669, N334, N312, N911);
nor NOR2 (N1672, N1657, N114);
xor XOR2 (N1673, N1668, N468);
not NOT1 (N1674, N1673);
xor XOR2 (N1675, N1664, N486);
nor NOR3 (N1676, N1659, N823, N453);
and AND2 (N1677, N1672, N956);
buf BUF1 (N1678, N1674);
and AND3 (N1679, N1649, N1177, N1308);
or OR3 (N1680, N1679, N173, N30);
and AND4 (N1681, N1676, N816, N1422, N519);
not NOT1 (N1682, N1681);
xor XOR2 (N1683, N1670, N865);
nor NOR2 (N1684, N1678, N427);
not NOT1 (N1685, N1675);
buf BUF1 (N1686, N1666);
nor NOR3 (N1687, N1654, N642, N1198);
nand NAND2 (N1688, N1682, N313);
buf BUF1 (N1689, N1687);
and AND4 (N1690, N1671, N185, N641, N1109);
nand NAND4 (N1691, N1680, N848, N1424, N225);
xor XOR2 (N1692, N1684, N143);
nor NOR4 (N1693, N1688, N636, N59, N426);
or OR3 (N1694, N1693, N941, N728);
buf BUF1 (N1695, N1677);
nand NAND2 (N1696, N1686, N34);
and AND3 (N1697, N1694, N43, N114);
not NOT1 (N1698, N1692);
not NOT1 (N1699, N1689);
not NOT1 (N1700, N1691);
nor NOR4 (N1701, N1697, N1331, N1266, N1558);
and AND3 (N1702, N1699, N934, N1686);
and AND4 (N1703, N1685, N195, N1626, N1286);
and AND4 (N1704, N1703, N632, N471, N355);
and AND4 (N1705, N1683, N422, N1419, N1038);
and AND4 (N1706, N1667, N280, N1630, N1267);
not NOT1 (N1707, N1698);
nand NAND2 (N1708, N1700, N418);
buf BUF1 (N1709, N1704);
not NOT1 (N1710, N1705);
xor XOR2 (N1711, N1708, N1293);
nand NAND3 (N1712, N1710, N1154, N1492);
or OR2 (N1713, N1701, N508);
buf BUF1 (N1714, N1706);
nand NAND2 (N1715, N1702, N772);
or OR4 (N1716, N1715, N1469, N1059, N628);
or OR4 (N1717, N1690, N1623, N384, N241);
buf BUF1 (N1718, N1695);
nand NAND2 (N1719, N1718, N533);
xor XOR2 (N1720, N1709, N914);
nand NAND4 (N1721, N1707, N75, N1707, N1261);
nor NOR4 (N1722, N1721, N1654, N1116, N1625);
xor XOR2 (N1723, N1714, N577);
not NOT1 (N1724, N1713);
xor XOR2 (N1725, N1716, N1121);
xor XOR2 (N1726, N1723, N1191);
nor NOR3 (N1727, N1726, N1193, N901);
buf BUF1 (N1728, N1727);
or OR2 (N1729, N1724, N700);
and AND4 (N1730, N1719, N126, N1198, N1660);
not NOT1 (N1731, N1712);
xor XOR2 (N1732, N1728, N216);
or OR3 (N1733, N1696, N1582, N249);
or OR2 (N1734, N1725, N1000);
nand NAND2 (N1735, N1717, N856);
xor XOR2 (N1736, N1734, N406);
or OR4 (N1737, N1729, N1381, N1600, N1630);
xor XOR2 (N1738, N1720, N1348);
not NOT1 (N1739, N1722);
nor NOR2 (N1740, N1733, N1181);
nor NOR4 (N1741, N1739, N180, N178, N1338);
or OR4 (N1742, N1730, N1102, N1319, N456);
or OR4 (N1743, N1711, N479, N677, N877);
and AND3 (N1744, N1736, N1648, N1466);
buf BUF1 (N1745, N1744);
buf BUF1 (N1746, N1740);
and AND3 (N1747, N1745, N290, N1286);
nor NOR4 (N1748, N1738, N269, N1239, N837);
buf BUF1 (N1749, N1741);
and AND4 (N1750, N1743, N406, N219, N45);
nand NAND3 (N1751, N1732, N1135, N1165);
buf BUF1 (N1752, N1742);
and AND4 (N1753, N1746, N204, N1322, N420);
nand NAND2 (N1754, N1752, N180);
and AND3 (N1755, N1747, N1409, N1081);
nand NAND2 (N1756, N1751, N389);
xor XOR2 (N1757, N1753, N1643);
nand NAND3 (N1758, N1755, N1192, N1202);
or OR2 (N1759, N1757, N1194);
and AND3 (N1760, N1754, N1177, N831);
and AND3 (N1761, N1760, N1225, N1295);
nand NAND4 (N1762, N1750, N227, N245, N322);
not NOT1 (N1763, N1735);
or OR2 (N1764, N1749, N1341);
and AND4 (N1765, N1756, N61, N1547, N271);
xor XOR2 (N1766, N1761, N735);
xor XOR2 (N1767, N1763, N858);
nand NAND4 (N1768, N1748, N325, N177, N721);
nor NOR3 (N1769, N1767, N863, N949);
or OR4 (N1770, N1765, N942, N643, N46);
or OR4 (N1771, N1766, N15, N1577, N1426);
not NOT1 (N1772, N1731);
and AND4 (N1773, N1758, N165, N98, N877);
not NOT1 (N1774, N1773);
nand NAND4 (N1775, N1774, N607, N1693, N1116);
nor NOR4 (N1776, N1762, N1626, N1230, N375);
and AND2 (N1777, N1768, N592);
not NOT1 (N1778, N1776);
buf BUF1 (N1779, N1759);
xor XOR2 (N1780, N1770, N1457);
nor NOR4 (N1781, N1737, N882, N1381, N1079);
xor XOR2 (N1782, N1780, N1321);
xor XOR2 (N1783, N1771, N1403);
and AND2 (N1784, N1775, N887);
or OR2 (N1785, N1769, N1154);
or OR3 (N1786, N1785, N59, N1562);
or OR2 (N1787, N1778, N625);
nand NAND4 (N1788, N1787, N4, N239, N120);
or OR4 (N1789, N1779, N1471, N1174, N1000);
and AND2 (N1790, N1777, N1009);
not NOT1 (N1791, N1789);
and AND4 (N1792, N1790, N1339, N175, N1447);
nand NAND4 (N1793, N1764, N706, N1699, N621);
and AND4 (N1794, N1786, N59, N440, N1747);
xor XOR2 (N1795, N1792, N482);
not NOT1 (N1796, N1781);
buf BUF1 (N1797, N1796);
and AND3 (N1798, N1783, N907, N729);
nand NAND4 (N1799, N1788, N509, N1103, N626);
or OR3 (N1800, N1784, N775, N393);
xor XOR2 (N1801, N1800, N1758);
buf BUF1 (N1802, N1798);
nor NOR4 (N1803, N1799, N1481, N943, N10);
nand NAND2 (N1804, N1782, N175);
not NOT1 (N1805, N1791);
nand NAND2 (N1806, N1805, N1456);
xor XOR2 (N1807, N1772, N1546);
not NOT1 (N1808, N1807);
and AND4 (N1809, N1801, N193, N1263, N1803);
or OR4 (N1810, N973, N791, N1420, N1417);
nor NOR3 (N1811, N1806, N1014, N585);
buf BUF1 (N1812, N1797);
buf BUF1 (N1813, N1795);
nor NOR2 (N1814, N1810, N1122);
or OR3 (N1815, N1814, N159, N172);
not NOT1 (N1816, N1815);
and AND2 (N1817, N1804, N533);
not NOT1 (N1818, N1813);
nor NOR3 (N1819, N1816, N1657, N1464);
xor XOR2 (N1820, N1809, N591);
or OR2 (N1821, N1802, N1489);
or OR4 (N1822, N1820, N722, N289, N1767);
buf BUF1 (N1823, N1821);
buf BUF1 (N1824, N1818);
xor XOR2 (N1825, N1793, N1799);
nor NOR2 (N1826, N1819, N839);
not NOT1 (N1827, N1823);
xor XOR2 (N1828, N1808, N1175);
nor NOR4 (N1829, N1812, N1358, N996, N776);
nand NAND3 (N1830, N1822, N1760, N521);
and AND2 (N1831, N1826, N474);
nand NAND2 (N1832, N1824, N1698);
xor XOR2 (N1833, N1829, N106);
not NOT1 (N1834, N1828);
or OR4 (N1835, N1794, N364, N1681, N1203);
not NOT1 (N1836, N1832);
nor NOR2 (N1837, N1835, N666);
nor NOR3 (N1838, N1834, N1404, N1393);
buf BUF1 (N1839, N1836);
buf BUF1 (N1840, N1817);
or OR3 (N1841, N1830, N1806, N156);
buf BUF1 (N1842, N1841);
nand NAND4 (N1843, N1811, N1426, N40, N1201);
not NOT1 (N1844, N1833);
and AND4 (N1845, N1838, N36, N421, N1487);
xor XOR2 (N1846, N1839, N1382);
buf BUF1 (N1847, N1846);
xor XOR2 (N1848, N1825, N885);
or OR3 (N1849, N1844, N1282, N519);
nor NOR4 (N1850, N1843, N765, N916, N1508);
xor XOR2 (N1851, N1840, N427);
nor NOR2 (N1852, N1842, N1050);
nand NAND4 (N1853, N1827, N1775, N1799, N1196);
or OR4 (N1854, N1847, N1471, N748, N370);
nor NOR4 (N1855, N1851, N1323, N1606, N870);
nor NOR2 (N1856, N1831, N1128);
nand NAND3 (N1857, N1856, N11, N20);
buf BUF1 (N1858, N1837);
nor NOR3 (N1859, N1857, N905, N1139);
not NOT1 (N1860, N1848);
nor NOR3 (N1861, N1852, N1042, N1045);
buf BUF1 (N1862, N1858);
and AND4 (N1863, N1845, N1533, N508, N523);
nand NAND4 (N1864, N1860, N1217, N1623, N1132);
nand NAND3 (N1865, N1850, N789, N1004);
and AND4 (N1866, N1854, N688, N1496, N697);
nand NAND4 (N1867, N1863, N261, N973, N747);
nand NAND2 (N1868, N1855, N1052);
not NOT1 (N1869, N1866);
xor XOR2 (N1870, N1861, N611);
buf BUF1 (N1871, N1865);
nor NOR4 (N1872, N1859, N262, N1702, N255);
nand NAND2 (N1873, N1864, N719);
buf BUF1 (N1874, N1849);
and AND3 (N1875, N1870, N1791, N116);
nand NAND4 (N1876, N1873, N168, N612, N1568);
buf BUF1 (N1877, N1869);
nor NOR2 (N1878, N1877, N1050);
not NOT1 (N1879, N1875);
nand NAND2 (N1880, N1867, N313);
or OR4 (N1881, N1874, N607, N1426, N240);
nand NAND3 (N1882, N1853, N1150, N1452);
nor NOR4 (N1883, N1876, N1776, N1036, N1683);
xor XOR2 (N1884, N1880, N1011);
nor NOR2 (N1885, N1878, N4);
or OR3 (N1886, N1884, N901, N623);
nor NOR4 (N1887, N1883, N840, N175, N1118);
buf BUF1 (N1888, N1872);
xor XOR2 (N1889, N1862, N193);
xor XOR2 (N1890, N1886, N1562);
and AND3 (N1891, N1871, N172, N892);
nand NAND3 (N1892, N1881, N1038, N1759);
or OR3 (N1893, N1889, N1125, N75);
buf BUF1 (N1894, N1892);
and AND3 (N1895, N1893, N894, N1390);
buf BUF1 (N1896, N1894);
nand NAND2 (N1897, N1891, N1642);
and AND3 (N1898, N1885, N969, N167);
or OR2 (N1899, N1895, N791);
not NOT1 (N1900, N1879);
not NOT1 (N1901, N1868);
buf BUF1 (N1902, N1898);
nand NAND2 (N1903, N1888, N347);
buf BUF1 (N1904, N1890);
nor NOR4 (N1905, N1901, N1724, N857, N160);
nor NOR3 (N1906, N1882, N617, N1585);
xor XOR2 (N1907, N1900, N737);
and AND4 (N1908, N1897, N1550, N1581, N19);
buf BUF1 (N1909, N1906);
not NOT1 (N1910, N1909);
xor XOR2 (N1911, N1907, N930);
or OR3 (N1912, N1902, N1773, N1910);
xor XOR2 (N1913, N1680, N1614);
nand NAND3 (N1914, N1887, N199, N411);
or OR2 (N1915, N1911, N1602);
nor NOR2 (N1916, N1908, N398);
xor XOR2 (N1917, N1903, N1915);
and AND2 (N1918, N992, N287);
or OR3 (N1919, N1913, N298, N1098);
nor NOR3 (N1920, N1905, N1751, N287);
not NOT1 (N1921, N1914);
xor XOR2 (N1922, N1921, N562);
xor XOR2 (N1923, N1919, N1140);
not NOT1 (N1924, N1923);
buf BUF1 (N1925, N1899);
xor XOR2 (N1926, N1920, N587);
xor XOR2 (N1927, N1918, N669);
buf BUF1 (N1928, N1925);
and AND3 (N1929, N1924, N989, N1159);
xor XOR2 (N1930, N1896, N1143);
nor NOR3 (N1931, N1927, N394, N406);
buf BUF1 (N1932, N1931);
and AND2 (N1933, N1928, N367);
xor XOR2 (N1934, N1926, N1141);
buf BUF1 (N1935, N1933);
or OR4 (N1936, N1917, N1756, N1906, N814);
nor NOR2 (N1937, N1932, N325);
nand NAND2 (N1938, N1934, N711);
or OR2 (N1939, N1938, N454);
xor XOR2 (N1940, N1939, N96);
or OR3 (N1941, N1937, N1226, N1922);
nor NOR2 (N1942, N1165, N546);
and AND4 (N1943, N1930, N165, N1466, N1794);
and AND3 (N1944, N1936, N1894, N1580);
and AND2 (N1945, N1944, N1293);
nand NAND3 (N1946, N1935, N1496, N1668);
nand NAND4 (N1947, N1945, N227, N980, N929);
xor XOR2 (N1948, N1946, N1223);
buf BUF1 (N1949, N1947);
or OR2 (N1950, N1916, N788);
xor XOR2 (N1951, N1940, N39);
or OR3 (N1952, N1929, N419, N1771);
buf BUF1 (N1953, N1904);
not NOT1 (N1954, N1952);
xor XOR2 (N1955, N1941, N1799);
buf BUF1 (N1956, N1954);
nor NOR4 (N1957, N1949, N717, N1937, N1557);
buf BUF1 (N1958, N1951);
or OR2 (N1959, N1957, N1932);
buf BUF1 (N1960, N1953);
nor NOR3 (N1961, N1942, N1776, N829);
not NOT1 (N1962, N1959);
xor XOR2 (N1963, N1962, N1822);
xor XOR2 (N1964, N1963, N1436);
buf BUF1 (N1965, N1912);
buf BUF1 (N1966, N1961);
or OR3 (N1967, N1956, N675, N375);
and AND2 (N1968, N1966, N280);
xor XOR2 (N1969, N1967, N1759);
nand NAND4 (N1970, N1958, N512, N1833, N765);
not NOT1 (N1971, N1964);
and AND4 (N1972, N1971, N1379, N126, N224);
nand NAND3 (N1973, N1960, N1626, N623);
buf BUF1 (N1974, N1970);
and AND4 (N1975, N1948, N818, N1398, N1094);
buf BUF1 (N1976, N1974);
buf BUF1 (N1977, N1969);
buf BUF1 (N1978, N1972);
or OR2 (N1979, N1975, N981);
not NOT1 (N1980, N1965);
and AND3 (N1981, N1950, N678, N709);
nor NOR3 (N1982, N1973, N371, N522);
buf BUF1 (N1983, N1979);
not NOT1 (N1984, N1955);
or OR2 (N1985, N1983, N147);
xor XOR2 (N1986, N1976, N1048);
nor NOR4 (N1987, N1986, N541, N1714, N142);
not NOT1 (N1988, N1982);
buf BUF1 (N1989, N1980);
xor XOR2 (N1990, N1985, N540);
xor XOR2 (N1991, N1990, N760);
xor XOR2 (N1992, N1968, N1756);
buf BUF1 (N1993, N1989);
nand NAND4 (N1994, N1991, N1941, N1032, N562);
buf BUF1 (N1995, N1993);
xor XOR2 (N1996, N1943, N1832);
buf BUF1 (N1997, N1987);
nor NOR2 (N1998, N1978, N599);
or OR2 (N1999, N1981, N1412);
xor XOR2 (N2000, N1984, N964);
or OR3 (N2001, N1994, N1740, N630);
or OR4 (N2002, N1992, N1607, N686, N753);
nor NOR4 (N2003, N1988, N1986, N877, N1225);
not NOT1 (N2004, N2002);
or OR4 (N2005, N1998, N1058, N1428, N30);
nor NOR3 (N2006, N2004, N38, N1471);
buf BUF1 (N2007, N1999);
buf BUF1 (N2008, N2001);
or OR2 (N2009, N2008, N226);
and AND2 (N2010, N1977, N1749);
nand NAND2 (N2011, N2003, N1537);
not NOT1 (N2012, N1996);
nand NAND2 (N2013, N2011, N500);
buf BUF1 (N2014, N1995);
nand NAND3 (N2015, N2005, N653, N1213);
and AND2 (N2016, N2015, N1946);
or OR3 (N2017, N2007, N415, N502);
not NOT1 (N2018, N1997);
buf BUF1 (N2019, N2012);
and AND2 (N2020, N2000, N758);
buf BUF1 (N2021, N2010);
or OR2 (N2022, N2009, N598);
or OR4 (N2023, N2006, N942, N1916, N1237);
nor NOR4 (N2024, N2022, N1353, N1395, N918);
xor XOR2 (N2025, N2020, N1808);
nor NOR4 (N2026, N2024, N454, N730, N935);
and AND4 (N2027, N2014, N1696, N528, N1314);
and AND4 (N2028, N2018, N626, N1406, N901);
and AND3 (N2029, N2019, N1694, N613);
buf BUF1 (N2030, N2028);
and AND3 (N2031, N2021, N547, N1865);
or OR3 (N2032, N2016, N1814, N620);
nor NOR4 (N2033, N2027, N1228, N1151, N1237);
not NOT1 (N2034, N2029);
not NOT1 (N2035, N2025);
not NOT1 (N2036, N2032);
nand NAND3 (N2037, N2036, N427, N813);
xor XOR2 (N2038, N2030, N1941);
not NOT1 (N2039, N2017);
nand NAND4 (N2040, N2039, N1069, N573, N1337);
or OR3 (N2041, N2031, N3, N378);
buf BUF1 (N2042, N2038);
or OR3 (N2043, N2023, N903, N1627);
and AND3 (N2044, N2037, N456, N669);
nor NOR4 (N2045, N2043, N821, N988, N1259);
nand NAND3 (N2046, N2041, N1047, N1612);
nand NAND2 (N2047, N2044, N1709);
buf BUF1 (N2048, N2042);
nor NOR4 (N2049, N2040, N1043, N994, N93);
or OR4 (N2050, N2026, N885, N858, N1329);
not NOT1 (N2051, N2034);
and AND3 (N2052, N2045, N326, N430);
not NOT1 (N2053, N2048);
buf BUF1 (N2054, N2051);
and AND2 (N2055, N2053, N656);
nand NAND2 (N2056, N2054, N1191);
xor XOR2 (N2057, N2033, N1006);
buf BUF1 (N2058, N2057);
and AND3 (N2059, N2055, N372, N1309);
nand NAND4 (N2060, N2050, N1727, N1326, N112);
xor XOR2 (N2061, N2056, N754);
not NOT1 (N2062, N2035);
buf BUF1 (N2063, N2062);
nand NAND2 (N2064, N2060, N1527);
buf BUF1 (N2065, N2052);
xor XOR2 (N2066, N2061, N1848);
or OR3 (N2067, N2066, N1539, N1530);
not NOT1 (N2068, N2064);
xor XOR2 (N2069, N2049, N11);
or OR4 (N2070, N2058, N1630, N575, N1343);
not NOT1 (N2071, N2013);
and AND3 (N2072, N2065, N1322, N313);
or OR2 (N2073, N2063, N1223);
or OR2 (N2074, N2072, N1840);
buf BUF1 (N2075, N2073);
nor NOR2 (N2076, N2047, N1164);
nor NOR4 (N2077, N2076, N172, N502, N133);
nand NAND2 (N2078, N2068, N3);
buf BUF1 (N2079, N2059);
or OR3 (N2080, N2069, N1302, N987);
xor XOR2 (N2081, N2080, N186);
and AND3 (N2082, N2077, N1700, N373);
and AND4 (N2083, N2082, N1835, N1332, N1785);
nand NAND2 (N2084, N2078, N448);
or OR3 (N2085, N2081, N1352, N169);
not NOT1 (N2086, N2079);
buf BUF1 (N2087, N2067);
or OR4 (N2088, N2074, N1533, N1675, N1337);
not NOT1 (N2089, N2088);
xor XOR2 (N2090, N2086, N1611);
nand NAND2 (N2091, N2083, N1190);
not NOT1 (N2092, N2084);
nand NAND2 (N2093, N2070, N497);
buf BUF1 (N2094, N2091);
or OR3 (N2095, N2093, N1747, N1537);
and AND3 (N2096, N2089, N1596, N387);
nor NOR2 (N2097, N2071, N2036);
not NOT1 (N2098, N2075);
xor XOR2 (N2099, N2098, N1473);
buf BUF1 (N2100, N2090);
not NOT1 (N2101, N2092);
and AND3 (N2102, N2096, N1548, N354);
and AND4 (N2103, N2094, N772, N2036, N1034);
nor NOR4 (N2104, N2097, N1052, N689, N1454);
buf BUF1 (N2105, N2085);
buf BUF1 (N2106, N2104);
buf BUF1 (N2107, N2103);
buf BUF1 (N2108, N2099);
buf BUF1 (N2109, N2108);
or OR2 (N2110, N2105, N1931);
nor NOR3 (N2111, N2109, N47, N1256);
buf BUF1 (N2112, N2111);
nor NOR4 (N2113, N2112, N1612, N1572, N948);
nor NOR4 (N2114, N2087, N2090, N1378, N204);
and AND2 (N2115, N2114, N1210);
xor XOR2 (N2116, N2046, N1467);
xor XOR2 (N2117, N2100, N1473);
nand NAND2 (N2118, N2101, N888);
and AND2 (N2119, N2117, N1311);
nor NOR2 (N2120, N2110, N135);
nor NOR3 (N2121, N2116, N863, N615);
and AND3 (N2122, N2120, N1308, N1243);
and AND2 (N2123, N2102, N1199);
nor NOR3 (N2124, N2106, N530, N2055);
nor NOR4 (N2125, N2115, N41, N205, N548);
or OR3 (N2126, N2113, N683, N942);
buf BUF1 (N2127, N2125);
and AND4 (N2128, N2124, N437, N1223, N823);
xor XOR2 (N2129, N2119, N1682);
buf BUF1 (N2130, N2129);
nand NAND4 (N2131, N2095, N1580, N318, N682);
buf BUF1 (N2132, N2118);
nor NOR4 (N2133, N2128, N1299, N397, N479);
xor XOR2 (N2134, N2121, N27);
or OR3 (N2135, N2133, N1812, N707);
nor NOR4 (N2136, N2126, N1214, N2030, N1931);
nor NOR2 (N2137, N2135, N1311);
buf BUF1 (N2138, N2130);
or OR4 (N2139, N2138, N301, N431, N1072);
buf BUF1 (N2140, N2107);
nand NAND3 (N2141, N2123, N420, N825);
or OR4 (N2142, N2139, N1311, N1351, N101);
or OR2 (N2143, N2132, N1283);
and AND2 (N2144, N2122, N1936);
or OR4 (N2145, N2137, N2102, N1712, N840);
and AND3 (N2146, N2144, N120, N956);
nand NAND3 (N2147, N2134, N1837, N30);
nor NOR2 (N2148, N2146, N558);
not NOT1 (N2149, N2145);
nand NAND2 (N2150, N2140, N97);
not NOT1 (N2151, N2127);
not NOT1 (N2152, N2150);
not NOT1 (N2153, N2143);
nor NOR3 (N2154, N2136, N283, N63);
and AND3 (N2155, N2147, N110, N1541);
nand NAND2 (N2156, N2148, N2010);
nand NAND2 (N2157, N2155, N765);
nor NOR3 (N2158, N2141, N1655, N690);
nor NOR4 (N2159, N2158, N366, N2093, N594);
nor NOR4 (N2160, N2151, N1318, N1225, N1225);
nand NAND3 (N2161, N2156, N81, N59);
not NOT1 (N2162, N2154);
not NOT1 (N2163, N2131);
nor NOR4 (N2164, N2162, N2013, N1761, N119);
xor XOR2 (N2165, N2160, N1879);
nor NOR2 (N2166, N2152, N1101);
not NOT1 (N2167, N2161);
nor NOR2 (N2168, N2149, N2075);
and AND3 (N2169, N2159, N954, N99);
not NOT1 (N2170, N2163);
or OR4 (N2171, N2157, N700, N1611, N852);
nor NOR3 (N2172, N2170, N1428, N2146);
not NOT1 (N2173, N2153);
nor NOR4 (N2174, N2169, N1290, N1209, N640);
nor NOR3 (N2175, N2168, N2014, N1812);
nand NAND3 (N2176, N2173, N1391, N1669);
xor XOR2 (N2177, N2174, N770);
or OR3 (N2178, N2166, N49, N538);
nor NOR4 (N2179, N2142, N37, N1226, N1408);
buf BUF1 (N2180, N2164);
not NOT1 (N2181, N2178);
nand NAND2 (N2182, N2180, N909);
nand NAND3 (N2183, N2175, N1940, N786);
or OR2 (N2184, N2181, N620);
nor NOR2 (N2185, N2172, N63);
xor XOR2 (N2186, N2184, N1548);
nor NOR4 (N2187, N2177, N263, N266, N1916);
buf BUF1 (N2188, N2179);
and AND3 (N2189, N2165, N1984, N1102);
nor NOR4 (N2190, N2183, N1041, N344, N1676);
buf BUF1 (N2191, N2182);
nor NOR3 (N2192, N2191, N131, N560);
and AND2 (N2193, N2190, N1189);
buf BUF1 (N2194, N2192);
or OR4 (N2195, N2176, N1604, N1330, N2115);
xor XOR2 (N2196, N2189, N892);
and AND3 (N2197, N2193, N212, N1169);
not NOT1 (N2198, N2167);
or OR3 (N2199, N2186, N1428, N1719);
xor XOR2 (N2200, N2185, N2177);
nand NAND4 (N2201, N2199, N783, N660, N1798);
not NOT1 (N2202, N2201);
and AND2 (N2203, N2197, N565);
not NOT1 (N2204, N2195);
xor XOR2 (N2205, N2188, N1380);
xor XOR2 (N2206, N2200, N1615);
nor NOR3 (N2207, N2196, N1421, N237);
not NOT1 (N2208, N2194);
or OR2 (N2209, N2202, N1678);
buf BUF1 (N2210, N2209);
or OR2 (N2211, N2205, N818);
nor NOR2 (N2212, N2198, N22);
xor XOR2 (N2213, N2187, N1943);
nor NOR3 (N2214, N2211, N2182, N578);
and AND3 (N2215, N2210, N306, N2161);
buf BUF1 (N2216, N2214);
nand NAND3 (N2217, N2213, N379, N1042);
xor XOR2 (N2218, N2217, N1377);
not NOT1 (N2219, N2208);
and AND2 (N2220, N2206, N1361);
nor NOR4 (N2221, N2220, N1837, N1216, N1960);
nor NOR2 (N2222, N2203, N393);
nor NOR4 (N2223, N2222, N174, N1902, N1271);
and AND4 (N2224, N2223, N1105, N2156, N775);
nand NAND3 (N2225, N2207, N1852, N796);
not NOT1 (N2226, N2212);
buf BUF1 (N2227, N2204);
or OR2 (N2228, N2226, N2123);
not NOT1 (N2229, N2219);
nor NOR4 (N2230, N2224, N1136, N2000, N1318);
or OR3 (N2231, N2227, N1615, N578);
not NOT1 (N2232, N2230);
nand NAND2 (N2233, N2221, N2193);
or OR3 (N2234, N2233, N499, N2110);
nand NAND2 (N2235, N2215, N89);
buf BUF1 (N2236, N2218);
nor NOR4 (N2237, N2171, N2175, N1971, N924);
and AND3 (N2238, N2228, N1004, N364);
buf BUF1 (N2239, N2216);
not NOT1 (N2240, N2234);
not NOT1 (N2241, N2229);
nor NOR2 (N2242, N2231, N1591);
not NOT1 (N2243, N2236);
not NOT1 (N2244, N2243);
buf BUF1 (N2245, N2232);
nor NOR2 (N2246, N2239, N65);
and AND2 (N2247, N2235, N131);
nand NAND4 (N2248, N2238, N2245, N879, N1412);
xor XOR2 (N2249, N552, N133);
not NOT1 (N2250, N2242);
not NOT1 (N2251, N2246);
and AND4 (N2252, N2244, N507, N137, N1920);
buf BUF1 (N2253, N2252);
or OR3 (N2254, N2237, N762, N623);
nand NAND4 (N2255, N2248, N1708, N611, N845);
and AND3 (N2256, N2255, N1519, N813);
or OR4 (N2257, N2241, N486, N679, N347);
nor NOR4 (N2258, N2256, N1205, N1359, N1572);
nor NOR4 (N2259, N2247, N1261, N1125, N215);
nand NAND3 (N2260, N2258, N394, N1757);
not NOT1 (N2261, N2254);
buf BUF1 (N2262, N2240);
or OR2 (N2263, N2259, N2240);
not NOT1 (N2264, N2250);
not NOT1 (N2265, N2253);
or OR4 (N2266, N2225, N808, N958, N219);
nand NAND2 (N2267, N2266, N2123);
not NOT1 (N2268, N2251);
xor XOR2 (N2269, N2261, N102);
not NOT1 (N2270, N2264);
and AND3 (N2271, N2257, N23, N2218);
xor XOR2 (N2272, N2260, N966);
and AND3 (N2273, N2271, N1508, N1270);
and AND4 (N2274, N2267, N313, N726, N1682);
and AND4 (N2275, N2274, N1429, N105, N959);
and AND4 (N2276, N2269, N218, N631, N603);
nand NAND2 (N2277, N2263, N1689);
or OR4 (N2278, N2277, N986, N79, N1470);
nor NOR2 (N2279, N2273, N473);
xor XOR2 (N2280, N2276, N1900);
not NOT1 (N2281, N2275);
not NOT1 (N2282, N2281);
buf BUF1 (N2283, N2278);
nor NOR3 (N2284, N2272, N2133, N380);
buf BUF1 (N2285, N2280);
buf BUF1 (N2286, N2249);
nand NAND3 (N2287, N2268, N204, N549);
nor NOR3 (N2288, N2287, N296, N454);
nand NAND2 (N2289, N2286, N1847);
not NOT1 (N2290, N2265);
nand NAND2 (N2291, N2262, N1800);
xor XOR2 (N2292, N2270, N1010);
nor NOR3 (N2293, N2283, N1386, N667);
or OR2 (N2294, N2293, N1706);
not NOT1 (N2295, N2290);
nor NOR4 (N2296, N2288, N1274, N530, N713);
buf BUF1 (N2297, N2294);
or OR2 (N2298, N2279, N1112);
nand NAND4 (N2299, N2289, N2129, N903, N1034);
and AND3 (N2300, N2285, N723, N1798);
not NOT1 (N2301, N2292);
or OR3 (N2302, N2297, N1565, N2161);
or OR2 (N2303, N2282, N403);
not NOT1 (N2304, N2303);
buf BUF1 (N2305, N2300);
nand NAND3 (N2306, N2301, N694, N1201);
nand NAND2 (N2307, N2295, N441);
and AND2 (N2308, N2298, N76);
and AND2 (N2309, N2308, N106);
nand NAND3 (N2310, N2284, N1205, N354);
nand NAND3 (N2311, N2304, N1738, N511);
nor NOR2 (N2312, N2299, N2112);
or OR2 (N2313, N2291, N1846);
not NOT1 (N2314, N2309);
and AND2 (N2315, N2312, N215);
and AND3 (N2316, N2307, N489, N790);
and AND4 (N2317, N2306, N50, N2211, N467);
buf BUF1 (N2318, N2317);
buf BUF1 (N2319, N2311);
buf BUF1 (N2320, N2319);
xor XOR2 (N2321, N2305, N1301);
xor XOR2 (N2322, N2296, N1976);
or OR2 (N2323, N2315, N1388);
and AND2 (N2324, N2318, N446);
buf BUF1 (N2325, N2322);
not NOT1 (N2326, N2324);
and AND4 (N2327, N2314, N2141, N15, N1069);
nand NAND3 (N2328, N2321, N960, N774);
nand NAND2 (N2329, N2302, N1869);
and AND3 (N2330, N2327, N619, N156);
not NOT1 (N2331, N2326);
nand NAND3 (N2332, N2329, N1884, N667);
or OR2 (N2333, N2323, N1421);
nand NAND2 (N2334, N2331, N1517);
not NOT1 (N2335, N2330);
and AND2 (N2336, N2335, N1605);
nor NOR3 (N2337, N2336, N1934, N1178);
nor NOR4 (N2338, N2310, N2174, N1534, N1005);
not NOT1 (N2339, N2328);
or OR3 (N2340, N2320, N2287, N187);
nand NAND3 (N2341, N2337, N2319, N490);
buf BUF1 (N2342, N2334);
or OR2 (N2343, N2325, N2233);
nor NOR2 (N2344, N2333, N1497);
and AND4 (N2345, N2338, N1445, N2086, N2228);
nor NOR4 (N2346, N2332, N809, N264, N2044);
nand NAND3 (N2347, N2342, N2250, N601);
nand NAND4 (N2348, N2341, N20, N552, N1757);
xor XOR2 (N2349, N2343, N2072);
and AND2 (N2350, N2349, N1412);
not NOT1 (N2351, N2313);
not NOT1 (N2352, N2316);
nand NAND2 (N2353, N2348, N368);
nor NOR4 (N2354, N2352, N1133, N2267, N1560);
buf BUF1 (N2355, N2347);
xor XOR2 (N2356, N2353, N518);
xor XOR2 (N2357, N2339, N1076);
nand NAND3 (N2358, N2345, N140, N76);
not NOT1 (N2359, N2354);
buf BUF1 (N2360, N2356);
xor XOR2 (N2361, N2351, N1334);
nand NAND4 (N2362, N2340, N1771, N152, N725);
buf BUF1 (N2363, N2359);
not NOT1 (N2364, N2358);
xor XOR2 (N2365, N2355, N1188);
xor XOR2 (N2366, N2363, N1236);
nand NAND2 (N2367, N2365, N1104);
or OR3 (N2368, N2360, N1295, N209);
not NOT1 (N2369, N2364);
xor XOR2 (N2370, N2362, N1568);
nand NAND3 (N2371, N2346, N1768, N1976);
or OR2 (N2372, N2350, N1539);
not NOT1 (N2373, N2371);
not NOT1 (N2374, N2344);
not NOT1 (N2375, N2370);
nor NOR2 (N2376, N2375, N2172);
or OR4 (N2377, N2372, N937, N1931, N1297);
or OR2 (N2378, N2377, N386);
nand NAND2 (N2379, N2369, N2083);
xor XOR2 (N2380, N2374, N166);
and AND4 (N2381, N2380, N1437, N267, N2200);
and AND2 (N2382, N2368, N350);
buf BUF1 (N2383, N2381);
nor NOR4 (N2384, N2367, N84, N243, N2162);
and AND2 (N2385, N2366, N750);
and AND2 (N2386, N2384, N198);
xor XOR2 (N2387, N2379, N862);
and AND2 (N2388, N2361, N925);
nand NAND3 (N2389, N2388, N881, N1774);
or OR2 (N2390, N2357, N813);
and AND2 (N2391, N2389, N1382);
nand NAND4 (N2392, N2378, N772, N954, N1502);
buf BUF1 (N2393, N2390);
buf BUF1 (N2394, N2385);
or OR3 (N2395, N2391, N1570, N267);
xor XOR2 (N2396, N2387, N1068);
or OR3 (N2397, N2394, N880, N2280);
or OR2 (N2398, N2386, N1754);
xor XOR2 (N2399, N2373, N652);
nor NOR2 (N2400, N2393, N447);
nor NOR4 (N2401, N2395, N598, N2210, N64);
and AND3 (N2402, N2383, N577, N1764);
nor NOR4 (N2403, N2398, N1594, N391, N1180);
and AND2 (N2404, N2396, N1828);
or OR4 (N2405, N2401, N1157, N77, N1220);
buf BUF1 (N2406, N2399);
xor XOR2 (N2407, N2392, N67);
not NOT1 (N2408, N2407);
buf BUF1 (N2409, N2402);
xor XOR2 (N2410, N2376, N1387);
or OR4 (N2411, N2400, N1182, N803, N989);
buf BUF1 (N2412, N2411);
nor NOR4 (N2413, N2382, N1416, N664, N156);
nor NOR3 (N2414, N2413, N1002, N2317);
nor NOR2 (N2415, N2409, N598);
nand NAND2 (N2416, N2397, N2112);
nand NAND2 (N2417, N2406, N1666);
or OR2 (N2418, N2414, N480);
nor NOR3 (N2419, N2415, N426, N1283);
nor NOR4 (N2420, N2416, N780, N1896, N62);
and AND2 (N2421, N2412, N81);
xor XOR2 (N2422, N2417, N2087);
nor NOR3 (N2423, N2418, N2351, N1614);
and AND3 (N2424, N2403, N464, N1734);
not NOT1 (N2425, N2421);
or OR3 (N2426, N2405, N1526, N254);
or OR3 (N2427, N2410, N225, N1149);
or OR3 (N2428, N2425, N515, N2036);
buf BUF1 (N2429, N2423);
xor XOR2 (N2430, N2408, N825);
and AND2 (N2431, N2428, N334);
buf BUF1 (N2432, N2430);
nor NOR2 (N2433, N2431, N1636);
nor NOR4 (N2434, N2419, N142, N585, N701);
xor XOR2 (N2435, N2427, N1791);
or OR4 (N2436, N2435, N2343, N336, N974);
not NOT1 (N2437, N2422);
not NOT1 (N2438, N2426);
nand NAND2 (N2439, N2434, N632);
nor NOR4 (N2440, N2433, N1709, N1804, N2204);
buf BUF1 (N2441, N2439);
and AND3 (N2442, N2432, N635, N1361);
nand NAND3 (N2443, N2437, N1268, N1459);
or OR4 (N2444, N2429, N934, N1612, N1461);
nand NAND4 (N2445, N2404, N1628, N1481, N1535);
xor XOR2 (N2446, N2438, N1230);
nor NOR2 (N2447, N2446, N640);
xor XOR2 (N2448, N2447, N137);
xor XOR2 (N2449, N2443, N1377);
buf BUF1 (N2450, N2441);
nand NAND2 (N2451, N2420, N966);
nor NOR3 (N2452, N2448, N2156, N1051);
and AND2 (N2453, N2451, N1742);
buf BUF1 (N2454, N2444);
nor NOR3 (N2455, N2445, N339, N1353);
xor XOR2 (N2456, N2453, N1744);
nor NOR4 (N2457, N2449, N3, N2070, N1726);
not NOT1 (N2458, N2436);
nor NOR4 (N2459, N2456, N2248, N998, N1989);
or OR3 (N2460, N2455, N28, N2059);
nand NAND2 (N2461, N2424, N1498);
nand NAND4 (N2462, N2459, N2173, N2113, N461);
or OR4 (N2463, N2457, N1626, N946, N2461);
or OR3 (N2464, N1946, N2297, N2355);
or OR2 (N2465, N2460, N1340);
nand NAND2 (N2466, N2452, N1954);
and AND3 (N2467, N2466, N757, N1372);
nor NOR4 (N2468, N2450, N1956, N1151, N149);
not NOT1 (N2469, N2463);
and AND2 (N2470, N2462, N1552);
and AND3 (N2471, N2458, N673, N1566);
xor XOR2 (N2472, N2471, N1709);
or OR4 (N2473, N2465, N1708, N19, N2172);
buf BUF1 (N2474, N2470);
buf BUF1 (N2475, N2464);
not NOT1 (N2476, N2473);
nand NAND3 (N2477, N2472, N551, N181);
nor NOR4 (N2478, N2469, N1255, N661, N987);
nor NOR3 (N2479, N2476, N147, N1325);
nor NOR2 (N2480, N2442, N527);
or OR2 (N2481, N2479, N2063);
or OR3 (N2482, N2475, N1282, N2145);
xor XOR2 (N2483, N2482, N1129);
or OR4 (N2484, N2478, N1842, N1991, N1083);
and AND3 (N2485, N2454, N450, N2025);
and AND2 (N2486, N2485, N2317);
nor NOR2 (N2487, N2481, N814);
nor NOR4 (N2488, N2467, N158, N2103, N300);
xor XOR2 (N2489, N2477, N1241);
xor XOR2 (N2490, N2488, N451);
and AND2 (N2491, N2487, N1999);
nor NOR3 (N2492, N2440, N2201, N800);
nand NAND2 (N2493, N2490, N966);
not NOT1 (N2494, N2484);
not NOT1 (N2495, N2492);
xor XOR2 (N2496, N2489, N1131);
buf BUF1 (N2497, N2494);
nand NAND3 (N2498, N2483, N10, N2447);
and AND3 (N2499, N2497, N40, N175);
or OR3 (N2500, N2493, N187, N2162);
nand NAND4 (N2501, N2499, N677, N2195, N2436);
xor XOR2 (N2502, N2500, N678);
xor XOR2 (N2503, N2468, N237);
or OR4 (N2504, N2496, N212, N1376, N1915);
xor XOR2 (N2505, N2498, N614);
nor NOR3 (N2506, N2486, N2114, N558);
or OR4 (N2507, N2506, N1214, N561, N377);
not NOT1 (N2508, N2480);
and AND3 (N2509, N2507, N1862, N1840);
or OR2 (N2510, N2503, N2020);
buf BUF1 (N2511, N2509);
or OR2 (N2512, N2505, N1477);
and AND4 (N2513, N2511, N1883, N2462, N1693);
not NOT1 (N2514, N2504);
xor XOR2 (N2515, N2495, N566);
buf BUF1 (N2516, N2513);
buf BUF1 (N2517, N2516);
and AND3 (N2518, N2491, N2011, N5);
buf BUF1 (N2519, N2515);
nand NAND3 (N2520, N2474, N1683, N1138);
and AND2 (N2521, N2518, N1160);
nor NOR4 (N2522, N2520, N1625, N743, N342);
nor NOR3 (N2523, N2501, N1475, N981);
nor NOR2 (N2524, N2523, N1969);
or OR3 (N2525, N2524, N456, N2470);
xor XOR2 (N2526, N2502, N2492);
nand NAND4 (N2527, N2526, N2400, N1914, N1721);
or OR3 (N2528, N2512, N1071, N1944);
nor NOR4 (N2529, N2510, N555, N1425, N1594);
nand NAND3 (N2530, N2519, N450, N1253);
buf BUF1 (N2531, N2527);
nor NOR4 (N2532, N2530, N1328, N205, N48);
and AND2 (N2533, N2508, N1459);
and AND4 (N2534, N2528, N1184, N289, N2023);
nor NOR4 (N2535, N2531, N1209, N1034, N681);
xor XOR2 (N2536, N2529, N89);
nor NOR4 (N2537, N2514, N2476, N742, N1547);
not NOT1 (N2538, N2532);
and AND3 (N2539, N2534, N2303, N1122);
buf BUF1 (N2540, N2533);
or OR2 (N2541, N2538, N1342);
not NOT1 (N2542, N2541);
or OR3 (N2543, N2522, N1815, N1087);
xor XOR2 (N2544, N2536, N1751);
and AND3 (N2545, N2517, N1388, N316);
xor XOR2 (N2546, N2537, N1358);
buf BUF1 (N2547, N2539);
not NOT1 (N2548, N2544);
nor NOR3 (N2549, N2542, N2214, N2275);
nand NAND3 (N2550, N2521, N1529, N552);
nor NOR3 (N2551, N2545, N99, N1590);
or OR2 (N2552, N2551, N443);
nor NOR2 (N2553, N2543, N844);
nand NAND4 (N2554, N2540, N1719, N67, N176);
not NOT1 (N2555, N2549);
not NOT1 (N2556, N2552);
and AND3 (N2557, N2553, N1130, N339);
xor XOR2 (N2558, N2556, N387);
buf BUF1 (N2559, N2554);
not NOT1 (N2560, N2548);
not NOT1 (N2561, N2550);
and AND2 (N2562, N2547, N723);
not NOT1 (N2563, N2562);
buf BUF1 (N2564, N2557);
and AND4 (N2565, N2560, N518, N2008, N1104);
and AND4 (N2566, N2561, N1504, N1786, N2105);
not NOT1 (N2567, N2565);
not NOT1 (N2568, N2564);
not NOT1 (N2569, N2568);
not NOT1 (N2570, N2546);
or OR3 (N2571, N2535, N1921, N1794);
buf BUF1 (N2572, N2571);
nand NAND3 (N2573, N2558, N1680, N1896);
nand NAND3 (N2574, N2573, N519, N625);
not NOT1 (N2575, N2525);
not NOT1 (N2576, N2559);
not NOT1 (N2577, N2555);
or OR4 (N2578, N2577, N527, N317, N2084);
or OR3 (N2579, N2566, N1649, N1307);
xor XOR2 (N2580, N2575, N1378);
nand NAND4 (N2581, N2574, N2048, N1806, N789);
not NOT1 (N2582, N2581);
nand NAND4 (N2583, N2576, N1218, N2412, N1549);
buf BUF1 (N2584, N2570);
nor NOR3 (N2585, N2582, N2580, N643);
not NOT1 (N2586, N490);
nor NOR4 (N2587, N2583, N1295, N2311, N1240);
nand NAND3 (N2588, N2563, N1485, N1726);
or OR3 (N2589, N2585, N896, N1755);
and AND4 (N2590, N2569, N1929, N1453, N2126);
buf BUF1 (N2591, N2584);
buf BUF1 (N2592, N2587);
xor XOR2 (N2593, N2592, N2280);
xor XOR2 (N2594, N2578, N1614);
not NOT1 (N2595, N2593);
nand NAND3 (N2596, N2586, N2337, N2395);
or OR3 (N2597, N2579, N1479, N460);
buf BUF1 (N2598, N2597);
and AND4 (N2599, N2594, N1860, N965, N1597);
nand NAND4 (N2600, N2590, N737, N657, N455);
or OR4 (N2601, N2595, N367, N1274, N1703);
not NOT1 (N2602, N2599);
buf BUF1 (N2603, N2567);
and AND2 (N2604, N2602, N1121);
nor NOR3 (N2605, N2603, N2278, N2479);
or OR3 (N2606, N2605, N809, N148);
nand NAND2 (N2607, N2601, N1865);
or OR4 (N2608, N2588, N1063, N228, N2290);
and AND3 (N2609, N2572, N170, N2193);
not NOT1 (N2610, N2606);
nor NOR4 (N2611, N2609, N242, N1090, N1147);
nor NOR2 (N2612, N2604, N1674);
and AND2 (N2613, N2607, N1045);
and AND2 (N2614, N2613, N1971);
nand NAND2 (N2615, N2612, N2344);
or OR2 (N2616, N2610, N1074);
xor XOR2 (N2617, N2598, N339);
nand NAND3 (N2618, N2591, N545, N2264);
xor XOR2 (N2619, N2617, N465);
buf BUF1 (N2620, N2619);
xor XOR2 (N2621, N2589, N4);
and AND2 (N2622, N2608, N640);
and AND4 (N2623, N2614, N10, N1692, N2388);
nand NAND3 (N2624, N2621, N1835, N1067);
not NOT1 (N2625, N2623);
and AND4 (N2626, N2596, N1271, N1376, N1120);
not NOT1 (N2627, N2625);
xor XOR2 (N2628, N2620, N13);
nand NAND4 (N2629, N2618, N1927, N1767, N2485);
xor XOR2 (N2630, N2622, N646);
buf BUF1 (N2631, N2600);
nand NAND3 (N2632, N2627, N699, N773);
buf BUF1 (N2633, N2628);
and AND3 (N2634, N2630, N1041, N615);
or OR4 (N2635, N2626, N534, N121, N422);
not NOT1 (N2636, N2611);
xor XOR2 (N2637, N2631, N1028);
buf BUF1 (N2638, N2629);
and AND2 (N2639, N2634, N2624);
nand NAND4 (N2640, N668, N2023, N2135, N1642);
and AND4 (N2641, N2636, N1372, N1208, N1118);
nor NOR2 (N2642, N2637, N2368);
nand NAND2 (N2643, N2615, N597);
nor NOR2 (N2644, N2643, N1068);
nor NOR3 (N2645, N2641, N160, N1337);
nor NOR3 (N2646, N2645, N2308, N635);
buf BUF1 (N2647, N2646);
buf BUF1 (N2648, N2640);
nor NOR2 (N2649, N2644, N694);
not NOT1 (N2650, N2638);
nand NAND4 (N2651, N2647, N772, N1588, N1769);
nor NOR2 (N2652, N2633, N2400);
nand NAND2 (N2653, N2639, N430);
not NOT1 (N2654, N2649);
not NOT1 (N2655, N2642);
not NOT1 (N2656, N2648);
nand NAND4 (N2657, N2650, N1029, N421, N2265);
buf BUF1 (N2658, N2657);
or OR2 (N2659, N2635, N994);
xor XOR2 (N2660, N2656, N1048);
nor NOR3 (N2661, N2616, N457, N575);
buf BUF1 (N2662, N2659);
xor XOR2 (N2663, N2662, N590);
nand NAND4 (N2664, N2651, N424, N2050, N1401);
nor NOR3 (N2665, N2664, N2029, N1940);
nor NOR2 (N2666, N2663, N1048);
buf BUF1 (N2667, N2653);
nand NAND4 (N2668, N2666, N74, N2132, N2206);
not NOT1 (N2669, N2667);
not NOT1 (N2670, N2669);
or OR4 (N2671, N2652, N1849, N1462, N544);
xor XOR2 (N2672, N2668, N1639);
not NOT1 (N2673, N2658);
xor XOR2 (N2674, N2670, N2133);
nand NAND3 (N2675, N2632, N370, N770);
buf BUF1 (N2676, N2660);
nor NOR4 (N2677, N2673, N1251, N1622, N692);
or OR2 (N2678, N2661, N2604);
xor XOR2 (N2679, N2672, N838);
xor XOR2 (N2680, N2679, N603);
xor XOR2 (N2681, N2678, N1080);
nand NAND3 (N2682, N2681, N941, N2133);
xor XOR2 (N2683, N2655, N391);
xor XOR2 (N2684, N2654, N1730);
and AND4 (N2685, N2680, N26, N2561, N2060);
and AND2 (N2686, N2674, N403);
nand NAND2 (N2687, N2686, N270);
and AND4 (N2688, N2685, N11, N1894, N2158);
buf BUF1 (N2689, N2688);
and AND3 (N2690, N2684, N501, N972);
or OR4 (N2691, N2676, N345, N1580, N2032);
buf BUF1 (N2692, N2683);
or OR2 (N2693, N2671, N672);
buf BUF1 (N2694, N2691);
buf BUF1 (N2695, N2687);
nor NOR4 (N2696, N2695, N763, N2336, N1462);
nor NOR3 (N2697, N2692, N1748, N1142);
not NOT1 (N2698, N2665);
nand NAND3 (N2699, N2697, N674, N313);
buf BUF1 (N2700, N2690);
or OR2 (N2701, N2693, N468);
and AND3 (N2702, N2696, N730, N1827);
not NOT1 (N2703, N2698);
buf BUF1 (N2704, N2675);
and AND4 (N2705, N2701, N694, N215, N662);
xor XOR2 (N2706, N2689, N1543);
nand NAND4 (N2707, N2702, N1822, N1655, N2548);
nand NAND3 (N2708, N2706, N1251, N1897);
not NOT1 (N2709, N2707);
buf BUF1 (N2710, N2700);
nor NOR3 (N2711, N2703, N529, N1096);
or OR2 (N2712, N2704, N220);
nand NAND2 (N2713, N2708, N669);
or OR2 (N2714, N2711, N2145);
nor NOR2 (N2715, N2710, N2622);
not NOT1 (N2716, N2682);
not NOT1 (N2717, N2716);
xor XOR2 (N2718, N2705, N1989);
or OR2 (N2719, N2694, N1448);
or OR4 (N2720, N2712, N1379, N1729, N1266);
nand NAND3 (N2721, N2709, N361, N511);
nor NOR4 (N2722, N2717, N478, N1473, N132);
nor NOR4 (N2723, N2720, N1022, N2637, N1327);
not NOT1 (N2724, N2721);
nand NAND2 (N2725, N2723, N533);
xor XOR2 (N2726, N2715, N850);
not NOT1 (N2727, N2718);
buf BUF1 (N2728, N2726);
not NOT1 (N2729, N2714);
buf BUF1 (N2730, N2722);
buf BUF1 (N2731, N2728);
xor XOR2 (N2732, N2724, N1198);
or OR4 (N2733, N2725, N2054, N378, N2282);
nor NOR2 (N2734, N2713, N2453);
or OR4 (N2735, N2730, N1455, N457, N1250);
nor NOR3 (N2736, N2727, N1303, N1812);
nor NOR4 (N2737, N2732, N1533, N1748, N2341);
xor XOR2 (N2738, N2699, N395);
xor XOR2 (N2739, N2729, N1583);
and AND4 (N2740, N2736, N961, N323, N2009);
not NOT1 (N2741, N2740);
not NOT1 (N2742, N2741);
nand NAND3 (N2743, N2735, N1742, N1072);
nand NAND3 (N2744, N2742, N2515, N1472);
nor NOR4 (N2745, N2677, N800, N19, N1265);
nor NOR2 (N2746, N2739, N342);
nor NOR4 (N2747, N2734, N2222, N499, N462);
or OR4 (N2748, N2743, N2184, N455, N2283);
nand NAND3 (N2749, N2731, N1571, N2102);
nor NOR4 (N2750, N2749, N23, N801, N235);
or OR3 (N2751, N2744, N1046, N2341);
buf BUF1 (N2752, N2748);
or OR4 (N2753, N2733, N2195, N1228, N987);
not NOT1 (N2754, N2737);
or OR3 (N2755, N2719, N292, N1640);
xor XOR2 (N2756, N2753, N567);
and AND3 (N2757, N2747, N1925, N1530);
nand NAND3 (N2758, N2738, N1042, N2644);
nand NAND4 (N2759, N2754, N1285, N1868, N708);
not NOT1 (N2760, N2757);
nor NOR3 (N2761, N2755, N1813, N1464);
xor XOR2 (N2762, N2759, N214);
and AND2 (N2763, N2752, N2109);
buf BUF1 (N2764, N2763);
nand NAND2 (N2765, N2758, N451);
buf BUF1 (N2766, N2751);
and AND2 (N2767, N2760, N401);
and AND4 (N2768, N2765, N978, N2304, N1295);
and AND3 (N2769, N2762, N27, N329);
xor XOR2 (N2770, N2745, N2013);
xor XOR2 (N2771, N2767, N1214);
buf BUF1 (N2772, N2761);
nand NAND4 (N2773, N2764, N2294, N1704, N686);
nor NOR3 (N2774, N2746, N770, N1264);
nor NOR4 (N2775, N2772, N1591, N250, N474);
nor NOR4 (N2776, N2773, N2321, N2721, N1437);
not NOT1 (N2777, N2768);
xor XOR2 (N2778, N2769, N253);
nor NOR4 (N2779, N2770, N2003, N2521, N554);
and AND3 (N2780, N2774, N451, N2470);
xor XOR2 (N2781, N2778, N2047);
and AND3 (N2782, N2781, N2259, N2419);
nand NAND3 (N2783, N2776, N105, N976);
buf BUF1 (N2784, N2783);
and AND3 (N2785, N2775, N999, N848);
xor XOR2 (N2786, N2756, N1961);
and AND3 (N2787, N2785, N1790, N491);
and AND3 (N2788, N2779, N2577, N1889);
or OR2 (N2789, N2750, N410);
buf BUF1 (N2790, N2784);
or OR2 (N2791, N2789, N2770);
xor XOR2 (N2792, N2786, N2338);
nand NAND2 (N2793, N2766, N2692);
buf BUF1 (N2794, N2787);
nor NOR2 (N2795, N2788, N2741);
nand NAND4 (N2796, N2780, N998, N1174, N715);
or OR3 (N2797, N2790, N1176, N1406);
or OR3 (N2798, N2771, N1548, N2232);
not NOT1 (N2799, N2796);
nor NOR3 (N2800, N2782, N2149, N746);
xor XOR2 (N2801, N2798, N48);
nand NAND3 (N2802, N2799, N657, N597);
and AND2 (N2803, N2802, N2470);
buf BUF1 (N2804, N2801);
nor NOR4 (N2805, N2791, N742, N1497, N1763);
buf BUF1 (N2806, N2800);
or OR2 (N2807, N2792, N1402);
or OR3 (N2808, N2777, N2376, N2513);
xor XOR2 (N2809, N2806, N1607);
and AND4 (N2810, N2808, N1746, N1461, N1052);
nand NAND2 (N2811, N2797, N1601);
and AND3 (N2812, N2805, N2151, N747);
or OR4 (N2813, N2809, N50, N1185, N1352);
nor NOR2 (N2814, N2795, N2102);
xor XOR2 (N2815, N2803, N1564);
and AND3 (N2816, N2815, N2408, N1194);
xor XOR2 (N2817, N2816, N2790);
not NOT1 (N2818, N2793);
nor NOR4 (N2819, N2811, N757, N1428, N201);
or OR4 (N2820, N2794, N346, N219, N873);
and AND3 (N2821, N2820, N1041, N2771);
or OR4 (N2822, N2804, N82, N32, N901);
nand NAND3 (N2823, N2822, N2118, N1904);
and AND3 (N2824, N2818, N849, N2311);
buf BUF1 (N2825, N2807);
or OR4 (N2826, N2812, N2589, N193, N2233);
buf BUF1 (N2827, N2813);
xor XOR2 (N2828, N2825, N2787);
buf BUF1 (N2829, N2819);
nand NAND2 (N2830, N2817, N636);
or OR2 (N2831, N2829, N944);
or OR2 (N2832, N2828, N780);
nand NAND3 (N2833, N2821, N565, N1679);
not NOT1 (N2834, N2824);
nor NOR3 (N2835, N2823, N1011, N33);
not NOT1 (N2836, N2827);
nand NAND2 (N2837, N2810, N370);
xor XOR2 (N2838, N2832, N698);
buf BUF1 (N2839, N2835);
nor NOR2 (N2840, N2826, N549);
nor NOR3 (N2841, N2834, N2390, N6);
nor NOR4 (N2842, N2840, N1347, N2544, N1097);
nand NAND3 (N2843, N2836, N1506, N2413);
buf BUF1 (N2844, N2841);
and AND4 (N2845, N2838, N2052, N1907, N2578);
nand NAND2 (N2846, N2833, N2453);
nand NAND3 (N2847, N2837, N1445, N632);
nand NAND4 (N2848, N2843, N560, N1759, N1338);
xor XOR2 (N2849, N2831, N1277);
or OR3 (N2850, N2814, N1264, N1001);
and AND4 (N2851, N2844, N1843, N541, N2809);
nor NOR4 (N2852, N2830, N1698, N1243, N1516);
buf BUF1 (N2853, N2851);
nor NOR4 (N2854, N2847, N2798, N590, N538);
and AND4 (N2855, N2839, N1472, N1639, N1739);
nor NOR4 (N2856, N2849, N856, N52, N837);
buf BUF1 (N2857, N2856);
nand NAND4 (N2858, N2854, N1767, N1429, N406);
nand NAND3 (N2859, N2852, N1620, N1648);
xor XOR2 (N2860, N2850, N378);
or OR3 (N2861, N2857, N2725, N126);
or OR3 (N2862, N2858, N1236, N589);
or OR3 (N2863, N2860, N2485, N2716);
nor NOR4 (N2864, N2861, N2207, N89, N463);
xor XOR2 (N2865, N2845, N1783);
buf BUF1 (N2866, N2865);
nand NAND4 (N2867, N2855, N693, N1180, N2701);
nand NAND4 (N2868, N2867, N2090, N2383, N2106);
nand NAND2 (N2869, N2853, N1274);
and AND2 (N2870, N2864, N1664);
nor NOR2 (N2871, N2848, N419);
or OR4 (N2872, N2846, N2047, N2379, N194);
and AND2 (N2873, N2863, N2239);
xor XOR2 (N2874, N2871, N109);
or OR2 (N2875, N2869, N828);
or OR2 (N2876, N2875, N848);
nor NOR3 (N2877, N2859, N2459, N2787);
xor XOR2 (N2878, N2842, N2755);
and AND4 (N2879, N2878, N1908, N320, N101);
not NOT1 (N2880, N2874);
or OR3 (N2881, N2862, N2237, N673);
buf BUF1 (N2882, N2880);
or OR2 (N2883, N2868, N2382);
xor XOR2 (N2884, N2870, N2863);
or OR4 (N2885, N2866, N1707, N790, N1137);
nand NAND2 (N2886, N2876, N773);
nor NOR3 (N2887, N2881, N2797, N1809);
and AND4 (N2888, N2884, N1055, N2611, N315);
buf BUF1 (N2889, N2877);
nand NAND4 (N2890, N2872, N1681, N33, N691);
xor XOR2 (N2891, N2886, N183);
and AND3 (N2892, N2888, N1480, N656);
buf BUF1 (N2893, N2890);
xor XOR2 (N2894, N2873, N367);
buf BUF1 (N2895, N2889);
and AND4 (N2896, N2883, N1306, N2476, N2867);
or OR3 (N2897, N2894, N2446, N55);
xor XOR2 (N2898, N2887, N1975);
nand NAND2 (N2899, N2891, N2292);
or OR3 (N2900, N2879, N53, N1309);
xor XOR2 (N2901, N2898, N756);
not NOT1 (N2902, N2896);
and AND3 (N2903, N2895, N200, N54);
nor NOR2 (N2904, N2902, N327);
not NOT1 (N2905, N2897);
and AND3 (N2906, N2904, N467, N1378);
buf BUF1 (N2907, N2893);
buf BUF1 (N2908, N2901);
and AND3 (N2909, N2899, N930, N946);
or OR4 (N2910, N2892, N1944, N2155, N878);
nor NOR2 (N2911, N2900, N1703);
or OR4 (N2912, N2882, N1209, N1159, N2892);
nor NOR4 (N2913, N2885, N1120, N2303, N1012);
and AND2 (N2914, N2903, N749);
nand NAND3 (N2915, N2908, N1952, N623);
buf BUF1 (N2916, N2913);
nor NOR4 (N2917, N2915, N317, N942, N1217);
buf BUF1 (N2918, N2912);
nand NAND3 (N2919, N2905, N1467, N2001);
nor NOR2 (N2920, N2906, N891);
buf BUF1 (N2921, N2910);
and AND3 (N2922, N2914, N569, N2911);
nor NOR3 (N2923, N1165, N2284, N1050);
and AND4 (N2924, N2907, N1749, N2662, N2262);
nand NAND3 (N2925, N2921, N853, N1800);
or OR4 (N2926, N2916, N1000, N1622, N1488);
buf BUF1 (N2927, N2925);
nor NOR4 (N2928, N2920, N2312, N2222, N668);
buf BUF1 (N2929, N2924);
and AND4 (N2930, N2917, N272, N1214, N106);
buf BUF1 (N2931, N2922);
xor XOR2 (N2932, N2923, N759);
not NOT1 (N2933, N2909);
nor NOR3 (N2934, N2929, N1857, N167);
not NOT1 (N2935, N2934);
nand NAND3 (N2936, N2930, N340, N2203);
nand NAND4 (N2937, N2935, N1217, N1726, N1048);
nor NOR2 (N2938, N2937, N335);
or OR4 (N2939, N2927, N574, N2899, N2910);
nor NOR2 (N2940, N2932, N1940);
and AND3 (N2941, N2938, N2099, N57);
not NOT1 (N2942, N2940);
xor XOR2 (N2943, N2928, N2542);
not NOT1 (N2944, N2942);
not NOT1 (N2945, N2944);
or OR4 (N2946, N2936, N2807, N2530, N640);
and AND3 (N2947, N2939, N1472, N304);
or OR2 (N2948, N2946, N310);
and AND2 (N2949, N2933, N2185);
xor XOR2 (N2950, N2945, N188);
nand NAND4 (N2951, N2941, N2710, N2656, N815);
nand NAND3 (N2952, N2950, N1692, N197);
nand NAND3 (N2953, N2943, N399, N588);
and AND4 (N2954, N2952, N580, N344, N399);
not NOT1 (N2955, N2931);
not NOT1 (N2956, N2926);
buf BUF1 (N2957, N2951);
and AND4 (N2958, N2948, N2848, N1611, N2008);
nand NAND3 (N2959, N2947, N1251, N2404);
xor XOR2 (N2960, N2956, N542);
and AND2 (N2961, N2918, N1595);
buf BUF1 (N2962, N2958);
or OR3 (N2963, N2959, N2251, N141);
or OR4 (N2964, N2963, N1451, N1748, N2697);
xor XOR2 (N2965, N2955, N254);
xor XOR2 (N2966, N2949, N365);
and AND2 (N2967, N2960, N2718);
or OR2 (N2968, N2953, N1859);
nand NAND2 (N2969, N2919, N1773);
nand NAND2 (N2970, N2967, N1726);
nor NOR2 (N2971, N2962, N1677);
nor NOR4 (N2972, N2961, N874, N66, N815);
buf BUF1 (N2973, N2966);
not NOT1 (N2974, N2954);
xor XOR2 (N2975, N2973, N1628);
buf BUF1 (N2976, N2970);
or OR4 (N2977, N2972, N1701, N762, N1686);
not NOT1 (N2978, N2957);
and AND2 (N2979, N2977, N2788);
xor XOR2 (N2980, N2976, N1057);
or OR2 (N2981, N2975, N2885);
and AND4 (N2982, N2969, N2827, N2723, N534);
nand NAND2 (N2983, N2968, N2796);
not NOT1 (N2984, N2978);
not NOT1 (N2985, N2974);
nand NAND2 (N2986, N2971, N735);
nand NAND4 (N2987, N2982, N1553, N1586, N1090);
nor NOR2 (N2988, N2983, N2746);
nand NAND4 (N2989, N2985, N1503, N1237, N2300);
xor XOR2 (N2990, N2965, N2480);
nand NAND4 (N2991, N2984, N227, N360, N283);
buf BUF1 (N2992, N2987);
nand NAND3 (N2993, N2992, N2694, N2622);
nand NAND4 (N2994, N2980, N1805, N1315, N2892);
nor NOR4 (N2995, N2989, N2272, N1969, N323);
not NOT1 (N2996, N2995);
not NOT1 (N2997, N2979);
or OR2 (N2998, N2981, N2923);
and AND4 (N2999, N2986, N2160, N1859, N899);
and AND2 (N3000, N2990, N2735);
nor NOR2 (N3001, N2988, N1767);
nor NOR4 (N3002, N2964, N1014, N2452, N986);
nand NAND3 (N3003, N2993, N456, N2380);
or OR3 (N3004, N2999, N2811, N171);
nand NAND4 (N3005, N3003, N1453, N888, N1095);
nor NOR2 (N3006, N2991, N2539);
nor NOR3 (N3007, N2997, N1950, N166);
nand NAND4 (N3008, N3005, N229, N506, N555);
nand NAND3 (N3009, N3004, N874, N1022);
or OR3 (N3010, N2996, N735, N2477);
nor NOR4 (N3011, N3008, N2853, N587, N2625);
buf BUF1 (N3012, N3009);
or OR3 (N3013, N3011, N969, N1181);
buf BUF1 (N3014, N2994);
buf BUF1 (N3015, N3002);
xor XOR2 (N3016, N3012, N1244);
xor XOR2 (N3017, N3015, N1395);
xor XOR2 (N3018, N3007, N1677);
or OR2 (N3019, N3000, N754);
not NOT1 (N3020, N3013);
buf BUF1 (N3021, N3006);
and AND4 (N3022, N3019, N2610, N1443, N2089);
nor NOR4 (N3023, N3010, N621, N994, N2157);
not NOT1 (N3024, N3023);
not NOT1 (N3025, N2998);
and AND2 (N3026, N3024, N2842);
not NOT1 (N3027, N3018);
not NOT1 (N3028, N3014);
nand NAND2 (N3029, N3020, N2578);
or OR3 (N3030, N3021, N522, N1676);
not NOT1 (N3031, N3026);
or OR3 (N3032, N3027, N2100, N2454);
nand NAND2 (N3033, N3029, N1697);
or OR4 (N3034, N3033, N1948, N797, N1040);
nor NOR2 (N3035, N3030, N1647);
not NOT1 (N3036, N3022);
or OR3 (N3037, N3025, N173, N439);
nor NOR4 (N3038, N3037, N1367, N2713, N2154);
nand NAND2 (N3039, N3035, N529);
or OR2 (N3040, N3034, N181);
or OR4 (N3041, N3040, N402, N139, N2817);
nor NOR4 (N3042, N3031, N1830, N894, N2794);
or OR4 (N3043, N3036, N2116, N1829, N2292);
or OR3 (N3044, N3001, N2541, N2736);
not NOT1 (N3045, N3044);
not NOT1 (N3046, N3041);
and AND4 (N3047, N3028, N959, N2814, N1847);
not NOT1 (N3048, N3017);
buf BUF1 (N3049, N3016);
xor XOR2 (N3050, N3042, N1079);
and AND2 (N3051, N3049, N1847);
not NOT1 (N3052, N3043);
or OR2 (N3053, N3045, N527);
xor XOR2 (N3054, N3050, N2162);
and AND3 (N3055, N3052, N782, N57);
not NOT1 (N3056, N3048);
nor NOR3 (N3057, N3051, N1615, N885);
xor XOR2 (N3058, N3053, N1937);
nand NAND3 (N3059, N3039, N1120, N1147);
xor XOR2 (N3060, N3038, N1681);
not NOT1 (N3061, N3060);
nand NAND3 (N3062, N3057, N397, N900);
buf BUF1 (N3063, N3062);
not NOT1 (N3064, N3059);
and AND3 (N3065, N3032, N1267, N236);
or OR4 (N3066, N3046, N1024, N756, N2428);
xor XOR2 (N3067, N3061, N1329);
and AND4 (N3068, N3065, N165, N2255, N401);
not NOT1 (N3069, N3055);
and AND4 (N3070, N3063, N1055, N1283, N402);
nor NOR3 (N3071, N3064, N715, N1842);
xor XOR2 (N3072, N3069, N1864);
not NOT1 (N3073, N3058);
nand NAND3 (N3074, N3068, N909, N2393);
not NOT1 (N3075, N3074);
nand NAND3 (N3076, N3071, N1658, N1510);
buf BUF1 (N3077, N3070);
buf BUF1 (N3078, N3056);
or OR3 (N3079, N3067, N3077, N2966);
buf BUF1 (N3080, N151);
not NOT1 (N3081, N3066);
nand NAND2 (N3082, N3081, N2854);
nand NAND2 (N3083, N3072, N2547);
nand NAND2 (N3084, N3054, N1472);
nor NOR2 (N3085, N3078, N2701);
or OR3 (N3086, N3085, N1224, N1937);
nand NAND3 (N3087, N3086, N2208, N2808);
and AND3 (N3088, N3082, N2322, N834);
not NOT1 (N3089, N3075);
nor NOR3 (N3090, N3089, N1878, N2095);
or OR2 (N3091, N3090, N2898);
not NOT1 (N3092, N3076);
xor XOR2 (N3093, N3079, N2902);
buf BUF1 (N3094, N3083);
and AND3 (N3095, N3080, N2491, N238);
or OR2 (N3096, N3093, N5);
or OR3 (N3097, N3088, N1265, N1390);
and AND2 (N3098, N3047, N2963);
not NOT1 (N3099, N3094);
xor XOR2 (N3100, N3099, N1759);
nor NOR2 (N3101, N3097, N136);
buf BUF1 (N3102, N3095);
or OR2 (N3103, N3087, N2502);
nor NOR3 (N3104, N3073, N429, N2472);
not NOT1 (N3105, N3098);
and AND4 (N3106, N3084, N1742, N701, N3071);
xor XOR2 (N3107, N3096, N1369);
or OR4 (N3108, N3101, N2387, N639, N1688);
buf BUF1 (N3109, N3091);
xor XOR2 (N3110, N3106, N61);
nor NOR2 (N3111, N3103, N1290);
and AND4 (N3112, N3111, N419, N2209, N2373);
buf BUF1 (N3113, N3109);
or OR4 (N3114, N3107, N2068, N2413, N2372);
buf BUF1 (N3115, N3105);
buf BUF1 (N3116, N3102);
nor NOR4 (N3117, N3115, N2568, N1476, N2227);
not NOT1 (N3118, N3113);
nand NAND4 (N3119, N3117, N2481, N108, N1567);
nor NOR2 (N3120, N3092, N553);
or OR4 (N3121, N3119, N2079, N2075, N2714);
nand NAND3 (N3122, N3104, N712, N120);
not NOT1 (N3123, N3110);
nand NAND3 (N3124, N3100, N1702, N2531);
xor XOR2 (N3125, N3122, N207);
xor XOR2 (N3126, N3123, N2486);
nor NOR4 (N3127, N3126, N2416, N313, N2956);
nand NAND4 (N3128, N3108, N2675, N620, N2318);
nand NAND3 (N3129, N3114, N2035, N414);
xor XOR2 (N3130, N3127, N1480);
xor XOR2 (N3131, N3125, N2012);
nor NOR2 (N3132, N3120, N1969);
not NOT1 (N3133, N3116);
nor NOR3 (N3134, N3133, N3068, N621);
not NOT1 (N3135, N3128);
and AND3 (N3136, N3130, N3062, N809);
buf BUF1 (N3137, N3132);
not NOT1 (N3138, N3118);
not NOT1 (N3139, N3134);
buf BUF1 (N3140, N3121);
or OR2 (N3141, N3138, N1982);
not NOT1 (N3142, N3131);
not NOT1 (N3143, N3141);
xor XOR2 (N3144, N3137, N1746);
nand NAND4 (N3145, N3124, N2965, N2190, N1232);
and AND3 (N3146, N3143, N2489, N1143);
xor XOR2 (N3147, N3146, N423);
nand NAND3 (N3148, N3142, N2082, N2707);
not NOT1 (N3149, N3139);
nand NAND2 (N3150, N3147, N3025);
nand NAND3 (N3151, N3144, N1209, N3119);
nor NOR3 (N3152, N3140, N653, N3059);
not NOT1 (N3153, N3152);
and AND2 (N3154, N3145, N2866);
and AND3 (N3155, N3149, N1563, N354);
buf BUF1 (N3156, N3129);
and AND4 (N3157, N3154, N366, N2228, N1314);
not NOT1 (N3158, N3155);
nor NOR4 (N3159, N3158, N2023, N1764, N806);
nor NOR3 (N3160, N3150, N2859, N239);
nor NOR4 (N3161, N3160, N550, N525, N734);
not NOT1 (N3162, N3157);
or OR3 (N3163, N3159, N1871, N306);
and AND4 (N3164, N3163, N909, N703, N1342);
or OR4 (N3165, N3164, N443, N1530, N31);
nand NAND4 (N3166, N3136, N431, N1752, N3062);
or OR3 (N3167, N3148, N1811, N1362);
or OR2 (N3168, N3165, N2368);
nand NAND4 (N3169, N3153, N842, N2281, N349);
or OR4 (N3170, N3156, N2777, N262, N2902);
nor NOR4 (N3171, N3135, N2932, N1226, N1669);
nand NAND3 (N3172, N3170, N1013, N595);
xor XOR2 (N3173, N3171, N2312);
nand NAND2 (N3174, N3161, N1294);
nand NAND3 (N3175, N3166, N2644, N2794);
not NOT1 (N3176, N3167);
nor NOR3 (N3177, N3151, N1431, N476);
not NOT1 (N3178, N3112);
nor NOR3 (N3179, N3175, N2781, N1890);
nand NAND4 (N3180, N3179, N1472, N2350, N53);
buf BUF1 (N3181, N3180);
not NOT1 (N3182, N3177);
and AND2 (N3183, N3162, N3087);
xor XOR2 (N3184, N3183, N1712);
or OR4 (N3185, N3176, N88, N911, N3008);
and AND2 (N3186, N3172, N2422);
nor NOR4 (N3187, N3173, N2963, N1905, N1134);
nand NAND3 (N3188, N3182, N1494, N64);
not NOT1 (N3189, N3184);
xor XOR2 (N3190, N3189, N1879);
nand NAND2 (N3191, N3181, N4);
or OR2 (N3192, N3186, N2011);
nand NAND4 (N3193, N3178, N858, N1379, N963);
and AND4 (N3194, N3174, N309, N1182, N888);
buf BUF1 (N3195, N3194);
or OR2 (N3196, N3193, N1192);
nand NAND4 (N3197, N3196, N890, N2163, N1841);
not NOT1 (N3198, N3191);
buf BUF1 (N3199, N3190);
and AND3 (N3200, N3192, N2163, N1047);
not NOT1 (N3201, N3188);
nor NOR3 (N3202, N3201, N2357, N509);
or OR2 (N3203, N3197, N1059);
xor XOR2 (N3204, N3202, N3194);
not NOT1 (N3205, N3200);
and AND2 (N3206, N3195, N318);
nand NAND4 (N3207, N3203, N1050, N1555, N3079);
buf BUF1 (N3208, N3198);
not NOT1 (N3209, N3187);
buf BUF1 (N3210, N3209);
and AND2 (N3211, N3206, N2847);
nor NOR4 (N3212, N3185, N1017, N2296, N2872);
not NOT1 (N3213, N3199);
nor NOR3 (N3214, N3204, N3026, N2374);
buf BUF1 (N3215, N3212);
buf BUF1 (N3216, N3213);
or OR4 (N3217, N3168, N1771, N3012, N3137);
or OR4 (N3218, N3205, N2963, N2112, N1596);
buf BUF1 (N3219, N3214);
buf BUF1 (N3220, N3207);
or OR2 (N3221, N3215, N2920);
nand NAND4 (N3222, N3219, N1251, N1824, N1464);
xor XOR2 (N3223, N3221, N2467);
or OR3 (N3224, N3222, N541, N235);
buf BUF1 (N3225, N3224);
or OR4 (N3226, N3217, N3212, N2690, N1431);
or OR4 (N3227, N3218, N2421, N1645, N1414);
nor NOR3 (N3228, N3216, N2924, N1104);
and AND3 (N3229, N3208, N1347, N2246);
xor XOR2 (N3230, N3220, N3025);
buf BUF1 (N3231, N3169);
nor NOR2 (N3232, N3225, N803);
and AND4 (N3233, N3232, N3002, N1950, N320);
buf BUF1 (N3234, N3210);
nor NOR4 (N3235, N3226, N2499, N1804, N2072);
and AND3 (N3236, N3227, N3005, N106);
nor NOR3 (N3237, N3233, N766, N2662);
nor NOR4 (N3238, N3223, N591, N1758, N444);
not NOT1 (N3239, N3234);
or OR2 (N3240, N3239, N252);
xor XOR2 (N3241, N3235, N2816);
and AND3 (N3242, N3211, N2850, N830);
nor NOR2 (N3243, N3230, N2528);
not NOT1 (N3244, N3242);
not NOT1 (N3245, N3244);
and AND2 (N3246, N3231, N1851);
not NOT1 (N3247, N3243);
xor XOR2 (N3248, N3237, N935);
and AND4 (N3249, N3246, N2214, N841, N3188);
nor NOR3 (N3250, N3240, N2171, N1390);
and AND2 (N3251, N3229, N2685);
not NOT1 (N3252, N3238);
nand NAND2 (N3253, N3247, N2595);
xor XOR2 (N3254, N3249, N2459);
xor XOR2 (N3255, N3228, N2503);
not NOT1 (N3256, N3236);
and AND4 (N3257, N3255, N2092, N364, N2963);
not NOT1 (N3258, N3254);
nor NOR2 (N3259, N3253, N2905);
xor XOR2 (N3260, N3241, N1685);
not NOT1 (N3261, N3257);
xor XOR2 (N3262, N3245, N2199);
nand NAND2 (N3263, N3259, N342);
or OR3 (N3264, N3261, N842, N1217);
buf BUF1 (N3265, N3252);
or OR2 (N3266, N3256, N536);
buf BUF1 (N3267, N3250);
xor XOR2 (N3268, N3248, N113);
not NOT1 (N3269, N3264);
or OR4 (N3270, N3266, N2712, N1034, N1127);
and AND3 (N3271, N3269, N157, N2206);
or OR4 (N3272, N3262, N1114, N613, N688);
nand NAND4 (N3273, N3272, N1063, N28, N1495);
and AND2 (N3274, N3258, N174);
nand NAND2 (N3275, N3270, N1434);
or OR2 (N3276, N3260, N3177);
nor NOR4 (N3277, N3275, N1766, N279, N2603);
or OR3 (N3278, N3263, N2130, N846);
not NOT1 (N3279, N3251);
nand NAND3 (N3280, N3277, N1993, N758);
xor XOR2 (N3281, N3273, N273);
buf BUF1 (N3282, N3271);
buf BUF1 (N3283, N3267);
xor XOR2 (N3284, N3265, N2302);
buf BUF1 (N3285, N3283);
nor NOR4 (N3286, N3274, N1907, N1843, N1039);
xor XOR2 (N3287, N3268, N1694);
and AND4 (N3288, N3281, N975, N2704, N1344);
xor XOR2 (N3289, N3279, N2520);
or OR4 (N3290, N3276, N761, N745, N1501);
nand NAND3 (N3291, N3288, N2824, N1845);
nor NOR4 (N3292, N3280, N2123, N627, N3018);
and AND4 (N3293, N3292, N2309, N1355, N1940);
and AND3 (N3294, N3278, N2773, N2801);
and AND4 (N3295, N3289, N2845, N3118, N916);
nor NOR4 (N3296, N3290, N3058, N627, N414);
not NOT1 (N3297, N3294);
or OR4 (N3298, N3297, N826, N1655, N466);
nor NOR4 (N3299, N3291, N291, N1268, N1107);
or OR3 (N3300, N3285, N1085, N585);
nand NAND4 (N3301, N3287, N3127, N828, N2020);
not NOT1 (N3302, N3284);
not NOT1 (N3303, N3293);
buf BUF1 (N3304, N3300);
or OR3 (N3305, N3302, N1944, N2162);
or OR4 (N3306, N3286, N3235, N1564, N2984);
buf BUF1 (N3307, N3306);
or OR4 (N3308, N3282, N2347, N2370, N1247);
not NOT1 (N3309, N3304);
nor NOR2 (N3310, N3307, N145);
xor XOR2 (N3311, N3310, N1051);
nor NOR3 (N3312, N3309, N2291, N2514);
xor XOR2 (N3313, N3299, N50);
not NOT1 (N3314, N3308);
and AND3 (N3315, N3296, N457, N2596);
xor XOR2 (N3316, N3298, N293);
or OR4 (N3317, N3295, N2880, N317, N1271);
or OR4 (N3318, N3317, N1277, N1581, N577);
and AND2 (N3319, N3301, N1128);
nor NOR3 (N3320, N3316, N165, N1488);
nand NAND4 (N3321, N3305, N2831, N2003, N2886);
xor XOR2 (N3322, N3318, N2843);
xor XOR2 (N3323, N3314, N2664);
nor NOR2 (N3324, N3311, N115);
or OR3 (N3325, N3313, N1866, N2268);
nand NAND4 (N3326, N3312, N11, N37, N583);
xor XOR2 (N3327, N3321, N380);
and AND3 (N3328, N3319, N297, N2423);
and AND2 (N3329, N3325, N81);
nand NAND2 (N3330, N3324, N1468);
and AND4 (N3331, N3326, N74, N1876, N91);
not NOT1 (N3332, N3320);
or OR3 (N3333, N3328, N1675, N2321);
buf BUF1 (N3334, N3331);
and AND4 (N3335, N3330, N1761, N1230, N51);
nor NOR4 (N3336, N3329, N1944, N3294, N2187);
and AND3 (N3337, N3335, N3289, N1981);
and AND3 (N3338, N3337, N1723, N852);
nand NAND2 (N3339, N3323, N2451);
xor XOR2 (N3340, N3336, N1686);
and AND2 (N3341, N3338, N1306);
or OR2 (N3342, N3327, N1114);
buf BUF1 (N3343, N3332);
xor XOR2 (N3344, N3334, N391);
xor XOR2 (N3345, N3315, N765);
and AND2 (N3346, N3340, N167);
buf BUF1 (N3347, N3341);
not NOT1 (N3348, N3303);
nand NAND4 (N3349, N3345, N1113, N2594, N2403);
buf BUF1 (N3350, N3339);
nor NOR3 (N3351, N3322, N188, N99);
nand NAND2 (N3352, N3343, N1189);
nand NAND2 (N3353, N3347, N2037);
or OR3 (N3354, N3333, N2995, N1186);
not NOT1 (N3355, N3352);
and AND3 (N3356, N3351, N948, N317);
nand NAND2 (N3357, N3356, N883);
nand NAND4 (N3358, N3354, N1574, N3222, N1202);
nand NAND4 (N3359, N3348, N2282, N554, N589);
xor XOR2 (N3360, N3349, N1706);
nor NOR3 (N3361, N3344, N2039, N2405);
and AND3 (N3362, N3359, N957, N2389);
nand NAND2 (N3363, N3350, N1250);
xor XOR2 (N3364, N3358, N2231);
nand NAND4 (N3365, N3364, N2475, N1798, N2044);
xor XOR2 (N3366, N3362, N3323);
nand NAND3 (N3367, N3355, N2394, N2994);
or OR3 (N3368, N3363, N3005, N821);
not NOT1 (N3369, N3357);
xor XOR2 (N3370, N3366, N956);
buf BUF1 (N3371, N3368);
buf BUF1 (N3372, N3369);
or OR3 (N3373, N3371, N2593, N880);
not NOT1 (N3374, N3353);
xor XOR2 (N3375, N3374, N838);
nor NOR4 (N3376, N3365, N997, N389, N1453);
nand NAND2 (N3377, N3373, N3241);
nand NAND3 (N3378, N3360, N1815, N141);
nand NAND4 (N3379, N3370, N2254, N910, N1788);
not NOT1 (N3380, N3379);
xor XOR2 (N3381, N3372, N2042);
not NOT1 (N3382, N3377);
nand NAND3 (N3383, N3376, N1930, N2063);
buf BUF1 (N3384, N3367);
nor NOR3 (N3385, N3382, N107, N377);
and AND4 (N3386, N3383, N2365, N2813, N1627);
or OR3 (N3387, N3380, N1441, N1274);
nor NOR4 (N3388, N3342, N2819, N2851, N411);
not NOT1 (N3389, N3375);
buf BUF1 (N3390, N3389);
buf BUF1 (N3391, N3384);
or OR2 (N3392, N3391, N2418);
or OR2 (N3393, N3387, N2419);
buf BUF1 (N3394, N3388);
not NOT1 (N3395, N3394);
xor XOR2 (N3396, N3386, N476);
not NOT1 (N3397, N3395);
not NOT1 (N3398, N3385);
not NOT1 (N3399, N3397);
xor XOR2 (N3400, N3390, N2346);
buf BUF1 (N3401, N3392);
not NOT1 (N3402, N3401);
xor XOR2 (N3403, N3361, N1034);
and AND2 (N3404, N3403, N144);
not NOT1 (N3405, N3396);
xor XOR2 (N3406, N3393, N3320);
nand NAND3 (N3407, N3346, N3252, N892);
buf BUF1 (N3408, N3402);
and AND2 (N3409, N3400, N2456);
xor XOR2 (N3410, N3407, N2807);
not NOT1 (N3411, N3405);
not NOT1 (N3412, N3381);
not NOT1 (N3413, N3378);
or OR4 (N3414, N3410, N2623, N2224, N567);
nor NOR4 (N3415, N3398, N2284, N2138, N2845);
xor XOR2 (N3416, N3414, N2573);
not NOT1 (N3417, N3399);
xor XOR2 (N3418, N3415, N2804);
nor NOR3 (N3419, N3412, N3085, N3019);
nor NOR4 (N3420, N3416, N2410, N1876, N1016);
xor XOR2 (N3421, N3413, N3074);
nand NAND2 (N3422, N3406, N2784);
and AND4 (N3423, N3409, N968, N1872, N2401);
nand NAND3 (N3424, N3417, N135, N623);
or OR4 (N3425, N3418, N2398, N674, N956);
buf BUF1 (N3426, N3420);
or OR2 (N3427, N3425, N1133);
buf BUF1 (N3428, N3411);
xor XOR2 (N3429, N3427, N1628);
and AND3 (N3430, N3404, N1688, N45);
or OR3 (N3431, N3424, N3415, N652);
nand NAND4 (N3432, N3421, N2140, N890, N458);
and AND3 (N3433, N3430, N1582, N418);
nor NOR2 (N3434, N3429, N1408);
and AND2 (N3435, N3434, N1790);
nand NAND3 (N3436, N3423, N1536, N1107);
nor NOR3 (N3437, N3435, N1224, N3011);
and AND3 (N3438, N3436, N973, N1283);
nor NOR3 (N3439, N3408, N369, N2485);
xor XOR2 (N3440, N3437, N2049);
or OR4 (N3441, N3438, N487, N2477, N3251);
not NOT1 (N3442, N3433);
or OR4 (N3443, N3428, N2428, N1329, N695);
buf BUF1 (N3444, N3432);
and AND2 (N3445, N3431, N726);
buf BUF1 (N3446, N3443);
nor NOR4 (N3447, N3446, N3044, N3124, N775);
nor NOR4 (N3448, N3444, N2848, N513, N978);
nand NAND2 (N3449, N3447, N240);
or OR4 (N3450, N3440, N337, N1433, N556);
buf BUF1 (N3451, N3448);
and AND3 (N3452, N3442, N1777, N1681);
nand NAND4 (N3453, N3452, N2307, N2050, N478);
buf BUF1 (N3454, N3439);
or OR2 (N3455, N3441, N2953);
buf BUF1 (N3456, N3419);
nor NOR4 (N3457, N3456, N1103, N531, N3350);
and AND3 (N3458, N3457, N2701, N1445);
and AND3 (N3459, N3426, N2370, N331);
xor XOR2 (N3460, N3422, N1926);
not NOT1 (N3461, N3453);
not NOT1 (N3462, N3449);
not NOT1 (N3463, N3451);
nor NOR4 (N3464, N3460, N1529, N1653, N3371);
xor XOR2 (N3465, N3462, N2215);
buf BUF1 (N3466, N3459);
buf BUF1 (N3467, N3463);
xor XOR2 (N3468, N3465, N264);
nand NAND4 (N3469, N3467, N1683, N1894, N1208);
buf BUF1 (N3470, N3450);
and AND2 (N3471, N3455, N3387);
nor NOR4 (N3472, N3471, N3035, N2375, N825);
or OR2 (N3473, N3472, N1598);
nand NAND4 (N3474, N3461, N2301, N1896, N422);
not NOT1 (N3475, N3458);
or OR2 (N3476, N3475, N741);
or OR4 (N3477, N3468, N1008, N1526, N3312);
and AND4 (N3478, N3464, N558, N3265, N1517);
buf BUF1 (N3479, N3473);
nor NOR3 (N3480, N3454, N3466, N1911);
or OR4 (N3481, N2100, N1838, N260, N2633);
nor NOR3 (N3482, N3480, N1129, N9);
not NOT1 (N3483, N3481);
not NOT1 (N3484, N3478);
nand NAND2 (N3485, N3484, N291);
nor NOR4 (N3486, N3469, N2860, N1790, N1072);
xor XOR2 (N3487, N3476, N1180);
not NOT1 (N3488, N3486);
nor NOR4 (N3489, N3485, N320, N2845, N380);
buf BUF1 (N3490, N3445);
and AND2 (N3491, N3474, N929);
xor XOR2 (N3492, N3488, N199);
buf BUF1 (N3493, N3470);
or OR3 (N3494, N3483, N631, N1334);
buf BUF1 (N3495, N3487);
buf BUF1 (N3496, N3482);
and AND4 (N3497, N3495, N2458, N2277, N2275);
xor XOR2 (N3498, N3497, N1422);
and AND3 (N3499, N3498, N2582, N2944);
nor NOR3 (N3500, N3491, N2653, N3298);
or OR2 (N3501, N3493, N3269);
and AND4 (N3502, N3500, N3348, N2172, N889);
nor NOR4 (N3503, N3496, N3452, N945, N3126);
not NOT1 (N3504, N3492);
buf BUF1 (N3505, N3490);
buf BUF1 (N3506, N3477);
xor XOR2 (N3507, N3504, N2876);
and AND2 (N3508, N3489, N2830);
not NOT1 (N3509, N3503);
nor NOR4 (N3510, N3479, N655, N774, N365);
nand NAND2 (N3511, N3505, N2106);
and AND2 (N3512, N3501, N2207);
xor XOR2 (N3513, N3506, N2102);
or OR3 (N3514, N3502, N2064, N935);
not NOT1 (N3515, N3507);
nor NOR2 (N3516, N3499, N2071);
buf BUF1 (N3517, N3516);
nor NOR4 (N3518, N3512, N680, N2358, N1757);
not NOT1 (N3519, N3510);
buf BUF1 (N3520, N3519);
xor XOR2 (N3521, N3494, N2005);
or OR3 (N3522, N3520, N2535, N1159);
or OR2 (N3523, N3515, N1498);
xor XOR2 (N3524, N3514, N1686);
xor XOR2 (N3525, N3518, N2895);
buf BUF1 (N3526, N3525);
or OR3 (N3527, N3517, N3133, N2589);
xor XOR2 (N3528, N3513, N3060);
xor XOR2 (N3529, N3521, N2683);
or OR3 (N3530, N3529, N2519, N3462);
xor XOR2 (N3531, N3508, N472);
nor NOR4 (N3532, N3531, N1589, N2286, N2689);
nand NAND3 (N3533, N3532, N1366, N1609);
or OR3 (N3534, N3509, N225, N2204);
nand NAND2 (N3535, N3522, N852);
not NOT1 (N3536, N3534);
nor NOR3 (N3537, N3528, N2079, N3479);
and AND4 (N3538, N3511, N1414, N1974, N3049);
nand NAND4 (N3539, N3537, N3056, N2640, N1303);
not NOT1 (N3540, N3523);
nor NOR4 (N3541, N3539, N1862, N2167, N1685);
nor NOR4 (N3542, N3533, N1312, N1431, N87);
nand NAND3 (N3543, N3526, N100, N2214);
buf BUF1 (N3544, N3527);
xor XOR2 (N3545, N3524, N903);
not NOT1 (N3546, N3544);
not NOT1 (N3547, N3546);
nor NOR4 (N3548, N3541, N485, N1506, N3394);
not NOT1 (N3549, N3536);
nand NAND4 (N3550, N3545, N3385, N1041, N653);
xor XOR2 (N3551, N3543, N1318);
and AND3 (N3552, N3535, N2890, N1935);
buf BUF1 (N3553, N3547);
nand NAND2 (N3554, N3540, N347);
xor XOR2 (N3555, N3538, N1597);
xor XOR2 (N3556, N3549, N1911);
and AND3 (N3557, N3542, N2321, N1178);
nor NOR2 (N3558, N3530, N2215);
or OR3 (N3559, N3556, N409, N2002);
or OR2 (N3560, N3553, N3220);
not NOT1 (N3561, N3559);
xor XOR2 (N3562, N3561, N3214);
not NOT1 (N3563, N3558);
nand NAND3 (N3564, N3563, N2992, N3427);
or OR3 (N3565, N3562, N962, N1493);
and AND2 (N3566, N3560, N1110);
xor XOR2 (N3567, N3550, N1589);
buf BUF1 (N3568, N3554);
or OR3 (N3569, N3567, N3219, N1047);
buf BUF1 (N3570, N3566);
buf BUF1 (N3571, N3570);
or OR2 (N3572, N3552, N154);
xor XOR2 (N3573, N3568, N2876);
and AND4 (N3574, N3557, N2587, N73, N550);
xor XOR2 (N3575, N3574, N2903);
nand NAND2 (N3576, N3564, N873);
not NOT1 (N3577, N3571);
xor XOR2 (N3578, N3577, N2087);
not NOT1 (N3579, N3572);
nand NAND4 (N3580, N3579, N3223, N310, N3356);
not NOT1 (N3581, N3548);
not NOT1 (N3582, N3578);
nor NOR4 (N3583, N3582, N1860, N1956, N3391);
not NOT1 (N3584, N3551);
not NOT1 (N3585, N3576);
nand NAND2 (N3586, N3581, N3182);
nor NOR3 (N3587, N3583, N3452, N2265);
or OR2 (N3588, N3575, N2541);
and AND3 (N3589, N3585, N365, N2421);
xor XOR2 (N3590, N3584, N1058);
buf BUF1 (N3591, N3586);
nor NOR2 (N3592, N3555, N1357);
or OR2 (N3593, N3569, N2814);
xor XOR2 (N3594, N3590, N2754);
nor NOR4 (N3595, N3591, N608, N287, N1909);
xor XOR2 (N3596, N3592, N1169);
nand NAND3 (N3597, N3587, N3323, N651);
xor XOR2 (N3598, N3573, N2227);
xor XOR2 (N3599, N3597, N1169);
nand NAND3 (N3600, N3589, N3585, N486);
nor NOR2 (N3601, N3595, N2027);
and AND4 (N3602, N3598, N1923, N1458, N2013);
nand NAND2 (N3603, N3594, N3189);
or OR2 (N3604, N3596, N2343);
nor NOR3 (N3605, N3593, N1314, N360);
and AND2 (N3606, N3600, N2619);
or OR2 (N3607, N3601, N3556);
xor XOR2 (N3608, N3604, N3065);
xor XOR2 (N3609, N3606, N3149);
xor XOR2 (N3610, N3603, N113);
nand NAND2 (N3611, N3610, N2505);
and AND4 (N3612, N3609, N2787, N3177, N885);
or OR4 (N3613, N3588, N582, N1469, N188);
nand NAND4 (N3614, N3565, N1242, N1805, N55);
nand NAND2 (N3615, N3608, N317);
not NOT1 (N3616, N3611);
not NOT1 (N3617, N3612);
nand NAND2 (N3618, N3605, N950);
not NOT1 (N3619, N3618);
nor NOR3 (N3620, N3580, N745, N2476);
or OR2 (N3621, N3617, N3307);
buf BUF1 (N3622, N3614);
or OR2 (N3623, N3599, N2760);
nand NAND4 (N3624, N3607, N590, N623, N271);
not NOT1 (N3625, N3616);
xor XOR2 (N3626, N3621, N2137);
not NOT1 (N3627, N3625);
xor XOR2 (N3628, N3623, N1738);
xor XOR2 (N3629, N3624, N3551);
nand NAND2 (N3630, N3602, N3070);
nor NOR4 (N3631, N3630, N512, N368, N3428);
buf BUF1 (N3632, N3613);
or OR3 (N3633, N3628, N2920, N3318);
nand NAND4 (N3634, N3620, N1772, N1753, N2693);
nand NAND3 (N3635, N3615, N779, N3566);
xor XOR2 (N3636, N3632, N482);
and AND2 (N3637, N3626, N3077);
nand NAND4 (N3638, N3634, N3091, N867, N123);
not NOT1 (N3639, N3629);
nand NAND2 (N3640, N3635, N315);
nor NOR4 (N3641, N3638, N2153, N1161, N1859);
buf BUF1 (N3642, N3640);
and AND4 (N3643, N3637, N1751, N2508, N1787);
nor NOR3 (N3644, N3642, N1830, N1330);
not NOT1 (N3645, N3639);
not NOT1 (N3646, N3631);
or OR2 (N3647, N3622, N187);
nor NOR3 (N3648, N3636, N2935, N3027);
nor NOR2 (N3649, N3645, N2996);
not NOT1 (N3650, N3648);
and AND2 (N3651, N3627, N103);
nand NAND2 (N3652, N3649, N1743);
or OR3 (N3653, N3646, N2672, N860);
and AND2 (N3654, N3641, N3129);
and AND4 (N3655, N3653, N1503, N3430, N1421);
and AND4 (N3656, N3643, N294, N1285, N861);
or OR2 (N3657, N3654, N2590);
xor XOR2 (N3658, N3633, N2983);
buf BUF1 (N3659, N3650);
buf BUF1 (N3660, N3655);
or OR2 (N3661, N3658, N1272);
nor NOR3 (N3662, N3661, N2788, N2196);
or OR4 (N3663, N3662, N2297, N530, N2682);
xor XOR2 (N3664, N3660, N423);
xor XOR2 (N3665, N3619, N1320);
and AND3 (N3666, N3651, N3458, N461);
xor XOR2 (N3667, N3663, N2308);
xor XOR2 (N3668, N3666, N2687);
nand NAND3 (N3669, N3665, N1898, N2358);
xor XOR2 (N3670, N3656, N1848);
not NOT1 (N3671, N3647);
or OR4 (N3672, N3652, N169, N70, N2993);
buf BUF1 (N3673, N3659);
not NOT1 (N3674, N3664);
and AND3 (N3675, N3673, N3147, N1229);
not NOT1 (N3676, N3671);
not NOT1 (N3677, N3668);
and AND4 (N3678, N3670, N1634, N351, N1513);
or OR4 (N3679, N3675, N2865, N3341, N2987);
and AND4 (N3680, N3669, N1932, N2523, N362);
or OR2 (N3681, N3679, N825);
xor XOR2 (N3682, N3677, N3034);
not NOT1 (N3683, N3667);
nor NOR4 (N3684, N3682, N2685, N352, N458);
buf BUF1 (N3685, N3681);
and AND4 (N3686, N3657, N1500, N1406, N1495);
buf BUF1 (N3687, N3644);
not NOT1 (N3688, N3680);
nor NOR3 (N3689, N3688, N520, N2018);
xor XOR2 (N3690, N3676, N263);
buf BUF1 (N3691, N3690);
nand NAND4 (N3692, N3684, N1429, N3015, N2164);
nand NAND2 (N3693, N3674, N460);
nor NOR4 (N3694, N3686, N1372, N1431, N1400);
buf BUF1 (N3695, N3687);
and AND3 (N3696, N3678, N1085, N1320);
xor XOR2 (N3697, N3672, N1083);
nand NAND2 (N3698, N3695, N2476);
or OR2 (N3699, N3691, N1477);
or OR2 (N3700, N3683, N2603);
xor XOR2 (N3701, N3689, N272);
and AND4 (N3702, N3697, N1651, N3701, N437);
nor NOR2 (N3703, N1652, N1447);
xor XOR2 (N3704, N3699, N1995);
nand NAND3 (N3705, N3700, N1116, N690);
nand NAND4 (N3706, N3702, N3258, N2813, N3121);
nor NOR4 (N3707, N3706, N300, N2625, N754);
nor NOR2 (N3708, N3692, N298);
and AND2 (N3709, N3705, N1964);
nand NAND2 (N3710, N3703, N2437);
or OR2 (N3711, N3693, N666);
nand NAND2 (N3712, N3710, N1776);
or OR2 (N3713, N3708, N130);
or OR3 (N3714, N3685, N2363, N990);
nor NOR4 (N3715, N3707, N756, N1260, N2138);
not NOT1 (N3716, N3694);
buf BUF1 (N3717, N3704);
nand NAND2 (N3718, N3717, N3297);
buf BUF1 (N3719, N3711);
xor XOR2 (N3720, N3712, N53);
and AND3 (N3721, N3714, N3079, N3237);
and AND3 (N3722, N3698, N1192, N1254);
xor XOR2 (N3723, N3721, N101);
nand NAND3 (N3724, N3715, N1441, N868);
not NOT1 (N3725, N3713);
nor NOR2 (N3726, N3724, N1161);
nor NOR4 (N3727, N3726, N40, N47, N16);
and AND4 (N3728, N3709, N2676, N2207, N1795);
nor NOR4 (N3729, N3716, N1215, N899, N1235);
not NOT1 (N3730, N3719);
xor XOR2 (N3731, N3696, N255);
buf BUF1 (N3732, N3730);
not NOT1 (N3733, N3720);
not NOT1 (N3734, N3733);
buf BUF1 (N3735, N3722);
xor XOR2 (N3736, N3727, N258);
buf BUF1 (N3737, N3735);
xor XOR2 (N3738, N3732, N1674);
buf BUF1 (N3739, N3736);
buf BUF1 (N3740, N3718);
nand NAND2 (N3741, N3725, N110);
and AND3 (N3742, N3723, N2667, N75);
xor XOR2 (N3743, N3731, N2987);
and AND3 (N3744, N3740, N2992, N785);
or OR4 (N3745, N3742, N489, N696, N3371);
and AND4 (N3746, N3739, N3406, N2224, N385);
buf BUF1 (N3747, N3738);
and AND2 (N3748, N3728, N2821);
buf BUF1 (N3749, N3737);
buf BUF1 (N3750, N3746);
xor XOR2 (N3751, N3743, N1951);
not NOT1 (N3752, N3745);
not NOT1 (N3753, N3744);
or OR3 (N3754, N3752, N3395, N2014);
and AND2 (N3755, N3748, N1140);
nor NOR4 (N3756, N3747, N1328, N2372, N2227);
or OR4 (N3757, N3729, N2644, N1672, N3555);
xor XOR2 (N3758, N3757, N1193);
or OR2 (N3759, N3756, N995);
and AND4 (N3760, N3758, N1509, N2169, N1958);
and AND3 (N3761, N3754, N792, N2185);
xor XOR2 (N3762, N3753, N1672);
nor NOR3 (N3763, N3761, N1423, N2454);
not NOT1 (N3764, N3734);
xor XOR2 (N3765, N3762, N2577);
buf BUF1 (N3766, N3741);
buf BUF1 (N3767, N3759);
and AND2 (N3768, N3767, N2083);
xor XOR2 (N3769, N3766, N2941);
buf BUF1 (N3770, N3751);
nor NOR4 (N3771, N3760, N1531, N70, N1464);
xor XOR2 (N3772, N3764, N3067);
nand NAND4 (N3773, N3763, N2050, N1730, N3244);
or OR4 (N3774, N3773, N910, N746, N1738);
not NOT1 (N3775, N3769);
xor XOR2 (N3776, N3750, N439);
nand NAND2 (N3777, N3771, N1881);
nor NOR2 (N3778, N3772, N25);
or OR3 (N3779, N3749, N1789, N945);
or OR4 (N3780, N3778, N3589, N3137, N3712);
or OR3 (N3781, N3768, N3009, N3429);
buf BUF1 (N3782, N3776);
xor XOR2 (N3783, N3781, N2437);
nand NAND4 (N3784, N3774, N239, N2844, N397);
and AND2 (N3785, N3783, N1589);
and AND3 (N3786, N3780, N299, N2626);
or OR2 (N3787, N3784, N2253);
and AND4 (N3788, N3785, N3201, N3744, N682);
not NOT1 (N3789, N3779);
xor XOR2 (N3790, N3789, N3198);
and AND3 (N3791, N3770, N356, N3515);
nand NAND3 (N3792, N3765, N823, N1774);
xor XOR2 (N3793, N3775, N1594);
xor XOR2 (N3794, N3793, N764);
xor XOR2 (N3795, N3777, N1186);
nor NOR3 (N3796, N3786, N2769, N1755);
nand NAND4 (N3797, N3790, N1886, N2721, N2531);
nor NOR2 (N3798, N3792, N475);
not NOT1 (N3799, N3797);
and AND2 (N3800, N3796, N2974);
and AND3 (N3801, N3800, N119, N1929);
or OR3 (N3802, N3798, N2111, N1352);
xor XOR2 (N3803, N3795, N319);
xor XOR2 (N3804, N3803, N3070);
or OR4 (N3805, N3782, N2167, N3768, N2450);
and AND2 (N3806, N3804, N2314);
and AND4 (N3807, N3755, N2714, N1337, N3749);
nand NAND3 (N3808, N3807, N2943, N2369);
nand NAND2 (N3809, N3788, N1867);
xor XOR2 (N3810, N3794, N126);
not NOT1 (N3811, N3809);
nor NOR4 (N3812, N3802, N2539, N555, N2772);
xor XOR2 (N3813, N3811, N3210);
nor NOR2 (N3814, N3813, N1257);
and AND2 (N3815, N3806, N2305);
or OR4 (N3816, N3791, N305, N3776, N70);
nor NOR2 (N3817, N3815, N776);
not NOT1 (N3818, N3799);
nand NAND3 (N3819, N3816, N3419, N1768);
nand NAND2 (N3820, N3814, N2410);
not NOT1 (N3821, N3820);
xor XOR2 (N3822, N3817, N3078);
and AND4 (N3823, N3801, N66, N2011, N1185);
nor NOR3 (N3824, N3808, N1056, N1568);
nor NOR3 (N3825, N3810, N1975, N2729);
nor NOR3 (N3826, N3805, N216, N2441);
nor NOR4 (N3827, N3826, N3503, N1829, N809);
xor XOR2 (N3828, N3827, N1034);
buf BUF1 (N3829, N3819);
not NOT1 (N3830, N3823);
and AND3 (N3831, N3825, N1169, N2065);
nor NOR4 (N3832, N3812, N2276, N1053, N1644);
nand NAND2 (N3833, N3831, N741);
and AND3 (N3834, N3821, N1285, N265);
buf BUF1 (N3835, N3824);
buf BUF1 (N3836, N3834);
nand NAND3 (N3837, N3829, N2753, N2456);
and AND2 (N3838, N3822, N1293);
nand NAND3 (N3839, N3828, N2384, N2356);
and AND3 (N3840, N3787, N3459, N3567);
not NOT1 (N3841, N3818);
nor NOR2 (N3842, N3830, N3829);
buf BUF1 (N3843, N3835);
nor NOR4 (N3844, N3842, N2052, N1551, N1384);
nor NOR2 (N3845, N3839, N1956);
buf BUF1 (N3846, N3841);
xor XOR2 (N3847, N3838, N3110);
buf BUF1 (N3848, N3836);
or OR3 (N3849, N3843, N1669, N2748);
xor XOR2 (N3850, N3848, N2083);
nand NAND4 (N3851, N3845, N1482, N498, N114);
nand NAND3 (N3852, N3847, N1427, N2829);
nor NOR4 (N3853, N3849, N2172, N2565, N958);
not NOT1 (N3854, N3844);
xor XOR2 (N3855, N3837, N2952);
and AND4 (N3856, N3833, N1299, N881, N3429);
or OR3 (N3857, N3853, N2785, N2579);
and AND4 (N3858, N3852, N2050, N2653, N3782);
not NOT1 (N3859, N3850);
nand NAND4 (N3860, N3856, N2498, N1370, N3256);
xor XOR2 (N3861, N3859, N3847);
buf BUF1 (N3862, N3851);
and AND4 (N3863, N3840, N1458, N1849, N3800);
nand NAND3 (N3864, N3854, N700, N983);
not NOT1 (N3865, N3832);
xor XOR2 (N3866, N3846, N2187);
nand NAND3 (N3867, N3857, N1751, N920);
xor XOR2 (N3868, N3860, N857);
or OR2 (N3869, N3855, N2837);
not NOT1 (N3870, N3867);
buf BUF1 (N3871, N3862);
nand NAND2 (N3872, N3863, N2186);
or OR3 (N3873, N3861, N2108, N1865);
and AND3 (N3874, N3868, N2645, N2488);
buf BUF1 (N3875, N3864);
and AND4 (N3876, N3870, N560, N3728, N1613);
buf BUF1 (N3877, N3872);
xor XOR2 (N3878, N3874, N3823);
not NOT1 (N3879, N3875);
nor NOR2 (N3880, N3877, N3237);
xor XOR2 (N3881, N3876, N1503);
nor NOR3 (N3882, N3858, N1363, N1148);
not NOT1 (N3883, N3881);
nor NOR2 (N3884, N3871, N2913);
buf BUF1 (N3885, N3866);
nand NAND4 (N3886, N3878, N1683, N2002, N546);
and AND2 (N3887, N3883, N1905);
buf BUF1 (N3888, N3886);
buf BUF1 (N3889, N3873);
not NOT1 (N3890, N3885);
buf BUF1 (N3891, N3890);
xor XOR2 (N3892, N3879, N553);
nor NOR2 (N3893, N3891, N2608);
not NOT1 (N3894, N3893);
buf BUF1 (N3895, N3869);
and AND2 (N3896, N3887, N1124);
or OR3 (N3897, N3880, N1763, N973);
or OR4 (N3898, N3895, N2378, N2349, N2945);
nand NAND2 (N3899, N3889, N1944);
nand NAND4 (N3900, N3897, N2663, N683, N2071);
xor XOR2 (N3901, N3899, N48);
or OR2 (N3902, N3882, N2714);
buf BUF1 (N3903, N3902);
xor XOR2 (N3904, N3900, N2316);
xor XOR2 (N3905, N3898, N191);
nor NOR2 (N3906, N3894, N2165);
not NOT1 (N3907, N3892);
nor NOR3 (N3908, N3884, N2078, N579);
and AND2 (N3909, N3908, N2021);
and AND3 (N3910, N3903, N178, N3632);
and AND3 (N3911, N3906, N41, N46);
and AND3 (N3912, N3901, N1417, N3711);
nand NAND3 (N3913, N3865, N1486, N2111);
or OR3 (N3914, N3912, N402, N2665);
buf BUF1 (N3915, N3909);
not NOT1 (N3916, N3911);
xor XOR2 (N3917, N3904, N2979);
or OR3 (N3918, N3913, N2704, N3332);
not NOT1 (N3919, N3917);
and AND3 (N3920, N3916, N1258, N3054);
nand NAND2 (N3921, N3914, N507);
nor NOR3 (N3922, N3888, N3573, N3724);
or OR4 (N3923, N3910, N2499, N3860, N1464);
and AND4 (N3924, N3918, N1653, N3223, N1253);
not NOT1 (N3925, N3919);
and AND4 (N3926, N3924, N3000, N1830, N2452);
nand NAND3 (N3927, N3921, N3280, N2827);
not NOT1 (N3928, N3927);
nand NAND2 (N3929, N3922, N1374);
or OR2 (N3930, N3925, N2231);
buf BUF1 (N3931, N3926);
nand NAND3 (N3932, N3923, N960, N2186);
nor NOR3 (N3933, N3905, N881, N1788);
buf BUF1 (N3934, N3928);
nor NOR3 (N3935, N3929, N712, N2073);
nor NOR4 (N3936, N3935, N3285, N3375, N2994);
and AND3 (N3937, N3933, N2788, N3609);
not NOT1 (N3938, N3907);
or OR2 (N3939, N3932, N432);
and AND3 (N3940, N3920, N680, N1452);
nor NOR4 (N3941, N3930, N3906, N2758, N3930);
buf BUF1 (N3942, N3938);
nand NAND4 (N3943, N3934, N1961, N1810, N1380);
or OR2 (N3944, N3939, N3672);
buf BUF1 (N3945, N3915);
nor NOR3 (N3946, N3943, N3831, N2988);
nand NAND2 (N3947, N3941, N223);
nand NAND2 (N3948, N3931, N3497);
nand NAND3 (N3949, N3940, N1712, N455);
nand NAND3 (N3950, N3948, N2183, N2416);
xor XOR2 (N3951, N3942, N618);
and AND4 (N3952, N3944, N3681, N3049, N1267);
nand NAND2 (N3953, N3945, N1766);
not NOT1 (N3954, N3947);
not NOT1 (N3955, N3896);
and AND2 (N3956, N3955, N662);
or OR2 (N3957, N3953, N3382);
and AND2 (N3958, N3936, N3663);
buf BUF1 (N3959, N3952);
nor NOR4 (N3960, N3946, N1815, N2359, N1160);
xor XOR2 (N3961, N3957, N849);
nor NOR4 (N3962, N3959, N3745, N1584, N3466);
and AND3 (N3963, N3949, N1788, N765);
nand NAND4 (N3964, N3951, N754, N2171, N2864);
and AND4 (N3965, N3954, N3110, N1409, N2522);
buf BUF1 (N3966, N3958);
nor NOR4 (N3967, N3956, N2419, N3180, N1567);
xor XOR2 (N3968, N3960, N172);
not NOT1 (N3969, N3937);
buf BUF1 (N3970, N3967);
xor XOR2 (N3971, N3968, N119);
xor XOR2 (N3972, N3964, N1863);
buf BUF1 (N3973, N3963);
nand NAND3 (N3974, N3961, N301, N1459);
nand NAND4 (N3975, N3974, N2210, N3004, N1126);
or OR4 (N3976, N3966, N140, N1304, N825);
xor XOR2 (N3977, N3972, N1375);
or OR3 (N3978, N3969, N1134, N2266);
or OR3 (N3979, N3950, N2904, N3223);
buf BUF1 (N3980, N3971);
nor NOR3 (N3981, N3979, N892, N3184);
buf BUF1 (N3982, N3978);
buf BUF1 (N3983, N3980);
and AND4 (N3984, N3982, N2674, N3620, N3290);
and AND2 (N3985, N3970, N1011);
xor XOR2 (N3986, N3975, N380);
buf BUF1 (N3987, N3985);
not NOT1 (N3988, N3973);
xor XOR2 (N3989, N3983, N1834);
nor NOR2 (N3990, N3962, N971);
or OR2 (N3991, N3986, N527);
and AND4 (N3992, N3989, N815, N2054, N2326);
buf BUF1 (N3993, N3984);
nand NAND3 (N3994, N3977, N818, N3698);
nand NAND2 (N3995, N3987, N2499);
nor NOR3 (N3996, N3988, N2488, N1086);
nand NAND2 (N3997, N3965, N1388);
and AND4 (N3998, N3997, N2470, N2674, N2471);
nor NOR2 (N3999, N3998, N1072);
nand NAND2 (N4000, N3981, N405);
nor NOR4 (N4001, N3992, N3968, N3014, N1985);
not NOT1 (N4002, N3996);
or OR4 (N4003, N4000, N1457, N3277, N3976);
nand NAND2 (N4004, N3451, N2412);
nand NAND3 (N4005, N4002, N817, N1926);
not NOT1 (N4006, N4005);
xor XOR2 (N4007, N3999, N2170);
and AND2 (N4008, N4004, N2370);
and AND4 (N4009, N4007, N3, N3714, N2839);
nand NAND4 (N4010, N3991, N3836, N2106, N4002);
xor XOR2 (N4011, N3990, N346);
not NOT1 (N4012, N4001);
and AND4 (N4013, N3994, N1144, N1674, N2567);
nand NAND2 (N4014, N3995, N738);
endmodule