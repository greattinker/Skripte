// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14;

output N711,N712,N713,N683,N706,N703,N709,N702,N707,N714;

nand NAND2 (N15, N13, N2);
nor NOR4 (N16, N2, N2, N8, N6);
xor XOR2 (N17, N14, N3);
or OR3 (N18, N3, N11, N6);
nor NOR4 (N19, N5, N13, N8, N6);
and AND3 (N20, N13, N14, N12);
or OR2 (N21, N17, N8);
nor NOR2 (N22, N9, N16);
and AND2 (N23, N13, N5);
buf BUF1 (N24, N13);
or OR4 (N25, N4, N11, N2, N24);
and AND4 (N26, N17, N18, N5, N17);
xor XOR2 (N27, N5, N3);
buf BUF1 (N28, N19);
buf BUF1 (N29, N7);
or OR3 (N30, N22, N5, N7);
buf BUF1 (N31, N20);
buf BUF1 (N32, N28);
or OR3 (N33, N25, N17, N8);
or OR3 (N34, N15, N4, N15);
and AND2 (N35, N34, N13);
buf BUF1 (N36, N33);
xor XOR2 (N37, N30, N27);
nor NOR3 (N38, N9, N24, N21);
and AND2 (N39, N30, N21);
not NOT1 (N40, N31);
not NOT1 (N41, N35);
nor NOR4 (N42, N40, N31, N6, N20);
buf BUF1 (N43, N26);
or OR3 (N44, N36, N39, N18);
not NOT1 (N45, N19);
and AND3 (N46, N29, N43, N32);
buf BUF1 (N47, N2);
and AND4 (N48, N7, N42, N31, N18);
nor NOR4 (N49, N2, N46, N17, N13);
buf BUF1 (N50, N5);
not NOT1 (N51, N41);
not NOT1 (N52, N50);
or OR4 (N53, N51, N35, N42, N31);
and AND4 (N54, N23, N49, N45, N6);
not NOT1 (N55, N33);
nand NAND4 (N56, N15, N26, N14, N37);
xor XOR2 (N57, N15, N16);
not NOT1 (N58, N56);
or OR2 (N59, N38, N58);
nor NOR3 (N60, N7, N23, N20);
or OR2 (N61, N55, N31);
not NOT1 (N62, N61);
nor NOR3 (N63, N48, N26, N29);
nor NOR2 (N64, N63, N2);
xor XOR2 (N65, N64, N21);
and AND4 (N66, N60, N11, N21, N33);
nand NAND4 (N67, N59, N6, N65, N51);
nand NAND4 (N68, N63, N14, N33, N41);
and AND3 (N69, N53, N7, N63);
xor XOR2 (N70, N57, N26);
and AND4 (N71, N54, N16, N27, N21);
and AND4 (N72, N44, N41, N18, N6);
not NOT1 (N73, N71);
and AND4 (N74, N47, N14, N4, N11);
buf BUF1 (N75, N70);
nor NOR4 (N76, N72, N56, N52, N63);
buf BUF1 (N77, N59);
xor XOR2 (N78, N75, N25);
nor NOR4 (N79, N76, N55, N14, N16);
xor XOR2 (N80, N73, N24);
or OR4 (N81, N67, N1, N71, N21);
nor NOR3 (N82, N74, N59, N54);
nor NOR2 (N83, N78, N40);
nor NOR3 (N84, N69, N46, N17);
and AND2 (N85, N79, N63);
not NOT1 (N86, N77);
nor NOR2 (N87, N82, N19);
xor XOR2 (N88, N86, N1);
xor XOR2 (N89, N62, N4);
and AND4 (N90, N84, N80, N78, N50);
and AND2 (N91, N14, N72);
and AND3 (N92, N90, N77, N14);
or OR2 (N93, N87, N8);
or OR3 (N94, N85, N42, N3);
buf BUF1 (N95, N81);
and AND3 (N96, N93, N64, N89);
xor XOR2 (N97, N96, N23);
buf BUF1 (N98, N56);
or OR2 (N99, N92, N80);
nor NOR2 (N100, N91, N14);
nor NOR3 (N101, N68, N25, N91);
or OR2 (N102, N83, N27);
and AND3 (N103, N88, N71, N41);
or OR2 (N104, N101, N21);
xor XOR2 (N105, N95, N26);
xor XOR2 (N106, N103, N24);
xor XOR2 (N107, N66, N22);
not NOT1 (N108, N97);
xor XOR2 (N109, N102, N10);
or OR2 (N110, N94, N93);
xor XOR2 (N111, N98, N59);
not NOT1 (N112, N100);
or OR4 (N113, N108, N100, N85, N100);
not NOT1 (N114, N104);
nand NAND3 (N115, N105, N66, N75);
or OR2 (N116, N107, N81);
buf BUF1 (N117, N106);
or OR2 (N118, N113, N33);
not NOT1 (N119, N110);
buf BUF1 (N120, N116);
nor NOR4 (N121, N112, N15, N117, N83);
and AND2 (N122, N117, N34);
and AND3 (N123, N99, N118, N104);
not NOT1 (N124, N11);
xor XOR2 (N125, N115, N54);
not NOT1 (N126, N111);
and AND4 (N127, N126, N81, N69, N50);
not NOT1 (N128, N119);
and AND4 (N129, N127, N105, N20, N72);
nand NAND4 (N130, N109, N27, N27, N100);
nor NOR4 (N131, N130, N95, N3, N122);
nor NOR3 (N132, N77, N6, N74);
nand NAND3 (N133, N128, N83, N2);
not NOT1 (N134, N132);
or OR2 (N135, N120, N105);
and AND2 (N136, N131, N15);
buf BUF1 (N137, N124);
nor NOR2 (N138, N129, N10);
buf BUF1 (N139, N121);
or OR3 (N140, N139, N10, N96);
xor XOR2 (N141, N114, N114);
xor XOR2 (N142, N134, N125);
nand NAND3 (N143, N45, N51, N77);
and AND2 (N144, N140, N115);
or OR4 (N145, N141, N38, N75, N51);
or OR2 (N146, N145, N39);
or OR3 (N147, N123, N146, N132);
or OR4 (N148, N5, N54, N51, N121);
nand NAND4 (N149, N143, N146, N13, N83);
buf BUF1 (N150, N148);
nor NOR4 (N151, N144, N20, N50, N69);
not NOT1 (N152, N151);
nand NAND2 (N153, N137, N30);
nand NAND2 (N154, N150, N80);
nor NOR3 (N155, N138, N114, N62);
not NOT1 (N156, N135);
not NOT1 (N157, N149);
nand NAND2 (N158, N136, N76);
or OR3 (N159, N153, N51, N18);
buf BUF1 (N160, N159);
xor XOR2 (N161, N154, N96);
not NOT1 (N162, N142);
and AND3 (N163, N155, N73, N113);
or OR2 (N164, N152, N120);
xor XOR2 (N165, N163, N150);
nor NOR3 (N166, N162, N24, N20);
and AND4 (N167, N160, N49, N98, N74);
and AND4 (N168, N166, N33, N57, N94);
nand NAND3 (N169, N167, N142, N163);
buf BUF1 (N170, N157);
not NOT1 (N171, N168);
buf BUF1 (N172, N147);
nor NOR4 (N173, N161, N37, N132, N83);
or OR4 (N174, N169, N156, N103, N4);
or OR4 (N175, N41, N87, N122, N172);
buf BUF1 (N176, N112);
not NOT1 (N177, N173);
not NOT1 (N178, N133);
or OR2 (N179, N171, N5);
xor XOR2 (N180, N170, N91);
and AND4 (N181, N165, N24, N125, N45);
xor XOR2 (N182, N179, N59);
not NOT1 (N183, N181);
buf BUF1 (N184, N175);
or OR2 (N185, N183, N113);
and AND4 (N186, N185, N116, N144, N42);
or OR4 (N187, N180, N168, N14, N165);
nand NAND4 (N188, N174, N102, N102, N26);
xor XOR2 (N189, N176, N98);
xor XOR2 (N190, N178, N74);
not NOT1 (N191, N189);
xor XOR2 (N192, N184, N65);
xor XOR2 (N193, N177, N21);
or OR3 (N194, N164, N107, N146);
and AND3 (N195, N193, N114, N77);
nor NOR4 (N196, N187, N73, N20, N71);
nand NAND2 (N197, N192, N10);
and AND4 (N198, N190, N165, N166, N108);
or OR2 (N199, N194, N193);
buf BUF1 (N200, N197);
not NOT1 (N201, N186);
nand NAND4 (N202, N200, N43, N74, N76);
and AND4 (N203, N191, N178, N114, N117);
or OR2 (N204, N158, N200);
or OR4 (N205, N201, N153, N107, N152);
xor XOR2 (N206, N196, N86);
nand NAND2 (N207, N182, N70);
buf BUF1 (N208, N202);
not NOT1 (N209, N206);
buf BUF1 (N210, N203);
and AND2 (N211, N208, N170);
or OR3 (N212, N207, N208, N151);
nor NOR4 (N213, N195, N111, N154, N207);
nor NOR2 (N214, N212, N83);
nor NOR4 (N215, N214, N41, N90, N152);
nand NAND3 (N216, N199, N82, N152);
not NOT1 (N217, N188);
and AND4 (N218, N216, N146, N155, N134);
buf BUF1 (N219, N209);
nor NOR2 (N220, N219, N144);
and AND2 (N221, N220, N61);
and AND4 (N222, N204, N152, N131, N1);
nand NAND2 (N223, N221, N201);
nand NAND4 (N224, N213, N125, N192, N131);
nor NOR4 (N225, N218, N48, N131, N14);
and AND4 (N226, N225, N70, N97, N35);
not NOT1 (N227, N198);
not NOT1 (N228, N210);
buf BUF1 (N229, N224);
and AND2 (N230, N229, N174);
xor XOR2 (N231, N227, N224);
buf BUF1 (N232, N228);
or OR2 (N233, N232, N207);
nor NOR2 (N234, N211, N118);
xor XOR2 (N235, N233, N212);
not NOT1 (N236, N231);
nor NOR3 (N237, N235, N109, N56);
buf BUF1 (N238, N222);
nand NAND2 (N239, N223, N237);
nor NOR3 (N240, N128, N199, N55);
buf BUF1 (N241, N226);
or OR3 (N242, N230, N90, N202);
or OR2 (N243, N242, N212);
nand NAND4 (N244, N238, N92, N224, N208);
xor XOR2 (N245, N217, N107);
not NOT1 (N246, N241);
and AND2 (N247, N240, N146);
nand NAND3 (N248, N234, N221, N80);
buf BUF1 (N249, N239);
not NOT1 (N250, N236);
xor XOR2 (N251, N244, N236);
xor XOR2 (N252, N215, N223);
xor XOR2 (N253, N252, N39);
or OR2 (N254, N205, N35);
xor XOR2 (N255, N254, N66);
xor XOR2 (N256, N247, N113);
nand NAND4 (N257, N243, N73, N239, N134);
or OR4 (N258, N245, N99, N206, N90);
nor NOR4 (N259, N246, N6, N86, N172);
and AND2 (N260, N259, N166);
nor NOR3 (N261, N256, N104, N199);
not NOT1 (N262, N249);
nand NAND3 (N263, N255, N34, N30);
nor NOR4 (N264, N248, N205, N103, N31);
nand NAND2 (N265, N261, N115);
or OR2 (N266, N262, N25);
not NOT1 (N267, N264);
nand NAND4 (N268, N260, N116, N63, N58);
or OR4 (N269, N263, N218, N27, N21);
nand NAND4 (N270, N258, N60, N179, N3);
nor NOR3 (N271, N269, N133, N64);
buf BUF1 (N272, N271);
buf BUF1 (N273, N267);
buf BUF1 (N274, N257);
buf BUF1 (N275, N272);
or OR4 (N276, N250, N181, N102, N181);
and AND3 (N277, N265, N123, N193);
or OR4 (N278, N268, N195, N54, N131);
buf BUF1 (N279, N274);
buf BUF1 (N280, N277);
nand NAND2 (N281, N280, N213);
and AND2 (N282, N279, N62);
nor NOR2 (N283, N273, N179);
not NOT1 (N284, N281);
nor NOR3 (N285, N266, N227, N146);
or OR3 (N286, N251, N226, N180);
and AND2 (N287, N286, N217);
or OR3 (N288, N285, N253, N108);
or OR4 (N289, N2, N36, N202, N48);
and AND4 (N290, N270, N165, N116, N44);
and AND2 (N291, N276, N25);
and AND3 (N292, N282, N120, N110);
nand NAND2 (N293, N292, N117);
nor NOR2 (N294, N289, N174);
not NOT1 (N295, N284);
and AND4 (N296, N295, N295, N187, N150);
or OR3 (N297, N288, N96, N75);
xor XOR2 (N298, N290, N85);
or OR3 (N299, N275, N267, N184);
xor XOR2 (N300, N296, N29);
nand NAND4 (N301, N291, N218, N64, N287);
buf BUF1 (N302, N99);
and AND3 (N303, N299, N230, N8);
and AND4 (N304, N294, N71, N25, N244);
nand NAND4 (N305, N301, N160, N90, N54);
nor NOR2 (N306, N305, N130);
not NOT1 (N307, N300);
nor NOR4 (N308, N298, N259, N22, N195);
nand NAND2 (N309, N283, N17);
not NOT1 (N310, N308);
nor NOR3 (N311, N297, N20, N9);
and AND4 (N312, N278, N134, N38, N252);
buf BUF1 (N313, N309);
not NOT1 (N314, N302);
not NOT1 (N315, N311);
nand NAND3 (N316, N304, N49, N179);
buf BUF1 (N317, N313);
buf BUF1 (N318, N303);
nor NOR3 (N319, N318, N166, N213);
or OR2 (N320, N319, N161);
nor NOR2 (N321, N316, N215);
buf BUF1 (N322, N314);
or OR2 (N323, N306, N269);
buf BUF1 (N324, N310);
nor NOR3 (N325, N321, N260, N62);
buf BUF1 (N326, N317);
not NOT1 (N327, N324);
nand NAND4 (N328, N322, N121, N80, N35);
nand NAND2 (N329, N323, N96);
not NOT1 (N330, N329);
nor NOR2 (N331, N327, N44);
nand NAND2 (N332, N326, N252);
buf BUF1 (N333, N315);
not NOT1 (N334, N307);
nor NOR2 (N335, N328, N311);
buf BUF1 (N336, N331);
nand NAND4 (N337, N333, N119, N243, N81);
buf BUF1 (N338, N312);
not NOT1 (N339, N330);
and AND2 (N340, N332, N109);
nand NAND4 (N341, N336, N40, N123, N8);
nand NAND3 (N342, N335, N85, N121);
or OR3 (N343, N342, N268, N34);
buf BUF1 (N344, N320);
buf BUF1 (N345, N343);
xor XOR2 (N346, N293, N210);
xor XOR2 (N347, N346, N306);
xor XOR2 (N348, N340, N139);
nand NAND4 (N349, N339, N124, N67, N289);
not NOT1 (N350, N325);
buf BUF1 (N351, N341);
xor XOR2 (N352, N334, N66);
not NOT1 (N353, N344);
nand NAND4 (N354, N338, N241, N288, N274);
xor XOR2 (N355, N350, N154);
nor NOR4 (N356, N351, N176, N217, N336);
xor XOR2 (N357, N345, N340);
not NOT1 (N358, N352);
not NOT1 (N359, N356);
and AND4 (N360, N354, N176, N339, N232);
and AND2 (N361, N349, N306);
buf BUF1 (N362, N357);
xor XOR2 (N363, N358, N5);
or OR3 (N364, N355, N204, N230);
buf BUF1 (N365, N360);
buf BUF1 (N366, N363);
nand NAND3 (N367, N362, N202, N82);
xor XOR2 (N368, N367, N329);
not NOT1 (N369, N366);
nand NAND3 (N370, N368, N22, N162);
not NOT1 (N371, N353);
not NOT1 (N372, N371);
nor NOR2 (N373, N337, N103);
xor XOR2 (N374, N372, N74);
buf BUF1 (N375, N361);
or OR4 (N376, N359, N58, N162, N309);
not NOT1 (N377, N374);
or OR2 (N378, N369, N304);
nand NAND4 (N379, N378, N236, N264, N315);
nor NOR3 (N380, N377, N54, N258);
nor NOR4 (N381, N365, N218, N263, N306);
xor XOR2 (N382, N379, N17);
and AND3 (N383, N376, N105, N108);
buf BUF1 (N384, N364);
buf BUF1 (N385, N375);
nand NAND3 (N386, N373, N233, N246);
nand NAND3 (N387, N382, N157, N363);
not NOT1 (N388, N347);
nand NAND3 (N389, N385, N359, N184);
buf BUF1 (N390, N389);
xor XOR2 (N391, N384, N316);
not NOT1 (N392, N348);
nor NOR2 (N393, N390, N327);
nand NAND2 (N394, N387, N151);
nor NOR2 (N395, N391, N368);
nand NAND4 (N396, N393, N230, N105, N281);
not NOT1 (N397, N395);
not NOT1 (N398, N380);
or OR4 (N399, N386, N323, N27, N341);
buf BUF1 (N400, N396);
buf BUF1 (N401, N397);
and AND2 (N402, N388, N187);
nand NAND2 (N403, N370, N52);
buf BUF1 (N404, N398);
nand NAND4 (N405, N394, N162, N76, N74);
not NOT1 (N406, N405);
nand NAND4 (N407, N401, N178, N290, N13);
nand NAND3 (N408, N392, N103, N278);
nor NOR2 (N409, N402, N26);
and AND2 (N410, N408, N406);
and AND2 (N411, N17, N176);
buf BUF1 (N412, N399);
buf BUF1 (N413, N410);
and AND2 (N414, N400, N348);
nand NAND4 (N415, N381, N226, N407, N18);
and AND3 (N416, N317, N390, N358);
or OR2 (N417, N414, N345);
xor XOR2 (N418, N403, N62);
not NOT1 (N419, N417);
xor XOR2 (N420, N416, N116);
or OR3 (N421, N383, N151, N289);
and AND4 (N422, N411, N121, N381, N180);
not NOT1 (N423, N421);
buf BUF1 (N424, N409);
and AND4 (N425, N422, N414, N247, N208);
nor NOR4 (N426, N419, N102, N297, N111);
not NOT1 (N427, N423);
not NOT1 (N428, N418);
nor NOR2 (N429, N413, N253);
not NOT1 (N430, N425);
nor NOR4 (N431, N404, N323, N315, N346);
nand NAND4 (N432, N430, N69, N251, N169);
and AND4 (N433, N429, N63, N355, N189);
or OR2 (N434, N420, N106);
or OR2 (N435, N434, N318);
nand NAND4 (N436, N426, N4, N373, N109);
nor NOR3 (N437, N432, N340, N269);
nor NOR4 (N438, N424, N3, N195, N282);
not NOT1 (N439, N415);
and AND4 (N440, N436, N354, N38, N157);
nand NAND3 (N441, N428, N280, N176);
nor NOR3 (N442, N441, N317, N308);
or OR3 (N443, N433, N333, N26);
xor XOR2 (N444, N443, N153);
not NOT1 (N445, N439);
nand NAND4 (N446, N442, N96, N260, N351);
or OR2 (N447, N412, N422);
not NOT1 (N448, N435);
nand NAND3 (N449, N445, N95, N30);
buf BUF1 (N450, N437);
and AND4 (N451, N446, N421, N273, N307);
nor NOR4 (N452, N449, N214, N385, N39);
xor XOR2 (N453, N452, N284);
or OR3 (N454, N450, N20, N218);
xor XOR2 (N455, N431, N208);
not NOT1 (N456, N447);
or OR2 (N457, N427, N64);
not NOT1 (N458, N440);
or OR4 (N459, N438, N285, N139, N170);
or OR4 (N460, N458, N74, N7, N440);
buf BUF1 (N461, N448);
nand NAND3 (N462, N451, N136, N453);
not NOT1 (N463, N352);
and AND4 (N464, N459, N17, N396, N434);
or OR3 (N465, N457, N54, N260);
nand NAND3 (N466, N460, N15, N97);
buf BUF1 (N467, N455);
not NOT1 (N468, N461);
and AND4 (N469, N468, N3, N229, N100);
or OR3 (N470, N454, N212, N323);
xor XOR2 (N471, N444, N141);
and AND3 (N472, N467, N333, N30);
or OR3 (N473, N465, N418, N413);
nand NAND4 (N474, N471, N345, N258, N80);
nand NAND2 (N475, N473, N254);
or OR4 (N476, N475, N103, N399, N34);
and AND2 (N477, N462, N208);
xor XOR2 (N478, N472, N137);
nor NOR4 (N479, N469, N301, N227, N89);
nor NOR2 (N480, N477, N43);
nor NOR4 (N481, N480, N83, N152, N295);
nand NAND3 (N482, N479, N174, N234);
or OR4 (N483, N456, N363, N99, N428);
buf BUF1 (N484, N476);
nand NAND4 (N485, N481, N80, N63, N410);
and AND2 (N486, N463, N293);
xor XOR2 (N487, N474, N78);
nor NOR3 (N488, N487, N204, N439);
nand NAND4 (N489, N484, N140, N269, N45);
nor NOR2 (N490, N483, N23);
xor XOR2 (N491, N470, N426);
nand NAND4 (N492, N466, N277, N146, N491);
or OR4 (N493, N397, N363, N461, N278);
and AND4 (N494, N493, N159, N437, N104);
xor XOR2 (N495, N489, N307);
or OR4 (N496, N485, N183, N74, N59);
nand NAND4 (N497, N494, N356, N281, N460);
buf BUF1 (N498, N482);
nand NAND4 (N499, N492, N494, N292, N29);
not NOT1 (N500, N490);
nand NAND2 (N501, N488, N120);
or OR2 (N502, N500, N393);
or OR2 (N503, N502, N58);
or OR3 (N504, N498, N277, N360);
nor NOR2 (N505, N495, N428);
nand NAND3 (N506, N496, N439, N154);
nor NOR4 (N507, N464, N283, N16, N271);
nor NOR4 (N508, N504, N448, N213, N370);
or OR4 (N509, N503, N405, N83, N16);
not NOT1 (N510, N497);
nor NOR2 (N511, N486, N222);
and AND3 (N512, N478, N308, N282);
not NOT1 (N513, N511);
nor NOR3 (N514, N501, N89, N173);
nor NOR3 (N515, N510, N224, N271);
nor NOR4 (N516, N509, N10, N476, N238);
and AND3 (N517, N506, N199, N75);
nor NOR4 (N518, N505, N58, N189, N59);
nand NAND2 (N519, N512, N458);
and AND4 (N520, N513, N492, N11, N71);
or OR3 (N521, N507, N484, N164);
buf BUF1 (N522, N515);
buf BUF1 (N523, N522);
and AND4 (N524, N514, N334, N168, N454);
nor NOR4 (N525, N508, N85, N179, N116);
or OR2 (N526, N523, N384);
nor NOR3 (N527, N526, N400, N355);
buf BUF1 (N528, N519);
not NOT1 (N529, N499);
and AND4 (N530, N527, N147, N202, N295);
nor NOR3 (N531, N524, N142, N310);
not NOT1 (N532, N516);
or OR4 (N533, N532, N465, N291, N331);
nand NAND2 (N534, N525, N501);
and AND4 (N535, N530, N330, N529, N372);
or OR3 (N536, N351, N257, N39);
and AND2 (N537, N534, N536);
and AND2 (N538, N325, N20);
nor NOR3 (N539, N538, N165, N149);
not NOT1 (N540, N518);
nor NOR2 (N541, N520, N136);
and AND2 (N542, N540, N451);
nor NOR2 (N543, N531, N338);
and AND4 (N544, N528, N413, N59, N399);
or OR3 (N545, N535, N68, N522);
xor XOR2 (N546, N544, N113);
nand NAND2 (N547, N545, N422);
or OR3 (N548, N546, N7, N13);
xor XOR2 (N549, N537, N453);
xor XOR2 (N550, N548, N72);
nand NAND2 (N551, N549, N161);
and AND3 (N552, N539, N380, N175);
xor XOR2 (N553, N521, N100);
xor XOR2 (N554, N542, N198);
nor NOR3 (N555, N547, N495, N228);
xor XOR2 (N556, N552, N49);
buf BUF1 (N557, N517);
and AND3 (N558, N555, N442, N133);
or OR4 (N559, N554, N349, N385, N515);
buf BUF1 (N560, N541);
xor XOR2 (N561, N559, N210);
nand NAND3 (N562, N533, N346, N10);
buf BUF1 (N563, N543);
or OR2 (N564, N558, N415);
nand NAND4 (N565, N560, N442, N54, N235);
nand NAND2 (N566, N563, N396);
and AND3 (N567, N557, N78, N525);
nor NOR4 (N568, N550, N297, N36, N567);
nor NOR3 (N569, N322, N431, N153);
or OR3 (N570, N562, N516, N336);
not NOT1 (N571, N566);
buf BUF1 (N572, N570);
not NOT1 (N573, N568);
not NOT1 (N574, N551);
and AND4 (N575, N569, N490, N153, N81);
xor XOR2 (N576, N574, N104);
xor XOR2 (N577, N575, N574);
buf BUF1 (N578, N571);
and AND4 (N579, N564, N346, N119, N313);
xor XOR2 (N580, N565, N378);
xor XOR2 (N581, N572, N417);
nand NAND2 (N582, N578, N222);
buf BUF1 (N583, N576);
xor XOR2 (N584, N579, N339);
not NOT1 (N585, N582);
buf BUF1 (N586, N585);
buf BUF1 (N587, N586);
or OR4 (N588, N581, N488, N322, N281);
nand NAND2 (N589, N556, N398);
nand NAND2 (N590, N583, N390);
and AND3 (N591, N584, N569, N450);
or OR3 (N592, N588, N52, N261);
or OR2 (N593, N553, N150);
nand NAND4 (N594, N573, N193, N376, N18);
not NOT1 (N595, N577);
nand NAND2 (N596, N595, N468);
not NOT1 (N597, N593);
buf BUF1 (N598, N597);
not NOT1 (N599, N589);
nand NAND3 (N600, N590, N517, N249);
and AND2 (N601, N599, N37);
xor XOR2 (N602, N587, N315);
xor XOR2 (N603, N591, N455);
nand NAND2 (N604, N601, N260);
or OR3 (N605, N600, N497, N100);
not NOT1 (N606, N561);
not NOT1 (N607, N603);
not NOT1 (N608, N580);
xor XOR2 (N609, N592, N435);
and AND2 (N610, N602, N300);
not NOT1 (N611, N610);
nor NOR4 (N612, N608, N164, N418, N597);
buf BUF1 (N613, N598);
not NOT1 (N614, N607);
xor XOR2 (N615, N613, N614);
or OR3 (N616, N15, N612, N547);
nand NAND2 (N617, N410, N442);
and AND2 (N618, N616, N223);
nor NOR2 (N619, N617, N572);
buf BUF1 (N620, N605);
nand NAND2 (N621, N604, N555);
or OR4 (N622, N619, N149, N148, N390);
and AND2 (N623, N622, N459);
not NOT1 (N624, N594);
not NOT1 (N625, N618);
and AND2 (N626, N623, N207);
xor XOR2 (N627, N624, N535);
not NOT1 (N628, N609);
nor NOR4 (N629, N627, N174, N563, N510);
xor XOR2 (N630, N606, N593);
buf BUF1 (N631, N611);
or OR3 (N632, N631, N233, N47);
or OR3 (N633, N620, N70, N590);
nand NAND2 (N634, N629, N547);
nor NOR4 (N635, N633, N383, N461, N393);
or OR3 (N636, N596, N40, N51);
nand NAND2 (N637, N630, N374);
not NOT1 (N638, N637);
xor XOR2 (N639, N634, N629);
xor XOR2 (N640, N628, N364);
xor XOR2 (N641, N621, N599);
nor NOR4 (N642, N632, N451, N318, N182);
not NOT1 (N643, N615);
and AND4 (N644, N643, N605, N508, N545);
xor XOR2 (N645, N639, N371);
buf BUF1 (N646, N645);
xor XOR2 (N647, N626, N234);
nand NAND4 (N648, N640, N51, N506, N355);
not NOT1 (N649, N648);
nand NAND2 (N650, N636, N56);
and AND2 (N651, N647, N150);
buf BUF1 (N652, N644);
nand NAND4 (N653, N625, N359, N68, N182);
or OR3 (N654, N650, N34, N514);
not NOT1 (N655, N649);
xor XOR2 (N656, N654, N421);
xor XOR2 (N657, N652, N488);
not NOT1 (N658, N656);
xor XOR2 (N659, N646, N436);
nor NOR3 (N660, N653, N214, N486);
or OR2 (N661, N655, N637);
xor XOR2 (N662, N638, N263);
buf BUF1 (N663, N651);
buf BUF1 (N664, N660);
nand NAND4 (N665, N658, N293, N661, N7);
xor XOR2 (N666, N344, N385);
and AND4 (N667, N657, N307, N224, N213);
nor NOR3 (N668, N662, N60, N655);
xor XOR2 (N669, N641, N283);
xor XOR2 (N670, N666, N325);
not NOT1 (N671, N635);
or OR3 (N672, N667, N114, N23);
buf BUF1 (N673, N642);
nor NOR3 (N674, N663, N269, N125);
nand NAND2 (N675, N665, N188);
xor XOR2 (N676, N675, N489);
and AND4 (N677, N668, N466, N432, N572);
nand NAND3 (N678, N672, N212, N151);
not NOT1 (N679, N674);
nand NAND2 (N680, N678, N149);
xor XOR2 (N681, N669, N581);
buf BUF1 (N682, N676);
or OR2 (N683, N682, N89);
buf BUF1 (N684, N664);
and AND3 (N685, N670, N513, N108);
buf BUF1 (N686, N671);
xor XOR2 (N687, N679, N519);
not NOT1 (N688, N681);
or OR4 (N689, N659, N251, N365, N195);
and AND3 (N690, N677, N60, N256);
or OR2 (N691, N684, N117);
nand NAND3 (N692, N688, N24, N474);
nand NAND4 (N693, N685, N321, N687, N547);
buf BUF1 (N694, N320);
buf BUF1 (N695, N680);
not NOT1 (N696, N690);
nand NAND2 (N697, N686, N142);
nor NOR2 (N698, N673, N679);
and AND4 (N699, N691, N284, N46, N512);
xor XOR2 (N700, N689, N648);
or OR4 (N701, N695, N479, N207, N359);
xor XOR2 (N702, N698, N189);
nor NOR3 (N703, N701, N302, N592);
or OR3 (N704, N692, N264, N591);
xor XOR2 (N705, N697, N378);
buf BUF1 (N706, N704);
or OR3 (N707, N696, N572, N65);
buf BUF1 (N708, N693);
nand NAND3 (N709, N694, N373, N198);
xor XOR2 (N710, N699, N296);
buf BUF1 (N711, N700);
and AND4 (N712, N710, N637, N139, N321);
xor XOR2 (N713, N705, N244);
nor NOR3 (N714, N708, N246, N353);
endmodule