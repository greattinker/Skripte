// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22;

output N4017,N4007,N4003,N4021,N4019,N4020,N4014,N4011,N4015,N4022;

nor NOR3 (N23, N1, N9, N20);
nand NAND2 (N24, N10, N9);
buf BUF1 (N25, N12);
xor XOR2 (N26, N2, N24);
or OR2 (N27, N23, N5);
buf BUF1 (N28, N21);
not NOT1 (N29, N5);
xor XOR2 (N30, N29, N25);
or OR2 (N31, N27, N25);
nor NOR2 (N32, N21, N18);
nor NOR2 (N33, N2, N6);
xor XOR2 (N34, N27, N19);
nor NOR3 (N35, N28, N10, N14);
xor XOR2 (N36, N6, N32);
or OR3 (N37, N21, N17, N21);
nand NAND2 (N38, N35, N14);
xor XOR2 (N39, N11, N37);
xor XOR2 (N40, N35, N23);
not NOT1 (N41, N24);
and AND3 (N42, N34, N38, N24);
nor NOR4 (N43, N37, N28, N34, N7);
nor NOR3 (N44, N36, N21, N31);
and AND4 (N45, N6, N28, N33, N44);
nor NOR4 (N46, N32, N32, N15, N2);
nand NAND3 (N47, N8, N9, N14);
xor XOR2 (N48, N26, N33);
xor XOR2 (N49, N47, N8);
nand NAND2 (N50, N46, N5);
nor NOR3 (N51, N50, N48, N46);
or OR3 (N52, N13, N45, N17);
not NOT1 (N53, N22);
buf BUF1 (N54, N41);
and AND4 (N55, N30, N54, N2, N26);
buf BUF1 (N56, N26);
xor XOR2 (N57, N55, N34);
nand NAND4 (N58, N57, N42, N16, N22);
nand NAND3 (N59, N52, N10, N49);
or OR4 (N60, N26, N58, N23, N8);
nand NAND3 (N61, N13, N5, N25);
xor XOR2 (N62, N42, N59);
nand NAND3 (N63, N38, N37, N40);
not NOT1 (N64, N42);
xor XOR2 (N65, N56, N50);
xor XOR2 (N66, N65, N55);
buf BUF1 (N67, N66);
nand NAND4 (N68, N60, N35, N5, N52);
xor XOR2 (N69, N63, N42);
buf BUF1 (N70, N51);
buf BUF1 (N71, N68);
not NOT1 (N72, N69);
and AND4 (N73, N43, N69, N27, N35);
buf BUF1 (N74, N39);
or OR2 (N75, N71, N35);
or OR2 (N76, N61, N23);
not NOT1 (N77, N74);
or OR4 (N78, N77, N37, N6, N66);
or OR3 (N79, N72, N37, N10);
or OR3 (N80, N75, N41, N46);
and AND4 (N81, N76, N45, N32, N1);
nor NOR2 (N82, N67, N40);
not NOT1 (N83, N80);
xor XOR2 (N84, N64, N46);
or OR2 (N85, N79, N45);
nand NAND4 (N86, N70, N67, N74, N41);
not NOT1 (N87, N73);
xor XOR2 (N88, N82, N11);
buf BUF1 (N89, N53);
and AND3 (N90, N84, N27, N25);
buf BUF1 (N91, N88);
xor XOR2 (N92, N62, N82);
xor XOR2 (N93, N78, N52);
xor XOR2 (N94, N81, N63);
or OR2 (N95, N86, N20);
xor XOR2 (N96, N87, N12);
nor NOR4 (N97, N96, N40, N3, N96);
not NOT1 (N98, N95);
and AND4 (N99, N92, N5, N59, N60);
not NOT1 (N100, N91);
nand NAND3 (N101, N93, N2, N41);
nor NOR3 (N102, N100, N30, N72);
nand NAND3 (N103, N102, N60, N96);
nor NOR4 (N104, N90, N16, N36, N83);
xor XOR2 (N105, N29, N46);
nor NOR2 (N106, N103, N52);
nor NOR2 (N107, N105, N104);
or OR2 (N108, N26, N94);
not NOT1 (N109, N80);
or OR4 (N110, N108, N34, N46, N51);
xor XOR2 (N111, N110, N90);
xor XOR2 (N112, N107, N18);
or OR3 (N113, N85, N9, N91);
nand NAND4 (N114, N99, N27, N79, N29);
and AND4 (N115, N106, N37, N57, N109);
buf BUF1 (N116, N105);
or OR4 (N117, N116, N91, N38, N97);
nand NAND3 (N118, N88, N34, N80);
or OR4 (N119, N112, N83, N44, N117);
or OR2 (N120, N38, N24);
not NOT1 (N121, N113);
or OR2 (N122, N89, N57);
not NOT1 (N123, N122);
xor XOR2 (N124, N101, N72);
buf BUF1 (N125, N121);
xor XOR2 (N126, N125, N9);
nor NOR3 (N127, N126, N110, N59);
not NOT1 (N128, N120);
nand NAND4 (N129, N118, N105, N64, N83);
or OR2 (N130, N124, N100);
and AND4 (N131, N123, N127, N114, N78);
nor NOR4 (N132, N109, N90, N98, N35);
or OR3 (N133, N95, N25, N41);
and AND3 (N134, N30, N109, N17);
and AND3 (N135, N128, N125, N19);
buf BUF1 (N136, N115);
not NOT1 (N137, N119);
not NOT1 (N138, N130);
not NOT1 (N139, N138);
or OR4 (N140, N136, N12, N61, N36);
and AND4 (N141, N129, N7, N93, N116);
nor NOR3 (N142, N139, N66, N128);
or OR4 (N143, N141, N134, N63, N54);
or OR4 (N144, N99, N89, N132, N115);
buf BUF1 (N145, N2);
nand NAND3 (N146, N135, N90, N18);
and AND3 (N147, N142, N110, N131);
nor NOR2 (N148, N123, N135);
and AND2 (N149, N137, N117);
nand NAND2 (N150, N146, N116);
nand NAND4 (N151, N148, N138, N71, N55);
not NOT1 (N152, N149);
nor NOR2 (N153, N145, N55);
not NOT1 (N154, N143);
xor XOR2 (N155, N111, N27);
or OR4 (N156, N150, N147, N64, N58);
or OR4 (N157, N75, N147, N6, N35);
xor XOR2 (N158, N154, N69);
buf BUF1 (N159, N155);
and AND4 (N160, N133, N34, N65, N52);
or OR2 (N161, N158, N21);
nand NAND3 (N162, N161, N69, N127);
not NOT1 (N163, N152);
or OR2 (N164, N144, N59);
nand NAND2 (N165, N162, N59);
nor NOR3 (N166, N160, N110, N15);
or OR3 (N167, N163, N94, N152);
not NOT1 (N168, N151);
and AND4 (N169, N153, N6, N70, N31);
and AND2 (N170, N140, N155);
and AND4 (N171, N159, N72, N52, N29);
nand NAND3 (N172, N165, N2, N127);
xor XOR2 (N173, N156, N58);
nor NOR3 (N174, N168, N92, N33);
or OR3 (N175, N170, N84, N5);
nand NAND2 (N176, N175, N170);
and AND3 (N177, N172, N79, N27);
nor NOR2 (N178, N174, N24);
or OR2 (N179, N166, N127);
or OR3 (N180, N171, N92, N18);
nor NOR4 (N181, N173, N81, N155, N106);
not NOT1 (N182, N167);
nor NOR4 (N183, N164, N163, N82, N132);
or OR4 (N184, N178, N125, N155, N111);
nor NOR2 (N185, N176, N76);
not NOT1 (N186, N180);
and AND3 (N187, N179, N174, N105);
and AND4 (N188, N183, N18, N53, N79);
xor XOR2 (N189, N186, N73);
xor XOR2 (N190, N189, N84);
xor XOR2 (N191, N181, N82);
not NOT1 (N192, N182);
and AND2 (N193, N187, N85);
or OR2 (N194, N157, N32);
and AND4 (N195, N193, N170, N139, N174);
not NOT1 (N196, N188);
nand NAND3 (N197, N196, N109, N32);
not NOT1 (N198, N185);
or OR4 (N199, N177, N103, N185, N126);
nand NAND3 (N200, N169, N162, N186);
buf BUF1 (N201, N199);
nor NOR3 (N202, N184, N98, N171);
or OR4 (N203, N191, N148, N127, N199);
and AND3 (N204, N190, N174, N118);
or OR3 (N205, N204, N195, N60);
or OR2 (N206, N7, N51);
or OR2 (N207, N205, N55);
or OR4 (N208, N197, N160, N150, N114);
nand NAND4 (N209, N207, N158, N181, N2);
not NOT1 (N210, N202);
and AND2 (N211, N203, N26);
and AND4 (N212, N206, N201, N187, N129);
buf BUF1 (N213, N136);
nor NOR3 (N214, N210, N167, N11);
and AND4 (N215, N198, N167, N112, N148);
buf BUF1 (N216, N209);
and AND4 (N217, N200, N191, N165, N21);
and AND3 (N218, N215, N201, N171);
buf BUF1 (N219, N208);
nand NAND3 (N220, N217, N147, N109);
xor XOR2 (N221, N194, N213);
not NOT1 (N222, N8);
and AND3 (N223, N214, N210, N147);
nand NAND4 (N224, N221, N26, N112, N52);
buf BUF1 (N225, N222);
xor XOR2 (N226, N192, N47);
or OR3 (N227, N219, N213, N175);
buf BUF1 (N228, N216);
nor NOR3 (N229, N223, N45, N131);
and AND2 (N230, N228, N151);
not NOT1 (N231, N229);
xor XOR2 (N232, N211, N78);
or OR4 (N233, N220, N157, N154, N186);
nor NOR3 (N234, N226, N7, N200);
not NOT1 (N235, N230);
xor XOR2 (N236, N232, N84);
buf BUF1 (N237, N225);
or OR2 (N238, N237, N67);
buf BUF1 (N239, N233);
xor XOR2 (N240, N238, N40);
buf BUF1 (N241, N236);
nand NAND2 (N242, N241, N145);
not NOT1 (N243, N242);
or OR2 (N244, N239, N67);
xor XOR2 (N245, N224, N102);
nor NOR3 (N246, N231, N146, N76);
xor XOR2 (N247, N244, N163);
buf BUF1 (N248, N245);
nor NOR4 (N249, N212, N134, N8, N133);
nand NAND4 (N250, N247, N143, N133, N45);
and AND2 (N251, N218, N234);
nand NAND2 (N252, N109, N52);
nand NAND2 (N253, N246, N66);
not NOT1 (N254, N251);
nand NAND3 (N255, N253, N221, N95);
and AND4 (N256, N252, N60, N105, N40);
not NOT1 (N257, N240);
nor NOR2 (N258, N249, N98);
buf BUF1 (N259, N258);
buf BUF1 (N260, N256);
nor NOR2 (N261, N248, N194);
nand NAND2 (N262, N235, N234);
nand NAND3 (N263, N260, N222, N168);
buf BUF1 (N264, N257);
buf BUF1 (N265, N259);
and AND3 (N266, N250, N150, N43);
and AND3 (N267, N262, N23, N160);
not NOT1 (N268, N264);
and AND2 (N269, N255, N64);
nor NOR3 (N270, N254, N107, N89);
xor XOR2 (N271, N268, N97);
buf BUF1 (N272, N263);
not NOT1 (N273, N267);
xor XOR2 (N274, N266, N24);
xor XOR2 (N275, N243, N259);
nor NOR2 (N276, N273, N33);
nor NOR3 (N277, N271, N251, N61);
buf BUF1 (N278, N274);
buf BUF1 (N279, N278);
nand NAND3 (N280, N261, N137, N140);
buf BUF1 (N281, N279);
and AND3 (N282, N280, N47, N176);
nand NAND4 (N283, N270, N202, N32, N196);
nor NOR4 (N284, N275, N128, N269, N84);
and AND4 (N285, N256, N26, N65, N159);
nor NOR4 (N286, N272, N235, N210, N79);
or OR3 (N287, N283, N276, N173);
xor XOR2 (N288, N186, N248);
not NOT1 (N289, N288);
buf BUF1 (N290, N227);
buf BUF1 (N291, N277);
not NOT1 (N292, N287);
xor XOR2 (N293, N289, N280);
or OR2 (N294, N291, N142);
xor XOR2 (N295, N284, N233);
xor XOR2 (N296, N281, N10);
or OR2 (N297, N282, N250);
or OR3 (N298, N293, N93, N9);
buf BUF1 (N299, N298);
buf BUF1 (N300, N285);
or OR3 (N301, N295, N44, N199);
not NOT1 (N302, N301);
not NOT1 (N303, N297);
not NOT1 (N304, N290);
xor XOR2 (N305, N286, N211);
buf BUF1 (N306, N299);
xor XOR2 (N307, N305, N153);
nand NAND2 (N308, N300, N121);
and AND2 (N309, N307, N138);
and AND4 (N310, N296, N221, N106, N176);
nor NOR4 (N311, N294, N112, N190, N284);
and AND4 (N312, N303, N65, N175, N158);
nor NOR4 (N313, N311, N196, N107, N41);
or OR3 (N314, N292, N111, N304);
and AND2 (N315, N201, N73);
nor NOR3 (N316, N306, N77, N11);
nand NAND4 (N317, N313, N277, N271, N156);
nor NOR4 (N318, N312, N8, N191, N311);
xor XOR2 (N319, N308, N169);
and AND3 (N320, N265, N147, N73);
nand NAND4 (N321, N315, N176, N89, N38);
xor XOR2 (N322, N321, N223);
and AND2 (N323, N310, N188);
buf BUF1 (N324, N314);
nor NOR2 (N325, N309, N94);
nand NAND3 (N326, N318, N154, N238);
nand NAND4 (N327, N302, N50, N207, N64);
not NOT1 (N328, N324);
and AND3 (N329, N328, N124, N18);
nor NOR2 (N330, N322, N54);
or OR2 (N331, N323, N183);
and AND4 (N332, N325, N81, N150, N278);
nand NAND2 (N333, N330, N108);
nand NAND2 (N334, N317, N53);
xor XOR2 (N335, N334, N70);
xor XOR2 (N336, N326, N79);
not NOT1 (N337, N320);
nand NAND3 (N338, N329, N128, N178);
nand NAND2 (N339, N338, N77);
not NOT1 (N340, N332);
and AND4 (N341, N333, N223, N10, N42);
and AND2 (N342, N337, N51);
not NOT1 (N343, N319);
nor NOR3 (N344, N339, N171, N181);
or OR4 (N345, N343, N334, N294, N335);
buf BUF1 (N346, N220);
xor XOR2 (N347, N346, N287);
or OR4 (N348, N327, N82, N195, N170);
or OR3 (N349, N336, N62, N222);
buf BUF1 (N350, N316);
buf BUF1 (N351, N347);
and AND4 (N352, N341, N195, N172, N7);
not NOT1 (N353, N350);
buf BUF1 (N354, N348);
or OR3 (N355, N340, N258, N308);
nor NOR2 (N356, N331, N286);
not NOT1 (N357, N355);
xor XOR2 (N358, N353, N88);
nor NOR3 (N359, N345, N330, N55);
not NOT1 (N360, N356);
nor NOR2 (N361, N352, N213);
or OR4 (N362, N360, N268, N26, N55);
or OR2 (N363, N354, N94);
buf BUF1 (N364, N358);
nand NAND2 (N365, N344, N90);
buf BUF1 (N366, N349);
nand NAND3 (N367, N359, N183, N349);
nand NAND3 (N368, N364, N125, N9);
xor XOR2 (N369, N368, N260);
or OR2 (N370, N342, N168);
xor XOR2 (N371, N357, N361);
buf BUF1 (N372, N56);
xor XOR2 (N373, N370, N22);
nor NOR3 (N374, N373, N151, N186);
or OR4 (N375, N372, N73, N351, N228);
or OR2 (N376, N184, N154);
not NOT1 (N377, N375);
not NOT1 (N378, N371);
not NOT1 (N379, N376);
nand NAND2 (N380, N367, N247);
nor NOR4 (N381, N377, N77, N342, N108);
buf BUF1 (N382, N374);
nor NOR2 (N383, N362, N198);
nand NAND3 (N384, N383, N67, N212);
buf BUF1 (N385, N382);
and AND3 (N386, N380, N378, N180);
xor XOR2 (N387, N293, N79);
xor XOR2 (N388, N381, N358);
not NOT1 (N389, N385);
and AND2 (N390, N387, N136);
and AND3 (N391, N389, N218, N389);
not NOT1 (N392, N365);
and AND4 (N393, N366, N92, N315, N49);
buf BUF1 (N394, N369);
not NOT1 (N395, N390);
or OR2 (N396, N379, N3);
nor NOR4 (N397, N388, N73, N379, N166);
buf BUF1 (N398, N394);
or OR3 (N399, N396, N381, N376);
and AND3 (N400, N399, N350, N39);
and AND2 (N401, N397, N29);
xor XOR2 (N402, N391, N315);
nor NOR4 (N403, N363, N323, N388, N194);
or OR2 (N404, N384, N112);
not NOT1 (N405, N403);
buf BUF1 (N406, N392);
buf BUF1 (N407, N401);
and AND3 (N408, N400, N28, N35);
nor NOR4 (N409, N393, N378, N386, N85);
xor XOR2 (N410, N37, N110);
nor NOR3 (N411, N407, N403, N17);
or OR3 (N412, N405, N403, N364);
nor NOR3 (N413, N409, N48, N257);
and AND4 (N414, N408, N240, N191, N223);
not NOT1 (N415, N404);
buf BUF1 (N416, N398);
nor NOR3 (N417, N412, N333, N137);
buf BUF1 (N418, N416);
and AND2 (N419, N411, N272);
and AND2 (N420, N410, N61);
not NOT1 (N421, N418);
and AND2 (N422, N417, N226);
or OR3 (N423, N395, N222, N213);
xor XOR2 (N424, N421, N137);
xor XOR2 (N425, N413, N338);
not NOT1 (N426, N423);
buf BUF1 (N427, N415);
or OR4 (N428, N419, N283, N252, N244);
and AND2 (N429, N426, N6);
nand NAND2 (N430, N420, N397);
not NOT1 (N431, N430);
or OR2 (N432, N425, N15);
nor NOR2 (N433, N414, N46);
xor XOR2 (N434, N402, N343);
not NOT1 (N435, N406);
xor XOR2 (N436, N424, N372);
and AND3 (N437, N431, N118, N151);
or OR3 (N438, N435, N433, N238);
xor XOR2 (N439, N419, N272);
or OR4 (N440, N432, N33, N272, N73);
not NOT1 (N441, N429);
nand NAND4 (N442, N440, N164, N108, N404);
nand NAND4 (N443, N442, N211, N67, N431);
or OR4 (N444, N428, N351, N209, N172);
not NOT1 (N445, N443);
xor XOR2 (N446, N437, N69);
buf BUF1 (N447, N446);
xor XOR2 (N448, N434, N87);
not NOT1 (N449, N444);
not NOT1 (N450, N438);
not NOT1 (N451, N441);
or OR2 (N452, N445, N130);
or OR3 (N453, N427, N139, N322);
xor XOR2 (N454, N451, N31);
not NOT1 (N455, N447);
nand NAND4 (N456, N450, N157, N198, N242);
not NOT1 (N457, N456);
xor XOR2 (N458, N455, N445);
nor NOR4 (N459, N452, N234, N424, N436);
nor NOR4 (N460, N104, N399, N404, N137);
xor XOR2 (N461, N457, N145);
or OR2 (N462, N439, N176);
buf BUF1 (N463, N449);
xor XOR2 (N464, N461, N14);
not NOT1 (N465, N459);
buf BUF1 (N466, N454);
nor NOR4 (N467, N463, N395, N337, N252);
xor XOR2 (N468, N464, N454);
nand NAND2 (N469, N460, N112);
xor XOR2 (N470, N469, N4);
nor NOR3 (N471, N453, N223, N83);
buf BUF1 (N472, N462);
buf BUF1 (N473, N467);
or OR2 (N474, N466, N272);
nor NOR4 (N475, N471, N59, N370, N165);
nor NOR3 (N476, N422, N373, N122);
nor NOR4 (N477, N476, N281, N313, N81);
buf BUF1 (N478, N474);
or OR3 (N479, N458, N197, N378);
not NOT1 (N480, N479);
nand NAND2 (N481, N478, N267);
nand NAND2 (N482, N448, N458);
xor XOR2 (N483, N470, N19);
or OR3 (N484, N483, N213, N168);
and AND4 (N485, N477, N454, N484, N275);
nor NOR2 (N486, N293, N396);
nor NOR3 (N487, N472, N298, N172);
xor XOR2 (N488, N468, N221);
xor XOR2 (N489, N485, N329);
or OR4 (N490, N481, N375, N246, N1);
nand NAND4 (N491, N486, N286, N1, N445);
nor NOR3 (N492, N475, N150, N63);
or OR2 (N493, N482, N98);
nor NOR4 (N494, N493, N352, N46, N386);
xor XOR2 (N495, N487, N403);
nand NAND3 (N496, N488, N44, N326);
xor XOR2 (N497, N491, N420);
not NOT1 (N498, N480);
nand NAND4 (N499, N490, N444, N394, N476);
or OR2 (N500, N494, N314);
and AND3 (N501, N497, N213, N324);
buf BUF1 (N502, N501);
nor NOR4 (N503, N502, N57, N377, N268);
nand NAND2 (N504, N499, N81);
nor NOR4 (N505, N504, N378, N392, N420);
buf BUF1 (N506, N473);
or OR4 (N507, N503, N480, N504, N451);
or OR3 (N508, N507, N219, N73);
xor XOR2 (N509, N465, N187);
nor NOR3 (N510, N492, N88, N141);
xor XOR2 (N511, N500, N82);
buf BUF1 (N512, N506);
buf BUF1 (N513, N489);
nor NOR3 (N514, N509, N348, N100);
not NOT1 (N515, N511);
buf BUF1 (N516, N498);
not NOT1 (N517, N516);
not NOT1 (N518, N495);
and AND4 (N519, N518, N81, N230, N392);
and AND2 (N520, N510, N334);
buf BUF1 (N521, N513);
xor XOR2 (N522, N517, N255);
buf BUF1 (N523, N519);
buf BUF1 (N524, N496);
nand NAND3 (N525, N521, N176, N371);
xor XOR2 (N526, N522, N359);
or OR3 (N527, N520, N307, N47);
nand NAND4 (N528, N512, N82, N93, N444);
not NOT1 (N529, N526);
xor XOR2 (N530, N524, N162);
not NOT1 (N531, N505);
nor NOR3 (N532, N525, N406, N451);
or OR4 (N533, N515, N125, N313, N331);
not NOT1 (N534, N533);
xor XOR2 (N535, N531, N409);
nor NOR3 (N536, N523, N417, N123);
or OR3 (N537, N532, N514, N386);
nand NAND2 (N538, N200, N261);
nor NOR4 (N539, N537, N182, N213, N306);
not NOT1 (N540, N535);
or OR4 (N541, N538, N209, N316, N155);
nand NAND4 (N542, N534, N515, N304, N365);
not NOT1 (N543, N527);
nor NOR4 (N544, N529, N176, N539, N245);
xor XOR2 (N545, N228, N253);
or OR4 (N546, N508, N206, N424, N402);
or OR2 (N547, N545, N193);
and AND4 (N548, N536, N237, N144, N505);
nand NAND2 (N549, N546, N213);
nand NAND3 (N550, N530, N29, N265);
xor XOR2 (N551, N540, N93);
or OR4 (N552, N548, N302, N308, N301);
and AND4 (N553, N550, N364, N244, N365);
or OR4 (N554, N544, N382, N442, N122);
xor XOR2 (N555, N549, N225);
and AND2 (N556, N528, N132);
xor XOR2 (N557, N547, N544);
nand NAND4 (N558, N555, N224, N83, N24);
nor NOR3 (N559, N543, N191, N59);
nor NOR4 (N560, N552, N553, N153, N87);
nand NAND4 (N561, N316, N218, N471, N197);
not NOT1 (N562, N541);
not NOT1 (N563, N551);
or OR2 (N564, N560, N411);
buf BUF1 (N565, N564);
xor XOR2 (N566, N559, N98);
not NOT1 (N567, N565);
buf BUF1 (N568, N542);
not NOT1 (N569, N568);
and AND4 (N570, N563, N85, N83, N171);
nand NAND4 (N571, N569, N294, N246, N62);
xor XOR2 (N572, N567, N195);
nand NAND4 (N573, N571, N352, N127, N411);
and AND3 (N574, N566, N187, N243);
buf BUF1 (N575, N574);
and AND2 (N576, N557, N390);
nand NAND4 (N577, N561, N157, N299, N169);
buf BUF1 (N578, N573);
not NOT1 (N579, N576);
nor NOR3 (N580, N575, N483, N439);
and AND4 (N581, N556, N101, N249, N97);
nand NAND3 (N582, N558, N284, N433);
nand NAND4 (N583, N562, N521, N388, N444);
xor XOR2 (N584, N577, N330);
not NOT1 (N585, N582);
buf BUF1 (N586, N554);
and AND2 (N587, N580, N232);
nor NOR3 (N588, N587, N519, N578);
not NOT1 (N589, N139);
not NOT1 (N590, N585);
not NOT1 (N591, N581);
xor XOR2 (N592, N588, N425);
and AND3 (N593, N592, N312, N395);
or OR4 (N594, N584, N262, N168, N234);
not NOT1 (N595, N589);
not NOT1 (N596, N595);
not NOT1 (N597, N579);
or OR4 (N598, N594, N123, N575, N337);
buf BUF1 (N599, N598);
nand NAND2 (N600, N596, N95);
nand NAND4 (N601, N583, N566, N569, N368);
nor NOR4 (N602, N601, N443, N52, N520);
nor NOR4 (N603, N586, N514, N388, N163);
nor NOR4 (N604, N572, N317, N506, N183);
not NOT1 (N605, N603);
xor XOR2 (N606, N590, N177);
or OR2 (N607, N602, N31);
buf BUF1 (N608, N570);
xor XOR2 (N609, N591, N77);
nor NOR3 (N610, N609, N549, N593);
xor XOR2 (N611, N466, N577);
and AND4 (N612, N605, N574, N276, N479);
buf BUF1 (N613, N612);
and AND4 (N614, N604, N394, N492, N542);
buf BUF1 (N615, N610);
xor XOR2 (N616, N614, N424);
nand NAND2 (N617, N615, N134);
not NOT1 (N618, N599);
nand NAND4 (N619, N617, N84, N328, N39);
or OR2 (N620, N618, N138);
and AND4 (N621, N600, N470, N118, N369);
or OR2 (N622, N616, N242);
nor NOR4 (N623, N606, N408, N406, N225);
and AND4 (N624, N613, N225, N100, N334);
nand NAND2 (N625, N621, N516);
xor XOR2 (N626, N622, N606);
buf BUF1 (N627, N619);
xor XOR2 (N628, N607, N160);
buf BUF1 (N629, N624);
and AND2 (N630, N627, N96);
buf BUF1 (N631, N630);
nand NAND2 (N632, N626, N529);
or OR4 (N633, N625, N387, N316, N7);
buf BUF1 (N634, N597);
not NOT1 (N635, N634);
and AND4 (N636, N623, N186, N230, N222);
and AND3 (N637, N620, N195, N284);
buf BUF1 (N638, N611);
or OR4 (N639, N635, N163, N12, N595);
nand NAND2 (N640, N629, N445);
or OR4 (N641, N633, N110, N172, N585);
xor XOR2 (N642, N641, N496);
xor XOR2 (N643, N632, N136);
buf BUF1 (N644, N643);
and AND2 (N645, N640, N546);
and AND4 (N646, N636, N227, N89, N642);
not NOT1 (N647, N110);
not NOT1 (N648, N646);
nand NAND3 (N649, N638, N109, N169);
and AND4 (N650, N631, N626, N342, N529);
xor XOR2 (N651, N628, N290);
nand NAND3 (N652, N650, N121, N274);
and AND3 (N653, N648, N121, N166);
or OR4 (N654, N651, N519, N289, N132);
nand NAND4 (N655, N649, N300, N548, N575);
nand NAND2 (N656, N608, N541);
xor XOR2 (N657, N654, N229);
nand NAND2 (N658, N647, N413);
nand NAND2 (N659, N657, N33);
nand NAND3 (N660, N653, N68, N194);
or OR2 (N661, N637, N463);
buf BUF1 (N662, N655);
or OR3 (N663, N644, N558, N178);
buf BUF1 (N664, N645);
and AND3 (N665, N662, N295, N324);
nand NAND2 (N666, N639, N416);
nand NAND2 (N667, N656, N142);
not NOT1 (N668, N652);
nand NAND2 (N669, N665, N607);
and AND4 (N670, N668, N216, N561, N361);
nor NOR3 (N671, N660, N552, N669);
not NOT1 (N672, N524);
buf BUF1 (N673, N659);
nor NOR4 (N674, N672, N404, N220, N290);
xor XOR2 (N675, N674, N286);
and AND4 (N676, N670, N160, N305, N665);
nand NAND4 (N677, N673, N370, N202, N477);
buf BUF1 (N678, N671);
xor XOR2 (N679, N675, N39);
buf BUF1 (N680, N677);
nand NAND2 (N681, N679, N464);
and AND2 (N682, N678, N28);
buf BUF1 (N683, N667);
and AND4 (N684, N663, N450, N346, N10);
xor XOR2 (N685, N683, N683);
xor XOR2 (N686, N685, N428);
nor NOR4 (N687, N681, N200, N32, N349);
not NOT1 (N688, N680);
buf BUF1 (N689, N664);
not NOT1 (N690, N684);
xor XOR2 (N691, N689, N131);
nand NAND2 (N692, N691, N123);
or OR3 (N693, N686, N448, N614);
buf BUF1 (N694, N693);
buf BUF1 (N695, N688);
xor XOR2 (N696, N687, N298);
not NOT1 (N697, N694);
xor XOR2 (N698, N690, N304);
or OR3 (N699, N696, N482, N578);
nor NOR4 (N700, N698, N648, N439, N638);
and AND2 (N701, N666, N528);
xor XOR2 (N702, N682, N246);
xor XOR2 (N703, N702, N365);
nand NAND4 (N704, N701, N380, N181, N397);
not NOT1 (N705, N658);
or OR2 (N706, N704, N277);
nand NAND3 (N707, N705, N485, N486);
or OR3 (N708, N699, N517, N379);
nand NAND4 (N709, N708, N300, N161, N637);
not NOT1 (N710, N695);
nand NAND3 (N711, N697, N31, N559);
or OR3 (N712, N676, N699, N673);
not NOT1 (N713, N700);
nand NAND3 (N714, N712, N591, N687);
nand NAND2 (N715, N661, N113);
nor NOR3 (N716, N707, N698, N60);
buf BUF1 (N717, N692);
and AND4 (N718, N716, N54, N652, N519);
not NOT1 (N719, N709);
nor NOR3 (N720, N706, N237, N222);
xor XOR2 (N721, N719, N159);
not NOT1 (N722, N703);
nand NAND4 (N723, N722, N446, N515, N459);
not NOT1 (N724, N713);
nand NAND2 (N725, N720, N323);
buf BUF1 (N726, N710);
not NOT1 (N727, N715);
and AND4 (N728, N718, N533, N572, N399);
nand NAND2 (N729, N727, N651);
or OR2 (N730, N714, N518);
or OR3 (N731, N711, N374, N378);
nor NOR3 (N732, N724, N406, N344);
nand NAND4 (N733, N731, N13, N8, N445);
nor NOR3 (N734, N729, N290, N247);
or OR4 (N735, N733, N660, N619, N114);
or OR4 (N736, N721, N98, N92, N1);
or OR2 (N737, N726, N403);
and AND4 (N738, N717, N273, N677, N565);
nor NOR4 (N739, N728, N57, N712, N185);
nand NAND2 (N740, N732, N155);
not NOT1 (N741, N739);
not NOT1 (N742, N723);
xor XOR2 (N743, N738, N670);
not NOT1 (N744, N737);
nor NOR2 (N745, N730, N83);
or OR3 (N746, N745, N270, N659);
or OR3 (N747, N740, N552, N308);
xor XOR2 (N748, N746, N280);
nand NAND3 (N749, N742, N453, N465);
not NOT1 (N750, N748);
xor XOR2 (N751, N725, N103);
or OR4 (N752, N736, N243, N488, N674);
not NOT1 (N753, N741);
or OR3 (N754, N749, N8, N532);
or OR4 (N755, N750, N715, N566, N723);
xor XOR2 (N756, N751, N121);
nor NOR4 (N757, N744, N666, N656, N731);
or OR3 (N758, N756, N256, N726);
not NOT1 (N759, N758);
nor NOR4 (N760, N754, N539, N215, N569);
nor NOR2 (N761, N760, N745);
not NOT1 (N762, N735);
nand NAND4 (N763, N755, N646, N720, N262);
or OR2 (N764, N753, N331);
buf BUF1 (N765, N761);
not NOT1 (N766, N757);
buf BUF1 (N767, N765);
xor XOR2 (N768, N752, N543);
nor NOR4 (N769, N743, N591, N63, N35);
not NOT1 (N770, N768);
and AND4 (N771, N769, N455, N178, N498);
nor NOR3 (N772, N734, N592, N715);
or OR3 (N773, N770, N273, N456);
nand NAND3 (N774, N764, N59, N71);
or OR3 (N775, N771, N298, N337);
and AND2 (N776, N767, N458);
not NOT1 (N777, N747);
nor NOR4 (N778, N777, N755, N290, N499);
xor XOR2 (N779, N772, N130);
nand NAND4 (N780, N776, N634, N203, N573);
nand NAND3 (N781, N766, N562, N749);
not NOT1 (N782, N780);
not NOT1 (N783, N773);
or OR2 (N784, N762, N538);
not NOT1 (N785, N784);
nand NAND2 (N786, N763, N429);
or OR2 (N787, N781, N363);
xor XOR2 (N788, N783, N49);
buf BUF1 (N789, N786);
not NOT1 (N790, N775);
nand NAND2 (N791, N789, N583);
xor XOR2 (N792, N759, N7);
or OR4 (N793, N785, N551, N313, N68);
and AND4 (N794, N779, N565, N543, N707);
nor NOR3 (N795, N774, N378, N110);
nor NOR2 (N796, N795, N265);
not NOT1 (N797, N778);
buf BUF1 (N798, N793);
buf BUF1 (N799, N794);
nor NOR2 (N800, N797, N794);
buf BUF1 (N801, N796);
not NOT1 (N802, N788);
and AND4 (N803, N791, N769, N260, N28);
buf BUF1 (N804, N802);
or OR3 (N805, N804, N521, N230);
nand NAND3 (N806, N803, N578, N607);
nand NAND3 (N807, N792, N478, N494);
buf BUF1 (N808, N799);
nand NAND4 (N809, N790, N393, N122, N72);
buf BUF1 (N810, N787);
xor XOR2 (N811, N798, N251);
or OR4 (N812, N810, N296, N519, N671);
buf BUF1 (N813, N812);
not NOT1 (N814, N806);
nor NOR3 (N815, N801, N321, N690);
xor XOR2 (N816, N800, N476);
nand NAND4 (N817, N816, N35, N524, N163);
not NOT1 (N818, N813);
xor XOR2 (N819, N805, N462);
nor NOR2 (N820, N782, N362);
and AND4 (N821, N818, N1, N253, N776);
and AND2 (N822, N811, N152);
nor NOR2 (N823, N814, N724);
nand NAND2 (N824, N807, N557);
not NOT1 (N825, N820);
xor XOR2 (N826, N817, N404);
buf BUF1 (N827, N821);
nand NAND2 (N828, N825, N296);
xor XOR2 (N829, N822, N516);
and AND3 (N830, N829, N296, N395);
not NOT1 (N831, N826);
not NOT1 (N832, N827);
nand NAND3 (N833, N831, N146, N48);
xor XOR2 (N834, N823, N347);
nand NAND3 (N835, N828, N448, N467);
buf BUF1 (N836, N819);
buf BUF1 (N837, N834);
not NOT1 (N838, N808);
not NOT1 (N839, N836);
nor NOR4 (N840, N832, N582, N2, N809);
not NOT1 (N841, N603);
or OR2 (N842, N835, N532);
not NOT1 (N843, N839);
nand NAND4 (N844, N840, N328, N438, N563);
nor NOR4 (N845, N815, N170, N422, N175);
nor NOR4 (N846, N841, N626, N584, N203);
buf BUF1 (N847, N843);
and AND2 (N848, N844, N518);
xor XOR2 (N849, N845, N410);
xor XOR2 (N850, N849, N633);
nor NOR2 (N851, N838, N282);
buf BUF1 (N852, N848);
buf BUF1 (N853, N837);
nor NOR2 (N854, N824, N490);
or OR3 (N855, N850, N270, N654);
nor NOR3 (N856, N854, N400, N578);
nor NOR3 (N857, N833, N796, N585);
nor NOR3 (N858, N851, N315, N106);
nand NAND2 (N859, N857, N857);
or OR2 (N860, N847, N47);
buf BUF1 (N861, N856);
and AND4 (N862, N861, N436, N716, N797);
nand NAND3 (N863, N846, N143, N719);
buf BUF1 (N864, N842);
or OR2 (N865, N860, N830);
or OR3 (N866, N125, N263, N650);
not NOT1 (N867, N862);
nor NOR2 (N868, N853, N804);
xor XOR2 (N869, N866, N858);
xor XOR2 (N870, N429, N423);
xor XOR2 (N871, N867, N19);
xor XOR2 (N872, N855, N106);
and AND3 (N873, N870, N678, N624);
not NOT1 (N874, N868);
nand NAND2 (N875, N869, N365);
nand NAND2 (N876, N872, N218);
buf BUF1 (N877, N873);
nand NAND2 (N878, N864, N161);
nand NAND3 (N879, N863, N400, N557);
or OR3 (N880, N878, N444, N394);
nand NAND4 (N881, N880, N782, N2, N668);
or OR4 (N882, N877, N672, N500, N277);
or OR4 (N883, N882, N794, N626, N234);
nor NOR3 (N884, N871, N771, N383);
and AND2 (N885, N884, N497);
and AND2 (N886, N879, N97);
and AND4 (N887, N875, N146, N547, N308);
not NOT1 (N888, N874);
buf BUF1 (N889, N852);
and AND3 (N890, N876, N162, N637);
buf BUF1 (N891, N885);
and AND4 (N892, N883, N476, N309, N279);
xor XOR2 (N893, N889, N644);
nand NAND2 (N894, N888, N474);
not NOT1 (N895, N881);
xor XOR2 (N896, N890, N273);
and AND4 (N897, N887, N287, N444, N461);
not NOT1 (N898, N892);
nand NAND3 (N899, N865, N25, N98);
xor XOR2 (N900, N886, N220);
buf BUF1 (N901, N896);
and AND3 (N902, N900, N768, N748);
nand NAND3 (N903, N894, N523, N197);
nand NAND2 (N904, N895, N457);
buf BUF1 (N905, N859);
not NOT1 (N906, N898);
buf BUF1 (N907, N905);
buf BUF1 (N908, N901);
not NOT1 (N909, N897);
buf BUF1 (N910, N903);
xor XOR2 (N911, N907, N601);
and AND2 (N912, N906, N477);
nor NOR2 (N913, N902, N665);
and AND3 (N914, N913, N404, N26);
or OR4 (N915, N908, N641, N434, N458);
nor NOR4 (N916, N914, N395, N730, N732);
nor NOR4 (N917, N916, N52, N384, N194);
nand NAND2 (N918, N893, N22);
and AND2 (N919, N904, N715);
and AND4 (N920, N919, N379, N205, N597);
or OR4 (N921, N918, N626, N872, N274);
nand NAND2 (N922, N899, N174);
nand NAND3 (N923, N922, N76, N914);
buf BUF1 (N924, N912);
or OR2 (N925, N921, N612);
not NOT1 (N926, N911);
and AND2 (N927, N925, N584);
and AND3 (N928, N927, N187, N147);
buf BUF1 (N929, N926);
and AND2 (N930, N923, N908);
buf BUF1 (N931, N920);
or OR2 (N932, N910, N412);
xor XOR2 (N933, N915, N142);
not NOT1 (N934, N933);
nor NOR3 (N935, N929, N220, N623);
xor XOR2 (N936, N909, N343);
and AND4 (N937, N928, N894, N272, N484);
and AND4 (N938, N917, N404, N394, N729);
not NOT1 (N939, N931);
nand NAND4 (N940, N939, N819, N457, N75);
or OR3 (N941, N930, N62, N397);
xor XOR2 (N942, N938, N612);
or OR3 (N943, N940, N299, N880);
and AND4 (N944, N934, N481, N838, N222);
buf BUF1 (N945, N936);
buf BUF1 (N946, N935);
or OR2 (N947, N937, N579);
xor XOR2 (N948, N947, N399);
and AND4 (N949, N932, N68, N364, N74);
buf BUF1 (N950, N924);
xor XOR2 (N951, N891, N726);
nor NOR2 (N952, N941, N305);
not NOT1 (N953, N944);
and AND4 (N954, N951, N238, N209, N898);
nand NAND4 (N955, N954, N191, N340, N863);
nor NOR4 (N956, N952, N212, N769, N884);
or OR2 (N957, N955, N306);
nor NOR4 (N958, N949, N819, N673, N802);
buf BUF1 (N959, N948);
not NOT1 (N960, N953);
xor XOR2 (N961, N945, N823);
nand NAND2 (N962, N946, N243);
and AND2 (N963, N956, N174);
nor NOR2 (N964, N942, N358);
not NOT1 (N965, N950);
xor XOR2 (N966, N963, N48);
and AND3 (N967, N961, N584, N779);
or OR2 (N968, N965, N73);
or OR4 (N969, N968, N481, N554, N670);
or OR2 (N970, N958, N197);
nand NAND2 (N971, N959, N855);
or OR3 (N972, N962, N688, N581);
or OR2 (N973, N969, N878);
not NOT1 (N974, N943);
not NOT1 (N975, N971);
nor NOR3 (N976, N973, N19, N309);
or OR2 (N977, N966, N962);
nand NAND4 (N978, N970, N540, N243, N947);
nor NOR4 (N979, N978, N675, N709, N126);
not NOT1 (N980, N976);
buf BUF1 (N981, N967);
buf BUF1 (N982, N975);
and AND3 (N983, N974, N164, N932);
and AND2 (N984, N980, N769);
and AND3 (N985, N972, N869, N21);
and AND2 (N986, N984, N439);
or OR3 (N987, N982, N452, N417);
not NOT1 (N988, N985);
not NOT1 (N989, N964);
not NOT1 (N990, N979);
or OR3 (N991, N986, N684, N420);
not NOT1 (N992, N989);
or OR3 (N993, N960, N567, N358);
nand NAND2 (N994, N983, N733);
buf BUF1 (N995, N957);
buf BUF1 (N996, N977);
and AND3 (N997, N991, N313, N794);
or OR3 (N998, N992, N797, N756);
and AND2 (N999, N997, N218);
nor NOR4 (N1000, N993, N235, N646, N956);
nor NOR4 (N1001, N1000, N309, N823, N632);
nand NAND4 (N1002, N988, N68, N859, N382);
buf BUF1 (N1003, N996);
or OR3 (N1004, N994, N207, N698);
or OR3 (N1005, N987, N895, N32);
and AND3 (N1006, N1002, N843, N64);
or OR4 (N1007, N1004, N957, N590, N255);
nor NOR3 (N1008, N999, N333, N115);
nor NOR4 (N1009, N990, N413, N673, N768);
buf BUF1 (N1010, N1006);
and AND3 (N1011, N981, N858, N803);
nand NAND4 (N1012, N1011, N733, N410, N100);
not NOT1 (N1013, N1001);
nand NAND3 (N1014, N1003, N788, N580);
nand NAND2 (N1015, N1014, N856);
nand NAND4 (N1016, N1007, N372, N214, N40);
nand NAND2 (N1017, N1009, N264);
not NOT1 (N1018, N1005);
xor XOR2 (N1019, N995, N304);
and AND4 (N1020, N998, N164, N461, N577);
not NOT1 (N1021, N1019);
or OR2 (N1022, N1010, N84);
nand NAND2 (N1023, N1018, N133);
and AND4 (N1024, N1022, N162, N575, N105);
xor XOR2 (N1025, N1013, N647);
not NOT1 (N1026, N1017);
xor XOR2 (N1027, N1008, N663);
and AND3 (N1028, N1020, N666, N437);
nor NOR3 (N1029, N1025, N607, N632);
not NOT1 (N1030, N1016);
not NOT1 (N1031, N1015);
nor NOR2 (N1032, N1021, N219);
nor NOR3 (N1033, N1032, N879, N810);
and AND4 (N1034, N1024, N829, N963, N334);
and AND3 (N1035, N1027, N905, N398);
xor XOR2 (N1036, N1033, N385);
buf BUF1 (N1037, N1028);
xor XOR2 (N1038, N1037, N896);
nand NAND4 (N1039, N1026, N676, N974, N531);
xor XOR2 (N1040, N1034, N1013);
nand NAND2 (N1041, N1023, N565);
buf BUF1 (N1042, N1030);
or OR2 (N1043, N1040, N237);
not NOT1 (N1044, N1029);
buf BUF1 (N1045, N1043);
nand NAND3 (N1046, N1044, N367, N701);
or OR3 (N1047, N1035, N324, N219);
buf BUF1 (N1048, N1041);
not NOT1 (N1049, N1036);
buf BUF1 (N1050, N1046);
and AND4 (N1051, N1038, N303, N344, N380);
nor NOR3 (N1052, N1045, N809, N684);
and AND3 (N1053, N1052, N584, N772);
nor NOR2 (N1054, N1049, N1039);
or OR3 (N1055, N753, N649, N471);
xor XOR2 (N1056, N1048, N338);
nand NAND2 (N1057, N1042, N561);
and AND2 (N1058, N1050, N424);
or OR2 (N1059, N1058, N922);
xor XOR2 (N1060, N1012, N86);
nor NOR3 (N1061, N1056, N779, N653);
and AND3 (N1062, N1031, N18, N583);
nor NOR2 (N1063, N1053, N212);
buf BUF1 (N1064, N1057);
xor XOR2 (N1065, N1063, N934);
xor XOR2 (N1066, N1064, N313);
nor NOR2 (N1067, N1065, N387);
xor XOR2 (N1068, N1067, N597);
not NOT1 (N1069, N1055);
buf BUF1 (N1070, N1061);
or OR4 (N1071, N1069, N270, N784, N829);
nand NAND3 (N1072, N1066, N771, N967);
nand NAND2 (N1073, N1054, N639);
nand NAND4 (N1074, N1073, N693, N365, N376);
nor NOR4 (N1075, N1074, N211, N117, N147);
or OR3 (N1076, N1070, N747, N667);
not NOT1 (N1077, N1071);
or OR4 (N1078, N1059, N675, N389, N952);
and AND3 (N1079, N1078, N644, N113);
or OR3 (N1080, N1047, N693, N242);
and AND3 (N1081, N1060, N1077, N522);
buf BUF1 (N1082, N144);
buf BUF1 (N1083, N1081);
not NOT1 (N1084, N1079);
not NOT1 (N1085, N1083);
and AND2 (N1086, N1051, N295);
buf BUF1 (N1087, N1068);
buf BUF1 (N1088, N1082);
xor XOR2 (N1089, N1084, N179);
not NOT1 (N1090, N1062);
nor NOR3 (N1091, N1085, N908, N57);
or OR3 (N1092, N1072, N670, N257);
or OR4 (N1093, N1087, N40, N1002, N192);
not NOT1 (N1094, N1092);
or OR3 (N1095, N1091, N724, N549);
buf BUF1 (N1096, N1095);
not NOT1 (N1097, N1080);
buf BUF1 (N1098, N1076);
or OR3 (N1099, N1075, N542, N388);
xor XOR2 (N1100, N1093, N957);
and AND4 (N1101, N1086, N649, N1024, N488);
and AND4 (N1102, N1101, N32, N818, N203);
or OR2 (N1103, N1096, N159);
xor XOR2 (N1104, N1098, N747);
and AND2 (N1105, N1088, N157);
buf BUF1 (N1106, N1104);
nand NAND2 (N1107, N1106, N650);
not NOT1 (N1108, N1097);
or OR2 (N1109, N1100, N141);
xor XOR2 (N1110, N1108, N949);
buf BUF1 (N1111, N1109);
not NOT1 (N1112, N1103);
and AND4 (N1113, N1102, N578, N74, N612);
not NOT1 (N1114, N1110);
not NOT1 (N1115, N1090);
or OR3 (N1116, N1113, N281, N270);
xor XOR2 (N1117, N1112, N144);
xor XOR2 (N1118, N1115, N616);
not NOT1 (N1119, N1089);
buf BUF1 (N1120, N1094);
or OR4 (N1121, N1116, N849, N70, N486);
nand NAND3 (N1122, N1111, N974, N1057);
and AND4 (N1123, N1119, N1114, N541, N321);
and AND2 (N1124, N704, N1094);
and AND2 (N1125, N1124, N539);
buf BUF1 (N1126, N1118);
nor NOR3 (N1127, N1125, N932, N217);
not NOT1 (N1128, N1122);
xor XOR2 (N1129, N1127, N912);
not NOT1 (N1130, N1105);
nand NAND2 (N1131, N1107, N414);
buf BUF1 (N1132, N1123);
and AND3 (N1133, N1126, N651, N1052);
xor XOR2 (N1134, N1132, N958);
xor XOR2 (N1135, N1120, N234);
or OR2 (N1136, N1129, N792);
buf BUF1 (N1137, N1117);
nor NOR3 (N1138, N1135, N529, N882);
or OR4 (N1139, N1133, N688, N280, N618);
nor NOR3 (N1140, N1138, N412, N582);
or OR2 (N1141, N1130, N115);
nand NAND2 (N1142, N1141, N760);
nor NOR2 (N1143, N1134, N10);
nor NOR3 (N1144, N1143, N619, N848);
buf BUF1 (N1145, N1128);
nor NOR4 (N1146, N1142, N279, N226, N460);
and AND4 (N1147, N1131, N527, N1002, N1070);
or OR3 (N1148, N1145, N1116, N486);
nand NAND2 (N1149, N1139, N504);
xor XOR2 (N1150, N1149, N678);
nand NAND4 (N1151, N1136, N1133, N174, N738);
xor XOR2 (N1152, N1137, N1106);
nor NOR4 (N1153, N1121, N241, N422, N803);
not NOT1 (N1154, N1150);
and AND2 (N1155, N1144, N148);
not NOT1 (N1156, N1151);
not NOT1 (N1157, N1148);
xor XOR2 (N1158, N1146, N193);
nor NOR2 (N1159, N1099, N97);
and AND3 (N1160, N1156, N568, N126);
or OR2 (N1161, N1155, N978);
nand NAND4 (N1162, N1157, N211, N1012, N52);
xor XOR2 (N1163, N1160, N83);
nand NAND4 (N1164, N1152, N101, N988, N570);
nand NAND2 (N1165, N1164, N277);
and AND2 (N1166, N1147, N768);
nor NOR2 (N1167, N1140, N94);
nand NAND2 (N1168, N1161, N593);
nor NOR3 (N1169, N1159, N554, N36);
and AND3 (N1170, N1167, N757, N224);
nand NAND2 (N1171, N1154, N99);
buf BUF1 (N1172, N1166);
nor NOR4 (N1173, N1168, N862, N1110, N687);
nand NAND2 (N1174, N1169, N561);
not NOT1 (N1175, N1170);
buf BUF1 (N1176, N1162);
buf BUF1 (N1177, N1174);
nand NAND4 (N1178, N1177, N581, N128, N526);
nor NOR4 (N1179, N1173, N764, N362, N32);
not NOT1 (N1180, N1172);
nand NAND4 (N1181, N1175, N725, N573, N129);
and AND4 (N1182, N1180, N837, N20, N323);
buf BUF1 (N1183, N1171);
or OR2 (N1184, N1176, N1137);
and AND3 (N1185, N1183, N2, N697);
nand NAND3 (N1186, N1185, N298, N115);
not NOT1 (N1187, N1158);
not NOT1 (N1188, N1186);
not NOT1 (N1189, N1178);
nor NOR2 (N1190, N1184, N337);
nand NAND3 (N1191, N1181, N824, N710);
xor XOR2 (N1192, N1179, N266);
or OR4 (N1193, N1182, N1119, N550, N1133);
nor NOR2 (N1194, N1189, N959);
nor NOR4 (N1195, N1194, N1021, N774, N710);
not NOT1 (N1196, N1195);
nand NAND2 (N1197, N1188, N745);
xor XOR2 (N1198, N1192, N792);
xor XOR2 (N1199, N1165, N809);
and AND2 (N1200, N1191, N146);
nor NOR4 (N1201, N1190, N24, N681, N224);
not NOT1 (N1202, N1187);
not NOT1 (N1203, N1197);
xor XOR2 (N1204, N1199, N963);
xor XOR2 (N1205, N1193, N240);
xor XOR2 (N1206, N1200, N1138);
nor NOR3 (N1207, N1204, N1147, N877);
nor NOR3 (N1208, N1201, N326, N190);
or OR3 (N1209, N1196, N401, N110);
nor NOR2 (N1210, N1203, N1001);
nor NOR3 (N1211, N1210, N864, N1123);
or OR3 (N1212, N1207, N770, N1078);
nor NOR2 (N1213, N1211, N588);
buf BUF1 (N1214, N1202);
nor NOR3 (N1215, N1214, N586, N165);
nor NOR3 (N1216, N1208, N631, N486);
or OR3 (N1217, N1206, N288, N924);
and AND3 (N1218, N1217, N781, N269);
buf BUF1 (N1219, N1212);
or OR2 (N1220, N1205, N432);
nand NAND2 (N1221, N1218, N88);
nor NOR2 (N1222, N1219, N1025);
or OR3 (N1223, N1222, N646, N779);
and AND4 (N1224, N1221, N711, N110, N731);
xor XOR2 (N1225, N1216, N990);
buf BUF1 (N1226, N1198);
not NOT1 (N1227, N1215);
not NOT1 (N1228, N1213);
nor NOR3 (N1229, N1224, N955, N439);
nor NOR3 (N1230, N1163, N1216, N777);
nor NOR2 (N1231, N1225, N839);
buf BUF1 (N1232, N1227);
and AND4 (N1233, N1228, N442, N640, N757);
or OR2 (N1234, N1231, N572);
or OR3 (N1235, N1232, N559, N751);
and AND2 (N1236, N1233, N340);
and AND3 (N1237, N1226, N123, N977);
and AND4 (N1238, N1220, N106, N923, N469);
and AND2 (N1239, N1236, N1153);
nor NOR3 (N1240, N641, N431, N709);
nand NAND2 (N1241, N1237, N864);
xor XOR2 (N1242, N1235, N327);
or OR4 (N1243, N1241, N838, N643, N948);
not NOT1 (N1244, N1209);
nor NOR4 (N1245, N1229, N1062, N221, N1000);
buf BUF1 (N1246, N1242);
nand NAND3 (N1247, N1246, N881, N620);
nor NOR2 (N1248, N1223, N368);
or OR4 (N1249, N1238, N999, N798, N162);
buf BUF1 (N1250, N1248);
buf BUF1 (N1251, N1243);
buf BUF1 (N1252, N1245);
or OR4 (N1253, N1249, N1033, N540, N785);
nor NOR4 (N1254, N1250, N1097, N278, N437);
or OR2 (N1255, N1254, N869);
buf BUF1 (N1256, N1244);
buf BUF1 (N1257, N1255);
not NOT1 (N1258, N1239);
buf BUF1 (N1259, N1258);
not NOT1 (N1260, N1253);
xor XOR2 (N1261, N1234, N1189);
not NOT1 (N1262, N1261);
xor XOR2 (N1263, N1260, N945);
or OR2 (N1264, N1252, N118);
nor NOR4 (N1265, N1259, N780, N144, N60);
buf BUF1 (N1266, N1251);
or OR3 (N1267, N1256, N628, N942);
and AND4 (N1268, N1266, N790, N992, N324);
xor XOR2 (N1269, N1240, N607);
or OR4 (N1270, N1268, N1139, N782, N477);
or OR2 (N1271, N1270, N612);
xor XOR2 (N1272, N1269, N1144);
nor NOR2 (N1273, N1265, N708);
nand NAND3 (N1274, N1271, N585, N24);
nor NOR3 (N1275, N1264, N242, N1258);
nand NAND3 (N1276, N1273, N101, N276);
buf BUF1 (N1277, N1262);
and AND2 (N1278, N1275, N892);
buf BUF1 (N1279, N1230);
and AND4 (N1280, N1267, N325, N1017, N44);
nand NAND3 (N1281, N1276, N1112, N635);
or OR2 (N1282, N1278, N268);
nor NOR4 (N1283, N1279, N743, N1217, N763);
not NOT1 (N1284, N1283);
not NOT1 (N1285, N1280);
nor NOR3 (N1286, N1247, N146, N885);
nor NOR4 (N1287, N1277, N683, N20, N1014);
nor NOR4 (N1288, N1257, N203, N1228, N815);
nand NAND4 (N1289, N1285, N725, N878, N1168);
nand NAND3 (N1290, N1284, N271, N1161);
nor NOR2 (N1291, N1263, N692);
not NOT1 (N1292, N1289);
nor NOR4 (N1293, N1274, N1182, N826, N942);
nand NAND2 (N1294, N1287, N1272);
nor NOR4 (N1295, N145, N224, N195, N529);
nand NAND4 (N1296, N1282, N66, N632, N1009);
nor NOR4 (N1297, N1294, N353, N87, N274);
and AND3 (N1298, N1286, N882, N389);
buf BUF1 (N1299, N1298);
buf BUF1 (N1300, N1281);
xor XOR2 (N1301, N1288, N582);
or OR4 (N1302, N1295, N456, N848, N452);
and AND3 (N1303, N1301, N313, N506);
not NOT1 (N1304, N1302);
or OR3 (N1305, N1292, N884, N1084);
buf BUF1 (N1306, N1296);
and AND4 (N1307, N1305, N238, N507, N862);
nor NOR4 (N1308, N1293, N249, N46, N75);
and AND4 (N1309, N1291, N628, N736, N857);
nand NAND4 (N1310, N1303, N864, N756, N962);
and AND2 (N1311, N1310, N13);
not NOT1 (N1312, N1306);
nor NOR2 (N1313, N1312, N274);
xor XOR2 (N1314, N1307, N957);
not NOT1 (N1315, N1308);
not NOT1 (N1316, N1313);
not NOT1 (N1317, N1300);
buf BUF1 (N1318, N1314);
xor XOR2 (N1319, N1311, N21);
not NOT1 (N1320, N1317);
or OR3 (N1321, N1315, N958, N135);
nand NAND4 (N1322, N1318, N763, N468, N224);
nor NOR4 (N1323, N1290, N347, N1053, N67);
not NOT1 (N1324, N1319);
buf BUF1 (N1325, N1320);
buf BUF1 (N1326, N1325);
xor XOR2 (N1327, N1326, N648);
nor NOR2 (N1328, N1309, N589);
nor NOR4 (N1329, N1323, N513, N397, N994);
and AND3 (N1330, N1316, N273, N822);
nand NAND2 (N1331, N1304, N803);
nand NAND2 (N1332, N1321, N312);
xor XOR2 (N1333, N1329, N698);
buf BUF1 (N1334, N1324);
xor XOR2 (N1335, N1332, N1052);
or OR2 (N1336, N1322, N406);
xor XOR2 (N1337, N1331, N720);
and AND3 (N1338, N1299, N1237, N643);
nor NOR4 (N1339, N1327, N1335, N385, N70);
not NOT1 (N1340, N314);
not NOT1 (N1341, N1334);
xor XOR2 (N1342, N1297, N24);
nand NAND4 (N1343, N1336, N1032, N1280, N127);
nand NAND4 (N1344, N1333, N463, N1292, N272);
and AND2 (N1345, N1339, N1043);
not NOT1 (N1346, N1330);
and AND4 (N1347, N1337, N808, N241, N527);
nand NAND2 (N1348, N1342, N262);
nand NAND2 (N1349, N1340, N367);
buf BUF1 (N1350, N1328);
buf BUF1 (N1351, N1350);
or OR4 (N1352, N1348, N1313, N1088, N47);
nor NOR4 (N1353, N1352, N509, N187, N346);
buf BUF1 (N1354, N1344);
xor XOR2 (N1355, N1341, N835);
buf BUF1 (N1356, N1355);
xor XOR2 (N1357, N1353, N1039);
buf BUF1 (N1358, N1354);
nor NOR2 (N1359, N1347, N1096);
not NOT1 (N1360, N1356);
not NOT1 (N1361, N1345);
buf BUF1 (N1362, N1361);
xor XOR2 (N1363, N1357, N1013);
or OR2 (N1364, N1338, N1340);
xor XOR2 (N1365, N1362, N494);
buf BUF1 (N1366, N1360);
or OR2 (N1367, N1364, N339);
not NOT1 (N1368, N1343);
xor XOR2 (N1369, N1346, N996);
not NOT1 (N1370, N1367);
buf BUF1 (N1371, N1359);
nor NOR2 (N1372, N1371, N481);
and AND3 (N1373, N1369, N172, N1107);
nand NAND2 (N1374, N1351, N213);
buf BUF1 (N1375, N1370);
nand NAND3 (N1376, N1375, N1158, N954);
and AND3 (N1377, N1374, N1369, N293);
not NOT1 (N1378, N1376);
xor XOR2 (N1379, N1378, N289);
xor XOR2 (N1380, N1379, N559);
or OR3 (N1381, N1377, N113, N896);
nor NOR3 (N1382, N1363, N926, N56);
xor XOR2 (N1383, N1381, N1009);
nand NAND4 (N1384, N1358, N474, N42, N596);
xor XOR2 (N1385, N1383, N43);
not NOT1 (N1386, N1384);
nand NAND4 (N1387, N1386, N296, N963, N669);
nand NAND2 (N1388, N1368, N68);
nor NOR4 (N1389, N1349, N983, N516, N1352);
and AND3 (N1390, N1382, N1007, N829);
nand NAND3 (N1391, N1389, N263, N1007);
not NOT1 (N1392, N1388);
nand NAND4 (N1393, N1373, N862, N520, N791);
nand NAND2 (N1394, N1366, N1239);
or OR2 (N1395, N1391, N493);
or OR2 (N1396, N1395, N362);
not NOT1 (N1397, N1393);
nand NAND4 (N1398, N1380, N1184, N1143, N1008);
and AND4 (N1399, N1385, N64, N202, N333);
or OR3 (N1400, N1397, N493, N834);
nor NOR2 (N1401, N1400, N892);
and AND2 (N1402, N1365, N364);
buf BUF1 (N1403, N1398);
buf BUF1 (N1404, N1392);
nor NOR4 (N1405, N1372, N1254, N1217, N770);
xor XOR2 (N1406, N1394, N569);
or OR2 (N1407, N1401, N1179);
xor XOR2 (N1408, N1402, N1255);
buf BUF1 (N1409, N1405);
xor XOR2 (N1410, N1387, N1180);
or OR4 (N1411, N1406, N1003, N206, N565);
nand NAND3 (N1412, N1410, N52, N960);
buf BUF1 (N1413, N1404);
and AND3 (N1414, N1412, N1275, N1066);
nor NOR3 (N1415, N1396, N923, N952);
nand NAND3 (N1416, N1415, N1303, N107);
xor XOR2 (N1417, N1390, N1166);
not NOT1 (N1418, N1411);
or OR3 (N1419, N1416, N734, N894);
and AND3 (N1420, N1407, N762, N316);
and AND4 (N1421, N1413, N509, N265, N919);
nor NOR4 (N1422, N1409, N1098, N162, N774);
nand NAND3 (N1423, N1420, N502, N643);
not NOT1 (N1424, N1423);
and AND4 (N1425, N1419, N771, N528, N470);
and AND3 (N1426, N1417, N368, N1304);
or OR4 (N1427, N1425, N161, N406, N1220);
and AND2 (N1428, N1426, N1117);
buf BUF1 (N1429, N1424);
buf BUF1 (N1430, N1408);
nand NAND2 (N1431, N1399, N1087);
not NOT1 (N1432, N1422);
or OR2 (N1433, N1421, N1321);
or OR3 (N1434, N1433, N700, N623);
nand NAND4 (N1435, N1418, N1250, N469, N1356);
or OR3 (N1436, N1427, N1185, N1025);
xor XOR2 (N1437, N1430, N788);
and AND4 (N1438, N1435, N1375, N1208, N1195);
or OR3 (N1439, N1434, N619, N115);
xor XOR2 (N1440, N1439, N1376);
xor XOR2 (N1441, N1436, N279);
nor NOR4 (N1442, N1414, N408, N314, N308);
xor XOR2 (N1443, N1432, N449);
buf BUF1 (N1444, N1431);
and AND4 (N1445, N1438, N484, N932, N608);
nand NAND4 (N1446, N1437, N298, N1152, N487);
or OR2 (N1447, N1443, N813);
xor XOR2 (N1448, N1447, N607);
and AND3 (N1449, N1441, N1352, N122);
nand NAND3 (N1450, N1444, N1083, N571);
nand NAND2 (N1451, N1448, N529);
not NOT1 (N1452, N1446);
or OR2 (N1453, N1449, N1383);
nor NOR4 (N1454, N1442, N928, N1043, N740);
nor NOR2 (N1455, N1429, N295);
or OR3 (N1456, N1454, N836, N134);
buf BUF1 (N1457, N1428);
buf BUF1 (N1458, N1403);
not NOT1 (N1459, N1440);
or OR4 (N1460, N1453, N773, N689, N1071);
or OR2 (N1461, N1450, N919);
nor NOR2 (N1462, N1456, N1354);
xor XOR2 (N1463, N1455, N446);
not NOT1 (N1464, N1461);
not NOT1 (N1465, N1464);
and AND3 (N1466, N1463, N245, N174);
or OR4 (N1467, N1458, N1374, N442, N658);
buf BUF1 (N1468, N1445);
xor XOR2 (N1469, N1465, N1097);
nand NAND4 (N1470, N1462, N762, N1149, N682);
buf BUF1 (N1471, N1467);
not NOT1 (N1472, N1470);
nor NOR3 (N1473, N1469, N1220, N680);
buf BUF1 (N1474, N1473);
not NOT1 (N1475, N1460);
nor NOR4 (N1476, N1471, N404, N1021, N647);
not NOT1 (N1477, N1457);
not NOT1 (N1478, N1474);
buf BUF1 (N1479, N1472);
and AND3 (N1480, N1451, N672, N967);
and AND2 (N1481, N1478, N1158);
or OR4 (N1482, N1459, N1270, N341, N1042);
nor NOR4 (N1483, N1476, N1089, N316, N109);
or OR4 (N1484, N1480, N726, N551, N442);
or OR2 (N1485, N1475, N519);
or OR2 (N1486, N1452, N516);
nand NAND4 (N1487, N1485, N772, N829, N480);
buf BUF1 (N1488, N1487);
buf BUF1 (N1489, N1483);
not NOT1 (N1490, N1466);
and AND4 (N1491, N1484, N1324, N898, N157);
nand NAND3 (N1492, N1491, N811, N910);
or OR4 (N1493, N1477, N1428, N1313, N336);
not NOT1 (N1494, N1490);
xor XOR2 (N1495, N1488, N406);
nand NAND3 (N1496, N1481, N170, N816);
not NOT1 (N1497, N1479);
buf BUF1 (N1498, N1495);
nor NOR2 (N1499, N1496, N210);
and AND4 (N1500, N1492, N571, N485, N223);
nor NOR2 (N1501, N1499, N1401);
not NOT1 (N1502, N1498);
buf BUF1 (N1503, N1500);
or OR4 (N1504, N1502, N554, N41, N791);
xor XOR2 (N1505, N1501, N1208);
and AND4 (N1506, N1494, N700, N1374, N33);
and AND2 (N1507, N1497, N888);
buf BUF1 (N1508, N1505);
or OR2 (N1509, N1489, N268);
nand NAND4 (N1510, N1493, N582, N1246, N1300);
xor XOR2 (N1511, N1503, N807);
not NOT1 (N1512, N1508);
not NOT1 (N1513, N1486);
not NOT1 (N1514, N1482);
buf BUF1 (N1515, N1511);
buf BUF1 (N1516, N1510);
xor XOR2 (N1517, N1506, N1238);
xor XOR2 (N1518, N1517, N382);
xor XOR2 (N1519, N1468, N367);
nor NOR2 (N1520, N1504, N838);
or OR2 (N1521, N1516, N12);
and AND4 (N1522, N1513, N317, N1236, N295);
buf BUF1 (N1523, N1520);
nor NOR4 (N1524, N1523, N1520, N420, N1287);
or OR2 (N1525, N1512, N763);
nor NOR3 (N1526, N1522, N1177, N96);
xor XOR2 (N1527, N1507, N921);
buf BUF1 (N1528, N1514);
buf BUF1 (N1529, N1518);
or OR3 (N1530, N1525, N66, N532);
or OR3 (N1531, N1530, N748, N1328);
nand NAND3 (N1532, N1519, N79, N138);
and AND2 (N1533, N1526, N782);
nand NAND2 (N1534, N1531, N1394);
not NOT1 (N1535, N1529);
or OR3 (N1536, N1533, N1256, N801);
or OR3 (N1537, N1534, N987, N1211);
and AND3 (N1538, N1536, N340, N1163);
xor XOR2 (N1539, N1509, N1431);
and AND4 (N1540, N1524, N971, N1180, N280);
buf BUF1 (N1541, N1527);
not NOT1 (N1542, N1515);
xor XOR2 (N1543, N1528, N1527);
nand NAND2 (N1544, N1538, N1527);
nor NOR2 (N1545, N1539, N1124);
not NOT1 (N1546, N1537);
not NOT1 (N1547, N1540);
xor XOR2 (N1548, N1521, N1451);
or OR4 (N1549, N1543, N1459, N1449, N136);
or OR3 (N1550, N1535, N622, N696);
and AND2 (N1551, N1550, N10);
buf BUF1 (N1552, N1544);
or OR3 (N1553, N1548, N1434, N163);
or OR2 (N1554, N1553, N1317);
or OR4 (N1555, N1547, N812, N47, N236);
not NOT1 (N1556, N1552);
xor XOR2 (N1557, N1541, N565);
nor NOR3 (N1558, N1554, N860, N601);
xor XOR2 (N1559, N1542, N104);
nand NAND3 (N1560, N1558, N372, N1127);
xor XOR2 (N1561, N1559, N53);
nor NOR3 (N1562, N1549, N551, N1210);
nand NAND4 (N1563, N1551, N1399, N317, N280);
buf BUF1 (N1564, N1555);
nor NOR3 (N1565, N1562, N1064, N132);
nor NOR4 (N1566, N1545, N1239, N1372, N1071);
nor NOR4 (N1567, N1565, N52, N253, N1208);
not NOT1 (N1568, N1561);
or OR2 (N1569, N1567, N717);
buf BUF1 (N1570, N1569);
and AND3 (N1571, N1532, N1376, N307);
nand NAND2 (N1572, N1560, N1123);
or OR4 (N1573, N1572, N742, N547, N1155);
or OR4 (N1574, N1563, N776, N957, N234);
buf BUF1 (N1575, N1568);
and AND4 (N1576, N1556, N572, N1445, N1242);
nand NAND3 (N1577, N1546, N1030, N121);
and AND4 (N1578, N1576, N40, N510, N740);
nand NAND2 (N1579, N1577, N1095);
buf BUF1 (N1580, N1573);
xor XOR2 (N1581, N1564, N1264);
nor NOR2 (N1582, N1566, N1018);
nor NOR4 (N1583, N1575, N373, N1450, N137);
and AND2 (N1584, N1557, N1296);
or OR3 (N1585, N1571, N539, N1427);
nor NOR4 (N1586, N1570, N1431, N1307, N1408);
and AND2 (N1587, N1574, N1226);
not NOT1 (N1588, N1587);
nor NOR2 (N1589, N1581, N1556);
xor XOR2 (N1590, N1586, N217);
nand NAND2 (N1591, N1580, N786);
buf BUF1 (N1592, N1590);
buf BUF1 (N1593, N1584);
and AND2 (N1594, N1589, N421);
and AND2 (N1595, N1583, N256);
xor XOR2 (N1596, N1588, N981);
and AND4 (N1597, N1592, N597, N880, N966);
xor XOR2 (N1598, N1582, N632);
not NOT1 (N1599, N1597);
or OR3 (N1600, N1579, N1216, N168);
not NOT1 (N1601, N1591);
nor NOR2 (N1602, N1596, N1489);
xor XOR2 (N1603, N1578, N484);
nand NAND4 (N1604, N1593, N343, N1475, N1051);
xor XOR2 (N1605, N1600, N821);
nor NOR4 (N1606, N1602, N35, N797, N744);
buf BUF1 (N1607, N1598);
and AND2 (N1608, N1585, N8);
or OR2 (N1609, N1601, N111);
nor NOR2 (N1610, N1603, N1190);
nand NAND3 (N1611, N1609, N253, N613);
nand NAND3 (N1612, N1610, N174, N1531);
not NOT1 (N1613, N1611);
xor XOR2 (N1614, N1595, N670);
nand NAND3 (N1615, N1607, N1123, N1297);
buf BUF1 (N1616, N1605);
buf BUF1 (N1617, N1594);
nand NAND3 (N1618, N1604, N737, N1434);
or OR4 (N1619, N1615, N1473, N677, N199);
not NOT1 (N1620, N1617);
and AND2 (N1621, N1599, N551);
not NOT1 (N1622, N1606);
xor XOR2 (N1623, N1614, N245);
nand NAND4 (N1624, N1612, N1595, N1528, N1364);
nor NOR2 (N1625, N1616, N1285);
and AND2 (N1626, N1618, N826);
nor NOR2 (N1627, N1626, N1519);
nor NOR3 (N1628, N1623, N1110, N1163);
or OR4 (N1629, N1619, N1093, N357, N1097);
not NOT1 (N1630, N1627);
xor XOR2 (N1631, N1630, N451);
and AND2 (N1632, N1613, N723);
and AND3 (N1633, N1608, N1327, N120);
not NOT1 (N1634, N1621);
buf BUF1 (N1635, N1633);
buf BUF1 (N1636, N1625);
buf BUF1 (N1637, N1635);
xor XOR2 (N1638, N1624, N1054);
or OR2 (N1639, N1620, N1102);
nor NOR2 (N1640, N1636, N98);
or OR3 (N1641, N1639, N681, N674);
not NOT1 (N1642, N1641);
or OR2 (N1643, N1634, N1008);
not NOT1 (N1644, N1640);
nand NAND2 (N1645, N1632, N1162);
not NOT1 (N1646, N1637);
nand NAND3 (N1647, N1628, N1116, N1019);
or OR4 (N1648, N1638, N363, N715, N1392);
nand NAND2 (N1649, N1645, N526);
xor XOR2 (N1650, N1642, N1105);
and AND3 (N1651, N1644, N86, N974);
and AND3 (N1652, N1629, N145, N607);
not NOT1 (N1653, N1649);
and AND2 (N1654, N1647, N223);
xor XOR2 (N1655, N1648, N633);
not NOT1 (N1656, N1655);
nand NAND3 (N1657, N1622, N1139, N1096);
buf BUF1 (N1658, N1654);
or OR4 (N1659, N1658, N808, N165, N1193);
buf BUF1 (N1660, N1643);
xor XOR2 (N1661, N1657, N1269);
buf BUF1 (N1662, N1659);
nor NOR2 (N1663, N1651, N291);
xor XOR2 (N1664, N1650, N1253);
xor XOR2 (N1665, N1662, N106);
buf BUF1 (N1666, N1656);
and AND2 (N1667, N1646, N1555);
xor XOR2 (N1668, N1660, N330);
not NOT1 (N1669, N1653);
buf BUF1 (N1670, N1668);
not NOT1 (N1671, N1664);
nand NAND4 (N1672, N1631, N1363, N164, N365);
or OR3 (N1673, N1670, N90, N734);
buf BUF1 (N1674, N1673);
nand NAND4 (N1675, N1666, N898, N1352, N180);
not NOT1 (N1676, N1672);
nand NAND4 (N1677, N1652, N558, N472, N763);
or OR2 (N1678, N1665, N956);
and AND3 (N1679, N1675, N7, N688);
buf BUF1 (N1680, N1671);
or OR2 (N1681, N1677, N66);
not NOT1 (N1682, N1678);
nand NAND2 (N1683, N1679, N425);
and AND4 (N1684, N1674, N433, N1232, N1439);
or OR3 (N1685, N1676, N1461, N117);
nand NAND2 (N1686, N1669, N1349);
and AND3 (N1687, N1663, N1686, N1499);
buf BUF1 (N1688, N1249);
buf BUF1 (N1689, N1685);
nand NAND4 (N1690, N1682, N296, N1655, N887);
not NOT1 (N1691, N1688);
and AND4 (N1692, N1689, N1402, N650, N1265);
not NOT1 (N1693, N1680);
not NOT1 (N1694, N1684);
and AND4 (N1695, N1661, N551, N235, N1597);
buf BUF1 (N1696, N1681);
nand NAND3 (N1697, N1691, N999, N689);
not NOT1 (N1698, N1696);
xor XOR2 (N1699, N1697, N457);
and AND2 (N1700, N1695, N573);
xor XOR2 (N1701, N1687, N990);
nand NAND4 (N1702, N1694, N1255, N416, N299);
or OR2 (N1703, N1698, N351);
nor NOR4 (N1704, N1701, N559, N142, N526);
nor NOR4 (N1705, N1703, N1575, N1473, N1425);
not NOT1 (N1706, N1700);
and AND2 (N1707, N1667, N1436);
not NOT1 (N1708, N1683);
nand NAND4 (N1709, N1706, N402, N1171, N601);
or OR4 (N1710, N1704, N1308, N1607, N63);
and AND4 (N1711, N1708, N1178, N1559, N25);
and AND3 (N1712, N1690, N1114, N283);
xor XOR2 (N1713, N1710, N1065);
not NOT1 (N1714, N1711);
or OR4 (N1715, N1699, N265, N212, N555);
not NOT1 (N1716, N1693);
nor NOR2 (N1717, N1707, N794);
nor NOR2 (N1718, N1716, N1540);
nor NOR3 (N1719, N1717, N106, N615);
nor NOR4 (N1720, N1705, N978, N659, N1216);
not NOT1 (N1721, N1702);
and AND4 (N1722, N1715, N808, N99, N93);
nand NAND3 (N1723, N1719, N421, N1008);
or OR3 (N1724, N1714, N1202, N564);
or OR2 (N1725, N1713, N1188);
or OR3 (N1726, N1709, N558, N875);
nor NOR3 (N1727, N1712, N1, N1195);
nor NOR4 (N1728, N1721, N233, N834, N439);
nand NAND2 (N1729, N1725, N1661);
not NOT1 (N1730, N1726);
buf BUF1 (N1731, N1722);
xor XOR2 (N1732, N1718, N441);
nor NOR2 (N1733, N1732, N1540);
buf BUF1 (N1734, N1720);
not NOT1 (N1735, N1727);
or OR2 (N1736, N1728, N389);
xor XOR2 (N1737, N1724, N1096);
nor NOR3 (N1738, N1734, N1356, N1488);
or OR4 (N1739, N1692, N1279, N566, N699);
or OR2 (N1740, N1729, N1217);
buf BUF1 (N1741, N1723);
and AND3 (N1742, N1741, N11, N659);
buf BUF1 (N1743, N1730);
nand NAND4 (N1744, N1733, N115, N912, N1019);
and AND3 (N1745, N1739, N1006, N1593);
nor NOR3 (N1746, N1745, N34, N812);
nand NAND4 (N1747, N1735, N1335, N453, N639);
or OR2 (N1748, N1740, N820);
not NOT1 (N1749, N1744);
or OR3 (N1750, N1747, N277, N1279);
xor XOR2 (N1751, N1746, N198);
not NOT1 (N1752, N1743);
not NOT1 (N1753, N1748);
and AND2 (N1754, N1753, N1666);
or OR3 (N1755, N1737, N448, N53);
xor XOR2 (N1756, N1755, N1685);
nand NAND3 (N1757, N1750, N771, N1294);
and AND3 (N1758, N1742, N1291, N635);
buf BUF1 (N1759, N1751);
buf BUF1 (N1760, N1754);
and AND2 (N1761, N1749, N953);
nor NOR2 (N1762, N1757, N1740);
buf BUF1 (N1763, N1756);
or OR3 (N1764, N1761, N1360, N549);
not NOT1 (N1765, N1736);
nor NOR2 (N1766, N1765, N229);
or OR2 (N1767, N1752, N1578);
or OR3 (N1768, N1731, N1415, N314);
buf BUF1 (N1769, N1768);
nor NOR3 (N1770, N1759, N59, N790);
and AND4 (N1771, N1738, N553, N1643, N519);
and AND3 (N1772, N1762, N1603, N1113);
not NOT1 (N1773, N1764);
not NOT1 (N1774, N1766);
nor NOR4 (N1775, N1763, N1731, N1567, N1169);
or OR4 (N1776, N1775, N754, N1172, N838);
and AND3 (N1777, N1769, N797, N1281);
nand NAND2 (N1778, N1758, N785);
xor XOR2 (N1779, N1771, N630);
nand NAND2 (N1780, N1770, N1583);
xor XOR2 (N1781, N1780, N982);
xor XOR2 (N1782, N1776, N837);
and AND4 (N1783, N1772, N444, N589, N1489);
nor NOR2 (N1784, N1774, N419);
buf BUF1 (N1785, N1773);
xor XOR2 (N1786, N1760, N954);
xor XOR2 (N1787, N1779, N1056);
and AND3 (N1788, N1781, N1550, N1467);
nor NOR4 (N1789, N1782, N606, N310, N166);
buf BUF1 (N1790, N1767);
or OR4 (N1791, N1787, N1340, N1523, N1611);
nor NOR2 (N1792, N1788, N916);
xor XOR2 (N1793, N1777, N576);
buf BUF1 (N1794, N1778);
or OR3 (N1795, N1791, N679, N247);
nor NOR2 (N1796, N1795, N101);
xor XOR2 (N1797, N1783, N720);
nor NOR2 (N1798, N1786, N319);
buf BUF1 (N1799, N1792);
not NOT1 (N1800, N1794);
xor XOR2 (N1801, N1789, N514);
nor NOR4 (N1802, N1785, N1171, N630, N1191);
nor NOR4 (N1803, N1799, N364, N1088, N1050);
nor NOR3 (N1804, N1802, N542, N1331);
buf BUF1 (N1805, N1800);
or OR3 (N1806, N1804, N1212, N25);
or OR4 (N1807, N1797, N1716, N79, N1781);
buf BUF1 (N1808, N1796);
and AND2 (N1809, N1807, N872);
and AND3 (N1810, N1808, N645, N1564);
or OR2 (N1811, N1784, N62);
and AND2 (N1812, N1810, N1779);
and AND4 (N1813, N1811, N1089, N199, N737);
buf BUF1 (N1814, N1790);
or OR4 (N1815, N1813, N453, N1775, N296);
nor NOR3 (N1816, N1801, N757, N434);
nor NOR2 (N1817, N1798, N700);
not NOT1 (N1818, N1805);
nor NOR2 (N1819, N1815, N1059);
or OR3 (N1820, N1803, N939, N576);
buf BUF1 (N1821, N1819);
nand NAND4 (N1822, N1816, N757, N1332, N231);
and AND4 (N1823, N1809, N381, N859, N1060);
xor XOR2 (N1824, N1823, N727);
xor XOR2 (N1825, N1806, N917);
or OR2 (N1826, N1793, N598);
or OR3 (N1827, N1822, N251, N371);
and AND4 (N1828, N1812, N900, N313, N1632);
buf BUF1 (N1829, N1821);
not NOT1 (N1830, N1825);
nor NOR4 (N1831, N1827, N325, N1507, N893);
nand NAND3 (N1832, N1818, N463, N1775);
nor NOR4 (N1833, N1826, N1747, N888, N935);
buf BUF1 (N1834, N1820);
not NOT1 (N1835, N1824);
and AND4 (N1836, N1834, N835, N1783, N286);
not NOT1 (N1837, N1817);
xor XOR2 (N1838, N1837, N1198);
and AND2 (N1839, N1828, N1553);
nor NOR3 (N1840, N1839, N1746, N225);
not NOT1 (N1841, N1833);
nor NOR3 (N1842, N1814, N489, N656);
xor XOR2 (N1843, N1836, N1763);
nor NOR4 (N1844, N1835, N515, N1731, N728);
nor NOR4 (N1845, N1830, N473, N57, N1657);
not NOT1 (N1846, N1832);
not NOT1 (N1847, N1845);
or OR4 (N1848, N1847, N1299, N775, N1422);
not NOT1 (N1849, N1829);
buf BUF1 (N1850, N1842);
xor XOR2 (N1851, N1840, N81);
not NOT1 (N1852, N1843);
nor NOR4 (N1853, N1851, N218, N1336, N1665);
not NOT1 (N1854, N1844);
xor XOR2 (N1855, N1852, N637);
or OR4 (N1856, N1846, N1836, N1223, N1757);
and AND2 (N1857, N1853, N824);
nor NOR2 (N1858, N1850, N1411);
or OR4 (N1859, N1841, N1720, N1722, N885);
not NOT1 (N1860, N1859);
nor NOR3 (N1861, N1860, N1761, N1743);
buf BUF1 (N1862, N1854);
and AND2 (N1863, N1838, N1054);
nand NAND2 (N1864, N1849, N1617);
or OR2 (N1865, N1856, N1752);
and AND2 (N1866, N1848, N1426);
xor XOR2 (N1867, N1861, N211);
nor NOR2 (N1868, N1831, N1788);
nor NOR3 (N1869, N1855, N1003, N491);
and AND3 (N1870, N1868, N1302, N143);
nand NAND2 (N1871, N1864, N1391);
and AND2 (N1872, N1858, N1549);
not NOT1 (N1873, N1863);
xor XOR2 (N1874, N1867, N1503);
or OR3 (N1875, N1869, N1397, N1317);
and AND4 (N1876, N1866, N1805, N87, N1079);
not NOT1 (N1877, N1865);
and AND3 (N1878, N1857, N169, N79);
buf BUF1 (N1879, N1875);
xor XOR2 (N1880, N1871, N1117);
not NOT1 (N1881, N1874);
not NOT1 (N1882, N1862);
buf BUF1 (N1883, N1878);
nor NOR3 (N1884, N1876, N1263, N425);
buf BUF1 (N1885, N1883);
buf BUF1 (N1886, N1873);
buf BUF1 (N1887, N1872);
buf BUF1 (N1888, N1886);
not NOT1 (N1889, N1884);
nor NOR2 (N1890, N1879, N1593);
nand NAND2 (N1891, N1890, N1447);
xor XOR2 (N1892, N1877, N923);
not NOT1 (N1893, N1888);
nand NAND4 (N1894, N1882, N1460, N1676, N1729);
nand NAND2 (N1895, N1891, N1776);
or OR2 (N1896, N1894, N1165);
nand NAND3 (N1897, N1870, N633, N1253);
buf BUF1 (N1898, N1897);
nor NOR2 (N1899, N1893, N705);
and AND3 (N1900, N1895, N1423, N1777);
buf BUF1 (N1901, N1881);
xor XOR2 (N1902, N1901, N1221);
and AND3 (N1903, N1892, N762, N954);
buf BUF1 (N1904, N1880);
nor NOR3 (N1905, N1896, N204, N838);
buf BUF1 (N1906, N1887);
xor XOR2 (N1907, N1905, N1328);
nor NOR2 (N1908, N1898, N1449);
and AND2 (N1909, N1903, N1781);
not NOT1 (N1910, N1904);
xor XOR2 (N1911, N1907, N1108);
nand NAND2 (N1912, N1910, N1547);
nor NOR3 (N1913, N1899, N1785, N22);
buf BUF1 (N1914, N1885);
nand NAND2 (N1915, N1889, N1601);
and AND3 (N1916, N1912, N757, N136);
nor NOR4 (N1917, N1914, N1518, N1708, N1572);
or OR2 (N1918, N1915, N1475);
or OR4 (N1919, N1906, N1705, N382, N494);
buf BUF1 (N1920, N1909);
nand NAND4 (N1921, N1902, N1209, N929, N799);
nand NAND3 (N1922, N1916, N517, N351);
or OR2 (N1923, N1921, N16);
or OR2 (N1924, N1923, N1671);
nand NAND2 (N1925, N1918, N1387);
nand NAND4 (N1926, N1919, N1258, N1436, N1320);
or OR3 (N1927, N1920, N293, N955);
not NOT1 (N1928, N1926);
and AND3 (N1929, N1922, N50, N1173);
nor NOR4 (N1930, N1908, N1690, N1599, N255);
xor XOR2 (N1931, N1924, N1385);
or OR2 (N1932, N1917, N1201);
and AND2 (N1933, N1900, N1357);
xor XOR2 (N1934, N1928, N512);
not NOT1 (N1935, N1911);
not NOT1 (N1936, N1925);
not NOT1 (N1937, N1935);
nand NAND4 (N1938, N1927, N1465, N1899, N1399);
xor XOR2 (N1939, N1931, N1663);
or OR4 (N1940, N1913, N363, N923, N711);
or OR2 (N1941, N1940, N1530);
buf BUF1 (N1942, N1939);
nor NOR2 (N1943, N1942, N426);
xor XOR2 (N1944, N1932, N1190);
and AND3 (N1945, N1938, N1754, N649);
xor XOR2 (N1946, N1934, N612);
not NOT1 (N1947, N1943);
and AND3 (N1948, N1941, N1085, N1899);
buf BUF1 (N1949, N1937);
and AND4 (N1950, N1947, N1267, N1574, N81);
or OR2 (N1951, N1948, N1127);
buf BUF1 (N1952, N1945);
xor XOR2 (N1953, N1933, N1537);
xor XOR2 (N1954, N1936, N1007);
or OR4 (N1955, N1930, N1395, N789, N391);
xor XOR2 (N1956, N1950, N603);
and AND4 (N1957, N1954, N186, N1218, N1057);
not NOT1 (N1958, N1955);
xor XOR2 (N1959, N1929, N1071);
nand NAND2 (N1960, N1957, N1039);
nand NAND4 (N1961, N1959, N753, N153, N645);
nor NOR2 (N1962, N1961, N945);
or OR4 (N1963, N1951, N671, N1736, N1385);
nand NAND3 (N1964, N1949, N1402, N1705);
or OR2 (N1965, N1962, N455);
or OR3 (N1966, N1952, N652, N1012);
nand NAND2 (N1967, N1958, N926);
nand NAND4 (N1968, N1967, N209, N484, N171);
and AND3 (N1969, N1964, N1188, N1693);
and AND3 (N1970, N1969, N689, N1793);
buf BUF1 (N1971, N1946);
or OR2 (N1972, N1960, N499);
xor XOR2 (N1973, N1963, N465);
buf BUF1 (N1974, N1956);
and AND2 (N1975, N1973, N152);
xor XOR2 (N1976, N1944, N959);
not NOT1 (N1977, N1970);
not NOT1 (N1978, N1953);
or OR4 (N1979, N1977, N1796, N1106, N528);
and AND3 (N1980, N1965, N710, N1343);
buf BUF1 (N1981, N1974);
or OR2 (N1982, N1971, N1550);
buf BUF1 (N1983, N1972);
xor XOR2 (N1984, N1968, N913);
not NOT1 (N1985, N1984);
buf BUF1 (N1986, N1966);
nand NAND3 (N1987, N1986, N1484, N121);
nor NOR2 (N1988, N1985, N740);
nand NAND2 (N1989, N1988, N473);
not NOT1 (N1990, N1979);
and AND2 (N1991, N1983, N706);
or OR3 (N1992, N1987, N1655, N676);
buf BUF1 (N1993, N1980);
nor NOR3 (N1994, N1978, N1378, N693);
nand NAND2 (N1995, N1991, N743);
not NOT1 (N1996, N1994);
not NOT1 (N1997, N1989);
not NOT1 (N1998, N1990);
and AND2 (N1999, N1975, N216);
xor XOR2 (N2000, N1982, N523);
xor XOR2 (N2001, N1999, N346);
not NOT1 (N2002, N2001);
or OR2 (N2003, N1997, N1833);
buf BUF1 (N2004, N2002);
not NOT1 (N2005, N1998);
and AND4 (N2006, N1996, N1281, N762, N1401);
xor XOR2 (N2007, N2006, N1075);
nor NOR4 (N2008, N1995, N336, N201, N113);
xor XOR2 (N2009, N1981, N17);
or OR3 (N2010, N2008, N814, N753);
nand NAND3 (N2011, N2007, N2001, N796);
and AND3 (N2012, N2004, N1452, N445);
nand NAND2 (N2013, N2010, N784);
buf BUF1 (N2014, N2009);
nand NAND2 (N2015, N2003, N1934);
nor NOR4 (N2016, N1976, N1099, N1227, N1696);
not NOT1 (N2017, N2012);
and AND3 (N2018, N2017, N736, N1871);
and AND4 (N2019, N1992, N1505, N1678, N127);
and AND3 (N2020, N2000, N1980, N702);
or OR4 (N2021, N2020, N1969, N202, N1755);
nor NOR2 (N2022, N2019, N1550);
xor XOR2 (N2023, N2018, N1937);
not NOT1 (N2024, N2014);
not NOT1 (N2025, N2022);
nand NAND2 (N2026, N2016, N1267);
and AND3 (N2027, N2025, N1393, N614);
or OR4 (N2028, N2027, N1119, N657, N1621);
nor NOR2 (N2029, N1993, N1853);
xor XOR2 (N2030, N2028, N1035);
nor NOR4 (N2031, N2023, N1536, N1677, N1955);
buf BUF1 (N2032, N2026);
nor NOR2 (N2033, N2013, N1039);
or OR3 (N2034, N2015, N1118, N1570);
and AND3 (N2035, N2005, N591, N378);
buf BUF1 (N2036, N2030);
buf BUF1 (N2037, N2035);
xor XOR2 (N2038, N2032, N1062);
nor NOR2 (N2039, N2034, N573);
buf BUF1 (N2040, N2011);
xor XOR2 (N2041, N2036, N1553);
not NOT1 (N2042, N2021);
xor XOR2 (N2043, N2039, N843);
buf BUF1 (N2044, N2038);
buf BUF1 (N2045, N2031);
or OR2 (N2046, N2045, N1671);
xor XOR2 (N2047, N2044, N1100);
xor XOR2 (N2048, N2047, N965);
or OR2 (N2049, N2029, N1242);
not NOT1 (N2050, N2040);
xor XOR2 (N2051, N2048, N333);
and AND4 (N2052, N2050, N672, N1134, N271);
or OR2 (N2053, N2033, N1456);
xor XOR2 (N2054, N2042, N234);
xor XOR2 (N2055, N2053, N1882);
not NOT1 (N2056, N2024);
not NOT1 (N2057, N2043);
nor NOR3 (N2058, N2057, N1015, N689);
not NOT1 (N2059, N2046);
not NOT1 (N2060, N2058);
buf BUF1 (N2061, N2059);
not NOT1 (N2062, N2037);
and AND2 (N2063, N2052, N64);
xor XOR2 (N2064, N2041, N1736);
buf BUF1 (N2065, N2054);
xor XOR2 (N2066, N2051, N2000);
xor XOR2 (N2067, N2066, N441);
or OR3 (N2068, N2063, N1977, N1280);
not NOT1 (N2069, N2067);
not NOT1 (N2070, N2056);
nand NAND2 (N2071, N2068, N1747);
and AND4 (N2072, N2065, N1988, N15, N835);
nand NAND2 (N2073, N2061, N821);
not NOT1 (N2074, N2070);
not NOT1 (N2075, N2064);
nor NOR2 (N2076, N2060, N6);
and AND4 (N2077, N2071, N1679, N1290, N1826);
and AND4 (N2078, N2077, N675, N1927, N1753);
buf BUF1 (N2079, N2072);
nand NAND4 (N2080, N2073, N1722, N1908, N1097);
nand NAND2 (N2081, N2079, N1721);
not NOT1 (N2082, N2049);
not NOT1 (N2083, N2069);
buf BUF1 (N2084, N2078);
and AND4 (N2085, N2075, N740, N1195, N542);
buf BUF1 (N2086, N2081);
not NOT1 (N2087, N2055);
or OR4 (N2088, N2076, N224, N731, N2002);
nor NOR2 (N2089, N2074, N685);
buf BUF1 (N2090, N2088);
and AND3 (N2091, N2090, N249, N1626);
not NOT1 (N2092, N2084);
and AND4 (N2093, N2062, N518, N881, N612);
nor NOR3 (N2094, N2082, N2032, N73);
xor XOR2 (N2095, N2089, N1396);
nor NOR2 (N2096, N2087, N2087);
nand NAND4 (N2097, N2095, N379, N910, N1868);
nand NAND3 (N2098, N2080, N1593, N1672);
buf BUF1 (N2099, N2098);
not NOT1 (N2100, N2097);
nand NAND4 (N2101, N2085, N1710, N1056, N823);
or OR4 (N2102, N2100, N1142, N1894, N793);
nand NAND2 (N2103, N2102, N880);
buf BUF1 (N2104, N2083);
buf BUF1 (N2105, N2091);
nand NAND4 (N2106, N2092, N9, N2101, N866);
xor XOR2 (N2107, N1141, N1140);
or OR2 (N2108, N2104, N1936);
not NOT1 (N2109, N2106);
xor XOR2 (N2110, N2094, N422);
nor NOR3 (N2111, N2108, N1144, N2063);
buf BUF1 (N2112, N2109);
xor XOR2 (N2113, N2111, N922);
nor NOR4 (N2114, N2103, N779, N2076, N1621);
buf BUF1 (N2115, N2105);
and AND4 (N2116, N2096, N1419, N684, N240);
nand NAND4 (N2117, N2115, N1353, N1464, N1851);
or OR4 (N2118, N2116, N1001, N1381, N738);
not NOT1 (N2119, N2113);
buf BUF1 (N2120, N2107);
xor XOR2 (N2121, N2099, N1128);
nor NOR2 (N2122, N2086, N2059);
xor XOR2 (N2123, N2110, N1722);
or OR2 (N2124, N2122, N739);
or OR2 (N2125, N2123, N1592);
not NOT1 (N2126, N2114);
nor NOR4 (N2127, N2124, N293, N79, N481);
nand NAND4 (N2128, N2119, N1663, N50, N1190);
or OR3 (N2129, N2093, N993, N168);
and AND2 (N2130, N2118, N1492);
and AND4 (N2131, N2121, N1962, N1706, N306);
xor XOR2 (N2132, N2125, N1531);
nand NAND2 (N2133, N2131, N1724);
nor NOR4 (N2134, N2129, N220, N2036, N959);
xor XOR2 (N2135, N2112, N1333);
and AND4 (N2136, N2135, N1092, N1163, N957);
not NOT1 (N2137, N2133);
xor XOR2 (N2138, N2130, N1390);
or OR4 (N2139, N2117, N1748, N834, N1614);
or OR4 (N2140, N2120, N888, N483, N2063);
nor NOR4 (N2141, N2137, N1270, N267, N207);
xor XOR2 (N2142, N2128, N1321);
xor XOR2 (N2143, N2136, N1617);
not NOT1 (N2144, N2126);
buf BUF1 (N2145, N2143);
or OR3 (N2146, N2132, N1082, N1943);
and AND3 (N2147, N2139, N914, N620);
xor XOR2 (N2148, N2145, N1573);
nor NOR2 (N2149, N2141, N797);
nand NAND4 (N2150, N2146, N958, N757, N1215);
or OR2 (N2151, N2144, N1213);
xor XOR2 (N2152, N2149, N252);
and AND2 (N2153, N2151, N603);
nor NOR2 (N2154, N2148, N1109);
and AND2 (N2155, N2138, N346);
or OR4 (N2156, N2147, N991, N33, N1116);
or OR4 (N2157, N2156, N1754, N1875, N1654);
nand NAND2 (N2158, N2140, N1332);
buf BUF1 (N2159, N2154);
or OR3 (N2160, N2155, N836, N1167);
nor NOR2 (N2161, N2160, N1787);
xor XOR2 (N2162, N2134, N1491);
nor NOR3 (N2163, N2161, N309, N1586);
xor XOR2 (N2164, N2157, N1686);
nor NOR4 (N2165, N2159, N1186, N720, N2107);
not NOT1 (N2166, N2158);
nand NAND2 (N2167, N2163, N192);
or OR2 (N2168, N2164, N1775);
nand NAND2 (N2169, N2127, N479);
buf BUF1 (N2170, N2165);
xor XOR2 (N2171, N2152, N1776);
nor NOR4 (N2172, N2168, N1893, N1493, N1793);
not NOT1 (N2173, N2170);
not NOT1 (N2174, N2171);
buf BUF1 (N2175, N2172);
or OR4 (N2176, N2162, N2094, N1435, N940);
and AND4 (N2177, N2167, N480, N924, N913);
buf BUF1 (N2178, N2175);
and AND4 (N2179, N2178, N2021, N2004, N1162);
nand NAND2 (N2180, N2166, N196);
not NOT1 (N2181, N2177);
xor XOR2 (N2182, N2142, N1707);
nor NOR4 (N2183, N2181, N1430, N2149, N1020);
not NOT1 (N2184, N2179);
and AND2 (N2185, N2176, N956);
nand NAND4 (N2186, N2153, N361, N2082, N854);
xor XOR2 (N2187, N2184, N1433);
buf BUF1 (N2188, N2182);
nor NOR3 (N2189, N2150, N554, N286);
buf BUF1 (N2190, N2169);
nand NAND4 (N2191, N2189, N1923, N501, N243);
nand NAND4 (N2192, N2180, N414, N2170, N1007);
not NOT1 (N2193, N2185);
nor NOR4 (N2194, N2190, N1822, N1398, N1754);
buf BUF1 (N2195, N2193);
nor NOR3 (N2196, N2192, N1360, N1118);
nand NAND4 (N2197, N2191, N327, N1992, N959);
nand NAND4 (N2198, N2196, N410, N930, N1356);
or OR4 (N2199, N2198, N837, N854, N1670);
xor XOR2 (N2200, N2174, N883);
nor NOR3 (N2201, N2173, N735, N80);
xor XOR2 (N2202, N2197, N2157);
not NOT1 (N2203, N2199);
nor NOR4 (N2204, N2188, N1136, N2130, N155);
nand NAND2 (N2205, N2200, N1595);
nor NOR4 (N2206, N2195, N1456, N1799, N1834);
not NOT1 (N2207, N2206);
nor NOR2 (N2208, N2201, N210);
nand NAND2 (N2209, N2208, N1111);
buf BUF1 (N2210, N2203);
not NOT1 (N2211, N2205);
buf BUF1 (N2212, N2183);
nor NOR4 (N2213, N2194, N934, N1915, N1);
nand NAND4 (N2214, N2207, N514, N682, N2129);
not NOT1 (N2215, N2204);
nand NAND2 (N2216, N2214, N588);
xor XOR2 (N2217, N2211, N493);
and AND2 (N2218, N2217, N981);
nand NAND2 (N2219, N2218, N1173);
nand NAND3 (N2220, N2210, N925, N1680);
nor NOR2 (N2221, N2219, N873);
or OR2 (N2222, N2209, N1592);
and AND4 (N2223, N2213, N1380, N85, N769);
xor XOR2 (N2224, N2186, N1410);
not NOT1 (N2225, N2220);
and AND4 (N2226, N2216, N1701, N835, N1481);
not NOT1 (N2227, N2187);
xor XOR2 (N2228, N2212, N813);
xor XOR2 (N2229, N2222, N1414);
nor NOR4 (N2230, N2202, N450, N462, N1055);
buf BUF1 (N2231, N2228);
nand NAND4 (N2232, N2221, N1116, N1137, N16);
not NOT1 (N2233, N2229);
or OR4 (N2234, N2233, N602, N89, N1804);
or OR2 (N2235, N2224, N483);
nand NAND2 (N2236, N2223, N1076);
or OR2 (N2237, N2231, N2093);
or OR3 (N2238, N2227, N2077, N583);
or OR2 (N2239, N2230, N1760);
not NOT1 (N2240, N2232);
not NOT1 (N2241, N2235);
xor XOR2 (N2242, N2239, N2200);
nand NAND4 (N2243, N2241, N2182, N1983, N297);
nand NAND3 (N2244, N2234, N2172, N1955);
nor NOR4 (N2245, N2238, N1692, N1281, N27);
xor XOR2 (N2246, N2237, N1056);
not NOT1 (N2247, N2236);
not NOT1 (N2248, N2242);
xor XOR2 (N2249, N2226, N2166);
or OR2 (N2250, N2215, N668);
buf BUF1 (N2251, N2247);
xor XOR2 (N2252, N2243, N579);
nand NAND3 (N2253, N2245, N1874, N371);
nor NOR4 (N2254, N2248, N1472, N1605, N904);
not NOT1 (N2255, N2250);
nor NOR3 (N2256, N2255, N807, N2093);
not NOT1 (N2257, N2253);
or OR4 (N2258, N2257, N1163, N868, N434);
nor NOR3 (N2259, N2244, N2198, N1711);
nor NOR3 (N2260, N2256, N1251, N170);
xor XOR2 (N2261, N2252, N133);
buf BUF1 (N2262, N2225);
and AND4 (N2263, N2251, N209, N862, N731);
xor XOR2 (N2264, N2262, N2039);
buf BUF1 (N2265, N2249);
nand NAND4 (N2266, N2254, N906, N93, N1953);
not NOT1 (N2267, N2265);
and AND2 (N2268, N2246, N1322);
and AND2 (N2269, N2268, N2225);
nand NAND3 (N2270, N2267, N1886, N1746);
nor NOR3 (N2271, N2259, N2256, N1359);
not NOT1 (N2272, N2269);
xor XOR2 (N2273, N2263, N418);
and AND2 (N2274, N2272, N1790);
buf BUF1 (N2275, N2264);
not NOT1 (N2276, N2240);
not NOT1 (N2277, N2274);
xor XOR2 (N2278, N2260, N1294);
xor XOR2 (N2279, N2271, N1460);
xor XOR2 (N2280, N2278, N2180);
nand NAND3 (N2281, N2258, N1113, N217);
xor XOR2 (N2282, N2277, N910);
nand NAND3 (N2283, N2261, N1048, N928);
nor NOR4 (N2284, N2276, N1974, N2196, N2062);
nor NOR3 (N2285, N2280, N205, N438);
not NOT1 (N2286, N2270);
buf BUF1 (N2287, N2281);
nor NOR3 (N2288, N2286, N449, N933);
buf BUF1 (N2289, N2273);
or OR2 (N2290, N2275, N1062);
and AND4 (N2291, N2266, N550, N253, N362);
nor NOR2 (N2292, N2283, N240);
nand NAND2 (N2293, N2285, N825);
buf BUF1 (N2294, N2282);
and AND2 (N2295, N2279, N2080);
and AND2 (N2296, N2291, N93);
buf BUF1 (N2297, N2290);
and AND3 (N2298, N2296, N1287, N1218);
and AND2 (N2299, N2292, N1566);
xor XOR2 (N2300, N2299, N1298);
buf BUF1 (N2301, N2284);
or OR3 (N2302, N2293, N1371, N1851);
nor NOR3 (N2303, N2294, N2149, N1608);
buf BUF1 (N2304, N2288);
nor NOR2 (N2305, N2304, N1036);
not NOT1 (N2306, N2303);
buf BUF1 (N2307, N2301);
buf BUF1 (N2308, N2297);
buf BUF1 (N2309, N2306);
not NOT1 (N2310, N2295);
nor NOR4 (N2311, N2300, N2013, N88, N2277);
buf BUF1 (N2312, N2302);
nand NAND2 (N2313, N2309, N1620);
nand NAND2 (N2314, N2307, N1370);
xor XOR2 (N2315, N2287, N383);
nor NOR3 (N2316, N2289, N2105, N1669);
buf BUF1 (N2317, N2298);
and AND2 (N2318, N2315, N455);
nor NOR2 (N2319, N2310, N600);
nand NAND2 (N2320, N2313, N1892);
nand NAND2 (N2321, N2312, N57);
buf BUF1 (N2322, N2308);
and AND3 (N2323, N2305, N695, N1578);
not NOT1 (N2324, N2320);
nor NOR2 (N2325, N2314, N2009);
or OR3 (N2326, N2318, N1322, N1853);
nor NOR4 (N2327, N2311, N474, N869, N763);
and AND4 (N2328, N2325, N885, N1940, N1751);
not NOT1 (N2329, N2323);
buf BUF1 (N2330, N2316);
buf BUF1 (N2331, N2324);
nor NOR2 (N2332, N2331, N1282);
nor NOR4 (N2333, N2329, N954, N34, N1887);
nand NAND4 (N2334, N2317, N1276, N2189, N1453);
not NOT1 (N2335, N2322);
nand NAND4 (N2336, N2333, N940, N1628, N2025);
nor NOR4 (N2337, N2321, N1217, N2316, N285);
and AND4 (N2338, N2330, N305, N308, N1818);
nor NOR3 (N2339, N2336, N1616, N1247);
or OR2 (N2340, N2339, N1222);
not NOT1 (N2341, N2327);
nor NOR4 (N2342, N2335, N699, N393, N340);
nand NAND2 (N2343, N2328, N1823);
nor NOR2 (N2344, N2319, N1529);
buf BUF1 (N2345, N2337);
or OR2 (N2346, N2344, N40);
xor XOR2 (N2347, N2341, N1893);
nand NAND4 (N2348, N2338, N2141, N474, N435);
not NOT1 (N2349, N2347);
nor NOR3 (N2350, N2332, N1361, N1147);
xor XOR2 (N2351, N2340, N1602);
and AND2 (N2352, N2345, N2336);
xor XOR2 (N2353, N2342, N1772);
and AND3 (N2354, N2351, N1261, N419);
buf BUF1 (N2355, N2343);
or OR3 (N2356, N2326, N2059, N216);
or OR2 (N2357, N2355, N728);
and AND4 (N2358, N2354, N496, N1352, N817);
nor NOR3 (N2359, N2356, N812, N1469);
not NOT1 (N2360, N2353);
not NOT1 (N2361, N2334);
not NOT1 (N2362, N2352);
buf BUF1 (N2363, N2349);
nor NOR3 (N2364, N2348, N1261, N2099);
xor XOR2 (N2365, N2350, N427);
buf BUF1 (N2366, N2361);
xor XOR2 (N2367, N2364, N2179);
nor NOR3 (N2368, N2346, N436, N2306);
and AND3 (N2369, N2366, N172, N784);
xor XOR2 (N2370, N2367, N436);
and AND2 (N2371, N2365, N730);
and AND3 (N2372, N2359, N39, N1151);
not NOT1 (N2373, N2371);
not NOT1 (N2374, N2357);
not NOT1 (N2375, N2372);
and AND3 (N2376, N2362, N553, N1499);
buf BUF1 (N2377, N2369);
buf BUF1 (N2378, N2376);
xor XOR2 (N2379, N2373, N587);
nand NAND3 (N2380, N2368, N1716, N594);
nor NOR3 (N2381, N2378, N1658, N557);
buf BUF1 (N2382, N2360);
and AND3 (N2383, N2370, N1628, N825);
xor XOR2 (N2384, N2374, N1910);
not NOT1 (N2385, N2363);
nand NAND2 (N2386, N2377, N2112);
buf BUF1 (N2387, N2384);
nor NOR3 (N2388, N2379, N327, N1565);
xor XOR2 (N2389, N2375, N2194);
xor XOR2 (N2390, N2386, N1466);
not NOT1 (N2391, N2383);
buf BUF1 (N2392, N2385);
and AND3 (N2393, N2380, N997, N1063);
not NOT1 (N2394, N2390);
and AND2 (N2395, N2393, N1115);
and AND3 (N2396, N2389, N2283, N635);
buf BUF1 (N2397, N2382);
buf BUF1 (N2398, N2387);
buf BUF1 (N2399, N2397);
and AND3 (N2400, N2394, N1679, N2205);
nand NAND2 (N2401, N2388, N1420);
not NOT1 (N2402, N2391);
nand NAND2 (N2403, N2396, N1590);
nand NAND3 (N2404, N2392, N468, N161);
not NOT1 (N2405, N2399);
or OR2 (N2406, N2398, N306);
nand NAND4 (N2407, N2404, N1994, N29, N808);
buf BUF1 (N2408, N2402);
or OR3 (N2409, N2395, N1948, N774);
nand NAND4 (N2410, N2405, N2303, N2098, N761);
nand NAND2 (N2411, N2410, N2261);
xor XOR2 (N2412, N2406, N2280);
nand NAND2 (N2413, N2407, N1903);
nor NOR4 (N2414, N2408, N236, N1638, N2404);
and AND3 (N2415, N2403, N1906, N822);
xor XOR2 (N2416, N2381, N1175);
nor NOR3 (N2417, N2413, N992, N2179);
or OR4 (N2418, N2411, N2046, N734, N844);
not NOT1 (N2419, N2401);
xor XOR2 (N2420, N2415, N302);
and AND4 (N2421, N2420, N419, N1562, N301);
not NOT1 (N2422, N2419);
or OR4 (N2423, N2416, N1553, N2133, N617);
nand NAND3 (N2424, N2400, N1742, N780);
not NOT1 (N2425, N2417);
and AND2 (N2426, N2421, N179);
and AND2 (N2427, N2426, N1542);
buf BUF1 (N2428, N2418);
nand NAND3 (N2429, N2423, N880, N120);
not NOT1 (N2430, N2425);
nand NAND4 (N2431, N2429, N1455, N1702, N1434);
and AND3 (N2432, N2427, N1643, N1256);
and AND4 (N2433, N2414, N366, N636, N1863);
not NOT1 (N2434, N2431);
nand NAND2 (N2435, N2409, N435);
and AND3 (N2436, N2432, N882, N1823);
and AND3 (N2437, N2435, N396, N733);
nand NAND3 (N2438, N2358, N348, N1885);
buf BUF1 (N2439, N2438);
not NOT1 (N2440, N2433);
xor XOR2 (N2441, N2434, N989);
nand NAND3 (N2442, N2412, N276, N2266);
xor XOR2 (N2443, N2430, N674);
nor NOR3 (N2444, N2422, N1341, N1673);
xor XOR2 (N2445, N2424, N640);
or OR3 (N2446, N2437, N1596, N463);
nand NAND4 (N2447, N2443, N1582, N622, N155);
nand NAND2 (N2448, N2436, N2352);
and AND4 (N2449, N2442, N481, N1293, N1878);
nand NAND4 (N2450, N2428, N2017, N1487, N1056);
xor XOR2 (N2451, N2446, N2037);
and AND3 (N2452, N2451, N273, N263);
nor NOR2 (N2453, N2447, N1925);
nand NAND3 (N2454, N2448, N1294, N2429);
nand NAND3 (N2455, N2450, N1203, N442);
buf BUF1 (N2456, N2455);
nand NAND4 (N2457, N2452, N552, N2419, N1447);
and AND2 (N2458, N2457, N2082);
or OR3 (N2459, N2458, N1327, N1993);
xor XOR2 (N2460, N2440, N2160);
nand NAND4 (N2461, N2439, N2433, N38, N1270);
and AND4 (N2462, N2449, N1338, N2159, N34);
not NOT1 (N2463, N2462);
and AND2 (N2464, N2441, N2340);
nor NOR4 (N2465, N2454, N655, N2097, N1677);
and AND3 (N2466, N2459, N2368, N778);
xor XOR2 (N2467, N2463, N1910);
nand NAND3 (N2468, N2453, N32, N2451);
nor NOR4 (N2469, N2460, N283, N2049, N1407);
nand NAND2 (N2470, N2468, N251);
nor NOR4 (N2471, N2467, N2262, N1811, N1241);
nand NAND2 (N2472, N2445, N119);
nor NOR2 (N2473, N2464, N2138);
nor NOR3 (N2474, N2470, N51, N1014);
buf BUF1 (N2475, N2466);
nor NOR3 (N2476, N2471, N2219, N340);
xor XOR2 (N2477, N2473, N143);
nand NAND3 (N2478, N2461, N1418, N1923);
or OR2 (N2479, N2465, N435);
nor NOR2 (N2480, N2479, N1010);
nor NOR2 (N2481, N2469, N1004);
nand NAND2 (N2482, N2478, N537);
nor NOR2 (N2483, N2472, N2237);
nand NAND4 (N2484, N2480, N2438, N2284, N2480);
not NOT1 (N2485, N2475);
and AND3 (N2486, N2444, N1187, N1358);
buf BUF1 (N2487, N2485);
and AND4 (N2488, N2486, N2203, N144, N160);
nor NOR3 (N2489, N2477, N1113, N878);
not NOT1 (N2490, N2488);
nand NAND4 (N2491, N2484, N415, N648, N2120);
or OR3 (N2492, N2476, N2131, N2022);
not NOT1 (N2493, N2492);
nand NAND4 (N2494, N2482, N2259, N1807, N477);
not NOT1 (N2495, N2487);
not NOT1 (N2496, N2489);
nand NAND4 (N2497, N2474, N196, N1147, N1399);
nand NAND2 (N2498, N2481, N252);
xor XOR2 (N2499, N2498, N192);
and AND4 (N2500, N2496, N147, N1675, N1042);
buf BUF1 (N2501, N2500);
nor NOR3 (N2502, N2456, N1034, N1735);
or OR2 (N2503, N2491, N1105);
buf BUF1 (N2504, N2497);
nor NOR3 (N2505, N2502, N1906, N1328);
and AND3 (N2506, N2503, N609, N468);
xor XOR2 (N2507, N2501, N389);
and AND2 (N2508, N2506, N256);
and AND4 (N2509, N2493, N968, N1328, N2188);
and AND2 (N2510, N2494, N1339);
and AND3 (N2511, N2510, N1112, N385);
or OR4 (N2512, N2505, N306, N2140, N1025);
nor NOR3 (N2513, N2507, N1106, N1551);
nand NAND2 (N2514, N2499, N336);
or OR2 (N2515, N2490, N2319);
and AND2 (N2516, N2515, N866);
buf BUF1 (N2517, N2513);
xor XOR2 (N2518, N2504, N2007);
xor XOR2 (N2519, N2483, N36);
and AND2 (N2520, N2512, N769);
or OR2 (N2521, N2511, N772);
nand NAND3 (N2522, N2519, N25, N2064);
buf BUF1 (N2523, N2509);
or OR4 (N2524, N2522, N2426, N1333, N16);
nor NOR2 (N2525, N2508, N1826);
nor NOR2 (N2526, N2520, N755);
nand NAND3 (N2527, N2524, N1845, N1482);
buf BUF1 (N2528, N2516);
not NOT1 (N2529, N2527);
nand NAND2 (N2530, N2529, N2170);
xor XOR2 (N2531, N2521, N2197);
or OR4 (N2532, N2517, N424, N570, N108);
buf BUF1 (N2533, N2532);
nand NAND4 (N2534, N2526, N2338, N2256, N2178);
or OR3 (N2535, N2523, N2415, N1775);
and AND4 (N2536, N2535, N2062, N295, N1657);
nor NOR4 (N2537, N2495, N806, N735, N1010);
not NOT1 (N2538, N2536);
or OR3 (N2539, N2530, N2494, N65);
not NOT1 (N2540, N2528);
nand NAND2 (N2541, N2538, N913);
nand NAND4 (N2542, N2541, N2229, N39, N1589);
nor NOR4 (N2543, N2539, N2263, N457, N2164);
or OR2 (N2544, N2531, N885);
nor NOR2 (N2545, N2537, N511);
and AND3 (N2546, N2543, N1130, N1880);
or OR4 (N2547, N2518, N1708, N1263, N285);
buf BUF1 (N2548, N2545);
or OR3 (N2549, N2544, N852, N2137);
buf BUF1 (N2550, N2546);
nor NOR2 (N2551, N2547, N365);
or OR4 (N2552, N2542, N1157, N1584, N1122);
buf BUF1 (N2553, N2533);
and AND4 (N2554, N2552, N493, N928, N372);
nor NOR4 (N2555, N2549, N1110, N1825, N16);
or OR4 (N2556, N2525, N1953, N210, N1854);
nand NAND3 (N2557, N2540, N979, N624);
and AND3 (N2558, N2556, N1234, N2143);
nor NOR4 (N2559, N2558, N2155, N833, N1677);
not NOT1 (N2560, N2557);
or OR3 (N2561, N2560, N834, N612);
and AND3 (N2562, N2548, N552, N1912);
nand NAND2 (N2563, N2554, N2129);
nor NOR2 (N2564, N2563, N1369);
nand NAND4 (N2565, N2555, N2390, N987, N810);
not NOT1 (N2566, N2553);
nor NOR3 (N2567, N2559, N558, N2063);
or OR4 (N2568, N2550, N905, N1143, N959);
and AND3 (N2569, N2565, N1668, N1332);
xor XOR2 (N2570, N2562, N1199);
buf BUF1 (N2571, N2569);
or OR4 (N2572, N2566, N37, N1323, N1861);
not NOT1 (N2573, N2514);
nand NAND3 (N2574, N2564, N2449, N25);
not NOT1 (N2575, N2534);
nand NAND3 (N2576, N2572, N725, N397);
and AND4 (N2577, N2571, N2522, N844, N978);
xor XOR2 (N2578, N2577, N2164);
or OR2 (N2579, N2561, N759);
buf BUF1 (N2580, N2574);
buf BUF1 (N2581, N2580);
xor XOR2 (N2582, N2568, N1356);
and AND3 (N2583, N2551, N1295, N2326);
not NOT1 (N2584, N2582);
xor XOR2 (N2585, N2584, N2380);
buf BUF1 (N2586, N2578);
or OR2 (N2587, N2573, N1511);
not NOT1 (N2588, N2587);
or OR4 (N2589, N2579, N2029, N1812, N1872);
nor NOR4 (N2590, N2567, N1049, N1072, N2484);
nand NAND2 (N2591, N2586, N1858);
buf BUF1 (N2592, N2581);
nor NOR3 (N2593, N2583, N2432, N509);
or OR3 (N2594, N2585, N898, N1842);
not NOT1 (N2595, N2590);
and AND2 (N2596, N2575, N1737);
nor NOR4 (N2597, N2588, N1303, N1354, N676);
buf BUF1 (N2598, N2589);
or OR3 (N2599, N2595, N2157, N1666);
not NOT1 (N2600, N2592);
nor NOR4 (N2601, N2576, N1042, N1895, N251);
nor NOR3 (N2602, N2593, N1396, N1598);
nor NOR2 (N2603, N2594, N2110);
nand NAND4 (N2604, N2603, N1550, N1035, N2283);
not NOT1 (N2605, N2604);
not NOT1 (N2606, N2599);
buf BUF1 (N2607, N2596);
not NOT1 (N2608, N2605);
nand NAND3 (N2609, N2608, N1283, N2577);
or OR3 (N2610, N2609, N1971, N330);
not NOT1 (N2611, N2570);
not NOT1 (N2612, N2597);
nand NAND2 (N2613, N2610, N145);
not NOT1 (N2614, N2606);
nor NOR3 (N2615, N2612, N604, N2318);
or OR2 (N2616, N2600, N2449);
and AND4 (N2617, N2601, N286, N1493, N102);
nor NOR4 (N2618, N2607, N941, N246, N947);
xor XOR2 (N2619, N2617, N2459);
xor XOR2 (N2620, N2618, N1727);
not NOT1 (N2621, N2616);
not NOT1 (N2622, N2615);
nand NAND3 (N2623, N2622, N1502, N2287);
not NOT1 (N2624, N2611);
nor NOR2 (N2625, N2624, N522);
nor NOR4 (N2626, N2602, N1827, N825, N511);
and AND3 (N2627, N2625, N2585, N1254);
nor NOR2 (N2628, N2620, N926);
or OR3 (N2629, N2623, N323, N365);
and AND4 (N2630, N2614, N2559, N631, N511);
nand NAND2 (N2631, N2626, N760);
buf BUF1 (N2632, N2619);
or OR3 (N2633, N2629, N431, N1116);
and AND2 (N2634, N2633, N1369);
not NOT1 (N2635, N2598);
buf BUF1 (N2636, N2621);
nand NAND2 (N2637, N2632, N1720);
nor NOR2 (N2638, N2634, N1794);
or OR3 (N2639, N2613, N1111, N1232);
not NOT1 (N2640, N2591);
nor NOR2 (N2641, N2627, N2307);
nor NOR4 (N2642, N2631, N2222, N1607, N1453);
xor XOR2 (N2643, N2642, N2093);
nor NOR2 (N2644, N2636, N2247);
not NOT1 (N2645, N2640);
buf BUF1 (N2646, N2639);
nor NOR4 (N2647, N2646, N1249, N1172, N748);
xor XOR2 (N2648, N2628, N988);
nor NOR3 (N2649, N2644, N686, N1013);
buf BUF1 (N2650, N2645);
xor XOR2 (N2651, N2638, N213);
not NOT1 (N2652, N2635);
xor XOR2 (N2653, N2637, N268);
xor XOR2 (N2654, N2643, N2105);
buf BUF1 (N2655, N2641);
nor NOR2 (N2656, N2648, N2545);
and AND3 (N2657, N2649, N1561, N2447);
buf BUF1 (N2658, N2651);
nor NOR4 (N2659, N2652, N1192, N1322, N1082);
xor XOR2 (N2660, N2659, N1610);
xor XOR2 (N2661, N2647, N2476);
nand NAND3 (N2662, N2660, N318, N912);
and AND3 (N2663, N2653, N2034, N690);
buf BUF1 (N2664, N2663);
nor NOR3 (N2665, N2630, N976, N159);
and AND3 (N2666, N2655, N637, N697);
nor NOR4 (N2667, N2661, N814, N2345, N795);
and AND3 (N2668, N2665, N734, N265);
not NOT1 (N2669, N2666);
buf BUF1 (N2670, N2657);
buf BUF1 (N2671, N2650);
buf BUF1 (N2672, N2667);
not NOT1 (N2673, N2662);
and AND3 (N2674, N2658, N1295, N2409);
xor XOR2 (N2675, N2674, N2572);
nor NOR4 (N2676, N2654, N1574, N1480, N975);
and AND4 (N2677, N2671, N699, N414, N841);
not NOT1 (N2678, N2672);
or OR3 (N2679, N2678, N1436, N1792);
nand NAND3 (N2680, N2673, N359, N2502);
not NOT1 (N2681, N2677);
not NOT1 (N2682, N2669);
nor NOR2 (N2683, N2680, N1498);
xor XOR2 (N2684, N2675, N2063);
not NOT1 (N2685, N2656);
xor XOR2 (N2686, N2664, N831);
xor XOR2 (N2687, N2682, N1206);
or OR2 (N2688, N2681, N660);
nand NAND3 (N2689, N2688, N1022, N531);
or OR3 (N2690, N2686, N1235, N517);
and AND4 (N2691, N2668, N863, N39, N2085);
xor XOR2 (N2692, N2691, N1377);
nor NOR4 (N2693, N2692, N134, N590, N1554);
and AND4 (N2694, N2676, N289, N685, N1067);
xor XOR2 (N2695, N2689, N1566);
xor XOR2 (N2696, N2679, N1585);
or OR4 (N2697, N2693, N1450, N2444, N2177);
xor XOR2 (N2698, N2694, N644);
buf BUF1 (N2699, N2697);
buf BUF1 (N2700, N2685);
xor XOR2 (N2701, N2698, N1140);
or OR2 (N2702, N2687, N1926);
buf BUF1 (N2703, N2702);
or OR3 (N2704, N2684, N174, N1012);
not NOT1 (N2705, N2683);
or OR4 (N2706, N2704, N1477, N2695, N2609);
or OR2 (N2707, N478, N1212);
or OR4 (N2708, N2699, N2182, N409, N1816);
nand NAND2 (N2709, N2707, N244);
nand NAND4 (N2710, N2696, N25, N1688, N266);
xor XOR2 (N2711, N2701, N1839);
and AND3 (N2712, N2705, N572, N485);
not NOT1 (N2713, N2708);
buf BUF1 (N2714, N2706);
or OR3 (N2715, N2713, N1536, N2424);
nor NOR4 (N2716, N2710, N166, N375, N2241);
buf BUF1 (N2717, N2711);
not NOT1 (N2718, N2714);
xor XOR2 (N2719, N2717, N899);
xor XOR2 (N2720, N2690, N936);
or OR2 (N2721, N2718, N387);
and AND2 (N2722, N2670, N1469);
or OR2 (N2723, N2709, N1288);
xor XOR2 (N2724, N2719, N1481);
nor NOR3 (N2725, N2720, N1287, N1235);
or OR3 (N2726, N2725, N2443, N81);
nor NOR4 (N2727, N2712, N191, N1194, N2445);
not NOT1 (N2728, N2715);
nand NAND3 (N2729, N2721, N1296, N2135);
or OR4 (N2730, N2726, N1457, N2478, N2435);
and AND3 (N2731, N2730, N1910, N1569);
and AND2 (N2732, N2731, N1604);
and AND2 (N2733, N2728, N1023);
nand NAND3 (N2734, N2729, N1858, N1863);
xor XOR2 (N2735, N2724, N1595);
xor XOR2 (N2736, N2733, N141);
buf BUF1 (N2737, N2732);
xor XOR2 (N2738, N2716, N2579);
or OR2 (N2739, N2703, N2345);
and AND3 (N2740, N2700, N1852, N2577);
not NOT1 (N2741, N2737);
buf BUF1 (N2742, N2734);
buf BUF1 (N2743, N2727);
buf BUF1 (N2744, N2743);
or OR4 (N2745, N2741, N1523, N431, N865);
not NOT1 (N2746, N2735);
xor XOR2 (N2747, N2739, N659);
xor XOR2 (N2748, N2740, N2532);
nor NOR4 (N2749, N2747, N2438, N1661, N447);
nand NAND3 (N2750, N2723, N588, N44);
xor XOR2 (N2751, N2738, N405);
and AND4 (N2752, N2749, N815, N505, N1645);
xor XOR2 (N2753, N2736, N2377);
xor XOR2 (N2754, N2744, N952);
nor NOR3 (N2755, N2722, N2585, N372);
or OR3 (N2756, N2742, N1949, N1737);
or OR4 (N2757, N2751, N202, N1751, N1349);
nand NAND4 (N2758, N2750, N1163, N1904, N2699);
buf BUF1 (N2759, N2755);
nor NOR4 (N2760, N2753, N1449, N1880, N199);
not NOT1 (N2761, N2746);
nor NOR3 (N2762, N2760, N474, N658);
buf BUF1 (N2763, N2748);
buf BUF1 (N2764, N2758);
nand NAND2 (N2765, N2759, N2333);
buf BUF1 (N2766, N2761);
nor NOR3 (N2767, N2766, N155, N811);
not NOT1 (N2768, N2754);
buf BUF1 (N2769, N2762);
xor XOR2 (N2770, N2757, N1185);
nand NAND2 (N2771, N2768, N1603);
and AND4 (N2772, N2769, N2211, N1581, N2046);
buf BUF1 (N2773, N2765);
nand NAND4 (N2774, N2773, N1871, N832, N2324);
or OR3 (N2775, N2774, N962, N2513);
not NOT1 (N2776, N2764);
nor NOR4 (N2777, N2775, N1120, N283, N359);
and AND2 (N2778, N2770, N1927);
xor XOR2 (N2779, N2772, N874);
and AND2 (N2780, N2777, N530);
or OR2 (N2781, N2780, N340);
nand NAND2 (N2782, N2767, N693);
nand NAND2 (N2783, N2779, N2703);
nor NOR2 (N2784, N2778, N1842);
buf BUF1 (N2785, N2752);
nor NOR2 (N2786, N2784, N2447);
xor XOR2 (N2787, N2782, N502);
and AND2 (N2788, N2785, N1462);
xor XOR2 (N2789, N2783, N2074);
or OR3 (N2790, N2771, N1273, N2529);
xor XOR2 (N2791, N2788, N1908);
nand NAND4 (N2792, N2787, N367, N1389, N275);
buf BUF1 (N2793, N2781);
xor XOR2 (N2794, N2763, N474);
xor XOR2 (N2795, N2790, N797);
nor NOR3 (N2796, N2786, N166, N2567);
or OR3 (N2797, N2791, N2473, N230);
and AND4 (N2798, N2789, N1301, N1298, N314);
nand NAND3 (N2799, N2793, N2120, N1463);
nand NAND2 (N2800, N2797, N630);
nor NOR3 (N2801, N2776, N892, N1790);
and AND3 (N2802, N2796, N1304, N1448);
xor XOR2 (N2803, N2801, N2732);
and AND4 (N2804, N2756, N561, N236, N246);
nand NAND4 (N2805, N2794, N573, N2479, N1082);
and AND3 (N2806, N2803, N1779, N1738);
not NOT1 (N2807, N2804);
not NOT1 (N2808, N2805);
and AND2 (N2809, N2745, N775);
and AND2 (N2810, N2795, N1384);
not NOT1 (N2811, N2802);
and AND2 (N2812, N2809, N1330);
xor XOR2 (N2813, N2811, N500);
xor XOR2 (N2814, N2812, N2626);
or OR3 (N2815, N2798, N291, N2223);
nand NAND2 (N2816, N2810, N1955);
not NOT1 (N2817, N2807);
or OR2 (N2818, N2799, N2242);
buf BUF1 (N2819, N2792);
not NOT1 (N2820, N2806);
and AND2 (N2821, N2800, N2316);
nor NOR2 (N2822, N2816, N1804);
nor NOR4 (N2823, N2813, N2163, N1173, N628);
buf BUF1 (N2824, N2819);
nor NOR2 (N2825, N2817, N873);
nor NOR4 (N2826, N2821, N2446, N631, N76);
nor NOR3 (N2827, N2815, N1219, N1072);
buf BUF1 (N2828, N2818);
not NOT1 (N2829, N2828);
xor XOR2 (N2830, N2820, N2571);
and AND3 (N2831, N2830, N1573, N1945);
or OR2 (N2832, N2824, N2063);
buf BUF1 (N2833, N2827);
buf BUF1 (N2834, N2831);
and AND3 (N2835, N2833, N1733, N2415);
or OR3 (N2836, N2808, N881, N1662);
not NOT1 (N2837, N2834);
xor XOR2 (N2838, N2825, N1495);
and AND4 (N2839, N2814, N2621, N1362, N2101);
or OR2 (N2840, N2837, N2696);
nor NOR2 (N2841, N2835, N15);
not NOT1 (N2842, N2840);
nand NAND2 (N2843, N2842, N1786);
not NOT1 (N2844, N2843);
or OR4 (N2845, N2836, N1604, N2707, N764);
nand NAND3 (N2846, N2832, N2192, N2016);
not NOT1 (N2847, N2844);
buf BUF1 (N2848, N2841);
xor XOR2 (N2849, N2839, N2587);
buf BUF1 (N2850, N2847);
xor XOR2 (N2851, N2848, N133);
xor XOR2 (N2852, N2850, N2246);
buf BUF1 (N2853, N2851);
nor NOR4 (N2854, N2852, N1698, N1062, N1404);
nor NOR2 (N2855, N2838, N1876);
and AND2 (N2856, N2855, N1930);
nand NAND4 (N2857, N2823, N833, N139, N1803);
not NOT1 (N2858, N2853);
not NOT1 (N2859, N2849);
nand NAND4 (N2860, N2856, N1870, N2733, N1065);
buf BUF1 (N2861, N2846);
xor XOR2 (N2862, N2822, N2085);
and AND4 (N2863, N2845, N246, N228, N84);
or OR2 (N2864, N2861, N662);
or OR2 (N2865, N2860, N1037);
nand NAND4 (N2866, N2854, N2253, N755, N119);
nor NOR2 (N2867, N2866, N280);
not NOT1 (N2868, N2857);
or OR3 (N2869, N2868, N1453, N1084);
not NOT1 (N2870, N2862);
xor XOR2 (N2871, N2829, N263);
or OR2 (N2872, N2867, N509);
and AND3 (N2873, N2858, N1578, N2251);
or OR2 (N2874, N2871, N848);
nand NAND4 (N2875, N2874, N1773, N648, N686);
nor NOR2 (N2876, N2869, N1492);
or OR3 (N2877, N2870, N2268, N77);
buf BUF1 (N2878, N2877);
and AND3 (N2879, N2878, N2807, N469);
xor XOR2 (N2880, N2826, N629);
nand NAND4 (N2881, N2872, N2747, N1210, N2488);
xor XOR2 (N2882, N2864, N816);
xor XOR2 (N2883, N2859, N1931);
not NOT1 (N2884, N2875);
xor XOR2 (N2885, N2879, N2780);
nor NOR2 (N2886, N2876, N40);
nand NAND2 (N2887, N2884, N2787);
nor NOR2 (N2888, N2881, N555);
or OR2 (N2889, N2873, N1314);
xor XOR2 (N2890, N2888, N1122);
or OR2 (N2891, N2887, N2551);
and AND3 (N2892, N2880, N2174, N879);
buf BUF1 (N2893, N2885);
nor NOR3 (N2894, N2892, N1693, N1646);
or OR4 (N2895, N2894, N1737, N1107, N1955);
or OR4 (N2896, N2883, N700, N217, N201);
not NOT1 (N2897, N2890);
and AND3 (N2898, N2886, N2728, N1011);
nor NOR3 (N2899, N2895, N2881, N1236);
not NOT1 (N2900, N2896);
nor NOR2 (N2901, N2897, N1028);
and AND3 (N2902, N2900, N411, N1870);
or OR3 (N2903, N2882, N137, N2703);
xor XOR2 (N2904, N2889, N1793);
nor NOR3 (N2905, N2893, N1760, N2470);
nor NOR3 (N2906, N2899, N2203, N2489);
nand NAND4 (N2907, N2901, N300, N1416, N665);
buf BUF1 (N2908, N2904);
nor NOR3 (N2909, N2908, N56, N1430);
xor XOR2 (N2910, N2902, N1613);
nand NAND2 (N2911, N2909, N2369);
nand NAND4 (N2912, N2898, N1033, N1938, N2272);
not NOT1 (N2913, N2891);
nor NOR3 (N2914, N2907, N2505, N1232);
nor NOR4 (N2915, N2914, N289, N1458, N2615);
or OR4 (N2916, N2910, N33, N298, N639);
or OR3 (N2917, N2903, N173, N2346);
nand NAND2 (N2918, N2905, N1599);
and AND3 (N2919, N2917, N1601, N2690);
or OR3 (N2920, N2913, N170, N2672);
xor XOR2 (N2921, N2919, N638);
xor XOR2 (N2922, N2912, N2227);
nor NOR3 (N2923, N2863, N2495, N496);
buf BUF1 (N2924, N2922);
nor NOR2 (N2925, N2911, N1086);
not NOT1 (N2926, N2916);
not NOT1 (N2927, N2906);
nor NOR2 (N2928, N2927, N2085);
buf BUF1 (N2929, N2926);
buf BUF1 (N2930, N2920);
and AND3 (N2931, N2918, N1092, N323);
buf BUF1 (N2932, N2921);
buf BUF1 (N2933, N2932);
xor XOR2 (N2934, N2923, N1588);
or OR2 (N2935, N2933, N1253);
and AND2 (N2936, N2924, N2247);
nand NAND3 (N2937, N2935, N1641, N930);
or OR2 (N2938, N2915, N570);
nand NAND3 (N2939, N2928, N733, N1133);
and AND4 (N2940, N2865, N2504, N2280, N2258);
nand NAND3 (N2941, N2940, N2398, N2769);
and AND4 (N2942, N2941, N224, N215, N1273);
xor XOR2 (N2943, N2930, N1869);
nor NOR3 (N2944, N2936, N1662, N2343);
buf BUF1 (N2945, N2937);
xor XOR2 (N2946, N2938, N434);
not NOT1 (N2947, N2931);
not NOT1 (N2948, N2934);
or OR4 (N2949, N2925, N835, N212, N2356);
nand NAND4 (N2950, N2944, N2593, N122, N1671);
nor NOR3 (N2951, N2942, N371, N1131);
buf BUF1 (N2952, N2950);
and AND2 (N2953, N2939, N466);
buf BUF1 (N2954, N2945);
or OR2 (N2955, N2946, N1019);
nand NAND3 (N2956, N2943, N856, N1571);
buf BUF1 (N2957, N2947);
nor NOR4 (N2958, N2952, N1432, N1137, N10);
not NOT1 (N2959, N2948);
nor NOR2 (N2960, N2957, N1715);
not NOT1 (N2961, N2951);
not NOT1 (N2962, N2929);
not NOT1 (N2963, N2962);
nand NAND4 (N2964, N2959, N342, N2411, N47);
nand NAND2 (N2965, N2955, N687);
xor XOR2 (N2966, N2964, N1270);
not NOT1 (N2967, N2954);
or OR4 (N2968, N2963, N1570, N195, N2787);
nand NAND3 (N2969, N2958, N801, N73);
not NOT1 (N2970, N2965);
and AND4 (N2971, N2960, N1758, N1177, N495);
and AND4 (N2972, N2953, N837, N960, N1936);
nand NAND3 (N2973, N2967, N1731, N2113);
xor XOR2 (N2974, N2973, N2805);
buf BUF1 (N2975, N2970);
buf BUF1 (N2976, N2974);
and AND2 (N2977, N2956, N565);
nor NOR4 (N2978, N2976, N565, N562, N1146);
not NOT1 (N2979, N2968);
buf BUF1 (N2980, N2971);
or OR2 (N2981, N2978, N2568);
nand NAND4 (N2982, N2972, N2962, N2824, N339);
xor XOR2 (N2983, N2979, N1155);
xor XOR2 (N2984, N2980, N334);
not NOT1 (N2985, N2983);
not NOT1 (N2986, N2961);
buf BUF1 (N2987, N2975);
nor NOR2 (N2988, N2987, N743);
not NOT1 (N2989, N2982);
nor NOR2 (N2990, N2949, N2324);
nor NOR2 (N2991, N2986, N455);
and AND3 (N2992, N2985, N441, N157);
and AND3 (N2993, N2966, N569, N474);
xor XOR2 (N2994, N2988, N589);
and AND2 (N2995, N2989, N880);
xor XOR2 (N2996, N2969, N2536);
nand NAND4 (N2997, N2977, N1330, N2357, N2701);
buf BUF1 (N2998, N2997);
buf BUF1 (N2999, N2993);
nand NAND4 (N3000, N2998, N1108, N904, N2775);
nor NOR3 (N3001, N2999, N420, N1539);
nand NAND2 (N3002, N2990, N270);
buf BUF1 (N3003, N3002);
buf BUF1 (N3004, N2996);
not NOT1 (N3005, N2992);
nand NAND4 (N3006, N3000, N609, N1956, N2033);
xor XOR2 (N3007, N3005, N1936);
xor XOR2 (N3008, N2981, N2321);
nor NOR3 (N3009, N2984, N796, N2565);
nand NAND3 (N3010, N3008, N1445, N101);
nor NOR3 (N3011, N3004, N519, N2724);
or OR2 (N3012, N3009, N1115);
nor NOR3 (N3013, N3003, N2108, N1720);
buf BUF1 (N3014, N3013);
and AND2 (N3015, N3011, N1108);
nor NOR2 (N3016, N3014, N1767);
nor NOR3 (N3017, N3010, N1158, N1341);
nand NAND3 (N3018, N3012, N1873, N2482);
xor XOR2 (N3019, N2995, N2309);
or OR2 (N3020, N2994, N2763);
and AND4 (N3021, N3016, N2248, N2443, N2750);
buf BUF1 (N3022, N3017);
buf BUF1 (N3023, N3001);
and AND3 (N3024, N3019, N1744, N2902);
xor XOR2 (N3025, N3020, N230);
and AND4 (N3026, N3018, N2345, N1762, N815);
and AND4 (N3027, N3024, N1924, N754, N1664);
and AND2 (N3028, N3025, N868);
xor XOR2 (N3029, N3028, N670);
or OR2 (N3030, N3021, N560);
xor XOR2 (N3031, N3027, N852);
and AND4 (N3032, N3023, N1784, N2189, N5);
buf BUF1 (N3033, N3006);
not NOT1 (N3034, N3007);
not NOT1 (N3035, N3030);
not NOT1 (N3036, N3015);
nand NAND2 (N3037, N3026, N1878);
or OR4 (N3038, N3032, N2670, N2171, N1883);
xor XOR2 (N3039, N2991, N2378);
buf BUF1 (N3040, N3039);
nand NAND4 (N3041, N3031, N1979, N1546, N2282);
and AND2 (N3042, N3022, N1182);
nand NAND4 (N3043, N3035, N747, N2618, N2895);
or OR4 (N3044, N3038, N913, N1853, N1396);
nor NOR4 (N3045, N3034, N2179, N1704, N1948);
or OR3 (N3046, N3033, N1243, N1550);
nor NOR2 (N3047, N3029, N532);
not NOT1 (N3048, N3045);
not NOT1 (N3049, N3041);
xor XOR2 (N3050, N3042, N1955);
or OR2 (N3051, N3046, N2433);
nand NAND3 (N3052, N3048, N501, N1637);
xor XOR2 (N3053, N3037, N1691);
xor XOR2 (N3054, N3036, N1428);
xor XOR2 (N3055, N3053, N970);
xor XOR2 (N3056, N3054, N2996);
xor XOR2 (N3057, N3056, N1833);
buf BUF1 (N3058, N3050);
xor XOR2 (N3059, N3055, N2576);
nand NAND2 (N3060, N3058, N1254);
nor NOR4 (N3061, N3044, N542, N2628, N2887);
or OR4 (N3062, N3052, N1223, N2199, N2796);
nand NAND2 (N3063, N3043, N1845);
nor NOR4 (N3064, N3060, N1446, N1619, N2658);
not NOT1 (N3065, N3061);
not NOT1 (N3066, N3049);
nor NOR3 (N3067, N3047, N1187, N822);
and AND4 (N3068, N3057, N91, N850, N1449);
xor XOR2 (N3069, N3068, N2858);
buf BUF1 (N3070, N3067);
nand NAND3 (N3071, N3064, N596, N1920);
not NOT1 (N3072, N3066);
nand NAND2 (N3073, N3051, N1038);
not NOT1 (N3074, N3040);
nor NOR4 (N3075, N3062, N2534, N2412, N1170);
nand NAND4 (N3076, N3070, N705, N3071, N1948);
not NOT1 (N3077, N268);
buf BUF1 (N3078, N3065);
xor XOR2 (N3079, N3078, N740);
not NOT1 (N3080, N3077);
buf BUF1 (N3081, N3073);
xor XOR2 (N3082, N3081, N1032);
not NOT1 (N3083, N3079);
xor XOR2 (N3084, N3083, N1558);
not NOT1 (N3085, N3072);
and AND3 (N3086, N3085, N2529, N1144);
or OR2 (N3087, N3076, N1410);
buf BUF1 (N3088, N3059);
and AND4 (N3089, N3087, N1633, N882, N386);
not NOT1 (N3090, N3089);
or OR2 (N3091, N3088, N733);
nor NOR4 (N3092, N3074, N1397, N2402, N65);
or OR3 (N3093, N3075, N556, N2413);
buf BUF1 (N3094, N3063);
or OR4 (N3095, N3092, N1118, N1174, N2607);
nand NAND2 (N3096, N3093, N1782);
or OR4 (N3097, N3091, N1125, N2408, N316);
and AND4 (N3098, N3094, N522, N1241, N2311);
not NOT1 (N3099, N3086);
buf BUF1 (N3100, N3098);
or OR4 (N3101, N3080, N828, N1312, N2379);
xor XOR2 (N3102, N3099, N2718);
buf BUF1 (N3103, N3096);
nand NAND4 (N3104, N3097, N3075, N1621, N1285);
and AND3 (N3105, N3084, N2123, N2209);
xor XOR2 (N3106, N3069, N2064);
buf BUF1 (N3107, N3104);
and AND2 (N3108, N3100, N762);
nand NAND2 (N3109, N3101, N2355);
nand NAND2 (N3110, N3095, N311);
nand NAND2 (N3111, N3108, N988);
buf BUF1 (N3112, N3105);
buf BUF1 (N3113, N3106);
buf BUF1 (N3114, N3102);
xor XOR2 (N3115, N3103, N1034);
and AND2 (N3116, N3110, N2567);
nor NOR3 (N3117, N3113, N797, N924);
and AND3 (N3118, N3111, N1048, N350);
not NOT1 (N3119, N3107);
xor XOR2 (N3120, N3112, N692);
not NOT1 (N3121, N3116);
not NOT1 (N3122, N3121);
nand NAND2 (N3123, N3119, N916);
nor NOR3 (N3124, N3114, N694, N1006);
or OR4 (N3125, N3090, N2980, N1840, N2074);
xor XOR2 (N3126, N3117, N2756);
nor NOR3 (N3127, N3123, N1647, N583);
nand NAND4 (N3128, N3122, N1332, N2361, N274);
not NOT1 (N3129, N3115);
xor XOR2 (N3130, N3109, N113);
nand NAND2 (N3131, N3126, N2323);
and AND2 (N3132, N3118, N2472);
not NOT1 (N3133, N3082);
not NOT1 (N3134, N3125);
buf BUF1 (N3135, N3133);
or OR3 (N3136, N3132, N2986, N2059);
not NOT1 (N3137, N3135);
or OR3 (N3138, N3137, N2282, N2938);
nor NOR2 (N3139, N3134, N567);
buf BUF1 (N3140, N3124);
xor XOR2 (N3141, N3138, N1235);
xor XOR2 (N3142, N3129, N595);
or OR3 (N3143, N3127, N814, N1038);
or OR3 (N3144, N3130, N733, N2777);
and AND4 (N3145, N3142, N3059, N2581, N673);
nand NAND2 (N3146, N3141, N2900);
nand NAND4 (N3147, N3140, N1425, N2182, N280);
xor XOR2 (N3148, N3145, N885);
not NOT1 (N3149, N3139);
and AND3 (N3150, N3120, N123, N1900);
or OR3 (N3151, N3136, N2575, N1224);
or OR4 (N3152, N3128, N46, N2825, N39);
xor XOR2 (N3153, N3151, N3025);
xor XOR2 (N3154, N3143, N706);
or OR2 (N3155, N3154, N2213);
xor XOR2 (N3156, N3153, N176);
not NOT1 (N3157, N3155);
not NOT1 (N3158, N3156);
or OR4 (N3159, N3149, N2045, N250, N1751);
not NOT1 (N3160, N3152);
nand NAND2 (N3161, N3131, N242);
or OR2 (N3162, N3150, N545);
and AND2 (N3163, N3146, N217);
nand NAND3 (N3164, N3159, N1791, N451);
and AND3 (N3165, N3160, N1045, N2100);
and AND3 (N3166, N3162, N748, N2002);
and AND2 (N3167, N3144, N547);
or OR2 (N3168, N3158, N1522);
xor XOR2 (N3169, N3161, N1749);
or OR2 (N3170, N3169, N2942);
or OR4 (N3171, N3163, N1510, N2787, N2044);
buf BUF1 (N3172, N3170);
not NOT1 (N3173, N3148);
and AND3 (N3174, N3165, N2129, N2803);
and AND2 (N3175, N3157, N343);
and AND3 (N3176, N3172, N2181, N1771);
xor XOR2 (N3177, N3167, N2760);
not NOT1 (N3178, N3147);
and AND2 (N3179, N3177, N749);
nor NOR4 (N3180, N3174, N681, N17, N2221);
nand NAND2 (N3181, N3176, N120);
nand NAND2 (N3182, N3178, N3104);
nor NOR3 (N3183, N3173, N1550, N1940);
or OR3 (N3184, N3175, N2683, N2488);
xor XOR2 (N3185, N3164, N2193);
buf BUF1 (N3186, N3184);
buf BUF1 (N3187, N3181);
nor NOR2 (N3188, N3166, N2348);
xor XOR2 (N3189, N3183, N2063);
xor XOR2 (N3190, N3179, N2077);
not NOT1 (N3191, N3189);
or OR3 (N3192, N3171, N435, N2607);
not NOT1 (N3193, N3190);
nand NAND4 (N3194, N3185, N685, N1965, N67);
buf BUF1 (N3195, N3192);
and AND3 (N3196, N3195, N2257, N1754);
xor XOR2 (N3197, N3182, N2454);
and AND4 (N3198, N3168, N1521, N982, N136);
or OR2 (N3199, N3187, N246);
or OR2 (N3200, N3186, N584);
or OR4 (N3201, N3180, N1821, N1268, N1234);
nor NOR2 (N3202, N3198, N3086);
nor NOR4 (N3203, N3202, N767, N3064, N529);
xor XOR2 (N3204, N3196, N2726);
xor XOR2 (N3205, N3191, N384);
buf BUF1 (N3206, N3205);
not NOT1 (N3207, N3194);
nor NOR4 (N3208, N3193, N1846, N1287, N941);
xor XOR2 (N3209, N3200, N3176);
or OR4 (N3210, N3199, N1093, N1883, N2526);
nor NOR3 (N3211, N3204, N860, N199);
and AND2 (N3212, N3208, N1928);
xor XOR2 (N3213, N3210, N3206);
xor XOR2 (N3214, N1881, N1390);
xor XOR2 (N3215, N3214, N1874);
nor NOR2 (N3216, N3197, N935);
or OR2 (N3217, N3209, N2769);
nand NAND3 (N3218, N3213, N1897, N2235);
buf BUF1 (N3219, N3188);
not NOT1 (N3220, N3207);
nor NOR2 (N3221, N3211, N1302);
nand NAND2 (N3222, N3218, N1463);
not NOT1 (N3223, N3215);
buf BUF1 (N3224, N3221);
nand NAND4 (N3225, N3219, N1767, N2309, N758);
xor XOR2 (N3226, N3220, N1574);
buf BUF1 (N3227, N3223);
and AND3 (N3228, N3216, N101, N308);
and AND3 (N3229, N3226, N2167, N281);
nand NAND2 (N3230, N3201, N2338);
and AND4 (N3231, N3230, N2879, N1205, N1085);
nor NOR2 (N3232, N3212, N1193);
nand NAND3 (N3233, N3229, N403, N1923);
buf BUF1 (N3234, N3222);
nand NAND4 (N3235, N3227, N331, N1972, N758);
not NOT1 (N3236, N3217);
or OR4 (N3237, N3203, N328, N2812, N3045);
buf BUF1 (N3238, N3233);
or OR2 (N3239, N3232, N1201);
buf BUF1 (N3240, N3237);
xor XOR2 (N3241, N3228, N1812);
nand NAND3 (N3242, N3234, N629, N2024);
buf BUF1 (N3243, N3238);
nand NAND4 (N3244, N3225, N2266, N1113, N1587);
nor NOR2 (N3245, N3231, N1360);
and AND4 (N3246, N3244, N2469, N3231, N1138);
not NOT1 (N3247, N3242);
nand NAND3 (N3248, N3235, N1763, N2505);
buf BUF1 (N3249, N3240);
nand NAND3 (N3250, N3239, N1835, N71);
not NOT1 (N3251, N3243);
xor XOR2 (N3252, N3224, N2281);
nand NAND3 (N3253, N3252, N683, N1100);
not NOT1 (N3254, N3236);
or OR2 (N3255, N3249, N1319);
xor XOR2 (N3256, N3245, N1963);
nor NOR4 (N3257, N3256, N2717, N3160, N2996);
nor NOR2 (N3258, N3247, N2460);
xor XOR2 (N3259, N3255, N1327);
xor XOR2 (N3260, N3259, N1911);
and AND2 (N3261, N3253, N1522);
nand NAND4 (N3262, N3257, N169, N667, N3104);
xor XOR2 (N3263, N3262, N1979);
xor XOR2 (N3264, N3248, N626);
nor NOR4 (N3265, N3251, N533, N1044, N1140);
buf BUF1 (N3266, N3241);
nand NAND3 (N3267, N3260, N3014, N2658);
nor NOR2 (N3268, N3263, N1297);
or OR2 (N3269, N3267, N2457);
buf BUF1 (N3270, N3246);
buf BUF1 (N3271, N3265);
or OR4 (N3272, N3269, N1935, N3055, N439);
nand NAND2 (N3273, N3270, N593);
nand NAND3 (N3274, N3261, N1819, N137);
nor NOR2 (N3275, N3264, N591);
or OR4 (N3276, N3254, N3013, N3025, N287);
xor XOR2 (N3277, N3266, N2659);
nor NOR4 (N3278, N3276, N1159, N2224, N2950);
not NOT1 (N3279, N3277);
not NOT1 (N3280, N3250);
not NOT1 (N3281, N3274);
nand NAND3 (N3282, N3275, N390, N1404);
xor XOR2 (N3283, N3258, N2886);
xor XOR2 (N3284, N3283, N1448);
buf BUF1 (N3285, N3280);
or OR2 (N3286, N3273, N4);
and AND2 (N3287, N3284, N2313);
and AND4 (N3288, N3285, N219, N241, N3046);
xor XOR2 (N3289, N3281, N2969);
nand NAND3 (N3290, N3282, N2757, N3083);
nor NOR4 (N3291, N3272, N468, N3213, N38);
xor XOR2 (N3292, N3290, N3285);
or OR4 (N3293, N3268, N999, N1600, N310);
buf BUF1 (N3294, N3289);
or OR2 (N3295, N3287, N2340);
buf BUF1 (N3296, N3286);
buf BUF1 (N3297, N3291);
or OR3 (N3298, N3278, N2039, N1880);
and AND4 (N3299, N3297, N3151, N1906, N443);
nor NOR2 (N3300, N3288, N217);
or OR4 (N3301, N3293, N2003, N65, N3245);
not NOT1 (N3302, N3296);
and AND2 (N3303, N3292, N3103);
nor NOR4 (N3304, N3298, N3166, N569, N1802);
not NOT1 (N3305, N3304);
not NOT1 (N3306, N3294);
not NOT1 (N3307, N3305);
not NOT1 (N3308, N3301);
nand NAND3 (N3309, N3307, N1117, N3187);
not NOT1 (N3310, N3302);
nor NOR3 (N3311, N3279, N3241, N616);
and AND2 (N3312, N3299, N1583);
nor NOR3 (N3313, N3308, N1187, N2092);
nand NAND2 (N3314, N3310, N1303);
buf BUF1 (N3315, N3312);
not NOT1 (N3316, N3295);
buf BUF1 (N3317, N3306);
nand NAND3 (N3318, N3311, N1446, N1040);
buf BUF1 (N3319, N3314);
and AND4 (N3320, N3315, N3173, N1949, N3132);
not NOT1 (N3321, N3319);
buf BUF1 (N3322, N3313);
buf BUF1 (N3323, N3320);
buf BUF1 (N3324, N3303);
nor NOR3 (N3325, N3316, N1406, N3057);
not NOT1 (N3326, N3317);
buf BUF1 (N3327, N3318);
or OR4 (N3328, N3326, N1501, N3032, N3109);
nor NOR4 (N3329, N3324, N2411, N447, N254);
nand NAND4 (N3330, N3271, N1233, N1862, N2382);
nand NAND4 (N3331, N3309, N1020, N3093, N1071);
and AND4 (N3332, N3322, N1398, N3147, N2600);
nand NAND2 (N3333, N3332, N1871);
nand NAND3 (N3334, N3327, N2017, N827);
not NOT1 (N3335, N3300);
and AND4 (N3336, N3335, N3252, N1627, N2567);
xor XOR2 (N3337, N3336, N1216);
not NOT1 (N3338, N3330);
and AND3 (N3339, N3333, N1300, N1085);
nand NAND3 (N3340, N3337, N18, N1774);
not NOT1 (N3341, N3329);
or OR2 (N3342, N3340, N1546);
nor NOR3 (N3343, N3334, N76, N3153);
nand NAND4 (N3344, N3343, N3258, N1721, N125);
or OR4 (N3345, N3342, N2851, N40, N733);
nand NAND2 (N3346, N3321, N1915);
nand NAND3 (N3347, N3331, N2944, N1514);
or OR2 (N3348, N3325, N2492);
buf BUF1 (N3349, N3346);
nand NAND3 (N3350, N3349, N3131, N857);
nand NAND2 (N3351, N3339, N2134);
not NOT1 (N3352, N3344);
xor XOR2 (N3353, N3350, N610);
xor XOR2 (N3354, N3353, N2172);
xor XOR2 (N3355, N3354, N1733);
not NOT1 (N3356, N3351);
buf BUF1 (N3357, N3355);
xor XOR2 (N3358, N3338, N114);
xor XOR2 (N3359, N3341, N2647);
not NOT1 (N3360, N3352);
not NOT1 (N3361, N3328);
xor XOR2 (N3362, N3356, N3257);
xor XOR2 (N3363, N3361, N2289);
nand NAND2 (N3364, N3359, N1737);
buf BUF1 (N3365, N3358);
and AND4 (N3366, N3365, N2773, N1475, N2070);
nand NAND4 (N3367, N3345, N3230, N1925, N2503);
buf BUF1 (N3368, N3366);
nor NOR3 (N3369, N3357, N3178, N310);
not NOT1 (N3370, N3360);
not NOT1 (N3371, N3367);
or OR3 (N3372, N3323, N3015, N3356);
nor NOR2 (N3373, N3369, N3342);
not NOT1 (N3374, N3372);
or OR2 (N3375, N3368, N2515);
not NOT1 (N3376, N3362);
or OR3 (N3377, N3363, N3010, N748);
nand NAND4 (N3378, N3377, N2970, N3099, N2746);
not NOT1 (N3379, N3348);
xor XOR2 (N3380, N3375, N1996);
or OR4 (N3381, N3364, N2165, N602, N1015);
buf BUF1 (N3382, N3374);
not NOT1 (N3383, N3381);
nand NAND2 (N3384, N3347, N3110);
or OR3 (N3385, N3382, N3, N1805);
xor XOR2 (N3386, N3371, N2296);
not NOT1 (N3387, N3379);
nand NAND2 (N3388, N3384, N30);
and AND2 (N3389, N3373, N1678);
buf BUF1 (N3390, N3386);
xor XOR2 (N3391, N3385, N2838);
or OR3 (N3392, N3378, N443, N662);
and AND4 (N3393, N3388, N2099, N2330, N950);
nor NOR2 (N3394, N3387, N324);
xor XOR2 (N3395, N3383, N2633);
or OR2 (N3396, N3370, N525);
and AND3 (N3397, N3393, N2112, N87);
buf BUF1 (N3398, N3392);
nand NAND2 (N3399, N3391, N621);
or OR2 (N3400, N3397, N1393);
and AND4 (N3401, N3400, N88, N943, N1028);
xor XOR2 (N3402, N3376, N3241);
and AND2 (N3403, N3389, N1246);
xor XOR2 (N3404, N3394, N609);
or OR2 (N3405, N3380, N3255);
xor XOR2 (N3406, N3390, N2182);
nor NOR2 (N3407, N3395, N2374);
nor NOR4 (N3408, N3405, N1759, N409, N2496);
and AND3 (N3409, N3399, N2345, N1658);
nor NOR4 (N3410, N3403, N2735, N3242, N2286);
nand NAND3 (N3411, N3408, N22, N1213);
or OR3 (N3412, N3401, N1641, N1704);
or OR3 (N3413, N3407, N3083, N3336);
nand NAND2 (N3414, N3410, N1741);
or OR3 (N3415, N3409, N2911, N3100);
nor NOR2 (N3416, N3398, N2141);
nand NAND3 (N3417, N3414, N2268, N98);
or OR3 (N3418, N3396, N23, N1891);
nor NOR3 (N3419, N3418, N879, N2508);
or OR4 (N3420, N3419, N440, N2512, N294);
nor NOR3 (N3421, N3406, N491, N792);
nand NAND3 (N3422, N3404, N3357, N627);
or OR4 (N3423, N3402, N2436, N2539, N2698);
nand NAND3 (N3424, N3422, N1009, N966);
xor XOR2 (N3425, N3417, N1383);
not NOT1 (N3426, N3420);
and AND4 (N3427, N3421, N698, N1328, N508);
and AND2 (N3428, N3425, N477);
nand NAND3 (N3429, N3424, N2413, N2381);
xor XOR2 (N3430, N3415, N2903);
nor NOR2 (N3431, N3416, N446);
nor NOR2 (N3432, N3431, N2883);
xor XOR2 (N3433, N3426, N745);
not NOT1 (N3434, N3413);
buf BUF1 (N3435, N3434);
not NOT1 (N3436, N3435);
nor NOR4 (N3437, N3429, N2628, N2607, N1159);
or OR3 (N3438, N3423, N2940, N2415);
nor NOR4 (N3439, N3430, N1787, N2072, N1403);
or OR3 (N3440, N3427, N1020, N586);
and AND4 (N3441, N3411, N2381, N1926, N1129);
nand NAND2 (N3442, N3438, N3215);
nand NAND4 (N3443, N3432, N3211, N2472, N2114);
xor XOR2 (N3444, N3436, N176);
not NOT1 (N3445, N3442);
or OR2 (N3446, N3445, N3198);
and AND2 (N3447, N3439, N3294);
buf BUF1 (N3448, N3447);
or OR4 (N3449, N3448, N584, N2348, N2414);
nand NAND2 (N3450, N3449, N1276);
xor XOR2 (N3451, N3446, N2183);
xor XOR2 (N3452, N3437, N2856);
buf BUF1 (N3453, N3450);
not NOT1 (N3454, N3444);
buf BUF1 (N3455, N3428);
buf BUF1 (N3456, N3441);
nand NAND2 (N3457, N3451, N514);
buf BUF1 (N3458, N3457);
nand NAND3 (N3459, N3456, N2185, N1293);
buf BUF1 (N3460, N3443);
and AND2 (N3461, N3459, N2828);
not NOT1 (N3462, N3454);
not NOT1 (N3463, N3455);
not NOT1 (N3464, N3461);
and AND2 (N3465, N3453, N558);
not NOT1 (N3466, N3465);
and AND3 (N3467, N3466, N2638, N1892);
nor NOR3 (N3468, N3460, N924, N3250);
nand NAND4 (N3469, N3452, N831, N2675, N672);
or OR4 (N3470, N3433, N1490, N3022, N3285);
buf BUF1 (N3471, N3458);
xor XOR2 (N3472, N3440, N1841);
buf BUF1 (N3473, N3463);
or OR4 (N3474, N3412, N356, N363, N3465);
and AND2 (N3475, N3468, N1996);
xor XOR2 (N3476, N3471, N307);
or OR3 (N3477, N3467, N3136, N2774);
not NOT1 (N3478, N3472);
xor XOR2 (N3479, N3473, N3007);
nor NOR3 (N3480, N3469, N770, N1123);
or OR2 (N3481, N3464, N2127);
not NOT1 (N3482, N3478);
or OR2 (N3483, N3476, N1392);
or OR3 (N3484, N3477, N2984, N1609);
not NOT1 (N3485, N3482);
nor NOR4 (N3486, N3484, N178, N2508, N870);
buf BUF1 (N3487, N3486);
nor NOR3 (N3488, N3470, N3312, N462);
and AND3 (N3489, N3474, N3053, N2617);
xor XOR2 (N3490, N3480, N2821);
or OR2 (N3491, N3489, N2963);
xor XOR2 (N3492, N3490, N942);
nand NAND2 (N3493, N3481, N847);
buf BUF1 (N3494, N3492);
nand NAND2 (N3495, N3475, N120);
and AND2 (N3496, N3488, N2896);
nor NOR4 (N3497, N3494, N1485, N1600, N3054);
buf BUF1 (N3498, N3497);
xor XOR2 (N3499, N3485, N2197);
buf BUF1 (N3500, N3487);
xor XOR2 (N3501, N3491, N861);
buf BUF1 (N3502, N3500);
nor NOR2 (N3503, N3495, N747);
nand NAND3 (N3504, N3483, N3336, N343);
nor NOR4 (N3505, N3499, N2285, N2868, N3365);
nand NAND3 (N3506, N3504, N124, N310);
not NOT1 (N3507, N3493);
and AND2 (N3508, N3462, N920);
buf BUF1 (N3509, N3505);
nand NAND3 (N3510, N3479, N443, N300);
nand NAND3 (N3511, N3510, N2325, N645);
not NOT1 (N3512, N3501);
and AND3 (N3513, N3496, N354, N1137);
or OR2 (N3514, N3511, N313);
buf BUF1 (N3515, N3509);
buf BUF1 (N3516, N3498);
nor NOR2 (N3517, N3508, N3303);
and AND2 (N3518, N3513, N2734);
xor XOR2 (N3519, N3518, N431);
and AND2 (N3520, N3519, N1423);
xor XOR2 (N3521, N3503, N1742);
nand NAND2 (N3522, N3502, N501);
buf BUF1 (N3523, N3516);
and AND3 (N3524, N3517, N2214, N24);
not NOT1 (N3525, N3524);
buf BUF1 (N3526, N3507);
or OR4 (N3527, N3525, N217, N2748, N3244);
buf BUF1 (N3528, N3512);
buf BUF1 (N3529, N3528);
or OR4 (N3530, N3522, N3383, N742, N3163);
or OR3 (N3531, N3526, N2046, N1219);
and AND3 (N3532, N3527, N194, N106);
xor XOR2 (N3533, N3523, N428);
nand NAND3 (N3534, N3520, N2742, N2730);
not NOT1 (N3535, N3534);
buf BUF1 (N3536, N3535);
or OR4 (N3537, N3536, N972, N3345, N215);
or OR2 (N3538, N3506, N761);
nor NOR3 (N3539, N3532, N1780, N2924);
nand NAND2 (N3540, N3538, N2177);
not NOT1 (N3541, N3540);
not NOT1 (N3542, N3530);
and AND4 (N3543, N3539, N3113, N20, N1160);
not NOT1 (N3544, N3542);
nor NOR3 (N3545, N3515, N379, N240);
or OR4 (N3546, N3533, N1814, N1106, N1910);
buf BUF1 (N3547, N3537);
xor XOR2 (N3548, N3544, N1904);
xor XOR2 (N3549, N3531, N2569);
or OR3 (N3550, N3548, N477, N2490);
or OR2 (N3551, N3545, N2165);
buf BUF1 (N3552, N3546);
nor NOR2 (N3553, N3529, N1090);
or OR2 (N3554, N3551, N1889);
nor NOR3 (N3555, N3554, N319, N1597);
nand NAND3 (N3556, N3555, N1558, N662);
nand NAND3 (N3557, N3552, N3055, N512);
nor NOR3 (N3558, N3556, N398, N2129);
buf BUF1 (N3559, N3549);
not NOT1 (N3560, N3550);
xor XOR2 (N3561, N3521, N3003);
buf BUF1 (N3562, N3547);
or OR2 (N3563, N3558, N1938);
nor NOR2 (N3564, N3514, N836);
or OR2 (N3565, N3564, N1611);
or OR3 (N3566, N3541, N1511, N632);
nand NAND3 (N3567, N3560, N1463, N1052);
not NOT1 (N3568, N3543);
xor XOR2 (N3569, N3557, N3238);
nor NOR2 (N3570, N3568, N187);
nor NOR4 (N3571, N3563, N1149, N291, N3488);
nand NAND3 (N3572, N3562, N3016, N2480);
not NOT1 (N3573, N3572);
and AND3 (N3574, N3559, N889, N774);
or OR2 (N3575, N3566, N1045);
and AND2 (N3576, N3570, N2400);
and AND2 (N3577, N3574, N2939);
not NOT1 (N3578, N3573);
buf BUF1 (N3579, N3553);
xor XOR2 (N3580, N3575, N2455);
nor NOR2 (N3581, N3561, N2730);
not NOT1 (N3582, N3581);
nor NOR3 (N3583, N3578, N1643, N3501);
nand NAND4 (N3584, N3567, N1349, N1369, N1714);
or OR2 (N3585, N3583, N230);
xor XOR2 (N3586, N3579, N2753);
nor NOR4 (N3587, N3586, N3480, N1332, N3337);
nand NAND2 (N3588, N3584, N3276);
nor NOR4 (N3589, N3587, N1665, N1836, N2566);
and AND4 (N3590, N3588, N2636, N1580, N3522);
not NOT1 (N3591, N3585);
not NOT1 (N3592, N3576);
nor NOR3 (N3593, N3589, N1267, N2864);
nand NAND2 (N3594, N3580, N1533);
not NOT1 (N3595, N3592);
and AND4 (N3596, N3594, N1574, N3251, N465);
xor XOR2 (N3597, N3593, N1518);
nand NAND3 (N3598, N3596, N1992, N800);
or OR3 (N3599, N3571, N796, N2050);
and AND2 (N3600, N3599, N1827);
and AND2 (N3601, N3600, N833);
and AND3 (N3602, N3598, N3451, N2677);
xor XOR2 (N3603, N3601, N1771);
or OR2 (N3604, N3595, N1117);
xor XOR2 (N3605, N3565, N3088);
nor NOR4 (N3606, N3604, N2160, N1507, N865);
not NOT1 (N3607, N3569);
and AND2 (N3608, N3590, N1349);
nand NAND3 (N3609, N3591, N2403, N3160);
buf BUF1 (N3610, N3606);
or OR2 (N3611, N3608, N2201);
or OR4 (N3612, N3610, N490, N23, N583);
not NOT1 (N3613, N3609);
buf BUF1 (N3614, N3602);
not NOT1 (N3615, N3607);
buf BUF1 (N3616, N3605);
not NOT1 (N3617, N3597);
xor XOR2 (N3618, N3613, N3060);
nor NOR4 (N3619, N3611, N1241, N705, N1397);
nand NAND4 (N3620, N3619, N2350, N3582, N574);
or OR3 (N3621, N389, N2002, N1215);
or OR3 (N3622, N3614, N2512, N1182);
not NOT1 (N3623, N3621);
and AND2 (N3624, N3623, N249);
not NOT1 (N3625, N3622);
and AND2 (N3626, N3603, N2156);
buf BUF1 (N3627, N3612);
or OR4 (N3628, N3618, N10, N3031, N498);
not NOT1 (N3629, N3617);
xor XOR2 (N3630, N3624, N3297);
nand NAND4 (N3631, N3630, N1500, N3520, N1410);
or OR2 (N3632, N3628, N3488);
nand NAND3 (N3633, N3615, N3400, N3171);
and AND2 (N3634, N3629, N383);
or OR4 (N3635, N3633, N3559, N299, N610);
not NOT1 (N3636, N3635);
not NOT1 (N3637, N3620);
buf BUF1 (N3638, N3626);
nor NOR2 (N3639, N3631, N1155);
nand NAND2 (N3640, N3639, N1897);
or OR4 (N3641, N3636, N1652, N1999, N2563);
nand NAND3 (N3642, N3638, N1164, N2329);
buf BUF1 (N3643, N3625);
xor XOR2 (N3644, N3640, N26);
buf BUF1 (N3645, N3616);
buf BUF1 (N3646, N3644);
xor XOR2 (N3647, N3646, N395);
nand NAND3 (N3648, N3643, N2188, N455);
buf BUF1 (N3649, N3627);
and AND3 (N3650, N3634, N1221, N1552);
nand NAND2 (N3651, N3577, N1641);
nor NOR3 (N3652, N3641, N1625, N1232);
nand NAND2 (N3653, N3652, N2745);
nor NOR3 (N3654, N3637, N1755, N2000);
nand NAND3 (N3655, N3642, N738, N946);
and AND3 (N3656, N3651, N3480, N2566);
nand NAND4 (N3657, N3656, N3627, N243, N1874);
buf BUF1 (N3658, N3655);
nor NOR2 (N3659, N3658, N3525);
xor XOR2 (N3660, N3632, N2145);
not NOT1 (N3661, N3650);
nand NAND3 (N3662, N3648, N1323, N1345);
xor XOR2 (N3663, N3659, N1125);
xor XOR2 (N3664, N3661, N2114);
nand NAND2 (N3665, N3654, N466);
buf BUF1 (N3666, N3647);
nor NOR4 (N3667, N3662, N178, N2899, N83);
nand NAND2 (N3668, N3645, N2990);
nand NAND4 (N3669, N3660, N1063, N1631, N586);
nor NOR2 (N3670, N3667, N3240);
buf BUF1 (N3671, N3663);
not NOT1 (N3672, N3666);
not NOT1 (N3673, N3668);
and AND2 (N3674, N3653, N1795);
nand NAND4 (N3675, N3670, N318, N2062, N817);
and AND2 (N3676, N3669, N173);
or OR3 (N3677, N3676, N7, N1008);
nor NOR4 (N3678, N3657, N1299, N5, N1272);
and AND4 (N3679, N3673, N2350, N2177, N1216);
nand NAND3 (N3680, N3678, N1982, N971);
xor XOR2 (N3681, N3649, N753);
not NOT1 (N3682, N3681);
xor XOR2 (N3683, N3682, N2858);
or OR4 (N3684, N3674, N2160, N2382, N279);
or OR4 (N3685, N3675, N3682, N1083, N1077);
buf BUF1 (N3686, N3677);
not NOT1 (N3687, N3684);
nand NAND4 (N3688, N3686, N3336, N1785, N1973);
xor XOR2 (N3689, N3685, N490);
not NOT1 (N3690, N3671);
not NOT1 (N3691, N3690);
not NOT1 (N3692, N3679);
buf BUF1 (N3693, N3680);
and AND4 (N3694, N3672, N1797, N2276, N941);
xor XOR2 (N3695, N3694, N426);
buf BUF1 (N3696, N3688);
not NOT1 (N3697, N3687);
not NOT1 (N3698, N3697);
buf BUF1 (N3699, N3693);
or OR4 (N3700, N3664, N3651, N2845, N1416);
and AND3 (N3701, N3695, N184, N243);
nor NOR4 (N3702, N3700, N1727, N3310, N1148);
buf BUF1 (N3703, N3689);
not NOT1 (N3704, N3692);
nor NOR3 (N3705, N3699, N2973, N350);
xor XOR2 (N3706, N3701, N1540);
or OR3 (N3707, N3705, N2952, N2761);
nand NAND4 (N3708, N3696, N1558, N577, N303);
not NOT1 (N3709, N3708);
or OR4 (N3710, N3702, N3272, N3348, N17);
or OR2 (N3711, N3709, N2891);
nor NOR4 (N3712, N3707, N1731, N291, N803);
xor XOR2 (N3713, N3703, N1250);
or OR2 (N3714, N3698, N2148);
buf BUF1 (N3715, N3665);
and AND2 (N3716, N3710, N1109);
nand NAND4 (N3717, N3711, N605, N3507, N1640);
buf BUF1 (N3718, N3704);
or OR3 (N3719, N3713, N3180, N2068);
and AND3 (N3720, N3718, N146, N2540);
nand NAND4 (N3721, N3706, N2206, N2238, N2681);
or OR4 (N3722, N3721, N738, N2602, N2576);
xor XOR2 (N3723, N3712, N2427);
xor XOR2 (N3724, N3715, N1532);
nor NOR2 (N3725, N3720, N162);
nand NAND2 (N3726, N3719, N545);
and AND4 (N3727, N3683, N861, N2356, N1883);
nor NOR4 (N3728, N3724, N2653, N414, N1551);
nor NOR2 (N3729, N3723, N1956);
xor XOR2 (N3730, N3725, N652);
or OR3 (N3731, N3729, N1305, N2385);
buf BUF1 (N3732, N3691);
not NOT1 (N3733, N3716);
nand NAND2 (N3734, N3731, N1026);
buf BUF1 (N3735, N3714);
xor XOR2 (N3736, N3734, N3358);
nor NOR4 (N3737, N3728, N3196, N1796, N528);
and AND4 (N3738, N3735, N2772, N1933, N2320);
and AND4 (N3739, N3726, N1521, N23, N3358);
not NOT1 (N3740, N3737);
buf BUF1 (N3741, N3732);
or OR4 (N3742, N3727, N1628, N1257, N3511);
or OR2 (N3743, N3740, N1192);
xor XOR2 (N3744, N3739, N1471);
or OR4 (N3745, N3736, N688, N2510, N2962);
xor XOR2 (N3746, N3742, N1587);
or OR2 (N3747, N3733, N3445);
not NOT1 (N3748, N3717);
buf BUF1 (N3749, N3744);
and AND3 (N3750, N3738, N2123, N3060);
xor XOR2 (N3751, N3722, N694);
and AND4 (N3752, N3748, N529, N938, N3125);
nand NAND2 (N3753, N3751, N2157);
or OR2 (N3754, N3752, N1416);
xor XOR2 (N3755, N3754, N2778);
and AND3 (N3756, N3750, N3214, N2769);
nand NAND3 (N3757, N3756, N2776, N939);
and AND2 (N3758, N3745, N610);
buf BUF1 (N3759, N3749);
nand NAND4 (N3760, N3758, N1877, N2645, N2788);
nand NAND2 (N3761, N3753, N3708);
or OR2 (N3762, N3747, N2869);
and AND4 (N3763, N3762, N1902, N137, N3661);
not NOT1 (N3764, N3761);
buf BUF1 (N3765, N3764);
xor XOR2 (N3766, N3763, N2075);
or OR2 (N3767, N3765, N724);
not NOT1 (N3768, N3767);
not NOT1 (N3769, N3730);
and AND4 (N3770, N3757, N3093, N729, N2446);
nor NOR3 (N3771, N3743, N3172, N2657);
xor XOR2 (N3772, N3769, N3409);
not NOT1 (N3773, N3755);
xor XOR2 (N3774, N3772, N2398);
or OR2 (N3775, N3768, N2843);
or OR2 (N3776, N3774, N1972);
and AND2 (N3777, N3759, N678);
nand NAND3 (N3778, N3741, N1656, N2276);
and AND3 (N3779, N3746, N1667, N2521);
and AND4 (N3780, N3771, N1628, N3665, N2061);
not NOT1 (N3781, N3776);
or OR2 (N3782, N3780, N2517);
or OR4 (N3783, N3766, N1160, N397, N236);
and AND3 (N3784, N3781, N2596, N2388);
xor XOR2 (N3785, N3775, N1162);
not NOT1 (N3786, N3779);
xor XOR2 (N3787, N3778, N3313);
buf BUF1 (N3788, N3787);
nand NAND4 (N3789, N3785, N1402, N1381, N3331);
buf BUF1 (N3790, N3777);
nand NAND3 (N3791, N3783, N3426, N537);
buf BUF1 (N3792, N3760);
nand NAND2 (N3793, N3770, N1143);
not NOT1 (N3794, N3782);
not NOT1 (N3795, N3788);
xor XOR2 (N3796, N3784, N3762);
not NOT1 (N3797, N3773);
xor XOR2 (N3798, N3791, N3550);
and AND4 (N3799, N3789, N1162, N317, N1299);
xor XOR2 (N3800, N3798, N87);
not NOT1 (N3801, N3790);
buf BUF1 (N3802, N3795);
buf BUF1 (N3803, N3800);
nand NAND3 (N3804, N3786, N2291, N127);
and AND3 (N3805, N3799, N673, N1423);
nand NAND3 (N3806, N3796, N3617, N1074);
nand NAND4 (N3807, N3802, N1965, N3166, N362);
xor XOR2 (N3808, N3797, N1996);
nand NAND3 (N3809, N3805, N3573, N3509);
xor XOR2 (N3810, N3792, N3338);
or OR4 (N3811, N3806, N3171, N2101, N337);
xor XOR2 (N3812, N3811, N2881);
xor XOR2 (N3813, N3804, N3471);
and AND3 (N3814, N3813, N3102, N2665);
not NOT1 (N3815, N3794);
and AND2 (N3816, N3810, N1618);
or OR3 (N3817, N3815, N1591, N1728);
not NOT1 (N3818, N3812);
buf BUF1 (N3819, N3808);
xor XOR2 (N3820, N3793, N805);
nor NOR4 (N3821, N3816, N1323, N1484, N9);
nand NAND3 (N3822, N3819, N1520, N3573);
nand NAND3 (N3823, N3822, N212, N3760);
not NOT1 (N3824, N3801);
or OR4 (N3825, N3820, N1910, N3129, N3706);
or OR3 (N3826, N3807, N1781, N6);
nor NOR4 (N3827, N3817, N2924, N668, N2189);
and AND2 (N3828, N3809, N985);
xor XOR2 (N3829, N3814, N2002);
nor NOR3 (N3830, N3821, N3091, N3004);
nor NOR2 (N3831, N3828, N3142);
buf BUF1 (N3832, N3803);
nand NAND3 (N3833, N3830, N1010, N1744);
and AND3 (N3834, N3831, N449, N701);
not NOT1 (N3835, N3833);
or OR2 (N3836, N3826, N656);
buf BUF1 (N3837, N3823);
buf BUF1 (N3838, N3836);
nor NOR4 (N3839, N3818, N1803, N1625, N1272);
or OR4 (N3840, N3827, N2818, N801, N752);
buf BUF1 (N3841, N3834);
nand NAND3 (N3842, N3839, N2344, N2401);
nor NOR4 (N3843, N3829, N440, N1716, N106);
or OR2 (N3844, N3824, N2887);
nand NAND4 (N3845, N3842, N2099, N2958, N2461);
buf BUF1 (N3846, N3835);
or OR4 (N3847, N3841, N3835, N2915, N1785);
nand NAND4 (N3848, N3832, N1203, N676, N3318);
or OR4 (N3849, N3848, N661, N1592, N2225);
nand NAND2 (N3850, N3847, N1836);
or OR4 (N3851, N3840, N605, N2072, N362);
or OR3 (N3852, N3851, N3442, N2565);
not NOT1 (N3853, N3837);
nand NAND3 (N3854, N3850, N3134, N2680);
buf BUF1 (N3855, N3838);
not NOT1 (N3856, N3843);
or OR3 (N3857, N3846, N263, N311);
nand NAND4 (N3858, N3854, N800, N883, N2578);
buf BUF1 (N3859, N3849);
nor NOR2 (N3860, N3845, N3002);
not NOT1 (N3861, N3856);
xor XOR2 (N3862, N3852, N3550);
and AND2 (N3863, N3853, N1618);
not NOT1 (N3864, N3855);
xor XOR2 (N3865, N3859, N479);
not NOT1 (N3866, N3844);
and AND3 (N3867, N3865, N1771, N2306);
buf BUF1 (N3868, N3862);
nor NOR2 (N3869, N3866, N3108);
not NOT1 (N3870, N3825);
buf BUF1 (N3871, N3861);
and AND2 (N3872, N3869, N2888);
xor XOR2 (N3873, N3871, N349);
not NOT1 (N3874, N3872);
nor NOR3 (N3875, N3870, N1073, N1936);
buf BUF1 (N3876, N3873);
nor NOR3 (N3877, N3868, N2603, N608);
not NOT1 (N3878, N3875);
nor NOR3 (N3879, N3874, N2736, N1619);
and AND2 (N3880, N3878, N2081);
nor NOR2 (N3881, N3880, N3055);
nor NOR4 (N3882, N3879, N2371, N2250, N3777);
nand NAND3 (N3883, N3857, N3868, N1889);
nor NOR4 (N3884, N3867, N2522, N3829, N3421);
nor NOR2 (N3885, N3858, N3694);
buf BUF1 (N3886, N3885);
buf BUF1 (N3887, N3864);
nand NAND3 (N3888, N3887, N2253, N3769);
and AND4 (N3889, N3876, N1440, N3501, N2624);
or OR2 (N3890, N3881, N1861);
xor XOR2 (N3891, N3890, N793);
not NOT1 (N3892, N3860);
xor XOR2 (N3893, N3882, N117);
or OR3 (N3894, N3883, N1681, N2829);
nand NAND2 (N3895, N3877, N1510);
buf BUF1 (N3896, N3884);
and AND2 (N3897, N3892, N2812);
buf BUF1 (N3898, N3895);
xor XOR2 (N3899, N3891, N2527);
nand NAND3 (N3900, N3899, N1331, N2107);
xor XOR2 (N3901, N3888, N1316);
buf BUF1 (N3902, N3894);
and AND4 (N3903, N3886, N2303, N2805, N2046);
buf BUF1 (N3904, N3893);
xor XOR2 (N3905, N3904, N2977);
nor NOR2 (N3906, N3901, N2596);
nor NOR3 (N3907, N3902, N1850, N78);
xor XOR2 (N3908, N3897, N1187);
nand NAND3 (N3909, N3896, N1075, N525);
or OR3 (N3910, N3905, N900, N662);
nor NOR3 (N3911, N3889, N1979, N3286);
buf BUF1 (N3912, N3910);
or OR3 (N3913, N3900, N3407, N2605);
nand NAND4 (N3914, N3911, N781, N672, N3473);
nor NOR3 (N3915, N3907, N3088, N306);
xor XOR2 (N3916, N3912, N3431);
buf BUF1 (N3917, N3903);
xor XOR2 (N3918, N3898, N2779);
and AND3 (N3919, N3906, N3305, N1041);
buf BUF1 (N3920, N3918);
nand NAND2 (N3921, N3913, N277);
nand NAND3 (N3922, N3921, N868, N3564);
nand NAND3 (N3923, N3922, N1248, N476);
nand NAND2 (N3924, N3909, N238);
and AND3 (N3925, N3919, N2734, N677);
nand NAND4 (N3926, N3863, N1916, N2208, N2479);
buf BUF1 (N3927, N3920);
nand NAND3 (N3928, N3924, N2425, N1667);
or OR3 (N3929, N3927, N172, N2933);
nand NAND4 (N3930, N3908, N3093, N1892, N450);
not NOT1 (N3931, N3930);
not NOT1 (N3932, N3914);
or OR3 (N3933, N3915, N3917, N1928);
not NOT1 (N3934, N996);
and AND2 (N3935, N3923, N1799);
xor XOR2 (N3936, N3916, N2002);
nor NOR4 (N3937, N3936, N599, N125, N749);
and AND4 (N3938, N3932, N1633, N344, N2549);
xor XOR2 (N3939, N3928, N517);
nor NOR2 (N3940, N3933, N3540);
not NOT1 (N3941, N3939);
xor XOR2 (N3942, N3925, N2355);
nor NOR3 (N3943, N3926, N3602, N3687);
nand NAND2 (N3944, N3942, N1665);
nand NAND2 (N3945, N3940, N409);
not NOT1 (N3946, N3931);
and AND2 (N3947, N3934, N2145);
or OR4 (N3948, N3938, N549, N509, N2394);
or OR2 (N3949, N3947, N856);
nand NAND2 (N3950, N3937, N74);
xor XOR2 (N3951, N3946, N1835);
nor NOR4 (N3952, N3943, N298, N1068, N58);
buf BUF1 (N3953, N3935);
or OR4 (N3954, N3945, N566, N88, N2196);
or OR2 (N3955, N3950, N1512);
buf BUF1 (N3956, N3951);
nor NOR4 (N3957, N3941, N2749, N1414, N1537);
or OR3 (N3958, N3956, N2003, N2740);
and AND3 (N3959, N3958, N418, N1203);
nand NAND2 (N3960, N3957, N3648);
and AND4 (N3961, N3952, N2900, N2229, N1118);
xor XOR2 (N3962, N3949, N1378);
nand NAND3 (N3963, N3955, N1450, N2603);
xor XOR2 (N3964, N3953, N534);
buf BUF1 (N3965, N3959);
and AND3 (N3966, N3954, N120, N1632);
xor XOR2 (N3967, N3963, N3230);
nand NAND2 (N3968, N3966, N1061);
or OR2 (N3969, N3944, N3521);
buf BUF1 (N3970, N3961);
or OR2 (N3971, N3965, N2461);
nand NAND4 (N3972, N3968, N2945, N225, N291);
nand NAND3 (N3973, N3962, N2154, N2696);
xor XOR2 (N3974, N3964, N2253);
xor XOR2 (N3975, N3967, N2523);
and AND3 (N3976, N3972, N1329, N1821);
xor XOR2 (N3977, N3960, N3512);
and AND4 (N3978, N3970, N2632, N604, N429);
not NOT1 (N3979, N3948);
nor NOR3 (N3980, N3976, N1032, N724);
nand NAND2 (N3981, N3969, N3192);
and AND3 (N3982, N3973, N2850, N1524);
nand NAND2 (N3983, N3978, N2947);
not NOT1 (N3984, N3983);
buf BUF1 (N3985, N3971);
nor NOR3 (N3986, N3975, N1394, N1659);
nand NAND3 (N3987, N3982, N421, N2832);
nor NOR3 (N3988, N3985, N319, N1730);
or OR2 (N3989, N3984, N2620);
buf BUF1 (N3990, N3980);
xor XOR2 (N3991, N3979, N3227);
nor NOR4 (N3992, N3987, N3329, N1316, N2252);
xor XOR2 (N3993, N3988, N2504);
not NOT1 (N3994, N3993);
xor XOR2 (N3995, N3990, N74);
xor XOR2 (N3996, N3994, N2749);
not NOT1 (N3997, N3929);
or OR3 (N3998, N3974, N1115, N1969);
and AND4 (N3999, N3995, N584, N25, N1986);
nand NAND4 (N4000, N3989, N3601, N3827, N106);
and AND3 (N4001, N3981, N332, N81);
nor NOR2 (N4002, N3999, N3643);
buf BUF1 (N4003, N3996);
nor NOR4 (N4004, N3991, N1122, N2598, N84);
buf BUF1 (N4005, N3997);
or OR4 (N4006, N4002, N147, N2078, N3914);
or OR2 (N4007, N4000, N1329);
nor NOR4 (N4008, N3977, N88, N2910, N3550);
not NOT1 (N4009, N3986);
nor NOR4 (N4010, N4004, N939, N1275, N834);
nand NAND2 (N4011, N4001, N3327);
or OR2 (N4012, N4006, N2898);
not NOT1 (N4013, N4009);
xor XOR2 (N4014, N4012, N182);
nand NAND3 (N4015, N4013, N1908, N992);
buf BUF1 (N4016, N3998);
xor XOR2 (N4017, N4016, N2160);
not NOT1 (N4018, N3992);
or OR4 (N4019, N4008, N3975, N592, N2622);
not NOT1 (N4020, N4005);
nor NOR4 (N4021, N4018, N1001, N2446, N982);
nor NOR2 (N4022, N4010, N3336);
endmodule