// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17;

output N8011,N8013,N8014,N8007,N8016,N8012,N7998,N8003,N8010,N8017;

nor NOR2 (N18, N14, N4);
nand NAND2 (N19, N5, N6);
xor XOR2 (N20, N1, N19);
nor NOR2 (N21, N16, N13);
xor XOR2 (N22, N2, N4);
xor XOR2 (N23, N7, N12);
buf BUF1 (N24, N17);
nand NAND3 (N25, N1, N24, N24);
xor XOR2 (N26, N11, N7);
nor NOR4 (N27, N20, N26, N11, N12);
buf BUF1 (N28, N10);
nand NAND3 (N29, N27, N26, N15);
buf BUF1 (N30, N26);
not NOT1 (N31, N13);
xor XOR2 (N32, N7, N2);
or OR4 (N33, N25, N11, N8, N17);
or OR2 (N34, N23, N32);
nor NOR2 (N35, N2, N10);
buf BUF1 (N36, N30);
and AND4 (N37, N28, N5, N26, N4);
xor XOR2 (N38, N34, N1);
or OR2 (N39, N22, N16);
or OR2 (N40, N37, N34);
nor NOR3 (N41, N31, N26, N10);
and AND4 (N42, N36, N31, N38, N25);
buf BUF1 (N43, N10);
not NOT1 (N44, N21);
xor XOR2 (N45, N42, N44);
buf BUF1 (N46, N35);
nand NAND3 (N47, N13, N5, N14);
buf BUF1 (N48, N39);
nor NOR2 (N49, N43, N3);
not NOT1 (N50, N29);
xor XOR2 (N51, N18, N1);
not NOT1 (N52, N33);
not NOT1 (N53, N41);
or OR4 (N54, N50, N50, N4, N17);
nor NOR3 (N55, N45, N44, N22);
nand NAND3 (N56, N53, N24, N45);
nor NOR2 (N57, N40, N24);
nand NAND4 (N58, N49, N49, N47, N51);
or OR3 (N59, N14, N20, N57);
xor XOR2 (N60, N31, N4);
not NOT1 (N61, N23);
buf BUF1 (N62, N58);
nor NOR2 (N63, N52, N30);
buf BUF1 (N64, N59);
not NOT1 (N65, N46);
nand NAND3 (N66, N55, N62, N3);
nand NAND4 (N67, N45, N62, N24, N41);
nand NAND4 (N68, N56, N25, N61, N7);
buf BUF1 (N69, N19);
or OR3 (N70, N65, N9, N16);
not NOT1 (N71, N48);
buf BUF1 (N72, N66);
nor NOR3 (N73, N63, N3, N64);
and AND3 (N74, N53, N40, N71);
and AND4 (N75, N10, N28, N58, N32);
nor NOR2 (N76, N72, N14);
and AND3 (N77, N54, N52, N36);
buf BUF1 (N78, N68);
nand NAND3 (N79, N60, N30, N55);
nor NOR3 (N80, N79, N5, N74);
not NOT1 (N81, N41);
nand NAND4 (N82, N69, N44, N27, N51);
not NOT1 (N83, N82);
xor XOR2 (N84, N75, N65);
and AND4 (N85, N80, N58, N19, N14);
nor NOR3 (N86, N81, N71, N65);
not NOT1 (N87, N70);
and AND2 (N88, N86, N15);
and AND3 (N89, N67, N66, N7);
and AND4 (N90, N84, N33, N69, N78);
and AND2 (N91, N36, N82);
buf BUF1 (N92, N83);
nand NAND4 (N93, N76, N36, N49, N16);
and AND4 (N94, N85, N32, N93, N72);
xor XOR2 (N95, N62, N83);
and AND2 (N96, N94, N6);
nand NAND4 (N97, N96, N42, N10, N4);
and AND3 (N98, N77, N97, N34);
xor XOR2 (N99, N51, N95);
or OR2 (N100, N3, N46);
and AND4 (N101, N88, N27, N79, N74);
nand NAND4 (N102, N98, N16, N69, N61);
nand NAND3 (N103, N101, N4, N32);
xor XOR2 (N104, N100, N43);
not NOT1 (N105, N99);
and AND4 (N106, N89, N84, N46, N64);
xor XOR2 (N107, N92, N22);
not NOT1 (N108, N106);
nor NOR3 (N109, N104, N30, N4);
and AND3 (N110, N87, N57, N71);
xor XOR2 (N111, N108, N90);
nand NAND3 (N112, N93, N58, N30);
not NOT1 (N113, N103);
buf BUF1 (N114, N109);
nand NAND3 (N115, N73, N71, N61);
or OR2 (N116, N102, N70);
or OR4 (N117, N91, N8, N46, N48);
nor NOR4 (N118, N111, N54, N58, N77);
not NOT1 (N119, N107);
and AND2 (N120, N105, N31);
nor NOR2 (N121, N112, N120);
or OR4 (N122, N54, N72, N22, N26);
xor XOR2 (N123, N110, N90);
not NOT1 (N124, N117);
nor NOR4 (N125, N115, N80, N110, N51);
buf BUF1 (N126, N124);
buf BUF1 (N127, N125);
not NOT1 (N128, N122);
buf BUF1 (N129, N127);
buf BUF1 (N130, N129);
not NOT1 (N131, N119);
nand NAND3 (N132, N121, N103, N43);
and AND2 (N133, N118, N120);
or OR3 (N134, N132, N14, N98);
or OR3 (N135, N130, N49, N30);
buf BUF1 (N136, N123);
or OR2 (N137, N113, N33);
buf BUF1 (N138, N137);
nor NOR3 (N139, N116, N17, N45);
and AND2 (N140, N138, N39);
xor XOR2 (N141, N128, N3);
not NOT1 (N142, N133);
buf BUF1 (N143, N140);
nor NOR2 (N144, N135, N43);
nor NOR2 (N145, N134, N130);
or OR4 (N146, N142, N11, N72, N125);
and AND4 (N147, N143, N51, N45, N82);
and AND4 (N148, N146, N12, N48, N74);
not NOT1 (N149, N145);
nor NOR4 (N150, N136, N33, N51, N86);
xor XOR2 (N151, N141, N46);
buf BUF1 (N152, N149);
and AND2 (N153, N131, N72);
nor NOR4 (N154, N126, N126, N20, N114);
nand NAND2 (N155, N55, N120);
or OR4 (N156, N154, N23, N96, N35);
buf BUF1 (N157, N148);
xor XOR2 (N158, N152, N58);
xor XOR2 (N159, N158, N113);
and AND4 (N160, N159, N84, N15, N100);
not NOT1 (N161, N155);
and AND2 (N162, N144, N153);
xor XOR2 (N163, N53, N39);
xor XOR2 (N164, N160, N33);
nor NOR2 (N165, N161, N44);
nor NOR2 (N166, N150, N117);
not NOT1 (N167, N157);
buf BUF1 (N168, N165);
xor XOR2 (N169, N147, N79);
nand NAND4 (N170, N151, N132, N108, N21);
xor XOR2 (N171, N170, N81);
or OR2 (N172, N166, N61);
or OR4 (N173, N171, N96, N81, N32);
or OR2 (N174, N167, N92);
buf BUF1 (N175, N173);
nor NOR3 (N176, N156, N52, N30);
xor XOR2 (N177, N162, N35);
buf BUF1 (N178, N175);
xor XOR2 (N179, N174, N114);
not NOT1 (N180, N163);
not NOT1 (N181, N177);
nor NOR2 (N182, N180, N81);
buf BUF1 (N183, N176);
buf BUF1 (N184, N164);
nand NAND3 (N185, N178, N138, N67);
nor NOR3 (N186, N139, N11, N9);
or OR4 (N187, N169, N24, N162, N60);
or OR4 (N188, N172, N103, N155, N24);
nand NAND3 (N189, N182, N152, N181);
nand NAND2 (N190, N178, N40);
not NOT1 (N191, N168);
and AND2 (N192, N184, N134);
and AND2 (N193, N191, N160);
or OR2 (N194, N187, N190);
nor NOR2 (N195, N106, N138);
buf BUF1 (N196, N194);
nor NOR4 (N197, N185, N77, N56, N7);
buf BUF1 (N198, N193);
nor NOR3 (N199, N179, N113, N56);
nor NOR2 (N200, N189, N17);
nor NOR2 (N201, N183, N191);
buf BUF1 (N202, N201);
xor XOR2 (N203, N192, N166);
nor NOR4 (N204, N202, N181, N176, N49);
nand NAND2 (N205, N188, N58);
and AND3 (N206, N195, N113, N119);
or OR4 (N207, N199, N80, N27, N173);
or OR4 (N208, N204, N16, N36, N169);
xor XOR2 (N209, N200, N16);
and AND4 (N210, N205, N172, N131, N195);
not NOT1 (N211, N196);
not NOT1 (N212, N206);
buf BUF1 (N213, N208);
or OR3 (N214, N198, N27, N179);
xor XOR2 (N215, N212, N61);
not NOT1 (N216, N197);
not NOT1 (N217, N216);
or OR3 (N218, N213, N56, N215);
xor XOR2 (N219, N77, N47);
nor NOR2 (N220, N186, N194);
or OR2 (N221, N211, N80);
not NOT1 (N222, N219);
and AND3 (N223, N221, N151, N17);
not NOT1 (N224, N207);
nor NOR2 (N225, N220, N108);
not NOT1 (N226, N209);
xor XOR2 (N227, N218, N208);
not NOT1 (N228, N210);
nand NAND4 (N229, N227, N42, N101, N143);
and AND4 (N230, N228, N116, N134, N14);
and AND3 (N231, N223, N109, N70);
not NOT1 (N232, N231);
xor XOR2 (N233, N226, N131);
or OR4 (N234, N203, N233, N172, N81);
nor NOR2 (N235, N216, N100);
not NOT1 (N236, N222);
xor XOR2 (N237, N217, N98);
not NOT1 (N238, N214);
nor NOR4 (N239, N235, N128, N77, N63);
not NOT1 (N240, N238);
or OR3 (N241, N224, N99, N52);
or OR3 (N242, N229, N44, N97);
not NOT1 (N243, N237);
buf BUF1 (N244, N240);
buf BUF1 (N245, N242);
buf BUF1 (N246, N239);
or OR3 (N247, N234, N238, N164);
nor NOR4 (N248, N247, N95, N14, N194);
nor NOR2 (N249, N244, N193);
or OR4 (N250, N243, N77, N115, N152);
not NOT1 (N251, N250);
xor XOR2 (N252, N245, N194);
buf BUF1 (N253, N236);
or OR2 (N254, N241, N129);
and AND3 (N255, N251, N25, N6);
and AND4 (N256, N248, N112, N115, N130);
buf BUF1 (N257, N256);
nand NAND3 (N258, N232, N239, N95);
buf BUF1 (N259, N257);
and AND2 (N260, N225, N209);
xor XOR2 (N261, N249, N169);
not NOT1 (N262, N253);
nor NOR2 (N263, N254, N237);
not NOT1 (N264, N255);
or OR3 (N265, N258, N235, N122);
xor XOR2 (N266, N264, N186);
xor XOR2 (N267, N260, N64);
nor NOR4 (N268, N263, N183, N229, N77);
or OR3 (N269, N268, N129, N179);
not NOT1 (N270, N267);
buf BUF1 (N271, N266);
not NOT1 (N272, N230);
and AND2 (N273, N270, N198);
and AND2 (N274, N246, N86);
buf BUF1 (N275, N271);
not NOT1 (N276, N252);
nor NOR2 (N277, N269, N84);
not NOT1 (N278, N274);
nand NAND4 (N279, N278, N125, N73, N134);
nor NOR2 (N280, N265, N185);
buf BUF1 (N281, N272);
buf BUF1 (N282, N261);
or OR3 (N283, N277, N103, N39);
nand NAND3 (N284, N283, N176, N97);
nor NOR2 (N285, N275, N227);
nand NAND3 (N286, N284, N101, N81);
nand NAND4 (N287, N280, N194, N178, N218);
and AND3 (N288, N287, N237, N110);
not NOT1 (N289, N259);
xor XOR2 (N290, N286, N75);
or OR3 (N291, N289, N94, N268);
nand NAND4 (N292, N288, N137, N188, N141);
and AND3 (N293, N292, N56, N11);
nor NOR4 (N294, N276, N200, N137, N138);
buf BUF1 (N295, N285);
not NOT1 (N296, N290);
and AND2 (N297, N295, N77);
buf BUF1 (N298, N293);
or OR4 (N299, N279, N277, N211, N157);
or OR4 (N300, N282, N228, N140, N56);
not NOT1 (N301, N262);
nand NAND3 (N302, N298, N270, N215);
or OR2 (N303, N301, N172);
or OR3 (N304, N291, N171, N210);
and AND2 (N305, N294, N101);
buf BUF1 (N306, N273);
buf BUF1 (N307, N297);
buf BUF1 (N308, N299);
buf BUF1 (N309, N303);
buf BUF1 (N310, N302);
xor XOR2 (N311, N309, N13);
nand NAND4 (N312, N311, N98, N25, N305);
not NOT1 (N313, N166);
xor XOR2 (N314, N313, N58);
not NOT1 (N315, N312);
nand NAND2 (N316, N307, N144);
or OR2 (N317, N304, N298);
and AND3 (N318, N315, N77, N76);
xor XOR2 (N319, N281, N52);
buf BUF1 (N320, N319);
and AND4 (N321, N318, N31, N208, N180);
not NOT1 (N322, N310);
and AND3 (N323, N321, N55, N252);
or OR4 (N324, N308, N149, N201, N131);
not NOT1 (N325, N296);
nor NOR4 (N326, N323, N197, N161, N152);
or OR3 (N327, N317, N232, N270);
buf BUF1 (N328, N300);
xor XOR2 (N329, N328, N61);
buf BUF1 (N330, N306);
nor NOR3 (N331, N322, N64, N229);
and AND2 (N332, N330, N159);
nor NOR3 (N333, N327, N151, N201);
nor NOR3 (N334, N316, N120, N180);
and AND3 (N335, N314, N246, N220);
xor XOR2 (N336, N324, N219);
buf BUF1 (N337, N332);
not NOT1 (N338, N333);
buf BUF1 (N339, N335);
nor NOR4 (N340, N336, N281, N68, N64);
nor NOR3 (N341, N320, N222, N2);
xor XOR2 (N342, N338, N8);
nor NOR3 (N343, N325, N107, N2);
nand NAND2 (N344, N340, N158);
nand NAND2 (N345, N331, N63);
nor NOR2 (N346, N326, N338);
buf BUF1 (N347, N344);
nand NAND4 (N348, N339, N20, N282, N164);
buf BUF1 (N349, N346);
or OR2 (N350, N329, N133);
xor XOR2 (N351, N347, N128);
buf BUF1 (N352, N348);
nor NOR3 (N353, N341, N270, N170);
or OR4 (N354, N349, N248, N84, N262);
nand NAND4 (N355, N352, N259, N109, N312);
and AND4 (N356, N334, N47, N72, N266);
not NOT1 (N357, N356);
or OR4 (N358, N350, N175, N289, N225);
not NOT1 (N359, N358);
buf BUF1 (N360, N343);
nor NOR2 (N361, N360, N85);
buf BUF1 (N362, N345);
or OR2 (N363, N359, N238);
nor NOR3 (N364, N342, N11, N344);
nand NAND2 (N365, N353, N185);
or OR2 (N366, N364, N234);
buf BUF1 (N367, N357);
nor NOR2 (N368, N363, N179);
or OR4 (N369, N365, N216, N105, N316);
nor NOR2 (N370, N354, N67);
not NOT1 (N371, N351);
buf BUF1 (N372, N355);
xor XOR2 (N373, N367, N199);
not NOT1 (N374, N371);
buf BUF1 (N375, N361);
and AND2 (N376, N362, N343);
nor NOR2 (N377, N368, N97);
not NOT1 (N378, N376);
and AND3 (N379, N374, N330, N45);
not NOT1 (N380, N373);
nand NAND3 (N381, N378, N184, N161);
xor XOR2 (N382, N379, N219);
not NOT1 (N383, N369);
xor XOR2 (N384, N381, N47);
not NOT1 (N385, N382);
and AND2 (N386, N384, N38);
nor NOR4 (N387, N377, N374, N333, N164);
nand NAND2 (N388, N337, N200);
buf BUF1 (N389, N388);
not NOT1 (N390, N366);
not NOT1 (N391, N387);
or OR4 (N392, N385, N194, N116, N391);
xor XOR2 (N393, N288, N176);
not NOT1 (N394, N386);
buf BUF1 (N395, N389);
or OR3 (N396, N392, N54, N158);
xor XOR2 (N397, N390, N200);
not NOT1 (N398, N396);
not NOT1 (N399, N370);
and AND2 (N400, N398, N274);
nor NOR3 (N401, N397, N258, N106);
or OR2 (N402, N401, N307);
nor NOR2 (N403, N393, N374);
xor XOR2 (N404, N380, N26);
nand NAND4 (N405, N394, N371, N370, N330);
or OR4 (N406, N403, N183, N397, N90);
and AND4 (N407, N402, N111, N179, N346);
nor NOR4 (N408, N383, N247, N272, N369);
nand NAND2 (N409, N407, N66);
xor XOR2 (N410, N400, N158);
xor XOR2 (N411, N406, N305);
buf BUF1 (N412, N395);
buf BUF1 (N413, N411);
or OR2 (N414, N408, N299);
xor XOR2 (N415, N399, N53);
buf BUF1 (N416, N409);
and AND4 (N417, N410, N58, N132, N64);
nor NOR2 (N418, N415, N231);
buf BUF1 (N419, N413);
not NOT1 (N420, N412);
nor NOR4 (N421, N414, N358, N166, N294);
buf BUF1 (N422, N372);
nand NAND4 (N423, N404, N171, N102, N304);
xor XOR2 (N424, N423, N139);
buf BUF1 (N425, N405);
buf BUF1 (N426, N422);
or OR2 (N427, N416, N400);
or OR3 (N428, N424, N97, N43);
xor XOR2 (N429, N419, N102);
nor NOR2 (N430, N418, N38);
nor NOR2 (N431, N425, N18);
nand NAND2 (N432, N427, N205);
nor NOR3 (N433, N420, N117, N312);
nand NAND2 (N434, N421, N150);
not NOT1 (N435, N428);
not NOT1 (N436, N426);
not NOT1 (N437, N431);
and AND2 (N438, N417, N240);
buf BUF1 (N439, N438);
nor NOR2 (N440, N433, N65);
and AND4 (N441, N375, N334, N338, N90);
and AND2 (N442, N435, N76);
and AND3 (N443, N432, N392, N389);
nand NAND2 (N444, N437, N243);
nand NAND4 (N445, N442, N404, N232, N361);
and AND2 (N446, N444, N350);
not NOT1 (N447, N446);
nor NOR3 (N448, N443, N444, N324);
and AND4 (N449, N429, N344, N260, N129);
not NOT1 (N450, N441);
not NOT1 (N451, N449);
not NOT1 (N452, N434);
not NOT1 (N453, N448);
and AND2 (N454, N439, N8);
and AND2 (N455, N453, N414);
xor XOR2 (N456, N447, N22);
xor XOR2 (N457, N454, N427);
nor NOR3 (N458, N450, N355, N65);
and AND3 (N459, N456, N413, N33);
nand NAND2 (N460, N451, N431);
buf BUF1 (N461, N430);
or OR4 (N462, N457, N411, N392, N336);
xor XOR2 (N463, N458, N255);
not NOT1 (N464, N459);
xor XOR2 (N465, N464, N330);
not NOT1 (N466, N460);
xor XOR2 (N467, N452, N90);
or OR4 (N468, N461, N108, N428, N421);
not NOT1 (N469, N462);
and AND2 (N470, N468, N438);
or OR2 (N471, N467, N233);
buf BUF1 (N472, N436);
xor XOR2 (N473, N465, N98);
nand NAND3 (N474, N469, N230, N152);
buf BUF1 (N475, N472);
nor NOR2 (N476, N440, N247);
xor XOR2 (N477, N455, N302);
nand NAND4 (N478, N445, N406, N74, N112);
buf BUF1 (N479, N475);
nor NOR4 (N480, N466, N130, N312, N385);
xor XOR2 (N481, N476, N32);
nor NOR4 (N482, N480, N354, N151, N157);
nor NOR2 (N483, N470, N105);
xor XOR2 (N484, N479, N94);
xor XOR2 (N485, N471, N396);
buf BUF1 (N486, N473);
buf BUF1 (N487, N477);
and AND4 (N488, N463, N232, N316, N350);
not NOT1 (N489, N486);
nor NOR4 (N490, N478, N236, N56, N333);
xor XOR2 (N491, N487, N199);
buf BUF1 (N492, N488);
nor NOR2 (N493, N490, N444);
nand NAND4 (N494, N481, N80, N377, N92);
nand NAND3 (N495, N492, N271, N350);
nand NAND3 (N496, N494, N263, N434);
buf BUF1 (N497, N484);
or OR2 (N498, N491, N157);
or OR3 (N499, N496, N173, N246);
xor XOR2 (N500, N489, N225);
and AND3 (N501, N482, N55, N311);
and AND2 (N502, N474, N191);
or OR2 (N503, N497, N103);
buf BUF1 (N504, N483);
not NOT1 (N505, N501);
nor NOR4 (N506, N502, N495, N409, N193);
xor XOR2 (N507, N119, N324);
xor XOR2 (N508, N503, N147);
buf BUF1 (N509, N493);
buf BUF1 (N510, N506);
nor NOR3 (N511, N485, N139, N130);
nand NAND2 (N512, N511, N39);
nand NAND2 (N513, N508, N260);
and AND4 (N514, N513, N432, N370, N143);
or OR3 (N515, N512, N375, N88);
or OR2 (N516, N509, N456);
xor XOR2 (N517, N515, N400);
xor XOR2 (N518, N505, N32);
not NOT1 (N519, N510);
nand NAND2 (N520, N500, N124);
or OR4 (N521, N504, N313, N439, N47);
nor NOR2 (N522, N498, N521);
xor XOR2 (N523, N403, N102);
not NOT1 (N524, N514);
nor NOR3 (N525, N516, N233, N445);
and AND2 (N526, N519, N502);
nor NOR3 (N527, N499, N24, N452);
or OR3 (N528, N526, N319, N509);
xor XOR2 (N529, N517, N5);
and AND3 (N530, N522, N349, N316);
not NOT1 (N531, N530);
not NOT1 (N532, N529);
or OR3 (N533, N528, N35, N389);
nand NAND4 (N534, N532, N229, N403, N49);
not NOT1 (N535, N525);
nand NAND4 (N536, N527, N294, N108, N214);
nand NAND4 (N537, N531, N404, N486, N337);
xor XOR2 (N538, N533, N14);
or OR4 (N539, N538, N211, N431, N166);
not NOT1 (N540, N534);
nor NOR2 (N541, N539, N441);
buf BUF1 (N542, N536);
xor XOR2 (N543, N540, N103);
not NOT1 (N544, N520);
xor XOR2 (N545, N523, N151);
nor NOR3 (N546, N537, N430, N199);
xor XOR2 (N547, N543, N147);
nor NOR3 (N548, N535, N146, N452);
or OR4 (N549, N524, N435, N422, N66);
and AND3 (N550, N546, N79, N228);
xor XOR2 (N551, N541, N36);
and AND3 (N552, N550, N465, N124);
nor NOR2 (N553, N549, N68);
not NOT1 (N554, N542);
buf BUF1 (N555, N545);
and AND2 (N556, N551, N14);
not NOT1 (N557, N554);
nand NAND3 (N558, N548, N217, N17);
nand NAND4 (N559, N556, N258, N536, N153);
nand NAND2 (N560, N552, N367);
and AND3 (N561, N558, N409, N442);
xor XOR2 (N562, N507, N85);
buf BUF1 (N563, N557);
or OR3 (N564, N563, N246, N66);
and AND2 (N565, N562, N336);
nand NAND2 (N566, N547, N49);
nand NAND4 (N567, N553, N546, N422, N205);
nor NOR4 (N568, N555, N116, N67, N485);
xor XOR2 (N569, N559, N517);
not NOT1 (N570, N565);
buf BUF1 (N571, N567);
nor NOR4 (N572, N566, N324, N416, N71);
xor XOR2 (N573, N568, N195);
or OR2 (N574, N570, N548);
nor NOR3 (N575, N518, N359, N165);
buf BUF1 (N576, N560);
nor NOR3 (N577, N544, N318, N489);
not NOT1 (N578, N571);
buf BUF1 (N579, N574);
not NOT1 (N580, N578);
buf BUF1 (N581, N580);
nor NOR3 (N582, N579, N144, N213);
nand NAND2 (N583, N572, N112);
nor NOR2 (N584, N581, N350);
or OR4 (N585, N582, N308, N166, N354);
not NOT1 (N586, N561);
nand NAND3 (N587, N585, N135, N483);
and AND2 (N588, N575, N69);
nor NOR3 (N589, N573, N212, N118);
xor XOR2 (N590, N584, N116);
or OR3 (N591, N590, N208, N496);
and AND2 (N592, N583, N475);
and AND2 (N593, N592, N225);
nand NAND2 (N594, N591, N565);
xor XOR2 (N595, N594, N299);
buf BUF1 (N596, N564);
or OR2 (N597, N593, N30);
buf BUF1 (N598, N588);
not NOT1 (N599, N598);
nor NOR2 (N600, N599, N577);
not NOT1 (N601, N232);
buf BUF1 (N602, N601);
or OR3 (N603, N589, N218, N213);
not NOT1 (N604, N569);
xor XOR2 (N605, N595, N216);
buf BUF1 (N606, N603);
nand NAND2 (N607, N596, N1);
or OR3 (N608, N604, N69, N97);
and AND2 (N609, N597, N474);
nand NAND2 (N610, N602, N121);
not NOT1 (N611, N608);
or OR2 (N612, N600, N393);
buf BUF1 (N613, N587);
nor NOR4 (N614, N605, N174, N385, N177);
xor XOR2 (N615, N606, N573);
or OR3 (N616, N586, N522, N148);
buf BUF1 (N617, N613);
or OR2 (N618, N612, N239);
or OR2 (N619, N618, N158);
xor XOR2 (N620, N619, N111);
xor XOR2 (N621, N615, N443);
nor NOR4 (N622, N609, N219, N293, N438);
xor XOR2 (N623, N617, N467);
xor XOR2 (N624, N620, N312);
buf BUF1 (N625, N576);
nand NAND4 (N626, N623, N177, N135, N518);
and AND4 (N627, N614, N264, N229, N322);
nor NOR4 (N628, N621, N386, N1, N496);
or OR3 (N629, N616, N478, N455);
xor XOR2 (N630, N626, N454);
buf BUF1 (N631, N627);
nor NOR2 (N632, N628, N149);
nor NOR4 (N633, N630, N330, N592, N108);
and AND3 (N634, N633, N547, N347);
buf BUF1 (N635, N625);
nor NOR3 (N636, N624, N272, N290);
xor XOR2 (N637, N636, N136);
nor NOR2 (N638, N607, N42);
buf BUF1 (N639, N634);
xor XOR2 (N640, N638, N47);
not NOT1 (N641, N622);
or OR4 (N642, N632, N538, N419, N396);
not NOT1 (N643, N631);
nand NAND4 (N644, N639, N570, N564, N607);
xor XOR2 (N645, N642, N507);
xor XOR2 (N646, N635, N528);
nor NOR3 (N647, N611, N278, N32);
xor XOR2 (N648, N629, N235);
buf BUF1 (N649, N640);
nor NOR3 (N650, N645, N641, N317);
buf BUF1 (N651, N86);
xor XOR2 (N652, N651, N86);
xor XOR2 (N653, N650, N46);
xor XOR2 (N654, N610, N582);
not NOT1 (N655, N646);
and AND4 (N656, N647, N543, N448, N368);
not NOT1 (N657, N655);
and AND2 (N658, N649, N642);
nor NOR3 (N659, N644, N340, N282);
xor XOR2 (N660, N648, N624);
or OR3 (N661, N659, N493, N641);
not NOT1 (N662, N653);
nand NAND2 (N663, N652, N322);
nor NOR3 (N664, N643, N129, N45);
nor NOR3 (N665, N658, N232, N90);
xor XOR2 (N666, N654, N488);
nand NAND2 (N667, N663, N264);
and AND2 (N668, N666, N102);
not NOT1 (N669, N665);
nand NAND3 (N670, N656, N229, N515);
xor XOR2 (N671, N668, N168);
and AND3 (N672, N664, N81, N545);
not NOT1 (N673, N671);
not NOT1 (N674, N667);
nor NOR2 (N675, N661, N507);
xor XOR2 (N676, N662, N63);
or OR4 (N677, N673, N327, N495, N19);
xor XOR2 (N678, N676, N93);
xor XOR2 (N679, N637, N444);
or OR3 (N680, N679, N451, N79);
and AND3 (N681, N675, N474, N397);
xor XOR2 (N682, N672, N359);
buf BUF1 (N683, N657);
xor XOR2 (N684, N670, N79);
nor NOR2 (N685, N677, N481);
nor NOR4 (N686, N678, N142, N52, N97);
not NOT1 (N687, N680);
or OR3 (N688, N686, N30, N245);
not NOT1 (N689, N685);
or OR2 (N690, N687, N86);
not NOT1 (N691, N689);
buf BUF1 (N692, N681);
or OR3 (N693, N682, N336, N625);
buf BUF1 (N694, N692);
or OR4 (N695, N691, N135, N691, N446);
nor NOR4 (N696, N694, N78, N386, N456);
buf BUF1 (N697, N688);
nor NOR2 (N698, N693, N682);
or OR3 (N699, N698, N645, N54);
not NOT1 (N700, N683);
and AND3 (N701, N669, N112, N399);
not NOT1 (N702, N700);
nand NAND2 (N703, N684, N287);
and AND3 (N704, N690, N410, N669);
not NOT1 (N705, N696);
not NOT1 (N706, N702);
or OR3 (N707, N704, N254, N384);
and AND4 (N708, N697, N112, N466, N167);
nor NOR4 (N709, N707, N156, N673, N75);
not NOT1 (N710, N705);
xor XOR2 (N711, N695, N395);
nand NAND2 (N712, N710, N40);
buf BUF1 (N713, N708);
nand NAND2 (N714, N709, N82);
and AND4 (N715, N699, N692, N287, N468);
xor XOR2 (N716, N701, N407);
nand NAND2 (N717, N706, N705);
buf BUF1 (N718, N717);
nor NOR2 (N719, N718, N349);
or OR4 (N720, N713, N602, N569, N470);
or OR2 (N721, N719, N698);
or OR4 (N722, N715, N152, N303, N274);
or OR3 (N723, N712, N280, N165);
nor NOR3 (N724, N723, N261, N395);
not NOT1 (N725, N720);
and AND4 (N726, N722, N401, N535, N647);
xor XOR2 (N727, N724, N85);
nand NAND3 (N728, N721, N141, N11);
or OR4 (N729, N727, N252, N263, N644);
buf BUF1 (N730, N714);
not NOT1 (N731, N729);
and AND4 (N732, N660, N635, N390, N380);
and AND2 (N733, N674, N636);
and AND2 (N734, N731, N89);
not NOT1 (N735, N734);
not NOT1 (N736, N725);
xor XOR2 (N737, N730, N247);
or OR2 (N738, N735, N571);
nor NOR3 (N739, N728, N297, N656);
xor XOR2 (N740, N737, N275);
or OR2 (N741, N711, N529);
xor XOR2 (N742, N738, N586);
and AND3 (N743, N726, N308, N12);
not NOT1 (N744, N742);
nor NOR2 (N745, N736, N44);
nand NAND3 (N746, N739, N375, N430);
nor NOR4 (N747, N746, N152, N536, N195);
xor XOR2 (N748, N744, N140);
not NOT1 (N749, N733);
not NOT1 (N750, N743);
not NOT1 (N751, N748);
or OR4 (N752, N750, N174, N258, N600);
buf BUF1 (N753, N703);
not NOT1 (N754, N753);
not NOT1 (N755, N749);
nor NOR3 (N756, N752, N237, N160);
xor XOR2 (N757, N745, N218);
not NOT1 (N758, N747);
not NOT1 (N759, N751);
nand NAND2 (N760, N716, N737);
xor XOR2 (N761, N758, N309);
and AND2 (N762, N732, N569);
nand NAND4 (N763, N762, N253, N635, N364);
nor NOR2 (N764, N757, N63);
buf BUF1 (N765, N764);
xor XOR2 (N766, N754, N187);
nor NOR4 (N767, N740, N162, N456, N93);
nor NOR3 (N768, N756, N14, N401);
nand NAND3 (N769, N759, N182, N211);
nand NAND3 (N770, N741, N192, N652);
nand NAND4 (N771, N768, N680, N622, N489);
not NOT1 (N772, N769);
not NOT1 (N773, N755);
and AND4 (N774, N772, N586, N132, N64);
or OR4 (N775, N761, N188, N476, N659);
and AND3 (N776, N766, N690, N132);
nand NAND2 (N777, N771, N79);
nor NOR3 (N778, N763, N769, N761);
not NOT1 (N779, N760);
nor NOR2 (N780, N775, N2);
nand NAND2 (N781, N779, N536);
buf BUF1 (N782, N781);
or OR2 (N783, N767, N411);
or OR2 (N784, N780, N163);
and AND3 (N785, N777, N45, N154);
and AND4 (N786, N774, N691, N423, N388);
and AND2 (N787, N786, N535);
not NOT1 (N788, N770);
nand NAND4 (N789, N776, N239, N546, N193);
xor XOR2 (N790, N783, N566);
xor XOR2 (N791, N765, N173);
not NOT1 (N792, N787);
and AND2 (N793, N792, N225);
buf BUF1 (N794, N784);
or OR4 (N795, N778, N257, N296, N162);
nand NAND3 (N796, N794, N648, N657);
not NOT1 (N797, N791);
or OR3 (N798, N793, N302, N461);
or OR4 (N799, N788, N385, N388, N246);
not NOT1 (N800, N799);
or OR2 (N801, N789, N793);
xor XOR2 (N802, N790, N257);
not NOT1 (N803, N801);
nor NOR3 (N804, N798, N195, N399);
nand NAND2 (N805, N796, N91);
not NOT1 (N806, N800);
nor NOR2 (N807, N797, N789);
nor NOR3 (N808, N795, N771, N574);
and AND2 (N809, N773, N711);
or OR4 (N810, N809, N748, N179, N128);
xor XOR2 (N811, N808, N497);
buf BUF1 (N812, N802);
xor XOR2 (N813, N803, N92);
or OR2 (N814, N807, N186);
or OR4 (N815, N806, N39, N727, N110);
nor NOR2 (N816, N810, N476);
or OR3 (N817, N782, N743, N642);
buf BUF1 (N818, N812);
nor NOR2 (N819, N815, N602);
nand NAND2 (N820, N805, N3);
buf BUF1 (N821, N813);
or OR2 (N822, N821, N806);
nand NAND4 (N823, N814, N466, N703, N462);
and AND4 (N824, N820, N762, N488, N778);
buf BUF1 (N825, N819);
and AND4 (N826, N817, N809, N390, N546);
and AND2 (N827, N825, N517);
buf BUF1 (N828, N827);
buf BUF1 (N829, N823);
xor XOR2 (N830, N785, N790);
nand NAND2 (N831, N830, N65);
not NOT1 (N832, N829);
or OR3 (N833, N818, N141, N61);
xor XOR2 (N834, N832, N721);
nand NAND4 (N835, N828, N316, N269, N432);
and AND4 (N836, N822, N285, N97, N369);
xor XOR2 (N837, N824, N71);
xor XOR2 (N838, N833, N650);
not NOT1 (N839, N835);
nand NAND4 (N840, N837, N380, N139, N100);
and AND2 (N841, N811, N558);
buf BUF1 (N842, N841);
or OR4 (N843, N840, N766, N554, N562);
buf BUF1 (N844, N843);
buf BUF1 (N845, N816);
and AND3 (N846, N838, N352, N225);
nor NOR3 (N847, N844, N370, N269);
not NOT1 (N848, N834);
and AND4 (N849, N836, N653, N485, N118);
buf BUF1 (N850, N848);
xor XOR2 (N851, N804, N233);
xor XOR2 (N852, N831, N722);
xor XOR2 (N853, N826, N709);
buf BUF1 (N854, N839);
buf BUF1 (N855, N846);
not NOT1 (N856, N845);
buf BUF1 (N857, N849);
nand NAND4 (N858, N855, N319, N733, N195);
not NOT1 (N859, N851);
nand NAND4 (N860, N852, N808, N357, N409);
nand NAND3 (N861, N859, N674, N805);
not NOT1 (N862, N847);
or OR4 (N863, N860, N838, N338, N772);
xor XOR2 (N864, N863, N536);
buf BUF1 (N865, N856);
buf BUF1 (N866, N864);
xor XOR2 (N867, N866, N666);
xor XOR2 (N868, N842, N693);
and AND3 (N869, N853, N339, N124);
nand NAND4 (N870, N865, N173, N238, N342);
xor XOR2 (N871, N867, N412);
xor XOR2 (N872, N857, N179);
and AND3 (N873, N871, N190, N66);
and AND2 (N874, N870, N848);
nor NOR3 (N875, N862, N591, N826);
xor XOR2 (N876, N872, N62);
nand NAND2 (N877, N869, N713);
nand NAND4 (N878, N858, N141, N746, N595);
buf BUF1 (N879, N850);
buf BUF1 (N880, N873);
xor XOR2 (N881, N861, N182);
and AND2 (N882, N875, N632);
or OR2 (N883, N854, N867);
and AND4 (N884, N876, N702, N772, N869);
or OR3 (N885, N878, N732, N516);
xor XOR2 (N886, N882, N675);
and AND3 (N887, N884, N527, N855);
nor NOR3 (N888, N881, N725, N752);
nand NAND2 (N889, N883, N866);
xor XOR2 (N890, N888, N144);
nand NAND4 (N891, N886, N519, N443, N268);
nand NAND4 (N892, N889, N777, N563, N840);
or OR3 (N893, N879, N874, N3);
and AND2 (N894, N684, N613);
or OR2 (N895, N894, N235);
nor NOR4 (N896, N895, N569, N573, N266);
not NOT1 (N897, N877);
buf BUF1 (N898, N892);
and AND2 (N899, N897, N875);
buf BUF1 (N900, N885);
xor XOR2 (N901, N900, N705);
nand NAND4 (N902, N868, N354, N518, N631);
xor XOR2 (N903, N898, N444);
nand NAND2 (N904, N899, N760);
nor NOR2 (N905, N887, N607);
and AND3 (N906, N891, N303, N6);
nand NAND4 (N907, N903, N573, N97, N634);
nand NAND4 (N908, N880, N394, N543, N517);
or OR3 (N909, N896, N729, N353);
not NOT1 (N910, N904);
not NOT1 (N911, N907);
and AND4 (N912, N911, N352, N206, N3);
or OR4 (N913, N893, N543, N500, N146);
nand NAND2 (N914, N901, N555);
or OR3 (N915, N912, N14, N157);
nand NAND4 (N916, N915, N323, N816, N882);
xor XOR2 (N917, N908, N41);
or OR4 (N918, N906, N705, N296, N397);
buf BUF1 (N919, N918);
xor XOR2 (N920, N917, N796);
or OR3 (N921, N902, N60, N729);
not NOT1 (N922, N913);
xor XOR2 (N923, N921, N51);
and AND2 (N924, N910, N301);
buf BUF1 (N925, N922);
and AND2 (N926, N924, N731);
xor XOR2 (N927, N926, N226);
or OR2 (N928, N925, N110);
not NOT1 (N929, N923);
nor NOR2 (N930, N916, N892);
not NOT1 (N931, N930);
not NOT1 (N932, N919);
buf BUF1 (N933, N928);
or OR2 (N934, N929, N177);
nand NAND2 (N935, N909, N306);
xor XOR2 (N936, N890, N692);
buf BUF1 (N937, N905);
xor XOR2 (N938, N914, N774);
or OR3 (N939, N932, N698, N162);
and AND4 (N940, N931, N427, N206, N132);
nand NAND2 (N941, N920, N911);
nand NAND2 (N942, N927, N785);
or OR4 (N943, N935, N841, N933, N124);
xor XOR2 (N944, N410, N730);
nor NOR3 (N945, N944, N630, N700);
xor XOR2 (N946, N943, N884);
and AND3 (N947, N942, N777, N602);
nand NAND2 (N948, N938, N938);
buf BUF1 (N949, N939);
and AND3 (N950, N948, N186, N127);
and AND2 (N951, N934, N845);
buf BUF1 (N952, N951);
buf BUF1 (N953, N941);
nor NOR3 (N954, N949, N710, N89);
xor XOR2 (N955, N950, N279);
nand NAND2 (N956, N946, N396);
buf BUF1 (N957, N955);
nand NAND2 (N958, N947, N168);
and AND2 (N959, N956, N420);
and AND2 (N960, N957, N355);
nand NAND4 (N961, N936, N129, N259, N924);
buf BUF1 (N962, N952);
nor NOR3 (N963, N940, N87, N277);
not NOT1 (N964, N954);
nor NOR3 (N965, N937, N404, N45);
or OR3 (N966, N960, N562, N940);
or OR3 (N967, N964, N682, N741);
nor NOR3 (N968, N959, N330, N304);
nand NAND4 (N969, N967, N721, N667, N767);
buf BUF1 (N970, N969);
buf BUF1 (N971, N945);
buf BUF1 (N972, N970);
or OR4 (N973, N958, N451, N838, N219);
not NOT1 (N974, N953);
or OR2 (N975, N965, N633);
not NOT1 (N976, N966);
or OR2 (N977, N973, N816);
nor NOR4 (N978, N961, N668, N410, N465);
nor NOR2 (N979, N963, N45);
buf BUF1 (N980, N975);
or OR4 (N981, N972, N592, N150, N583);
and AND4 (N982, N971, N424, N75, N849);
and AND3 (N983, N979, N611, N177);
nor NOR2 (N984, N977, N76);
xor XOR2 (N985, N980, N939);
nor NOR2 (N986, N982, N207);
xor XOR2 (N987, N986, N257);
buf BUF1 (N988, N962);
nand NAND3 (N989, N987, N694, N845);
buf BUF1 (N990, N984);
xor XOR2 (N991, N988, N841);
and AND2 (N992, N985, N800);
buf BUF1 (N993, N992);
not NOT1 (N994, N989);
buf BUF1 (N995, N983);
and AND3 (N996, N976, N760, N379);
or OR3 (N997, N978, N348, N9);
nor NOR2 (N998, N995, N250);
nand NAND4 (N999, N974, N294, N926, N783);
and AND4 (N1000, N981, N884, N638, N542);
nor NOR2 (N1001, N990, N577);
nand NAND3 (N1002, N993, N920, N937);
xor XOR2 (N1003, N1002, N588);
buf BUF1 (N1004, N1003);
xor XOR2 (N1005, N1001, N422);
nor NOR2 (N1006, N991, N9);
nor NOR2 (N1007, N1006, N215);
or OR2 (N1008, N1007, N540);
buf BUF1 (N1009, N994);
and AND2 (N1010, N1004, N920);
not NOT1 (N1011, N996);
nor NOR3 (N1012, N1009, N337, N247);
xor XOR2 (N1013, N997, N547);
xor XOR2 (N1014, N1005, N437);
nand NAND2 (N1015, N1011, N100);
and AND2 (N1016, N1010, N197);
xor XOR2 (N1017, N968, N440);
buf BUF1 (N1018, N1008);
xor XOR2 (N1019, N1016, N908);
nand NAND2 (N1020, N1018, N874);
not NOT1 (N1021, N999);
or OR2 (N1022, N1012, N802);
nand NAND4 (N1023, N1015, N32, N376, N936);
not NOT1 (N1024, N1017);
nand NAND3 (N1025, N1022, N132, N236);
xor XOR2 (N1026, N1014, N77);
not NOT1 (N1027, N1024);
xor XOR2 (N1028, N1020, N716);
and AND4 (N1029, N1026, N714, N712, N288);
xor XOR2 (N1030, N1029, N387);
buf BUF1 (N1031, N1025);
not NOT1 (N1032, N1021);
xor XOR2 (N1033, N1030, N812);
and AND4 (N1034, N1023, N320, N148, N430);
xor XOR2 (N1035, N1027, N958);
nand NAND3 (N1036, N1019, N732, N684);
nor NOR4 (N1037, N1013, N181, N871, N475);
nand NAND3 (N1038, N1034, N513, N463);
and AND3 (N1039, N1036, N890, N170);
not NOT1 (N1040, N1039);
or OR2 (N1041, N1032, N180);
not NOT1 (N1042, N1028);
buf BUF1 (N1043, N1037);
not NOT1 (N1044, N1042);
buf BUF1 (N1045, N1044);
and AND2 (N1046, N1031, N662);
not NOT1 (N1047, N998);
nor NOR2 (N1048, N1047, N893);
xor XOR2 (N1049, N1040, N708);
or OR3 (N1050, N1041, N31, N807);
nand NAND2 (N1051, N1046, N917);
nand NAND2 (N1052, N1000, N427);
buf BUF1 (N1053, N1045);
nor NOR3 (N1054, N1038, N35, N880);
and AND3 (N1055, N1043, N1022, N734);
nor NOR2 (N1056, N1051, N339);
or OR4 (N1057, N1052, N418, N292, N179);
nand NAND3 (N1058, N1049, N404, N828);
xor XOR2 (N1059, N1058, N1046);
or OR4 (N1060, N1048, N159, N108, N546);
nand NAND4 (N1061, N1057, N588, N599, N722);
nand NAND2 (N1062, N1033, N168);
or OR3 (N1063, N1059, N563, N69);
buf BUF1 (N1064, N1054);
xor XOR2 (N1065, N1053, N1058);
and AND2 (N1066, N1060, N399);
or OR3 (N1067, N1065, N244, N1030);
or OR4 (N1068, N1064, N492, N990, N572);
not NOT1 (N1069, N1061);
or OR4 (N1070, N1035, N407, N1063, N343);
nand NAND3 (N1071, N763, N624, N841);
not NOT1 (N1072, N1056);
nand NAND3 (N1073, N1055, N601, N275);
nor NOR3 (N1074, N1067, N778, N908);
nand NAND4 (N1075, N1068, N412, N853, N407);
or OR2 (N1076, N1070, N791);
or OR4 (N1077, N1062, N659, N808, N486);
or OR4 (N1078, N1075, N1010, N863, N482);
nor NOR3 (N1079, N1073, N563, N456);
nor NOR2 (N1080, N1079, N26);
or OR2 (N1081, N1066, N258);
not NOT1 (N1082, N1050);
xor XOR2 (N1083, N1072, N402);
and AND3 (N1084, N1077, N117, N376);
not NOT1 (N1085, N1069);
or OR2 (N1086, N1084, N850);
and AND3 (N1087, N1080, N168, N235);
buf BUF1 (N1088, N1071);
xor XOR2 (N1089, N1082, N268);
xor XOR2 (N1090, N1085, N508);
not NOT1 (N1091, N1090);
and AND4 (N1092, N1087, N446, N930, N517);
nand NAND4 (N1093, N1083, N389, N985, N619);
buf BUF1 (N1094, N1086);
and AND2 (N1095, N1094, N9);
and AND4 (N1096, N1074, N148, N918, N254);
and AND4 (N1097, N1096, N667, N909, N985);
and AND2 (N1098, N1081, N1090);
buf BUF1 (N1099, N1093);
not NOT1 (N1100, N1097);
xor XOR2 (N1101, N1100, N730);
xor XOR2 (N1102, N1101, N1085);
xor XOR2 (N1103, N1088, N438);
not NOT1 (N1104, N1092);
and AND3 (N1105, N1095, N1035, N746);
and AND2 (N1106, N1089, N394);
nor NOR3 (N1107, N1098, N192, N696);
nand NAND4 (N1108, N1078, N228, N760, N685);
and AND2 (N1109, N1099, N1013);
and AND4 (N1110, N1104, N797, N262, N194);
nand NAND3 (N1111, N1091, N740, N298);
buf BUF1 (N1112, N1111);
buf BUF1 (N1113, N1109);
xor XOR2 (N1114, N1106, N308);
xor XOR2 (N1115, N1076, N118);
xor XOR2 (N1116, N1114, N362);
xor XOR2 (N1117, N1110, N389);
buf BUF1 (N1118, N1107);
and AND2 (N1119, N1102, N135);
xor XOR2 (N1120, N1119, N388);
xor XOR2 (N1121, N1108, N260);
or OR4 (N1122, N1116, N511, N45, N466);
xor XOR2 (N1123, N1120, N138);
buf BUF1 (N1124, N1123);
nand NAND4 (N1125, N1124, N829, N278, N870);
nand NAND2 (N1126, N1113, N145);
nor NOR3 (N1127, N1122, N822, N454);
nor NOR3 (N1128, N1125, N799, N464);
not NOT1 (N1129, N1112);
or OR4 (N1130, N1103, N429, N465, N152);
nor NOR3 (N1131, N1105, N943, N321);
buf BUF1 (N1132, N1131);
nand NAND4 (N1133, N1127, N403, N277, N954);
buf BUF1 (N1134, N1115);
nor NOR3 (N1135, N1134, N1015, N702);
buf BUF1 (N1136, N1121);
nand NAND2 (N1137, N1133, N214);
not NOT1 (N1138, N1118);
and AND4 (N1139, N1138, N593, N122, N646);
and AND4 (N1140, N1135, N387, N736, N597);
not NOT1 (N1141, N1132);
and AND2 (N1142, N1136, N610);
or OR2 (N1143, N1142, N72);
xor XOR2 (N1144, N1139, N485);
buf BUF1 (N1145, N1143);
buf BUF1 (N1146, N1140);
or OR4 (N1147, N1130, N901, N1068, N910);
not NOT1 (N1148, N1146);
buf BUF1 (N1149, N1117);
nand NAND4 (N1150, N1129, N902, N672, N272);
xor XOR2 (N1151, N1141, N355);
or OR4 (N1152, N1149, N1054, N343, N746);
and AND3 (N1153, N1150, N779, N498);
or OR4 (N1154, N1151, N783, N885, N241);
or OR4 (N1155, N1147, N371, N80, N820);
and AND3 (N1156, N1144, N682, N971);
nand NAND4 (N1157, N1154, N710, N801, N878);
and AND4 (N1158, N1145, N87, N890, N353);
nand NAND2 (N1159, N1137, N607);
nand NAND3 (N1160, N1158, N824, N530);
xor XOR2 (N1161, N1156, N918);
nand NAND4 (N1162, N1153, N706, N951, N111);
or OR2 (N1163, N1162, N771);
or OR3 (N1164, N1126, N148, N786);
nor NOR2 (N1165, N1157, N1013);
xor XOR2 (N1166, N1160, N837);
and AND4 (N1167, N1128, N122, N199, N669);
nand NAND2 (N1168, N1164, N163);
buf BUF1 (N1169, N1159);
nand NAND2 (N1170, N1168, N210);
xor XOR2 (N1171, N1148, N370);
xor XOR2 (N1172, N1166, N383);
and AND2 (N1173, N1163, N132);
buf BUF1 (N1174, N1169);
xor XOR2 (N1175, N1165, N997);
or OR4 (N1176, N1170, N542, N687, N847);
nand NAND2 (N1177, N1175, N2);
and AND2 (N1178, N1176, N665);
and AND2 (N1179, N1171, N391);
or OR3 (N1180, N1152, N764, N751);
or OR3 (N1181, N1179, N921, N828);
nand NAND2 (N1182, N1155, N58);
xor XOR2 (N1183, N1174, N1105);
or OR3 (N1184, N1177, N200, N725);
buf BUF1 (N1185, N1180);
buf BUF1 (N1186, N1178);
buf BUF1 (N1187, N1182);
nand NAND4 (N1188, N1173, N904, N179, N1151);
not NOT1 (N1189, N1185);
or OR3 (N1190, N1188, N670, N835);
buf BUF1 (N1191, N1190);
buf BUF1 (N1192, N1184);
nor NOR2 (N1193, N1192, N18);
and AND2 (N1194, N1193, N265);
nor NOR3 (N1195, N1189, N709, N47);
nand NAND4 (N1196, N1167, N803, N887, N466);
or OR2 (N1197, N1186, N952);
nor NOR2 (N1198, N1194, N1098);
xor XOR2 (N1199, N1198, N454);
nor NOR4 (N1200, N1196, N505, N169, N687);
not NOT1 (N1201, N1183);
nor NOR2 (N1202, N1195, N91);
buf BUF1 (N1203, N1187);
not NOT1 (N1204, N1197);
xor XOR2 (N1205, N1200, N265);
buf BUF1 (N1206, N1203);
buf BUF1 (N1207, N1161);
xor XOR2 (N1208, N1205, N360);
and AND3 (N1209, N1201, N968, N260);
nand NAND3 (N1210, N1208, N840, N985);
buf BUF1 (N1211, N1172);
or OR4 (N1212, N1202, N99, N867, N100);
not NOT1 (N1213, N1212);
nand NAND4 (N1214, N1199, N336, N82, N337);
and AND4 (N1215, N1213, N1152, N9, N991);
nand NAND3 (N1216, N1207, N837, N166);
nand NAND4 (N1217, N1210, N1041, N973, N1205);
nor NOR2 (N1218, N1216, N1151);
nor NOR3 (N1219, N1204, N536, N514);
or OR2 (N1220, N1214, N879);
nor NOR2 (N1221, N1215, N444);
xor XOR2 (N1222, N1211, N593);
not NOT1 (N1223, N1209);
nand NAND3 (N1224, N1221, N568, N686);
nor NOR3 (N1225, N1224, N1018, N668);
nand NAND2 (N1226, N1225, N43);
xor XOR2 (N1227, N1219, N674);
xor XOR2 (N1228, N1222, N38);
or OR2 (N1229, N1218, N856);
buf BUF1 (N1230, N1229);
buf BUF1 (N1231, N1206);
xor XOR2 (N1232, N1227, N905);
and AND2 (N1233, N1230, N960);
and AND2 (N1234, N1191, N99);
xor XOR2 (N1235, N1233, N687);
nand NAND4 (N1236, N1226, N861, N452, N200);
xor XOR2 (N1237, N1231, N850);
not NOT1 (N1238, N1234);
not NOT1 (N1239, N1238);
or OR3 (N1240, N1228, N1187, N201);
buf BUF1 (N1241, N1220);
and AND3 (N1242, N1236, N669, N820);
buf BUF1 (N1243, N1242);
and AND3 (N1244, N1181, N1190, N587);
not NOT1 (N1245, N1237);
nand NAND3 (N1246, N1245, N307, N126);
not NOT1 (N1247, N1244);
or OR2 (N1248, N1232, N399);
and AND2 (N1249, N1240, N1101);
not NOT1 (N1250, N1243);
and AND4 (N1251, N1249, N328, N98, N828);
xor XOR2 (N1252, N1223, N680);
not NOT1 (N1253, N1247);
nor NOR3 (N1254, N1246, N1187, N314);
nor NOR2 (N1255, N1253, N161);
nand NAND2 (N1256, N1241, N460);
not NOT1 (N1257, N1255);
nand NAND2 (N1258, N1250, N844);
not NOT1 (N1259, N1254);
and AND2 (N1260, N1239, N928);
not NOT1 (N1261, N1259);
nand NAND2 (N1262, N1252, N718);
xor XOR2 (N1263, N1235, N248);
buf BUF1 (N1264, N1262);
and AND2 (N1265, N1258, N1067);
nand NAND3 (N1266, N1264, N1083, N314);
or OR3 (N1267, N1251, N432, N930);
buf BUF1 (N1268, N1260);
buf BUF1 (N1269, N1217);
or OR2 (N1270, N1267, N590);
nor NOR4 (N1271, N1256, N188, N1152, N1105);
nand NAND3 (N1272, N1248, N30, N1199);
nor NOR3 (N1273, N1269, N436, N102);
not NOT1 (N1274, N1261);
buf BUF1 (N1275, N1272);
or OR2 (N1276, N1263, N1035);
nand NAND2 (N1277, N1271, N448);
xor XOR2 (N1278, N1276, N613);
not NOT1 (N1279, N1274);
xor XOR2 (N1280, N1265, N528);
and AND2 (N1281, N1270, N929);
xor XOR2 (N1282, N1279, N588);
or OR4 (N1283, N1273, N403, N807, N628);
or OR4 (N1284, N1278, N210, N1139, N114);
not NOT1 (N1285, N1257);
xor XOR2 (N1286, N1284, N990);
or OR4 (N1287, N1282, N826, N554, N1128);
xor XOR2 (N1288, N1268, N901);
not NOT1 (N1289, N1288);
xor XOR2 (N1290, N1280, N155);
buf BUF1 (N1291, N1281);
nand NAND3 (N1292, N1291, N37, N856);
nor NOR3 (N1293, N1287, N5, N120);
not NOT1 (N1294, N1277);
xor XOR2 (N1295, N1289, N689);
xor XOR2 (N1296, N1290, N1277);
not NOT1 (N1297, N1286);
nand NAND4 (N1298, N1285, N198, N491, N1088);
not NOT1 (N1299, N1298);
nor NOR4 (N1300, N1296, N281, N243, N555);
buf BUF1 (N1301, N1299);
nor NOR2 (N1302, N1295, N845);
nand NAND4 (N1303, N1297, N1289, N1121, N434);
not NOT1 (N1304, N1294);
or OR3 (N1305, N1301, N645, N231);
or OR4 (N1306, N1293, N228, N600, N524);
and AND4 (N1307, N1300, N81, N1107, N559);
and AND2 (N1308, N1283, N453);
or OR4 (N1309, N1303, N452, N803, N55);
buf BUF1 (N1310, N1308);
or OR4 (N1311, N1310, N67, N632, N1255);
or OR2 (N1312, N1266, N813);
not NOT1 (N1313, N1311);
nand NAND2 (N1314, N1305, N421);
nand NAND2 (N1315, N1309, N808);
or OR4 (N1316, N1312, N1103, N628, N587);
not NOT1 (N1317, N1306);
xor XOR2 (N1318, N1292, N517);
or OR2 (N1319, N1304, N1218);
xor XOR2 (N1320, N1307, N283);
or OR4 (N1321, N1316, N498, N928, N650);
not NOT1 (N1322, N1319);
xor XOR2 (N1323, N1275, N345);
nand NAND3 (N1324, N1313, N1189, N1024);
and AND2 (N1325, N1320, N742);
or OR2 (N1326, N1317, N465);
xor XOR2 (N1327, N1322, N28);
nand NAND3 (N1328, N1325, N76, N115);
not NOT1 (N1329, N1328);
xor XOR2 (N1330, N1314, N1320);
and AND2 (N1331, N1318, N1035);
or OR4 (N1332, N1321, N295, N902, N592);
xor XOR2 (N1333, N1332, N1030);
buf BUF1 (N1334, N1324);
nand NAND4 (N1335, N1327, N703, N167, N1105);
nor NOR3 (N1336, N1335, N922, N475);
nor NOR4 (N1337, N1334, N944, N998, N655);
or OR4 (N1338, N1302, N181, N1033, N404);
nand NAND2 (N1339, N1315, N968);
and AND3 (N1340, N1331, N637, N665);
and AND3 (N1341, N1329, N1292, N845);
and AND3 (N1342, N1333, N1143, N789);
not NOT1 (N1343, N1339);
buf BUF1 (N1344, N1341);
nand NAND4 (N1345, N1340, N566, N637, N857);
nor NOR2 (N1346, N1344, N682);
nand NAND2 (N1347, N1346, N727);
nor NOR4 (N1348, N1330, N1195, N568, N1155);
xor XOR2 (N1349, N1348, N189);
xor XOR2 (N1350, N1345, N138);
nand NAND2 (N1351, N1323, N803);
xor XOR2 (N1352, N1343, N959);
or OR4 (N1353, N1350, N99, N821, N795);
or OR2 (N1354, N1349, N918);
xor XOR2 (N1355, N1336, N931);
or OR4 (N1356, N1354, N714, N1038, N884);
not NOT1 (N1357, N1338);
not NOT1 (N1358, N1337);
nand NAND3 (N1359, N1342, N771, N726);
nand NAND3 (N1360, N1358, N251, N247);
xor XOR2 (N1361, N1353, N756);
and AND2 (N1362, N1359, N531);
xor XOR2 (N1363, N1362, N53);
nand NAND4 (N1364, N1356, N705, N277, N418);
and AND3 (N1365, N1360, N854, N1331);
nand NAND4 (N1366, N1352, N1274, N11, N403);
or OR2 (N1367, N1326, N604);
nor NOR4 (N1368, N1367, N132, N646, N1039);
buf BUF1 (N1369, N1357);
not NOT1 (N1370, N1355);
or OR4 (N1371, N1364, N1068, N1163, N64);
not NOT1 (N1372, N1368);
xor XOR2 (N1373, N1369, N1240);
nand NAND3 (N1374, N1373, N68, N1245);
buf BUF1 (N1375, N1370);
xor XOR2 (N1376, N1365, N275);
not NOT1 (N1377, N1347);
nand NAND3 (N1378, N1361, N610, N1299);
nand NAND3 (N1379, N1376, N80, N118);
buf BUF1 (N1380, N1366);
nor NOR2 (N1381, N1371, N827);
xor XOR2 (N1382, N1351, N1312);
and AND3 (N1383, N1380, N275, N500);
nor NOR3 (N1384, N1363, N449, N91);
and AND3 (N1385, N1384, N1089, N1024);
or OR2 (N1386, N1379, N618);
nand NAND3 (N1387, N1377, N81, N1158);
xor XOR2 (N1388, N1374, N360);
buf BUF1 (N1389, N1383);
not NOT1 (N1390, N1378);
nor NOR3 (N1391, N1389, N1239, N908);
buf BUF1 (N1392, N1388);
xor XOR2 (N1393, N1391, N1218);
buf BUF1 (N1394, N1386);
and AND2 (N1395, N1392, N1281);
buf BUF1 (N1396, N1394);
not NOT1 (N1397, N1375);
or OR4 (N1398, N1381, N1179, N389, N576);
not NOT1 (N1399, N1390);
or OR2 (N1400, N1393, N1384);
nand NAND4 (N1401, N1372, N979, N1363, N170);
or OR4 (N1402, N1382, N1263, N551, N462);
nor NOR2 (N1403, N1385, N873);
xor XOR2 (N1404, N1399, N812);
not NOT1 (N1405, N1398);
nand NAND4 (N1406, N1405, N928, N1090, N1047);
not NOT1 (N1407, N1402);
and AND2 (N1408, N1401, N73);
nand NAND4 (N1409, N1395, N382, N472, N968);
buf BUF1 (N1410, N1400);
nor NOR4 (N1411, N1410, N646, N1243, N82);
nand NAND3 (N1412, N1411, N669, N623);
xor XOR2 (N1413, N1387, N213);
or OR3 (N1414, N1408, N1095, N737);
nand NAND4 (N1415, N1407, N1008, N990, N1208);
or OR4 (N1416, N1415, N910, N1407, N1323);
nand NAND2 (N1417, N1416, N1135);
not NOT1 (N1418, N1406);
or OR4 (N1419, N1417, N341, N702, N49);
and AND4 (N1420, N1409, N1328, N349, N520);
nor NOR2 (N1421, N1414, N766);
or OR3 (N1422, N1420, N233, N1265);
buf BUF1 (N1423, N1422);
and AND3 (N1424, N1418, N1002, N303);
nor NOR2 (N1425, N1419, N214);
nor NOR3 (N1426, N1421, N680, N1383);
or OR2 (N1427, N1404, N691);
buf BUF1 (N1428, N1423);
nor NOR4 (N1429, N1428, N197, N293, N1269);
xor XOR2 (N1430, N1413, N978);
xor XOR2 (N1431, N1396, N524);
xor XOR2 (N1432, N1403, N1065);
not NOT1 (N1433, N1425);
not NOT1 (N1434, N1431);
or OR2 (N1435, N1426, N1097);
not NOT1 (N1436, N1397);
xor XOR2 (N1437, N1432, N946);
buf BUF1 (N1438, N1433);
xor XOR2 (N1439, N1424, N619);
nand NAND2 (N1440, N1430, N898);
not NOT1 (N1441, N1440);
or OR2 (N1442, N1437, N996);
xor XOR2 (N1443, N1427, N242);
nand NAND3 (N1444, N1429, N831, N109);
and AND4 (N1445, N1444, N240, N707, N101);
xor XOR2 (N1446, N1435, N375);
not NOT1 (N1447, N1412);
nor NOR3 (N1448, N1442, N1163, N914);
or OR4 (N1449, N1436, N210, N229, N1430);
and AND3 (N1450, N1443, N917, N1141);
and AND4 (N1451, N1448, N1332, N401, N48);
nor NOR3 (N1452, N1439, N367, N1432);
or OR4 (N1453, N1441, N1192, N503, N1036);
xor XOR2 (N1454, N1449, N2);
buf BUF1 (N1455, N1453);
and AND4 (N1456, N1450, N967, N1055, N856);
nand NAND4 (N1457, N1438, N455, N1071, N423);
or OR4 (N1458, N1454, N498, N868, N126);
nor NOR2 (N1459, N1452, N989);
or OR2 (N1460, N1457, N1064);
xor XOR2 (N1461, N1445, N1094);
nand NAND4 (N1462, N1455, N215, N1136, N1299);
and AND4 (N1463, N1446, N719, N512, N824);
nor NOR4 (N1464, N1458, N855, N104, N1038);
buf BUF1 (N1465, N1434);
and AND4 (N1466, N1464, N851, N839, N725);
not NOT1 (N1467, N1459);
nor NOR2 (N1468, N1456, N1295);
and AND4 (N1469, N1468, N228, N1321, N945);
and AND4 (N1470, N1461, N66, N223, N484);
buf BUF1 (N1471, N1451);
nand NAND4 (N1472, N1466, N424, N704, N36);
nor NOR3 (N1473, N1460, N557, N1237);
or OR4 (N1474, N1447, N477, N340, N15);
or OR4 (N1475, N1473, N795, N904, N214);
nand NAND3 (N1476, N1463, N902, N856);
nand NAND3 (N1477, N1472, N272, N1083);
and AND2 (N1478, N1465, N1244);
or OR2 (N1479, N1471, N1042);
xor XOR2 (N1480, N1462, N635);
nor NOR4 (N1481, N1479, N971, N44, N1190);
nand NAND2 (N1482, N1478, N1183);
not NOT1 (N1483, N1475);
nor NOR4 (N1484, N1482, N55, N1110, N394);
nand NAND3 (N1485, N1470, N33, N811);
xor XOR2 (N1486, N1485, N122);
nand NAND4 (N1487, N1480, N63, N211, N1261);
or OR3 (N1488, N1487, N1262, N652);
and AND2 (N1489, N1484, N12);
buf BUF1 (N1490, N1489);
and AND2 (N1491, N1490, N148);
not NOT1 (N1492, N1488);
and AND4 (N1493, N1477, N132, N68, N134);
buf BUF1 (N1494, N1483);
xor XOR2 (N1495, N1494, N850);
and AND2 (N1496, N1481, N659);
xor XOR2 (N1497, N1467, N540);
and AND2 (N1498, N1491, N167);
and AND4 (N1499, N1495, N59, N1094, N910);
buf BUF1 (N1500, N1469);
and AND3 (N1501, N1493, N1275, N449);
buf BUF1 (N1502, N1501);
and AND2 (N1503, N1498, N24);
and AND4 (N1504, N1502, N1116, N690, N1444);
nor NOR2 (N1505, N1500, N208);
xor XOR2 (N1506, N1505, N1142);
and AND2 (N1507, N1496, N5);
or OR4 (N1508, N1506, N1129, N557, N274);
or OR3 (N1509, N1499, N1008, N232);
not NOT1 (N1510, N1486);
xor XOR2 (N1511, N1503, N1441);
buf BUF1 (N1512, N1492);
not NOT1 (N1513, N1508);
or OR4 (N1514, N1474, N225, N152, N413);
and AND4 (N1515, N1511, N400, N33, N224);
not NOT1 (N1516, N1507);
nor NOR2 (N1517, N1509, N1040);
not NOT1 (N1518, N1510);
nor NOR4 (N1519, N1515, N1161, N177, N210);
not NOT1 (N1520, N1518);
or OR4 (N1521, N1512, N1290, N631, N168);
xor XOR2 (N1522, N1517, N1438);
xor XOR2 (N1523, N1497, N315);
nand NAND2 (N1524, N1520, N1055);
xor XOR2 (N1525, N1524, N1272);
and AND3 (N1526, N1476, N522, N10);
nor NOR2 (N1527, N1514, N706);
and AND4 (N1528, N1522, N1260, N353, N807);
not NOT1 (N1529, N1513);
xor XOR2 (N1530, N1521, N105);
xor XOR2 (N1531, N1516, N307);
nor NOR2 (N1532, N1519, N1360);
buf BUF1 (N1533, N1526);
xor XOR2 (N1534, N1532, N418);
and AND3 (N1535, N1534, N1094, N1309);
xor XOR2 (N1536, N1531, N336);
and AND2 (N1537, N1533, N718);
nand NAND3 (N1538, N1528, N804, N1268);
and AND2 (N1539, N1530, N1080);
not NOT1 (N1540, N1527);
xor XOR2 (N1541, N1537, N1178);
not NOT1 (N1542, N1541);
buf BUF1 (N1543, N1536);
nand NAND4 (N1544, N1543, N597, N278, N833);
and AND3 (N1545, N1538, N1096, N523);
nor NOR4 (N1546, N1523, N566, N1485, N1531);
or OR3 (N1547, N1540, N84, N1409);
nand NAND4 (N1548, N1545, N902, N654, N306);
buf BUF1 (N1549, N1539);
and AND4 (N1550, N1542, N318, N578, N920);
nor NOR2 (N1551, N1550, N904);
and AND3 (N1552, N1547, N39, N1141);
nand NAND2 (N1553, N1546, N1483);
xor XOR2 (N1554, N1535, N871);
buf BUF1 (N1555, N1551);
buf BUF1 (N1556, N1553);
or OR3 (N1557, N1555, N318, N1263);
and AND3 (N1558, N1504, N1088, N614);
buf BUF1 (N1559, N1556);
not NOT1 (N1560, N1549);
nand NAND4 (N1561, N1529, N832, N892, N496);
and AND3 (N1562, N1561, N177, N1217);
nand NAND4 (N1563, N1562, N894, N1365, N163);
buf BUF1 (N1564, N1560);
nand NAND3 (N1565, N1559, N131, N117);
nor NOR4 (N1566, N1548, N372, N709, N373);
not NOT1 (N1567, N1558);
xor XOR2 (N1568, N1552, N430);
not NOT1 (N1569, N1564);
nand NAND4 (N1570, N1566, N1078, N219, N322);
xor XOR2 (N1571, N1565, N522);
and AND4 (N1572, N1563, N191, N1290, N1146);
buf BUF1 (N1573, N1557);
not NOT1 (N1574, N1544);
nor NOR3 (N1575, N1572, N44, N82);
and AND3 (N1576, N1554, N672, N258);
and AND3 (N1577, N1525, N130, N468);
nand NAND2 (N1578, N1574, N613);
not NOT1 (N1579, N1576);
or OR2 (N1580, N1579, N853);
or OR2 (N1581, N1578, N994);
and AND3 (N1582, N1573, N371, N514);
and AND4 (N1583, N1582, N123, N239, N1196);
or OR3 (N1584, N1581, N53, N5);
xor XOR2 (N1585, N1580, N20);
or OR2 (N1586, N1568, N656);
nand NAND3 (N1587, N1570, N1391, N692);
or OR2 (N1588, N1577, N361);
buf BUF1 (N1589, N1571);
or OR3 (N1590, N1575, N658, N213);
or OR3 (N1591, N1567, N757, N447);
or OR3 (N1592, N1587, N381, N323);
xor XOR2 (N1593, N1592, N96);
or OR4 (N1594, N1584, N1370, N1593, N1168);
nor NOR4 (N1595, N920, N671, N507, N1410);
nand NAND2 (N1596, N1595, N339);
not NOT1 (N1597, N1569);
or OR3 (N1598, N1597, N1243, N1537);
nor NOR2 (N1599, N1586, N6);
and AND4 (N1600, N1598, N579, N986, N1173);
nand NAND2 (N1601, N1599, N905);
buf BUF1 (N1602, N1601);
or OR4 (N1603, N1600, N960, N874, N1365);
xor XOR2 (N1604, N1594, N1135);
xor XOR2 (N1605, N1603, N986);
nand NAND2 (N1606, N1590, N297);
nor NOR4 (N1607, N1585, N1376, N277, N799);
nor NOR3 (N1608, N1583, N490, N81);
nand NAND2 (N1609, N1588, N258);
nand NAND2 (N1610, N1606, N1308);
nand NAND3 (N1611, N1591, N761, N1290);
nor NOR2 (N1612, N1602, N712);
nor NOR4 (N1613, N1607, N1336, N1258, N194);
and AND2 (N1614, N1611, N1388);
and AND4 (N1615, N1608, N1036, N773, N1148);
not NOT1 (N1616, N1604);
nand NAND4 (N1617, N1596, N172, N169, N114);
buf BUF1 (N1618, N1614);
not NOT1 (N1619, N1617);
and AND3 (N1620, N1613, N13, N947);
or OR2 (N1621, N1589, N1169);
xor XOR2 (N1622, N1621, N1364);
nand NAND4 (N1623, N1622, N810, N509, N1368);
and AND2 (N1624, N1609, N1500);
nor NOR2 (N1625, N1619, N1058);
nand NAND4 (N1626, N1605, N254, N1398, N848);
or OR3 (N1627, N1615, N1258, N1296);
and AND3 (N1628, N1620, N16, N685);
nor NOR3 (N1629, N1623, N1178, N376);
buf BUF1 (N1630, N1610);
not NOT1 (N1631, N1616);
not NOT1 (N1632, N1627);
buf BUF1 (N1633, N1618);
and AND2 (N1634, N1628, N345);
not NOT1 (N1635, N1631);
nor NOR3 (N1636, N1625, N854, N96);
and AND4 (N1637, N1624, N291, N1526, N1092);
nand NAND2 (N1638, N1634, N912);
xor XOR2 (N1639, N1612, N351);
and AND3 (N1640, N1636, N1629, N4);
not NOT1 (N1641, N1013);
buf BUF1 (N1642, N1637);
nor NOR2 (N1643, N1635, N1370);
nand NAND3 (N1644, N1639, N1524, N595);
nor NOR4 (N1645, N1626, N1049, N819, N83);
xor XOR2 (N1646, N1641, N788);
buf BUF1 (N1647, N1642);
nor NOR2 (N1648, N1646, N1081);
nor NOR3 (N1649, N1643, N208, N1155);
and AND2 (N1650, N1644, N1644);
or OR4 (N1651, N1633, N647, N737, N596);
buf BUF1 (N1652, N1632);
nand NAND4 (N1653, N1647, N100, N745, N778);
or OR3 (N1654, N1651, N853, N1176);
and AND4 (N1655, N1638, N1132, N1120, N1255);
not NOT1 (N1656, N1650);
and AND2 (N1657, N1656, N1577);
or OR2 (N1658, N1640, N82);
nor NOR4 (N1659, N1652, N946, N527, N730);
buf BUF1 (N1660, N1648);
xor XOR2 (N1661, N1660, N1345);
buf BUF1 (N1662, N1649);
nor NOR4 (N1663, N1630, N1177, N381, N593);
xor XOR2 (N1664, N1645, N73);
xor XOR2 (N1665, N1664, N874);
buf BUF1 (N1666, N1655);
and AND3 (N1667, N1657, N236, N405);
buf BUF1 (N1668, N1666);
and AND4 (N1669, N1662, N202, N113, N1506);
nor NOR4 (N1670, N1654, N1065, N1466, N12);
nor NOR2 (N1671, N1665, N1035);
xor XOR2 (N1672, N1661, N741);
or OR4 (N1673, N1670, N385, N493, N504);
and AND2 (N1674, N1668, N319);
or OR4 (N1675, N1669, N556, N1172, N1433);
and AND3 (N1676, N1663, N1470, N769);
nor NOR3 (N1677, N1659, N1540, N867);
not NOT1 (N1678, N1653);
buf BUF1 (N1679, N1658);
nand NAND4 (N1680, N1674, N1525, N1600, N1360);
or OR4 (N1681, N1676, N59, N1526, N772);
xor XOR2 (N1682, N1680, N1411);
and AND4 (N1683, N1681, N1181, N29, N778);
xor XOR2 (N1684, N1679, N1031);
nor NOR4 (N1685, N1677, N1013, N246, N429);
nand NAND3 (N1686, N1675, N783, N306);
nor NOR3 (N1687, N1667, N316, N1660);
nor NOR2 (N1688, N1672, N611);
or OR3 (N1689, N1683, N1573, N1174);
and AND3 (N1690, N1684, N936, N827);
and AND4 (N1691, N1671, N1312, N1053, N1007);
buf BUF1 (N1692, N1690);
or OR4 (N1693, N1682, N1289, N474, N1282);
nor NOR3 (N1694, N1678, N190, N1108);
and AND4 (N1695, N1691, N1303, N631, N1626);
not NOT1 (N1696, N1687);
xor XOR2 (N1697, N1693, N662);
xor XOR2 (N1698, N1692, N1168);
and AND2 (N1699, N1696, N327);
or OR3 (N1700, N1698, N1278, N922);
xor XOR2 (N1701, N1697, N487);
xor XOR2 (N1702, N1699, N1389);
or OR3 (N1703, N1701, N365, N1689);
nor NOR2 (N1704, N1234, N1378);
nor NOR4 (N1705, N1694, N1373, N896, N1515);
nor NOR2 (N1706, N1704, N1673);
nand NAND2 (N1707, N615, N1585);
nand NAND2 (N1708, N1686, N374);
nand NAND4 (N1709, N1685, N531, N342, N803);
buf BUF1 (N1710, N1706);
xor XOR2 (N1711, N1700, N220);
nand NAND3 (N1712, N1711, N73, N699);
and AND4 (N1713, N1709, N652, N787, N1056);
xor XOR2 (N1714, N1702, N145);
buf BUF1 (N1715, N1710);
and AND2 (N1716, N1714, N4);
and AND4 (N1717, N1713, N1297, N411, N979);
not NOT1 (N1718, N1717);
buf BUF1 (N1719, N1718);
and AND2 (N1720, N1705, N1705);
xor XOR2 (N1721, N1688, N790);
nand NAND4 (N1722, N1719, N1468, N851, N1117);
nand NAND2 (N1723, N1703, N1442);
not NOT1 (N1724, N1712);
nand NAND2 (N1725, N1716, N1456);
nor NOR3 (N1726, N1723, N120, N1684);
xor XOR2 (N1727, N1722, N1725);
buf BUF1 (N1728, N741);
not NOT1 (N1729, N1721);
and AND4 (N1730, N1715, N739, N1159, N221);
and AND2 (N1731, N1728, N1162);
xor XOR2 (N1732, N1720, N934);
nor NOR2 (N1733, N1731, N18);
nor NOR3 (N1734, N1729, N561, N506);
and AND3 (N1735, N1730, N101, N10);
or OR3 (N1736, N1734, N1470, N1107);
buf BUF1 (N1737, N1695);
or OR3 (N1738, N1707, N1459, N1236);
nor NOR2 (N1739, N1727, N343);
nor NOR2 (N1740, N1724, N558);
xor XOR2 (N1741, N1726, N1212);
nand NAND2 (N1742, N1740, N1402);
buf BUF1 (N1743, N1733);
nor NOR3 (N1744, N1743, N953, N1027);
buf BUF1 (N1745, N1736);
and AND4 (N1746, N1735, N917, N100, N1523);
not NOT1 (N1747, N1739);
nand NAND3 (N1748, N1747, N73, N491);
or OR2 (N1749, N1741, N236);
and AND3 (N1750, N1742, N1189, N806);
and AND4 (N1751, N1744, N613, N199, N866);
or OR2 (N1752, N1738, N999);
nand NAND4 (N1753, N1746, N1055, N276, N779);
not NOT1 (N1754, N1708);
nand NAND2 (N1755, N1732, N990);
xor XOR2 (N1756, N1752, N175);
buf BUF1 (N1757, N1737);
buf BUF1 (N1758, N1756);
buf BUF1 (N1759, N1758);
and AND4 (N1760, N1750, N307, N1182, N747);
and AND4 (N1761, N1753, N282, N853, N118);
nand NAND2 (N1762, N1759, N1415);
not NOT1 (N1763, N1754);
not NOT1 (N1764, N1760);
not NOT1 (N1765, N1745);
not NOT1 (N1766, N1757);
nor NOR4 (N1767, N1764, N1354, N1238, N1062);
buf BUF1 (N1768, N1751);
xor XOR2 (N1769, N1763, N671);
and AND2 (N1770, N1768, N195);
or OR2 (N1771, N1765, N1070);
and AND4 (N1772, N1770, N1700, N1190, N1014);
and AND3 (N1773, N1749, N726, N1491);
nor NOR2 (N1774, N1773, N161);
buf BUF1 (N1775, N1769);
xor XOR2 (N1776, N1755, N392);
buf BUF1 (N1777, N1774);
nand NAND2 (N1778, N1762, N1600);
buf BUF1 (N1779, N1761);
and AND2 (N1780, N1777, N766);
not NOT1 (N1781, N1748);
and AND2 (N1782, N1780, N1444);
buf BUF1 (N1783, N1771);
or OR3 (N1784, N1775, N1020, N712);
or OR4 (N1785, N1778, N487, N1733, N1322);
nor NOR4 (N1786, N1776, N1590, N717, N363);
xor XOR2 (N1787, N1781, N92);
nor NOR4 (N1788, N1767, N627, N1127, N1105);
not NOT1 (N1789, N1783);
xor XOR2 (N1790, N1784, N783);
nand NAND4 (N1791, N1786, N101, N1319, N1162);
nor NOR2 (N1792, N1791, N965);
or OR3 (N1793, N1792, N1679, N1724);
xor XOR2 (N1794, N1790, N787);
or OR4 (N1795, N1772, N844, N47, N1475);
buf BUF1 (N1796, N1789);
nor NOR4 (N1797, N1793, N1088, N325, N188);
and AND3 (N1798, N1796, N1388, N78);
not NOT1 (N1799, N1798);
buf BUF1 (N1800, N1787);
nor NOR2 (N1801, N1785, N954);
nand NAND2 (N1802, N1782, N358);
or OR4 (N1803, N1766, N590, N573, N944);
nor NOR3 (N1804, N1801, N917, N1772);
or OR2 (N1805, N1804, N592);
xor XOR2 (N1806, N1799, N1055);
or OR3 (N1807, N1803, N1566, N164);
and AND2 (N1808, N1800, N999);
not NOT1 (N1809, N1788);
nor NOR4 (N1810, N1808, N253, N1195, N43);
nand NAND2 (N1811, N1807, N1782);
or OR3 (N1812, N1794, N37, N1809);
or OR2 (N1813, N635, N1634);
not NOT1 (N1814, N1812);
nand NAND2 (N1815, N1805, N1562);
buf BUF1 (N1816, N1795);
xor XOR2 (N1817, N1802, N1164);
nand NAND4 (N1818, N1813, N341, N1780, N1308);
nand NAND4 (N1819, N1815, N1801, N1596, N106);
and AND4 (N1820, N1810, N418, N1721, N508);
buf BUF1 (N1821, N1818);
and AND2 (N1822, N1817, N252);
buf BUF1 (N1823, N1806);
xor XOR2 (N1824, N1819, N1258);
nand NAND2 (N1825, N1822, N1612);
nor NOR3 (N1826, N1814, N1115, N786);
nor NOR2 (N1827, N1824, N1598);
nor NOR4 (N1828, N1823, N859, N163, N446);
xor XOR2 (N1829, N1820, N62);
nor NOR2 (N1830, N1779, N1144);
or OR4 (N1831, N1816, N136, N252, N349);
xor XOR2 (N1832, N1829, N1377);
nand NAND2 (N1833, N1811, N921);
or OR4 (N1834, N1833, N696, N76, N1130);
xor XOR2 (N1835, N1830, N1123);
not NOT1 (N1836, N1835);
nand NAND3 (N1837, N1834, N1655, N1103);
nand NAND3 (N1838, N1837, N991, N89);
nand NAND4 (N1839, N1831, N924, N239, N1336);
or OR3 (N1840, N1832, N1452, N875);
nor NOR4 (N1841, N1840, N1710, N1458, N1335);
nor NOR2 (N1842, N1827, N1457);
nor NOR3 (N1843, N1836, N660, N1461);
xor XOR2 (N1844, N1825, N892);
nor NOR3 (N1845, N1838, N407, N1289);
nor NOR4 (N1846, N1844, N1811, N805, N1637);
and AND3 (N1847, N1821, N800, N1096);
xor XOR2 (N1848, N1826, N31);
or OR2 (N1849, N1797, N1702);
nand NAND2 (N1850, N1846, N2);
xor XOR2 (N1851, N1843, N330);
buf BUF1 (N1852, N1849);
buf BUF1 (N1853, N1842);
and AND4 (N1854, N1853, N92, N746, N570);
nand NAND2 (N1855, N1848, N1675);
or OR3 (N1856, N1855, N1088, N1217);
nor NOR2 (N1857, N1856, N569);
xor XOR2 (N1858, N1841, N45);
or OR4 (N1859, N1857, N1485, N86, N1086);
xor XOR2 (N1860, N1847, N1190);
not NOT1 (N1861, N1851);
and AND2 (N1862, N1861, N1177);
and AND2 (N1863, N1852, N1628);
nor NOR2 (N1864, N1858, N739);
xor XOR2 (N1865, N1839, N917);
and AND2 (N1866, N1850, N424);
xor XOR2 (N1867, N1854, N132);
not NOT1 (N1868, N1866);
or OR4 (N1869, N1867, N878, N93, N1533);
nor NOR4 (N1870, N1863, N1102, N1810, N1866);
not NOT1 (N1871, N1828);
buf BUF1 (N1872, N1868);
or OR4 (N1873, N1860, N719, N1152, N338);
nand NAND2 (N1874, N1869, N1601);
nor NOR3 (N1875, N1862, N1153, N1833);
nand NAND2 (N1876, N1845, N1514);
buf BUF1 (N1877, N1874);
and AND4 (N1878, N1873, N632, N985, N1493);
xor XOR2 (N1879, N1865, N1222);
nor NOR2 (N1880, N1870, N1582);
xor XOR2 (N1881, N1859, N1754);
xor XOR2 (N1882, N1876, N1554);
buf BUF1 (N1883, N1872);
nor NOR3 (N1884, N1877, N1361, N552);
and AND3 (N1885, N1871, N129, N888);
xor XOR2 (N1886, N1881, N559);
nor NOR3 (N1887, N1875, N1796, N1872);
and AND4 (N1888, N1864, N131, N30, N481);
or OR4 (N1889, N1886, N1819, N1486, N247);
or OR4 (N1890, N1878, N563, N868, N380);
and AND2 (N1891, N1880, N1047);
not NOT1 (N1892, N1888);
xor XOR2 (N1893, N1885, N1257);
xor XOR2 (N1894, N1887, N1577);
xor XOR2 (N1895, N1884, N764);
and AND4 (N1896, N1890, N1118, N595, N779);
and AND4 (N1897, N1893, N527, N430, N1801);
buf BUF1 (N1898, N1879);
nand NAND2 (N1899, N1895, N380);
and AND3 (N1900, N1883, N1491, N53);
nor NOR3 (N1901, N1898, N197, N1471);
not NOT1 (N1902, N1896);
not NOT1 (N1903, N1900);
or OR2 (N1904, N1882, N268);
nand NAND4 (N1905, N1904, N90, N188, N1630);
buf BUF1 (N1906, N1897);
not NOT1 (N1907, N1892);
nand NAND2 (N1908, N1894, N81);
not NOT1 (N1909, N1891);
nand NAND4 (N1910, N1899, N172, N246, N18);
nand NAND3 (N1911, N1909, N584, N1625);
nor NOR4 (N1912, N1902, N1242, N810, N1834);
and AND2 (N1913, N1903, N1343);
xor XOR2 (N1914, N1912, N715);
or OR2 (N1915, N1901, N587);
and AND4 (N1916, N1907, N223, N529, N1617);
not NOT1 (N1917, N1914);
nor NOR2 (N1918, N1905, N1375);
nor NOR4 (N1919, N1906, N744, N867, N1887);
and AND3 (N1920, N1913, N1841, N730);
not NOT1 (N1921, N1917);
and AND4 (N1922, N1918, N1767, N1661, N101);
or OR2 (N1923, N1889, N608);
and AND2 (N1924, N1915, N1233);
and AND4 (N1925, N1908, N224, N1219, N277);
buf BUF1 (N1926, N1919);
nand NAND2 (N1927, N1920, N309);
nand NAND4 (N1928, N1927, N79, N387, N546);
or OR4 (N1929, N1910, N1898, N1518, N1733);
nand NAND3 (N1930, N1921, N132, N464);
buf BUF1 (N1931, N1922);
buf BUF1 (N1932, N1929);
xor XOR2 (N1933, N1911, N548);
xor XOR2 (N1934, N1925, N1872);
nor NOR4 (N1935, N1928, N87, N18, N1384);
and AND2 (N1936, N1931, N923);
nor NOR2 (N1937, N1935, N996);
nor NOR4 (N1938, N1916, N859, N1625, N966);
not NOT1 (N1939, N1924);
not NOT1 (N1940, N1937);
nand NAND3 (N1941, N1938, N712, N723);
nor NOR4 (N1942, N1932, N1114, N1870, N112);
and AND3 (N1943, N1941, N952, N1741);
xor XOR2 (N1944, N1933, N519);
nand NAND4 (N1945, N1942, N737, N434, N1674);
and AND2 (N1946, N1926, N1759);
xor XOR2 (N1947, N1946, N197);
xor XOR2 (N1948, N1943, N153);
buf BUF1 (N1949, N1944);
and AND4 (N1950, N1949, N1886, N1004, N1389);
nor NOR4 (N1951, N1945, N504, N1243, N851);
and AND3 (N1952, N1947, N648, N1337);
or OR4 (N1953, N1951, N1441, N1854, N238);
xor XOR2 (N1954, N1948, N1482);
xor XOR2 (N1955, N1934, N193);
or OR3 (N1956, N1936, N1544, N53);
not NOT1 (N1957, N1955);
nand NAND2 (N1958, N1930, N126);
buf BUF1 (N1959, N1954);
not NOT1 (N1960, N1958);
or OR2 (N1961, N1923, N1773);
and AND3 (N1962, N1960, N1932, N904);
buf BUF1 (N1963, N1956);
xor XOR2 (N1964, N1939, N1320);
not NOT1 (N1965, N1964);
xor XOR2 (N1966, N1953, N1832);
nor NOR2 (N1967, N1961, N892);
buf BUF1 (N1968, N1950);
not NOT1 (N1969, N1957);
and AND2 (N1970, N1969, N1168);
nor NOR2 (N1971, N1965, N234);
nand NAND4 (N1972, N1959, N69, N766, N65);
not NOT1 (N1973, N1968);
and AND4 (N1974, N1973, N197, N1952, N325);
or OR3 (N1975, N455, N264, N721);
xor XOR2 (N1976, N1971, N6);
not NOT1 (N1977, N1967);
xor XOR2 (N1978, N1977, N1820);
or OR4 (N1979, N1963, N1484, N1406, N755);
nand NAND4 (N1980, N1962, N291, N123, N943);
xor XOR2 (N1981, N1978, N1742);
and AND3 (N1982, N1975, N487, N1860);
not NOT1 (N1983, N1940);
not NOT1 (N1984, N1980);
xor XOR2 (N1985, N1979, N349);
not NOT1 (N1986, N1981);
and AND2 (N1987, N1966, N1134);
or OR3 (N1988, N1972, N272, N1488);
not NOT1 (N1989, N1988);
and AND2 (N1990, N1986, N1682);
nand NAND3 (N1991, N1983, N126, N935);
and AND2 (N1992, N1991, N1132);
not NOT1 (N1993, N1990);
and AND2 (N1994, N1974, N1443);
and AND4 (N1995, N1987, N1910, N360, N1216);
nor NOR3 (N1996, N1995, N405, N982);
not NOT1 (N1997, N1989);
and AND4 (N1998, N1997, N928, N1946, N1468);
not NOT1 (N1999, N1982);
xor XOR2 (N2000, N1999, N626);
or OR4 (N2001, N1992, N1887, N1549, N421);
nor NOR4 (N2002, N1994, N1519, N1751, N133);
and AND4 (N2003, N2000, N1561, N1577, N1408);
and AND4 (N2004, N1998, N1152, N833, N1025);
not NOT1 (N2005, N1993);
xor XOR2 (N2006, N2004, N1501);
or OR4 (N2007, N1976, N1734, N1524, N1733);
and AND4 (N2008, N2002, N879, N1423, N1747);
nor NOR2 (N2009, N1996, N200);
buf BUF1 (N2010, N1985);
and AND4 (N2011, N2001, N220, N1514, N1598);
nand NAND3 (N2012, N2010, N1207, N86);
not NOT1 (N2013, N2008);
buf BUF1 (N2014, N2003);
and AND3 (N2015, N2012, N404, N1264);
or OR2 (N2016, N2013, N1085);
not NOT1 (N2017, N2009);
or OR3 (N2018, N2014, N210, N1183);
nor NOR2 (N2019, N2017, N1512);
nor NOR4 (N2020, N2011, N1801, N1789, N82);
and AND2 (N2021, N2007, N737);
and AND2 (N2022, N2021, N535);
nand NAND3 (N2023, N2015, N1299, N546);
nor NOR2 (N2024, N2022, N268);
not NOT1 (N2025, N2018);
xor XOR2 (N2026, N1984, N726);
xor XOR2 (N2027, N2006, N541);
and AND4 (N2028, N2023, N1534, N526, N1363);
or OR3 (N2029, N2025, N800, N707);
not NOT1 (N2030, N2019);
and AND4 (N2031, N2024, N476, N1106, N1858);
or OR4 (N2032, N2027, N209, N949, N1144);
nor NOR2 (N2033, N2032, N1740);
nor NOR4 (N2034, N2020, N1005, N464, N1600);
nor NOR4 (N2035, N2033, N1913, N1315, N976);
buf BUF1 (N2036, N2030);
or OR2 (N2037, N2005, N1707);
not NOT1 (N2038, N2016);
nor NOR2 (N2039, N2038, N566);
not NOT1 (N2040, N2031);
buf BUF1 (N2041, N1970);
buf BUF1 (N2042, N2037);
nand NAND2 (N2043, N2039, N218);
xor XOR2 (N2044, N2036, N775);
nor NOR2 (N2045, N2029, N1842);
xor XOR2 (N2046, N2044, N1521);
and AND3 (N2047, N2034, N609, N103);
nand NAND2 (N2048, N2043, N1689);
xor XOR2 (N2049, N2042, N459);
nand NAND2 (N2050, N2046, N2005);
or OR3 (N2051, N2040, N758, N1763);
and AND4 (N2052, N2051, N1755, N375, N346);
xor XOR2 (N2053, N2041, N1607);
nor NOR2 (N2054, N2050, N508);
nand NAND3 (N2055, N2048, N791, N879);
or OR2 (N2056, N2049, N263);
and AND2 (N2057, N2053, N886);
nand NAND2 (N2058, N2052, N1102);
and AND4 (N2059, N2045, N600, N1848, N1674);
not NOT1 (N2060, N2057);
nor NOR2 (N2061, N2056, N620);
not NOT1 (N2062, N2028);
xor XOR2 (N2063, N2035, N1268);
or OR2 (N2064, N2060, N488);
nand NAND3 (N2065, N2055, N2019, N1346);
or OR4 (N2066, N2065, N682, N1324, N300);
not NOT1 (N2067, N2064);
buf BUF1 (N2068, N2067);
not NOT1 (N2069, N2063);
nand NAND3 (N2070, N2062, N1790, N713);
xor XOR2 (N2071, N2059, N1307);
nand NAND4 (N2072, N2070, N1902, N478, N2039);
xor XOR2 (N2073, N2061, N1925);
buf BUF1 (N2074, N2026);
and AND2 (N2075, N2072, N1072);
not NOT1 (N2076, N2058);
and AND3 (N2077, N2069, N676, N1389);
and AND4 (N2078, N2068, N699, N1233, N40);
not NOT1 (N2079, N2054);
nor NOR4 (N2080, N2077, N540, N1012, N490);
nor NOR3 (N2081, N2080, N176, N495);
not NOT1 (N2082, N2075);
or OR2 (N2083, N2047, N1691);
buf BUF1 (N2084, N2079);
nand NAND2 (N2085, N2081, N208);
nor NOR2 (N2086, N2083, N1812);
nor NOR2 (N2087, N2082, N806);
nor NOR3 (N2088, N2076, N361, N478);
nor NOR2 (N2089, N2066, N39);
nand NAND2 (N2090, N2074, N353);
buf BUF1 (N2091, N2086);
buf BUF1 (N2092, N2090);
nand NAND2 (N2093, N2089, N181);
xor XOR2 (N2094, N2073, N81);
nor NOR3 (N2095, N2093, N1962, N793);
nor NOR4 (N2096, N2088, N544, N2074, N973);
and AND4 (N2097, N2087, N1343, N1668, N872);
not NOT1 (N2098, N2095);
nand NAND3 (N2099, N2097, N1648, N2090);
xor XOR2 (N2100, N2071, N2088);
and AND4 (N2101, N2085, N1826, N1244, N1644);
or OR3 (N2102, N2091, N179, N1604);
not NOT1 (N2103, N2084);
nand NAND4 (N2104, N2100, N725, N276, N1517);
nand NAND2 (N2105, N2096, N1674);
and AND2 (N2106, N2101, N60);
nand NAND2 (N2107, N2105, N98);
nand NAND2 (N2108, N2102, N30);
or OR4 (N2109, N2107, N1927, N132, N1121);
buf BUF1 (N2110, N2106);
nor NOR2 (N2111, N2103, N331);
nor NOR3 (N2112, N2099, N1245, N752);
and AND4 (N2113, N2110, N2014, N295, N421);
not NOT1 (N2114, N2108);
nor NOR4 (N2115, N2104, N584, N1055, N195);
xor XOR2 (N2116, N2094, N225);
or OR2 (N2117, N2115, N1703);
not NOT1 (N2118, N2112);
nor NOR2 (N2119, N2114, N282);
and AND3 (N2120, N2119, N1090, N1383);
not NOT1 (N2121, N2118);
not NOT1 (N2122, N2092);
not NOT1 (N2123, N2111);
nor NOR2 (N2124, N2117, N864);
nand NAND3 (N2125, N2122, N317, N822);
nor NOR3 (N2126, N2098, N1756, N765);
nand NAND3 (N2127, N2116, N973, N768);
buf BUF1 (N2128, N2123);
and AND4 (N2129, N2121, N1911, N958, N311);
and AND2 (N2130, N2109, N414);
not NOT1 (N2131, N2129);
and AND2 (N2132, N2124, N1353);
not NOT1 (N2133, N2126);
nand NAND2 (N2134, N2125, N1108);
not NOT1 (N2135, N2133);
not NOT1 (N2136, N2127);
nor NOR3 (N2137, N2130, N2077, N1385);
and AND3 (N2138, N2132, N855, N1122);
not NOT1 (N2139, N2137);
nand NAND3 (N2140, N2135, N851, N1853);
buf BUF1 (N2141, N2113);
nand NAND4 (N2142, N2078, N1016, N2138, N328);
not NOT1 (N2143, N171);
xor XOR2 (N2144, N2142, N1647);
nand NAND3 (N2145, N2134, N675, N1684);
not NOT1 (N2146, N2139);
nand NAND3 (N2147, N2145, N2103, N57);
buf BUF1 (N2148, N2147);
nor NOR4 (N2149, N2140, N1595, N1643, N934);
nand NAND4 (N2150, N2148, N1229, N411, N513);
nand NAND3 (N2151, N2120, N1288, N1683);
buf BUF1 (N2152, N2151);
nor NOR2 (N2153, N2149, N1075);
buf BUF1 (N2154, N2150);
buf BUF1 (N2155, N2154);
xor XOR2 (N2156, N2131, N1449);
not NOT1 (N2157, N2146);
nand NAND4 (N2158, N2152, N399, N909, N2133);
nand NAND3 (N2159, N2158, N830, N1718);
and AND2 (N2160, N2136, N503);
nand NAND2 (N2161, N2159, N318);
nor NOR3 (N2162, N2161, N899, N195);
or OR4 (N2163, N2162, N2059, N34, N293);
nor NOR3 (N2164, N2128, N449, N275);
and AND4 (N2165, N2143, N2015, N765, N1035);
nor NOR2 (N2166, N2163, N745);
and AND4 (N2167, N2165, N1482, N531, N1063);
nor NOR4 (N2168, N2156, N928, N2035, N1845);
not NOT1 (N2169, N2141);
not NOT1 (N2170, N2160);
and AND2 (N2171, N2144, N444);
xor XOR2 (N2172, N2167, N1886);
not NOT1 (N2173, N2166);
nor NOR4 (N2174, N2170, N739, N44, N1872);
or OR2 (N2175, N2169, N321);
not NOT1 (N2176, N2155);
and AND3 (N2177, N2172, N53, N318);
and AND3 (N2178, N2164, N57, N1755);
or OR2 (N2179, N2153, N2054);
nor NOR4 (N2180, N2174, N992, N709, N1239);
or OR4 (N2181, N2171, N1611, N2049, N1159);
or OR4 (N2182, N2168, N785, N931, N542);
and AND4 (N2183, N2181, N180, N241, N1089);
buf BUF1 (N2184, N2173);
and AND2 (N2185, N2177, N492);
nand NAND4 (N2186, N2184, N1840, N1425, N850);
xor XOR2 (N2187, N2183, N1390);
or OR2 (N2188, N2176, N665);
and AND2 (N2189, N2175, N1884);
buf BUF1 (N2190, N2180);
xor XOR2 (N2191, N2178, N1728);
xor XOR2 (N2192, N2185, N1752);
or OR4 (N2193, N2179, N105, N1443, N1179);
and AND3 (N2194, N2187, N1088, N1662);
buf BUF1 (N2195, N2157);
and AND4 (N2196, N2192, N1824, N881, N837);
xor XOR2 (N2197, N2190, N621);
nand NAND4 (N2198, N2191, N2181, N360, N1431);
not NOT1 (N2199, N2198);
or OR2 (N2200, N2189, N1916);
nor NOR2 (N2201, N2194, N1289);
and AND2 (N2202, N2197, N2129);
nor NOR4 (N2203, N2195, N1483, N1828, N967);
nor NOR3 (N2204, N2200, N1865, N1488);
xor XOR2 (N2205, N2193, N120);
nor NOR3 (N2206, N2196, N260, N432);
or OR3 (N2207, N2182, N1313, N868);
xor XOR2 (N2208, N2186, N45);
buf BUF1 (N2209, N2204);
and AND3 (N2210, N2188, N837, N880);
and AND3 (N2211, N2205, N452, N612);
not NOT1 (N2212, N2203);
nand NAND2 (N2213, N2206, N1360);
or OR4 (N2214, N2201, N43, N394, N749);
or OR4 (N2215, N2208, N1378, N933, N1547);
nand NAND4 (N2216, N2202, N1234, N1886, N513);
or OR3 (N2217, N2211, N1444, N911);
or OR2 (N2218, N2216, N1737);
and AND2 (N2219, N2209, N1632);
xor XOR2 (N2220, N2219, N946);
nor NOR3 (N2221, N2218, N223, N1116);
nand NAND3 (N2222, N2220, N1759, N1903);
nor NOR2 (N2223, N2212, N2125);
and AND4 (N2224, N2223, N1297, N1150, N2109);
not NOT1 (N2225, N2213);
nor NOR4 (N2226, N2215, N1404, N690, N280);
and AND4 (N2227, N2207, N463, N1581, N91);
nor NOR4 (N2228, N2224, N768, N836, N748);
xor XOR2 (N2229, N2222, N386);
xor XOR2 (N2230, N2221, N1854);
and AND3 (N2231, N2229, N2217, N1724);
xor XOR2 (N2232, N1885, N1220);
and AND2 (N2233, N2227, N34);
nand NAND3 (N2234, N2232, N2194, N247);
nor NOR2 (N2235, N2226, N36);
buf BUF1 (N2236, N2234);
not NOT1 (N2237, N2228);
not NOT1 (N2238, N2225);
not NOT1 (N2239, N2235);
nor NOR2 (N2240, N2239, N1508);
nor NOR4 (N2241, N2199, N1370, N609, N1793);
buf BUF1 (N2242, N2214);
and AND2 (N2243, N2237, N1835);
and AND2 (N2244, N2231, N2172);
and AND3 (N2245, N2233, N1736, N2031);
buf BUF1 (N2246, N2244);
nand NAND3 (N2247, N2210, N435, N1394);
buf BUF1 (N2248, N2245);
or OR2 (N2249, N2243, N1805);
or OR4 (N2250, N2230, N62, N372, N2142);
nand NAND3 (N2251, N2247, N777, N1434);
nor NOR3 (N2252, N2242, N1823, N1314);
or OR4 (N2253, N2248, N1484, N252, N408);
nor NOR4 (N2254, N2250, N1812, N1803, N447);
or OR3 (N2255, N2251, N652, N1213);
nor NOR4 (N2256, N2240, N1259, N488, N1664);
nand NAND3 (N2257, N2241, N235, N968);
buf BUF1 (N2258, N2249);
and AND2 (N2259, N2252, N1720);
buf BUF1 (N2260, N2253);
or OR3 (N2261, N2256, N442, N46);
xor XOR2 (N2262, N2259, N1711);
buf BUF1 (N2263, N2257);
or OR4 (N2264, N2254, N1155, N1910, N1738);
buf BUF1 (N2265, N2264);
nand NAND2 (N2266, N2261, N370);
or OR2 (N2267, N2265, N1697);
xor XOR2 (N2268, N2255, N1493);
nand NAND4 (N2269, N2258, N1883, N1348, N1402);
not NOT1 (N2270, N2246);
and AND2 (N2271, N2263, N894);
nor NOR2 (N2272, N2268, N2143);
or OR2 (N2273, N2272, N1574);
nor NOR2 (N2274, N2260, N1998);
not NOT1 (N2275, N2266);
nand NAND4 (N2276, N2274, N301, N234, N2196);
nand NAND3 (N2277, N2270, N1105, N571);
nand NAND3 (N2278, N2269, N1587, N1381);
or OR3 (N2279, N2238, N2041, N1531);
nor NOR2 (N2280, N2273, N184);
nor NOR4 (N2281, N2275, N1608, N757, N1279);
nor NOR2 (N2282, N2236, N353);
buf BUF1 (N2283, N2282);
buf BUF1 (N2284, N2262);
or OR4 (N2285, N2267, N1436, N2284, N2280);
buf BUF1 (N2286, N272);
xor XOR2 (N2287, N1636, N1490);
and AND2 (N2288, N2287, N1408);
xor XOR2 (N2289, N2285, N1871);
buf BUF1 (N2290, N2278);
or OR3 (N2291, N2289, N1943, N2269);
not NOT1 (N2292, N2288);
or OR3 (N2293, N2291, N880, N2076);
nand NAND2 (N2294, N2281, N1201);
xor XOR2 (N2295, N2277, N2202);
not NOT1 (N2296, N2279);
not NOT1 (N2297, N2294);
nor NOR4 (N2298, N2296, N1011, N95, N2146);
and AND2 (N2299, N2297, N625);
nand NAND3 (N2300, N2295, N939, N561);
not NOT1 (N2301, N2271);
xor XOR2 (N2302, N2300, N2053);
or OR2 (N2303, N2286, N2102);
or OR2 (N2304, N2303, N189);
or OR2 (N2305, N2301, N1162);
nand NAND2 (N2306, N2292, N1230);
nand NAND2 (N2307, N2304, N356);
xor XOR2 (N2308, N2307, N1293);
not NOT1 (N2309, N2290);
and AND4 (N2310, N2306, N2138, N1034, N2208);
buf BUF1 (N2311, N2276);
nand NAND4 (N2312, N2305, N1406, N974, N1977);
nor NOR4 (N2313, N2310, N340, N458, N1094);
and AND2 (N2314, N2283, N289);
or OR3 (N2315, N2308, N883, N1176);
nor NOR3 (N2316, N2299, N490, N155);
nor NOR4 (N2317, N2298, N1550, N1595, N2235);
nor NOR3 (N2318, N2311, N902, N1994);
or OR3 (N2319, N2318, N190, N1606);
and AND3 (N2320, N2317, N1685, N2048);
xor XOR2 (N2321, N2319, N97);
and AND4 (N2322, N2302, N360, N989, N1220);
xor XOR2 (N2323, N2322, N1316);
or OR4 (N2324, N2316, N1646, N1421, N1457);
not NOT1 (N2325, N2313);
nor NOR4 (N2326, N2323, N1211, N1521, N1509);
nand NAND3 (N2327, N2312, N357, N2172);
or OR4 (N2328, N2325, N891, N536, N1750);
and AND3 (N2329, N2320, N323, N791);
xor XOR2 (N2330, N2309, N475);
xor XOR2 (N2331, N2321, N1829);
not NOT1 (N2332, N2293);
and AND4 (N2333, N2314, N1306, N382, N1482);
nand NAND3 (N2334, N2331, N1151, N1766);
buf BUF1 (N2335, N2329);
or OR4 (N2336, N2332, N716, N1710, N2234);
xor XOR2 (N2337, N2330, N2011);
buf BUF1 (N2338, N2324);
not NOT1 (N2339, N2333);
buf BUF1 (N2340, N2335);
nor NOR4 (N2341, N2326, N1345, N992, N2046);
or OR2 (N2342, N2337, N767);
nand NAND4 (N2343, N2315, N1114, N538, N1194);
buf BUF1 (N2344, N2328);
not NOT1 (N2345, N2336);
xor XOR2 (N2346, N2343, N788);
nand NAND2 (N2347, N2327, N1644);
nand NAND4 (N2348, N2347, N1965, N878, N1462);
nor NOR3 (N2349, N2340, N94, N2067);
nor NOR4 (N2350, N2348, N1542, N1254, N1665);
or OR4 (N2351, N2341, N2219, N913, N250);
xor XOR2 (N2352, N2351, N710);
not NOT1 (N2353, N2344);
not NOT1 (N2354, N2345);
or OR4 (N2355, N2346, N504, N1444, N1588);
xor XOR2 (N2356, N2353, N897);
or OR4 (N2357, N2354, N2087, N1604, N1394);
nor NOR3 (N2358, N2342, N1460, N604);
xor XOR2 (N2359, N2356, N1209);
nor NOR2 (N2360, N2350, N1626);
buf BUF1 (N2361, N2355);
nand NAND4 (N2362, N2359, N791, N655, N1443);
nor NOR4 (N2363, N2339, N1388, N1419, N1496);
and AND4 (N2364, N2360, N754, N1805, N858);
or OR3 (N2365, N2358, N556, N1172);
nor NOR2 (N2366, N2363, N791);
or OR4 (N2367, N2352, N417, N1204, N349);
nor NOR2 (N2368, N2361, N1725);
nor NOR3 (N2369, N2349, N191, N2285);
buf BUF1 (N2370, N2338);
buf BUF1 (N2371, N2367);
buf BUF1 (N2372, N2368);
buf BUF1 (N2373, N2366);
xor XOR2 (N2374, N2362, N798);
or OR3 (N2375, N2370, N1391, N1370);
nand NAND2 (N2376, N2373, N617);
buf BUF1 (N2377, N2364);
xor XOR2 (N2378, N2374, N2258);
or OR2 (N2379, N2378, N2147);
not NOT1 (N2380, N2371);
nor NOR3 (N2381, N2357, N1992, N1979);
nor NOR4 (N2382, N2380, N2063, N572, N263);
nor NOR4 (N2383, N2334, N218, N997, N1019);
and AND4 (N2384, N2365, N2079, N695, N48);
buf BUF1 (N2385, N2382);
nand NAND2 (N2386, N2377, N1475);
nor NOR4 (N2387, N2379, N107, N858, N1280);
nor NOR2 (N2388, N2386, N58);
and AND2 (N2389, N2384, N981);
xor XOR2 (N2390, N2388, N274);
or OR4 (N2391, N2381, N508, N2340, N1411);
nand NAND2 (N2392, N2376, N1509);
nor NOR3 (N2393, N2391, N210, N1547);
nand NAND4 (N2394, N2369, N2029, N996, N117);
nand NAND4 (N2395, N2394, N1540, N1952, N942);
buf BUF1 (N2396, N2387);
or OR4 (N2397, N2375, N1380, N1161, N1570);
nand NAND3 (N2398, N2383, N1122, N1499);
nor NOR3 (N2399, N2397, N2204, N648);
and AND2 (N2400, N2389, N2048);
buf BUF1 (N2401, N2385);
nor NOR3 (N2402, N2400, N683, N119);
nor NOR4 (N2403, N2392, N850, N1053, N495);
and AND4 (N2404, N2403, N1399, N2206, N405);
or OR4 (N2405, N2401, N1730, N1140, N687);
nor NOR2 (N2406, N2404, N2056);
or OR3 (N2407, N2405, N2075, N1069);
buf BUF1 (N2408, N2402);
and AND4 (N2409, N2372, N1987, N565, N755);
and AND2 (N2410, N2408, N654);
buf BUF1 (N2411, N2396);
not NOT1 (N2412, N2409);
nor NOR3 (N2413, N2390, N1954, N325);
not NOT1 (N2414, N2407);
nor NOR4 (N2415, N2412, N977, N862, N373);
buf BUF1 (N2416, N2393);
and AND3 (N2417, N2414, N501, N902);
or OR3 (N2418, N2417, N527, N998);
nand NAND2 (N2419, N2395, N1299);
xor XOR2 (N2420, N2410, N962);
nor NOR4 (N2421, N2406, N1868, N593, N1989);
xor XOR2 (N2422, N2416, N374);
buf BUF1 (N2423, N2421);
nor NOR2 (N2424, N2420, N624);
buf BUF1 (N2425, N2399);
nand NAND3 (N2426, N2418, N1846, N716);
or OR3 (N2427, N2415, N689, N291);
buf BUF1 (N2428, N2398);
nand NAND3 (N2429, N2425, N64, N1082);
nand NAND2 (N2430, N2426, N673);
nor NOR2 (N2431, N2427, N1661);
buf BUF1 (N2432, N2422);
not NOT1 (N2433, N2432);
xor XOR2 (N2434, N2428, N1848);
and AND4 (N2435, N2424, N1953, N613, N2104);
xor XOR2 (N2436, N2435, N1884);
not NOT1 (N2437, N2423);
and AND2 (N2438, N2429, N751);
or OR3 (N2439, N2438, N1095, N1075);
not NOT1 (N2440, N2434);
nor NOR3 (N2441, N2440, N47, N2176);
not NOT1 (N2442, N2436);
xor XOR2 (N2443, N2433, N2278);
nand NAND3 (N2444, N2443, N1724, N428);
xor XOR2 (N2445, N2430, N2374);
or OR3 (N2446, N2441, N378, N449);
and AND3 (N2447, N2411, N1141, N566);
and AND3 (N2448, N2419, N2017, N1644);
xor XOR2 (N2449, N2413, N859);
nor NOR2 (N2450, N2437, N1269);
or OR2 (N2451, N2446, N2330);
not NOT1 (N2452, N2431);
xor XOR2 (N2453, N2448, N2112);
not NOT1 (N2454, N2449);
xor XOR2 (N2455, N2444, N446);
not NOT1 (N2456, N2445);
nor NOR2 (N2457, N2450, N748);
nor NOR3 (N2458, N2455, N1318, N1722);
buf BUF1 (N2459, N2454);
xor XOR2 (N2460, N2447, N2050);
nand NAND2 (N2461, N2453, N680);
not NOT1 (N2462, N2452);
not NOT1 (N2463, N2442);
not NOT1 (N2464, N2458);
xor XOR2 (N2465, N2439, N2210);
nor NOR4 (N2466, N2457, N1319, N939, N1611);
nand NAND4 (N2467, N2451, N1060, N728, N1174);
or OR4 (N2468, N2462, N2118, N604, N2395);
nand NAND2 (N2469, N2466, N1727);
or OR2 (N2470, N2465, N1010);
or OR3 (N2471, N2459, N783, N440);
buf BUF1 (N2472, N2456);
not NOT1 (N2473, N2471);
or OR2 (N2474, N2464, N1923);
or OR2 (N2475, N2468, N1005);
nand NAND4 (N2476, N2475, N1865, N2058, N1115);
xor XOR2 (N2477, N2467, N1868);
or OR3 (N2478, N2477, N638, N1416);
xor XOR2 (N2479, N2463, N454);
nor NOR3 (N2480, N2461, N534, N1106);
nand NAND2 (N2481, N2472, N1702);
xor XOR2 (N2482, N2481, N857);
nor NOR3 (N2483, N2473, N219, N1326);
or OR3 (N2484, N2482, N2476, N441);
nor NOR3 (N2485, N1036, N41, N532);
not NOT1 (N2486, N2479);
and AND3 (N2487, N2480, N625, N508);
and AND2 (N2488, N2460, N1408);
buf BUF1 (N2489, N2488);
buf BUF1 (N2490, N2474);
nor NOR4 (N2491, N2484, N1553, N1853, N1821);
xor XOR2 (N2492, N2478, N2344);
or OR4 (N2493, N2485, N1464, N563, N2149);
nor NOR2 (N2494, N2489, N1977);
xor XOR2 (N2495, N2486, N1995);
xor XOR2 (N2496, N2469, N1297);
not NOT1 (N2497, N2487);
xor XOR2 (N2498, N2491, N1960);
buf BUF1 (N2499, N2470);
nand NAND2 (N2500, N2496, N938);
not NOT1 (N2501, N2494);
nor NOR2 (N2502, N2495, N443);
and AND4 (N2503, N2499, N122, N1950, N2351);
nor NOR2 (N2504, N2503, N2085);
and AND2 (N2505, N2493, N1071);
or OR2 (N2506, N2504, N181);
nor NOR4 (N2507, N2500, N2293, N623, N1775);
buf BUF1 (N2508, N2490);
nor NOR2 (N2509, N2497, N1460);
and AND4 (N2510, N2509, N1342, N1677, N1806);
buf BUF1 (N2511, N2507);
nor NOR3 (N2512, N2511, N1800, N2186);
nor NOR3 (N2513, N2483, N207, N1572);
nor NOR2 (N2514, N2501, N1180);
nor NOR3 (N2515, N2506, N400, N814);
and AND3 (N2516, N2505, N2079, N1776);
nand NAND3 (N2517, N2510, N613, N1329);
xor XOR2 (N2518, N2516, N1712);
xor XOR2 (N2519, N2513, N45);
and AND4 (N2520, N2512, N69, N703, N1400);
nand NAND2 (N2521, N2520, N223);
nor NOR2 (N2522, N2519, N2256);
and AND2 (N2523, N2498, N489);
buf BUF1 (N2524, N2508);
nor NOR4 (N2525, N2523, N426, N1741, N2037);
nand NAND3 (N2526, N2502, N1764, N1501);
not NOT1 (N2527, N2518);
nand NAND3 (N2528, N2525, N1149, N669);
not NOT1 (N2529, N2515);
buf BUF1 (N2530, N2529);
xor XOR2 (N2531, N2527, N2458);
or OR2 (N2532, N2522, N105);
xor XOR2 (N2533, N2526, N38);
buf BUF1 (N2534, N2517);
nor NOR2 (N2535, N2531, N619);
or OR4 (N2536, N2530, N133, N838, N2242);
xor XOR2 (N2537, N2534, N2394);
and AND2 (N2538, N2536, N1083);
not NOT1 (N2539, N2492);
buf BUF1 (N2540, N2539);
not NOT1 (N2541, N2521);
buf BUF1 (N2542, N2540);
or OR2 (N2543, N2535, N1437);
buf BUF1 (N2544, N2514);
nand NAND3 (N2545, N2538, N1935, N723);
xor XOR2 (N2546, N2542, N1469);
not NOT1 (N2547, N2543);
xor XOR2 (N2548, N2544, N1488);
and AND4 (N2549, N2528, N1142, N1164, N2326);
nand NAND2 (N2550, N2533, N663);
buf BUF1 (N2551, N2549);
or OR4 (N2552, N2546, N1662, N992, N837);
xor XOR2 (N2553, N2551, N2122);
or OR2 (N2554, N2547, N1087);
and AND4 (N2555, N2554, N1072, N599, N436);
or OR2 (N2556, N2555, N743);
and AND2 (N2557, N2532, N1849);
or OR4 (N2558, N2541, N1101, N452, N2390);
buf BUF1 (N2559, N2556);
xor XOR2 (N2560, N2545, N851);
nor NOR3 (N2561, N2550, N1796, N1223);
or OR4 (N2562, N2558, N2362, N1211, N594);
not NOT1 (N2563, N2562);
buf BUF1 (N2564, N2553);
and AND4 (N2565, N2524, N1116, N1146, N2053);
nand NAND3 (N2566, N2537, N1054, N2489);
nor NOR2 (N2567, N2560, N1928);
and AND2 (N2568, N2563, N1532);
or OR4 (N2569, N2561, N1567, N2438, N528);
or OR3 (N2570, N2567, N471, N2558);
not NOT1 (N2571, N2570);
xor XOR2 (N2572, N2566, N1452);
xor XOR2 (N2573, N2565, N2037);
or OR2 (N2574, N2559, N1615);
or OR4 (N2575, N2574, N2160, N1742, N452);
and AND3 (N2576, N2557, N2500, N727);
xor XOR2 (N2577, N2575, N518);
and AND4 (N2578, N2571, N1639, N2572, N13);
nor NOR4 (N2579, N716, N150, N2251, N2125);
nand NAND4 (N2580, N2577, N1654, N419, N592);
nor NOR4 (N2581, N2552, N876, N1138, N114);
buf BUF1 (N2582, N2564);
not NOT1 (N2583, N2568);
buf BUF1 (N2584, N2580);
nand NAND3 (N2585, N2581, N866, N2195);
buf BUF1 (N2586, N2579);
xor XOR2 (N2587, N2578, N1527);
and AND4 (N2588, N2582, N355, N1934, N1846);
nor NOR2 (N2589, N2583, N2583);
xor XOR2 (N2590, N2584, N525);
nand NAND3 (N2591, N2585, N35, N1602);
buf BUF1 (N2592, N2590);
xor XOR2 (N2593, N2576, N791);
or OR3 (N2594, N2593, N1796, N757);
nor NOR3 (N2595, N2548, N1265, N1332);
and AND4 (N2596, N2592, N2045, N1199, N2437);
and AND3 (N2597, N2569, N1153, N1669);
not NOT1 (N2598, N2591);
not NOT1 (N2599, N2589);
buf BUF1 (N2600, N2573);
nor NOR2 (N2601, N2594, N1821);
or OR2 (N2602, N2588, N1505);
xor XOR2 (N2603, N2598, N806);
and AND3 (N2604, N2586, N287, N1106);
or OR3 (N2605, N2587, N2239, N2390);
nand NAND2 (N2606, N2600, N1483);
or OR2 (N2607, N2606, N2329);
or OR2 (N2608, N2599, N1558);
and AND2 (N2609, N2595, N1514);
or OR3 (N2610, N2607, N9, N1192);
buf BUF1 (N2611, N2609);
nand NAND3 (N2612, N2604, N1541, N2447);
or OR4 (N2613, N2597, N2199, N1767, N1853);
nand NAND2 (N2614, N2601, N2405);
not NOT1 (N2615, N2608);
buf BUF1 (N2616, N2603);
not NOT1 (N2617, N2602);
buf BUF1 (N2618, N2610);
nor NOR3 (N2619, N2617, N1421, N1837);
xor XOR2 (N2620, N2618, N597);
nand NAND2 (N2621, N2596, N29);
or OR4 (N2622, N2621, N1518, N2232, N104);
nand NAND4 (N2623, N2614, N1867, N1756, N1226);
or OR4 (N2624, N2612, N301, N922, N1483);
and AND4 (N2625, N2611, N1623, N1406, N1051);
nor NOR4 (N2626, N2613, N816, N244, N1443);
buf BUF1 (N2627, N2616);
nor NOR4 (N2628, N2624, N1642, N267, N1609);
nor NOR2 (N2629, N2623, N517);
not NOT1 (N2630, N2620);
nor NOR4 (N2631, N2619, N1257, N882, N1585);
buf BUF1 (N2632, N2629);
xor XOR2 (N2633, N2625, N289);
buf BUF1 (N2634, N2633);
xor XOR2 (N2635, N2628, N2260);
nor NOR4 (N2636, N2631, N1047, N2631, N683);
xor XOR2 (N2637, N2632, N495);
buf BUF1 (N2638, N2627);
nor NOR2 (N2639, N2635, N1699);
nor NOR4 (N2640, N2626, N2204, N399, N1940);
buf BUF1 (N2641, N2634);
buf BUF1 (N2642, N2640);
not NOT1 (N2643, N2639);
or OR3 (N2644, N2642, N1484, N490);
buf BUF1 (N2645, N2637);
buf BUF1 (N2646, N2622);
nor NOR3 (N2647, N2645, N2435, N1922);
and AND2 (N2648, N2641, N2145);
buf BUF1 (N2649, N2636);
nand NAND2 (N2650, N2643, N464);
buf BUF1 (N2651, N2648);
nand NAND2 (N2652, N2647, N1444);
and AND4 (N2653, N2638, N189, N149, N2168);
nand NAND4 (N2654, N2650, N1927, N1087, N1548);
and AND4 (N2655, N2644, N1936, N1789, N992);
not NOT1 (N2656, N2651);
not NOT1 (N2657, N2615);
and AND3 (N2658, N2652, N2194, N2238);
buf BUF1 (N2659, N2653);
not NOT1 (N2660, N2658);
or OR4 (N2661, N2646, N2125, N1877, N1917);
or OR3 (N2662, N2660, N2383, N81);
and AND3 (N2663, N2661, N844, N348);
nand NAND4 (N2664, N2657, N580, N958, N873);
buf BUF1 (N2665, N2649);
and AND4 (N2666, N2665, N709, N1057, N543);
nor NOR3 (N2667, N2630, N334, N938);
nor NOR2 (N2668, N2662, N784);
or OR4 (N2669, N2659, N262, N2427, N221);
not NOT1 (N2670, N2668);
and AND3 (N2671, N2666, N885, N1189);
nor NOR2 (N2672, N2605, N1340);
xor XOR2 (N2673, N2672, N227);
or OR4 (N2674, N2663, N2572, N2161, N1973);
xor XOR2 (N2675, N2667, N1837);
buf BUF1 (N2676, N2671);
buf BUF1 (N2677, N2670);
buf BUF1 (N2678, N2664);
and AND4 (N2679, N2677, N1729, N2672, N337);
and AND3 (N2680, N2656, N1936, N1566);
and AND2 (N2681, N2679, N93);
buf BUF1 (N2682, N2674);
nor NOR2 (N2683, N2673, N1775);
xor XOR2 (N2684, N2654, N1101);
nand NAND2 (N2685, N2675, N724);
or OR4 (N2686, N2682, N1637, N1911, N1706);
or OR3 (N2687, N2678, N2611, N573);
nor NOR4 (N2688, N2685, N1166, N958, N1682);
not NOT1 (N2689, N2683);
nand NAND2 (N2690, N2689, N782);
or OR4 (N2691, N2686, N618, N1429, N242);
nor NOR4 (N2692, N2691, N515, N2619, N429);
not NOT1 (N2693, N2688);
not NOT1 (N2694, N2693);
nand NAND2 (N2695, N2690, N809);
not NOT1 (N2696, N2692);
buf BUF1 (N2697, N2695);
nand NAND4 (N2698, N2655, N2039, N790, N836);
nor NOR2 (N2699, N2676, N329);
buf BUF1 (N2700, N2698);
or OR2 (N2701, N2697, N478);
not NOT1 (N2702, N2694);
and AND3 (N2703, N2702, N2406, N1563);
and AND3 (N2704, N2701, N2652, N1815);
or OR3 (N2705, N2696, N789, N561);
nor NOR2 (N2706, N2700, N696);
not NOT1 (N2707, N2703);
nand NAND4 (N2708, N2684, N1532, N1938, N923);
and AND3 (N2709, N2687, N138, N817);
xor XOR2 (N2710, N2709, N2083);
not NOT1 (N2711, N2707);
xor XOR2 (N2712, N2708, N1520);
or OR2 (N2713, N2681, N2375);
not NOT1 (N2714, N2712);
nor NOR4 (N2715, N2669, N2620, N471, N1820);
or OR3 (N2716, N2706, N92, N1725);
nand NAND3 (N2717, N2699, N2375, N1790);
nand NAND3 (N2718, N2710, N1539, N1405);
or OR3 (N2719, N2716, N1981, N2052);
not NOT1 (N2720, N2711);
not NOT1 (N2721, N2717);
and AND4 (N2722, N2705, N1609, N824, N1773);
buf BUF1 (N2723, N2722);
not NOT1 (N2724, N2714);
not NOT1 (N2725, N2680);
nor NOR2 (N2726, N2718, N694);
and AND2 (N2727, N2720, N1383);
nor NOR2 (N2728, N2724, N745);
nand NAND2 (N2729, N2727, N2682);
buf BUF1 (N2730, N2728);
and AND2 (N2731, N2715, N1486);
xor XOR2 (N2732, N2726, N1174);
nor NOR4 (N2733, N2732, N638, N2374, N1863);
or OR4 (N2734, N2731, N1060, N2432, N1195);
or OR3 (N2735, N2729, N322, N1631);
and AND4 (N2736, N2719, N815, N1870, N2567);
buf BUF1 (N2737, N2735);
buf BUF1 (N2738, N2733);
nand NAND2 (N2739, N2736, N2327);
buf BUF1 (N2740, N2721);
not NOT1 (N2741, N2739);
or OR2 (N2742, N2737, N1928);
and AND4 (N2743, N2738, N279, N2025, N1266);
and AND4 (N2744, N2730, N612, N975, N2227);
nand NAND2 (N2745, N2734, N372);
xor XOR2 (N2746, N2704, N1255);
xor XOR2 (N2747, N2744, N2204);
not NOT1 (N2748, N2742);
nor NOR3 (N2749, N2748, N2400, N655);
nand NAND4 (N2750, N2749, N1120, N2298, N1261);
not NOT1 (N2751, N2725);
and AND4 (N2752, N2741, N1772, N1826, N2148);
buf BUF1 (N2753, N2750);
not NOT1 (N2754, N2747);
nor NOR3 (N2755, N2743, N68, N1811);
buf BUF1 (N2756, N2745);
not NOT1 (N2757, N2752);
xor XOR2 (N2758, N2755, N2305);
and AND4 (N2759, N2746, N85, N199, N1541);
buf BUF1 (N2760, N2758);
buf BUF1 (N2761, N2754);
xor XOR2 (N2762, N2753, N2498);
buf BUF1 (N2763, N2757);
and AND2 (N2764, N2762, N213);
nand NAND2 (N2765, N2759, N474);
buf BUF1 (N2766, N2765);
and AND2 (N2767, N2713, N1782);
nand NAND4 (N2768, N2766, N1173, N1065, N1914);
buf BUF1 (N2769, N2740);
xor XOR2 (N2770, N2723, N1965);
xor XOR2 (N2771, N2769, N2250);
nor NOR4 (N2772, N2756, N68, N2617, N490);
nor NOR3 (N2773, N2751, N426, N2585);
or OR2 (N2774, N2763, N536);
buf BUF1 (N2775, N2771);
or OR3 (N2776, N2761, N193, N1875);
not NOT1 (N2777, N2764);
xor XOR2 (N2778, N2772, N2277);
or OR4 (N2779, N2760, N1392, N1131, N871);
and AND2 (N2780, N2777, N2689);
not NOT1 (N2781, N2774);
nor NOR3 (N2782, N2776, N577, N1057);
buf BUF1 (N2783, N2781);
xor XOR2 (N2784, N2768, N1862);
nand NAND4 (N2785, N2784, N2420, N2446, N21);
or OR4 (N2786, N2785, N1347, N871, N1813);
buf BUF1 (N2787, N2775);
buf BUF1 (N2788, N2773);
nor NOR2 (N2789, N2783, N1500);
or OR3 (N2790, N2786, N1604, N2480);
buf BUF1 (N2791, N2780);
nor NOR2 (N2792, N2782, N753);
xor XOR2 (N2793, N2787, N961);
not NOT1 (N2794, N2770);
or OR3 (N2795, N2793, N2033, N1202);
not NOT1 (N2796, N2778);
or OR2 (N2797, N2790, N1430);
nor NOR2 (N2798, N2797, N2024);
buf BUF1 (N2799, N2789);
or OR3 (N2800, N2792, N1035, N277);
and AND2 (N2801, N2795, N2463);
and AND4 (N2802, N2767, N2398, N1940, N1172);
or OR4 (N2803, N2779, N1260, N83, N2156);
and AND4 (N2804, N2800, N2704, N784, N2082);
and AND3 (N2805, N2798, N1723, N574);
xor XOR2 (N2806, N2803, N2736);
buf BUF1 (N2807, N2794);
buf BUF1 (N2808, N2788);
xor XOR2 (N2809, N2805, N449);
not NOT1 (N2810, N2804);
or OR3 (N2811, N2796, N2448, N2166);
buf BUF1 (N2812, N2811);
xor XOR2 (N2813, N2812, N1499);
nand NAND3 (N2814, N2806, N1133, N492);
nand NAND2 (N2815, N2801, N414);
buf BUF1 (N2816, N2815);
nand NAND3 (N2817, N2808, N289, N895);
buf BUF1 (N2818, N2817);
and AND2 (N2819, N2802, N918);
and AND2 (N2820, N2816, N1913);
not NOT1 (N2821, N2813);
not NOT1 (N2822, N2820);
and AND4 (N2823, N2822, N1352, N2815, N1184);
not NOT1 (N2824, N2814);
and AND3 (N2825, N2809, N1277, N2335);
nand NAND3 (N2826, N2818, N285, N1124);
buf BUF1 (N2827, N2799);
or OR2 (N2828, N2827, N2492);
xor XOR2 (N2829, N2791, N50);
or OR2 (N2830, N2826, N2541);
buf BUF1 (N2831, N2825);
and AND2 (N2832, N2821, N1273);
or OR3 (N2833, N2823, N2783, N2666);
nor NOR2 (N2834, N2810, N392);
not NOT1 (N2835, N2831);
not NOT1 (N2836, N2807);
buf BUF1 (N2837, N2830);
not NOT1 (N2838, N2834);
buf BUF1 (N2839, N2836);
xor XOR2 (N2840, N2829, N1542);
and AND4 (N2841, N2828, N881, N2620, N1993);
and AND2 (N2842, N2837, N575);
or OR3 (N2843, N2835, N639, N763);
buf BUF1 (N2844, N2838);
buf BUF1 (N2845, N2840);
xor XOR2 (N2846, N2844, N2677);
nor NOR4 (N2847, N2846, N704, N2452, N2729);
nand NAND3 (N2848, N2839, N2475, N1927);
and AND4 (N2849, N2848, N2601, N1614, N2003);
and AND2 (N2850, N2833, N956);
xor XOR2 (N2851, N2850, N1570);
and AND2 (N2852, N2841, N868);
nor NOR3 (N2853, N2851, N149, N918);
buf BUF1 (N2854, N2832);
xor XOR2 (N2855, N2819, N2505);
buf BUF1 (N2856, N2824);
xor XOR2 (N2857, N2855, N1346);
not NOT1 (N2858, N2856);
not NOT1 (N2859, N2845);
or OR3 (N2860, N2859, N1543, N541);
and AND2 (N2861, N2853, N276);
nand NAND4 (N2862, N2847, N1447, N164, N1647);
nand NAND4 (N2863, N2862, N1559, N2528, N2441);
not NOT1 (N2864, N2860);
xor XOR2 (N2865, N2843, N754);
xor XOR2 (N2866, N2861, N2529);
buf BUF1 (N2867, N2854);
buf BUF1 (N2868, N2842);
buf BUF1 (N2869, N2865);
nand NAND2 (N2870, N2867, N1925);
buf BUF1 (N2871, N2849);
nor NOR3 (N2872, N2863, N2089, N21);
nand NAND3 (N2873, N2858, N638, N2754);
not NOT1 (N2874, N2864);
buf BUF1 (N2875, N2873);
xor XOR2 (N2876, N2868, N117);
and AND2 (N2877, N2866, N980);
or OR4 (N2878, N2874, N1510, N1930, N2723);
buf BUF1 (N2879, N2871);
not NOT1 (N2880, N2878);
nor NOR4 (N2881, N2879, N828, N2043, N150);
and AND4 (N2882, N2881, N2421, N777, N934);
nand NAND2 (N2883, N2877, N2255);
or OR3 (N2884, N2870, N510, N2303);
not NOT1 (N2885, N2872);
xor XOR2 (N2886, N2852, N1782);
xor XOR2 (N2887, N2857, N757);
buf BUF1 (N2888, N2886);
nand NAND4 (N2889, N2869, N545, N1129, N2533);
nand NAND4 (N2890, N2885, N226, N1637, N2666);
xor XOR2 (N2891, N2884, N2759);
xor XOR2 (N2892, N2890, N2104);
or OR2 (N2893, N2880, N1134);
and AND2 (N2894, N2891, N1584);
or OR3 (N2895, N2894, N2076, N673);
nand NAND2 (N2896, N2887, N2331);
xor XOR2 (N2897, N2876, N803);
buf BUF1 (N2898, N2883);
or OR3 (N2899, N2895, N2795, N594);
nor NOR2 (N2900, N2899, N1210);
and AND2 (N2901, N2900, N536);
nand NAND3 (N2902, N2892, N1454, N2468);
and AND3 (N2903, N2897, N729, N2166);
and AND4 (N2904, N2902, N970, N1026, N1535);
buf BUF1 (N2905, N2901);
buf BUF1 (N2906, N2875);
or OR4 (N2907, N2896, N82, N581, N689);
nor NOR4 (N2908, N2907, N1585, N741, N1713);
not NOT1 (N2909, N2893);
buf BUF1 (N2910, N2908);
and AND4 (N2911, N2888, N967, N1871, N1213);
nor NOR3 (N2912, N2906, N1414, N176);
nand NAND2 (N2913, N2904, N2292);
or OR4 (N2914, N2898, N243, N1592, N2563);
nand NAND3 (N2915, N2889, N1244, N594);
nand NAND2 (N2916, N2910, N1098);
nor NOR2 (N2917, N2912, N354);
and AND2 (N2918, N2913, N2664);
and AND3 (N2919, N2909, N1010, N1532);
or OR4 (N2920, N2882, N1183, N2674, N2291);
xor XOR2 (N2921, N2917, N1770);
nor NOR4 (N2922, N2919, N480, N794, N79);
and AND3 (N2923, N2921, N2316, N579);
or OR2 (N2924, N2915, N2243);
and AND3 (N2925, N2905, N286, N1080);
xor XOR2 (N2926, N2924, N681);
not NOT1 (N2927, N2918);
buf BUF1 (N2928, N2911);
not NOT1 (N2929, N2922);
not NOT1 (N2930, N2903);
nand NAND2 (N2931, N2930, N2115);
not NOT1 (N2932, N2914);
or OR3 (N2933, N2931, N2519, N1326);
nand NAND4 (N2934, N2920, N1327, N1143, N1068);
nand NAND2 (N2935, N2925, N1413);
xor XOR2 (N2936, N2928, N214);
nand NAND4 (N2937, N2929, N594, N1810, N2163);
buf BUF1 (N2938, N2927);
buf BUF1 (N2939, N2933);
xor XOR2 (N2940, N2926, N1375);
xor XOR2 (N2941, N2934, N864);
xor XOR2 (N2942, N2938, N1728);
buf BUF1 (N2943, N2939);
nand NAND3 (N2944, N2916, N1539, N2899);
nand NAND4 (N2945, N2937, N1500, N2699, N2941);
not NOT1 (N2946, N1141);
and AND3 (N2947, N2935, N1640, N2788);
nand NAND3 (N2948, N2945, N2824, N2405);
nand NAND3 (N2949, N2932, N2771, N1884);
not NOT1 (N2950, N2936);
and AND2 (N2951, N2940, N490);
not NOT1 (N2952, N2947);
xor XOR2 (N2953, N2942, N738);
or OR2 (N2954, N2923, N2676);
nor NOR4 (N2955, N2952, N1299, N1268, N1272);
not NOT1 (N2956, N2949);
nor NOR4 (N2957, N2944, N1931, N310, N2391);
buf BUF1 (N2958, N2955);
nor NOR4 (N2959, N2953, N573, N836, N1101);
xor XOR2 (N2960, N2948, N1299);
xor XOR2 (N2961, N2957, N438);
nor NOR3 (N2962, N2951, N499, N1222);
buf BUF1 (N2963, N2962);
nor NOR4 (N2964, N2946, N2379, N1261, N2460);
buf BUF1 (N2965, N2954);
and AND3 (N2966, N2943, N2831, N594);
and AND3 (N2967, N2961, N878, N265);
not NOT1 (N2968, N2959);
and AND3 (N2969, N2950, N1363, N2548);
not NOT1 (N2970, N2963);
xor XOR2 (N2971, N2965, N125);
not NOT1 (N2972, N2956);
nand NAND2 (N2973, N2958, N1461);
nand NAND3 (N2974, N2960, N2878, N830);
xor XOR2 (N2975, N2967, N2686);
buf BUF1 (N2976, N2968);
nor NOR2 (N2977, N2970, N751);
nand NAND2 (N2978, N2973, N2200);
xor XOR2 (N2979, N2976, N1403);
xor XOR2 (N2980, N2975, N247);
or OR3 (N2981, N2974, N2225, N103);
nand NAND2 (N2982, N2979, N890);
xor XOR2 (N2983, N2972, N2622);
not NOT1 (N2984, N2980);
nor NOR4 (N2985, N2983, N1309, N2243, N2774);
buf BUF1 (N2986, N2985);
xor XOR2 (N2987, N2977, N695);
nand NAND2 (N2988, N2987, N577);
or OR4 (N2989, N2984, N820, N594, N1712);
not NOT1 (N2990, N2966);
nor NOR4 (N2991, N2988, N1946, N969, N2463);
buf BUF1 (N2992, N2978);
not NOT1 (N2993, N2971);
nor NOR2 (N2994, N2982, N744);
xor XOR2 (N2995, N2969, N2619);
nand NAND4 (N2996, N2989, N2501, N208, N2450);
not NOT1 (N2997, N2996);
xor XOR2 (N2998, N2992, N958);
xor XOR2 (N2999, N2994, N1702);
and AND4 (N3000, N2986, N1996, N500, N1613);
and AND3 (N3001, N2993, N1099, N1513);
nand NAND2 (N3002, N2995, N1535);
nor NOR4 (N3003, N2964, N776, N2076, N2295);
or OR4 (N3004, N3001, N1679, N2641, N493);
buf BUF1 (N3005, N2981);
and AND2 (N3006, N2997, N538);
buf BUF1 (N3007, N3004);
or OR4 (N3008, N2990, N204, N1660, N2274);
buf BUF1 (N3009, N3007);
and AND2 (N3010, N3006, N1838);
nor NOR2 (N3011, N2999, N46);
and AND3 (N3012, N3010, N2069, N2499);
buf BUF1 (N3013, N3008);
buf BUF1 (N3014, N3012);
buf BUF1 (N3015, N2991);
nand NAND3 (N3016, N3011, N1961, N358);
nand NAND4 (N3017, N3009, N168, N1659, N1862);
xor XOR2 (N3018, N3000, N2327);
xor XOR2 (N3019, N3018, N2840);
and AND3 (N3020, N3002, N2716, N1214);
buf BUF1 (N3021, N3003);
nand NAND3 (N3022, N3005, N1371, N646);
and AND4 (N3023, N3017, N969, N1370, N483);
xor XOR2 (N3024, N3022, N2280);
not NOT1 (N3025, N3021);
or OR2 (N3026, N3014, N776);
nor NOR3 (N3027, N3013, N2637, N832);
not NOT1 (N3028, N3023);
buf BUF1 (N3029, N3020);
nand NAND3 (N3030, N3025, N437, N152);
xor XOR2 (N3031, N3026, N2771);
nand NAND4 (N3032, N3028, N1811, N1827, N395);
xor XOR2 (N3033, N3019, N1913);
buf BUF1 (N3034, N3033);
and AND3 (N3035, N3015, N2500, N1688);
or OR3 (N3036, N3030, N1285, N1785);
nand NAND3 (N3037, N3029, N1615, N1170);
or OR3 (N3038, N3034, N2180, N413);
and AND4 (N3039, N3035, N2090, N792, N634);
nand NAND3 (N3040, N3038, N750, N2401);
and AND2 (N3041, N3016, N871);
buf BUF1 (N3042, N3036);
nand NAND2 (N3043, N3027, N2125);
xor XOR2 (N3044, N3040, N1038);
nor NOR2 (N3045, N2998, N2685);
xor XOR2 (N3046, N3037, N389);
xor XOR2 (N3047, N3045, N1518);
and AND4 (N3048, N3031, N2409, N303, N1687);
xor XOR2 (N3049, N3042, N1207);
buf BUF1 (N3050, N3048);
not NOT1 (N3051, N3047);
or OR2 (N3052, N3032, N2840);
xor XOR2 (N3053, N3043, N1762);
nor NOR4 (N3054, N3053, N1205, N1510, N2510);
not NOT1 (N3055, N3054);
nor NOR3 (N3056, N3050, N1291, N1348);
or OR2 (N3057, N3039, N1288);
xor XOR2 (N3058, N3024, N226);
not NOT1 (N3059, N3058);
or OR2 (N3060, N3046, N1897);
buf BUF1 (N3061, N3055);
and AND2 (N3062, N3057, N2974);
not NOT1 (N3063, N3056);
nor NOR3 (N3064, N3059, N1766, N619);
not NOT1 (N3065, N3049);
xor XOR2 (N3066, N3065, N1079);
buf BUF1 (N3067, N3061);
and AND3 (N3068, N3064, N170, N1641);
and AND3 (N3069, N3060, N1203, N1673);
nand NAND2 (N3070, N3066, N1881);
buf BUF1 (N3071, N3068);
not NOT1 (N3072, N3071);
nand NAND2 (N3073, N3052, N1645);
nand NAND4 (N3074, N3073, N1077, N2741, N2021);
nor NOR3 (N3075, N3067, N2474, N2881);
nor NOR4 (N3076, N3074, N977, N1364, N224);
and AND3 (N3077, N3069, N2749, N155);
buf BUF1 (N3078, N3070);
not NOT1 (N3079, N3075);
nor NOR3 (N3080, N3077, N2121, N595);
and AND4 (N3081, N3041, N2452, N3020, N1576);
nor NOR3 (N3082, N3051, N1834, N2568);
nor NOR2 (N3083, N3079, N232);
not NOT1 (N3084, N3078);
and AND3 (N3085, N3082, N563, N1463);
nand NAND2 (N3086, N3062, N957);
buf BUF1 (N3087, N3072);
nor NOR2 (N3088, N3085, N2470);
nor NOR4 (N3089, N3076, N2798, N851, N2999);
nand NAND3 (N3090, N3088, N1157, N2465);
or OR2 (N3091, N3090, N2117);
not NOT1 (N3092, N3084);
and AND3 (N3093, N3091, N1535, N989);
xor XOR2 (N3094, N3086, N2126);
buf BUF1 (N3095, N3093);
xor XOR2 (N3096, N3080, N1398);
nand NAND4 (N3097, N3096, N2184, N1959, N369);
nor NOR4 (N3098, N3097, N113, N2740, N1884);
not NOT1 (N3099, N3092);
xor XOR2 (N3100, N3089, N230);
xor XOR2 (N3101, N3099, N1553);
or OR4 (N3102, N3101, N979, N1431, N193);
nor NOR2 (N3103, N3102, N2089);
or OR3 (N3104, N3098, N1211, N47);
buf BUF1 (N3105, N3087);
xor XOR2 (N3106, N3083, N2418);
xor XOR2 (N3107, N3095, N2880);
nand NAND2 (N3108, N3104, N1981);
or OR2 (N3109, N3044, N602);
nand NAND4 (N3110, N3107, N1098, N157, N1512);
buf BUF1 (N3111, N3103);
not NOT1 (N3112, N3109);
and AND2 (N3113, N3081, N2398);
buf BUF1 (N3114, N3100);
xor XOR2 (N3115, N3106, N341);
buf BUF1 (N3116, N3094);
or OR2 (N3117, N3110, N2859);
nor NOR2 (N3118, N3116, N2620);
nand NAND4 (N3119, N3117, N1116, N1441, N243);
nand NAND2 (N3120, N3111, N2911);
and AND2 (N3121, N3113, N520);
xor XOR2 (N3122, N3114, N2666);
nor NOR3 (N3123, N3122, N2560, N1194);
buf BUF1 (N3124, N3123);
nor NOR2 (N3125, N3108, N464);
not NOT1 (N3126, N3063);
xor XOR2 (N3127, N3125, N1475);
nor NOR4 (N3128, N3127, N2018, N1314, N593);
and AND2 (N3129, N3124, N183);
nor NOR4 (N3130, N3119, N798, N1438, N1767);
buf BUF1 (N3131, N3130);
and AND3 (N3132, N3128, N1221, N3105);
nand NAND2 (N3133, N769, N912);
xor XOR2 (N3134, N3121, N1250);
buf BUF1 (N3135, N3120);
nand NAND3 (N3136, N3133, N1545, N607);
buf BUF1 (N3137, N3136);
nor NOR4 (N3138, N3126, N61, N2563, N4);
buf BUF1 (N3139, N3137);
nor NOR2 (N3140, N3135, N1447);
nand NAND3 (N3141, N3139, N2719, N2401);
and AND3 (N3142, N3138, N680, N2461);
xor XOR2 (N3143, N3129, N3104);
buf BUF1 (N3144, N3141);
nor NOR3 (N3145, N3118, N2774, N175);
nand NAND3 (N3146, N3115, N2760, N2626);
nand NAND2 (N3147, N3144, N1833);
buf BUF1 (N3148, N3143);
buf BUF1 (N3149, N3142);
and AND2 (N3150, N3132, N1785);
buf BUF1 (N3151, N3148);
nor NOR3 (N3152, N3149, N905, N1507);
xor XOR2 (N3153, N3152, N1168);
and AND4 (N3154, N3134, N33, N2813, N2170);
nand NAND2 (N3155, N3150, N1676);
nor NOR3 (N3156, N3145, N2010, N1469);
not NOT1 (N3157, N3154);
or OR2 (N3158, N3155, N617);
not NOT1 (N3159, N3146);
not NOT1 (N3160, N3147);
nor NOR2 (N3161, N3151, N2692);
buf BUF1 (N3162, N3131);
xor XOR2 (N3163, N3112, N308);
xor XOR2 (N3164, N3160, N2827);
not NOT1 (N3165, N3159);
and AND4 (N3166, N3161, N2171, N1523, N2786);
nand NAND3 (N3167, N3166, N187, N2274);
and AND3 (N3168, N3156, N2050, N891);
nor NOR4 (N3169, N3164, N117, N269, N2506);
nand NAND3 (N3170, N3153, N540, N295);
and AND2 (N3171, N3165, N2383);
or OR3 (N3172, N3163, N2583, N391);
or OR4 (N3173, N3167, N976, N2704, N1868);
not NOT1 (N3174, N3171);
xor XOR2 (N3175, N3170, N878);
nand NAND3 (N3176, N3174, N667, N1369);
not NOT1 (N3177, N3172);
nand NAND2 (N3178, N3162, N1339);
nor NOR2 (N3179, N3169, N1411);
not NOT1 (N3180, N3158);
nand NAND3 (N3181, N3157, N2288, N93);
not NOT1 (N3182, N3180);
nor NOR4 (N3183, N3173, N137, N1481, N1274);
nor NOR4 (N3184, N3179, N2615, N545, N1182);
and AND4 (N3185, N3182, N404, N294, N2455);
or OR4 (N3186, N3176, N1379, N2859, N913);
and AND2 (N3187, N3175, N427);
nor NOR2 (N3188, N3187, N2832);
xor XOR2 (N3189, N3183, N1095);
buf BUF1 (N3190, N3186);
or OR4 (N3191, N3177, N2757, N936, N1021);
or OR3 (N3192, N3188, N2217, N586);
xor XOR2 (N3193, N3189, N1986);
nor NOR3 (N3194, N3192, N1722, N2346);
not NOT1 (N3195, N3168);
and AND2 (N3196, N3181, N3083);
or OR3 (N3197, N3195, N419, N2230);
or OR2 (N3198, N3185, N2756);
or OR2 (N3199, N3193, N1761);
not NOT1 (N3200, N3199);
not NOT1 (N3201, N3140);
not NOT1 (N3202, N3190);
not NOT1 (N3203, N3196);
xor XOR2 (N3204, N3184, N2414);
or OR3 (N3205, N3194, N224, N2735);
or OR4 (N3206, N3205, N563, N1099, N742);
not NOT1 (N3207, N3203);
nor NOR2 (N3208, N3178, N1257);
nand NAND3 (N3209, N3202, N1425, N2745);
nand NAND2 (N3210, N3209, N470);
not NOT1 (N3211, N3208);
and AND4 (N3212, N3210, N296, N1385, N1427);
buf BUF1 (N3213, N3212);
not NOT1 (N3214, N3198);
buf BUF1 (N3215, N3214);
or OR4 (N3216, N3215, N3006, N2146, N1388);
or OR4 (N3217, N3216, N3173, N432, N1184);
or OR2 (N3218, N3201, N2525);
or OR2 (N3219, N3218, N2634);
xor XOR2 (N3220, N3213, N2707);
buf BUF1 (N3221, N3191);
buf BUF1 (N3222, N3207);
and AND2 (N3223, N3200, N37);
xor XOR2 (N3224, N3197, N1301);
buf BUF1 (N3225, N3223);
or OR3 (N3226, N3221, N2938, N963);
buf BUF1 (N3227, N3220);
xor XOR2 (N3228, N3206, N1021);
nand NAND2 (N3229, N3219, N3087);
nor NOR3 (N3230, N3217, N3196, N2514);
xor XOR2 (N3231, N3211, N2860);
or OR2 (N3232, N3226, N2370);
xor XOR2 (N3233, N3225, N2131);
xor XOR2 (N3234, N3227, N462);
and AND2 (N3235, N3233, N761);
buf BUF1 (N3236, N3229);
and AND3 (N3237, N3224, N1249, N1723);
or OR3 (N3238, N3232, N1873, N1994);
or OR4 (N3239, N3238, N2648, N2156, N357);
nand NAND3 (N3240, N3204, N1487, N1645);
nor NOR2 (N3241, N3230, N1161);
xor XOR2 (N3242, N3239, N2470);
xor XOR2 (N3243, N3237, N2103);
or OR2 (N3244, N3234, N2450);
buf BUF1 (N3245, N3231);
buf BUF1 (N3246, N3228);
buf BUF1 (N3247, N3236);
and AND4 (N3248, N3247, N502, N3039, N585);
not NOT1 (N3249, N3222);
nand NAND4 (N3250, N3244, N744, N2918, N2973);
xor XOR2 (N3251, N3242, N3227);
buf BUF1 (N3252, N3241);
buf BUF1 (N3253, N3252);
xor XOR2 (N3254, N3248, N417);
nor NOR2 (N3255, N3240, N2070);
and AND3 (N3256, N3245, N9, N2470);
or OR4 (N3257, N3256, N2597, N2418, N1012);
and AND4 (N3258, N3257, N2722, N1184, N1723);
not NOT1 (N3259, N3251);
buf BUF1 (N3260, N3255);
not NOT1 (N3261, N3260);
buf BUF1 (N3262, N3254);
buf BUF1 (N3263, N3235);
xor XOR2 (N3264, N3258, N1507);
nor NOR3 (N3265, N3253, N765, N3197);
not NOT1 (N3266, N3243);
not NOT1 (N3267, N3266);
and AND2 (N3268, N3246, N176);
xor XOR2 (N3269, N3261, N673);
xor XOR2 (N3270, N3269, N1653);
nor NOR4 (N3271, N3268, N1513, N2117, N2503);
nand NAND2 (N3272, N3263, N730);
or OR4 (N3273, N3250, N326, N2949, N1435);
buf BUF1 (N3274, N3249);
xor XOR2 (N3275, N3274, N104);
or OR3 (N3276, N3264, N800, N3274);
nor NOR4 (N3277, N3273, N765, N1552, N2473);
and AND2 (N3278, N3265, N2430);
xor XOR2 (N3279, N3272, N3238);
xor XOR2 (N3280, N3277, N2773);
not NOT1 (N3281, N3267);
not NOT1 (N3282, N3279);
and AND3 (N3283, N3281, N2993, N2259);
or OR4 (N3284, N3271, N1951, N1188, N933);
nor NOR2 (N3285, N3270, N465);
or OR4 (N3286, N3278, N1362, N1783, N3247);
or OR2 (N3287, N3262, N699);
nor NOR4 (N3288, N3275, N1779, N2911, N611);
nor NOR4 (N3289, N3283, N2244, N2956, N157);
or OR4 (N3290, N3282, N2875, N976, N1220);
nand NAND3 (N3291, N3280, N2884, N1385);
xor XOR2 (N3292, N3289, N3211);
not NOT1 (N3293, N3259);
buf BUF1 (N3294, N3285);
nor NOR3 (N3295, N3288, N2387, N1967);
or OR2 (N3296, N3286, N817);
xor XOR2 (N3297, N3292, N1525);
xor XOR2 (N3298, N3293, N2980);
and AND4 (N3299, N3291, N453, N3004, N550);
or OR4 (N3300, N3287, N1599, N942, N2155);
buf BUF1 (N3301, N3299);
nand NAND4 (N3302, N3284, N2756, N472, N2885);
or OR4 (N3303, N3294, N534, N662, N2368);
xor XOR2 (N3304, N3298, N2822);
nor NOR2 (N3305, N3296, N2185);
not NOT1 (N3306, N3295);
xor XOR2 (N3307, N3303, N2671);
or OR3 (N3308, N3297, N210, N1510);
nand NAND3 (N3309, N3300, N3220, N578);
xor XOR2 (N3310, N3301, N67);
xor XOR2 (N3311, N3309, N2690);
nor NOR4 (N3312, N3305, N2889, N2584, N1962);
nand NAND4 (N3313, N3304, N1583, N1846, N438);
xor XOR2 (N3314, N3307, N1498);
buf BUF1 (N3315, N3302);
nand NAND2 (N3316, N3312, N829);
buf BUF1 (N3317, N3313);
buf BUF1 (N3318, N3310);
buf BUF1 (N3319, N3290);
not NOT1 (N3320, N3319);
xor XOR2 (N3321, N3316, N271);
nand NAND3 (N3322, N3321, N496, N1293);
nand NAND2 (N3323, N3317, N3025);
buf BUF1 (N3324, N3322);
xor XOR2 (N3325, N3315, N2692);
xor XOR2 (N3326, N3325, N2962);
xor XOR2 (N3327, N3326, N3112);
buf BUF1 (N3328, N3314);
or OR4 (N3329, N3311, N2064, N733, N984);
not NOT1 (N3330, N3318);
xor XOR2 (N3331, N3327, N2731);
and AND4 (N3332, N3323, N1709, N2125, N2303);
or OR2 (N3333, N3330, N113);
nor NOR3 (N3334, N3328, N2007, N2003);
not NOT1 (N3335, N3276);
not NOT1 (N3336, N3334);
xor XOR2 (N3337, N3308, N2103);
nand NAND2 (N3338, N3320, N825);
and AND3 (N3339, N3332, N108, N2029);
nor NOR4 (N3340, N3331, N477, N235, N2168);
not NOT1 (N3341, N3336);
or OR4 (N3342, N3306, N767, N587, N1188);
xor XOR2 (N3343, N3340, N612);
nor NOR4 (N3344, N3333, N1520, N2005, N1981);
buf BUF1 (N3345, N3343);
buf BUF1 (N3346, N3344);
and AND3 (N3347, N3329, N2416, N2461);
and AND3 (N3348, N3341, N942, N2531);
and AND4 (N3349, N3337, N2915, N2212, N857);
xor XOR2 (N3350, N3342, N2556);
not NOT1 (N3351, N3339);
or OR4 (N3352, N3338, N1674, N3298, N1297);
not NOT1 (N3353, N3347);
xor XOR2 (N3354, N3352, N1410);
xor XOR2 (N3355, N3348, N2086);
nand NAND2 (N3356, N3345, N3125);
xor XOR2 (N3357, N3353, N1623);
xor XOR2 (N3358, N3324, N1275);
buf BUF1 (N3359, N3351);
or OR2 (N3360, N3354, N1172);
and AND4 (N3361, N3356, N368, N3312, N602);
not NOT1 (N3362, N3346);
or OR2 (N3363, N3349, N1307);
nand NAND2 (N3364, N3363, N1472);
not NOT1 (N3365, N3362);
xor XOR2 (N3366, N3357, N1463);
or OR3 (N3367, N3355, N2542, N2464);
xor XOR2 (N3368, N3366, N1359);
nand NAND4 (N3369, N3365, N1771, N4, N1134);
and AND2 (N3370, N3335, N721);
xor XOR2 (N3371, N3361, N1692);
or OR2 (N3372, N3358, N106);
buf BUF1 (N3373, N3350);
nor NOR2 (N3374, N3367, N358);
buf BUF1 (N3375, N3364);
or OR4 (N3376, N3369, N2976, N1416, N2327);
nor NOR3 (N3377, N3368, N1458, N1972);
buf BUF1 (N3378, N3373);
nand NAND3 (N3379, N3371, N2599, N508);
nor NOR3 (N3380, N3377, N2739, N902);
nand NAND3 (N3381, N3378, N2308, N182);
and AND3 (N3382, N3380, N1829, N2028);
and AND3 (N3383, N3381, N1010, N940);
nor NOR3 (N3384, N3360, N2485, N1766);
not NOT1 (N3385, N3376);
not NOT1 (N3386, N3359);
and AND3 (N3387, N3370, N714, N2147);
buf BUF1 (N3388, N3385);
not NOT1 (N3389, N3382);
and AND4 (N3390, N3384, N2063, N768, N2752);
not NOT1 (N3391, N3379);
buf BUF1 (N3392, N3388);
nor NOR3 (N3393, N3389, N314, N3006);
not NOT1 (N3394, N3383);
or OR2 (N3395, N3390, N1004);
or OR3 (N3396, N3387, N967, N2362);
not NOT1 (N3397, N3392);
xor XOR2 (N3398, N3372, N160);
not NOT1 (N3399, N3391);
or OR4 (N3400, N3396, N515, N3066, N2168);
buf BUF1 (N3401, N3374);
and AND4 (N3402, N3386, N1431, N2378, N382);
buf BUF1 (N3403, N3395);
nor NOR2 (N3404, N3402, N2746);
not NOT1 (N3405, N3404);
and AND4 (N3406, N3398, N2724, N1467, N774);
nand NAND4 (N3407, N3405, N3164, N2752, N1896);
nand NAND3 (N3408, N3406, N759, N443);
nor NOR4 (N3409, N3403, N2798, N827, N2185);
xor XOR2 (N3410, N3409, N810);
or OR4 (N3411, N3375, N969, N1265, N1594);
buf BUF1 (N3412, N3410);
not NOT1 (N3413, N3393);
buf BUF1 (N3414, N3408);
xor XOR2 (N3415, N3399, N1003);
nand NAND3 (N3416, N3413, N2281, N412);
and AND3 (N3417, N3412, N1752, N3007);
not NOT1 (N3418, N3417);
buf BUF1 (N3419, N3414);
nand NAND4 (N3420, N3419, N2028, N2380, N495);
nor NOR3 (N3421, N3400, N2560, N3150);
xor XOR2 (N3422, N3415, N689);
and AND2 (N3423, N3401, N1807);
not NOT1 (N3424, N3407);
xor XOR2 (N3425, N3420, N3005);
nand NAND4 (N3426, N3397, N2457, N2500, N1230);
not NOT1 (N3427, N3426);
or OR4 (N3428, N3394, N2384, N2899, N3318);
nand NAND3 (N3429, N3424, N3190, N1052);
or OR3 (N3430, N3421, N742, N1704);
nand NAND2 (N3431, N3422, N2153);
xor XOR2 (N3432, N3423, N106);
or OR3 (N3433, N3411, N3183, N1019);
xor XOR2 (N3434, N3416, N1190);
xor XOR2 (N3435, N3429, N319);
buf BUF1 (N3436, N3428);
or OR3 (N3437, N3431, N3128, N3340);
and AND3 (N3438, N3436, N1671, N1159);
or OR4 (N3439, N3425, N93, N169, N1899);
nor NOR3 (N3440, N3433, N3311, N2840);
nand NAND2 (N3441, N3435, N1393);
nor NOR4 (N3442, N3418, N395, N3156, N3381);
buf BUF1 (N3443, N3441);
not NOT1 (N3444, N3437);
nand NAND2 (N3445, N3430, N178);
xor XOR2 (N3446, N3427, N753);
nand NAND3 (N3447, N3446, N2238, N2206);
or OR4 (N3448, N3434, N1015, N1130, N2548);
nand NAND4 (N3449, N3443, N2207, N1931, N2973);
xor XOR2 (N3450, N3448, N2335);
xor XOR2 (N3451, N3444, N2129);
buf BUF1 (N3452, N3445);
nand NAND4 (N3453, N3452, N3274, N2332, N1573);
nand NAND4 (N3454, N3439, N446, N500, N1688);
buf BUF1 (N3455, N3447);
nand NAND4 (N3456, N3454, N2232, N99, N3238);
buf BUF1 (N3457, N3442);
or OR4 (N3458, N3438, N2907, N2591, N32);
and AND4 (N3459, N3440, N3116, N305, N545);
xor XOR2 (N3460, N3451, N309);
xor XOR2 (N3461, N3432, N433);
xor XOR2 (N3462, N3461, N2048);
not NOT1 (N3463, N3453);
or OR4 (N3464, N3455, N2430, N1462, N926);
nor NOR2 (N3465, N3456, N2239);
and AND3 (N3466, N3460, N102, N2208);
and AND3 (N3467, N3462, N1155, N952);
nor NOR4 (N3468, N3458, N2093, N247, N608);
or OR3 (N3469, N3466, N1948, N3104);
nor NOR3 (N3470, N3465, N2118, N977);
and AND4 (N3471, N3464, N2895, N3237, N662);
buf BUF1 (N3472, N3470);
nand NAND2 (N3473, N3457, N1626);
buf BUF1 (N3474, N3473);
xor XOR2 (N3475, N3472, N2029);
nor NOR2 (N3476, N3475, N1998);
nor NOR3 (N3477, N3468, N2323, N747);
and AND4 (N3478, N3471, N2324, N3382, N2806);
buf BUF1 (N3479, N3459);
not NOT1 (N3480, N3463);
not NOT1 (N3481, N3478);
nor NOR3 (N3482, N3449, N2029, N1009);
not NOT1 (N3483, N3479);
not NOT1 (N3484, N3480);
and AND4 (N3485, N3467, N2163, N2944, N3096);
or OR2 (N3486, N3476, N700);
or OR3 (N3487, N3474, N514, N1478);
buf BUF1 (N3488, N3450);
and AND3 (N3489, N3484, N1283, N1630);
not NOT1 (N3490, N3486);
not NOT1 (N3491, N3481);
xor XOR2 (N3492, N3488, N1726);
buf BUF1 (N3493, N3490);
nor NOR4 (N3494, N3477, N1892, N728, N3430);
not NOT1 (N3495, N3492);
or OR4 (N3496, N3489, N1715, N1810, N2889);
buf BUF1 (N3497, N3495);
not NOT1 (N3498, N3493);
and AND4 (N3499, N3485, N1437, N491, N1420);
or OR2 (N3500, N3469, N2152);
xor XOR2 (N3501, N3496, N2810);
nand NAND2 (N3502, N3482, N1654);
and AND4 (N3503, N3498, N2116, N1382, N543);
and AND2 (N3504, N3487, N1803);
nand NAND2 (N3505, N3500, N1343);
xor XOR2 (N3506, N3491, N874);
or OR4 (N3507, N3506, N3030, N947, N499);
nand NAND2 (N3508, N3507, N3409);
buf BUF1 (N3509, N3502);
not NOT1 (N3510, N3504);
buf BUF1 (N3511, N3494);
not NOT1 (N3512, N3508);
not NOT1 (N3513, N3499);
or OR4 (N3514, N3501, N215, N3059, N2170);
and AND3 (N3515, N3513, N2510, N55);
or OR3 (N3516, N3510, N168, N983);
and AND2 (N3517, N3509, N2939);
buf BUF1 (N3518, N3517);
not NOT1 (N3519, N3518);
buf BUF1 (N3520, N3519);
xor XOR2 (N3521, N3512, N818);
xor XOR2 (N3522, N3511, N1016);
and AND4 (N3523, N3497, N199, N3396, N2418);
xor XOR2 (N3524, N3516, N1378);
not NOT1 (N3525, N3523);
not NOT1 (N3526, N3524);
buf BUF1 (N3527, N3520);
not NOT1 (N3528, N3483);
or OR4 (N3529, N3505, N1365, N493, N293);
nand NAND4 (N3530, N3526, N418, N1357, N2315);
not NOT1 (N3531, N3530);
buf BUF1 (N3532, N3528);
buf BUF1 (N3533, N3529);
xor XOR2 (N3534, N3522, N1334);
nor NOR3 (N3535, N3533, N628, N367);
xor XOR2 (N3536, N3527, N948);
not NOT1 (N3537, N3515);
or OR4 (N3538, N3503, N190, N1393, N1318);
xor XOR2 (N3539, N3532, N869);
xor XOR2 (N3540, N3537, N2821);
not NOT1 (N3541, N3538);
buf BUF1 (N3542, N3514);
buf BUF1 (N3543, N3521);
buf BUF1 (N3544, N3525);
xor XOR2 (N3545, N3541, N337);
not NOT1 (N3546, N3545);
nand NAND2 (N3547, N3542, N3036);
not NOT1 (N3548, N3547);
nor NOR3 (N3549, N3544, N1941, N1096);
or OR4 (N3550, N3534, N128, N1711, N1689);
nor NOR4 (N3551, N3536, N1612, N121, N428);
not NOT1 (N3552, N3540);
and AND2 (N3553, N3531, N845);
or OR4 (N3554, N3550, N3423, N2544, N3294);
xor XOR2 (N3555, N3551, N2708);
or OR2 (N3556, N3549, N985);
xor XOR2 (N3557, N3546, N2636);
xor XOR2 (N3558, N3552, N1332);
not NOT1 (N3559, N3548);
nand NAND4 (N3560, N3559, N413, N181, N367);
xor XOR2 (N3561, N3539, N90);
nor NOR2 (N3562, N3557, N3474);
nand NAND2 (N3563, N3554, N1506);
nor NOR3 (N3564, N3543, N1161, N3350);
not NOT1 (N3565, N3535);
buf BUF1 (N3566, N3562);
nor NOR3 (N3567, N3561, N862, N7);
nor NOR3 (N3568, N3566, N1979, N1467);
nand NAND2 (N3569, N3568, N3454);
buf BUF1 (N3570, N3563);
xor XOR2 (N3571, N3564, N1770);
buf BUF1 (N3572, N3571);
buf BUF1 (N3573, N3572);
and AND4 (N3574, N3556, N2112, N805, N675);
or OR2 (N3575, N3570, N1200);
not NOT1 (N3576, N3574);
not NOT1 (N3577, N3553);
and AND3 (N3578, N3567, N1126, N1150);
not NOT1 (N3579, N3560);
nand NAND3 (N3580, N3558, N274, N2420);
xor XOR2 (N3581, N3565, N873);
and AND3 (N3582, N3555, N3548, N2931);
or OR4 (N3583, N3582, N2058, N1054, N2225);
not NOT1 (N3584, N3573);
or OR3 (N3585, N3577, N951, N716);
nor NOR4 (N3586, N3569, N3245, N2405, N2856);
xor XOR2 (N3587, N3575, N899);
and AND3 (N3588, N3579, N2182, N3484);
nor NOR4 (N3589, N3576, N46, N994, N2835);
or OR2 (N3590, N3587, N933);
nand NAND2 (N3591, N3584, N2854);
or OR3 (N3592, N3583, N692, N596);
xor XOR2 (N3593, N3588, N2019);
and AND4 (N3594, N3593, N1728, N159, N651);
and AND3 (N3595, N3589, N766, N1412);
and AND2 (N3596, N3580, N2466);
or OR3 (N3597, N3594, N447, N3054);
xor XOR2 (N3598, N3591, N3556);
nor NOR2 (N3599, N3578, N2883);
and AND3 (N3600, N3595, N1436, N3210);
xor XOR2 (N3601, N3597, N2977);
buf BUF1 (N3602, N3590);
not NOT1 (N3603, N3586);
nor NOR2 (N3604, N3585, N671);
or OR3 (N3605, N3601, N204, N1697);
xor XOR2 (N3606, N3605, N3328);
or OR3 (N3607, N3598, N2893, N3106);
xor XOR2 (N3608, N3599, N1048);
or OR3 (N3609, N3596, N2630, N2353);
buf BUF1 (N3610, N3602);
and AND2 (N3611, N3592, N2196);
or OR3 (N3612, N3604, N1660, N539);
not NOT1 (N3613, N3600);
buf BUF1 (N3614, N3606);
buf BUF1 (N3615, N3607);
not NOT1 (N3616, N3610);
nand NAND2 (N3617, N3609, N3041);
buf BUF1 (N3618, N3581);
and AND3 (N3619, N3611, N946, N2909);
or OR4 (N3620, N3608, N3456, N2110, N3472);
not NOT1 (N3621, N3619);
and AND2 (N3622, N3621, N2835);
buf BUF1 (N3623, N3620);
nand NAND4 (N3624, N3616, N447, N88, N1300);
or OR2 (N3625, N3622, N1142);
or OR3 (N3626, N3603, N2066, N3228);
and AND2 (N3627, N3612, N1778);
or OR2 (N3628, N3613, N2022);
nand NAND3 (N3629, N3628, N3617, N71);
nand NAND2 (N3630, N2797, N3107);
nand NAND2 (N3631, N3625, N2203);
or OR2 (N3632, N3630, N620);
and AND4 (N3633, N3618, N1459, N1128, N3066);
or OR3 (N3634, N3623, N3, N2730);
buf BUF1 (N3635, N3632);
buf BUF1 (N3636, N3627);
nor NOR2 (N3637, N3615, N654);
nor NOR2 (N3638, N3633, N1020);
nand NAND2 (N3639, N3624, N134);
not NOT1 (N3640, N3638);
xor XOR2 (N3641, N3640, N3245);
nor NOR2 (N3642, N3634, N3320);
not NOT1 (N3643, N3631);
nand NAND2 (N3644, N3641, N2514);
nand NAND2 (N3645, N3643, N680);
or OR3 (N3646, N3637, N1606, N1709);
nor NOR2 (N3647, N3635, N1080);
buf BUF1 (N3648, N3639);
not NOT1 (N3649, N3648);
and AND2 (N3650, N3649, N343);
or OR2 (N3651, N3646, N2064);
nor NOR2 (N3652, N3651, N1440);
xor XOR2 (N3653, N3645, N3544);
nand NAND4 (N3654, N3644, N2213, N2246, N2916);
or OR4 (N3655, N3614, N3463, N2388, N11);
nor NOR3 (N3656, N3647, N2164, N2465);
or OR4 (N3657, N3626, N1239, N662, N468);
nor NOR4 (N3658, N3636, N449, N87, N1524);
xor XOR2 (N3659, N3653, N1828);
nand NAND4 (N3660, N3650, N1058, N1612, N369);
nor NOR2 (N3661, N3658, N1524);
buf BUF1 (N3662, N3642);
buf BUF1 (N3663, N3654);
xor XOR2 (N3664, N3629, N2389);
not NOT1 (N3665, N3661);
nor NOR2 (N3666, N3663, N1542);
and AND3 (N3667, N3655, N1450, N361);
or OR2 (N3668, N3666, N2099);
xor XOR2 (N3669, N3668, N1548);
and AND2 (N3670, N3669, N3606);
and AND4 (N3671, N3660, N2654, N1035, N282);
not NOT1 (N3672, N3656);
nand NAND3 (N3673, N3657, N790, N3445);
nor NOR3 (N3674, N3662, N2282, N3630);
nor NOR2 (N3675, N3674, N3235);
and AND4 (N3676, N3665, N3106, N1958, N3403);
nor NOR4 (N3677, N3675, N993, N489, N3657);
and AND4 (N3678, N3667, N2948, N2544, N1077);
buf BUF1 (N3679, N3677);
and AND4 (N3680, N3664, N1668, N274, N2809);
and AND2 (N3681, N3652, N884);
nand NAND2 (N3682, N3670, N1);
and AND3 (N3683, N3680, N1562, N1476);
nand NAND2 (N3684, N3683, N1102);
or OR4 (N3685, N3659, N1270, N2902, N2537);
not NOT1 (N3686, N3679);
and AND2 (N3687, N3684, N732);
nand NAND2 (N3688, N3686, N103);
xor XOR2 (N3689, N3673, N2567);
or OR3 (N3690, N3689, N1112, N225);
nand NAND4 (N3691, N3687, N665, N703, N1389);
or OR3 (N3692, N3676, N535, N1017);
xor XOR2 (N3693, N3690, N2204);
or OR4 (N3694, N3681, N3432, N3040, N227);
nand NAND3 (N3695, N3694, N1586, N1855);
or OR4 (N3696, N3672, N326, N852, N1168);
nand NAND3 (N3697, N3696, N3138, N3695);
buf BUF1 (N3698, N463);
nand NAND3 (N3699, N3693, N410, N1606);
nand NAND4 (N3700, N3697, N3532, N1561, N558);
or OR2 (N3701, N3691, N642);
nor NOR2 (N3702, N3678, N1858);
nor NOR2 (N3703, N3685, N582);
not NOT1 (N3704, N3692);
not NOT1 (N3705, N3701);
or OR4 (N3706, N3702, N745, N529, N3065);
xor XOR2 (N3707, N3705, N2240);
nor NOR3 (N3708, N3699, N2005, N576);
buf BUF1 (N3709, N3704);
nor NOR2 (N3710, N3688, N815);
nor NOR3 (N3711, N3709, N2024, N79);
buf BUF1 (N3712, N3707);
buf BUF1 (N3713, N3682);
xor XOR2 (N3714, N3703, N729);
buf BUF1 (N3715, N3671);
not NOT1 (N3716, N3700);
and AND4 (N3717, N3716, N644, N2042, N165);
not NOT1 (N3718, N3715);
or OR4 (N3719, N3712, N1742, N3591, N348);
xor XOR2 (N3720, N3710, N2134);
buf BUF1 (N3721, N3719);
nor NOR2 (N3722, N3698, N555);
xor XOR2 (N3723, N3711, N3080);
and AND4 (N3724, N3708, N2593, N1224, N1762);
not NOT1 (N3725, N3718);
not NOT1 (N3726, N3723);
nand NAND2 (N3727, N3724, N3040);
buf BUF1 (N3728, N3722);
or OR2 (N3729, N3726, N2485);
and AND2 (N3730, N3717, N3133);
or OR4 (N3731, N3727, N2460, N311, N2976);
or OR2 (N3732, N3729, N2216);
or OR4 (N3733, N3714, N2791, N856, N2785);
nand NAND4 (N3734, N3730, N504, N2998, N1820);
xor XOR2 (N3735, N3732, N577);
and AND2 (N3736, N3725, N1428);
and AND3 (N3737, N3735, N1342, N3296);
nand NAND4 (N3738, N3733, N351, N1914, N3161);
not NOT1 (N3739, N3731);
nor NOR3 (N3740, N3734, N3275, N54);
buf BUF1 (N3741, N3728);
buf BUF1 (N3742, N3720);
and AND4 (N3743, N3742, N2039, N293, N2628);
xor XOR2 (N3744, N3706, N2058);
nor NOR4 (N3745, N3721, N3600, N2866, N1022);
buf BUF1 (N3746, N3744);
and AND2 (N3747, N3743, N3708);
nand NAND2 (N3748, N3739, N3331);
nor NOR4 (N3749, N3747, N139, N1650, N1544);
nor NOR3 (N3750, N3713, N983, N2284);
nor NOR2 (N3751, N3737, N285);
nand NAND3 (N3752, N3738, N3400, N1304);
nor NOR2 (N3753, N3736, N3752);
not NOT1 (N3754, N3613);
and AND2 (N3755, N3741, N101);
nor NOR3 (N3756, N3750, N1619, N2913);
not NOT1 (N3757, N3745);
and AND4 (N3758, N3746, N1182, N275, N2852);
and AND4 (N3759, N3757, N859, N1637, N1061);
xor XOR2 (N3760, N3748, N579);
buf BUF1 (N3761, N3749);
and AND3 (N3762, N3755, N3331, N2380);
or OR4 (N3763, N3761, N2145, N3132, N1612);
and AND2 (N3764, N3758, N1817);
buf BUF1 (N3765, N3762);
nand NAND4 (N3766, N3740, N809, N261, N1161);
not NOT1 (N3767, N3751);
xor XOR2 (N3768, N3753, N1734);
not NOT1 (N3769, N3764);
not NOT1 (N3770, N3756);
xor XOR2 (N3771, N3763, N3675);
buf BUF1 (N3772, N3771);
or OR2 (N3773, N3772, N3587);
not NOT1 (N3774, N3773);
and AND4 (N3775, N3774, N1418, N1675, N1168);
and AND3 (N3776, N3765, N332, N515);
nor NOR4 (N3777, N3770, N404, N2841, N939);
nand NAND3 (N3778, N3768, N1862, N1084);
nand NAND3 (N3779, N3759, N1519, N3133);
or OR3 (N3780, N3769, N3635, N1469);
xor XOR2 (N3781, N3754, N160);
not NOT1 (N3782, N3778);
nor NOR2 (N3783, N3782, N3146);
nand NAND3 (N3784, N3783, N708, N3116);
nand NAND3 (N3785, N3767, N435, N102);
nand NAND3 (N3786, N3784, N1982, N3574);
nand NAND2 (N3787, N3760, N1951);
xor XOR2 (N3788, N3779, N150);
not NOT1 (N3789, N3785);
nor NOR4 (N3790, N3777, N3264, N2106, N1729);
nand NAND2 (N3791, N3787, N3270);
or OR4 (N3792, N3776, N1405, N243, N408);
or OR3 (N3793, N3791, N1353, N1743);
or OR3 (N3794, N3780, N2932, N405);
or OR2 (N3795, N3766, N1327);
buf BUF1 (N3796, N3794);
or OR3 (N3797, N3775, N1390, N590);
nor NOR4 (N3798, N3781, N2874, N375, N1783);
buf BUF1 (N3799, N3792);
and AND2 (N3800, N3788, N1439);
buf BUF1 (N3801, N3798);
nor NOR4 (N3802, N3799, N2759, N1809, N2226);
nor NOR4 (N3803, N3786, N1215, N3305, N103);
nor NOR3 (N3804, N3800, N2227, N1701);
buf BUF1 (N3805, N3801);
or OR3 (N3806, N3802, N958, N213);
not NOT1 (N3807, N3789);
not NOT1 (N3808, N3795);
nand NAND4 (N3809, N3803, N2044, N3073, N3210);
nand NAND3 (N3810, N3796, N2068, N1680);
or OR4 (N3811, N3809, N3634, N534, N822);
not NOT1 (N3812, N3797);
or OR3 (N3813, N3812, N1862, N266);
not NOT1 (N3814, N3810);
nand NAND4 (N3815, N3808, N1463, N2897, N377);
nand NAND3 (N3816, N3814, N3015, N493);
and AND3 (N3817, N3815, N2489, N3774);
nand NAND2 (N3818, N3816, N2351);
xor XOR2 (N3819, N3818, N123);
or OR4 (N3820, N3806, N2084, N1011, N3311);
and AND4 (N3821, N3819, N3038, N2659, N3566);
not NOT1 (N3822, N3811);
buf BUF1 (N3823, N3804);
nand NAND2 (N3824, N3813, N2815);
buf BUF1 (N3825, N3821);
buf BUF1 (N3826, N3823);
or OR3 (N3827, N3817, N909, N1341);
xor XOR2 (N3828, N3825, N3280);
xor XOR2 (N3829, N3805, N626);
nor NOR2 (N3830, N3807, N2459);
nor NOR4 (N3831, N3829, N2566, N1170, N2771);
nor NOR3 (N3832, N3830, N2393, N2649);
buf BUF1 (N3833, N3793);
nor NOR4 (N3834, N3831, N3033, N423, N2981);
nor NOR4 (N3835, N3828, N805, N1835, N2404);
and AND3 (N3836, N3822, N2561, N2076);
nand NAND2 (N3837, N3835, N2880);
buf BUF1 (N3838, N3832);
buf BUF1 (N3839, N3833);
buf BUF1 (N3840, N3837);
nor NOR3 (N3841, N3840, N2409, N191);
or OR4 (N3842, N3838, N3571, N455, N1728);
nor NOR4 (N3843, N3834, N2206, N3694, N996);
not NOT1 (N3844, N3824);
nor NOR2 (N3845, N3820, N1061);
or OR4 (N3846, N3844, N2288, N3401, N3195);
nor NOR2 (N3847, N3841, N1532);
nor NOR4 (N3848, N3836, N2074, N1381, N2806);
not NOT1 (N3849, N3790);
not NOT1 (N3850, N3827);
nand NAND2 (N3851, N3849, N2425);
xor XOR2 (N3852, N3851, N574);
not NOT1 (N3853, N3847);
xor XOR2 (N3854, N3853, N1220);
buf BUF1 (N3855, N3850);
not NOT1 (N3856, N3843);
buf BUF1 (N3857, N3842);
xor XOR2 (N3858, N3856, N1389);
xor XOR2 (N3859, N3826, N3664);
and AND4 (N3860, N3858, N862, N1685, N507);
buf BUF1 (N3861, N3848);
nand NAND4 (N3862, N3857, N1129, N1100, N3409);
nor NOR4 (N3863, N3859, N1196, N2335, N258);
or OR3 (N3864, N3846, N756, N3002);
xor XOR2 (N3865, N3861, N1281);
buf BUF1 (N3866, N3854);
not NOT1 (N3867, N3852);
not NOT1 (N3868, N3865);
nor NOR2 (N3869, N3866, N1467);
or OR3 (N3870, N3845, N1249, N1070);
not NOT1 (N3871, N3839);
and AND4 (N3872, N3870, N2826, N2393, N2046);
nand NAND4 (N3873, N3860, N2004, N704, N1815);
buf BUF1 (N3874, N3873);
nand NAND4 (N3875, N3869, N3819, N1925, N3469);
and AND4 (N3876, N3874, N2665, N1262, N2770);
or OR2 (N3877, N3867, N1064);
not NOT1 (N3878, N3855);
buf BUF1 (N3879, N3872);
nor NOR3 (N3880, N3864, N798, N400);
and AND2 (N3881, N3880, N629);
xor XOR2 (N3882, N3879, N3546);
not NOT1 (N3883, N3876);
and AND4 (N3884, N3877, N3575, N256, N1850);
not NOT1 (N3885, N3862);
or OR3 (N3886, N3883, N2329, N699);
and AND2 (N3887, N3881, N2152);
xor XOR2 (N3888, N3886, N2625);
not NOT1 (N3889, N3868);
not NOT1 (N3890, N3889);
not NOT1 (N3891, N3884);
not NOT1 (N3892, N3888);
buf BUF1 (N3893, N3882);
buf BUF1 (N3894, N3863);
nor NOR4 (N3895, N3871, N1225, N3367, N315);
nor NOR2 (N3896, N3894, N3483);
nand NAND2 (N3897, N3892, N437);
not NOT1 (N3898, N3878);
buf BUF1 (N3899, N3895);
and AND4 (N3900, N3899, N243, N963, N2228);
not NOT1 (N3901, N3887);
or OR3 (N3902, N3885, N1651, N2550);
nand NAND3 (N3903, N3900, N3294, N1112);
nand NAND2 (N3904, N3891, N710);
not NOT1 (N3905, N3903);
and AND3 (N3906, N3896, N1562, N1713);
xor XOR2 (N3907, N3906, N3739);
or OR4 (N3908, N3901, N2782, N525, N3762);
xor XOR2 (N3909, N3902, N1027);
and AND4 (N3910, N3875, N1480, N3695, N1137);
nand NAND2 (N3911, N3898, N2323);
and AND4 (N3912, N3910, N3549, N727, N3455);
xor XOR2 (N3913, N3904, N2351);
nand NAND2 (N3914, N3893, N3134);
nor NOR2 (N3915, N3911, N3844);
nand NAND3 (N3916, N3897, N1197, N605);
nor NOR3 (N3917, N3909, N3478, N3482);
nor NOR2 (N3918, N3905, N271);
and AND3 (N3919, N3914, N1568, N1830);
or OR4 (N3920, N3919, N815, N3238, N1253);
nor NOR2 (N3921, N3890, N721);
and AND2 (N3922, N3907, N3344);
xor XOR2 (N3923, N3921, N2731);
or OR3 (N3924, N3923, N2273, N2032);
not NOT1 (N3925, N3916);
nor NOR4 (N3926, N3922, N1297, N2307, N2281);
xor XOR2 (N3927, N3908, N1588);
nor NOR2 (N3928, N3924, N3910);
nor NOR3 (N3929, N3917, N2792, N3042);
xor XOR2 (N3930, N3918, N3280);
and AND3 (N3931, N3926, N3858, N2989);
or OR2 (N3932, N3927, N1294);
and AND3 (N3933, N3913, N146, N3645);
buf BUF1 (N3934, N3920);
nor NOR4 (N3935, N3915, N1802, N3517, N2297);
buf BUF1 (N3936, N3935);
nor NOR3 (N3937, N3929, N1745, N198);
buf BUF1 (N3938, N3933);
nor NOR2 (N3939, N3934, N235);
and AND3 (N3940, N3912, N1573, N908);
or OR2 (N3941, N3940, N1183);
and AND2 (N3942, N3932, N518);
xor XOR2 (N3943, N3931, N69);
nand NAND2 (N3944, N3939, N1515);
xor XOR2 (N3945, N3925, N276);
not NOT1 (N3946, N3945);
xor XOR2 (N3947, N3928, N3796);
nor NOR2 (N3948, N3936, N2232);
buf BUF1 (N3949, N3947);
or OR2 (N3950, N3949, N986);
xor XOR2 (N3951, N3942, N3655);
and AND4 (N3952, N3948, N2328, N3714, N1117);
nor NOR4 (N3953, N3941, N3288, N262, N3324);
nand NAND3 (N3954, N3937, N2964, N1419);
xor XOR2 (N3955, N3950, N183);
not NOT1 (N3956, N3955);
and AND2 (N3957, N3954, N3570);
and AND3 (N3958, N3946, N1947, N1767);
buf BUF1 (N3959, N3952);
not NOT1 (N3960, N3956);
nor NOR4 (N3961, N3938, N558, N1917, N1841);
nand NAND4 (N3962, N3961, N3164, N800, N1698);
nor NOR2 (N3963, N3957, N2046);
not NOT1 (N3964, N3943);
and AND3 (N3965, N3953, N1315, N3711);
not NOT1 (N3966, N3963);
and AND4 (N3967, N3966, N551, N1063, N2222);
xor XOR2 (N3968, N3951, N3340);
and AND2 (N3969, N3958, N3393);
buf BUF1 (N3970, N3964);
xor XOR2 (N3971, N3959, N1012);
xor XOR2 (N3972, N3970, N2455);
xor XOR2 (N3973, N3965, N648);
and AND2 (N3974, N3930, N3406);
nor NOR3 (N3975, N3944, N3272, N1740);
not NOT1 (N3976, N3962);
and AND4 (N3977, N3976, N3113, N1471, N3960);
not NOT1 (N3978, N2261);
nand NAND2 (N3979, N3973, N322);
xor XOR2 (N3980, N3971, N2532);
or OR3 (N3981, N3975, N114, N671);
xor XOR2 (N3982, N3980, N2951);
nand NAND3 (N3983, N3979, N1527, N2866);
and AND2 (N3984, N3983, N978);
nand NAND3 (N3985, N3981, N1417, N3383);
xor XOR2 (N3986, N3969, N3861);
xor XOR2 (N3987, N3982, N863);
nor NOR4 (N3988, N3987, N530, N3805, N2285);
not NOT1 (N3989, N3977);
nand NAND3 (N3990, N3986, N1978, N3852);
nor NOR2 (N3991, N3978, N2969);
nor NOR2 (N3992, N3991, N908);
nor NOR3 (N3993, N3967, N3109, N3961);
xor XOR2 (N3994, N3993, N1833);
nor NOR3 (N3995, N3972, N260, N1864);
xor XOR2 (N3996, N3988, N75);
buf BUF1 (N3997, N3985);
buf BUF1 (N3998, N3992);
or OR2 (N3999, N3968, N582);
buf BUF1 (N4000, N3990);
not NOT1 (N4001, N3998);
not NOT1 (N4002, N3999);
xor XOR2 (N4003, N3997, N211);
or OR3 (N4004, N4003, N3816, N2504);
and AND4 (N4005, N3995, N881, N2043, N1046);
nand NAND4 (N4006, N4004, N3355, N2324, N805);
nor NOR4 (N4007, N4001, N347, N3359, N21);
and AND4 (N4008, N4007, N1822, N3637, N3854);
nand NAND4 (N4009, N3984, N2804, N3617, N2011);
xor XOR2 (N4010, N3994, N2296);
and AND3 (N4011, N3989, N3301, N1840);
nor NOR2 (N4012, N4011, N664);
and AND2 (N4013, N4009, N3810);
and AND3 (N4014, N3974, N2887, N3392);
and AND2 (N4015, N4013, N3699);
or OR2 (N4016, N4002, N3156);
nand NAND2 (N4017, N4015, N874);
and AND2 (N4018, N4006, N3075);
xor XOR2 (N4019, N4000, N3087);
buf BUF1 (N4020, N4014);
and AND3 (N4021, N4005, N2208, N2789);
or OR2 (N4022, N4018, N2758);
and AND4 (N4023, N3996, N1186, N658, N1831);
not NOT1 (N4024, N4023);
not NOT1 (N4025, N4022);
nor NOR2 (N4026, N4019, N795);
not NOT1 (N4027, N4010);
or OR3 (N4028, N4026, N32, N764);
and AND4 (N4029, N4016, N2769, N3950, N1170);
and AND2 (N4030, N4017, N2792);
xor XOR2 (N4031, N4024, N1859);
nor NOR2 (N4032, N4025, N1864);
xor XOR2 (N4033, N4020, N166);
or OR2 (N4034, N4031, N35);
and AND4 (N4035, N4021, N2447, N3881, N234);
not NOT1 (N4036, N4030);
or OR2 (N4037, N4027, N913);
nor NOR2 (N4038, N4036, N411);
not NOT1 (N4039, N4035);
xor XOR2 (N4040, N4038, N1631);
and AND3 (N4041, N4008, N638, N2387);
nor NOR4 (N4042, N4037, N3483, N2994, N747);
not NOT1 (N4043, N4028);
buf BUF1 (N4044, N4012);
or OR4 (N4045, N4039, N3587, N1638, N3448);
not NOT1 (N4046, N4043);
buf BUF1 (N4047, N4034);
nor NOR3 (N4048, N4044, N3528, N2453);
xor XOR2 (N4049, N4040, N228);
not NOT1 (N4050, N4049);
and AND2 (N4051, N4045, N136);
and AND4 (N4052, N4051, N294, N3064, N418);
nor NOR3 (N4053, N4033, N3807, N906);
buf BUF1 (N4054, N4050);
nand NAND3 (N4055, N4052, N482, N2384);
xor XOR2 (N4056, N4047, N1898);
and AND3 (N4057, N4041, N176, N2854);
and AND3 (N4058, N4042, N2378, N2950);
nor NOR4 (N4059, N4057, N1697, N887, N2419);
xor XOR2 (N4060, N4032, N1940);
xor XOR2 (N4061, N4046, N102);
nor NOR2 (N4062, N4029, N1354);
and AND2 (N4063, N4062, N415);
or OR2 (N4064, N4059, N1732);
or OR4 (N4065, N4054, N3428, N219, N49);
not NOT1 (N4066, N4064);
xor XOR2 (N4067, N4065, N4013);
not NOT1 (N4068, N4053);
nand NAND4 (N4069, N4066, N3490, N1928, N3442);
xor XOR2 (N4070, N4067, N1861);
nor NOR4 (N4071, N4061, N786, N3758, N3186);
or OR4 (N4072, N4048, N3061, N592, N3509);
and AND4 (N4073, N4068, N3003, N1276, N2062);
xor XOR2 (N4074, N4055, N2700);
or OR4 (N4075, N4063, N2598, N1228, N49);
nor NOR3 (N4076, N4069, N781, N2601);
nand NAND3 (N4077, N4074, N2142, N290);
nor NOR2 (N4078, N4058, N1258);
xor XOR2 (N4079, N4076, N792);
xor XOR2 (N4080, N4056, N59);
not NOT1 (N4081, N4070);
and AND2 (N4082, N4072, N2663);
nor NOR3 (N4083, N4071, N3616, N710);
and AND2 (N4084, N4073, N867);
not NOT1 (N4085, N4082);
not NOT1 (N4086, N4081);
not NOT1 (N4087, N4080);
nand NAND2 (N4088, N4060, N2246);
buf BUF1 (N4089, N4088);
buf BUF1 (N4090, N4084);
and AND4 (N4091, N4075, N560, N3126, N697);
nand NAND2 (N4092, N4077, N3754);
nor NOR2 (N4093, N4078, N3610);
buf BUF1 (N4094, N4093);
and AND4 (N4095, N4094, N2868, N1174, N1460);
nor NOR4 (N4096, N4095, N2461, N1651, N3777);
not NOT1 (N4097, N4090);
or OR2 (N4098, N4092, N3907);
xor XOR2 (N4099, N4083, N647);
buf BUF1 (N4100, N4087);
buf BUF1 (N4101, N4085);
or OR2 (N4102, N4079, N3243);
or OR2 (N4103, N4089, N2389);
and AND4 (N4104, N4098, N359, N3592, N2793);
nor NOR2 (N4105, N4103, N621);
nand NAND2 (N4106, N4091, N2047);
not NOT1 (N4107, N4099);
nand NAND2 (N4108, N4105, N174);
nor NOR4 (N4109, N4101, N1666, N2647, N196);
xor XOR2 (N4110, N4096, N759);
buf BUF1 (N4111, N4110);
nor NOR2 (N4112, N4104, N3535);
and AND4 (N4113, N4100, N2858, N1162, N640);
nand NAND4 (N4114, N4111, N2387, N2800, N3687);
nand NAND3 (N4115, N4113, N368, N713);
buf BUF1 (N4116, N4108);
xor XOR2 (N4117, N4109, N2532);
or OR4 (N4118, N4115, N1802, N1073, N3429);
or OR4 (N4119, N4116, N3241, N3321, N112);
nor NOR3 (N4120, N4112, N1112, N3549);
buf BUF1 (N4121, N4107);
and AND2 (N4122, N4114, N2115);
nor NOR2 (N4123, N4119, N1826);
xor XOR2 (N4124, N4097, N3737);
buf BUF1 (N4125, N4102);
buf BUF1 (N4126, N4086);
not NOT1 (N4127, N4126);
xor XOR2 (N4128, N4117, N3077);
nand NAND4 (N4129, N4122, N3649, N391, N2705);
xor XOR2 (N4130, N4121, N2944);
xor XOR2 (N4131, N4123, N3990);
or OR2 (N4132, N4127, N2563);
buf BUF1 (N4133, N4129);
and AND3 (N4134, N4118, N3180, N3669);
not NOT1 (N4135, N4130);
nand NAND3 (N4136, N4135, N2892, N447);
xor XOR2 (N4137, N4128, N885);
buf BUF1 (N4138, N4132);
and AND4 (N4139, N4125, N1532, N543, N3945);
and AND2 (N4140, N4137, N4123);
nor NOR2 (N4141, N4134, N2304);
nand NAND3 (N4142, N4136, N3470, N1170);
and AND4 (N4143, N4120, N1432, N1146, N1105);
nand NAND3 (N4144, N4141, N3889, N3090);
xor XOR2 (N4145, N4139, N2033);
not NOT1 (N4146, N4145);
xor XOR2 (N4147, N4138, N2890);
not NOT1 (N4148, N4131);
xor XOR2 (N4149, N4144, N349);
and AND4 (N4150, N4143, N427, N482, N3494);
or OR2 (N4151, N4133, N2019);
and AND3 (N4152, N4142, N3415, N1804);
nor NOR3 (N4153, N4146, N594, N2370);
xor XOR2 (N4154, N4124, N2820);
and AND2 (N4155, N4151, N167);
nor NOR2 (N4156, N4149, N2723);
and AND2 (N4157, N4147, N3674);
nor NOR4 (N4158, N4154, N475, N3587, N755);
not NOT1 (N4159, N4140);
xor XOR2 (N4160, N4148, N3819);
xor XOR2 (N4161, N4158, N3788);
nor NOR3 (N4162, N4155, N150, N4116);
nand NAND3 (N4163, N4106, N268, N760);
buf BUF1 (N4164, N4157);
buf BUF1 (N4165, N4162);
nand NAND2 (N4166, N4160, N2659);
and AND2 (N4167, N4165, N3563);
buf BUF1 (N4168, N4153);
nor NOR4 (N4169, N4161, N4018, N2036, N1031);
nand NAND3 (N4170, N4159, N258, N3419);
not NOT1 (N4171, N4152);
and AND4 (N4172, N4156, N2020, N3662, N3521);
nand NAND4 (N4173, N4163, N2742, N1246, N2723);
not NOT1 (N4174, N4166);
buf BUF1 (N4175, N4167);
xor XOR2 (N4176, N4175, N3202);
or OR4 (N4177, N4168, N2182, N3813, N307);
nand NAND3 (N4178, N4171, N2509, N3353);
nor NOR3 (N4179, N4170, N4135, N3146);
and AND4 (N4180, N4177, N4010, N2692, N3886);
nor NOR4 (N4181, N4172, N2821, N1550, N3623);
and AND2 (N4182, N4178, N1026);
nor NOR3 (N4183, N4176, N2113, N1001);
buf BUF1 (N4184, N4169);
buf BUF1 (N4185, N4183);
and AND2 (N4186, N4150, N2222);
xor XOR2 (N4187, N4174, N2856);
nor NOR2 (N4188, N4181, N3484);
not NOT1 (N4189, N4187);
and AND2 (N4190, N4189, N820);
not NOT1 (N4191, N4173);
not NOT1 (N4192, N4188);
and AND2 (N4193, N4184, N3653);
not NOT1 (N4194, N4185);
nor NOR2 (N4195, N4193, N422);
nor NOR3 (N4196, N4192, N3610, N1744);
xor XOR2 (N4197, N4194, N2114);
nand NAND4 (N4198, N4179, N3524, N775, N3508);
or OR2 (N4199, N4196, N1816);
nand NAND2 (N4200, N4180, N3827);
not NOT1 (N4201, N4198);
not NOT1 (N4202, N4186);
nand NAND3 (N4203, N4197, N3046, N2963);
nor NOR2 (N4204, N4195, N799);
or OR2 (N4205, N4200, N807);
nor NOR4 (N4206, N4203, N2024, N3649, N1184);
and AND2 (N4207, N4199, N2500);
nor NOR4 (N4208, N4182, N2895, N237, N2638);
not NOT1 (N4209, N4190);
nor NOR2 (N4210, N4204, N50);
nand NAND4 (N4211, N4191, N3249, N1121, N2250);
buf BUF1 (N4212, N4201);
nor NOR2 (N4213, N4207, N1348);
xor XOR2 (N4214, N4211, N1294);
xor XOR2 (N4215, N4210, N434);
xor XOR2 (N4216, N4212, N3166);
and AND3 (N4217, N4206, N2267, N595);
and AND2 (N4218, N4213, N2555);
xor XOR2 (N4219, N4214, N3152);
nand NAND3 (N4220, N4164, N3429, N1879);
nor NOR4 (N4221, N4215, N2684, N2284, N1271);
nand NAND2 (N4222, N4216, N3147);
buf BUF1 (N4223, N4217);
or OR4 (N4224, N4209, N2261, N3054, N2640);
nand NAND3 (N4225, N4220, N1260, N3063);
xor XOR2 (N4226, N4225, N1383);
xor XOR2 (N4227, N4221, N3960);
nand NAND2 (N4228, N4223, N1209);
or OR2 (N4229, N4218, N242);
or OR4 (N4230, N4208, N2799, N1023, N3378);
not NOT1 (N4231, N4202);
and AND4 (N4232, N4231, N1851, N1636, N3195);
not NOT1 (N4233, N4219);
buf BUF1 (N4234, N4229);
buf BUF1 (N4235, N4230);
and AND4 (N4236, N4222, N4133, N3282, N4039);
buf BUF1 (N4237, N4234);
buf BUF1 (N4238, N4237);
nand NAND2 (N4239, N4224, N3240);
and AND4 (N4240, N4235, N1541, N2138, N463);
xor XOR2 (N4241, N4228, N98);
or OR2 (N4242, N4227, N3032);
or OR4 (N4243, N4226, N456, N3736, N2880);
and AND3 (N4244, N4236, N1844, N4211);
buf BUF1 (N4245, N4232);
nor NOR3 (N4246, N4240, N1977, N2240);
not NOT1 (N4247, N4205);
or OR4 (N4248, N4239, N1704, N3000, N3768);
nand NAND3 (N4249, N4241, N1339, N4218);
and AND3 (N4250, N4243, N1774, N2380);
buf BUF1 (N4251, N4233);
not NOT1 (N4252, N4251);
buf BUF1 (N4253, N4238);
nand NAND3 (N4254, N4250, N1035, N883);
not NOT1 (N4255, N4245);
buf BUF1 (N4256, N4249);
buf BUF1 (N4257, N4248);
not NOT1 (N4258, N4257);
not NOT1 (N4259, N4258);
nand NAND4 (N4260, N4247, N276, N1770, N3868);
xor XOR2 (N4261, N4260, N1126);
and AND2 (N4262, N4259, N2003);
buf BUF1 (N4263, N4262);
and AND2 (N4264, N4242, N3370);
and AND2 (N4265, N4261, N2718);
buf BUF1 (N4266, N4265);
nand NAND3 (N4267, N4255, N4152, N2710);
not NOT1 (N4268, N4267);
nand NAND3 (N4269, N4254, N2962, N1556);
nand NAND4 (N4270, N4264, N875, N2929, N813);
buf BUF1 (N4271, N4266);
nand NAND2 (N4272, N4256, N424);
and AND2 (N4273, N4246, N137);
or OR3 (N4274, N4273, N2034, N2994);
and AND4 (N4275, N4244, N689, N2965, N2044);
buf BUF1 (N4276, N4268);
or OR4 (N4277, N4274, N3919, N1755, N715);
nand NAND4 (N4278, N4263, N2670, N3431, N1364);
nor NOR4 (N4279, N4276, N2497, N229, N2876);
not NOT1 (N4280, N4278);
nor NOR4 (N4281, N4252, N3902, N3154, N3993);
nand NAND2 (N4282, N4270, N260);
xor XOR2 (N4283, N4280, N2029);
or OR3 (N4284, N4275, N3373, N4057);
xor XOR2 (N4285, N4282, N2851);
xor XOR2 (N4286, N4253, N1387);
or OR3 (N4287, N4279, N1795, N2491);
buf BUF1 (N4288, N4285);
xor XOR2 (N4289, N4288, N4265);
or OR4 (N4290, N4277, N641, N3218, N4267);
xor XOR2 (N4291, N4283, N1168);
not NOT1 (N4292, N4289);
xor XOR2 (N4293, N4269, N1409);
xor XOR2 (N4294, N4292, N2578);
or OR4 (N4295, N4281, N3772, N3869, N2902);
xor XOR2 (N4296, N4284, N3902);
nor NOR3 (N4297, N4295, N1678, N403);
or OR4 (N4298, N4290, N3883, N2105, N944);
nor NOR3 (N4299, N4296, N1382, N4179);
xor XOR2 (N4300, N4272, N4030);
xor XOR2 (N4301, N4300, N3050);
not NOT1 (N4302, N4297);
and AND4 (N4303, N4294, N4130, N2240, N1080);
or OR4 (N4304, N4286, N3879, N1512, N355);
not NOT1 (N4305, N4291);
and AND2 (N4306, N4271, N3100);
nor NOR3 (N4307, N4306, N1731, N3562);
or OR3 (N4308, N4307, N4278, N443);
xor XOR2 (N4309, N4303, N1799);
nor NOR4 (N4310, N4298, N2078, N2380, N3534);
nand NAND4 (N4311, N4304, N4021, N148, N3642);
nand NAND2 (N4312, N4311, N1082);
and AND2 (N4313, N4293, N3332);
xor XOR2 (N4314, N4310, N2643);
nor NOR2 (N4315, N4312, N1153);
and AND2 (N4316, N4299, N3648);
xor XOR2 (N4317, N4302, N172);
or OR3 (N4318, N4316, N1319, N3743);
buf BUF1 (N4319, N4305);
xor XOR2 (N4320, N4317, N1899);
or OR2 (N4321, N4314, N4246);
xor XOR2 (N4322, N4321, N4013);
or OR3 (N4323, N4322, N1393, N2834);
and AND3 (N4324, N4320, N1998, N2662);
and AND3 (N4325, N4308, N1877, N866);
buf BUF1 (N4326, N4324);
and AND3 (N4327, N4287, N1466, N2633);
nand NAND3 (N4328, N4309, N1388, N824);
xor XOR2 (N4329, N4315, N924);
nand NAND3 (N4330, N4301, N2327, N1087);
and AND3 (N4331, N4319, N2685, N3128);
buf BUF1 (N4332, N4327);
and AND3 (N4333, N4332, N2013, N3680);
xor XOR2 (N4334, N4333, N4007);
nand NAND2 (N4335, N4325, N359);
nor NOR4 (N4336, N4326, N1229, N164, N2146);
and AND2 (N4337, N4329, N2123);
buf BUF1 (N4338, N4336);
not NOT1 (N4339, N4323);
nand NAND3 (N4340, N4335, N4221, N2021);
and AND3 (N4341, N4339, N327, N3497);
or OR2 (N4342, N4330, N1933);
or OR3 (N4343, N4340, N1268, N1030);
xor XOR2 (N4344, N4342, N3129);
not NOT1 (N4345, N4331);
nor NOR2 (N4346, N4337, N929);
buf BUF1 (N4347, N4318);
or OR3 (N4348, N4328, N2552, N29);
buf BUF1 (N4349, N4345);
not NOT1 (N4350, N4341);
xor XOR2 (N4351, N4349, N3351);
nor NOR4 (N4352, N4344, N1323, N3122, N2951);
or OR3 (N4353, N4343, N3309, N2450);
nor NOR2 (N4354, N4334, N3865);
buf BUF1 (N4355, N4353);
nand NAND4 (N4356, N4338, N206, N1117, N198);
or OR4 (N4357, N4313, N3221, N1242, N3370);
xor XOR2 (N4358, N4351, N983);
not NOT1 (N4359, N4350);
nand NAND3 (N4360, N4355, N427, N3668);
nor NOR2 (N4361, N4352, N804);
nor NOR2 (N4362, N4360, N874);
or OR3 (N4363, N4348, N770, N519);
nor NOR2 (N4364, N4363, N1844);
not NOT1 (N4365, N4359);
nand NAND3 (N4366, N4362, N956, N391);
or OR3 (N4367, N4347, N4005, N3127);
nor NOR3 (N4368, N4354, N1292, N4031);
nor NOR4 (N4369, N4366, N3697, N2940, N1751);
not NOT1 (N4370, N4367);
buf BUF1 (N4371, N4357);
or OR2 (N4372, N4365, N3046);
not NOT1 (N4373, N4361);
not NOT1 (N4374, N4373);
nor NOR4 (N4375, N4371, N1477, N671, N2433);
or OR2 (N4376, N4364, N1503);
xor XOR2 (N4377, N4372, N4017);
nor NOR3 (N4378, N4376, N3836, N183);
buf BUF1 (N4379, N4368);
nor NOR2 (N4380, N4346, N4136);
and AND4 (N4381, N4369, N2869, N741, N1200);
nand NAND4 (N4382, N4381, N649, N4101, N651);
xor XOR2 (N4383, N4377, N3246);
nand NAND4 (N4384, N4378, N1916, N4081, N4288);
not NOT1 (N4385, N4379);
nor NOR3 (N4386, N4356, N1753, N768);
nor NOR2 (N4387, N4358, N3678);
nor NOR4 (N4388, N4375, N1977, N2776, N2894);
buf BUF1 (N4389, N4384);
not NOT1 (N4390, N4380);
buf BUF1 (N4391, N4374);
nor NOR2 (N4392, N4370, N205);
nor NOR3 (N4393, N4385, N4127, N2349);
nand NAND4 (N4394, N4383, N703, N3112, N3253);
nand NAND3 (N4395, N4392, N4137, N299);
xor XOR2 (N4396, N4391, N2215);
and AND4 (N4397, N4393, N569, N4209, N891);
or OR3 (N4398, N4387, N1240, N3406);
and AND3 (N4399, N4398, N1026, N3445);
buf BUF1 (N4400, N4382);
buf BUF1 (N4401, N4386);
or OR3 (N4402, N4394, N4164, N487);
buf BUF1 (N4403, N4388);
nand NAND3 (N4404, N4396, N1958, N2854);
nand NAND2 (N4405, N4404, N2729);
xor XOR2 (N4406, N4389, N4362);
buf BUF1 (N4407, N4402);
nand NAND4 (N4408, N4400, N4208, N3157, N1826);
buf BUF1 (N4409, N4406);
and AND2 (N4410, N4390, N1825);
nor NOR3 (N4411, N4408, N966, N3709);
not NOT1 (N4412, N4410);
nand NAND2 (N4413, N4399, N1361);
not NOT1 (N4414, N4409);
and AND2 (N4415, N4411, N305);
not NOT1 (N4416, N4412);
not NOT1 (N4417, N4416);
or OR2 (N4418, N4397, N277);
xor XOR2 (N4419, N4405, N1916);
or OR4 (N4420, N4403, N4104, N2809, N3493);
and AND2 (N4421, N4413, N172);
and AND2 (N4422, N4415, N2798);
buf BUF1 (N4423, N4395);
buf BUF1 (N4424, N4421);
buf BUF1 (N4425, N4424);
nor NOR4 (N4426, N4425, N2317, N617, N219);
nor NOR3 (N4427, N4423, N2216, N184);
or OR4 (N4428, N4426, N3115, N3359, N414);
nor NOR4 (N4429, N4427, N24, N4285, N3777);
xor XOR2 (N4430, N4422, N1710);
xor XOR2 (N4431, N4418, N1110);
and AND2 (N4432, N4420, N1933);
buf BUF1 (N4433, N4401);
not NOT1 (N4434, N4433);
and AND3 (N4435, N4430, N309, N3189);
xor XOR2 (N4436, N4434, N4313);
nor NOR2 (N4437, N4431, N1588);
or OR2 (N4438, N4414, N1784);
not NOT1 (N4439, N4417);
nand NAND3 (N4440, N4419, N1253, N1188);
or OR2 (N4441, N4429, N1333);
nand NAND3 (N4442, N4435, N2469, N3788);
or OR3 (N4443, N4440, N1871, N2283);
xor XOR2 (N4444, N4438, N313);
nand NAND2 (N4445, N4444, N3562);
buf BUF1 (N4446, N4437);
and AND4 (N4447, N4445, N214, N2917, N2711);
nor NOR2 (N4448, N4436, N446);
nor NOR3 (N4449, N4448, N1160, N1650);
nand NAND3 (N4450, N4432, N1976, N1258);
buf BUF1 (N4451, N4450);
or OR4 (N4452, N4451, N750, N1868, N3900);
nor NOR3 (N4453, N4452, N3642, N1421);
xor XOR2 (N4454, N4439, N2834);
or OR2 (N4455, N4446, N469);
buf BUF1 (N4456, N4441);
xor XOR2 (N4457, N4456, N800);
and AND4 (N4458, N4447, N2828, N3214, N535);
not NOT1 (N4459, N4458);
buf BUF1 (N4460, N4443);
xor XOR2 (N4461, N4428, N695);
buf BUF1 (N4462, N4449);
not NOT1 (N4463, N4454);
buf BUF1 (N4464, N4442);
buf BUF1 (N4465, N4462);
or OR3 (N4466, N4457, N1165, N954);
or OR2 (N4467, N4465, N2913);
xor XOR2 (N4468, N4466, N1193);
nand NAND3 (N4469, N4467, N3295, N4224);
and AND4 (N4470, N4469, N1921, N1962, N4210);
and AND2 (N4471, N4460, N2518);
buf BUF1 (N4472, N4470);
buf BUF1 (N4473, N4453);
nor NOR2 (N4474, N4473, N3498);
buf BUF1 (N4475, N4455);
xor XOR2 (N4476, N4461, N3154);
nand NAND2 (N4477, N4459, N940);
buf BUF1 (N4478, N4463);
not NOT1 (N4479, N4478);
xor XOR2 (N4480, N4476, N1716);
xor XOR2 (N4481, N4407, N1637);
nand NAND4 (N4482, N4480, N3251, N2255, N1983);
buf BUF1 (N4483, N4481);
nor NOR4 (N4484, N4472, N2158, N2137, N1227);
and AND2 (N4485, N4484, N2543);
xor XOR2 (N4486, N4477, N3140);
xor XOR2 (N4487, N4485, N480);
not NOT1 (N4488, N4471);
nor NOR4 (N4489, N4486, N3713, N1380, N4036);
not NOT1 (N4490, N4482);
nor NOR2 (N4491, N4483, N2460);
xor XOR2 (N4492, N4487, N1372);
buf BUF1 (N4493, N4492);
buf BUF1 (N4494, N4489);
and AND2 (N4495, N4475, N4319);
and AND3 (N4496, N4491, N4406, N4338);
and AND4 (N4497, N4490, N3637, N4307, N3562);
not NOT1 (N4498, N4464);
nor NOR4 (N4499, N4496, N1201, N2327, N1355);
buf BUF1 (N4500, N4494);
and AND4 (N4501, N4468, N1679, N430, N1557);
nand NAND4 (N4502, N4493, N419, N3028, N782);
nor NOR2 (N4503, N4499, N2198);
and AND3 (N4504, N4474, N2147, N2663);
nand NAND3 (N4505, N4479, N1569, N3151);
and AND3 (N4506, N4502, N405, N4271);
buf BUF1 (N4507, N4488);
buf BUF1 (N4508, N4495);
and AND3 (N4509, N4504, N1989, N415);
nand NAND3 (N4510, N4497, N1178, N3021);
xor XOR2 (N4511, N4507, N1369);
and AND4 (N4512, N4511, N3316, N1595, N2791);
buf BUF1 (N4513, N4501);
not NOT1 (N4514, N4506);
xor XOR2 (N4515, N4508, N2324);
xor XOR2 (N4516, N4510, N3738);
not NOT1 (N4517, N4512);
or OR2 (N4518, N4513, N2972);
nor NOR3 (N4519, N4514, N1927, N2547);
buf BUF1 (N4520, N4503);
or OR3 (N4521, N4515, N1556, N146);
not NOT1 (N4522, N4519);
buf BUF1 (N4523, N4516);
xor XOR2 (N4524, N4517, N4256);
xor XOR2 (N4525, N4509, N1921);
xor XOR2 (N4526, N4518, N3192);
nor NOR2 (N4527, N4505, N1316);
buf BUF1 (N4528, N4500);
or OR2 (N4529, N4498, N2781);
not NOT1 (N4530, N4526);
xor XOR2 (N4531, N4527, N1489);
nand NAND3 (N4532, N4530, N2142, N391);
and AND2 (N4533, N4523, N764);
or OR3 (N4534, N4528, N732, N3779);
or OR4 (N4535, N4533, N3264, N3665, N2325);
buf BUF1 (N4536, N4521);
xor XOR2 (N4537, N4534, N1724);
nor NOR2 (N4538, N4536, N462);
buf BUF1 (N4539, N4524);
nand NAND2 (N4540, N4529, N3621);
and AND4 (N4541, N4525, N1211, N713, N2461);
or OR2 (N4542, N4537, N1926);
not NOT1 (N4543, N4532);
and AND4 (N4544, N4542, N4519, N3564, N1706);
xor XOR2 (N4545, N4539, N2154);
and AND2 (N4546, N4520, N4455);
and AND2 (N4547, N4541, N635);
or OR4 (N4548, N4531, N1613, N3293, N407);
xor XOR2 (N4549, N4522, N3653);
nor NOR4 (N4550, N4545, N2517, N2806, N2335);
nand NAND2 (N4551, N4547, N3738);
nor NOR3 (N4552, N4546, N2583, N4325);
not NOT1 (N4553, N4549);
xor XOR2 (N4554, N4543, N2335);
buf BUF1 (N4555, N4553);
xor XOR2 (N4556, N4552, N3699);
not NOT1 (N4557, N4555);
buf BUF1 (N4558, N4556);
not NOT1 (N4559, N4540);
nand NAND3 (N4560, N4558, N36, N3709);
buf BUF1 (N4561, N4551);
xor XOR2 (N4562, N4561, N2386);
xor XOR2 (N4563, N4559, N4014);
nand NAND4 (N4564, N4548, N342, N3700, N3913);
xor XOR2 (N4565, N4557, N2209);
buf BUF1 (N4566, N4563);
not NOT1 (N4567, N4564);
xor XOR2 (N4568, N4544, N3744);
xor XOR2 (N4569, N4538, N1909);
nor NOR2 (N4570, N4560, N3643);
and AND4 (N4571, N4566, N184, N4281, N3626);
and AND3 (N4572, N4567, N2726, N347);
or OR2 (N4573, N4572, N1182);
or OR4 (N4574, N4571, N590, N4441, N2534);
xor XOR2 (N4575, N4565, N1139);
not NOT1 (N4576, N4568);
or OR3 (N4577, N4554, N3453, N1883);
nand NAND3 (N4578, N4574, N658, N786);
xor XOR2 (N4579, N4578, N2595);
xor XOR2 (N4580, N4570, N3706);
not NOT1 (N4581, N4550);
not NOT1 (N4582, N4579);
nand NAND2 (N4583, N4582, N1273);
xor XOR2 (N4584, N4580, N2691);
or OR2 (N4585, N4584, N3454);
nand NAND3 (N4586, N4581, N2894, N1855);
not NOT1 (N4587, N4573);
xor XOR2 (N4588, N4562, N4029);
nand NAND4 (N4589, N4588, N811, N1047, N163);
buf BUF1 (N4590, N4535);
xor XOR2 (N4591, N4589, N218);
or OR2 (N4592, N4585, N2553);
and AND4 (N4593, N4569, N3882, N1367, N3945);
buf BUF1 (N4594, N4577);
buf BUF1 (N4595, N4583);
xor XOR2 (N4596, N4590, N2420);
nand NAND2 (N4597, N4596, N767);
buf BUF1 (N4598, N4587);
buf BUF1 (N4599, N4586);
buf BUF1 (N4600, N4598);
xor XOR2 (N4601, N4599, N1736);
or OR4 (N4602, N4600, N313, N3900, N1261);
xor XOR2 (N4603, N4602, N3437);
and AND3 (N4604, N4592, N817, N4165);
not NOT1 (N4605, N4594);
or OR4 (N4606, N4591, N3928, N1145, N604);
not NOT1 (N4607, N4603);
buf BUF1 (N4608, N4606);
not NOT1 (N4609, N4593);
buf BUF1 (N4610, N4576);
nand NAND2 (N4611, N4597, N1447);
and AND3 (N4612, N4601, N457, N434);
nand NAND2 (N4613, N4611, N2108);
nor NOR4 (N4614, N4605, N4326, N2842, N1100);
not NOT1 (N4615, N4604);
nand NAND2 (N4616, N4613, N1121);
nand NAND4 (N4617, N4575, N3889, N2338, N77);
or OR3 (N4618, N4607, N2969, N1142);
and AND2 (N4619, N4615, N2241);
or OR4 (N4620, N4609, N2239, N1910, N599);
or OR3 (N4621, N4612, N1546, N423);
and AND3 (N4622, N4617, N3436, N921);
xor XOR2 (N4623, N4595, N4201);
not NOT1 (N4624, N4622);
buf BUF1 (N4625, N4608);
or OR2 (N4626, N4620, N2265);
or OR4 (N4627, N4614, N3322, N2280, N514);
nor NOR2 (N4628, N4618, N1077);
or OR2 (N4629, N4621, N3428);
buf BUF1 (N4630, N4628);
or OR2 (N4631, N4630, N1836);
buf BUF1 (N4632, N4631);
buf BUF1 (N4633, N4610);
buf BUF1 (N4634, N4629);
and AND4 (N4635, N4624, N1937, N3219, N3186);
or OR3 (N4636, N4634, N1473, N4212);
or OR3 (N4637, N4616, N1926, N1368);
xor XOR2 (N4638, N4636, N2630);
nor NOR4 (N4639, N4637, N2208, N3305, N517);
xor XOR2 (N4640, N4632, N3692);
nand NAND4 (N4641, N4638, N2247, N1536, N4597);
and AND4 (N4642, N4626, N173, N2082, N634);
and AND3 (N4643, N4639, N2345, N2078);
and AND3 (N4644, N4635, N1146, N1259);
buf BUF1 (N4645, N4627);
not NOT1 (N4646, N4641);
nor NOR2 (N4647, N4644, N1393);
nand NAND4 (N4648, N4623, N1736, N2958, N425);
not NOT1 (N4649, N4643);
buf BUF1 (N4650, N4649);
xor XOR2 (N4651, N4633, N3398);
or OR3 (N4652, N4642, N4127, N174);
nor NOR4 (N4653, N4619, N2182, N654, N177);
not NOT1 (N4654, N4647);
buf BUF1 (N4655, N4625);
buf BUF1 (N4656, N4653);
and AND2 (N4657, N4652, N4635);
nand NAND2 (N4658, N4650, N852);
not NOT1 (N4659, N4656);
buf BUF1 (N4660, N4654);
xor XOR2 (N4661, N4657, N4158);
nor NOR3 (N4662, N4661, N3664, N2086);
or OR2 (N4663, N4645, N2838);
not NOT1 (N4664, N4655);
buf BUF1 (N4665, N4646);
nand NAND4 (N4666, N4664, N4044, N4291, N1359);
nand NAND2 (N4667, N4666, N2086);
and AND4 (N4668, N4663, N4266, N780, N4453);
nand NAND4 (N4669, N4667, N3922, N1163, N1666);
nand NAND3 (N4670, N4660, N2690, N3995);
and AND2 (N4671, N4670, N2733);
not NOT1 (N4672, N4658);
nand NAND3 (N4673, N4668, N570, N2103);
xor XOR2 (N4674, N4671, N1321);
not NOT1 (N4675, N4659);
xor XOR2 (N4676, N4674, N2781);
not NOT1 (N4677, N4651);
and AND4 (N4678, N4676, N930, N1507, N1923);
or OR2 (N4679, N4677, N2110);
not NOT1 (N4680, N4673);
xor XOR2 (N4681, N4665, N2860);
buf BUF1 (N4682, N4675);
nand NAND3 (N4683, N4680, N796, N8);
buf BUF1 (N4684, N4672);
and AND3 (N4685, N4648, N3403, N2468);
nor NOR2 (N4686, N4685, N1962);
buf BUF1 (N4687, N4678);
buf BUF1 (N4688, N4684);
not NOT1 (N4689, N4669);
and AND2 (N4690, N4681, N2774);
xor XOR2 (N4691, N4640, N3872);
nand NAND2 (N4692, N4689, N3911);
nor NOR3 (N4693, N4662, N2702, N4012);
buf BUF1 (N4694, N4688);
or OR2 (N4695, N4687, N1387);
and AND4 (N4696, N4692, N3747, N2954, N795);
buf BUF1 (N4697, N4693);
and AND3 (N4698, N4696, N1365, N3673);
not NOT1 (N4699, N4686);
nor NOR3 (N4700, N4699, N2712, N2265);
nor NOR3 (N4701, N4679, N1064, N2322);
not NOT1 (N4702, N4690);
xor XOR2 (N4703, N4697, N1250);
or OR3 (N4704, N4700, N4360, N2309);
xor XOR2 (N4705, N4682, N1935);
nand NAND3 (N4706, N4683, N1952, N1891);
xor XOR2 (N4707, N4698, N2728);
buf BUF1 (N4708, N4707);
buf BUF1 (N4709, N4695);
and AND4 (N4710, N4705, N1184, N3617, N1632);
buf BUF1 (N4711, N4691);
xor XOR2 (N4712, N4703, N4633);
not NOT1 (N4713, N4704);
buf BUF1 (N4714, N4702);
not NOT1 (N4715, N4713);
not NOT1 (N4716, N4715);
nor NOR4 (N4717, N4710, N123, N4102, N2948);
buf BUF1 (N4718, N4706);
xor XOR2 (N4719, N4717, N2650);
buf BUF1 (N4720, N4714);
xor XOR2 (N4721, N4694, N2521);
or OR4 (N4722, N4701, N4335, N2101, N3768);
buf BUF1 (N4723, N4711);
nand NAND4 (N4724, N4712, N1672, N614, N1002);
xor XOR2 (N4725, N4719, N3372);
not NOT1 (N4726, N4722);
xor XOR2 (N4727, N4724, N891);
and AND3 (N4728, N4708, N1196, N2755);
or OR4 (N4729, N4725, N1617, N3150, N2777);
or OR3 (N4730, N4720, N1330, N1152);
not NOT1 (N4731, N4709);
and AND2 (N4732, N4730, N1079);
and AND4 (N4733, N4718, N4681, N1876, N2048);
not NOT1 (N4734, N4727);
buf BUF1 (N4735, N4732);
xor XOR2 (N4736, N4716, N2019);
nor NOR2 (N4737, N4731, N2198);
nor NOR4 (N4738, N4728, N2585, N4650, N2658);
buf BUF1 (N4739, N4734);
and AND2 (N4740, N4726, N3800);
nor NOR2 (N4741, N4737, N1948);
xor XOR2 (N4742, N4735, N783);
not NOT1 (N4743, N4721);
or OR2 (N4744, N4736, N3897);
not NOT1 (N4745, N4738);
nor NOR2 (N4746, N4741, N4443);
or OR4 (N4747, N4740, N1375, N3891, N4468);
and AND4 (N4748, N4745, N2235, N3819, N3670);
nand NAND3 (N4749, N4747, N2994, N923);
or OR3 (N4750, N4739, N1132, N722);
or OR3 (N4751, N4748, N3335, N3107);
and AND2 (N4752, N4723, N4685);
xor XOR2 (N4753, N4749, N3793);
not NOT1 (N4754, N4742);
or OR2 (N4755, N4754, N21);
or OR2 (N4756, N4753, N2316);
nand NAND4 (N4757, N4744, N277, N679, N1361);
buf BUF1 (N4758, N4750);
buf BUF1 (N4759, N4729);
buf BUF1 (N4760, N4759);
and AND4 (N4761, N4758, N1149, N3215, N4074);
not NOT1 (N4762, N4757);
xor XOR2 (N4763, N4752, N4151);
or OR4 (N4764, N4756, N4499, N3659, N512);
not NOT1 (N4765, N4743);
xor XOR2 (N4766, N4746, N2080);
xor XOR2 (N4767, N4760, N1688);
buf BUF1 (N4768, N4733);
not NOT1 (N4769, N4765);
buf BUF1 (N4770, N4751);
buf BUF1 (N4771, N4755);
buf BUF1 (N4772, N4769);
not NOT1 (N4773, N4770);
not NOT1 (N4774, N4762);
buf BUF1 (N4775, N4764);
or OR4 (N4776, N4772, N3891, N2668, N2932);
or OR4 (N4777, N4776, N1480, N2097, N890);
not NOT1 (N4778, N4775);
and AND2 (N4779, N4766, N1207);
not NOT1 (N4780, N4768);
not NOT1 (N4781, N4780);
xor XOR2 (N4782, N4781, N3181);
buf BUF1 (N4783, N4771);
nand NAND2 (N4784, N4774, N561);
buf BUF1 (N4785, N4763);
buf BUF1 (N4786, N4784);
nand NAND4 (N4787, N4773, N2385, N2158, N247);
or OR3 (N4788, N4767, N111, N1733);
nand NAND3 (N4789, N4786, N1974, N283);
and AND4 (N4790, N4777, N3695, N4369, N3252);
buf BUF1 (N4791, N4789);
nand NAND2 (N4792, N4761, N457);
nand NAND2 (N4793, N4783, N4207);
nand NAND4 (N4794, N4785, N2117, N4592, N4483);
nand NAND4 (N4795, N4794, N252, N3992, N3510);
nand NAND3 (N4796, N4787, N4124, N4692);
or OR3 (N4797, N4795, N4584, N2348);
or OR3 (N4798, N4793, N3890, N232);
nor NOR2 (N4799, N4790, N3842);
and AND4 (N4800, N4779, N1189, N919, N1484);
nand NAND4 (N4801, N4800, N4115, N461, N2391);
buf BUF1 (N4802, N4791);
not NOT1 (N4803, N4796);
nor NOR4 (N4804, N4798, N2045, N3923, N4496);
or OR2 (N4805, N4801, N4215);
buf BUF1 (N4806, N4802);
xor XOR2 (N4807, N4799, N1535);
buf BUF1 (N4808, N4807);
not NOT1 (N4809, N4804);
buf BUF1 (N4810, N4809);
and AND2 (N4811, N4805, N1471);
buf BUF1 (N4812, N4808);
not NOT1 (N4813, N4792);
nor NOR4 (N4814, N4813, N1841, N778, N2105);
buf BUF1 (N4815, N4778);
not NOT1 (N4816, N4814);
and AND3 (N4817, N4811, N2158, N1533);
nor NOR2 (N4818, N4788, N2671);
buf BUF1 (N4819, N4815);
nand NAND2 (N4820, N4782, N1122);
buf BUF1 (N4821, N4816);
xor XOR2 (N4822, N4821, N596);
and AND4 (N4823, N4797, N4396, N605, N3437);
nor NOR2 (N4824, N4810, N574);
xor XOR2 (N4825, N4822, N582);
nor NOR2 (N4826, N4820, N4667);
and AND2 (N4827, N4826, N3715);
or OR3 (N4828, N4825, N2421, N1961);
nor NOR2 (N4829, N4817, N490);
nand NAND3 (N4830, N4829, N4359, N2137);
or OR4 (N4831, N4828, N4407, N3758, N2985);
not NOT1 (N4832, N4823);
xor XOR2 (N4833, N4803, N3601);
xor XOR2 (N4834, N4812, N2080);
and AND3 (N4835, N4806, N3957, N4358);
nor NOR2 (N4836, N4827, N2685);
nor NOR3 (N4837, N4819, N2869, N1197);
not NOT1 (N4838, N4831);
and AND2 (N4839, N4838, N3605);
nor NOR2 (N4840, N4834, N378);
and AND3 (N4841, N4835, N951, N4464);
nor NOR2 (N4842, N4837, N139);
xor XOR2 (N4843, N4836, N3433);
or OR2 (N4844, N4832, N3607);
and AND3 (N4845, N4841, N3902, N2252);
nor NOR3 (N4846, N4844, N3354, N4717);
xor XOR2 (N4847, N4830, N1229);
buf BUF1 (N4848, N4840);
not NOT1 (N4849, N4818);
buf BUF1 (N4850, N4839);
nor NOR4 (N4851, N4850, N785, N80, N2219);
nand NAND4 (N4852, N4847, N2959, N2817, N4010);
buf BUF1 (N4853, N4845);
buf BUF1 (N4854, N4833);
nor NOR2 (N4855, N4846, N4057);
xor XOR2 (N4856, N4854, N1491);
nor NOR2 (N4857, N4851, N4257);
nand NAND2 (N4858, N4852, N403);
or OR3 (N4859, N4853, N4736, N4442);
and AND4 (N4860, N4857, N1939, N4546, N3046);
buf BUF1 (N4861, N4849);
or OR2 (N4862, N4842, N736);
nand NAND2 (N4863, N4860, N4531);
xor XOR2 (N4864, N4861, N1367);
xor XOR2 (N4865, N4824, N2751);
nor NOR4 (N4866, N4848, N1261, N3544, N3349);
not NOT1 (N4867, N4866);
xor XOR2 (N4868, N4862, N2198);
not NOT1 (N4869, N4859);
nor NOR3 (N4870, N4843, N4867, N3161);
nand NAND3 (N4871, N2461, N1979, N4459);
and AND4 (N4872, N4856, N4790, N4190, N1904);
not NOT1 (N4873, N4871);
nor NOR2 (N4874, N4858, N4440);
buf BUF1 (N4875, N4864);
and AND4 (N4876, N4855, N1318, N214, N818);
nor NOR2 (N4877, N4863, N3259);
xor XOR2 (N4878, N4865, N2133);
or OR2 (N4879, N4869, N606);
or OR3 (N4880, N4876, N584, N2753);
nand NAND3 (N4881, N4873, N154, N2001);
nand NAND3 (N4882, N4872, N82, N2169);
nor NOR4 (N4883, N4882, N1731, N2118, N1791);
nand NAND4 (N4884, N4881, N2643, N2305, N1491);
or OR3 (N4885, N4880, N2653, N2424);
nor NOR2 (N4886, N4870, N2379);
not NOT1 (N4887, N4877);
or OR2 (N4888, N4878, N4628);
not NOT1 (N4889, N4887);
xor XOR2 (N4890, N4874, N97);
or OR2 (N4891, N4879, N2160);
or OR4 (N4892, N4875, N3645, N3292, N864);
xor XOR2 (N4893, N4885, N4027);
buf BUF1 (N4894, N4892);
not NOT1 (N4895, N4889);
or OR2 (N4896, N4893, N2089);
buf BUF1 (N4897, N4891);
xor XOR2 (N4898, N4883, N644);
and AND3 (N4899, N4896, N4574, N1253);
buf BUF1 (N4900, N4897);
or OR3 (N4901, N4900, N3930, N3303);
nor NOR3 (N4902, N4899, N987, N2309);
buf BUF1 (N4903, N4894);
not NOT1 (N4904, N4901);
not NOT1 (N4905, N4886);
or OR3 (N4906, N4902, N1114, N1950);
buf BUF1 (N4907, N4898);
not NOT1 (N4908, N4895);
and AND4 (N4909, N4888, N696, N4043, N523);
xor XOR2 (N4910, N4868, N2539);
buf BUF1 (N4911, N4908);
nand NAND4 (N4912, N4907, N1899, N3176, N3733);
or OR3 (N4913, N4905, N3695, N4220);
nand NAND2 (N4914, N4890, N3639);
buf BUF1 (N4915, N4903);
and AND2 (N4916, N4909, N4309);
or OR3 (N4917, N4904, N3376, N1931);
and AND4 (N4918, N4917, N2532, N3341, N1229);
not NOT1 (N4919, N4915);
nor NOR4 (N4920, N4916, N900, N1174, N4598);
buf BUF1 (N4921, N4914);
or OR3 (N4922, N4910, N51, N1566);
not NOT1 (N4923, N4922);
nor NOR2 (N4924, N4911, N2034);
and AND3 (N4925, N4913, N1694, N4882);
nor NOR4 (N4926, N4924, N3013, N4693, N4284);
buf BUF1 (N4927, N4925);
xor XOR2 (N4928, N4919, N240);
and AND2 (N4929, N4928, N3809);
xor XOR2 (N4930, N4926, N1006);
nand NAND4 (N4931, N4921, N3406, N4595, N1799);
nand NAND2 (N4932, N4930, N2512);
buf BUF1 (N4933, N4929);
and AND3 (N4934, N4933, N3302, N611);
nand NAND2 (N4935, N4906, N4364);
or OR2 (N4936, N4912, N3945);
xor XOR2 (N4937, N4920, N1378);
nand NAND2 (N4938, N4884, N3160);
xor XOR2 (N4939, N4927, N4209);
not NOT1 (N4940, N4936);
and AND4 (N4941, N4918, N1770, N550, N146);
and AND2 (N4942, N4937, N2401);
and AND4 (N4943, N4931, N115, N2978, N4460);
and AND2 (N4944, N4942, N3381);
not NOT1 (N4945, N4940);
not NOT1 (N4946, N4934);
or OR4 (N4947, N4923, N4545, N4243, N1882);
buf BUF1 (N4948, N4944);
nand NAND3 (N4949, N4945, N4656, N3562);
buf BUF1 (N4950, N4946);
buf BUF1 (N4951, N4939);
and AND4 (N4952, N4932, N1024, N1367, N359);
xor XOR2 (N4953, N4943, N1123);
buf BUF1 (N4954, N4950);
xor XOR2 (N4955, N4938, N4402);
buf BUF1 (N4956, N4948);
and AND2 (N4957, N4953, N3502);
and AND4 (N4958, N4941, N1659, N3449, N176);
nand NAND2 (N4959, N4935, N773);
nand NAND3 (N4960, N4958, N1352, N1364);
or OR3 (N4961, N4951, N3361, N4600);
or OR2 (N4962, N4957, N2479);
and AND3 (N4963, N4962, N1064, N539);
not NOT1 (N4964, N4960);
xor XOR2 (N4965, N4963, N3656);
not NOT1 (N4966, N4952);
or OR3 (N4967, N4959, N1816, N2743);
and AND4 (N4968, N4949, N2924, N2233, N3982);
buf BUF1 (N4969, N4961);
or OR4 (N4970, N4955, N964, N2394, N2196);
xor XOR2 (N4971, N4954, N1156);
buf BUF1 (N4972, N4970);
xor XOR2 (N4973, N4968, N4957);
buf BUF1 (N4974, N4967);
nor NOR4 (N4975, N4964, N4177, N4315, N919);
buf BUF1 (N4976, N4956);
nor NOR3 (N4977, N4976, N3916, N2125);
nand NAND3 (N4978, N4965, N2260, N4406);
not NOT1 (N4979, N4977);
buf BUF1 (N4980, N4974);
buf BUF1 (N4981, N4978);
nand NAND2 (N4982, N4966, N1652);
not NOT1 (N4983, N4973);
nand NAND4 (N4984, N4983, N1308, N2747, N2901);
not NOT1 (N4985, N4980);
buf BUF1 (N4986, N4984);
not NOT1 (N4987, N4981);
xor XOR2 (N4988, N4947, N1079);
not NOT1 (N4989, N4972);
nand NAND4 (N4990, N4985, N525, N2539, N1323);
or OR3 (N4991, N4986, N2291, N2140);
not NOT1 (N4992, N4988);
xor XOR2 (N4993, N4991, N1745);
xor XOR2 (N4994, N4992, N3923);
xor XOR2 (N4995, N4979, N2338);
nand NAND3 (N4996, N4975, N3587, N4061);
not NOT1 (N4997, N4971);
buf BUF1 (N4998, N4987);
nand NAND2 (N4999, N4969, N3983);
nor NOR4 (N5000, N4996, N1316, N4522, N431);
or OR4 (N5001, N4990, N2302, N24, N1533);
nor NOR3 (N5002, N4999, N1348, N4012);
nor NOR3 (N5003, N4995, N4629, N171);
nor NOR4 (N5004, N5000, N4622, N4136, N1949);
not NOT1 (N5005, N4989);
and AND2 (N5006, N5003, N4896);
nor NOR3 (N5007, N5002, N1334, N3078);
nand NAND3 (N5008, N5001, N2649, N4555);
nand NAND4 (N5009, N5004, N4487, N4968, N2617);
not NOT1 (N5010, N4998);
not NOT1 (N5011, N5006);
buf BUF1 (N5012, N5005);
nor NOR3 (N5013, N5010, N3920, N1901);
xor XOR2 (N5014, N4993, N3536);
buf BUF1 (N5015, N5011);
nor NOR4 (N5016, N5013, N3466, N3895, N1423);
buf BUF1 (N5017, N5014);
and AND2 (N5018, N5015, N2065);
not NOT1 (N5019, N5007);
xor XOR2 (N5020, N4997, N4838);
and AND3 (N5021, N5019, N3011, N4113);
xor XOR2 (N5022, N5012, N4737);
xor XOR2 (N5023, N5020, N328);
not NOT1 (N5024, N4994);
buf BUF1 (N5025, N5008);
nor NOR2 (N5026, N5025, N1670);
and AND2 (N5027, N5009, N3690);
or OR4 (N5028, N5024, N2831, N4266, N1879);
xor XOR2 (N5029, N5022, N1716);
not NOT1 (N5030, N5029);
and AND4 (N5031, N5018, N3636, N3196, N4102);
nand NAND2 (N5032, N5030, N3256);
xor XOR2 (N5033, N4982, N3939);
and AND2 (N5034, N5017, N1956);
and AND3 (N5035, N5023, N4352, N1391);
xor XOR2 (N5036, N5026, N1970);
not NOT1 (N5037, N5031);
or OR2 (N5038, N5027, N1830);
and AND3 (N5039, N5028, N2000, N928);
xor XOR2 (N5040, N5038, N2452);
not NOT1 (N5041, N5039);
not NOT1 (N5042, N5021);
nand NAND3 (N5043, N5041, N907, N2967);
and AND2 (N5044, N5043, N2684);
not NOT1 (N5045, N5016);
or OR4 (N5046, N5040, N1974, N2860, N3);
nor NOR3 (N5047, N5037, N2319, N3856);
xor XOR2 (N5048, N5045, N3775);
nand NAND2 (N5049, N5047, N3467);
nor NOR4 (N5050, N5049, N4085, N394, N4437);
buf BUF1 (N5051, N5034);
not NOT1 (N5052, N5036);
and AND4 (N5053, N5044, N4473, N2573, N4557);
not NOT1 (N5054, N5048);
or OR4 (N5055, N5052, N960, N3472, N390);
or OR4 (N5056, N5053, N5043, N2659, N3873);
nand NAND2 (N5057, N5042, N1995);
buf BUF1 (N5058, N5054);
or OR2 (N5059, N5046, N4401);
not NOT1 (N5060, N5057);
buf BUF1 (N5061, N5035);
xor XOR2 (N5062, N5056, N458);
not NOT1 (N5063, N5061);
nand NAND3 (N5064, N5058, N3888, N4738);
not NOT1 (N5065, N5032);
xor XOR2 (N5066, N5059, N3467);
not NOT1 (N5067, N5055);
or OR2 (N5068, N5033, N3946);
xor XOR2 (N5069, N5065, N746);
buf BUF1 (N5070, N5069);
and AND4 (N5071, N5063, N1580, N4335, N1687);
or OR3 (N5072, N5050, N3450, N1392);
buf BUF1 (N5073, N5068);
and AND3 (N5074, N5070, N4385, N1957);
buf BUF1 (N5075, N5060);
nand NAND3 (N5076, N5062, N554, N611);
nand NAND2 (N5077, N5076, N1606);
nor NOR4 (N5078, N5066, N571, N897, N3461);
or OR3 (N5079, N5073, N3037, N4359);
buf BUF1 (N5080, N5051);
nand NAND4 (N5081, N5067, N4082, N459, N1655);
nor NOR3 (N5082, N5064, N617, N274);
nor NOR2 (N5083, N5078, N1680);
xor XOR2 (N5084, N5072, N845);
not NOT1 (N5085, N5082);
xor XOR2 (N5086, N5085, N19);
or OR3 (N5087, N5075, N4508, N3320);
or OR3 (N5088, N5074, N2243, N1836);
buf BUF1 (N5089, N5087);
nand NAND4 (N5090, N5081, N1031, N2571, N3116);
xor XOR2 (N5091, N5083, N4472);
xor XOR2 (N5092, N5084, N4883);
nor NOR3 (N5093, N5089, N4609, N76);
xor XOR2 (N5094, N5088, N413);
and AND4 (N5095, N5077, N4570, N2446, N2398);
not NOT1 (N5096, N5079);
nor NOR4 (N5097, N5086, N4163, N1371, N1169);
or OR2 (N5098, N5095, N1785);
nor NOR2 (N5099, N5097, N4951);
buf BUF1 (N5100, N5098);
or OR3 (N5101, N5094, N55, N3175);
nor NOR4 (N5102, N5080, N3871, N3189, N1332);
nand NAND4 (N5103, N5090, N4413, N2027, N411);
nor NOR3 (N5104, N5103, N817, N4582);
nor NOR3 (N5105, N5092, N1468, N3151);
not NOT1 (N5106, N5100);
nor NOR3 (N5107, N5105, N1568, N1023);
or OR2 (N5108, N5096, N337);
or OR4 (N5109, N5107, N2599, N4562, N2218);
nor NOR4 (N5110, N5108, N3236, N3347, N4413);
buf BUF1 (N5111, N5102);
or OR2 (N5112, N5104, N1246);
nand NAND3 (N5113, N5093, N3365, N2207);
xor XOR2 (N5114, N5112, N1701);
xor XOR2 (N5115, N5099, N2156);
or OR4 (N5116, N5114, N4402, N5003, N2802);
or OR4 (N5117, N5113, N2897, N2521, N4709);
xor XOR2 (N5118, N5091, N3034);
nand NAND3 (N5119, N5115, N86, N526);
nand NAND3 (N5120, N5106, N2211, N4306);
nand NAND4 (N5121, N5118, N3687, N3769, N1072);
nand NAND2 (N5122, N5101, N731);
and AND4 (N5123, N5110, N3486, N3232, N1327);
and AND3 (N5124, N5120, N1851, N1313);
and AND2 (N5125, N5124, N4043);
not NOT1 (N5126, N5119);
xor XOR2 (N5127, N5123, N4964);
xor XOR2 (N5128, N5127, N384);
nor NOR2 (N5129, N5071, N2003);
and AND4 (N5130, N5109, N3804, N3676, N1085);
buf BUF1 (N5131, N5121);
xor XOR2 (N5132, N5130, N2400);
or OR3 (N5133, N5126, N2420, N2462);
buf BUF1 (N5134, N5117);
nand NAND3 (N5135, N5116, N3607, N4151);
nor NOR2 (N5136, N5131, N2672);
xor XOR2 (N5137, N5111, N849);
xor XOR2 (N5138, N5133, N932);
not NOT1 (N5139, N5138);
not NOT1 (N5140, N5132);
buf BUF1 (N5141, N5134);
or OR2 (N5142, N5137, N2094);
or OR2 (N5143, N5122, N2998);
buf BUF1 (N5144, N5125);
or OR4 (N5145, N5141, N207, N2215, N1674);
nor NOR2 (N5146, N5139, N2797);
or OR4 (N5147, N5144, N4799, N1299, N2533);
and AND3 (N5148, N5136, N2037, N2713);
buf BUF1 (N5149, N5145);
nor NOR4 (N5150, N5143, N1210, N3339, N3484);
or OR2 (N5151, N5147, N5100);
nor NOR4 (N5152, N5150, N808, N4890, N1155);
or OR4 (N5153, N5142, N3923, N2635, N2144);
buf BUF1 (N5154, N5148);
nand NAND2 (N5155, N5152, N256);
not NOT1 (N5156, N5128);
nand NAND4 (N5157, N5140, N2574, N2009, N897);
nor NOR3 (N5158, N5146, N3955, N3152);
xor XOR2 (N5159, N5158, N5114);
not NOT1 (N5160, N5156);
buf BUF1 (N5161, N5160);
buf BUF1 (N5162, N5135);
or OR4 (N5163, N5151, N4938, N61, N4530);
xor XOR2 (N5164, N5162, N2599);
nand NAND2 (N5165, N5155, N359);
and AND3 (N5166, N5164, N2409, N1583);
not NOT1 (N5167, N5153);
not NOT1 (N5168, N5154);
xor XOR2 (N5169, N5166, N4925);
or OR2 (N5170, N5165, N3066);
or OR2 (N5171, N5167, N2677);
not NOT1 (N5172, N5163);
nor NOR3 (N5173, N5168, N2323, N1557);
and AND2 (N5174, N5172, N2815);
buf BUF1 (N5175, N5170);
and AND3 (N5176, N5157, N4127, N1821);
or OR2 (N5177, N5129, N2273);
buf BUF1 (N5178, N5169);
buf BUF1 (N5179, N5174);
and AND4 (N5180, N5179, N5169, N1743, N4802);
xor XOR2 (N5181, N5173, N3765);
xor XOR2 (N5182, N5149, N1360);
and AND4 (N5183, N5178, N2515, N3515, N3864);
nor NOR4 (N5184, N5181, N4089, N1539, N4578);
xor XOR2 (N5185, N5176, N1439);
nand NAND2 (N5186, N5185, N1254);
and AND4 (N5187, N5182, N3261, N2324, N936);
buf BUF1 (N5188, N5183);
or OR4 (N5189, N5175, N3465, N845, N2138);
or OR4 (N5190, N5189, N5148, N2766, N4340);
and AND4 (N5191, N5190, N4474, N2819, N3306);
xor XOR2 (N5192, N5161, N2836);
nand NAND2 (N5193, N5188, N5123);
nand NAND2 (N5194, N5187, N4813);
nand NAND2 (N5195, N5171, N1769);
not NOT1 (N5196, N5193);
xor XOR2 (N5197, N5186, N1327);
or OR2 (N5198, N5197, N1071);
xor XOR2 (N5199, N5194, N2803);
nand NAND3 (N5200, N5199, N4967, N5167);
and AND2 (N5201, N5196, N2579);
nor NOR3 (N5202, N5177, N4153, N2151);
or OR2 (N5203, N5192, N1698);
buf BUF1 (N5204, N5200);
nand NAND3 (N5205, N5180, N3461, N3743);
buf BUF1 (N5206, N5203);
not NOT1 (N5207, N5184);
or OR3 (N5208, N5206, N1446, N1269);
nand NAND3 (N5209, N5191, N2074, N4212);
xor XOR2 (N5210, N5207, N4231);
xor XOR2 (N5211, N5210, N3114);
and AND2 (N5212, N5201, N2835);
nand NAND2 (N5213, N5195, N4987);
nand NAND3 (N5214, N5211, N175, N4901);
and AND2 (N5215, N5214, N3505);
not NOT1 (N5216, N5213);
not NOT1 (N5217, N5198);
or OR3 (N5218, N5212, N3779, N1206);
and AND4 (N5219, N5159, N1175, N1112, N1779);
nand NAND2 (N5220, N5219, N2942);
nor NOR2 (N5221, N5205, N4048);
and AND2 (N5222, N5208, N1898);
nand NAND2 (N5223, N5218, N4533);
or OR4 (N5224, N5223, N1948, N4128, N2461);
nor NOR3 (N5225, N5202, N1430, N3933);
or OR4 (N5226, N5215, N4241, N2517, N3868);
nor NOR3 (N5227, N5226, N511, N4767);
or OR3 (N5228, N5216, N1668, N1426);
nor NOR4 (N5229, N5222, N682, N4719, N2073);
or OR4 (N5230, N5209, N3939, N3136, N4052);
or OR4 (N5231, N5220, N4837, N4812, N4117);
and AND3 (N5232, N5217, N876, N1872);
buf BUF1 (N5233, N5224);
nor NOR2 (N5234, N5231, N1589);
nor NOR2 (N5235, N5227, N3613);
buf BUF1 (N5236, N5234);
and AND3 (N5237, N5230, N3843, N1963);
nand NAND4 (N5238, N5233, N2912, N3385, N990);
buf BUF1 (N5239, N5232);
not NOT1 (N5240, N5228);
buf BUF1 (N5241, N5221);
nor NOR4 (N5242, N5229, N913, N2105, N1622);
not NOT1 (N5243, N5240);
or OR3 (N5244, N5237, N4693, N4052);
or OR3 (N5245, N5243, N995, N3812);
buf BUF1 (N5246, N5225);
nor NOR3 (N5247, N5235, N3702, N3117);
or OR2 (N5248, N5244, N4197);
nand NAND2 (N5249, N5247, N1579);
nand NAND3 (N5250, N5248, N706, N4840);
xor XOR2 (N5251, N5250, N3990);
xor XOR2 (N5252, N5242, N5070);
and AND2 (N5253, N5238, N1155);
xor XOR2 (N5254, N5245, N3383);
and AND2 (N5255, N5253, N3831);
not NOT1 (N5256, N5255);
xor XOR2 (N5257, N5204, N5194);
buf BUF1 (N5258, N5236);
and AND4 (N5259, N5251, N2093, N4483, N4028);
buf BUF1 (N5260, N5259);
and AND4 (N5261, N5254, N4278, N940, N3605);
or OR4 (N5262, N5256, N4833, N2563, N4739);
xor XOR2 (N5263, N5249, N614);
not NOT1 (N5264, N5252);
not NOT1 (N5265, N5261);
nor NOR2 (N5266, N5246, N4463);
and AND3 (N5267, N5262, N821, N4435);
and AND2 (N5268, N5264, N53);
nand NAND2 (N5269, N5267, N5248);
buf BUF1 (N5270, N5241);
and AND2 (N5271, N5269, N1171);
or OR3 (N5272, N5257, N4011, N3619);
not NOT1 (N5273, N5260);
nor NOR2 (N5274, N5266, N4091);
nand NAND2 (N5275, N5268, N1198);
nor NOR2 (N5276, N5274, N402);
or OR3 (N5277, N5275, N3894, N3120);
nand NAND2 (N5278, N5270, N1848);
xor XOR2 (N5279, N5276, N1829);
buf BUF1 (N5280, N5277);
buf BUF1 (N5281, N5239);
nor NOR3 (N5282, N5272, N3677, N1584);
or OR3 (N5283, N5280, N4756, N540);
and AND4 (N5284, N5279, N3896, N2685, N1860);
nand NAND3 (N5285, N5281, N1593, N1043);
and AND3 (N5286, N5273, N4938, N5283);
buf BUF1 (N5287, N2544);
nand NAND4 (N5288, N5265, N494, N191, N3979);
buf BUF1 (N5289, N5286);
or OR4 (N5290, N5258, N2185, N3380, N3789);
or OR4 (N5291, N5285, N1247, N3440, N1923);
and AND2 (N5292, N5287, N4414);
not NOT1 (N5293, N5290);
buf BUF1 (N5294, N5288);
xor XOR2 (N5295, N5294, N1923);
and AND3 (N5296, N5284, N4671, N2758);
or OR2 (N5297, N5292, N5024);
nor NOR3 (N5298, N5289, N5260, N1895);
buf BUF1 (N5299, N5282);
and AND3 (N5300, N5291, N4924, N1562);
buf BUF1 (N5301, N5295);
not NOT1 (N5302, N5301);
nor NOR3 (N5303, N5297, N189, N1128);
not NOT1 (N5304, N5263);
buf BUF1 (N5305, N5296);
nor NOR2 (N5306, N5300, N253);
nor NOR2 (N5307, N5293, N3831);
and AND3 (N5308, N5302, N1316, N211);
nand NAND4 (N5309, N5298, N4339, N1751, N5115);
or OR4 (N5310, N5306, N5124, N1387, N3157);
buf BUF1 (N5311, N5308);
nor NOR4 (N5312, N5278, N674, N275, N1981);
or OR2 (N5313, N5312, N4480);
or OR3 (N5314, N5309, N3650, N4825);
buf BUF1 (N5315, N5313);
nor NOR3 (N5316, N5310, N4151, N1441);
xor XOR2 (N5317, N5314, N2106);
not NOT1 (N5318, N5317);
xor XOR2 (N5319, N5307, N1088);
nor NOR2 (N5320, N5305, N1106);
nor NOR2 (N5321, N5318, N2726);
nand NAND3 (N5322, N5315, N3957, N3555);
or OR4 (N5323, N5322, N3775, N794, N192);
and AND2 (N5324, N5316, N3252);
or OR2 (N5325, N5320, N4497);
and AND2 (N5326, N5324, N4902);
nand NAND2 (N5327, N5321, N4182);
and AND2 (N5328, N5311, N1376);
or OR3 (N5329, N5323, N5003, N1954);
or OR4 (N5330, N5325, N3878, N3739, N1893);
xor XOR2 (N5331, N5299, N5161);
nor NOR2 (N5332, N5304, N5268);
xor XOR2 (N5333, N5331, N1329);
or OR2 (N5334, N5328, N3725);
or OR2 (N5335, N5330, N3975);
buf BUF1 (N5336, N5303);
not NOT1 (N5337, N5329);
nand NAND3 (N5338, N5333, N3673, N2317);
or OR4 (N5339, N5336, N3567, N3759, N1797);
or OR4 (N5340, N5338, N2561, N3983, N4887);
buf BUF1 (N5341, N5340);
or OR3 (N5342, N5332, N793, N2013);
xor XOR2 (N5343, N5342, N818);
xor XOR2 (N5344, N5271, N4219);
nor NOR3 (N5345, N5335, N2347, N4440);
not NOT1 (N5346, N5341);
nand NAND3 (N5347, N5339, N1839, N1651);
nand NAND3 (N5348, N5334, N730, N2554);
or OR4 (N5349, N5319, N1396, N3891, N3602);
xor XOR2 (N5350, N5344, N2444);
nand NAND3 (N5351, N5343, N637, N3346);
nor NOR2 (N5352, N5348, N4155);
buf BUF1 (N5353, N5350);
and AND3 (N5354, N5345, N4746, N2608);
and AND4 (N5355, N5347, N3294, N5190, N3009);
buf BUF1 (N5356, N5327);
nand NAND3 (N5357, N5349, N5154, N221);
not NOT1 (N5358, N5352);
or OR4 (N5359, N5355, N3448, N4148, N3984);
nor NOR4 (N5360, N5337, N4709, N2763, N1114);
and AND2 (N5361, N5356, N4757);
and AND2 (N5362, N5360, N1125);
not NOT1 (N5363, N5361);
nor NOR3 (N5364, N5358, N3500, N1180);
or OR3 (N5365, N5357, N4525, N1589);
xor XOR2 (N5366, N5353, N1051);
buf BUF1 (N5367, N5346);
not NOT1 (N5368, N5359);
nor NOR2 (N5369, N5326, N4526);
or OR2 (N5370, N5368, N1443);
xor XOR2 (N5371, N5362, N648);
or OR3 (N5372, N5369, N3308, N2698);
nor NOR3 (N5373, N5367, N1418, N1947);
xor XOR2 (N5374, N5354, N1685);
not NOT1 (N5375, N5373);
buf BUF1 (N5376, N5351);
or OR2 (N5377, N5376, N2311);
or OR3 (N5378, N5377, N3122, N3349);
nand NAND3 (N5379, N5371, N3850, N2716);
xor XOR2 (N5380, N5372, N2805);
nand NAND3 (N5381, N5380, N1630, N4786);
and AND3 (N5382, N5370, N2594, N3396);
and AND2 (N5383, N5378, N280);
xor XOR2 (N5384, N5382, N179);
not NOT1 (N5385, N5374);
nor NOR2 (N5386, N5365, N3363);
not NOT1 (N5387, N5364);
nor NOR2 (N5388, N5383, N4153);
nor NOR3 (N5389, N5387, N691, N2500);
or OR3 (N5390, N5386, N4511, N3580);
xor XOR2 (N5391, N5388, N2823);
nor NOR2 (N5392, N5389, N1560);
nand NAND3 (N5393, N5385, N5229, N2686);
nand NAND3 (N5394, N5379, N1817, N224);
nand NAND3 (N5395, N5394, N4249, N1632);
buf BUF1 (N5396, N5390);
or OR4 (N5397, N5391, N3803, N1355, N4434);
or OR4 (N5398, N5396, N507, N2688, N3001);
or OR2 (N5399, N5366, N3371);
xor XOR2 (N5400, N5399, N2321);
nor NOR4 (N5401, N5392, N965, N4416, N431);
not NOT1 (N5402, N5384);
nor NOR3 (N5403, N5393, N4070, N4342);
buf BUF1 (N5404, N5375);
buf BUF1 (N5405, N5402);
and AND4 (N5406, N5400, N4594, N3547, N1834);
buf BUF1 (N5407, N5363);
nor NOR3 (N5408, N5398, N2689, N2730);
not NOT1 (N5409, N5381);
and AND3 (N5410, N5405, N5106, N2617);
or OR2 (N5411, N5401, N4650);
nand NAND4 (N5412, N5407, N5281, N2054, N1484);
buf BUF1 (N5413, N5404);
buf BUF1 (N5414, N5395);
nand NAND4 (N5415, N5413, N683, N1863, N3369);
nor NOR2 (N5416, N5412, N4018);
and AND3 (N5417, N5409, N3060, N5329);
or OR4 (N5418, N5397, N3325, N4330, N5014);
xor XOR2 (N5419, N5408, N79);
or OR3 (N5420, N5417, N4409, N3501);
buf BUF1 (N5421, N5418);
and AND2 (N5422, N5421, N598);
nand NAND2 (N5423, N5415, N3486);
nand NAND4 (N5424, N5423, N596, N2024, N786);
or OR2 (N5425, N5403, N4906);
xor XOR2 (N5426, N5425, N4937);
or OR2 (N5427, N5411, N5192);
nand NAND4 (N5428, N5420, N158, N4008, N4059);
and AND4 (N5429, N5410, N2070, N2977, N4935);
buf BUF1 (N5430, N5424);
not NOT1 (N5431, N5427);
nand NAND3 (N5432, N5422, N4525, N4537);
not NOT1 (N5433, N5430);
buf BUF1 (N5434, N5429);
nor NOR4 (N5435, N5416, N1051, N2935, N4613);
or OR2 (N5436, N5414, N4599);
not NOT1 (N5437, N5431);
nand NAND3 (N5438, N5419, N2263, N1520);
and AND2 (N5439, N5426, N255);
xor XOR2 (N5440, N5434, N3472);
and AND2 (N5441, N5432, N3667);
and AND3 (N5442, N5406, N390, N4158);
nor NOR3 (N5443, N5435, N1112, N1623);
xor XOR2 (N5444, N5433, N2620);
nand NAND2 (N5445, N5442, N1283);
nand NAND4 (N5446, N5438, N147, N1832, N947);
not NOT1 (N5447, N5441);
nor NOR2 (N5448, N5428, N4841);
xor XOR2 (N5449, N5437, N1805);
not NOT1 (N5450, N5446);
xor XOR2 (N5451, N5445, N5362);
not NOT1 (N5452, N5450);
nand NAND2 (N5453, N5443, N3934);
buf BUF1 (N5454, N5453);
or OR4 (N5455, N5436, N5092, N5013, N4689);
buf BUF1 (N5456, N5454);
and AND4 (N5457, N5444, N4566, N3808, N4093);
or OR3 (N5458, N5439, N736, N966);
buf BUF1 (N5459, N5449);
or OR3 (N5460, N5447, N2922, N1298);
not NOT1 (N5461, N5458);
xor XOR2 (N5462, N5455, N125);
xor XOR2 (N5463, N5462, N2748);
nand NAND4 (N5464, N5461, N3099, N3266, N5391);
not NOT1 (N5465, N5459);
and AND3 (N5466, N5456, N1076, N345);
and AND2 (N5467, N5451, N1117);
and AND4 (N5468, N5467, N1895, N629, N2020);
not NOT1 (N5469, N5466);
or OR4 (N5470, N5457, N4036, N89, N4597);
not NOT1 (N5471, N5465);
buf BUF1 (N5472, N5448);
or OR2 (N5473, N5471, N331);
buf BUF1 (N5474, N5440);
nor NOR3 (N5475, N5473, N3588, N4764);
or OR2 (N5476, N5475, N2846);
not NOT1 (N5477, N5460);
or OR3 (N5478, N5472, N2331, N357);
buf BUF1 (N5479, N5470);
xor XOR2 (N5480, N5464, N5279);
xor XOR2 (N5481, N5479, N4393);
and AND2 (N5482, N5452, N4859);
or OR2 (N5483, N5468, N3338);
and AND2 (N5484, N5482, N5121);
not NOT1 (N5485, N5484);
nor NOR3 (N5486, N5485, N2036, N3084);
nor NOR2 (N5487, N5476, N3693);
or OR2 (N5488, N5481, N4286);
or OR4 (N5489, N5463, N1544, N5075, N1553);
or OR2 (N5490, N5487, N3026);
and AND3 (N5491, N5480, N84, N4869);
or OR3 (N5492, N5491, N2372, N419);
xor XOR2 (N5493, N5488, N3886);
buf BUF1 (N5494, N5478);
or OR4 (N5495, N5494, N396, N342, N393);
or OR3 (N5496, N5489, N5022, N3911);
xor XOR2 (N5497, N5486, N2918);
nor NOR4 (N5498, N5490, N4501, N1176, N5158);
nand NAND4 (N5499, N5498, N3143, N946, N755);
and AND4 (N5500, N5477, N4073, N464, N1727);
nor NOR3 (N5501, N5469, N3789, N4084);
nand NAND4 (N5502, N5497, N3181, N66, N1321);
not NOT1 (N5503, N5474);
buf BUF1 (N5504, N5503);
nand NAND2 (N5505, N5492, N4897);
not NOT1 (N5506, N5499);
xor XOR2 (N5507, N5483, N233);
nor NOR2 (N5508, N5495, N4323);
and AND3 (N5509, N5501, N4081, N1124);
or OR2 (N5510, N5506, N1036);
nor NOR2 (N5511, N5496, N1998);
nor NOR2 (N5512, N5507, N2740);
not NOT1 (N5513, N5508);
or OR2 (N5514, N5504, N4910);
and AND3 (N5515, N5514, N4755, N1250);
not NOT1 (N5516, N5500);
xor XOR2 (N5517, N5502, N2318);
or OR4 (N5518, N5512, N2124, N2070, N5301);
buf BUF1 (N5519, N5505);
nand NAND2 (N5520, N5509, N4841);
buf BUF1 (N5521, N5519);
buf BUF1 (N5522, N5521);
not NOT1 (N5523, N5511);
not NOT1 (N5524, N5523);
not NOT1 (N5525, N5524);
or OR3 (N5526, N5513, N2023, N3228);
not NOT1 (N5527, N5516);
xor XOR2 (N5528, N5517, N743);
and AND3 (N5529, N5518, N4121, N4589);
or OR3 (N5530, N5520, N2097, N1331);
not NOT1 (N5531, N5522);
nor NOR3 (N5532, N5529, N3846, N2606);
nor NOR3 (N5533, N5530, N3262, N565);
nand NAND3 (N5534, N5515, N2709, N4845);
nand NAND3 (N5535, N5527, N4133, N1756);
nor NOR3 (N5536, N5531, N1472, N873);
xor XOR2 (N5537, N5526, N2644);
and AND3 (N5538, N5528, N623, N4622);
and AND4 (N5539, N5537, N1924, N186, N1212);
nor NOR2 (N5540, N5510, N1163);
not NOT1 (N5541, N5493);
xor XOR2 (N5542, N5541, N5123);
nand NAND4 (N5543, N5535, N2952, N3176, N2420);
nor NOR4 (N5544, N5542, N826, N2529, N2171);
xor XOR2 (N5545, N5534, N115);
nor NOR3 (N5546, N5538, N2210, N3661);
nand NAND3 (N5547, N5546, N1105, N3756);
buf BUF1 (N5548, N5536);
nor NOR2 (N5549, N5544, N4136);
nand NAND4 (N5550, N5532, N320, N3252, N2580);
nand NAND2 (N5551, N5525, N483);
not NOT1 (N5552, N5550);
nand NAND4 (N5553, N5540, N100, N5447, N3195);
or OR4 (N5554, N5551, N3149, N4406, N2495);
or OR4 (N5555, N5543, N557, N1919, N4196);
nand NAND4 (N5556, N5553, N1794, N5194, N98);
and AND3 (N5557, N5533, N4858, N3323);
nor NOR4 (N5558, N5547, N355, N5314, N3285);
xor XOR2 (N5559, N5545, N4488);
not NOT1 (N5560, N5549);
nand NAND2 (N5561, N5558, N1663);
xor XOR2 (N5562, N5556, N3854);
nand NAND4 (N5563, N5561, N5200, N615, N3676);
and AND3 (N5564, N5539, N1259, N3423);
or OR2 (N5565, N5555, N5332);
buf BUF1 (N5566, N5562);
not NOT1 (N5567, N5557);
not NOT1 (N5568, N5566);
not NOT1 (N5569, N5552);
nand NAND4 (N5570, N5563, N4748, N2540, N938);
nor NOR3 (N5571, N5559, N217, N3961);
xor XOR2 (N5572, N5548, N3001);
xor XOR2 (N5573, N5564, N3542);
nor NOR3 (N5574, N5573, N1256, N882);
and AND2 (N5575, N5574, N2282);
xor XOR2 (N5576, N5568, N53);
not NOT1 (N5577, N5560);
not NOT1 (N5578, N5575);
and AND2 (N5579, N5577, N4204);
xor XOR2 (N5580, N5554, N3417);
nor NOR3 (N5581, N5567, N2170, N4712);
nor NOR4 (N5582, N5581, N3914, N4024, N2950);
or OR4 (N5583, N5582, N872, N1446, N1655);
buf BUF1 (N5584, N5580);
buf BUF1 (N5585, N5584);
buf BUF1 (N5586, N5571);
nor NOR3 (N5587, N5565, N3585, N3725);
nor NOR4 (N5588, N5586, N2055, N4529, N2691);
not NOT1 (N5589, N5576);
or OR3 (N5590, N5569, N3984, N4683);
and AND3 (N5591, N5587, N4917, N4745);
nor NOR4 (N5592, N5590, N158, N3274, N2482);
xor XOR2 (N5593, N5579, N2167);
xor XOR2 (N5594, N5570, N5107);
or OR2 (N5595, N5593, N1788);
xor XOR2 (N5596, N5591, N1889);
nor NOR4 (N5597, N5595, N797, N4615, N785);
or OR4 (N5598, N5594, N4208, N1510, N4069);
buf BUF1 (N5599, N5592);
nor NOR2 (N5600, N5578, N767);
and AND4 (N5601, N5589, N1610, N3554, N4384);
not NOT1 (N5602, N5599);
not NOT1 (N5603, N5597);
and AND4 (N5604, N5602, N250, N3677, N2288);
or OR4 (N5605, N5600, N3709, N3368, N4033);
xor XOR2 (N5606, N5585, N1603);
nand NAND3 (N5607, N5603, N220, N4222);
buf BUF1 (N5608, N5596);
or OR3 (N5609, N5583, N385, N231);
or OR4 (N5610, N5605, N4691, N2158, N4147);
or OR2 (N5611, N5604, N2373);
buf BUF1 (N5612, N5607);
nor NOR4 (N5613, N5612, N4567, N3767, N3432);
and AND3 (N5614, N5610, N2871, N4611);
or OR2 (N5615, N5613, N343);
nand NAND2 (N5616, N5608, N4251);
nand NAND4 (N5617, N5616, N3286, N3909, N5412);
nor NOR3 (N5618, N5588, N2597, N1782);
buf BUF1 (N5619, N5598);
and AND2 (N5620, N5611, N287);
nand NAND2 (N5621, N5601, N2937);
and AND4 (N5622, N5617, N2866, N4179, N2517);
or OR4 (N5623, N5622, N2036, N4281, N3568);
not NOT1 (N5624, N5619);
and AND4 (N5625, N5623, N3940, N2444, N1275);
and AND4 (N5626, N5625, N4843, N1638, N3030);
nand NAND4 (N5627, N5621, N2330, N4269, N573);
nand NAND2 (N5628, N5615, N1711);
nor NOR4 (N5629, N5572, N724, N3348, N5479);
not NOT1 (N5630, N5614);
xor XOR2 (N5631, N5624, N5535);
not NOT1 (N5632, N5631);
buf BUF1 (N5633, N5627);
and AND4 (N5634, N5633, N5321, N1102, N1912);
not NOT1 (N5635, N5618);
not NOT1 (N5636, N5629);
nand NAND3 (N5637, N5635, N1103, N367);
xor XOR2 (N5638, N5632, N2220);
and AND4 (N5639, N5630, N1339, N3055, N2117);
buf BUF1 (N5640, N5626);
buf BUF1 (N5641, N5634);
not NOT1 (N5642, N5609);
buf BUF1 (N5643, N5639);
buf BUF1 (N5644, N5641);
xor XOR2 (N5645, N5642, N544);
or OR2 (N5646, N5636, N4019);
nand NAND2 (N5647, N5637, N2623);
xor XOR2 (N5648, N5606, N4364);
buf BUF1 (N5649, N5646);
and AND2 (N5650, N5638, N5501);
nor NOR2 (N5651, N5645, N1332);
buf BUF1 (N5652, N5649);
nor NOR3 (N5653, N5644, N784, N503);
buf BUF1 (N5654, N5653);
nand NAND3 (N5655, N5647, N3941, N2376);
or OR2 (N5656, N5651, N2216);
nand NAND2 (N5657, N5650, N1877);
xor XOR2 (N5658, N5643, N4404);
xor XOR2 (N5659, N5654, N397);
nand NAND3 (N5660, N5640, N58, N923);
buf BUF1 (N5661, N5655);
and AND3 (N5662, N5659, N3746, N5521);
xor XOR2 (N5663, N5661, N3146);
nand NAND4 (N5664, N5662, N2648, N5534, N1913);
nor NOR2 (N5665, N5620, N3931);
not NOT1 (N5666, N5660);
nand NAND4 (N5667, N5648, N5455, N5165, N5386);
or OR3 (N5668, N5657, N1622, N4847);
not NOT1 (N5669, N5668);
nand NAND3 (N5670, N5658, N560, N129);
nor NOR3 (N5671, N5670, N342, N2097);
or OR2 (N5672, N5666, N5169);
xor XOR2 (N5673, N5628, N36);
not NOT1 (N5674, N5652);
nand NAND2 (N5675, N5673, N2185);
buf BUF1 (N5676, N5675);
xor XOR2 (N5677, N5665, N2053);
xor XOR2 (N5678, N5672, N1508);
buf BUF1 (N5679, N5663);
nand NAND3 (N5680, N5656, N2530, N4374);
not NOT1 (N5681, N5679);
buf BUF1 (N5682, N5680);
and AND4 (N5683, N5682, N4780, N5546, N3239);
or OR4 (N5684, N5664, N2820, N1811, N244);
or OR3 (N5685, N5676, N4221, N3814);
not NOT1 (N5686, N5674);
or OR3 (N5687, N5686, N1798, N3476);
buf BUF1 (N5688, N5683);
nor NOR2 (N5689, N5684, N5570);
nand NAND4 (N5690, N5677, N2884, N2652, N3328);
and AND4 (N5691, N5685, N80, N1828, N44);
buf BUF1 (N5692, N5678);
or OR4 (N5693, N5681, N2479, N4423, N5166);
nand NAND4 (N5694, N5691, N4389, N5008, N1842);
buf BUF1 (N5695, N5690);
nor NOR3 (N5696, N5667, N4050, N1539);
nor NOR3 (N5697, N5696, N966, N1372);
xor XOR2 (N5698, N5671, N5005);
nor NOR3 (N5699, N5695, N1642, N3758);
buf BUF1 (N5700, N5669);
or OR3 (N5701, N5694, N1645, N1409);
nand NAND4 (N5702, N5689, N1115, N3941, N1403);
xor XOR2 (N5703, N5702, N1663);
nor NOR2 (N5704, N5703, N4064);
or OR2 (N5705, N5701, N4369);
or OR2 (N5706, N5688, N2387);
nand NAND3 (N5707, N5687, N5394, N3897);
nor NOR4 (N5708, N5705, N4834, N744, N409);
or OR2 (N5709, N5697, N4434);
not NOT1 (N5710, N5708);
nand NAND3 (N5711, N5707, N5353, N5274);
xor XOR2 (N5712, N5700, N4709);
buf BUF1 (N5713, N5699);
and AND2 (N5714, N5693, N3095);
or OR4 (N5715, N5706, N863, N4855, N3100);
xor XOR2 (N5716, N5713, N3283);
buf BUF1 (N5717, N5698);
not NOT1 (N5718, N5704);
xor XOR2 (N5719, N5709, N5017);
and AND4 (N5720, N5711, N5364, N2882, N4412);
buf BUF1 (N5721, N5719);
or OR2 (N5722, N5720, N1021);
nor NOR3 (N5723, N5718, N5269, N2932);
xor XOR2 (N5724, N5714, N2685);
or OR4 (N5725, N5692, N2002, N4136, N1994);
or OR3 (N5726, N5717, N5217, N2121);
xor XOR2 (N5727, N5715, N1279);
nor NOR2 (N5728, N5725, N3104);
nor NOR4 (N5729, N5728, N2141, N2416, N4145);
not NOT1 (N5730, N5724);
nand NAND2 (N5731, N5723, N1822);
not NOT1 (N5732, N5722);
nor NOR4 (N5733, N5731, N3223, N122, N1975);
buf BUF1 (N5734, N5726);
and AND4 (N5735, N5716, N733, N4583, N1400);
nor NOR4 (N5736, N5727, N3208, N4054, N3131);
nor NOR3 (N5737, N5730, N3503, N3911);
xor XOR2 (N5738, N5729, N1309);
and AND2 (N5739, N5721, N3649);
xor XOR2 (N5740, N5734, N2459);
nand NAND3 (N5741, N5740, N1043, N807);
buf BUF1 (N5742, N5735);
buf BUF1 (N5743, N5737);
not NOT1 (N5744, N5743);
or OR3 (N5745, N5738, N993, N2372);
and AND3 (N5746, N5732, N5368, N781);
xor XOR2 (N5747, N5733, N1888);
nand NAND3 (N5748, N5746, N1458, N3177);
not NOT1 (N5749, N5739);
not NOT1 (N5750, N5712);
or OR4 (N5751, N5750, N3766, N4388, N4399);
buf BUF1 (N5752, N5744);
not NOT1 (N5753, N5752);
nand NAND4 (N5754, N5753, N3678, N5040, N3856);
nor NOR4 (N5755, N5736, N1942, N5388, N56);
nor NOR3 (N5756, N5742, N889, N5121);
and AND2 (N5757, N5751, N614);
not NOT1 (N5758, N5745);
xor XOR2 (N5759, N5748, N92);
and AND2 (N5760, N5755, N239);
nand NAND4 (N5761, N5710, N2633, N3638, N412);
or OR2 (N5762, N5741, N2367);
or OR3 (N5763, N5759, N999, N5669);
nand NAND4 (N5764, N5757, N929, N257, N1622);
and AND4 (N5765, N5747, N4808, N3561, N3003);
xor XOR2 (N5766, N5763, N3920);
xor XOR2 (N5767, N5756, N2418);
or OR4 (N5768, N5762, N1578, N5534, N3818);
nor NOR2 (N5769, N5767, N2471);
nand NAND2 (N5770, N5764, N4117);
xor XOR2 (N5771, N5749, N1653);
not NOT1 (N5772, N5761);
and AND2 (N5773, N5758, N5058);
buf BUF1 (N5774, N5760);
and AND4 (N5775, N5754, N1621, N1932, N842);
nor NOR4 (N5776, N5772, N3715, N3514, N3068);
nor NOR4 (N5777, N5776, N4424, N1909, N4214);
xor XOR2 (N5778, N5771, N4439);
not NOT1 (N5779, N5777);
or OR3 (N5780, N5778, N3779, N2403);
nand NAND4 (N5781, N5768, N3844, N4506, N2821);
nor NOR3 (N5782, N5769, N4131, N4581);
buf BUF1 (N5783, N5782);
not NOT1 (N5784, N5781);
nand NAND3 (N5785, N5783, N4991, N5323);
and AND3 (N5786, N5773, N2704, N5460);
not NOT1 (N5787, N5770);
xor XOR2 (N5788, N5780, N4716);
nand NAND3 (N5789, N5779, N4572, N5365);
or OR4 (N5790, N5775, N2487, N1844, N487);
not NOT1 (N5791, N5790);
xor XOR2 (N5792, N5765, N5027);
buf BUF1 (N5793, N5785);
nor NOR4 (N5794, N5789, N1663, N1517, N3089);
xor XOR2 (N5795, N5786, N3920);
and AND3 (N5796, N5791, N5666, N2154);
not NOT1 (N5797, N5795);
nor NOR3 (N5798, N5788, N2059, N5585);
buf BUF1 (N5799, N5784);
not NOT1 (N5800, N5796);
nor NOR2 (N5801, N5774, N731);
nand NAND3 (N5802, N5793, N823, N3094);
buf BUF1 (N5803, N5794);
buf BUF1 (N5804, N5799);
and AND2 (N5805, N5800, N1127);
buf BUF1 (N5806, N5792);
and AND3 (N5807, N5805, N3452, N327);
xor XOR2 (N5808, N5807, N485);
buf BUF1 (N5809, N5801);
and AND3 (N5810, N5798, N5585, N1157);
and AND4 (N5811, N5766, N4717, N294, N5205);
not NOT1 (N5812, N5804);
nand NAND2 (N5813, N5803, N1526);
and AND2 (N5814, N5811, N81);
not NOT1 (N5815, N5808);
buf BUF1 (N5816, N5802);
buf BUF1 (N5817, N5787);
buf BUF1 (N5818, N5817);
or OR4 (N5819, N5816, N966, N2226, N1436);
not NOT1 (N5820, N5797);
not NOT1 (N5821, N5813);
buf BUF1 (N5822, N5812);
buf BUF1 (N5823, N5806);
and AND3 (N5824, N5810, N2962, N4518);
nand NAND4 (N5825, N5818, N2290, N1187, N1956);
not NOT1 (N5826, N5819);
xor XOR2 (N5827, N5815, N2969);
nor NOR4 (N5828, N5823, N1086, N2197, N14);
and AND3 (N5829, N5827, N3636, N2064);
or OR2 (N5830, N5826, N4431);
nand NAND3 (N5831, N5828, N311, N2491);
nor NOR2 (N5832, N5831, N5045);
and AND2 (N5833, N5825, N2310);
buf BUF1 (N5834, N5821);
nor NOR4 (N5835, N5809, N4059, N705, N3672);
and AND3 (N5836, N5814, N4858, N746);
nor NOR4 (N5837, N5822, N2190, N753, N4864);
not NOT1 (N5838, N5829);
nor NOR3 (N5839, N5835, N4047, N4660);
or OR2 (N5840, N5838, N4773);
nor NOR2 (N5841, N5839, N793);
xor XOR2 (N5842, N5836, N5578);
not NOT1 (N5843, N5833);
xor XOR2 (N5844, N5843, N11);
nand NAND2 (N5845, N5840, N4291);
not NOT1 (N5846, N5842);
not NOT1 (N5847, N5830);
buf BUF1 (N5848, N5841);
and AND4 (N5849, N5847, N4654, N2620, N1352);
or OR4 (N5850, N5834, N234, N3796, N647);
nand NAND2 (N5851, N5824, N5165);
nand NAND4 (N5852, N5845, N2304, N4517, N3069);
or OR3 (N5853, N5849, N723, N3344);
xor XOR2 (N5854, N5848, N4637);
not NOT1 (N5855, N5850);
or OR2 (N5856, N5846, N1295);
and AND3 (N5857, N5855, N3711, N2127);
xor XOR2 (N5858, N5854, N1429);
buf BUF1 (N5859, N5844);
and AND2 (N5860, N5859, N3052);
xor XOR2 (N5861, N5858, N546);
and AND4 (N5862, N5837, N3789, N516, N5516);
or OR2 (N5863, N5861, N4755);
or OR4 (N5864, N5851, N2969, N3840, N3165);
or OR3 (N5865, N5862, N1769, N3224);
nand NAND3 (N5866, N5865, N718, N457);
buf BUF1 (N5867, N5820);
xor XOR2 (N5868, N5864, N2848);
xor XOR2 (N5869, N5868, N4268);
nor NOR4 (N5870, N5863, N2527, N3455, N3113);
not NOT1 (N5871, N5866);
and AND2 (N5872, N5871, N2822);
nand NAND3 (N5873, N5852, N1459, N2196);
or OR4 (N5874, N5873, N3992, N3401, N5581);
or OR4 (N5875, N5856, N1910, N1633, N3154);
xor XOR2 (N5876, N5869, N5074);
and AND4 (N5877, N5853, N4757, N1067, N4498);
nand NAND4 (N5878, N5867, N4320, N1137, N1395);
not NOT1 (N5879, N5870);
nand NAND4 (N5880, N5860, N3121, N1751, N537);
or OR2 (N5881, N5832, N1558);
and AND2 (N5882, N5881, N3371);
or OR2 (N5883, N5874, N2007);
xor XOR2 (N5884, N5857, N2233);
xor XOR2 (N5885, N5880, N2413);
or OR3 (N5886, N5876, N1359, N801);
not NOT1 (N5887, N5877);
not NOT1 (N5888, N5886);
buf BUF1 (N5889, N5875);
buf BUF1 (N5890, N5883);
xor XOR2 (N5891, N5890, N2711);
nand NAND4 (N5892, N5885, N1546, N734, N3045);
buf BUF1 (N5893, N5888);
nor NOR4 (N5894, N5887, N3195, N2443, N2870);
or OR2 (N5895, N5889, N1996);
and AND4 (N5896, N5893, N1905, N3670, N214);
or OR4 (N5897, N5895, N212, N3468, N4169);
nor NOR2 (N5898, N5884, N4669);
nand NAND3 (N5899, N5892, N3546, N1381);
nor NOR4 (N5900, N5879, N3156, N1795, N1780);
xor XOR2 (N5901, N5891, N5462);
buf BUF1 (N5902, N5901);
buf BUF1 (N5903, N5878);
xor XOR2 (N5904, N5894, N4159);
xor XOR2 (N5905, N5882, N2312);
xor XOR2 (N5906, N5897, N5719);
and AND4 (N5907, N5904, N3713, N2213, N3357);
nor NOR4 (N5908, N5898, N1307, N4829, N5235);
nor NOR2 (N5909, N5896, N2016);
nor NOR3 (N5910, N5900, N5384, N3883);
nor NOR2 (N5911, N5910, N2023);
and AND2 (N5912, N5905, N620);
buf BUF1 (N5913, N5872);
and AND3 (N5914, N5902, N836, N4947);
buf BUF1 (N5915, N5912);
or OR3 (N5916, N5908, N3037, N4032);
xor XOR2 (N5917, N5914, N3492);
and AND2 (N5918, N5899, N5621);
buf BUF1 (N5919, N5917);
or OR3 (N5920, N5903, N4428, N1511);
buf BUF1 (N5921, N5919);
nand NAND3 (N5922, N5907, N5323, N2190);
and AND3 (N5923, N5915, N99, N3591);
buf BUF1 (N5924, N5913);
xor XOR2 (N5925, N5909, N5668);
nor NOR2 (N5926, N5924, N4170);
nor NOR3 (N5927, N5916, N5299, N5032);
xor XOR2 (N5928, N5921, N136);
or OR2 (N5929, N5927, N4838);
or OR2 (N5930, N5911, N4766);
not NOT1 (N5931, N5918);
or OR3 (N5932, N5923, N3669, N1004);
xor XOR2 (N5933, N5922, N5166);
not NOT1 (N5934, N5925);
or OR3 (N5935, N5928, N4098, N2803);
nor NOR3 (N5936, N5906, N442, N891);
nand NAND3 (N5937, N5936, N1392, N1344);
and AND2 (N5938, N5935, N1275);
not NOT1 (N5939, N5931);
xor XOR2 (N5940, N5929, N626);
nand NAND2 (N5941, N5932, N1381);
or OR2 (N5942, N5941, N3411);
xor XOR2 (N5943, N5933, N553);
not NOT1 (N5944, N5938);
or OR3 (N5945, N5920, N3679, N3949);
buf BUF1 (N5946, N5945);
xor XOR2 (N5947, N5940, N4702);
xor XOR2 (N5948, N5937, N3639);
buf BUF1 (N5949, N5943);
and AND3 (N5950, N5947, N4144, N4783);
xor XOR2 (N5951, N5939, N4571);
and AND4 (N5952, N5949, N1160, N1943, N1233);
nor NOR3 (N5953, N5948, N4863, N5494);
and AND3 (N5954, N5942, N4085, N1321);
not NOT1 (N5955, N5946);
buf BUF1 (N5956, N5954);
nor NOR2 (N5957, N5952, N4839);
and AND4 (N5958, N5951, N1144, N2448, N2913);
or OR2 (N5959, N5930, N2002);
not NOT1 (N5960, N5934);
or OR4 (N5961, N5950, N4239, N4047, N5289);
or OR4 (N5962, N5961, N4427, N4231, N1640);
and AND2 (N5963, N5960, N2615);
nand NAND2 (N5964, N5926, N376);
buf BUF1 (N5965, N5964);
xor XOR2 (N5966, N5953, N1960);
nand NAND3 (N5967, N5955, N1142, N5707);
buf BUF1 (N5968, N5957);
and AND3 (N5969, N5963, N1682, N2846);
not NOT1 (N5970, N5968);
nor NOR3 (N5971, N5962, N1900, N4856);
or OR4 (N5972, N5959, N2131, N1519, N3459);
xor XOR2 (N5973, N5958, N5391);
and AND4 (N5974, N5973, N70, N4899, N1216);
nand NAND2 (N5975, N5967, N3414);
buf BUF1 (N5976, N5972);
or OR3 (N5977, N5974, N1758, N97);
and AND3 (N5978, N5944, N2717, N5742);
xor XOR2 (N5979, N5978, N5457);
or OR2 (N5980, N5965, N1672);
buf BUF1 (N5981, N5956);
and AND4 (N5982, N5975, N3380, N2130, N3992);
nor NOR4 (N5983, N5970, N1314, N989, N2198);
not NOT1 (N5984, N5979);
buf BUF1 (N5985, N5969);
nor NOR2 (N5986, N5984, N1887);
nand NAND2 (N5987, N5971, N2276);
and AND3 (N5988, N5976, N551, N3493);
not NOT1 (N5989, N5986);
and AND2 (N5990, N5988, N4446);
or OR3 (N5991, N5982, N5630, N4978);
xor XOR2 (N5992, N5977, N1010);
xor XOR2 (N5993, N5981, N4067);
and AND2 (N5994, N5991, N3389);
xor XOR2 (N5995, N5992, N2240);
not NOT1 (N5996, N5985);
not NOT1 (N5997, N5993);
not NOT1 (N5998, N5994);
and AND2 (N5999, N5980, N4916);
buf BUF1 (N6000, N5990);
nor NOR3 (N6001, N5989, N2796, N5397);
nand NAND4 (N6002, N6000, N2125, N2897, N5398);
xor XOR2 (N6003, N5996, N613);
buf BUF1 (N6004, N5999);
not NOT1 (N6005, N6003);
buf BUF1 (N6006, N6005);
nand NAND2 (N6007, N6006, N2683);
or OR4 (N6008, N5997, N1657, N1170, N130);
buf BUF1 (N6009, N5966);
buf BUF1 (N6010, N6001);
or OR4 (N6011, N6007, N2463, N5453, N1645);
xor XOR2 (N6012, N6008, N4981);
and AND3 (N6013, N5987, N2068, N3477);
and AND3 (N6014, N5983, N2928, N4390);
nor NOR2 (N6015, N6004, N3266);
buf BUF1 (N6016, N6013);
nor NOR4 (N6017, N5995, N1714, N5753, N4004);
xor XOR2 (N6018, N6011, N333);
not NOT1 (N6019, N6014);
buf BUF1 (N6020, N6009);
not NOT1 (N6021, N6016);
or OR3 (N6022, N6017, N3774, N3579);
nor NOR3 (N6023, N6019, N5744, N3787);
nand NAND3 (N6024, N6002, N3181, N2462);
and AND3 (N6025, N6023, N3486, N533);
or OR3 (N6026, N6025, N1789, N3646);
or OR2 (N6027, N6015, N910);
nand NAND4 (N6028, N5998, N1627, N5764, N6017);
not NOT1 (N6029, N6026);
nand NAND4 (N6030, N6029, N2055, N246, N2354);
nand NAND2 (N6031, N6022, N3853);
xor XOR2 (N6032, N6028, N4579);
nand NAND2 (N6033, N6030, N474);
or OR4 (N6034, N6021, N3299, N1092, N3070);
xor XOR2 (N6035, N6012, N2576);
nand NAND4 (N6036, N6018, N2581, N2275, N4179);
and AND4 (N6037, N6010, N5840, N4435, N4433);
or OR3 (N6038, N6024, N2499, N162);
nand NAND4 (N6039, N6034, N2641, N3064, N5696);
not NOT1 (N6040, N6039);
nor NOR3 (N6041, N6033, N2822, N2772);
xor XOR2 (N6042, N6032, N5974);
not NOT1 (N6043, N6038);
buf BUF1 (N6044, N6027);
buf BUF1 (N6045, N6035);
nand NAND3 (N6046, N6040, N3750, N2742);
buf BUF1 (N6047, N6031);
nor NOR4 (N6048, N6036, N4630, N4200, N498);
or OR2 (N6049, N6043, N2732);
nand NAND2 (N6050, N6049, N2976);
xor XOR2 (N6051, N6047, N1977);
nand NAND2 (N6052, N6050, N4632);
buf BUF1 (N6053, N6052);
buf BUF1 (N6054, N6046);
or OR3 (N6055, N6045, N3058, N5266);
nor NOR3 (N6056, N6054, N3091, N4337);
nand NAND4 (N6057, N6041, N962, N4326, N464);
or OR4 (N6058, N6044, N4091, N1531, N1776);
not NOT1 (N6059, N6057);
xor XOR2 (N6060, N6020, N2544);
and AND4 (N6061, N6048, N395, N1948, N723);
and AND3 (N6062, N6037, N270, N3629);
or OR4 (N6063, N6053, N3863, N5511, N5501);
not NOT1 (N6064, N6051);
nand NAND3 (N6065, N6060, N3841, N2775);
nor NOR3 (N6066, N6062, N1516, N1335);
nand NAND3 (N6067, N6042, N4416, N2312);
nor NOR4 (N6068, N6066, N246, N4349, N2192);
or OR2 (N6069, N6061, N5185);
and AND3 (N6070, N6058, N1663, N5326);
buf BUF1 (N6071, N6055);
nand NAND2 (N6072, N6069, N4159);
or OR2 (N6073, N6070, N194);
xor XOR2 (N6074, N6071, N583);
and AND3 (N6075, N6059, N2958, N3270);
nand NAND4 (N6076, N6063, N1028, N205, N4422);
buf BUF1 (N6077, N6064);
buf BUF1 (N6078, N6074);
nor NOR2 (N6079, N6072, N3580);
nor NOR4 (N6080, N6077, N5251, N1392, N1101);
or OR4 (N6081, N6079, N4661, N5807, N3320);
nand NAND3 (N6082, N6076, N4755, N604);
xor XOR2 (N6083, N6080, N2020);
xor XOR2 (N6084, N6068, N5970);
and AND3 (N6085, N6082, N5244, N5008);
nor NOR4 (N6086, N6085, N316, N3544, N3462);
not NOT1 (N6087, N6078);
buf BUF1 (N6088, N6056);
nand NAND3 (N6089, N6088, N3340, N2282);
and AND2 (N6090, N6067, N2714);
nor NOR3 (N6091, N6086, N5293, N1560);
nand NAND4 (N6092, N6090, N2474, N1921, N615);
or OR3 (N6093, N6087, N1762, N5135);
or OR3 (N6094, N6093, N3691, N114);
nor NOR4 (N6095, N6081, N5844, N4913, N1274);
nor NOR4 (N6096, N6089, N321, N3172, N92);
nor NOR2 (N6097, N6065, N3274);
and AND3 (N6098, N6092, N3447, N3255);
not NOT1 (N6099, N6096);
nor NOR4 (N6100, N6098, N552, N2189, N1219);
nand NAND2 (N6101, N6075, N1691);
and AND2 (N6102, N6101, N3872);
nor NOR3 (N6103, N6095, N1445, N2489);
xor XOR2 (N6104, N6091, N688);
nor NOR4 (N6105, N6073, N4433, N3782, N974);
nor NOR3 (N6106, N6097, N3789, N5262);
nor NOR3 (N6107, N6100, N5971, N2668);
xor XOR2 (N6108, N6084, N5925);
nand NAND4 (N6109, N6105, N1002, N2483, N1490);
nor NOR3 (N6110, N6109, N2714, N1358);
or OR4 (N6111, N6102, N2, N3030, N5878);
buf BUF1 (N6112, N6110);
and AND4 (N6113, N6094, N394, N5706, N3198);
xor XOR2 (N6114, N6099, N5412);
nor NOR2 (N6115, N6108, N5365);
nor NOR3 (N6116, N6104, N2873, N2984);
or OR4 (N6117, N6111, N4049, N4773, N4405);
buf BUF1 (N6118, N6116);
xor XOR2 (N6119, N6115, N4615);
buf BUF1 (N6120, N6103);
nand NAND2 (N6121, N6113, N470);
nand NAND2 (N6122, N6083, N4376);
or OR3 (N6123, N6106, N1812, N4264);
nor NOR3 (N6124, N6114, N79, N4580);
buf BUF1 (N6125, N6123);
nand NAND3 (N6126, N6119, N3275, N5377);
nand NAND4 (N6127, N6121, N3244, N3826, N5442);
xor XOR2 (N6128, N6124, N4636);
and AND3 (N6129, N6118, N5156, N4257);
nor NOR4 (N6130, N6117, N504, N5828, N2524);
nand NAND4 (N6131, N6128, N487, N2897, N1070);
or OR2 (N6132, N6130, N2726);
not NOT1 (N6133, N6125);
not NOT1 (N6134, N6132);
nand NAND4 (N6135, N6133, N2865, N1327, N4178);
nand NAND2 (N6136, N6126, N4608);
xor XOR2 (N6137, N6107, N6074);
and AND3 (N6138, N6131, N4992, N1069);
not NOT1 (N6139, N6120);
not NOT1 (N6140, N6122);
not NOT1 (N6141, N6139);
xor XOR2 (N6142, N6129, N4941);
xor XOR2 (N6143, N6138, N3222);
buf BUF1 (N6144, N6112);
nand NAND3 (N6145, N6144, N358, N4372);
nor NOR3 (N6146, N6140, N5904, N2510);
xor XOR2 (N6147, N6141, N2172);
and AND3 (N6148, N6146, N3151, N2141);
nor NOR2 (N6149, N6136, N3176);
or OR4 (N6150, N6143, N2622, N3573, N1023);
nand NAND3 (N6151, N6145, N285, N2027);
and AND3 (N6152, N6150, N169, N6002);
xor XOR2 (N6153, N6151, N1335);
not NOT1 (N6154, N6148);
nor NOR2 (N6155, N6154, N2217);
xor XOR2 (N6156, N6127, N2585);
not NOT1 (N6157, N6149);
not NOT1 (N6158, N6142);
nor NOR4 (N6159, N6135, N5148, N3280, N6061);
nor NOR4 (N6160, N6157, N6006, N4528, N2811);
nand NAND4 (N6161, N6153, N2207, N2152, N4796);
xor XOR2 (N6162, N6159, N5604);
and AND2 (N6163, N6161, N5704);
and AND4 (N6164, N6158, N182, N627, N3182);
or OR2 (N6165, N6134, N1750);
or OR2 (N6166, N6147, N1489);
nand NAND2 (N6167, N6156, N3622);
and AND2 (N6168, N6162, N625);
and AND2 (N6169, N6155, N1152);
and AND4 (N6170, N6137, N4233, N3080, N2498);
nand NAND4 (N6171, N6166, N5642, N2488, N933);
or OR3 (N6172, N6167, N2728, N3663);
or OR4 (N6173, N6172, N301, N5432, N1180);
not NOT1 (N6174, N6160);
xor XOR2 (N6175, N6163, N2969);
not NOT1 (N6176, N6173);
not NOT1 (N6177, N6168);
nor NOR4 (N6178, N6165, N2959, N3136, N2168);
not NOT1 (N6179, N6178);
xor XOR2 (N6180, N6175, N2313);
nor NOR2 (N6181, N6164, N4262);
not NOT1 (N6182, N6171);
nand NAND3 (N6183, N6182, N6148, N3888);
buf BUF1 (N6184, N6176);
buf BUF1 (N6185, N6170);
nor NOR3 (N6186, N6180, N530, N4061);
buf BUF1 (N6187, N6185);
nand NAND4 (N6188, N6152, N4090, N3371, N5600);
or OR4 (N6189, N6187, N1403, N4083, N5421);
nand NAND4 (N6190, N6189, N437, N5249, N3696);
nand NAND4 (N6191, N6184, N3339, N5772, N359);
not NOT1 (N6192, N6177);
not NOT1 (N6193, N6174);
nand NAND4 (N6194, N6192, N2784, N2312, N3614);
xor XOR2 (N6195, N6181, N2137);
buf BUF1 (N6196, N6194);
xor XOR2 (N6197, N6186, N2518);
and AND4 (N6198, N6195, N2298, N3991, N750);
or OR3 (N6199, N6179, N5088, N2428);
or OR3 (N6200, N6196, N3239, N2664);
nor NOR2 (N6201, N6169, N1101);
and AND2 (N6202, N6200, N5099);
or OR4 (N6203, N6198, N2210, N1442, N1270);
nand NAND2 (N6204, N6197, N635);
or OR2 (N6205, N6188, N5813);
nand NAND4 (N6206, N6183, N337, N3283, N5302);
not NOT1 (N6207, N6205);
buf BUF1 (N6208, N6203);
buf BUF1 (N6209, N6202);
not NOT1 (N6210, N6193);
xor XOR2 (N6211, N6201, N4443);
or OR2 (N6212, N6208, N1243);
nor NOR3 (N6213, N6191, N5744, N3842);
nor NOR4 (N6214, N6211, N512, N4289, N4603);
nand NAND4 (N6215, N6212, N5783, N4319, N2966);
nand NAND4 (N6216, N6199, N1182, N1360, N3969);
or OR2 (N6217, N6213, N1144);
and AND4 (N6218, N6206, N2990, N5589, N2554);
buf BUF1 (N6219, N6207);
buf BUF1 (N6220, N6218);
not NOT1 (N6221, N6210);
and AND4 (N6222, N6219, N2536, N5867, N573);
nand NAND2 (N6223, N6214, N4766);
nor NOR2 (N6224, N6216, N326);
buf BUF1 (N6225, N6224);
and AND2 (N6226, N6204, N3718);
or OR2 (N6227, N6222, N5651);
xor XOR2 (N6228, N6220, N924);
and AND3 (N6229, N6225, N4311, N1090);
and AND3 (N6230, N6209, N6072, N6045);
nand NAND3 (N6231, N6217, N3548, N2768);
nor NOR4 (N6232, N6229, N2423, N4474, N4610);
and AND3 (N6233, N6226, N5772, N4174);
nor NOR3 (N6234, N6230, N1431, N2463);
buf BUF1 (N6235, N6228);
buf BUF1 (N6236, N6223);
and AND3 (N6237, N6234, N769, N563);
xor XOR2 (N6238, N6236, N1893);
nand NAND3 (N6239, N6238, N1930, N5668);
nand NAND2 (N6240, N6190, N2331);
nor NOR3 (N6241, N6231, N1102, N4543);
buf BUF1 (N6242, N6233);
nor NOR4 (N6243, N6242, N1259, N4148, N2692);
nor NOR3 (N6244, N6237, N4940, N3478);
not NOT1 (N6245, N6244);
buf BUF1 (N6246, N6232);
nand NAND4 (N6247, N6221, N1258, N5205, N1965);
buf BUF1 (N6248, N6246);
not NOT1 (N6249, N6239);
and AND4 (N6250, N6240, N4920, N132, N4567);
or OR2 (N6251, N6247, N5703);
xor XOR2 (N6252, N6235, N368);
not NOT1 (N6253, N6249);
xor XOR2 (N6254, N6253, N4807);
not NOT1 (N6255, N6248);
nand NAND3 (N6256, N6255, N3052, N3831);
not NOT1 (N6257, N6215);
buf BUF1 (N6258, N6251);
or OR2 (N6259, N6241, N2860);
and AND4 (N6260, N6227, N4112, N45, N3298);
not NOT1 (N6261, N6259);
and AND3 (N6262, N6252, N2799, N6126);
buf BUF1 (N6263, N6256);
not NOT1 (N6264, N6250);
xor XOR2 (N6265, N6258, N5191);
or OR4 (N6266, N6254, N2486, N505, N4995);
nand NAND2 (N6267, N6265, N2148);
nand NAND4 (N6268, N6267, N2335, N4083, N5144);
xor XOR2 (N6269, N6257, N448);
not NOT1 (N6270, N6243);
or OR4 (N6271, N6264, N5007, N2626, N3972);
or OR4 (N6272, N6245, N3302, N5266, N2769);
nor NOR3 (N6273, N6266, N2759, N2479);
not NOT1 (N6274, N6263);
xor XOR2 (N6275, N6271, N3994);
and AND3 (N6276, N6272, N4389, N3513);
nor NOR3 (N6277, N6269, N4183, N525);
buf BUF1 (N6278, N6273);
xor XOR2 (N6279, N6277, N6051);
or OR4 (N6280, N6274, N3861, N314, N4689);
xor XOR2 (N6281, N6275, N719);
or OR3 (N6282, N6276, N428, N193);
or OR4 (N6283, N6262, N550, N679, N5780);
and AND2 (N6284, N6260, N896);
nand NAND4 (N6285, N6280, N2505, N1772, N3565);
and AND3 (N6286, N6270, N1970, N1932);
nand NAND2 (N6287, N6278, N2794);
nand NAND3 (N6288, N6282, N1086, N3469);
or OR3 (N6289, N6283, N2547, N5307);
xor XOR2 (N6290, N6289, N821);
xor XOR2 (N6291, N6286, N3024);
and AND4 (N6292, N6261, N4429, N4501, N4846);
buf BUF1 (N6293, N6268);
or OR4 (N6294, N6287, N2047, N2674, N1320);
xor XOR2 (N6295, N6285, N1703);
or OR4 (N6296, N6295, N5214, N285, N1669);
or OR2 (N6297, N6288, N2834);
not NOT1 (N6298, N6291);
or OR3 (N6299, N6293, N148, N3031);
buf BUF1 (N6300, N6279);
not NOT1 (N6301, N6300);
nand NAND3 (N6302, N6290, N2119, N6059);
or OR2 (N6303, N6284, N4108);
xor XOR2 (N6304, N6292, N5811);
not NOT1 (N6305, N6296);
not NOT1 (N6306, N6299);
buf BUF1 (N6307, N6302);
or OR3 (N6308, N6297, N454, N298);
or OR2 (N6309, N6307, N2684);
nand NAND3 (N6310, N6301, N2122, N4422);
and AND2 (N6311, N6303, N5698);
nand NAND3 (N6312, N6308, N6064, N956);
and AND4 (N6313, N6304, N4878, N2454, N5485);
xor XOR2 (N6314, N6298, N220);
not NOT1 (N6315, N6310);
and AND2 (N6316, N6313, N1833);
buf BUF1 (N6317, N6305);
or OR3 (N6318, N6316, N2379, N2800);
buf BUF1 (N6319, N6294);
or OR2 (N6320, N6281, N2377);
nor NOR4 (N6321, N6312, N2769, N5290, N2647);
not NOT1 (N6322, N6321);
and AND3 (N6323, N6306, N4735, N4265);
and AND4 (N6324, N6317, N950, N3730, N3462);
nor NOR4 (N6325, N6315, N2226, N1592, N587);
xor XOR2 (N6326, N6325, N1242);
nand NAND4 (N6327, N6309, N6114, N5051, N87);
nor NOR4 (N6328, N6327, N1316, N61, N1769);
nor NOR3 (N6329, N6322, N1349, N5437);
nor NOR4 (N6330, N6329, N1368, N2892, N4032);
or OR2 (N6331, N6330, N4385);
or OR3 (N6332, N6331, N923, N5932);
nor NOR4 (N6333, N6323, N1032, N3214, N1155);
nor NOR4 (N6334, N6332, N291, N1786, N4421);
xor XOR2 (N6335, N6320, N1051);
xor XOR2 (N6336, N6333, N901);
not NOT1 (N6337, N6334);
buf BUF1 (N6338, N6336);
or OR2 (N6339, N6319, N4030);
not NOT1 (N6340, N6339);
or OR2 (N6341, N6311, N1043);
xor XOR2 (N6342, N6335, N167);
xor XOR2 (N6343, N6318, N4070);
nand NAND3 (N6344, N6328, N2410, N2351);
nand NAND2 (N6345, N6341, N3204);
nor NOR2 (N6346, N6340, N5673);
and AND3 (N6347, N6326, N5408, N3199);
nand NAND4 (N6348, N6342, N3770, N2683, N2237);
nand NAND4 (N6349, N6337, N4566, N892, N2470);
and AND2 (N6350, N6347, N4297);
or OR2 (N6351, N6346, N3932);
or OR2 (N6352, N6348, N3721);
not NOT1 (N6353, N6345);
or OR3 (N6354, N6349, N4592, N3989);
xor XOR2 (N6355, N6343, N736);
xor XOR2 (N6356, N6350, N1133);
buf BUF1 (N6357, N6356);
and AND2 (N6358, N6355, N224);
or OR4 (N6359, N6358, N406, N5372, N3433);
nor NOR3 (N6360, N6344, N1406, N536);
buf BUF1 (N6361, N6353);
xor XOR2 (N6362, N6351, N599);
and AND4 (N6363, N6352, N3172, N5913, N4298);
nand NAND4 (N6364, N6357, N5853, N2151, N2878);
nor NOR2 (N6365, N6359, N2413);
nand NAND2 (N6366, N6338, N3940);
nand NAND2 (N6367, N6354, N2802);
buf BUF1 (N6368, N6324);
and AND2 (N6369, N6367, N2338);
and AND2 (N6370, N6365, N6100);
or OR3 (N6371, N6361, N100, N4979);
buf BUF1 (N6372, N6364);
and AND3 (N6373, N6366, N5498, N2750);
or OR3 (N6374, N6369, N1859, N1508);
nor NOR4 (N6375, N6372, N2778, N4358, N4397);
buf BUF1 (N6376, N6314);
and AND3 (N6377, N6374, N4653, N1250);
and AND2 (N6378, N6363, N1413);
xor XOR2 (N6379, N6362, N4210);
not NOT1 (N6380, N6370);
nand NAND4 (N6381, N6360, N4110, N2978, N1703);
and AND2 (N6382, N6380, N6161);
buf BUF1 (N6383, N6373);
nand NAND3 (N6384, N6383, N3345, N3150);
xor XOR2 (N6385, N6384, N2856);
or OR3 (N6386, N6378, N4807, N1429);
not NOT1 (N6387, N6375);
nor NOR3 (N6388, N6379, N5890, N3726);
nand NAND2 (N6389, N6377, N2095);
nor NOR2 (N6390, N6382, N3418);
buf BUF1 (N6391, N6376);
or OR3 (N6392, N6381, N1604, N1451);
or OR2 (N6393, N6385, N1690);
buf BUF1 (N6394, N6389);
and AND2 (N6395, N6390, N1302);
xor XOR2 (N6396, N6393, N1388);
nand NAND3 (N6397, N6368, N4348, N4722);
or OR2 (N6398, N6396, N5077);
not NOT1 (N6399, N6397);
not NOT1 (N6400, N6395);
not NOT1 (N6401, N6387);
nand NAND3 (N6402, N6398, N5253, N5353);
buf BUF1 (N6403, N6402);
nand NAND3 (N6404, N6371, N4671, N2901);
and AND2 (N6405, N6403, N6042);
not NOT1 (N6406, N6386);
nor NOR4 (N6407, N6399, N1770, N988, N3834);
or OR4 (N6408, N6391, N5276, N2852, N5783);
or OR2 (N6409, N6392, N945);
and AND3 (N6410, N6408, N275, N597);
or OR4 (N6411, N6404, N3153, N1025, N2931);
xor XOR2 (N6412, N6406, N4759);
and AND2 (N6413, N6400, N6185);
nor NOR4 (N6414, N6409, N5482, N2585, N970);
nor NOR4 (N6415, N6413, N438, N2889, N4886);
or OR4 (N6416, N6410, N4366, N838, N3765);
nand NAND2 (N6417, N6412, N5698);
xor XOR2 (N6418, N6407, N6157);
not NOT1 (N6419, N6405);
not NOT1 (N6420, N6388);
nor NOR4 (N6421, N6394, N5956, N3043, N716);
not NOT1 (N6422, N6418);
not NOT1 (N6423, N6416);
buf BUF1 (N6424, N6422);
nand NAND4 (N6425, N6411, N4206, N3597, N2021);
xor XOR2 (N6426, N6417, N474);
buf BUF1 (N6427, N6425);
or OR3 (N6428, N6426, N6334, N1398);
or OR3 (N6429, N6423, N3860, N6044);
or OR3 (N6430, N6414, N4029, N2102);
and AND4 (N6431, N6427, N3533, N4413, N92);
or OR3 (N6432, N6415, N1601, N1876);
xor XOR2 (N6433, N6421, N5849);
or OR2 (N6434, N6430, N4258);
xor XOR2 (N6435, N6434, N1283);
nand NAND3 (N6436, N6419, N1095, N4215);
and AND4 (N6437, N6429, N1118, N342, N4410);
and AND2 (N6438, N6401, N2361);
nor NOR3 (N6439, N6438, N4641, N3543);
nor NOR3 (N6440, N6428, N5582, N2635);
not NOT1 (N6441, N6435);
nand NAND2 (N6442, N6437, N3023);
or OR3 (N6443, N6420, N1327, N2648);
or OR4 (N6444, N6424, N6, N4334, N2069);
not NOT1 (N6445, N6443);
buf BUF1 (N6446, N6431);
xor XOR2 (N6447, N6440, N848);
not NOT1 (N6448, N6447);
buf BUF1 (N6449, N6433);
buf BUF1 (N6450, N6448);
nor NOR4 (N6451, N6439, N249, N563, N4550);
xor XOR2 (N6452, N6432, N3187);
or OR2 (N6453, N6436, N6375);
and AND2 (N6454, N6450, N230);
not NOT1 (N6455, N6451);
and AND3 (N6456, N6444, N4207, N4794);
and AND2 (N6457, N6441, N1730);
and AND4 (N6458, N6457, N722, N1184, N799);
and AND2 (N6459, N6456, N1569);
and AND2 (N6460, N6458, N3121);
or OR4 (N6461, N6459, N5431, N6417, N3558);
not NOT1 (N6462, N6446);
nand NAND4 (N6463, N6453, N1663, N2874, N1276);
xor XOR2 (N6464, N6442, N3577);
xor XOR2 (N6465, N6463, N4880);
xor XOR2 (N6466, N6460, N1197);
buf BUF1 (N6467, N6455);
or OR3 (N6468, N6465, N4712, N3248);
and AND3 (N6469, N6452, N1412, N1583);
nand NAND3 (N6470, N6449, N5369, N3286);
and AND4 (N6471, N6445, N5463, N4184, N2897);
buf BUF1 (N6472, N6469);
xor XOR2 (N6473, N6461, N6113);
xor XOR2 (N6474, N6454, N3669);
or OR2 (N6475, N6468, N6343);
not NOT1 (N6476, N6466);
nand NAND3 (N6477, N6472, N3429, N34);
xor XOR2 (N6478, N6470, N188);
buf BUF1 (N6479, N6476);
and AND2 (N6480, N6462, N5136);
nand NAND4 (N6481, N6477, N3295, N4078, N1195);
or OR2 (N6482, N6481, N475);
buf BUF1 (N6483, N6479);
nor NOR3 (N6484, N6480, N4547, N94);
nor NOR2 (N6485, N6478, N428);
nor NOR2 (N6486, N6475, N2107);
buf BUF1 (N6487, N6471);
not NOT1 (N6488, N6482);
xor XOR2 (N6489, N6485, N6395);
not NOT1 (N6490, N6467);
nand NAND2 (N6491, N6488, N5519);
buf BUF1 (N6492, N6484);
or OR4 (N6493, N6483, N1246, N4275, N507);
nor NOR4 (N6494, N6487, N6119, N6135, N1749);
xor XOR2 (N6495, N6490, N304);
or OR3 (N6496, N6494, N5586, N1040);
xor XOR2 (N6497, N6474, N789);
buf BUF1 (N6498, N6497);
not NOT1 (N6499, N6496);
or OR4 (N6500, N6498, N775, N6454, N759);
buf BUF1 (N6501, N6491);
xor XOR2 (N6502, N6492, N2749);
and AND3 (N6503, N6473, N3697, N2203);
and AND2 (N6504, N6489, N1589);
or OR4 (N6505, N6499, N5579, N3421, N1441);
buf BUF1 (N6506, N6505);
not NOT1 (N6507, N6486);
nand NAND4 (N6508, N6500, N5472, N2899, N3069);
xor XOR2 (N6509, N6501, N431);
buf BUF1 (N6510, N6502);
xor XOR2 (N6511, N6508, N2297);
or OR4 (N6512, N6506, N1457, N740, N1803);
nor NOR2 (N6513, N6464, N6127);
xor XOR2 (N6514, N6510, N4107);
nor NOR2 (N6515, N6503, N1915);
xor XOR2 (N6516, N6493, N5941);
or OR4 (N6517, N6507, N3014, N5855, N2766);
not NOT1 (N6518, N6495);
nor NOR2 (N6519, N6509, N2698);
not NOT1 (N6520, N6504);
nor NOR3 (N6521, N6514, N5193, N2304);
nor NOR4 (N6522, N6517, N5195, N2066, N1367);
nor NOR2 (N6523, N6513, N1638);
and AND3 (N6524, N6520, N4508, N6513);
or OR4 (N6525, N6524, N6190, N1058, N4190);
and AND2 (N6526, N6522, N4181);
and AND3 (N6527, N6512, N2246, N451);
xor XOR2 (N6528, N6527, N4703);
and AND2 (N6529, N6526, N5307);
nand NAND2 (N6530, N6525, N4237);
and AND2 (N6531, N6523, N4691);
not NOT1 (N6532, N6511);
and AND4 (N6533, N6515, N573, N6522, N2334);
nor NOR3 (N6534, N6516, N993, N3870);
nor NOR2 (N6535, N6529, N5269);
xor XOR2 (N6536, N6533, N3295);
nand NAND2 (N6537, N6521, N1437);
xor XOR2 (N6538, N6532, N2747);
nand NAND4 (N6539, N6534, N3511, N3200, N1233);
not NOT1 (N6540, N6536);
buf BUF1 (N6541, N6518);
buf BUF1 (N6542, N6541);
buf BUF1 (N6543, N6540);
and AND3 (N6544, N6542, N2967, N2731);
not NOT1 (N6545, N6544);
not NOT1 (N6546, N6528);
and AND3 (N6547, N6535, N4065, N6543);
buf BUF1 (N6548, N4191);
buf BUF1 (N6549, N6547);
buf BUF1 (N6550, N6519);
buf BUF1 (N6551, N6531);
and AND2 (N6552, N6537, N832);
or OR2 (N6553, N6546, N3655);
and AND3 (N6554, N6552, N3585, N2381);
or OR2 (N6555, N6545, N6479);
xor XOR2 (N6556, N6554, N1103);
buf BUF1 (N6557, N6556);
buf BUF1 (N6558, N6555);
nand NAND4 (N6559, N6538, N1042, N639, N6420);
and AND2 (N6560, N6530, N5341);
nor NOR2 (N6561, N6548, N169);
xor XOR2 (N6562, N6549, N6167);
not NOT1 (N6563, N6560);
buf BUF1 (N6564, N6563);
not NOT1 (N6565, N6553);
buf BUF1 (N6566, N6557);
or OR4 (N6567, N6558, N4131, N2556, N6345);
nand NAND3 (N6568, N6566, N2100, N2086);
or OR4 (N6569, N6539, N2956, N5463, N3719);
and AND4 (N6570, N6561, N4964, N5364, N5839);
not NOT1 (N6571, N6567);
nand NAND4 (N6572, N6568, N2056, N2892, N2921);
and AND4 (N6573, N6571, N793, N1245, N2322);
buf BUF1 (N6574, N6570);
buf BUF1 (N6575, N6564);
not NOT1 (N6576, N6569);
buf BUF1 (N6577, N6551);
not NOT1 (N6578, N6577);
xor XOR2 (N6579, N6559, N1101);
and AND3 (N6580, N6578, N937, N5032);
nand NAND2 (N6581, N6573, N4997);
not NOT1 (N6582, N6576);
buf BUF1 (N6583, N6581);
not NOT1 (N6584, N6550);
nor NOR3 (N6585, N6580, N9, N859);
xor XOR2 (N6586, N6582, N1057);
and AND3 (N6587, N6583, N723, N2109);
xor XOR2 (N6588, N6562, N6124);
xor XOR2 (N6589, N6572, N2600);
or OR2 (N6590, N6586, N2984);
xor XOR2 (N6591, N6589, N2083);
nor NOR3 (N6592, N6590, N880, N2470);
xor XOR2 (N6593, N6592, N2436);
xor XOR2 (N6594, N6588, N303);
not NOT1 (N6595, N6594);
not NOT1 (N6596, N6579);
and AND4 (N6597, N6587, N79, N5793, N5905);
xor XOR2 (N6598, N6585, N4558);
xor XOR2 (N6599, N6565, N6260);
buf BUF1 (N6600, N6575);
not NOT1 (N6601, N6597);
nand NAND3 (N6602, N6598, N3629, N5929);
and AND4 (N6603, N6599, N1015, N5260, N2661);
and AND4 (N6604, N6596, N2675, N3418, N4172);
or OR3 (N6605, N6600, N2751, N4631);
not NOT1 (N6606, N6593);
nor NOR3 (N6607, N6603, N1430, N2382);
or OR3 (N6608, N6601, N6402, N2016);
and AND4 (N6609, N6607, N1857, N2706, N5060);
buf BUF1 (N6610, N6574);
not NOT1 (N6611, N6605);
and AND2 (N6612, N6604, N2419);
not NOT1 (N6613, N6608);
xor XOR2 (N6614, N6611, N948);
xor XOR2 (N6615, N6591, N5505);
nand NAND2 (N6616, N6609, N4287);
xor XOR2 (N6617, N6615, N872);
and AND4 (N6618, N6614, N71, N315, N1253);
not NOT1 (N6619, N6606);
or OR4 (N6620, N6612, N1791, N6184, N6324);
xor XOR2 (N6621, N6617, N3993);
xor XOR2 (N6622, N6619, N711);
xor XOR2 (N6623, N6618, N3317);
nor NOR3 (N6624, N6621, N852, N1851);
or OR2 (N6625, N6610, N159);
and AND2 (N6626, N6595, N2138);
and AND4 (N6627, N6616, N1260, N4342, N4552);
not NOT1 (N6628, N6613);
nor NOR3 (N6629, N6622, N829, N1322);
buf BUF1 (N6630, N6627);
nand NAND2 (N6631, N6584, N2617);
not NOT1 (N6632, N6602);
buf BUF1 (N6633, N6625);
and AND4 (N6634, N6629, N1770, N2689, N4738);
nor NOR4 (N6635, N6630, N251, N3037, N3014);
nor NOR2 (N6636, N6631, N3236);
nand NAND2 (N6637, N6623, N2025);
nand NAND3 (N6638, N6626, N3528, N6372);
nor NOR4 (N6639, N6638, N4891, N3150, N4553);
not NOT1 (N6640, N6635);
buf BUF1 (N6641, N6632);
and AND3 (N6642, N6633, N4876, N4568);
nor NOR4 (N6643, N6640, N2783, N5843, N1511);
or OR2 (N6644, N6642, N5494);
nor NOR4 (N6645, N6644, N3598, N2650, N1397);
not NOT1 (N6646, N6643);
not NOT1 (N6647, N6620);
or OR4 (N6648, N6637, N1806, N4609, N4967);
or OR4 (N6649, N6641, N1731, N4034, N4509);
or OR2 (N6650, N6624, N3759);
and AND3 (N6651, N6646, N6640, N165);
nand NAND2 (N6652, N6628, N1480);
not NOT1 (N6653, N6648);
or OR4 (N6654, N6653, N3812, N5842, N6509);
xor XOR2 (N6655, N6636, N2548);
nand NAND3 (N6656, N6654, N401, N2948);
buf BUF1 (N6657, N6651);
not NOT1 (N6658, N6645);
xor XOR2 (N6659, N6658, N4630);
or OR3 (N6660, N6656, N4797, N833);
nor NOR4 (N6661, N6655, N1440, N4444, N5112);
nand NAND2 (N6662, N6650, N1017);
not NOT1 (N6663, N6659);
xor XOR2 (N6664, N6647, N3073);
not NOT1 (N6665, N6649);
nand NAND4 (N6666, N6657, N3949, N2268, N3097);
and AND3 (N6667, N6666, N1047, N4189);
nor NOR3 (N6668, N6665, N1427, N6339);
xor XOR2 (N6669, N6664, N3777);
not NOT1 (N6670, N6667);
buf BUF1 (N6671, N6668);
and AND4 (N6672, N6670, N5240, N3928, N4752);
or OR2 (N6673, N6660, N4953);
not NOT1 (N6674, N6669);
or OR4 (N6675, N6672, N355, N942, N6607);
nor NOR4 (N6676, N6673, N1602, N2688, N740);
and AND2 (N6677, N6675, N5752);
not NOT1 (N6678, N6676);
buf BUF1 (N6679, N6639);
nand NAND4 (N6680, N6678, N3087, N3657, N1292);
not NOT1 (N6681, N6679);
or OR3 (N6682, N6652, N3878, N5717);
and AND2 (N6683, N6663, N1279);
not NOT1 (N6684, N6661);
buf BUF1 (N6685, N6683);
nand NAND2 (N6686, N6680, N231);
or OR3 (N6687, N6684, N4761, N2792);
or OR2 (N6688, N6686, N3500);
or OR2 (N6689, N6685, N3822);
and AND3 (N6690, N6682, N5620, N79);
and AND4 (N6691, N6689, N5219, N1296, N2622);
buf BUF1 (N6692, N6671);
nor NOR2 (N6693, N6674, N614);
buf BUF1 (N6694, N6691);
xor XOR2 (N6695, N6692, N1724);
buf BUF1 (N6696, N6693);
not NOT1 (N6697, N6688);
or OR3 (N6698, N6662, N1220, N5284);
or OR4 (N6699, N6697, N6460, N457, N760);
nand NAND4 (N6700, N6677, N5704, N3821, N4895);
nor NOR4 (N6701, N6696, N322, N2025, N6208);
xor XOR2 (N6702, N6695, N3815);
xor XOR2 (N6703, N6702, N6468);
xor XOR2 (N6704, N6690, N4709);
nor NOR3 (N6705, N6704, N1072, N5283);
nor NOR2 (N6706, N6694, N6367);
not NOT1 (N6707, N6703);
buf BUF1 (N6708, N6705);
not NOT1 (N6709, N6681);
buf BUF1 (N6710, N6687);
nor NOR3 (N6711, N6699, N2453, N2453);
buf BUF1 (N6712, N6707);
buf BUF1 (N6713, N6698);
or OR4 (N6714, N6701, N4149, N122, N587);
xor XOR2 (N6715, N6712, N5819);
and AND3 (N6716, N6708, N776, N5881);
nor NOR3 (N6717, N6713, N4906, N5213);
nor NOR2 (N6718, N6717, N4189);
or OR4 (N6719, N6634, N3245, N1986, N5741);
and AND4 (N6720, N6700, N1680, N2206, N150);
nor NOR2 (N6721, N6711, N2645);
and AND2 (N6722, N6715, N3507);
or OR4 (N6723, N6718, N4567, N3157, N4902);
not NOT1 (N6724, N6721);
and AND4 (N6725, N6724, N4057, N6703, N1055);
nor NOR2 (N6726, N6719, N5935);
nor NOR2 (N6727, N6720, N2951);
nor NOR4 (N6728, N6723, N1699, N3789, N748);
nand NAND3 (N6729, N6725, N945, N3253);
nand NAND4 (N6730, N6706, N6128, N1415, N2579);
xor XOR2 (N6731, N6727, N1620);
xor XOR2 (N6732, N6714, N3056);
not NOT1 (N6733, N6732);
and AND3 (N6734, N6729, N4318, N813);
or OR2 (N6735, N6733, N269);
nor NOR4 (N6736, N6709, N5640, N5161, N6614);
buf BUF1 (N6737, N6726);
xor XOR2 (N6738, N6736, N6054);
not NOT1 (N6739, N6710);
nor NOR3 (N6740, N6730, N1118, N3295);
and AND2 (N6741, N6737, N3463);
not NOT1 (N6742, N6722);
and AND4 (N6743, N6738, N616, N2356, N3097);
or OR3 (N6744, N6716, N2699, N2181);
not NOT1 (N6745, N6734);
not NOT1 (N6746, N6735);
not NOT1 (N6747, N6743);
nand NAND4 (N6748, N6740, N2973, N1239, N3509);
nand NAND2 (N6749, N6739, N5267);
or OR2 (N6750, N6731, N3722);
xor XOR2 (N6751, N6728, N1046);
or OR2 (N6752, N6746, N3811);
nor NOR4 (N6753, N6750, N6268, N1535, N2082);
nand NAND3 (N6754, N6751, N2516, N5071);
xor XOR2 (N6755, N6745, N5410);
nor NOR4 (N6756, N6744, N2917, N4911, N997);
xor XOR2 (N6757, N6741, N4134);
not NOT1 (N6758, N6752);
xor XOR2 (N6759, N6753, N3520);
buf BUF1 (N6760, N6756);
not NOT1 (N6761, N6748);
buf BUF1 (N6762, N6760);
or OR3 (N6763, N6742, N1693, N3915);
or OR3 (N6764, N6758, N2730, N2530);
or OR2 (N6765, N6761, N2809);
and AND3 (N6766, N6757, N4877, N2887);
nor NOR4 (N6767, N6765, N2546, N267, N2761);
or OR3 (N6768, N6755, N772, N5080);
buf BUF1 (N6769, N6762);
not NOT1 (N6770, N6759);
not NOT1 (N6771, N6767);
buf BUF1 (N6772, N6754);
and AND4 (N6773, N6771, N2907, N4015, N570);
nor NOR3 (N6774, N6747, N2899, N3017);
buf BUF1 (N6775, N6773);
and AND4 (N6776, N6749, N4003, N5786, N739);
xor XOR2 (N6777, N6774, N1324);
or OR3 (N6778, N6764, N4901, N309);
nor NOR3 (N6779, N6775, N6253, N2433);
not NOT1 (N6780, N6769);
or OR2 (N6781, N6778, N6012);
not NOT1 (N6782, N6780);
nor NOR2 (N6783, N6766, N5813);
or OR4 (N6784, N6782, N3231, N317, N6264);
or OR3 (N6785, N6768, N1037, N3876);
xor XOR2 (N6786, N6781, N705);
and AND4 (N6787, N6779, N5151, N285, N3220);
not NOT1 (N6788, N6776);
nor NOR3 (N6789, N6763, N3830, N3558);
buf BUF1 (N6790, N6788);
nand NAND2 (N6791, N6772, N3421);
nand NAND4 (N6792, N6785, N2916, N2089, N2936);
or OR2 (N6793, N6783, N33);
xor XOR2 (N6794, N6770, N3608);
not NOT1 (N6795, N6793);
and AND3 (N6796, N6794, N410, N851);
buf BUF1 (N6797, N6786);
or OR2 (N6798, N6784, N3130);
nand NAND2 (N6799, N6795, N796);
not NOT1 (N6800, N6791);
nand NAND2 (N6801, N6799, N3532);
or OR4 (N6802, N6800, N3301, N258, N1672);
buf BUF1 (N6803, N6796);
nor NOR2 (N6804, N6798, N4918);
not NOT1 (N6805, N6777);
and AND4 (N6806, N6787, N2520, N5516, N2908);
nand NAND4 (N6807, N6801, N1636, N6315, N4209);
not NOT1 (N6808, N6805);
not NOT1 (N6809, N6790);
buf BUF1 (N6810, N6808);
not NOT1 (N6811, N6797);
nand NAND3 (N6812, N6807, N2291, N4080);
and AND2 (N6813, N6810, N1610);
or OR2 (N6814, N6813, N4468);
xor XOR2 (N6815, N6806, N3792);
and AND4 (N6816, N6815, N3094, N2898, N5064);
xor XOR2 (N6817, N6812, N506);
nand NAND2 (N6818, N6811, N2643);
nand NAND4 (N6819, N6803, N6079, N3780, N997);
nor NOR2 (N6820, N6802, N3619);
or OR4 (N6821, N6789, N1947, N6307, N2454);
and AND3 (N6822, N6809, N1929, N5685);
or OR2 (N6823, N6818, N1864);
nor NOR4 (N6824, N6817, N1648, N6772, N4567);
buf BUF1 (N6825, N6804);
not NOT1 (N6826, N6792);
buf BUF1 (N6827, N6826);
nor NOR3 (N6828, N6827, N2777, N2373);
xor XOR2 (N6829, N6823, N5432);
and AND4 (N6830, N6821, N1937, N1254, N2511);
buf BUF1 (N6831, N6816);
and AND2 (N6832, N6822, N3500);
xor XOR2 (N6833, N6819, N1816);
buf BUF1 (N6834, N6829);
nand NAND4 (N6835, N6830, N1008, N1301, N2820);
buf BUF1 (N6836, N6820);
buf BUF1 (N6837, N6832);
xor XOR2 (N6838, N6814, N486);
xor XOR2 (N6839, N6833, N3184);
xor XOR2 (N6840, N6825, N1659);
and AND4 (N6841, N6838, N3367, N4075, N4814);
buf BUF1 (N6842, N6837);
xor XOR2 (N6843, N6835, N1419);
or OR2 (N6844, N6839, N996);
or OR2 (N6845, N6843, N5588);
nand NAND4 (N6846, N6841, N4879, N1157, N143);
or OR2 (N6847, N6844, N2411);
or OR3 (N6848, N6831, N4775, N2806);
nand NAND2 (N6849, N6834, N4290);
buf BUF1 (N6850, N6846);
or OR2 (N6851, N6849, N4780);
buf BUF1 (N6852, N6850);
nand NAND2 (N6853, N6840, N1471);
and AND2 (N6854, N6836, N1839);
and AND2 (N6855, N6851, N4245);
xor XOR2 (N6856, N6842, N6568);
not NOT1 (N6857, N6848);
nor NOR3 (N6858, N6857, N2437, N6188);
not NOT1 (N6859, N6847);
nand NAND4 (N6860, N6824, N6227, N959, N2919);
buf BUF1 (N6861, N6858);
nand NAND3 (N6862, N6828, N1308, N2268);
buf BUF1 (N6863, N6854);
xor XOR2 (N6864, N6863, N4679);
nor NOR4 (N6865, N6852, N1023, N300, N6122);
or OR3 (N6866, N6861, N5602, N2593);
xor XOR2 (N6867, N6859, N4761);
nand NAND3 (N6868, N6864, N5763, N5493);
not NOT1 (N6869, N6862);
and AND2 (N6870, N6855, N2026);
buf BUF1 (N6871, N6868);
buf BUF1 (N6872, N6871);
not NOT1 (N6873, N6856);
or OR3 (N6874, N6853, N5213, N3391);
or OR3 (N6875, N6870, N5552, N5735);
or OR2 (N6876, N6875, N5894);
nand NAND2 (N6877, N6865, N3465);
nand NAND3 (N6878, N6869, N6081, N410);
buf BUF1 (N6879, N6876);
nor NOR4 (N6880, N6867, N6075, N1556, N6652);
nand NAND2 (N6881, N6845, N5720);
not NOT1 (N6882, N6879);
xor XOR2 (N6883, N6880, N343);
xor XOR2 (N6884, N6866, N2502);
nor NOR2 (N6885, N6872, N6608);
nand NAND4 (N6886, N6885, N6826, N1129, N4085);
nand NAND2 (N6887, N6882, N2699);
not NOT1 (N6888, N6884);
not NOT1 (N6889, N6873);
or OR3 (N6890, N6860, N3206, N766);
buf BUF1 (N6891, N6886);
nor NOR3 (N6892, N6877, N1133, N6647);
xor XOR2 (N6893, N6881, N1427);
buf BUF1 (N6894, N6892);
not NOT1 (N6895, N6894);
xor XOR2 (N6896, N6888, N6868);
or OR3 (N6897, N6889, N1677, N5996);
and AND2 (N6898, N6896, N2406);
buf BUF1 (N6899, N6891);
and AND3 (N6900, N6899, N6309, N5015);
buf BUF1 (N6901, N6900);
not NOT1 (N6902, N6878);
nand NAND2 (N6903, N6874, N3560);
buf BUF1 (N6904, N6898);
not NOT1 (N6905, N6895);
not NOT1 (N6906, N6890);
not NOT1 (N6907, N6901);
nand NAND3 (N6908, N6897, N3165, N5441);
or OR3 (N6909, N6908, N2828, N6737);
and AND3 (N6910, N6905, N4452, N163);
xor XOR2 (N6911, N6907, N6475);
buf BUF1 (N6912, N6906);
nor NOR2 (N6913, N6910, N912);
and AND4 (N6914, N6893, N4520, N1400, N682);
nand NAND2 (N6915, N6911, N5888);
buf BUF1 (N6916, N6903);
or OR2 (N6917, N6915, N695);
buf BUF1 (N6918, N6904);
and AND2 (N6919, N6902, N5345);
buf BUF1 (N6920, N6916);
not NOT1 (N6921, N6917);
or OR3 (N6922, N6919, N1171, N296);
nand NAND2 (N6923, N6920, N152);
nand NAND4 (N6924, N6913, N2471, N4602, N5665);
nand NAND3 (N6925, N6883, N4118, N3651);
buf BUF1 (N6926, N6918);
xor XOR2 (N6927, N6887, N6206);
not NOT1 (N6928, N6924);
not NOT1 (N6929, N6921);
and AND3 (N6930, N6909, N333, N5704);
or OR2 (N6931, N6927, N2785);
or OR3 (N6932, N6928, N3707, N5135);
nor NOR4 (N6933, N6912, N5845, N5089, N4735);
or OR4 (N6934, N6925, N5842, N6331, N2677);
or OR4 (N6935, N6923, N6506, N6431, N6881);
or OR4 (N6936, N6932, N4594, N5657, N23);
nand NAND2 (N6937, N6935, N5238);
or OR2 (N6938, N6936, N4407);
or OR2 (N6939, N6934, N1218);
buf BUF1 (N6940, N6929);
and AND3 (N6941, N6931, N3700, N4268);
buf BUF1 (N6942, N6922);
nor NOR2 (N6943, N6926, N5246);
nor NOR4 (N6944, N6930, N3314, N6240, N6486);
xor XOR2 (N6945, N6939, N1108);
not NOT1 (N6946, N6942);
xor XOR2 (N6947, N6943, N1409);
or OR2 (N6948, N6914, N5807);
buf BUF1 (N6949, N6933);
nand NAND2 (N6950, N6949, N5716);
not NOT1 (N6951, N6941);
nand NAND2 (N6952, N6938, N4800);
xor XOR2 (N6953, N6940, N5122);
xor XOR2 (N6954, N6944, N1877);
not NOT1 (N6955, N6947);
xor XOR2 (N6956, N6946, N6835);
xor XOR2 (N6957, N6953, N5522);
nor NOR3 (N6958, N6948, N4772, N2938);
buf BUF1 (N6959, N6950);
or OR2 (N6960, N6952, N730);
nand NAND2 (N6961, N6955, N2343);
or OR4 (N6962, N6957, N4094, N1254, N5018);
not NOT1 (N6963, N6962);
xor XOR2 (N6964, N6959, N6907);
and AND3 (N6965, N6945, N6186, N3367);
or OR4 (N6966, N6960, N299, N2253, N1028);
xor XOR2 (N6967, N6958, N4968);
not NOT1 (N6968, N6965);
nand NAND2 (N6969, N6963, N6124);
or OR3 (N6970, N6954, N3947, N3710);
buf BUF1 (N6971, N6951);
and AND4 (N6972, N6966, N5494, N5342, N1086);
nor NOR2 (N6973, N6969, N1472);
buf BUF1 (N6974, N6971);
or OR2 (N6975, N6973, N3825);
or OR2 (N6976, N6964, N3343);
or OR3 (N6977, N6976, N1142, N1376);
nand NAND3 (N6978, N6968, N349, N1757);
nor NOR4 (N6979, N6937, N5454, N2499, N1384);
and AND4 (N6980, N6967, N5525, N898, N1364);
and AND2 (N6981, N6972, N78);
or OR3 (N6982, N6978, N6962, N8);
nor NOR4 (N6983, N6974, N2908, N3069, N5999);
buf BUF1 (N6984, N6981);
buf BUF1 (N6985, N6980);
nand NAND4 (N6986, N6979, N6650, N3508, N4646);
buf BUF1 (N6987, N6961);
buf BUF1 (N6988, N6983);
xor XOR2 (N6989, N6988, N829);
buf BUF1 (N6990, N6986);
not NOT1 (N6991, N6956);
nand NAND2 (N6992, N6984, N2501);
not NOT1 (N6993, N6985);
not NOT1 (N6994, N6970);
buf BUF1 (N6995, N6994);
nand NAND3 (N6996, N6993, N756, N164);
nand NAND2 (N6997, N6989, N2817);
and AND2 (N6998, N6996, N5267);
not NOT1 (N6999, N6992);
nand NAND2 (N7000, N6991, N2253);
not NOT1 (N7001, N6982);
and AND3 (N7002, N6990, N766, N5608);
xor XOR2 (N7003, N6977, N3955);
nor NOR4 (N7004, N6997, N3292, N5900, N2688);
and AND4 (N7005, N6998, N495, N1644, N2420);
not NOT1 (N7006, N6975);
buf BUF1 (N7007, N7003);
or OR3 (N7008, N7004, N1239, N1586);
or OR4 (N7009, N7005, N1845, N2876, N1915);
buf BUF1 (N7010, N7008);
or OR4 (N7011, N6999, N4372, N2144, N4026);
and AND4 (N7012, N7007, N5175, N3194, N3619);
xor XOR2 (N7013, N6995, N3611);
and AND4 (N7014, N7011, N1118, N2785, N2217);
or OR2 (N7015, N7006, N1863);
or OR4 (N7016, N7001, N3145, N755, N1686);
nand NAND4 (N7017, N7000, N4622, N4553, N1485);
buf BUF1 (N7018, N7010);
and AND3 (N7019, N7015, N2233, N2431);
and AND4 (N7020, N7018, N1667, N2271, N6576);
not NOT1 (N7021, N7009);
not NOT1 (N7022, N7021);
or OR3 (N7023, N7013, N133, N6320);
not NOT1 (N7024, N7002);
or OR3 (N7025, N7016, N2006, N1478);
and AND3 (N7026, N7025, N6889, N2378);
nand NAND3 (N7027, N7012, N1220, N3855);
xor XOR2 (N7028, N7022, N4711);
or OR3 (N7029, N7019, N1510, N4841);
and AND3 (N7030, N7028, N6883, N3341);
nand NAND4 (N7031, N7014, N467, N5670, N5319);
or OR3 (N7032, N7017, N6511, N6997);
nor NOR2 (N7033, N7031, N4066);
nand NAND2 (N7034, N7032, N5562);
nor NOR2 (N7035, N7024, N4639);
not NOT1 (N7036, N7035);
not NOT1 (N7037, N7026);
or OR2 (N7038, N7036, N3111);
nor NOR2 (N7039, N7027, N5363);
or OR3 (N7040, N7037, N7023, N844);
and AND2 (N7041, N413, N5827);
not NOT1 (N7042, N7030);
buf BUF1 (N7043, N7039);
nand NAND2 (N7044, N7029, N3041);
buf BUF1 (N7045, N7038);
xor XOR2 (N7046, N7044, N3671);
and AND2 (N7047, N7040, N3678);
xor XOR2 (N7048, N7033, N4387);
nor NOR3 (N7049, N7046, N5532, N5529);
xor XOR2 (N7050, N7047, N5065);
buf BUF1 (N7051, N6987);
or OR2 (N7052, N7050, N3559);
nand NAND3 (N7053, N7049, N2600, N1549);
nand NAND3 (N7054, N7020, N5329, N3031);
not NOT1 (N7055, N7054);
not NOT1 (N7056, N7034);
or OR4 (N7057, N7041, N3031, N5384, N4104);
nor NOR4 (N7058, N7056, N1472, N2347, N6003);
nor NOR4 (N7059, N7053, N1732, N5924, N2326);
nor NOR4 (N7060, N7043, N6213, N3833, N5741);
xor XOR2 (N7061, N7059, N3894);
or OR4 (N7062, N7060, N1531, N1621, N6814);
or OR2 (N7063, N7062, N2607);
buf BUF1 (N7064, N7063);
not NOT1 (N7065, N7055);
not NOT1 (N7066, N7051);
buf BUF1 (N7067, N7066);
nor NOR4 (N7068, N7058, N4802, N6799, N5033);
and AND4 (N7069, N7057, N6319, N6292, N4739);
or OR3 (N7070, N7067, N6820, N211);
or OR3 (N7071, N7070, N3659, N1712);
xor XOR2 (N7072, N7061, N1327);
nand NAND2 (N7073, N7068, N5053);
not NOT1 (N7074, N7069);
buf BUF1 (N7075, N7074);
and AND3 (N7076, N7045, N3772, N5776);
nor NOR3 (N7077, N7042, N4856, N3609);
xor XOR2 (N7078, N7076, N4257);
and AND3 (N7079, N7064, N3155, N6406);
and AND2 (N7080, N7052, N1838);
buf BUF1 (N7081, N7077);
xor XOR2 (N7082, N7065, N2931);
nand NAND4 (N7083, N7072, N4201, N1842, N350);
buf BUF1 (N7084, N7080);
nor NOR2 (N7085, N7079, N6630);
or OR3 (N7086, N7082, N1959, N4883);
buf BUF1 (N7087, N7085);
buf BUF1 (N7088, N7073);
xor XOR2 (N7089, N7071, N2135);
xor XOR2 (N7090, N7089, N655);
xor XOR2 (N7091, N7078, N5579);
nand NAND3 (N7092, N7084, N6809, N1726);
and AND3 (N7093, N7092, N1921, N1053);
nand NAND3 (N7094, N7081, N3747, N3873);
xor XOR2 (N7095, N7088, N6780);
xor XOR2 (N7096, N7086, N698);
or OR2 (N7097, N7075, N154);
nand NAND2 (N7098, N7097, N1438);
buf BUF1 (N7099, N7048);
not NOT1 (N7100, N7095);
buf BUF1 (N7101, N7096);
or OR4 (N7102, N7090, N2621, N5728, N5999);
xor XOR2 (N7103, N7099, N6086);
or OR2 (N7104, N7100, N6529);
xor XOR2 (N7105, N7094, N996);
nand NAND2 (N7106, N7105, N3474);
buf BUF1 (N7107, N7098);
nand NAND3 (N7108, N7093, N4623, N2534);
buf BUF1 (N7109, N7106);
xor XOR2 (N7110, N7101, N4635);
xor XOR2 (N7111, N7104, N2168);
not NOT1 (N7112, N7087);
xor XOR2 (N7113, N7083, N6938);
xor XOR2 (N7114, N7107, N7000);
nor NOR3 (N7115, N7091, N790, N6608);
buf BUF1 (N7116, N7110);
buf BUF1 (N7117, N7111);
not NOT1 (N7118, N7109);
xor XOR2 (N7119, N7115, N6469);
nor NOR3 (N7120, N7118, N1774, N3150);
nor NOR3 (N7121, N7112, N5422, N3726);
nand NAND2 (N7122, N7120, N1944);
not NOT1 (N7123, N7114);
or OR2 (N7124, N7116, N123);
nand NAND3 (N7125, N7102, N1631, N7034);
not NOT1 (N7126, N7108);
not NOT1 (N7127, N7122);
not NOT1 (N7128, N7127);
and AND4 (N7129, N7128, N4889, N406, N5292);
buf BUF1 (N7130, N7113);
and AND3 (N7131, N7121, N1077, N897);
nor NOR3 (N7132, N7130, N6129, N4156);
not NOT1 (N7133, N7103);
or OR2 (N7134, N7131, N6384);
or OR3 (N7135, N7123, N5626, N2020);
xor XOR2 (N7136, N7133, N5457);
not NOT1 (N7137, N7136);
nand NAND3 (N7138, N7137, N6382, N3248);
nor NOR2 (N7139, N7129, N2472);
xor XOR2 (N7140, N7124, N3009);
or OR3 (N7141, N7140, N3742, N180);
not NOT1 (N7142, N7134);
buf BUF1 (N7143, N7119);
and AND3 (N7144, N7139, N5847, N7085);
or OR2 (N7145, N7138, N258);
buf BUF1 (N7146, N7132);
and AND2 (N7147, N7144, N5530);
or OR2 (N7148, N7147, N1790);
nor NOR4 (N7149, N7125, N55, N6060, N5242);
not NOT1 (N7150, N7143);
nor NOR4 (N7151, N7149, N2473, N3030, N6542);
not NOT1 (N7152, N7146);
or OR2 (N7153, N7150, N4400);
or OR3 (N7154, N7151, N2624, N3457);
nand NAND4 (N7155, N7117, N5248, N3014, N6307);
and AND3 (N7156, N7142, N6345, N393);
xor XOR2 (N7157, N7152, N1000);
or OR2 (N7158, N7148, N3832);
and AND4 (N7159, N7158, N5047, N2991, N993);
nor NOR4 (N7160, N7154, N5989, N5132, N6626);
not NOT1 (N7161, N7156);
nor NOR2 (N7162, N7155, N6210);
nor NOR4 (N7163, N7135, N4540, N6483, N4897);
nor NOR2 (N7164, N7161, N4539);
and AND4 (N7165, N7160, N1628, N3852, N3035);
nand NAND4 (N7166, N7141, N5189, N460, N6932);
nor NOR3 (N7167, N7166, N5881, N2051);
buf BUF1 (N7168, N7153);
not NOT1 (N7169, N7126);
nor NOR3 (N7170, N7157, N6796, N6992);
or OR2 (N7171, N7162, N1096);
nand NAND2 (N7172, N7145, N3447);
and AND3 (N7173, N7171, N728, N4668);
buf BUF1 (N7174, N7164);
buf BUF1 (N7175, N7167);
nand NAND2 (N7176, N7172, N5493);
buf BUF1 (N7177, N7170);
and AND3 (N7178, N7163, N1440, N4369);
and AND3 (N7179, N7169, N1361, N5328);
nand NAND2 (N7180, N7168, N6454);
and AND2 (N7181, N7174, N410);
buf BUF1 (N7182, N7178);
xor XOR2 (N7183, N7176, N1213);
and AND2 (N7184, N7181, N1090);
nand NAND2 (N7185, N7175, N6411);
buf BUF1 (N7186, N7185);
not NOT1 (N7187, N7186);
buf BUF1 (N7188, N7159);
buf BUF1 (N7189, N7187);
not NOT1 (N7190, N7183);
nor NOR2 (N7191, N7180, N3220);
xor XOR2 (N7192, N7191, N7017);
not NOT1 (N7193, N7182);
xor XOR2 (N7194, N7184, N5126);
nand NAND2 (N7195, N7189, N6827);
not NOT1 (N7196, N7190);
nor NOR3 (N7197, N7196, N2161, N1044);
or OR2 (N7198, N7193, N4571);
buf BUF1 (N7199, N7188);
or OR3 (N7200, N7198, N878, N2317);
xor XOR2 (N7201, N7195, N3868);
xor XOR2 (N7202, N7177, N3001);
or OR3 (N7203, N7197, N5684, N217);
nand NAND2 (N7204, N7179, N3392);
or OR4 (N7205, N7192, N2592, N3582, N6593);
nor NOR2 (N7206, N7201, N3419);
and AND3 (N7207, N7200, N4147, N666);
buf BUF1 (N7208, N7203);
xor XOR2 (N7209, N7206, N5969);
nand NAND4 (N7210, N7202, N5792, N376, N2772);
xor XOR2 (N7211, N7207, N458);
or OR2 (N7212, N7205, N4914);
or OR4 (N7213, N7165, N7167, N2681, N4013);
and AND3 (N7214, N7213, N1249, N1938);
nor NOR4 (N7215, N7209, N2580, N3760, N6296);
nand NAND3 (N7216, N7212, N4579, N805);
not NOT1 (N7217, N7211);
nor NOR3 (N7218, N7215, N12, N5977);
buf BUF1 (N7219, N7214);
nor NOR2 (N7220, N7208, N4639);
not NOT1 (N7221, N7220);
or OR2 (N7222, N7194, N3260);
and AND4 (N7223, N7173, N1340, N2798, N4852);
xor XOR2 (N7224, N7216, N2325);
and AND3 (N7225, N7221, N3712, N4480);
xor XOR2 (N7226, N7210, N364);
xor XOR2 (N7227, N7217, N2276);
nand NAND2 (N7228, N7225, N5471);
or OR2 (N7229, N7227, N4783);
xor XOR2 (N7230, N7204, N2075);
and AND4 (N7231, N7199, N4943, N2664, N1298);
not NOT1 (N7232, N7219);
nor NOR4 (N7233, N7232, N893, N2947, N4361);
nor NOR2 (N7234, N7223, N2292);
or OR4 (N7235, N7229, N143, N2698, N3068);
xor XOR2 (N7236, N7230, N3729);
buf BUF1 (N7237, N7234);
and AND3 (N7238, N7235, N6038, N2592);
and AND2 (N7239, N7231, N441);
or OR3 (N7240, N7233, N6364, N284);
buf BUF1 (N7241, N7224);
not NOT1 (N7242, N7238);
nor NOR4 (N7243, N7240, N2077, N6345, N7095);
not NOT1 (N7244, N7218);
nor NOR3 (N7245, N7222, N5003, N282);
xor XOR2 (N7246, N7236, N2309);
xor XOR2 (N7247, N7228, N4391);
buf BUF1 (N7248, N7245);
nand NAND2 (N7249, N7247, N4626);
nor NOR3 (N7250, N7243, N6916, N2021);
and AND4 (N7251, N7246, N4089, N732, N6649);
or OR2 (N7252, N7244, N2463);
not NOT1 (N7253, N7237);
nor NOR2 (N7254, N7251, N3658);
and AND2 (N7255, N7241, N871);
nand NAND4 (N7256, N7226, N1015, N2472, N4921);
not NOT1 (N7257, N7249);
not NOT1 (N7258, N7254);
nor NOR4 (N7259, N7242, N7037, N6064, N4650);
xor XOR2 (N7260, N7257, N4518);
or OR4 (N7261, N7259, N6056, N5949, N697);
not NOT1 (N7262, N7261);
buf BUF1 (N7263, N7262);
buf BUF1 (N7264, N7258);
buf BUF1 (N7265, N7264);
or OR3 (N7266, N7260, N6815, N5673);
xor XOR2 (N7267, N7256, N6888);
not NOT1 (N7268, N7250);
and AND4 (N7269, N7239, N1092, N5268, N5711);
buf BUF1 (N7270, N7265);
and AND2 (N7271, N7268, N3512);
nor NOR4 (N7272, N7270, N6969, N7177, N2070);
and AND2 (N7273, N7263, N5361);
buf BUF1 (N7274, N7266);
or OR4 (N7275, N7271, N2194, N6390, N4420);
nand NAND4 (N7276, N7267, N2106, N5148, N1864);
or OR2 (N7277, N7248, N294);
and AND3 (N7278, N7253, N633, N904);
xor XOR2 (N7279, N7276, N4119);
and AND2 (N7280, N7274, N6458);
or OR4 (N7281, N7272, N1991, N6071, N4508);
not NOT1 (N7282, N7275);
not NOT1 (N7283, N7277);
xor XOR2 (N7284, N7273, N2854);
nor NOR3 (N7285, N7252, N2821, N6158);
buf BUF1 (N7286, N7279);
or OR4 (N7287, N7281, N4781, N1765, N2458);
buf BUF1 (N7288, N7284);
buf BUF1 (N7289, N7283);
buf BUF1 (N7290, N7289);
not NOT1 (N7291, N7282);
nor NOR3 (N7292, N7290, N876, N852);
buf BUF1 (N7293, N7255);
not NOT1 (N7294, N7288);
nor NOR4 (N7295, N7278, N785, N2053, N857);
and AND3 (N7296, N7295, N109, N1154);
nor NOR3 (N7297, N7293, N5392, N7243);
and AND4 (N7298, N7296, N7030, N3117, N5051);
or OR4 (N7299, N7269, N143, N3733, N4253);
xor XOR2 (N7300, N7292, N5348);
and AND3 (N7301, N7298, N6607, N5122);
and AND4 (N7302, N7299, N4979, N1378, N2802);
nand NAND2 (N7303, N7280, N4082);
xor XOR2 (N7304, N7297, N7256);
and AND3 (N7305, N7286, N2357, N1486);
nand NAND3 (N7306, N7285, N3833, N11);
buf BUF1 (N7307, N7302);
or OR2 (N7308, N7305, N5442);
or OR3 (N7309, N7304, N6356, N1621);
xor XOR2 (N7310, N7294, N6563);
nor NOR2 (N7311, N7309, N3739);
buf BUF1 (N7312, N7291);
not NOT1 (N7313, N7300);
xor XOR2 (N7314, N7310, N3879);
and AND4 (N7315, N7313, N7226, N3229, N1943);
nand NAND2 (N7316, N7308, N5938);
nand NAND2 (N7317, N7314, N5451);
or OR2 (N7318, N7306, N5878);
nand NAND2 (N7319, N7311, N247);
or OR4 (N7320, N7287, N740, N3233, N3803);
xor XOR2 (N7321, N7317, N4263);
nand NAND4 (N7322, N7303, N3063, N3739, N5724);
buf BUF1 (N7323, N7322);
buf BUF1 (N7324, N7301);
or OR4 (N7325, N7321, N1030, N4509, N303);
and AND4 (N7326, N7312, N169, N6869, N4266);
not NOT1 (N7327, N7307);
nand NAND4 (N7328, N7324, N919, N2760, N6976);
buf BUF1 (N7329, N7318);
nor NOR2 (N7330, N7315, N4813);
and AND4 (N7331, N7327, N4915, N2653, N1706);
and AND4 (N7332, N7326, N2294, N4026, N4377);
and AND3 (N7333, N7332, N1693, N5175);
not NOT1 (N7334, N7330);
not NOT1 (N7335, N7334);
buf BUF1 (N7336, N7320);
nor NOR3 (N7337, N7336, N2874, N5357);
nor NOR4 (N7338, N7337, N5076, N5389, N2244);
and AND4 (N7339, N7328, N3340, N6646, N3595);
buf BUF1 (N7340, N7333);
not NOT1 (N7341, N7325);
or OR4 (N7342, N7329, N4793, N6752, N6450);
not NOT1 (N7343, N7341);
or OR2 (N7344, N7343, N6990);
not NOT1 (N7345, N7344);
or OR4 (N7346, N7342, N2277, N1887, N7107);
xor XOR2 (N7347, N7331, N7046);
not NOT1 (N7348, N7338);
not NOT1 (N7349, N7323);
and AND3 (N7350, N7346, N168, N171);
xor XOR2 (N7351, N7348, N3497);
nor NOR4 (N7352, N7345, N7308, N6464, N3006);
nand NAND3 (N7353, N7316, N5957, N6202);
not NOT1 (N7354, N7351);
nand NAND2 (N7355, N7354, N3668);
and AND4 (N7356, N7347, N6830, N1397, N4428);
not NOT1 (N7357, N7349);
and AND4 (N7358, N7339, N3855, N43, N5844);
nor NOR2 (N7359, N7356, N3289);
nor NOR2 (N7360, N7358, N4157);
xor XOR2 (N7361, N7360, N784);
nand NAND4 (N7362, N7359, N1017, N6759, N5199);
xor XOR2 (N7363, N7353, N6865);
not NOT1 (N7364, N7319);
not NOT1 (N7365, N7355);
xor XOR2 (N7366, N7350, N3184);
and AND2 (N7367, N7364, N2250);
not NOT1 (N7368, N7363);
not NOT1 (N7369, N7352);
nor NOR2 (N7370, N7362, N5206);
buf BUF1 (N7371, N7361);
nand NAND4 (N7372, N7357, N2537, N5137, N3731);
and AND4 (N7373, N7372, N4507, N3154, N6767);
xor XOR2 (N7374, N7365, N7093);
and AND2 (N7375, N7366, N1407);
nor NOR2 (N7376, N7371, N4928);
and AND2 (N7377, N7369, N3232);
nand NAND4 (N7378, N7375, N2464, N3993, N1195);
not NOT1 (N7379, N7335);
not NOT1 (N7380, N7378);
and AND3 (N7381, N7380, N6337, N1156);
not NOT1 (N7382, N7370);
nand NAND4 (N7383, N7381, N5845, N5550, N1728);
xor XOR2 (N7384, N7373, N6057);
not NOT1 (N7385, N7368);
nor NOR4 (N7386, N7377, N3804, N4401, N4766);
xor XOR2 (N7387, N7340, N3853);
and AND3 (N7388, N7382, N4458, N356);
nand NAND3 (N7389, N7384, N7340, N5192);
nand NAND4 (N7390, N7389, N4438, N3538, N540);
nor NOR4 (N7391, N7388, N6046, N571, N1128);
xor XOR2 (N7392, N7391, N2682);
or OR3 (N7393, N7379, N6158, N737);
and AND2 (N7394, N7386, N4422);
and AND2 (N7395, N7387, N2407);
not NOT1 (N7396, N7376);
or OR3 (N7397, N7367, N1800, N777);
or OR2 (N7398, N7374, N4888);
or OR4 (N7399, N7392, N3432, N7188, N1483);
or OR3 (N7400, N7395, N569, N5889);
nor NOR3 (N7401, N7385, N5650, N5722);
xor XOR2 (N7402, N7396, N2952);
and AND4 (N7403, N7390, N4094, N5412, N3735);
not NOT1 (N7404, N7383);
nand NAND4 (N7405, N7393, N5340, N178, N7065);
buf BUF1 (N7406, N7394);
and AND2 (N7407, N7400, N5605);
nand NAND3 (N7408, N7397, N827, N2649);
nor NOR4 (N7409, N7408, N3940, N4713, N4728);
xor XOR2 (N7410, N7409, N6398);
buf BUF1 (N7411, N7405);
xor XOR2 (N7412, N7403, N3093);
nor NOR2 (N7413, N7402, N6201);
buf BUF1 (N7414, N7413);
and AND2 (N7415, N7401, N3233);
and AND3 (N7416, N7411, N6746, N3208);
xor XOR2 (N7417, N7407, N6104);
xor XOR2 (N7418, N7410, N3018);
and AND4 (N7419, N7417, N4124, N3535, N305);
xor XOR2 (N7420, N7412, N2875);
not NOT1 (N7421, N7414);
xor XOR2 (N7422, N7418, N5743);
not NOT1 (N7423, N7420);
buf BUF1 (N7424, N7415);
nor NOR2 (N7425, N7419, N4311);
nor NOR4 (N7426, N7399, N3918, N4672, N1929);
nand NAND2 (N7427, N7421, N2237);
buf BUF1 (N7428, N7425);
nand NAND2 (N7429, N7422, N3735);
not NOT1 (N7430, N7404);
buf BUF1 (N7431, N7429);
buf BUF1 (N7432, N7416);
and AND4 (N7433, N7406, N5521, N2398, N111);
not NOT1 (N7434, N7423);
nand NAND3 (N7435, N7428, N5099, N4467);
and AND2 (N7436, N7432, N5790);
and AND3 (N7437, N7426, N2293, N6542);
buf BUF1 (N7438, N7430);
xor XOR2 (N7439, N7431, N6817);
not NOT1 (N7440, N7434);
not NOT1 (N7441, N7424);
not NOT1 (N7442, N7439);
xor XOR2 (N7443, N7437, N5680);
or OR4 (N7444, N7440, N6993, N2715, N6581);
nor NOR3 (N7445, N7438, N178, N677);
xor XOR2 (N7446, N7435, N3532);
buf BUF1 (N7447, N7398);
nand NAND2 (N7448, N7447, N2273);
nor NOR4 (N7449, N7427, N3411, N6809, N4024);
xor XOR2 (N7450, N7433, N6934);
buf BUF1 (N7451, N7442);
and AND4 (N7452, N7451, N7077, N3997, N7107);
nand NAND2 (N7453, N7450, N3311);
nor NOR3 (N7454, N7444, N483, N5214);
or OR4 (N7455, N7454, N623, N5687, N6479);
or OR2 (N7456, N7452, N7454);
not NOT1 (N7457, N7456);
not NOT1 (N7458, N7441);
or OR3 (N7459, N7436, N3253, N6482);
xor XOR2 (N7460, N7445, N499);
or OR4 (N7461, N7453, N5575, N936, N4675);
or OR2 (N7462, N7446, N5526);
nor NOR2 (N7463, N7462, N7066);
buf BUF1 (N7464, N7449);
buf BUF1 (N7465, N7464);
buf BUF1 (N7466, N7443);
buf BUF1 (N7467, N7459);
not NOT1 (N7468, N7461);
buf BUF1 (N7469, N7458);
and AND3 (N7470, N7468, N1163, N3709);
buf BUF1 (N7471, N7455);
and AND4 (N7472, N7457, N5341, N3688, N4645);
or OR3 (N7473, N7467, N6402, N3087);
nor NOR3 (N7474, N7463, N3019, N3893);
nand NAND4 (N7475, N7448, N3499, N1916, N7060);
nand NAND4 (N7476, N7466, N6724, N5208, N4499);
buf BUF1 (N7477, N7473);
and AND3 (N7478, N7460, N1364, N5531);
buf BUF1 (N7479, N7476);
or OR4 (N7480, N7471, N6215, N3109, N569);
and AND3 (N7481, N7472, N2094, N2226);
or OR3 (N7482, N7474, N3680, N2056);
or OR4 (N7483, N7475, N4548, N5820, N3076);
nor NOR2 (N7484, N7465, N3532);
xor XOR2 (N7485, N7469, N1455);
buf BUF1 (N7486, N7477);
nand NAND3 (N7487, N7483, N5040, N1712);
and AND4 (N7488, N7478, N2124, N2710, N237);
and AND2 (N7489, N7485, N7070);
or OR3 (N7490, N7470, N6353, N864);
buf BUF1 (N7491, N7480);
buf BUF1 (N7492, N7479);
or OR3 (N7493, N7490, N835, N6951);
and AND4 (N7494, N7491, N3807, N4242, N4573);
or OR4 (N7495, N7484, N6400, N3709, N139);
nor NOR4 (N7496, N7481, N4479, N5929, N55);
not NOT1 (N7497, N7492);
not NOT1 (N7498, N7494);
or OR2 (N7499, N7498, N2298);
buf BUF1 (N7500, N7496);
nor NOR4 (N7501, N7495, N4055, N394, N1994);
nand NAND4 (N7502, N7499, N7283, N5996, N2805);
and AND2 (N7503, N7487, N3418);
or OR4 (N7504, N7502, N2003, N1540, N5729);
nor NOR2 (N7505, N7482, N1828);
not NOT1 (N7506, N7493);
buf BUF1 (N7507, N7501);
buf BUF1 (N7508, N7488);
nand NAND4 (N7509, N7486, N3053, N4171, N2390);
nand NAND3 (N7510, N7503, N5353, N492);
xor XOR2 (N7511, N7504, N7391);
nand NAND4 (N7512, N7505, N6650, N498, N2222);
nand NAND4 (N7513, N7506, N4900, N4055, N6768);
or OR4 (N7514, N7513, N6259, N4064, N1088);
and AND2 (N7515, N7497, N1438);
not NOT1 (N7516, N7514);
or OR3 (N7517, N7509, N6282, N1859);
and AND3 (N7518, N7510, N6305, N6763);
xor XOR2 (N7519, N7500, N3594);
nor NOR4 (N7520, N7508, N686, N6354, N2374);
not NOT1 (N7521, N7507);
xor XOR2 (N7522, N7520, N7332);
nor NOR4 (N7523, N7521, N6050, N4298, N4256);
xor XOR2 (N7524, N7515, N1456);
nor NOR3 (N7525, N7516, N2536, N6645);
nand NAND2 (N7526, N7522, N7002);
and AND2 (N7527, N7524, N6068);
or OR3 (N7528, N7527, N3461, N4261);
or OR2 (N7529, N7511, N2987);
not NOT1 (N7530, N7517);
buf BUF1 (N7531, N7529);
nor NOR2 (N7532, N7530, N1225);
and AND4 (N7533, N7489, N1580, N5244, N7357);
not NOT1 (N7534, N7523);
nor NOR2 (N7535, N7533, N2443);
xor XOR2 (N7536, N7528, N2875);
and AND2 (N7537, N7518, N3550);
buf BUF1 (N7538, N7535);
buf BUF1 (N7539, N7536);
nand NAND4 (N7540, N7532, N3951, N3016, N2557);
xor XOR2 (N7541, N7537, N4540);
not NOT1 (N7542, N7525);
and AND3 (N7543, N7526, N2130, N585);
buf BUF1 (N7544, N7542);
nor NOR3 (N7545, N7543, N4641, N2396);
nor NOR4 (N7546, N7534, N2931, N2843, N6581);
xor XOR2 (N7547, N7544, N4189);
or OR3 (N7548, N7531, N4670, N2002);
nor NOR3 (N7549, N7545, N4718, N636);
nor NOR2 (N7550, N7546, N2732);
and AND3 (N7551, N7547, N1104, N5432);
nand NAND3 (N7552, N7519, N3522, N2544);
not NOT1 (N7553, N7548);
or OR2 (N7554, N7549, N4694);
nand NAND2 (N7555, N7554, N1178);
and AND4 (N7556, N7540, N120, N5364, N4252);
and AND4 (N7557, N7553, N5810, N2688, N1719);
nor NOR3 (N7558, N7538, N6337, N3606);
or OR3 (N7559, N7550, N3695, N1106);
or OR4 (N7560, N7556, N6208, N449, N4107);
or OR2 (N7561, N7551, N5801);
nor NOR2 (N7562, N7557, N3519);
and AND3 (N7563, N7541, N739, N2949);
xor XOR2 (N7564, N7512, N2368);
nor NOR4 (N7565, N7561, N2930, N6457, N1681);
nor NOR4 (N7566, N7552, N3404, N6958, N1464);
nand NAND2 (N7567, N7566, N4508);
nor NOR2 (N7568, N7563, N1513);
buf BUF1 (N7569, N7568);
buf BUF1 (N7570, N7539);
not NOT1 (N7571, N7555);
nand NAND4 (N7572, N7559, N5357, N5076, N3244);
nand NAND3 (N7573, N7570, N6397, N2068);
and AND3 (N7574, N7571, N3371, N1670);
and AND4 (N7575, N7573, N850, N3856, N4364);
and AND3 (N7576, N7575, N5874, N7327);
xor XOR2 (N7577, N7560, N751);
nand NAND4 (N7578, N7572, N7290, N1120, N1759);
and AND2 (N7579, N7558, N561);
and AND2 (N7580, N7567, N583);
and AND2 (N7581, N7562, N6389);
xor XOR2 (N7582, N7579, N4370);
and AND3 (N7583, N7565, N4236, N6737);
nand NAND3 (N7584, N7564, N2697, N1362);
nor NOR4 (N7585, N7574, N5004, N6502, N5660);
or OR2 (N7586, N7569, N4694);
nor NOR3 (N7587, N7582, N6746, N7539);
or OR3 (N7588, N7586, N5796, N3262);
not NOT1 (N7589, N7581);
and AND2 (N7590, N7589, N3064);
xor XOR2 (N7591, N7580, N5662);
or OR4 (N7592, N7583, N5749, N86, N875);
or OR2 (N7593, N7592, N114);
nand NAND4 (N7594, N7577, N6573, N2475, N5326);
nand NAND4 (N7595, N7578, N4343, N7294, N6374);
and AND4 (N7596, N7590, N2059, N7324, N2851);
not NOT1 (N7597, N7596);
nand NAND3 (N7598, N7597, N4510, N665);
nor NOR3 (N7599, N7593, N3840, N5457);
or OR2 (N7600, N7587, N5802);
buf BUF1 (N7601, N7584);
not NOT1 (N7602, N7585);
nor NOR3 (N7603, N7598, N474, N6392);
and AND3 (N7604, N7594, N6119, N2647);
not NOT1 (N7605, N7600);
nor NOR3 (N7606, N7603, N6920, N3909);
buf BUF1 (N7607, N7591);
xor XOR2 (N7608, N7607, N4965);
and AND2 (N7609, N7604, N6787);
not NOT1 (N7610, N7605);
nor NOR4 (N7611, N7606, N6413, N4289, N6395);
nand NAND4 (N7612, N7602, N7588, N500, N1891);
xor XOR2 (N7613, N4399, N6049);
xor XOR2 (N7614, N7576, N1855);
nand NAND3 (N7615, N7599, N3844, N5534);
buf BUF1 (N7616, N7614);
nor NOR2 (N7617, N7609, N4721);
xor XOR2 (N7618, N7612, N6252);
or OR3 (N7619, N7618, N1138, N1199);
nand NAND3 (N7620, N7611, N3255, N2142);
or OR4 (N7621, N7615, N4459, N1445, N6791);
nor NOR2 (N7622, N7595, N4706);
buf BUF1 (N7623, N7601);
buf BUF1 (N7624, N7610);
nand NAND2 (N7625, N7608, N2168);
or OR2 (N7626, N7621, N4894);
or OR3 (N7627, N7620, N3462, N538);
buf BUF1 (N7628, N7623);
nor NOR4 (N7629, N7626, N3544, N1793, N2596);
and AND2 (N7630, N7625, N3999);
or OR2 (N7631, N7630, N139);
or OR4 (N7632, N7631, N2456, N3034, N1660);
nand NAND4 (N7633, N7624, N6138, N7566, N2914);
xor XOR2 (N7634, N7632, N4405);
or OR2 (N7635, N7628, N6043);
or OR4 (N7636, N7616, N7331, N6167, N3853);
and AND3 (N7637, N7634, N4838, N4760);
xor XOR2 (N7638, N7637, N3310);
nand NAND4 (N7639, N7638, N4912, N1872, N3077);
xor XOR2 (N7640, N7633, N5636);
nand NAND3 (N7641, N7636, N2839, N1040);
or OR3 (N7642, N7640, N3695, N734);
and AND2 (N7643, N7641, N32);
not NOT1 (N7644, N7635);
not NOT1 (N7645, N7639);
or OR3 (N7646, N7619, N7351, N6464);
nand NAND3 (N7647, N7646, N7094, N5798);
nand NAND3 (N7648, N7627, N3163, N1341);
not NOT1 (N7649, N7642);
buf BUF1 (N7650, N7648);
or OR4 (N7651, N7645, N3221, N1227, N2168);
nor NOR3 (N7652, N7629, N1300, N1902);
nand NAND3 (N7653, N7652, N2676, N1510);
or OR2 (N7654, N7651, N4782);
or OR2 (N7655, N7622, N4113);
and AND3 (N7656, N7644, N6072, N1374);
buf BUF1 (N7657, N7647);
not NOT1 (N7658, N7653);
and AND4 (N7659, N7654, N1737, N554, N189);
nand NAND2 (N7660, N7643, N4435);
and AND3 (N7661, N7659, N914, N7110);
nand NAND2 (N7662, N7617, N659);
xor XOR2 (N7663, N7662, N3795);
and AND4 (N7664, N7650, N4006, N759, N5841);
and AND3 (N7665, N7664, N5918, N2879);
nand NAND3 (N7666, N7655, N7009, N830);
and AND3 (N7667, N7665, N1090, N4146);
buf BUF1 (N7668, N7657);
or OR3 (N7669, N7661, N5725, N1955);
not NOT1 (N7670, N7668);
or OR2 (N7671, N7666, N3493);
and AND4 (N7672, N7667, N1998, N1074, N3161);
and AND3 (N7673, N7670, N6046, N1696);
buf BUF1 (N7674, N7663);
xor XOR2 (N7675, N7649, N3335);
and AND4 (N7676, N7658, N4387, N2261, N3194);
nor NOR3 (N7677, N7674, N215, N6176);
and AND4 (N7678, N7660, N1644, N1267, N6404);
or OR4 (N7679, N7672, N7467, N1828, N819);
and AND3 (N7680, N7671, N807, N4681);
and AND2 (N7681, N7673, N2381);
buf BUF1 (N7682, N7680);
not NOT1 (N7683, N7678);
or OR3 (N7684, N7676, N4150, N665);
or OR2 (N7685, N7679, N42);
and AND3 (N7686, N7684, N4998, N2021);
buf BUF1 (N7687, N7669);
nor NOR2 (N7688, N7681, N3121);
xor XOR2 (N7689, N7613, N2623);
xor XOR2 (N7690, N7675, N5905);
and AND4 (N7691, N7677, N7660, N743, N3084);
nor NOR3 (N7692, N7688, N2961, N3345);
buf BUF1 (N7693, N7686);
and AND2 (N7694, N7693, N2591);
buf BUF1 (N7695, N7689);
xor XOR2 (N7696, N7692, N1551);
nor NOR4 (N7697, N7695, N5505, N3766, N5241);
nand NAND3 (N7698, N7687, N6294, N2999);
nor NOR3 (N7699, N7696, N7412, N5825);
not NOT1 (N7700, N7683);
nand NAND4 (N7701, N7691, N3568, N3104, N404);
and AND4 (N7702, N7700, N6772, N2034, N7066);
nand NAND2 (N7703, N7685, N1036);
buf BUF1 (N7704, N7697);
nand NAND3 (N7705, N7690, N4027, N4063);
or OR2 (N7706, N7682, N5527);
not NOT1 (N7707, N7704);
xor XOR2 (N7708, N7698, N3406);
nor NOR3 (N7709, N7706, N1103, N1026);
buf BUF1 (N7710, N7656);
or OR2 (N7711, N7701, N7442);
nand NAND3 (N7712, N7707, N7101, N1469);
nor NOR2 (N7713, N7699, N5229);
buf BUF1 (N7714, N7710);
xor XOR2 (N7715, N7713, N1835);
and AND4 (N7716, N7694, N2353, N3722, N3121);
not NOT1 (N7717, N7711);
nand NAND2 (N7718, N7717, N3589);
nand NAND4 (N7719, N7718, N3284, N5587, N1135);
nor NOR4 (N7720, N7709, N813, N6887, N3009);
not NOT1 (N7721, N7705);
nor NOR3 (N7722, N7702, N4413, N1681);
and AND3 (N7723, N7719, N628, N5153);
not NOT1 (N7724, N7722);
or OR2 (N7725, N7715, N7163);
buf BUF1 (N7726, N7725);
nand NAND2 (N7727, N7708, N5222);
nor NOR2 (N7728, N7716, N7702);
buf BUF1 (N7729, N7727);
nor NOR4 (N7730, N7729, N2486, N3511, N5719);
not NOT1 (N7731, N7721);
buf BUF1 (N7732, N7730);
buf BUF1 (N7733, N7703);
not NOT1 (N7734, N7724);
buf BUF1 (N7735, N7723);
not NOT1 (N7736, N7735);
nand NAND2 (N7737, N7726, N4697);
xor XOR2 (N7738, N7733, N2473);
and AND3 (N7739, N7714, N2102, N3487);
or OR3 (N7740, N7734, N6185, N7275);
or OR4 (N7741, N7738, N6097, N7178, N5422);
nand NAND4 (N7742, N7739, N3911, N5712, N3580);
xor XOR2 (N7743, N7736, N1300);
or OR2 (N7744, N7741, N4701);
buf BUF1 (N7745, N7720);
nor NOR3 (N7746, N7740, N7271, N3853);
nor NOR3 (N7747, N7737, N6307, N5933);
xor XOR2 (N7748, N7742, N7593);
not NOT1 (N7749, N7728);
nor NOR3 (N7750, N7743, N6725, N6964);
or OR3 (N7751, N7749, N5835, N2303);
not NOT1 (N7752, N7731);
xor XOR2 (N7753, N7712, N3264);
or OR2 (N7754, N7751, N1976);
or OR4 (N7755, N7744, N1524, N4182, N2096);
nor NOR3 (N7756, N7748, N2648, N3779);
or OR4 (N7757, N7753, N800, N4701, N554);
buf BUF1 (N7758, N7747);
xor XOR2 (N7759, N7750, N3149);
nand NAND3 (N7760, N7746, N903, N4429);
buf BUF1 (N7761, N7754);
buf BUF1 (N7762, N7732);
buf BUF1 (N7763, N7756);
xor XOR2 (N7764, N7759, N7332);
nand NAND2 (N7765, N7758, N667);
or OR2 (N7766, N7755, N331);
not NOT1 (N7767, N7766);
and AND4 (N7768, N7763, N1755, N5160, N332);
buf BUF1 (N7769, N7757);
xor XOR2 (N7770, N7760, N1779);
not NOT1 (N7771, N7761);
not NOT1 (N7772, N7768);
and AND2 (N7773, N7752, N2170);
not NOT1 (N7774, N7770);
xor XOR2 (N7775, N7765, N7130);
nand NAND4 (N7776, N7774, N5702, N4486, N7713);
not NOT1 (N7777, N7776);
nand NAND3 (N7778, N7762, N5680, N7112);
xor XOR2 (N7779, N7767, N6172);
nand NAND3 (N7780, N7772, N5175, N150);
or OR2 (N7781, N7771, N3645);
buf BUF1 (N7782, N7775);
buf BUF1 (N7783, N7764);
xor XOR2 (N7784, N7777, N5574);
nand NAND4 (N7785, N7782, N315, N1203, N6018);
buf BUF1 (N7786, N7785);
nand NAND4 (N7787, N7779, N5036, N2561, N4730);
xor XOR2 (N7788, N7745, N6758);
or OR3 (N7789, N7784, N5798, N3884);
not NOT1 (N7790, N7786);
and AND2 (N7791, N7769, N1205);
nand NAND2 (N7792, N7789, N2278);
not NOT1 (N7793, N7792);
nand NAND2 (N7794, N7790, N6546);
xor XOR2 (N7795, N7781, N365);
nand NAND4 (N7796, N7778, N6675, N59, N3366);
buf BUF1 (N7797, N7795);
nor NOR2 (N7798, N7783, N1616);
buf BUF1 (N7799, N7787);
buf BUF1 (N7800, N7773);
xor XOR2 (N7801, N7797, N5589);
nor NOR3 (N7802, N7780, N5855, N2510);
nor NOR3 (N7803, N7799, N6252, N3124);
nand NAND2 (N7804, N7794, N1261);
or OR2 (N7805, N7802, N5019);
and AND3 (N7806, N7796, N4512, N7313);
buf BUF1 (N7807, N7798);
buf BUF1 (N7808, N7791);
and AND3 (N7809, N7806, N6380, N6406);
nor NOR2 (N7810, N7809, N648);
or OR2 (N7811, N7808, N4589);
buf BUF1 (N7812, N7810);
not NOT1 (N7813, N7793);
and AND3 (N7814, N7788, N2620, N1436);
nor NOR4 (N7815, N7800, N2784, N3193, N1342);
nand NAND4 (N7816, N7815, N2582, N5742, N2473);
xor XOR2 (N7817, N7814, N6110);
nor NOR2 (N7818, N7804, N6780);
or OR3 (N7819, N7807, N6935, N67);
buf BUF1 (N7820, N7817);
buf BUF1 (N7821, N7811);
or OR2 (N7822, N7803, N5087);
and AND3 (N7823, N7822, N4029, N2925);
nor NOR4 (N7824, N7813, N2547, N1518, N4433);
nand NAND2 (N7825, N7819, N576);
xor XOR2 (N7826, N7825, N948);
and AND2 (N7827, N7818, N2904);
nand NAND2 (N7828, N7816, N7602);
and AND2 (N7829, N7821, N3096);
nand NAND2 (N7830, N7829, N7141);
nand NAND2 (N7831, N7828, N5390);
not NOT1 (N7832, N7805);
buf BUF1 (N7833, N7820);
not NOT1 (N7834, N7833);
nand NAND3 (N7835, N7830, N1828, N5066);
not NOT1 (N7836, N7831);
not NOT1 (N7837, N7823);
and AND4 (N7838, N7824, N5310, N2226, N1070);
buf BUF1 (N7839, N7801);
and AND2 (N7840, N7834, N6013);
buf BUF1 (N7841, N7838);
nor NOR2 (N7842, N7837, N2932);
nor NOR2 (N7843, N7832, N7612);
and AND2 (N7844, N7835, N4925);
buf BUF1 (N7845, N7812);
and AND3 (N7846, N7839, N3063, N1283);
nand NAND3 (N7847, N7846, N4924, N3264);
and AND2 (N7848, N7841, N1944);
not NOT1 (N7849, N7842);
xor XOR2 (N7850, N7849, N3340);
not NOT1 (N7851, N7845);
buf BUF1 (N7852, N7827);
and AND3 (N7853, N7852, N742, N89);
nand NAND2 (N7854, N7844, N3374);
and AND4 (N7855, N7843, N4578, N6869, N3681);
buf BUF1 (N7856, N7826);
buf BUF1 (N7857, N7854);
not NOT1 (N7858, N7857);
not NOT1 (N7859, N7856);
nand NAND2 (N7860, N7859, N4232);
nand NAND4 (N7861, N7847, N3224, N3509, N7307);
or OR4 (N7862, N7858, N3208, N30, N2759);
or OR4 (N7863, N7850, N5808, N5324, N3191);
xor XOR2 (N7864, N7855, N2616);
not NOT1 (N7865, N7860);
nor NOR2 (N7866, N7836, N5428);
nand NAND2 (N7867, N7851, N3300);
nand NAND2 (N7868, N7861, N1089);
or OR4 (N7869, N7862, N897, N5869, N893);
or OR4 (N7870, N7868, N2569, N3668, N2831);
or OR2 (N7871, N7869, N2547);
xor XOR2 (N7872, N7848, N1244);
buf BUF1 (N7873, N7866);
and AND2 (N7874, N7873, N2997);
nor NOR4 (N7875, N7871, N1566, N5989, N2266);
not NOT1 (N7876, N7853);
buf BUF1 (N7877, N7863);
and AND3 (N7878, N7874, N6084, N3748);
or OR4 (N7879, N7867, N3107, N159, N6319);
nor NOR4 (N7880, N7872, N3597, N7756, N2649);
xor XOR2 (N7881, N7877, N5544);
or OR3 (N7882, N7840, N901, N1072);
nand NAND4 (N7883, N7865, N6011, N7320, N3837);
buf BUF1 (N7884, N7864);
or OR2 (N7885, N7883, N7634);
or OR3 (N7886, N7880, N6073, N4432);
not NOT1 (N7887, N7882);
xor XOR2 (N7888, N7870, N7693);
buf BUF1 (N7889, N7886);
not NOT1 (N7890, N7878);
nand NAND2 (N7891, N7875, N4341);
and AND2 (N7892, N7881, N7434);
or OR2 (N7893, N7888, N729);
or OR2 (N7894, N7876, N4388);
nor NOR2 (N7895, N7887, N902);
nand NAND2 (N7896, N7893, N5659);
or OR3 (N7897, N7885, N5515, N2188);
buf BUF1 (N7898, N7890);
xor XOR2 (N7899, N7891, N6683);
not NOT1 (N7900, N7897);
xor XOR2 (N7901, N7884, N1901);
nand NAND2 (N7902, N7900, N2507);
buf BUF1 (N7903, N7892);
and AND2 (N7904, N7889, N6318);
not NOT1 (N7905, N7879);
or OR3 (N7906, N7898, N3474, N1214);
and AND4 (N7907, N7899, N4077, N442, N6303);
nand NAND2 (N7908, N7901, N5058);
not NOT1 (N7909, N7905);
nor NOR4 (N7910, N7902, N4013, N6389, N1371);
nor NOR4 (N7911, N7896, N2974, N177, N1464);
and AND4 (N7912, N7904, N7682, N7409, N7178);
not NOT1 (N7913, N7903);
nor NOR4 (N7914, N7911, N165, N3003, N578);
xor XOR2 (N7915, N7909, N6248);
xor XOR2 (N7916, N7906, N1224);
buf BUF1 (N7917, N7916);
not NOT1 (N7918, N7915);
buf BUF1 (N7919, N7912);
xor XOR2 (N7920, N7894, N1309);
or OR4 (N7921, N7919, N4541, N4743, N4970);
buf BUF1 (N7922, N7913);
and AND2 (N7923, N7918, N2529);
nor NOR2 (N7924, N7920, N7205);
nand NAND3 (N7925, N7908, N5053, N3854);
nand NAND2 (N7926, N7921, N320);
not NOT1 (N7927, N7923);
not NOT1 (N7928, N7895);
not NOT1 (N7929, N7910);
buf BUF1 (N7930, N7907);
not NOT1 (N7931, N7927);
and AND4 (N7932, N7930, N1907, N7310, N5810);
or OR4 (N7933, N7917, N7203, N329, N6402);
and AND4 (N7934, N7926, N2234, N904, N1647);
not NOT1 (N7935, N7933);
nor NOR4 (N7936, N7924, N5180, N6222, N548);
and AND2 (N7937, N7929, N5801);
nand NAND3 (N7938, N7932, N2331, N514);
xor XOR2 (N7939, N7934, N7885);
buf BUF1 (N7940, N7935);
not NOT1 (N7941, N7928);
or OR2 (N7942, N7925, N1451);
nor NOR2 (N7943, N7938, N6565);
buf BUF1 (N7944, N7941);
not NOT1 (N7945, N7943);
nand NAND2 (N7946, N7945, N3458);
nor NOR3 (N7947, N7939, N2754, N3365);
nor NOR4 (N7948, N7940, N6782, N3756, N869);
or OR4 (N7949, N7944, N4213, N1909, N3797);
nand NAND2 (N7950, N7937, N4171);
xor XOR2 (N7951, N7948, N6686);
or OR3 (N7952, N7946, N7948, N2245);
and AND3 (N7953, N7942, N4937, N7605);
buf BUF1 (N7954, N7950);
and AND4 (N7955, N7947, N3652, N4019, N1919);
buf BUF1 (N7956, N7931);
buf BUF1 (N7957, N7952);
xor XOR2 (N7958, N7949, N3745);
nand NAND2 (N7959, N7954, N2564);
not NOT1 (N7960, N7914);
or OR4 (N7961, N7960, N7105, N5739, N866);
not NOT1 (N7962, N7922);
nand NAND3 (N7963, N7951, N7532, N7724);
xor XOR2 (N7964, N7961, N2556);
nand NAND2 (N7965, N7963, N7518);
nor NOR4 (N7966, N7958, N7690, N506, N4290);
not NOT1 (N7967, N7959);
and AND4 (N7968, N7955, N52, N4546, N1407);
xor XOR2 (N7969, N7956, N3497);
xor XOR2 (N7970, N7965, N4613);
and AND2 (N7971, N7936, N2460);
not NOT1 (N7972, N7969);
not NOT1 (N7973, N7966);
and AND4 (N7974, N7973, N1627, N509, N5035);
nand NAND4 (N7975, N7970, N3334, N2707, N1604);
or OR2 (N7976, N7972, N2592);
nor NOR2 (N7977, N7976, N2124);
or OR2 (N7978, N7962, N15);
or OR2 (N7979, N7975, N523);
nand NAND4 (N7980, N7971, N2201, N7956, N5175);
nor NOR4 (N7981, N7967, N7551, N3871, N6384);
or OR3 (N7982, N7957, N1290, N6751);
nor NOR3 (N7983, N7953, N167, N6785);
buf BUF1 (N7984, N7978);
and AND4 (N7985, N7981, N6262, N6559, N5153);
nor NOR4 (N7986, N7980, N6121, N3653, N5);
or OR4 (N7987, N7974, N3894, N5824, N7355);
buf BUF1 (N7988, N7983);
not NOT1 (N7989, N7982);
or OR4 (N7990, N7986, N2372, N4320, N4026);
xor XOR2 (N7991, N7987, N846);
nand NAND4 (N7992, N7984, N5391, N303, N7198);
and AND3 (N7993, N7968, N4598, N3411);
nand NAND2 (N7994, N7979, N4357);
and AND2 (N7995, N7964, N568);
not NOT1 (N7996, N7992);
and AND4 (N7997, N7988, N4, N6469, N7931);
and AND3 (N7998, N7997, N7747, N668);
or OR4 (N7999, N7996, N2102, N6226, N5506);
xor XOR2 (N8000, N7977, N100);
buf BUF1 (N8001, N7994);
nand NAND4 (N8002, N7989, N6377, N878, N7243);
and AND2 (N8003, N7985, N411);
or OR3 (N8004, N7999, N4460, N7312);
not NOT1 (N8005, N7990);
and AND2 (N8006, N8005, N7040);
and AND4 (N8007, N8006, N7225, N1226, N7143);
or OR3 (N8008, N7991, N646, N6931);
buf BUF1 (N8009, N7993);
nand NAND2 (N8010, N8000, N1738);
not NOT1 (N8011, N8004);
xor XOR2 (N8012, N8009, N2083);
xor XOR2 (N8013, N8001, N4734);
not NOT1 (N8014, N8008);
not NOT1 (N8015, N8002);
nand NAND2 (N8016, N7995, N7373);
buf BUF1 (N8017, N8015);
endmodule