// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19;

output N8010,N8013,N8017,N7999,N8014,N7987,N8008,N8018,N8016,N8019;

nor NOR4 (N20, N17, N5, N1, N12);
not NOT1 (N21, N11);
and AND2 (N22, N14, N11);
and AND3 (N23, N12, N8, N3);
nor NOR4 (N24, N7, N2, N4, N23);
nand NAND3 (N25, N4, N23, N16);
nor NOR4 (N26, N8, N20, N23, N4);
buf BUF1 (N27, N20);
and AND3 (N28, N18, N8, N19);
nor NOR3 (N29, N26, N22, N18);
nand NAND3 (N30, N26, N29, N8);
or OR2 (N31, N25, N15);
buf BUF1 (N32, N27);
buf BUF1 (N33, N4);
and AND2 (N34, N20, N7);
nor NOR2 (N35, N26, N31);
nand NAND3 (N36, N25, N16, N6);
xor XOR2 (N37, N8, N28);
or OR3 (N38, N4, N7, N14);
buf BUF1 (N39, N36);
nor NOR3 (N40, N32, N26, N30);
not NOT1 (N41, N39);
nor NOR4 (N42, N30, N25, N18, N5);
xor XOR2 (N43, N35, N25);
nor NOR4 (N44, N34, N33, N6, N17);
buf BUF1 (N45, N35);
nor NOR2 (N46, N40, N34);
xor XOR2 (N47, N46, N2);
buf BUF1 (N48, N44);
buf BUF1 (N49, N38);
nor NOR3 (N50, N37, N29, N49);
not NOT1 (N51, N31);
buf BUF1 (N52, N42);
and AND3 (N53, N50, N44, N25);
and AND4 (N54, N21, N48, N14, N30);
nor NOR3 (N55, N53, N5, N6);
buf BUF1 (N56, N52);
or OR4 (N57, N50, N5, N18, N8);
buf BUF1 (N58, N55);
xor XOR2 (N59, N45, N12);
not NOT1 (N60, N59);
xor XOR2 (N61, N56, N26);
xor XOR2 (N62, N43, N2);
and AND3 (N63, N24, N29, N44);
or OR4 (N64, N60, N22, N24, N18);
buf BUF1 (N65, N57);
nor NOR4 (N66, N62, N29, N21, N54);
not NOT1 (N67, N2);
buf BUF1 (N68, N61);
xor XOR2 (N69, N63, N26);
nand NAND2 (N70, N58, N26);
nor NOR4 (N71, N67, N28, N37, N53);
nand NAND2 (N72, N66, N67);
buf BUF1 (N73, N68);
buf BUF1 (N74, N72);
or OR3 (N75, N47, N20, N47);
nor NOR3 (N76, N71, N66, N5);
nand NAND3 (N77, N76, N58, N32);
not NOT1 (N78, N64);
nand NAND3 (N79, N51, N78, N31);
xor XOR2 (N80, N75, N22);
nand NAND2 (N81, N3, N41);
nand NAND3 (N82, N43, N47, N48);
xor XOR2 (N83, N65, N32);
or OR4 (N84, N79, N14, N77, N48);
nand NAND4 (N85, N42, N80, N81, N55);
or OR3 (N86, N84, N10, N9);
xor XOR2 (N87, N52, N52);
or OR3 (N88, N4, N64, N25);
xor XOR2 (N89, N85, N54);
buf BUF1 (N90, N74);
xor XOR2 (N91, N83, N80);
buf BUF1 (N92, N73);
nor NOR2 (N93, N88, N9);
and AND3 (N94, N93, N69, N86);
not NOT1 (N95, N21);
not NOT1 (N96, N64);
nand NAND4 (N97, N96, N15, N10, N47);
nand NAND2 (N98, N89, N24);
xor XOR2 (N99, N98, N37);
or OR2 (N100, N95, N74);
or OR3 (N101, N90, N71, N34);
nor NOR4 (N102, N94, N39, N45, N75);
nor NOR2 (N103, N97, N92);
nand NAND3 (N104, N44, N35, N99);
nor NOR3 (N105, N22, N11, N83);
buf BUF1 (N106, N104);
buf BUF1 (N107, N106);
not NOT1 (N108, N107);
not NOT1 (N109, N108);
buf BUF1 (N110, N105);
nor NOR4 (N111, N101, N96, N61, N25);
or OR2 (N112, N70, N101);
nand NAND2 (N113, N82, N64);
nand NAND4 (N114, N87, N75, N16, N79);
nand NAND4 (N115, N111, N2, N62, N13);
or OR2 (N116, N109, N16);
buf BUF1 (N117, N102);
or OR3 (N118, N117, N28, N106);
nor NOR4 (N119, N116, N106, N87, N5);
not NOT1 (N120, N103);
buf BUF1 (N121, N100);
buf BUF1 (N122, N113);
buf BUF1 (N123, N120);
not NOT1 (N124, N112);
xor XOR2 (N125, N124, N92);
or OR3 (N126, N110, N119, N119);
not NOT1 (N127, N112);
nor NOR3 (N128, N125, N15, N72);
buf BUF1 (N129, N121);
or OR2 (N130, N126, N4);
nand NAND2 (N131, N129, N54);
xor XOR2 (N132, N130, N113);
nor NOR4 (N133, N91, N45, N30, N129);
or OR4 (N134, N127, N69, N109, N89);
or OR3 (N135, N133, N115, N105);
or OR4 (N136, N50, N10, N37, N100);
buf BUF1 (N137, N123);
buf BUF1 (N138, N131);
or OR3 (N139, N136, N84, N29);
or OR4 (N140, N135, N126, N130, N29);
not NOT1 (N141, N134);
nor NOR3 (N142, N140, N137, N79);
or OR3 (N143, N98, N17, N131);
or OR4 (N144, N132, N117, N42, N15);
and AND3 (N145, N144, N25, N67);
buf BUF1 (N146, N141);
or OR4 (N147, N114, N123, N50, N65);
buf BUF1 (N148, N139);
not NOT1 (N149, N147);
xor XOR2 (N150, N143, N112);
buf BUF1 (N151, N128);
not NOT1 (N152, N122);
not NOT1 (N153, N142);
and AND4 (N154, N153, N128, N44, N61);
or OR3 (N155, N118, N54, N33);
nand NAND3 (N156, N151, N116, N102);
nor NOR3 (N157, N156, N58, N51);
or OR4 (N158, N157, N130, N45, N87);
xor XOR2 (N159, N154, N92);
or OR4 (N160, N150, N44, N17, N11);
xor XOR2 (N161, N155, N97);
or OR2 (N162, N146, N77);
buf BUF1 (N163, N162);
nand NAND3 (N164, N152, N88, N125);
not NOT1 (N165, N148);
nor NOR2 (N166, N163, N162);
buf BUF1 (N167, N164);
xor XOR2 (N168, N145, N100);
or OR2 (N169, N159, N127);
nor NOR3 (N170, N168, N38, N14);
buf BUF1 (N171, N138);
buf BUF1 (N172, N170);
xor XOR2 (N173, N169, N26);
or OR3 (N174, N172, N25, N7);
and AND2 (N175, N166, N132);
or OR2 (N176, N167, N133);
xor XOR2 (N177, N165, N78);
or OR2 (N178, N161, N164);
nor NOR4 (N179, N178, N21, N65, N111);
nand NAND4 (N180, N177, N167, N47, N112);
nand NAND2 (N181, N149, N104);
or OR2 (N182, N179, N168);
or OR3 (N183, N171, N141, N10);
xor XOR2 (N184, N174, N25);
nor NOR2 (N185, N181, N160);
and AND2 (N186, N51, N92);
xor XOR2 (N187, N185, N100);
nor NOR2 (N188, N173, N139);
and AND4 (N189, N188, N76, N120, N133);
or OR2 (N190, N186, N29);
and AND4 (N191, N184, N64, N134, N154);
or OR3 (N192, N175, N19, N93);
not NOT1 (N193, N158);
xor XOR2 (N194, N190, N99);
xor XOR2 (N195, N192, N58);
not NOT1 (N196, N191);
nand NAND4 (N197, N189, N189, N148, N149);
or OR3 (N198, N197, N8, N38);
nand NAND3 (N199, N182, N107, N4);
or OR3 (N200, N194, N88, N94);
buf BUF1 (N201, N176);
buf BUF1 (N202, N200);
buf BUF1 (N203, N196);
and AND2 (N204, N203, N136);
not NOT1 (N205, N180);
and AND2 (N206, N183, N19);
or OR3 (N207, N206, N60, N48);
nand NAND3 (N208, N205, N170, N22);
xor XOR2 (N209, N207, N175);
nand NAND4 (N210, N209, N123, N145, N75);
buf BUF1 (N211, N202);
and AND2 (N212, N208, N105);
not NOT1 (N213, N195);
nor NOR3 (N214, N199, N115, N125);
or OR4 (N215, N193, N214, N53, N209);
nor NOR3 (N216, N121, N165, N177);
nor NOR4 (N217, N216, N137, N105, N121);
nor NOR4 (N218, N212, N92, N140, N62);
xor XOR2 (N219, N218, N93);
not NOT1 (N220, N219);
xor XOR2 (N221, N211, N200);
or OR3 (N222, N198, N93, N151);
nor NOR3 (N223, N217, N200, N31);
and AND4 (N224, N221, N32, N66, N207);
nor NOR3 (N225, N201, N49, N186);
not NOT1 (N226, N220);
buf BUF1 (N227, N224);
buf BUF1 (N228, N226);
nand NAND3 (N229, N210, N184, N101);
xor XOR2 (N230, N223, N71);
xor XOR2 (N231, N222, N92);
xor XOR2 (N232, N231, N218);
or OR3 (N233, N213, N29, N24);
nor NOR4 (N234, N229, N57, N159, N73);
xor XOR2 (N235, N228, N71);
nand NAND2 (N236, N227, N155);
nor NOR4 (N237, N235, N167, N77, N195);
nor NOR2 (N238, N233, N94);
not NOT1 (N239, N230);
nor NOR2 (N240, N225, N108);
buf BUF1 (N241, N238);
nand NAND3 (N242, N215, N59, N28);
xor XOR2 (N243, N239, N115);
and AND3 (N244, N237, N235, N126);
and AND2 (N245, N241, N73);
not NOT1 (N246, N240);
and AND4 (N247, N234, N185, N208, N181);
buf BUF1 (N248, N232);
nor NOR4 (N249, N187, N205, N113, N165);
nand NAND2 (N250, N245, N91);
nand NAND4 (N251, N242, N66, N8, N11);
and AND4 (N252, N246, N9, N126, N184);
nor NOR2 (N253, N236, N97);
not NOT1 (N254, N248);
or OR2 (N255, N204, N225);
nand NAND2 (N256, N244, N209);
xor XOR2 (N257, N243, N112);
nor NOR4 (N258, N250, N128, N39, N38);
not NOT1 (N259, N249);
nor NOR2 (N260, N254, N97);
nor NOR3 (N261, N247, N221, N257);
nand NAND3 (N262, N84, N29, N261);
or OR3 (N263, N89, N153, N166);
xor XOR2 (N264, N262, N69);
not NOT1 (N265, N258);
or OR2 (N266, N255, N134);
or OR3 (N267, N256, N105, N143);
buf BUF1 (N268, N251);
and AND2 (N269, N267, N153);
nand NAND3 (N270, N268, N81, N130);
nor NOR3 (N271, N253, N66, N123);
nor NOR3 (N272, N271, N226, N224);
or OR4 (N273, N272, N105, N230, N229);
not NOT1 (N274, N259);
nor NOR4 (N275, N260, N60, N166, N59);
or OR4 (N276, N264, N151, N181, N193);
nor NOR4 (N277, N269, N19, N131, N164);
and AND2 (N278, N273, N215);
not NOT1 (N279, N278);
or OR3 (N280, N263, N189, N7);
or OR2 (N281, N279, N251);
buf BUF1 (N282, N277);
and AND3 (N283, N280, N1, N165);
or OR3 (N284, N275, N85, N229);
buf BUF1 (N285, N281);
and AND3 (N286, N265, N170, N107);
nand NAND2 (N287, N284, N245);
nand NAND2 (N288, N252, N249);
nor NOR3 (N289, N274, N214, N77);
not NOT1 (N290, N287);
or OR4 (N291, N276, N179, N155, N205);
or OR4 (N292, N266, N36, N94, N17);
or OR4 (N293, N292, N160, N188, N75);
not NOT1 (N294, N288);
buf BUF1 (N295, N294);
xor XOR2 (N296, N290, N10);
buf BUF1 (N297, N295);
nor NOR4 (N298, N289, N216, N89, N181);
or OR4 (N299, N285, N32, N25, N160);
not NOT1 (N300, N286);
not NOT1 (N301, N296);
and AND4 (N302, N301, N242, N232, N287);
and AND2 (N303, N282, N43);
not NOT1 (N304, N303);
or OR2 (N305, N299, N279);
buf BUF1 (N306, N305);
xor XOR2 (N307, N297, N56);
and AND3 (N308, N304, N141, N203);
xor XOR2 (N309, N308, N211);
buf BUF1 (N310, N302);
xor XOR2 (N311, N309, N55);
nand NAND2 (N312, N311, N28);
nor NOR2 (N313, N270, N231);
and AND3 (N314, N300, N138, N104);
nand NAND4 (N315, N314, N183, N81, N234);
nand NAND4 (N316, N283, N250, N208, N198);
or OR3 (N317, N310, N295, N176);
nand NAND3 (N318, N317, N151, N268);
buf BUF1 (N319, N306);
buf BUF1 (N320, N313);
nor NOR2 (N321, N291, N137);
or OR3 (N322, N298, N119, N258);
not NOT1 (N323, N320);
buf BUF1 (N324, N307);
nor NOR2 (N325, N324, N3);
xor XOR2 (N326, N319, N8);
and AND4 (N327, N325, N102, N285, N31);
nor NOR3 (N328, N327, N11, N312);
buf BUF1 (N329, N185);
nor NOR2 (N330, N293, N178);
buf BUF1 (N331, N316);
nand NAND4 (N332, N329, N238, N124, N166);
or OR2 (N333, N322, N158);
xor XOR2 (N334, N321, N197);
nor NOR3 (N335, N318, N158, N51);
nand NAND2 (N336, N330, N226);
or OR2 (N337, N334, N141);
nand NAND4 (N338, N328, N172, N205, N96);
not NOT1 (N339, N338);
and AND2 (N340, N331, N180);
buf BUF1 (N341, N332);
nor NOR4 (N342, N335, N128, N196, N84);
nand NAND3 (N343, N326, N179, N126);
and AND3 (N344, N340, N218, N245);
or OR4 (N345, N339, N251, N73, N234);
buf BUF1 (N346, N315);
and AND2 (N347, N343, N210);
buf BUF1 (N348, N342);
xor XOR2 (N349, N341, N256);
and AND4 (N350, N336, N305, N163, N149);
nor NOR3 (N351, N337, N221, N152);
nor NOR4 (N352, N351, N216, N23, N5);
and AND3 (N353, N352, N281, N36);
or OR2 (N354, N349, N117);
xor XOR2 (N355, N354, N10);
and AND3 (N356, N344, N81, N278);
and AND2 (N357, N345, N95);
xor XOR2 (N358, N323, N345);
and AND3 (N359, N350, N316, N51);
nor NOR2 (N360, N347, N254);
nand NAND2 (N361, N346, N322);
and AND2 (N362, N353, N228);
not NOT1 (N363, N348);
nand NAND2 (N364, N360, N239);
nor NOR2 (N365, N362, N46);
nor NOR3 (N366, N359, N286, N242);
or OR2 (N367, N364, N250);
or OR2 (N368, N367, N82);
or OR3 (N369, N358, N59, N248);
or OR2 (N370, N361, N366);
and AND2 (N371, N178, N354);
and AND2 (N372, N355, N58);
and AND3 (N373, N333, N304, N295);
nor NOR4 (N374, N373, N148, N326, N153);
nand NAND2 (N375, N374, N360);
nand NAND4 (N376, N365, N240, N90, N203);
not NOT1 (N377, N356);
or OR4 (N378, N377, N171, N8, N338);
or OR2 (N379, N372, N1);
buf BUF1 (N380, N371);
and AND2 (N381, N368, N126);
xor XOR2 (N382, N379, N161);
nor NOR2 (N383, N375, N100);
or OR2 (N384, N369, N298);
nand NAND4 (N385, N381, N268, N139, N380);
nor NOR4 (N386, N374, N204, N45, N144);
buf BUF1 (N387, N363);
or OR4 (N388, N357, N78, N59, N94);
and AND3 (N389, N383, N192, N13);
nor NOR2 (N390, N385, N183);
or OR4 (N391, N370, N288, N58, N338);
and AND2 (N392, N389, N251);
buf BUF1 (N393, N388);
nor NOR4 (N394, N392, N100, N366, N293);
nor NOR4 (N395, N376, N342, N332, N37);
nand NAND3 (N396, N382, N295, N304);
and AND2 (N397, N391, N185);
not NOT1 (N398, N386);
and AND2 (N399, N396, N125);
xor XOR2 (N400, N394, N353);
and AND2 (N401, N387, N276);
and AND4 (N402, N397, N144, N27, N283);
nor NOR2 (N403, N401, N305);
not NOT1 (N404, N399);
nand NAND3 (N405, N384, N306, N281);
buf BUF1 (N406, N400);
buf BUF1 (N407, N406);
xor XOR2 (N408, N390, N117);
nand NAND2 (N409, N395, N134);
buf BUF1 (N410, N408);
not NOT1 (N411, N403);
nand NAND4 (N412, N402, N96, N67, N136);
not NOT1 (N413, N412);
xor XOR2 (N414, N378, N223);
buf BUF1 (N415, N405);
and AND4 (N416, N415, N229, N78, N76);
and AND4 (N417, N411, N375, N120, N63);
nor NOR3 (N418, N410, N189, N173);
buf BUF1 (N419, N414);
buf BUF1 (N420, N419);
xor XOR2 (N421, N407, N232);
not NOT1 (N422, N404);
or OR4 (N423, N418, N184, N190, N386);
buf BUF1 (N424, N409);
buf BUF1 (N425, N421);
nor NOR3 (N426, N420, N100, N193);
or OR3 (N427, N423, N113, N228);
nor NOR2 (N428, N427, N172);
nor NOR2 (N429, N416, N204);
nor NOR2 (N430, N429, N373);
xor XOR2 (N431, N426, N56);
not NOT1 (N432, N422);
or OR4 (N433, N413, N102, N425, N410);
nand NAND3 (N434, N75, N411, N334);
or OR3 (N435, N430, N225, N241);
nor NOR4 (N436, N417, N87, N283, N347);
not NOT1 (N437, N398);
and AND3 (N438, N432, N9, N113);
or OR2 (N439, N437, N219);
nand NAND2 (N440, N393, N318);
xor XOR2 (N441, N424, N278);
and AND2 (N442, N438, N350);
buf BUF1 (N443, N441);
buf BUF1 (N444, N434);
nor NOR2 (N445, N435, N267);
buf BUF1 (N446, N428);
xor XOR2 (N447, N431, N138);
buf BUF1 (N448, N446);
buf BUF1 (N449, N433);
nor NOR3 (N450, N440, N227, N216);
or OR3 (N451, N443, N314, N291);
xor XOR2 (N452, N442, N197);
not NOT1 (N453, N448);
buf BUF1 (N454, N451);
buf BUF1 (N455, N447);
and AND2 (N456, N449, N391);
or OR3 (N457, N454, N368, N35);
nand NAND3 (N458, N445, N80, N352);
not NOT1 (N459, N452);
nor NOR4 (N460, N436, N342, N352, N109);
xor XOR2 (N461, N453, N235);
and AND4 (N462, N455, N333, N316, N284);
or OR2 (N463, N456, N293);
buf BUF1 (N464, N463);
xor XOR2 (N465, N458, N245);
xor XOR2 (N466, N460, N307);
or OR4 (N467, N450, N223, N156, N248);
nand NAND4 (N468, N444, N421, N307, N379);
buf BUF1 (N469, N462);
buf BUF1 (N470, N468);
nand NAND3 (N471, N461, N208, N308);
or OR3 (N472, N471, N24, N362);
or OR3 (N473, N467, N223, N159);
or OR4 (N474, N439, N73, N153, N290);
and AND4 (N475, N473, N357, N13, N232);
xor XOR2 (N476, N475, N249);
nor NOR3 (N477, N464, N196, N428);
not NOT1 (N478, N459);
nor NOR2 (N479, N476, N444);
nor NOR2 (N480, N457, N342);
and AND4 (N481, N469, N79, N51, N29);
xor XOR2 (N482, N477, N240);
or OR3 (N483, N478, N211, N364);
xor XOR2 (N484, N480, N50);
or OR4 (N485, N479, N143, N126, N337);
and AND4 (N486, N482, N338, N422, N92);
not NOT1 (N487, N484);
or OR4 (N488, N472, N387, N245, N375);
xor XOR2 (N489, N474, N176);
buf BUF1 (N490, N489);
nand NAND4 (N491, N483, N380, N50, N291);
not NOT1 (N492, N485);
xor XOR2 (N493, N491, N200);
buf BUF1 (N494, N481);
nand NAND3 (N495, N465, N257, N469);
and AND3 (N496, N466, N253, N212);
nor NOR4 (N497, N488, N144, N114, N246);
nand NAND2 (N498, N494, N57);
buf BUF1 (N499, N492);
and AND2 (N500, N498, N419);
xor XOR2 (N501, N497, N379);
nand NAND4 (N502, N486, N392, N352, N224);
and AND2 (N503, N470, N117);
nand NAND3 (N504, N503, N255, N198);
nand NAND3 (N505, N490, N431, N446);
nand NAND4 (N506, N505, N260, N481, N225);
and AND2 (N507, N487, N157);
not NOT1 (N508, N501);
buf BUF1 (N509, N495);
or OR3 (N510, N506, N72, N339);
or OR4 (N511, N499, N114, N286, N149);
not NOT1 (N512, N496);
buf BUF1 (N513, N493);
buf BUF1 (N514, N511);
or OR4 (N515, N513, N314, N440, N105);
nand NAND2 (N516, N502, N447);
buf BUF1 (N517, N507);
not NOT1 (N518, N508);
xor XOR2 (N519, N500, N437);
xor XOR2 (N520, N516, N278);
and AND4 (N521, N520, N10, N368, N228);
and AND2 (N522, N517, N291);
buf BUF1 (N523, N512);
xor XOR2 (N524, N515, N408);
not NOT1 (N525, N521);
buf BUF1 (N526, N522);
and AND2 (N527, N518, N145);
and AND3 (N528, N526, N453, N419);
nand NAND2 (N529, N514, N363);
not NOT1 (N530, N524);
xor XOR2 (N531, N504, N373);
or OR4 (N532, N519, N508, N179, N93);
xor XOR2 (N533, N510, N302);
xor XOR2 (N534, N532, N419);
xor XOR2 (N535, N527, N374);
nand NAND2 (N536, N535, N172);
nor NOR3 (N537, N531, N3, N150);
or OR3 (N538, N536, N386, N136);
buf BUF1 (N539, N523);
nor NOR2 (N540, N537, N320);
buf BUF1 (N541, N528);
xor XOR2 (N542, N539, N67);
nor NOR3 (N543, N540, N124, N32);
or OR3 (N544, N533, N472, N74);
and AND2 (N545, N530, N493);
not NOT1 (N546, N529);
not NOT1 (N547, N543);
nand NAND2 (N548, N534, N527);
nor NOR3 (N549, N544, N157, N276);
nand NAND4 (N550, N509, N442, N531, N171);
and AND2 (N551, N549, N542);
buf BUF1 (N552, N159);
or OR4 (N553, N538, N435, N55, N280);
buf BUF1 (N554, N553);
xor XOR2 (N555, N545, N328);
and AND2 (N556, N525, N273);
buf BUF1 (N557, N541);
and AND4 (N558, N547, N246, N37, N467);
xor XOR2 (N559, N557, N453);
or OR3 (N560, N559, N434, N412);
xor XOR2 (N561, N556, N514);
xor XOR2 (N562, N546, N431);
or OR2 (N563, N558, N121);
xor XOR2 (N564, N551, N18);
buf BUF1 (N565, N564);
nand NAND2 (N566, N563, N233);
buf BUF1 (N567, N550);
not NOT1 (N568, N561);
not NOT1 (N569, N560);
or OR4 (N570, N555, N280, N355, N106);
and AND2 (N571, N569, N366);
nor NOR2 (N572, N565, N186);
nand NAND4 (N573, N566, N491, N231, N298);
or OR4 (N574, N573, N468, N50, N568);
and AND4 (N575, N11, N170, N73, N316);
and AND4 (N576, N552, N429, N76, N349);
nand NAND2 (N577, N562, N264);
xor XOR2 (N578, N577, N332);
not NOT1 (N579, N576);
and AND3 (N580, N548, N539, N336);
nor NOR2 (N581, N572, N13);
and AND4 (N582, N578, N84, N383, N461);
nand NAND4 (N583, N582, N436, N440, N131);
buf BUF1 (N584, N575);
not NOT1 (N585, N570);
and AND4 (N586, N584, N340, N261, N330);
xor XOR2 (N587, N583, N78);
not NOT1 (N588, N579);
and AND3 (N589, N586, N271, N91);
nand NAND3 (N590, N585, N246, N165);
not NOT1 (N591, N587);
or OR2 (N592, N590, N3);
or OR4 (N593, N580, N120, N50, N513);
nor NOR3 (N594, N588, N60, N340);
and AND2 (N595, N592, N164);
xor XOR2 (N596, N567, N325);
nand NAND3 (N597, N554, N336, N453);
xor XOR2 (N598, N581, N428);
not NOT1 (N599, N594);
not NOT1 (N600, N596);
and AND4 (N601, N593, N166, N274, N360);
not NOT1 (N602, N595);
buf BUF1 (N603, N571);
and AND3 (N604, N600, N290, N59);
and AND3 (N605, N597, N116, N283);
and AND4 (N606, N602, N228, N35, N46);
buf BUF1 (N607, N598);
not NOT1 (N608, N589);
nand NAND2 (N609, N604, N9);
nand NAND2 (N610, N601, N464);
or OR2 (N611, N608, N183);
and AND3 (N612, N574, N588, N606);
xor XOR2 (N613, N466, N290);
not NOT1 (N614, N591);
nor NOR2 (N615, N611, N144);
nand NAND3 (N616, N605, N393, N172);
xor XOR2 (N617, N614, N32);
nand NAND3 (N618, N612, N226, N173);
buf BUF1 (N619, N613);
not NOT1 (N620, N615);
and AND2 (N621, N599, N437);
not NOT1 (N622, N621);
or OR2 (N623, N607, N567);
not NOT1 (N624, N619);
not NOT1 (N625, N603);
nor NOR2 (N626, N616, N614);
not NOT1 (N627, N617);
xor XOR2 (N628, N624, N478);
or OR4 (N629, N609, N448, N105, N332);
or OR3 (N630, N620, N343, N456);
and AND4 (N631, N630, N83, N74, N352);
buf BUF1 (N632, N625);
buf BUF1 (N633, N631);
xor XOR2 (N634, N627, N17);
or OR2 (N635, N623, N515);
nor NOR3 (N636, N629, N8, N257);
and AND4 (N637, N633, N499, N4, N394);
and AND3 (N638, N635, N187, N54);
buf BUF1 (N639, N638);
and AND4 (N640, N639, N16, N342, N534);
not NOT1 (N641, N622);
buf BUF1 (N642, N641);
buf BUF1 (N643, N642);
buf BUF1 (N644, N632);
nand NAND3 (N645, N628, N65, N8);
xor XOR2 (N646, N636, N422);
or OR2 (N647, N644, N53);
or OR2 (N648, N637, N585);
not NOT1 (N649, N646);
nand NAND4 (N650, N618, N425, N391, N52);
and AND4 (N651, N645, N63, N597, N626);
and AND2 (N652, N567, N626);
nand NAND3 (N653, N650, N337, N200);
buf BUF1 (N654, N634);
nor NOR3 (N655, N649, N432, N61);
or OR3 (N656, N655, N224, N216);
nor NOR3 (N657, N647, N27, N455);
nand NAND4 (N658, N652, N511, N491, N474);
xor XOR2 (N659, N654, N638);
nand NAND4 (N660, N656, N315, N501, N128);
nand NAND4 (N661, N653, N577, N132, N323);
buf BUF1 (N662, N661);
not NOT1 (N663, N640);
nor NOR4 (N664, N643, N260, N433, N603);
nand NAND2 (N665, N610, N237);
xor XOR2 (N666, N648, N317);
not NOT1 (N667, N660);
nand NAND3 (N668, N657, N662, N328);
xor XOR2 (N669, N635, N141);
xor XOR2 (N670, N663, N472);
xor XOR2 (N671, N665, N495);
buf BUF1 (N672, N658);
or OR2 (N673, N669, N211);
nand NAND3 (N674, N671, N648, N152);
and AND4 (N675, N651, N533, N130, N433);
or OR4 (N676, N668, N319, N15, N192);
and AND3 (N677, N670, N488, N29);
xor XOR2 (N678, N674, N196);
buf BUF1 (N679, N673);
not NOT1 (N680, N675);
or OR2 (N681, N679, N351);
nand NAND4 (N682, N666, N41, N358, N609);
or OR4 (N683, N682, N195, N235, N39);
not NOT1 (N684, N683);
or OR3 (N685, N664, N323, N124);
buf BUF1 (N686, N676);
xor XOR2 (N687, N680, N123);
buf BUF1 (N688, N677);
and AND3 (N689, N688, N520, N162);
xor XOR2 (N690, N689, N371);
nor NOR3 (N691, N659, N355, N238);
and AND3 (N692, N687, N575, N203);
and AND2 (N693, N685, N326);
not NOT1 (N694, N678);
not NOT1 (N695, N681);
and AND4 (N696, N694, N216, N68, N595);
nor NOR3 (N697, N686, N294, N617);
nand NAND3 (N698, N667, N353, N275);
and AND4 (N699, N697, N342, N388, N415);
and AND3 (N700, N690, N644, N97);
xor XOR2 (N701, N691, N438);
nor NOR3 (N702, N692, N464, N39);
xor XOR2 (N703, N699, N72);
xor XOR2 (N704, N672, N480);
nor NOR4 (N705, N696, N252, N181, N203);
and AND4 (N706, N703, N427, N123, N436);
buf BUF1 (N707, N704);
nand NAND3 (N708, N695, N200, N341);
and AND2 (N709, N698, N27);
and AND3 (N710, N708, N408, N46);
xor XOR2 (N711, N702, N62);
nor NOR3 (N712, N707, N276, N43);
nor NOR3 (N713, N701, N67, N392);
nor NOR2 (N714, N706, N649);
not NOT1 (N715, N684);
or OR2 (N716, N693, N59);
xor XOR2 (N717, N711, N238);
not NOT1 (N718, N715);
buf BUF1 (N719, N713);
and AND4 (N720, N712, N215, N304, N350);
xor XOR2 (N721, N717, N114);
not NOT1 (N722, N714);
nand NAND4 (N723, N722, N256, N434, N343);
buf BUF1 (N724, N720);
buf BUF1 (N725, N721);
xor XOR2 (N726, N719, N263);
and AND2 (N727, N705, N315);
or OR4 (N728, N726, N306, N181, N77);
buf BUF1 (N729, N724);
not NOT1 (N730, N710);
nand NAND2 (N731, N730, N268);
buf BUF1 (N732, N723);
xor XOR2 (N733, N727, N369);
nand NAND3 (N734, N732, N438, N187);
not NOT1 (N735, N718);
nand NAND4 (N736, N725, N15, N83, N635);
buf BUF1 (N737, N709);
nor NOR2 (N738, N729, N102);
xor XOR2 (N739, N737, N346);
nand NAND2 (N740, N738, N442);
buf BUF1 (N741, N734);
xor XOR2 (N742, N733, N239);
buf BUF1 (N743, N735);
nand NAND3 (N744, N731, N562, N144);
or OR4 (N745, N739, N89, N502, N706);
xor XOR2 (N746, N728, N365);
nand NAND3 (N747, N716, N489, N547);
buf BUF1 (N748, N747);
buf BUF1 (N749, N741);
and AND4 (N750, N746, N40, N600, N3);
nand NAND4 (N751, N748, N596, N471, N81);
xor XOR2 (N752, N700, N545);
and AND3 (N753, N743, N445, N48);
xor XOR2 (N754, N753, N365);
and AND3 (N755, N752, N91, N160);
nor NOR3 (N756, N749, N5, N594);
and AND3 (N757, N736, N194, N409);
nor NOR2 (N758, N740, N683);
not NOT1 (N759, N744);
and AND3 (N760, N759, N720, N111);
or OR4 (N761, N760, N213, N467, N263);
xor XOR2 (N762, N757, N508);
nand NAND4 (N763, N756, N507, N604, N703);
nand NAND2 (N764, N763, N431);
buf BUF1 (N765, N742);
nand NAND4 (N766, N755, N108, N647, N25);
xor XOR2 (N767, N761, N410);
buf BUF1 (N768, N764);
not NOT1 (N769, N750);
nor NOR2 (N770, N745, N636);
or OR4 (N771, N762, N419, N547, N28);
and AND4 (N772, N770, N571, N740, N105);
not NOT1 (N773, N751);
or OR4 (N774, N773, N421, N370, N192);
xor XOR2 (N775, N758, N189);
nor NOR3 (N776, N775, N179, N314);
buf BUF1 (N777, N767);
nor NOR3 (N778, N769, N722, N30);
xor XOR2 (N779, N776, N586);
nor NOR3 (N780, N766, N741, N632);
and AND4 (N781, N778, N320, N48, N248);
not NOT1 (N782, N781);
or OR3 (N783, N780, N310, N227);
nand NAND3 (N784, N779, N541, N383);
or OR4 (N785, N783, N347, N428, N513);
or OR2 (N786, N754, N475);
or OR3 (N787, N768, N700, N241);
xor XOR2 (N788, N786, N708);
nand NAND3 (N789, N782, N620, N275);
not NOT1 (N790, N771);
or OR4 (N791, N784, N470, N80, N534);
xor XOR2 (N792, N765, N105);
buf BUF1 (N793, N789);
buf BUF1 (N794, N791);
not NOT1 (N795, N785);
and AND3 (N796, N793, N69, N487);
xor XOR2 (N797, N796, N151);
not NOT1 (N798, N777);
or OR4 (N799, N788, N302, N180, N499);
nor NOR3 (N800, N799, N569, N594);
or OR3 (N801, N798, N345, N426);
not NOT1 (N802, N795);
nand NAND2 (N803, N787, N410);
nand NAND2 (N804, N801, N786);
nand NAND4 (N805, N792, N275, N368, N712);
nand NAND4 (N806, N802, N764, N113, N359);
or OR3 (N807, N804, N406, N165);
xor XOR2 (N808, N806, N415);
nor NOR2 (N809, N800, N12);
buf BUF1 (N810, N805);
xor XOR2 (N811, N810, N472);
buf BUF1 (N812, N807);
nor NOR4 (N813, N790, N181, N640, N97);
or OR2 (N814, N794, N742);
xor XOR2 (N815, N774, N551);
buf BUF1 (N816, N772);
not NOT1 (N817, N811);
not NOT1 (N818, N817);
xor XOR2 (N819, N809, N543);
buf BUF1 (N820, N819);
nor NOR2 (N821, N803, N643);
nand NAND2 (N822, N797, N102);
xor XOR2 (N823, N814, N602);
xor XOR2 (N824, N821, N689);
nor NOR2 (N825, N823, N295);
nand NAND2 (N826, N816, N78);
not NOT1 (N827, N825);
and AND4 (N828, N813, N196, N636, N640);
xor XOR2 (N829, N828, N502);
xor XOR2 (N830, N822, N748);
not NOT1 (N831, N824);
buf BUF1 (N832, N830);
not NOT1 (N833, N832);
and AND4 (N834, N815, N608, N310, N788);
nand NAND2 (N835, N812, N97);
and AND2 (N836, N829, N615);
or OR2 (N837, N820, N327);
not NOT1 (N838, N836);
xor XOR2 (N839, N833, N609);
and AND2 (N840, N835, N36);
xor XOR2 (N841, N808, N838);
buf BUF1 (N842, N44);
buf BUF1 (N843, N827);
buf BUF1 (N844, N843);
xor XOR2 (N845, N844, N411);
buf BUF1 (N846, N837);
not NOT1 (N847, N841);
nand NAND4 (N848, N842, N775, N758, N257);
or OR4 (N849, N834, N372, N571, N539);
buf BUF1 (N850, N847);
xor XOR2 (N851, N839, N399);
and AND4 (N852, N848, N116, N123, N406);
and AND2 (N853, N851, N82);
nor NOR2 (N854, N845, N137);
nor NOR3 (N855, N854, N685, N634);
or OR3 (N856, N831, N376, N646);
buf BUF1 (N857, N855);
not NOT1 (N858, N852);
nor NOR3 (N859, N857, N279, N155);
nor NOR2 (N860, N859, N625);
nand NAND3 (N861, N826, N140, N159);
not NOT1 (N862, N846);
not NOT1 (N863, N853);
not NOT1 (N864, N863);
or OR4 (N865, N840, N154, N394, N373);
or OR2 (N866, N849, N767);
and AND2 (N867, N864, N69);
xor XOR2 (N868, N860, N100);
or OR2 (N869, N850, N797);
nor NOR2 (N870, N861, N768);
xor XOR2 (N871, N818, N538);
nand NAND4 (N872, N871, N422, N332, N481);
nand NAND2 (N873, N862, N150);
xor XOR2 (N874, N867, N28);
and AND4 (N875, N858, N72, N147, N216);
nand NAND4 (N876, N874, N625, N56, N805);
not NOT1 (N877, N866);
buf BUF1 (N878, N868);
buf BUF1 (N879, N875);
or OR3 (N880, N856, N561, N223);
buf BUF1 (N881, N878);
not NOT1 (N882, N881);
or OR4 (N883, N869, N573, N32, N200);
not NOT1 (N884, N865);
nand NAND2 (N885, N884, N42);
nor NOR3 (N886, N879, N8, N315);
xor XOR2 (N887, N885, N297);
or OR2 (N888, N876, N123);
buf BUF1 (N889, N872);
or OR2 (N890, N880, N603);
and AND3 (N891, N883, N765, N574);
and AND3 (N892, N877, N148, N28);
xor XOR2 (N893, N890, N89);
and AND4 (N894, N893, N626, N315, N725);
buf BUF1 (N895, N894);
not NOT1 (N896, N873);
not NOT1 (N897, N882);
and AND4 (N898, N886, N735, N313, N302);
and AND2 (N899, N891, N71);
nand NAND2 (N900, N896, N571);
buf BUF1 (N901, N898);
nor NOR4 (N902, N889, N468, N184, N137);
nand NAND2 (N903, N899, N686);
not NOT1 (N904, N903);
or OR3 (N905, N870, N786, N648);
and AND4 (N906, N897, N104, N686, N186);
nor NOR4 (N907, N902, N69, N837, N574);
and AND3 (N908, N905, N580, N601);
buf BUF1 (N909, N904);
or OR4 (N910, N895, N490, N654, N694);
and AND4 (N911, N888, N505, N160, N258);
nand NAND3 (N912, N901, N853, N796);
buf BUF1 (N913, N907);
buf BUF1 (N914, N910);
not NOT1 (N915, N913);
buf BUF1 (N916, N912);
nand NAND3 (N917, N916, N414, N692);
or OR4 (N918, N917, N712, N906, N775);
buf BUF1 (N919, N271);
not NOT1 (N920, N887);
and AND3 (N921, N892, N617, N224);
nand NAND4 (N922, N918, N827, N85, N262);
not NOT1 (N923, N911);
xor XOR2 (N924, N920, N75);
nor NOR2 (N925, N924, N178);
nor NOR4 (N926, N908, N45, N11, N800);
buf BUF1 (N927, N921);
nor NOR4 (N928, N915, N29, N127, N515);
nand NAND3 (N929, N926, N548, N555);
nand NAND2 (N930, N919, N850);
and AND2 (N931, N925, N700);
buf BUF1 (N932, N923);
nand NAND2 (N933, N909, N722);
xor XOR2 (N934, N933, N84);
xor XOR2 (N935, N922, N869);
xor XOR2 (N936, N927, N489);
buf BUF1 (N937, N935);
nor NOR3 (N938, N931, N30, N33);
xor XOR2 (N939, N900, N596);
xor XOR2 (N940, N928, N867);
buf BUF1 (N941, N938);
nor NOR2 (N942, N914, N112);
not NOT1 (N943, N934);
and AND3 (N944, N942, N603, N838);
nand NAND2 (N945, N936, N902);
nor NOR3 (N946, N945, N42, N824);
buf BUF1 (N947, N944);
not NOT1 (N948, N946);
nand NAND2 (N949, N947, N641);
nor NOR2 (N950, N937, N369);
or OR4 (N951, N940, N536, N728, N12);
xor XOR2 (N952, N948, N268);
nand NAND2 (N953, N950, N331);
xor XOR2 (N954, N932, N708);
or OR3 (N955, N941, N342, N404);
xor XOR2 (N956, N929, N296);
buf BUF1 (N957, N943);
or OR2 (N958, N949, N936);
and AND3 (N959, N939, N60, N771);
and AND4 (N960, N958, N34, N939, N704);
not NOT1 (N961, N952);
buf BUF1 (N962, N953);
nor NOR2 (N963, N956, N491);
nor NOR3 (N964, N961, N258, N775);
nor NOR2 (N965, N962, N881);
and AND3 (N966, N930, N374, N519);
nor NOR2 (N967, N951, N29);
or OR2 (N968, N957, N701);
buf BUF1 (N969, N954);
xor XOR2 (N970, N969, N301);
and AND4 (N971, N959, N506, N772, N208);
or OR4 (N972, N968, N302, N345, N537);
not NOT1 (N973, N971);
nand NAND3 (N974, N955, N71, N184);
not NOT1 (N975, N973);
or OR2 (N976, N960, N512);
xor XOR2 (N977, N974, N112);
or OR4 (N978, N970, N790, N631, N330);
and AND4 (N979, N967, N946, N396, N452);
nor NOR4 (N980, N976, N972, N846, N604);
and AND2 (N981, N604, N28);
nor NOR4 (N982, N978, N973, N538, N968);
xor XOR2 (N983, N980, N207);
and AND3 (N984, N964, N943, N189);
or OR3 (N985, N966, N139, N436);
nor NOR3 (N986, N981, N516, N648);
or OR2 (N987, N985, N402);
nand NAND3 (N988, N982, N245, N952);
not NOT1 (N989, N975);
nand NAND2 (N990, N987, N860);
nand NAND2 (N991, N979, N60);
buf BUF1 (N992, N984);
nor NOR2 (N993, N986, N728);
xor XOR2 (N994, N990, N809);
not NOT1 (N995, N988);
or OR2 (N996, N965, N130);
or OR2 (N997, N995, N879);
nand NAND4 (N998, N991, N475, N59, N700);
and AND3 (N999, N998, N534, N831);
or OR3 (N1000, N996, N338, N326);
buf BUF1 (N1001, N997);
buf BUF1 (N1002, N999);
nor NOR3 (N1003, N977, N640, N402);
buf BUF1 (N1004, N989);
and AND2 (N1005, N1000, N917);
nand NAND4 (N1006, N1001, N260, N638, N41);
nand NAND2 (N1007, N994, N986);
xor XOR2 (N1008, N1004, N678);
not NOT1 (N1009, N1003);
nand NAND3 (N1010, N993, N718, N239);
nor NOR4 (N1011, N963, N956, N193, N897);
or OR2 (N1012, N1008, N180);
or OR3 (N1013, N992, N791, N441);
and AND3 (N1014, N1005, N82, N849);
buf BUF1 (N1015, N983);
not NOT1 (N1016, N1002);
nand NAND2 (N1017, N1011, N141);
buf BUF1 (N1018, N1010);
nor NOR2 (N1019, N1014, N432);
xor XOR2 (N1020, N1009, N927);
nand NAND4 (N1021, N1020, N303, N264, N725);
nor NOR2 (N1022, N1007, N716);
and AND3 (N1023, N1018, N193, N42);
or OR3 (N1024, N1012, N821, N88);
xor XOR2 (N1025, N1016, N319);
nand NAND2 (N1026, N1019, N885);
not NOT1 (N1027, N1006);
not NOT1 (N1028, N1021);
buf BUF1 (N1029, N1026);
buf BUF1 (N1030, N1023);
nor NOR3 (N1031, N1030, N752, N687);
and AND2 (N1032, N1022, N398);
nand NAND4 (N1033, N1025, N594, N503, N461);
or OR3 (N1034, N1033, N250, N35);
nand NAND3 (N1035, N1024, N835, N835);
buf BUF1 (N1036, N1032);
or OR4 (N1037, N1035, N840, N453, N515);
nor NOR4 (N1038, N1028, N744, N34, N627);
not NOT1 (N1039, N1015);
nand NAND4 (N1040, N1036, N322, N273, N1027);
not NOT1 (N1041, N539);
buf BUF1 (N1042, N1029);
nor NOR4 (N1043, N1038, N66, N338, N294);
nand NAND2 (N1044, N1013, N156);
or OR2 (N1045, N1041, N144);
or OR2 (N1046, N1034, N709);
nand NAND4 (N1047, N1042, N611, N902, N918);
buf BUF1 (N1048, N1039);
not NOT1 (N1049, N1048);
or OR4 (N1050, N1040, N998, N179, N75);
buf BUF1 (N1051, N1049);
and AND2 (N1052, N1043, N156);
xor XOR2 (N1053, N1017, N84);
xor XOR2 (N1054, N1053, N1031);
buf BUF1 (N1055, N139);
nor NOR2 (N1056, N1050, N858);
buf BUF1 (N1057, N1052);
xor XOR2 (N1058, N1046, N1);
xor XOR2 (N1059, N1051, N464);
buf BUF1 (N1060, N1059);
or OR3 (N1061, N1057, N291, N480);
buf BUF1 (N1062, N1045);
not NOT1 (N1063, N1044);
xor XOR2 (N1064, N1058, N13);
buf BUF1 (N1065, N1054);
buf BUF1 (N1066, N1063);
and AND2 (N1067, N1037, N482);
nor NOR3 (N1068, N1055, N890, N674);
not NOT1 (N1069, N1047);
or OR3 (N1070, N1066, N910, N292);
nand NAND4 (N1071, N1069, N968, N263, N957);
and AND4 (N1072, N1061, N441, N104, N56);
buf BUF1 (N1073, N1060);
xor XOR2 (N1074, N1072, N434);
or OR4 (N1075, N1070, N402, N212, N1026);
nand NAND3 (N1076, N1074, N751, N734);
nor NOR2 (N1077, N1073, N20);
xor XOR2 (N1078, N1056, N351);
nor NOR3 (N1079, N1075, N959, N320);
nor NOR3 (N1080, N1079, N1033, N212);
and AND4 (N1081, N1064, N227, N33, N973);
nand NAND2 (N1082, N1071, N772);
buf BUF1 (N1083, N1077);
buf BUF1 (N1084, N1068);
nor NOR4 (N1085, N1081, N556, N848, N466);
xor XOR2 (N1086, N1085, N562);
not NOT1 (N1087, N1086);
buf BUF1 (N1088, N1083);
and AND2 (N1089, N1084, N192);
not NOT1 (N1090, N1076);
or OR3 (N1091, N1089, N100, N903);
nor NOR4 (N1092, N1090, N628, N981, N52);
or OR2 (N1093, N1062, N194);
nand NAND4 (N1094, N1091, N1035, N989, N285);
nand NAND4 (N1095, N1093, N1075, N1012, N333);
and AND2 (N1096, N1092, N882);
xor XOR2 (N1097, N1095, N43);
nor NOR3 (N1098, N1094, N133, N12);
and AND2 (N1099, N1067, N918);
xor XOR2 (N1100, N1087, N867);
xor XOR2 (N1101, N1080, N635);
nor NOR3 (N1102, N1097, N437, N49);
nand NAND4 (N1103, N1099, N586, N647, N799);
nor NOR2 (N1104, N1096, N308);
and AND4 (N1105, N1104, N11, N388, N366);
and AND4 (N1106, N1100, N630, N911, N73);
xor XOR2 (N1107, N1102, N402);
nand NAND2 (N1108, N1101, N239);
xor XOR2 (N1109, N1108, N784);
nor NOR2 (N1110, N1082, N787);
xor XOR2 (N1111, N1106, N927);
not NOT1 (N1112, N1078);
nand NAND4 (N1113, N1098, N738, N468, N607);
or OR3 (N1114, N1103, N809, N60);
nand NAND2 (N1115, N1111, N244);
not NOT1 (N1116, N1105);
nand NAND4 (N1117, N1114, N744, N281, N819);
nand NAND2 (N1118, N1065, N366);
and AND4 (N1119, N1107, N495, N778, N338);
and AND2 (N1120, N1110, N430);
not NOT1 (N1121, N1113);
or OR2 (N1122, N1088, N87);
nor NOR3 (N1123, N1120, N143, N181);
xor XOR2 (N1124, N1117, N176);
nand NAND3 (N1125, N1116, N710, N248);
or OR4 (N1126, N1109, N1120, N1112, N1067);
nor NOR4 (N1127, N238, N939, N985, N903);
xor XOR2 (N1128, N1125, N283);
not NOT1 (N1129, N1124);
nor NOR2 (N1130, N1128, N847);
not NOT1 (N1131, N1123);
or OR2 (N1132, N1122, N519);
or OR3 (N1133, N1132, N376, N152);
nor NOR3 (N1134, N1130, N1097, N48);
not NOT1 (N1135, N1131);
nand NAND4 (N1136, N1129, N1093, N182, N1033);
not NOT1 (N1137, N1127);
nor NOR2 (N1138, N1115, N793);
buf BUF1 (N1139, N1118);
or OR3 (N1140, N1126, N108, N755);
buf BUF1 (N1141, N1119);
not NOT1 (N1142, N1137);
and AND3 (N1143, N1136, N642, N592);
xor XOR2 (N1144, N1141, N1087);
not NOT1 (N1145, N1144);
buf BUF1 (N1146, N1138);
nor NOR2 (N1147, N1140, N181);
nand NAND2 (N1148, N1139, N230);
nand NAND4 (N1149, N1135, N450, N865, N231);
or OR3 (N1150, N1134, N570, N199);
nor NOR2 (N1151, N1145, N1040);
nor NOR4 (N1152, N1151, N942, N339, N985);
xor XOR2 (N1153, N1150, N466);
nand NAND3 (N1154, N1133, N211, N992);
not NOT1 (N1155, N1121);
buf BUF1 (N1156, N1147);
buf BUF1 (N1157, N1153);
not NOT1 (N1158, N1142);
buf BUF1 (N1159, N1154);
not NOT1 (N1160, N1158);
xor XOR2 (N1161, N1160, N502);
not NOT1 (N1162, N1146);
or OR4 (N1163, N1152, N868, N794, N434);
nor NOR2 (N1164, N1163, N75);
or OR4 (N1165, N1155, N734, N848, N1027);
nor NOR3 (N1166, N1161, N481, N593);
buf BUF1 (N1167, N1159);
nor NOR3 (N1168, N1162, N61, N556);
not NOT1 (N1169, N1165);
nor NOR4 (N1170, N1169, N161, N1106, N1015);
nor NOR2 (N1171, N1167, N1059);
nor NOR4 (N1172, N1157, N224, N629, N878);
xor XOR2 (N1173, N1170, N815);
or OR3 (N1174, N1172, N791, N475);
not NOT1 (N1175, N1174);
nor NOR2 (N1176, N1166, N883);
buf BUF1 (N1177, N1143);
and AND2 (N1178, N1175, N623);
and AND4 (N1179, N1171, N790, N497, N953);
nor NOR2 (N1180, N1149, N1085);
nor NOR2 (N1181, N1164, N701);
xor XOR2 (N1182, N1181, N1093);
not NOT1 (N1183, N1178);
nor NOR3 (N1184, N1156, N1013, N519);
and AND2 (N1185, N1176, N817);
and AND2 (N1186, N1173, N931);
nand NAND4 (N1187, N1179, N447, N169, N296);
and AND4 (N1188, N1187, N245, N546, N698);
or OR4 (N1189, N1184, N395, N325, N240);
not NOT1 (N1190, N1186);
buf BUF1 (N1191, N1148);
and AND2 (N1192, N1182, N1029);
nand NAND2 (N1193, N1185, N251);
nand NAND4 (N1194, N1193, N443, N744, N409);
buf BUF1 (N1195, N1194);
and AND4 (N1196, N1168, N629, N775, N694);
not NOT1 (N1197, N1180);
or OR2 (N1198, N1191, N398);
nor NOR3 (N1199, N1177, N951, N601);
not NOT1 (N1200, N1197);
or OR4 (N1201, N1195, N1047, N1193, N548);
and AND3 (N1202, N1188, N20, N243);
xor XOR2 (N1203, N1202, N437);
nor NOR2 (N1204, N1198, N938);
nand NAND3 (N1205, N1199, N276, N704);
or OR3 (N1206, N1190, N894, N292);
not NOT1 (N1207, N1206);
buf BUF1 (N1208, N1196);
not NOT1 (N1209, N1201);
or OR4 (N1210, N1205, N986, N92, N578);
xor XOR2 (N1211, N1189, N1110);
nand NAND4 (N1212, N1209, N765, N1204, N744);
not NOT1 (N1213, N483);
and AND4 (N1214, N1213, N292, N1088, N1123);
buf BUF1 (N1215, N1211);
or OR4 (N1216, N1200, N964, N109, N519);
buf BUF1 (N1217, N1214);
buf BUF1 (N1218, N1207);
not NOT1 (N1219, N1216);
buf BUF1 (N1220, N1219);
or OR3 (N1221, N1192, N649, N273);
buf BUF1 (N1222, N1217);
buf BUF1 (N1223, N1203);
or OR3 (N1224, N1220, N232, N855);
nand NAND4 (N1225, N1224, N1044, N946, N289);
buf BUF1 (N1226, N1210);
or OR3 (N1227, N1183, N1135, N1146);
buf BUF1 (N1228, N1212);
not NOT1 (N1229, N1208);
nor NOR2 (N1230, N1223, N1138);
xor XOR2 (N1231, N1222, N288);
nand NAND3 (N1232, N1231, N747, N23);
nand NAND2 (N1233, N1218, N870);
nand NAND4 (N1234, N1233, N664, N1154, N832);
nand NAND2 (N1235, N1227, N82);
xor XOR2 (N1236, N1225, N746);
nor NOR4 (N1237, N1236, N966, N239, N823);
xor XOR2 (N1238, N1215, N626);
or OR3 (N1239, N1229, N257, N1093);
buf BUF1 (N1240, N1234);
xor XOR2 (N1241, N1230, N32);
xor XOR2 (N1242, N1232, N1009);
buf BUF1 (N1243, N1237);
nor NOR3 (N1244, N1240, N412, N713);
xor XOR2 (N1245, N1242, N33);
nor NOR4 (N1246, N1235, N63, N2, N1129);
or OR2 (N1247, N1228, N591);
buf BUF1 (N1248, N1239);
nand NAND4 (N1249, N1221, N622, N756, N140);
and AND4 (N1250, N1247, N6, N637, N758);
or OR4 (N1251, N1245, N194, N958, N23);
xor XOR2 (N1252, N1244, N555);
nand NAND2 (N1253, N1249, N512);
buf BUF1 (N1254, N1252);
xor XOR2 (N1255, N1248, N1094);
buf BUF1 (N1256, N1255);
nor NOR2 (N1257, N1253, N349);
nor NOR4 (N1258, N1257, N632, N315, N879);
xor XOR2 (N1259, N1238, N500);
nor NOR3 (N1260, N1259, N1113, N829);
and AND3 (N1261, N1250, N26, N114);
and AND2 (N1262, N1241, N47);
xor XOR2 (N1263, N1262, N514);
xor XOR2 (N1264, N1260, N566);
not NOT1 (N1265, N1251);
buf BUF1 (N1266, N1264);
nand NAND4 (N1267, N1266, N766, N825, N364);
xor XOR2 (N1268, N1226, N805);
or OR3 (N1269, N1243, N1189, N489);
xor XOR2 (N1270, N1267, N156);
and AND2 (N1271, N1263, N425);
nand NAND3 (N1272, N1271, N502, N19);
or OR2 (N1273, N1269, N613);
nor NOR2 (N1274, N1246, N1040);
or OR4 (N1275, N1274, N754, N20, N848);
not NOT1 (N1276, N1261);
buf BUF1 (N1277, N1256);
buf BUF1 (N1278, N1254);
not NOT1 (N1279, N1275);
not NOT1 (N1280, N1276);
nor NOR4 (N1281, N1270, N909, N1267, N133);
and AND2 (N1282, N1277, N40);
and AND4 (N1283, N1282, N480, N189, N178);
nand NAND3 (N1284, N1273, N370, N824);
nor NOR3 (N1285, N1268, N1201, N1037);
and AND2 (N1286, N1265, N749);
not NOT1 (N1287, N1279);
not NOT1 (N1288, N1284);
nor NOR3 (N1289, N1286, N488, N170);
nand NAND2 (N1290, N1278, N697);
and AND4 (N1291, N1287, N1040, N1211, N1132);
xor XOR2 (N1292, N1291, N625);
buf BUF1 (N1293, N1280);
nand NAND4 (N1294, N1288, N664, N568, N721);
nand NAND4 (N1295, N1289, N1293, N1072, N1261);
xor XOR2 (N1296, N322, N1236);
xor XOR2 (N1297, N1285, N358);
nand NAND3 (N1298, N1290, N353, N391);
buf BUF1 (N1299, N1295);
buf BUF1 (N1300, N1297);
and AND2 (N1301, N1299, N1295);
nor NOR4 (N1302, N1281, N103, N232, N676);
xor XOR2 (N1303, N1258, N242);
and AND2 (N1304, N1292, N658);
buf BUF1 (N1305, N1298);
and AND4 (N1306, N1303, N1199, N1302, N1255);
and AND3 (N1307, N975, N944, N597);
not NOT1 (N1308, N1301);
and AND3 (N1309, N1305, N1086, N156);
nand NAND4 (N1310, N1283, N1050, N160, N710);
xor XOR2 (N1311, N1308, N1093);
nand NAND2 (N1312, N1300, N860);
and AND3 (N1313, N1309, N96, N80);
or OR2 (N1314, N1313, N291);
or OR2 (N1315, N1304, N39);
not NOT1 (N1316, N1314);
xor XOR2 (N1317, N1311, N1315);
and AND4 (N1318, N752, N482, N1008, N191);
xor XOR2 (N1319, N1312, N1066);
xor XOR2 (N1320, N1316, N1267);
nand NAND3 (N1321, N1306, N741, N683);
nor NOR4 (N1322, N1296, N488, N783, N157);
buf BUF1 (N1323, N1272);
xor XOR2 (N1324, N1322, N1173);
nand NAND3 (N1325, N1307, N783, N646);
and AND2 (N1326, N1318, N788);
not NOT1 (N1327, N1325);
and AND4 (N1328, N1320, N1110, N656, N112);
and AND4 (N1329, N1324, N424, N95, N1025);
nand NAND3 (N1330, N1294, N408, N1182);
or OR3 (N1331, N1329, N409, N173);
nor NOR2 (N1332, N1319, N1242);
not NOT1 (N1333, N1327);
or OR3 (N1334, N1317, N1312, N756);
and AND3 (N1335, N1321, N17, N559);
and AND3 (N1336, N1323, N12, N642);
nor NOR4 (N1337, N1330, N1131, N198, N756);
nor NOR3 (N1338, N1337, N945, N1220);
or OR2 (N1339, N1335, N867);
nand NAND3 (N1340, N1336, N1170, N1078);
buf BUF1 (N1341, N1334);
xor XOR2 (N1342, N1328, N330);
nor NOR2 (N1343, N1340, N647);
xor XOR2 (N1344, N1338, N782);
buf BUF1 (N1345, N1310);
buf BUF1 (N1346, N1342);
or OR4 (N1347, N1345, N195, N1229, N199);
and AND3 (N1348, N1347, N30, N1041);
and AND4 (N1349, N1348, N588, N588, N730);
nor NOR3 (N1350, N1346, N1289, N1212);
nand NAND3 (N1351, N1339, N570, N415);
and AND4 (N1352, N1341, N881, N878, N876);
not NOT1 (N1353, N1351);
xor XOR2 (N1354, N1350, N593);
buf BUF1 (N1355, N1354);
not NOT1 (N1356, N1353);
and AND4 (N1357, N1349, N695, N102, N1254);
nor NOR3 (N1358, N1332, N1054, N1067);
or OR4 (N1359, N1343, N61, N568, N123);
buf BUF1 (N1360, N1357);
not NOT1 (N1361, N1356);
nor NOR2 (N1362, N1355, N672);
nor NOR2 (N1363, N1361, N787);
nor NOR2 (N1364, N1359, N322);
buf BUF1 (N1365, N1333);
nor NOR2 (N1366, N1360, N1281);
or OR3 (N1367, N1331, N1058, N4);
xor XOR2 (N1368, N1358, N324);
nor NOR3 (N1369, N1362, N740, N528);
xor XOR2 (N1370, N1365, N893);
and AND4 (N1371, N1352, N51, N14, N107);
nor NOR2 (N1372, N1344, N1080);
buf BUF1 (N1373, N1366);
buf BUF1 (N1374, N1369);
nand NAND2 (N1375, N1374, N559);
xor XOR2 (N1376, N1326, N153);
nor NOR4 (N1377, N1373, N182, N1089, N931);
nor NOR2 (N1378, N1377, N1200);
nand NAND3 (N1379, N1378, N1030, N950);
or OR2 (N1380, N1370, N554);
not NOT1 (N1381, N1372);
nand NAND2 (N1382, N1364, N333);
nand NAND3 (N1383, N1382, N1035, N1177);
nor NOR2 (N1384, N1367, N1113);
nor NOR4 (N1385, N1371, N127, N602, N543);
buf BUF1 (N1386, N1383);
or OR4 (N1387, N1376, N1359, N477, N236);
buf BUF1 (N1388, N1368);
not NOT1 (N1389, N1386);
xor XOR2 (N1390, N1380, N1349);
xor XOR2 (N1391, N1363, N1218);
and AND2 (N1392, N1389, N840);
nand NAND2 (N1393, N1390, N753);
xor XOR2 (N1394, N1379, N1194);
nand NAND3 (N1395, N1394, N1271, N976);
nand NAND3 (N1396, N1395, N914, N205);
or OR3 (N1397, N1387, N4, N775);
or OR2 (N1398, N1397, N344);
and AND3 (N1399, N1393, N397, N499);
and AND3 (N1400, N1375, N13, N1098);
xor XOR2 (N1401, N1391, N107);
nand NAND2 (N1402, N1398, N423);
nor NOR4 (N1403, N1388, N905, N28, N35);
xor XOR2 (N1404, N1396, N227);
or OR4 (N1405, N1402, N424, N588, N1348);
buf BUF1 (N1406, N1403);
xor XOR2 (N1407, N1405, N1384);
or OR3 (N1408, N682, N765, N21);
and AND4 (N1409, N1392, N819, N72, N49);
xor XOR2 (N1410, N1407, N678);
nand NAND3 (N1411, N1400, N183, N1048);
and AND3 (N1412, N1410, N1262, N974);
nor NOR3 (N1413, N1399, N1407, N972);
not NOT1 (N1414, N1413);
and AND3 (N1415, N1409, N1246, N187);
not NOT1 (N1416, N1385);
xor XOR2 (N1417, N1401, N1293);
nand NAND2 (N1418, N1412, N862);
or OR4 (N1419, N1417, N679, N1287, N120);
buf BUF1 (N1420, N1408);
or OR2 (N1421, N1406, N12);
xor XOR2 (N1422, N1418, N921);
or OR2 (N1423, N1420, N1215);
buf BUF1 (N1424, N1411);
or OR3 (N1425, N1423, N463, N1326);
nand NAND3 (N1426, N1421, N365, N1367);
nor NOR4 (N1427, N1424, N1191, N1094, N1080);
and AND2 (N1428, N1415, N1088);
nand NAND4 (N1429, N1427, N90, N474, N135);
and AND2 (N1430, N1429, N83);
nand NAND3 (N1431, N1381, N1161, N148);
and AND2 (N1432, N1422, N735);
or OR3 (N1433, N1416, N450, N186);
not NOT1 (N1434, N1414);
and AND3 (N1435, N1434, N775, N535);
or OR2 (N1436, N1425, N150);
not NOT1 (N1437, N1419);
xor XOR2 (N1438, N1433, N671);
nor NOR4 (N1439, N1435, N958, N248, N838);
nor NOR2 (N1440, N1431, N1339);
not NOT1 (N1441, N1436);
nor NOR3 (N1442, N1440, N551, N1418);
nand NAND2 (N1443, N1438, N1302);
or OR2 (N1444, N1432, N61);
not NOT1 (N1445, N1439);
xor XOR2 (N1446, N1437, N144);
nand NAND2 (N1447, N1430, N821);
not NOT1 (N1448, N1442);
and AND3 (N1449, N1444, N1035, N928);
nand NAND2 (N1450, N1426, N313);
nand NAND3 (N1451, N1447, N107, N1181);
nand NAND3 (N1452, N1404, N449, N49);
xor XOR2 (N1453, N1446, N835);
not NOT1 (N1454, N1452);
buf BUF1 (N1455, N1443);
or OR4 (N1456, N1451, N475, N1260, N139);
nand NAND2 (N1457, N1455, N826);
nor NOR3 (N1458, N1457, N904, N1269);
buf BUF1 (N1459, N1453);
buf BUF1 (N1460, N1448);
or OR3 (N1461, N1460, N729, N481);
xor XOR2 (N1462, N1456, N1209);
buf BUF1 (N1463, N1445);
buf BUF1 (N1464, N1450);
or OR3 (N1465, N1441, N327, N1135);
nand NAND3 (N1466, N1459, N82, N129);
not NOT1 (N1467, N1464);
nor NOR3 (N1468, N1462, N1048, N921);
xor XOR2 (N1469, N1449, N1333);
nand NAND4 (N1470, N1465, N241, N44, N51);
not NOT1 (N1471, N1469);
nand NAND4 (N1472, N1466, N1340, N659, N269);
xor XOR2 (N1473, N1454, N1306);
xor XOR2 (N1474, N1458, N1391);
or OR3 (N1475, N1470, N1099, N817);
not NOT1 (N1476, N1471);
xor XOR2 (N1477, N1463, N750);
or OR2 (N1478, N1475, N709);
buf BUF1 (N1479, N1477);
nor NOR3 (N1480, N1476, N223, N580);
and AND4 (N1481, N1474, N30, N511, N1086);
xor XOR2 (N1482, N1480, N1412);
and AND3 (N1483, N1478, N775, N8);
nand NAND3 (N1484, N1479, N1235, N161);
xor XOR2 (N1485, N1461, N774);
not NOT1 (N1486, N1428);
not NOT1 (N1487, N1482);
nand NAND4 (N1488, N1481, N964, N237, N557);
xor XOR2 (N1489, N1483, N80);
nand NAND4 (N1490, N1467, N467, N451, N823);
buf BUF1 (N1491, N1472);
not NOT1 (N1492, N1489);
or OR2 (N1493, N1484, N1077);
nand NAND2 (N1494, N1488, N580);
and AND2 (N1495, N1468, N62);
not NOT1 (N1496, N1490);
buf BUF1 (N1497, N1492);
not NOT1 (N1498, N1486);
not NOT1 (N1499, N1495);
xor XOR2 (N1500, N1493, N764);
buf BUF1 (N1501, N1499);
nor NOR4 (N1502, N1500, N513, N1482, N1068);
or OR2 (N1503, N1491, N117);
not NOT1 (N1504, N1487);
and AND3 (N1505, N1485, N696, N1396);
and AND4 (N1506, N1497, N75, N184, N1485);
not NOT1 (N1507, N1503);
not NOT1 (N1508, N1507);
nor NOR3 (N1509, N1504, N914, N1075);
and AND3 (N1510, N1498, N996, N379);
or OR4 (N1511, N1508, N972, N1199, N1265);
nor NOR2 (N1512, N1506, N33);
or OR3 (N1513, N1502, N1508, N561);
buf BUF1 (N1514, N1496);
buf BUF1 (N1515, N1512);
xor XOR2 (N1516, N1505, N1430);
nor NOR3 (N1517, N1494, N1228, N421);
nand NAND4 (N1518, N1501, N789, N296, N889);
xor XOR2 (N1519, N1516, N520);
nand NAND4 (N1520, N1519, N347, N1201, N1356);
not NOT1 (N1521, N1514);
and AND4 (N1522, N1518, N1149, N689, N1435);
nand NAND2 (N1523, N1515, N1146);
buf BUF1 (N1524, N1522);
not NOT1 (N1525, N1524);
nor NOR4 (N1526, N1509, N263, N992, N677);
and AND2 (N1527, N1473, N219);
buf BUF1 (N1528, N1520);
not NOT1 (N1529, N1527);
xor XOR2 (N1530, N1511, N30);
nand NAND3 (N1531, N1510, N1315, N1094);
xor XOR2 (N1532, N1517, N1312);
or OR2 (N1533, N1531, N1311);
not NOT1 (N1534, N1526);
nor NOR2 (N1535, N1523, N41);
nor NOR3 (N1536, N1529, N774, N421);
and AND2 (N1537, N1525, N698);
and AND3 (N1538, N1528, N373, N558);
nand NAND3 (N1539, N1530, N465, N744);
buf BUF1 (N1540, N1521);
xor XOR2 (N1541, N1532, N147);
not NOT1 (N1542, N1513);
not NOT1 (N1543, N1534);
xor XOR2 (N1544, N1541, N531);
buf BUF1 (N1545, N1543);
not NOT1 (N1546, N1533);
buf BUF1 (N1547, N1542);
or OR3 (N1548, N1539, N1544, N740);
and AND3 (N1549, N380, N12, N671);
nor NOR2 (N1550, N1538, N1162);
nor NOR3 (N1551, N1547, N215, N1298);
not NOT1 (N1552, N1550);
and AND2 (N1553, N1551, N908);
not NOT1 (N1554, N1546);
nor NOR2 (N1555, N1549, N1375);
buf BUF1 (N1556, N1554);
nor NOR3 (N1557, N1537, N1232, N82);
or OR4 (N1558, N1552, N1288, N700, N1391);
not NOT1 (N1559, N1536);
nor NOR4 (N1560, N1540, N769, N314, N308);
nor NOR2 (N1561, N1560, N871);
not NOT1 (N1562, N1553);
or OR3 (N1563, N1557, N1140, N821);
xor XOR2 (N1564, N1535, N1212);
buf BUF1 (N1565, N1545);
xor XOR2 (N1566, N1548, N146);
and AND3 (N1567, N1558, N188, N1011);
nor NOR3 (N1568, N1566, N739, N554);
xor XOR2 (N1569, N1565, N1496);
or OR3 (N1570, N1569, N1381, N1348);
buf BUF1 (N1571, N1568);
xor XOR2 (N1572, N1555, N1256);
and AND2 (N1573, N1564, N228);
nand NAND2 (N1574, N1571, N1075);
nor NOR3 (N1575, N1561, N680, N1442);
xor XOR2 (N1576, N1575, N816);
buf BUF1 (N1577, N1574);
xor XOR2 (N1578, N1576, N291);
not NOT1 (N1579, N1578);
nand NAND3 (N1580, N1570, N1025, N72);
nor NOR4 (N1581, N1567, N1303, N865, N1453);
xor XOR2 (N1582, N1579, N420);
and AND3 (N1583, N1559, N158, N752);
buf BUF1 (N1584, N1582);
or OR2 (N1585, N1581, N1443);
nand NAND3 (N1586, N1572, N1582, N1045);
nand NAND2 (N1587, N1585, N109);
not NOT1 (N1588, N1577);
nor NOR2 (N1589, N1556, N976);
or OR2 (N1590, N1587, N1069);
nor NOR3 (N1591, N1590, N258, N1167);
and AND4 (N1592, N1589, N756, N1014, N1124);
xor XOR2 (N1593, N1586, N1511);
nand NAND3 (N1594, N1592, N363, N156);
and AND3 (N1595, N1583, N1403, N375);
and AND4 (N1596, N1594, N868, N808, N1393);
and AND2 (N1597, N1588, N764);
or OR4 (N1598, N1584, N1205, N107, N886);
nor NOR3 (N1599, N1563, N537, N149);
nand NAND2 (N1600, N1597, N938);
nor NOR4 (N1601, N1600, N1279, N1600, N925);
xor XOR2 (N1602, N1593, N1464);
buf BUF1 (N1603, N1573);
nor NOR3 (N1604, N1602, N78, N202);
buf BUF1 (N1605, N1595);
buf BUF1 (N1606, N1603);
buf BUF1 (N1607, N1604);
xor XOR2 (N1608, N1606, N1548);
buf BUF1 (N1609, N1607);
or OR3 (N1610, N1591, N1115, N1096);
nor NOR2 (N1611, N1609, N466);
xor XOR2 (N1612, N1611, N295);
buf BUF1 (N1613, N1580);
nor NOR4 (N1614, N1608, N573, N1310, N209);
xor XOR2 (N1615, N1601, N1238);
xor XOR2 (N1616, N1613, N744);
or OR3 (N1617, N1616, N1207, N7);
or OR2 (N1618, N1614, N1006);
and AND2 (N1619, N1612, N1590);
nor NOR2 (N1620, N1605, N439);
nand NAND2 (N1621, N1615, N449);
buf BUF1 (N1622, N1562);
xor XOR2 (N1623, N1618, N581);
or OR3 (N1624, N1620, N348, N323);
xor XOR2 (N1625, N1622, N1080);
or OR2 (N1626, N1596, N466);
and AND3 (N1627, N1623, N867, N138);
nand NAND3 (N1628, N1598, N937, N1532);
and AND4 (N1629, N1624, N977, N1385, N170);
or OR2 (N1630, N1621, N1240);
and AND4 (N1631, N1628, N1368, N855, N939);
xor XOR2 (N1632, N1626, N262);
and AND2 (N1633, N1630, N669);
buf BUF1 (N1634, N1627);
and AND4 (N1635, N1625, N670, N1140, N196);
xor XOR2 (N1636, N1633, N973);
buf BUF1 (N1637, N1610);
or OR2 (N1638, N1637, N1049);
nor NOR3 (N1639, N1619, N701, N1470);
not NOT1 (N1640, N1639);
and AND2 (N1641, N1634, N777);
nor NOR4 (N1642, N1629, N1377, N1273, N831);
not NOT1 (N1643, N1640);
buf BUF1 (N1644, N1642);
nand NAND4 (N1645, N1636, N299, N650, N342);
and AND3 (N1646, N1643, N1254, N630);
and AND4 (N1647, N1635, N440, N1218, N622);
not NOT1 (N1648, N1617);
and AND2 (N1649, N1631, N1480);
not NOT1 (N1650, N1648);
xor XOR2 (N1651, N1644, N513);
and AND4 (N1652, N1649, N1383, N1095, N164);
not NOT1 (N1653, N1650);
and AND4 (N1654, N1632, N523, N1624, N118);
or OR3 (N1655, N1653, N629, N1367);
or OR3 (N1656, N1655, N1048, N195);
nor NOR2 (N1657, N1641, N757);
or OR2 (N1658, N1654, N811);
and AND2 (N1659, N1599, N1614);
xor XOR2 (N1660, N1647, N666);
not NOT1 (N1661, N1660);
nand NAND2 (N1662, N1638, N477);
not NOT1 (N1663, N1657);
nand NAND3 (N1664, N1659, N1359, N810);
not NOT1 (N1665, N1656);
nor NOR3 (N1666, N1665, N1205, N1184);
buf BUF1 (N1667, N1646);
or OR3 (N1668, N1664, N414, N316);
buf BUF1 (N1669, N1666);
nand NAND4 (N1670, N1663, N593, N1103, N1668);
nand NAND4 (N1671, N731, N1379, N695, N1648);
and AND4 (N1672, N1651, N633, N658, N810);
not NOT1 (N1673, N1661);
and AND2 (N1674, N1645, N1005);
or OR4 (N1675, N1674, N59, N340, N779);
nor NOR3 (N1676, N1673, N1385, N915);
xor XOR2 (N1677, N1671, N681);
or OR4 (N1678, N1667, N1552, N1574, N649);
nor NOR3 (N1679, N1678, N222, N1511);
or OR3 (N1680, N1675, N1160, N1323);
or OR2 (N1681, N1658, N820);
not NOT1 (N1682, N1680);
and AND4 (N1683, N1672, N1436, N1350, N656);
or OR4 (N1684, N1669, N1292, N152, N1517);
xor XOR2 (N1685, N1679, N492);
nand NAND4 (N1686, N1685, N1643, N729, N301);
buf BUF1 (N1687, N1652);
nor NOR3 (N1688, N1662, N1090, N1579);
nor NOR2 (N1689, N1684, N1529);
buf BUF1 (N1690, N1686);
nand NAND2 (N1691, N1677, N982);
nor NOR3 (N1692, N1670, N1565, N477);
nor NOR3 (N1693, N1689, N1510, N336);
nand NAND2 (N1694, N1692, N569);
and AND2 (N1695, N1693, N1680);
buf BUF1 (N1696, N1681);
nor NOR3 (N1697, N1676, N1068, N1045);
nor NOR2 (N1698, N1687, N1184);
and AND3 (N1699, N1683, N233, N1553);
nor NOR4 (N1700, N1691, N335, N1653, N1425);
nor NOR3 (N1701, N1694, N140, N110);
xor XOR2 (N1702, N1699, N472);
xor XOR2 (N1703, N1682, N461);
and AND3 (N1704, N1695, N1576, N1565);
or OR2 (N1705, N1697, N1293);
buf BUF1 (N1706, N1701);
or OR3 (N1707, N1698, N1281, N693);
buf BUF1 (N1708, N1700);
or OR2 (N1709, N1708, N888);
or OR3 (N1710, N1703, N190, N1515);
nand NAND2 (N1711, N1709, N1158);
buf BUF1 (N1712, N1690);
nand NAND3 (N1713, N1696, N155, N1062);
nor NOR2 (N1714, N1713, N925);
or OR2 (N1715, N1706, N1212);
nand NAND2 (N1716, N1711, N1238);
and AND3 (N1717, N1715, N1200, N1126);
not NOT1 (N1718, N1705);
nor NOR4 (N1719, N1714, N998, N1146, N1062);
nor NOR3 (N1720, N1717, N1569, N576);
and AND4 (N1721, N1716, N948, N540, N362);
buf BUF1 (N1722, N1712);
not NOT1 (N1723, N1702);
and AND3 (N1724, N1721, N1419, N1626);
nor NOR4 (N1725, N1688, N778, N357, N878);
or OR2 (N1726, N1704, N416);
not NOT1 (N1727, N1723);
and AND2 (N1728, N1727, N823);
and AND3 (N1729, N1728, N641, N249);
nand NAND3 (N1730, N1725, N386, N1325);
not NOT1 (N1731, N1719);
nor NOR2 (N1732, N1718, N1390);
nor NOR4 (N1733, N1722, N299, N1169, N1250);
buf BUF1 (N1734, N1724);
nand NAND4 (N1735, N1733, N921, N656, N1589);
not NOT1 (N1736, N1729);
or OR3 (N1737, N1731, N1677, N146);
nand NAND3 (N1738, N1736, N1, N1271);
and AND3 (N1739, N1730, N573, N922);
and AND2 (N1740, N1737, N772);
and AND4 (N1741, N1710, N856, N370, N1180);
buf BUF1 (N1742, N1739);
and AND4 (N1743, N1720, N1628, N238, N1001);
buf BUF1 (N1744, N1735);
and AND4 (N1745, N1734, N1218, N1683, N1304);
nand NAND4 (N1746, N1745, N345, N705, N337);
not NOT1 (N1747, N1746);
not NOT1 (N1748, N1707);
and AND3 (N1749, N1726, N840, N1004);
nand NAND4 (N1750, N1738, N1545, N1427, N634);
xor XOR2 (N1751, N1750, N1467);
xor XOR2 (N1752, N1742, N535);
nand NAND3 (N1753, N1740, N765, N1731);
not NOT1 (N1754, N1748);
not NOT1 (N1755, N1754);
or OR4 (N1756, N1732, N178, N1615, N246);
or OR2 (N1757, N1753, N1523);
nor NOR2 (N1758, N1752, N1684);
nand NAND2 (N1759, N1756, N1509);
buf BUF1 (N1760, N1759);
or OR4 (N1761, N1741, N162, N400, N1340);
not NOT1 (N1762, N1751);
buf BUF1 (N1763, N1762);
and AND4 (N1764, N1760, N1396, N1092, N707);
xor XOR2 (N1765, N1747, N584);
nor NOR3 (N1766, N1749, N870, N1508);
buf BUF1 (N1767, N1764);
nand NAND2 (N1768, N1767, N1573);
xor XOR2 (N1769, N1765, N1695);
nand NAND2 (N1770, N1757, N116);
or OR4 (N1771, N1744, N103, N687, N871);
and AND3 (N1772, N1758, N579, N1164);
or OR2 (N1773, N1771, N894);
not NOT1 (N1774, N1755);
nand NAND4 (N1775, N1770, N1161, N609, N1079);
buf BUF1 (N1776, N1766);
and AND3 (N1777, N1773, N66, N240);
not NOT1 (N1778, N1769);
nand NAND4 (N1779, N1763, N1701, N264, N1124);
not NOT1 (N1780, N1775);
xor XOR2 (N1781, N1780, N1323);
buf BUF1 (N1782, N1778);
not NOT1 (N1783, N1776);
buf BUF1 (N1784, N1743);
nand NAND3 (N1785, N1772, N125, N1340);
nand NAND4 (N1786, N1783, N1519, N1431, N484);
buf BUF1 (N1787, N1782);
xor XOR2 (N1788, N1784, N855);
xor XOR2 (N1789, N1781, N331);
nor NOR4 (N1790, N1777, N1694, N695, N363);
buf BUF1 (N1791, N1785);
buf BUF1 (N1792, N1790);
or OR2 (N1793, N1792, N442);
or OR2 (N1794, N1793, N1698);
buf BUF1 (N1795, N1788);
xor XOR2 (N1796, N1786, N404);
xor XOR2 (N1797, N1794, N162);
or OR4 (N1798, N1797, N1718, N1135, N554);
and AND3 (N1799, N1789, N150, N1058);
nand NAND3 (N1800, N1768, N501, N954);
buf BUF1 (N1801, N1800);
nand NAND2 (N1802, N1761, N1508);
buf BUF1 (N1803, N1774);
nand NAND3 (N1804, N1787, N363, N210);
or OR2 (N1805, N1779, N934);
and AND3 (N1806, N1804, N510, N493);
nand NAND3 (N1807, N1798, N513, N856);
not NOT1 (N1808, N1801);
nor NOR2 (N1809, N1803, N451);
and AND3 (N1810, N1791, N547, N1494);
nand NAND3 (N1811, N1799, N1651, N964);
not NOT1 (N1812, N1802);
or OR2 (N1813, N1808, N10);
nor NOR3 (N1814, N1809, N1028, N1083);
nor NOR2 (N1815, N1806, N1420);
xor XOR2 (N1816, N1811, N1479);
buf BUF1 (N1817, N1813);
and AND4 (N1818, N1807, N700, N1729, N462);
xor XOR2 (N1819, N1815, N1016);
not NOT1 (N1820, N1795);
and AND2 (N1821, N1816, N1730);
nand NAND2 (N1822, N1810, N328);
xor XOR2 (N1823, N1817, N589);
xor XOR2 (N1824, N1818, N1767);
buf BUF1 (N1825, N1812);
and AND4 (N1826, N1823, N764, N980, N1654);
nor NOR3 (N1827, N1826, N494, N535);
buf BUF1 (N1828, N1825);
and AND4 (N1829, N1819, N1532, N439, N283);
and AND3 (N1830, N1821, N349, N512);
or OR2 (N1831, N1829, N151);
buf BUF1 (N1832, N1796);
or OR3 (N1833, N1824, N582, N803);
buf BUF1 (N1834, N1827);
nand NAND4 (N1835, N1828, N384, N1480, N655);
nor NOR4 (N1836, N1833, N1584, N562, N1223);
nor NOR4 (N1837, N1814, N1096, N329, N1438);
nand NAND3 (N1838, N1831, N1075, N1407);
or OR3 (N1839, N1830, N1357, N61);
nand NAND4 (N1840, N1836, N627, N614, N320);
and AND3 (N1841, N1839, N946, N615);
xor XOR2 (N1842, N1838, N1567);
buf BUF1 (N1843, N1841);
or OR2 (N1844, N1834, N635);
and AND2 (N1845, N1842, N1268);
not NOT1 (N1846, N1805);
not NOT1 (N1847, N1837);
nor NOR4 (N1848, N1843, N1009, N1417, N80);
nand NAND3 (N1849, N1847, N548, N959);
and AND4 (N1850, N1835, N1165, N1286, N287);
or OR4 (N1851, N1848, N1096, N1207, N364);
nand NAND4 (N1852, N1846, N1117, N637, N665);
xor XOR2 (N1853, N1840, N91);
and AND4 (N1854, N1850, N292, N1781, N63);
buf BUF1 (N1855, N1844);
not NOT1 (N1856, N1851);
and AND4 (N1857, N1852, N122, N1650, N992);
xor XOR2 (N1858, N1854, N836);
not NOT1 (N1859, N1858);
not NOT1 (N1860, N1853);
not NOT1 (N1861, N1822);
not NOT1 (N1862, N1845);
not NOT1 (N1863, N1849);
not NOT1 (N1864, N1832);
or OR3 (N1865, N1862, N1233, N565);
and AND4 (N1866, N1863, N534, N1350, N1708);
or OR4 (N1867, N1820, N817, N1213, N1539);
nor NOR2 (N1868, N1867, N619);
not NOT1 (N1869, N1864);
or OR3 (N1870, N1857, N1083, N1717);
not NOT1 (N1871, N1855);
nor NOR4 (N1872, N1865, N1540, N1365, N300);
or OR3 (N1873, N1856, N24, N577);
nand NAND4 (N1874, N1860, N1578, N1396, N1399);
xor XOR2 (N1875, N1874, N1421);
nand NAND3 (N1876, N1861, N1696, N1108);
or OR3 (N1877, N1859, N1666, N1364);
xor XOR2 (N1878, N1876, N825);
and AND2 (N1879, N1870, N1875);
nand NAND2 (N1880, N923, N1583);
or OR4 (N1881, N1877, N189, N1475, N990);
xor XOR2 (N1882, N1872, N1222);
and AND2 (N1883, N1869, N846);
nor NOR3 (N1884, N1879, N811, N263);
not NOT1 (N1885, N1882);
xor XOR2 (N1886, N1881, N1358);
xor XOR2 (N1887, N1868, N1189);
nor NOR2 (N1888, N1886, N439);
buf BUF1 (N1889, N1871);
nor NOR2 (N1890, N1888, N805);
and AND4 (N1891, N1890, N729, N435, N1658);
xor XOR2 (N1892, N1873, N918);
nor NOR2 (N1893, N1884, N1414);
and AND4 (N1894, N1891, N1775, N1427, N180);
not NOT1 (N1895, N1878);
nor NOR2 (N1896, N1885, N1004);
and AND2 (N1897, N1893, N405);
and AND2 (N1898, N1866, N1081);
buf BUF1 (N1899, N1887);
and AND4 (N1900, N1897, N776, N107, N1437);
buf BUF1 (N1901, N1895);
buf BUF1 (N1902, N1892);
xor XOR2 (N1903, N1900, N1881);
buf BUF1 (N1904, N1880);
xor XOR2 (N1905, N1904, N1528);
nand NAND2 (N1906, N1899, N1384);
nand NAND4 (N1907, N1898, N885, N1069, N371);
xor XOR2 (N1908, N1889, N384);
and AND2 (N1909, N1883, N1075);
nor NOR2 (N1910, N1907, N649);
nand NAND2 (N1911, N1909, N143);
or OR3 (N1912, N1906, N1891, N1775);
nor NOR3 (N1913, N1894, N1378, N1223);
buf BUF1 (N1914, N1912);
not NOT1 (N1915, N1914);
xor XOR2 (N1916, N1910, N989);
and AND3 (N1917, N1911, N818, N1817);
nor NOR4 (N1918, N1903, N1664, N1161, N774);
and AND4 (N1919, N1918, N1104, N647, N460);
not NOT1 (N1920, N1908);
and AND2 (N1921, N1915, N1017);
nor NOR4 (N1922, N1902, N1920, N51, N1864);
buf BUF1 (N1923, N252);
not NOT1 (N1924, N1919);
nand NAND3 (N1925, N1923, N150, N115);
nor NOR3 (N1926, N1921, N402, N590);
and AND3 (N1927, N1926, N436, N1174);
not NOT1 (N1928, N1896);
and AND4 (N1929, N1922, N1089, N262, N830);
nor NOR3 (N1930, N1901, N1593, N1439);
nor NOR4 (N1931, N1930, N1442, N202, N1344);
and AND3 (N1932, N1917, N1064, N1019);
xor XOR2 (N1933, N1931, N989);
not NOT1 (N1934, N1932);
and AND4 (N1935, N1905, N1864, N1730, N254);
nor NOR4 (N1936, N1934, N194, N721, N1666);
buf BUF1 (N1937, N1928);
not NOT1 (N1938, N1924);
not NOT1 (N1939, N1925);
not NOT1 (N1940, N1939);
and AND3 (N1941, N1935, N1437, N1526);
and AND3 (N1942, N1938, N292, N1935);
and AND3 (N1943, N1916, N1377, N715);
nand NAND2 (N1944, N1943, N1622);
nor NOR4 (N1945, N1944, N36, N1669, N1785);
and AND4 (N1946, N1937, N667, N1527, N287);
and AND2 (N1947, N1941, N77);
nor NOR4 (N1948, N1933, N198, N328, N139);
and AND4 (N1949, N1940, N186, N1902, N1835);
and AND2 (N1950, N1949, N484);
nor NOR2 (N1951, N1945, N182);
nand NAND3 (N1952, N1948, N1828, N1615);
not NOT1 (N1953, N1913);
nor NOR3 (N1954, N1952, N686, N172);
buf BUF1 (N1955, N1950);
or OR3 (N1956, N1946, N610, N173);
xor XOR2 (N1957, N1951, N778);
or OR4 (N1958, N1955, N1578, N43, N1126);
not NOT1 (N1959, N1953);
xor XOR2 (N1960, N1958, N1820);
xor XOR2 (N1961, N1927, N1078);
buf BUF1 (N1962, N1954);
not NOT1 (N1963, N1936);
and AND4 (N1964, N1963, N416, N525, N458);
or OR3 (N1965, N1929, N1866, N1909);
xor XOR2 (N1966, N1964, N584);
nor NOR4 (N1967, N1942, N1545, N1711, N308);
or OR3 (N1968, N1961, N339, N723);
buf BUF1 (N1969, N1966);
or OR4 (N1970, N1962, N980, N1360, N1953);
nand NAND2 (N1971, N1959, N1297);
and AND2 (N1972, N1965, N1484);
not NOT1 (N1973, N1972);
buf BUF1 (N1974, N1969);
or OR2 (N1975, N1974, N352);
not NOT1 (N1976, N1956);
and AND3 (N1977, N1967, N10, N73);
xor XOR2 (N1978, N1973, N404);
nor NOR2 (N1979, N1960, N1074);
not NOT1 (N1980, N1979);
or OR2 (N1981, N1978, N1295);
nor NOR4 (N1982, N1977, N1140, N950, N1592);
nor NOR3 (N1983, N1957, N1404, N14);
not NOT1 (N1984, N1975);
and AND4 (N1985, N1947, N526, N1567, N32);
nor NOR3 (N1986, N1970, N535, N386);
and AND4 (N1987, N1982, N1005, N1754, N553);
nand NAND4 (N1988, N1968, N1815, N268, N1237);
buf BUF1 (N1989, N1971);
nor NOR2 (N1990, N1983, N1137);
and AND3 (N1991, N1988, N347, N1434);
and AND2 (N1992, N1985, N1473);
or OR4 (N1993, N1989, N964, N1905, N860);
nand NAND2 (N1994, N1987, N1521);
nor NOR3 (N1995, N1991, N1219, N887);
not NOT1 (N1996, N1994);
and AND3 (N1997, N1980, N1990, N921);
not NOT1 (N1998, N1859);
and AND3 (N1999, N1986, N606, N1239);
or OR3 (N2000, N1992, N184, N521);
not NOT1 (N2001, N1981);
or OR4 (N2002, N1998, N136, N1217, N9);
and AND3 (N2003, N1984, N535, N132);
or OR3 (N2004, N2001, N1880, N778);
or OR4 (N2005, N1995, N1403, N347, N1644);
not NOT1 (N2006, N1993);
not NOT1 (N2007, N2002);
nor NOR3 (N2008, N2007, N1792, N582);
nor NOR2 (N2009, N1996, N1584);
nor NOR3 (N2010, N2003, N575, N903);
and AND4 (N2011, N2004, N1828, N1488, N1571);
nand NAND4 (N2012, N2011, N1851, N1044, N1556);
and AND2 (N2013, N2009, N93);
not NOT1 (N2014, N2013);
and AND2 (N2015, N2000, N1209);
or OR2 (N2016, N2015, N656);
and AND3 (N2017, N2008, N821, N844);
buf BUF1 (N2018, N1999);
nand NAND4 (N2019, N2010, N1450, N236, N1892);
or OR4 (N2020, N2016, N355, N1073, N1378);
or OR3 (N2021, N2012, N1148, N1171);
xor XOR2 (N2022, N2017, N538);
buf BUF1 (N2023, N2019);
buf BUF1 (N2024, N2023);
or OR2 (N2025, N2006, N1793);
xor XOR2 (N2026, N2014, N1311);
not NOT1 (N2027, N2024);
nand NAND3 (N2028, N2021, N720, N1284);
buf BUF1 (N2029, N2028);
xor XOR2 (N2030, N2027, N80);
xor XOR2 (N2031, N2005, N831);
or OR3 (N2032, N2022, N263, N1929);
nor NOR2 (N2033, N2029, N509);
nor NOR2 (N2034, N2025, N1523);
buf BUF1 (N2035, N2034);
nand NAND4 (N2036, N1976, N448, N124, N1629);
nand NAND4 (N2037, N2026, N122, N816, N1407);
nand NAND2 (N2038, N1997, N1287);
or OR2 (N2039, N2036, N266);
and AND2 (N2040, N2035, N572);
xor XOR2 (N2041, N2038, N2039);
not NOT1 (N2042, N1384);
buf BUF1 (N2043, N2041);
nor NOR4 (N2044, N2033, N165, N327, N1678);
or OR4 (N2045, N2042, N959, N1539, N1458);
xor XOR2 (N2046, N2031, N1801);
nor NOR2 (N2047, N2037, N1551);
nor NOR4 (N2048, N2046, N1518, N1203, N80);
or OR4 (N2049, N2040, N1755, N169, N1961);
and AND2 (N2050, N2048, N1923);
or OR4 (N2051, N2049, N168, N142, N1603);
not NOT1 (N2052, N2044);
buf BUF1 (N2053, N2045);
nor NOR3 (N2054, N2047, N908, N298);
xor XOR2 (N2055, N2032, N1903);
nor NOR2 (N2056, N2051, N621);
and AND3 (N2057, N2050, N1736, N1539);
nand NAND3 (N2058, N2052, N1953, N421);
buf BUF1 (N2059, N2054);
buf BUF1 (N2060, N2057);
nand NAND4 (N2061, N2030, N1170, N1466, N1364);
not NOT1 (N2062, N2061);
buf BUF1 (N2063, N2055);
nand NAND2 (N2064, N2059, N2062);
nor NOR2 (N2065, N1339, N1451);
and AND2 (N2066, N2043, N348);
buf BUF1 (N2067, N2058);
nor NOR4 (N2068, N2053, N971, N344, N719);
xor XOR2 (N2069, N2056, N1057);
and AND3 (N2070, N2068, N436, N1957);
nor NOR2 (N2071, N2065, N1262);
or OR4 (N2072, N2069, N156, N1513, N1991);
buf BUF1 (N2073, N2060);
buf BUF1 (N2074, N2073);
xor XOR2 (N2075, N2067, N1172);
nand NAND2 (N2076, N2074, N223);
buf BUF1 (N2077, N2071);
not NOT1 (N2078, N2072);
or OR3 (N2079, N2076, N1087, N925);
or OR2 (N2080, N2077, N1803);
or OR3 (N2081, N2070, N1930, N499);
nor NOR4 (N2082, N2020, N96, N1644, N1462);
xor XOR2 (N2083, N2064, N2031);
nor NOR2 (N2084, N2080, N995);
and AND2 (N2085, N2081, N826);
not NOT1 (N2086, N2063);
not NOT1 (N2087, N2075);
nor NOR3 (N2088, N2083, N948, N2000);
not NOT1 (N2089, N2066);
and AND2 (N2090, N2078, N85);
not NOT1 (N2091, N2088);
buf BUF1 (N2092, N2084);
not NOT1 (N2093, N2087);
or OR4 (N2094, N2079, N933, N1150, N1402);
and AND2 (N2095, N2093, N1917);
xor XOR2 (N2096, N2091, N653);
and AND4 (N2097, N2094, N407, N297, N443);
and AND2 (N2098, N2018, N1402);
nand NAND2 (N2099, N2096, N1188);
or OR4 (N2100, N2092, N949, N515, N1680);
or OR2 (N2101, N2097, N1379);
nand NAND3 (N2102, N2099, N1494, N1365);
buf BUF1 (N2103, N2101);
nor NOR3 (N2104, N2095, N1148, N1906);
nand NAND2 (N2105, N2098, N1196);
and AND4 (N2106, N2090, N918, N1471, N1209);
or OR2 (N2107, N2085, N1099);
buf BUF1 (N2108, N2104);
not NOT1 (N2109, N2086);
buf BUF1 (N2110, N2106);
not NOT1 (N2111, N2107);
nor NOR3 (N2112, N2108, N104, N282);
nor NOR2 (N2113, N2111, N561);
and AND4 (N2114, N2105, N1448, N1545, N1667);
nor NOR2 (N2115, N2114, N1731);
and AND4 (N2116, N2103, N1491, N1583, N823);
nand NAND3 (N2117, N2112, N846, N1664);
and AND3 (N2118, N2082, N167, N1983);
or OR4 (N2119, N2100, N701, N34, N1761);
xor XOR2 (N2120, N2119, N381);
not NOT1 (N2121, N2110);
nor NOR4 (N2122, N2121, N1458, N876, N703);
nor NOR2 (N2123, N2122, N1297);
and AND4 (N2124, N2118, N1080, N677, N194);
xor XOR2 (N2125, N2115, N1533);
xor XOR2 (N2126, N2116, N1381);
xor XOR2 (N2127, N2117, N150);
and AND4 (N2128, N2089, N1389, N879, N1617);
nand NAND3 (N2129, N2124, N282, N1591);
xor XOR2 (N2130, N2125, N1652);
xor XOR2 (N2131, N2130, N1330);
xor XOR2 (N2132, N2126, N690);
not NOT1 (N2133, N2120);
and AND3 (N2134, N2109, N137, N2099);
buf BUF1 (N2135, N2113);
nor NOR4 (N2136, N2129, N1761, N1883, N153);
or OR3 (N2137, N2132, N633, N2058);
nor NOR3 (N2138, N2123, N1356, N1160);
nor NOR2 (N2139, N2102, N1594);
xor XOR2 (N2140, N2134, N438);
nand NAND2 (N2141, N2131, N459);
nor NOR4 (N2142, N2133, N1236, N1168, N1011);
nand NAND2 (N2143, N2138, N2128);
xor XOR2 (N2144, N1836, N699);
nor NOR2 (N2145, N2140, N1965);
nor NOR2 (N2146, N2142, N601);
and AND2 (N2147, N2145, N1664);
buf BUF1 (N2148, N2137);
buf BUF1 (N2149, N2135);
buf BUF1 (N2150, N2146);
and AND4 (N2151, N2139, N918, N833, N1026);
xor XOR2 (N2152, N2136, N2102);
or OR2 (N2153, N2143, N622);
buf BUF1 (N2154, N2148);
nor NOR4 (N2155, N2147, N1813, N1381, N1903);
or OR3 (N2156, N2151, N640, N908);
not NOT1 (N2157, N2150);
buf BUF1 (N2158, N2141);
or OR2 (N2159, N2158, N1359);
and AND2 (N2160, N2149, N1404);
buf BUF1 (N2161, N2159);
or OR4 (N2162, N2155, N22, N1185, N302);
not NOT1 (N2163, N2154);
buf BUF1 (N2164, N2156);
nand NAND2 (N2165, N2161, N1157);
not NOT1 (N2166, N2153);
xor XOR2 (N2167, N2127, N417);
nand NAND3 (N2168, N2164, N1036, N2079);
buf BUF1 (N2169, N2157);
nor NOR2 (N2170, N2168, N1087);
or OR3 (N2171, N2166, N11, N1253);
nor NOR4 (N2172, N2170, N669, N866, N1083);
or OR3 (N2173, N2160, N1362, N710);
nor NOR2 (N2174, N2172, N2112);
buf BUF1 (N2175, N2173);
xor XOR2 (N2176, N2167, N630);
buf BUF1 (N2177, N2169);
and AND4 (N2178, N2162, N2175, N1307, N934);
xor XOR2 (N2179, N2092, N1641);
or OR3 (N2180, N2174, N1053, N80);
nand NAND3 (N2181, N2178, N284, N1946);
not NOT1 (N2182, N2181);
nand NAND4 (N2183, N2177, N1948, N1254, N1861);
nor NOR4 (N2184, N2176, N747, N934, N1382);
not NOT1 (N2185, N2163);
not NOT1 (N2186, N2144);
not NOT1 (N2187, N2179);
buf BUF1 (N2188, N2186);
not NOT1 (N2189, N2165);
nor NOR4 (N2190, N2180, N398, N1276, N1030);
not NOT1 (N2191, N2183);
buf BUF1 (N2192, N2190);
or OR4 (N2193, N2191, N1172, N1645, N1675);
xor XOR2 (N2194, N2189, N445);
nand NAND2 (N2195, N2152, N1204);
nor NOR2 (N2196, N2187, N1829);
and AND4 (N2197, N2194, N843, N1706, N1398);
buf BUF1 (N2198, N2193);
nand NAND3 (N2199, N2192, N1299, N560);
nand NAND4 (N2200, N2197, N681, N1256, N2019);
nand NAND4 (N2201, N2182, N1543, N1365, N1517);
nor NOR3 (N2202, N2200, N700, N2195);
or OR2 (N2203, N1247, N1634);
or OR4 (N2204, N2185, N1364, N21, N513);
buf BUF1 (N2205, N2184);
nor NOR3 (N2206, N2171, N497, N1977);
xor XOR2 (N2207, N2205, N537);
buf BUF1 (N2208, N2203);
or OR3 (N2209, N2196, N801, N492);
buf BUF1 (N2210, N2188);
nand NAND2 (N2211, N2210, N388);
xor XOR2 (N2212, N2201, N536);
nor NOR2 (N2213, N2207, N1820);
buf BUF1 (N2214, N2209);
and AND3 (N2215, N2208, N1023, N1774);
buf BUF1 (N2216, N2198);
buf BUF1 (N2217, N2199);
not NOT1 (N2218, N2204);
not NOT1 (N2219, N2215);
nor NOR4 (N2220, N2218, N1229, N1276, N1142);
or OR3 (N2221, N2206, N198, N1921);
nor NOR4 (N2222, N2214, N1839, N1736, N720);
not NOT1 (N2223, N2217);
nand NAND2 (N2224, N2220, N1624);
not NOT1 (N2225, N2222);
or OR2 (N2226, N2216, N1169);
nand NAND4 (N2227, N2221, N827, N1785, N199);
xor XOR2 (N2228, N2219, N273);
and AND4 (N2229, N2227, N1807, N1663, N1800);
nor NOR4 (N2230, N2212, N2212, N1145, N1808);
xor XOR2 (N2231, N2225, N1761);
nand NAND4 (N2232, N2224, N276, N1116, N2158);
nand NAND3 (N2233, N2213, N516, N2143);
buf BUF1 (N2234, N2231);
nor NOR2 (N2235, N2234, N1888);
not NOT1 (N2236, N2211);
or OR3 (N2237, N2226, N1608, N460);
not NOT1 (N2238, N2232);
not NOT1 (N2239, N2236);
and AND4 (N2240, N2228, N1959, N2066, N1628);
and AND3 (N2241, N2239, N557, N1726);
nor NOR2 (N2242, N2235, N2042);
or OR4 (N2243, N2241, N489, N101, N1889);
nor NOR2 (N2244, N2230, N1909);
xor XOR2 (N2245, N2202, N372);
nand NAND2 (N2246, N2229, N514);
nor NOR2 (N2247, N2240, N549);
or OR3 (N2248, N2223, N1980, N284);
nand NAND2 (N2249, N2247, N2128);
buf BUF1 (N2250, N2238);
xor XOR2 (N2251, N2250, N2209);
and AND3 (N2252, N2233, N258, N150);
nor NOR2 (N2253, N2242, N1759);
nand NAND2 (N2254, N2245, N1899);
nor NOR2 (N2255, N2237, N1981);
nor NOR2 (N2256, N2249, N801);
or OR4 (N2257, N2254, N1913, N1446, N45);
or OR4 (N2258, N2248, N593, N1552, N1065);
not NOT1 (N2259, N2255);
or OR2 (N2260, N2244, N1087);
nor NOR3 (N2261, N2256, N333, N1114);
not NOT1 (N2262, N2258);
nand NAND3 (N2263, N2261, N366, N492);
xor XOR2 (N2264, N2263, N1652);
xor XOR2 (N2265, N2251, N720);
or OR3 (N2266, N2264, N309, N2193);
or OR3 (N2267, N2262, N1045, N514);
or OR2 (N2268, N2257, N1388);
nand NAND2 (N2269, N2265, N1922);
not NOT1 (N2270, N2259);
buf BUF1 (N2271, N2269);
not NOT1 (N2272, N2266);
and AND2 (N2273, N2243, N90);
or OR4 (N2274, N2252, N1127, N2178, N1203);
xor XOR2 (N2275, N2260, N407);
xor XOR2 (N2276, N2275, N746);
xor XOR2 (N2277, N2273, N210);
xor XOR2 (N2278, N2274, N1378);
and AND2 (N2279, N2271, N1318);
not NOT1 (N2280, N2279);
nand NAND2 (N2281, N2253, N623);
not NOT1 (N2282, N2281);
and AND4 (N2283, N2282, N711, N1983, N1389);
buf BUF1 (N2284, N2278);
not NOT1 (N2285, N2270);
not NOT1 (N2286, N2267);
or OR3 (N2287, N2268, N1328, N663);
not NOT1 (N2288, N2283);
nor NOR2 (N2289, N2276, N1507);
or OR4 (N2290, N2280, N2093, N1788, N1143);
not NOT1 (N2291, N2277);
xor XOR2 (N2292, N2285, N147);
buf BUF1 (N2293, N2292);
xor XOR2 (N2294, N2290, N199);
or OR4 (N2295, N2284, N1780, N1767, N554);
or OR2 (N2296, N2293, N1957);
not NOT1 (N2297, N2294);
or OR3 (N2298, N2272, N924, N1357);
not NOT1 (N2299, N2288);
nor NOR3 (N2300, N2298, N160, N1029);
not NOT1 (N2301, N2296);
nor NOR3 (N2302, N2301, N769, N2256);
xor XOR2 (N2303, N2286, N1914);
xor XOR2 (N2304, N2300, N2267);
nor NOR4 (N2305, N2303, N1794, N367, N148);
nand NAND2 (N2306, N2246, N1301);
xor XOR2 (N2307, N2304, N43);
and AND3 (N2308, N2306, N1375, N1903);
and AND2 (N2309, N2302, N1716);
xor XOR2 (N2310, N2309, N2099);
buf BUF1 (N2311, N2305);
not NOT1 (N2312, N2297);
nand NAND2 (N2313, N2289, N99);
and AND3 (N2314, N2295, N803, N1482);
nor NOR2 (N2315, N2313, N2028);
buf BUF1 (N2316, N2310);
buf BUF1 (N2317, N2287);
nand NAND3 (N2318, N2316, N963, N926);
nor NOR2 (N2319, N2291, N1842);
and AND3 (N2320, N2319, N610, N1082);
nor NOR2 (N2321, N2315, N1093);
buf BUF1 (N2322, N2318);
buf BUF1 (N2323, N2321);
xor XOR2 (N2324, N2322, N2262);
xor XOR2 (N2325, N2311, N242);
not NOT1 (N2326, N2317);
buf BUF1 (N2327, N2314);
not NOT1 (N2328, N2324);
buf BUF1 (N2329, N2328);
buf BUF1 (N2330, N2327);
not NOT1 (N2331, N2323);
nor NOR2 (N2332, N2312, N114);
nand NAND3 (N2333, N2308, N2180, N2263);
buf BUF1 (N2334, N2307);
xor XOR2 (N2335, N2325, N1946);
xor XOR2 (N2336, N2335, N1759);
nand NAND4 (N2337, N2326, N1425, N1066, N2093);
xor XOR2 (N2338, N2329, N1730);
buf BUF1 (N2339, N2320);
nand NAND3 (N2340, N2333, N2076, N1483);
and AND4 (N2341, N2339, N1187, N167, N2281);
and AND2 (N2342, N2338, N1847);
buf BUF1 (N2343, N2330);
nor NOR4 (N2344, N2343, N1979, N1479, N1908);
buf BUF1 (N2345, N2340);
xor XOR2 (N2346, N2299, N1736);
not NOT1 (N2347, N2332);
buf BUF1 (N2348, N2341);
nor NOR3 (N2349, N2342, N1554, N1113);
buf BUF1 (N2350, N2345);
or OR4 (N2351, N2349, N659, N2166, N1166);
or OR4 (N2352, N2337, N1655, N528, N847);
nor NOR4 (N2353, N2336, N2150, N1340, N289);
nand NAND4 (N2354, N2353, N753, N1798, N1328);
xor XOR2 (N2355, N2351, N1090);
or OR4 (N2356, N2348, N267, N2330, N504);
not NOT1 (N2357, N2352);
xor XOR2 (N2358, N2357, N427);
xor XOR2 (N2359, N2347, N449);
and AND2 (N2360, N2354, N308);
buf BUF1 (N2361, N2360);
or OR2 (N2362, N2334, N1514);
buf BUF1 (N2363, N2346);
buf BUF1 (N2364, N2358);
nand NAND4 (N2365, N2363, N727, N2170, N1973);
xor XOR2 (N2366, N2356, N1069);
buf BUF1 (N2367, N2331);
buf BUF1 (N2368, N2355);
and AND2 (N2369, N2364, N527);
nand NAND4 (N2370, N2366, N2217, N1011, N2177);
nor NOR3 (N2371, N2362, N335, N2147);
not NOT1 (N2372, N2371);
buf BUF1 (N2373, N2359);
xor XOR2 (N2374, N2373, N1889);
buf BUF1 (N2375, N2367);
nand NAND4 (N2376, N2361, N1771, N220, N866);
xor XOR2 (N2377, N2370, N2224);
buf BUF1 (N2378, N2376);
nor NOR2 (N2379, N2378, N1312);
buf BUF1 (N2380, N2377);
buf BUF1 (N2381, N2380);
buf BUF1 (N2382, N2369);
nand NAND3 (N2383, N2368, N599, N646);
not NOT1 (N2384, N2383);
nand NAND3 (N2385, N2384, N1608, N1653);
buf BUF1 (N2386, N2385);
buf BUF1 (N2387, N2350);
and AND4 (N2388, N2379, N957, N1874, N2165);
buf BUF1 (N2389, N2344);
buf BUF1 (N2390, N2365);
buf BUF1 (N2391, N2375);
and AND2 (N2392, N2391, N2132);
nand NAND4 (N2393, N2387, N990, N228, N1077);
or OR3 (N2394, N2386, N1657, N696);
buf BUF1 (N2395, N2389);
not NOT1 (N2396, N2388);
and AND4 (N2397, N2393, N1956, N865, N1962);
or OR2 (N2398, N2372, N156);
and AND3 (N2399, N2394, N821, N735);
nor NOR2 (N2400, N2392, N1611);
and AND3 (N2401, N2395, N1566, N1905);
and AND4 (N2402, N2396, N557, N703, N1495);
not NOT1 (N2403, N2399);
or OR3 (N2404, N2398, N744, N1741);
nor NOR2 (N2405, N2404, N396);
xor XOR2 (N2406, N2381, N997);
and AND2 (N2407, N2390, N1999);
buf BUF1 (N2408, N2397);
nor NOR3 (N2409, N2374, N2261, N2393);
xor XOR2 (N2410, N2409, N2087);
and AND3 (N2411, N2406, N832, N1536);
not NOT1 (N2412, N2401);
or OR4 (N2413, N2402, N677, N2147, N1004);
buf BUF1 (N2414, N2382);
buf BUF1 (N2415, N2407);
buf BUF1 (N2416, N2414);
nand NAND2 (N2417, N2412, N2167);
or OR2 (N2418, N2415, N10);
not NOT1 (N2419, N2410);
nor NOR4 (N2420, N2413, N2163, N1820, N1527);
nor NOR4 (N2421, N2403, N2124, N1067, N833);
xor XOR2 (N2422, N2417, N1107);
nor NOR3 (N2423, N2420, N187, N1731);
not NOT1 (N2424, N2416);
buf BUF1 (N2425, N2422);
nand NAND3 (N2426, N2423, N416, N1247);
xor XOR2 (N2427, N2419, N865);
not NOT1 (N2428, N2408);
nand NAND2 (N2429, N2400, N229);
buf BUF1 (N2430, N2405);
buf BUF1 (N2431, N2421);
buf BUF1 (N2432, N2431);
xor XOR2 (N2433, N2427, N2351);
buf BUF1 (N2434, N2428);
not NOT1 (N2435, N2429);
nand NAND3 (N2436, N2434, N451, N2146);
nand NAND4 (N2437, N2432, N1214, N2380, N613);
xor XOR2 (N2438, N2425, N1646);
or OR3 (N2439, N2418, N1340, N1163);
not NOT1 (N2440, N2433);
nor NOR4 (N2441, N2424, N1178, N463, N1845);
buf BUF1 (N2442, N2411);
not NOT1 (N2443, N2437);
buf BUF1 (N2444, N2442);
buf BUF1 (N2445, N2439);
or OR3 (N2446, N2444, N750, N237);
not NOT1 (N2447, N2445);
and AND2 (N2448, N2435, N1703);
nor NOR3 (N2449, N2446, N2273, N1463);
nand NAND2 (N2450, N2426, N1000);
nor NOR2 (N2451, N2449, N1032);
nor NOR4 (N2452, N2447, N514, N910, N1506);
xor XOR2 (N2453, N2438, N1979);
or OR2 (N2454, N2452, N1235);
xor XOR2 (N2455, N2443, N2031);
not NOT1 (N2456, N2450);
or OR2 (N2457, N2441, N133);
not NOT1 (N2458, N2451);
and AND4 (N2459, N2457, N960, N1012, N1511);
and AND3 (N2460, N2459, N209, N2009);
and AND2 (N2461, N2454, N1814);
buf BUF1 (N2462, N2430);
nor NOR4 (N2463, N2455, N148, N1471, N1389);
not NOT1 (N2464, N2456);
or OR3 (N2465, N2464, N285, N529);
xor XOR2 (N2466, N2448, N1301);
nor NOR2 (N2467, N2460, N2229);
xor XOR2 (N2468, N2467, N837);
and AND2 (N2469, N2440, N1819);
nand NAND4 (N2470, N2458, N605, N326, N1116);
nor NOR3 (N2471, N2465, N126, N2200);
not NOT1 (N2472, N2469);
not NOT1 (N2473, N2472);
or OR2 (N2474, N2466, N943);
or OR3 (N2475, N2436, N1580, N857);
or OR2 (N2476, N2463, N2116);
nand NAND2 (N2477, N2471, N578);
buf BUF1 (N2478, N2477);
or OR3 (N2479, N2474, N2215, N2377);
nand NAND3 (N2480, N2453, N213, N314);
nor NOR3 (N2481, N2461, N2257, N99);
and AND4 (N2482, N2480, N269, N864, N515);
and AND4 (N2483, N2482, N437, N2058, N9);
buf BUF1 (N2484, N2483);
and AND3 (N2485, N2479, N2351, N1919);
or OR3 (N2486, N2470, N743, N1922);
xor XOR2 (N2487, N2473, N2127);
nand NAND2 (N2488, N2481, N1291);
nand NAND3 (N2489, N2468, N732, N1474);
not NOT1 (N2490, N2462);
not NOT1 (N2491, N2478);
nor NOR2 (N2492, N2490, N1598);
not NOT1 (N2493, N2486);
xor XOR2 (N2494, N2492, N1901);
and AND4 (N2495, N2485, N1636, N160, N262);
or OR3 (N2496, N2491, N2119, N867);
nand NAND3 (N2497, N2495, N358, N677);
xor XOR2 (N2498, N2489, N1601);
or OR2 (N2499, N2476, N2002);
not NOT1 (N2500, N2499);
xor XOR2 (N2501, N2498, N767);
not NOT1 (N2502, N2488);
nand NAND2 (N2503, N2494, N1105);
and AND3 (N2504, N2487, N1743, N225);
xor XOR2 (N2505, N2484, N2341);
or OR3 (N2506, N2502, N76, N1955);
xor XOR2 (N2507, N2501, N486);
nor NOR4 (N2508, N2505, N589, N390, N742);
or OR4 (N2509, N2506, N641, N959, N1000);
or OR4 (N2510, N2508, N1655, N2404, N1128);
nand NAND3 (N2511, N2510, N8, N143);
or OR4 (N2512, N2500, N1549, N1244, N2375);
not NOT1 (N2513, N2512);
or OR4 (N2514, N2507, N1222, N1784, N904);
xor XOR2 (N2515, N2475, N453);
buf BUF1 (N2516, N2509);
nand NAND2 (N2517, N2515, N594);
nor NOR4 (N2518, N2504, N508, N2364, N1874);
nand NAND3 (N2519, N2513, N1698, N938);
buf BUF1 (N2520, N2503);
and AND3 (N2521, N2516, N990, N100);
nor NOR2 (N2522, N2520, N686);
nor NOR3 (N2523, N2497, N597, N1708);
buf BUF1 (N2524, N2518);
nor NOR3 (N2525, N2522, N1594, N2008);
xor XOR2 (N2526, N2511, N1250);
nor NOR4 (N2527, N2496, N2245, N2209, N972);
not NOT1 (N2528, N2493);
not NOT1 (N2529, N2525);
xor XOR2 (N2530, N2514, N2204);
or OR3 (N2531, N2517, N1825, N1771);
xor XOR2 (N2532, N2530, N1649);
xor XOR2 (N2533, N2532, N717);
nand NAND2 (N2534, N2519, N751);
and AND2 (N2535, N2529, N48);
nor NOR4 (N2536, N2523, N1021, N572, N1890);
nand NAND2 (N2537, N2531, N1989);
nand NAND4 (N2538, N2537, N2075, N2350, N627);
and AND2 (N2539, N2524, N471);
and AND4 (N2540, N2536, N949, N2458, N283);
not NOT1 (N2541, N2539);
not NOT1 (N2542, N2540);
xor XOR2 (N2543, N2533, N1960);
or OR4 (N2544, N2543, N1709, N1613, N1285);
and AND3 (N2545, N2534, N358, N2032);
buf BUF1 (N2546, N2535);
buf BUF1 (N2547, N2545);
nor NOR4 (N2548, N2547, N70, N2002, N1199);
buf BUF1 (N2549, N2544);
buf BUF1 (N2550, N2521);
nand NAND2 (N2551, N2549, N941);
buf BUF1 (N2552, N2526);
nand NAND3 (N2553, N2538, N791, N542);
nor NOR4 (N2554, N2546, N210, N1247, N1058);
buf BUF1 (N2555, N2528);
and AND4 (N2556, N2527, N190, N1068, N530);
buf BUF1 (N2557, N2550);
xor XOR2 (N2558, N2555, N882);
buf BUF1 (N2559, N2553);
and AND3 (N2560, N2554, N563, N2314);
buf BUF1 (N2561, N2557);
or OR4 (N2562, N2561, N1057, N1738, N1569);
not NOT1 (N2563, N2541);
nor NOR2 (N2564, N2542, N523);
xor XOR2 (N2565, N2564, N1457);
xor XOR2 (N2566, N2562, N282);
xor XOR2 (N2567, N2563, N1541);
xor XOR2 (N2568, N2551, N1789);
buf BUF1 (N2569, N2567);
buf BUF1 (N2570, N2566);
and AND3 (N2571, N2556, N2220, N1628);
and AND4 (N2572, N2548, N2296, N1454, N1094);
nor NOR4 (N2573, N2571, N2019, N1589, N174);
or OR4 (N2574, N2559, N1366, N959, N133);
buf BUF1 (N2575, N2569);
xor XOR2 (N2576, N2558, N653);
and AND4 (N2577, N2565, N763, N2364, N46);
nor NOR4 (N2578, N2552, N881, N851, N134);
nor NOR2 (N2579, N2568, N190);
buf BUF1 (N2580, N2575);
xor XOR2 (N2581, N2570, N1009);
and AND3 (N2582, N2574, N2087, N971);
buf BUF1 (N2583, N2579);
xor XOR2 (N2584, N2578, N1409);
xor XOR2 (N2585, N2560, N1113);
xor XOR2 (N2586, N2582, N1580);
buf BUF1 (N2587, N2581);
nor NOR4 (N2588, N2580, N1783, N1256, N2073);
or OR2 (N2589, N2588, N291);
nand NAND3 (N2590, N2585, N2516, N1997);
and AND2 (N2591, N2583, N1057);
xor XOR2 (N2592, N2587, N1244);
and AND3 (N2593, N2586, N515, N1219);
or OR3 (N2594, N2584, N1628, N1756);
or OR4 (N2595, N2594, N2574, N493, N1668);
xor XOR2 (N2596, N2589, N880);
or OR4 (N2597, N2595, N1963, N572, N268);
or OR4 (N2598, N2597, N31, N2408, N1927);
nor NOR4 (N2599, N2576, N1994, N541, N2149);
nand NAND2 (N2600, N2599, N1445);
nor NOR3 (N2601, N2591, N2049, N1617);
or OR4 (N2602, N2596, N2572, N1225, N379);
not NOT1 (N2603, N773);
buf BUF1 (N2604, N2598);
or OR2 (N2605, N2600, N1818);
and AND4 (N2606, N2601, N35, N602, N90);
or OR4 (N2607, N2603, N1790, N1195, N929);
xor XOR2 (N2608, N2592, N613);
not NOT1 (N2609, N2577);
nand NAND4 (N2610, N2604, N1236, N2543, N2082);
not NOT1 (N2611, N2606);
xor XOR2 (N2612, N2602, N1306);
not NOT1 (N2613, N2573);
buf BUF1 (N2614, N2593);
and AND3 (N2615, N2612, N2528, N331);
not NOT1 (N2616, N2615);
or OR3 (N2617, N2607, N2196, N1448);
xor XOR2 (N2618, N2613, N2117);
or OR3 (N2619, N2605, N1996, N543);
and AND4 (N2620, N2609, N107, N1360, N2312);
nor NOR3 (N2621, N2620, N273, N905);
or OR4 (N2622, N2611, N2365, N1031, N857);
or OR2 (N2623, N2616, N1936);
nor NOR4 (N2624, N2610, N2009, N1175, N1443);
buf BUF1 (N2625, N2617);
not NOT1 (N2626, N2590);
buf BUF1 (N2627, N2624);
not NOT1 (N2628, N2614);
and AND2 (N2629, N2628, N794);
nand NAND4 (N2630, N2626, N2465, N1687, N1402);
not NOT1 (N2631, N2608);
buf BUF1 (N2632, N2631);
xor XOR2 (N2633, N2630, N2177);
not NOT1 (N2634, N2619);
buf BUF1 (N2635, N2627);
xor XOR2 (N2636, N2625, N564);
and AND2 (N2637, N2629, N1273);
or OR4 (N2638, N2632, N1461, N599, N2608);
and AND3 (N2639, N2622, N345, N2366);
or OR2 (N2640, N2635, N2211);
or OR3 (N2641, N2618, N249, N802);
or OR4 (N2642, N2639, N784, N1509, N173);
xor XOR2 (N2643, N2640, N1318);
buf BUF1 (N2644, N2636);
xor XOR2 (N2645, N2621, N1061);
nor NOR4 (N2646, N2643, N1157, N2534, N1820);
or OR2 (N2647, N2645, N2059);
nand NAND4 (N2648, N2634, N78, N1229, N1650);
or OR2 (N2649, N2648, N184);
buf BUF1 (N2650, N2641);
and AND4 (N2651, N2650, N746, N1607, N2059);
xor XOR2 (N2652, N2637, N963);
buf BUF1 (N2653, N2633);
buf BUF1 (N2654, N2623);
and AND3 (N2655, N2644, N1609, N1855);
nand NAND4 (N2656, N2655, N1598, N2349, N874);
buf BUF1 (N2657, N2647);
not NOT1 (N2658, N2642);
nand NAND4 (N2659, N2652, N758, N275, N227);
nand NAND3 (N2660, N2654, N285, N1254);
xor XOR2 (N2661, N2656, N147);
xor XOR2 (N2662, N2658, N322);
nor NOR4 (N2663, N2661, N1003, N232, N1828);
nor NOR3 (N2664, N2662, N308, N1527);
not NOT1 (N2665, N2659);
xor XOR2 (N2666, N2649, N1425);
xor XOR2 (N2667, N2660, N1733);
or OR3 (N2668, N2665, N1804, N644);
and AND3 (N2669, N2638, N1652, N15);
nor NOR3 (N2670, N2653, N12, N1312);
and AND2 (N2671, N2667, N37);
nand NAND2 (N2672, N2666, N2652);
and AND2 (N2673, N2670, N2509);
nand NAND4 (N2674, N2657, N2265, N673, N531);
or OR2 (N2675, N2669, N1242);
nand NAND2 (N2676, N2672, N1858);
xor XOR2 (N2677, N2646, N680);
nor NOR4 (N2678, N2677, N690, N2157, N1864);
nand NAND4 (N2679, N2651, N1465, N2545, N435);
nand NAND2 (N2680, N2664, N783);
nor NOR3 (N2681, N2679, N15, N43);
and AND4 (N2682, N2680, N1181, N319, N965);
xor XOR2 (N2683, N2663, N1389);
and AND2 (N2684, N2676, N1614);
not NOT1 (N2685, N2684);
buf BUF1 (N2686, N2671);
and AND3 (N2687, N2681, N2624, N1669);
not NOT1 (N2688, N2678);
and AND2 (N2689, N2683, N2182);
nor NOR4 (N2690, N2689, N383, N1727, N625);
nand NAND4 (N2691, N2682, N2633, N2488, N2657);
nor NOR3 (N2692, N2685, N489, N1947);
nor NOR4 (N2693, N2686, N932, N934, N1825);
not NOT1 (N2694, N2675);
nor NOR3 (N2695, N2694, N405, N2443);
xor XOR2 (N2696, N2692, N1152);
nand NAND2 (N2697, N2696, N516);
or OR2 (N2698, N2668, N2585);
xor XOR2 (N2699, N2673, N2177);
buf BUF1 (N2700, N2693);
nand NAND2 (N2701, N2674, N1146);
buf BUF1 (N2702, N2695);
and AND2 (N2703, N2699, N1478);
and AND2 (N2704, N2698, N1047);
nor NOR2 (N2705, N2690, N1154);
and AND3 (N2706, N2705, N496, N944);
nand NAND2 (N2707, N2701, N1059);
buf BUF1 (N2708, N2687);
and AND3 (N2709, N2702, N222, N1812);
and AND3 (N2710, N2697, N889, N1634);
nand NAND3 (N2711, N2710, N436, N2002);
xor XOR2 (N2712, N2711, N126);
xor XOR2 (N2713, N2707, N149);
nand NAND3 (N2714, N2713, N1165, N591);
buf BUF1 (N2715, N2714);
buf BUF1 (N2716, N2691);
and AND3 (N2717, N2712, N493, N1767);
not NOT1 (N2718, N2704);
nor NOR4 (N2719, N2700, N1013, N2137, N1391);
nand NAND3 (N2720, N2703, N818, N1665);
buf BUF1 (N2721, N2720);
and AND2 (N2722, N2715, N99);
xor XOR2 (N2723, N2721, N461);
not NOT1 (N2724, N2706);
buf BUF1 (N2725, N2716);
xor XOR2 (N2726, N2725, N282);
nor NOR4 (N2727, N2719, N956, N737, N2415);
or OR2 (N2728, N2708, N2430);
and AND2 (N2729, N2722, N1596);
buf BUF1 (N2730, N2724);
not NOT1 (N2731, N2728);
nand NAND4 (N2732, N2729, N1787, N2456, N302);
not NOT1 (N2733, N2717);
not NOT1 (N2734, N2732);
and AND3 (N2735, N2723, N2200, N1721);
buf BUF1 (N2736, N2709);
buf BUF1 (N2737, N2736);
nor NOR2 (N2738, N2730, N922);
and AND2 (N2739, N2688, N8);
and AND4 (N2740, N2727, N684, N2044, N1511);
xor XOR2 (N2741, N2734, N1856);
nor NOR2 (N2742, N2735, N1396);
xor XOR2 (N2743, N2740, N938);
xor XOR2 (N2744, N2739, N1833);
nand NAND3 (N2745, N2741, N2082, N844);
xor XOR2 (N2746, N2743, N1982);
xor XOR2 (N2747, N2745, N1456);
not NOT1 (N2748, N2742);
and AND3 (N2749, N2748, N455, N1682);
not NOT1 (N2750, N2726);
not NOT1 (N2751, N2733);
and AND2 (N2752, N2744, N2312);
not NOT1 (N2753, N2750);
or OR4 (N2754, N2746, N1196, N831, N880);
and AND2 (N2755, N2738, N2304);
and AND3 (N2756, N2718, N1016, N2594);
nor NOR3 (N2757, N2747, N1438, N2693);
or OR3 (N2758, N2755, N1023, N916);
or OR4 (N2759, N2749, N579, N1333, N2290);
buf BUF1 (N2760, N2754);
or OR3 (N2761, N2753, N1197, N189);
and AND2 (N2762, N2761, N1095);
nor NOR2 (N2763, N2752, N2174);
nor NOR4 (N2764, N2760, N1800, N2209, N1386);
xor XOR2 (N2765, N2757, N295);
buf BUF1 (N2766, N2758);
xor XOR2 (N2767, N2763, N1105);
xor XOR2 (N2768, N2766, N1747);
not NOT1 (N2769, N2764);
xor XOR2 (N2770, N2751, N702);
not NOT1 (N2771, N2762);
not NOT1 (N2772, N2759);
nor NOR3 (N2773, N2768, N9, N1848);
not NOT1 (N2774, N2770);
xor XOR2 (N2775, N2767, N1078);
xor XOR2 (N2776, N2772, N2356);
nor NOR2 (N2777, N2774, N1649);
not NOT1 (N2778, N2775);
xor XOR2 (N2779, N2771, N854);
or OR3 (N2780, N2777, N2498, N1963);
or OR3 (N2781, N2765, N1305, N2307);
and AND2 (N2782, N2756, N1840);
xor XOR2 (N2783, N2776, N427);
not NOT1 (N2784, N2781);
nor NOR2 (N2785, N2783, N2564);
not NOT1 (N2786, N2780);
nand NAND2 (N2787, N2737, N2180);
buf BUF1 (N2788, N2784);
not NOT1 (N2789, N2787);
buf BUF1 (N2790, N2773);
buf BUF1 (N2791, N2779);
not NOT1 (N2792, N2789);
nor NOR2 (N2793, N2790, N717);
and AND3 (N2794, N2731, N202, N2124);
and AND2 (N2795, N2769, N677);
nor NOR3 (N2796, N2785, N362, N1631);
xor XOR2 (N2797, N2782, N36);
or OR4 (N2798, N2791, N1525, N1106, N1562);
or OR4 (N2799, N2794, N113, N2185, N609);
buf BUF1 (N2800, N2793);
or OR3 (N2801, N2792, N650, N2207);
buf BUF1 (N2802, N2800);
xor XOR2 (N2803, N2795, N1611);
and AND2 (N2804, N2799, N654);
nor NOR3 (N2805, N2786, N1534, N2544);
or OR4 (N2806, N2796, N2548, N1764, N1230);
buf BUF1 (N2807, N2804);
and AND4 (N2808, N2807, N858, N1666, N2507);
xor XOR2 (N2809, N2797, N183);
xor XOR2 (N2810, N2788, N977);
nand NAND4 (N2811, N2810, N1679, N2384, N1403);
and AND2 (N2812, N2798, N396);
or OR2 (N2813, N2806, N1723);
and AND4 (N2814, N2811, N2001, N1117, N1609);
nor NOR3 (N2815, N2778, N2678, N512);
xor XOR2 (N2816, N2809, N1301);
xor XOR2 (N2817, N2808, N1777);
buf BUF1 (N2818, N2814);
nor NOR4 (N2819, N2805, N1235, N1187, N865);
or OR2 (N2820, N2817, N774);
nor NOR2 (N2821, N2801, N1127);
xor XOR2 (N2822, N2815, N746);
and AND2 (N2823, N2812, N1012);
nand NAND4 (N2824, N2819, N2501, N2526, N2359);
and AND2 (N2825, N2813, N841);
nor NOR2 (N2826, N2818, N916);
and AND3 (N2827, N2802, N1729, N132);
buf BUF1 (N2828, N2824);
nor NOR3 (N2829, N2821, N627, N1050);
nand NAND2 (N2830, N2827, N1773);
xor XOR2 (N2831, N2820, N283);
nand NAND3 (N2832, N2829, N2588, N955);
not NOT1 (N2833, N2816);
not NOT1 (N2834, N2826);
buf BUF1 (N2835, N2823);
and AND4 (N2836, N2830, N2227, N2449, N5);
and AND3 (N2837, N2833, N538, N795);
and AND2 (N2838, N2835, N1441);
and AND3 (N2839, N2828, N300, N2605);
and AND3 (N2840, N2837, N2652, N1855);
not NOT1 (N2841, N2838);
or OR2 (N2842, N2834, N2071);
not NOT1 (N2843, N2836);
nor NOR2 (N2844, N2831, N1340);
xor XOR2 (N2845, N2841, N480);
xor XOR2 (N2846, N2803, N2278);
nand NAND4 (N2847, N2842, N1861, N2687, N2388);
buf BUF1 (N2848, N2822);
and AND3 (N2849, N2846, N413, N770);
buf BUF1 (N2850, N2825);
nand NAND4 (N2851, N2848, N2293, N1823, N2627);
nand NAND2 (N2852, N2843, N112);
xor XOR2 (N2853, N2852, N576);
nand NAND3 (N2854, N2839, N1030, N990);
nor NOR4 (N2855, N2847, N1913, N674, N2087);
xor XOR2 (N2856, N2840, N2374);
or OR4 (N2857, N2845, N2524, N833, N626);
or OR4 (N2858, N2857, N192, N112, N1769);
and AND4 (N2859, N2855, N1128, N1271, N1140);
and AND4 (N2860, N2849, N318, N560, N2674);
xor XOR2 (N2861, N2858, N1022);
xor XOR2 (N2862, N2844, N455);
or OR4 (N2863, N2860, N2379, N2635, N739);
xor XOR2 (N2864, N2863, N2271);
and AND2 (N2865, N2853, N2213);
or OR3 (N2866, N2859, N447, N470);
buf BUF1 (N2867, N2856);
not NOT1 (N2868, N2861);
xor XOR2 (N2869, N2867, N77);
nor NOR3 (N2870, N2854, N1693, N2058);
and AND3 (N2871, N2850, N153, N446);
not NOT1 (N2872, N2862);
or OR4 (N2873, N2832, N92, N1228, N2442);
and AND4 (N2874, N2869, N1508, N1766, N850);
buf BUF1 (N2875, N2874);
xor XOR2 (N2876, N2851, N2821);
not NOT1 (N2877, N2864);
not NOT1 (N2878, N2876);
or OR2 (N2879, N2872, N1157);
and AND4 (N2880, N2873, N2754, N1685, N2391);
not NOT1 (N2881, N2866);
not NOT1 (N2882, N2871);
buf BUF1 (N2883, N2870);
buf BUF1 (N2884, N2868);
and AND4 (N2885, N2883, N1630, N2017, N1545);
or OR3 (N2886, N2865, N87, N2499);
xor XOR2 (N2887, N2878, N2817);
and AND3 (N2888, N2879, N2634, N1717);
xor XOR2 (N2889, N2877, N2109);
or OR3 (N2890, N2888, N1934, N2085);
nand NAND4 (N2891, N2875, N636, N1550, N1637);
and AND4 (N2892, N2881, N2288, N2270, N556);
nor NOR3 (N2893, N2886, N424, N630);
not NOT1 (N2894, N2891);
not NOT1 (N2895, N2885);
xor XOR2 (N2896, N2890, N2670);
nor NOR2 (N2897, N2882, N2699);
nor NOR3 (N2898, N2895, N1419, N2585);
nor NOR4 (N2899, N2887, N2882, N1537, N2111);
not NOT1 (N2900, N2899);
and AND4 (N2901, N2898, N1105, N1858, N1670);
nand NAND3 (N2902, N2892, N2048, N1068);
nand NAND4 (N2903, N2894, N119, N2546, N1677);
not NOT1 (N2904, N2889);
nand NAND4 (N2905, N2884, N734, N1186, N1260);
not NOT1 (N2906, N2897);
nor NOR2 (N2907, N2902, N1647);
or OR3 (N2908, N2906, N2617, N701);
nor NOR3 (N2909, N2900, N2694, N110);
nor NOR3 (N2910, N2904, N1448, N2210);
or OR3 (N2911, N2893, N470, N2079);
or OR4 (N2912, N2880, N2017, N2066, N1911);
xor XOR2 (N2913, N2901, N2770);
and AND4 (N2914, N2910, N1524, N1456, N2676);
nand NAND3 (N2915, N2912, N1924, N38);
and AND2 (N2916, N2907, N54);
buf BUF1 (N2917, N2913);
not NOT1 (N2918, N2896);
or OR3 (N2919, N2911, N1627, N1637);
and AND4 (N2920, N2918, N496, N847, N1308);
xor XOR2 (N2921, N2920, N1013);
nor NOR4 (N2922, N2917, N2768, N179, N2788);
xor XOR2 (N2923, N2921, N1351);
xor XOR2 (N2924, N2903, N835);
and AND4 (N2925, N2916, N427, N506, N1237);
nor NOR4 (N2926, N2909, N2199, N2463, N1131);
nand NAND4 (N2927, N2914, N2023, N1341, N788);
nor NOR3 (N2928, N2927, N2819, N214);
nor NOR3 (N2929, N2905, N2077, N2288);
or OR2 (N2930, N2929, N215);
nand NAND2 (N2931, N2925, N2645);
buf BUF1 (N2932, N2908);
or OR2 (N2933, N2924, N930);
buf BUF1 (N2934, N2933);
buf BUF1 (N2935, N2919);
not NOT1 (N2936, N2932);
or OR3 (N2937, N2936, N1323, N2207);
buf BUF1 (N2938, N2937);
buf BUF1 (N2939, N2934);
nand NAND4 (N2940, N2926, N1346, N1295, N38);
buf BUF1 (N2941, N2923);
buf BUF1 (N2942, N2935);
nand NAND3 (N2943, N2939, N157, N200);
and AND3 (N2944, N2931, N2108, N1942);
and AND3 (N2945, N2941, N1483, N2575);
xor XOR2 (N2946, N2945, N2702);
and AND2 (N2947, N2942, N715);
not NOT1 (N2948, N2938);
nand NAND3 (N2949, N2922, N1291, N917);
or OR3 (N2950, N2928, N887, N406);
buf BUF1 (N2951, N2915);
nor NOR3 (N2952, N2930, N2097, N2606);
nor NOR3 (N2953, N2950, N1098, N2916);
nor NOR3 (N2954, N2953, N2483, N2558);
nand NAND2 (N2955, N2948, N2032);
nor NOR3 (N2956, N2949, N69, N1223);
nand NAND2 (N2957, N2955, N253);
buf BUF1 (N2958, N2954);
and AND2 (N2959, N2943, N2726);
nor NOR2 (N2960, N2959, N2400);
buf BUF1 (N2961, N2952);
buf BUF1 (N2962, N2951);
or OR4 (N2963, N2961, N2153, N2315, N2095);
nor NOR4 (N2964, N2957, N1503, N2308, N2931);
not NOT1 (N2965, N2960);
and AND2 (N2966, N2944, N152);
nand NAND3 (N2967, N2963, N136, N2520);
nand NAND3 (N2968, N2947, N2311, N333);
or OR2 (N2969, N2962, N784);
or OR4 (N2970, N2969, N413, N119, N2017);
nor NOR2 (N2971, N2966, N119);
nor NOR3 (N2972, N2958, N1839, N71);
and AND3 (N2973, N2956, N2056, N1668);
nor NOR2 (N2974, N2946, N2742);
not NOT1 (N2975, N2940);
xor XOR2 (N2976, N2965, N359);
buf BUF1 (N2977, N2972);
xor XOR2 (N2978, N2973, N1466);
not NOT1 (N2979, N2971);
not NOT1 (N2980, N2967);
and AND4 (N2981, N2968, N547, N466, N1406);
or OR2 (N2982, N2970, N1945);
nor NOR4 (N2983, N2974, N1299, N7, N2814);
or OR3 (N2984, N2978, N2720, N2107);
not NOT1 (N2985, N2979);
xor XOR2 (N2986, N2982, N245);
xor XOR2 (N2987, N2983, N2229);
buf BUF1 (N2988, N2984);
not NOT1 (N2989, N2977);
nand NAND3 (N2990, N2988, N2286, N1284);
xor XOR2 (N2991, N2981, N1647);
nor NOR2 (N2992, N2989, N2868);
and AND4 (N2993, N2986, N1648, N2048, N1099);
nand NAND2 (N2994, N2991, N2979);
xor XOR2 (N2995, N2964, N1354);
not NOT1 (N2996, N2990);
or OR2 (N2997, N2985, N2818);
and AND2 (N2998, N2997, N403);
nor NOR2 (N2999, N2995, N2122);
not NOT1 (N3000, N2998);
and AND3 (N3001, N2992, N1286, N1904);
buf BUF1 (N3002, N2975);
and AND4 (N3003, N3002, N151, N1344, N1956);
buf BUF1 (N3004, N3000);
xor XOR2 (N3005, N3001, N690);
buf BUF1 (N3006, N3004);
buf BUF1 (N3007, N2996);
not NOT1 (N3008, N3003);
not NOT1 (N3009, N2980);
and AND3 (N3010, N3008, N1345, N2976);
not NOT1 (N3011, N1563);
and AND4 (N3012, N3006, N2177, N2754, N2315);
nor NOR3 (N3013, N3007, N1854, N968);
and AND2 (N3014, N3010, N502);
nand NAND3 (N3015, N3013, N378, N581);
not NOT1 (N3016, N3005);
or OR4 (N3017, N3011, N1729, N1870, N2903);
xor XOR2 (N3018, N3016, N2720);
nor NOR2 (N3019, N3015, N2930);
buf BUF1 (N3020, N2999);
nand NAND4 (N3021, N2994, N54, N2460, N1541);
or OR4 (N3022, N2987, N528, N1805, N2406);
and AND3 (N3023, N3012, N1429, N2179);
nand NAND2 (N3024, N3023, N755);
or OR2 (N3025, N3021, N749);
and AND3 (N3026, N3020, N1238, N2089);
buf BUF1 (N3027, N3025);
buf BUF1 (N3028, N3017);
buf BUF1 (N3029, N3024);
and AND4 (N3030, N3019, N1933, N965, N1003);
buf BUF1 (N3031, N3029);
nand NAND3 (N3032, N3028, N2, N2334);
not NOT1 (N3033, N3009);
not NOT1 (N3034, N3022);
xor XOR2 (N3035, N3031, N29);
nand NAND4 (N3036, N3027, N2806, N1705, N2748);
buf BUF1 (N3037, N3026);
nor NOR2 (N3038, N3033, N523);
not NOT1 (N3039, N3030);
not NOT1 (N3040, N3039);
nand NAND4 (N3041, N3040, N1924, N954, N1673);
buf BUF1 (N3042, N3037);
nand NAND4 (N3043, N3036, N2018, N1716, N844);
and AND4 (N3044, N3018, N470, N2757, N1949);
nand NAND2 (N3045, N3044, N2146);
nand NAND3 (N3046, N3034, N1221, N2922);
nor NOR2 (N3047, N3032, N2696);
buf BUF1 (N3048, N3042);
nand NAND2 (N3049, N3041, N482);
and AND2 (N3050, N3014, N1510);
or OR2 (N3051, N3035, N2895);
nor NOR2 (N3052, N3048, N1791);
buf BUF1 (N3053, N3050);
nor NOR3 (N3054, N3047, N386, N2706);
and AND3 (N3055, N3046, N1363, N1950);
nand NAND4 (N3056, N3052, N2399, N2431, N597);
nor NOR4 (N3057, N2993, N73, N2913, N1773);
buf BUF1 (N3058, N3045);
and AND2 (N3059, N3056, N292);
xor XOR2 (N3060, N3051, N1008);
buf BUF1 (N3061, N3060);
xor XOR2 (N3062, N3057, N1371);
nand NAND4 (N3063, N3058, N408, N242, N2346);
and AND2 (N3064, N3038, N270);
and AND3 (N3065, N3053, N308, N766);
and AND2 (N3066, N3054, N1504);
buf BUF1 (N3067, N3066);
nand NAND2 (N3068, N3063, N3064);
or OR3 (N3069, N165, N1935, N2958);
nand NAND2 (N3070, N3059, N826);
xor XOR2 (N3071, N3055, N832);
not NOT1 (N3072, N3062);
or OR2 (N3073, N3068, N684);
and AND3 (N3074, N3072, N1992, N1656);
xor XOR2 (N3075, N3061, N881);
xor XOR2 (N3076, N3070, N507);
or OR2 (N3077, N3065, N1095);
nor NOR4 (N3078, N3074, N890, N428, N405);
nand NAND4 (N3079, N3043, N453, N2145, N653);
nor NOR3 (N3080, N3078, N852, N1520);
nand NAND2 (N3081, N3076, N950);
nor NOR2 (N3082, N3069, N1673);
xor XOR2 (N3083, N3075, N966);
nand NAND4 (N3084, N3082, N1813, N2244, N1957);
xor XOR2 (N3085, N3083, N2691);
and AND3 (N3086, N3067, N2974, N2449);
xor XOR2 (N3087, N3084, N1712);
or OR3 (N3088, N3087, N255, N929);
nor NOR2 (N3089, N3049, N1581);
or OR3 (N3090, N3085, N1342, N2789);
not NOT1 (N3091, N3071);
nor NOR4 (N3092, N3081, N760, N2362, N2467);
or OR3 (N3093, N3073, N1397, N1805);
buf BUF1 (N3094, N3091);
or OR4 (N3095, N3093, N1504, N1006, N2317);
buf BUF1 (N3096, N3086);
and AND3 (N3097, N3095, N1216, N2046);
nor NOR2 (N3098, N3088, N1348);
buf BUF1 (N3099, N3090);
buf BUF1 (N3100, N3080);
or OR3 (N3101, N3098, N953, N3037);
not NOT1 (N3102, N3099);
nand NAND3 (N3103, N3101, N1232, N3027);
nand NAND4 (N3104, N3079, N2377, N2244, N1531);
nor NOR4 (N3105, N3097, N2531, N1901, N2263);
and AND2 (N3106, N3094, N1507);
nand NAND2 (N3107, N3077, N1054);
or OR3 (N3108, N3105, N2164, N738);
buf BUF1 (N3109, N3107);
nand NAND3 (N3110, N3109, N3066, N1991);
or OR2 (N3111, N3092, N1022);
or OR4 (N3112, N3111, N1606, N2313, N3099);
or OR3 (N3113, N3106, N882, N1464);
not NOT1 (N3114, N3108);
nand NAND3 (N3115, N3112, N427, N2454);
buf BUF1 (N3116, N3115);
nor NOR2 (N3117, N3100, N2694);
or OR3 (N3118, N3116, N633, N2301);
not NOT1 (N3119, N3113);
nand NAND3 (N3120, N3117, N3100, N2260);
nor NOR3 (N3121, N3114, N83, N2407);
xor XOR2 (N3122, N3102, N2635);
buf BUF1 (N3123, N3104);
or OR2 (N3124, N3120, N865);
and AND2 (N3125, N3124, N2162);
not NOT1 (N3126, N3110);
and AND3 (N3127, N3126, N2941, N2408);
xor XOR2 (N3128, N3096, N3011);
xor XOR2 (N3129, N3103, N591);
not NOT1 (N3130, N3122);
or OR3 (N3131, N3128, N511, N1540);
or OR4 (N3132, N3121, N1025, N1305, N472);
nor NOR3 (N3133, N3089, N2383, N1376);
nand NAND3 (N3134, N3129, N41, N2812);
or OR2 (N3135, N3130, N1738);
and AND3 (N3136, N3133, N52, N2646);
nor NOR3 (N3137, N3134, N2249, N618);
buf BUF1 (N3138, N3136);
not NOT1 (N3139, N3138);
buf BUF1 (N3140, N3139);
xor XOR2 (N3141, N3125, N2568);
nor NOR3 (N3142, N3140, N2402, N500);
buf BUF1 (N3143, N3118);
buf BUF1 (N3144, N3142);
buf BUF1 (N3145, N3143);
nand NAND3 (N3146, N3131, N1073, N2096);
nor NOR4 (N3147, N3123, N1556, N2428, N1453);
xor XOR2 (N3148, N3132, N1513);
xor XOR2 (N3149, N3119, N1054);
or OR2 (N3150, N3137, N592);
not NOT1 (N3151, N3148);
or OR2 (N3152, N3135, N1972);
nor NOR4 (N3153, N3144, N15, N1438, N601);
or OR3 (N3154, N3153, N1212, N493);
or OR3 (N3155, N3145, N1174, N2416);
nand NAND3 (N3156, N3155, N867, N1359);
or OR2 (N3157, N3127, N48);
buf BUF1 (N3158, N3152);
not NOT1 (N3159, N3157);
nor NOR4 (N3160, N3146, N644, N892, N1956);
xor XOR2 (N3161, N3159, N2613);
and AND4 (N3162, N3161, N395, N1996, N2048);
xor XOR2 (N3163, N3149, N1975);
xor XOR2 (N3164, N3160, N2725);
nor NOR3 (N3165, N3141, N1201, N510);
not NOT1 (N3166, N3150);
or OR4 (N3167, N3165, N1535, N496, N2787);
and AND3 (N3168, N3163, N477, N3093);
nand NAND4 (N3169, N3162, N2341, N1519, N2903);
or OR2 (N3170, N3169, N1278);
nor NOR2 (N3171, N3168, N219);
xor XOR2 (N3172, N3170, N2169);
buf BUF1 (N3173, N3151);
not NOT1 (N3174, N3167);
or OR3 (N3175, N3164, N1113, N2872);
xor XOR2 (N3176, N3174, N1337);
not NOT1 (N3177, N3154);
nand NAND2 (N3178, N3173, N1766);
and AND4 (N3179, N3166, N2650, N438, N1599);
not NOT1 (N3180, N3158);
or OR4 (N3181, N3178, N521, N2194, N1415);
not NOT1 (N3182, N3177);
nand NAND2 (N3183, N3175, N1140);
nand NAND3 (N3184, N3180, N1390, N1199);
not NOT1 (N3185, N3156);
or OR4 (N3186, N3185, N2124, N1218, N2761);
not NOT1 (N3187, N3184);
nor NOR2 (N3188, N3183, N143);
nand NAND4 (N3189, N3179, N2978, N849, N846);
nand NAND2 (N3190, N3186, N2321);
xor XOR2 (N3191, N3182, N2938);
and AND2 (N3192, N3172, N1410);
xor XOR2 (N3193, N3176, N2510);
buf BUF1 (N3194, N3188);
not NOT1 (N3195, N3191);
not NOT1 (N3196, N3147);
and AND3 (N3197, N3181, N2006, N878);
nor NOR2 (N3198, N3171, N807);
and AND3 (N3199, N3197, N648, N493);
nand NAND4 (N3200, N3193, N1957, N3091, N2935);
xor XOR2 (N3201, N3194, N318);
nand NAND4 (N3202, N3198, N2823, N376, N166);
or OR3 (N3203, N3200, N2187, N629);
nand NAND2 (N3204, N3189, N495);
nand NAND3 (N3205, N3192, N3024, N1267);
nor NOR3 (N3206, N3199, N2857, N2208);
or OR4 (N3207, N3201, N2253, N149, N1263);
nor NOR4 (N3208, N3190, N1241, N1310, N2978);
xor XOR2 (N3209, N3204, N1747);
nor NOR4 (N3210, N3202, N2391, N2500, N3004);
not NOT1 (N3211, N3207);
buf BUF1 (N3212, N3211);
nand NAND3 (N3213, N3187, N1930, N809);
buf BUF1 (N3214, N3208);
and AND3 (N3215, N3195, N1054, N3083);
buf BUF1 (N3216, N3196);
buf BUF1 (N3217, N3210);
buf BUF1 (N3218, N3217);
and AND3 (N3219, N3209, N2479, N89);
or OR3 (N3220, N3212, N1267, N280);
buf BUF1 (N3221, N3205);
and AND2 (N3222, N3203, N369);
not NOT1 (N3223, N3218);
nand NAND3 (N3224, N3215, N720, N1097);
nand NAND3 (N3225, N3224, N633, N1112);
and AND2 (N3226, N3219, N1078);
not NOT1 (N3227, N3225);
or OR2 (N3228, N3226, N1081);
nor NOR4 (N3229, N3216, N2074, N2502, N1674);
or OR2 (N3230, N3222, N1038);
nand NAND2 (N3231, N3230, N198);
not NOT1 (N3232, N3223);
nor NOR2 (N3233, N3220, N2946);
and AND4 (N3234, N3229, N2819, N2466, N677);
buf BUF1 (N3235, N3227);
not NOT1 (N3236, N3234);
xor XOR2 (N3237, N3235, N2807);
and AND2 (N3238, N3231, N506);
nor NOR3 (N3239, N3221, N896, N204);
buf BUF1 (N3240, N3213);
buf BUF1 (N3241, N3238);
nand NAND3 (N3242, N3233, N2988, N2058);
xor XOR2 (N3243, N3237, N1227);
nand NAND2 (N3244, N3242, N396);
nor NOR4 (N3245, N3240, N1473, N399, N1414);
nor NOR2 (N3246, N3228, N2537);
buf BUF1 (N3247, N3239);
buf BUF1 (N3248, N3244);
not NOT1 (N3249, N3248);
and AND4 (N3250, N3206, N3012, N2237, N301);
not NOT1 (N3251, N3250);
not NOT1 (N3252, N3251);
and AND4 (N3253, N3232, N3, N1663, N43);
not NOT1 (N3254, N3245);
or OR2 (N3255, N3252, N397);
nand NAND3 (N3256, N3254, N1340, N1121);
not NOT1 (N3257, N3246);
nor NOR2 (N3258, N3241, N2751);
nor NOR3 (N3259, N3255, N1177, N2881);
buf BUF1 (N3260, N3236);
nand NAND3 (N3261, N3256, N654, N1774);
or OR2 (N3262, N3259, N2175);
not NOT1 (N3263, N3257);
xor XOR2 (N3264, N3263, N3167);
not NOT1 (N3265, N3247);
and AND4 (N3266, N3264, N1378, N498, N1721);
not NOT1 (N3267, N3266);
buf BUF1 (N3268, N3253);
or OR3 (N3269, N3243, N3082, N494);
xor XOR2 (N3270, N3261, N1107);
and AND4 (N3271, N3260, N2405, N1212, N826);
nor NOR3 (N3272, N3214, N2752, N2053);
xor XOR2 (N3273, N3249, N569);
and AND2 (N3274, N3269, N28);
nand NAND3 (N3275, N3273, N2819, N1276);
nand NAND4 (N3276, N3258, N613, N3023, N1591);
xor XOR2 (N3277, N3268, N1694);
xor XOR2 (N3278, N3277, N1473);
and AND3 (N3279, N3278, N105, N269);
not NOT1 (N3280, N3272);
nor NOR3 (N3281, N3267, N424, N670);
and AND3 (N3282, N3276, N1504, N156);
nand NAND4 (N3283, N3271, N1344, N2999, N2108);
xor XOR2 (N3284, N3274, N1174);
buf BUF1 (N3285, N3282);
buf BUF1 (N3286, N3270);
xor XOR2 (N3287, N3265, N1402);
nand NAND3 (N3288, N3283, N2212, N3204);
xor XOR2 (N3289, N3285, N1833);
nand NAND2 (N3290, N3279, N1205);
buf BUF1 (N3291, N3288);
not NOT1 (N3292, N3275);
xor XOR2 (N3293, N3287, N2609);
buf BUF1 (N3294, N3291);
not NOT1 (N3295, N3286);
nand NAND4 (N3296, N3292, N1792, N3168, N3211);
not NOT1 (N3297, N3281);
nand NAND3 (N3298, N3294, N921, N2575);
or OR2 (N3299, N3284, N1968);
or OR2 (N3300, N3295, N97);
nand NAND4 (N3301, N3299, N137, N849, N2123);
nand NAND4 (N3302, N3301, N343, N2431, N904);
xor XOR2 (N3303, N3298, N663);
or OR3 (N3304, N3297, N491, N2360);
not NOT1 (N3305, N3293);
and AND4 (N3306, N3289, N652, N3013, N1803);
not NOT1 (N3307, N3262);
buf BUF1 (N3308, N3306);
nand NAND2 (N3309, N3280, N956);
and AND4 (N3310, N3307, N420, N1915, N2051);
nor NOR2 (N3311, N3310, N2474);
buf BUF1 (N3312, N3305);
buf BUF1 (N3313, N3308);
buf BUF1 (N3314, N3313);
nor NOR2 (N3315, N3311, N1619);
or OR2 (N3316, N3304, N1301);
xor XOR2 (N3317, N3302, N2097);
or OR4 (N3318, N3303, N2294, N3222, N2073);
nand NAND2 (N3319, N3318, N1486);
buf BUF1 (N3320, N3309);
nor NOR3 (N3321, N3315, N424, N2420);
nor NOR4 (N3322, N3319, N3127, N1444, N2567);
or OR2 (N3323, N3290, N547);
nand NAND2 (N3324, N3322, N1345);
buf BUF1 (N3325, N3314);
nor NOR4 (N3326, N3312, N761, N619, N2806);
nor NOR4 (N3327, N3300, N1072, N2791, N2112);
buf BUF1 (N3328, N3323);
xor XOR2 (N3329, N3326, N1142);
or OR4 (N3330, N3329, N779, N62, N2293);
buf BUF1 (N3331, N3325);
not NOT1 (N3332, N3327);
not NOT1 (N3333, N3328);
or OR4 (N3334, N3296, N43, N2613, N2739);
nor NOR2 (N3335, N3331, N1536);
nor NOR4 (N3336, N3321, N2525, N383, N2731);
nor NOR2 (N3337, N3330, N2162);
buf BUF1 (N3338, N3334);
or OR2 (N3339, N3338, N3332);
and AND2 (N3340, N1259, N863);
nand NAND2 (N3341, N3339, N1891);
nor NOR2 (N3342, N3324, N2812);
or OR3 (N3343, N3341, N2324, N136);
or OR3 (N3344, N3320, N3202, N2052);
not NOT1 (N3345, N3333);
not NOT1 (N3346, N3345);
and AND2 (N3347, N3340, N2412);
and AND3 (N3348, N3336, N1459, N441);
and AND2 (N3349, N3347, N520);
nand NAND3 (N3350, N3346, N361, N679);
buf BUF1 (N3351, N3337);
not NOT1 (N3352, N3343);
nor NOR4 (N3353, N3351, N2878, N1599, N1654);
and AND2 (N3354, N3349, N2661);
not NOT1 (N3355, N3316);
and AND2 (N3356, N3317, N2248);
or OR2 (N3357, N3348, N1802);
not NOT1 (N3358, N3355);
xor XOR2 (N3359, N3354, N1810);
not NOT1 (N3360, N3335);
or OR3 (N3361, N3358, N1784, N547);
not NOT1 (N3362, N3353);
xor XOR2 (N3363, N3362, N2156);
nor NOR3 (N3364, N3356, N1658, N1773);
buf BUF1 (N3365, N3360);
and AND3 (N3366, N3352, N2594, N2583);
and AND3 (N3367, N3365, N2330, N1614);
buf BUF1 (N3368, N3363);
nor NOR2 (N3369, N3350, N548);
not NOT1 (N3370, N3368);
xor XOR2 (N3371, N3369, N371);
nor NOR3 (N3372, N3344, N1091, N2381);
and AND3 (N3373, N3372, N2295, N1745);
nor NOR4 (N3374, N3364, N1967, N2692, N3116);
xor XOR2 (N3375, N3366, N122);
nor NOR2 (N3376, N3370, N1817);
and AND3 (N3377, N3374, N2601, N2648);
buf BUF1 (N3378, N3359);
nor NOR2 (N3379, N3377, N2826);
buf BUF1 (N3380, N3376);
nand NAND3 (N3381, N3373, N2049, N1335);
nor NOR3 (N3382, N3378, N1265, N3199);
not NOT1 (N3383, N3361);
and AND2 (N3384, N3371, N3105);
buf BUF1 (N3385, N3384);
and AND4 (N3386, N3379, N3092, N1811, N1646);
or OR3 (N3387, N3386, N655, N999);
xor XOR2 (N3388, N3387, N705);
nor NOR4 (N3389, N3367, N3093, N1025, N2082);
or OR2 (N3390, N3389, N1079);
nor NOR4 (N3391, N3383, N2258, N3122, N1020);
xor XOR2 (N3392, N3391, N3238);
buf BUF1 (N3393, N3342);
and AND3 (N3394, N3357, N2754, N513);
xor XOR2 (N3395, N3375, N830);
nand NAND3 (N3396, N3381, N1807, N2157);
buf BUF1 (N3397, N3392);
buf BUF1 (N3398, N3393);
and AND3 (N3399, N3380, N554, N1326);
nor NOR4 (N3400, N3399, N3007, N3117, N194);
not NOT1 (N3401, N3400);
buf BUF1 (N3402, N3401);
buf BUF1 (N3403, N3385);
nand NAND2 (N3404, N3395, N1879);
or OR2 (N3405, N3382, N433);
xor XOR2 (N3406, N3405, N1071);
buf BUF1 (N3407, N3390);
nor NOR4 (N3408, N3404, N2975, N2974, N188);
and AND3 (N3409, N3408, N3054, N588);
not NOT1 (N3410, N3396);
nor NOR2 (N3411, N3403, N782);
xor XOR2 (N3412, N3407, N115);
not NOT1 (N3413, N3406);
or OR3 (N3414, N3388, N54, N654);
or OR2 (N3415, N3411, N1247);
or OR4 (N3416, N3409, N373, N858, N632);
not NOT1 (N3417, N3414);
buf BUF1 (N3418, N3402);
xor XOR2 (N3419, N3415, N3170);
and AND4 (N3420, N3418, N435, N2691, N3234);
or OR4 (N3421, N3394, N785, N2033, N3181);
or OR2 (N3422, N3420, N729);
xor XOR2 (N3423, N3413, N1323);
nor NOR2 (N3424, N3398, N1685);
or OR4 (N3425, N3423, N816, N2768, N1802);
nand NAND4 (N3426, N3416, N987, N3087, N226);
nand NAND3 (N3427, N3422, N711, N412);
not NOT1 (N3428, N3424);
and AND4 (N3429, N3425, N2241, N2556, N3085);
or OR2 (N3430, N3397, N1774);
and AND4 (N3431, N3428, N1795, N1463, N2201);
or OR3 (N3432, N3412, N595, N3014);
not NOT1 (N3433, N3430);
and AND4 (N3434, N3410, N1148, N2416, N1055);
or OR3 (N3435, N3419, N2860, N1861);
nor NOR2 (N3436, N3434, N2278);
not NOT1 (N3437, N3432);
not NOT1 (N3438, N3433);
or OR4 (N3439, N3429, N903, N1903, N2866);
nand NAND2 (N3440, N3439, N2216);
xor XOR2 (N3441, N3417, N666);
nand NAND3 (N3442, N3427, N1886, N1031);
nor NOR2 (N3443, N3421, N2500);
or OR2 (N3444, N3426, N2946);
nand NAND3 (N3445, N3438, N2032, N1593);
or OR3 (N3446, N3443, N1067, N1627);
nor NOR3 (N3447, N3437, N2422, N2176);
nand NAND2 (N3448, N3446, N1742);
and AND2 (N3449, N3447, N1508);
not NOT1 (N3450, N3431);
and AND3 (N3451, N3435, N2851, N2901);
nand NAND3 (N3452, N3440, N1607, N658);
nand NAND4 (N3453, N3444, N2113, N590, N50);
buf BUF1 (N3454, N3453);
not NOT1 (N3455, N3436);
xor XOR2 (N3456, N3452, N2965);
nor NOR4 (N3457, N3449, N3446, N1262, N3401);
or OR4 (N3458, N3456, N515, N1565, N1932);
buf BUF1 (N3459, N3450);
nor NOR2 (N3460, N3448, N1360);
and AND2 (N3461, N3451, N1537);
nand NAND2 (N3462, N3442, N1797);
nand NAND3 (N3463, N3461, N44, N2980);
and AND3 (N3464, N3460, N1361, N1761);
nor NOR4 (N3465, N3441, N1973, N1626, N895);
xor XOR2 (N3466, N3445, N2029);
buf BUF1 (N3467, N3463);
xor XOR2 (N3468, N3465, N356);
or OR3 (N3469, N3464, N293, N1389);
not NOT1 (N3470, N3454);
nand NAND3 (N3471, N3469, N1875, N2653);
nand NAND4 (N3472, N3455, N1631, N1554, N672);
nand NAND2 (N3473, N3466, N2887);
nor NOR2 (N3474, N3473, N1612);
or OR2 (N3475, N3471, N2114);
nand NAND2 (N3476, N3475, N3423);
nand NAND2 (N3477, N3472, N2097);
nand NAND2 (N3478, N3474, N3434);
xor XOR2 (N3479, N3468, N5);
and AND3 (N3480, N3476, N3030, N3312);
xor XOR2 (N3481, N3457, N1895);
nand NAND2 (N3482, N3462, N2651);
xor XOR2 (N3483, N3478, N173);
and AND2 (N3484, N3458, N832);
nor NOR3 (N3485, N3477, N2229, N1826);
nand NAND4 (N3486, N3470, N107, N2442, N1773);
or OR3 (N3487, N3482, N2931, N2704);
buf BUF1 (N3488, N3467);
or OR2 (N3489, N3481, N292);
buf BUF1 (N3490, N3483);
xor XOR2 (N3491, N3480, N1334);
xor XOR2 (N3492, N3486, N746);
or OR2 (N3493, N3484, N2719);
nor NOR3 (N3494, N3479, N63, N3207);
or OR2 (N3495, N3492, N1742);
or OR3 (N3496, N3490, N107, N446);
or OR3 (N3497, N3493, N1975, N2029);
nand NAND3 (N3498, N3497, N822, N2979);
or OR4 (N3499, N3485, N1030, N1097, N519);
or OR2 (N3500, N3487, N635);
not NOT1 (N3501, N3498);
nand NAND3 (N3502, N3488, N858, N1261);
buf BUF1 (N3503, N3499);
buf BUF1 (N3504, N3494);
buf BUF1 (N3505, N3489);
and AND4 (N3506, N3459, N3162, N1268, N1984);
not NOT1 (N3507, N3505);
and AND2 (N3508, N3502, N2448);
nor NOR3 (N3509, N3508, N2900, N2819);
and AND3 (N3510, N3507, N2609, N1412);
buf BUF1 (N3511, N3500);
nor NOR4 (N3512, N3495, N2444, N872, N166);
nand NAND3 (N3513, N3506, N2707, N2620);
and AND4 (N3514, N3491, N1799, N3425, N2557);
or OR2 (N3515, N3504, N203);
and AND3 (N3516, N3510, N2476, N1236);
nor NOR4 (N3517, N3509, N877, N682, N1058);
xor XOR2 (N3518, N3517, N3458);
or OR3 (N3519, N3516, N3048, N2845);
nand NAND3 (N3520, N3513, N2468, N3431);
buf BUF1 (N3521, N3496);
or OR3 (N3522, N3501, N1367, N3330);
or OR2 (N3523, N3521, N2543);
or OR3 (N3524, N3519, N1195, N198);
not NOT1 (N3525, N3515);
not NOT1 (N3526, N3503);
nand NAND2 (N3527, N3511, N1822);
and AND3 (N3528, N3525, N1825, N328);
nand NAND3 (N3529, N3514, N1569, N1694);
not NOT1 (N3530, N3524);
not NOT1 (N3531, N3530);
nand NAND4 (N3532, N3527, N1969, N3005, N2567);
nand NAND4 (N3533, N3526, N3283, N2305, N921);
and AND4 (N3534, N3523, N2303, N2874, N2061);
buf BUF1 (N3535, N3520);
and AND2 (N3536, N3534, N52);
and AND4 (N3537, N3529, N1298, N3129, N823);
buf BUF1 (N3538, N3528);
and AND2 (N3539, N3537, N1733);
and AND4 (N3540, N3532, N1358, N519, N3517);
and AND2 (N3541, N3540, N839);
buf BUF1 (N3542, N3536);
or OR4 (N3543, N3512, N1867, N2989, N1500);
xor XOR2 (N3544, N3535, N1316);
and AND4 (N3545, N3522, N1511, N2161, N1371);
not NOT1 (N3546, N3542);
xor XOR2 (N3547, N3545, N971);
and AND4 (N3548, N3533, N2440, N671, N2145);
and AND2 (N3549, N3546, N1098);
and AND3 (N3550, N3541, N2331, N1850);
nor NOR3 (N3551, N3538, N2328, N3440);
nand NAND2 (N3552, N3547, N2668);
not NOT1 (N3553, N3539);
or OR2 (N3554, N3548, N1679);
xor XOR2 (N3555, N3550, N210);
not NOT1 (N3556, N3553);
not NOT1 (N3557, N3554);
and AND4 (N3558, N3544, N2705, N1681, N38);
not NOT1 (N3559, N3543);
or OR3 (N3560, N3557, N3318, N2187);
and AND3 (N3561, N3555, N1882, N866);
and AND2 (N3562, N3551, N2457);
buf BUF1 (N3563, N3562);
nand NAND4 (N3564, N3561, N630, N2059, N3441);
nor NOR2 (N3565, N3559, N1549);
nor NOR4 (N3566, N3531, N1475, N716, N98);
or OR4 (N3567, N3552, N740, N3209, N3110);
nor NOR4 (N3568, N3560, N2678, N102, N2787);
and AND3 (N3569, N3549, N855, N1785);
and AND4 (N3570, N3567, N1361, N1632, N2091);
buf BUF1 (N3571, N3568);
and AND2 (N3572, N3558, N470);
xor XOR2 (N3573, N3572, N333);
xor XOR2 (N3574, N3518, N284);
not NOT1 (N3575, N3571);
and AND3 (N3576, N3556, N1431, N1659);
or OR4 (N3577, N3575, N2466, N380, N1087);
xor XOR2 (N3578, N3565, N1309);
buf BUF1 (N3579, N3576);
xor XOR2 (N3580, N3578, N725);
buf BUF1 (N3581, N3566);
and AND2 (N3582, N3573, N1373);
xor XOR2 (N3583, N3579, N539);
or OR4 (N3584, N3582, N3009, N2106, N3159);
not NOT1 (N3585, N3563);
buf BUF1 (N3586, N3569);
and AND2 (N3587, N3581, N2377);
buf BUF1 (N3588, N3577);
xor XOR2 (N3589, N3583, N834);
and AND2 (N3590, N3585, N914);
buf BUF1 (N3591, N3588);
nor NOR3 (N3592, N3580, N64, N3034);
or OR4 (N3593, N3574, N256, N684, N1680);
nand NAND2 (N3594, N3592, N1390);
xor XOR2 (N3595, N3584, N1028);
and AND2 (N3596, N3590, N498);
buf BUF1 (N3597, N3595);
xor XOR2 (N3598, N3589, N956);
and AND2 (N3599, N3586, N2170);
not NOT1 (N3600, N3564);
nor NOR4 (N3601, N3593, N3018, N2503, N3329);
nand NAND3 (N3602, N3570, N1978, N3112);
or OR3 (N3603, N3591, N2476, N3223);
nor NOR2 (N3604, N3587, N97);
not NOT1 (N3605, N3594);
or OR3 (N3606, N3598, N570, N479);
nor NOR4 (N3607, N3604, N1483, N78, N2040);
not NOT1 (N3608, N3603);
not NOT1 (N3609, N3597);
buf BUF1 (N3610, N3608);
buf BUF1 (N3611, N3606);
buf BUF1 (N3612, N3609);
not NOT1 (N3613, N3602);
and AND2 (N3614, N3611, N946);
nand NAND4 (N3615, N3614, N1336, N1820, N2762);
nor NOR4 (N3616, N3613, N1899, N1315, N2239);
buf BUF1 (N3617, N3605);
and AND4 (N3618, N3616, N1702, N1075, N1219);
xor XOR2 (N3619, N3615, N3493);
xor XOR2 (N3620, N3607, N2178);
and AND3 (N3621, N3601, N1075, N3211);
or OR4 (N3622, N3617, N309, N3205, N1179);
nand NAND4 (N3623, N3599, N2916, N2819, N2544);
or OR3 (N3624, N3618, N823, N2519);
not NOT1 (N3625, N3612);
buf BUF1 (N3626, N3619);
not NOT1 (N3627, N3623);
or OR4 (N3628, N3620, N3443, N501, N642);
xor XOR2 (N3629, N3610, N2013);
or OR4 (N3630, N3596, N160, N697, N2007);
not NOT1 (N3631, N3629);
or OR3 (N3632, N3627, N784, N171);
and AND3 (N3633, N3625, N329, N3415);
not NOT1 (N3634, N3628);
not NOT1 (N3635, N3624);
not NOT1 (N3636, N3634);
nand NAND3 (N3637, N3631, N201, N1443);
xor XOR2 (N3638, N3637, N52);
or OR2 (N3639, N3636, N2041);
and AND2 (N3640, N3600, N1492);
nand NAND2 (N3641, N3626, N2465);
not NOT1 (N3642, N3641);
nand NAND4 (N3643, N3635, N2298, N1544, N184);
and AND2 (N3644, N3632, N932);
nand NAND3 (N3645, N3638, N3096, N3420);
or OR3 (N3646, N3645, N2456, N3573);
nand NAND3 (N3647, N3644, N2865, N3629);
or OR4 (N3648, N3647, N3485, N1872, N3202);
not NOT1 (N3649, N3648);
nor NOR3 (N3650, N3621, N1319, N2505);
xor XOR2 (N3651, N3640, N512);
buf BUF1 (N3652, N3630);
xor XOR2 (N3653, N3650, N397);
or OR4 (N3654, N3651, N3424, N3555, N2270);
xor XOR2 (N3655, N3649, N1075);
nand NAND2 (N3656, N3652, N3101);
not NOT1 (N3657, N3639);
xor XOR2 (N3658, N3643, N1815);
not NOT1 (N3659, N3622);
nor NOR4 (N3660, N3658, N327, N2303, N753);
and AND2 (N3661, N3656, N656);
xor XOR2 (N3662, N3655, N1019);
nor NOR3 (N3663, N3653, N47, N267);
nand NAND2 (N3664, N3646, N1921);
and AND2 (N3665, N3663, N3494);
and AND4 (N3666, N3665, N1872, N589, N447);
not NOT1 (N3667, N3633);
xor XOR2 (N3668, N3661, N3441);
nor NOR3 (N3669, N3664, N589, N457);
not NOT1 (N3670, N3668);
or OR2 (N3671, N3666, N260);
nor NOR4 (N3672, N3667, N3552, N1388, N3583);
and AND3 (N3673, N3671, N681, N3349);
not NOT1 (N3674, N3659);
and AND3 (N3675, N3660, N2890, N2768);
xor XOR2 (N3676, N3654, N1232);
not NOT1 (N3677, N3670);
nor NOR3 (N3678, N3669, N3579, N3281);
not NOT1 (N3679, N3672);
nand NAND2 (N3680, N3679, N1429);
nor NOR4 (N3681, N3642, N1535, N1760, N506);
buf BUF1 (N3682, N3657);
and AND4 (N3683, N3673, N3496, N1020, N3646);
or OR4 (N3684, N3677, N765, N1658, N556);
and AND4 (N3685, N3675, N437, N25, N3361);
and AND2 (N3686, N3681, N1798);
nor NOR4 (N3687, N3682, N1871, N3664, N239);
xor XOR2 (N3688, N3662, N2108);
xor XOR2 (N3689, N3674, N2287);
not NOT1 (N3690, N3687);
buf BUF1 (N3691, N3684);
nor NOR3 (N3692, N3690, N1358, N3065);
nor NOR4 (N3693, N3680, N3285, N3561, N1651);
buf BUF1 (N3694, N3692);
and AND4 (N3695, N3683, N1222, N30, N3250);
buf BUF1 (N3696, N3693);
xor XOR2 (N3697, N3696, N2821);
nand NAND4 (N3698, N3688, N1963, N1303, N1435);
or OR2 (N3699, N3694, N286);
and AND4 (N3700, N3699, N936, N1872, N339);
nand NAND2 (N3701, N3697, N594);
not NOT1 (N3702, N3698);
nor NOR3 (N3703, N3689, N1, N1774);
nor NOR2 (N3704, N3702, N2085);
not NOT1 (N3705, N3676);
or OR3 (N3706, N3685, N2901, N1775);
not NOT1 (N3707, N3704);
or OR3 (N3708, N3701, N2992, N2947);
not NOT1 (N3709, N3678);
buf BUF1 (N3710, N3706);
not NOT1 (N3711, N3709);
xor XOR2 (N3712, N3707, N3404);
buf BUF1 (N3713, N3708);
not NOT1 (N3714, N3695);
or OR2 (N3715, N3711, N1261);
nor NOR4 (N3716, N3703, N986, N2663, N3135);
or OR2 (N3717, N3691, N3632);
nor NOR4 (N3718, N3713, N3505, N1776, N1098);
not NOT1 (N3719, N3700);
xor XOR2 (N3720, N3716, N3304);
xor XOR2 (N3721, N3712, N1242);
and AND3 (N3722, N3715, N15, N2733);
nand NAND2 (N3723, N3722, N1665);
nor NOR2 (N3724, N3718, N2649);
nor NOR3 (N3725, N3719, N1936, N858);
nor NOR4 (N3726, N3720, N1441, N1323, N2842);
xor XOR2 (N3727, N3721, N594);
nor NOR4 (N3728, N3717, N917, N2706, N117);
not NOT1 (N3729, N3723);
nor NOR2 (N3730, N3714, N2955);
buf BUF1 (N3731, N3705);
nor NOR4 (N3732, N3710, N3447, N2592, N458);
nor NOR4 (N3733, N3726, N1346, N439, N1446);
and AND2 (N3734, N3731, N1720);
buf BUF1 (N3735, N3725);
nand NAND3 (N3736, N3730, N1684, N241);
nand NAND4 (N3737, N3736, N685, N970, N3200);
buf BUF1 (N3738, N3686);
nor NOR3 (N3739, N3738, N1486, N3335);
and AND4 (N3740, N3728, N542, N2088, N3001);
and AND3 (N3741, N3734, N2357, N244);
or OR4 (N3742, N3739, N2560, N24, N2287);
or OR4 (N3743, N3740, N162, N3057, N2072);
and AND2 (N3744, N3724, N2641);
nor NOR2 (N3745, N3742, N644);
xor XOR2 (N3746, N3743, N2680);
xor XOR2 (N3747, N3745, N3355);
buf BUF1 (N3748, N3746);
nand NAND3 (N3749, N3741, N1094, N2184);
and AND2 (N3750, N3748, N63);
and AND2 (N3751, N3729, N3500);
nand NAND3 (N3752, N3747, N3669, N2009);
or OR2 (N3753, N3751, N1178);
nor NOR3 (N3754, N3737, N1234, N308);
buf BUF1 (N3755, N3733);
buf BUF1 (N3756, N3735);
buf BUF1 (N3757, N3755);
not NOT1 (N3758, N3732);
or OR3 (N3759, N3752, N214, N2911);
xor XOR2 (N3760, N3756, N2953);
or OR3 (N3761, N3759, N2136, N1917);
and AND2 (N3762, N3757, N3282);
buf BUF1 (N3763, N3727);
nand NAND3 (N3764, N3762, N3123, N471);
not NOT1 (N3765, N3749);
and AND3 (N3766, N3763, N939, N1603);
and AND2 (N3767, N3764, N3443);
or OR4 (N3768, N3750, N1862, N987, N2882);
buf BUF1 (N3769, N3761);
buf BUF1 (N3770, N3758);
buf BUF1 (N3771, N3765);
buf BUF1 (N3772, N3769);
or OR2 (N3773, N3771, N666);
or OR2 (N3774, N3760, N2590);
nand NAND3 (N3775, N3744, N2464, N557);
nor NOR2 (N3776, N3753, N2941);
nor NOR3 (N3777, N3767, N2382, N2708);
xor XOR2 (N3778, N3774, N1912);
or OR4 (N3779, N3775, N2201, N1460, N1032);
buf BUF1 (N3780, N3772);
nor NOR4 (N3781, N3776, N4, N2041, N1056);
and AND4 (N3782, N3781, N3570, N2791, N283);
nor NOR2 (N3783, N3780, N265);
or OR3 (N3784, N3754, N1468, N2535);
nand NAND4 (N3785, N3782, N60, N2022, N721);
not NOT1 (N3786, N3766);
nor NOR4 (N3787, N3777, N1581, N2679, N2795);
xor XOR2 (N3788, N3778, N1445);
and AND3 (N3789, N3786, N2233, N3441);
not NOT1 (N3790, N3783);
nor NOR4 (N3791, N3789, N3223, N2893, N1583);
xor XOR2 (N3792, N3790, N3380);
or OR4 (N3793, N3784, N3423, N506, N3641);
xor XOR2 (N3794, N3773, N2898);
xor XOR2 (N3795, N3770, N501);
not NOT1 (N3796, N3787);
nand NAND4 (N3797, N3779, N636, N2577, N2030);
or OR2 (N3798, N3785, N3642);
not NOT1 (N3799, N3797);
xor XOR2 (N3800, N3768, N2281);
nand NAND4 (N3801, N3794, N905, N3096, N3761);
and AND4 (N3802, N3800, N3644, N378, N2128);
xor XOR2 (N3803, N3792, N761);
not NOT1 (N3804, N3796);
buf BUF1 (N3805, N3788);
and AND4 (N3806, N3798, N3110, N1664, N139);
buf BUF1 (N3807, N3805);
buf BUF1 (N3808, N3806);
nand NAND4 (N3809, N3791, N2900, N2722, N941);
xor XOR2 (N3810, N3804, N3648);
buf BUF1 (N3811, N3809);
or OR4 (N3812, N3811, N1479, N2391, N46);
and AND2 (N3813, N3807, N3707);
or OR3 (N3814, N3803, N566, N2212);
not NOT1 (N3815, N3814);
or OR3 (N3816, N3795, N2476, N1513);
or OR4 (N3817, N3812, N735, N1175, N1187);
not NOT1 (N3818, N3813);
nand NAND3 (N3819, N3816, N270, N164);
buf BUF1 (N3820, N3810);
or OR4 (N3821, N3815, N2277, N2703, N935);
not NOT1 (N3822, N3793);
and AND2 (N3823, N3818, N1464);
buf BUF1 (N3824, N3799);
xor XOR2 (N3825, N3801, N3465);
and AND3 (N3826, N3822, N1786, N941);
and AND3 (N3827, N3802, N1891, N3475);
and AND4 (N3828, N3808, N1453, N3753, N1812);
nand NAND4 (N3829, N3827, N1112, N2804, N3264);
nor NOR4 (N3830, N3826, N855, N625, N2926);
not NOT1 (N3831, N3830);
buf BUF1 (N3832, N3817);
xor XOR2 (N3833, N3825, N3301);
buf BUF1 (N3834, N3823);
xor XOR2 (N3835, N3829, N1085);
nor NOR4 (N3836, N3828, N1515, N3343, N2469);
buf BUF1 (N3837, N3824);
xor XOR2 (N3838, N3820, N3701);
or OR2 (N3839, N3833, N706);
nand NAND2 (N3840, N3834, N2992);
nor NOR4 (N3841, N3839, N2084, N683, N732);
xor XOR2 (N3842, N3831, N2094);
nor NOR2 (N3843, N3837, N2984);
not NOT1 (N3844, N3841);
and AND2 (N3845, N3843, N3696);
not NOT1 (N3846, N3845);
nor NOR3 (N3847, N3844, N3744, N3142);
or OR3 (N3848, N3842, N1078, N3572);
not NOT1 (N3849, N3821);
and AND3 (N3850, N3832, N1909, N1406);
or OR4 (N3851, N3847, N947, N1443, N1380);
nor NOR4 (N3852, N3819, N902, N185, N2830);
not NOT1 (N3853, N3851);
nor NOR2 (N3854, N3850, N1660);
and AND3 (N3855, N3835, N514, N988);
not NOT1 (N3856, N3846);
nand NAND2 (N3857, N3854, N2457);
or OR2 (N3858, N3852, N1744);
xor XOR2 (N3859, N3848, N2053);
and AND4 (N3860, N3853, N2246, N2054, N3539);
or OR2 (N3861, N3856, N1569);
nor NOR3 (N3862, N3861, N603, N1782);
buf BUF1 (N3863, N3840);
not NOT1 (N3864, N3838);
nor NOR2 (N3865, N3863, N1552);
buf BUF1 (N3866, N3858);
buf BUF1 (N3867, N3860);
buf BUF1 (N3868, N3857);
nor NOR3 (N3869, N3862, N2549, N3726);
or OR2 (N3870, N3865, N207);
and AND2 (N3871, N3870, N1706);
nor NOR2 (N3872, N3859, N2574);
nor NOR3 (N3873, N3872, N3790, N1583);
nor NOR2 (N3874, N3871, N3469);
nor NOR3 (N3875, N3864, N2358, N2163);
nand NAND4 (N3876, N3874, N2101, N2956, N1033);
and AND3 (N3877, N3876, N1721, N769);
xor XOR2 (N3878, N3869, N588);
nor NOR4 (N3879, N3868, N3510, N3318, N2161);
and AND3 (N3880, N3875, N3006, N1527);
xor XOR2 (N3881, N3855, N2452);
not NOT1 (N3882, N3877);
or OR4 (N3883, N3880, N287, N984, N697);
nor NOR2 (N3884, N3836, N1383);
xor XOR2 (N3885, N3867, N3777);
nor NOR4 (N3886, N3849, N1460, N2922, N466);
nand NAND3 (N3887, N3883, N712, N2776);
not NOT1 (N3888, N3882);
or OR4 (N3889, N3873, N520, N1185, N2082);
nor NOR2 (N3890, N3887, N455);
not NOT1 (N3891, N3885);
nor NOR4 (N3892, N3866, N882, N224, N426);
nor NOR2 (N3893, N3891, N223);
xor XOR2 (N3894, N3881, N3090);
nor NOR2 (N3895, N3888, N2487);
buf BUF1 (N3896, N3879);
and AND4 (N3897, N3892, N3541, N1267, N3780);
or OR2 (N3898, N3884, N3281);
xor XOR2 (N3899, N3886, N3351);
or OR2 (N3900, N3894, N2500);
or OR2 (N3901, N3900, N3774);
or OR2 (N3902, N3889, N118);
not NOT1 (N3903, N3897);
nand NAND4 (N3904, N3899, N2139, N1844, N3468);
and AND2 (N3905, N3903, N1213);
buf BUF1 (N3906, N3895);
or OR3 (N3907, N3890, N1945, N1545);
buf BUF1 (N3908, N3905);
and AND2 (N3909, N3901, N3425);
buf BUF1 (N3910, N3878);
xor XOR2 (N3911, N3898, N2229);
nand NAND4 (N3912, N3910, N2055, N3433, N2019);
not NOT1 (N3913, N3908);
buf BUF1 (N3914, N3893);
and AND4 (N3915, N3914, N2538, N2992, N2686);
or OR4 (N3916, N3915, N2116, N2616, N2366);
nand NAND2 (N3917, N3896, N1290);
or OR3 (N3918, N3913, N675, N2137);
nand NAND3 (N3919, N3912, N3777, N953);
nor NOR4 (N3920, N3907, N376, N1722, N2413);
and AND3 (N3921, N3909, N3022, N2580);
and AND3 (N3922, N3917, N1647, N776);
not NOT1 (N3923, N3906);
not NOT1 (N3924, N3923);
or OR4 (N3925, N3920, N770, N2897, N3323);
not NOT1 (N3926, N3904);
not NOT1 (N3927, N3916);
nor NOR2 (N3928, N3921, N3054);
nand NAND3 (N3929, N3927, N3697, N1887);
nor NOR4 (N3930, N3918, N1649, N571, N479);
and AND2 (N3931, N3929, N2821);
nor NOR3 (N3932, N3930, N1144, N2505);
or OR4 (N3933, N3931, N1376, N2480, N2078);
not NOT1 (N3934, N3926);
and AND2 (N3935, N3911, N2392);
or OR2 (N3936, N3902, N3806);
xor XOR2 (N3937, N3933, N41);
and AND4 (N3938, N3937, N87, N199, N2997);
and AND4 (N3939, N3922, N3906, N1708, N2068);
not NOT1 (N3940, N3928);
and AND4 (N3941, N3925, N1136, N693, N2331);
not NOT1 (N3942, N3924);
not NOT1 (N3943, N3932);
or OR3 (N3944, N3943, N1990, N2160);
nand NAND2 (N3945, N3938, N1101);
not NOT1 (N3946, N3942);
nand NAND3 (N3947, N3939, N3853, N1847);
or OR2 (N3948, N3945, N3531);
and AND3 (N3949, N3941, N1091, N699);
not NOT1 (N3950, N3947);
nand NAND2 (N3951, N3944, N2441);
buf BUF1 (N3952, N3919);
not NOT1 (N3953, N3952);
or OR4 (N3954, N3949, N3691, N2621, N1780);
not NOT1 (N3955, N3954);
xor XOR2 (N3956, N3953, N579);
not NOT1 (N3957, N3948);
nor NOR4 (N3958, N3957, N2034, N2118, N2950);
not NOT1 (N3959, N3955);
and AND4 (N3960, N3946, N1566, N3449, N472);
buf BUF1 (N3961, N3935);
nor NOR2 (N3962, N3951, N2417);
and AND3 (N3963, N3959, N2924, N2129);
nor NOR4 (N3964, N3956, N1946, N2347, N3110);
and AND3 (N3965, N3934, N3125, N1742);
or OR4 (N3966, N3940, N2761, N3540, N2188);
buf BUF1 (N3967, N3936);
xor XOR2 (N3968, N3966, N3337);
buf BUF1 (N3969, N3965);
nand NAND2 (N3970, N3958, N3685);
nand NAND3 (N3971, N3970, N473, N2738);
not NOT1 (N3972, N3968);
or OR2 (N3973, N3963, N2237);
or OR4 (N3974, N3969, N2199, N1816, N167);
nor NOR4 (N3975, N3962, N2194, N2499, N317);
xor XOR2 (N3976, N3964, N1697);
nor NOR2 (N3977, N3961, N3414);
not NOT1 (N3978, N3977);
xor XOR2 (N3979, N3967, N76);
nand NAND3 (N3980, N3972, N3435, N608);
nor NOR3 (N3981, N3978, N134, N2527);
not NOT1 (N3982, N3981);
nand NAND3 (N3983, N3950, N20, N127);
buf BUF1 (N3984, N3974);
buf BUF1 (N3985, N3973);
nor NOR3 (N3986, N3984, N495, N3385);
or OR3 (N3987, N3971, N1345, N1009);
buf BUF1 (N3988, N3983);
or OR4 (N3989, N3986, N1210, N2927, N320);
nor NOR4 (N3990, N3960, N2369, N3898, N1251);
xor XOR2 (N3991, N3988, N2314);
nand NAND4 (N3992, N3987, N3871, N2173, N333);
or OR4 (N3993, N3992, N837, N2719, N1783);
and AND4 (N3994, N3976, N154, N1700, N1841);
nand NAND3 (N3995, N3979, N1685, N251);
not NOT1 (N3996, N3990);
or OR3 (N3997, N3980, N570, N547);
or OR4 (N3998, N3994, N1510, N2388, N361);
xor XOR2 (N3999, N3993, N1219);
and AND3 (N4000, N3982, N1693, N3020);
and AND3 (N4001, N3975, N3130, N2988);
not NOT1 (N4002, N3995);
buf BUF1 (N4003, N3996);
and AND4 (N4004, N4000, N2004, N1491, N2151);
nand NAND3 (N4005, N3989, N3421, N3042);
or OR3 (N4006, N4003, N1909, N2427);
or OR3 (N4007, N3985, N1865, N2219);
and AND2 (N4008, N4002, N3549);
buf BUF1 (N4009, N4007);
nand NAND4 (N4010, N4001, N2, N1128, N1384);
and AND2 (N4011, N4008, N1057);
nand NAND2 (N4012, N3997, N4003);
xor XOR2 (N4013, N4009, N2020);
or OR2 (N4014, N3991, N2691);
nor NOR4 (N4015, N4004, N1720, N2929, N1265);
xor XOR2 (N4016, N4005, N138);
buf BUF1 (N4017, N4010);
nor NOR2 (N4018, N4015, N1781);
or OR3 (N4019, N4013, N3319, N458);
or OR2 (N4020, N4006, N385);
and AND3 (N4021, N4012, N3298, N3471);
and AND4 (N4022, N4014, N1565, N2764, N2302);
buf BUF1 (N4023, N4017);
and AND2 (N4024, N4023, N2251);
xor XOR2 (N4025, N4021, N3142);
nand NAND3 (N4026, N3999, N1712, N2443);
nand NAND2 (N4027, N3998, N4025);
and AND3 (N4028, N2153, N1782, N2671);
or OR4 (N4029, N4028, N1039, N591, N1108);
nand NAND2 (N4030, N4024, N3004);
nand NAND2 (N4031, N4020, N823);
buf BUF1 (N4032, N4029);
buf BUF1 (N4033, N4018);
nand NAND3 (N4034, N4027, N1732, N274);
not NOT1 (N4035, N4022);
xor XOR2 (N4036, N4035, N2063);
or OR3 (N4037, N4019, N1556, N2121);
buf BUF1 (N4038, N4011);
xor XOR2 (N4039, N4038, N1664);
not NOT1 (N4040, N4016);
nand NAND4 (N4041, N4036, N769, N1837, N1798);
or OR3 (N4042, N4041, N1190, N3646);
buf BUF1 (N4043, N4037);
nand NAND4 (N4044, N4032, N2570, N3232, N300);
nor NOR4 (N4045, N4039, N1349, N2942, N3304);
buf BUF1 (N4046, N4033);
and AND4 (N4047, N4031, N472, N3098, N3506);
nor NOR2 (N4048, N4040, N1538);
buf BUF1 (N4049, N4030);
nor NOR2 (N4050, N4046, N2724);
or OR2 (N4051, N4026, N3365);
buf BUF1 (N4052, N4049);
or OR4 (N4053, N4044, N151, N3773, N1089);
buf BUF1 (N4054, N4042);
and AND2 (N4055, N4043, N2790);
or OR2 (N4056, N4045, N1721);
buf BUF1 (N4057, N4054);
and AND2 (N4058, N4052, N3684);
buf BUF1 (N4059, N4056);
buf BUF1 (N4060, N4059);
and AND4 (N4061, N4058, N3267, N840, N1475);
xor XOR2 (N4062, N4051, N2947);
and AND2 (N4063, N4034, N1043);
buf BUF1 (N4064, N4057);
nor NOR4 (N4065, N4063, N1010, N2714, N2506);
or OR3 (N4066, N4050, N4058, N59);
and AND3 (N4067, N4064, N1570, N2404);
nand NAND2 (N4068, N4047, N4041);
xor XOR2 (N4069, N4053, N3539);
and AND3 (N4070, N4068, N1385, N952);
buf BUF1 (N4071, N4061);
nor NOR3 (N4072, N4055, N3798, N2088);
or OR2 (N4073, N4072, N1044);
or OR4 (N4074, N4071, N2232, N833, N32);
and AND2 (N4075, N4065, N535);
xor XOR2 (N4076, N4073, N3624);
not NOT1 (N4077, N4075);
or OR4 (N4078, N4048, N50, N415, N1534);
buf BUF1 (N4079, N4074);
nor NOR4 (N4080, N4060, N3791, N61, N4037);
buf BUF1 (N4081, N4080);
or OR3 (N4082, N4077, N3752, N1081);
buf BUF1 (N4083, N4076);
xor XOR2 (N4084, N4083, N181);
not NOT1 (N4085, N4066);
not NOT1 (N4086, N4079);
and AND3 (N4087, N4069, N25, N1480);
nor NOR4 (N4088, N4078, N2271, N688, N3512);
buf BUF1 (N4089, N4082);
nor NOR4 (N4090, N4086, N2932, N683, N2308);
nor NOR2 (N4091, N4062, N225);
nor NOR4 (N4092, N4081, N3569, N3881, N1394);
nor NOR2 (N4093, N4087, N1464);
xor XOR2 (N4094, N4090, N53);
and AND2 (N4095, N4091, N1702);
nor NOR3 (N4096, N4088, N4045, N3770);
nor NOR2 (N4097, N4084, N422);
and AND3 (N4098, N4096, N1333, N554);
xor XOR2 (N4099, N4092, N1424);
or OR3 (N4100, N4085, N2359, N3614);
and AND2 (N4101, N4098, N3767);
or OR3 (N4102, N4097, N1931, N1736);
buf BUF1 (N4103, N4067);
and AND2 (N4104, N4095, N2352);
not NOT1 (N4105, N4100);
and AND4 (N4106, N4094, N2730, N126, N3889);
nor NOR3 (N4107, N4070, N3679, N3349);
and AND4 (N4108, N4106, N2080, N75, N2840);
and AND2 (N4109, N4093, N566);
buf BUF1 (N4110, N4089);
not NOT1 (N4111, N4105);
buf BUF1 (N4112, N4107);
not NOT1 (N4113, N4112);
nand NAND2 (N4114, N4108, N2857);
not NOT1 (N4115, N4104);
buf BUF1 (N4116, N4102);
not NOT1 (N4117, N4099);
nor NOR2 (N4118, N4117, N446);
xor XOR2 (N4119, N4115, N1540);
not NOT1 (N4120, N4116);
nor NOR2 (N4121, N4118, N3624);
xor XOR2 (N4122, N4113, N1559);
not NOT1 (N4123, N4114);
or OR4 (N4124, N4111, N1961, N2187, N1113);
xor XOR2 (N4125, N4123, N1641);
buf BUF1 (N4126, N4109);
xor XOR2 (N4127, N4101, N3846);
nand NAND3 (N4128, N4120, N1212, N835);
xor XOR2 (N4129, N4128, N2915);
not NOT1 (N4130, N4121);
nor NOR3 (N4131, N4125, N334, N3467);
xor XOR2 (N4132, N4110, N4054);
and AND2 (N4133, N4129, N1896);
nand NAND2 (N4134, N4131, N3491);
xor XOR2 (N4135, N4119, N2349);
buf BUF1 (N4136, N4132);
xor XOR2 (N4137, N4127, N4112);
buf BUF1 (N4138, N4133);
xor XOR2 (N4139, N4103, N3433);
or OR4 (N4140, N4136, N1890, N2411, N1217);
buf BUF1 (N4141, N4139);
nor NOR3 (N4142, N4141, N1841, N2246);
buf BUF1 (N4143, N4140);
xor XOR2 (N4144, N4137, N3417);
nand NAND2 (N4145, N4143, N1633);
not NOT1 (N4146, N4122);
and AND4 (N4147, N4138, N1551, N3121, N2676);
nand NAND3 (N4148, N4134, N503, N19);
nand NAND2 (N4149, N4124, N3696);
not NOT1 (N4150, N4130);
or OR3 (N4151, N4135, N2497, N1059);
or OR4 (N4152, N4148, N1133, N613, N1223);
and AND3 (N4153, N4146, N844, N1440);
and AND3 (N4154, N4144, N1096, N848);
and AND4 (N4155, N4147, N319, N2749, N1363);
buf BUF1 (N4156, N4149);
or OR4 (N4157, N4156, N2950, N928, N1092);
nand NAND4 (N4158, N4142, N4062, N377, N3594);
nand NAND2 (N4159, N4155, N4156);
nand NAND4 (N4160, N4126, N3253, N3867, N3736);
buf BUF1 (N4161, N4159);
or OR2 (N4162, N4153, N795);
or OR3 (N4163, N4150, N2583, N2552);
not NOT1 (N4164, N4151);
not NOT1 (N4165, N4161);
nor NOR4 (N4166, N4163, N2339, N2753, N1011);
nor NOR2 (N4167, N4166, N1426);
nand NAND2 (N4168, N4152, N1766);
buf BUF1 (N4169, N4157);
or OR2 (N4170, N4158, N3382);
xor XOR2 (N4171, N4145, N1585);
nor NOR3 (N4172, N4171, N3067, N1788);
buf BUF1 (N4173, N4169);
buf BUF1 (N4174, N4172);
nand NAND2 (N4175, N4174, N2288);
xor XOR2 (N4176, N4170, N1442);
and AND4 (N4177, N4162, N3247, N459, N3088);
xor XOR2 (N4178, N4173, N2405);
or OR4 (N4179, N4164, N2393, N1234, N3076);
or OR2 (N4180, N4160, N2537);
nand NAND3 (N4181, N4180, N1304, N4081);
nand NAND4 (N4182, N4167, N2777, N3056, N1975);
xor XOR2 (N4183, N4175, N1376);
or OR2 (N4184, N4154, N2349);
nor NOR3 (N4185, N4179, N131, N2970);
nor NOR2 (N4186, N4185, N3239);
and AND2 (N4187, N4165, N2795);
buf BUF1 (N4188, N4178);
buf BUF1 (N4189, N4168);
and AND4 (N4190, N4187, N2627, N4096, N2998);
nand NAND4 (N4191, N4182, N3530, N3690, N1652);
nand NAND4 (N4192, N4183, N865, N3113, N4168);
or OR3 (N4193, N4176, N2987, N3770);
or OR2 (N4194, N4191, N100);
xor XOR2 (N4195, N4194, N2497);
buf BUF1 (N4196, N4189);
or OR2 (N4197, N4181, N2413);
buf BUF1 (N4198, N4188);
nor NOR4 (N4199, N4197, N2591, N1380, N206);
buf BUF1 (N4200, N4193);
and AND4 (N4201, N4186, N2469, N2200, N1208);
buf BUF1 (N4202, N4200);
buf BUF1 (N4203, N4199);
or OR2 (N4204, N4196, N334);
and AND4 (N4205, N4192, N1588, N2043, N124);
nor NOR4 (N4206, N4204, N154, N930, N953);
nor NOR2 (N4207, N4205, N4013);
buf BUF1 (N4208, N4203);
nor NOR3 (N4209, N4201, N126, N289);
not NOT1 (N4210, N4195);
and AND2 (N4211, N4206, N3230);
or OR3 (N4212, N4207, N1492, N1640);
nand NAND3 (N4213, N4184, N3299, N886);
and AND2 (N4214, N4190, N2446);
xor XOR2 (N4215, N4202, N502);
nor NOR3 (N4216, N4214, N4018, N1101);
nand NAND3 (N4217, N4210, N2331, N2879);
not NOT1 (N4218, N4215);
not NOT1 (N4219, N4218);
buf BUF1 (N4220, N4198);
nand NAND4 (N4221, N4217, N1567, N1825, N2889);
xor XOR2 (N4222, N4208, N1314);
nand NAND4 (N4223, N4219, N2457, N3640, N1479);
and AND4 (N4224, N4221, N2984, N4216, N46);
nor NOR4 (N4225, N3081, N1809, N980, N2242);
nor NOR3 (N4226, N4223, N3723, N3255);
not NOT1 (N4227, N4220);
buf BUF1 (N4228, N4209);
nor NOR4 (N4229, N4227, N1956, N1782, N2218);
nor NOR3 (N4230, N4212, N1699, N2742);
buf BUF1 (N4231, N4222);
nand NAND3 (N4232, N4230, N2098, N2546);
or OR3 (N4233, N4228, N2090, N3458);
nor NOR3 (N4234, N4177, N2841, N4107);
nand NAND2 (N4235, N4229, N1913);
not NOT1 (N4236, N4235);
nand NAND3 (N4237, N4224, N3325, N1054);
buf BUF1 (N4238, N4236);
nand NAND3 (N4239, N4226, N637, N2810);
not NOT1 (N4240, N4232);
xor XOR2 (N4241, N4231, N511);
and AND2 (N4242, N4234, N302);
and AND3 (N4243, N4237, N2903, N1199);
and AND2 (N4244, N4241, N2251);
and AND3 (N4245, N4242, N3833, N3509);
not NOT1 (N4246, N4233);
nor NOR2 (N4247, N4238, N3240);
nor NOR4 (N4248, N4245, N3910, N3218, N3435);
not NOT1 (N4249, N4246);
xor XOR2 (N4250, N4239, N3078);
buf BUF1 (N4251, N4240);
nor NOR4 (N4252, N4211, N3884, N206, N2474);
xor XOR2 (N4253, N4251, N2771);
nor NOR3 (N4254, N4253, N3103, N2829);
xor XOR2 (N4255, N4244, N912);
and AND3 (N4256, N4254, N3318, N3323);
and AND2 (N4257, N4225, N1119);
or OR3 (N4258, N4256, N145, N4036);
not NOT1 (N4259, N4249);
and AND4 (N4260, N4257, N2311, N3716, N660);
or OR3 (N4261, N4247, N4175, N2216);
or OR2 (N4262, N4252, N1463);
and AND2 (N4263, N4250, N1199);
buf BUF1 (N4264, N4260);
buf BUF1 (N4265, N4262);
not NOT1 (N4266, N4263);
xor XOR2 (N4267, N4265, N2901);
not NOT1 (N4268, N4243);
nor NOR2 (N4269, N4266, N1550);
nand NAND3 (N4270, N4259, N3980, N715);
and AND2 (N4271, N4264, N3930);
xor XOR2 (N4272, N4213, N3598);
nor NOR4 (N4273, N4267, N4160, N3770, N3236);
nor NOR2 (N4274, N4272, N1178);
nor NOR3 (N4275, N4248, N729, N324);
or OR2 (N4276, N4271, N322);
nand NAND2 (N4277, N4273, N2125);
or OR2 (N4278, N4258, N903);
or OR2 (N4279, N4276, N2370);
nand NAND3 (N4280, N4268, N3973, N3716);
or OR4 (N4281, N4261, N3632, N4159, N454);
xor XOR2 (N4282, N4274, N2886);
not NOT1 (N4283, N4277);
nand NAND2 (N4284, N4255, N45);
nand NAND3 (N4285, N4275, N3534, N3868);
buf BUF1 (N4286, N4280);
or OR3 (N4287, N4269, N202, N4016);
and AND3 (N4288, N4286, N428, N2738);
nand NAND2 (N4289, N4284, N7);
and AND4 (N4290, N4282, N111, N4181, N2118);
nor NOR3 (N4291, N4290, N127, N1808);
buf BUF1 (N4292, N4285);
nand NAND3 (N4293, N4278, N2501, N3130);
and AND2 (N4294, N4288, N1072);
or OR2 (N4295, N4279, N3130);
not NOT1 (N4296, N4294);
not NOT1 (N4297, N4291);
and AND2 (N4298, N4270, N776);
not NOT1 (N4299, N4287);
buf BUF1 (N4300, N4296);
not NOT1 (N4301, N4293);
not NOT1 (N4302, N4298);
not NOT1 (N4303, N4301);
or OR2 (N4304, N4295, N1994);
buf BUF1 (N4305, N4299);
xor XOR2 (N4306, N4283, N1212);
nor NOR2 (N4307, N4304, N2330);
buf BUF1 (N4308, N4281);
nand NAND2 (N4309, N4307, N336);
nor NOR3 (N4310, N4297, N649, N2987);
or OR3 (N4311, N4306, N483, N887);
buf BUF1 (N4312, N4292);
nand NAND3 (N4313, N4310, N853, N3154);
not NOT1 (N4314, N4300);
not NOT1 (N4315, N4302);
nor NOR2 (N4316, N4309, N1925);
nand NAND2 (N4317, N4308, N3012);
nor NOR4 (N4318, N4311, N3161, N545, N561);
nor NOR3 (N4319, N4314, N1430, N377);
buf BUF1 (N4320, N4313);
nand NAND3 (N4321, N4318, N4276, N4099);
nor NOR3 (N4322, N4305, N3085, N829);
or OR3 (N4323, N4321, N4127, N3181);
xor XOR2 (N4324, N4322, N3915);
nand NAND2 (N4325, N4316, N3670);
or OR3 (N4326, N4312, N1248, N416);
xor XOR2 (N4327, N4323, N2214);
or OR3 (N4328, N4315, N2323, N33);
not NOT1 (N4329, N4320);
or OR2 (N4330, N4319, N2468);
buf BUF1 (N4331, N4327);
buf BUF1 (N4332, N4317);
nand NAND3 (N4333, N4303, N1678, N4193);
and AND3 (N4334, N4289, N3011, N3460);
and AND3 (N4335, N4330, N1091, N2643);
or OR2 (N4336, N4326, N193);
nand NAND3 (N4337, N4333, N1720, N3502);
nor NOR2 (N4338, N4336, N3785);
or OR4 (N4339, N4325, N2722, N1275, N1311);
nand NAND3 (N4340, N4324, N2565, N663);
xor XOR2 (N4341, N4339, N2873);
buf BUF1 (N4342, N4332);
and AND2 (N4343, N4338, N1584);
or OR4 (N4344, N4337, N3747, N2326, N3029);
or OR3 (N4345, N4328, N13, N3422);
nand NAND2 (N4346, N4344, N1985);
buf BUF1 (N4347, N4343);
nand NAND2 (N4348, N4340, N3039);
nor NOR4 (N4349, N4329, N2460, N307, N1342);
and AND3 (N4350, N4335, N1649, N756);
not NOT1 (N4351, N4350);
not NOT1 (N4352, N4334);
or OR2 (N4353, N4345, N4257);
or OR3 (N4354, N4342, N3587, N3424);
buf BUF1 (N4355, N4348);
not NOT1 (N4356, N4349);
xor XOR2 (N4357, N4347, N3272);
not NOT1 (N4358, N4355);
nand NAND2 (N4359, N4353, N2196);
not NOT1 (N4360, N4359);
nand NAND3 (N4361, N4341, N3612, N3935);
xor XOR2 (N4362, N4354, N2968);
buf BUF1 (N4363, N4346);
nand NAND3 (N4364, N4356, N4049, N4070);
buf BUF1 (N4365, N4362);
not NOT1 (N4366, N4361);
and AND3 (N4367, N4331, N1268, N3947);
buf BUF1 (N4368, N4367);
buf BUF1 (N4369, N4364);
or OR2 (N4370, N4360, N1989);
buf BUF1 (N4371, N4370);
not NOT1 (N4372, N4369);
nor NOR2 (N4373, N4352, N713);
buf BUF1 (N4374, N4368);
nor NOR3 (N4375, N4365, N1452, N4374);
not NOT1 (N4376, N2708);
nor NOR4 (N4377, N4363, N2070, N2212, N2457);
or OR2 (N4378, N4357, N210);
nand NAND3 (N4379, N4366, N2105, N1217);
and AND2 (N4380, N4376, N2199);
and AND2 (N4381, N4375, N3649);
buf BUF1 (N4382, N4378);
and AND2 (N4383, N4377, N4251);
nor NOR4 (N4384, N4372, N1205, N1427, N46);
nor NOR4 (N4385, N4371, N1723, N3028, N2558);
not NOT1 (N4386, N4351);
nor NOR4 (N4387, N4380, N2528, N2491, N2605);
buf BUF1 (N4388, N4358);
buf BUF1 (N4389, N4386);
and AND3 (N4390, N4385, N1833, N3252);
and AND2 (N4391, N4379, N73);
xor XOR2 (N4392, N4390, N1627);
xor XOR2 (N4393, N4373, N1861);
nor NOR3 (N4394, N4381, N711, N3099);
buf BUF1 (N4395, N4389);
nor NOR2 (N4396, N4392, N3944);
or OR2 (N4397, N4395, N406);
nand NAND2 (N4398, N4383, N1666);
buf BUF1 (N4399, N4391);
and AND4 (N4400, N4384, N2474, N2126, N286);
nand NAND2 (N4401, N4388, N1371);
buf BUF1 (N4402, N4397);
not NOT1 (N4403, N4396);
nand NAND2 (N4404, N4382, N964);
nand NAND2 (N4405, N4402, N2564);
not NOT1 (N4406, N4401);
xor XOR2 (N4407, N4393, N1057);
xor XOR2 (N4408, N4404, N111);
xor XOR2 (N4409, N4408, N1161);
xor XOR2 (N4410, N4405, N1066);
or OR3 (N4411, N4399, N1091, N641);
or OR2 (N4412, N4398, N1661);
not NOT1 (N4413, N4412);
or OR4 (N4414, N4406, N2042, N1651, N3067);
xor XOR2 (N4415, N4400, N461);
xor XOR2 (N4416, N4411, N621);
nor NOR3 (N4417, N4394, N4185, N1593);
xor XOR2 (N4418, N4403, N1080);
nand NAND3 (N4419, N4410, N3331, N3368);
nand NAND2 (N4420, N4387, N514);
and AND2 (N4421, N4420, N3505);
buf BUF1 (N4422, N4417);
buf BUF1 (N4423, N4409);
nor NOR4 (N4424, N4418, N1489, N2141, N2838);
nor NOR4 (N4425, N4415, N4208, N139, N3328);
nand NAND2 (N4426, N4419, N147);
and AND3 (N4427, N4407, N3035, N1286);
or OR4 (N4428, N4414, N540, N344, N2988);
or OR3 (N4429, N4428, N1571, N2137);
xor XOR2 (N4430, N4422, N5);
xor XOR2 (N4431, N4423, N876);
nand NAND4 (N4432, N4413, N305, N4003, N434);
nor NOR3 (N4433, N4426, N2520, N1411);
buf BUF1 (N4434, N4433);
and AND3 (N4435, N4431, N2273, N2602);
or OR3 (N4436, N4424, N1250, N2603);
and AND3 (N4437, N4436, N1273, N4276);
nor NOR4 (N4438, N4435, N1386, N4240, N974);
and AND3 (N4439, N4427, N3353, N1399);
xor XOR2 (N4440, N4425, N2257);
buf BUF1 (N4441, N4439);
nor NOR4 (N4442, N4437, N2378, N2807, N70);
nand NAND4 (N4443, N4416, N669, N2906, N619);
xor XOR2 (N4444, N4442, N3409);
buf BUF1 (N4445, N4430);
and AND2 (N4446, N4441, N1132);
not NOT1 (N4447, N4432);
xor XOR2 (N4448, N4421, N3190);
or OR2 (N4449, N4443, N1793);
not NOT1 (N4450, N4444);
or OR2 (N4451, N4446, N3684);
xor XOR2 (N4452, N4445, N607);
or OR4 (N4453, N4429, N2935, N3719, N113);
or OR2 (N4454, N4451, N1601);
buf BUF1 (N4455, N4438);
not NOT1 (N4456, N4448);
nor NOR2 (N4457, N4453, N1220);
not NOT1 (N4458, N4440);
and AND4 (N4459, N4449, N1307, N3869, N2113);
buf BUF1 (N4460, N4454);
not NOT1 (N4461, N4450);
nand NAND4 (N4462, N4452, N2576, N2958, N740);
buf BUF1 (N4463, N4462);
buf BUF1 (N4464, N4434);
and AND2 (N4465, N4460, N3845);
not NOT1 (N4466, N4457);
or OR2 (N4467, N4461, N1163);
xor XOR2 (N4468, N4466, N2091);
not NOT1 (N4469, N4468);
xor XOR2 (N4470, N4465, N2062);
or OR3 (N4471, N4456, N3121, N1381);
nand NAND2 (N4472, N4470, N448);
and AND2 (N4473, N4469, N3703);
xor XOR2 (N4474, N4458, N2296);
nor NOR2 (N4475, N4471, N2789);
or OR4 (N4476, N4455, N4216, N360, N3582);
not NOT1 (N4477, N4473);
buf BUF1 (N4478, N4475);
and AND4 (N4479, N4477, N2637, N2045, N866);
and AND3 (N4480, N4467, N1443, N1759);
xor XOR2 (N4481, N4447, N1096);
nand NAND4 (N4482, N4479, N727, N57, N786);
and AND4 (N4483, N4464, N1191, N273, N1103);
xor XOR2 (N4484, N4483, N854);
nor NOR2 (N4485, N4474, N3794);
xor XOR2 (N4486, N4482, N3960);
or OR3 (N4487, N4484, N1855, N2304);
not NOT1 (N4488, N4487);
nor NOR2 (N4489, N4472, N372);
or OR2 (N4490, N4489, N3227);
nand NAND2 (N4491, N4480, N56);
nand NAND3 (N4492, N4476, N1494, N3664);
xor XOR2 (N4493, N4478, N3009);
xor XOR2 (N4494, N4490, N661);
buf BUF1 (N4495, N4481);
nand NAND3 (N4496, N4493, N3317, N1587);
and AND4 (N4497, N4488, N3293, N4213, N960);
or OR2 (N4498, N4497, N187);
and AND3 (N4499, N4492, N4139, N1541);
and AND3 (N4500, N4491, N3567, N3200);
nand NAND3 (N4501, N4499, N3530, N4364);
not NOT1 (N4502, N4500);
or OR2 (N4503, N4496, N3307);
nand NAND2 (N4504, N4501, N3042);
xor XOR2 (N4505, N4486, N2598);
not NOT1 (N4506, N4502);
not NOT1 (N4507, N4503);
nand NAND2 (N4508, N4485, N1876);
nor NOR4 (N4509, N4494, N607, N3595, N2814);
and AND2 (N4510, N4498, N329);
or OR3 (N4511, N4463, N1724, N2648);
nor NOR3 (N4512, N4509, N2887, N143);
buf BUF1 (N4513, N4506);
not NOT1 (N4514, N4459);
xor XOR2 (N4515, N4514, N3525);
nand NAND4 (N4516, N4505, N3809, N33, N697);
and AND4 (N4517, N4511, N813, N3385, N2812);
xor XOR2 (N4518, N4513, N3816);
nor NOR2 (N4519, N4504, N4100);
xor XOR2 (N4520, N4512, N1743);
nand NAND4 (N4521, N4507, N3161, N2464, N4357);
and AND2 (N4522, N4519, N366);
nor NOR2 (N4523, N4515, N2309);
nor NOR4 (N4524, N4508, N677, N4301, N3931);
nor NOR2 (N4525, N4518, N3651);
buf BUF1 (N4526, N4510);
buf BUF1 (N4527, N4520);
buf BUF1 (N4528, N4521);
xor XOR2 (N4529, N4528, N1127);
buf BUF1 (N4530, N4527);
nor NOR4 (N4531, N4524, N1820, N2694, N3201);
xor XOR2 (N4532, N4522, N2754);
nor NOR4 (N4533, N4526, N247, N1, N3849);
nor NOR4 (N4534, N4532, N1614, N1156, N1224);
or OR2 (N4535, N4523, N640);
nor NOR4 (N4536, N4531, N3116, N2124, N3884);
and AND3 (N4537, N4533, N3425, N1404);
nor NOR4 (N4538, N4537, N4171, N503, N880);
xor XOR2 (N4539, N4529, N3905);
buf BUF1 (N4540, N4516);
or OR4 (N4541, N4517, N1309, N436, N2249);
nor NOR2 (N4542, N4538, N1413);
xor XOR2 (N4543, N4534, N1913);
nand NAND4 (N4544, N4540, N266, N778, N1981);
and AND4 (N4545, N4536, N1234, N635, N2448);
nor NOR3 (N4546, N4535, N3100, N1238);
buf BUF1 (N4547, N4541);
nor NOR4 (N4548, N4543, N2357, N2285, N4154);
or OR2 (N4549, N4495, N701);
buf BUF1 (N4550, N4539);
xor XOR2 (N4551, N4525, N3714);
buf BUF1 (N4552, N4547);
or OR4 (N4553, N4544, N1488, N4381, N3036);
or OR4 (N4554, N4550, N1824, N3245, N2925);
buf BUF1 (N4555, N4549);
and AND4 (N4556, N4530, N3265, N1118, N1964);
not NOT1 (N4557, N4556);
buf BUF1 (N4558, N4548);
buf BUF1 (N4559, N4546);
not NOT1 (N4560, N4542);
buf BUF1 (N4561, N4553);
or OR3 (N4562, N4561, N4421, N379);
buf BUF1 (N4563, N4555);
nand NAND4 (N4564, N4545, N3786, N2615, N2469);
not NOT1 (N4565, N4559);
xor XOR2 (N4566, N4562, N1326);
nor NOR3 (N4567, N4552, N926, N2195);
xor XOR2 (N4568, N4566, N1139);
buf BUF1 (N4569, N4563);
and AND3 (N4570, N4567, N637, N4067);
buf BUF1 (N4571, N4560);
nand NAND4 (N4572, N4568, N539, N2512, N2395);
or OR3 (N4573, N4557, N1998, N4503);
xor XOR2 (N4574, N4565, N227);
nor NOR3 (N4575, N4551, N1971, N2095);
and AND2 (N4576, N4574, N225);
nand NAND3 (N4577, N4573, N1815, N1725);
and AND2 (N4578, N4558, N816);
and AND3 (N4579, N4578, N3587, N3020);
buf BUF1 (N4580, N4564);
buf BUF1 (N4581, N4554);
and AND3 (N4582, N4580, N2017, N2854);
or OR2 (N4583, N4572, N670);
nor NOR3 (N4584, N4569, N109, N1646);
nor NOR2 (N4585, N4577, N3775);
and AND4 (N4586, N4570, N414, N1133, N1748);
and AND4 (N4587, N4585, N2020, N1937, N2589);
not NOT1 (N4588, N4587);
nand NAND3 (N4589, N4584, N2213, N3017);
buf BUF1 (N4590, N4583);
not NOT1 (N4591, N4588);
buf BUF1 (N4592, N4579);
buf BUF1 (N4593, N4589);
xor XOR2 (N4594, N4576, N1638);
nor NOR4 (N4595, N4586, N3369, N3490, N3047);
xor XOR2 (N4596, N4594, N2710);
and AND4 (N4597, N4596, N2574, N3081, N497);
or OR3 (N4598, N4590, N253, N2775);
and AND2 (N4599, N4593, N2368);
not NOT1 (N4600, N4591);
or OR4 (N4601, N4592, N2980, N3132, N2306);
and AND3 (N4602, N4597, N655, N3738);
or OR4 (N4603, N4581, N2804, N4116, N1579);
nor NOR2 (N4604, N4571, N3312);
and AND2 (N4605, N4603, N3812);
or OR3 (N4606, N4595, N3779, N3883);
and AND2 (N4607, N4582, N3095);
nand NAND2 (N4608, N4601, N3072);
and AND4 (N4609, N4607, N834, N3791, N3815);
nand NAND2 (N4610, N4605, N2777);
buf BUF1 (N4611, N4606);
buf BUF1 (N4612, N4604);
and AND3 (N4613, N4598, N1227, N4581);
buf BUF1 (N4614, N4575);
or OR4 (N4615, N4611, N2610, N1380, N3515);
or OR3 (N4616, N4609, N86, N3108);
xor XOR2 (N4617, N4600, N3709);
and AND3 (N4618, N4615, N532, N3122);
xor XOR2 (N4619, N4616, N4321);
buf BUF1 (N4620, N4619);
or OR2 (N4621, N4599, N1570);
xor XOR2 (N4622, N4620, N473);
xor XOR2 (N4623, N4622, N78);
nand NAND4 (N4624, N4623, N4109, N3766, N851);
nand NAND4 (N4625, N4610, N3815, N2763, N1491);
buf BUF1 (N4626, N4624);
nand NAND4 (N4627, N4617, N2436, N3750, N2645);
nor NOR2 (N4628, N4602, N3850);
and AND3 (N4629, N4626, N4010, N3185);
or OR2 (N4630, N4618, N2839);
and AND2 (N4631, N4614, N1035);
and AND4 (N4632, N4630, N2989, N1978, N2936);
and AND3 (N4633, N4621, N397, N3129);
nand NAND3 (N4634, N4628, N2459, N4498);
nor NOR2 (N4635, N4612, N356);
nand NAND3 (N4636, N4627, N3871, N712);
nor NOR4 (N4637, N4631, N2606, N4635, N4133);
xor XOR2 (N4638, N1863, N3493);
or OR4 (N4639, N4633, N2935, N4340, N2862);
and AND3 (N4640, N4629, N883, N1119);
and AND3 (N4641, N4632, N3356, N2783);
nor NOR4 (N4642, N4634, N3698, N1448, N4569);
nand NAND4 (N4643, N4613, N1990, N245, N2148);
and AND2 (N4644, N4625, N934);
not NOT1 (N4645, N4642);
buf BUF1 (N4646, N4645);
nor NOR3 (N4647, N4641, N3816, N1913);
or OR3 (N4648, N4636, N4351, N2908);
buf BUF1 (N4649, N4638);
xor XOR2 (N4650, N4640, N3694);
and AND2 (N4651, N4647, N1718);
buf BUF1 (N4652, N4639);
buf BUF1 (N4653, N4644);
and AND4 (N4654, N4608, N163, N2761, N4122);
or OR2 (N4655, N4652, N4450);
not NOT1 (N4656, N4654);
not NOT1 (N4657, N4653);
not NOT1 (N4658, N4651);
not NOT1 (N4659, N4643);
xor XOR2 (N4660, N4658, N4021);
and AND2 (N4661, N4650, N926);
or OR2 (N4662, N4649, N2429);
or OR3 (N4663, N4637, N1523, N3960);
not NOT1 (N4664, N4648);
and AND4 (N4665, N4663, N10, N3078, N4559);
xor XOR2 (N4666, N4662, N4046);
not NOT1 (N4667, N4665);
nor NOR3 (N4668, N4656, N3906, N2664);
and AND4 (N4669, N4655, N3199, N1308, N4491);
buf BUF1 (N4670, N4667);
or OR3 (N4671, N4670, N1003, N1770);
or OR4 (N4672, N4669, N1270, N1238, N380);
buf BUF1 (N4673, N4646);
or OR3 (N4674, N4660, N2727, N1695);
nand NAND3 (N4675, N4671, N4453, N2992);
and AND3 (N4676, N4657, N3403, N4207);
buf BUF1 (N4677, N4666);
and AND4 (N4678, N4673, N4274, N1014, N2435);
or OR4 (N4679, N4664, N1849, N164, N3477);
nor NOR2 (N4680, N4679, N2411);
buf BUF1 (N4681, N4680);
or OR3 (N4682, N4676, N2732, N2345);
xor XOR2 (N4683, N4675, N572);
or OR3 (N4684, N4682, N1458, N2281);
nor NOR3 (N4685, N4668, N3408, N4104);
or OR2 (N4686, N4677, N1556);
not NOT1 (N4687, N4674);
or OR3 (N4688, N4683, N3906, N1139);
xor XOR2 (N4689, N4672, N1961);
nor NOR4 (N4690, N4659, N3718, N3934, N4089);
nor NOR3 (N4691, N4685, N2448, N1948);
not NOT1 (N4692, N4690);
xor XOR2 (N4693, N4681, N2524);
nand NAND2 (N4694, N4684, N4228);
nand NAND4 (N4695, N4689, N4335, N735, N1495);
nor NOR3 (N4696, N4693, N4257, N892);
and AND4 (N4697, N4678, N882, N3220, N3876);
or OR4 (N4698, N4695, N93, N1939, N3198);
or OR3 (N4699, N4694, N834, N591);
not NOT1 (N4700, N4688);
and AND2 (N4701, N4696, N3212);
buf BUF1 (N4702, N4691);
or OR4 (N4703, N4661, N3614, N4611, N3203);
xor XOR2 (N4704, N4702, N4036);
not NOT1 (N4705, N4703);
xor XOR2 (N4706, N4705, N1217);
xor XOR2 (N4707, N4697, N4100);
not NOT1 (N4708, N4707);
buf BUF1 (N4709, N4706);
and AND2 (N4710, N4708, N4434);
nor NOR3 (N4711, N4704, N2168, N3337);
xor XOR2 (N4712, N4686, N660);
not NOT1 (N4713, N4700);
nand NAND2 (N4714, N4711, N4538);
not NOT1 (N4715, N4710);
not NOT1 (N4716, N4698);
and AND4 (N4717, N4692, N2161, N2975, N4367);
and AND2 (N4718, N4701, N1241);
nand NAND3 (N4719, N4687, N3740, N4423);
or OR2 (N4720, N4719, N405);
xor XOR2 (N4721, N4717, N269);
and AND4 (N4722, N4715, N4287, N4490, N4013);
and AND2 (N4723, N4720, N3150);
xor XOR2 (N4724, N4721, N1546);
not NOT1 (N4725, N4709);
nand NAND3 (N4726, N4723, N291, N4069);
not NOT1 (N4727, N4699);
nand NAND3 (N4728, N4713, N2465, N420);
buf BUF1 (N4729, N4722);
or OR3 (N4730, N4724, N2727, N4695);
nor NOR4 (N4731, N4725, N2601, N2292, N2119);
nand NAND3 (N4732, N4730, N1251, N1140);
nand NAND2 (N4733, N4714, N3278);
or OR4 (N4734, N4728, N2690, N3551, N2545);
not NOT1 (N4735, N4734);
not NOT1 (N4736, N4729);
or OR2 (N4737, N4731, N2575);
buf BUF1 (N4738, N4716);
nand NAND2 (N4739, N4712, N4121);
nor NOR4 (N4740, N4739, N1743, N572, N4495);
nand NAND4 (N4741, N4727, N914, N2396, N3167);
xor XOR2 (N4742, N4726, N3442);
nand NAND4 (N4743, N4735, N2138, N1390, N2393);
xor XOR2 (N4744, N4742, N1251);
and AND3 (N4745, N4740, N4638, N937);
buf BUF1 (N4746, N4745);
buf BUF1 (N4747, N4733);
and AND4 (N4748, N4732, N2984, N4547, N1509);
xor XOR2 (N4749, N4743, N3476);
not NOT1 (N4750, N4718);
not NOT1 (N4751, N4749);
or OR3 (N4752, N4746, N228, N558);
or OR3 (N4753, N4747, N3969, N1652);
not NOT1 (N4754, N4753);
nor NOR3 (N4755, N4750, N4651, N3806);
or OR2 (N4756, N4752, N1762);
xor XOR2 (N4757, N4754, N1932);
xor XOR2 (N4758, N4755, N3590);
and AND3 (N4759, N4741, N4022, N2942);
or OR3 (N4760, N4757, N739, N3395);
nor NOR4 (N4761, N4760, N1124, N899, N557);
nor NOR2 (N4762, N4738, N295);
buf BUF1 (N4763, N4756);
nor NOR4 (N4764, N4761, N1242, N309, N965);
nor NOR3 (N4765, N4751, N879, N1920);
buf BUF1 (N4766, N4748);
nor NOR3 (N4767, N4758, N2808, N3473);
not NOT1 (N4768, N4764);
xor XOR2 (N4769, N4759, N1574);
buf BUF1 (N4770, N4744);
nand NAND3 (N4771, N4769, N3570, N2012);
nor NOR2 (N4772, N4765, N1393);
nand NAND2 (N4773, N4762, N3053);
nor NOR3 (N4774, N4737, N992, N1368);
nand NAND2 (N4775, N4767, N1276);
buf BUF1 (N4776, N4771);
or OR4 (N4777, N4770, N623, N2725, N1473);
or OR3 (N4778, N4763, N1983, N2303);
buf BUF1 (N4779, N4777);
not NOT1 (N4780, N4775);
or OR2 (N4781, N4779, N3150);
and AND2 (N4782, N4778, N2300);
not NOT1 (N4783, N4773);
nand NAND3 (N4784, N4774, N210, N4006);
nand NAND4 (N4785, N4780, N2182, N128, N2810);
and AND3 (N4786, N4785, N2662, N3406);
or OR2 (N4787, N4776, N4672);
and AND4 (N4788, N4772, N2724, N1377, N4782);
nand NAND2 (N4789, N1430, N4644);
and AND3 (N4790, N4781, N682, N260);
buf BUF1 (N4791, N4784);
buf BUF1 (N4792, N4787);
buf BUF1 (N4793, N4790);
nand NAND4 (N4794, N4791, N2901, N4280, N1360);
xor XOR2 (N4795, N4766, N661);
not NOT1 (N4796, N4768);
nor NOR2 (N4797, N4786, N3089);
xor XOR2 (N4798, N4788, N1970);
nand NAND2 (N4799, N4798, N2327);
not NOT1 (N4800, N4736);
nand NAND4 (N4801, N4800, N3192, N1048, N3034);
buf BUF1 (N4802, N4795);
nor NOR4 (N4803, N4799, N3842, N3463, N3528);
nand NAND2 (N4804, N4797, N536);
not NOT1 (N4805, N4794);
buf BUF1 (N4806, N4805);
or OR2 (N4807, N4803, N2521);
and AND2 (N4808, N4807, N4096);
nand NAND3 (N4809, N4804, N3035, N3864);
xor XOR2 (N4810, N4809, N3362);
xor XOR2 (N4811, N4806, N1962);
buf BUF1 (N4812, N4801);
or OR2 (N4813, N4792, N1370);
not NOT1 (N4814, N4796);
or OR3 (N4815, N4813, N3986, N2239);
nand NAND2 (N4816, N4814, N1863);
xor XOR2 (N4817, N4808, N1268);
and AND3 (N4818, N4815, N1119, N4375);
xor XOR2 (N4819, N4811, N3874);
nand NAND3 (N4820, N4789, N2037, N2149);
xor XOR2 (N4821, N4812, N4150);
xor XOR2 (N4822, N4817, N2437);
buf BUF1 (N4823, N4818);
nor NOR3 (N4824, N4802, N3308, N4691);
not NOT1 (N4825, N4822);
or OR2 (N4826, N4823, N3245);
xor XOR2 (N4827, N4793, N954);
nor NOR3 (N4828, N4810, N3728, N4202);
xor XOR2 (N4829, N4819, N3727);
buf BUF1 (N4830, N4816);
xor XOR2 (N4831, N4826, N984);
not NOT1 (N4832, N4828);
nand NAND3 (N4833, N4827, N2257, N1568);
xor XOR2 (N4834, N4829, N3627);
nand NAND2 (N4835, N4832, N255);
buf BUF1 (N4836, N4834);
and AND4 (N4837, N4783, N1702, N4076, N3964);
nand NAND4 (N4838, N4830, N242, N4006, N4185);
nand NAND4 (N4839, N4833, N1039, N4738, N3285);
buf BUF1 (N4840, N4824);
and AND4 (N4841, N4821, N290, N477, N3609);
or OR2 (N4842, N4836, N633);
not NOT1 (N4843, N4831);
buf BUF1 (N4844, N4825);
nand NAND4 (N4845, N4820, N2418, N335, N1072);
nor NOR2 (N4846, N4842, N4514);
nor NOR2 (N4847, N4840, N161);
not NOT1 (N4848, N4835);
nor NOR3 (N4849, N4839, N3756, N2729);
buf BUF1 (N4850, N4837);
nand NAND3 (N4851, N4849, N1151, N727);
nand NAND2 (N4852, N4848, N4538);
buf BUF1 (N4853, N4851);
nand NAND2 (N4854, N4853, N4291);
or OR3 (N4855, N4854, N1121, N3330);
nor NOR3 (N4856, N4850, N2053, N1388);
or OR2 (N4857, N4844, N3758);
xor XOR2 (N4858, N4841, N1859);
buf BUF1 (N4859, N4852);
xor XOR2 (N4860, N4843, N1932);
nand NAND2 (N4861, N4860, N1874);
nand NAND4 (N4862, N4859, N2774, N3218, N3031);
and AND3 (N4863, N4856, N524, N4014);
not NOT1 (N4864, N4838);
nor NOR3 (N4865, N4864, N1772, N869);
or OR4 (N4866, N4862, N2541, N3228, N236);
and AND3 (N4867, N4845, N595, N4753);
not NOT1 (N4868, N4866);
and AND4 (N4869, N4867, N899, N4149, N548);
not NOT1 (N4870, N4863);
nand NAND2 (N4871, N4865, N3957);
xor XOR2 (N4872, N4847, N3151);
nand NAND3 (N4873, N4855, N2857, N3517);
and AND2 (N4874, N4870, N3965);
or OR4 (N4875, N4872, N1285, N1801, N3560);
not NOT1 (N4876, N4869);
xor XOR2 (N4877, N4871, N2249);
nor NOR2 (N4878, N4858, N4403);
nand NAND4 (N4879, N4868, N2819, N1587, N2651);
xor XOR2 (N4880, N4846, N3664);
buf BUF1 (N4881, N4877);
nor NOR4 (N4882, N4878, N1908, N835, N1481);
and AND3 (N4883, N4875, N280, N2615);
not NOT1 (N4884, N4876);
nand NAND2 (N4885, N4857, N1156);
nand NAND4 (N4886, N4879, N1842, N1089, N2808);
not NOT1 (N4887, N4886);
not NOT1 (N4888, N4880);
xor XOR2 (N4889, N4884, N1943);
xor XOR2 (N4890, N4887, N4780);
and AND3 (N4891, N4874, N391, N4105);
buf BUF1 (N4892, N4861);
or OR4 (N4893, N4888, N819, N4617, N4620);
or OR4 (N4894, N4892, N1759, N1844, N2233);
buf BUF1 (N4895, N4893);
nor NOR2 (N4896, N4885, N2272);
or OR3 (N4897, N4891, N1967, N172);
nor NOR4 (N4898, N4895, N2416, N1612, N335);
or OR2 (N4899, N4897, N2274);
and AND3 (N4900, N4899, N4726, N4629);
nor NOR2 (N4901, N4900, N17);
not NOT1 (N4902, N4883);
buf BUF1 (N4903, N4882);
nand NAND2 (N4904, N4898, N3773);
or OR3 (N4905, N4903, N1737, N1831);
or OR3 (N4906, N4901, N2504, N1884);
and AND2 (N4907, N4896, N2485);
nor NOR3 (N4908, N4906, N453, N3547);
nor NOR4 (N4909, N4908, N2455, N3438, N2494);
nand NAND2 (N4910, N4907, N3385);
nor NOR3 (N4911, N4873, N246, N3649);
nor NOR4 (N4912, N4905, N4080, N162, N1248);
or OR4 (N4913, N4890, N3579, N1476, N2066);
not NOT1 (N4914, N4904);
xor XOR2 (N4915, N4902, N1943);
nand NAND4 (N4916, N4913, N290, N2414, N37);
or OR4 (N4917, N4894, N1789, N3482, N3333);
nand NAND3 (N4918, N4915, N3926, N3641);
nand NAND3 (N4919, N4881, N832, N2409);
xor XOR2 (N4920, N4916, N4851);
nand NAND4 (N4921, N4917, N922, N513, N1906);
nand NAND3 (N4922, N4911, N373, N2572);
nand NAND2 (N4923, N4921, N1394);
buf BUF1 (N4924, N4918);
xor XOR2 (N4925, N4889, N4048);
not NOT1 (N4926, N4919);
and AND3 (N4927, N4909, N1403, N4020);
not NOT1 (N4928, N4926);
nand NAND4 (N4929, N4923, N1141, N403, N3388);
nor NOR3 (N4930, N4924, N2624, N1824);
nor NOR2 (N4931, N4920, N3273);
and AND2 (N4932, N4929, N2408);
not NOT1 (N4933, N4932);
nor NOR3 (N4934, N4910, N2336, N2071);
buf BUF1 (N4935, N4925);
nand NAND2 (N4936, N4912, N64);
nor NOR4 (N4937, N4927, N3055, N2238, N894);
not NOT1 (N4938, N4922);
nand NAND3 (N4939, N4934, N2328, N2544);
or OR4 (N4940, N4931, N97, N2494, N3351);
nand NAND4 (N4941, N4930, N1691, N875, N3552);
and AND4 (N4942, N4935, N3959, N2136, N1494);
buf BUF1 (N4943, N4928);
xor XOR2 (N4944, N4938, N2366);
xor XOR2 (N4945, N4942, N224);
xor XOR2 (N4946, N4939, N891);
or OR2 (N4947, N4945, N3542);
not NOT1 (N4948, N4940);
not NOT1 (N4949, N4937);
nand NAND3 (N4950, N4944, N662, N1167);
nand NAND4 (N4951, N4936, N2791, N3297, N926);
not NOT1 (N4952, N4948);
buf BUF1 (N4953, N4949);
buf BUF1 (N4954, N4943);
nor NOR2 (N4955, N4950, N4512);
nor NOR4 (N4956, N4953, N3894, N4914, N2679);
not NOT1 (N4957, N2508);
and AND2 (N4958, N4946, N4002);
or OR2 (N4959, N4955, N1457);
xor XOR2 (N4960, N4956, N1763);
or OR3 (N4961, N4947, N4750, N393);
or OR2 (N4962, N4958, N224);
or OR4 (N4963, N4962, N4951, N2970, N4462);
buf BUF1 (N4964, N4146);
not NOT1 (N4965, N4963);
not NOT1 (N4966, N4960);
buf BUF1 (N4967, N4957);
not NOT1 (N4968, N4952);
xor XOR2 (N4969, N4964, N13);
nor NOR2 (N4970, N4966, N511);
or OR4 (N4971, N4941, N4620, N1709, N4068);
not NOT1 (N4972, N4968);
nand NAND3 (N4973, N4971, N3451, N932);
nor NOR3 (N4974, N4954, N2912, N4300);
and AND3 (N4975, N4959, N95, N3951);
nor NOR2 (N4976, N4972, N1722);
not NOT1 (N4977, N4975);
or OR3 (N4978, N4965, N3329, N1141);
nor NOR4 (N4979, N4969, N1710, N4027, N1113);
and AND3 (N4980, N4961, N3286, N1489);
buf BUF1 (N4981, N4979);
nor NOR3 (N4982, N4933, N431, N505);
nand NAND3 (N4983, N4982, N310, N4982);
buf BUF1 (N4984, N4976);
nand NAND2 (N4985, N4984, N4806);
buf BUF1 (N4986, N4978);
not NOT1 (N4987, N4970);
and AND2 (N4988, N4985, N3221);
xor XOR2 (N4989, N4974, N4208);
not NOT1 (N4990, N4983);
not NOT1 (N4991, N4977);
or OR2 (N4992, N4988, N3245);
not NOT1 (N4993, N4992);
buf BUF1 (N4994, N4986);
or OR2 (N4995, N4990, N346);
xor XOR2 (N4996, N4967, N4993);
xor XOR2 (N4997, N2064, N4728);
and AND2 (N4998, N4989, N2389);
not NOT1 (N4999, N4973);
or OR2 (N5000, N4980, N3783);
or OR2 (N5001, N4999, N3623);
buf BUF1 (N5002, N4996);
buf BUF1 (N5003, N4998);
nor NOR3 (N5004, N5003, N4408, N919);
buf BUF1 (N5005, N4981);
nor NOR3 (N5006, N4991, N1450, N3292);
nand NAND2 (N5007, N5001, N1574);
not NOT1 (N5008, N5007);
xor XOR2 (N5009, N4995, N3450);
buf BUF1 (N5010, N5009);
nand NAND2 (N5011, N5010, N3420);
xor XOR2 (N5012, N5002, N502);
and AND3 (N5013, N5006, N127, N4859);
not NOT1 (N5014, N4997);
or OR3 (N5015, N5011, N4885, N4967);
and AND4 (N5016, N5012, N1467, N549, N1643);
nor NOR4 (N5017, N5000, N2096, N4913, N790);
buf BUF1 (N5018, N5013);
or OR2 (N5019, N5016, N2320);
not NOT1 (N5020, N5004);
buf BUF1 (N5021, N5005);
nand NAND2 (N5022, N4987, N1922);
not NOT1 (N5023, N5021);
and AND3 (N5024, N5020, N1798, N2471);
xor XOR2 (N5025, N5017, N2869);
or OR3 (N5026, N5025, N4164, N2286);
not NOT1 (N5027, N5014);
not NOT1 (N5028, N5023);
nor NOR4 (N5029, N5022, N3311, N1882, N4716);
xor XOR2 (N5030, N4994, N4008);
buf BUF1 (N5031, N5029);
xor XOR2 (N5032, N5019, N3647);
nor NOR4 (N5033, N5018, N3552, N3318, N3732);
and AND2 (N5034, N5026, N4478);
nand NAND2 (N5035, N5032, N3289);
not NOT1 (N5036, N5024);
or OR4 (N5037, N5035, N370, N4788, N1687);
nand NAND4 (N5038, N5037, N2430, N4558, N235);
xor XOR2 (N5039, N5031, N984);
xor XOR2 (N5040, N5036, N4526);
or OR3 (N5041, N5008, N2253, N4040);
or OR4 (N5042, N5041, N935, N1082, N2552);
or OR3 (N5043, N5015, N1165, N762);
nor NOR3 (N5044, N5034, N159, N2936);
nor NOR4 (N5045, N5043, N4983, N2261, N2291);
buf BUF1 (N5046, N5038);
nand NAND4 (N5047, N5040, N3014, N4013, N2640);
not NOT1 (N5048, N5045);
nand NAND3 (N5049, N5039, N362, N4929);
and AND4 (N5050, N5049, N674, N4971, N1088);
and AND3 (N5051, N5046, N1427, N613);
nand NAND3 (N5052, N5030, N2805, N771);
and AND2 (N5053, N5028, N640);
nand NAND4 (N5054, N5052, N748, N860, N3592);
or OR4 (N5055, N5042, N4024, N2215, N4139);
not NOT1 (N5056, N5054);
nand NAND4 (N5057, N5033, N4884, N1330, N5018);
nand NAND4 (N5058, N5051, N747, N3222, N2158);
and AND4 (N5059, N5048, N2290, N4653, N5043);
or OR3 (N5060, N5059, N573, N541);
buf BUF1 (N5061, N5050);
nor NOR2 (N5062, N5055, N1176);
xor XOR2 (N5063, N5061, N2531);
or OR4 (N5064, N5062, N1595, N2651, N147);
and AND3 (N5065, N5044, N2376, N4048);
buf BUF1 (N5066, N5056);
nor NOR2 (N5067, N5053, N3048);
buf BUF1 (N5068, N5060);
nand NAND3 (N5069, N5064, N3947, N1611);
nand NAND3 (N5070, N5067, N3922, N62);
nand NAND4 (N5071, N5068, N795, N2872, N1311);
and AND4 (N5072, N5071, N4719, N3743, N2308);
buf BUF1 (N5073, N5066);
not NOT1 (N5074, N5063);
nor NOR4 (N5075, N5072, N4242, N3958, N651);
nand NAND2 (N5076, N5073, N540);
nand NAND2 (N5077, N5065, N4377);
and AND2 (N5078, N5058, N2491);
xor XOR2 (N5079, N5077, N5019);
or OR4 (N5080, N5075, N2763, N1937, N153);
xor XOR2 (N5081, N5069, N1447);
or OR3 (N5082, N5027, N578, N681);
buf BUF1 (N5083, N5047);
nor NOR2 (N5084, N5074, N3883);
nand NAND2 (N5085, N5076, N3981);
and AND3 (N5086, N5079, N4825, N4448);
nand NAND4 (N5087, N5082, N2991, N2857, N898);
buf BUF1 (N5088, N5083);
not NOT1 (N5089, N5086);
nor NOR4 (N5090, N5078, N244, N117, N4762);
or OR2 (N5091, N5088, N3388);
buf BUF1 (N5092, N5084);
buf BUF1 (N5093, N5070);
not NOT1 (N5094, N5090);
xor XOR2 (N5095, N5091, N1952);
xor XOR2 (N5096, N5093, N366);
not NOT1 (N5097, N5089);
nor NOR3 (N5098, N5094, N173, N4999);
buf BUF1 (N5099, N5080);
or OR4 (N5100, N5098, N5013, N4984, N2751);
not NOT1 (N5101, N5092);
and AND3 (N5102, N5096, N4658, N589);
or OR2 (N5103, N5085, N3048);
xor XOR2 (N5104, N5081, N3067);
not NOT1 (N5105, N5099);
nor NOR2 (N5106, N5102, N4315);
or OR4 (N5107, N5095, N1866, N4387, N1650);
nand NAND2 (N5108, N5107, N1315);
not NOT1 (N5109, N5087);
nor NOR3 (N5110, N5097, N2999, N3984);
and AND2 (N5111, N5057, N4067);
and AND3 (N5112, N5100, N4702, N2753);
buf BUF1 (N5113, N5104);
and AND3 (N5114, N5103, N2839, N4545);
buf BUF1 (N5115, N5110);
buf BUF1 (N5116, N5108);
not NOT1 (N5117, N5109);
or OR4 (N5118, N5116, N3652, N1811, N4458);
buf BUF1 (N5119, N5117);
or OR2 (N5120, N5119, N3649);
not NOT1 (N5121, N5111);
and AND2 (N5122, N5120, N1337);
xor XOR2 (N5123, N5106, N1804);
xor XOR2 (N5124, N5113, N2721);
or OR3 (N5125, N5114, N3446, N514);
or OR4 (N5126, N5122, N2959, N2342, N4029);
nor NOR2 (N5127, N5123, N2775);
and AND2 (N5128, N5121, N331);
nor NOR2 (N5129, N5124, N2423);
nor NOR3 (N5130, N5125, N1500, N3492);
and AND4 (N5131, N5118, N3118, N4785, N3388);
nand NAND2 (N5132, N5127, N2800);
or OR2 (N5133, N5126, N1648);
nor NOR2 (N5134, N5129, N3871);
not NOT1 (N5135, N5105);
nor NOR2 (N5136, N5130, N4918);
not NOT1 (N5137, N5133);
or OR3 (N5138, N5136, N1217, N212);
nand NAND4 (N5139, N5101, N657, N158, N1883);
nor NOR3 (N5140, N5134, N706, N1900);
nand NAND4 (N5141, N5132, N2676, N4679, N1533);
xor XOR2 (N5142, N5115, N3324);
not NOT1 (N5143, N5131);
buf BUF1 (N5144, N5128);
nand NAND4 (N5145, N5139, N2524, N3002, N977);
and AND3 (N5146, N5144, N2564, N22);
nor NOR4 (N5147, N5138, N3205, N2031, N4645);
or OR2 (N5148, N5143, N932);
nand NAND4 (N5149, N5145, N2265, N3466, N1064);
buf BUF1 (N5150, N5149);
nor NOR2 (N5151, N5148, N3329);
nand NAND2 (N5152, N5140, N390);
or OR2 (N5153, N5142, N2847);
and AND2 (N5154, N5146, N78);
nor NOR3 (N5155, N5141, N4376, N2975);
buf BUF1 (N5156, N5153);
not NOT1 (N5157, N5156);
nor NOR4 (N5158, N5155, N3915, N163, N4728);
and AND3 (N5159, N5154, N3308, N1606);
xor XOR2 (N5160, N5150, N3656);
or OR4 (N5161, N5159, N125, N3842, N2185);
nor NOR4 (N5162, N5112, N2973, N1062, N1833);
nor NOR4 (N5163, N5162, N3332, N2086, N2728);
and AND4 (N5164, N5161, N1518, N968, N1162);
not NOT1 (N5165, N5158);
not NOT1 (N5166, N5147);
not NOT1 (N5167, N5164);
xor XOR2 (N5168, N5137, N2358);
buf BUF1 (N5169, N5167);
or OR4 (N5170, N5168, N1260, N2463, N1442);
nor NOR2 (N5171, N5169, N1527);
and AND2 (N5172, N5166, N4103);
nor NOR3 (N5173, N5135, N2316, N3810);
and AND4 (N5174, N5160, N5021, N1797, N1710);
or OR3 (N5175, N5173, N1157, N5156);
or OR3 (N5176, N5157, N2275, N690);
xor XOR2 (N5177, N5152, N1736);
not NOT1 (N5178, N5176);
or OR4 (N5179, N5170, N69, N560, N3624);
nand NAND3 (N5180, N5172, N3952, N3012);
and AND4 (N5181, N5151, N1819, N3322, N3501);
nand NAND4 (N5182, N5179, N3550, N713, N4631);
or OR3 (N5183, N5163, N4810, N114);
not NOT1 (N5184, N5180);
nor NOR4 (N5185, N5171, N3647, N622, N132);
nor NOR4 (N5186, N5178, N3129, N1707, N474);
and AND3 (N5187, N5181, N2688, N1494);
not NOT1 (N5188, N5187);
nand NAND2 (N5189, N5185, N3205);
nand NAND4 (N5190, N5175, N3622, N3323, N3910);
buf BUF1 (N5191, N5177);
nand NAND2 (N5192, N5186, N4487);
nor NOR4 (N5193, N5182, N4788, N2948, N1456);
buf BUF1 (N5194, N5189);
buf BUF1 (N5195, N5192);
nor NOR4 (N5196, N5191, N4244, N3201, N2636);
nand NAND2 (N5197, N5194, N947);
and AND4 (N5198, N5190, N3234, N588, N481);
nand NAND3 (N5199, N5193, N2217, N5068);
nand NAND3 (N5200, N5199, N4210, N432);
nand NAND4 (N5201, N5197, N4905, N4526, N2475);
nor NOR2 (N5202, N5196, N2782);
not NOT1 (N5203, N5165);
and AND2 (N5204, N5195, N1564);
nor NOR3 (N5205, N5183, N1101, N4444);
and AND3 (N5206, N5203, N1064, N2584);
nand NAND3 (N5207, N5204, N3596, N3191);
not NOT1 (N5208, N5198);
not NOT1 (N5209, N5188);
buf BUF1 (N5210, N5174);
buf BUF1 (N5211, N5207);
nor NOR4 (N5212, N5205, N4802, N643, N1823);
nor NOR4 (N5213, N5212, N1435, N5098, N4685);
not NOT1 (N5214, N5201);
or OR3 (N5215, N5211, N1746, N271);
and AND3 (N5216, N5209, N3452, N246);
not NOT1 (N5217, N5210);
nand NAND4 (N5218, N5216, N4250, N3342, N2120);
nand NAND4 (N5219, N5214, N424, N2226, N682);
xor XOR2 (N5220, N5208, N727);
not NOT1 (N5221, N5219);
xor XOR2 (N5222, N5221, N3848);
and AND4 (N5223, N5215, N2548, N3535, N1106);
and AND4 (N5224, N5220, N2446, N4478, N4024);
xor XOR2 (N5225, N5206, N4841);
not NOT1 (N5226, N5222);
xor XOR2 (N5227, N5184, N2165);
buf BUF1 (N5228, N5226);
nand NAND3 (N5229, N5218, N2739, N3008);
or OR4 (N5230, N5213, N4920, N4724, N3016);
xor XOR2 (N5231, N5230, N1259);
or OR2 (N5232, N5225, N2962);
not NOT1 (N5233, N5228);
not NOT1 (N5234, N5223);
xor XOR2 (N5235, N5231, N4829);
or OR4 (N5236, N5229, N1882, N4580, N577);
and AND4 (N5237, N5236, N2256, N2211, N475);
xor XOR2 (N5238, N5202, N1212);
buf BUF1 (N5239, N5217);
buf BUF1 (N5240, N5200);
nand NAND3 (N5241, N5234, N3905, N3546);
nand NAND4 (N5242, N5235, N1784, N1383, N3177);
not NOT1 (N5243, N5237);
nor NOR3 (N5244, N5239, N1053, N1282);
nor NOR4 (N5245, N5240, N1473, N1976, N337);
nor NOR2 (N5246, N5224, N4185);
nor NOR3 (N5247, N5245, N4431, N363);
nor NOR4 (N5248, N5244, N4729, N4722, N3050);
and AND4 (N5249, N5238, N2428, N360, N4309);
and AND2 (N5250, N5241, N3730);
nand NAND2 (N5251, N5233, N1108);
and AND4 (N5252, N5232, N2414, N1767, N1929);
buf BUF1 (N5253, N5249);
xor XOR2 (N5254, N5243, N5217);
and AND2 (N5255, N5252, N2831);
buf BUF1 (N5256, N5227);
xor XOR2 (N5257, N5253, N3435);
not NOT1 (N5258, N5246);
or OR4 (N5259, N5247, N1148, N5152, N3154);
nor NOR4 (N5260, N5250, N453, N3580, N3640);
buf BUF1 (N5261, N5258);
xor XOR2 (N5262, N5242, N4916);
and AND2 (N5263, N5261, N4803);
xor XOR2 (N5264, N5255, N5026);
nor NOR2 (N5265, N5264, N4628);
and AND4 (N5266, N5265, N3491, N1082, N4393);
nand NAND4 (N5267, N5263, N4024, N1146, N2800);
not NOT1 (N5268, N5254);
xor XOR2 (N5269, N5257, N1769);
nor NOR3 (N5270, N5268, N846, N2881);
buf BUF1 (N5271, N5259);
or OR4 (N5272, N5271, N3363, N638, N1604);
or OR2 (N5273, N5266, N5265);
nor NOR3 (N5274, N5269, N3050, N355);
or OR2 (N5275, N5274, N308);
and AND2 (N5276, N5260, N1972);
nand NAND4 (N5277, N5256, N184, N1413, N3611);
nand NAND3 (N5278, N5273, N4233, N5014);
and AND4 (N5279, N5267, N5029, N1370, N1260);
not NOT1 (N5280, N5270);
xor XOR2 (N5281, N5276, N3876);
xor XOR2 (N5282, N5277, N1516);
xor XOR2 (N5283, N5251, N1824);
not NOT1 (N5284, N5282);
not NOT1 (N5285, N5272);
not NOT1 (N5286, N5281);
not NOT1 (N5287, N5283);
nand NAND2 (N5288, N5262, N649);
buf BUF1 (N5289, N5285);
and AND2 (N5290, N5275, N4289);
xor XOR2 (N5291, N5287, N1994);
nor NOR2 (N5292, N5280, N2057);
nand NAND4 (N5293, N5290, N2576, N159, N735);
buf BUF1 (N5294, N5289);
not NOT1 (N5295, N5292);
or OR3 (N5296, N5295, N4114, N1042);
nand NAND3 (N5297, N5293, N5174, N1603);
nor NOR4 (N5298, N5291, N13, N3661, N2667);
nand NAND2 (N5299, N5294, N528);
xor XOR2 (N5300, N5299, N4322);
and AND4 (N5301, N5278, N2694, N108, N3507);
buf BUF1 (N5302, N5286);
nand NAND3 (N5303, N5297, N4616, N4346);
and AND4 (N5304, N5279, N5043, N74, N4216);
nand NAND3 (N5305, N5301, N564, N4836);
and AND2 (N5306, N5302, N1216);
and AND3 (N5307, N5303, N5, N4603);
not NOT1 (N5308, N5248);
buf BUF1 (N5309, N5305);
and AND2 (N5310, N5307, N3061);
or OR2 (N5311, N5309, N4450);
and AND2 (N5312, N5311, N1329);
and AND3 (N5313, N5288, N4975, N2679);
not NOT1 (N5314, N5296);
and AND2 (N5315, N5284, N4313);
not NOT1 (N5316, N5304);
nor NOR4 (N5317, N5313, N850, N334, N4602);
or OR2 (N5318, N5310, N2902);
buf BUF1 (N5319, N5312);
xor XOR2 (N5320, N5306, N1736);
or OR2 (N5321, N5316, N5170);
and AND3 (N5322, N5315, N432, N1840);
or OR2 (N5323, N5300, N344);
or OR3 (N5324, N5319, N3900, N3351);
nor NOR2 (N5325, N5314, N4388);
xor XOR2 (N5326, N5317, N1432);
and AND3 (N5327, N5326, N3509, N385);
nor NOR2 (N5328, N5324, N4289);
xor XOR2 (N5329, N5328, N5051);
or OR4 (N5330, N5320, N1954, N404, N1557);
and AND4 (N5331, N5325, N2213, N1782, N2761);
buf BUF1 (N5332, N5330);
buf BUF1 (N5333, N5327);
and AND4 (N5334, N5318, N5019, N3904, N2964);
and AND2 (N5335, N5333, N3259);
nand NAND3 (N5336, N5335, N4995, N2517);
and AND3 (N5337, N5308, N592, N4475);
nand NAND3 (N5338, N5334, N3596, N4282);
xor XOR2 (N5339, N5298, N2142);
xor XOR2 (N5340, N5332, N5003);
and AND2 (N5341, N5331, N2453);
and AND3 (N5342, N5323, N4295, N1645);
nand NAND3 (N5343, N5321, N3944, N5062);
buf BUF1 (N5344, N5340);
or OR2 (N5345, N5342, N2158);
nand NAND2 (N5346, N5345, N4066);
and AND3 (N5347, N5346, N5336, N4035);
nand NAND4 (N5348, N2704, N4628, N4510, N5340);
xor XOR2 (N5349, N5338, N472);
or OR2 (N5350, N5343, N419);
buf BUF1 (N5351, N5339);
and AND4 (N5352, N5329, N4245, N1791, N4651);
and AND3 (N5353, N5341, N3111, N3776);
and AND3 (N5354, N5344, N5155, N3258);
not NOT1 (N5355, N5350);
buf BUF1 (N5356, N5354);
nor NOR2 (N5357, N5352, N1054);
buf BUF1 (N5358, N5347);
not NOT1 (N5359, N5353);
xor XOR2 (N5360, N5349, N1358);
not NOT1 (N5361, N5322);
or OR2 (N5362, N5357, N5166);
nand NAND4 (N5363, N5359, N2796, N135, N1329);
and AND4 (N5364, N5360, N3519, N1649, N64);
nand NAND3 (N5365, N5355, N4784, N1096);
nor NOR3 (N5366, N5364, N1582, N3888);
not NOT1 (N5367, N5365);
buf BUF1 (N5368, N5366);
or OR2 (N5369, N5368, N3362);
nor NOR4 (N5370, N5363, N1158, N3421, N5351);
xor XOR2 (N5371, N2377, N716);
xor XOR2 (N5372, N5370, N4539);
nor NOR3 (N5373, N5369, N2253, N3852);
nand NAND4 (N5374, N5362, N1140, N1186, N805);
nand NAND2 (N5375, N5361, N282);
nor NOR4 (N5376, N5373, N3058, N2441, N1020);
or OR3 (N5377, N5337, N3630, N3651);
not NOT1 (N5378, N5356);
and AND4 (N5379, N5358, N2149, N1429, N207);
nor NOR3 (N5380, N5378, N2998, N233);
nand NAND4 (N5381, N5377, N4995, N3163, N3956);
xor XOR2 (N5382, N5367, N3076);
nor NOR2 (N5383, N5381, N3726);
nand NAND3 (N5384, N5382, N106, N4112);
nor NOR2 (N5385, N5379, N2464);
nor NOR4 (N5386, N5375, N3450, N4815, N2068);
xor XOR2 (N5387, N5372, N3945);
not NOT1 (N5388, N5385);
nor NOR4 (N5389, N5380, N3253, N3727, N4350);
and AND2 (N5390, N5383, N436);
and AND4 (N5391, N5384, N98, N101, N4370);
or OR3 (N5392, N5374, N2156, N3979);
not NOT1 (N5393, N5391);
xor XOR2 (N5394, N5389, N4185);
and AND3 (N5395, N5393, N3981, N2866);
buf BUF1 (N5396, N5386);
not NOT1 (N5397, N5388);
buf BUF1 (N5398, N5396);
xor XOR2 (N5399, N5395, N3903);
and AND2 (N5400, N5371, N2673);
or OR2 (N5401, N5400, N82);
buf BUF1 (N5402, N5376);
nand NAND4 (N5403, N5392, N2675, N3673, N3474);
xor XOR2 (N5404, N5402, N4226);
xor XOR2 (N5405, N5387, N4395);
and AND4 (N5406, N5348, N3347, N3970, N4304);
xor XOR2 (N5407, N5405, N5046);
or OR4 (N5408, N5401, N4084, N4762, N4247);
buf BUF1 (N5409, N5394);
nor NOR2 (N5410, N5407, N4060);
nand NAND2 (N5411, N5403, N3323);
and AND4 (N5412, N5406, N5115, N3028, N1731);
xor XOR2 (N5413, N5399, N2470);
and AND4 (N5414, N5412, N2217, N4916, N787);
nand NAND2 (N5415, N5413, N891);
nor NOR3 (N5416, N5390, N2215, N1096);
and AND4 (N5417, N5415, N719, N3415, N2457);
not NOT1 (N5418, N5398);
xor XOR2 (N5419, N5409, N2743);
nor NOR2 (N5420, N5419, N3257);
buf BUF1 (N5421, N5404);
not NOT1 (N5422, N5414);
nand NAND2 (N5423, N5422, N2379);
not NOT1 (N5424, N5416);
nand NAND4 (N5425, N5423, N1905, N4674, N3942);
buf BUF1 (N5426, N5425);
nand NAND2 (N5427, N5420, N3896);
and AND3 (N5428, N5418, N56, N3308);
nor NOR4 (N5429, N5408, N2443, N5050, N4621);
xor XOR2 (N5430, N5421, N981);
buf BUF1 (N5431, N5410);
nand NAND3 (N5432, N5417, N5091, N5129);
nor NOR4 (N5433, N5397, N1640, N2232, N1206);
nor NOR3 (N5434, N5432, N4453, N1293);
or OR2 (N5435, N5429, N3120);
buf BUF1 (N5436, N5426);
and AND4 (N5437, N5433, N536, N295, N4624);
and AND3 (N5438, N5436, N20, N2528);
and AND4 (N5439, N5438, N855, N1960, N3286);
and AND3 (N5440, N5424, N85, N1404);
nand NAND4 (N5441, N5428, N1609, N1040, N3827);
nor NOR4 (N5442, N5439, N379, N4397, N2802);
xor XOR2 (N5443, N5434, N3704);
buf BUF1 (N5444, N5411);
xor XOR2 (N5445, N5441, N2043);
nand NAND3 (N5446, N5445, N3454, N4964);
nand NAND4 (N5447, N5427, N4533, N5407, N3330);
nand NAND4 (N5448, N5442, N1993, N4470, N992);
xor XOR2 (N5449, N5430, N4062);
not NOT1 (N5450, N5443);
or OR4 (N5451, N5447, N1030, N3674, N4042);
not NOT1 (N5452, N5449);
and AND3 (N5453, N5450, N27, N2301);
nor NOR3 (N5454, N5448, N4806, N1010);
buf BUF1 (N5455, N5437);
xor XOR2 (N5456, N5444, N1265);
buf BUF1 (N5457, N5455);
nor NOR3 (N5458, N5451, N904, N1705);
or OR3 (N5459, N5458, N1437, N5110);
or OR3 (N5460, N5459, N3082, N2543);
xor XOR2 (N5461, N5460, N981);
and AND3 (N5462, N5440, N1307, N657);
and AND3 (N5463, N5456, N357, N1408);
nor NOR2 (N5464, N5457, N4077);
buf BUF1 (N5465, N5453);
or OR4 (N5466, N5465, N4726, N1585, N4383);
nor NOR2 (N5467, N5431, N1114);
and AND3 (N5468, N5463, N354, N4945);
or OR2 (N5469, N5468, N2266);
nand NAND2 (N5470, N5469, N1150);
and AND2 (N5471, N5446, N939);
xor XOR2 (N5472, N5461, N2510);
and AND2 (N5473, N5467, N4855);
nand NAND4 (N5474, N5454, N2880, N1954, N4540);
not NOT1 (N5475, N5473);
and AND2 (N5476, N5464, N5473);
nand NAND3 (N5477, N5462, N4743, N4742);
not NOT1 (N5478, N5475);
buf BUF1 (N5479, N5452);
buf BUF1 (N5480, N5476);
not NOT1 (N5481, N5477);
not NOT1 (N5482, N5478);
and AND4 (N5483, N5474, N68, N5419, N3143);
nand NAND3 (N5484, N5435, N3820, N3074);
or OR2 (N5485, N5482, N4541);
not NOT1 (N5486, N5481);
nand NAND2 (N5487, N5486, N4588);
nor NOR3 (N5488, N5470, N4095, N1197);
buf BUF1 (N5489, N5471);
nand NAND4 (N5490, N5479, N4993, N4732, N1069);
nand NAND3 (N5491, N5480, N1376, N2260);
xor XOR2 (N5492, N5483, N2773);
xor XOR2 (N5493, N5488, N4798);
xor XOR2 (N5494, N5485, N1431);
and AND2 (N5495, N5466, N2271);
or OR2 (N5496, N5490, N1092);
or OR4 (N5497, N5496, N2571, N563, N2660);
nand NAND2 (N5498, N5495, N1473);
nor NOR2 (N5499, N5487, N2191);
nand NAND4 (N5500, N5491, N4927, N4177, N2990);
not NOT1 (N5501, N5489);
buf BUF1 (N5502, N5484);
and AND4 (N5503, N5492, N1927, N2971, N3633);
not NOT1 (N5504, N5497);
nor NOR4 (N5505, N5498, N5431, N2097, N371);
xor XOR2 (N5506, N5504, N4781);
and AND4 (N5507, N5494, N705, N4790, N2846);
nand NAND4 (N5508, N5500, N2339, N4419, N1631);
or OR4 (N5509, N5499, N3830, N1048, N5289);
buf BUF1 (N5510, N5508);
nand NAND4 (N5511, N5510, N2937, N1523, N5285);
and AND2 (N5512, N5509, N5006);
or OR4 (N5513, N5501, N3474, N1405, N633);
not NOT1 (N5514, N5505);
nor NOR3 (N5515, N5472, N956, N3560);
nor NOR4 (N5516, N5502, N1095, N5109, N1230);
buf BUF1 (N5517, N5512);
nand NAND3 (N5518, N5493, N4942, N2460);
xor XOR2 (N5519, N5517, N2336);
and AND3 (N5520, N5518, N3260, N2894);
nand NAND3 (N5521, N5519, N694, N394);
nand NAND3 (N5522, N5521, N675, N2379);
xor XOR2 (N5523, N5522, N3991);
not NOT1 (N5524, N5523);
buf BUF1 (N5525, N5514);
nand NAND2 (N5526, N5525, N3809);
not NOT1 (N5527, N5513);
nand NAND4 (N5528, N5511, N4678, N758, N337);
buf BUF1 (N5529, N5515);
buf BUF1 (N5530, N5516);
nor NOR4 (N5531, N5530, N3475, N3739, N3515);
buf BUF1 (N5532, N5527);
and AND2 (N5533, N5524, N1171);
and AND2 (N5534, N5526, N3953);
xor XOR2 (N5535, N5506, N4655);
xor XOR2 (N5536, N5534, N561);
and AND3 (N5537, N5535, N4702, N1749);
nor NOR4 (N5538, N5533, N3166, N2826, N5390);
or OR2 (N5539, N5531, N841);
buf BUF1 (N5540, N5528);
buf BUF1 (N5541, N5507);
nor NOR2 (N5542, N5539, N2534);
and AND2 (N5543, N5538, N4832);
xor XOR2 (N5544, N5520, N3048);
nand NAND2 (N5545, N5536, N3656);
nor NOR3 (N5546, N5541, N745, N4279);
nand NAND4 (N5547, N5545, N4161, N2927, N626);
nand NAND4 (N5548, N5546, N4778, N276, N2882);
buf BUF1 (N5549, N5540);
not NOT1 (N5550, N5542);
and AND4 (N5551, N5532, N3436, N1751, N4993);
xor XOR2 (N5552, N5550, N3852);
nor NOR2 (N5553, N5529, N3611);
nand NAND3 (N5554, N5503, N3358, N3116);
buf BUF1 (N5555, N5554);
or OR4 (N5556, N5552, N2842, N285, N3090);
and AND4 (N5557, N5556, N1063, N2097, N697);
nand NAND2 (N5558, N5553, N1531);
or OR2 (N5559, N5549, N1981);
buf BUF1 (N5560, N5558);
or OR2 (N5561, N5551, N3740);
buf BUF1 (N5562, N5547);
nand NAND4 (N5563, N5562, N4484, N1229, N1786);
or OR3 (N5564, N5555, N2982, N4587);
nand NAND3 (N5565, N5544, N3134, N3481);
buf BUF1 (N5566, N5537);
or OR4 (N5567, N5548, N4170, N458, N2661);
nor NOR4 (N5568, N5563, N3584, N5357, N704);
nor NOR4 (N5569, N5567, N327, N4719, N1833);
or OR4 (N5570, N5565, N446, N2890, N3230);
and AND3 (N5571, N5561, N2039, N1312);
and AND2 (N5572, N5559, N2275);
nand NAND4 (N5573, N5568, N1473, N4423, N3102);
buf BUF1 (N5574, N5557);
xor XOR2 (N5575, N5571, N3726);
buf BUF1 (N5576, N5564);
xor XOR2 (N5577, N5573, N1119);
or OR4 (N5578, N5576, N1969, N946, N2856);
not NOT1 (N5579, N5543);
nand NAND3 (N5580, N5560, N208, N2126);
xor XOR2 (N5581, N5578, N5204);
nand NAND2 (N5582, N5574, N3780);
nor NOR4 (N5583, N5581, N3199, N2259, N1429);
buf BUF1 (N5584, N5575);
buf BUF1 (N5585, N5580);
buf BUF1 (N5586, N5569);
buf BUF1 (N5587, N5586);
not NOT1 (N5588, N5566);
buf BUF1 (N5589, N5583);
nor NOR2 (N5590, N5572, N3363);
xor XOR2 (N5591, N5577, N2981);
xor XOR2 (N5592, N5570, N2299);
buf BUF1 (N5593, N5589);
nor NOR2 (N5594, N5584, N2270);
xor XOR2 (N5595, N5587, N977);
buf BUF1 (N5596, N5595);
not NOT1 (N5597, N5593);
or OR2 (N5598, N5590, N24);
not NOT1 (N5599, N5591);
not NOT1 (N5600, N5594);
xor XOR2 (N5601, N5582, N583);
not NOT1 (N5602, N5601);
and AND4 (N5603, N5600, N495, N1481, N1055);
nand NAND2 (N5604, N5603, N1561);
xor XOR2 (N5605, N5588, N863);
xor XOR2 (N5606, N5604, N1703);
buf BUF1 (N5607, N5598);
not NOT1 (N5608, N5585);
nand NAND3 (N5609, N5597, N2919, N199);
or OR2 (N5610, N5596, N946);
nor NOR2 (N5611, N5605, N4738);
nand NAND2 (N5612, N5610, N1166);
not NOT1 (N5613, N5609);
buf BUF1 (N5614, N5599);
xor XOR2 (N5615, N5602, N2987);
and AND2 (N5616, N5615, N4926);
buf BUF1 (N5617, N5592);
buf BUF1 (N5618, N5608);
not NOT1 (N5619, N5618);
xor XOR2 (N5620, N5611, N5396);
buf BUF1 (N5621, N5579);
nor NOR4 (N5622, N5617, N3232, N2789, N1360);
nand NAND2 (N5623, N5619, N1820);
and AND3 (N5624, N5616, N1379, N4681);
or OR2 (N5625, N5613, N4238);
or OR3 (N5626, N5625, N5333, N2458);
nor NOR2 (N5627, N5612, N4980);
xor XOR2 (N5628, N5620, N2806);
not NOT1 (N5629, N5623);
nor NOR3 (N5630, N5626, N4745, N3165);
or OR3 (N5631, N5621, N1912, N1344);
or OR2 (N5632, N5630, N2805);
and AND4 (N5633, N5614, N1619, N1198, N503);
buf BUF1 (N5634, N5606);
xor XOR2 (N5635, N5627, N1957);
xor XOR2 (N5636, N5629, N4405);
and AND4 (N5637, N5631, N479, N3338, N4710);
nand NAND3 (N5638, N5636, N5467, N2535);
or OR3 (N5639, N5635, N4166, N1452);
or OR3 (N5640, N5622, N4890, N3619);
nand NAND3 (N5641, N5624, N4422, N3952);
buf BUF1 (N5642, N5628);
buf BUF1 (N5643, N5639);
or OR2 (N5644, N5634, N5401);
buf BUF1 (N5645, N5633);
or OR4 (N5646, N5640, N4429, N154, N2988);
not NOT1 (N5647, N5637);
not NOT1 (N5648, N5641);
or OR4 (N5649, N5645, N3996, N536, N4465);
xor XOR2 (N5650, N5638, N1070);
xor XOR2 (N5651, N5632, N2111);
nor NOR3 (N5652, N5650, N3615, N2644);
not NOT1 (N5653, N5652);
buf BUF1 (N5654, N5644);
nand NAND2 (N5655, N5654, N2167);
nor NOR4 (N5656, N5651, N4144, N4133, N1925);
nor NOR2 (N5657, N5655, N1805);
or OR2 (N5658, N5642, N4488);
buf BUF1 (N5659, N5657);
xor XOR2 (N5660, N5648, N4316);
not NOT1 (N5661, N5658);
xor XOR2 (N5662, N5607, N5073);
nor NOR3 (N5663, N5659, N1442, N752);
and AND3 (N5664, N5653, N3322, N2959);
and AND3 (N5665, N5660, N3759, N2191);
nor NOR3 (N5666, N5663, N4339, N2464);
nor NOR3 (N5667, N5656, N4509, N1516);
buf BUF1 (N5668, N5647);
nor NOR2 (N5669, N5643, N3046);
nand NAND3 (N5670, N5646, N3025, N4957);
buf BUF1 (N5671, N5665);
and AND2 (N5672, N5670, N3904);
and AND3 (N5673, N5661, N2886, N4794);
not NOT1 (N5674, N5667);
buf BUF1 (N5675, N5664);
or OR3 (N5676, N5673, N3707, N1486);
or OR2 (N5677, N5668, N275);
xor XOR2 (N5678, N5677, N5618);
nand NAND2 (N5679, N5671, N496);
and AND4 (N5680, N5669, N4917, N5110, N1145);
buf BUF1 (N5681, N5666);
and AND3 (N5682, N5649, N459, N246);
nor NOR3 (N5683, N5678, N29, N626);
nor NOR4 (N5684, N5674, N4367, N3434, N4335);
xor XOR2 (N5685, N5672, N3292);
not NOT1 (N5686, N5662);
nor NOR3 (N5687, N5676, N263, N1279);
nor NOR4 (N5688, N5685, N3561, N2768, N1628);
nand NAND3 (N5689, N5683, N2622, N5196);
not NOT1 (N5690, N5675);
and AND3 (N5691, N5680, N1772, N4274);
or OR2 (N5692, N5689, N3026);
nor NOR3 (N5693, N5679, N3044, N842);
nor NOR4 (N5694, N5692, N5629, N5369, N444);
buf BUF1 (N5695, N5688);
not NOT1 (N5696, N5694);
or OR3 (N5697, N5686, N5147, N2260);
xor XOR2 (N5698, N5695, N3073);
or OR4 (N5699, N5684, N1684, N4023, N4819);
xor XOR2 (N5700, N5699, N1869);
buf BUF1 (N5701, N5696);
not NOT1 (N5702, N5701);
buf BUF1 (N5703, N5690);
buf BUF1 (N5704, N5691);
nand NAND2 (N5705, N5697, N3641);
nor NOR4 (N5706, N5702, N1869, N5062, N5126);
not NOT1 (N5707, N5700);
or OR4 (N5708, N5707, N4551, N1294, N261);
nand NAND2 (N5709, N5698, N2512);
nor NOR2 (N5710, N5704, N504);
not NOT1 (N5711, N5705);
and AND2 (N5712, N5687, N656);
nor NOR3 (N5713, N5693, N542, N3325);
nand NAND4 (N5714, N5682, N128, N5266, N2583);
nor NOR3 (N5715, N5703, N333, N4390);
nand NAND2 (N5716, N5712, N1868);
nor NOR2 (N5717, N5716, N4699);
buf BUF1 (N5718, N5708);
nand NAND3 (N5719, N5718, N424, N4244);
not NOT1 (N5720, N5710);
buf BUF1 (N5721, N5711);
xor XOR2 (N5722, N5720, N3668);
nor NOR4 (N5723, N5713, N4783, N4010, N5543);
or OR3 (N5724, N5723, N1847, N4634);
and AND3 (N5725, N5722, N407, N148);
and AND4 (N5726, N5714, N5550, N3997, N111);
nor NOR2 (N5727, N5726, N3881);
xor XOR2 (N5728, N5725, N4144);
nor NOR2 (N5729, N5709, N143);
nor NOR3 (N5730, N5721, N3036, N214);
xor XOR2 (N5731, N5719, N1888);
xor XOR2 (N5732, N5731, N4288);
buf BUF1 (N5733, N5729);
not NOT1 (N5734, N5733);
and AND2 (N5735, N5728, N4062);
not NOT1 (N5736, N5681);
xor XOR2 (N5737, N5706, N1933);
xor XOR2 (N5738, N5715, N1274);
nor NOR2 (N5739, N5730, N5276);
buf BUF1 (N5740, N5735);
not NOT1 (N5741, N5724);
xor XOR2 (N5742, N5741, N1229);
nand NAND2 (N5743, N5738, N4156);
or OR4 (N5744, N5734, N3099, N5379, N5646);
buf BUF1 (N5745, N5732);
nor NOR2 (N5746, N5736, N44);
buf BUF1 (N5747, N5744);
or OR2 (N5748, N5740, N5518);
buf BUF1 (N5749, N5747);
nor NOR3 (N5750, N5745, N2400, N2774);
and AND4 (N5751, N5748, N878, N3057, N740);
and AND3 (N5752, N5750, N3727, N5633);
not NOT1 (N5753, N5746);
or OR4 (N5754, N5752, N4271, N969, N3856);
or OR2 (N5755, N5742, N4157);
nand NAND2 (N5756, N5727, N63);
or OR2 (N5757, N5739, N375);
not NOT1 (N5758, N5755);
and AND2 (N5759, N5758, N171);
and AND3 (N5760, N5717, N4570, N4369);
not NOT1 (N5761, N5737);
or OR3 (N5762, N5754, N2001, N4722);
or OR3 (N5763, N5757, N212, N1319);
nor NOR2 (N5764, N5762, N2328);
buf BUF1 (N5765, N5753);
not NOT1 (N5766, N5764);
and AND3 (N5767, N5760, N2826, N501);
nand NAND3 (N5768, N5767, N1264, N970);
or OR4 (N5769, N5751, N2209, N2471, N3115);
xor XOR2 (N5770, N5743, N5204);
nor NOR2 (N5771, N5763, N4261);
or OR2 (N5772, N5766, N2073);
nor NOR2 (N5773, N5765, N680);
and AND3 (N5774, N5769, N1598, N5398);
buf BUF1 (N5775, N5773);
nor NOR4 (N5776, N5749, N3493, N4928, N2585);
nor NOR2 (N5777, N5771, N3718);
nand NAND2 (N5778, N5756, N967);
nand NAND2 (N5779, N5778, N1);
and AND3 (N5780, N5776, N2975, N463);
nor NOR4 (N5781, N5759, N4552, N2035, N5373);
buf BUF1 (N5782, N5761);
or OR3 (N5783, N5774, N459, N5484);
buf BUF1 (N5784, N5779);
not NOT1 (N5785, N5772);
or OR2 (N5786, N5784, N178);
nor NOR3 (N5787, N5781, N3402, N2205);
not NOT1 (N5788, N5775);
buf BUF1 (N5789, N5768);
or OR4 (N5790, N5777, N2144, N3751, N5786);
not NOT1 (N5791, N2624);
buf BUF1 (N5792, N5770);
buf BUF1 (N5793, N5789);
nor NOR3 (N5794, N5791, N2197, N4961);
xor XOR2 (N5795, N5787, N1998);
nor NOR2 (N5796, N5790, N628);
nor NOR4 (N5797, N5780, N1312, N4180, N4021);
buf BUF1 (N5798, N5783);
nand NAND4 (N5799, N5794, N1729, N3222, N4247);
buf BUF1 (N5800, N5799);
nor NOR3 (N5801, N5792, N4643, N3364);
buf BUF1 (N5802, N5800);
buf BUF1 (N5803, N5798);
nor NOR2 (N5804, N5793, N2966);
nor NOR2 (N5805, N5785, N3716);
buf BUF1 (N5806, N5782);
or OR4 (N5807, N5804, N2537, N1830, N3593);
not NOT1 (N5808, N5797);
or OR2 (N5809, N5795, N1239);
xor XOR2 (N5810, N5806, N1178);
not NOT1 (N5811, N5801);
or OR2 (N5812, N5802, N1764);
buf BUF1 (N5813, N5805);
nand NAND4 (N5814, N5812, N4440, N3575, N5381);
nand NAND2 (N5815, N5809, N1705);
not NOT1 (N5816, N5813);
buf BUF1 (N5817, N5816);
buf BUF1 (N5818, N5814);
not NOT1 (N5819, N5818);
and AND4 (N5820, N5803, N3308, N4724, N2822);
buf BUF1 (N5821, N5811);
or OR3 (N5822, N5808, N1069, N3880);
nor NOR2 (N5823, N5822, N717);
nand NAND4 (N5824, N5817, N2382, N5057, N3874);
and AND4 (N5825, N5819, N3037, N3683, N1109);
buf BUF1 (N5826, N5821);
and AND4 (N5827, N5810, N192, N5423, N3186);
not NOT1 (N5828, N5820);
nor NOR3 (N5829, N5815, N1469, N2399);
not NOT1 (N5830, N5796);
and AND3 (N5831, N5825, N1873, N5479);
and AND2 (N5832, N5823, N923);
buf BUF1 (N5833, N5788);
buf BUF1 (N5834, N5826);
and AND4 (N5835, N5828, N5430, N4486, N5760);
and AND3 (N5836, N5833, N801, N2984);
buf BUF1 (N5837, N5831);
nor NOR3 (N5838, N5829, N6, N4732);
and AND3 (N5839, N5827, N3, N5029);
buf BUF1 (N5840, N5837);
nor NOR3 (N5841, N5834, N5732, N1119);
xor XOR2 (N5842, N5835, N1583);
nand NAND2 (N5843, N5832, N644);
nor NOR2 (N5844, N5840, N3652);
xor XOR2 (N5845, N5838, N608);
nor NOR2 (N5846, N5844, N4339);
nor NOR4 (N5847, N5830, N850, N4102, N621);
and AND4 (N5848, N5824, N3435, N3831, N5645);
buf BUF1 (N5849, N5843);
not NOT1 (N5850, N5836);
and AND4 (N5851, N5848, N2714, N3420, N5481);
nor NOR4 (N5852, N5849, N576, N2733, N3890);
or OR3 (N5853, N5851, N3726, N1158);
or OR4 (N5854, N5807, N3862, N4015, N2502);
nand NAND3 (N5855, N5850, N687, N418);
not NOT1 (N5856, N5842);
or OR2 (N5857, N5839, N3464);
or OR2 (N5858, N5852, N4021);
and AND4 (N5859, N5855, N1473, N5040, N35);
and AND4 (N5860, N5857, N2293, N1907, N2634);
buf BUF1 (N5861, N5847);
nand NAND2 (N5862, N5858, N21);
nor NOR2 (N5863, N5841, N5286);
not NOT1 (N5864, N5845);
nor NOR2 (N5865, N5856, N4540);
and AND2 (N5866, N5854, N4981);
nor NOR4 (N5867, N5846, N4922, N3323, N855);
not NOT1 (N5868, N5864);
and AND2 (N5869, N5861, N5481);
xor XOR2 (N5870, N5860, N3705);
xor XOR2 (N5871, N5869, N2259);
nor NOR4 (N5872, N5867, N983, N5193, N3729);
nand NAND2 (N5873, N5866, N4824);
nor NOR3 (N5874, N5865, N1438, N4663);
and AND3 (N5875, N5872, N2914, N1719);
not NOT1 (N5876, N5874);
buf BUF1 (N5877, N5859);
not NOT1 (N5878, N5870);
nand NAND2 (N5879, N5853, N2376);
or OR2 (N5880, N5877, N2507);
nand NAND2 (N5881, N5873, N2108);
buf BUF1 (N5882, N5862);
xor XOR2 (N5883, N5878, N1190);
not NOT1 (N5884, N5879);
nand NAND4 (N5885, N5881, N2796, N4333, N4717);
and AND3 (N5886, N5885, N787, N2365);
nor NOR3 (N5887, N5880, N2792, N2155);
or OR4 (N5888, N5883, N2042, N1172, N2083);
nor NOR3 (N5889, N5875, N4717, N1277);
buf BUF1 (N5890, N5887);
buf BUF1 (N5891, N5889);
nand NAND4 (N5892, N5886, N3811, N4189, N5529);
nand NAND3 (N5893, N5882, N4557, N990);
xor XOR2 (N5894, N5888, N113);
xor XOR2 (N5895, N5892, N2955);
not NOT1 (N5896, N5893);
nand NAND2 (N5897, N5890, N2411);
nand NAND3 (N5898, N5863, N226, N5136);
and AND2 (N5899, N5895, N3797);
xor XOR2 (N5900, N5899, N4785);
or OR3 (N5901, N5896, N236, N1311);
buf BUF1 (N5902, N5868);
buf BUF1 (N5903, N5884);
buf BUF1 (N5904, N5891);
nor NOR3 (N5905, N5897, N2290, N3315);
and AND3 (N5906, N5900, N4691, N2685);
buf BUF1 (N5907, N5894);
xor XOR2 (N5908, N5876, N3847);
not NOT1 (N5909, N5903);
or OR4 (N5910, N5904, N1005, N180, N4964);
nor NOR4 (N5911, N5901, N3448, N2650, N4466);
nor NOR2 (N5912, N5910, N5559);
nor NOR2 (N5913, N5907, N2155);
and AND3 (N5914, N5908, N1274, N4248);
nand NAND3 (N5915, N5911, N1237, N5756);
and AND3 (N5916, N5905, N1191, N4452);
or OR4 (N5917, N5916, N828, N4982, N4411);
and AND3 (N5918, N5917, N1280, N2711);
nand NAND4 (N5919, N5912, N3304, N3872, N5224);
xor XOR2 (N5920, N5914, N466);
and AND4 (N5921, N5919, N2363, N3951, N2813);
not NOT1 (N5922, N5902);
xor XOR2 (N5923, N5906, N5182);
nand NAND4 (N5924, N5871, N1791, N3728, N3631);
buf BUF1 (N5925, N5915);
nor NOR2 (N5926, N5913, N1771);
or OR2 (N5927, N5920, N3863);
nor NOR2 (N5928, N5927, N3472);
and AND2 (N5929, N5925, N951);
xor XOR2 (N5930, N5928, N5244);
or OR3 (N5931, N5926, N2263, N3073);
nor NOR3 (N5932, N5931, N4768, N2686);
not NOT1 (N5933, N5909);
and AND3 (N5934, N5930, N3314, N2295);
nor NOR2 (N5935, N5924, N3011);
not NOT1 (N5936, N5934);
not NOT1 (N5937, N5936);
or OR2 (N5938, N5918, N4689);
nand NAND3 (N5939, N5929, N803, N4571);
xor XOR2 (N5940, N5938, N5035);
buf BUF1 (N5941, N5932);
nor NOR3 (N5942, N5921, N846, N1902);
not NOT1 (N5943, N5941);
or OR2 (N5944, N5922, N2475);
buf BUF1 (N5945, N5944);
not NOT1 (N5946, N5923);
nand NAND2 (N5947, N5942, N998);
buf BUF1 (N5948, N5945);
or OR4 (N5949, N5943, N1474, N3715, N5533);
xor XOR2 (N5950, N5935, N3658);
buf BUF1 (N5951, N5946);
nand NAND3 (N5952, N5933, N3175, N1010);
not NOT1 (N5953, N5949);
nor NOR2 (N5954, N5950, N1263);
not NOT1 (N5955, N5937);
and AND2 (N5956, N5951, N2300);
or OR4 (N5957, N5948, N1402, N4655, N1978);
xor XOR2 (N5958, N5939, N3447);
or OR3 (N5959, N5955, N3334, N1605);
not NOT1 (N5960, N5947);
and AND4 (N5961, N5952, N2031, N1782, N5112);
xor XOR2 (N5962, N5959, N2499);
nor NOR2 (N5963, N5961, N220);
xor XOR2 (N5964, N5962, N1772);
nand NAND3 (N5965, N5898, N5265, N5272);
nor NOR2 (N5966, N5956, N4493);
nand NAND4 (N5967, N5957, N4185, N3387, N50);
nand NAND3 (N5968, N5954, N3600, N1778);
nor NOR2 (N5969, N5953, N5464);
and AND3 (N5970, N5969, N5769, N2856);
xor XOR2 (N5971, N5940, N4085);
or OR2 (N5972, N5968, N2563);
nor NOR2 (N5973, N5966, N5554);
and AND2 (N5974, N5963, N1920);
buf BUF1 (N5975, N5970);
or OR2 (N5976, N5958, N1778);
not NOT1 (N5977, N5972);
buf BUF1 (N5978, N5976);
nand NAND2 (N5979, N5978, N922);
xor XOR2 (N5980, N5975, N211);
and AND3 (N5981, N5960, N5354, N4580);
nor NOR4 (N5982, N5973, N1888, N5209, N2778);
nor NOR3 (N5983, N5971, N2223, N452);
nand NAND3 (N5984, N5983, N5378, N2773);
or OR3 (N5985, N5965, N1678, N3778);
and AND2 (N5986, N5984, N4131);
not NOT1 (N5987, N5985);
not NOT1 (N5988, N5982);
xor XOR2 (N5989, N5964, N4829);
nor NOR4 (N5990, N5989, N1176, N1640, N4296);
buf BUF1 (N5991, N5977);
buf BUF1 (N5992, N5986);
not NOT1 (N5993, N5974);
nand NAND3 (N5994, N5992, N2352, N882);
xor XOR2 (N5995, N5980, N407);
and AND4 (N5996, N5990, N3329, N2104, N4753);
nand NAND3 (N5997, N5987, N3330, N4936);
nand NAND3 (N5998, N5997, N498, N3080);
or OR2 (N5999, N5998, N4499);
nor NOR2 (N6000, N5994, N3356);
xor XOR2 (N6001, N5979, N4756);
nand NAND3 (N6002, N5999, N920, N3526);
and AND4 (N6003, N5995, N5374, N4554, N4832);
or OR4 (N6004, N6000, N313, N2843, N3222);
and AND4 (N6005, N6002, N4044, N1659, N4921);
nand NAND2 (N6006, N5967, N4362);
nor NOR4 (N6007, N6006, N5919, N1220, N2596);
nand NAND2 (N6008, N6001, N5882);
xor XOR2 (N6009, N6004, N2568);
nor NOR3 (N6010, N5993, N1101, N4127);
buf BUF1 (N6011, N6005);
nand NAND3 (N6012, N5991, N95, N5176);
nand NAND4 (N6013, N6010, N3498, N5256, N1765);
nand NAND2 (N6014, N6009, N4192);
buf BUF1 (N6015, N6013);
buf BUF1 (N6016, N5981);
xor XOR2 (N6017, N6008, N3029);
buf BUF1 (N6018, N6015);
and AND2 (N6019, N6012, N3347);
xor XOR2 (N6020, N6003, N1680);
or OR4 (N6021, N6019, N2496, N3463, N3611);
nand NAND4 (N6022, N5988, N1477, N2036, N4272);
and AND4 (N6023, N6020, N4506, N108, N4365);
and AND3 (N6024, N6007, N4001, N5279);
nand NAND4 (N6025, N6011, N1433, N5405, N3594);
buf BUF1 (N6026, N6024);
nor NOR4 (N6027, N6018, N5884, N3648, N1245);
nand NAND2 (N6028, N6021, N2089);
and AND4 (N6029, N6022, N4486, N3189, N1229);
and AND2 (N6030, N5996, N1617);
xor XOR2 (N6031, N6030, N5262);
nor NOR3 (N6032, N6026, N588, N3469);
not NOT1 (N6033, N6031);
nand NAND2 (N6034, N6017, N5919);
or OR4 (N6035, N6014, N3559, N1407, N1154);
and AND3 (N6036, N6029, N2091, N4493);
nor NOR3 (N6037, N6025, N179, N5842);
xor XOR2 (N6038, N6034, N1520);
or OR3 (N6039, N6033, N3545, N3227);
buf BUF1 (N6040, N6032);
nor NOR4 (N6041, N6037, N1615, N3738, N5172);
or OR2 (N6042, N6016, N1138);
not NOT1 (N6043, N6041);
nor NOR3 (N6044, N6038, N5330, N2920);
nor NOR2 (N6045, N6040, N5501);
buf BUF1 (N6046, N6039);
nand NAND3 (N6047, N6023, N4631, N5915);
or OR2 (N6048, N6045, N1562);
xor XOR2 (N6049, N6035, N4367);
buf BUF1 (N6050, N6028);
not NOT1 (N6051, N6043);
buf BUF1 (N6052, N6036);
nand NAND3 (N6053, N6049, N714, N4263);
and AND2 (N6054, N6053, N1785);
xor XOR2 (N6055, N6048, N230);
or OR3 (N6056, N6051, N5466, N2320);
nand NAND4 (N6057, N6046, N2273, N2266, N6009);
and AND2 (N6058, N6055, N530);
xor XOR2 (N6059, N6054, N184);
nand NAND3 (N6060, N6027, N1461, N1016);
nor NOR4 (N6061, N6042, N4651, N2119, N1795);
and AND3 (N6062, N6057, N4153, N3181);
nand NAND2 (N6063, N6059, N1686);
not NOT1 (N6064, N6063);
and AND2 (N6065, N6058, N4956);
buf BUF1 (N6066, N6050);
xor XOR2 (N6067, N6065, N2533);
not NOT1 (N6068, N6064);
not NOT1 (N6069, N6068);
and AND2 (N6070, N6067, N5582);
xor XOR2 (N6071, N6047, N2789);
xor XOR2 (N6072, N6061, N782);
or OR3 (N6073, N6069, N62, N903);
and AND2 (N6074, N6066, N4686);
xor XOR2 (N6075, N6073, N4913);
or OR3 (N6076, N6074, N3819, N3006);
xor XOR2 (N6077, N6060, N2212);
and AND4 (N6078, N6062, N316, N5453, N3963);
buf BUF1 (N6079, N6077);
or OR4 (N6080, N6052, N5686, N3691, N5802);
nand NAND2 (N6081, N6056, N126);
not NOT1 (N6082, N6076);
nor NOR2 (N6083, N6080, N6082);
buf BUF1 (N6084, N3886);
buf BUF1 (N6085, N6071);
not NOT1 (N6086, N6079);
and AND2 (N6087, N6083, N5125);
and AND4 (N6088, N6084, N302, N1676, N3757);
nand NAND4 (N6089, N6081, N4206, N3751, N4804);
xor XOR2 (N6090, N6044, N1521);
nor NOR4 (N6091, N6075, N2574, N2934, N786);
and AND3 (N6092, N6088, N2301, N6067);
not NOT1 (N6093, N6092);
buf BUF1 (N6094, N6091);
not NOT1 (N6095, N6085);
and AND3 (N6096, N6078, N4519, N327);
nor NOR2 (N6097, N6086, N5473);
nor NOR4 (N6098, N6089, N2148, N790, N2822);
or OR4 (N6099, N6095, N2075, N5636, N544);
xor XOR2 (N6100, N6087, N1683);
and AND3 (N6101, N6094, N4880, N491);
nor NOR3 (N6102, N6072, N5539, N275);
and AND2 (N6103, N6102, N4782);
or OR4 (N6104, N6097, N389, N1584, N6001);
nor NOR4 (N6105, N6090, N2040, N2975, N3032);
nor NOR2 (N6106, N6101, N5367);
xor XOR2 (N6107, N6103, N401);
nor NOR3 (N6108, N6105, N2742, N5253);
not NOT1 (N6109, N6099);
not NOT1 (N6110, N6108);
not NOT1 (N6111, N6093);
not NOT1 (N6112, N6104);
and AND4 (N6113, N6100, N2693, N4591, N2981);
nand NAND3 (N6114, N6113, N4563, N5793);
nor NOR4 (N6115, N6107, N2044, N5465, N3462);
buf BUF1 (N6116, N6070);
or OR3 (N6117, N6111, N4271, N3262);
nand NAND3 (N6118, N6106, N893, N6041);
nor NOR3 (N6119, N6109, N932, N2773);
buf BUF1 (N6120, N6110);
nor NOR2 (N6121, N6114, N3071);
buf BUF1 (N6122, N6117);
not NOT1 (N6123, N6115);
nand NAND2 (N6124, N6121, N5722);
nor NOR2 (N6125, N6124, N2217);
or OR4 (N6126, N6125, N2039, N4472, N3088);
not NOT1 (N6127, N6126);
and AND4 (N6128, N6123, N4698, N1841, N2906);
or OR3 (N6129, N6098, N611, N1509);
xor XOR2 (N6130, N6122, N2891);
nand NAND4 (N6131, N6120, N2755, N5198, N1297);
nand NAND3 (N6132, N6112, N1575, N3162);
xor XOR2 (N6133, N6096, N4535);
not NOT1 (N6134, N6127);
not NOT1 (N6135, N6128);
or OR4 (N6136, N6119, N1745, N3056, N4619);
xor XOR2 (N6137, N6131, N158);
or OR2 (N6138, N6132, N2148);
or OR3 (N6139, N6118, N3062, N5292);
nor NOR2 (N6140, N6138, N5804);
nand NAND2 (N6141, N6135, N433);
xor XOR2 (N6142, N6137, N5400);
buf BUF1 (N6143, N6142);
xor XOR2 (N6144, N6140, N5490);
nand NAND4 (N6145, N6139, N1830, N748, N2871);
nor NOR2 (N6146, N6141, N5530);
xor XOR2 (N6147, N6143, N2086);
or OR2 (N6148, N6133, N5873);
xor XOR2 (N6149, N6130, N996);
not NOT1 (N6150, N6148);
buf BUF1 (N6151, N6147);
and AND2 (N6152, N6146, N4508);
nand NAND3 (N6153, N6136, N4220, N3929);
nor NOR2 (N6154, N6151, N4490);
and AND4 (N6155, N6152, N4707, N2131, N3704);
not NOT1 (N6156, N6129);
or OR4 (N6157, N6145, N1356, N5403, N2847);
nand NAND2 (N6158, N6155, N1322);
not NOT1 (N6159, N6153);
nor NOR3 (N6160, N6144, N4169, N1027);
nor NOR2 (N6161, N6150, N3879);
nor NOR2 (N6162, N6134, N1186);
and AND4 (N6163, N6154, N3179, N4390, N5727);
xor XOR2 (N6164, N6157, N1900);
nor NOR3 (N6165, N6161, N5568, N1332);
nand NAND3 (N6166, N6160, N202, N5076);
nor NOR4 (N6167, N6156, N2192, N574, N3511);
not NOT1 (N6168, N6167);
nand NAND3 (N6169, N6162, N2217, N1244);
nor NOR4 (N6170, N6169, N3592, N4108, N3427);
nor NOR3 (N6171, N6168, N2912, N4225);
or OR2 (N6172, N6164, N561);
nor NOR4 (N6173, N6149, N3409, N3932, N4297);
buf BUF1 (N6174, N6166);
xor XOR2 (N6175, N6170, N1063);
xor XOR2 (N6176, N6159, N690);
nor NOR4 (N6177, N6174, N1976, N2963, N4171);
and AND2 (N6178, N6116, N120);
not NOT1 (N6179, N6172);
or OR2 (N6180, N6179, N5478);
nor NOR4 (N6181, N6171, N5514, N5018, N1553);
xor XOR2 (N6182, N6176, N682);
buf BUF1 (N6183, N6173);
and AND2 (N6184, N6182, N3037);
buf BUF1 (N6185, N6181);
nor NOR3 (N6186, N6158, N2823, N3321);
xor XOR2 (N6187, N6165, N3458);
nor NOR3 (N6188, N6180, N394, N131);
xor XOR2 (N6189, N6175, N2451);
or OR3 (N6190, N6178, N3816, N1993);
nand NAND3 (N6191, N6177, N4897, N253);
not NOT1 (N6192, N6184);
nor NOR4 (N6193, N6185, N3973, N2721, N620);
or OR4 (N6194, N6191, N6045, N6104, N2089);
not NOT1 (N6195, N6193);
and AND3 (N6196, N6190, N2176, N2638);
xor XOR2 (N6197, N6163, N6097);
nor NOR3 (N6198, N6195, N6038, N1120);
nand NAND3 (N6199, N6186, N6090, N5591);
not NOT1 (N6200, N6189);
or OR3 (N6201, N6194, N3978, N4549);
and AND4 (N6202, N6199, N174, N1485, N5853);
not NOT1 (N6203, N6192);
nor NOR2 (N6204, N6203, N1483);
xor XOR2 (N6205, N6200, N2583);
nand NAND4 (N6206, N6197, N3324, N5021, N4453);
nor NOR4 (N6207, N6188, N3787, N4829, N2554);
not NOT1 (N6208, N6205);
not NOT1 (N6209, N6207);
buf BUF1 (N6210, N6202);
or OR2 (N6211, N6210, N2385);
and AND3 (N6212, N6211, N5090, N2687);
not NOT1 (N6213, N6187);
and AND3 (N6214, N6208, N3635, N5862);
xor XOR2 (N6215, N6213, N4128);
or OR4 (N6216, N6198, N3513, N1231, N1176);
nand NAND4 (N6217, N6209, N217, N2063, N4289);
and AND4 (N6218, N6215, N5153, N2343, N2844);
and AND3 (N6219, N6204, N5326, N4560);
or OR3 (N6220, N6212, N1428, N2516);
buf BUF1 (N6221, N6214);
and AND4 (N6222, N6201, N2624, N112, N987);
and AND3 (N6223, N6196, N3053, N4328);
buf BUF1 (N6224, N6220);
xor XOR2 (N6225, N6217, N1834);
nand NAND2 (N6226, N6183, N1445);
buf BUF1 (N6227, N6218);
xor XOR2 (N6228, N6227, N4294);
nor NOR2 (N6229, N6226, N4387);
not NOT1 (N6230, N6228);
not NOT1 (N6231, N6225);
nand NAND3 (N6232, N6222, N4231, N2596);
xor XOR2 (N6233, N6231, N2260);
xor XOR2 (N6234, N6221, N1276);
not NOT1 (N6235, N6206);
nor NOR4 (N6236, N6230, N2251, N529, N1882);
nor NOR3 (N6237, N6216, N5530, N2568);
buf BUF1 (N6238, N6219);
nand NAND2 (N6239, N6234, N5085);
xor XOR2 (N6240, N6235, N5857);
or OR3 (N6241, N6240, N1085, N4854);
nor NOR2 (N6242, N6232, N1683);
nor NOR4 (N6243, N6229, N1803, N5143, N4086);
xor XOR2 (N6244, N6239, N6026);
nand NAND4 (N6245, N6241, N84, N5203, N3865);
or OR4 (N6246, N6236, N5327, N4063, N1316);
nand NAND3 (N6247, N6243, N4230, N6079);
nand NAND2 (N6248, N6245, N3974);
and AND4 (N6249, N6248, N2737, N6108, N1291);
or OR2 (N6250, N6249, N5543);
and AND4 (N6251, N6237, N6214, N1571, N6127);
nor NOR3 (N6252, N6233, N296, N3892);
buf BUF1 (N6253, N6252);
nand NAND3 (N6254, N6238, N5436, N3606);
xor XOR2 (N6255, N6246, N1573);
or OR3 (N6256, N6255, N1172, N874);
buf BUF1 (N6257, N6251);
nor NOR2 (N6258, N6250, N2018);
and AND3 (N6259, N6242, N1707, N1576);
not NOT1 (N6260, N6223);
xor XOR2 (N6261, N6259, N3343);
nand NAND4 (N6262, N6247, N35, N3130, N6186);
xor XOR2 (N6263, N6224, N1399);
buf BUF1 (N6264, N6244);
nor NOR4 (N6265, N6263, N1290, N5217, N5250);
or OR2 (N6266, N6258, N2218);
nor NOR4 (N6267, N6253, N5572, N736, N2365);
buf BUF1 (N6268, N6264);
xor XOR2 (N6269, N6261, N5873);
not NOT1 (N6270, N6269);
and AND4 (N6271, N6256, N4565, N6024, N3933);
buf BUF1 (N6272, N6257);
not NOT1 (N6273, N6260);
and AND3 (N6274, N6273, N977, N5860);
buf BUF1 (N6275, N6266);
and AND2 (N6276, N6271, N4335);
or OR2 (N6277, N6276, N2108);
not NOT1 (N6278, N6274);
xor XOR2 (N6279, N6278, N5605);
nand NAND2 (N6280, N6267, N3607);
and AND3 (N6281, N6272, N453, N4663);
nand NAND3 (N6282, N6279, N3543, N2536);
not NOT1 (N6283, N6282);
or OR3 (N6284, N6277, N5541, N2231);
xor XOR2 (N6285, N6262, N4381);
and AND3 (N6286, N6281, N3153, N2261);
and AND2 (N6287, N6265, N3614);
nor NOR4 (N6288, N6254, N2300, N29, N2405);
not NOT1 (N6289, N6287);
xor XOR2 (N6290, N6275, N5589);
and AND3 (N6291, N6290, N3051, N849);
xor XOR2 (N6292, N6286, N3070);
buf BUF1 (N6293, N6283);
nand NAND2 (N6294, N6268, N6042);
xor XOR2 (N6295, N6294, N757);
buf BUF1 (N6296, N6292);
buf BUF1 (N6297, N6295);
and AND4 (N6298, N6296, N1881, N1885, N755);
buf BUF1 (N6299, N6284);
not NOT1 (N6300, N6298);
not NOT1 (N6301, N6288);
and AND2 (N6302, N6280, N5976);
not NOT1 (N6303, N6270);
buf BUF1 (N6304, N6285);
or OR4 (N6305, N6289, N2220, N734, N5540);
and AND2 (N6306, N6304, N5684);
buf BUF1 (N6307, N6297);
and AND3 (N6308, N6302, N2675, N5724);
buf BUF1 (N6309, N6308);
xor XOR2 (N6310, N6300, N5607);
buf BUF1 (N6311, N6303);
nor NOR4 (N6312, N6291, N1031, N2601, N3160);
not NOT1 (N6313, N6299);
not NOT1 (N6314, N6310);
nor NOR2 (N6315, N6309, N5416);
or OR4 (N6316, N6315, N3454, N4159, N77);
not NOT1 (N6317, N6305);
nor NOR2 (N6318, N6317, N5936);
nand NAND3 (N6319, N6311, N2646, N4220);
or OR4 (N6320, N6301, N3724, N5980, N2808);
xor XOR2 (N6321, N6293, N1116);
xor XOR2 (N6322, N6314, N5331);
not NOT1 (N6323, N6307);
nand NAND4 (N6324, N6318, N3921, N2517, N5897);
or OR3 (N6325, N6322, N3135, N2923);
or OR3 (N6326, N6323, N4091, N2677);
buf BUF1 (N6327, N6321);
or OR3 (N6328, N6316, N2639, N5785);
buf BUF1 (N6329, N6327);
nand NAND4 (N6330, N6325, N1403, N5413, N73);
buf BUF1 (N6331, N6330);
and AND3 (N6332, N6326, N5565, N1183);
or OR2 (N6333, N6331, N5622);
not NOT1 (N6334, N6306);
or OR4 (N6335, N6312, N3853, N5601, N5795);
buf BUF1 (N6336, N6332);
xor XOR2 (N6337, N6333, N4787);
xor XOR2 (N6338, N6334, N460);
nand NAND4 (N6339, N6338, N340, N5865, N5792);
not NOT1 (N6340, N6328);
xor XOR2 (N6341, N6336, N697);
not NOT1 (N6342, N6340);
xor XOR2 (N6343, N6341, N626);
not NOT1 (N6344, N6335);
nand NAND3 (N6345, N6342, N6139, N457);
nor NOR4 (N6346, N6320, N3369, N3961, N3398);
nor NOR3 (N6347, N6343, N4474, N4901);
not NOT1 (N6348, N6346);
nand NAND2 (N6349, N6344, N789);
or OR4 (N6350, N6348, N1560, N1547, N1614);
or OR2 (N6351, N6324, N4737);
buf BUF1 (N6352, N6339);
nand NAND3 (N6353, N6329, N2102, N2985);
or OR4 (N6354, N6352, N3021, N3099, N504);
nor NOR4 (N6355, N6345, N2494, N3002, N4750);
nor NOR4 (N6356, N6337, N5105, N383, N5230);
xor XOR2 (N6357, N6319, N1438);
or OR3 (N6358, N6356, N5318, N2116);
or OR3 (N6359, N6349, N6169, N5996);
and AND2 (N6360, N6357, N22);
xor XOR2 (N6361, N6354, N2597);
nor NOR2 (N6362, N6359, N106);
nor NOR2 (N6363, N6351, N2069);
and AND3 (N6364, N6355, N4667, N2871);
buf BUF1 (N6365, N6347);
nand NAND2 (N6366, N6365, N4329);
not NOT1 (N6367, N6361);
nor NOR2 (N6368, N6313, N5334);
buf BUF1 (N6369, N6366);
nor NOR3 (N6370, N6362, N3058, N4777);
or OR4 (N6371, N6368, N292, N763, N5892);
nand NAND2 (N6372, N6363, N5883);
xor XOR2 (N6373, N6371, N137);
nand NAND3 (N6374, N6353, N5751, N5034);
nor NOR2 (N6375, N6373, N5186);
buf BUF1 (N6376, N6364);
nor NOR4 (N6377, N6374, N3505, N1283, N1433);
nor NOR3 (N6378, N6370, N5350, N2642);
not NOT1 (N6379, N6375);
or OR3 (N6380, N6379, N4447, N5533);
or OR3 (N6381, N6367, N3153, N1567);
or OR4 (N6382, N6376, N5236, N6011, N5925);
xor XOR2 (N6383, N6369, N6100);
or OR4 (N6384, N6377, N1650, N3755, N631);
buf BUF1 (N6385, N6381);
and AND3 (N6386, N6385, N344, N1088);
nor NOR4 (N6387, N6383, N3240, N1174, N5443);
buf BUF1 (N6388, N6358);
nor NOR2 (N6389, N6360, N4709);
not NOT1 (N6390, N6382);
buf BUF1 (N6391, N6389);
nor NOR2 (N6392, N6391, N4252);
and AND3 (N6393, N6386, N1067, N4915);
not NOT1 (N6394, N6393);
nor NOR3 (N6395, N6394, N6090, N2671);
or OR4 (N6396, N6350, N6233, N3153, N6385);
buf BUF1 (N6397, N6384);
and AND2 (N6398, N6380, N823);
or OR2 (N6399, N6398, N470);
not NOT1 (N6400, N6387);
xor XOR2 (N6401, N6397, N3618);
nand NAND4 (N6402, N6378, N68, N4206, N1557);
buf BUF1 (N6403, N6392);
buf BUF1 (N6404, N6395);
or OR3 (N6405, N6399, N5696, N2829);
and AND2 (N6406, N6390, N3272);
nand NAND3 (N6407, N6372, N6227, N423);
nand NAND2 (N6408, N6405, N5031);
nor NOR3 (N6409, N6403, N4954, N3042);
or OR3 (N6410, N6388, N4540, N4462);
and AND4 (N6411, N6410, N3427, N4231, N4736);
nor NOR2 (N6412, N6409, N5375);
and AND2 (N6413, N6407, N686);
nand NAND4 (N6414, N6400, N4178, N2293, N2228);
nand NAND3 (N6415, N6413, N3238, N3341);
and AND2 (N6416, N6415, N2841);
nand NAND2 (N6417, N6412, N3126);
buf BUF1 (N6418, N6416);
buf BUF1 (N6419, N6411);
buf BUF1 (N6420, N6414);
and AND3 (N6421, N6420, N6095, N1357);
not NOT1 (N6422, N6418);
xor XOR2 (N6423, N6401, N3206);
not NOT1 (N6424, N6419);
not NOT1 (N6425, N6406);
buf BUF1 (N6426, N6396);
nand NAND2 (N6427, N6408, N3182);
and AND3 (N6428, N6404, N5146, N4786);
xor XOR2 (N6429, N6424, N5934);
nor NOR2 (N6430, N6427, N1079);
or OR2 (N6431, N6423, N5886);
nand NAND2 (N6432, N6431, N4785);
nand NAND3 (N6433, N6430, N4431, N4735);
xor XOR2 (N6434, N6433, N2444);
or OR4 (N6435, N6426, N6175, N4201, N965);
nor NOR4 (N6436, N6434, N2597, N3952, N255);
nand NAND4 (N6437, N6432, N196, N5330, N2750);
xor XOR2 (N6438, N6421, N4991);
nand NAND3 (N6439, N6417, N3161, N988);
nand NAND3 (N6440, N6402, N140, N939);
or OR2 (N6441, N6438, N3181);
nand NAND2 (N6442, N6428, N3308);
not NOT1 (N6443, N6437);
nor NOR4 (N6444, N6425, N822, N201, N3514);
and AND4 (N6445, N6444, N1291, N4183, N5653);
xor XOR2 (N6446, N6441, N1420);
nand NAND4 (N6447, N6440, N3103, N1546, N2753);
not NOT1 (N6448, N6439);
or OR2 (N6449, N6446, N210);
nor NOR3 (N6450, N6429, N3936, N881);
buf BUF1 (N6451, N6443);
xor XOR2 (N6452, N6451, N5591);
not NOT1 (N6453, N6435);
buf BUF1 (N6454, N6447);
not NOT1 (N6455, N6454);
buf BUF1 (N6456, N6453);
buf BUF1 (N6457, N6442);
or OR3 (N6458, N6452, N1634, N5395);
not NOT1 (N6459, N6448);
not NOT1 (N6460, N6457);
nand NAND2 (N6461, N6445, N1696);
and AND4 (N6462, N6458, N1533, N1479, N4494);
or OR3 (N6463, N6460, N2794, N3728);
or OR3 (N6464, N6463, N739, N1791);
buf BUF1 (N6465, N6456);
xor XOR2 (N6466, N6461, N1889);
nor NOR4 (N6467, N6422, N895, N3494, N1200);
nand NAND4 (N6468, N6467, N5168, N2122, N3117);
buf BUF1 (N6469, N6464);
nor NOR2 (N6470, N6450, N6338);
not NOT1 (N6471, N6466);
and AND3 (N6472, N6436, N1865, N314);
and AND2 (N6473, N6469, N5078);
nor NOR3 (N6474, N6473, N1692, N4765);
nand NAND2 (N6475, N6465, N754);
nor NOR4 (N6476, N6468, N4065, N2992, N2278);
and AND3 (N6477, N6455, N5105, N1624);
not NOT1 (N6478, N6472);
and AND2 (N6479, N6474, N2865);
nor NOR4 (N6480, N6479, N5077, N5879, N5884);
buf BUF1 (N6481, N6449);
buf BUF1 (N6482, N6480);
not NOT1 (N6483, N6470);
and AND3 (N6484, N6476, N2449, N623);
and AND4 (N6485, N6459, N380, N5161, N3231);
not NOT1 (N6486, N6477);
nand NAND2 (N6487, N6471, N3601);
not NOT1 (N6488, N6487);
not NOT1 (N6489, N6485);
not NOT1 (N6490, N6462);
not NOT1 (N6491, N6475);
buf BUF1 (N6492, N6482);
not NOT1 (N6493, N6492);
xor XOR2 (N6494, N6483, N4750);
nor NOR3 (N6495, N6486, N388, N1250);
nand NAND4 (N6496, N6484, N3030, N847, N2533);
or OR2 (N6497, N6490, N4357);
buf BUF1 (N6498, N6489);
or OR2 (N6499, N6495, N6473);
buf BUF1 (N6500, N6488);
buf BUF1 (N6501, N6481);
buf BUF1 (N6502, N6496);
nor NOR2 (N6503, N6478, N4581);
nor NOR3 (N6504, N6502, N4706, N4192);
or OR4 (N6505, N6499, N4391, N3564, N6054);
not NOT1 (N6506, N6501);
not NOT1 (N6507, N6493);
not NOT1 (N6508, N6504);
buf BUF1 (N6509, N6508);
xor XOR2 (N6510, N6491, N4023);
nor NOR4 (N6511, N6503, N542, N4543, N5968);
nand NAND4 (N6512, N6507, N2596, N3038, N2938);
not NOT1 (N6513, N6497);
or OR4 (N6514, N6498, N4729, N4080, N839);
and AND3 (N6515, N6506, N972, N3068);
and AND4 (N6516, N6513, N4757, N2802, N4412);
not NOT1 (N6517, N6512);
not NOT1 (N6518, N6500);
and AND2 (N6519, N6518, N5846);
not NOT1 (N6520, N6515);
and AND3 (N6521, N6509, N4676, N2669);
nor NOR4 (N6522, N6521, N2448, N119, N6352);
not NOT1 (N6523, N6522);
and AND3 (N6524, N6519, N3067, N2962);
buf BUF1 (N6525, N6511);
not NOT1 (N6526, N6523);
xor XOR2 (N6527, N6524, N219);
not NOT1 (N6528, N6520);
or OR3 (N6529, N6494, N2274, N4253);
and AND2 (N6530, N6529, N5025);
nand NAND2 (N6531, N6526, N2607);
nand NAND3 (N6532, N6505, N626, N2807);
or OR4 (N6533, N6516, N1080, N2675, N2389);
or OR3 (N6534, N6510, N1662, N1193);
not NOT1 (N6535, N6530);
nor NOR3 (N6536, N6535, N3491, N5311);
and AND4 (N6537, N6531, N3469, N1019, N1426);
not NOT1 (N6538, N6537);
nand NAND2 (N6539, N6525, N6318);
and AND2 (N6540, N6514, N4116);
xor XOR2 (N6541, N6534, N202);
or OR2 (N6542, N6532, N3124);
or OR2 (N6543, N6541, N677);
and AND4 (N6544, N6538, N292, N925, N238);
and AND2 (N6545, N6536, N1961);
nor NOR4 (N6546, N6542, N2149, N3190, N680);
nor NOR3 (N6547, N6543, N5887, N1665);
xor XOR2 (N6548, N6546, N2991);
nor NOR4 (N6549, N6544, N4806, N3048, N426);
and AND3 (N6550, N6539, N3253, N6386);
nor NOR2 (N6551, N6550, N4277);
not NOT1 (N6552, N6548);
nor NOR2 (N6553, N6517, N5596);
buf BUF1 (N6554, N6545);
buf BUF1 (N6555, N6553);
or OR4 (N6556, N6540, N2528, N1565, N1065);
nor NOR4 (N6557, N6556, N4033, N2645, N6237);
xor XOR2 (N6558, N6554, N5548);
xor XOR2 (N6559, N6547, N1116);
nand NAND3 (N6560, N6549, N2252, N261);
nor NOR4 (N6561, N6552, N36, N5910, N761);
or OR2 (N6562, N6551, N5896);
not NOT1 (N6563, N6562);
xor XOR2 (N6564, N6561, N1390);
and AND2 (N6565, N6564, N3268);
not NOT1 (N6566, N6527);
nor NOR2 (N6567, N6558, N3039);
buf BUF1 (N6568, N6560);
buf BUF1 (N6569, N6533);
nor NOR2 (N6570, N6559, N4715);
or OR2 (N6571, N6567, N3427);
nand NAND2 (N6572, N6565, N2947);
nand NAND2 (N6573, N6572, N3280);
xor XOR2 (N6574, N6557, N4345);
nor NOR4 (N6575, N6563, N1962, N3740, N5739);
nor NOR4 (N6576, N6568, N6053, N4929, N4935);
or OR4 (N6577, N6571, N2970, N1529, N5029);
nand NAND2 (N6578, N6528, N1645);
not NOT1 (N6579, N6555);
xor XOR2 (N6580, N6573, N163);
nand NAND2 (N6581, N6579, N4912);
not NOT1 (N6582, N6577);
nand NAND3 (N6583, N6574, N699, N687);
or OR3 (N6584, N6569, N369, N3604);
or OR2 (N6585, N6566, N5265);
nand NAND3 (N6586, N6582, N5173, N3129);
xor XOR2 (N6587, N6581, N1243);
and AND3 (N6588, N6585, N504, N3473);
xor XOR2 (N6589, N6580, N462);
nor NOR4 (N6590, N6575, N4320, N44, N2191);
xor XOR2 (N6591, N6583, N92);
buf BUF1 (N6592, N6578);
not NOT1 (N6593, N6587);
buf BUF1 (N6594, N6570);
xor XOR2 (N6595, N6589, N2621);
buf BUF1 (N6596, N6590);
nor NOR4 (N6597, N6586, N1657, N4787, N632);
or OR2 (N6598, N6594, N6188);
buf BUF1 (N6599, N6593);
or OR3 (N6600, N6599, N3769, N3);
or OR4 (N6601, N6596, N1568, N1244, N1055);
nor NOR3 (N6602, N6584, N2336, N5108);
or OR2 (N6603, N6598, N3527);
not NOT1 (N6604, N6597);
or OR4 (N6605, N6600, N3682, N1200, N5982);
nand NAND3 (N6606, N6604, N1267, N5229);
nand NAND2 (N6607, N6591, N5320);
xor XOR2 (N6608, N6606, N1464);
and AND3 (N6609, N6601, N1367, N6182);
nor NOR4 (N6610, N6595, N1994, N2924, N2850);
and AND2 (N6611, N6592, N4315);
not NOT1 (N6612, N6588);
buf BUF1 (N6613, N6603);
nor NOR2 (N6614, N6608, N1847);
xor XOR2 (N6615, N6614, N3736);
and AND4 (N6616, N6576, N5623, N2521, N3282);
nor NOR2 (N6617, N6602, N33);
not NOT1 (N6618, N6611);
nor NOR2 (N6619, N6605, N6208);
xor XOR2 (N6620, N6618, N853);
nor NOR2 (N6621, N6610, N6162);
and AND4 (N6622, N6616, N6337, N5530, N82);
nand NAND3 (N6623, N6609, N5129, N1408);
not NOT1 (N6624, N6617);
nor NOR4 (N6625, N6607, N6398, N6203, N4048);
xor XOR2 (N6626, N6623, N3147);
and AND3 (N6627, N6624, N253, N821);
nor NOR2 (N6628, N6627, N1017);
buf BUF1 (N6629, N6622);
not NOT1 (N6630, N6615);
nand NAND4 (N6631, N6612, N4924, N2238, N1215);
buf BUF1 (N6632, N6620);
nor NOR3 (N6633, N6628, N4491, N5530);
not NOT1 (N6634, N6621);
nand NAND4 (N6635, N6619, N1119, N2104, N6522);
buf BUF1 (N6636, N6625);
not NOT1 (N6637, N6629);
or OR4 (N6638, N6630, N3321, N3374, N348);
xor XOR2 (N6639, N6632, N1752);
not NOT1 (N6640, N6637);
or OR3 (N6641, N6636, N6383, N305);
or OR2 (N6642, N6631, N2634);
or OR4 (N6643, N6638, N3915, N5992, N5365);
not NOT1 (N6644, N6633);
buf BUF1 (N6645, N6613);
or OR3 (N6646, N6645, N2331, N1808);
xor XOR2 (N6647, N6635, N2310);
not NOT1 (N6648, N6634);
xor XOR2 (N6649, N6647, N4182);
or OR2 (N6650, N6639, N213);
not NOT1 (N6651, N6641);
xor XOR2 (N6652, N6643, N4848);
nand NAND3 (N6653, N6642, N2013, N1205);
nand NAND3 (N6654, N6651, N2004, N1476);
or OR4 (N6655, N6646, N3233, N3620, N4254);
xor XOR2 (N6656, N6640, N47);
xor XOR2 (N6657, N6648, N5802);
or OR4 (N6658, N6657, N192, N6576, N4328);
or OR2 (N6659, N6644, N1878);
buf BUF1 (N6660, N6626);
and AND4 (N6661, N6655, N3617, N1922, N5607);
or OR2 (N6662, N6661, N5220);
xor XOR2 (N6663, N6659, N1417);
or OR4 (N6664, N6649, N5966, N601, N4811);
xor XOR2 (N6665, N6660, N6274);
xor XOR2 (N6666, N6650, N5299);
not NOT1 (N6667, N6658);
not NOT1 (N6668, N6665);
nor NOR4 (N6669, N6653, N1639, N4049, N4877);
and AND2 (N6670, N6668, N1167);
or OR2 (N6671, N6670, N2918);
buf BUF1 (N6672, N6664);
buf BUF1 (N6673, N6669);
not NOT1 (N6674, N6666);
and AND3 (N6675, N6663, N4335, N4652);
or OR3 (N6676, N6671, N2876, N1995);
not NOT1 (N6677, N6676);
or OR3 (N6678, N6672, N3080, N4452);
and AND2 (N6679, N6675, N1135);
and AND2 (N6680, N6652, N4425);
xor XOR2 (N6681, N6662, N1774);
not NOT1 (N6682, N6667);
and AND4 (N6683, N6674, N1872, N6480, N3375);
xor XOR2 (N6684, N6683, N4272);
xor XOR2 (N6685, N6682, N5762);
nand NAND2 (N6686, N6679, N4730);
or OR4 (N6687, N6678, N198, N172, N4781);
nor NOR3 (N6688, N6677, N1376, N3227);
nand NAND4 (N6689, N6681, N5465, N1448, N4705);
buf BUF1 (N6690, N6689);
buf BUF1 (N6691, N6688);
buf BUF1 (N6692, N6691);
and AND4 (N6693, N6685, N255, N3899, N563);
not NOT1 (N6694, N6656);
not NOT1 (N6695, N6690);
buf BUF1 (N6696, N6684);
not NOT1 (N6697, N6696);
or OR4 (N6698, N6680, N1699, N2178, N6370);
xor XOR2 (N6699, N6697, N5438);
and AND4 (N6700, N6686, N6380, N6412, N1125);
and AND4 (N6701, N6693, N2202, N5677, N3326);
not NOT1 (N6702, N6673);
buf BUF1 (N6703, N6699);
or OR2 (N6704, N6687, N5819);
not NOT1 (N6705, N6700);
and AND3 (N6706, N6705, N3573, N4346);
buf BUF1 (N6707, N6698);
and AND2 (N6708, N6692, N6546);
xor XOR2 (N6709, N6654, N2447);
and AND4 (N6710, N6708, N2731, N3349, N2113);
buf BUF1 (N6711, N6694);
xor XOR2 (N6712, N6707, N5115);
xor XOR2 (N6713, N6701, N1327);
nand NAND4 (N6714, N6713, N3252, N1599, N2890);
nand NAND2 (N6715, N6710, N3253);
nand NAND3 (N6716, N6712, N2044, N1656);
nor NOR3 (N6717, N6715, N803, N4289);
buf BUF1 (N6718, N6695);
xor XOR2 (N6719, N6714, N593);
nand NAND2 (N6720, N6719, N1853);
xor XOR2 (N6721, N6720, N2270);
nor NOR3 (N6722, N6718, N761, N542);
nor NOR2 (N6723, N6702, N6071);
not NOT1 (N6724, N6722);
nand NAND2 (N6725, N6711, N3879);
nor NOR3 (N6726, N6725, N506, N4972);
buf BUF1 (N6727, N6721);
xor XOR2 (N6728, N6716, N4145);
and AND2 (N6729, N6709, N6344);
buf BUF1 (N6730, N6717);
and AND3 (N6731, N6723, N1961, N2560);
not NOT1 (N6732, N6703);
and AND4 (N6733, N6732, N6552, N4287, N2635);
xor XOR2 (N6734, N6733, N101);
or OR4 (N6735, N6734, N6330, N3775, N4723);
nand NAND4 (N6736, N6704, N2177, N5451, N5806);
nor NOR2 (N6737, N6736, N1022);
nor NOR4 (N6738, N6706, N5138, N6216, N33);
nand NAND3 (N6739, N6730, N1923, N4794);
buf BUF1 (N6740, N6737);
buf BUF1 (N6741, N6726);
nor NOR3 (N6742, N6729, N4690, N5671);
nand NAND4 (N6743, N6724, N1011, N4206, N3221);
not NOT1 (N6744, N6727);
nor NOR3 (N6745, N6741, N3318, N236);
xor XOR2 (N6746, N6735, N4516);
and AND2 (N6747, N6745, N4806);
or OR3 (N6748, N6738, N1100, N179);
and AND4 (N6749, N6728, N488, N5228, N5210);
nor NOR3 (N6750, N6748, N4726, N6690);
nand NAND4 (N6751, N6749, N5629, N4476, N19);
not NOT1 (N6752, N6751);
nor NOR3 (N6753, N6750, N5542, N4267);
nand NAND4 (N6754, N6746, N2145, N6072, N6457);
buf BUF1 (N6755, N6742);
nand NAND4 (N6756, N6740, N3920, N161, N5009);
and AND3 (N6757, N6753, N2894, N3216);
and AND4 (N6758, N6757, N3430, N5491, N3413);
buf BUF1 (N6759, N6758);
buf BUF1 (N6760, N6752);
or OR2 (N6761, N6756, N2462);
buf BUF1 (N6762, N6754);
xor XOR2 (N6763, N6759, N266);
or OR3 (N6764, N6761, N3517, N2046);
xor XOR2 (N6765, N6755, N1783);
not NOT1 (N6766, N6731);
not NOT1 (N6767, N6744);
not NOT1 (N6768, N6760);
not NOT1 (N6769, N6767);
nand NAND4 (N6770, N6765, N1039, N6458, N2976);
xor XOR2 (N6771, N6770, N1324);
or OR4 (N6772, N6762, N5983, N6167, N5918);
buf BUF1 (N6773, N6743);
xor XOR2 (N6774, N6773, N1678);
nand NAND2 (N6775, N6772, N4604);
not NOT1 (N6776, N6739);
or OR2 (N6777, N6769, N5229);
or OR3 (N6778, N6777, N2819, N6265);
xor XOR2 (N6779, N6764, N5789);
nor NOR3 (N6780, N6775, N5851, N1388);
and AND3 (N6781, N6747, N4341, N518);
and AND2 (N6782, N6778, N2739);
not NOT1 (N6783, N6766);
xor XOR2 (N6784, N6771, N1822);
and AND4 (N6785, N6768, N1655, N6510, N2833);
not NOT1 (N6786, N6780);
not NOT1 (N6787, N6785);
or OR3 (N6788, N6776, N5944, N1031);
xor XOR2 (N6789, N6781, N3681);
or OR4 (N6790, N6787, N2306, N4164, N6194);
xor XOR2 (N6791, N6779, N5840);
and AND2 (N6792, N6784, N6507);
not NOT1 (N6793, N6790);
buf BUF1 (N6794, N6791);
nand NAND4 (N6795, N6792, N2095, N2348, N6204);
nand NAND2 (N6796, N6782, N3627);
and AND4 (N6797, N6788, N3463, N6523, N522);
xor XOR2 (N6798, N6797, N6335);
buf BUF1 (N6799, N6774);
xor XOR2 (N6800, N6763, N1010);
buf BUF1 (N6801, N6800);
and AND2 (N6802, N6798, N6149);
nand NAND3 (N6803, N6796, N3823, N3125);
and AND2 (N6804, N6789, N1849);
nor NOR2 (N6805, N6793, N2625);
buf BUF1 (N6806, N6805);
buf BUF1 (N6807, N6806);
not NOT1 (N6808, N6795);
nor NOR4 (N6809, N6799, N3333, N5113, N876);
buf BUF1 (N6810, N6808);
buf BUF1 (N6811, N6783);
or OR4 (N6812, N6807, N5520, N3731, N1069);
not NOT1 (N6813, N6812);
nor NOR2 (N6814, N6786, N301);
nand NAND2 (N6815, N6814, N6172);
and AND2 (N6816, N6813, N4007);
not NOT1 (N6817, N6815);
xor XOR2 (N6818, N6794, N530);
or OR4 (N6819, N6817, N3185, N6764, N2063);
or OR4 (N6820, N6810, N736, N6721, N5019);
not NOT1 (N6821, N6820);
buf BUF1 (N6822, N6804);
nand NAND4 (N6823, N6816, N1946, N5192, N5240);
buf BUF1 (N6824, N6801);
or OR4 (N6825, N6822, N1210, N6248, N758);
not NOT1 (N6826, N6819);
and AND4 (N6827, N6823, N4897, N6240, N2524);
not NOT1 (N6828, N6826);
buf BUF1 (N6829, N6828);
not NOT1 (N6830, N6825);
and AND3 (N6831, N6830, N6501, N131);
nor NOR4 (N6832, N6803, N2346, N4475, N5453);
and AND4 (N6833, N6832, N1613, N3559, N2094);
not NOT1 (N6834, N6829);
nor NOR3 (N6835, N6824, N3117, N6825);
and AND3 (N6836, N6821, N3736, N3982);
buf BUF1 (N6837, N6834);
or OR3 (N6838, N6811, N4590, N2225);
or OR3 (N6839, N6837, N3282, N1297);
nor NOR3 (N6840, N6827, N3974, N4894);
nor NOR3 (N6841, N6839, N5413, N4696);
not NOT1 (N6842, N6833);
nand NAND2 (N6843, N6838, N6757);
nand NAND3 (N6844, N6842, N18, N2506);
buf BUF1 (N6845, N6818);
or OR4 (N6846, N6845, N3046, N2975, N6398);
buf BUF1 (N6847, N6844);
buf BUF1 (N6848, N6841);
xor XOR2 (N6849, N6802, N2538);
and AND3 (N6850, N6843, N3180, N2787);
buf BUF1 (N6851, N6849);
not NOT1 (N6852, N6850);
or OR3 (N6853, N6831, N4726, N5068);
not NOT1 (N6854, N6848);
or OR2 (N6855, N6852, N1420);
nor NOR2 (N6856, N6846, N6667);
nor NOR3 (N6857, N6851, N2408, N2285);
nand NAND2 (N6858, N6840, N2444);
and AND4 (N6859, N6857, N2015, N1497, N2088);
or OR3 (N6860, N6809, N5416, N4135);
xor XOR2 (N6861, N6859, N2610);
not NOT1 (N6862, N6836);
or OR2 (N6863, N6847, N4909);
not NOT1 (N6864, N6860);
buf BUF1 (N6865, N6856);
nor NOR4 (N6866, N6858, N521, N5959, N4368);
nor NOR3 (N6867, N6863, N662, N6390);
xor XOR2 (N6868, N6864, N1015);
not NOT1 (N6869, N6865);
or OR3 (N6870, N6868, N2668, N5035);
buf BUF1 (N6871, N6855);
and AND2 (N6872, N6867, N230);
nor NOR3 (N6873, N6861, N5961, N2942);
nand NAND2 (N6874, N6853, N3613);
or OR2 (N6875, N6862, N6333);
xor XOR2 (N6876, N6835, N2196);
and AND2 (N6877, N6870, N6107);
nand NAND4 (N6878, N6872, N4706, N5591, N6399);
not NOT1 (N6879, N6866);
xor XOR2 (N6880, N6873, N2876);
and AND4 (N6881, N6871, N803, N482, N6686);
nor NOR3 (N6882, N6869, N1446, N2166);
buf BUF1 (N6883, N6878);
nor NOR4 (N6884, N6876, N2323, N3743, N533);
buf BUF1 (N6885, N6854);
nand NAND4 (N6886, N6884, N4639, N6200, N1549);
xor XOR2 (N6887, N6881, N2147);
not NOT1 (N6888, N6887);
buf BUF1 (N6889, N6875);
not NOT1 (N6890, N6889);
and AND2 (N6891, N6885, N422);
or OR3 (N6892, N6883, N5684, N6531);
buf BUF1 (N6893, N6879);
nand NAND3 (N6894, N6880, N114, N3201);
nor NOR3 (N6895, N6893, N3676, N2952);
not NOT1 (N6896, N6874);
nand NAND3 (N6897, N6895, N6779, N883);
not NOT1 (N6898, N6877);
not NOT1 (N6899, N6892);
nor NOR4 (N6900, N6888, N5095, N6645, N5163);
or OR2 (N6901, N6891, N6632);
buf BUF1 (N6902, N6890);
xor XOR2 (N6903, N6898, N4622);
or OR4 (N6904, N6903, N5955, N3657, N4082);
nor NOR2 (N6905, N6894, N5689);
and AND3 (N6906, N6897, N2078, N3742);
not NOT1 (N6907, N6896);
nand NAND2 (N6908, N6907, N3561);
xor XOR2 (N6909, N6901, N4978);
xor XOR2 (N6910, N6906, N1020);
and AND2 (N6911, N6905, N4316);
not NOT1 (N6912, N6910);
not NOT1 (N6913, N6882);
nand NAND4 (N6914, N6899, N2405, N2215, N338);
buf BUF1 (N6915, N6900);
nand NAND4 (N6916, N6904, N5645, N594, N2659);
xor XOR2 (N6917, N6913, N189);
buf BUF1 (N6918, N6917);
and AND2 (N6919, N6908, N4985);
and AND3 (N6920, N6918, N2419, N4990);
nor NOR2 (N6921, N6886, N5441);
nand NAND2 (N6922, N6911, N5330);
and AND2 (N6923, N6916, N5690);
or OR2 (N6924, N6919, N5821);
nand NAND4 (N6925, N6924, N3732, N3211, N4206);
not NOT1 (N6926, N6915);
or OR3 (N6927, N6922, N742, N5948);
nand NAND3 (N6928, N6912, N855, N6701);
nor NOR4 (N6929, N6920, N777, N4805, N4728);
nand NAND4 (N6930, N6921, N3988, N1547, N2557);
or OR4 (N6931, N6925, N5004, N419, N4188);
not NOT1 (N6932, N6929);
and AND2 (N6933, N6914, N4004);
nor NOR4 (N6934, N6902, N6308, N1826, N6532);
nor NOR3 (N6935, N6931, N1066, N3275);
not NOT1 (N6936, N6934);
nand NAND4 (N6937, N6932, N4850, N3820, N780);
not NOT1 (N6938, N6937);
nor NOR2 (N6939, N6927, N4917);
not NOT1 (N6940, N6923);
xor XOR2 (N6941, N6926, N1970);
nand NAND4 (N6942, N6938, N40, N1548, N6272);
buf BUF1 (N6943, N6933);
and AND3 (N6944, N6936, N4843, N392);
or OR2 (N6945, N6939, N3498);
and AND4 (N6946, N6943, N1465, N2115, N200);
nor NOR2 (N6947, N6945, N3554);
and AND3 (N6948, N6935, N5957, N1224);
and AND3 (N6949, N6930, N3146, N826);
not NOT1 (N6950, N6947);
nand NAND2 (N6951, N6948, N4157);
nand NAND2 (N6952, N6946, N5009);
not NOT1 (N6953, N6952);
xor XOR2 (N6954, N6942, N4953);
or OR4 (N6955, N6909, N4714, N1222, N4626);
and AND2 (N6956, N6951, N4885);
and AND2 (N6957, N6955, N4523);
nor NOR2 (N6958, N6941, N6679);
xor XOR2 (N6959, N6949, N2473);
or OR2 (N6960, N6953, N328);
and AND4 (N6961, N6944, N6649, N4086, N1491);
and AND4 (N6962, N6940, N3562, N62, N5393);
nand NAND4 (N6963, N6928, N5902, N2594, N4519);
xor XOR2 (N6964, N6956, N4108);
or OR3 (N6965, N6962, N6710, N2676);
nor NOR4 (N6966, N6954, N201, N6392, N5780);
and AND4 (N6967, N6964, N6155, N3166, N2583);
buf BUF1 (N6968, N6957);
or OR3 (N6969, N6960, N2705, N699);
xor XOR2 (N6970, N6958, N2712);
buf BUF1 (N6971, N6950);
nor NOR2 (N6972, N6967, N171);
or OR2 (N6973, N6971, N2180);
not NOT1 (N6974, N6965);
nor NOR4 (N6975, N6973, N5646, N3014, N4799);
nor NOR4 (N6976, N6970, N2888, N5515, N3046);
nand NAND3 (N6977, N6976, N2201, N4321);
and AND2 (N6978, N6966, N718);
and AND4 (N6979, N6978, N5427, N4172, N4460);
buf BUF1 (N6980, N6961);
xor XOR2 (N6981, N6963, N1697);
buf BUF1 (N6982, N6977);
nand NAND3 (N6983, N6959, N920, N1012);
and AND2 (N6984, N6980, N4301);
nor NOR3 (N6985, N6974, N5843, N3476);
xor XOR2 (N6986, N6982, N1595);
not NOT1 (N6987, N6979);
nor NOR3 (N6988, N6987, N5735, N5535);
not NOT1 (N6989, N6981);
xor XOR2 (N6990, N6968, N2851);
and AND4 (N6991, N6975, N6914, N855, N6300);
xor XOR2 (N6992, N6989, N3909);
nand NAND3 (N6993, N6983, N1322, N5740);
buf BUF1 (N6994, N6991);
xor XOR2 (N6995, N6969, N68);
and AND4 (N6996, N6972, N2820, N4480, N4605);
or OR2 (N6997, N6992, N1531);
nand NAND3 (N6998, N6995, N628, N3518);
buf BUF1 (N6999, N6986);
nand NAND2 (N7000, N6998, N3997);
or OR4 (N7001, N7000, N6245, N3568, N1956);
and AND3 (N7002, N6996, N4745, N349);
and AND4 (N7003, N7001, N4060, N4620, N2129);
nand NAND3 (N7004, N6999, N3862, N3150);
or OR2 (N7005, N6993, N6573);
nor NOR4 (N7006, N6994, N2293, N6127, N3666);
buf BUF1 (N7007, N7006);
and AND2 (N7008, N6997, N1183);
or OR3 (N7009, N7007, N1739, N4626);
buf BUF1 (N7010, N7005);
nand NAND4 (N7011, N6988, N1168, N2325, N3572);
buf BUF1 (N7012, N7009);
nand NAND2 (N7013, N7010, N4811);
nor NOR2 (N7014, N7011, N2072);
buf BUF1 (N7015, N7004);
nand NAND2 (N7016, N7012, N3995);
nor NOR4 (N7017, N6990, N1911, N3653, N4003);
xor XOR2 (N7018, N6984, N5619);
or OR2 (N7019, N7008, N3562);
and AND4 (N7020, N7016, N1956, N4722, N1936);
or OR2 (N7021, N7013, N3142);
nor NOR4 (N7022, N7003, N5032, N5083, N1957);
not NOT1 (N7023, N7021);
or OR4 (N7024, N7018, N3227, N6904, N5276);
nor NOR3 (N7025, N7002, N180, N2951);
not NOT1 (N7026, N7022);
buf BUF1 (N7027, N7017);
nand NAND4 (N7028, N7025, N6199, N3398, N4573);
or OR4 (N7029, N7024, N805, N3054, N1926);
buf BUF1 (N7030, N7014);
xor XOR2 (N7031, N7019, N1609);
xor XOR2 (N7032, N7030, N6373);
not NOT1 (N7033, N7026);
nor NOR4 (N7034, N7032, N1660, N6901, N3983);
and AND3 (N7035, N7023, N881, N2266);
not NOT1 (N7036, N7035);
nand NAND2 (N7037, N7029, N5980);
nor NOR3 (N7038, N7031, N6916, N677);
xor XOR2 (N7039, N7028, N1000);
nand NAND3 (N7040, N7015, N3757, N1320);
buf BUF1 (N7041, N6985);
and AND3 (N7042, N7040, N3027, N1828);
nand NAND4 (N7043, N7033, N6367, N6034, N4155);
nand NAND2 (N7044, N7043, N2537);
nand NAND2 (N7045, N7020, N699);
nand NAND3 (N7046, N7027, N3870, N4371);
xor XOR2 (N7047, N7041, N591);
or OR2 (N7048, N7045, N3494);
xor XOR2 (N7049, N7047, N2033);
and AND3 (N7050, N7038, N448, N5643);
and AND4 (N7051, N7039, N4167, N6355, N6949);
not NOT1 (N7052, N7049);
and AND3 (N7053, N7034, N2062, N5717);
and AND2 (N7054, N7048, N4719);
and AND3 (N7055, N7042, N4825, N4492);
xor XOR2 (N7056, N7046, N1059);
and AND3 (N7057, N7051, N3239, N198);
nand NAND3 (N7058, N7053, N3451, N2570);
buf BUF1 (N7059, N7050);
nand NAND3 (N7060, N7036, N1192, N4791);
and AND2 (N7061, N7044, N2139);
and AND3 (N7062, N7060, N5175, N6674);
or OR3 (N7063, N7059, N5600, N3401);
nand NAND4 (N7064, N7056, N2050, N6087, N2222);
nand NAND4 (N7065, N7057, N1774, N3455, N419);
xor XOR2 (N7066, N7054, N3376);
xor XOR2 (N7067, N7064, N3139);
or OR2 (N7068, N7065, N3896);
or OR3 (N7069, N7066, N1377, N1176);
or OR3 (N7070, N7055, N1375, N2363);
buf BUF1 (N7071, N7069);
not NOT1 (N7072, N7063);
nor NOR2 (N7073, N7062, N3971);
and AND2 (N7074, N7061, N4273);
not NOT1 (N7075, N7073);
or OR4 (N7076, N7067, N3000, N4015, N3531);
not NOT1 (N7077, N7052);
nand NAND3 (N7078, N7058, N3542, N6945);
or OR4 (N7079, N7074, N983, N6, N737);
buf BUF1 (N7080, N7078);
and AND2 (N7081, N7075, N2106);
xor XOR2 (N7082, N7081, N2056);
or OR4 (N7083, N7037, N1289, N6600, N6826);
nor NOR3 (N7084, N7077, N3160, N2062);
nand NAND4 (N7085, N7079, N6764, N954, N5011);
or OR2 (N7086, N7076, N1619);
not NOT1 (N7087, N7085);
not NOT1 (N7088, N7086);
nor NOR2 (N7089, N7080, N982);
and AND4 (N7090, N7068, N7069, N5916, N2033);
not NOT1 (N7091, N7083);
nor NOR4 (N7092, N7090, N56, N1171, N2579);
nand NAND3 (N7093, N7071, N4428, N2438);
buf BUF1 (N7094, N7072);
buf BUF1 (N7095, N7082);
nand NAND4 (N7096, N7084, N5076, N2789, N6840);
or OR2 (N7097, N7070, N5490);
and AND4 (N7098, N7091, N4171, N4627, N889);
or OR2 (N7099, N7092, N1226);
xor XOR2 (N7100, N7098, N5066);
or OR2 (N7101, N7096, N6834);
xor XOR2 (N7102, N7088, N2062);
not NOT1 (N7103, N7099);
or OR3 (N7104, N7095, N2790, N4096);
and AND2 (N7105, N7089, N4062);
not NOT1 (N7106, N7104);
and AND3 (N7107, N7105, N2718, N5754);
and AND3 (N7108, N7094, N5498, N3255);
or OR3 (N7109, N7102, N6875, N452);
or OR3 (N7110, N7109, N3198, N2748);
xor XOR2 (N7111, N7101, N7106);
nor NOR2 (N7112, N1238, N2239);
buf BUF1 (N7113, N7112);
nor NOR4 (N7114, N7100, N1963, N4974, N5176);
and AND4 (N7115, N7107, N3176, N2017, N1238);
nor NOR2 (N7116, N7093, N3914);
xor XOR2 (N7117, N7108, N6013);
nand NAND2 (N7118, N7087, N6179);
nor NOR3 (N7119, N7103, N724, N1278);
buf BUF1 (N7120, N7113);
or OR3 (N7121, N7120, N4851, N6854);
and AND2 (N7122, N7118, N2481);
buf BUF1 (N7123, N7097);
nand NAND3 (N7124, N7115, N5809, N2139);
nor NOR3 (N7125, N7114, N3462, N5710);
buf BUF1 (N7126, N7119);
buf BUF1 (N7127, N7116);
or OR4 (N7128, N7125, N2208, N762, N2839);
and AND2 (N7129, N7111, N948);
or OR4 (N7130, N7123, N4383, N3945, N1421);
and AND4 (N7131, N7126, N904, N4510, N763);
nand NAND3 (N7132, N7124, N6998, N2985);
nand NAND4 (N7133, N7127, N1491, N6419, N580);
buf BUF1 (N7134, N7110);
not NOT1 (N7135, N7121);
buf BUF1 (N7136, N7130);
nand NAND4 (N7137, N7122, N3042, N3508, N5187);
nand NAND3 (N7138, N7132, N5638, N3537);
and AND2 (N7139, N7135, N3808);
and AND4 (N7140, N7137, N6970, N5111, N578);
xor XOR2 (N7141, N7117, N6744);
not NOT1 (N7142, N7133);
nor NOR3 (N7143, N7140, N4019, N84);
nor NOR4 (N7144, N7131, N328, N5599, N3607);
buf BUF1 (N7145, N7144);
buf BUF1 (N7146, N7138);
or OR2 (N7147, N7141, N2784);
nor NOR4 (N7148, N7134, N2302, N4577, N5074);
and AND3 (N7149, N7143, N2193, N115);
not NOT1 (N7150, N7142);
buf BUF1 (N7151, N7128);
and AND3 (N7152, N7151, N7077, N6778);
or OR2 (N7153, N7139, N5660);
and AND4 (N7154, N7148, N2064, N5689, N6328);
and AND2 (N7155, N7147, N1057);
or OR2 (N7156, N7145, N2038);
and AND3 (N7157, N7156, N5741, N1736);
nor NOR4 (N7158, N7149, N3591, N4391, N3487);
nand NAND2 (N7159, N7136, N3417);
buf BUF1 (N7160, N7155);
or OR4 (N7161, N7158, N5672, N3015, N220);
not NOT1 (N7162, N7152);
buf BUF1 (N7163, N7161);
and AND3 (N7164, N7157, N2710, N109);
and AND2 (N7165, N7160, N373);
or OR4 (N7166, N7150, N3384, N4536, N956);
not NOT1 (N7167, N7159);
buf BUF1 (N7168, N7163);
not NOT1 (N7169, N7129);
buf BUF1 (N7170, N7165);
nand NAND2 (N7171, N7146, N6537);
nand NAND4 (N7172, N7162, N4037, N2609, N1447);
xor XOR2 (N7173, N7167, N4563);
or OR4 (N7174, N7164, N5199, N21, N1948);
buf BUF1 (N7175, N7170);
buf BUF1 (N7176, N7173);
xor XOR2 (N7177, N7174, N3727);
nor NOR2 (N7178, N7153, N2523);
nand NAND4 (N7179, N7168, N1658, N3487, N1761);
nand NAND4 (N7180, N7154, N6745, N4630, N6334);
not NOT1 (N7181, N7172);
and AND2 (N7182, N7175, N3186);
buf BUF1 (N7183, N7169);
or OR3 (N7184, N7181, N4825, N2865);
buf BUF1 (N7185, N7176);
and AND4 (N7186, N7182, N6434, N6915, N6610);
or OR4 (N7187, N7178, N5231, N5058, N1796);
not NOT1 (N7188, N7180);
not NOT1 (N7189, N7186);
or OR2 (N7190, N7187, N2313);
xor XOR2 (N7191, N7188, N4105);
nand NAND2 (N7192, N7185, N2199);
not NOT1 (N7193, N7171);
nand NAND4 (N7194, N7177, N908, N3095, N6647);
not NOT1 (N7195, N7183);
or OR2 (N7196, N7189, N3227);
and AND2 (N7197, N7193, N2702);
buf BUF1 (N7198, N7192);
or OR4 (N7199, N7179, N4272, N6242, N3006);
buf BUF1 (N7200, N7191);
not NOT1 (N7201, N7199);
xor XOR2 (N7202, N7190, N1916);
and AND4 (N7203, N7166, N3380, N127, N1733);
buf BUF1 (N7204, N7184);
or OR2 (N7205, N7204, N4389);
buf BUF1 (N7206, N7201);
xor XOR2 (N7207, N7202, N5276);
nor NOR4 (N7208, N7203, N6595, N3064, N2799);
xor XOR2 (N7209, N7194, N1521);
nor NOR4 (N7210, N7207, N1845, N6420, N3453);
buf BUF1 (N7211, N7206);
and AND4 (N7212, N7209, N5369, N1433, N4799);
nand NAND2 (N7213, N7211, N4566);
nor NOR4 (N7214, N7197, N5623, N817, N3497);
buf BUF1 (N7215, N7195);
nor NOR2 (N7216, N7215, N2611);
nor NOR3 (N7217, N7216, N3244, N2981);
xor XOR2 (N7218, N7200, N6458);
nor NOR2 (N7219, N7217, N2541);
or OR3 (N7220, N7210, N3884, N1791);
not NOT1 (N7221, N7214);
nand NAND2 (N7222, N7208, N2029);
nand NAND4 (N7223, N7219, N4926, N2165, N7200);
nand NAND3 (N7224, N7218, N4392, N777);
and AND2 (N7225, N7222, N2583);
or OR4 (N7226, N7205, N419, N6518, N5110);
xor XOR2 (N7227, N7225, N2788);
not NOT1 (N7228, N7212);
not NOT1 (N7229, N7213);
buf BUF1 (N7230, N7221);
xor XOR2 (N7231, N7230, N1833);
buf BUF1 (N7232, N7198);
and AND4 (N7233, N7232, N6603, N4843, N5852);
not NOT1 (N7234, N7231);
nor NOR3 (N7235, N7234, N6935, N4632);
nor NOR4 (N7236, N7224, N3340, N2858, N536);
and AND4 (N7237, N7226, N362, N1113, N2802);
or OR4 (N7238, N7233, N3676, N41, N7057);
not NOT1 (N7239, N7229);
nor NOR2 (N7240, N7227, N1322);
xor XOR2 (N7241, N7238, N2348);
not NOT1 (N7242, N7241);
nor NOR2 (N7243, N7196, N3712);
buf BUF1 (N7244, N7243);
nor NOR2 (N7245, N7239, N1493);
nor NOR2 (N7246, N7242, N6378);
nor NOR3 (N7247, N7240, N7142, N6870);
buf BUF1 (N7248, N7236);
and AND2 (N7249, N7237, N2148);
buf BUF1 (N7250, N7247);
nand NAND3 (N7251, N7249, N6546, N667);
not NOT1 (N7252, N7223);
buf BUF1 (N7253, N7251);
and AND3 (N7254, N7235, N1264, N4930);
and AND2 (N7255, N7245, N3225);
xor XOR2 (N7256, N7246, N5638);
buf BUF1 (N7257, N7252);
and AND3 (N7258, N7253, N1549, N2082);
nand NAND3 (N7259, N7256, N74, N7258);
or OR2 (N7260, N5199, N6490);
nand NAND2 (N7261, N7255, N4873);
nor NOR3 (N7262, N7220, N2048, N4092);
xor XOR2 (N7263, N7250, N3948);
xor XOR2 (N7264, N7259, N3952);
buf BUF1 (N7265, N7244);
nor NOR3 (N7266, N7248, N38, N5723);
nand NAND3 (N7267, N7265, N906, N3438);
not NOT1 (N7268, N7263);
not NOT1 (N7269, N7264);
nand NAND2 (N7270, N7262, N4204);
nand NAND3 (N7271, N7261, N3457, N6767);
and AND3 (N7272, N7254, N2146, N5428);
nand NAND3 (N7273, N7272, N4818, N4016);
or OR4 (N7274, N7228, N1456, N4235, N710);
buf BUF1 (N7275, N7267);
or OR4 (N7276, N7271, N6085, N5673, N855);
and AND4 (N7277, N7276, N2926, N3069, N3651);
or OR3 (N7278, N7277, N4883, N3146);
xor XOR2 (N7279, N7270, N4007);
nor NOR2 (N7280, N7269, N6199);
buf BUF1 (N7281, N7268);
or OR4 (N7282, N7279, N2827, N2189, N4966);
nand NAND2 (N7283, N7275, N2086);
xor XOR2 (N7284, N7273, N3802);
buf BUF1 (N7285, N7260);
buf BUF1 (N7286, N7285);
nand NAND4 (N7287, N7283, N1900, N4153, N3844);
buf BUF1 (N7288, N7281);
nand NAND3 (N7289, N7278, N4368, N5478);
not NOT1 (N7290, N7266);
xor XOR2 (N7291, N7284, N4424);
nor NOR3 (N7292, N7287, N113, N1057);
and AND2 (N7293, N7292, N5930);
and AND3 (N7294, N7290, N3671, N815);
xor XOR2 (N7295, N7282, N3239);
not NOT1 (N7296, N7280);
buf BUF1 (N7297, N7274);
not NOT1 (N7298, N7295);
nor NOR3 (N7299, N7294, N3007, N5295);
xor XOR2 (N7300, N7257, N3053);
and AND4 (N7301, N7297, N2525, N3929, N6118);
or OR4 (N7302, N7299, N2142, N5055, N3124);
or OR2 (N7303, N7296, N1760);
nand NAND2 (N7304, N7293, N3444);
or OR4 (N7305, N7303, N7101, N4416, N1826);
nor NOR4 (N7306, N7298, N5689, N407, N4202);
buf BUF1 (N7307, N7302);
nor NOR4 (N7308, N7307, N566, N1147, N7217);
buf BUF1 (N7309, N7304);
not NOT1 (N7310, N7308);
and AND3 (N7311, N7300, N6663, N5323);
xor XOR2 (N7312, N7311, N1194);
buf BUF1 (N7313, N7288);
and AND3 (N7314, N7301, N7288, N2955);
and AND4 (N7315, N7309, N2092, N2157, N4203);
buf BUF1 (N7316, N7306);
nor NOR3 (N7317, N7286, N4016, N2015);
nor NOR4 (N7318, N7312, N3530, N3775, N767);
not NOT1 (N7319, N7316);
and AND4 (N7320, N7315, N420, N3770, N421);
and AND3 (N7321, N7310, N7154, N2052);
nor NOR3 (N7322, N7318, N6208, N4577);
or OR3 (N7323, N7321, N2799, N1021);
and AND2 (N7324, N7317, N5106);
not NOT1 (N7325, N7320);
nand NAND3 (N7326, N7322, N6102, N4235);
and AND3 (N7327, N7323, N4067, N5860);
and AND2 (N7328, N7324, N5468);
nand NAND3 (N7329, N7319, N3510, N5077);
buf BUF1 (N7330, N7326);
and AND4 (N7331, N7328, N654, N4705, N6157);
nor NOR4 (N7332, N7289, N4226, N6300, N5823);
and AND2 (N7333, N7325, N3039);
buf BUF1 (N7334, N7313);
and AND3 (N7335, N7333, N4445, N890);
nor NOR2 (N7336, N7291, N5893);
xor XOR2 (N7337, N7330, N5941);
nand NAND2 (N7338, N7337, N3089);
xor XOR2 (N7339, N7332, N2794);
or OR4 (N7340, N7336, N6585, N901, N4018);
nand NAND3 (N7341, N7334, N1473, N554);
nor NOR4 (N7342, N7340, N5464, N5893, N1106);
and AND2 (N7343, N7342, N5481);
and AND3 (N7344, N7331, N5984, N6652);
buf BUF1 (N7345, N7305);
or OR4 (N7346, N7338, N2164, N2995, N4724);
buf BUF1 (N7347, N7343);
nand NAND2 (N7348, N7341, N2126);
not NOT1 (N7349, N7344);
buf BUF1 (N7350, N7329);
not NOT1 (N7351, N7347);
and AND3 (N7352, N7327, N1012, N2646);
nor NOR3 (N7353, N7348, N2209, N3289);
nor NOR2 (N7354, N7314, N6756);
xor XOR2 (N7355, N7352, N3474);
nor NOR4 (N7356, N7351, N7120, N515, N2884);
and AND4 (N7357, N7355, N3805, N6760, N1210);
nor NOR4 (N7358, N7350, N7118, N2246, N4501);
nand NAND2 (N7359, N7349, N7071);
nor NOR2 (N7360, N7353, N1421);
buf BUF1 (N7361, N7345);
nand NAND4 (N7362, N7346, N3984, N6303, N6844);
nand NAND4 (N7363, N7361, N718, N2670, N3445);
and AND3 (N7364, N7354, N6860, N6782);
or OR4 (N7365, N7335, N6687, N5178, N6426);
nor NOR3 (N7366, N7356, N2641, N39);
not NOT1 (N7367, N7339);
or OR3 (N7368, N7364, N6910, N58);
xor XOR2 (N7369, N7365, N108);
and AND3 (N7370, N7362, N609, N5285);
not NOT1 (N7371, N7368);
nand NAND3 (N7372, N7357, N5577, N3252);
not NOT1 (N7373, N7366);
buf BUF1 (N7374, N7370);
or OR4 (N7375, N7369, N6504, N2917, N2053);
buf BUF1 (N7376, N7367);
and AND3 (N7377, N7359, N4316, N2816);
nor NOR3 (N7378, N7375, N3180, N5951);
buf BUF1 (N7379, N7363);
and AND4 (N7380, N7358, N6731, N4140, N4606);
and AND2 (N7381, N7374, N3158);
and AND2 (N7382, N7377, N577);
and AND3 (N7383, N7373, N4176, N2842);
buf BUF1 (N7384, N7380);
buf BUF1 (N7385, N7381);
and AND3 (N7386, N7360, N4735, N4188);
and AND3 (N7387, N7371, N2619, N3109);
buf BUF1 (N7388, N7372);
nand NAND2 (N7389, N7386, N428);
or OR3 (N7390, N7388, N7190, N5672);
not NOT1 (N7391, N7384);
not NOT1 (N7392, N7390);
nor NOR2 (N7393, N7379, N6923);
or OR2 (N7394, N7383, N1465);
buf BUF1 (N7395, N7376);
and AND3 (N7396, N7394, N1046, N7284);
not NOT1 (N7397, N7393);
nor NOR2 (N7398, N7392, N102);
buf BUF1 (N7399, N7389);
or OR2 (N7400, N7396, N1657);
not NOT1 (N7401, N7391);
not NOT1 (N7402, N7387);
or OR3 (N7403, N7399, N5584, N6093);
nor NOR4 (N7404, N7397, N4351, N4137, N4894);
buf BUF1 (N7405, N7395);
nor NOR3 (N7406, N7401, N705, N3264);
or OR3 (N7407, N7382, N6104, N3754);
not NOT1 (N7408, N7403);
xor XOR2 (N7409, N7385, N4929);
not NOT1 (N7410, N7408);
nor NOR2 (N7411, N7398, N4087);
or OR4 (N7412, N7406, N6526, N1313, N3607);
buf BUF1 (N7413, N7404);
buf BUF1 (N7414, N7413);
or OR4 (N7415, N7405, N1535, N4716, N7055);
not NOT1 (N7416, N7410);
nor NOR4 (N7417, N7411, N3142, N3556, N6314);
nor NOR3 (N7418, N7412, N453, N1525);
not NOT1 (N7419, N7415);
and AND4 (N7420, N7416, N5265, N6842, N3634);
or OR4 (N7421, N7420, N4688, N6593, N4232);
not NOT1 (N7422, N7400);
or OR4 (N7423, N7418, N5344, N3720, N3064);
nand NAND4 (N7424, N7378, N6111, N3343, N6519);
nand NAND3 (N7425, N7417, N3915, N6252);
and AND3 (N7426, N7425, N6478, N5475);
and AND3 (N7427, N7426, N126, N315);
nor NOR3 (N7428, N7414, N6263, N5370);
nand NAND2 (N7429, N7427, N5853);
not NOT1 (N7430, N7402);
not NOT1 (N7431, N7409);
nand NAND2 (N7432, N7428, N2628);
not NOT1 (N7433, N7431);
not NOT1 (N7434, N7429);
xor XOR2 (N7435, N7432, N2884);
or OR4 (N7436, N7430, N6175, N7121, N4920);
not NOT1 (N7437, N7407);
not NOT1 (N7438, N7421);
xor XOR2 (N7439, N7424, N3464);
xor XOR2 (N7440, N7438, N1799);
not NOT1 (N7441, N7423);
nor NOR4 (N7442, N7441, N1957, N4486, N860);
and AND2 (N7443, N7437, N6513);
xor XOR2 (N7444, N7435, N5395);
nor NOR3 (N7445, N7443, N2378, N4619);
not NOT1 (N7446, N7433);
xor XOR2 (N7447, N7444, N208);
nor NOR4 (N7448, N7446, N6244, N2478, N1353);
buf BUF1 (N7449, N7436);
buf BUF1 (N7450, N7439);
and AND3 (N7451, N7447, N1841, N3741);
and AND3 (N7452, N7434, N4392, N2055);
xor XOR2 (N7453, N7419, N2355);
not NOT1 (N7454, N7453);
and AND2 (N7455, N7442, N6896);
nor NOR4 (N7456, N7450, N6153, N3606, N2982);
not NOT1 (N7457, N7456);
nand NAND3 (N7458, N7448, N4864, N7386);
buf BUF1 (N7459, N7454);
nor NOR4 (N7460, N7440, N7038, N761, N7332);
not NOT1 (N7461, N7459);
nor NOR3 (N7462, N7452, N4609, N5419);
nor NOR2 (N7463, N7462, N1582);
nor NOR3 (N7464, N7457, N332, N1001);
nor NOR4 (N7465, N7449, N6744, N3564, N2276);
not NOT1 (N7466, N7465);
nand NAND3 (N7467, N7422, N38, N963);
buf BUF1 (N7468, N7460);
or OR3 (N7469, N7464, N4141, N3556);
not NOT1 (N7470, N7461);
nor NOR2 (N7471, N7467, N4952);
and AND2 (N7472, N7471, N3769);
buf BUF1 (N7473, N7472);
or OR3 (N7474, N7451, N3, N4016);
xor XOR2 (N7475, N7445, N648);
buf BUF1 (N7476, N7473);
nand NAND2 (N7477, N7476, N1642);
nand NAND4 (N7478, N7475, N4060, N6759, N3166);
buf BUF1 (N7479, N7470);
nand NAND2 (N7480, N7458, N2513);
and AND4 (N7481, N7477, N2361, N2748, N4969);
xor XOR2 (N7482, N7480, N4395);
nor NOR2 (N7483, N7474, N1198);
xor XOR2 (N7484, N7481, N1393);
or OR4 (N7485, N7463, N1902, N1449, N1636);
xor XOR2 (N7486, N7469, N6601);
or OR2 (N7487, N7455, N799);
buf BUF1 (N7488, N7478);
nor NOR4 (N7489, N7484, N5088, N3624, N4246);
not NOT1 (N7490, N7483);
or OR2 (N7491, N7490, N6203);
nand NAND4 (N7492, N7486, N7267, N7161, N3694);
xor XOR2 (N7493, N7492, N3773);
and AND3 (N7494, N7482, N1507, N1948);
and AND4 (N7495, N7466, N5248, N4436, N3591);
nor NOR3 (N7496, N7494, N2256, N7486);
buf BUF1 (N7497, N7491);
nor NOR2 (N7498, N7495, N4612);
or OR4 (N7499, N7488, N876, N4597, N1309);
and AND3 (N7500, N7489, N6449, N592);
and AND4 (N7501, N7498, N700, N2713, N534);
not NOT1 (N7502, N7499);
xor XOR2 (N7503, N7468, N6125);
or OR3 (N7504, N7502, N3049, N4139);
not NOT1 (N7505, N7504);
not NOT1 (N7506, N7503);
and AND4 (N7507, N7500, N1331, N3031, N303);
nand NAND2 (N7508, N7507, N4799);
xor XOR2 (N7509, N7508, N3781);
nor NOR2 (N7510, N7493, N764);
buf BUF1 (N7511, N7505);
xor XOR2 (N7512, N7510, N503);
not NOT1 (N7513, N7479);
buf BUF1 (N7514, N7511);
nand NAND4 (N7515, N7514, N4948, N6469, N4944);
nor NOR2 (N7516, N7512, N2207);
nor NOR2 (N7517, N7485, N1769);
or OR4 (N7518, N7501, N6812, N1701, N7201);
buf BUF1 (N7519, N7496);
not NOT1 (N7520, N7516);
or OR4 (N7521, N7497, N6194, N4452, N1907);
or OR4 (N7522, N7506, N3761, N725, N1687);
not NOT1 (N7523, N7517);
buf BUF1 (N7524, N7518);
or OR4 (N7525, N7523, N1887, N1527, N400);
not NOT1 (N7526, N7525);
or OR2 (N7527, N7487, N3368);
nor NOR4 (N7528, N7519, N6190, N5360, N2595);
nand NAND4 (N7529, N7520, N7026, N1906, N3564);
nand NAND2 (N7530, N7529, N5211);
xor XOR2 (N7531, N7528, N6352);
nor NOR3 (N7532, N7524, N2450, N6598);
xor XOR2 (N7533, N7521, N4398);
and AND3 (N7534, N7530, N5465, N2980);
not NOT1 (N7535, N7527);
nor NOR3 (N7536, N7535, N6946, N4037);
and AND3 (N7537, N7513, N1795, N2438);
or OR2 (N7538, N7526, N2120);
and AND2 (N7539, N7536, N4020);
or OR3 (N7540, N7537, N4837, N6629);
not NOT1 (N7541, N7531);
and AND3 (N7542, N7509, N598, N1190);
not NOT1 (N7543, N7542);
buf BUF1 (N7544, N7522);
buf BUF1 (N7545, N7541);
nand NAND2 (N7546, N7532, N4521);
nor NOR4 (N7547, N7544, N3372, N822, N1420);
nand NAND2 (N7548, N7539, N5759);
nor NOR3 (N7549, N7534, N6328, N7413);
not NOT1 (N7550, N7547);
xor XOR2 (N7551, N7515, N2074);
not NOT1 (N7552, N7548);
and AND3 (N7553, N7533, N5954, N1242);
nor NOR4 (N7554, N7546, N2729, N2444, N4026);
buf BUF1 (N7555, N7552);
xor XOR2 (N7556, N7551, N490);
or OR4 (N7557, N7550, N6455, N1804, N5265);
and AND4 (N7558, N7556, N5896, N3207, N2866);
buf BUF1 (N7559, N7549);
xor XOR2 (N7560, N7543, N347);
xor XOR2 (N7561, N7553, N4132);
nor NOR2 (N7562, N7560, N2306);
buf BUF1 (N7563, N7559);
xor XOR2 (N7564, N7545, N1153);
nor NOR2 (N7565, N7562, N3540);
or OR2 (N7566, N7561, N716);
xor XOR2 (N7567, N7538, N2546);
nand NAND3 (N7568, N7563, N5361, N1936);
xor XOR2 (N7569, N7564, N7562);
not NOT1 (N7570, N7568);
and AND3 (N7571, N7569, N2179, N4397);
nor NOR4 (N7572, N7570, N3872, N7280, N7318);
buf BUF1 (N7573, N7540);
nand NAND2 (N7574, N7571, N6161);
nor NOR3 (N7575, N7566, N6506, N3939);
xor XOR2 (N7576, N7574, N2095);
nand NAND3 (N7577, N7567, N7334, N6230);
not NOT1 (N7578, N7577);
or OR4 (N7579, N7573, N6177, N3591, N6643);
and AND2 (N7580, N7576, N6401);
xor XOR2 (N7581, N7578, N3229);
xor XOR2 (N7582, N7565, N1877);
nor NOR4 (N7583, N7582, N1531, N2450, N3090);
or OR2 (N7584, N7579, N4384);
and AND3 (N7585, N7557, N580, N4158);
xor XOR2 (N7586, N7581, N5423);
not NOT1 (N7587, N7572);
nand NAND3 (N7588, N7555, N5422, N6292);
and AND4 (N7589, N7580, N3939, N626, N2284);
buf BUF1 (N7590, N7558);
xor XOR2 (N7591, N7584, N1531);
and AND3 (N7592, N7591, N1318, N3587);
or OR4 (N7593, N7586, N693, N5864, N4014);
or OR3 (N7594, N7585, N3748, N1316);
xor XOR2 (N7595, N7554, N4327);
not NOT1 (N7596, N7587);
nor NOR3 (N7597, N7583, N2884, N290);
and AND4 (N7598, N7589, N1231, N7296, N5580);
buf BUF1 (N7599, N7596);
and AND2 (N7600, N7592, N6624);
or OR2 (N7601, N7600, N3251);
nor NOR2 (N7602, N7590, N2218);
buf BUF1 (N7603, N7593);
xor XOR2 (N7604, N7595, N7010);
nor NOR2 (N7605, N7598, N4945);
xor XOR2 (N7606, N7594, N1399);
and AND4 (N7607, N7575, N1699, N1753, N4177);
not NOT1 (N7608, N7605);
xor XOR2 (N7609, N7599, N3565);
and AND3 (N7610, N7606, N1233, N2002);
buf BUF1 (N7611, N7602);
not NOT1 (N7612, N7611);
buf BUF1 (N7613, N7607);
and AND4 (N7614, N7604, N3483, N7271, N4741);
nor NOR3 (N7615, N7612, N2552, N2190);
xor XOR2 (N7616, N7597, N333);
not NOT1 (N7617, N7613);
or OR4 (N7618, N7614, N2778, N3409, N5733);
or OR3 (N7619, N7603, N3736, N4216);
or OR2 (N7620, N7609, N620);
not NOT1 (N7621, N7601);
nor NOR2 (N7622, N7610, N7419);
nor NOR3 (N7623, N7619, N6023, N7195);
xor XOR2 (N7624, N7588, N5788);
buf BUF1 (N7625, N7622);
nand NAND4 (N7626, N7623, N1807, N5198, N7344);
or OR2 (N7627, N7618, N256);
nand NAND3 (N7628, N7608, N3230, N3323);
xor XOR2 (N7629, N7615, N3064);
buf BUF1 (N7630, N7616);
or OR2 (N7631, N7627, N1556);
and AND2 (N7632, N7631, N5600);
nor NOR2 (N7633, N7624, N6662);
nand NAND4 (N7634, N7626, N2867, N6555, N2170);
and AND4 (N7635, N7621, N10, N797, N334);
nand NAND2 (N7636, N7629, N6233);
buf BUF1 (N7637, N7632);
buf BUF1 (N7638, N7630);
or OR4 (N7639, N7617, N3694, N3827, N6255);
buf BUF1 (N7640, N7637);
not NOT1 (N7641, N7636);
or OR3 (N7642, N7639, N5724, N3921);
and AND2 (N7643, N7633, N3395);
nand NAND2 (N7644, N7620, N2842);
and AND4 (N7645, N7635, N6114, N2175, N3815);
or OR3 (N7646, N7634, N5680, N2889);
not NOT1 (N7647, N7628);
nand NAND2 (N7648, N7642, N7012);
or OR4 (N7649, N7643, N6785, N1085, N2861);
or OR3 (N7650, N7625, N3604, N1570);
nand NAND3 (N7651, N7640, N2653, N5286);
not NOT1 (N7652, N7638);
xor XOR2 (N7653, N7641, N595);
or OR4 (N7654, N7652, N2043, N4316, N3330);
nor NOR4 (N7655, N7650, N2026, N5687, N5128);
nor NOR3 (N7656, N7648, N410, N4492);
and AND2 (N7657, N7654, N1178);
buf BUF1 (N7658, N7656);
and AND2 (N7659, N7651, N708);
or OR3 (N7660, N7644, N6924, N1302);
or OR4 (N7661, N7655, N3699, N2823, N1473);
or OR4 (N7662, N7661, N6354, N4369, N2628);
and AND4 (N7663, N7658, N5212, N5389, N7070);
and AND4 (N7664, N7647, N6584, N7514, N2743);
not NOT1 (N7665, N7663);
xor XOR2 (N7666, N7649, N5026);
nand NAND3 (N7667, N7662, N1871, N2145);
nor NOR4 (N7668, N7653, N6194, N4005, N3344);
xor XOR2 (N7669, N7646, N6952);
and AND4 (N7670, N7667, N6113, N7305, N5140);
nand NAND2 (N7671, N7666, N2941);
xor XOR2 (N7672, N7664, N2921);
and AND2 (N7673, N7657, N1606);
nor NOR3 (N7674, N7659, N5679, N6399);
buf BUF1 (N7675, N7670);
nor NOR2 (N7676, N7660, N411);
nand NAND4 (N7677, N7669, N4849, N718, N5727);
nand NAND4 (N7678, N7668, N3349, N6660, N7389);
nand NAND3 (N7679, N7671, N5211, N4298);
or OR4 (N7680, N7677, N3438, N5263, N1596);
not NOT1 (N7681, N7680);
or OR4 (N7682, N7665, N2669, N6432, N2772);
xor XOR2 (N7683, N7682, N2711);
nor NOR3 (N7684, N7676, N4899, N637);
xor XOR2 (N7685, N7675, N192);
not NOT1 (N7686, N7684);
nand NAND4 (N7687, N7683, N2779, N2009, N1174);
not NOT1 (N7688, N7674);
or OR4 (N7689, N7672, N333, N7268, N4850);
nor NOR2 (N7690, N7685, N4667);
nand NAND3 (N7691, N7688, N4333, N4997);
nor NOR3 (N7692, N7686, N5248, N1671);
nor NOR4 (N7693, N7691, N6474, N5580, N4386);
not NOT1 (N7694, N7681);
not NOT1 (N7695, N7692);
xor XOR2 (N7696, N7678, N5663);
not NOT1 (N7697, N7693);
and AND3 (N7698, N7645, N3076, N6042);
or OR2 (N7699, N7690, N983);
not NOT1 (N7700, N7698);
buf BUF1 (N7701, N7696);
and AND3 (N7702, N7689, N517, N1271);
buf BUF1 (N7703, N7673);
and AND4 (N7704, N7699, N526, N4686, N4716);
nand NAND3 (N7705, N7695, N2615, N7458);
not NOT1 (N7706, N7702);
nor NOR3 (N7707, N7706, N5580, N6312);
and AND2 (N7708, N7707, N1037);
nor NOR2 (N7709, N7703, N7490);
and AND4 (N7710, N7697, N597, N7080, N3055);
or OR3 (N7711, N7710, N1716, N5756);
or OR2 (N7712, N7694, N136);
or OR3 (N7713, N7711, N6264, N3229);
not NOT1 (N7714, N7705);
nand NAND4 (N7715, N7679, N1175, N4037, N3209);
or OR2 (N7716, N7704, N7);
xor XOR2 (N7717, N7700, N1567);
and AND2 (N7718, N7701, N5167);
xor XOR2 (N7719, N7714, N1299);
nand NAND2 (N7720, N7712, N4121);
xor XOR2 (N7721, N7717, N4653);
nand NAND4 (N7722, N7721, N4070, N1406, N2637);
xor XOR2 (N7723, N7718, N5949);
not NOT1 (N7724, N7708);
nor NOR3 (N7725, N7722, N7659, N3308);
nand NAND4 (N7726, N7687, N1371, N7549, N6362);
not NOT1 (N7727, N7724);
nor NOR4 (N7728, N7715, N2615, N1770, N2635);
nand NAND2 (N7729, N7719, N6605);
buf BUF1 (N7730, N7720);
and AND3 (N7731, N7713, N2838, N3316);
or OR2 (N7732, N7716, N1518);
nand NAND2 (N7733, N7725, N653);
nand NAND4 (N7734, N7723, N6376, N7404, N5545);
nor NOR2 (N7735, N7730, N106);
and AND3 (N7736, N7726, N3684, N4372);
nor NOR3 (N7737, N7709, N2214, N1534);
or OR4 (N7738, N7734, N994, N952, N2510);
nand NAND3 (N7739, N7729, N6577, N5833);
nor NOR2 (N7740, N7728, N2345);
xor XOR2 (N7741, N7733, N4779);
buf BUF1 (N7742, N7740);
and AND2 (N7743, N7738, N1659);
nor NOR2 (N7744, N7731, N504);
nor NOR2 (N7745, N7727, N5198);
and AND2 (N7746, N7743, N3303);
xor XOR2 (N7747, N7736, N1145);
or OR4 (N7748, N7739, N4378, N1828, N5169);
xor XOR2 (N7749, N7732, N2878);
and AND4 (N7750, N7744, N6536, N3289, N5057);
xor XOR2 (N7751, N7746, N4508);
xor XOR2 (N7752, N7748, N2238);
nor NOR2 (N7753, N7735, N6713);
not NOT1 (N7754, N7749);
nand NAND2 (N7755, N7750, N5849);
or OR2 (N7756, N7742, N386);
buf BUF1 (N7757, N7747);
not NOT1 (N7758, N7756);
xor XOR2 (N7759, N7758, N953);
and AND2 (N7760, N7752, N3892);
and AND2 (N7761, N7759, N630);
nor NOR4 (N7762, N7741, N2971, N6391, N4545);
or OR4 (N7763, N7754, N3125, N742, N4715);
nor NOR3 (N7764, N7763, N7253, N5106);
and AND3 (N7765, N7753, N7017, N2410);
or OR4 (N7766, N7762, N2646, N4934, N4286);
nor NOR3 (N7767, N7760, N1206, N5723);
nand NAND3 (N7768, N7761, N4675, N6038);
nand NAND4 (N7769, N7766, N6276, N2280, N5306);
nand NAND4 (N7770, N7764, N5607, N3563, N4261);
and AND3 (N7771, N7767, N397, N3220);
buf BUF1 (N7772, N7757);
not NOT1 (N7773, N7751);
or OR3 (N7774, N7773, N1379, N6391);
and AND3 (N7775, N7770, N7005, N4620);
xor XOR2 (N7776, N7775, N3267);
nand NAND3 (N7777, N7755, N2788, N1330);
nand NAND2 (N7778, N7772, N2787);
xor XOR2 (N7779, N7745, N6122);
nand NAND3 (N7780, N7778, N3085, N283);
nor NOR3 (N7781, N7777, N2667, N1687);
and AND3 (N7782, N7765, N5897, N5743);
and AND2 (N7783, N7782, N3207);
buf BUF1 (N7784, N7779);
nand NAND2 (N7785, N7780, N6738);
xor XOR2 (N7786, N7768, N5922);
not NOT1 (N7787, N7785);
buf BUF1 (N7788, N7771);
buf BUF1 (N7789, N7787);
and AND2 (N7790, N7776, N2562);
buf BUF1 (N7791, N7781);
xor XOR2 (N7792, N7784, N5745);
nor NOR4 (N7793, N7791, N3743, N4352, N3114);
xor XOR2 (N7794, N7792, N2197);
xor XOR2 (N7795, N7774, N4176);
xor XOR2 (N7796, N7786, N6725);
not NOT1 (N7797, N7769);
buf BUF1 (N7798, N7796);
or OR3 (N7799, N7737, N7202, N5680);
not NOT1 (N7800, N7797);
buf BUF1 (N7801, N7793);
nor NOR4 (N7802, N7790, N791, N7618, N5019);
or OR3 (N7803, N7789, N414, N735);
xor XOR2 (N7804, N7799, N1974);
and AND3 (N7805, N7800, N3651, N1131);
nor NOR4 (N7806, N7801, N1360, N2558, N6335);
nor NOR4 (N7807, N7794, N1083, N2873, N5417);
or OR2 (N7808, N7788, N484);
nor NOR2 (N7809, N7783, N5875);
and AND3 (N7810, N7798, N248, N4468);
and AND2 (N7811, N7804, N5145);
nor NOR2 (N7812, N7803, N4068);
and AND4 (N7813, N7806, N3907, N6394, N4974);
or OR4 (N7814, N7805, N2807, N3231, N7369);
or OR3 (N7815, N7811, N4327, N5596);
xor XOR2 (N7816, N7815, N7039);
xor XOR2 (N7817, N7813, N2103);
nor NOR3 (N7818, N7814, N7053, N3894);
nand NAND4 (N7819, N7817, N5087, N2597, N3055);
xor XOR2 (N7820, N7818, N3894);
nand NAND2 (N7821, N7810, N5095);
not NOT1 (N7822, N7820);
buf BUF1 (N7823, N7808);
nor NOR3 (N7824, N7821, N6103, N4727);
nor NOR2 (N7825, N7795, N4295);
or OR4 (N7826, N7809, N7019, N2300, N1691);
nand NAND3 (N7827, N7812, N5970, N3042);
not NOT1 (N7828, N7827);
or OR2 (N7829, N7802, N1242);
and AND4 (N7830, N7828, N5190, N670, N457);
or OR4 (N7831, N7823, N5416, N4744, N225);
nor NOR3 (N7832, N7831, N674, N5637);
nor NOR2 (N7833, N7819, N6626);
nor NOR2 (N7834, N7816, N7187);
or OR3 (N7835, N7807, N1923, N5949);
nor NOR2 (N7836, N7830, N4008);
nand NAND3 (N7837, N7826, N7758, N4571);
nor NOR4 (N7838, N7822, N2482, N2405, N4497);
or OR3 (N7839, N7824, N3217, N7575);
and AND4 (N7840, N7829, N1968, N5596, N392);
buf BUF1 (N7841, N7838);
nand NAND4 (N7842, N7840, N849, N2438, N7023);
and AND3 (N7843, N7836, N3681, N926);
nor NOR4 (N7844, N7825, N6270, N179, N709);
and AND4 (N7845, N7839, N6390, N6020, N7687);
nand NAND3 (N7846, N7842, N5646, N4614);
buf BUF1 (N7847, N7841);
nand NAND2 (N7848, N7837, N5510);
buf BUF1 (N7849, N7846);
nand NAND4 (N7850, N7834, N901, N5332, N6854);
xor XOR2 (N7851, N7844, N7625);
nand NAND4 (N7852, N7832, N4050, N2905, N6562);
nand NAND3 (N7853, N7835, N23, N2219);
nand NAND3 (N7854, N7850, N3129, N1762);
and AND2 (N7855, N7847, N4172);
buf BUF1 (N7856, N7852);
not NOT1 (N7857, N7843);
nand NAND3 (N7858, N7848, N2123, N3121);
and AND3 (N7859, N7858, N6145, N5676);
not NOT1 (N7860, N7845);
nand NAND4 (N7861, N7859, N1137, N4291, N2737);
not NOT1 (N7862, N7853);
nor NOR3 (N7863, N7862, N2511, N664);
not NOT1 (N7864, N7861);
nand NAND4 (N7865, N7857, N6866, N7505, N1051);
and AND2 (N7866, N7856, N5810);
nor NOR2 (N7867, N7865, N6573);
nand NAND3 (N7868, N7855, N3900, N7448);
and AND2 (N7869, N7860, N1567);
buf BUF1 (N7870, N7854);
xor XOR2 (N7871, N7863, N758);
nor NOR2 (N7872, N7851, N4314);
nor NOR3 (N7873, N7869, N5237, N1353);
nand NAND4 (N7874, N7870, N7152, N5356, N6612);
not NOT1 (N7875, N7868);
buf BUF1 (N7876, N7873);
buf BUF1 (N7877, N7875);
buf BUF1 (N7878, N7874);
and AND4 (N7879, N7833, N5410, N2660, N7361);
not NOT1 (N7880, N7849);
nor NOR3 (N7881, N7864, N3636, N834);
and AND4 (N7882, N7879, N6608, N1741, N1451);
buf BUF1 (N7883, N7866);
xor XOR2 (N7884, N7881, N5896);
buf BUF1 (N7885, N7884);
not NOT1 (N7886, N7871);
nand NAND4 (N7887, N7882, N3854, N6873, N6798);
xor XOR2 (N7888, N7885, N4544);
nand NAND2 (N7889, N7888, N5969);
or OR4 (N7890, N7883, N2566, N4538, N6313);
xor XOR2 (N7891, N7872, N3624);
nand NAND3 (N7892, N7877, N5349, N6742);
nor NOR4 (N7893, N7890, N1715, N1142, N2719);
xor XOR2 (N7894, N7867, N1370);
buf BUF1 (N7895, N7893);
not NOT1 (N7896, N7891);
nand NAND4 (N7897, N7892, N997, N1694, N78);
not NOT1 (N7898, N7887);
not NOT1 (N7899, N7876);
not NOT1 (N7900, N7895);
not NOT1 (N7901, N7898);
or OR2 (N7902, N7886, N2794);
buf BUF1 (N7903, N7889);
xor XOR2 (N7904, N7880, N1629);
not NOT1 (N7905, N7900);
nor NOR3 (N7906, N7899, N6183, N2828);
xor XOR2 (N7907, N7905, N3001);
nand NAND4 (N7908, N7904, N3326, N1043, N5214);
buf BUF1 (N7909, N7897);
or OR2 (N7910, N7909, N3994);
buf BUF1 (N7911, N7878);
and AND2 (N7912, N7911, N5882);
nor NOR2 (N7913, N7906, N7007);
and AND4 (N7914, N7908, N521, N4685, N759);
nor NOR3 (N7915, N7894, N2832, N4043);
or OR2 (N7916, N7914, N5537);
or OR2 (N7917, N7913, N2810);
nand NAND4 (N7918, N7915, N7169, N3656, N7428);
or OR2 (N7919, N7918, N6007);
nand NAND2 (N7920, N7912, N4218);
or OR3 (N7921, N7907, N6851, N4741);
xor XOR2 (N7922, N7921, N6297);
and AND3 (N7923, N7910, N1091, N3972);
not NOT1 (N7924, N7896);
or OR4 (N7925, N7922, N2836, N2701, N2148);
nor NOR4 (N7926, N7916, N984, N6613, N1147);
xor XOR2 (N7927, N7924, N6368);
xor XOR2 (N7928, N7925, N4847);
buf BUF1 (N7929, N7919);
xor XOR2 (N7930, N7901, N2604);
and AND3 (N7931, N7903, N6210, N1484);
or OR3 (N7932, N7917, N5065, N7677);
xor XOR2 (N7933, N7923, N5152);
nand NAND3 (N7934, N7929, N6108, N5274);
nor NOR4 (N7935, N7931, N1056, N1811, N878);
not NOT1 (N7936, N7930);
or OR4 (N7937, N7933, N1849, N5543, N1183);
not NOT1 (N7938, N7926);
not NOT1 (N7939, N7932);
xor XOR2 (N7940, N7920, N7287);
and AND4 (N7941, N7939, N3217, N6328, N6739);
not NOT1 (N7942, N7936);
xor XOR2 (N7943, N7928, N7776);
and AND4 (N7944, N7941, N4938, N3250, N1518);
nor NOR4 (N7945, N7902, N2548, N4362, N642);
buf BUF1 (N7946, N7943);
nand NAND2 (N7947, N7938, N4286);
not NOT1 (N7948, N7946);
and AND2 (N7949, N7944, N911);
and AND2 (N7950, N7942, N578);
nand NAND4 (N7951, N7937, N7139, N841, N229);
nand NAND4 (N7952, N7951, N7322, N3419, N4850);
buf BUF1 (N7953, N7945);
and AND3 (N7954, N7953, N5542, N1099);
xor XOR2 (N7955, N7935, N3389);
xor XOR2 (N7956, N7948, N1919);
and AND3 (N7957, N7950, N1941, N1118);
nand NAND4 (N7958, N7927, N585, N4462, N161);
buf BUF1 (N7959, N7949);
nand NAND3 (N7960, N7934, N6623, N874);
nand NAND3 (N7961, N7947, N6145, N1868);
and AND2 (N7962, N7961, N1896);
not NOT1 (N7963, N7958);
and AND4 (N7964, N7940, N4023, N2746, N2955);
and AND2 (N7965, N7960, N5375);
buf BUF1 (N7966, N7959);
and AND4 (N7967, N7955, N5993, N7904, N6203);
not NOT1 (N7968, N7954);
and AND4 (N7969, N7952, N1573, N3986, N7422);
xor XOR2 (N7970, N7957, N117);
nand NAND4 (N7971, N7966, N1923, N6709, N6193);
nand NAND2 (N7972, N7971, N2234);
nor NOR2 (N7973, N7963, N6891);
nand NAND2 (N7974, N7964, N1485);
nor NOR4 (N7975, N7973, N5814, N7621, N4253);
or OR4 (N7976, N7967, N1086, N5457, N5795);
not NOT1 (N7977, N7968);
nand NAND3 (N7978, N7962, N3354, N5551);
or OR4 (N7979, N7965, N7030, N5009, N5511);
nand NAND4 (N7980, N7979, N1892, N393, N7831);
or OR3 (N7981, N7974, N3107, N2835);
not NOT1 (N7982, N7977);
buf BUF1 (N7983, N7980);
or OR3 (N7984, N7972, N6841, N1154);
or OR2 (N7985, N7975, N7635);
not NOT1 (N7986, N7978);
not NOT1 (N7987, N7984);
or OR2 (N7988, N7982, N2302);
xor XOR2 (N7989, N7969, N2521);
buf BUF1 (N7990, N7983);
nor NOR4 (N7991, N7956, N6439, N2750, N5512);
and AND2 (N7992, N7985, N4563);
and AND2 (N7993, N7991, N1055);
not NOT1 (N7994, N7976);
buf BUF1 (N7995, N7994);
and AND4 (N7996, N7988, N5217, N6164, N7366);
not NOT1 (N7997, N7996);
xor XOR2 (N7998, N7970, N6942);
nor NOR3 (N7999, N7997, N4196, N299);
nor NOR3 (N8000, N7995, N6160, N3157);
or OR4 (N8001, N7998, N6507, N5660, N419);
nand NAND4 (N8002, N7992, N5906, N5664, N4028);
not NOT1 (N8003, N8000);
and AND4 (N8004, N7981, N3665, N4415, N7691);
nor NOR4 (N8005, N7989, N721, N2681, N2786);
xor XOR2 (N8006, N8002, N2284);
and AND2 (N8007, N7993, N6832);
and AND3 (N8008, N8001, N6211, N1624);
nand NAND4 (N8009, N8004, N7921, N4834, N2145);
and AND2 (N8010, N8009, N358);
nand NAND2 (N8011, N8005, N5870);
or OR3 (N8012, N7986, N3547, N4889);
nor NOR4 (N8013, N8012, N6492, N471, N3066);
buf BUF1 (N8014, N8007);
and AND3 (N8015, N8006, N1526, N7521);
and AND3 (N8016, N8011, N3564, N3554);
or OR4 (N8017, N7990, N3180, N2213, N4881);
nor NOR4 (N8018, N8003, N4868, N6218, N7019);
and AND2 (N8019, N8015, N1924);
endmodule