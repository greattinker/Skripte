// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15;

output N25606,N25613,N25611,N25610,N25603,N25608,N25595,N25614,N25612,N25615;

nor NOR3 (N16, N1, N1, N14);
xor XOR2 (N17, N15, N15);
or OR3 (N18, N16, N13, N3);
not NOT1 (N19, N18);
not NOT1 (N20, N6);
not NOT1 (N21, N6);
and AND4 (N22, N9, N7, N6, N7);
and AND2 (N23, N7, N15);
nand NAND4 (N24, N15, N23, N8, N23);
xor XOR2 (N25, N12, N8);
and AND2 (N26, N23, N9);
nor NOR3 (N27, N15, N15, N14);
nand NAND3 (N28, N7, N26, N20);
not NOT1 (N29, N6);
or OR2 (N30, N12, N23);
buf BUF1 (N31, N30);
or OR3 (N32, N29, N2, N3);
or OR3 (N33, N19, N10, N12);
or OR3 (N34, N32, N18, N2);
xor XOR2 (N35, N24, N32);
or OR3 (N36, N27, N18, N32);
buf BUF1 (N37, N36);
and AND3 (N38, N28, N28, N4);
or OR4 (N39, N25, N32, N26, N32);
nand NAND3 (N40, N21, N27, N31);
buf BUF1 (N41, N22);
nand NAND4 (N42, N19, N38, N40, N10);
nor NOR2 (N43, N9, N16);
and AND3 (N44, N30, N33, N11);
xor XOR2 (N45, N8, N4);
not NOT1 (N46, N17);
nor NOR2 (N47, N39, N5);
or OR2 (N48, N47, N23);
or OR2 (N49, N41, N41);
nand NAND3 (N50, N46, N23, N14);
nor NOR4 (N51, N50, N32, N14, N22);
not NOT1 (N52, N51);
not NOT1 (N53, N35);
and AND4 (N54, N52, N47, N24, N24);
and AND2 (N55, N48, N31);
nor NOR4 (N56, N53, N24, N55, N49);
not NOT1 (N57, N12);
not NOT1 (N58, N34);
nor NOR3 (N59, N32, N35, N48);
nor NOR3 (N60, N56, N33, N17);
nand NAND4 (N61, N43, N43, N9, N47);
buf BUF1 (N62, N57);
buf BUF1 (N63, N58);
and AND4 (N64, N60, N37, N46, N48);
nor NOR4 (N65, N17, N44, N32, N50);
nor NOR3 (N66, N28, N5, N53);
not NOT1 (N67, N65);
or OR2 (N68, N54, N47);
buf BUF1 (N69, N62);
not NOT1 (N70, N69);
xor XOR2 (N71, N61, N22);
or OR4 (N72, N66, N52, N5, N5);
xor XOR2 (N73, N63, N63);
or OR3 (N74, N72, N53, N16);
and AND3 (N75, N42, N71, N8);
not NOT1 (N76, N25);
or OR3 (N77, N70, N3, N73);
nand NAND2 (N78, N52, N9);
or OR4 (N79, N74, N35, N67, N30);
not NOT1 (N80, N20);
not NOT1 (N81, N75);
xor XOR2 (N82, N45, N59);
not NOT1 (N83, N62);
or OR2 (N84, N77, N58);
buf BUF1 (N85, N82);
not NOT1 (N86, N80);
or OR4 (N87, N68, N10, N12, N29);
buf BUF1 (N88, N79);
buf BUF1 (N89, N87);
nand NAND4 (N90, N76, N9, N24, N71);
nor NOR2 (N91, N83, N62);
nand NAND2 (N92, N89, N48);
not NOT1 (N93, N78);
and AND4 (N94, N93, N66, N43, N14);
buf BUF1 (N95, N86);
not NOT1 (N96, N95);
buf BUF1 (N97, N92);
nor NOR3 (N98, N81, N86, N16);
not NOT1 (N99, N91);
xor XOR2 (N100, N85, N7);
not NOT1 (N101, N98);
and AND4 (N102, N101, N46, N9, N33);
nand NAND2 (N103, N97, N66);
nand NAND3 (N104, N99, N61, N47);
and AND3 (N105, N64, N34, N48);
nand NAND4 (N106, N104, N88, N19, N76);
nor NOR4 (N107, N1, N23, N91, N11);
buf BUF1 (N108, N100);
nor NOR4 (N109, N105, N49, N91, N26);
nor NOR4 (N110, N96, N101, N92, N55);
nand NAND3 (N111, N102, N92, N71);
nor NOR3 (N112, N84, N67, N111);
xor XOR2 (N113, N73, N97);
not NOT1 (N114, N110);
not NOT1 (N115, N114);
nand NAND3 (N116, N107, N80, N51);
and AND4 (N117, N109, N91, N77, N89);
or OR4 (N118, N90, N34, N103, N44);
not NOT1 (N119, N66);
not NOT1 (N120, N115);
and AND2 (N121, N112, N58);
not NOT1 (N122, N118);
xor XOR2 (N123, N94, N102);
xor XOR2 (N124, N113, N15);
nor NOR3 (N125, N121, N98, N57);
and AND4 (N126, N120, N79, N99, N120);
xor XOR2 (N127, N116, N116);
buf BUF1 (N128, N127);
xor XOR2 (N129, N128, N16);
buf BUF1 (N130, N129);
nand NAND3 (N131, N119, N91, N103);
and AND3 (N132, N131, N106, N77);
or OR3 (N133, N113, N117, N10);
not NOT1 (N134, N43);
and AND3 (N135, N123, N19, N49);
buf BUF1 (N136, N130);
and AND4 (N137, N125, N117, N84, N40);
nor NOR3 (N138, N136, N88, N30);
nor NOR2 (N139, N133, N2);
xor XOR2 (N140, N139, N10);
buf BUF1 (N141, N132);
buf BUF1 (N142, N124);
xor XOR2 (N143, N140, N86);
nor NOR4 (N144, N135, N54, N47, N42);
and AND2 (N145, N144, N104);
xor XOR2 (N146, N138, N9);
xor XOR2 (N147, N126, N93);
xor XOR2 (N148, N142, N125);
and AND3 (N149, N147, N137, N102);
nand NAND2 (N150, N117, N16);
not NOT1 (N151, N108);
or OR3 (N152, N143, N124, N81);
or OR2 (N153, N134, N110);
nor NOR3 (N154, N145, N99, N150);
nor NOR4 (N155, N43, N4, N78, N122);
not NOT1 (N156, N20);
xor XOR2 (N157, N149, N56);
and AND4 (N158, N156, N135, N96, N71);
and AND2 (N159, N141, N85);
nor NOR2 (N160, N146, N72);
nand NAND3 (N161, N153, N127, N28);
nor NOR4 (N162, N159, N91, N50, N114);
or OR3 (N163, N155, N82, N75);
buf BUF1 (N164, N161);
or OR3 (N165, N154, N63, N5);
nor NOR3 (N166, N158, N98, N165);
or OR2 (N167, N159, N125);
nor NOR3 (N168, N148, N72, N82);
xor XOR2 (N169, N163, N160);
nor NOR2 (N170, N148, N164);
or OR3 (N171, N13, N149, N57);
or OR2 (N172, N169, N113);
nor NOR2 (N173, N167, N19);
buf BUF1 (N174, N171);
or OR3 (N175, N172, N165, N66);
buf BUF1 (N176, N170);
xor XOR2 (N177, N152, N33);
xor XOR2 (N178, N176, N102);
not NOT1 (N179, N174);
xor XOR2 (N180, N157, N148);
and AND4 (N181, N151, N115, N104, N171);
and AND2 (N182, N168, N46);
or OR4 (N183, N173, N102, N101, N133);
or OR2 (N184, N162, N108);
and AND3 (N185, N181, N159, N178);
not NOT1 (N186, N153);
and AND2 (N187, N185, N31);
not NOT1 (N188, N166);
nand NAND3 (N189, N179, N138, N163);
xor XOR2 (N190, N183, N156);
xor XOR2 (N191, N182, N92);
nand NAND3 (N192, N187, N139, N50);
xor XOR2 (N193, N190, N115);
or OR2 (N194, N177, N94);
not NOT1 (N195, N188);
and AND4 (N196, N192, N147, N122, N6);
xor XOR2 (N197, N180, N192);
xor XOR2 (N198, N197, N134);
xor XOR2 (N199, N193, N95);
xor XOR2 (N200, N195, N98);
buf BUF1 (N201, N199);
xor XOR2 (N202, N184, N126);
not NOT1 (N203, N200);
or OR3 (N204, N175, N150, N81);
and AND4 (N205, N189, N191, N42, N150);
xor XOR2 (N206, N69, N169);
or OR4 (N207, N206, N81, N27, N184);
xor XOR2 (N208, N205, N34);
not NOT1 (N209, N207);
nand NAND3 (N210, N204, N114, N131);
or OR4 (N211, N186, N183, N92, N7);
xor XOR2 (N212, N202, N69);
buf BUF1 (N213, N203);
nand NAND3 (N214, N209, N194, N162);
or OR2 (N215, N67, N53);
xor XOR2 (N216, N198, N214);
nor NOR3 (N217, N103, N113, N67);
and AND4 (N218, N217, N181, N110, N56);
nand NAND3 (N219, N196, N106, N214);
or OR3 (N220, N201, N134, N16);
or OR4 (N221, N213, N163, N127, N145);
not NOT1 (N222, N211);
xor XOR2 (N223, N212, N63);
not NOT1 (N224, N219);
buf BUF1 (N225, N220);
not NOT1 (N226, N225);
buf BUF1 (N227, N221);
not NOT1 (N228, N223);
nand NAND2 (N229, N216, N80);
buf BUF1 (N230, N227);
nand NAND3 (N231, N230, N42, N28);
nor NOR4 (N232, N208, N164, N147, N139);
xor XOR2 (N233, N231, N159);
not NOT1 (N234, N226);
or OR2 (N235, N218, N40);
not NOT1 (N236, N234);
buf BUF1 (N237, N210);
buf BUF1 (N238, N228);
buf BUF1 (N239, N238);
nor NOR2 (N240, N224, N126);
xor XOR2 (N241, N215, N190);
buf BUF1 (N242, N222);
nand NAND4 (N243, N233, N190, N126, N186);
buf BUF1 (N244, N237);
nand NAND3 (N245, N244, N83, N120);
or OR4 (N246, N245, N140, N94, N14);
or OR3 (N247, N242, N151, N60);
nor NOR4 (N248, N239, N12, N113, N190);
and AND3 (N249, N246, N75, N100);
not NOT1 (N250, N236);
nand NAND3 (N251, N243, N67, N124);
nand NAND3 (N252, N251, N115, N39);
nor NOR2 (N253, N229, N124);
buf BUF1 (N254, N253);
nand NAND4 (N255, N232, N188, N89, N181);
nor NOR4 (N256, N240, N46, N51, N198);
buf BUF1 (N257, N249);
and AND2 (N258, N254, N243);
not NOT1 (N259, N235);
nand NAND3 (N260, N250, N256, N157);
xor XOR2 (N261, N8, N107);
buf BUF1 (N262, N255);
buf BUF1 (N263, N252);
or OR3 (N264, N262, N34, N133);
nand NAND4 (N265, N258, N176, N29, N254);
nor NOR3 (N266, N263, N158, N200);
and AND4 (N267, N261, N111, N169, N125);
not NOT1 (N268, N260);
not NOT1 (N269, N268);
nor NOR4 (N270, N267, N66, N3, N215);
not NOT1 (N271, N265);
and AND4 (N272, N264, N246, N118, N185);
not NOT1 (N273, N272);
not NOT1 (N274, N266);
xor XOR2 (N275, N271, N51);
and AND2 (N276, N247, N112);
or OR4 (N277, N276, N227, N129, N250);
nor NOR3 (N278, N277, N170, N198);
or OR2 (N279, N241, N18);
and AND2 (N280, N270, N279);
or OR3 (N281, N198, N23, N75);
and AND3 (N282, N278, N169, N29);
buf BUF1 (N283, N282);
not NOT1 (N284, N274);
and AND4 (N285, N280, N31, N94, N6);
not NOT1 (N286, N284);
xor XOR2 (N287, N259, N49);
xor XOR2 (N288, N248, N168);
and AND2 (N289, N283, N72);
and AND4 (N290, N285, N190, N173, N65);
or OR4 (N291, N286, N280, N57, N164);
buf BUF1 (N292, N273);
nor NOR2 (N293, N281, N227);
buf BUF1 (N294, N293);
buf BUF1 (N295, N269);
not NOT1 (N296, N287);
nor NOR4 (N297, N288, N215, N101, N37);
nor NOR4 (N298, N290, N175, N2, N159);
not NOT1 (N299, N294);
or OR2 (N300, N291, N27);
nand NAND4 (N301, N300, N2, N120, N206);
or OR3 (N302, N296, N69, N117);
not NOT1 (N303, N302);
nor NOR4 (N304, N303, N143, N115, N178);
buf BUF1 (N305, N301);
xor XOR2 (N306, N297, N265);
xor XOR2 (N307, N295, N3);
not NOT1 (N308, N299);
buf BUF1 (N309, N307);
or OR2 (N310, N306, N36);
nor NOR4 (N311, N309, N176, N39, N21);
nor NOR3 (N312, N304, N26, N274);
nor NOR3 (N313, N311, N60, N278);
or OR4 (N314, N305, N74, N14, N216);
and AND2 (N315, N313, N240);
and AND3 (N316, N257, N291, N24);
nand NAND2 (N317, N289, N311);
not NOT1 (N318, N292);
buf BUF1 (N319, N318);
buf BUF1 (N320, N312);
nand NAND4 (N321, N315, N68, N213, N2);
nor NOR4 (N322, N275, N291, N110, N132);
or OR2 (N323, N317, N319);
xor XOR2 (N324, N204, N270);
nor NOR4 (N325, N322, N151, N321, N201);
nand NAND4 (N326, N268, N156, N2, N101);
and AND4 (N327, N320, N61, N5, N183);
and AND3 (N328, N325, N249, N144);
or OR2 (N329, N327, N137);
and AND4 (N330, N328, N33, N124, N277);
nand NAND3 (N331, N324, N247, N168);
xor XOR2 (N332, N331, N153);
or OR2 (N333, N323, N69);
buf BUF1 (N334, N308);
xor XOR2 (N335, N310, N43);
or OR3 (N336, N298, N319, N165);
xor XOR2 (N337, N329, N173);
xor XOR2 (N338, N330, N18);
buf BUF1 (N339, N316);
nand NAND3 (N340, N326, N311, N252);
nand NAND4 (N341, N334, N232, N160, N340);
nand NAND3 (N342, N172, N63, N237);
nand NAND4 (N343, N332, N134, N231, N318);
buf BUF1 (N344, N341);
xor XOR2 (N345, N336, N245);
buf BUF1 (N346, N342);
nand NAND4 (N347, N337, N176, N145, N275);
xor XOR2 (N348, N339, N209);
not NOT1 (N349, N348);
xor XOR2 (N350, N333, N328);
nand NAND3 (N351, N344, N193, N293);
buf BUF1 (N352, N343);
not NOT1 (N353, N350);
nor NOR3 (N354, N338, N301, N316);
xor XOR2 (N355, N353, N12);
not NOT1 (N356, N352);
or OR3 (N357, N354, N225, N144);
and AND3 (N358, N355, N289, N194);
xor XOR2 (N359, N346, N281);
nand NAND3 (N360, N347, N265, N176);
buf BUF1 (N361, N358);
xor XOR2 (N362, N361, N3);
or OR2 (N363, N349, N36);
and AND4 (N364, N356, N161, N224, N32);
xor XOR2 (N365, N314, N127);
and AND3 (N366, N335, N40, N244);
nor NOR3 (N367, N366, N295, N245);
or OR3 (N368, N345, N236, N2);
nor NOR3 (N369, N351, N10, N199);
xor XOR2 (N370, N367, N278);
nor NOR3 (N371, N368, N321, N136);
buf BUF1 (N372, N359);
or OR3 (N373, N364, N21, N68);
xor XOR2 (N374, N372, N42);
and AND3 (N375, N369, N264, N76);
or OR2 (N376, N362, N131);
nand NAND4 (N377, N360, N243, N157, N304);
not NOT1 (N378, N371);
nor NOR4 (N379, N375, N240, N200, N173);
nor NOR3 (N380, N378, N128, N176);
and AND3 (N381, N380, N10, N5);
not NOT1 (N382, N363);
and AND2 (N383, N373, N237);
and AND2 (N384, N379, N279);
buf BUF1 (N385, N384);
not NOT1 (N386, N377);
buf BUF1 (N387, N381);
nor NOR4 (N388, N376, N180, N127, N251);
buf BUF1 (N389, N370);
nand NAND3 (N390, N385, N291, N189);
not NOT1 (N391, N374);
buf BUF1 (N392, N387);
not NOT1 (N393, N391);
or OR3 (N394, N390, N24, N221);
not NOT1 (N395, N393);
or OR4 (N396, N386, N368, N151, N120);
nor NOR3 (N397, N392, N270, N129);
buf BUF1 (N398, N382);
nand NAND3 (N399, N365, N374, N335);
and AND4 (N400, N396, N174, N306, N372);
nand NAND4 (N401, N389, N236, N246, N211);
xor XOR2 (N402, N395, N320);
not NOT1 (N403, N400);
buf BUF1 (N404, N397);
not NOT1 (N405, N404);
nor NOR4 (N406, N357, N40, N216, N297);
nand NAND4 (N407, N399, N134, N280, N208);
not NOT1 (N408, N403);
buf BUF1 (N409, N383);
nor NOR3 (N410, N407, N202, N192);
buf BUF1 (N411, N388);
xor XOR2 (N412, N401, N39);
and AND3 (N413, N406, N127, N321);
and AND2 (N414, N394, N171);
nand NAND4 (N415, N414, N204, N54, N399);
xor XOR2 (N416, N409, N185);
xor XOR2 (N417, N402, N18);
and AND3 (N418, N408, N308, N75);
nand NAND3 (N419, N398, N151, N267);
xor XOR2 (N420, N417, N323);
or OR4 (N421, N416, N231, N107, N157);
or OR2 (N422, N415, N328);
or OR4 (N423, N419, N400, N144, N178);
not NOT1 (N424, N413);
buf BUF1 (N425, N424);
nand NAND2 (N426, N410, N355);
xor XOR2 (N427, N425, N270);
nand NAND4 (N428, N420, N376, N423, N214);
nor NOR2 (N429, N162, N338);
or OR3 (N430, N428, N43, N369);
and AND3 (N431, N426, N104, N268);
or OR3 (N432, N418, N383, N79);
and AND2 (N433, N421, N296);
and AND2 (N434, N429, N211);
nor NOR2 (N435, N430, N88);
buf BUF1 (N436, N433);
not NOT1 (N437, N432);
not NOT1 (N438, N437);
or OR3 (N439, N411, N181, N401);
nor NOR2 (N440, N436, N127);
nor NOR4 (N441, N412, N331, N331, N147);
buf BUF1 (N442, N441);
nor NOR4 (N443, N427, N407, N397, N328);
or OR4 (N444, N431, N199, N316, N109);
not NOT1 (N445, N405);
buf BUF1 (N446, N443);
buf BUF1 (N447, N435);
or OR3 (N448, N442, N177, N146);
not NOT1 (N449, N446);
or OR4 (N450, N445, N55, N441, N192);
buf BUF1 (N451, N449);
or OR3 (N452, N434, N142, N307);
or OR4 (N453, N444, N98, N94, N250);
buf BUF1 (N454, N447);
nand NAND3 (N455, N448, N415, N78);
or OR4 (N456, N454, N364, N47, N384);
xor XOR2 (N457, N439, N389);
not NOT1 (N458, N457);
xor XOR2 (N459, N455, N428);
nand NAND3 (N460, N452, N285, N207);
and AND2 (N461, N458, N88);
nor NOR3 (N462, N422, N272, N400);
nor NOR3 (N463, N461, N234, N442);
buf BUF1 (N464, N453);
xor XOR2 (N465, N459, N367);
or OR2 (N466, N463, N441);
buf BUF1 (N467, N465);
and AND4 (N468, N450, N342, N277, N400);
and AND3 (N469, N451, N92, N27);
nor NOR2 (N470, N466, N263);
or OR3 (N471, N467, N7, N463);
buf BUF1 (N472, N471);
xor XOR2 (N473, N468, N50);
nor NOR2 (N474, N438, N10);
nand NAND2 (N475, N470, N316);
or OR3 (N476, N472, N131, N379);
or OR3 (N477, N469, N190, N356);
xor XOR2 (N478, N477, N277);
or OR3 (N479, N440, N73, N312);
nand NAND2 (N480, N460, N289);
xor XOR2 (N481, N456, N59);
not NOT1 (N482, N474);
nor NOR3 (N483, N482, N415, N464);
not NOT1 (N484, N243);
nand NAND3 (N485, N480, N179, N295);
xor XOR2 (N486, N483, N195);
xor XOR2 (N487, N484, N482);
and AND4 (N488, N487, N194, N255, N205);
buf BUF1 (N489, N486);
xor XOR2 (N490, N485, N138);
buf BUF1 (N491, N475);
buf BUF1 (N492, N488);
or OR3 (N493, N481, N110, N320);
not NOT1 (N494, N491);
or OR3 (N495, N492, N146, N490);
not NOT1 (N496, N115);
buf BUF1 (N497, N495);
buf BUF1 (N498, N462);
nor NOR4 (N499, N479, N436, N325, N334);
and AND4 (N500, N497, N207, N252, N216);
buf BUF1 (N501, N476);
nand NAND3 (N502, N501, N305, N368);
nor NOR3 (N503, N494, N20, N73);
nor NOR3 (N504, N496, N345, N285);
nor NOR2 (N505, N503, N38);
or OR2 (N506, N500, N465);
or OR4 (N507, N489, N162, N412, N25);
xor XOR2 (N508, N478, N190);
nor NOR3 (N509, N504, N444, N41);
not NOT1 (N510, N502);
xor XOR2 (N511, N473, N12);
or OR3 (N512, N493, N291, N113);
nand NAND4 (N513, N510, N418, N41, N72);
or OR2 (N514, N509, N472);
or OR3 (N515, N508, N74, N158);
buf BUF1 (N516, N498);
xor XOR2 (N517, N513, N466);
buf BUF1 (N518, N516);
not NOT1 (N519, N514);
nor NOR3 (N520, N515, N126, N94);
not NOT1 (N521, N505);
nand NAND3 (N522, N512, N297, N450);
not NOT1 (N523, N506);
nor NOR2 (N524, N521, N228);
nor NOR3 (N525, N522, N375, N266);
or OR2 (N526, N499, N191);
nor NOR4 (N527, N517, N222, N492, N261);
or OR2 (N528, N519, N414);
not NOT1 (N529, N518);
nor NOR2 (N530, N528, N463);
not NOT1 (N531, N507);
xor XOR2 (N532, N524, N388);
nand NAND2 (N533, N523, N329);
not NOT1 (N534, N520);
and AND3 (N535, N534, N214, N457);
or OR4 (N536, N527, N209, N433, N313);
nand NAND3 (N537, N530, N362, N344);
nand NAND4 (N538, N536, N435, N481, N510);
nand NAND2 (N539, N532, N377);
xor XOR2 (N540, N529, N477);
nand NAND4 (N541, N539, N151, N362, N151);
not NOT1 (N542, N535);
nor NOR3 (N543, N511, N457, N462);
not NOT1 (N544, N533);
buf BUF1 (N545, N526);
nand NAND4 (N546, N541, N147, N242, N53);
nand NAND4 (N547, N537, N476, N345, N250);
and AND2 (N548, N531, N86);
not NOT1 (N549, N540);
not NOT1 (N550, N544);
or OR3 (N551, N525, N96, N286);
not NOT1 (N552, N542);
buf BUF1 (N553, N538);
or OR2 (N554, N545, N178);
or OR2 (N555, N549, N63);
or OR3 (N556, N543, N506, N415);
nand NAND3 (N557, N553, N61, N23);
buf BUF1 (N558, N550);
nor NOR2 (N559, N556, N504);
xor XOR2 (N560, N551, N246);
nand NAND3 (N561, N547, N180, N536);
xor XOR2 (N562, N558, N534);
or OR4 (N563, N559, N171, N33, N305);
not NOT1 (N564, N548);
buf BUF1 (N565, N552);
nand NAND3 (N566, N564, N13, N108);
not NOT1 (N567, N546);
or OR3 (N568, N557, N41, N176);
nand NAND2 (N569, N562, N447);
xor XOR2 (N570, N567, N36);
nor NOR4 (N571, N560, N49, N41, N252);
nor NOR4 (N572, N563, N507, N153, N103);
or OR4 (N573, N571, N158, N179, N4);
nor NOR3 (N574, N555, N568, N21);
nor NOR3 (N575, N318, N426, N466);
not NOT1 (N576, N566);
nand NAND4 (N577, N573, N180, N79, N394);
xor XOR2 (N578, N574, N549);
xor XOR2 (N579, N565, N435);
or OR3 (N580, N561, N512, N206);
nand NAND4 (N581, N576, N255, N301, N438);
nor NOR2 (N582, N554, N521);
buf BUF1 (N583, N575);
nand NAND4 (N584, N577, N435, N407, N238);
or OR2 (N585, N580, N19);
nand NAND4 (N586, N584, N557, N379, N403);
or OR2 (N587, N585, N336);
nand NAND3 (N588, N570, N110, N410);
or OR3 (N589, N587, N205, N506);
buf BUF1 (N590, N569);
and AND3 (N591, N583, N189, N438);
and AND3 (N592, N578, N173, N254);
xor XOR2 (N593, N589, N99);
xor XOR2 (N594, N579, N371);
nor NOR2 (N595, N590, N46);
and AND4 (N596, N586, N289, N43, N11);
not NOT1 (N597, N588);
xor XOR2 (N598, N596, N88);
and AND3 (N599, N592, N250, N302);
not NOT1 (N600, N591);
buf BUF1 (N601, N581);
and AND2 (N602, N572, N517);
and AND2 (N603, N582, N490);
not NOT1 (N604, N594);
and AND3 (N605, N595, N553, N110);
or OR3 (N606, N604, N121, N9);
buf BUF1 (N607, N597);
or OR2 (N608, N601, N274);
buf BUF1 (N609, N600);
nand NAND4 (N610, N607, N258, N594, N375);
and AND2 (N611, N606, N143);
buf BUF1 (N612, N603);
and AND3 (N613, N608, N87, N294);
buf BUF1 (N614, N602);
nand NAND4 (N615, N609, N327, N590, N563);
buf BUF1 (N616, N610);
not NOT1 (N617, N614);
or OR4 (N618, N593, N213, N126, N431);
xor XOR2 (N619, N613, N389);
not NOT1 (N620, N599);
nand NAND4 (N621, N616, N114, N450, N159);
and AND3 (N622, N615, N293, N566);
nor NOR2 (N623, N611, N595);
nand NAND2 (N624, N617, N144);
buf BUF1 (N625, N618);
buf BUF1 (N626, N598);
not NOT1 (N627, N621);
and AND2 (N628, N612, N38);
buf BUF1 (N629, N605);
not NOT1 (N630, N628);
and AND4 (N631, N630, N534, N235, N208);
or OR4 (N632, N622, N138, N171, N104);
buf BUF1 (N633, N625);
xor XOR2 (N634, N632, N238);
and AND4 (N635, N634, N459, N561, N172);
or OR4 (N636, N624, N520, N454, N549);
xor XOR2 (N637, N627, N73);
not NOT1 (N638, N635);
or OR3 (N639, N619, N314, N490);
nor NOR3 (N640, N620, N356, N532);
or OR4 (N641, N640, N347, N634, N29);
or OR2 (N642, N631, N352);
buf BUF1 (N643, N636);
or OR3 (N644, N623, N66, N149);
nand NAND4 (N645, N626, N69, N423, N478);
buf BUF1 (N646, N629);
or OR3 (N647, N644, N609, N137);
buf BUF1 (N648, N643);
and AND2 (N649, N641, N265);
nand NAND2 (N650, N647, N277);
nand NAND4 (N651, N648, N171, N336, N73);
and AND4 (N652, N649, N56, N522, N298);
or OR3 (N653, N650, N98, N311);
nand NAND2 (N654, N638, N244);
xor XOR2 (N655, N653, N98);
buf BUF1 (N656, N639);
or OR2 (N657, N656, N404);
nor NOR2 (N658, N646, N256);
or OR3 (N659, N645, N481, N431);
xor XOR2 (N660, N652, N510);
buf BUF1 (N661, N659);
not NOT1 (N662, N657);
or OR4 (N663, N633, N560, N40, N212);
nor NOR3 (N664, N637, N606, N464);
and AND2 (N665, N660, N603);
nor NOR3 (N666, N661, N335, N125);
or OR2 (N667, N665, N613);
nand NAND3 (N668, N642, N514, N613);
xor XOR2 (N669, N668, N72);
not NOT1 (N670, N664);
not NOT1 (N671, N670);
nor NOR4 (N672, N651, N278, N455, N651);
not NOT1 (N673, N672);
and AND2 (N674, N663, N334);
not NOT1 (N675, N658);
buf BUF1 (N676, N674);
not NOT1 (N677, N671);
nor NOR4 (N678, N667, N620, N428, N175);
buf BUF1 (N679, N676);
buf BUF1 (N680, N673);
xor XOR2 (N681, N678, N422);
nand NAND2 (N682, N679, N524);
nor NOR2 (N683, N654, N119);
nand NAND3 (N684, N666, N405, N429);
xor XOR2 (N685, N662, N64);
nor NOR4 (N686, N685, N511, N241, N468);
buf BUF1 (N687, N655);
not NOT1 (N688, N683);
and AND4 (N689, N682, N437, N257, N559);
nand NAND2 (N690, N680, N23);
or OR3 (N691, N688, N196, N411);
or OR3 (N692, N684, N510, N179);
nand NAND4 (N693, N677, N668, N414, N257);
and AND4 (N694, N681, N494, N464, N253);
buf BUF1 (N695, N675);
or OR4 (N696, N669, N597, N118, N328);
nand NAND4 (N697, N692, N206, N592, N142);
nand NAND3 (N698, N695, N74, N54);
or OR4 (N699, N693, N372, N220, N576);
buf BUF1 (N700, N696);
buf BUF1 (N701, N689);
xor XOR2 (N702, N697, N509);
nand NAND2 (N703, N699, N255);
or OR2 (N704, N690, N400);
nand NAND4 (N705, N701, N22, N610, N351);
nand NAND2 (N706, N691, N299);
buf BUF1 (N707, N694);
xor XOR2 (N708, N703, N228);
xor XOR2 (N709, N706, N575);
xor XOR2 (N710, N708, N676);
or OR2 (N711, N704, N441);
nor NOR3 (N712, N705, N559, N305);
or OR2 (N713, N700, N534);
not NOT1 (N714, N709);
or OR4 (N715, N712, N108, N335, N704);
or OR4 (N716, N707, N689, N27, N417);
nand NAND3 (N717, N714, N38, N471);
nand NAND4 (N718, N710, N696, N522, N643);
not NOT1 (N719, N718);
not NOT1 (N720, N715);
buf BUF1 (N721, N698);
and AND3 (N722, N716, N55, N613);
buf BUF1 (N723, N687);
and AND3 (N724, N711, N294, N423);
not NOT1 (N725, N724);
and AND2 (N726, N720, N77);
or OR3 (N727, N702, N513, N469);
nand NAND2 (N728, N725, N483);
buf BUF1 (N729, N717);
nand NAND2 (N730, N713, N101);
or OR3 (N731, N719, N273, N48);
buf BUF1 (N732, N728);
or OR3 (N733, N730, N240, N304);
or OR2 (N734, N733, N665);
and AND3 (N735, N726, N253, N351);
xor XOR2 (N736, N686, N629);
xor XOR2 (N737, N721, N286);
and AND2 (N738, N723, N158);
buf BUF1 (N739, N735);
xor XOR2 (N740, N729, N1);
nand NAND4 (N741, N732, N19, N206, N192);
nor NOR2 (N742, N722, N95);
not NOT1 (N743, N731);
not NOT1 (N744, N738);
buf BUF1 (N745, N741);
or OR2 (N746, N737, N50);
nor NOR4 (N747, N727, N131, N181, N435);
nor NOR2 (N748, N746, N586);
nand NAND3 (N749, N734, N414, N151);
or OR4 (N750, N742, N405, N40, N679);
or OR4 (N751, N750, N494, N447, N77);
buf BUF1 (N752, N736);
xor XOR2 (N753, N744, N188);
and AND3 (N754, N751, N468, N528);
buf BUF1 (N755, N739);
or OR2 (N756, N754, N332);
nor NOR3 (N757, N755, N147, N350);
buf BUF1 (N758, N753);
xor XOR2 (N759, N757, N481);
nor NOR2 (N760, N758, N85);
not NOT1 (N761, N756);
xor XOR2 (N762, N752, N748);
not NOT1 (N763, N570);
not NOT1 (N764, N760);
buf BUF1 (N765, N740);
or OR3 (N766, N762, N233, N596);
and AND3 (N767, N759, N580, N765);
or OR2 (N768, N542, N598);
not NOT1 (N769, N768);
not NOT1 (N770, N743);
nand NAND4 (N771, N769, N685, N44, N270);
xor XOR2 (N772, N749, N621);
nand NAND3 (N773, N764, N96, N41);
nand NAND2 (N774, N771, N669);
and AND2 (N775, N772, N613);
not NOT1 (N776, N770);
and AND2 (N777, N766, N477);
nand NAND2 (N778, N745, N14);
not NOT1 (N779, N777);
nand NAND3 (N780, N747, N428, N500);
nand NAND4 (N781, N780, N731, N244, N540);
nand NAND4 (N782, N773, N622, N383, N99);
not NOT1 (N783, N767);
nor NOR2 (N784, N779, N26);
not NOT1 (N785, N774);
buf BUF1 (N786, N763);
xor XOR2 (N787, N775, N573);
not NOT1 (N788, N782);
buf BUF1 (N789, N776);
nor NOR4 (N790, N761, N738, N203, N288);
nor NOR3 (N791, N790, N270, N769);
xor XOR2 (N792, N783, N287);
buf BUF1 (N793, N778);
buf BUF1 (N794, N785);
not NOT1 (N795, N791);
xor XOR2 (N796, N792, N559);
xor XOR2 (N797, N795, N443);
not NOT1 (N798, N793);
or OR2 (N799, N796, N322);
or OR3 (N800, N784, N293, N755);
buf BUF1 (N801, N789);
nand NAND3 (N802, N799, N290, N785);
or OR2 (N803, N787, N713);
and AND2 (N804, N801, N599);
and AND3 (N805, N794, N193, N242);
not NOT1 (N806, N804);
or OR4 (N807, N803, N98, N13, N370);
or OR3 (N808, N788, N423, N148);
nor NOR2 (N809, N808, N597);
nand NAND2 (N810, N786, N414);
and AND2 (N811, N800, N563);
buf BUF1 (N812, N806);
or OR3 (N813, N810, N419, N761);
buf BUF1 (N814, N813);
or OR3 (N815, N812, N567, N272);
nor NOR4 (N816, N814, N683, N550, N488);
xor XOR2 (N817, N802, N218);
or OR4 (N818, N816, N349, N400, N85);
buf BUF1 (N819, N807);
buf BUF1 (N820, N805);
xor XOR2 (N821, N820, N664);
and AND2 (N822, N818, N634);
or OR3 (N823, N781, N381, N11);
and AND3 (N824, N797, N501, N510);
buf BUF1 (N825, N811);
nor NOR4 (N826, N821, N99, N251, N144);
not NOT1 (N827, N809);
nor NOR4 (N828, N825, N398, N191, N770);
not NOT1 (N829, N817);
not NOT1 (N830, N798);
nand NAND4 (N831, N824, N109, N355, N499);
and AND3 (N832, N819, N762, N290);
or OR2 (N833, N830, N579);
nand NAND3 (N834, N833, N425, N303);
and AND4 (N835, N822, N205, N439, N769);
and AND2 (N836, N834, N279);
nand NAND3 (N837, N829, N362, N503);
and AND4 (N838, N837, N559, N780, N688);
not NOT1 (N839, N832);
nor NOR3 (N840, N826, N254, N372);
nor NOR4 (N841, N828, N248, N657, N438);
xor XOR2 (N842, N838, N294);
xor XOR2 (N843, N842, N696);
nand NAND4 (N844, N827, N792, N611, N120);
and AND2 (N845, N839, N693);
nand NAND4 (N846, N841, N229, N682, N314);
not NOT1 (N847, N845);
or OR2 (N848, N840, N171);
and AND3 (N849, N815, N625, N524);
or OR3 (N850, N849, N42, N136);
buf BUF1 (N851, N847);
nor NOR3 (N852, N846, N391, N720);
xor XOR2 (N853, N836, N372);
nor NOR4 (N854, N853, N185, N695, N849);
or OR2 (N855, N848, N298);
buf BUF1 (N856, N835);
and AND2 (N857, N855, N321);
or OR2 (N858, N856, N485);
nand NAND2 (N859, N843, N467);
not NOT1 (N860, N858);
nand NAND4 (N861, N851, N94, N750, N784);
xor XOR2 (N862, N831, N646);
buf BUF1 (N863, N859);
nor NOR3 (N864, N860, N182, N88);
buf BUF1 (N865, N850);
nor NOR4 (N866, N864, N83, N191, N45);
xor XOR2 (N867, N852, N612);
buf BUF1 (N868, N823);
xor XOR2 (N869, N863, N189);
nor NOR4 (N870, N866, N830, N145, N482);
nand NAND2 (N871, N867, N12);
and AND4 (N872, N868, N861, N784, N454);
or OR3 (N873, N469, N517, N31);
or OR4 (N874, N857, N505, N707, N237);
buf BUF1 (N875, N869);
not NOT1 (N876, N862);
nor NOR3 (N877, N876, N706, N35);
nor NOR3 (N878, N875, N876, N187);
and AND2 (N879, N871, N233);
not NOT1 (N880, N854);
and AND2 (N881, N870, N610);
nor NOR3 (N882, N880, N563, N115);
xor XOR2 (N883, N882, N539);
and AND2 (N884, N877, N735);
nor NOR3 (N885, N878, N657, N452);
nor NOR3 (N886, N844, N200, N736);
or OR2 (N887, N879, N789);
or OR4 (N888, N881, N542, N793, N810);
nor NOR4 (N889, N888, N693, N673, N197);
nor NOR2 (N890, N874, N204);
nor NOR3 (N891, N865, N198, N421);
or OR2 (N892, N887, N469);
nand NAND2 (N893, N886, N89);
or OR3 (N894, N885, N567, N549);
not NOT1 (N895, N892);
or OR2 (N896, N891, N535);
nor NOR2 (N897, N873, N712);
nor NOR4 (N898, N883, N741, N653, N202);
nand NAND4 (N899, N872, N895, N583, N230);
nor NOR3 (N900, N755, N489, N764);
and AND4 (N901, N896, N571, N149, N40);
and AND3 (N902, N893, N736, N873);
or OR4 (N903, N902, N644, N875, N326);
nand NAND4 (N904, N897, N228, N331, N307);
nand NAND3 (N905, N899, N262, N608);
nand NAND3 (N906, N903, N626, N138);
nand NAND4 (N907, N898, N811, N890, N873);
nor NOR4 (N908, N253, N436, N813, N574);
or OR2 (N909, N908, N443);
and AND3 (N910, N907, N349, N552);
or OR3 (N911, N905, N339, N138);
buf BUF1 (N912, N906);
nand NAND4 (N913, N884, N453, N699, N716);
buf BUF1 (N914, N900);
nor NOR2 (N915, N904, N682);
or OR2 (N916, N894, N433);
nand NAND3 (N917, N910, N746, N106);
or OR3 (N918, N889, N391, N481);
and AND3 (N919, N909, N56, N419);
nand NAND4 (N920, N911, N387, N371, N503);
nor NOR2 (N921, N901, N869);
not NOT1 (N922, N916);
nor NOR3 (N923, N921, N819, N158);
nor NOR2 (N924, N914, N127);
and AND4 (N925, N918, N521, N201, N110);
nand NAND3 (N926, N920, N362, N743);
or OR2 (N927, N925, N42);
and AND4 (N928, N924, N267, N759, N907);
and AND4 (N929, N927, N261, N296, N105);
nand NAND4 (N930, N926, N787, N864, N347);
or OR3 (N931, N919, N452, N786);
xor XOR2 (N932, N931, N519);
or OR2 (N933, N929, N342);
xor XOR2 (N934, N922, N230);
buf BUF1 (N935, N932);
nor NOR3 (N936, N930, N885, N475);
nand NAND4 (N937, N923, N426, N178, N620);
not NOT1 (N938, N935);
not NOT1 (N939, N913);
and AND4 (N940, N937, N763, N567, N161);
buf BUF1 (N941, N934);
and AND2 (N942, N939, N386);
and AND2 (N943, N912, N366);
xor XOR2 (N944, N915, N861);
or OR3 (N945, N936, N321, N139);
not NOT1 (N946, N917);
and AND3 (N947, N945, N885, N182);
nand NAND2 (N948, N941, N132);
not NOT1 (N949, N947);
nand NAND2 (N950, N938, N586);
buf BUF1 (N951, N942);
or OR4 (N952, N943, N641, N388, N688);
and AND3 (N953, N928, N174, N493);
buf BUF1 (N954, N948);
nand NAND2 (N955, N949, N648);
not NOT1 (N956, N950);
buf BUF1 (N957, N951);
not NOT1 (N958, N940);
xor XOR2 (N959, N944, N40);
nand NAND4 (N960, N946, N610, N182, N782);
buf BUF1 (N961, N953);
buf BUF1 (N962, N933);
nor NOR4 (N963, N954, N957, N943, N767);
nor NOR4 (N964, N580, N704, N350, N744);
xor XOR2 (N965, N958, N15);
not NOT1 (N966, N952);
buf BUF1 (N967, N963);
nor NOR3 (N968, N965, N900, N143);
or OR3 (N969, N967, N46, N364);
and AND3 (N970, N969, N484, N322);
nor NOR2 (N971, N956, N951);
buf BUF1 (N972, N962);
not NOT1 (N973, N960);
nor NOR4 (N974, N968, N197, N896, N392);
nor NOR3 (N975, N974, N530, N735);
nand NAND3 (N976, N975, N755, N871);
xor XOR2 (N977, N972, N282);
nand NAND3 (N978, N964, N817, N736);
buf BUF1 (N979, N973);
xor XOR2 (N980, N970, N473);
and AND4 (N981, N966, N44, N133, N956);
not NOT1 (N982, N971);
not NOT1 (N983, N977);
nor NOR3 (N984, N982, N344, N217);
or OR3 (N985, N984, N564, N643);
or OR3 (N986, N955, N874, N827);
or OR4 (N987, N959, N233, N914, N607);
not NOT1 (N988, N980);
buf BUF1 (N989, N985);
or OR4 (N990, N978, N374, N863, N500);
not NOT1 (N991, N981);
or OR2 (N992, N976, N902);
nor NOR3 (N993, N987, N185, N518);
xor XOR2 (N994, N992, N118);
or OR3 (N995, N988, N485, N684);
not NOT1 (N996, N961);
buf BUF1 (N997, N986);
nor NOR4 (N998, N996, N730, N435, N765);
nor NOR3 (N999, N991, N303, N83);
or OR4 (N1000, N993, N122, N396, N558);
nand NAND2 (N1001, N1000, N25);
nand NAND3 (N1002, N983, N898, N690);
or OR4 (N1003, N1001, N280, N874, N178);
or OR3 (N1004, N995, N198, N555);
xor XOR2 (N1005, N999, N476);
nand NAND3 (N1006, N998, N818, N263);
not NOT1 (N1007, N989);
xor XOR2 (N1008, N1003, N21);
xor XOR2 (N1009, N990, N264);
and AND3 (N1010, N1007, N932, N671);
buf BUF1 (N1011, N1008);
not NOT1 (N1012, N1002);
or OR4 (N1013, N994, N409, N1, N270);
nand NAND2 (N1014, N1005, N688);
nand NAND4 (N1015, N1010, N444, N835, N671);
xor XOR2 (N1016, N1009, N797);
nand NAND2 (N1017, N997, N512);
xor XOR2 (N1018, N979, N673);
nor NOR4 (N1019, N1011, N65, N483, N85);
nor NOR4 (N1020, N1004, N779, N97, N100);
nor NOR2 (N1021, N1018, N626);
nor NOR4 (N1022, N1020, N337, N560, N806);
xor XOR2 (N1023, N1014, N39);
and AND2 (N1024, N1012, N848);
or OR2 (N1025, N1024, N416);
nand NAND2 (N1026, N1025, N940);
or OR3 (N1027, N1021, N573, N390);
not NOT1 (N1028, N1023);
not NOT1 (N1029, N1013);
nand NAND2 (N1030, N1028, N808);
buf BUF1 (N1031, N1015);
not NOT1 (N1032, N1006);
buf BUF1 (N1033, N1016);
and AND4 (N1034, N1027, N131, N113, N49);
and AND3 (N1035, N1026, N215, N123);
nor NOR2 (N1036, N1029, N1016);
and AND4 (N1037, N1030, N492, N792, N163);
xor XOR2 (N1038, N1031, N986);
xor XOR2 (N1039, N1022, N290);
not NOT1 (N1040, N1038);
and AND4 (N1041, N1037, N793, N58, N12);
and AND4 (N1042, N1032, N1021, N152, N378);
xor XOR2 (N1043, N1042, N307);
or OR3 (N1044, N1035, N360, N724);
xor XOR2 (N1045, N1017, N264);
xor XOR2 (N1046, N1033, N536);
nand NAND4 (N1047, N1034, N218, N527, N54);
or OR3 (N1048, N1040, N460, N387);
and AND2 (N1049, N1036, N234);
xor XOR2 (N1050, N1044, N409);
nand NAND3 (N1051, N1041, N389, N842);
nor NOR2 (N1052, N1050, N684);
or OR3 (N1053, N1039, N16, N557);
nand NAND4 (N1054, N1051, N231, N501, N302);
not NOT1 (N1055, N1049);
not NOT1 (N1056, N1048);
nand NAND3 (N1057, N1046, N875, N78);
not NOT1 (N1058, N1057);
xor XOR2 (N1059, N1047, N260);
xor XOR2 (N1060, N1053, N57);
not NOT1 (N1061, N1054);
buf BUF1 (N1062, N1056);
xor XOR2 (N1063, N1052, N576);
or OR3 (N1064, N1043, N449, N128);
and AND2 (N1065, N1055, N878);
nor NOR3 (N1066, N1058, N940, N382);
buf BUF1 (N1067, N1060);
nor NOR4 (N1068, N1067, N207, N299, N664);
nand NAND3 (N1069, N1068, N301, N161);
or OR3 (N1070, N1065, N364, N25);
and AND3 (N1071, N1066, N810, N732);
or OR3 (N1072, N1061, N395, N233);
nand NAND4 (N1073, N1064, N112, N147, N888);
or OR2 (N1074, N1019, N458);
nand NAND2 (N1075, N1062, N627);
buf BUF1 (N1076, N1045);
nand NAND3 (N1077, N1069, N538, N789);
or OR4 (N1078, N1059, N762, N403, N704);
nand NAND4 (N1079, N1073, N446, N985, N930);
or OR4 (N1080, N1076, N1016, N827, N928);
or OR2 (N1081, N1072, N844);
xor XOR2 (N1082, N1078, N246);
not NOT1 (N1083, N1063);
nand NAND2 (N1084, N1079, N625);
nor NOR4 (N1085, N1077, N989, N211, N1021);
not NOT1 (N1086, N1083);
nand NAND3 (N1087, N1074, N443, N1034);
or OR3 (N1088, N1085, N537, N84);
or OR3 (N1089, N1080, N955, N767);
or OR3 (N1090, N1071, N147, N795);
or OR3 (N1091, N1075, N277, N737);
or OR3 (N1092, N1091, N236, N225);
nor NOR3 (N1093, N1092, N738, N846);
or OR4 (N1094, N1081, N44, N837, N542);
and AND3 (N1095, N1088, N368, N25);
not NOT1 (N1096, N1094);
or OR3 (N1097, N1084, N1026, N130);
nand NAND4 (N1098, N1096, N444, N971, N709);
buf BUF1 (N1099, N1089);
or OR2 (N1100, N1087, N781);
or OR3 (N1101, N1099, N151, N1079);
nor NOR3 (N1102, N1093, N674, N942);
buf BUF1 (N1103, N1090);
nor NOR2 (N1104, N1098, N1017);
buf BUF1 (N1105, N1082);
nand NAND3 (N1106, N1103, N732, N431);
not NOT1 (N1107, N1105);
or OR4 (N1108, N1106, N541, N1025, N616);
not NOT1 (N1109, N1070);
nor NOR2 (N1110, N1097, N786);
not NOT1 (N1111, N1109);
nand NAND3 (N1112, N1095, N600, N232);
not NOT1 (N1113, N1111);
buf BUF1 (N1114, N1112);
or OR3 (N1115, N1086, N902, N776);
not NOT1 (N1116, N1115);
or OR4 (N1117, N1108, N907, N639, N919);
buf BUF1 (N1118, N1107);
buf BUF1 (N1119, N1100);
nor NOR4 (N1120, N1119, N88, N334, N876);
nor NOR2 (N1121, N1102, N61);
buf BUF1 (N1122, N1113);
buf BUF1 (N1123, N1122);
not NOT1 (N1124, N1101);
not NOT1 (N1125, N1110);
nand NAND3 (N1126, N1123, N678, N279);
nor NOR2 (N1127, N1104, N411);
buf BUF1 (N1128, N1117);
and AND2 (N1129, N1126, N595);
not NOT1 (N1130, N1127);
and AND3 (N1131, N1118, N359, N541);
and AND2 (N1132, N1124, N462);
buf BUF1 (N1133, N1114);
xor XOR2 (N1134, N1129, N738);
not NOT1 (N1135, N1121);
or OR4 (N1136, N1132, N72, N796, N419);
not NOT1 (N1137, N1135);
or OR3 (N1138, N1116, N461, N72);
nor NOR4 (N1139, N1133, N181, N78, N826);
nand NAND4 (N1140, N1125, N883, N1022, N15);
not NOT1 (N1141, N1136);
nor NOR3 (N1142, N1140, N939, N556);
not NOT1 (N1143, N1134);
nor NOR4 (N1144, N1130, N696, N1084, N708);
nand NAND3 (N1145, N1139, N213, N621);
buf BUF1 (N1146, N1120);
buf BUF1 (N1147, N1128);
buf BUF1 (N1148, N1146);
buf BUF1 (N1149, N1131);
xor XOR2 (N1150, N1138, N691);
buf BUF1 (N1151, N1137);
buf BUF1 (N1152, N1147);
and AND2 (N1153, N1150, N375);
xor XOR2 (N1154, N1145, N226);
or OR4 (N1155, N1148, N695, N491, N977);
or OR2 (N1156, N1142, N821);
not NOT1 (N1157, N1143);
xor XOR2 (N1158, N1151, N585);
or OR3 (N1159, N1156, N65, N997);
buf BUF1 (N1160, N1154);
nor NOR3 (N1161, N1155, N816, N390);
nand NAND2 (N1162, N1158, N281);
xor XOR2 (N1163, N1144, N1057);
nor NOR4 (N1164, N1152, N299, N965, N156);
and AND3 (N1165, N1153, N713, N113);
or OR4 (N1166, N1163, N739, N667, N551);
not NOT1 (N1167, N1166);
xor XOR2 (N1168, N1149, N1054);
not NOT1 (N1169, N1159);
xor XOR2 (N1170, N1168, N281);
buf BUF1 (N1171, N1169);
nor NOR4 (N1172, N1161, N331, N1164, N446);
xor XOR2 (N1173, N312, N55);
and AND4 (N1174, N1171, N28, N648, N526);
nand NAND4 (N1175, N1141, N350, N169, N307);
nor NOR2 (N1176, N1170, N916);
not NOT1 (N1177, N1157);
xor XOR2 (N1178, N1167, N350);
or OR2 (N1179, N1176, N790);
nor NOR4 (N1180, N1178, N850, N709, N222);
not NOT1 (N1181, N1162);
not NOT1 (N1182, N1177);
not NOT1 (N1183, N1173);
buf BUF1 (N1184, N1180);
or OR2 (N1185, N1172, N1040);
nor NOR4 (N1186, N1182, N744, N1185, N188);
not NOT1 (N1187, N797);
nand NAND2 (N1188, N1181, N1011);
not NOT1 (N1189, N1160);
nor NOR3 (N1190, N1174, N861, N909);
nand NAND4 (N1191, N1187, N93, N671, N205);
nor NOR3 (N1192, N1190, N530, N477);
buf BUF1 (N1193, N1184);
nor NOR2 (N1194, N1165, N26);
nand NAND4 (N1195, N1188, N915, N831, N58);
buf BUF1 (N1196, N1189);
and AND4 (N1197, N1179, N71, N32, N86);
nand NAND4 (N1198, N1192, N1044, N528, N1156);
nor NOR2 (N1199, N1175, N637);
or OR4 (N1200, N1198, N865, N715, N345);
nor NOR3 (N1201, N1197, N375, N633);
nor NOR4 (N1202, N1194, N168, N4, N1195);
buf BUF1 (N1203, N395);
and AND3 (N1204, N1186, N649, N86);
not NOT1 (N1205, N1196);
buf BUF1 (N1206, N1200);
nor NOR2 (N1207, N1202, N1016);
not NOT1 (N1208, N1206);
nor NOR4 (N1209, N1193, N103, N248, N672);
nand NAND2 (N1210, N1208, N789);
and AND4 (N1211, N1205, N249, N499, N1195);
buf BUF1 (N1212, N1210);
buf BUF1 (N1213, N1204);
xor XOR2 (N1214, N1199, N694);
nand NAND4 (N1215, N1207, N597, N261, N326);
buf BUF1 (N1216, N1203);
or OR4 (N1217, N1191, N595, N52, N800);
nand NAND3 (N1218, N1209, N792, N137);
buf BUF1 (N1219, N1215);
not NOT1 (N1220, N1211);
xor XOR2 (N1221, N1220, N268);
buf BUF1 (N1222, N1214);
and AND4 (N1223, N1221, N559, N946, N941);
or OR3 (N1224, N1216, N924, N179);
not NOT1 (N1225, N1183);
nor NOR4 (N1226, N1219, N1060, N1077, N874);
or OR4 (N1227, N1201, N155, N739, N667);
not NOT1 (N1228, N1226);
and AND4 (N1229, N1217, N555, N1197, N732);
nor NOR2 (N1230, N1229, N401);
and AND4 (N1231, N1228, N612, N111, N560);
not NOT1 (N1232, N1230);
nor NOR4 (N1233, N1223, N349, N396, N432);
nand NAND3 (N1234, N1212, N554, N224);
or OR3 (N1235, N1213, N360, N1145);
buf BUF1 (N1236, N1234);
nand NAND2 (N1237, N1227, N102);
nand NAND2 (N1238, N1231, N336);
not NOT1 (N1239, N1233);
nor NOR3 (N1240, N1237, N22, N819);
xor XOR2 (N1241, N1218, N62);
xor XOR2 (N1242, N1239, N903);
and AND2 (N1243, N1225, N581);
nand NAND2 (N1244, N1238, N834);
and AND2 (N1245, N1242, N124);
nand NAND3 (N1246, N1240, N869, N656);
and AND3 (N1247, N1222, N804, N381);
not NOT1 (N1248, N1236);
nand NAND3 (N1249, N1235, N294, N832);
xor XOR2 (N1250, N1246, N942);
nor NOR2 (N1251, N1245, N261);
buf BUF1 (N1252, N1232);
nand NAND3 (N1253, N1224, N551, N333);
and AND2 (N1254, N1248, N984);
xor XOR2 (N1255, N1244, N543);
and AND3 (N1256, N1241, N863, N224);
not NOT1 (N1257, N1251);
not NOT1 (N1258, N1249);
nand NAND4 (N1259, N1255, N143, N331, N739);
nor NOR4 (N1260, N1250, N810, N546, N267);
not NOT1 (N1261, N1252);
buf BUF1 (N1262, N1257);
nand NAND4 (N1263, N1262, N1071, N860, N198);
buf BUF1 (N1264, N1253);
or OR4 (N1265, N1261, N187, N1246, N261);
not NOT1 (N1266, N1247);
buf BUF1 (N1267, N1258);
nand NAND2 (N1268, N1267, N1055);
and AND2 (N1269, N1254, N574);
and AND3 (N1270, N1266, N241, N518);
nor NOR3 (N1271, N1268, N802, N1042);
xor XOR2 (N1272, N1269, N55);
buf BUF1 (N1273, N1271);
or OR2 (N1274, N1259, N873);
buf BUF1 (N1275, N1274);
buf BUF1 (N1276, N1270);
or OR4 (N1277, N1264, N999, N380, N423);
or OR3 (N1278, N1243, N1155, N1161);
or OR3 (N1279, N1275, N892, N1220);
not NOT1 (N1280, N1278);
not NOT1 (N1281, N1272);
xor XOR2 (N1282, N1256, N10);
or OR2 (N1283, N1276, N659);
or OR4 (N1284, N1273, N117, N325, N403);
buf BUF1 (N1285, N1277);
or OR4 (N1286, N1260, N1013, N457, N96);
buf BUF1 (N1287, N1280);
and AND4 (N1288, N1265, N733, N571, N676);
and AND2 (N1289, N1279, N341);
or OR2 (N1290, N1287, N1249);
not NOT1 (N1291, N1290);
nor NOR2 (N1292, N1291, N403);
or OR2 (N1293, N1288, N820);
buf BUF1 (N1294, N1289);
buf BUF1 (N1295, N1285);
nor NOR3 (N1296, N1286, N331, N1238);
or OR4 (N1297, N1293, N708, N625, N901);
xor XOR2 (N1298, N1297, N343);
xor XOR2 (N1299, N1295, N335);
xor XOR2 (N1300, N1263, N1232);
not NOT1 (N1301, N1283);
nand NAND4 (N1302, N1301, N341, N651, N214);
not NOT1 (N1303, N1302);
xor XOR2 (N1304, N1292, N343);
nor NOR4 (N1305, N1304, N1135, N454, N1134);
and AND2 (N1306, N1296, N891);
xor XOR2 (N1307, N1298, N608);
buf BUF1 (N1308, N1294);
and AND2 (N1309, N1281, N1155);
xor XOR2 (N1310, N1300, N581);
nor NOR3 (N1311, N1303, N819, N878);
nand NAND4 (N1312, N1299, N264, N975, N302);
and AND3 (N1313, N1282, N1177, N961);
buf BUF1 (N1314, N1308);
or OR4 (N1315, N1311, N749, N463, N1013);
or OR3 (N1316, N1306, N1028, N1187);
nand NAND4 (N1317, N1314, N823, N1288, N1021);
not NOT1 (N1318, N1317);
nor NOR3 (N1319, N1307, N529, N337);
nor NOR2 (N1320, N1312, N1259);
and AND2 (N1321, N1316, N332);
not NOT1 (N1322, N1309);
buf BUF1 (N1323, N1321);
nor NOR3 (N1324, N1323, N318, N937);
or OR3 (N1325, N1319, N1067, N322);
or OR3 (N1326, N1325, N900, N1012);
nor NOR3 (N1327, N1305, N1186, N978);
and AND3 (N1328, N1318, N1265, N1283);
xor XOR2 (N1329, N1322, N932);
buf BUF1 (N1330, N1324);
and AND2 (N1331, N1313, N610);
buf BUF1 (N1332, N1327);
and AND3 (N1333, N1329, N550, N717);
nand NAND3 (N1334, N1320, N662, N221);
not NOT1 (N1335, N1332);
or OR2 (N1336, N1334, N132);
and AND3 (N1337, N1328, N1084, N1213);
not NOT1 (N1338, N1336);
not NOT1 (N1339, N1331);
nand NAND4 (N1340, N1326, N1308, N627, N32);
nand NAND4 (N1341, N1284, N1244, N1022, N810);
nor NOR3 (N1342, N1340, N122, N785);
nand NAND2 (N1343, N1338, N993);
buf BUF1 (N1344, N1335);
nor NOR3 (N1345, N1343, N497, N608);
buf BUF1 (N1346, N1315);
nand NAND3 (N1347, N1344, N640, N495);
buf BUF1 (N1348, N1310);
and AND3 (N1349, N1333, N309, N363);
buf BUF1 (N1350, N1349);
nand NAND2 (N1351, N1346, N354);
nand NAND3 (N1352, N1351, N721, N735);
not NOT1 (N1353, N1348);
nor NOR2 (N1354, N1350, N162);
buf BUF1 (N1355, N1353);
nand NAND3 (N1356, N1342, N1337, N1184);
nand NAND3 (N1357, N684, N288, N1356);
buf BUF1 (N1358, N1317);
xor XOR2 (N1359, N1341, N1291);
and AND4 (N1360, N1358, N999, N1140, N1014);
or OR2 (N1361, N1359, N31);
buf BUF1 (N1362, N1361);
xor XOR2 (N1363, N1362, N350);
or OR3 (N1364, N1339, N170, N147);
xor XOR2 (N1365, N1360, N720);
nand NAND3 (N1366, N1347, N389, N1344);
xor XOR2 (N1367, N1366, N1364);
xor XOR2 (N1368, N1272, N944);
xor XOR2 (N1369, N1354, N153);
not NOT1 (N1370, N1355);
not NOT1 (N1371, N1345);
and AND3 (N1372, N1369, N422, N991);
and AND4 (N1373, N1371, N640, N825, N414);
and AND4 (N1374, N1363, N1278, N188, N760);
buf BUF1 (N1375, N1372);
not NOT1 (N1376, N1330);
nand NAND4 (N1377, N1357, N833, N1299, N1285);
not NOT1 (N1378, N1370);
or OR3 (N1379, N1367, N710, N43);
and AND2 (N1380, N1352, N912);
or OR3 (N1381, N1379, N390, N884);
or OR4 (N1382, N1376, N890, N1181, N1277);
nor NOR2 (N1383, N1368, N576);
and AND3 (N1384, N1377, N124, N841);
and AND3 (N1385, N1373, N1343, N1176);
or OR2 (N1386, N1383, N1224);
and AND3 (N1387, N1378, N418, N326);
and AND2 (N1388, N1375, N646);
xor XOR2 (N1389, N1385, N1251);
buf BUF1 (N1390, N1381);
xor XOR2 (N1391, N1384, N132);
not NOT1 (N1392, N1391);
buf BUF1 (N1393, N1390);
buf BUF1 (N1394, N1393);
xor XOR2 (N1395, N1387, N1378);
not NOT1 (N1396, N1389);
nand NAND4 (N1397, N1394, N816, N453, N773);
and AND2 (N1398, N1386, N757);
or OR4 (N1399, N1397, N487, N1063, N1124);
xor XOR2 (N1400, N1399, N725);
nor NOR4 (N1401, N1380, N367, N1258, N1213);
buf BUF1 (N1402, N1365);
nand NAND4 (N1403, N1395, N1300, N837, N610);
or OR4 (N1404, N1402, N1185, N131, N663);
or OR3 (N1405, N1404, N1125, N300);
xor XOR2 (N1406, N1405, N1269);
buf BUF1 (N1407, N1401);
not NOT1 (N1408, N1396);
xor XOR2 (N1409, N1388, N844);
nor NOR3 (N1410, N1403, N1078, N296);
buf BUF1 (N1411, N1374);
nor NOR2 (N1412, N1411, N1146);
buf BUF1 (N1413, N1407);
xor XOR2 (N1414, N1408, N550);
nor NOR2 (N1415, N1409, N1183);
nand NAND3 (N1416, N1415, N200, N100);
nand NAND4 (N1417, N1414, N624, N1400, N171);
buf BUF1 (N1418, N908);
buf BUF1 (N1419, N1410);
nand NAND3 (N1420, N1419, N1017, N475);
nand NAND2 (N1421, N1418, N243);
nand NAND4 (N1422, N1420, N768, N929, N741);
nand NAND2 (N1423, N1422, N446);
xor XOR2 (N1424, N1417, N462);
nor NOR3 (N1425, N1412, N714, N1050);
and AND3 (N1426, N1398, N846, N909);
nand NAND3 (N1427, N1425, N603, N867);
xor XOR2 (N1428, N1413, N980);
not NOT1 (N1429, N1421);
or OR4 (N1430, N1428, N1066, N98, N1194);
not NOT1 (N1431, N1426);
buf BUF1 (N1432, N1424);
xor XOR2 (N1433, N1432, N749);
or OR4 (N1434, N1382, N1230, N1266, N1190);
buf BUF1 (N1435, N1423);
xor XOR2 (N1436, N1430, N1165);
nor NOR2 (N1437, N1434, N304);
xor XOR2 (N1438, N1429, N243);
nor NOR4 (N1439, N1438, N1240, N1229, N38);
not NOT1 (N1440, N1439);
nand NAND2 (N1441, N1431, N139);
buf BUF1 (N1442, N1440);
and AND4 (N1443, N1406, N647, N1106, N390);
not NOT1 (N1444, N1441);
xor XOR2 (N1445, N1444, N101);
nand NAND2 (N1446, N1433, N553);
and AND2 (N1447, N1427, N218);
nand NAND4 (N1448, N1437, N777, N1315, N518);
buf BUF1 (N1449, N1446);
and AND4 (N1450, N1445, N1031, N165, N1405);
xor XOR2 (N1451, N1449, N1436);
or OR4 (N1452, N911, N1028, N709, N258);
nor NOR4 (N1453, N1435, N1135, N1260, N1062);
nand NAND2 (N1454, N1447, N1436);
buf BUF1 (N1455, N1450);
and AND4 (N1456, N1452, N1265, N881, N1326);
xor XOR2 (N1457, N1416, N409);
not NOT1 (N1458, N1457);
or OR2 (N1459, N1454, N462);
not NOT1 (N1460, N1392);
or OR2 (N1461, N1442, N823);
xor XOR2 (N1462, N1455, N129);
not NOT1 (N1463, N1458);
nor NOR3 (N1464, N1462, N800, N36);
nand NAND4 (N1465, N1460, N1211, N554, N1240);
xor XOR2 (N1466, N1448, N323);
nor NOR3 (N1467, N1465, N324, N1432);
xor XOR2 (N1468, N1464, N540);
not NOT1 (N1469, N1467);
nor NOR2 (N1470, N1469, N508);
buf BUF1 (N1471, N1451);
not NOT1 (N1472, N1466);
xor XOR2 (N1473, N1463, N84);
nand NAND2 (N1474, N1468, N1156);
not NOT1 (N1475, N1459);
and AND2 (N1476, N1453, N903);
buf BUF1 (N1477, N1461);
nand NAND2 (N1478, N1471, N594);
not NOT1 (N1479, N1470);
nor NOR2 (N1480, N1456, N1439);
buf BUF1 (N1481, N1476);
buf BUF1 (N1482, N1472);
nor NOR4 (N1483, N1480, N561, N392, N928);
not NOT1 (N1484, N1481);
not NOT1 (N1485, N1483);
not NOT1 (N1486, N1484);
xor XOR2 (N1487, N1443, N783);
not NOT1 (N1488, N1479);
nor NOR4 (N1489, N1473, N308, N999, N112);
buf BUF1 (N1490, N1477);
nor NOR3 (N1491, N1478, N367, N1251);
not NOT1 (N1492, N1482);
or OR2 (N1493, N1474, N1112);
xor XOR2 (N1494, N1492, N686);
not NOT1 (N1495, N1488);
nor NOR3 (N1496, N1485, N942, N146);
nor NOR3 (N1497, N1494, N828, N1048);
or OR4 (N1498, N1491, N784, N1305, N103);
or OR3 (N1499, N1487, N556, N520);
nand NAND2 (N1500, N1493, N1120);
or OR3 (N1501, N1486, N1146, N270);
not NOT1 (N1502, N1496);
nand NAND2 (N1503, N1475, N1384);
or OR4 (N1504, N1498, N409, N271, N225);
xor XOR2 (N1505, N1495, N1318);
and AND2 (N1506, N1489, N1378);
buf BUF1 (N1507, N1503);
nor NOR4 (N1508, N1506, N429, N1039, N452);
not NOT1 (N1509, N1501);
or OR3 (N1510, N1505, N1460, N59);
and AND3 (N1511, N1502, N1414, N30);
and AND4 (N1512, N1500, N853, N974, N97);
or OR2 (N1513, N1490, N895);
xor XOR2 (N1514, N1499, N198);
xor XOR2 (N1515, N1512, N967);
and AND3 (N1516, N1507, N5, N537);
nor NOR4 (N1517, N1516, N542, N886, N903);
buf BUF1 (N1518, N1513);
nor NOR2 (N1519, N1511, N1340);
or OR3 (N1520, N1518, N462, N1414);
nand NAND4 (N1521, N1504, N388, N77, N873);
buf BUF1 (N1522, N1509);
nor NOR4 (N1523, N1519, N1201, N239, N495);
or OR4 (N1524, N1521, N1114, N1484, N1357);
nand NAND4 (N1525, N1514, N676, N38, N1389);
nor NOR3 (N1526, N1522, N424, N117);
nand NAND4 (N1527, N1525, N805, N233, N1267);
nor NOR2 (N1528, N1508, N171);
buf BUF1 (N1529, N1527);
not NOT1 (N1530, N1526);
and AND2 (N1531, N1497, N1516);
not NOT1 (N1532, N1517);
or OR2 (N1533, N1531, N869);
nand NAND3 (N1534, N1533, N1353, N1419);
nor NOR3 (N1535, N1529, N226, N1419);
and AND3 (N1536, N1515, N616, N117);
or OR2 (N1537, N1524, N1145);
nand NAND3 (N1538, N1535, N605, N854);
or OR3 (N1539, N1534, N568, N312);
not NOT1 (N1540, N1528);
not NOT1 (N1541, N1510);
xor XOR2 (N1542, N1537, N903);
xor XOR2 (N1543, N1540, N624);
nor NOR3 (N1544, N1543, N717, N106);
and AND4 (N1545, N1541, N625, N873, N901);
not NOT1 (N1546, N1544);
nor NOR4 (N1547, N1530, N158, N956, N258);
not NOT1 (N1548, N1520);
not NOT1 (N1549, N1548);
nand NAND2 (N1550, N1536, N372);
not NOT1 (N1551, N1532);
or OR3 (N1552, N1547, N1100, N309);
and AND2 (N1553, N1551, N617);
xor XOR2 (N1554, N1546, N1343);
nand NAND3 (N1555, N1542, N1058, N403);
buf BUF1 (N1556, N1545);
or OR4 (N1557, N1555, N443, N1056, N607);
or OR4 (N1558, N1556, N751, N484, N949);
or OR2 (N1559, N1558, N478);
nor NOR4 (N1560, N1523, N319, N352, N1196);
xor XOR2 (N1561, N1557, N928);
xor XOR2 (N1562, N1559, N477);
or OR2 (N1563, N1538, N1452);
not NOT1 (N1564, N1562);
nand NAND4 (N1565, N1553, N560, N301, N1172);
not NOT1 (N1566, N1560);
nand NAND3 (N1567, N1566, N438, N1151);
xor XOR2 (N1568, N1549, N801);
and AND2 (N1569, N1564, N1194);
or OR4 (N1570, N1568, N1395, N1341, N660);
and AND3 (N1571, N1554, N1477, N294);
nand NAND3 (N1572, N1539, N422, N1444);
xor XOR2 (N1573, N1563, N845);
not NOT1 (N1574, N1567);
nand NAND3 (N1575, N1565, N862, N648);
xor XOR2 (N1576, N1572, N129);
not NOT1 (N1577, N1576);
buf BUF1 (N1578, N1573);
xor XOR2 (N1579, N1571, N413);
and AND4 (N1580, N1569, N1505, N290, N1257);
and AND2 (N1581, N1580, N186);
or OR3 (N1582, N1577, N28, N384);
not NOT1 (N1583, N1552);
nand NAND3 (N1584, N1550, N549, N356);
nand NAND3 (N1585, N1581, N1150, N1123);
nand NAND2 (N1586, N1570, N1285);
nand NAND2 (N1587, N1586, N451);
nand NAND2 (N1588, N1579, N1106);
or OR2 (N1589, N1588, N616);
not NOT1 (N1590, N1585);
buf BUF1 (N1591, N1584);
nor NOR4 (N1592, N1583, N1468, N1087, N1456);
nand NAND3 (N1593, N1590, N325, N886);
and AND3 (N1594, N1593, N131, N172);
and AND4 (N1595, N1591, N1225, N1167, N1);
nand NAND2 (N1596, N1574, N1231);
nor NOR3 (N1597, N1582, N1409, N205);
xor XOR2 (N1598, N1594, N1302);
buf BUF1 (N1599, N1592);
xor XOR2 (N1600, N1597, N1148);
nand NAND4 (N1601, N1575, N1262, N75, N656);
or OR4 (N1602, N1600, N713, N1547, N857);
nand NAND4 (N1603, N1601, N239, N1177, N1122);
not NOT1 (N1604, N1599);
not NOT1 (N1605, N1587);
and AND3 (N1606, N1589, N651, N1061);
nor NOR3 (N1607, N1605, N1523, N1103);
or OR2 (N1608, N1607, N1052);
and AND4 (N1609, N1598, N382, N1130, N971);
buf BUF1 (N1610, N1603);
not NOT1 (N1611, N1561);
or OR2 (N1612, N1604, N594);
nand NAND3 (N1613, N1608, N407, N1123);
xor XOR2 (N1614, N1613, N819);
not NOT1 (N1615, N1595);
xor XOR2 (N1616, N1610, N1507);
and AND2 (N1617, N1578, N1094);
nand NAND2 (N1618, N1616, N1025);
and AND2 (N1619, N1606, N1267);
xor XOR2 (N1620, N1619, N363);
nor NOR4 (N1621, N1612, N1066, N1203, N1434);
nand NAND3 (N1622, N1602, N348, N499);
nand NAND3 (N1623, N1618, N857, N1439);
or OR3 (N1624, N1611, N62, N1577);
buf BUF1 (N1625, N1623);
or OR2 (N1626, N1617, N639);
not NOT1 (N1627, N1609);
buf BUF1 (N1628, N1622);
nand NAND2 (N1629, N1615, N555);
and AND2 (N1630, N1627, N271);
nor NOR2 (N1631, N1596, N874);
xor XOR2 (N1632, N1628, N1121);
and AND2 (N1633, N1614, N1277);
buf BUF1 (N1634, N1631);
or OR4 (N1635, N1629, N413, N1527, N586);
or OR3 (N1636, N1625, N8, N280);
nand NAND4 (N1637, N1630, N1457, N1371, N1120);
not NOT1 (N1638, N1620);
buf BUF1 (N1639, N1633);
buf BUF1 (N1640, N1639);
and AND2 (N1641, N1638, N35);
not NOT1 (N1642, N1635);
and AND4 (N1643, N1624, N817, N200, N85);
not NOT1 (N1644, N1626);
buf BUF1 (N1645, N1642);
and AND4 (N1646, N1644, N633, N570, N353);
nor NOR4 (N1647, N1621, N510, N1498, N85);
buf BUF1 (N1648, N1637);
nor NOR3 (N1649, N1648, N238, N1159);
nand NAND4 (N1650, N1649, N493, N87, N1616);
or OR4 (N1651, N1650, N60, N154, N881);
xor XOR2 (N1652, N1634, N748);
buf BUF1 (N1653, N1647);
xor XOR2 (N1654, N1640, N861);
buf BUF1 (N1655, N1645);
not NOT1 (N1656, N1632);
or OR3 (N1657, N1653, N897, N994);
xor XOR2 (N1658, N1655, N259);
not NOT1 (N1659, N1641);
and AND4 (N1660, N1656, N1229, N66, N1127);
buf BUF1 (N1661, N1652);
or OR4 (N1662, N1651, N101, N1633, N471);
and AND4 (N1663, N1636, N1097, N1017, N489);
or OR3 (N1664, N1654, N902, N126);
not NOT1 (N1665, N1662);
nand NAND2 (N1666, N1663, N975);
not NOT1 (N1667, N1664);
buf BUF1 (N1668, N1659);
nor NOR4 (N1669, N1665, N777, N123, N571);
and AND4 (N1670, N1643, N1347, N832, N1202);
nor NOR2 (N1671, N1658, N434);
or OR4 (N1672, N1666, N1369, N1632, N152);
buf BUF1 (N1673, N1671);
or OR4 (N1674, N1670, N1251, N827, N1373);
nor NOR2 (N1675, N1674, N1584);
and AND2 (N1676, N1669, N617);
nand NAND2 (N1677, N1661, N41);
nand NAND3 (N1678, N1676, N1195, N1591);
nor NOR2 (N1679, N1678, N1603);
or OR4 (N1680, N1677, N1476, N1024, N1286);
buf BUF1 (N1681, N1646);
nand NAND3 (N1682, N1660, N1439, N1085);
xor XOR2 (N1683, N1657, N542);
buf BUF1 (N1684, N1679);
nor NOR3 (N1685, N1673, N1252, N227);
or OR3 (N1686, N1684, N9, N1408);
not NOT1 (N1687, N1686);
not NOT1 (N1688, N1667);
not NOT1 (N1689, N1682);
nand NAND3 (N1690, N1672, N162, N31);
xor XOR2 (N1691, N1685, N1084);
nor NOR4 (N1692, N1683, N243, N981, N1392);
nor NOR2 (N1693, N1687, N621);
or OR2 (N1694, N1691, N554);
nor NOR2 (N1695, N1694, N1300);
and AND3 (N1696, N1668, N286, N247);
and AND3 (N1697, N1688, N1405, N572);
xor XOR2 (N1698, N1689, N923);
nand NAND2 (N1699, N1697, N705);
or OR2 (N1700, N1692, N1222);
or OR2 (N1701, N1680, N348);
nor NOR4 (N1702, N1681, N532, N1228, N905);
nor NOR4 (N1703, N1690, N896, N630, N369);
nand NAND2 (N1704, N1700, N1686);
nor NOR2 (N1705, N1693, N1452);
and AND4 (N1706, N1696, N1181, N172, N900);
not NOT1 (N1707, N1698);
and AND4 (N1708, N1706, N200, N112, N1285);
and AND3 (N1709, N1703, N170, N1457);
buf BUF1 (N1710, N1702);
and AND2 (N1711, N1704, N527);
buf BUF1 (N1712, N1705);
buf BUF1 (N1713, N1699);
nor NOR2 (N1714, N1707, N1018);
buf BUF1 (N1715, N1710);
buf BUF1 (N1716, N1715);
nor NOR3 (N1717, N1695, N391, N1263);
nand NAND2 (N1718, N1701, N1505);
nor NOR3 (N1719, N1718, N645, N859);
nor NOR3 (N1720, N1675, N1093, N1310);
or OR4 (N1721, N1709, N658, N374, N1594);
and AND2 (N1722, N1714, N1337);
nand NAND4 (N1723, N1708, N1644, N609, N373);
xor XOR2 (N1724, N1720, N947);
or OR3 (N1725, N1717, N4, N475);
not NOT1 (N1726, N1721);
nand NAND3 (N1727, N1719, N1719, N738);
xor XOR2 (N1728, N1724, N614);
and AND2 (N1729, N1716, N267);
nor NOR4 (N1730, N1727, N672, N45, N693);
nand NAND3 (N1731, N1725, N1411, N543);
buf BUF1 (N1732, N1723);
or OR3 (N1733, N1732, N590, N39);
or OR3 (N1734, N1731, N843, N640);
nand NAND3 (N1735, N1729, N317, N1323);
xor XOR2 (N1736, N1711, N566);
not NOT1 (N1737, N1726);
nand NAND2 (N1738, N1722, N273);
or OR4 (N1739, N1737, N1680, N920, N280);
buf BUF1 (N1740, N1730);
buf BUF1 (N1741, N1734);
or OR2 (N1742, N1740, N718);
or OR3 (N1743, N1742, N1638, N784);
nor NOR2 (N1744, N1735, N292);
not NOT1 (N1745, N1713);
nand NAND4 (N1746, N1743, N497, N1554, N1209);
buf BUF1 (N1747, N1736);
nor NOR4 (N1748, N1746, N1686, N293, N289);
buf BUF1 (N1749, N1744);
nand NAND3 (N1750, N1745, N407, N439);
nand NAND3 (N1751, N1748, N926, N556);
or OR3 (N1752, N1739, N1234, N1418);
nand NAND3 (N1753, N1750, N1271, N1598);
buf BUF1 (N1754, N1751);
or OR2 (N1755, N1733, N289);
nand NAND3 (N1756, N1741, N21, N1141);
buf BUF1 (N1757, N1712);
xor XOR2 (N1758, N1728, N1025);
and AND4 (N1759, N1754, N1509, N509, N1589);
nand NAND2 (N1760, N1757, N1523);
or OR2 (N1761, N1759, N952);
not NOT1 (N1762, N1758);
buf BUF1 (N1763, N1753);
nand NAND2 (N1764, N1763, N1658);
nand NAND3 (N1765, N1764, N649, N1233);
nor NOR4 (N1766, N1752, N273, N904, N1038);
nor NOR3 (N1767, N1765, N1193, N68);
xor XOR2 (N1768, N1756, N1201);
buf BUF1 (N1769, N1762);
nor NOR2 (N1770, N1755, N1762);
or OR3 (N1771, N1760, N1442, N1190);
nand NAND2 (N1772, N1768, N1259);
xor XOR2 (N1773, N1769, N1326);
or OR4 (N1774, N1738, N746, N1514, N358);
buf BUF1 (N1775, N1771);
xor XOR2 (N1776, N1749, N842);
or OR4 (N1777, N1772, N263, N642, N322);
or OR4 (N1778, N1773, N1631, N1643, N183);
not NOT1 (N1779, N1774);
nor NOR2 (N1780, N1766, N428);
nand NAND2 (N1781, N1767, N1091);
buf BUF1 (N1782, N1780);
nor NOR3 (N1783, N1777, N250, N365);
or OR3 (N1784, N1779, N571, N1448);
buf BUF1 (N1785, N1776);
and AND4 (N1786, N1778, N1087, N89, N364);
xor XOR2 (N1787, N1747, N934);
and AND2 (N1788, N1784, N257);
and AND3 (N1789, N1785, N992, N1218);
nor NOR4 (N1790, N1775, N534, N8, N1482);
nand NAND2 (N1791, N1770, N483);
xor XOR2 (N1792, N1788, N645);
not NOT1 (N1793, N1761);
or OR4 (N1794, N1789, N62, N447, N1373);
xor XOR2 (N1795, N1792, N1404);
nand NAND3 (N1796, N1781, N896, N852);
not NOT1 (N1797, N1782);
and AND3 (N1798, N1786, N107, N1332);
or OR4 (N1799, N1787, N946, N1373, N63);
and AND4 (N1800, N1783, N650, N949, N1542);
xor XOR2 (N1801, N1794, N993);
buf BUF1 (N1802, N1793);
nor NOR3 (N1803, N1800, N1014, N1215);
and AND4 (N1804, N1802, N320, N1491, N169);
nand NAND2 (N1805, N1803, N1463);
buf BUF1 (N1806, N1801);
and AND4 (N1807, N1795, N966, N1777, N752);
nor NOR3 (N1808, N1791, N694, N351);
buf BUF1 (N1809, N1797);
nor NOR4 (N1810, N1790, N1428, N67, N1558);
not NOT1 (N1811, N1799);
not NOT1 (N1812, N1808);
and AND4 (N1813, N1806, N755, N1436, N412);
xor XOR2 (N1814, N1809, N604);
and AND2 (N1815, N1796, N1804);
xor XOR2 (N1816, N1269, N851);
xor XOR2 (N1817, N1810, N1326);
nor NOR4 (N1818, N1807, N1683, N1756, N976);
nor NOR2 (N1819, N1814, N219);
nand NAND3 (N1820, N1812, N1738, N359);
xor XOR2 (N1821, N1819, N665);
and AND3 (N1822, N1817, N1115, N1075);
and AND4 (N1823, N1821, N472, N708, N136);
buf BUF1 (N1824, N1816);
and AND3 (N1825, N1822, N615, N1582);
nand NAND2 (N1826, N1818, N1450);
nand NAND2 (N1827, N1811, N779);
buf BUF1 (N1828, N1815);
and AND3 (N1829, N1824, N989, N788);
nand NAND3 (N1830, N1798, N737, N203);
xor XOR2 (N1831, N1813, N506);
or OR2 (N1832, N1825, N1683);
nand NAND2 (N1833, N1829, N1503);
and AND3 (N1834, N1820, N1454, N228);
not NOT1 (N1835, N1823);
or OR2 (N1836, N1833, N1152);
or OR2 (N1837, N1835, N993);
not NOT1 (N1838, N1832);
or OR4 (N1839, N1805, N754, N505, N27);
nor NOR2 (N1840, N1830, N649);
and AND3 (N1841, N1836, N359, N977);
nor NOR4 (N1842, N1838, N1815, N1745, N668);
and AND4 (N1843, N1840, N134, N1671, N806);
or OR2 (N1844, N1828, N361);
nor NOR3 (N1845, N1831, N1769, N953);
xor XOR2 (N1846, N1834, N1313);
and AND2 (N1847, N1839, N1599);
nor NOR3 (N1848, N1847, N302, N974);
or OR4 (N1849, N1837, N618, N703, N614);
and AND4 (N1850, N1842, N648, N572, N721);
xor XOR2 (N1851, N1845, N1785);
xor XOR2 (N1852, N1846, N1564);
not NOT1 (N1853, N1844);
nor NOR4 (N1854, N1848, N468, N181, N323);
and AND4 (N1855, N1827, N1019, N699, N225);
not NOT1 (N1856, N1849);
buf BUF1 (N1857, N1855);
nand NAND4 (N1858, N1826, N857, N514, N882);
nand NAND4 (N1859, N1854, N1600, N1600, N1025);
or OR3 (N1860, N1850, N884, N1785);
not NOT1 (N1861, N1859);
buf BUF1 (N1862, N1856);
nand NAND4 (N1863, N1843, N620, N620, N1424);
and AND2 (N1864, N1857, N1861);
nand NAND4 (N1865, N822, N1542, N1167, N518);
and AND3 (N1866, N1865, N643, N856);
buf BUF1 (N1867, N1858);
nand NAND4 (N1868, N1841, N886, N331, N206);
buf BUF1 (N1869, N1867);
nor NOR3 (N1870, N1863, N422, N606);
not NOT1 (N1871, N1862);
not NOT1 (N1872, N1852);
nand NAND2 (N1873, N1869, N1612);
nand NAND2 (N1874, N1864, N442);
buf BUF1 (N1875, N1871);
or OR3 (N1876, N1860, N66, N15);
buf BUF1 (N1877, N1876);
and AND3 (N1878, N1870, N520, N950);
nand NAND4 (N1879, N1853, N1085, N103, N589);
nand NAND4 (N1880, N1866, N60, N926, N499);
xor XOR2 (N1881, N1878, N1240);
nor NOR2 (N1882, N1879, N581);
not NOT1 (N1883, N1875);
nand NAND3 (N1884, N1882, N1093, N716);
not NOT1 (N1885, N1851);
xor XOR2 (N1886, N1880, N693);
xor XOR2 (N1887, N1873, N979);
nand NAND2 (N1888, N1881, N167);
or OR2 (N1889, N1885, N687);
not NOT1 (N1890, N1874);
nor NOR4 (N1891, N1868, N531, N1646, N312);
nor NOR4 (N1892, N1877, N1392, N158, N1877);
nand NAND4 (N1893, N1872, N184, N1658, N903);
nand NAND3 (N1894, N1884, N631, N1879);
nor NOR2 (N1895, N1887, N1081);
and AND3 (N1896, N1889, N537, N109);
nor NOR4 (N1897, N1886, N264, N1230, N1736);
xor XOR2 (N1898, N1891, N1169);
or OR4 (N1899, N1897, N478, N1626, N179);
and AND2 (N1900, N1895, N1534);
or OR4 (N1901, N1883, N1516, N1570, N1841);
or OR4 (N1902, N1892, N1468, N945, N380);
and AND2 (N1903, N1900, N88);
xor XOR2 (N1904, N1898, N1884);
buf BUF1 (N1905, N1890);
not NOT1 (N1906, N1904);
nor NOR2 (N1907, N1896, N469);
not NOT1 (N1908, N1893);
and AND3 (N1909, N1894, N1171, N1597);
buf BUF1 (N1910, N1899);
buf BUF1 (N1911, N1909);
nor NOR3 (N1912, N1906, N142, N171);
nand NAND3 (N1913, N1888, N1744, N290);
buf BUF1 (N1914, N1902);
xor XOR2 (N1915, N1908, N89);
nand NAND4 (N1916, N1901, N1827, N155, N1201);
nand NAND4 (N1917, N1912, N441, N1581, N834);
nor NOR3 (N1918, N1914, N609, N1247);
not NOT1 (N1919, N1918);
and AND2 (N1920, N1911, N531);
nand NAND3 (N1921, N1907, N1724, N940);
nor NOR3 (N1922, N1910, N627, N1633);
nor NOR2 (N1923, N1921, N965);
xor XOR2 (N1924, N1916, N1475);
nor NOR3 (N1925, N1905, N1232, N1371);
nor NOR3 (N1926, N1923, N1669, N76);
not NOT1 (N1927, N1917);
nand NAND4 (N1928, N1927, N315, N502, N1842);
xor XOR2 (N1929, N1913, N830);
nand NAND4 (N1930, N1903, N1661, N1653, N156);
nor NOR4 (N1931, N1924, N1302, N533, N1841);
not NOT1 (N1932, N1931);
xor XOR2 (N1933, N1926, N530);
or OR2 (N1934, N1932, N795);
and AND2 (N1935, N1920, N789);
not NOT1 (N1936, N1934);
and AND4 (N1937, N1936, N125, N950, N1053);
and AND3 (N1938, N1933, N881, N1733);
and AND3 (N1939, N1938, N710, N342);
nand NAND4 (N1940, N1915, N1491, N273, N417);
and AND3 (N1941, N1928, N994, N1559);
nand NAND4 (N1942, N1922, N569, N250, N393);
and AND4 (N1943, N1939, N1677, N1516, N1709);
nand NAND3 (N1944, N1941, N1469, N88);
buf BUF1 (N1945, N1942);
and AND4 (N1946, N1944, N1225, N1870, N65);
buf BUF1 (N1947, N1943);
not NOT1 (N1948, N1947);
and AND2 (N1949, N1919, N839);
and AND2 (N1950, N1949, N267);
nor NOR4 (N1951, N1950, N1005, N226, N429);
buf BUF1 (N1952, N1935);
and AND2 (N1953, N1930, N584);
nand NAND3 (N1954, N1948, N1620, N1264);
or OR4 (N1955, N1951, N48, N653, N1171);
not NOT1 (N1956, N1937);
nor NOR2 (N1957, N1955, N1659);
buf BUF1 (N1958, N1945);
nor NOR2 (N1959, N1946, N138);
and AND2 (N1960, N1957, N487);
or OR2 (N1961, N1953, N1471);
not NOT1 (N1962, N1954);
nor NOR4 (N1963, N1956, N1956, N1627, N1760);
or OR3 (N1964, N1925, N1034, N1565);
or OR3 (N1965, N1959, N1769, N293);
and AND3 (N1966, N1958, N1243, N1275);
nor NOR2 (N1967, N1961, N1497);
nor NOR4 (N1968, N1964, N316, N1688, N1667);
not NOT1 (N1969, N1952);
not NOT1 (N1970, N1962);
xor XOR2 (N1971, N1963, N952);
or OR4 (N1972, N1929, N1484, N1797, N1082);
xor XOR2 (N1973, N1960, N210);
xor XOR2 (N1974, N1971, N547);
xor XOR2 (N1975, N1940, N311);
not NOT1 (N1976, N1972);
nand NAND3 (N1977, N1975, N1791, N1656);
or OR2 (N1978, N1966, N267);
xor XOR2 (N1979, N1977, N1474);
and AND4 (N1980, N1969, N1475, N177, N1283);
nor NOR3 (N1981, N1973, N1022, N238);
or OR3 (N1982, N1979, N1343, N472);
or OR4 (N1983, N1968, N396, N181, N245);
xor XOR2 (N1984, N1983, N355);
buf BUF1 (N1985, N1967);
xor XOR2 (N1986, N1976, N1063);
and AND3 (N1987, N1965, N1940, N1802);
xor XOR2 (N1988, N1981, N1849);
or OR4 (N1989, N1985, N1180, N1826, N499);
nand NAND4 (N1990, N1987, N265, N1884, N1810);
nor NOR4 (N1991, N1974, N178, N1773, N231);
not NOT1 (N1992, N1978);
not NOT1 (N1993, N1990);
nor NOR3 (N1994, N1988, N1922, N1113);
xor XOR2 (N1995, N1994, N527);
nor NOR3 (N1996, N1995, N807, N1548);
not NOT1 (N1997, N1986);
nor NOR2 (N1998, N1997, N613);
and AND2 (N1999, N1998, N966);
and AND3 (N2000, N1999, N1441, N1172);
or OR2 (N2001, N1980, N948);
nand NAND3 (N2002, N2001, N1853, N1937);
xor XOR2 (N2003, N1984, N1036);
buf BUF1 (N2004, N2000);
not NOT1 (N2005, N2004);
buf BUF1 (N2006, N2005);
buf BUF1 (N2007, N1996);
not NOT1 (N2008, N1982);
nor NOR3 (N2009, N1993, N1237, N1733);
nor NOR2 (N2010, N1991, N1829);
buf BUF1 (N2011, N1992);
buf BUF1 (N2012, N2002);
nor NOR2 (N2013, N1970, N1747);
nor NOR4 (N2014, N2008, N371, N71, N789);
xor XOR2 (N2015, N2007, N789);
buf BUF1 (N2016, N2012);
and AND3 (N2017, N2010, N759, N413);
buf BUF1 (N2018, N2013);
nand NAND3 (N2019, N2017, N943, N869);
xor XOR2 (N2020, N2011, N1648);
nand NAND3 (N2021, N2018, N1164, N515);
nand NAND3 (N2022, N2021, N1927, N667);
buf BUF1 (N2023, N2019);
and AND4 (N2024, N2022, N1141, N224, N103);
not NOT1 (N2025, N2020);
buf BUF1 (N2026, N2003);
nand NAND4 (N2027, N2015, N1851, N1271, N1562);
and AND2 (N2028, N2014, N164);
or OR3 (N2029, N1989, N1921, N234);
not NOT1 (N2030, N2027);
or OR2 (N2031, N2026, N914);
and AND2 (N2032, N2030, N1846);
or OR4 (N2033, N2006, N833, N520, N2016);
and AND2 (N2034, N104, N337);
nand NAND4 (N2035, N2028, N1709, N645, N809);
buf BUF1 (N2036, N2023);
not NOT1 (N2037, N2025);
buf BUF1 (N2038, N2035);
xor XOR2 (N2039, N2037, N771);
xor XOR2 (N2040, N2036, N1688);
nor NOR4 (N2041, N2032, N694, N818, N1593);
not NOT1 (N2042, N2009);
buf BUF1 (N2043, N2039);
nand NAND2 (N2044, N2041, N2);
buf BUF1 (N2045, N2042);
not NOT1 (N2046, N2034);
not NOT1 (N2047, N2043);
xor XOR2 (N2048, N2044, N1629);
buf BUF1 (N2049, N2040);
buf BUF1 (N2050, N2033);
nand NAND4 (N2051, N2045, N430, N1547, N1691);
and AND2 (N2052, N2024, N1273);
and AND3 (N2053, N2051, N614, N1359);
and AND2 (N2054, N2038, N1881);
buf BUF1 (N2055, N2029);
and AND2 (N2056, N2050, N732);
buf BUF1 (N2057, N2031);
xor XOR2 (N2058, N2056, N923);
and AND2 (N2059, N2048, N1796);
nor NOR4 (N2060, N2046, N541, N968, N1258);
or OR2 (N2061, N2052, N192);
buf BUF1 (N2062, N2057);
or OR4 (N2063, N2054, N1891, N1137, N766);
not NOT1 (N2064, N2060);
and AND4 (N2065, N2055, N526, N1988, N878);
xor XOR2 (N2066, N2063, N956);
not NOT1 (N2067, N2065);
nand NAND4 (N2068, N2067, N890, N1279, N1215);
xor XOR2 (N2069, N2059, N435);
nor NOR2 (N2070, N2068, N533);
nor NOR4 (N2071, N2047, N1940, N649, N1964);
nor NOR2 (N2072, N2062, N585);
or OR2 (N2073, N2066, N701);
nand NAND3 (N2074, N2072, N199, N1437);
and AND2 (N2075, N2064, N875);
and AND4 (N2076, N2071, N1015, N1832, N1406);
nand NAND2 (N2077, N2069, N1312);
and AND4 (N2078, N2061, N1627, N1010, N1068);
and AND4 (N2079, N2070, N1091, N101, N1764);
buf BUF1 (N2080, N2077);
nand NAND3 (N2081, N2049, N1956, N1933);
buf BUF1 (N2082, N2074);
and AND3 (N2083, N2075, N1731, N557);
not NOT1 (N2084, N2082);
buf BUF1 (N2085, N2058);
buf BUF1 (N2086, N2085);
or OR2 (N2087, N2079, N557);
and AND4 (N2088, N2084, N654, N1541, N1090);
and AND3 (N2089, N2087, N746, N213);
and AND4 (N2090, N2078, N2077, N1573, N1414);
nor NOR2 (N2091, N2086, N1306);
nor NOR4 (N2092, N2073, N1301, N1450, N331);
not NOT1 (N2093, N2053);
xor XOR2 (N2094, N2089, N209);
xor XOR2 (N2095, N2083, N481);
not NOT1 (N2096, N2091);
nor NOR2 (N2097, N2090, N1743);
nor NOR3 (N2098, N2095, N2021, N1891);
and AND3 (N2099, N2088, N1638, N980);
and AND3 (N2100, N2096, N1556, N1562);
not NOT1 (N2101, N2093);
not NOT1 (N2102, N2094);
and AND2 (N2103, N2099, N1320);
buf BUF1 (N2104, N2097);
nand NAND3 (N2105, N2092, N1684, N1061);
nor NOR3 (N2106, N2100, N1079, N26);
nand NAND4 (N2107, N2103, N1125, N1256, N1471);
nand NAND4 (N2108, N2105, N1174, N1086, N1833);
and AND3 (N2109, N2080, N264, N1787);
buf BUF1 (N2110, N2081);
not NOT1 (N2111, N2108);
nor NOR4 (N2112, N2076, N505, N236, N1548);
buf BUF1 (N2113, N2111);
xor XOR2 (N2114, N2112, N1691);
buf BUF1 (N2115, N2101);
nor NOR2 (N2116, N2107, N988);
and AND4 (N2117, N2115, N1799, N1977, N336);
nor NOR2 (N2118, N2116, N1283);
and AND3 (N2119, N2117, N1360, N1300);
xor XOR2 (N2120, N2113, N1475);
nor NOR2 (N2121, N2104, N413);
nand NAND4 (N2122, N2118, N1271, N169, N1192);
nor NOR3 (N2123, N2102, N260, N7);
nand NAND2 (N2124, N2120, N441);
or OR2 (N2125, N2109, N2038);
or OR3 (N2126, N2106, N1163, N2021);
buf BUF1 (N2127, N2123);
and AND4 (N2128, N2127, N792, N155, N629);
nand NAND2 (N2129, N2110, N2055);
nand NAND3 (N2130, N2125, N273, N1400);
nor NOR2 (N2131, N2119, N939);
nor NOR2 (N2132, N2129, N637);
nor NOR4 (N2133, N2130, N906, N50, N1273);
and AND4 (N2134, N2131, N856, N641, N163);
buf BUF1 (N2135, N2124);
nor NOR2 (N2136, N2135, N1147);
nand NAND3 (N2137, N2136, N1751, N1051);
nor NOR3 (N2138, N2134, N1306, N1776);
not NOT1 (N2139, N2098);
or OR2 (N2140, N2137, N480);
and AND4 (N2141, N2114, N1232, N1969, N708);
not NOT1 (N2142, N2140);
xor XOR2 (N2143, N2122, N1524);
xor XOR2 (N2144, N2141, N764);
not NOT1 (N2145, N2132);
buf BUF1 (N2146, N2121);
nand NAND4 (N2147, N2145, N1464, N456, N565);
or OR2 (N2148, N2128, N324);
nor NOR2 (N2149, N2138, N306);
and AND3 (N2150, N2148, N798, N210);
and AND3 (N2151, N2149, N1619, N1738);
nand NAND4 (N2152, N2144, N515, N932, N2110);
nor NOR4 (N2153, N2143, N1248, N278, N1251);
buf BUF1 (N2154, N2126);
and AND2 (N2155, N2142, N1313);
xor XOR2 (N2156, N2146, N1604);
or OR3 (N2157, N2152, N1908, N1739);
not NOT1 (N2158, N2156);
buf BUF1 (N2159, N2158);
nand NAND4 (N2160, N2157, N1593, N2157, N182);
nand NAND3 (N2161, N2159, N902, N1033);
nand NAND3 (N2162, N2139, N675, N1947);
or OR4 (N2163, N2155, N1143, N1643, N810);
xor XOR2 (N2164, N2163, N1718);
and AND4 (N2165, N2164, N17, N1827, N800);
nor NOR4 (N2166, N2133, N1426, N95, N1502);
or OR2 (N2167, N2153, N2053);
xor XOR2 (N2168, N2147, N2107);
buf BUF1 (N2169, N2150);
not NOT1 (N2170, N2168);
buf BUF1 (N2171, N2160);
and AND2 (N2172, N2154, N701);
buf BUF1 (N2173, N2171);
and AND4 (N2174, N2167, N270, N601, N1065);
buf BUF1 (N2175, N2173);
xor XOR2 (N2176, N2175, N1530);
or OR2 (N2177, N2174, N556);
nor NOR4 (N2178, N2176, N1816, N2117, N1333);
buf BUF1 (N2179, N2170);
or OR2 (N2180, N2172, N1721);
not NOT1 (N2181, N2151);
and AND2 (N2182, N2161, N333);
not NOT1 (N2183, N2182);
buf BUF1 (N2184, N2183);
or OR2 (N2185, N2178, N941);
xor XOR2 (N2186, N2185, N651);
buf BUF1 (N2187, N2177);
nor NOR4 (N2188, N2187, N522, N190, N26);
xor XOR2 (N2189, N2188, N85);
nor NOR3 (N2190, N2179, N432, N1391);
nand NAND4 (N2191, N2181, N1612, N1264, N1695);
not NOT1 (N2192, N2165);
and AND3 (N2193, N2192, N2148, N671);
and AND4 (N2194, N2189, N372, N1543, N744);
not NOT1 (N2195, N2180);
not NOT1 (N2196, N2169);
xor XOR2 (N2197, N2193, N2154);
or OR3 (N2198, N2166, N1243, N1032);
or OR3 (N2199, N2186, N1220, N508);
nor NOR3 (N2200, N2184, N1777, N1127);
nor NOR4 (N2201, N2198, N2056, N1446, N2037);
or OR4 (N2202, N2197, N1738, N399, N449);
buf BUF1 (N2203, N2202);
nand NAND4 (N2204, N2191, N323, N1344, N1325);
nand NAND3 (N2205, N2204, N1769, N645);
or OR2 (N2206, N2200, N1820);
nand NAND3 (N2207, N2201, N2108, N1385);
nor NOR4 (N2208, N2195, N1811, N2182, N804);
or OR4 (N2209, N2190, N1915, N708, N2097);
or OR4 (N2210, N2207, N1213, N1446, N1139);
nor NOR3 (N2211, N2210, N1910, N1083);
buf BUF1 (N2212, N2205);
xor XOR2 (N2213, N2196, N1752);
nor NOR3 (N2214, N2208, N34, N1723);
xor XOR2 (N2215, N2194, N631);
xor XOR2 (N2216, N2213, N2115);
or OR4 (N2217, N2162, N1940, N1160, N2063);
nor NOR4 (N2218, N2215, N917, N1230, N1236);
or OR2 (N2219, N2209, N1521);
not NOT1 (N2220, N2206);
and AND2 (N2221, N2199, N942);
nor NOR2 (N2222, N2203, N539);
or OR2 (N2223, N2211, N1459);
nand NAND2 (N2224, N2216, N767);
and AND3 (N2225, N2224, N558, N1785);
nand NAND4 (N2226, N2225, N18, N1528, N1598);
not NOT1 (N2227, N2220);
nor NOR4 (N2228, N2221, N256, N1700, N831);
nor NOR3 (N2229, N2223, N1500, N392);
and AND3 (N2230, N2218, N1485, N1245);
xor XOR2 (N2231, N2214, N1918);
and AND4 (N2232, N2217, N1174, N2155, N1434);
buf BUF1 (N2233, N2212);
buf BUF1 (N2234, N2219);
nand NAND2 (N2235, N2234, N303);
and AND4 (N2236, N2226, N854, N1722, N702);
buf BUF1 (N2237, N2222);
or OR3 (N2238, N2235, N1827, N1705);
not NOT1 (N2239, N2233);
buf BUF1 (N2240, N2227);
buf BUF1 (N2241, N2240);
nand NAND2 (N2242, N2236, N472);
buf BUF1 (N2243, N2238);
buf BUF1 (N2244, N2229);
or OR2 (N2245, N2243, N1685);
nor NOR2 (N2246, N2232, N1665);
not NOT1 (N2247, N2246);
buf BUF1 (N2248, N2241);
or OR4 (N2249, N2239, N2191, N103, N1814);
and AND3 (N2250, N2228, N1472, N1736);
or OR3 (N2251, N2245, N2236, N1006);
and AND3 (N2252, N2248, N256, N398);
nand NAND4 (N2253, N2251, N1354, N1938, N2025);
not NOT1 (N2254, N2242);
nor NOR3 (N2255, N2237, N939, N624);
xor XOR2 (N2256, N2252, N1850);
xor XOR2 (N2257, N2244, N1073);
buf BUF1 (N2258, N2253);
or OR2 (N2259, N2249, N1647);
nand NAND4 (N2260, N2255, N789, N828, N811);
nand NAND3 (N2261, N2258, N509, N52);
not NOT1 (N2262, N2259);
not NOT1 (N2263, N2247);
nor NOR4 (N2264, N2230, N1060, N819, N844);
and AND3 (N2265, N2260, N1383, N458);
nand NAND4 (N2266, N2265, N906, N118, N1514);
not NOT1 (N2267, N2256);
or OR4 (N2268, N2263, N1079, N1311, N1491);
nor NOR4 (N2269, N2268, N1809, N1706, N542);
nor NOR4 (N2270, N2250, N43, N606, N1556);
buf BUF1 (N2271, N2267);
not NOT1 (N2272, N2266);
xor XOR2 (N2273, N2270, N600);
buf BUF1 (N2274, N2261);
buf BUF1 (N2275, N2262);
and AND2 (N2276, N2271, N411);
not NOT1 (N2277, N2254);
or OR3 (N2278, N2264, N1480, N491);
nor NOR3 (N2279, N2272, N104, N531);
nand NAND2 (N2280, N2275, N1187);
and AND3 (N2281, N2276, N632, N1353);
nand NAND4 (N2282, N2231, N1175, N207, N895);
or OR2 (N2283, N2257, N1071);
buf BUF1 (N2284, N2280);
xor XOR2 (N2285, N2281, N84);
buf BUF1 (N2286, N2277);
buf BUF1 (N2287, N2278);
buf BUF1 (N2288, N2284);
nand NAND3 (N2289, N2287, N1126, N786);
buf BUF1 (N2290, N2273);
nor NOR3 (N2291, N2290, N270, N1833);
nor NOR3 (N2292, N2269, N317, N1488);
buf BUF1 (N2293, N2289);
nor NOR3 (N2294, N2285, N1609, N239);
or OR3 (N2295, N2293, N1154, N382);
nor NOR3 (N2296, N2292, N223, N1083);
not NOT1 (N2297, N2279);
xor XOR2 (N2298, N2286, N559);
nor NOR2 (N2299, N2295, N1856);
xor XOR2 (N2300, N2291, N439);
nor NOR4 (N2301, N2294, N1997, N1561, N1895);
xor XOR2 (N2302, N2283, N1888);
buf BUF1 (N2303, N2274);
or OR2 (N2304, N2282, N2162);
nand NAND4 (N2305, N2299, N447, N844, N1033);
or OR4 (N2306, N2303, N1833, N397, N1576);
buf BUF1 (N2307, N2306);
buf BUF1 (N2308, N2302);
or OR4 (N2309, N2307, N1652, N37, N1438);
and AND2 (N2310, N2301, N2088);
and AND4 (N2311, N2310, N1965, N1869, N1048);
nor NOR3 (N2312, N2309, N2150, N531);
nand NAND4 (N2313, N2308, N1229, N1665, N378);
and AND4 (N2314, N2312, N1569, N1267, N902);
buf BUF1 (N2315, N2288);
nand NAND3 (N2316, N2313, N776, N630);
nor NOR3 (N2317, N2304, N732, N2109);
xor XOR2 (N2318, N2311, N442);
nand NAND2 (N2319, N2296, N386);
nor NOR3 (N2320, N2316, N1358, N1973);
xor XOR2 (N2321, N2318, N1494);
nor NOR3 (N2322, N2314, N1488, N2031);
and AND3 (N2323, N2300, N1319, N109);
buf BUF1 (N2324, N2315);
or OR4 (N2325, N2319, N491, N989, N157);
xor XOR2 (N2326, N2320, N1126);
nand NAND3 (N2327, N2321, N1169, N1251);
or OR4 (N2328, N2327, N1718, N1055, N687);
nor NOR4 (N2329, N2322, N2106, N873, N793);
and AND3 (N2330, N2317, N1611, N1424);
buf BUF1 (N2331, N2324);
buf BUF1 (N2332, N2329);
not NOT1 (N2333, N2326);
not NOT1 (N2334, N2298);
nand NAND2 (N2335, N2334, N2188);
xor XOR2 (N2336, N2331, N2188);
or OR2 (N2337, N2323, N1947);
or OR4 (N2338, N2297, N1753, N1166, N2021);
nand NAND4 (N2339, N2328, N82, N1522, N2037);
and AND3 (N2340, N2338, N641, N1134);
xor XOR2 (N2341, N2333, N1275);
nand NAND2 (N2342, N2330, N49);
nor NOR2 (N2343, N2340, N1945);
or OR2 (N2344, N2335, N1935);
or OR3 (N2345, N2339, N1106, N708);
nor NOR3 (N2346, N2337, N2115, N410);
not NOT1 (N2347, N2336);
xor XOR2 (N2348, N2305, N1135);
or OR3 (N2349, N2347, N1555, N489);
not NOT1 (N2350, N2345);
not NOT1 (N2351, N2348);
xor XOR2 (N2352, N2344, N918);
and AND4 (N2353, N2343, N1136, N1072, N1393);
xor XOR2 (N2354, N2342, N1886);
buf BUF1 (N2355, N2349);
or OR4 (N2356, N2325, N608, N1576, N931);
nand NAND2 (N2357, N2353, N1479);
nor NOR3 (N2358, N2350, N965, N771);
xor XOR2 (N2359, N2355, N674);
nor NOR4 (N2360, N2357, N1773, N809, N1203);
nor NOR2 (N2361, N2360, N14);
not NOT1 (N2362, N2332);
nand NAND2 (N2363, N2346, N1221);
not NOT1 (N2364, N2358);
nand NAND3 (N2365, N2363, N1839, N278);
and AND2 (N2366, N2351, N1331);
xor XOR2 (N2367, N2362, N301);
nand NAND2 (N2368, N2352, N1308);
buf BUF1 (N2369, N2368);
not NOT1 (N2370, N2364);
xor XOR2 (N2371, N2369, N1653);
or OR4 (N2372, N2370, N295, N559, N218);
nand NAND4 (N2373, N2341, N1411, N85, N109);
nand NAND4 (N2374, N2359, N1260, N69, N1731);
nand NAND4 (N2375, N2372, N1927, N1085, N255);
nand NAND3 (N2376, N2354, N1768, N889);
not NOT1 (N2377, N2373);
buf BUF1 (N2378, N2356);
xor XOR2 (N2379, N2371, N4);
or OR2 (N2380, N2366, N1551);
and AND2 (N2381, N2378, N1917);
or OR3 (N2382, N2367, N1385, N2247);
not NOT1 (N2383, N2381);
or OR2 (N2384, N2361, N2163);
buf BUF1 (N2385, N2374);
nand NAND2 (N2386, N2376, N1466);
not NOT1 (N2387, N2375);
nand NAND2 (N2388, N2386, N1630);
not NOT1 (N2389, N2385);
nor NOR2 (N2390, N2389, N154);
or OR2 (N2391, N2365, N1112);
nor NOR2 (N2392, N2382, N1875);
buf BUF1 (N2393, N2391);
or OR2 (N2394, N2387, N1462);
nand NAND3 (N2395, N2393, N2149, N781);
and AND4 (N2396, N2395, N1529, N2074, N1121);
xor XOR2 (N2397, N2390, N681);
and AND4 (N2398, N2388, N781, N957, N2183);
and AND4 (N2399, N2396, N1966, N996, N319);
buf BUF1 (N2400, N2392);
nor NOR4 (N2401, N2399, N368, N2032, N60);
or OR3 (N2402, N2384, N1743, N2372);
nand NAND4 (N2403, N2377, N2101, N2240, N2092);
buf BUF1 (N2404, N2379);
or OR2 (N2405, N2380, N613);
nand NAND4 (N2406, N2405, N1581, N140, N490);
and AND3 (N2407, N2397, N132, N2311);
nor NOR2 (N2408, N2401, N926);
or OR4 (N2409, N2404, N694, N422, N1560);
xor XOR2 (N2410, N2408, N337);
not NOT1 (N2411, N2406);
xor XOR2 (N2412, N2400, N312);
nand NAND4 (N2413, N2398, N69, N618, N584);
and AND4 (N2414, N2411, N1153, N1612, N1037);
nand NAND2 (N2415, N2413, N1787);
and AND3 (N2416, N2410, N1542, N15);
nand NAND2 (N2417, N2394, N585);
or OR2 (N2418, N2415, N1627);
nand NAND4 (N2419, N2417, N1594, N1772, N970);
nand NAND2 (N2420, N2383, N1412);
and AND2 (N2421, N2419, N291);
and AND4 (N2422, N2403, N444, N479, N123);
xor XOR2 (N2423, N2421, N323);
and AND2 (N2424, N2416, N1083);
buf BUF1 (N2425, N2420);
not NOT1 (N2426, N2414);
nand NAND2 (N2427, N2409, N720);
xor XOR2 (N2428, N2427, N516);
xor XOR2 (N2429, N2418, N625);
nand NAND3 (N2430, N2424, N853, N1946);
buf BUF1 (N2431, N2407);
or OR3 (N2432, N2429, N1615, N2369);
nor NOR2 (N2433, N2426, N205);
buf BUF1 (N2434, N2433);
nand NAND4 (N2435, N2422, N4, N1805, N127);
xor XOR2 (N2436, N2430, N1467);
not NOT1 (N2437, N2402);
xor XOR2 (N2438, N2434, N458);
and AND4 (N2439, N2436, N908, N1974, N1332);
not NOT1 (N2440, N2432);
not NOT1 (N2441, N2412);
and AND4 (N2442, N2437, N1303, N66, N1590);
xor XOR2 (N2443, N2435, N2020);
xor XOR2 (N2444, N2442, N1176);
nand NAND4 (N2445, N2439, N566, N2289, N2314);
nor NOR2 (N2446, N2425, N1953);
buf BUF1 (N2447, N2446);
xor XOR2 (N2448, N2438, N1873);
buf BUF1 (N2449, N2443);
and AND4 (N2450, N2449, N595, N1906, N219);
not NOT1 (N2451, N2431);
not NOT1 (N2452, N2423);
or OR4 (N2453, N2452, N907, N904, N1201);
not NOT1 (N2454, N2445);
or OR4 (N2455, N2453, N112, N1668, N1406);
buf BUF1 (N2456, N2440);
buf BUF1 (N2457, N2447);
xor XOR2 (N2458, N2454, N223);
nor NOR3 (N2459, N2457, N2021, N1452);
xor XOR2 (N2460, N2441, N2397);
and AND2 (N2461, N2459, N518);
or OR2 (N2462, N2444, N572);
nand NAND4 (N2463, N2428, N1189, N963, N1551);
or OR4 (N2464, N2451, N1850, N556, N1210);
buf BUF1 (N2465, N2450);
nand NAND3 (N2466, N2465, N1080, N994);
or OR3 (N2467, N2461, N1069, N988);
xor XOR2 (N2468, N2460, N599);
buf BUF1 (N2469, N2458);
not NOT1 (N2470, N2462);
xor XOR2 (N2471, N2466, N2346);
not NOT1 (N2472, N2468);
nor NOR2 (N2473, N2470, N1992);
or OR4 (N2474, N2455, N931, N484, N2001);
buf BUF1 (N2475, N2456);
nor NOR4 (N2476, N2473, N400, N1359, N1725);
and AND2 (N2477, N2475, N238);
xor XOR2 (N2478, N2469, N1627);
and AND2 (N2479, N2477, N1630);
buf BUF1 (N2480, N2472);
nand NAND4 (N2481, N2479, N1131, N910, N1267);
not NOT1 (N2482, N2471);
buf BUF1 (N2483, N2464);
or OR3 (N2484, N2476, N1322, N1644);
nand NAND2 (N2485, N2448, N233);
xor XOR2 (N2486, N2478, N1952);
and AND3 (N2487, N2480, N53, N249);
buf BUF1 (N2488, N2474);
or OR2 (N2489, N2487, N2214);
and AND2 (N2490, N2488, N2091);
or OR4 (N2491, N2489, N948, N1958, N305);
xor XOR2 (N2492, N2467, N596);
nand NAND3 (N2493, N2463, N526, N358);
buf BUF1 (N2494, N2486);
nor NOR3 (N2495, N2483, N1480, N564);
buf BUF1 (N2496, N2485);
nor NOR2 (N2497, N2496, N2036);
xor XOR2 (N2498, N2495, N1250);
buf BUF1 (N2499, N2493);
not NOT1 (N2500, N2481);
buf BUF1 (N2501, N2491);
and AND2 (N2502, N2497, N510);
buf BUF1 (N2503, N2499);
nand NAND3 (N2504, N2484, N1944, N2020);
buf BUF1 (N2505, N2494);
and AND4 (N2506, N2482, N1223, N907, N1918);
and AND3 (N2507, N2502, N1816, N1180);
nor NOR2 (N2508, N2505, N1785);
and AND3 (N2509, N2506, N2386, N2125);
buf BUF1 (N2510, N2498);
nor NOR4 (N2511, N2510, N1349, N2061, N2403);
nand NAND4 (N2512, N2503, N872, N1062, N651);
not NOT1 (N2513, N2490);
nor NOR3 (N2514, N2507, N719, N1459);
xor XOR2 (N2515, N2508, N2480);
nor NOR2 (N2516, N2512, N2272);
nand NAND2 (N2517, N2516, N1292);
nand NAND2 (N2518, N2513, N317);
nor NOR3 (N2519, N2517, N1295, N735);
xor XOR2 (N2520, N2509, N1634);
buf BUF1 (N2521, N2501);
nand NAND2 (N2522, N2511, N364);
nand NAND2 (N2523, N2514, N1964);
nor NOR4 (N2524, N2500, N29, N1017, N1501);
and AND2 (N2525, N2523, N902);
not NOT1 (N2526, N2524);
xor XOR2 (N2527, N2515, N784);
nor NOR2 (N2528, N2520, N1620);
xor XOR2 (N2529, N2492, N1245);
nand NAND2 (N2530, N2519, N1348);
buf BUF1 (N2531, N2530);
and AND3 (N2532, N2518, N159, N1657);
nand NAND4 (N2533, N2522, N1082, N151, N1530);
not NOT1 (N2534, N2521);
not NOT1 (N2535, N2531);
nor NOR3 (N2536, N2527, N1533, N2108);
nand NAND4 (N2537, N2526, N2522, N1601, N2087);
buf BUF1 (N2538, N2533);
nand NAND4 (N2539, N2504, N1189, N2268, N929);
and AND4 (N2540, N2532, N78, N328, N1985);
not NOT1 (N2541, N2536);
xor XOR2 (N2542, N2529, N1392);
not NOT1 (N2543, N2541);
or OR4 (N2544, N2525, N579, N740, N2296);
and AND3 (N2545, N2539, N1889, N1738);
nor NOR2 (N2546, N2540, N1334);
or OR3 (N2547, N2528, N440, N528);
nand NAND3 (N2548, N2534, N333, N1455);
xor XOR2 (N2549, N2535, N812);
xor XOR2 (N2550, N2543, N2297);
buf BUF1 (N2551, N2548);
buf BUF1 (N2552, N2545);
nand NAND3 (N2553, N2542, N1520, N759);
not NOT1 (N2554, N2550);
not NOT1 (N2555, N2538);
nor NOR3 (N2556, N2553, N1949, N949);
and AND2 (N2557, N2552, N648);
and AND2 (N2558, N2556, N1669);
or OR4 (N2559, N2547, N640, N2120, N1606);
buf BUF1 (N2560, N2546);
and AND3 (N2561, N2549, N1699, N1365);
nor NOR2 (N2562, N2537, N1161);
xor XOR2 (N2563, N2544, N1516);
and AND3 (N2564, N2559, N1025, N710);
or OR3 (N2565, N2564, N1794, N154);
and AND4 (N2566, N2560, N2163, N9, N88);
nand NAND2 (N2567, N2555, N1043);
nor NOR2 (N2568, N2561, N183);
buf BUF1 (N2569, N2567);
not NOT1 (N2570, N2565);
nor NOR2 (N2571, N2563, N2269);
nand NAND2 (N2572, N2570, N2367);
and AND2 (N2573, N2558, N289);
or OR2 (N2574, N2562, N2334);
and AND4 (N2575, N2571, N907, N1308, N1835);
and AND2 (N2576, N2551, N367);
and AND2 (N2577, N2574, N1270);
buf BUF1 (N2578, N2576);
buf BUF1 (N2579, N2569);
nor NOR2 (N2580, N2578, N1859);
nor NOR3 (N2581, N2579, N1004, N1488);
buf BUF1 (N2582, N2566);
not NOT1 (N2583, N2554);
not NOT1 (N2584, N2581);
xor XOR2 (N2585, N2584, N1577);
nand NAND3 (N2586, N2557, N2216, N2572);
nand NAND4 (N2587, N451, N966, N598, N1895);
not NOT1 (N2588, N2586);
or OR4 (N2589, N2585, N145, N1935, N1746);
xor XOR2 (N2590, N2582, N2020);
and AND3 (N2591, N2573, N763, N127);
nor NOR2 (N2592, N2587, N576);
or OR4 (N2593, N2588, N2467, N126, N443);
not NOT1 (N2594, N2580);
buf BUF1 (N2595, N2592);
xor XOR2 (N2596, N2583, N2366);
and AND3 (N2597, N2595, N187, N665);
nor NOR2 (N2598, N2594, N1153);
or OR3 (N2599, N2591, N1189, N1493);
xor XOR2 (N2600, N2596, N2394);
buf BUF1 (N2601, N2599);
buf BUF1 (N2602, N2593);
nand NAND3 (N2603, N2589, N2173, N2279);
nor NOR3 (N2604, N2602, N936, N1672);
and AND2 (N2605, N2590, N2292);
nor NOR4 (N2606, N2604, N2471, N2447, N1845);
buf BUF1 (N2607, N2600);
nor NOR2 (N2608, N2597, N2507);
xor XOR2 (N2609, N2568, N2543);
xor XOR2 (N2610, N2603, N527);
nand NAND4 (N2611, N2577, N2329, N1797, N561);
nand NAND4 (N2612, N2575, N2528, N1810, N1685);
nor NOR3 (N2613, N2609, N1357, N58);
not NOT1 (N2614, N2608);
or OR2 (N2615, N2605, N890);
xor XOR2 (N2616, N2607, N1972);
not NOT1 (N2617, N2598);
or OR3 (N2618, N2615, N2050, N125);
xor XOR2 (N2619, N2618, N215);
xor XOR2 (N2620, N2619, N748);
not NOT1 (N2621, N2612);
and AND3 (N2622, N2601, N882, N1319);
buf BUF1 (N2623, N2616);
not NOT1 (N2624, N2620);
or OR2 (N2625, N2624, N232);
buf BUF1 (N2626, N2617);
xor XOR2 (N2627, N2622, N1843);
nor NOR3 (N2628, N2611, N2624, N739);
xor XOR2 (N2629, N2614, N1056);
xor XOR2 (N2630, N2613, N1694);
buf BUF1 (N2631, N2623);
xor XOR2 (N2632, N2629, N1842);
and AND2 (N2633, N2632, N2322);
xor XOR2 (N2634, N2606, N604);
and AND4 (N2635, N2626, N1170, N305, N2075);
or OR2 (N2636, N2635, N1094);
and AND3 (N2637, N2628, N2195, N304);
nand NAND4 (N2638, N2627, N2561, N760, N1209);
not NOT1 (N2639, N2638);
nor NOR4 (N2640, N2639, N454, N1932, N309);
not NOT1 (N2641, N2610);
buf BUF1 (N2642, N2636);
and AND4 (N2643, N2625, N1487, N696, N1334);
xor XOR2 (N2644, N2641, N489);
nand NAND4 (N2645, N2633, N269, N2163, N2);
xor XOR2 (N2646, N2637, N1255);
nand NAND2 (N2647, N2644, N1643);
not NOT1 (N2648, N2634);
xor XOR2 (N2649, N2621, N472);
and AND2 (N2650, N2630, N1170);
not NOT1 (N2651, N2650);
or OR3 (N2652, N2646, N1056, N1615);
nand NAND4 (N2653, N2640, N1944, N872, N2305);
xor XOR2 (N2654, N2651, N419);
not NOT1 (N2655, N2631);
nor NOR3 (N2656, N2652, N1374, N628);
buf BUF1 (N2657, N2642);
nor NOR4 (N2658, N2655, N646, N698, N238);
buf BUF1 (N2659, N2649);
buf BUF1 (N2660, N2654);
nor NOR4 (N2661, N2657, N1391, N120, N1862);
not NOT1 (N2662, N2653);
buf BUF1 (N2663, N2662);
buf BUF1 (N2664, N2647);
and AND4 (N2665, N2648, N442, N1881, N23);
buf BUF1 (N2666, N2658);
buf BUF1 (N2667, N2664);
buf BUF1 (N2668, N2659);
nand NAND2 (N2669, N2656, N1170);
nand NAND3 (N2670, N2665, N2370, N202);
nor NOR2 (N2671, N2670, N2040);
not NOT1 (N2672, N2643);
xor XOR2 (N2673, N2669, N2457);
xor XOR2 (N2674, N2666, N917);
not NOT1 (N2675, N2674);
or OR4 (N2676, N2673, N842, N982, N1139);
nor NOR4 (N2677, N2676, N689, N2271, N1265);
and AND2 (N2678, N2667, N1173);
nand NAND3 (N2679, N2645, N461, N1848);
buf BUF1 (N2680, N2679);
xor XOR2 (N2681, N2660, N2458);
xor XOR2 (N2682, N2671, N1100);
xor XOR2 (N2683, N2668, N612);
buf BUF1 (N2684, N2683);
xor XOR2 (N2685, N2663, N1136);
nand NAND2 (N2686, N2680, N1564);
nand NAND4 (N2687, N2681, N2109, N1192, N2237);
xor XOR2 (N2688, N2677, N520);
or OR4 (N2689, N2687, N2582, N55, N131);
xor XOR2 (N2690, N2675, N207);
nor NOR2 (N2691, N2678, N403);
nor NOR3 (N2692, N2691, N1834, N295);
xor XOR2 (N2693, N2661, N38);
nand NAND2 (N2694, N2686, N1225);
xor XOR2 (N2695, N2672, N1262);
buf BUF1 (N2696, N2684);
buf BUF1 (N2697, N2694);
or OR4 (N2698, N2690, N2695, N1112, N805);
or OR3 (N2699, N1119, N234, N2246);
buf BUF1 (N2700, N2693);
not NOT1 (N2701, N2688);
nor NOR3 (N2702, N2697, N1146, N2169);
not NOT1 (N2703, N2682);
not NOT1 (N2704, N2700);
or OR3 (N2705, N2703, N2124, N1430);
or OR2 (N2706, N2692, N178);
not NOT1 (N2707, N2689);
nor NOR2 (N2708, N2707, N1036);
xor XOR2 (N2709, N2696, N360);
nor NOR4 (N2710, N2701, N56, N2600, N1708);
buf BUF1 (N2711, N2705);
not NOT1 (N2712, N2710);
nor NOR4 (N2713, N2702, N1290, N2662, N784);
xor XOR2 (N2714, N2685, N1126);
or OR4 (N2715, N2709, N2426, N2068, N1801);
and AND4 (N2716, N2711, N1892, N154, N1212);
buf BUF1 (N2717, N2714);
and AND4 (N2718, N2699, N379, N1776, N723);
and AND3 (N2719, N2712, N1822, N2034);
nor NOR2 (N2720, N2719, N1992);
xor XOR2 (N2721, N2720, N980);
or OR2 (N2722, N2718, N1453);
nor NOR2 (N2723, N2698, N753);
buf BUF1 (N2724, N2716);
and AND3 (N2725, N2717, N2680, N1683);
xor XOR2 (N2726, N2724, N1141);
buf BUF1 (N2727, N2721);
xor XOR2 (N2728, N2713, N1900);
nor NOR4 (N2729, N2726, N2232, N1186, N270);
or OR4 (N2730, N2723, N807, N925, N302);
not NOT1 (N2731, N2706);
and AND4 (N2732, N2731, N9, N193, N393);
nor NOR3 (N2733, N2715, N1178, N742);
buf BUF1 (N2734, N2728);
and AND2 (N2735, N2733, N1226);
or OR3 (N2736, N2732, N2017, N2040);
and AND4 (N2737, N2722, N1970, N976, N1227);
not NOT1 (N2738, N2704);
nand NAND3 (N2739, N2736, N91, N2326);
or OR2 (N2740, N2730, N2632);
and AND3 (N2741, N2727, N311, N2154);
nor NOR4 (N2742, N2741, N1057, N2129, N1742);
nand NAND4 (N2743, N2735, N106, N1195, N2449);
or OR2 (N2744, N2725, N2703);
not NOT1 (N2745, N2740);
or OR4 (N2746, N2739, N623, N1797, N1983);
not NOT1 (N2747, N2743);
buf BUF1 (N2748, N2742);
nor NOR4 (N2749, N2747, N110, N2183, N2110);
or OR2 (N2750, N2729, N246);
buf BUF1 (N2751, N2750);
xor XOR2 (N2752, N2734, N1261);
nand NAND4 (N2753, N2751, N1840, N1528, N1918);
or OR3 (N2754, N2708, N1552, N2071);
not NOT1 (N2755, N2744);
or OR3 (N2756, N2752, N302, N1626);
nand NAND4 (N2757, N2748, N416, N676, N2423);
buf BUF1 (N2758, N2746);
not NOT1 (N2759, N2749);
or OR3 (N2760, N2737, N52, N2290);
nor NOR2 (N2761, N2754, N911);
and AND3 (N2762, N2758, N2596, N853);
not NOT1 (N2763, N2760);
or OR3 (N2764, N2755, N1624, N1397);
buf BUF1 (N2765, N2759);
buf BUF1 (N2766, N2763);
xor XOR2 (N2767, N2765, N2672);
nor NOR4 (N2768, N2766, N757, N1540, N2027);
nor NOR2 (N2769, N2767, N59);
buf BUF1 (N2770, N2756);
not NOT1 (N2771, N2738);
nand NAND3 (N2772, N2771, N1173, N2298);
and AND3 (N2773, N2770, N1700, N1132);
not NOT1 (N2774, N2769);
xor XOR2 (N2775, N2762, N1281);
nor NOR2 (N2776, N2757, N509);
buf BUF1 (N2777, N2761);
buf BUF1 (N2778, N2775);
and AND2 (N2779, N2745, N1031);
nor NOR2 (N2780, N2773, N161);
not NOT1 (N2781, N2753);
or OR4 (N2782, N2778, N2348, N1883, N2687);
nor NOR3 (N2783, N2777, N315, N1325);
xor XOR2 (N2784, N2783, N1216);
and AND2 (N2785, N2781, N1573);
and AND2 (N2786, N2774, N146);
nor NOR4 (N2787, N2776, N366, N32, N1491);
not NOT1 (N2788, N2786);
xor XOR2 (N2789, N2788, N238);
xor XOR2 (N2790, N2785, N1754);
and AND2 (N2791, N2780, N1600);
not NOT1 (N2792, N2791);
buf BUF1 (N2793, N2772);
and AND3 (N2794, N2792, N1237, N430);
xor XOR2 (N2795, N2787, N752);
buf BUF1 (N2796, N2789);
buf BUF1 (N2797, N2794);
not NOT1 (N2798, N2768);
and AND4 (N2799, N2797, N1457, N707, N524);
xor XOR2 (N2800, N2793, N1247);
or OR2 (N2801, N2790, N2000);
buf BUF1 (N2802, N2796);
and AND2 (N2803, N2784, N2130);
or OR3 (N2804, N2764, N2676, N1030);
nand NAND4 (N2805, N2782, N2563, N1792, N606);
not NOT1 (N2806, N2795);
xor XOR2 (N2807, N2779, N2598);
nand NAND4 (N2808, N2804, N617, N1423, N1368);
nand NAND2 (N2809, N2806, N560);
not NOT1 (N2810, N2807);
or OR3 (N2811, N2809, N600, N535);
nand NAND3 (N2812, N2800, N2523, N1112);
buf BUF1 (N2813, N2808);
nor NOR3 (N2814, N2803, N2164, N588);
xor XOR2 (N2815, N2802, N135);
and AND3 (N2816, N2801, N737, N1848);
nand NAND3 (N2817, N2813, N291, N691);
nand NAND4 (N2818, N2814, N6, N494, N743);
or OR4 (N2819, N2811, N931, N2675, N1036);
xor XOR2 (N2820, N2805, N907);
buf BUF1 (N2821, N2815);
nand NAND3 (N2822, N2799, N2046, N2383);
and AND4 (N2823, N2821, N2712, N159, N2350);
xor XOR2 (N2824, N2819, N1512);
nand NAND3 (N2825, N2818, N1871, N357);
buf BUF1 (N2826, N2820);
buf BUF1 (N2827, N2817);
nor NOR2 (N2828, N2810, N2668);
buf BUF1 (N2829, N2825);
and AND4 (N2830, N2826, N2466, N1655, N2278);
nand NAND3 (N2831, N2823, N1470, N2325);
and AND3 (N2832, N2822, N1766, N1525);
not NOT1 (N2833, N2824);
buf BUF1 (N2834, N2833);
not NOT1 (N2835, N2830);
xor XOR2 (N2836, N2834, N2305);
and AND4 (N2837, N2828, N2147, N893, N246);
buf BUF1 (N2838, N2829);
nor NOR3 (N2839, N2798, N2591, N2584);
nor NOR4 (N2840, N2812, N1874, N2761, N1649);
and AND4 (N2841, N2838, N670, N1283, N1050);
buf BUF1 (N2842, N2837);
nand NAND2 (N2843, N2816, N1610);
or OR4 (N2844, N2836, N225, N1671, N612);
nand NAND4 (N2845, N2843, N2631, N337, N195);
nand NAND4 (N2846, N2841, N501, N2121, N441);
and AND3 (N2847, N2842, N1317, N1657);
and AND2 (N2848, N2846, N832);
nor NOR2 (N2849, N2840, N1942);
and AND2 (N2850, N2832, N1223);
not NOT1 (N2851, N2849);
or OR2 (N2852, N2848, N1430);
nand NAND3 (N2853, N2850, N1045, N1671);
nand NAND4 (N2854, N2831, N1793, N501, N541);
or OR2 (N2855, N2847, N1813);
nand NAND3 (N2856, N2851, N1969, N410);
not NOT1 (N2857, N2853);
nand NAND3 (N2858, N2839, N286, N2670);
nand NAND2 (N2859, N2854, N849);
nand NAND2 (N2860, N2855, N1262);
nor NOR3 (N2861, N2857, N1108, N778);
buf BUF1 (N2862, N2835);
and AND4 (N2863, N2860, N2300, N2073, N903);
not NOT1 (N2864, N2827);
nand NAND4 (N2865, N2858, N511, N305, N843);
buf BUF1 (N2866, N2845);
nor NOR4 (N2867, N2859, N1240, N2514, N1101);
xor XOR2 (N2868, N2865, N832);
not NOT1 (N2869, N2856);
nand NAND2 (N2870, N2861, N760);
and AND4 (N2871, N2844, N1556, N450, N1087);
or OR3 (N2872, N2871, N193, N554);
not NOT1 (N2873, N2872);
and AND4 (N2874, N2867, N1011, N267, N1228);
buf BUF1 (N2875, N2864);
nand NAND2 (N2876, N2873, N2164);
not NOT1 (N2877, N2852);
and AND2 (N2878, N2876, N2046);
xor XOR2 (N2879, N2866, N2828);
not NOT1 (N2880, N2868);
xor XOR2 (N2881, N2870, N2076);
not NOT1 (N2882, N2878);
xor XOR2 (N2883, N2877, N1942);
not NOT1 (N2884, N2882);
xor XOR2 (N2885, N2880, N811);
nor NOR2 (N2886, N2883, N2159);
and AND2 (N2887, N2874, N2441);
not NOT1 (N2888, N2881);
buf BUF1 (N2889, N2863);
nand NAND2 (N2890, N2889, N1575);
buf BUF1 (N2891, N2862);
not NOT1 (N2892, N2891);
buf BUF1 (N2893, N2887);
buf BUF1 (N2894, N2875);
xor XOR2 (N2895, N2888, N1599);
buf BUF1 (N2896, N2884);
nand NAND4 (N2897, N2896, N1420, N1498, N2028);
buf BUF1 (N2898, N2892);
buf BUF1 (N2899, N2885);
not NOT1 (N2900, N2886);
or OR3 (N2901, N2893, N1622, N1003);
not NOT1 (N2902, N2901);
nor NOR4 (N2903, N2898, N2620, N2233, N2082);
or OR4 (N2904, N2897, N1793, N1872, N2248);
xor XOR2 (N2905, N2899, N1375);
xor XOR2 (N2906, N2895, N531);
nand NAND2 (N2907, N2905, N2342);
xor XOR2 (N2908, N2902, N434);
not NOT1 (N2909, N2879);
and AND2 (N2910, N2909, N1268);
nor NOR4 (N2911, N2904, N90, N2713, N1345);
xor XOR2 (N2912, N2911, N1957);
or OR4 (N2913, N2910, N1129, N553, N940);
xor XOR2 (N2914, N2906, N2404);
nor NOR3 (N2915, N2900, N169, N43);
nand NAND4 (N2916, N2914, N751, N709, N454);
nand NAND4 (N2917, N2907, N2590, N1947, N983);
and AND2 (N2918, N2917, N2455);
or OR2 (N2919, N2912, N2218);
xor XOR2 (N2920, N2908, N2840);
xor XOR2 (N2921, N2894, N973);
nand NAND2 (N2922, N2916, N293);
nand NAND2 (N2923, N2903, N1508);
nor NOR3 (N2924, N2918, N1895, N396);
nor NOR4 (N2925, N2922, N723, N1041, N1739);
xor XOR2 (N2926, N2869, N765);
buf BUF1 (N2927, N2921);
buf BUF1 (N2928, N2925);
xor XOR2 (N2929, N2913, N82);
nand NAND3 (N2930, N2928, N1126, N2693);
xor XOR2 (N2931, N2923, N285);
not NOT1 (N2932, N2924);
buf BUF1 (N2933, N2890);
buf BUF1 (N2934, N2926);
buf BUF1 (N2935, N2929);
xor XOR2 (N2936, N2935, N2439);
and AND3 (N2937, N2919, N900, N232);
xor XOR2 (N2938, N2934, N678);
and AND2 (N2939, N2927, N1536);
not NOT1 (N2940, N2920);
or OR2 (N2941, N2939, N2566);
xor XOR2 (N2942, N2932, N2628);
and AND4 (N2943, N2936, N2280, N1866, N329);
and AND2 (N2944, N2930, N622);
nor NOR3 (N2945, N2937, N547, N2580);
and AND4 (N2946, N2944, N2393, N1646, N1658);
not NOT1 (N2947, N2933);
xor XOR2 (N2948, N2946, N2915);
nor NOR3 (N2949, N2055, N1599, N125);
nor NOR3 (N2950, N2942, N2200, N2020);
xor XOR2 (N2951, N2931, N630);
xor XOR2 (N2952, N2947, N2728);
xor XOR2 (N2953, N2940, N1323);
or OR3 (N2954, N2943, N183, N1826);
or OR2 (N2955, N2938, N1492);
or OR2 (N2956, N2953, N2418);
nand NAND4 (N2957, N2949, N2719, N23, N558);
not NOT1 (N2958, N2951);
or OR2 (N2959, N2954, N923);
nand NAND2 (N2960, N2948, N422);
nand NAND4 (N2961, N2958, N1375, N2023, N1462);
or OR2 (N2962, N2952, N2533);
and AND4 (N2963, N2941, N675, N1460, N1086);
xor XOR2 (N2964, N2957, N2871);
nand NAND2 (N2965, N2960, N1857);
nor NOR4 (N2966, N2955, N873, N1268, N730);
and AND2 (N2967, N2964, N2940);
nand NAND3 (N2968, N2950, N2890, N2306);
buf BUF1 (N2969, N2961);
buf BUF1 (N2970, N2965);
xor XOR2 (N2971, N2962, N2903);
xor XOR2 (N2972, N2970, N1960);
xor XOR2 (N2973, N2959, N133);
not NOT1 (N2974, N2967);
xor XOR2 (N2975, N2945, N1393);
and AND2 (N2976, N2956, N1079);
and AND4 (N2977, N2972, N563, N423, N440);
nand NAND4 (N2978, N2971, N216, N1661, N1894);
xor XOR2 (N2979, N2963, N369);
buf BUF1 (N2980, N2968);
nand NAND3 (N2981, N2969, N2265, N2374);
buf BUF1 (N2982, N2977);
nor NOR4 (N2983, N2973, N1690, N818, N582);
not NOT1 (N2984, N2980);
xor XOR2 (N2985, N2983, N1565);
buf BUF1 (N2986, N2974);
or OR4 (N2987, N2982, N600, N2583, N1803);
xor XOR2 (N2988, N2976, N866);
or OR4 (N2989, N2978, N2214, N2760, N70);
xor XOR2 (N2990, N2966, N308);
xor XOR2 (N2991, N2985, N411);
xor XOR2 (N2992, N2981, N1250);
or OR3 (N2993, N2990, N1514, N2935);
not NOT1 (N2994, N2992);
or OR4 (N2995, N2991, N1898, N2374, N506);
and AND2 (N2996, N2986, N1809);
and AND4 (N2997, N2996, N686, N76, N2307);
nand NAND2 (N2998, N2995, N1937);
xor XOR2 (N2999, N2997, N2373);
nor NOR2 (N3000, N2993, N130);
not NOT1 (N3001, N2989);
not NOT1 (N3002, N3001);
not NOT1 (N3003, N3002);
nor NOR3 (N3004, N3003, N2331, N2903);
and AND4 (N3005, N2979, N1674, N1291, N1359);
and AND4 (N3006, N2987, N2070, N2610, N1539);
or OR3 (N3007, N2975, N1629, N237);
nand NAND2 (N3008, N3006, N2890);
or OR2 (N3009, N2984, N1090);
xor XOR2 (N3010, N2988, N193);
buf BUF1 (N3011, N3007);
xor XOR2 (N3012, N3005, N1424);
not NOT1 (N3013, N3004);
xor XOR2 (N3014, N3000, N156);
not NOT1 (N3015, N3014);
nor NOR4 (N3016, N3010, N2062, N2967, N1388);
xor XOR2 (N3017, N3016, N1871);
nand NAND3 (N3018, N3012, N2751, N1391);
not NOT1 (N3019, N2998);
nor NOR2 (N3020, N3009, N2593);
or OR4 (N3021, N3011, N1606, N1808, N1653);
and AND2 (N3022, N3021, N2120);
or OR3 (N3023, N3013, N1407, N2262);
nand NAND2 (N3024, N3015, N2393);
nor NOR2 (N3025, N3008, N1220);
nand NAND3 (N3026, N3019, N908, N567);
xor XOR2 (N3027, N3017, N1589);
not NOT1 (N3028, N3027);
not NOT1 (N3029, N3026);
buf BUF1 (N3030, N3029);
not NOT1 (N3031, N3030);
nand NAND4 (N3032, N3023, N1937, N2551, N1408);
buf BUF1 (N3033, N2999);
or OR2 (N3034, N3032, N1979);
nor NOR2 (N3035, N3020, N800);
not NOT1 (N3036, N3034);
xor XOR2 (N3037, N3022, N1962);
nand NAND4 (N3038, N3033, N1616, N1112, N892);
nand NAND2 (N3039, N3025, N1877);
nand NAND4 (N3040, N3024, N1183, N1403, N2949);
or OR3 (N3041, N3036, N569, N436);
not NOT1 (N3042, N3041);
xor XOR2 (N3043, N3038, N124);
buf BUF1 (N3044, N3042);
xor XOR2 (N3045, N3037, N1626);
or OR2 (N3046, N3028, N1333);
or OR2 (N3047, N3046, N1633);
and AND3 (N3048, N3018, N427, N1275);
nand NAND2 (N3049, N3044, N1132);
and AND3 (N3050, N3049, N1999, N73);
nand NAND4 (N3051, N2994, N609, N603, N2753);
buf BUF1 (N3052, N3035);
and AND3 (N3053, N3047, N1697, N936);
and AND4 (N3054, N3031, N2107, N2938, N2126);
xor XOR2 (N3055, N3040, N1971);
nand NAND4 (N3056, N3050, N2334, N2836, N127);
and AND4 (N3057, N3053, N2890, N1106, N2839);
and AND4 (N3058, N3057, N2974, N1112, N189);
not NOT1 (N3059, N3054);
and AND4 (N3060, N3059, N1340, N371, N2803);
xor XOR2 (N3061, N3055, N1633);
not NOT1 (N3062, N3043);
not NOT1 (N3063, N3061);
not NOT1 (N3064, N3052);
or OR3 (N3065, N3056, N910, N1886);
nor NOR2 (N3066, N3058, N2828);
not NOT1 (N3067, N3064);
and AND4 (N3068, N3065, N3041, N3059, N711);
not NOT1 (N3069, N3067);
not NOT1 (N3070, N3039);
nand NAND4 (N3071, N3062, N2692, N1383, N2631);
xor XOR2 (N3072, N3051, N3061);
buf BUF1 (N3073, N3069);
not NOT1 (N3074, N3070);
or OR4 (N3075, N3063, N2790, N520, N156);
nand NAND3 (N3076, N3071, N2049, N469);
not NOT1 (N3077, N3068);
and AND3 (N3078, N3077, N2419, N2683);
or OR3 (N3079, N3073, N2512, N2008);
xor XOR2 (N3080, N3078, N2490);
nor NOR3 (N3081, N3066, N2651, N362);
not NOT1 (N3082, N3076);
xor XOR2 (N3083, N3060, N2976);
nand NAND3 (N3084, N3072, N794, N821);
nor NOR4 (N3085, N3074, N2470, N2677, N40);
nand NAND2 (N3086, N3081, N937);
not NOT1 (N3087, N3084);
nor NOR2 (N3088, N3085, N1535);
or OR3 (N3089, N3088, N1391, N774);
buf BUF1 (N3090, N3080);
buf BUF1 (N3091, N3045);
or OR4 (N3092, N3075, N978, N2101, N2333);
or OR3 (N3093, N3048, N2724, N278);
or OR3 (N3094, N3091, N2859, N446);
nor NOR2 (N3095, N3087, N2147);
nor NOR3 (N3096, N3090, N1634, N1513);
xor XOR2 (N3097, N3086, N1801);
nand NAND2 (N3098, N3079, N1516);
and AND3 (N3099, N3082, N2120, N2893);
buf BUF1 (N3100, N3099);
xor XOR2 (N3101, N3098, N755);
nor NOR4 (N3102, N3097, N2516, N945, N2768);
xor XOR2 (N3103, N3095, N637);
xor XOR2 (N3104, N3101, N387);
nand NAND2 (N3105, N3103, N1175);
not NOT1 (N3106, N3094);
and AND2 (N3107, N3092, N266);
nand NAND4 (N3108, N3093, N2491, N2467, N2015);
buf BUF1 (N3109, N3106);
and AND4 (N3110, N3105, N307, N1764, N625);
nand NAND2 (N3111, N3096, N3060);
nand NAND4 (N3112, N3104, N728, N2091, N704);
nor NOR3 (N3113, N3112, N769, N2278);
buf BUF1 (N3114, N3089);
nor NOR3 (N3115, N3111, N2328, N1108);
xor XOR2 (N3116, N3083, N1840);
xor XOR2 (N3117, N3110, N2655);
not NOT1 (N3118, N3102);
buf BUF1 (N3119, N3117);
xor XOR2 (N3120, N3113, N1677);
buf BUF1 (N3121, N3115);
or OR2 (N3122, N3100, N646);
not NOT1 (N3123, N3109);
and AND2 (N3124, N3116, N88);
not NOT1 (N3125, N3123);
buf BUF1 (N3126, N3107);
xor XOR2 (N3127, N3108, N1979);
not NOT1 (N3128, N3126);
xor XOR2 (N3129, N3121, N1043);
and AND3 (N3130, N3118, N593, N181);
buf BUF1 (N3131, N3130);
or OR3 (N3132, N3120, N2759, N933);
buf BUF1 (N3133, N3129);
and AND2 (N3134, N3128, N1811);
xor XOR2 (N3135, N3127, N882);
not NOT1 (N3136, N3125);
buf BUF1 (N3137, N3134);
or OR3 (N3138, N3136, N2615, N941);
and AND2 (N3139, N3133, N1694);
xor XOR2 (N3140, N3135, N1077);
nand NAND3 (N3141, N3119, N458, N1898);
xor XOR2 (N3142, N3114, N1626);
not NOT1 (N3143, N3140);
nor NOR3 (N3144, N3142, N2358, N463);
nand NAND2 (N3145, N3131, N470);
xor XOR2 (N3146, N3139, N258);
xor XOR2 (N3147, N3145, N3062);
not NOT1 (N3148, N3141);
or OR2 (N3149, N3147, N2296);
xor XOR2 (N3150, N3148, N2313);
or OR2 (N3151, N3124, N3104);
nor NOR3 (N3152, N3150, N804, N730);
not NOT1 (N3153, N3152);
and AND2 (N3154, N3132, N1727);
not NOT1 (N3155, N3151);
and AND4 (N3156, N3138, N2620, N2492, N2669);
nand NAND3 (N3157, N3156, N535, N2762);
not NOT1 (N3158, N3154);
nor NOR2 (N3159, N3153, N2983);
buf BUF1 (N3160, N3146);
xor XOR2 (N3161, N3122, N2671);
nand NAND3 (N3162, N3143, N24, N2683);
and AND4 (N3163, N3155, N2381, N2398, N1830);
not NOT1 (N3164, N3157);
xor XOR2 (N3165, N3160, N308);
not NOT1 (N3166, N3165);
nand NAND2 (N3167, N3162, N2597);
or OR2 (N3168, N3166, N2167);
xor XOR2 (N3169, N3161, N2816);
and AND4 (N3170, N3158, N2893, N3105, N1291);
not NOT1 (N3171, N3149);
or OR2 (N3172, N3170, N2736);
or OR3 (N3173, N3144, N1319, N405);
or OR3 (N3174, N3171, N69, N1662);
buf BUF1 (N3175, N3137);
and AND3 (N3176, N3172, N3072, N2545);
nor NOR4 (N3177, N3168, N2331, N623, N3052);
and AND3 (N3178, N3169, N1834, N1736);
nor NOR3 (N3179, N3173, N220, N1012);
buf BUF1 (N3180, N3179);
and AND3 (N3181, N3176, N2285, N1535);
not NOT1 (N3182, N3174);
and AND4 (N3183, N3182, N1775, N2947, N1965);
xor XOR2 (N3184, N3183, N1628);
or OR3 (N3185, N3178, N2853, N2712);
nor NOR4 (N3186, N3164, N8, N255, N2608);
nand NAND2 (N3187, N3185, N1269);
nand NAND2 (N3188, N3184, N2977);
xor XOR2 (N3189, N3159, N523);
nand NAND2 (N3190, N3167, N2755);
not NOT1 (N3191, N3187);
nand NAND2 (N3192, N3163, N1553);
xor XOR2 (N3193, N3191, N268);
nor NOR2 (N3194, N3188, N47);
or OR4 (N3195, N3189, N1735, N3119, N180);
xor XOR2 (N3196, N3175, N2704);
nand NAND4 (N3197, N3177, N2756, N663, N380);
nand NAND4 (N3198, N3194, N2513, N2216, N1908);
or OR4 (N3199, N3190, N563, N2907, N565);
xor XOR2 (N3200, N3192, N289);
nor NOR3 (N3201, N3199, N3001, N3110);
nor NOR3 (N3202, N3197, N2305, N1393);
xor XOR2 (N3203, N3193, N2662);
buf BUF1 (N3204, N3180);
nor NOR3 (N3205, N3186, N2427, N1212);
and AND2 (N3206, N3196, N2208);
not NOT1 (N3207, N3198);
nand NAND3 (N3208, N3200, N2416, N1597);
nor NOR3 (N3209, N3208, N2623, N52);
nand NAND4 (N3210, N3201, N1433, N2026, N678);
not NOT1 (N3211, N3204);
nand NAND2 (N3212, N3209, N973);
and AND3 (N3213, N3181, N1122, N1313);
nand NAND4 (N3214, N3207, N1787, N651, N2013);
or OR2 (N3215, N3210, N2661);
not NOT1 (N3216, N3203);
and AND2 (N3217, N3214, N1607);
or OR4 (N3218, N3212, N66, N2937, N1446);
nand NAND3 (N3219, N3206, N267, N2921);
buf BUF1 (N3220, N3216);
buf BUF1 (N3221, N3213);
not NOT1 (N3222, N3220);
and AND2 (N3223, N3215, N3120);
not NOT1 (N3224, N3219);
nor NOR3 (N3225, N3221, N2595, N2192);
nor NOR4 (N3226, N3223, N1552, N844, N1199);
buf BUF1 (N3227, N3211);
nor NOR4 (N3228, N3224, N925, N1200, N292);
buf BUF1 (N3229, N3228);
nor NOR3 (N3230, N3218, N2724, N903);
and AND2 (N3231, N3195, N1065);
or OR3 (N3232, N3227, N2804, N2573);
buf BUF1 (N3233, N3230);
nand NAND4 (N3234, N3205, N1252, N3005, N1182);
not NOT1 (N3235, N3222);
nand NAND4 (N3236, N3234, N171, N1342, N3218);
xor XOR2 (N3237, N3236, N1730);
xor XOR2 (N3238, N3202, N906);
or OR4 (N3239, N3237, N1202, N2145, N1072);
nand NAND3 (N3240, N3225, N2474, N2307);
nor NOR3 (N3241, N3235, N152, N2987);
nor NOR2 (N3242, N3241, N844);
nor NOR2 (N3243, N3217, N2407);
not NOT1 (N3244, N3243);
buf BUF1 (N3245, N3240);
xor XOR2 (N3246, N3233, N2721);
nand NAND3 (N3247, N3231, N1495, N1047);
nand NAND4 (N3248, N3229, N1291, N2315, N106);
not NOT1 (N3249, N3244);
xor XOR2 (N3250, N3249, N1142);
and AND2 (N3251, N3226, N566);
xor XOR2 (N3252, N3250, N1233);
buf BUF1 (N3253, N3232);
or OR2 (N3254, N3247, N792);
and AND2 (N3255, N3253, N2640);
and AND3 (N3256, N3246, N771, N2960);
not NOT1 (N3257, N3252);
xor XOR2 (N3258, N3257, N806);
nand NAND2 (N3259, N3255, N868);
nand NAND2 (N3260, N3251, N1149);
buf BUF1 (N3261, N3238);
or OR2 (N3262, N3245, N1844);
nor NOR2 (N3263, N3256, N2673);
or OR3 (N3264, N3239, N912, N1012);
nor NOR2 (N3265, N3258, N2932);
nor NOR3 (N3266, N3248, N1697, N1507);
and AND2 (N3267, N3259, N2070);
and AND3 (N3268, N3267, N2753, N2326);
nand NAND3 (N3269, N3268, N625, N2123);
and AND4 (N3270, N3260, N481, N1185, N1936);
not NOT1 (N3271, N3254);
xor XOR2 (N3272, N3271, N1755);
nand NAND3 (N3273, N3242, N1007, N37);
buf BUF1 (N3274, N3262);
not NOT1 (N3275, N3274);
nand NAND3 (N3276, N3266, N133, N285);
or OR2 (N3277, N3275, N2837);
not NOT1 (N3278, N3272);
buf BUF1 (N3279, N3278);
xor XOR2 (N3280, N3273, N1249);
not NOT1 (N3281, N3269);
nand NAND4 (N3282, N3265, N3007, N211, N2760);
buf BUF1 (N3283, N3270);
or OR3 (N3284, N3263, N131, N3213);
xor XOR2 (N3285, N3277, N507);
nor NOR3 (N3286, N3283, N56, N2513);
and AND3 (N3287, N3276, N269, N1981);
not NOT1 (N3288, N3279);
xor XOR2 (N3289, N3280, N1477);
nor NOR3 (N3290, N3264, N1680, N3205);
or OR4 (N3291, N3289, N3236, N1237, N2191);
nor NOR2 (N3292, N3281, N2355);
buf BUF1 (N3293, N3261);
or OR2 (N3294, N3287, N2882);
xor XOR2 (N3295, N3282, N1228);
xor XOR2 (N3296, N3295, N1644);
xor XOR2 (N3297, N3285, N1565);
nand NAND2 (N3298, N3286, N2025);
xor XOR2 (N3299, N3290, N1983);
nor NOR2 (N3300, N3291, N1639);
xor XOR2 (N3301, N3300, N3047);
nand NAND4 (N3302, N3288, N2282, N686, N603);
not NOT1 (N3303, N3302);
nand NAND4 (N3304, N3294, N97, N1458, N3292);
and AND4 (N3305, N1976, N2857, N2566, N3056);
or OR3 (N3306, N3293, N3019, N389);
nor NOR3 (N3307, N3297, N2558, N2772);
nand NAND2 (N3308, N3304, N197);
xor XOR2 (N3309, N3308, N1833);
xor XOR2 (N3310, N3307, N3216);
buf BUF1 (N3311, N3309);
buf BUF1 (N3312, N3311);
or OR4 (N3313, N3299, N1765, N3102, N917);
buf BUF1 (N3314, N3296);
nor NOR3 (N3315, N3312, N2056, N787);
nor NOR2 (N3316, N3301, N2063);
and AND3 (N3317, N3306, N1739, N810);
and AND3 (N3318, N3303, N2657, N3296);
or OR4 (N3319, N3310, N2900, N1555, N1383);
nand NAND3 (N3320, N3318, N2664, N1258);
and AND3 (N3321, N3284, N953, N1099);
buf BUF1 (N3322, N3315);
buf BUF1 (N3323, N3298);
buf BUF1 (N3324, N3314);
or OR3 (N3325, N3322, N3108, N2671);
not NOT1 (N3326, N3319);
nor NOR2 (N3327, N3324, N454);
nand NAND2 (N3328, N3316, N885);
buf BUF1 (N3329, N3323);
buf BUF1 (N3330, N3327);
nand NAND4 (N3331, N3320, N611, N591, N2057);
and AND4 (N3332, N3313, N3219, N952, N1999);
or OR2 (N3333, N3305, N1549);
xor XOR2 (N3334, N3326, N2769);
xor XOR2 (N3335, N3330, N1742);
buf BUF1 (N3336, N3333);
or OR2 (N3337, N3329, N2983);
or OR2 (N3338, N3334, N2990);
nor NOR2 (N3339, N3317, N2254);
or OR2 (N3340, N3331, N42);
nand NAND2 (N3341, N3328, N1474);
not NOT1 (N3342, N3332);
nor NOR3 (N3343, N3340, N2788, N3092);
or OR4 (N3344, N3341, N773, N135, N2335);
or OR4 (N3345, N3325, N1185, N468, N2754);
not NOT1 (N3346, N3336);
not NOT1 (N3347, N3345);
nand NAND3 (N3348, N3347, N3143, N2037);
and AND3 (N3349, N3342, N56, N287);
and AND2 (N3350, N3321, N1345);
buf BUF1 (N3351, N3349);
buf BUF1 (N3352, N3348);
nor NOR2 (N3353, N3335, N596);
nor NOR3 (N3354, N3337, N1333, N2581);
xor XOR2 (N3355, N3343, N120);
not NOT1 (N3356, N3351);
buf BUF1 (N3357, N3338);
and AND3 (N3358, N3356, N867, N1256);
and AND3 (N3359, N3352, N1544, N2457);
or OR3 (N3360, N3350, N3231, N759);
xor XOR2 (N3361, N3355, N2713);
nor NOR4 (N3362, N3359, N1631, N2720, N3353);
nand NAND3 (N3363, N2219, N90, N1269);
nor NOR2 (N3364, N3357, N1885);
nor NOR2 (N3365, N3354, N467);
and AND3 (N3366, N3339, N2551, N241);
xor XOR2 (N3367, N3344, N1153);
xor XOR2 (N3368, N3366, N794);
buf BUF1 (N3369, N3364);
not NOT1 (N3370, N3346);
or OR2 (N3371, N3363, N1680);
xor XOR2 (N3372, N3360, N1124);
buf BUF1 (N3373, N3371);
not NOT1 (N3374, N3368);
not NOT1 (N3375, N3374);
not NOT1 (N3376, N3372);
xor XOR2 (N3377, N3367, N104);
nor NOR2 (N3378, N3362, N3082);
or OR2 (N3379, N3369, N2603);
xor XOR2 (N3380, N3358, N271);
and AND4 (N3381, N3370, N1098, N2091, N327);
xor XOR2 (N3382, N3361, N151);
not NOT1 (N3383, N3380);
or OR2 (N3384, N3365, N417);
not NOT1 (N3385, N3379);
nor NOR2 (N3386, N3385, N2796);
buf BUF1 (N3387, N3386);
nor NOR3 (N3388, N3376, N1014, N198);
xor XOR2 (N3389, N3375, N1081);
xor XOR2 (N3390, N3388, N696);
buf BUF1 (N3391, N3383);
nor NOR4 (N3392, N3373, N2297, N3337, N2971);
not NOT1 (N3393, N3390);
buf BUF1 (N3394, N3393);
not NOT1 (N3395, N3377);
nor NOR4 (N3396, N3378, N454, N547, N551);
xor XOR2 (N3397, N3387, N1424);
or OR4 (N3398, N3384, N1153, N2013, N1688);
buf BUF1 (N3399, N3395);
or OR3 (N3400, N3397, N3141, N2284);
xor XOR2 (N3401, N3399, N1866);
or OR2 (N3402, N3396, N596);
buf BUF1 (N3403, N3401);
or OR3 (N3404, N3381, N4, N2781);
xor XOR2 (N3405, N3382, N2704);
or OR4 (N3406, N3400, N358, N2720, N2626);
and AND3 (N3407, N3394, N3095, N3006);
nor NOR2 (N3408, N3404, N2958);
nor NOR3 (N3409, N3403, N1310, N2879);
and AND2 (N3410, N3391, N2838);
buf BUF1 (N3411, N3410);
buf BUF1 (N3412, N3398);
or OR2 (N3413, N3402, N3103);
nor NOR3 (N3414, N3413, N3058, N1483);
nand NAND2 (N3415, N3405, N837);
nor NOR4 (N3416, N3409, N2093, N1565, N510);
xor XOR2 (N3417, N3412, N2632);
or OR2 (N3418, N3417, N186);
nand NAND2 (N3419, N3411, N1652);
not NOT1 (N3420, N3406);
nor NOR4 (N3421, N3407, N2292, N2810, N307);
or OR4 (N3422, N3419, N131, N973, N1999);
buf BUF1 (N3423, N3408);
or OR2 (N3424, N3421, N958);
xor XOR2 (N3425, N3415, N2570);
xor XOR2 (N3426, N3389, N457);
nand NAND4 (N3427, N3420, N2723, N2119, N1819);
nand NAND3 (N3428, N3426, N2530, N2270);
or OR2 (N3429, N3392, N2277);
or OR3 (N3430, N3416, N3305, N737);
and AND2 (N3431, N3424, N1055);
xor XOR2 (N3432, N3425, N2474);
nand NAND2 (N3433, N3431, N573);
or OR3 (N3434, N3418, N2519, N1880);
xor XOR2 (N3435, N3433, N1971);
nand NAND3 (N3436, N3427, N955, N1433);
and AND3 (N3437, N3430, N3031, N599);
not NOT1 (N3438, N3414);
not NOT1 (N3439, N3435);
not NOT1 (N3440, N3422);
xor XOR2 (N3441, N3429, N3019);
buf BUF1 (N3442, N3428);
buf BUF1 (N3443, N3436);
not NOT1 (N3444, N3437);
or OR4 (N3445, N3439, N1601, N1511, N1343);
buf BUF1 (N3446, N3445);
xor XOR2 (N3447, N3442, N1582);
and AND3 (N3448, N3446, N761, N3396);
nor NOR3 (N3449, N3441, N1822, N2092);
nand NAND3 (N3450, N3440, N1571, N2753);
buf BUF1 (N3451, N3447);
nand NAND4 (N3452, N3451, N1658, N1407, N46);
nor NOR3 (N3453, N3423, N1487, N2305);
not NOT1 (N3454, N3448);
and AND2 (N3455, N3434, N3399);
or OR3 (N3456, N3444, N68, N1748);
not NOT1 (N3457, N3456);
or OR2 (N3458, N3443, N1383);
and AND4 (N3459, N3458, N2270, N811, N3323);
nor NOR3 (N3460, N3450, N1209, N3066);
buf BUF1 (N3461, N3457);
and AND4 (N3462, N3461, N3332, N2440, N983);
not NOT1 (N3463, N3459);
nor NOR3 (N3464, N3460, N3370, N720);
or OR3 (N3465, N3462, N2788, N335);
nand NAND2 (N3466, N3438, N961);
not NOT1 (N3467, N3455);
nand NAND2 (N3468, N3465, N1142);
nor NOR3 (N3469, N3468, N2828, N1045);
nor NOR2 (N3470, N3464, N502);
buf BUF1 (N3471, N3469);
and AND2 (N3472, N3454, N2098);
and AND2 (N3473, N3453, N692);
buf BUF1 (N3474, N3471);
nor NOR2 (N3475, N3474, N3098);
not NOT1 (N3476, N3470);
nor NOR4 (N3477, N3466, N1308, N997, N3083);
xor XOR2 (N3478, N3432, N3098);
not NOT1 (N3479, N3463);
nand NAND2 (N3480, N3452, N3069);
nand NAND3 (N3481, N3477, N2323, N2815);
nor NOR4 (N3482, N3472, N838, N3445, N575);
nand NAND2 (N3483, N3476, N774);
not NOT1 (N3484, N3449);
xor XOR2 (N3485, N3479, N2211);
nand NAND4 (N3486, N3484, N351, N58, N2076);
and AND4 (N3487, N3475, N2595, N819, N350);
nand NAND2 (N3488, N3485, N592);
or OR4 (N3489, N3478, N452, N1145, N3285);
or OR2 (N3490, N3489, N2548);
not NOT1 (N3491, N3481);
xor XOR2 (N3492, N3482, N1209);
xor XOR2 (N3493, N3473, N1801);
nand NAND3 (N3494, N3491, N2678, N1126);
and AND4 (N3495, N3490, N2797, N1270, N1224);
or OR3 (N3496, N3480, N480, N621);
and AND3 (N3497, N3493, N2713, N1213);
or OR4 (N3498, N3483, N2681, N3098, N2799);
or OR2 (N3499, N3492, N682);
not NOT1 (N3500, N3499);
nor NOR2 (N3501, N3500, N765);
buf BUF1 (N3502, N3467);
or OR3 (N3503, N3487, N2685, N2641);
buf BUF1 (N3504, N3502);
nand NAND3 (N3505, N3497, N3208, N2678);
or OR4 (N3506, N3501, N3183, N1658, N2407);
xor XOR2 (N3507, N3498, N2288);
buf BUF1 (N3508, N3486);
nor NOR2 (N3509, N3496, N394);
nor NOR4 (N3510, N3504, N1932, N3279, N2987);
buf BUF1 (N3511, N3495);
nor NOR2 (N3512, N3488, N2051);
not NOT1 (N3513, N3510);
not NOT1 (N3514, N3513);
nor NOR4 (N3515, N3503, N1411, N1746, N1685);
and AND4 (N3516, N3506, N278, N2549, N976);
xor XOR2 (N3517, N3505, N1263);
nand NAND2 (N3518, N3511, N2651);
nand NAND3 (N3519, N3507, N354, N529);
nand NAND4 (N3520, N3516, N112, N3253, N2544);
not NOT1 (N3521, N3515);
and AND2 (N3522, N3519, N2942);
and AND3 (N3523, N3518, N379, N747);
and AND2 (N3524, N3512, N2671);
not NOT1 (N3525, N3508);
nor NOR4 (N3526, N3520, N1090, N611, N1598);
xor XOR2 (N3527, N3526, N851);
nor NOR3 (N3528, N3527, N3159, N2926);
nand NAND2 (N3529, N3494, N2632);
buf BUF1 (N3530, N3523);
buf BUF1 (N3531, N3530);
nand NAND4 (N3532, N3531, N2905, N2533, N1638);
not NOT1 (N3533, N3509);
buf BUF1 (N3534, N3514);
xor XOR2 (N3535, N3529, N461);
and AND4 (N3536, N3532, N3216, N911, N2618);
xor XOR2 (N3537, N3533, N974);
buf BUF1 (N3538, N3525);
and AND4 (N3539, N3517, N2001, N686, N889);
buf BUF1 (N3540, N3534);
xor XOR2 (N3541, N3522, N1996);
and AND4 (N3542, N3538, N1371, N3036, N1276);
nor NOR4 (N3543, N3536, N496, N3390, N1015);
xor XOR2 (N3544, N3535, N2250);
not NOT1 (N3545, N3542);
nand NAND3 (N3546, N3541, N2020, N1471);
xor XOR2 (N3547, N3543, N3150);
nand NAND4 (N3548, N3540, N1602, N2494, N48);
xor XOR2 (N3549, N3544, N2733);
not NOT1 (N3550, N3537);
xor XOR2 (N3551, N3528, N1217);
not NOT1 (N3552, N3539);
xor XOR2 (N3553, N3552, N2685);
nand NAND3 (N3554, N3548, N3112, N1014);
not NOT1 (N3555, N3545);
and AND3 (N3556, N3546, N1812, N894);
not NOT1 (N3557, N3524);
or OR4 (N3558, N3521, N1589, N2707, N3013);
or OR3 (N3559, N3553, N545, N1117);
or OR3 (N3560, N3549, N2905, N1050);
nor NOR3 (N3561, N3559, N3532, N1558);
nand NAND4 (N3562, N3550, N485, N833, N2088);
not NOT1 (N3563, N3562);
nor NOR3 (N3564, N3560, N2931, N3086);
or OR3 (N3565, N3561, N3297, N137);
nor NOR2 (N3566, N3555, N670);
nor NOR3 (N3567, N3566, N1339, N613);
buf BUF1 (N3568, N3567);
nor NOR4 (N3569, N3557, N1560, N1501, N107);
nand NAND3 (N3570, N3563, N1855, N546);
and AND3 (N3571, N3554, N2137, N2349);
and AND3 (N3572, N3551, N2503, N225);
nand NAND3 (N3573, N3558, N841, N291);
and AND3 (N3574, N3568, N133, N2641);
nor NOR4 (N3575, N3570, N266, N1007, N373);
nand NAND4 (N3576, N3556, N2568, N843, N15);
not NOT1 (N3577, N3574);
nand NAND4 (N3578, N3575, N371, N2374, N272);
and AND4 (N3579, N3564, N1116, N2923, N212);
not NOT1 (N3580, N3573);
nor NOR2 (N3581, N3547, N1520);
nand NAND2 (N3582, N3569, N1018);
and AND3 (N3583, N3577, N2899, N2224);
buf BUF1 (N3584, N3579);
xor XOR2 (N3585, N3580, N754);
nand NAND2 (N3586, N3585, N3138);
and AND3 (N3587, N3583, N431, N60);
nand NAND3 (N3588, N3572, N1638, N1388);
buf BUF1 (N3589, N3586);
not NOT1 (N3590, N3589);
nand NAND4 (N3591, N3587, N999, N508, N416);
or OR3 (N3592, N3590, N659, N2610);
xor XOR2 (N3593, N3576, N267);
not NOT1 (N3594, N3584);
or OR4 (N3595, N3591, N2771, N1065, N719);
not NOT1 (N3596, N3578);
not NOT1 (N3597, N3594);
or OR2 (N3598, N3593, N1991);
not NOT1 (N3599, N3592);
nand NAND2 (N3600, N3582, N1176);
or OR4 (N3601, N3599, N3219, N3263, N3366);
xor XOR2 (N3602, N3597, N2716);
not NOT1 (N3603, N3598);
buf BUF1 (N3604, N3596);
nor NOR2 (N3605, N3603, N2003);
and AND2 (N3606, N3588, N1912);
nand NAND2 (N3607, N3571, N878);
nand NAND4 (N3608, N3604, N3484, N1615, N336);
or OR4 (N3609, N3606, N1908, N1088, N2363);
nand NAND4 (N3610, N3595, N3004, N452, N3339);
and AND4 (N3611, N3608, N2718, N1931, N1534);
and AND2 (N3612, N3600, N1805);
buf BUF1 (N3613, N3565);
nor NOR4 (N3614, N3609, N1325, N1898, N56);
not NOT1 (N3615, N3613);
nor NOR4 (N3616, N3612, N2173, N2627, N565);
buf BUF1 (N3617, N3605);
or OR2 (N3618, N3601, N1562);
and AND2 (N3619, N3611, N2864);
buf BUF1 (N3620, N3617);
and AND4 (N3621, N3614, N776, N3068, N2176);
nand NAND3 (N3622, N3620, N2988, N724);
not NOT1 (N3623, N3610);
nor NOR4 (N3624, N3607, N3434, N3029, N365);
not NOT1 (N3625, N3615);
or OR2 (N3626, N3624, N2530);
or OR3 (N3627, N3602, N550, N1789);
xor XOR2 (N3628, N3621, N3485);
buf BUF1 (N3629, N3628);
xor XOR2 (N3630, N3618, N692);
nor NOR3 (N3631, N3619, N3115, N1516);
and AND4 (N3632, N3616, N1896, N3599, N2537);
nand NAND4 (N3633, N3629, N1942, N1808, N2810);
xor XOR2 (N3634, N3633, N1125);
and AND4 (N3635, N3626, N2005, N2347, N1662);
nand NAND2 (N3636, N3581, N511);
not NOT1 (N3637, N3634);
not NOT1 (N3638, N3625);
buf BUF1 (N3639, N3630);
nor NOR3 (N3640, N3627, N1386, N3070);
and AND2 (N3641, N3639, N362);
nor NOR3 (N3642, N3622, N1108, N932);
not NOT1 (N3643, N3623);
nand NAND4 (N3644, N3640, N2643, N272, N525);
xor XOR2 (N3645, N3637, N3491);
not NOT1 (N3646, N3631);
nand NAND3 (N3647, N3641, N72, N3004);
not NOT1 (N3648, N3632);
not NOT1 (N3649, N3645);
nand NAND4 (N3650, N3644, N2407, N742, N1270);
nor NOR4 (N3651, N3647, N2203, N137, N1386);
xor XOR2 (N3652, N3636, N3176);
or OR4 (N3653, N3650, N2639, N1747, N2492);
nor NOR4 (N3654, N3642, N292, N1116, N2157);
nor NOR4 (N3655, N3649, N2544, N1951, N2205);
not NOT1 (N3656, N3653);
buf BUF1 (N3657, N3655);
nor NOR2 (N3658, N3651, N1243);
not NOT1 (N3659, N3657);
nor NOR3 (N3660, N3638, N3116, N1111);
nor NOR2 (N3661, N3654, N1921);
not NOT1 (N3662, N3646);
not NOT1 (N3663, N3635);
buf BUF1 (N3664, N3661);
not NOT1 (N3665, N3663);
and AND2 (N3666, N3664, N2716);
or OR4 (N3667, N3643, N1224, N1001, N2504);
or OR2 (N3668, N3652, N2158);
nor NOR3 (N3669, N3666, N250, N1578);
nor NOR3 (N3670, N3660, N1318, N2922);
buf BUF1 (N3671, N3667);
and AND2 (N3672, N3648, N2830);
nand NAND4 (N3673, N3662, N3171, N2415, N208);
buf BUF1 (N3674, N3673);
nor NOR2 (N3675, N3658, N274);
nor NOR3 (N3676, N3668, N2985, N1327);
not NOT1 (N3677, N3656);
not NOT1 (N3678, N3677);
not NOT1 (N3679, N3669);
and AND2 (N3680, N3675, N727);
or OR3 (N3681, N3679, N884, N970);
nand NAND4 (N3682, N3678, N2329, N2888, N3161);
or OR3 (N3683, N3672, N1783, N410);
nor NOR4 (N3684, N3671, N239, N618, N2951);
and AND3 (N3685, N3670, N669, N3363);
not NOT1 (N3686, N3681);
buf BUF1 (N3687, N3659);
xor XOR2 (N3688, N3687, N1509);
nand NAND2 (N3689, N3674, N2290);
or OR3 (N3690, N3676, N643, N2114);
nor NOR2 (N3691, N3690, N911);
nand NAND3 (N3692, N3688, N2180, N2911);
nor NOR4 (N3693, N3689, N3107, N2281, N2252);
or OR3 (N3694, N3683, N2146, N2397);
nand NAND2 (N3695, N3691, N3130);
buf BUF1 (N3696, N3665);
and AND4 (N3697, N3686, N2800, N2985, N30);
buf BUF1 (N3698, N3695);
nand NAND4 (N3699, N3697, N752, N1370, N164);
and AND4 (N3700, N3680, N1895, N211, N642);
and AND3 (N3701, N3685, N63, N70);
buf BUF1 (N3702, N3698);
xor XOR2 (N3703, N3699, N1468);
nand NAND4 (N3704, N3702, N446, N326, N3167);
nor NOR3 (N3705, N3701, N3560, N3268);
buf BUF1 (N3706, N3696);
or OR4 (N3707, N3706, N546, N3610, N1591);
not NOT1 (N3708, N3703);
or OR2 (N3709, N3708, N3605);
buf BUF1 (N3710, N3704);
nand NAND4 (N3711, N3694, N1713, N3016, N1154);
xor XOR2 (N3712, N3709, N3314);
buf BUF1 (N3713, N3707);
buf BUF1 (N3714, N3713);
or OR4 (N3715, N3714, N1028, N263, N2260);
xor XOR2 (N3716, N3693, N563);
nand NAND2 (N3717, N3712, N2240);
or OR2 (N3718, N3710, N1064);
nor NOR2 (N3719, N3692, N3302);
and AND2 (N3720, N3700, N583);
nand NAND3 (N3721, N3717, N2886, N857);
or OR3 (N3722, N3705, N1236, N2177);
buf BUF1 (N3723, N3721);
nand NAND4 (N3724, N3718, N3059, N1242, N680);
or OR2 (N3725, N3716, N1145);
not NOT1 (N3726, N3715);
nor NOR3 (N3727, N3722, N1137, N305);
not NOT1 (N3728, N3723);
xor XOR2 (N3729, N3711, N981);
and AND2 (N3730, N3719, N1105);
and AND2 (N3731, N3729, N1091);
or OR4 (N3732, N3682, N1416, N2684, N3229);
nand NAND2 (N3733, N3684, N1268);
xor XOR2 (N3734, N3726, N361);
nand NAND3 (N3735, N3725, N141, N2231);
or OR4 (N3736, N3730, N1064, N1106, N3319);
or OR3 (N3737, N3727, N1366, N949);
nor NOR3 (N3738, N3733, N3633, N70);
or OR4 (N3739, N3734, N624, N1357, N376);
and AND2 (N3740, N3731, N3437);
nor NOR2 (N3741, N3728, N2709);
and AND2 (N3742, N3724, N2151);
or OR2 (N3743, N3737, N2208);
and AND3 (N3744, N3743, N1815, N809);
or OR2 (N3745, N3720, N2210);
or OR2 (N3746, N3742, N326);
and AND4 (N3747, N3739, N30, N805, N1708);
and AND4 (N3748, N3741, N351, N2049, N3602);
nand NAND3 (N3749, N3736, N2346, N3298);
and AND4 (N3750, N3745, N776, N1395, N2475);
buf BUF1 (N3751, N3750);
not NOT1 (N3752, N3735);
and AND2 (N3753, N3749, N2784);
nand NAND2 (N3754, N3751, N1344);
xor XOR2 (N3755, N3738, N1223);
not NOT1 (N3756, N3732);
nand NAND2 (N3757, N3746, N996);
nand NAND2 (N3758, N3744, N480);
nor NOR3 (N3759, N3747, N3291, N1308);
xor XOR2 (N3760, N3740, N1721);
xor XOR2 (N3761, N3755, N944);
buf BUF1 (N3762, N3752);
nand NAND4 (N3763, N3762, N3664, N3033, N2023);
or OR3 (N3764, N3754, N3348, N394);
and AND4 (N3765, N3763, N3760, N1175, N743);
nor NOR2 (N3766, N3114, N3706);
not NOT1 (N3767, N3748);
buf BUF1 (N3768, N3759);
xor XOR2 (N3769, N3756, N1446);
nand NAND2 (N3770, N3769, N1391);
or OR4 (N3771, N3753, N2339, N1714, N1916);
xor XOR2 (N3772, N3764, N2496);
buf BUF1 (N3773, N3771);
nor NOR4 (N3774, N3767, N258, N439, N280);
nor NOR2 (N3775, N3766, N49);
and AND4 (N3776, N3757, N2804, N3685, N3700);
nor NOR4 (N3777, N3765, N1925, N3701, N3595);
and AND4 (N3778, N3768, N985, N136, N1027);
nand NAND3 (N3779, N3777, N237, N871);
buf BUF1 (N3780, N3761);
buf BUF1 (N3781, N3776);
nor NOR4 (N3782, N3779, N2, N299, N803);
nand NAND4 (N3783, N3780, N1131, N3607, N964);
not NOT1 (N3784, N3774);
buf BUF1 (N3785, N3773);
buf BUF1 (N3786, N3781);
or OR3 (N3787, N3772, N763, N527);
nand NAND2 (N3788, N3787, N2130);
or OR4 (N3789, N3785, N144, N1590, N3334);
nand NAND3 (N3790, N3770, N1043, N2802);
buf BUF1 (N3791, N3786);
or OR2 (N3792, N3790, N2808);
buf BUF1 (N3793, N3789);
or OR3 (N3794, N3793, N3435, N79);
nand NAND4 (N3795, N3775, N959, N2377, N175);
buf BUF1 (N3796, N3794);
buf BUF1 (N3797, N3784);
not NOT1 (N3798, N3792);
and AND3 (N3799, N3778, N1131, N901);
nand NAND2 (N3800, N3788, N3235);
nand NAND3 (N3801, N3797, N627, N2030);
xor XOR2 (N3802, N3758, N1546);
buf BUF1 (N3803, N3799);
xor XOR2 (N3804, N3803, N3199);
nand NAND2 (N3805, N3804, N541);
not NOT1 (N3806, N3805);
nor NOR4 (N3807, N3806, N456, N846, N1362);
or OR2 (N3808, N3795, N3191);
buf BUF1 (N3809, N3801);
nand NAND3 (N3810, N3800, N1402, N3630);
not NOT1 (N3811, N3807);
or OR3 (N3812, N3791, N556, N1396);
or OR4 (N3813, N3783, N664, N803, N2469);
not NOT1 (N3814, N3809);
not NOT1 (N3815, N3814);
nor NOR3 (N3816, N3813, N922, N2590);
nand NAND3 (N3817, N3810, N2521, N3226);
not NOT1 (N3818, N3802);
xor XOR2 (N3819, N3796, N3104);
buf BUF1 (N3820, N3812);
not NOT1 (N3821, N3820);
and AND4 (N3822, N3819, N943, N121, N2577);
and AND3 (N3823, N3811, N1168, N1337);
and AND3 (N3824, N3815, N2556, N2752);
or OR2 (N3825, N3818, N2168);
xor XOR2 (N3826, N3823, N1267);
and AND4 (N3827, N3817, N1535, N1080, N32);
or OR4 (N3828, N3826, N1474, N3487, N3819);
buf BUF1 (N3829, N3798);
nand NAND4 (N3830, N3827, N2553, N1947, N2682);
or OR2 (N3831, N3828, N1102);
nand NAND4 (N3832, N3816, N1600, N2768, N1098);
or OR4 (N3833, N3821, N3719, N465, N2678);
or OR3 (N3834, N3825, N1575, N3619);
buf BUF1 (N3835, N3829);
buf BUF1 (N3836, N3834);
and AND3 (N3837, N3835, N1132, N661);
or OR2 (N3838, N3824, N283);
and AND3 (N3839, N3808, N587, N1270);
xor XOR2 (N3840, N3831, N2164);
and AND4 (N3841, N3836, N954, N2249, N2430);
xor XOR2 (N3842, N3837, N166);
not NOT1 (N3843, N3839);
or OR2 (N3844, N3832, N528);
buf BUF1 (N3845, N3841);
and AND3 (N3846, N3822, N3394, N2985);
and AND3 (N3847, N3838, N3493, N2072);
and AND2 (N3848, N3840, N1853);
nor NOR4 (N3849, N3848, N2761, N2767, N2490);
xor XOR2 (N3850, N3845, N2197);
xor XOR2 (N3851, N3833, N537);
not NOT1 (N3852, N3843);
and AND3 (N3853, N3842, N505, N3385);
or OR2 (N3854, N3851, N2573);
not NOT1 (N3855, N3846);
not NOT1 (N3856, N3850);
or OR4 (N3857, N3855, N369, N2071, N2049);
buf BUF1 (N3858, N3782);
buf BUF1 (N3859, N3844);
nand NAND4 (N3860, N3853, N250, N1570, N2967);
nand NAND3 (N3861, N3849, N1549, N2631);
nor NOR4 (N3862, N3859, N2719, N495, N2005);
and AND2 (N3863, N3854, N145);
not NOT1 (N3864, N3847);
or OR3 (N3865, N3860, N1468, N3358);
xor XOR2 (N3866, N3858, N1021);
xor XOR2 (N3867, N3862, N2203);
or OR4 (N3868, N3867, N1196, N1153, N2036);
buf BUF1 (N3869, N3861);
not NOT1 (N3870, N3864);
xor XOR2 (N3871, N3868, N147);
nor NOR3 (N3872, N3856, N2389, N1798);
buf BUF1 (N3873, N3870);
and AND3 (N3874, N3863, N296, N1296);
xor XOR2 (N3875, N3871, N1384);
not NOT1 (N3876, N3857);
and AND3 (N3877, N3865, N1503, N3577);
or OR4 (N3878, N3872, N1552, N3048, N2609);
and AND4 (N3879, N3873, N397, N2014, N476);
not NOT1 (N3880, N3877);
nand NAND4 (N3881, N3879, N3605, N3198, N2940);
xor XOR2 (N3882, N3852, N2946);
or OR3 (N3883, N3882, N1209, N1069);
buf BUF1 (N3884, N3830);
xor XOR2 (N3885, N3874, N1241);
buf BUF1 (N3886, N3883);
buf BUF1 (N3887, N3881);
nor NOR3 (N3888, N3866, N1256, N2414);
xor XOR2 (N3889, N3887, N708);
and AND2 (N3890, N3875, N3429);
not NOT1 (N3891, N3869);
nor NOR2 (N3892, N3878, N1647);
xor XOR2 (N3893, N3876, N3361);
nor NOR2 (N3894, N3890, N3620);
nor NOR2 (N3895, N3891, N1590);
xor XOR2 (N3896, N3888, N1179);
buf BUF1 (N3897, N3894);
nand NAND4 (N3898, N3889, N3477, N225, N1967);
nand NAND3 (N3899, N3897, N2325, N3569);
xor XOR2 (N3900, N3896, N867);
not NOT1 (N3901, N3899);
buf BUF1 (N3902, N3880);
and AND2 (N3903, N3900, N508);
buf BUF1 (N3904, N3885);
xor XOR2 (N3905, N3892, N2225);
nand NAND4 (N3906, N3903, N729, N47, N2191);
nand NAND3 (N3907, N3902, N1563, N59);
nor NOR3 (N3908, N3904, N2271, N2161);
xor XOR2 (N3909, N3884, N2938);
buf BUF1 (N3910, N3906);
or OR4 (N3911, N3907, N2896, N2432, N323);
not NOT1 (N3912, N3905);
nand NAND4 (N3913, N3895, N2891, N1793, N1157);
not NOT1 (N3914, N3886);
buf BUF1 (N3915, N3898);
or OR3 (N3916, N3901, N785, N3591);
not NOT1 (N3917, N3916);
not NOT1 (N3918, N3913);
nand NAND2 (N3919, N3915, N2952);
buf BUF1 (N3920, N3909);
buf BUF1 (N3921, N3918);
or OR2 (N3922, N3914, N434);
not NOT1 (N3923, N3922);
nand NAND4 (N3924, N3908, N579, N1968, N1401);
or OR3 (N3925, N3910, N1944, N3817);
xor XOR2 (N3926, N3923, N541);
or OR2 (N3927, N3919, N3503);
nor NOR3 (N3928, N3920, N520, N924);
or OR3 (N3929, N3926, N3908, N2036);
buf BUF1 (N3930, N3893);
xor XOR2 (N3931, N3929, N1947);
nand NAND2 (N3932, N3928, N1768);
not NOT1 (N3933, N3925);
buf BUF1 (N3934, N3931);
not NOT1 (N3935, N3927);
nand NAND3 (N3936, N3917, N3778, N2390);
xor XOR2 (N3937, N3935, N173);
not NOT1 (N3938, N3911);
not NOT1 (N3939, N3930);
nor NOR4 (N3940, N3934, N647, N615, N3352);
nand NAND3 (N3941, N3939, N543, N80);
nor NOR3 (N3942, N3912, N3744, N3815);
or OR4 (N3943, N3932, N1614, N475, N1691);
nand NAND2 (N3944, N3941, N3861);
nor NOR4 (N3945, N3942, N3515, N918, N44);
buf BUF1 (N3946, N3921);
nor NOR2 (N3947, N3933, N1506);
or OR3 (N3948, N3947, N2275, N1040);
not NOT1 (N3949, N3944);
or OR2 (N3950, N3946, N1262);
xor XOR2 (N3951, N3924, N3621);
and AND3 (N3952, N3948, N3407, N2529);
not NOT1 (N3953, N3952);
or OR4 (N3954, N3937, N1084, N3231, N1771);
and AND4 (N3955, N3949, N1476, N3893, N1977);
not NOT1 (N3956, N3945);
and AND2 (N3957, N3936, N701);
not NOT1 (N3958, N3951);
not NOT1 (N3959, N3938);
or OR2 (N3960, N3940, N2469);
not NOT1 (N3961, N3953);
and AND2 (N3962, N3950, N1533);
nor NOR4 (N3963, N3955, N1305, N730, N504);
or OR2 (N3964, N3954, N590);
or OR2 (N3965, N3959, N3521);
not NOT1 (N3966, N3963);
nand NAND4 (N3967, N3957, N3549, N3677, N3063);
buf BUF1 (N3968, N3958);
nor NOR2 (N3969, N3967, N2139);
nand NAND3 (N3970, N3943, N1845, N1350);
xor XOR2 (N3971, N3964, N2729);
xor XOR2 (N3972, N3956, N2279);
nand NAND4 (N3973, N3968, N2008, N1868, N1976);
nand NAND2 (N3974, N3965, N3526);
nand NAND2 (N3975, N3966, N3679);
nor NOR2 (N3976, N3970, N419);
not NOT1 (N3977, N3969);
or OR3 (N3978, N3974, N3445, N2857);
not NOT1 (N3979, N3972);
not NOT1 (N3980, N3975);
nor NOR4 (N3981, N3978, N2824, N1118, N336);
or OR3 (N3982, N3979, N2289, N639);
nand NAND2 (N3983, N3961, N8);
nand NAND2 (N3984, N3977, N2842);
nor NOR4 (N3985, N3962, N3619, N894, N591);
buf BUF1 (N3986, N3971);
buf BUF1 (N3987, N3984);
buf BUF1 (N3988, N3985);
nand NAND4 (N3989, N3960, N74, N1122, N2229);
nor NOR4 (N3990, N3981, N289, N2503, N3722);
nor NOR4 (N3991, N3990, N2363, N3430, N84);
nor NOR4 (N3992, N3991, N2934, N259, N3973);
and AND2 (N3993, N3347, N3722);
nand NAND3 (N3994, N3986, N328, N2398);
nand NAND3 (N3995, N3992, N2931, N2384);
and AND4 (N3996, N3993, N2696, N2124, N1633);
nand NAND3 (N3997, N3994, N301, N1906);
and AND3 (N3998, N3995, N3032, N3382);
or OR3 (N3999, N3996, N1512, N2376);
or OR4 (N4000, N3982, N2096, N3089, N3499);
and AND3 (N4001, N3976, N2811, N2250);
xor XOR2 (N4002, N3983, N3856);
nand NAND2 (N4003, N4000, N1883);
xor XOR2 (N4004, N3980, N2098);
or OR2 (N4005, N3997, N358);
not NOT1 (N4006, N4004);
and AND3 (N4007, N4002, N2862, N1728);
nand NAND3 (N4008, N3999, N2877, N3925);
nand NAND2 (N4009, N4007, N3001);
buf BUF1 (N4010, N4001);
buf BUF1 (N4011, N3988);
and AND4 (N4012, N4006, N2870, N2699, N572);
nand NAND3 (N4013, N4012, N1120, N2980);
buf BUF1 (N4014, N4011);
not NOT1 (N4015, N4003);
nand NAND4 (N4016, N3987, N3074, N3353, N974);
not NOT1 (N4017, N3989);
nor NOR3 (N4018, N4014, N1018, N2863);
buf BUF1 (N4019, N4005);
xor XOR2 (N4020, N4010, N992);
xor XOR2 (N4021, N4013, N293);
not NOT1 (N4022, N4019);
nor NOR4 (N4023, N4018, N510, N2874, N1717);
or OR3 (N4024, N4008, N1270, N3541);
xor XOR2 (N4025, N4017, N2967);
nand NAND4 (N4026, N4016, N2982, N1027, N1657);
nand NAND4 (N4027, N4021, N3275, N841, N3077);
xor XOR2 (N4028, N4023, N2090);
buf BUF1 (N4029, N4020);
xor XOR2 (N4030, N4028, N1216);
or OR2 (N4031, N4029, N1629);
xor XOR2 (N4032, N4027, N1753);
nor NOR2 (N4033, N4022, N386);
or OR2 (N4034, N4033, N3394);
not NOT1 (N4035, N4026);
not NOT1 (N4036, N4034);
nor NOR2 (N4037, N4031, N3347);
buf BUF1 (N4038, N4037);
nand NAND4 (N4039, N4009, N3474, N713, N2979);
nand NAND4 (N4040, N4025, N258, N1768, N550);
xor XOR2 (N4041, N4039, N2759);
and AND3 (N4042, N4036, N3075, N94);
nor NOR3 (N4043, N4040, N3178, N2317);
nand NAND4 (N4044, N4024, N1040, N1397, N995);
and AND4 (N4045, N4030, N3256, N2083, N3898);
buf BUF1 (N4046, N4042);
nand NAND2 (N4047, N4044, N2585);
nand NAND4 (N4048, N4043, N3110, N3220, N2898);
nor NOR4 (N4049, N4041, N2181, N2643, N3455);
and AND2 (N4050, N3998, N1639);
or OR2 (N4051, N4035, N3614);
or OR2 (N4052, N4038, N1822);
not NOT1 (N4053, N4046);
buf BUF1 (N4054, N4050);
or OR4 (N4055, N4045, N704, N3262, N1934);
nand NAND3 (N4056, N4015, N691, N603);
and AND3 (N4057, N4049, N2048, N436);
and AND4 (N4058, N4052, N2548, N3097, N376);
not NOT1 (N4059, N4048);
or OR4 (N4060, N4053, N1873, N174, N1873);
buf BUF1 (N4061, N4047);
not NOT1 (N4062, N4060);
or OR2 (N4063, N4062, N1831);
xor XOR2 (N4064, N4056, N301);
and AND4 (N4065, N4058, N3804, N460, N1735);
buf BUF1 (N4066, N4051);
xor XOR2 (N4067, N4063, N993);
nand NAND2 (N4068, N4054, N51);
and AND2 (N4069, N4068, N1195);
nand NAND3 (N4070, N4032, N2439, N1063);
nor NOR2 (N4071, N4069, N3432);
and AND4 (N4072, N4057, N2515, N425, N1964);
nand NAND2 (N4073, N4064, N3733);
or OR2 (N4074, N4061, N3605);
nor NOR3 (N4075, N4055, N3359, N3957);
or OR2 (N4076, N4065, N272);
buf BUF1 (N4077, N4071);
or OR3 (N4078, N4059, N3010, N3139);
buf BUF1 (N4079, N4066);
nand NAND2 (N4080, N4074, N3360);
buf BUF1 (N4081, N4070);
nand NAND4 (N4082, N4079, N2672, N479, N620);
nand NAND4 (N4083, N4082, N3772, N2749, N568);
and AND2 (N4084, N4072, N4050);
buf BUF1 (N4085, N4075);
nand NAND4 (N4086, N4078, N727, N3094, N3286);
xor XOR2 (N4087, N4084, N1323);
xor XOR2 (N4088, N4077, N2964);
nand NAND3 (N4089, N4076, N2007, N3746);
xor XOR2 (N4090, N4073, N3619);
or OR2 (N4091, N4086, N1723);
not NOT1 (N4092, N4081);
nand NAND4 (N4093, N4092, N3537, N3320, N3226);
xor XOR2 (N4094, N4090, N3972);
nor NOR2 (N4095, N4083, N3074);
nand NAND2 (N4096, N4094, N185);
buf BUF1 (N4097, N4095);
nand NAND2 (N4098, N4097, N3092);
nor NOR2 (N4099, N4087, N1044);
and AND2 (N4100, N4085, N2326);
not NOT1 (N4101, N4096);
or OR2 (N4102, N4100, N664);
nand NAND4 (N4103, N4088, N1849, N1487, N217);
nor NOR3 (N4104, N4099, N2740, N340);
nor NOR4 (N4105, N4101, N2050, N541, N2266);
buf BUF1 (N4106, N4103);
nand NAND3 (N4107, N4080, N2107, N41);
not NOT1 (N4108, N4106);
nand NAND3 (N4109, N4067, N61, N324);
nor NOR3 (N4110, N4105, N2459, N600);
nor NOR3 (N4111, N4108, N2991, N4081);
nand NAND4 (N4112, N4104, N1166, N2189, N4011);
nor NOR3 (N4113, N4093, N2464, N3575);
nor NOR3 (N4114, N4109, N866, N3404);
xor XOR2 (N4115, N4102, N2198);
not NOT1 (N4116, N4091);
not NOT1 (N4117, N4116);
or OR3 (N4118, N4113, N913, N2231);
buf BUF1 (N4119, N4118);
and AND4 (N4120, N4107, N724, N3348, N732);
nand NAND2 (N4121, N4110, N3875);
buf BUF1 (N4122, N4121);
not NOT1 (N4123, N4117);
nand NAND2 (N4124, N4114, N454);
nand NAND3 (N4125, N4089, N3520, N1956);
nor NOR2 (N4126, N4123, N120);
nand NAND3 (N4127, N4120, N2292, N1654);
xor XOR2 (N4128, N4126, N1592);
nand NAND3 (N4129, N4111, N21, N2221);
and AND4 (N4130, N4112, N1427, N858, N2535);
nor NOR4 (N4131, N4127, N1949, N3615, N2354);
or OR3 (N4132, N4115, N1827, N1301);
nand NAND2 (N4133, N4124, N4121);
not NOT1 (N4134, N4131);
not NOT1 (N4135, N4130);
nand NAND2 (N4136, N4119, N924);
or OR4 (N4137, N4132, N1594, N2458, N1759);
xor XOR2 (N4138, N4125, N1683);
buf BUF1 (N4139, N4136);
xor XOR2 (N4140, N4139, N1108);
xor XOR2 (N4141, N4133, N3611);
and AND2 (N4142, N4138, N2285);
and AND4 (N4143, N4140, N458, N3964, N3015);
and AND3 (N4144, N4122, N2853, N2421);
xor XOR2 (N4145, N4142, N2532);
nand NAND4 (N4146, N4098, N2309, N581, N2790);
nand NAND3 (N4147, N4128, N3602, N157);
and AND4 (N4148, N4137, N657, N4126, N3654);
xor XOR2 (N4149, N4148, N2103);
nor NOR4 (N4150, N4135, N2855, N860, N2283);
nor NOR2 (N4151, N4144, N1371);
or OR4 (N4152, N4151, N3094, N1700, N2639);
or OR3 (N4153, N4141, N232, N4078);
buf BUF1 (N4154, N4146);
buf BUF1 (N4155, N4129);
buf BUF1 (N4156, N4150);
buf BUF1 (N4157, N4153);
nand NAND4 (N4158, N4155, N3578, N3153, N2474);
and AND2 (N4159, N4145, N707);
or OR2 (N4160, N4149, N4107);
or OR2 (N4161, N4158, N1731);
not NOT1 (N4162, N4160);
nand NAND3 (N4163, N4152, N1331, N1550);
not NOT1 (N4164, N4159);
not NOT1 (N4165, N4162);
buf BUF1 (N4166, N4134);
or OR2 (N4167, N4154, N2628);
not NOT1 (N4168, N4156);
nor NOR2 (N4169, N4147, N2580);
or OR2 (N4170, N4169, N3451);
nand NAND4 (N4171, N4161, N3278, N1917, N45);
nor NOR3 (N4172, N4167, N2006, N3889);
buf BUF1 (N4173, N4143);
xor XOR2 (N4174, N4171, N3549);
or OR3 (N4175, N4157, N123, N2536);
not NOT1 (N4176, N4172);
nand NAND3 (N4177, N4168, N1520, N1097);
nand NAND2 (N4178, N4164, N2672);
buf BUF1 (N4179, N4178);
and AND3 (N4180, N4179, N2097, N3857);
buf BUF1 (N4181, N4177);
xor XOR2 (N4182, N4175, N1871);
nand NAND4 (N4183, N4163, N3982, N1390, N2563);
not NOT1 (N4184, N4170);
and AND2 (N4185, N4176, N508);
xor XOR2 (N4186, N4182, N3202);
buf BUF1 (N4187, N4183);
and AND4 (N4188, N4165, N574, N3878, N2158);
nor NOR3 (N4189, N4166, N1982, N3867);
not NOT1 (N4190, N4187);
nand NAND2 (N4191, N4184, N1244);
nand NAND3 (N4192, N4188, N3275, N1221);
buf BUF1 (N4193, N4190);
and AND2 (N4194, N4174, N383);
buf BUF1 (N4195, N4181);
nor NOR3 (N4196, N4195, N2495, N3138);
nand NAND3 (N4197, N4180, N3350, N3203);
buf BUF1 (N4198, N4189);
and AND2 (N4199, N4193, N433);
buf BUF1 (N4200, N4185);
buf BUF1 (N4201, N4199);
nor NOR4 (N4202, N4201, N3170, N864, N3447);
nor NOR2 (N4203, N4197, N2673);
nand NAND2 (N4204, N4194, N3661);
and AND4 (N4205, N4186, N4002, N615, N3122);
xor XOR2 (N4206, N4173, N3458);
not NOT1 (N4207, N4203);
not NOT1 (N4208, N4196);
nand NAND4 (N4209, N4200, N2801, N2082, N3838);
or OR3 (N4210, N4202, N3505, N2405);
xor XOR2 (N4211, N4204, N1506);
xor XOR2 (N4212, N4208, N288);
buf BUF1 (N4213, N4205);
xor XOR2 (N4214, N4209, N929);
and AND3 (N4215, N4191, N591, N3526);
not NOT1 (N4216, N4214);
xor XOR2 (N4217, N4215, N1259);
buf BUF1 (N4218, N4210);
and AND4 (N4219, N4198, N3525, N3777, N3995);
nand NAND2 (N4220, N4192, N3029);
nor NOR2 (N4221, N4217, N300);
or OR4 (N4222, N4206, N1050, N1264, N2965);
buf BUF1 (N4223, N4213);
and AND3 (N4224, N4216, N3561, N1354);
xor XOR2 (N4225, N4220, N2288);
or OR4 (N4226, N4224, N2001, N2346, N1894);
not NOT1 (N4227, N4222);
or OR4 (N4228, N4211, N2553, N1920, N3167);
not NOT1 (N4229, N4225);
buf BUF1 (N4230, N4212);
not NOT1 (N4231, N4221);
nand NAND4 (N4232, N4229, N1446, N1452, N3294);
and AND3 (N4233, N4232, N2485, N2692);
nor NOR4 (N4234, N4233, N1535, N450, N685);
xor XOR2 (N4235, N4234, N11);
not NOT1 (N4236, N4230);
not NOT1 (N4237, N4236);
or OR4 (N4238, N4207, N420, N1899, N3289);
and AND4 (N4239, N4227, N389, N2460, N2782);
xor XOR2 (N4240, N4231, N1873);
xor XOR2 (N4241, N4223, N3389);
buf BUF1 (N4242, N4226);
nand NAND3 (N4243, N4237, N3257, N601);
or OR2 (N4244, N4240, N2086);
nor NOR2 (N4245, N4238, N29);
and AND2 (N4246, N4243, N1271);
xor XOR2 (N4247, N4244, N3040);
nand NAND2 (N4248, N4239, N633);
and AND3 (N4249, N4219, N1737, N1921);
and AND4 (N4250, N4241, N1879, N1498, N1065);
nor NOR3 (N4251, N4245, N4197, N2696);
and AND4 (N4252, N4218, N3195, N1281, N4025);
nand NAND3 (N4253, N4247, N1022, N3918);
and AND3 (N4254, N4249, N3486, N3987);
nand NAND2 (N4255, N4250, N3365);
buf BUF1 (N4256, N4251);
or OR4 (N4257, N4254, N204, N580, N643);
buf BUF1 (N4258, N4228);
and AND3 (N4259, N4257, N3626, N294);
or OR2 (N4260, N4252, N4001);
not NOT1 (N4261, N4256);
nand NAND4 (N4262, N4261, N3601, N673, N3018);
not NOT1 (N4263, N4258);
buf BUF1 (N4264, N4260);
not NOT1 (N4265, N4255);
xor XOR2 (N4266, N4263, N987);
or OR4 (N4267, N4259, N2825, N1109, N459);
nand NAND3 (N4268, N4262, N3324, N1807);
and AND4 (N4269, N4242, N1538, N1042, N2177);
nand NAND2 (N4270, N4265, N3448);
nor NOR3 (N4271, N4253, N3059, N2225);
buf BUF1 (N4272, N4248);
not NOT1 (N4273, N4271);
nand NAND2 (N4274, N4246, N2414);
and AND2 (N4275, N4267, N4001);
buf BUF1 (N4276, N4268);
not NOT1 (N4277, N4266);
xor XOR2 (N4278, N4270, N84);
buf BUF1 (N4279, N4275);
buf BUF1 (N4280, N4235);
buf BUF1 (N4281, N4279);
or OR4 (N4282, N4281, N1566, N2641, N184);
nand NAND2 (N4283, N4269, N4139);
and AND2 (N4284, N4272, N3254);
or OR3 (N4285, N4278, N389, N2992);
nand NAND3 (N4286, N4284, N2216, N1116);
not NOT1 (N4287, N4286);
or OR3 (N4288, N4287, N1441, N1593);
and AND3 (N4289, N4288, N1947, N3006);
and AND4 (N4290, N4276, N764, N976, N2041);
nor NOR3 (N4291, N4264, N3660, N1489);
xor XOR2 (N4292, N4282, N3272);
buf BUF1 (N4293, N4290);
not NOT1 (N4294, N4273);
and AND2 (N4295, N4293, N915);
or OR2 (N4296, N4274, N901);
buf BUF1 (N4297, N4283);
nand NAND2 (N4298, N4280, N1740);
not NOT1 (N4299, N4277);
buf BUF1 (N4300, N4285);
or OR4 (N4301, N4292, N2653, N3061, N2976);
nor NOR2 (N4302, N4300, N2909);
and AND4 (N4303, N4296, N1601, N4182, N1206);
nor NOR4 (N4304, N4289, N3476, N3737, N1845);
nand NAND2 (N4305, N4291, N4203);
not NOT1 (N4306, N4297);
xor XOR2 (N4307, N4306, N420);
nand NAND4 (N4308, N4304, N869, N3318, N191);
nor NOR4 (N4309, N4307, N2328, N3558, N160);
nor NOR2 (N4310, N4302, N3182);
and AND4 (N4311, N4303, N842, N4207, N2348);
buf BUF1 (N4312, N4311);
and AND4 (N4313, N4299, N1489, N320, N3125);
buf BUF1 (N4314, N4298);
nand NAND4 (N4315, N4301, N2867, N3492, N2826);
and AND2 (N4316, N4313, N2972);
xor XOR2 (N4317, N4305, N1653);
and AND4 (N4318, N4315, N532, N2951, N3153);
nand NAND3 (N4319, N4308, N1808, N967);
or OR4 (N4320, N4316, N845, N166, N2256);
xor XOR2 (N4321, N4318, N2417);
or OR2 (N4322, N4314, N2263);
or OR3 (N4323, N4295, N4161, N2685);
nand NAND4 (N4324, N4322, N1009, N950, N1701);
xor XOR2 (N4325, N4312, N3410);
or OR2 (N4326, N4294, N3326);
buf BUF1 (N4327, N4320);
not NOT1 (N4328, N4326);
or OR2 (N4329, N4324, N1786);
or OR4 (N4330, N4323, N2595, N2305, N2382);
nor NOR3 (N4331, N4327, N548, N2152);
or OR2 (N4332, N4329, N60);
buf BUF1 (N4333, N4309);
xor XOR2 (N4334, N4333, N1541);
not NOT1 (N4335, N4325);
and AND4 (N4336, N4335, N2340, N1712, N3491);
not NOT1 (N4337, N4319);
not NOT1 (N4338, N4337);
and AND2 (N4339, N4331, N1839);
or OR2 (N4340, N4317, N3701);
or OR4 (N4341, N4332, N881, N2126, N3436);
not NOT1 (N4342, N4338);
or OR4 (N4343, N4339, N3771, N2014, N2020);
buf BUF1 (N4344, N4340);
buf BUF1 (N4345, N4343);
not NOT1 (N4346, N4334);
nor NOR4 (N4347, N4345, N2514, N2900, N1066);
or OR4 (N4348, N4336, N4167, N1587, N1498);
and AND3 (N4349, N4321, N1054, N2059);
buf BUF1 (N4350, N4310);
buf BUF1 (N4351, N4348);
xor XOR2 (N4352, N4347, N2237);
nand NAND3 (N4353, N4341, N438, N2535);
nand NAND3 (N4354, N4349, N2817, N147);
or OR2 (N4355, N4352, N2538);
xor XOR2 (N4356, N4355, N2787);
nand NAND3 (N4357, N4351, N1369, N3723);
or OR3 (N4358, N4350, N2228, N1427);
nor NOR3 (N4359, N4357, N2309, N3675);
not NOT1 (N4360, N4353);
not NOT1 (N4361, N4354);
nor NOR4 (N4362, N4358, N2792, N3133, N2046);
buf BUF1 (N4363, N4328);
not NOT1 (N4364, N4359);
xor XOR2 (N4365, N4346, N3223);
nand NAND2 (N4366, N4364, N1021);
or OR3 (N4367, N4365, N1996, N1808);
or OR3 (N4368, N4362, N3746, N2542);
or OR2 (N4369, N4360, N3486);
xor XOR2 (N4370, N4368, N2107);
and AND4 (N4371, N4370, N545, N1842, N4108);
and AND4 (N4372, N4356, N2836, N2491, N4001);
and AND2 (N4373, N4344, N2176);
not NOT1 (N4374, N4363);
xor XOR2 (N4375, N4373, N3807);
not NOT1 (N4376, N4372);
or OR4 (N4377, N4330, N3830, N2869, N2850);
buf BUF1 (N4378, N4374);
xor XOR2 (N4379, N4367, N4099);
and AND3 (N4380, N4378, N1896, N3402);
xor XOR2 (N4381, N4375, N3133);
or OR2 (N4382, N4377, N1595);
xor XOR2 (N4383, N4342, N3050);
not NOT1 (N4384, N4379);
buf BUF1 (N4385, N4381);
not NOT1 (N4386, N4376);
buf BUF1 (N4387, N4384);
and AND4 (N4388, N4366, N4199, N2378, N1528);
nor NOR2 (N4389, N4387, N2174);
xor XOR2 (N4390, N4361, N3448);
not NOT1 (N4391, N4369);
nor NOR4 (N4392, N4388, N3568, N1763, N2186);
or OR3 (N4393, N4385, N1820, N3641);
or OR3 (N4394, N4382, N167, N2463);
xor XOR2 (N4395, N4393, N2899);
or OR4 (N4396, N4394, N1780, N2160, N3022);
buf BUF1 (N4397, N4380);
nor NOR3 (N4398, N4383, N1237, N265);
nor NOR3 (N4399, N4389, N217, N4276);
buf BUF1 (N4400, N4396);
or OR4 (N4401, N4400, N259, N2170, N4238);
nand NAND3 (N4402, N4399, N1077, N1443);
buf BUF1 (N4403, N4401);
and AND2 (N4404, N4398, N1679);
not NOT1 (N4405, N4397);
nand NAND3 (N4406, N4392, N204, N1213);
nor NOR4 (N4407, N4406, N1671, N1425, N1812);
not NOT1 (N4408, N4371);
buf BUF1 (N4409, N4404);
nor NOR3 (N4410, N4405, N2432, N842);
not NOT1 (N4411, N4410);
not NOT1 (N4412, N4407);
not NOT1 (N4413, N4403);
xor XOR2 (N4414, N4411, N4256);
nor NOR2 (N4415, N4386, N3320);
or OR4 (N4416, N4408, N3754, N316, N1503);
or OR2 (N4417, N4415, N4125);
not NOT1 (N4418, N4414);
xor XOR2 (N4419, N4390, N491);
nand NAND3 (N4420, N4402, N2442, N225);
or OR2 (N4421, N4391, N2116);
nor NOR4 (N4422, N4417, N3672, N2630, N1878);
xor XOR2 (N4423, N4418, N3796);
or OR3 (N4424, N4416, N609, N3903);
xor XOR2 (N4425, N4409, N3438);
or OR2 (N4426, N4421, N1921);
or OR2 (N4427, N4419, N2838);
buf BUF1 (N4428, N4427);
nor NOR4 (N4429, N4426, N4351, N3433, N588);
nor NOR2 (N4430, N4412, N517);
nand NAND3 (N4431, N4429, N2603, N3645);
nand NAND3 (N4432, N4395, N2809, N4186);
xor XOR2 (N4433, N4431, N1638);
or OR4 (N4434, N4424, N4181, N1580, N1387);
buf BUF1 (N4435, N4434);
nand NAND4 (N4436, N4425, N1772, N1269, N3655);
nand NAND3 (N4437, N4433, N348, N3125);
not NOT1 (N4438, N4413);
and AND4 (N4439, N4437, N3146, N2325, N4266);
or OR4 (N4440, N4439, N1226, N2058, N847);
xor XOR2 (N4441, N4420, N1740);
or OR4 (N4442, N4423, N3182, N4166, N1623);
not NOT1 (N4443, N4430);
xor XOR2 (N4444, N4422, N1736);
or OR3 (N4445, N4444, N1417, N2533);
nor NOR2 (N4446, N4436, N3912);
xor XOR2 (N4447, N4446, N4126);
nor NOR4 (N4448, N4428, N2835, N1704, N1664);
buf BUF1 (N4449, N4443);
nor NOR2 (N4450, N4449, N1701);
not NOT1 (N4451, N4435);
xor XOR2 (N4452, N4441, N1692);
nor NOR3 (N4453, N4440, N3261, N2143);
nor NOR3 (N4454, N4447, N4180, N2775);
not NOT1 (N4455, N4453);
xor XOR2 (N4456, N4451, N1853);
nand NAND4 (N4457, N4452, N2437, N2208, N4416);
nor NOR3 (N4458, N4448, N3910, N1748);
or OR4 (N4459, N4438, N2312, N3117, N957);
nand NAND3 (N4460, N4455, N1715, N1568);
nor NOR4 (N4461, N4459, N3670, N439, N2218);
nand NAND3 (N4462, N4458, N2263, N3828);
or OR2 (N4463, N4461, N1585);
nand NAND3 (N4464, N4457, N3221, N2719);
xor XOR2 (N4465, N4464, N1265);
and AND4 (N4466, N4463, N3622, N2952, N3207);
nor NOR3 (N4467, N4454, N1552, N4031);
nor NOR2 (N4468, N4460, N3260);
buf BUF1 (N4469, N4465);
nor NOR4 (N4470, N4456, N4233, N1061, N1596);
nand NAND4 (N4471, N4468, N1854, N2999, N3207);
nor NOR3 (N4472, N4469, N2000, N1154);
or OR4 (N4473, N4442, N3912, N1124, N2350);
or OR3 (N4474, N4432, N760, N1551);
xor XOR2 (N4475, N4472, N111);
not NOT1 (N4476, N4471);
buf BUF1 (N4477, N4450);
or OR3 (N4478, N4475, N4128, N929);
nor NOR4 (N4479, N4474, N742, N1396, N506);
buf BUF1 (N4480, N4470);
nand NAND4 (N4481, N4477, N2463, N2824, N3517);
buf BUF1 (N4482, N4476);
xor XOR2 (N4483, N4478, N2064);
and AND2 (N4484, N4480, N1980);
not NOT1 (N4485, N4462);
nor NOR2 (N4486, N4483, N2243);
buf BUF1 (N4487, N4473);
buf BUF1 (N4488, N4484);
not NOT1 (N4489, N4488);
or OR4 (N4490, N4479, N624, N4063, N696);
buf BUF1 (N4491, N4487);
xor XOR2 (N4492, N4481, N849);
or OR2 (N4493, N4445, N874);
not NOT1 (N4494, N4493);
not NOT1 (N4495, N4485);
not NOT1 (N4496, N4466);
or OR4 (N4497, N4489, N1210, N2910, N3480);
xor XOR2 (N4498, N4467, N58);
nor NOR2 (N4499, N4495, N3257);
nor NOR2 (N4500, N4497, N3444);
not NOT1 (N4501, N4500);
nor NOR3 (N4502, N4492, N472, N1586);
nand NAND2 (N4503, N4499, N2649);
nand NAND4 (N4504, N4491, N2752, N1097, N4380);
not NOT1 (N4505, N4498);
buf BUF1 (N4506, N4504);
buf BUF1 (N4507, N4502);
and AND3 (N4508, N4506, N1570, N607);
not NOT1 (N4509, N4503);
or OR4 (N4510, N4501, N1779, N2670, N3153);
and AND2 (N4511, N4508, N3032);
buf BUF1 (N4512, N4511);
buf BUF1 (N4513, N4486);
nand NAND4 (N4514, N4507, N1391, N455, N2885);
nor NOR4 (N4515, N4512, N4149, N2418, N4435);
not NOT1 (N4516, N4515);
or OR4 (N4517, N4514, N661, N644, N1154);
and AND2 (N4518, N4517, N3105);
nor NOR4 (N4519, N4490, N2477, N2220, N2883);
nand NAND3 (N4520, N4516, N3218, N734);
xor XOR2 (N4521, N4505, N1927);
not NOT1 (N4522, N4482);
buf BUF1 (N4523, N4513);
not NOT1 (N4524, N4496);
or OR4 (N4525, N4520, N2600, N2245, N2160);
not NOT1 (N4526, N4523);
nor NOR4 (N4527, N4522, N2312, N2957, N2817);
and AND4 (N4528, N4524, N1507, N4, N3622);
nor NOR3 (N4529, N4518, N3409, N4143);
or OR4 (N4530, N4527, N3208, N7, N4390);
and AND2 (N4531, N4510, N1196);
xor XOR2 (N4532, N4531, N1131);
or OR4 (N4533, N4509, N2137, N4479, N3569);
nand NAND4 (N4534, N4528, N2770, N2877, N1081);
xor XOR2 (N4535, N4533, N187);
xor XOR2 (N4536, N4534, N3985);
xor XOR2 (N4537, N4536, N4338);
nand NAND4 (N4538, N4535, N1452, N3706, N1178);
or OR4 (N4539, N4494, N3812, N2742, N1458);
nor NOR4 (N4540, N4532, N1079, N758, N4512);
and AND3 (N4541, N4519, N198, N4003);
or OR4 (N4542, N4538, N2831, N2175, N2677);
xor XOR2 (N4543, N4530, N1838);
nand NAND2 (N4544, N4541, N1633);
or OR4 (N4545, N4543, N4391, N1836, N3212);
buf BUF1 (N4546, N4542);
and AND3 (N4547, N4544, N1246, N3327);
not NOT1 (N4548, N4540);
buf BUF1 (N4549, N4548);
not NOT1 (N4550, N4549);
not NOT1 (N4551, N4526);
nor NOR3 (N4552, N4547, N2448, N1060);
or OR2 (N4553, N4529, N1857);
or OR3 (N4554, N4552, N1783, N2851);
or OR2 (N4555, N4537, N1087);
and AND4 (N4556, N4521, N4258, N3054, N62);
buf BUF1 (N4557, N4525);
not NOT1 (N4558, N4539);
xor XOR2 (N4559, N4557, N3943);
xor XOR2 (N4560, N4551, N3432);
nand NAND4 (N4561, N4545, N1990, N715, N2723);
nand NAND4 (N4562, N4556, N3076, N461, N871);
nand NAND2 (N4563, N4558, N718);
not NOT1 (N4564, N4546);
xor XOR2 (N4565, N4563, N1276);
and AND4 (N4566, N4561, N1673, N1757, N2932);
nor NOR4 (N4567, N4550, N489, N2976, N2787);
buf BUF1 (N4568, N4567);
buf BUF1 (N4569, N4562);
and AND3 (N4570, N4555, N869, N1906);
xor XOR2 (N4571, N4570, N3762);
and AND4 (N4572, N4564, N3170, N1465, N3740);
nor NOR4 (N4573, N4559, N942, N4360, N2304);
and AND3 (N4574, N4572, N149, N2718);
xor XOR2 (N4575, N4553, N1891);
nor NOR2 (N4576, N4575, N2573);
not NOT1 (N4577, N4566);
nand NAND2 (N4578, N4574, N3286);
and AND2 (N4579, N4577, N2520);
nand NAND4 (N4580, N4568, N2403, N3173, N338);
not NOT1 (N4581, N4578);
not NOT1 (N4582, N4576);
not NOT1 (N4583, N4573);
nand NAND3 (N4584, N4581, N2651, N3123);
and AND3 (N4585, N4583, N3795, N1800);
or OR3 (N4586, N4585, N3659, N704);
nand NAND2 (N4587, N4569, N160);
xor XOR2 (N4588, N4584, N2210);
and AND4 (N4589, N4560, N2601, N4540, N2944);
and AND2 (N4590, N4571, N2304);
nor NOR3 (N4591, N4554, N3263, N2762);
buf BUF1 (N4592, N4579);
not NOT1 (N4593, N4590);
buf BUF1 (N4594, N4592);
buf BUF1 (N4595, N4582);
buf BUF1 (N4596, N4594);
nand NAND3 (N4597, N4586, N3108, N3259);
not NOT1 (N4598, N4589);
or OR3 (N4599, N4597, N2679, N3182);
or OR3 (N4600, N4588, N4184, N1939);
or OR2 (N4601, N4593, N795);
buf BUF1 (N4602, N4601);
not NOT1 (N4603, N4596);
and AND3 (N4604, N4602, N1632, N335);
and AND4 (N4605, N4580, N3283, N682, N1048);
buf BUF1 (N4606, N4587);
buf BUF1 (N4607, N4598);
nor NOR2 (N4608, N4599, N3501);
not NOT1 (N4609, N4565);
buf BUF1 (N4610, N4600);
or OR3 (N4611, N4606, N640, N599);
and AND3 (N4612, N4591, N2573, N3799);
nand NAND2 (N4613, N4595, N132);
xor XOR2 (N4614, N4611, N3847);
and AND2 (N4615, N4603, N3237);
not NOT1 (N4616, N4609);
and AND2 (N4617, N4615, N3138);
and AND2 (N4618, N4614, N1919);
or OR2 (N4619, N4610, N354);
buf BUF1 (N4620, N4616);
not NOT1 (N4621, N4620);
buf BUF1 (N4622, N4604);
or OR2 (N4623, N4608, N3846);
not NOT1 (N4624, N4617);
not NOT1 (N4625, N4612);
xor XOR2 (N4626, N4625, N2218);
buf BUF1 (N4627, N4619);
not NOT1 (N4628, N4607);
or OR3 (N4629, N4624, N209, N2880);
buf BUF1 (N4630, N4618);
or OR4 (N4631, N4628, N470, N252, N2228);
and AND4 (N4632, N4626, N872, N2659, N1961);
and AND4 (N4633, N4630, N606, N555, N1266);
nor NOR3 (N4634, N4621, N1429, N2178);
nand NAND3 (N4635, N4629, N2116, N4035);
not NOT1 (N4636, N4631);
and AND2 (N4637, N4633, N3015);
or OR2 (N4638, N4635, N3196);
or OR3 (N4639, N4638, N2896, N4550);
nand NAND3 (N4640, N4623, N2134, N644);
and AND2 (N4641, N4640, N4534);
nand NAND3 (N4642, N4632, N3039, N2325);
buf BUF1 (N4643, N4637);
nor NOR2 (N4644, N4641, N1435);
not NOT1 (N4645, N4634);
buf BUF1 (N4646, N4613);
buf BUF1 (N4647, N4646);
or OR4 (N4648, N4627, N21, N38, N2039);
nand NAND2 (N4649, N4636, N4566);
xor XOR2 (N4650, N4622, N4246);
xor XOR2 (N4651, N4639, N2555);
not NOT1 (N4652, N4647);
nor NOR3 (N4653, N4643, N1648, N4095);
buf BUF1 (N4654, N4648);
or OR4 (N4655, N4650, N3871, N867, N1994);
nor NOR3 (N4656, N4605, N2870, N2695);
nand NAND3 (N4657, N4653, N1974, N869);
nor NOR4 (N4658, N4656, N3954, N1521, N1659);
or OR4 (N4659, N4645, N509, N2039, N2615);
and AND3 (N4660, N4644, N1053, N3542);
buf BUF1 (N4661, N4651);
xor XOR2 (N4662, N4658, N4193);
xor XOR2 (N4663, N4655, N4092);
not NOT1 (N4664, N4659);
nand NAND4 (N4665, N4649, N705, N58, N2763);
not NOT1 (N4666, N4642);
nor NOR3 (N4667, N4666, N215, N566);
or OR3 (N4668, N4667, N499, N3453);
nor NOR3 (N4669, N4664, N3579, N3158);
nor NOR4 (N4670, N4657, N3118, N3206, N1569);
not NOT1 (N4671, N4665);
xor XOR2 (N4672, N4652, N2135);
buf BUF1 (N4673, N4660);
not NOT1 (N4674, N4654);
not NOT1 (N4675, N4673);
nand NAND3 (N4676, N4671, N3112, N510);
or OR4 (N4677, N4669, N1524, N2652, N1393);
nor NOR2 (N4678, N4674, N4268);
and AND3 (N4679, N4662, N389, N3513);
buf BUF1 (N4680, N4677);
buf BUF1 (N4681, N4680);
buf BUF1 (N4682, N4668);
nor NOR2 (N4683, N4676, N2803);
or OR4 (N4684, N4682, N2916, N3095, N2684);
nand NAND3 (N4685, N4678, N481, N1220);
and AND2 (N4686, N4663, N3350);
not NOT1 (N4687, N4686);
nand NAND2 (N4688, N4685, N1936);
and AND2 (N4689, N4670, N4388);
nor NOR4 (N4690, N4689, N4635, N3396, N3444);
nor NOR4 (N4691, N4690, N4557, N1092, N182);
and AND3 (N4692, N4687, N501, N3007);
and AND2 (N4693, N4661, N607);
nor NOR2 (N4694, N4692, N2061);
xor XOR2 (N4695, N4679, N1166);
nand NAND4 (N4696, N4675, N3688, N3494, N2497);
xor XOR2 (N4697, N4693, N1618);
buf BUF1 (N4698, N4695);
or OR4 (N4699, N4696, N3366, N2495, N2731);
nand NAND3 (N4700, N4691, N3529, N949);
or OR2 (N4701, N4694, N957);
and AND3 (N4702, N4681, N1913, N703);
nand NAND3 (N4703, N4702, N3197, N4066);
buf BUF1 (N4704, N4703);
not NOT1 (N4705, N4697);
xor XOR2 (N4706, N4672, N1558);
nor NOR2 (N4707, N4704, N3273);
not NOT1 (N4708, N4700);
nand NAND2 (N4709, N4701, N2784);
not NOT1 (N4710, N4705);
xor XOR2 (N4711, N4708, N2829);
not NOT1 (N4712, N4684);
or OR4 (N4713, N4709, N3146, N4595, N3777);
not NOT1 (N4714, N4713);
and AND4 (N4715, N4706, N3502, N4159, N3632);
buf BUF1 (N4716, N4712);
and AND4 (N4717, N4698, N4356, N2155, N847);
xor XOR2 (N4718, N4717, N154);
and AND3 (N4719, N4715, N4490, N2015);
and AND2 (N4720, N4707, N949);
or OR2 (N4721, N4688, N2337);
or OR2 (N4722, N4714, N2146);
xor XOR2 (N4723, N4722, N3987);
nand NAND2 (N4724, N4683, N1980);
or OR4 (N4725, N4711, N2979, N240, N469);
buf BUF1 (N4726, N4699);
buf BUF1 (N4727, N4710);
and AND4 (N4728, N4719, N2125, N1365, N4446);
xor XOR2 (N4729, N4716, N1240);
xor XOR2 (N4730, N4723, N2458);
buf BUF1 (N4731, N4728);
nor NOR4 (N4732, N4729, N1954, N3158, N4287);
not NOT1 (N4733, N4727);
nand NAND3 (N4734, N4730, N3837, N3865);
and AND3 (N4735, N4725, N3015, N3828);
not NOT1 (N4736, N4735);
not NOT1 (N4737, N4731);
and AND3 (N4738, N4737, N641, N972);
nor NOR4 (N4739, N4733, N2082, N2633, N3415);
nand NAND2 (N4740, N4718, N1641);
and AND4 (N4741, N4726, N4466, N3498, N2790);
not NOT1 (N4742, N4740);
and AND4 (N4743, N4721, N2877, N3603, N2074);
not NOT1 (N4744, N4732);
buf BUF1 (N4745, N4720);
not NOT1 (N4746, N4743);
xor XOR2 (N4747, N4742, N117);
nor NOR2 (N4748, N4738, N1486);
nand NAND3 (N4749, N4739, N1415, N3898);
and AND2 (N4750, N4745, N2344);
nor NOR3 (N4751, N4724, N1034, N4722);
or OR3 (N4752, N4749, N1565, N1806);
or OR3 (N4753, N4741, N1332, N4582);
nor NOR2 (N4754, N4753, N1533);
nand NAND3 (N4755, N4752, N2588, N3749);
nor NOR3 (N4756, N4750, N3841, N962);
nor NOR2 (N4757, N4748, N1122);
or OR4 (N4758, N4757, N4750, N2869, N253);
nand NAND4 (N4759, N4746, N3103, N3071, N935);
nand NAND3 (N4760, N4756, N2652, N3375);
not NOT1 (N4761, N4734);
or OR3 (N4762, N4754, N4632, N3194);
or OR3 (N4763, N4760, N4603, N3397);
or OR3 (N4764, N4758, N3603, N1083);
buf BUF1 (N4765, N4759);
xor XOR2 (N4766, N4765, N2809);
nor NOR4 (N4767, N4755, N1987, N1399, N1674);
or OR2 (N4768, N4762, N2962);
and AND2 (N4769, N4768, N2338);
or OR4 (N4770, N4751, N3308, N15, N217);
not NOT1 (N4771, N4770);
or OR4 (N4772, N4769, N3669, N661, N4529);
or OR4 (N4773, N4763, N1059, N1836, N4699);
or OR4 (N4774, N4744, N1402, N3373, N1270);
not NOT1 (N4775, N4774);
nor NOR3 (N4776, N4771, N1820, N2086);
not NOT1 (N4777, N4747);
xor XOR2 (N4778, N4772, N1311);
and AND3 (N4779, N4778, N1235, N1772);
nand NAND4 (N4780, N4766, N1426, N1419, N2551);
and AND4 (N4781, N4736, N724, N1039, N2959);
nand NAND3 (N4782, N4764, N1727, N1799);
or OR2 (N4783, N4781, N909);
nor NOR2 (N4784, N4767, N4093);
buf BUF1 (N4785, N4773);
nand NAND3 (N4786, N4780, N3249, N1822);
and AND2 (N4787, N4782, N3284);
xor XOR2 (N4788, N4776, N3743);
and AND4 (N4789, N4761, N3058, N1829, N76);
xor XOR2 (N4790, N4784, N378);
nand NAND3 (N4791, N4789, N2031, N4725);
buf BUF1 (N4792, N4779);
nor NOR2 (N4793, N4787, N233);
nand NAND3 (N4794, N4790, N2233, N4515);
xor XOR2 (N4795, N4791, N2627);
and AND2 (N4796, N4788, N2091);
not NOT1 (N4797, N4796);
and AND3 (N4798, N4786, N4263, N1591);
nand NAND2 (N4799, N4777, N2123);
and AND2 (N4800, N4783, N4433);
nor NOR3 (N4801, N4775, N1316, N3185);
and AND3 (N4802, N4800, N2061, N3151);
not NOT1 (N4803, N4801);
nand NAND4 (N4804, N4797, N190, N4748, N4224);
nor NOR2 (N4805, N4798, N3536);
xor XOR2 (N4806, N4792, N2543);
and AND2 (N4807, N4802, N3505);
buf BUF1 (N4808, N4806);
xor XOR2 (N4809, N4804, N182);
nor NOR3 (N4810, N4795, N4279, N1870);
buf BUF1 (N4811, N4809);
or OR4 (N4812, N4793, N1469, N1283, N578);
or OR3 (N4813, N4807, N1677, N4477);
or OR4 (N4814, N4803, N2635, N3237, N3282);
xor XOR2 (N4815, N4808, N929);
buf BUF1 (N4816, N4814);
nor NOR3 (N4817, N4812, N1499, N4294);
and AND3 (N4818, N4794, N3432, N2601);
xor XOR2 (N4819, N4815, N2076);
and AND3 (N4820, N4811, N1503, N4132);
and AND3 (N4821, N4818, N4578, N1444);
and AND3 (N4822, N4819, N2647, N4345);
nor NOR3 (N4823, N4785, N4421, N3988);
xor XOR2 (N4824, N4822, N1018);
or OR4 (N4825, N4823, N3094, N4467, N2410);
or OR4 (N4826, N4824, N3967, N2450, N2452);
nand NAND4 (N4827, N4799, N4183, N3699, N4065);
nor NOR3 (N4828, N4827, N3284, N498);
not NOT1 (N4829, N4828);
or OR4 (N4830, N4820, N4009, N2534, N1494);
or OR4 (N4831, N4817, N4605, N2997, N2037);
nor NOR4 (N4832, N4816, N3319, N2171, N1308);
buf BUF1 (N4833, N4832);
xor XOR2 (N4834, N4829, N334);
nor NOR4 (N4835, N4831, N3312, N1202, N4011);
and AND2 (N4836, N4825, N522);
or OR2 (N4837, N4821, N1087);
buf BUF1 (N4838, N4805);
xor XOR2 (N4839, N4837, N3418);
not NOT1 (N4840, N4836);
nor NOR4 (N4841, N4813, N461, N1653, N3783);
buf BUF1 (N4842, N4830);
and AND3 (N4843, N4835, N176, N2418);
nor NOR2 (N4844, N4834, N2112);
not NOT1 (N4845, N4833);
nor NOR4 (N4846, N4838, N26, N2225, N2157);
buf BUF1 (N4847, N4844);
nor NOR4 (N4848, N4826, N2730, N4302, N1463);
not NOT1 (N4849, N4843);
xor XOR2 (N4850, N4810, N2953);
xor XOR2 (N4851, N4848, N1356);
buf BUF1 (N4852, N4840);
nand NAND3 (N4853, N4852, N3685, N652);
and AND4 (N4854, N4853, N3374, N1568, N3564);
xor XOR2 (N4855, N4839, N2157);
not NOT1 (N4856, N4845);
and AND4 (N4857, N4851, N2693, N1549, N3162);
and AND2 (N4858, N4841, N1857);
not NOT1 (N4859, N4855);
and AND4 (N4860, N4846, N1950, N893, N4306);
buf BUF1 (N4861, N4847);
nand NAND4 (N4862, N4854, N4101, N1549, N1501);
nor NOR2 (N4863, N4842, N489);
and AND4 (N4864, N4861, N2343, N394, N2916);
or OR2 (N4865, N4849, N3412);
and AND2 (N4866, N4864, N3908);
not NOT1 (N4867, N4850);
buf BUF1 (N4868, N4862);
nand NAND2 (N4869, N4866, N3652);
and AND4 (N4870, N4858, N4816, N4268, N4414);
nor NOR2 (N4871, N4869, N892);
nor NOR3 (N4872, N4868, N140, N3571);
nor NOR2 (N4873, N4871, N2889);
or OR2 (N4874, N4857, N2591);
not NOT1 (N4875, N4856);
and AND2 (N4876, N4873, N2280);
nor NOR4 (N4877, N4874, N3884, N1766, N1658);
and AND4 (N4878, N4876, N866, N1449, N4178);
buf BUF1 (N4879, N4875);
nand NAND2 (N4880, N4863, N4026);
xor XOR2 (N4881, N4860, N1952);
xor XOR2 (N4882, N4867, N2045);
or OR2 (N4883, N4870, N4791);
not NOT1 (N4884, N4859);
not NOT1 (N4885, N4878);
buf BUF1 (N4886, N4882);
not NOT1 (N4887, N4872);
nand NAND4 (N4888, N4881, N2358, N2848, N4638);
and AND4 (N4889, N4865, N1280, N512, N4527);
not NOT1 (N4890, N4887);
not NOT1 (N4891, N4883);
nand NAND4 (N4892, N4886, N4417, N102, N648);
and AND4 (N4893, N4884, N1224, N2881, N209);
buf BUF1 (N4894, N4893);
or OR4 (N4895, N4879, N4357, N937, N3198);
and AND4 (N4896, N4895, N395, N2133, N235);
or OR2 (N4897, N4877, N521);
xor XOR2 (N4898, N4894, N955);
and AND4 (N4899, N4891, N3347, N223, N3765);
not NOT1 (N4900, N4890);
not NOT1 (N4901, N4900);
nand NAND3 (N4902, N4889, N3172, N114);
nor NOR4 (N4903, N4880, N427, N2687, N4398);
nor NOR3 (N4904, N4898, N1137, N3854);
nor NOR4 (N4905, N4903, N4359, N4450, N1656);
not NOT1 (N4906, N4899);
xor XOR2 (N4907, N4897, N4453);
or OR3 (N4908, N4902, N3735, N711);
or OR3 (N4909, N4892, N2543, N29);
nand NAND4 (N4910, N4896, N4242, N450, N1840);
nor NOR2 (N4911, N4910, N1375);
buf BUF1 (N4912, N4885);
buf BUF1 (N4913, N4901);
nand NAND3 (N4914, N4908, N2137, N4818);
nand NAND2 (N4915, N4905, N86);
not NOT1 (N4916, N4907);
nor NOR2 (N4917, N4912, N989);
buf BUF1 (N4918, N4909);
or OR2 (N4919, N4918, N3057);
xor XOR2 (N4920, N4917, N4756);
nor NOR3 (N4921, N4920, N3164, N556);
nor NOR2 (N4922, N4921, N353);
nor NOR4 (N4923, N4888, N1005, N687, N1267);
and AND4 (N4924, N4904, N391, N679, N2768);
and AND2 (N4925, N4906, N4109);
and AND4 (N4926, N4924, N4347, N4367, N3572);
nor NOR3 (N4927, N4926, N2336, N251);
or OR3 (N4928, N4915, N341, N2825);
and AND3 (N4929, N4911, N199, N2567);
and AND2 (N4930, N4922, N4772);
or OR2 (N4931, N4916, N2996);
nand NAND2 (N4932, N4923, N1970);
xor XOR2 (N4933, N4930, N1411);
buf BUF1 (N4934, N4932);
nor NOR2 (N4935, N4925, N958);
buf BUF1 (N4936, N4929);
buf BUF1 (N4937, N4927);
or OR3 (N4938, N4914, N3614, N2491);
xor XOR2 (N4939, N4928, N3800);
nand NAND4 (N4940, N4935, N4643, N1516, N2537);
xor XOR2 (N4941, N4938, N1674);
and AND3 (N4942, N4933, N3575, N1463);
nand NAND2 (N4943, N4913, N1571);
or OR3 (N4944, N4919, N3066, N1497);
not NOT1 (N4945, N4934);
nand NAND3 (N4946, N4944, N4259, N2115);
not NOT1 (N4947, N4931);
and AND3 (N4948, N4942, N764, N44);
or OR4 (N4949, N4941, N3560, N3207, N1579);
and AND4 (N4950, N4940, N4448, N4524, N362);
not NOT1 (N4951, N4943);
and AND3 (N4952, N4936, N347, N161);
not NOT1 (N4953, N4937);
xor XOR2 (N4954, N4949, N4261);
nand NAND2 (N4955, N4952, N3262);
not NOT1 (N4956, N4953);
buf BUF1 (N4957, N4955);
nand NAND4 (N4958, N4954, N4875, N4166, N3984);
nor NOR3 (N4959, N4947, N2190, N61);
nand NAND2 (N4960, N4939, N3219);
or OR2 (N4961, N4957, N3720);
or OR4 (N4962, N4960, N476, N4337, N613);
nor NOR3 (N4963, N4958, N1318, N3777);
xor XOR2 (N4964, N4951, N2896);
and AND2 (N4965, N4962, N4309);
xor XOR2 (N4966, N4961, N3536);
xor XOR2 (N4967, N4959, N387);
or OR3 (N4968, N4967, N4603, N1490);
nand NAND2 (N4969, N4948, N3301);
xor XOR2 (N4970, N4969, N1099);
not NOT1 (N4971, N4970);
xor XOR2 (N4972, N4956, N3047);
nand NAND3 (N4973, N4968, N2290, N4095);
and AND2 (N4974, N4946, N3051);
buf BUF1 (N4975, N4971);
nor NOR2 (N4976, N4975, N2700);
buf BUF1 (N4977, N4974);
buf BUF1 (N4978, N4976);
not NOT1 (N4979, N4973);
nand NAND2 (N4980, N4950, N159);
and AND2 (N4981, N4966, N1258);
and AND4 (N4982, N4977, N544, N1451, N750);
nand NAND4 (N4983, N4979, N4152, N3977, N832);
xor XOR2 (N4984, N4964, N2180);
and AND3 (N4985, N4980, N853, N58);
nand NAND4 (N4986, N4984, N3059, N1904, N1611);
or OR4 (N4987, N4965, N2089, N2596, N1243);
nand NAND4 (N4988, N4978, N3816, N580, N1146);
and AND2 (N4989, N4987, N2897);
not NOT1 (N4990, N4989);
and AND3 (N4991, N4963, N442, N3792);
nor NOR3 (N4992, N4985, N2411, N4898);
nor NOR2 (N4993, N4992, N2328);
buf BUF1 (N4994, N4982);
nor NOR3 (N4995, N4972, N2549, N4612);
nor NOR2 (N4996, N4994, N341);
buf BUF1 (N4997, N4990);
or OR3 (N4998, N4988, N720, N4252);
and AND3 (N4999, N4983, N1537, N3062);
nand NAND4 (N5000, N4995, N813, N778, N55);
and AND2 (N5001, N4981, N1340);
and AND3 (N5002, N4996, N2535, N1085);
nor NOR2 (N5003, N4945, N291);
xor XOR2 (N5004, N4997, N103);
buf BUF1 (N5005, N5002);
and AND4 (N5006, N5003, N3455, N4513, N2254);
and AND4 (N5007, N5005, N125, N287, N4590);
buf BUF1 (N5008, N5004);
buf BUF1 (N5009, N4999);
nor NOR4 (N5010, N5008, N4711, N1792, N1954);
nand NAND3 (N5011, N5006, N4898, N383);
nor NOR4 (N5012, N4991, N596, N68, N187);
nor NOR2 (N5013, N5009, N1707);
nor NOR2 (N5014, N4986, N4981);
and AND3 (N5015, N5010, N4022, N2250);
nand NAND4 (N5016, N4998, N2352, N574, N3719);
buf BUF1 (N5017, N5016);
and AND4 (N5018, N5007, N947, N938, N4339);
and AND4 (N5019, N5001, N765, N401, N4971);
xor XOR2 (N5020, N5013, N4701);
and AND3 (N5021, N5000, N4813, N95);
and AND3 (N5022, N5018, N2966, N1473);
nor NOR2 (N5023, N5021, N705);
nor NOR4 (N5024, N5015, N1011, N2203, N1995);
not NOT1 (N5025, N5014);
not NOT1 (N5026, N5024);
nor NOR4 (N5027, N5023, N1609, N1277, N192);
or OR2 (N5028, N5022, N3493);
xor XOR2 (N5029, N5026, N722);
xor XOR2 (N5030, N5017, N1363);
nand NAND4 (N5031, N5030, N3517, N978, N2600);
nand NAND2 (N5032, N5011, N111);
nand NAND2 (N5033, N5020, N117);
nand NAND3 (N5034, N5032, N2768, N2503);
nor NOR4 (N5035, N5029, N4917, N3919, N3099);
and AND3 (N5036, N5027, N648, N1807);
or OR3 (N5037, N5036, N150, N238);
not NOT1 (N5038, N5033);
nand NAND3 (N5039, N5019, N3819, N4046);
nor NOR3 (N5040, N5038, N2829, N1459);
and AND2 (N5041, N5034, N3559);
buf BUF1 (N5042, N5037);
buf BUF1 (N5043, N5040);
nor NOR3 (N5044, N5031, N3244, N1368);
and AND4 (N5045, N5042, N165, N3237, N3882);
xor XOR2 (N5046, N5012, N3086);
nand NAND2 (N5047, N5045, N4831);
nor NOR4 (N5048, N5043, N2793, N1383, N4902);
not NOT1 (N5049, N5035);
and AND2 (N5050, N5028, N2599);
nor NOR4 (N5051, N4993, N4253, N2849, N2878);
or OR2 (N5052, N5041, N33);
nor NOR3 (N5053, N5025, N3862, N490);
or OR2 (N5054, N5051, N1564);
nand NAND3 (N5055, N5048, N1346, N1961);
not NOT1 (N5056, N5044);
nor NOR4 (N5057, N5050, N1772, N2543, N518);
buf BUF1 (N5058, N5039);
nor NOR3 (N5059, N5054, N3191, N971);
buf BUF1 (N5060, N5056);
and AND2 (N5061, N5046, N2970);
and AND2 (N5062, N5047, N762);
or OR4 (N5063, N5049, N2076, N1125, N3169);
and AND3 (N5064, N5059, N950, N4015);
or OR4 (N5065, N5055, N3822, N3436, N4547);
nor NOR2 (N5066, N5060, N3913);
not NOT1 (N5067, N5064);
nor NOR4 (N5068, N5053, N1263, N1281, N277);
nor NOR2 (N5069, N5067, N1215);
nor NOR2 (N5070, N5052, N2273);
buf BUF1 (N5071, N5063);
not NOT1 (N5072, N5070);
nand NAND4 (N5073, N5065, N4217, N2556, N594);
not NOT1 (N5074, N5061);
nor NOR4 (N5075, N5068, N2661, N2381, N1596);
or OR3 (N5076, N5073, N4187, N4499);
or OR3 (N5077, N5066, N1335, N3698);
buf BUF1 (N5078, N5071);
xor XOR2 (N5079, N5072, N78);
and AND3 (N5080, N5078, N1233, N3783);
nor NOR4 (N5081, N5057, N4484, N4845, N2951);
buf BUF1 (N5082, N5062);
nor NOR3 (N5083, N5058, N4293, N4254);
nor NOR2 (N5084, N5080, N2597);
xor XOR2 (N5085, N5079, N1);
nor NOR3 (N5086, N5083, N555, N4627);
buf BUF1 (N5087, N5082);
nand NAND2 (N5088, N5087, N833);
nand NAND3 (N5089, N5077, N1934, N1943);
and AND3 (N5090, N5069, N788, N2547);
and AND3 (N5091, N5089, N1355, N1912);
buf BUF1 (N5092, N5085);
nor NOR3 (N5093, N5075, N4980, N4354);
nand NAND4 (N5094, N5093, N2484, N2500, N4491);
or OR3 (N5095, N5094, N4390, N3713);
buf BUF1 (N5096, N5092);
xor XOR2 (N5097, N5091, N777);
nand NAND2 (N5098, N5074, N117);
or OR4 (N5099, N5086, N4723, N2013, N2254);
and AND2 (N5100, N5088, N894);
buf BUF1 (N5101, N5098);
or OR4 (N5102, N5100, N1349, N2661, N4417);
nor NOR4 (N5103, N5084, N3528, N2161, N3405);
and AND3 (N5104, N5102, N2462, N1793);
nor NOR4 (N5105, N5103, N212, N4021, N1225);
nand NAND2 (N5106, N5096, N2200);
not NOT1 (N5107, N5081);
or OR2 (N5108, N5107, N618);
nand NAND2 (N5109, N5095, N4279);
nor NOR2 (N5110, N5106, N3748);
buf BUF1 (N5111, N5108);
nand NAND3 (N5112, N5109, N2782, N634);
buf BUF1 (N5113, N5076);
xor XOR2 (N5114, N5105, N2013);
xor XOR2 (N5115, N5101, N897);
not NOT1 (N5116, N5104);
or OR2 (N5117, N5099, N5045);
buf BUF1 (N5118, N5114);
buf BUF1 (N5119, N5118);
xor XOR2 (N5120, N5115, N2275);
nor NOR3 (N5121, N5117, N1922, N245);
not NOT1 (N5122, N5113);
or OR2 (N5123, N5116, N3965);
or OR3 (N5124, N5097, N2134, N4605);
nor NOR4 (N5125, N5122, N4387, N1859, N1379);
buf BUF1 (N5126, N5124);
buf BUF1 (N5127, N5120);
not NOT1 (N5128, N5123);
nor NOR2 (N5129, N5126, N1190);
and AND3 (N5130, N5127, N1964, N517);
and AND4 (N5131, N5119, N1678, N2070, N1394);
not NOT1 (N5132, N5131);
buf BUF1 (N5133, N5121);
xor XOR2 (N5134, N5125, N3207);
not NOT1 (N5135, N5129);
and AND3 (N5136, N5128, N2918, N1501);
xor XOR2 (N5137, N5132, N123);
buf BUF1 (N5138, N5134);
nand NAND4 (N5139, N5138, N4996, N5104, N1896);
not NOT1 (N5140, N5133);
nand NAND2 (N5141, N5090, N3507);
buf BUF1 (N5142, N5137);
nor NOR2 (N5143, N5111, N774);
or OR4 (N5144, N5141, N5014, N4609, N2567);
or OR2 (N5145, N5135, N2986);
or OR2 (N5146, N5139, N1641);
xor XOR2 (N5147, N5146, N4122);
nor NOR2 (N5148, N5136, N4948);
nand NAND2 (N5149, N5148, N2521);
and AND2 (N5150, N5140, N1868);
nor NOR2 (N5151, N5147, N3642);
not NOT1 (N5152, N5151);
buf BUF1 (N5153, N5145);
and AND3 (N5154, N5152, N5034, N3633);
and AND3 (N5155, N5112, N4083, N1300);
xor XOR2 (N5156, N5153, N4654);
and AND3 (N5157, N5155, N238, N821);
nor NOR3 (N5158, N5154, N4026, N3880);
nor NOR3 (N5159, N5110, N3707, N1690);
nand NAND2 (N5160, N5143, N3668);
nor NOR3 (N5161, N5157, N3293, N3758);
nor NOR3 (N5162, N5149, N2199, N740);
nand NAND3 (N5163, N5150, N1972, N3943);
or OR4 (N5164, N5144, N4127, N4263, N1099);
and AND3 (N5165, N5163, N3335, N3172);
buf BUF1 (N5166, N5156);
not NOT1 (N5167, N5160);
nand NAND2 (N5168, N5164, N28);
not NOT1 (N5169, N5162);
or OR4 (N5170, N5158, N3145, N491, N5120);
nand NAND2 (N5171, N5130, N186);
nand NAND2 (N5172, N5169, N3754);
not NOT1 (N5173, N5161);
nand NAND2 (N5174, N5172, N3461);
nand NAND4 (N5175, N5174, N123, N3295, N3364);
nor NOR2 (N5176, N5173, N4768);
and AND3 (N5177, N5167, N2968, N3318);
nor NOR4 (N5178, N5166, N788, N2600, N2379);
and AND3 (N5179, N5170, N2392, N1040);
nand NAND2 (N5180, N5177, N5054);
buf BUF1 (N5181, N5142);
nand NAND2 (N5182, N5178, N4898);
nand NAND3 (N5183, N5181, N2939, N796);
not NOT1 (N5184, N5180);
or OR3 (N5185, N5159, N4523, N2050);
not NOT1 (N5186, N5179);
or OR2 (N5187, N5184, N3376);
nor NOR2 (N5188, N5183, N2003);
nand NAND2 (N5189, N5187, N1026);
buf BUF1 (N5190, N5189);
or OR3 (N5191, N5182, N2626, N2346);
and AND3 (N5192, N5175, N3754, N1045);
nand NAND3 (N5193, N5186, N2253, N124);
xor XOR2 (N5194, N5165, N1504);
or OR2 (N5195, N5171, N3042);
buf BUF1 (N5196, N5195);
buf BUF1 (N5197, N5191);
or OR4 (N5198, N5194, N3616, N2216, N4001);
nor NOR2 (N5199, N5197, N800);
not NOT1 (N5200, N5196);
xor XOR2 (N5201, N5185, N887);
not NOT1 (N5202, N5190);
and AND3 (N5203, N5168, N2695, N3106);
nand NAND2 (N5204, N5200, N4305);
buf BUF1 (N5205, N5192);
buf BUF1 (N5206, N5193);
nor NOR4 (N5207, N5188, N3570, N1852, N4418);
xor XOR2 (N5208, N5176, N4534);
nor NOR3 (N5209, N5208, N905, N1134);
nor NOR3 (N5210, N5204, N4251, N4067);
not NOT1 (N5211, N5205);
xor XOR2 (N5212, N5198, N1127);
nor NOR2 (N5213, N5199, N3879);
buf BUF1 (N5214, N5212);
or OR4 (N5215, N5211, N2396, N4539, N2379);
buf BUF1 (N5216, N5201);
nor NOR4 (N5217, N5207, N1089, N3363, N3223);
and AND4 (N5218, N5213, N2778, N4922, N2517);
or OR4 (N5219, N5214, N4902, N5000, N449);
or OR3 (N5220, N5209, N4201, N3542);
nand NAND2 (N5221, N5220, N2764);
xor XOR2 (N5222, N5217, N1093);
buf BUF1 (N5223, N5210);
nand NAND4 (N5224, N5216, N4821, N3853, N3761);
not NOT1 (N5225, N5215);
and AND2 (N5226, N5223, N2076);
nor NOR4 (N5227, N5222, N2774, N2359, N806);
xor XOR2 (N5228, N5203, N5156);
nand NAND2 (N5229, N5228, N4541);
buf BUF1 (N5230, N5227);
nand NAND4 (N5231, N5206, N3939, N552, N3550);
xor XOR2 (N5232, N5230, N628);
not NOT1 (N5233, N5225);
not NOT1 (N5234, N5202);
nor NOR4 (N5235, N5231, N1414, N3873, N4936);
nor NOR4 (N5236, N5224, N99, N4875, N3982);
or OR3 (N5237, N5229, N682, N5024);
and AND2 (N5238, N5219, N3886);
or OR4 (N5239, N5234, N4333, N5194, N1719);
buf BUF1 (N5240, N5218);
not NOT1 (N5241, N5232);
and AND3 (N5242, N5240, N3943, N225);
and AND4 (N5243, N5226, N753, N4479, N1100);
buf BUF1 (N5244, N5242);
and AND4 (N5245, N5243, N1106, N4442, N1087);
nand NAND4 (N5246, N5238, N3536, N4031, N426);
buf BUF1 (N5247, N5246);
buf BUF1 (N5248, N5237);
xor XOR2 (N5249, N5236, N4896);
buf BUF1 (N5250, N5247);
buf BUF1 (N5251, N5239);
buf BUF1 (N5252, N5244);
or OR4 (N5253, N5248, N1318, N640, N4854);
nand NAND2 (N5254, N5250, N4513);
nor NOR2 (N5255, N5252, N2708);
not NOT1 (N5256, N5255);
buf BUF1 (N5257, N5254);
and AND2 (N5258, N5235, N2785);
or OR2 (N5259, N5245, N3424);
not NOT1 (N5260, N5221);
and AND2 (N5261, N5260, N1292);
buf BUF1 (N5262, N5258);
not NOT1 (N5263, N5253);
xor XOR2 (N5264, N5262, N4090);
or OR3 (N5265, N5233, N4444, N652);
and AND4 (N5266, N5251, N2517, N521, N4506);
nand NAND2 (N5267, N5257, N3961);
not NOT1 (N5268, N5241);
not NOT1 (N5269, N5267);
not NOT1 (N5270, N5263);
xor XOR2 (N5271, N5259, N4967);
or OR2 (N5272, N5261, N42);
not NOT1 (N5273, N5270);
nand NAND2 (N5274, N5272, N1828);
nand NAND2 (N5275, N5256, N5074);
nor NOR2 (N5276, N5273, N4299);
not NOT1 (N5277, N5276);
nor NOR3 (N5278, N5274, N3722, N2149);
xor XOR2 (N5279, N5266, N938);
xor XOR2 (N5280, N5277, N69);
and AND4 (N5281, N5278, N1264, N4635, N3009);
and AND3 (N5282, N5271, N2766, N1462);
buf BUF1 (N5283, N5282);
xor XOR2 (N5284, N5264, N428);
nor NOR2 (N5285, N5275, N619);
nand NAND4 (N5286, N5265, N4028, N318, N4726);
not NOT1 (N5287, N5268);
xor XOR2 (N5288, N5279, N3921);
buf BUF1 (N5289, N5288);
and AND3 (N5290, N5280, N1086, N518);
nand NAND3 (N5291, N5281, N880, N1307);
xor XOR2 (N5292, N5291, N870);
nor NOR2 (N5293, N5284, N2426);
nor NOR2 (N5294, N5283, N3707);
buf BUF1 (N5295, N5286);
nor NOR4 (N5296, N5285, N4245, N1879, N618);
buf BUF1 (N5297, N5287);
xor XOR2 (N5298, N5295, N1074);
xor XOR2 (N5299, N5298, N3696);
buf BUF1 (N5300, N5297);
not NOT1 (N5301, N5290);
nand NAND2 (N5302, N5296, N2581);
nand NAND3 (N5303, N5249, N2107, N4692);
xor XOR2 (N5304, N5302, N3538);
xor XOR2 (N5305, N5289, N3682);
and AND4 (N5306, N5294, N2614, N1694, N4745);
xor XOR2 (N5307, N5293, N2497);
nor NOR4 (N5308, N5305, N2127, N753, N3720);
and AND4 (N5309, N5299, N2978, N2244, N1435);
buf BUF1 (N5310, N5308);
buf BUF1 (N5311, N5304);
nor NOR3 (N5312, N5292, N1725, N3413);
not NOT1 (N5313, N5306);
xor XOR2 (N5314, N5303, N5168);
or OR4 (N5315, N5300, N4961, N274, N1559);
not NOT1 (N5316, N5310);
xor XOR2 (N5317, N5313, N2276);
and AND4 (N5318, N5311, N2460, N5148, N3858);
not NOT1 (N5319, N5318);
and AND2 (N5320, N5269, N3357);
xor XOR2 (N5321, N5312, N3407);
or OR4 (N5322, N5321, N2501, N1057, N5265);
nor NOR3 (N5323, N5301, N4314, N496);
nor NOR2 (N5324, N5307, N3719);
not NOT1 (N5325, N5319);
and AND2 (N5326, N5323, N4734);
or OR4 (N5327, N5322, N4896, N2290, N4680);
nor NOR2 (N5328, N5317, N4608);
not NOT1 (N5329, N5316);
xor XOR2 (N5330, N5325, N4422);
buf BUF1 (N5331, N5314);
nand NAND2 (N5332, N5320, N3192);
xor XOR2 (N5333, N5326, N3079);
and AND4 (N5334, N5324, N1884, N3990, N4557);
xor XOR2 (N5335, N5330, N4861);
buf BUF1 (N5336, N5327);
nor NOR2 (N5337, N5332, N3402);
or OR3 (N5338, N5309, N3505, N4615);
xor XOR2 (N5339, N5334, N1286);
and AND2 (N5340, N5337, N3634);
nand NAND3 (N5341, N5333, N3786, N5056);
buf BUF1 (N5342, N5336);
nand NAND3 (N5343, N5340, N1661, N2537);
nand NAND3 (N5344, N5329, N642, N4958);
nand NAND4 (N5345, N5315, N1264, N827, N1637);
buf BUF1 (N5346, N5331);
nor NOR3 (N5347, N5338, N4559, N4457);
xor XOR2 (N5348, N5339, N3590);
not NOT1 (N5349, N5346);
or OR4 (N5350, N5341, N4312, N2928, N1517);
or OR2 (N5351, N5342, N1114);
not NOT1 (N5352, N5351);
not NOT1 (N5353, N5343);
or OR3 (N5354, N5350, N2467, N513);
not NOT1 (N5355, N5352);
nand NAND4 (N5356, N5344, N1235, N986, N4048);
and AND3 (N5357, N5347, N596, N4948);
nor NOR4 (N5358, N5349, N2668, N4044, N3760);
nand NAND3 (N5359, N5328, N3980, N1852);
nor NOR2 (N5360, N5357, N1083);
xor XOR2 (N5361, N5356, N3493);
xor XOR2 (N5362, N5355, N461);
nand NAND2 (N5363, N5358, N1751);
nand NAND2 (N5364, N5348, N2126);
nor NOR2 (N5365, N5361, N667);
not NOT1 (N5366, N5364);
and AND2 (N5367, N5360, N4416);
not NOT1 (N5368, N5335);
xor XOR2 (N5369, N5368, N2228);
nand NAND2 (N5370, N5367, N4848);
not NOT1 (N5371, N5369);
nor NOR3 (N5372, N5370, N1716, N2365);
xor XOR2 (N5373, N5371, N339);
nor NOR2 (N5374, N5372, N1680);
nor NOR4 (N5375, N5359, N3311, N2048, N3282);
xor XOR2 (N5376, N5375, N4628);
buf BUF1 (N5377, N5353);
nor NOR3 (N5378, N5374, N1515, N2412);
or OR3 (N5379, N5363, N2666, N3684);
and AND3 (N5380, N5345, N3912, N1750);
buf BUF1 (N5381, N5365);
and AND2 (N5382, N5376, N3155);
buf BUF1 (N5383, N5378);
and AND3 (N5384, N5362, N726, N2426);
not NOT1 (N5385, N5379);
not NOT1 (N5386, N5383);
nand NAND4 (N5387, N5373, N4473, N3869, N4255);
nor NOR4 (N5388, N5387, N354, N4724, N5118);
and AND3 (N5389, N5354, N87, N4241);
or OR2 (N5390, N5384, N5162);
or OR4 (N5391, N5389, N3234, N4965, N4794);
buf BUF1 (N5392, N5388);
nand NAND3 (N5393, N5386, N1705, N3785);
nand NAND2 (N5394, N5366, N3823);
or OR4 (N5395, N5391, N3010, N504, N2445);
and AND2 (N5396, N5393, N178);
or OR3 (N5397, N5380, N4695, N2701);
nor NOR3 (N5398, N5395, N4860, N2468);
or OR2 (N5399, N5385, N3742);
and AND3 (N5400, N5382, N3887, N5027);
xor XOR2 (N5401, N5400, N2650);
and AND3 (N5402, N5398, N2602, N3767);
and AND2 (N5403, N5394, N5136);
not NOT1 (N5404, N5397);
or OR2 (N5405, N5390, N3194);
not NOT1 (N5406, N5377);
and AND3 (N5407, N5406, N1097, N55);
and AND4 (N5408, N5399, N2684, N5003, N395);
xor XOR2 (N5409, N5401, N1272);
nor NOR2 (N5410, N5407, N4808);
nor NOR2 (N5411, N5381, N157);
nand NAND4 (N5412, N5405, N1049, N3031, N2049);
nand NAND4 (N5413, N5408, N2558, N3443, N3922);
nor NOR2 (N5414, N5404, N5294);
or OR2 (N5415, N5411, N2668);
not NOT1 (N5416, N5410);
and AND4 (N5417, N5403, N1515, N2323, N2192);
xor XOR2 (N5418, N5415, N3316);
nor NOR3 (N5419, N5417, N2759, N5265);
buf BUF1 (N5420, N5396);
buf BUF1 (N5421, N5409);
buf BUF1 (N5422, N5420);
buf BUF1 (N5423, N5419);
and AND4 (N5424, N5423, N315, N5105, N3375);
buf BUF1 (N5425, N5414);
nor NOR3 (N5426, N5392, N4437, N4014);
nand NAND2 (N5427, N5425, N2100);
xor XOR2 (N5428, N5416, N5187);
buf BUF1 (N5429, N5413);
or OR4 (N5430, N5412, N5084, N1189, N1247);
nand NAND3 (N5431, N5427, N2644, N3294);
nor NOR3 (N5432, N5431, N2236, N981);
not NOT1 (N5433, N5430);
xor XOR2 (N5434, N5424, N854);
xor XOR2 (N5435, N5432, N816);
nor NOR3 (N5436, N5421, N2392, N2551);
and AND2 (N5437, N5426, N375);
xor XOR2 (N5438, N5418, N5348);
and AND4 (N5439, N5438, N2731, N3515, N3018);
not NOT1 (N5440, N5434);
and AND2 (N5441, N5436, N326);
nand NAND3 (N5442, N5433, N1955, N3570);
or OR2 (N5443, N5439, N5063);
and AND2 (N5444, N5442, N5250);
or OR4 (N5445, N5441, N624, N3381, N3989);
nor NOR2 (N5446, N5445, N3484);
buf BUF1 (N5447, N5440);
buf BUF1 (N5448, N5429);
and AND2 (N5449, N5447, N5113);
buf BUF1 (N5450, N5449);
xor XOR2 (N5451, N5443, N2728);
buf BUF1 (N5452, N5437);
buf BUF1 (N5453, N5448);
nand NAND4 (N5454, N5453, N725, N4894, N2080);
nor NOR2 (N5455, N5454, N3015);
buf BUF1 (N5456, N5446);
nand NAND4 (N5457, N5422, N1202, N242, N2231);
xor XOR2 (N5458, N5435, N1192);
not NOT1 (N5459, N5428);
buf BUF1 (N5460, N5456);
or OR4 (N5461, N5452, N1449, N3184, N4712);
buf BUF1 (N5462, N5455);
nor NOR2 (N5463, N5461, N4170);
not NOT1 (N5464, N5402);
not NOT1 (N5465, N5459);
nand NAND3 (N5466, N5457, N4231, N3820);
nand NAND2 (N5467, N5464, N4581);
or OR3 (N5468, N5450, N5132, N4638);
xor XOR2 (N5469, N5463, N897);
nor NOR2 (N5470, N5469, N2621);
buf BUF1 (N5471, N5468);
buf BUF1 (N5472, N5460);
and AND3 (N5473, N5467, N3108, N690);
and AND4 (N5474, N5472, N4288, N3783, N4691);
nand NAND3 (N5475, N5451, N3287, N4630);
and AND3 (N5476, N5444, N5332, N2421);
nor NOR3 (N5477, N5470, N3419, N985);
nand NAND2 (N5478, N5471, N5331);
nor NOR4 (N5479, N5478, N2775, N2801, N4613);
xor XOR2 (N5480, N5466, N339);
or OR3 (N5481, N5476, N831, N2465);
and AND3 (N5482, N5473, N588, N3495);
not NOT1 (N5483, N5477);
nand NAND4 (N5484, N5479, N4916, N2303, N3082);
not NOT1 (N5485, N5474);
or OR3 (N5486, N5480, N3490, N4360);
nand NAND3 (N5487, N5465, N58, N2589);
nand NAND2 (N5488, N5482, N354);
and AND2 (N5489, N5483, N2684);
or OR2 (N5490, N5486, N1153);
nor NOR2 (N5491, N5490, N1619);
not NOT1 (N5492, N5475);
and AND4 (N5493, N5488, N5013, N4090, N4132);
nor NOR4 (N5494, N5487, N1238, N2103, N1060);
buf BUF1 (N5495, N5481);
nand NAND4 (N5496, N5494, N1174, N3937, N3358);
and AND4 (N5497, N5491, N3150, N3361, N3365);
buf BUF1 (N5498, N5485);
xor XOR2 (N5499, N5458, N3612);
buf BUF1 (N5500, N5495);
and AND3 (N5501, N5500, N2133, N4834);
and AND3 (N5502, N5462, N1235, N5305);
and AND4 (N5503, N5496, N1711, N957, N5477);
or OR2 (N5504, N5502, N160);
buf BUF1 (N5505, N5493);
not NOT1 (N5506, N5492);
and AND4 (N5507, N5505, N3886, N4622, N3238);
and AND4 (N5508, N5484, N2816, N642, N913);
nand NAND3 (N5509, N5498, N2643, N3509);
or OR3 (N5510, N5509, N423, N3183);
xor XOR2 (N5511, N5504, N5371);
or OR3 (N5512, N5489, N3003, N3825);
xor XOR2 (N5513, N5501, N4262);
xor XOR2 (N5514, N5503, N5168);
not NOT1 (N5515, N5508);
nand NAND4 (N5516, N5511, N2479, N2552, N4389);
xor XOR2 (N5517, N5515, N1835);
buf BUF1 (N5518, N5517);
buf BUF1 (N5519, N5516);
buf BUF1 (N5520, N5497);
not NOT1 (N5521, N5506);
xor XOR2 (N5522, N5521, N1990);
not NOT1 (N5523, N5499);
not NOT1 (N5524, N5513);
buf BUF1 (N5525, N5512);
xor XOR2 (N5526, N5523, N163);
or OR3 (N5527, N5518, N1413, N2934);
and AND3 (N5528, N5525, N4524, N928);
and AND3 (N5529, N5507, N5355, N1334);
or OR3 (N5530, N5522, N3985, N1725);
and AND2 (N5531, N5519, N1546);
not NOT1 (N5532, N5510);
or OR3 (N5533, N5520, N174, N3834);
and AND3 (N5534, N5530, N524, N4918);
xor XOR2 (N5535, N5532, N2574);
and AND3 (N5536, N5524, N759, N1326);
buf BUF1 (N5537, N5536);
xor XOR2 (N5538, N5526, N310);
nor NOR2 (N5539, N5531, N2700);
not NOT1 (N5540, N5528);
nor NOR2 (N5541, N5535, N4264);
or OR4 (N5542, N5527, N5490, N4791, N2179);
nor NOR3 (N5543, N5534, N450, N4767);
or OR4 (N5544, N5514, N318, N5124, N1314);
not NOT1 (N5545, N5543);
xor XOR2 (N5546, N5533, N4543);
xor XOR2 (N5547, N5541, N297);
and AND4 (N5548, N5529, N925, N2140, N1917);
buf BUF1 (N5549, N5540);
buf BUF1 (N5550, N5549);
not NOT1 (N5551, N5538);
nand NAND4 (N5552, N5545, N1333, N4095, N5542);
xor XOR2 (N5553, N14, N4528);
nand NAND2 (N5554, N5539, N3155);
not NOT1 (N5555, N5550);
and AND4 (N5556, N5552, N960, N316, N3891);
buf BUF1 (N5557, N5548);
xor XOR2 (N5558, N5537, N2125);
not NOT1 (N5559, N5556);
and AND3 (N5560, N5554, N3834, N5142);
xor XOR2 (N5561, N5560, N3034);
and AND2 (N5562, N5547, N3939);
nand NAND4 (N5563, N5562, N3086, N3964, N4518);
xor XOR2 (N5564, N5563, N1908);
not NOT1 (N5565, N5553);
nor NOR3 (N5566, N5564, N1510, N3237);
or OR4 (N5567, N5561, N1159, N749, N3988);
and AND2 (N5568, N5559, N3665);
buf BUF1 (N5569, N5567);
buf BUF1 (N5570, N5546);
not NOT1 (N5571, N5544);
not NOT1 (N5572, N5569);
not NOT1 (N5573, N5557);
xor XOR2 (N5574, N5558, N2853);
xor XOR2 (N5575, N5551, N4811);
buf BUF1 (N5576, N5574);
nor NOR4 (N5577, N5565, N3529, N1019, N1338);
and AND2 (N5578, N5572, N3506);
not NOT1 (N5579, N5566);
buf BUF1 (N5580, N5571);
xor XOR2 (N5581, N5573, N5318);
nor NOR4 (N5582, N5581, N4192, N490, N2820);
nand NAND4 (N5583, N5582, N2547, N58, N2770);
or OR2 (N5584, N5577, N5274);
nor NOR2 (N5585, N5583, N4917);
xor XOR2 (N5586, N5584, N901);
buf BUF1 (N5587, N5579);
and AND4 (N5588, N5587, N1397, N4577, N2191);
buf BUF1 (N5589, N5578);
nor NOR3 (N5590, N5589, N1908, N1534);
nand NAND4 (N5591, N5588, N5155, N2874, N4291);
nand NAND3 (N5592, N5570, N5310, N2828);
buf BUF1 (N5593, N5568);
and AND3 (N5594, N5590, N4308, N1815);
nand NAND2 (N5595, N5580, N567);
or OR3 (N5596, N5591, N3818, N1289);
and AND2 (N5597, N5586, N3529);
not NOT1 (N5598, N5595);
nand NAND3 (N5599, N5593, N2445, N3210);
not NOT1 (N5600, N5592);
nand NAND3 (N5601, N5598, N4101, N2556);
and AND2 (N5602, N5555, N5303);
and AND2 (N5603, N5576, N257);
not NOT1 (N5604, N5585);
xor XOR2 (N5605, N5602, N915);
and AND2 (N5606, N5600, N2390);
not NOT1 (N5607, N5604);
or OR3 (N5608, N5605, N209, N4540);
or OR3 (N5609, N5603, N4344, N610);
buf BUF1 (N5610, N5601);
nand NAND3 (N5611, N5607, N3002, N2582);
or OR4 (N5612, N5610, N1501, N2618, N4190);
not NOT1 (N5613, N5611);
not NOT1 (N5614, N5613);
and AND4 (N5615, N5599, N4402, N2533, N3056);
buf BUF1 (N5616, N5606);
nand NAND3 (N5617, N5608, N2969, N2352);
xor XOR2 (N5618, N5575, N4489);
xor XOR2 (N5619, N5617, N527);
not NOT1 (N5620, N5618);
xor XOR2 (N5621, N5615, N1583);
xor XOR2 (N5622, N5612, N2294);
or OR4 (N5623, N5597, N1242, N2191, N4507);
nor NOR4 (N5624, N5609, N589, N1978, N5394);
and AND4 (N5625, N5594, N1919, N4772, N1462);
not NOT1 (N5626, N5623);
and AND3 (N5627, N5625, N320, N1108);
nor NOR4 (N5628, N5619, N791, N1620, N1151);
buf BUF1 (N5629, N5622);
xor XOR2 (N5630, N5628, N873);
nand NAND2 (N5631, N5626, N4502);
not NOT1 (N5632, N5630);
nor NOR3 (N5633, N5624, N5293, N1041);
and AND2 (N5634, N5629, N299);
nor NOR4 (N5635, N5631, N3370, N2646, N2536);
or OR2 (N5636, N5635, N2653);
xor XOR2 (N5637, N5616, N4038);
or OR3 (N5638, N5633, N2975, N4631);
buf BUF1 (N5639, N5614);
or OR4 (N5640, N5637, N1899, N2294, N934);
nand NAND3 (N5641, N5639, N3124, N3945);
buf BUF1 (N5642, N5627);
not NOT1 (N5643, N5634);
xor XOR2 (N5644, N5638, N2960);
xor XOR2 (N5645, N5640, N3077);
not NOT1 (N5646, N5620);
and AND4 (N5647, N5643, N3657, N2681, N3285);
nand NAND2 (N5648, N5645, N1590);
nand NAND2 (N5649, N5646, N4370);
not NOT1 (N5650, N5621);
or OR2 (N5651, N5596, N4439);
nand NAND4 (N5652, N5636, N3203, N5259, N732);
nand NAND3 (N5653, N5644, N3106, N239);
nor NOR4 (N5654, N5649, N2870, N3745, N4332);
nor NOR3 (N5655, N5648, N3166, N3123);
or OR2 (N5656, N5655, N3460);
not NOT1 (N5657, N5641);
buf BUF1 (N5658, N5650);
nand NAND2 (N5659, N5654, N420);
or OR3 (N5660, N5652, N1436, N3320);
not NOT1 (N5661, N5660);
nand NAND2 (N5662, N5653, N1731);
or OR4 (N5663, N5657, N4390, N3282, N2737);
or OR2 (N5664, N5659, N1973);
xor XOR2 (N5665, N5651, N1428);
buf BUF1 (N5666, N5665);
or OR4 (N5667, N5664, N692, N2334, N1563);
xor XOR2 (N5668, N5656, N1018);
nor NOR2 (N5669, N5661, N233);
buf BUF1 (N5670, N5662);
nand NAND3 (N5671, N5670, N1239, N1512);
or OR2 (N5672, N5668, N5176);
nand NAND4 (N5673, N5647, N2396, N3737, N185);
and AND4 (N5674, N5658, N2315, N1130, N1618);
or OR3 (N5675, N5674, N3855, N4588);
nand NAND2 (N5676, N5666, N1005);
and AND3 (N5677, N5671, N1215, N1037);
and AND3 (N5678, N5676, N3138, N4584);
or OR3 (N5679, N5675, N2599, N1793);
nand NAND3 (N5680, N5669, N595, N4055);
buf BUF1 (N5681, N5679);
and AND3 (N5682, N5678, N656, N4487);
nor NOR4 (N5683, N5673, N1766, N2362, N3892);
not NOT1 (N5684, N5677);
nor NOR4 (N5685, N5667, N4941, N2901, N871);
nand NAND4 (N5686, N5683, N211, N2388, N1646);
xor XOR2 (N5687, N5672, N3857);
and AND3 (N5688, N5685, N914, N2077);
nor NOR4 (N5689, N5686, N1455, N4327, N1970);
nand NAND4 (N5690, N5687, N4209, N640, N1120);
or OR3 (N5691, N5688, N113, N1174);
or OR2 (N5692, N5684, N4214);
or OR3 (N5693, N5663, N3677, N602);
and AND3 (N5694, N5632, N5692, N5660);
xor XOR2 (N5695, N367, N3237);
buf BUF1 (N5696, N5682);
and AND2 (N5697, N5693, N4316);
not NOT1 (N5698, N5697);
nor NOR3 (N5699, N5698, N434, N4079);
and AND3 (N5700, N5696, N2950, N1338);
nand NAND4 (N5701, N5695, N2930, N2836, N4910);
and AND3 (N5702, N5691, N1358, N2165);
nand NAND4 (N5703, N5701, N933, N2239, N2329);
nor NOR4 (N5704, N5690, N1228, N1006, N90);
or OR4 (N5705, N5642, N4226, N769, N313);
or OR2 (N5706, N5700, N1891);
not NOT1 (N5707, N5681);
not NOT1 (N5708, N5705);
xor XOR2 (N5709, N5702, N3581);
xor XOR2 (N5710, N5708, N515);
buf BUF1 (N5711, N5694);
nand NAND4 (N5712, N5704, N356, N4240, N1235);
not NOT1 (N5713, N5712);
xor XOR2 (N5714, N5713, N2885);
not NOT1 (N5715, N5710);
nand NAND3 (N5716, N5714, N4002, N4936);
nand NAND2 (N5717, N5716, N4671);
nor NOR4 (N5718, N5680, N101, N4492, N5313);
xor XOR2 (N5719, N5718, N4940);
buf BUF1 (N5720, N5719);
or OR4 (N5721, N5720, N910, N90, N4262);
or OR4 (N5722, N5721, N4381, N4213, N4492);
not NOT1 (N5723, N5717);
nor NOR4 (N5724, N5707, N4101, N4355, N3189);
xor XOR2 (N5725, N5723, N647);
nor NOR4 (N5726, N5711, N2444, N3953, N5315);
not NOT1 (N5727, N5722);
not NOT1 (N5728, N5689);
buf BUF1 (N5729, N5727);
nor NOR2 (N5730, N5725, N3304);
and AND2 (N5731, N5706, N783);
xor XOR2 (N5732, N5703, N5337);
nor NOR3 (N5733, N5715, N450, N2397);
buf BUF1 (N5734, N5728);
nand NAND3 (N5735, N5699, N780, N3534);
xor XOR2 (N5736, N5731, N2576);
or OR4 (N5737, N5734, N5060, N5331, N3270);
and AND3 (N5738, N5724, N1466, N464);
nand NAND4 (N5739, N5737, N5579, N855, N416);
xor XOR2 (N5740, N5729, N1171);
not NOT1 (N5741, N5733);
nor NOR3 (N5742, N5739, N1301, N5737);
nor NOR4 (N5743, N5709, N2966, N1488, N4327);
not NOT1 (N5744, N5735);
and AND4 (N5745, N5736, N848, N2540, N3814);
buf BUF1 (N5746, N5740);
nand NAND2 (N5747, N5741, N4007);
or OR3 (N5748, N5746, N2581, N2099);
and AND4 (N5749, N5738, N3569, N4834, N5519);
nor NOR2 (N5750, N5730, N5670);
nor NOR4 (N5751, N5726, N4133, N5344, N4579);
nand NAND4 (N5752, N5732, N1929, N4466, N553);
and AND2 (N5753, N5742, N2911);
buf BUF1 (N5754, N5743);
buf BUF1 (N5755, N5744);
xor XOR2 (N5756, N5753, N2939);
and AND2 (N5757, N5754, N342);
not NOT1 (N5758, N5752);
and AND4 (N5759, N5751, N1476, N588, N4815);
not NOT1 (N5760, N5757);
or OR3 (N5761, N5747, N958, N2484);
nand NAND3 (N5762, N5760, N1376, N2634);
or OR4 (N5763, N5755, N5201, N1387, N5203);
or OR4 (N5764, N5749, N4716, N3257, N3082);
xor XOR2 (N5765, N5763, N4608);
not NOT1 (N5766, N5745);
nand NAND3 (N5767, N5750, N1809, N5516);
not NOT1 (N5768, N5767);
buf BUF1 (N5769, N5762);
xor XOR2 (N5770, N5765, N5496);
and AND3 (N5771, N5756, N1559, N1846);
buf BUF1 (N5772, N5768);
and AND4 (N5773, N5771, N3658, N3089, N4455);
or OR2 (N5774, N5761, N4622);
or OR3 (N5775, N5758, N2198, N2692);
xor XOR2 (N5776, N5769, N2102);
or OR3 (N5777, N5772, N4048, N5346);
buf BUF1 (N5778, N5777);
nand NAND2 (N5779, N5759, N1855);
nor NOR3 (N5780, N5766, N3378, N1935);
not NOT1 (N5781, N5775);
xor XOR2 (N5782, N5748, N3781);
nor NOR2 (N5783, N5781, N664);
nand NAND4 (N5784, N5778, N2873, N5704, N1684);
or OR3 (N5785, N5784, N1891, N1914);
buf BUF1 (N5786, N5779);
not NOT1 (N5787, N5780);
nand NAND3 (N5788, N5774, N3575, N3501);
nand NAND4 (N5789, N5776, N5215, N3328, N184);
nor NOR3 (N5790, N5773, N4759, N4936);
nand NAND4 (N5791, N5786, N561, N4081, N4183);
not NOT1 (N5792, N5783);
and AND4 (N5793, N5788, N1814, N3334, N5003);
buf BUF1 (N5794, N5770);
not NOT1 (N5795, N5790);
and AND3 (N5796, N5787, N1019, N3632);
nor NOR4 (N5797, N5782, N3484, N3097, N4792);
xor XOR2 (N5798, N5793, N5654);
nand NAND2 (N5799, N5785, N2762);
xor XOR2 (N5800, N5799, N5730);
nand NAND3 (N5801, N5764, N610, N5771);
nor NOR3 (N5802, N5791, N2198, N4858);
and AND2 (N5803, N5792, N5086);
buf BUF1 (N5804, N5789);
or OR2 (N5805, N5801, N3509);
nand NAND2 (N5806, N5797, N955);
xor XOR2 (N5807, N5794, N3446);
or OR3 (N5808, N5804, N4683, N5463);
xor XOR2 (N5809, N5802, N4428);
and AND2 (N5810, N5809, N5026);
and AND4 (N5811, N5803, N1270, N461, N679);
and AND2 (N5812, N5798, N5267);
xor XOR2 (N5813, N5808, N5394);
or OR3 (N5814, N5810, N969, N5315);
and AND2 (N5815, N5811, N2476);
and AND4 (N5816, N5806, N3631, N4481, N5324);
and AND4 (N5817, N5807, N3234, N3925, N4269);
not NOT1 (N5818, N5795);
xor XOR2 (N5819, N5814, N5415);
nor NOR4 (N5820, N5819, N3816, N303, N45);
nor NOR2 (N5821, N5818, N1367);
and AND2 (N5822, N5812, N5427);
nor NOR4 (N5823, N5805, N4486, N3675, N3172);
not NOT1 (N5824, N5796);
buf BUF1 (N5825, N5800);
xor XOR2 (N5826, N5821, N3758);
xor XOR2 (N5827, N5820, N81);
nand NAND2 (N5828, N5822, N3186);
nor NOR4 (N5829, N5826, N4513, N5394, N3501);
not NOT1 (N5830, N5813);
not NOT1 (N5831, N5823);
nor NOR4 (N5832, N5824, N3201, N3330, N5641);
nor NOR3 (N5833, N5825, N3748, N1831);
buf BUF1 (N5834, N5829);
buf BUF1 (N5835, N5817);
nand NAND4 (N5836, N5833, N1792, N1739, N1574);
xor XOR2 (N5837, N5816, N2303);
not NOT1 (N5838, N5830);
not NOT1 (N5839, N5834);
not NOT1 (N5840, N5835);
nand NAND3 (N5841, N5831, N4135, N1971);
and AND3 (N5842, N5827, N306, N293);
and AND4 (N5843, N5842, N1992, N2050, N5317);
and AND3 (N5844, N5838, N1961, N37);
xor XOR2 (N5845, N5828, N448);
xor XOR2 (N5846, N5832, N2401);
not NOT1 (N5847, N5841);
or OR3 (N5848, N5844, N4020, N1109);
buf BUF1 (N5849, N5836);
or OR2 (N5850, N5837, N5386);
or OR3 (N5851, N5847, N4284, N1259);
not NOT1 (N5852, N5850);
and AND4 (N5853, N5845, N1765, N3440, N4514);
not NOT1 (N5854, N5839);
and AND4 (N5855, N5843, N5800, N2144, N5514);
and AND2 (N5856, N5848, N1998);
nor NOR2 (N5857, N5840, N2088);
buf BUF1 (N5858, N5856);
buf BUF1 (N5859, N5855);
or OR3 (N5860, N5815, N4496, N6);
and AND4 (N5861, N5860, N2499, N565, N393);
buf BUF1 (N5862, N5857);
xor XOR2 (N5863, N5854, N2611);
buf BUF1 (N5864, N5846);
nor NOR3 (N5865, N5864, N4552, N4234);
not NOT1 (N5866, N5859);
buf BUF1 (N5867, N5862);
or OR3 (N5868, N5853, N1513, N5139);
buf BUF1 (N5869, N5867);
not NOT1 (N5870, N5851);
xor XOR2 (N5871, N5849, N1799);
or OR2 (N5872, N5870, N2767);
nand NAND3 (N5873, N5872, N5688, N1935);
nand NAND2 (N5874, N5858, N4679);
or OR3 (N5875, N5874, N2430, N2291);
xor XOR2 (N5876, N5852, N5824);
buf BUF1 (N5877, N5876);
nand NAND4 (N5878, N5868, N5295, N3233, N3372);
xor XOR2 (N5879, N5877, N351);
not NOT1 (N5880, N5875);
not NOT1 (N5881, N5879);
not NOT1 (N5882, N5863);
and AND2 (N5883, N5861, N2161);
buf BUF1 (N5884, N5869);
buf BUF1 (N5885, N5873);
buf BUF1 (N5886, N5866);
xor XOR2 (N5887, N5878, N5219);
nand NAND3 (N5888, N5871, N1183, N2991);
and AND3 (N5889, N5865, N938, N3848);
not NOT1 (N5890, N5886);
nor NOR4 (N5891, N5880, N2728, N3972, N2804);
nand NAND2 (N5892, N5890, N1751);
nor NOR4 (N5893, N5892, N5083, N1787, N13);
buf BUF1 (N5894, N5882);
and AND3 (N5895, N5889, N4427, N4619);
xor XOR2 (N5896, N5884, N4389);
nor NOR3 (N5897, N5893, N152, N293);
not NOT1 (N5898, N5891);
xor XOR2 (N5899, N5887, N589);
not NOT1 (N5900, N5888);
nand NAND3 (N5901, N5897, N600, N1829);
and AND3 (N5902, N5895, N35, N336);
nand NAND4 (N5903, N5899, N231, N3297, N254);
nand NAND4 (N5904, N5901, N541, N3853, N4366);
and AND4 (N5905, N5883, N5703, N4783, N4448);
xor XOR2 (N5906, N5905, N2082);
xor XOR2 (N5907, N5885, N866);
nand NAND4 (N5908, N5903, N4870, N3718, N5345);
not NOT1 (N5909, N5896);
and AND3 (N5910, N5881, N4370, N4960);
not NOT1 (N5911, N5909);
and AND4 (N5912, N5908, N5632, N671, N2503);
xor XOR2 (N5913, N5910, N1237);
not NOT1 (N5914, N5906);
nor NOR3 (N5915, N5911, N2112, N5745);
buf BUF1 (N5916, N5915);
buf BUF1 (N5917, N5898);
not NOT1 (N5918, N5917);
xor XOR2 (N5919, N5916, N463);
or OR4 (N5920, N5918, N115, N4837, N1328);
xor XOR2 (N5921, N5913, N2788);
nor NOR2 (N5922, N5902, N5002);
and AND2 (N5923, N5922, N2107);
buf BUF1 (N5924, N5923);
nand NAND2 (N5925, N5907, N5823);
nand NAND2 (N5926, N5921, N1298);
nand NAND2 (N5927, N5925, N2118);
and AND3 (N5928, N5900, N1650, N5443);
and AND2 (N5929, N5928, N3253);
not NOT1 (N5930, N5919);
xor XOR2 (N5931, N5920, N5308);
nand NAND3 (N5932, N5894, N4035, N1101);
xor XOR2 (N5933, N5932, N2141);
xor XOR2 (N5934, N5904, N5139);
or OR3 (N5935, N5926, N5546, N3683);
buf BUF1 (N5936, N5929);
not NOT1 (N5937, N5924);
nor NOR4 (N5938, N5937, N2377, N721, N122);
or OR3 (N5939, N5930, N670, N1656);
not NOT1 (N5940, N5939);
buf BUF1 (N5941, N5914);
not NOT1 (N5942, N5941);
not NOT1 (N5943, N5938);
and AND2 (N5944, N5940, N2361);
and AND3 (N5945, N5931, N4048, N4941);
xor XOR2 (N5946, N5936, N1367);
and AND3 (N5947, N5927, N2606, N1016);
xor XOR2 (N5948, N5912, N1582);
buf BUF1 (N5949, N5948);
xor XOR2 (N5950, N5935, N1356);
nand NAND3 (N5951, N5934, N4994, N14);
buf BUF1 (N5952, N5944);
buf BUF1 (N5953, N5952);
or OR4 (N5954, N5945, N5276, N5074, N5048);
or OR4 (N5955, N5951, N5906, N2421, N1224);
nor NOR3 (N5956, N5950, N1341, N4269);
nand NAND3 (N5957, N5954, N4803, N1851);
or OR4 (N5958, N5947, N3325, N1747, N5276);
nand NAND3 (N5959, N5949, N1989, N245);
nand NAND4 (N5960, N5959, N2595, N742, N3537);
xor XOR2 (N5961, N5957, N3175);
buf BUF1 (N5962, N5956);
or OR2 (N5963, N5955, N5071);
buf BUF1 (N5964, N5943);
or OR3 (N5965, N5962, N3086, N1030);
nand NAND2 (N5966, N5953, N3165);
xor XOR2 (N5967, N5965, N5603);
and AND3 (N5968, N5961, N889, N1376);
nand NAND4 (N5969, N5960, N4054, N5446, N3982);
and AND2 (N5970, N5963, N2886);
and AND2 (N5971, N5933, N3048);
and AND4 (N5972, N5969, N3056, N5929, N5482);
nor NOR4 (N5973, N5966, N599, N5940, N4649);
or OR2 (N5974, N5942, N1697);
nor NOR2 (N5975, N5973, N5895);
nand NAND2 (N5976, N5971, N731);
xor XOR2 (N5977, N5968, N1391);
or OR4 (N5978, N5974, N1239, N1549, N5229);
and AND3 (N5979, N5975, N969, N4525);
nand NAND3 (N5980, N5970, N5639, N5677);
xor XOR2 (N5981, N5980, N4107);
and AND3 (N5982, N5946, N2820, N3373);
nand NAND4 (N5983, N5958, N5446, N1317, N4398);
and AND3 (N5984, N5977, N4141, N2177);
and AND3 (N5985, N5981, N3826, N2228);
nand NAND2 (N5986, N5967, N1030);
nor NOR4 (N5987, N5983, N1746, N739, N1402);
xor XOR2 (N5988, N5976, N864);
not NOT1 (N5989, N5982);
buf BUF1 (N5990, N5985);
or OR4 (N5991, N5989, N1155, N309, N4492);
nand NAND3 (N5992, N5990, N4120, N410);
nand NAND2 (N5993, N5988, N3198);
buf BUF1 (N5994, N5972);
or OR4 (N5995, N5987, N1704, N3426, N1192);
nand NAND3 (N5996, N5978, N4769, N1140);
or OR3 (N5997, N5994, N2867, N977);
nand NAND3 (N5998, N5996, N3308, N4125);
buf BUF1 (N5999, N5991);
or OR3 (N6000, N5979, N2554, N4991);
not NOT1 (N6001, N5984);
nand NAND4 (N6002, N5997, N4755, N866, N2192);
not NOT1 (N6003, N5999);
buf BUF1 (N6004, N6003);
nor NOR3 (N6005, N5986, N4272, N1154);
nor NOR3 (N6006, N6004, N2675, N4055);
nor NOR3 (N6007, N6002, N970, N1357);
nor NOR3 (N6008, N6006, N1085, N101);
or OR2 (N6009, N5993, N2618);
nand NAND3 (N6010, N6009, N550, N4985);
or OR2 (N6011, N5992, N1328);
nor NOR4 (N6012, N5998, N1964, N613, N4273);
or OR4 (N6013, N6007, N2897, N5308, N4849);
nor NOR3 (N6014, N6001, N4781, N3168);
nand NAND3 (N6015, N6000, N5068, N1187);
buf BUF1 (N6016, N6013);
xor XOR2 (N6017, N6016, N4907);
and AND2 (N6018, N6008, N4890);
not NOT1 (N6019, N6015);
not NOT1 (N6020, N6014);
nor NOR4 (N6021, N6020, N5676, N2019, N1937);
xor XOR2 (N6022, N6017, N4961);
not NOT1 (N6023, N6005);
and AND4 (N6024, N5995, N5025, N789, N469);
xor XOR2 (N6025, N6018, N1798);
nor NOR2 (N6026, N5964, N4290);
or OR4 (N6027, N6026, N697, N530, N3106);
xor XOR2 (N6028, N6023, N5683);
nor NOR3 (N6029, N6022, N4110, N1028);
nand NAND3 (N6030, N6027, N2276, N4603);
not NOT1 (N6031, N6024);
xor XOR2 (N6032, N6029, N2894);
not NOT1 (N6033, N6019);
not NOT1 (N6034, N6033);
and AND4 (N6035, N6032, N4282, N1905, N2886);
or OR4 (N6036, N6011, N1391, N4805, N5842);
or OR2 (N6037, N6021, N2280);
or OR3 (N6038, N6037, N2865, N4260);
nand NAND4 (N6039, N6034, N3776, N4696, N1918);
nor NOR2 (N6040, N6010, N3271);
not NOT1 (N6041, N6031);
not NOT1 (N6042, N6041);
and AND3 (N6043, N6038, N3585, N3165);
not NOT1 (N6044, N6040);
nor NOR4 (N6045, N6012, N1544, N5849, N3107);
nand NAND3 (N6046, N6045, N4785, N1411);
and AND4 (N6047, N6044, N747, N3237, N2187);
not NOT1 (N6048, N6047);
xor XOR2 (N6049, N6042, N5380);
nand NAND3 (N6050, N6039, N3311, N2593);
nor NOR4 (N6051, N6028, N80, N2688, N2239);
not NOT1 (N6052, N6051);
nand NAND4 (N6053, N6049, N4991, N5363, N3633);
xor XOR2 (N6054, N6053, N3984);
nand NAND3 (N6055, N6048, N2193, N4607);
xor XOR2 (N6056, N6035, N5865);
and AND3 (N6057, N6055, N4369, N5642);
or OR4 (N6058, N6043, N3811, N2629, N1328);
and AND3 (N6059, N6052, N2624, N5495);
and AND2 (N6060, N6046, N4828);
and AND3 (N6061, N6054, N265, N4164);
nor NOR2 (N6062, N6036, N3274);
not NOT1 (N6063, N6056);
nor NOR4 (N6064, N6062, N5018, N5608, N358);
or OR4 (N6065, N6058, N2819, N1400, N2958);
or OR3 (N6066, N6030, N4182, N5348);
and AND2 (N6067, N6059, N3490);
and AND2 (N6068, N6064, N2621);
xor XOR2 (N6069, N6063, N2328);
or OR2 (N6070, N6068, N254);
and AND2 (N6071, N6066, N3772);
not NOT1 (N6072, N6057);
buf BUF1 (N6073, N6065);
or OR4 (N6074, N6025, N2456, N2983, N1494);
buf BUF1 (N6075, N6061);
and AND4 (N6076, N6067, N3791, N4631, N5353);
or OR3 (N6077, N6050, N3831, N3630);
or OR2 (N6078, N6077, N4537);
and AND3 (N6079, N6074, N1893, N2856);
buf BUF1 (N6080, N6069);
nand NAND4 (N6081, N6072, N2581, N2135, N4996);
nor NOR4 (N6082, N6073, N5412, N5160, N3744);
nand NAND2 (N6083, N6075, N4411);
and AND2 (N6084, N6080, N3194);
xor XOR2 (N6085, N6084, N3583);
xor XOR2 (N6086, N6079, N1987);
nand NAND4 (N6087, N6076, N5680, N5983, N4933);
nand NAND3 (N6088, N6071, N1423, N5511);
buf BUF1 (N6089, N6085);
xor XOR2 (N6090, N6086, N3539);
nand NAND2 (N6091, N6088, N5975);
or OR2 (N6092, N6090, N5312);
buf BUF1 (N6093, N6092);
and AND2 (N6094, N6060, N2968);
nand NAND4 (N6095, N6094, N5990, N2769, N4102);
nor NOR2 (N6096, N6089, N1199);
nor NOR3 (N6097, N6095, N2127, N3243);
nand NAND3 (N6098, N6093, N4431, N3550);
buf BUF1 (N6099, N6083);
xor XOR2 (N6100, N6078, N3629);
and AND4 (N6101, N6096, N3425, N3891, N4968);
not NOT1 (N6102, N6070);
nand NAND2 (N6103, N6099, N4003);
xor XOR2 (N6104, N6082, N5387);
nand NAND3 (N6105, N6102, N437, N5463);
nor NOR3 (N6106, N6098, N3953, N2590);
and AND2 (N6107, N6100, N4129);
or OR3 (N6108, N6087, N2063, N1229);
or OR4 (N6109, N6097, N1655, N5783, N2548);
xor XOR2 (N6110, N6101, N2082);
and AND4 (N6111, N6110, N3986, N1365, N2823);
xor XOR2 (N6112, N6081, N5224);
nand NAND3 (N6113, N6105, N3951, N5929);
not NOT1 (N6114, N6109);
xor XOR2 (N6115, N6113, N5280);
nand NAND3 (N6116, N6103, N1743, N5272);
buf BUF1 (N6117, N6115);
or OR3 (N6118, N6111, N4747, N4723);
buf BUF1 (N6119, N6091);
nor NOR2 (N6120, N6119, N3766);
nand NAND4 (N6121, N6112, N1281, N5552, N3998);
buf BUF1 (N6122, N6118);
xor XOR2 (N6123, N6120, N6054);
or OR4 (N6124, N6122, N6114, N2034, N1243);
and AND3 (N6125, N1165, N4268, N4219);
and AND3 (N6126, N6107, N4323, N5589);
or OR3 (N6127, N6108, N4512, N1894);
not NOT1 (N6128, N6117);
not NOT1 (N6129, N6116);
xor XOR2 (N6130, N6121, N2279);
nor NOR2 (N6131, N6125, N3130);
and AND4 (N6132, N6127, N2087, N3410, N4395);
nand NAND4 (N6133, N6132, N1701, N3428, N4909);
nor NOR4 (N6134, N6104, N980, N4863, N2116);
or OR4 (N6135, N6106, N331, N401, N5478);
xor XOR2 (N6136, N6123, N854);
buf BUF1 (N6137, N6135);
and AND2 (N6138, N6130, N3033);
nand NAND4 (N6139, N6136, N5272, N3356, N1187);
xor XOR2 (N6140, N6139, N2505);
or OR2 (N6141, N6124, N1721);
and AND4 (N6142, N6140, N514, N3009, N961);
buf BUF1 (N6143, N6134);
and AND2 (N6144, N6142, N886);
nor NOR4 (N6145, N6138, N5305, N5923, N4110);
nor NOR3 (N6146, N6141, N3385, N2543);
buf BUF1 (N6147, N6131);
xor XOR2 (N6148, N6144, N2036);
xor XOR2 (N6149, N6128, N898);
or OR2 (N6150, N6126, N1968);
nor NOR2 (N6151, N6148, N3226);
nand NAND3 (N6152, N6150, N3291, N2012);
nand NAND2 (N6153, N6137, N1222);
xor XOR2 (N6154, N6149, N4249);
xor XOR2 (N6155, N6129, N4286);
buf BUF1 (N6156, N6143);
and AND2 (N6157, N6145, N1587);
xor XOR2 (N6158, N6154, N3066);
and AND4 (N6159, N6147, N2716, N5542, N4132);
nor NOR4 (N6160, N6133, N6150, N3068, N4105);
or OR2 (N6161, N6158, N2220);
nor NOR2 (N6162, N6161, N1570);
xor XOR2 (N6163, N6155, N5589);
xor XOR2 (N6164, N6153, N5109);
nor NOR3 (N6165, N6157, N2481, N3005);
not NOT1 (N6166, N6146);
not NOT1 (N6167, N6159);
nor NOR3 (N6168, N6164, N1763, N5467);
xor XOR2 (N6169, N6152, N3634);
not NOT1 (N6170, N6168);
xor XOR2 (N6171, N6170, N3267);
nor NOR3 (N6172, N6160, N4798, N5742);
or OR3 (N6173, N6167, N4479, N5991);
nand NAND2 (N6174, N6172, N1104);
buf BUF1 (N6175, N6151);
nor NOR4 (N6176, N6162, N3175, N4331, N1579);
nand NAND4 (N6177, N6165, N3339, N3649, N1065);
nand NAND2 (N6178, N6176, N2272);
xor XOR2 (N6179, N6174, N1443);
and AND2 (N6180, N6169, N3656);
buf BUF1 (N6181, N6163);
xor XOR2 (N6182, N6156, N1467);
nand NAND4 (N6183, N6178, N3917, N6171, N5813);
or OR2 (N6184, N4949, N1687);
and AND4 (N6185, N6183, N5634, N4234, N1740);
or OR4 (N6186, N6177, N3550, N4806, N446);
not NOT1 (N6187, N6181);
not NOT1 (N6188, N6175);
nand NAND4 (N6189, N6186, N48, N5198, N1826);
or OR2 (N6190, N6185, N5677);
not NOT1 (N6191, N6180);
buf BUF1 (N6192, N6187);
or OR2 (N6193, N6188, N3973);
and AND4 (N6194, N6173, N4902, N2309, N3927);
or OR3 (N6195, N6190, N6024, N2705);
nor NOR2 (N6196, N6182, N3006);
or OR4 (N6197, N6166, N4375, N1456, N2823);
not NOT1 (N6198, N6191);
buf BUF1 (N6199, N6198);
xor XOR2 (N6200, N6196, N1983);
buf BUF1 (N6201, N6199);
nand NAND4 (N6202, N6184, N1980, N4620, N4450);
buf BUF1 (N6203, N6200);
xor XOR2 (N6204, N6197, N552);
nand NAND2 (N6205, N6192, N3781);
or OR3 (N6206, N6193, N401, N1550);
and AND3 (N6207, N6195, N1978, N3719);
nand NAND2 (N6208, N6201, N2986);
and AND3 (N6209, N6204, N1950, N1198);
or OR4 (N6210, N6209, N5807, N2160, N1953);
xor XOR2 (N6211, N6208, N1498);
not NOT1 (N6212, N6210);
and AND2 (N6213, N6189, N54);
and AND3 (N6214, N6179, N2775, N237);
nand NAND2 (N6215, N6212, N3365);
not NOT1 (N6216, N6194);
or OR4 (N6217, N6205, N6095, N1108, N2803);
xor XOR2 (N6218, N6203, N5916);
buf BUF1 (N6219, N6216);
nand NAND2 (N6220, N6218, N4305);
or OR4 (N6221, N6217, N5197, N3671, N876);
xor XOR2 (N6222, N6220, N3611);
buf BUF1 (N6223, N6211);
nand NAND4 (N6224, N6213, N5912, N2542, N908);
nand NAND2 (N6225, N6219, N6103);
nor NOR3 (N6226, N6221, N240, N1476);
nor NOR4 (N6227, N6215, N1705, N6139, N3662);
buf BUF1 (N6228, N6223);
nor NOR4 (N6229, N6222, N5101, N56, N5984);
not NOT1 (N6230, N6225);
not NOT1 (N6231, N6207);
not NOT1 (N6232, N6202);
xor XOR2 (N6233, N6227, N654);
and AND2 (N6234, N6226, N5815);
xor XOR2 (N6235, N6234, N4722);
and AND4 (N6236, N6206, N775, N4291, N2377);
xor XOR2 (N6237, N6229, N2544);
nand NAND2 (N6238, N6224, N64);
not NOT1 (N6239, N6237);
or OR3 (N6240, N6233, N5078, N629);
or OR3 (N6241, N6235, N4425, N4652);
buf BUF1 (N6242, N6228);
buf BUF1 (N6243, N6239);
and AND2 (N6244, N6236, N5850);
buf BUF1 (N6245, N6244);
nand NAND4 (N6246, N6232, N4580, N1578, N5264);
buf BUF1 (N6247, N6246);
not NOT1 (N6248, N6214);
nand NAND4 (N6249, N6245, N5428, N5873, N1765);
or OR3 (N6250, N6238, N2378, N1962);
or OR2 (N6251, N6247, N529);
or OR4 (N6252, N6251, N1818, N1370, N2363);
not NOT1 (N6253, N6248);
buf BUF1 (N6254, N6249);
or OR2 (N6255, N6250, N4185);
nand NAND4 (N6256, N6254, N1671, N5029, N3966);
nor NOR4 (N6257, N6255, N2860, N4389, N4940);
nand NAND2 (N6258, N6241, N5382);
and AND4 (N6259, N6253, N459, N1010, N1925);
buf BUF1 (N6260, N6256);
buf BUF1 (N6261, N6231);
nand NAND2 (N6262, N6230, N2674);
xor XOR2 (N6263, N6240, N1727);
nor NOR4 (N6264, N6260, N2742, N6206, N2941);
nor NOR4 (N6265, N6252, N5708, N2664, N1684);
not NOT1 (N6266, N6243);
buf BUF1 (N6267, N6265);
xor XOR2 (N6268, N6262, N5711);
buf BUF1 (N6269, N6258);
or OR4 (N6270, N6263, N5430, N3194, N4330);
nand NAND2 (N6271, N6267, N3324);
and AND3 (N6272, N6261, N3323, N1340);
and AND2 (N6273, N6269, N770);
not NOT1 (N6274, N6266);
and AND2 (N6275, N6259, N6150);
and AND2 (N6276, N6271, N3625);
or OR3 (N6277, N6276, N5093, N3006);
not NOT1 (N6278, N6268);
nor NOR3 (N6279, N6278, N4630, N5238);
buf BUF1 (N6280, N6273);
xor XOR2 (N6281, N6279, N4635);
xor XOR2 (N6282, N6280, N4491);
buf BUF1 (N6283, N6282);
nand NAND4 (N6284, N6264, N1876, N395, N5015);
and AND3 (N6285, N6281, N4551, N360);
and AND4 (N6286, N6242, N162, N3934, N1217);
nor NOR3 (N6287, N6257, N6227, N3549);
xor XOR2 (N6288, N6272, N4847);
nor NOR3 (N6289, N6284, N1176, N3459);
nand NAND3 (N6290, N6277, N1057, N2260);
xor XOR2 (N6291, N6275, N4412);
nand NAND4 (N6292, N6270, N4152, N2086, N496);
xor XOR2 (N6293, N6285, N5294);
or OR4 (N6294, N6291, N4023, N1482, N4757);
or OR4 (N6295, N6288, N3460, N6167, N3468);
nor NOR2 (N6296, N6287, N5615);
or OR2 (N6297, N6290, N2896);
buf BUF1 (N6298, N6297);
nor NOR2 (N6299, N6296, N2229);
or OR4 (N6300, N6289, N4781, N4901, N5668);
not NOT1 (N6301, N6294);
or OR4 (N6302, N6298, N5510, N3613, N602);
buf BUF1 (N6303, N6274);
or OR2 (N6304, N6299, N2836);
nor NOR3 (N6305, N6301, N645, N1769);
and AND3 (N6306, N6283, N1809, N1719);
xor XOR2 (N6307, N6303, N427);
not NOT1 (N6308, N6295);
and AND4 (N6309, N6307, N1887, N4083, N2721);
nand NAND2 (N6310, N6292, N1701);
nand NAND3 (N6311, N6302, N5756, N2891);
or OR2 (N6312, N6305, N175);
nand NAND2 (N6313, N6309, N911);
not NOT1 (N6314, N6286);
buf BUF1 (N6315, N6313);
or OR2 (N6316, N6304, N3709);
not NOT1 (N6317, N6316);
nand NAND4 (N6318, N6312, N3838, N5887, N2993);
xor XOR2 (N6319, N6308, N1594);
nand NAND4 (N6320, N6317, N4519, N490, N5639);
nor NOR3 (N6321, N6310, N1541, N3475);
not NOT1 (N6322, N6311);
or OR3 (N6323, N6300, N4442, N563);
nand NAND4 (N6324, N6306, N2541, N3880, N1932);
nand NAND3 (N6325, N6319, N2324, N816);
nor NOR2 (N6326, N6322, N1753);
not NOT1 (N6327, N6325);
xor XOR2 (N6328, N6324, N6309);
nor NOR4 (N6329, N6326, N5554, N1900, N1499);
nand NAND4 (N6330, N6321, N2873, N1887, N1221);
nor NOR4 (N6331, N6330, N1312, N2518, N3480);
nor NOR3 (N6332, N6293, N5864, N5310);
not NOT1 (N6333, N6327);
and AND3 (N6334, N6320, N5426, N4688);
xor XOR2 (N6335, N6331, N1417);
not NOT1 (N6336, N6318);
nor NOR4 (N6337, N6314, N3541, N3805, N5496);
not NOT1 (N6338, N6334);
buf BUF1 (N6339, N6328);
buf BUF1 (N6340, N6337);
xor XOR2 (N6341, N6329, N4398);
nor NOR3 (N6342, N6339, N3422, N948);
buf BUF1 (N6343, N6332);
buf BUF1 (N6344, N6315);
xor XOR2 (N6345, N6338, N3142);
and AND2 (N6346, N6343, N3138);
not NOT1 (N6347, N6336);
nor NOR3 (N6348, N6333, N584, N3006);
or OR4 (N6349, N6345, N4707, N762, N3746);
nand NAND2 (N6350, N6348, N5135);
not NOT1 (N6351, N6323);
xor XOR2 (N6352, N6347, N2834);
nor NOR4 (N6353, N6352, N5642, N2261, N677);
buf BUF1 (N6354, N6340);
xor XOR2 (N6355, N6346, N3782);
xor XOR2 (N6356, N6341, N2422);
and AND3 (N6357, N6350, N2443, N3599);
nand NAND3 (N6358, N6356, N108, N1673);
nand NAND3 (N6359, N6355, N4855, N5694);
and AND2 (N6360, N6349, N3450);
nand NAND4 (N6361, N6351, N4382, N4889, N6295);
or OR3 (N6362, N6361, N4772, N6076);
xor XOR2 (N6363, N6344, N1489);
nand NAND3 (N6364, N6362, N1619, N4521);
and AND3 (N6365, N6364, N4825, N1650);
or OR4 (N6366, N6342, N2819, N1236, N4349);
buf BUF1 (N6367, N6360);
xor XOR2 (N6368, N6366, N4939);
buf BUF1 (N6369, N6359);
buf BUF1 (N6370, N6357);
and AND4 (N6371, N6365, N5264, N3476, N5375);
nor NOR4 (N6372, N6368, N23, N855, N5471);
buf BUF1 (N6373, N6353);
nand NAND4 (N6374, N6363, N5327, N1066, N3102);
nand NAND2 (N6375, N6335, N4387);
not NOT1 (N6376, N6354);
nor NOR2 (N6377, N6374, N269);
and AND2 (N6378, N6370, N5780);
buf BUF1 (N6379, N6372);
nor NOR3 (N6380, N6379, N780, N575);
nand NAND4 (N6381, N6375, N3962, N4598, N4145);
not NOT1 (N6382, N6369);
nand NAND4 (N6383, N6358, N2076, N2059, N3552);
nand NAND3 (N6384, N6380, N3109, N4936);
and AND2 (N6385, N6382, N5884);
and AND3 (N6386, N6378, N6281, N1824);
or OR3 (N6387, N6385, N4127, N1640);
xor XOR2 (N6388, N6381, N1499);
nor NOR3 (N6389, N6377, N2280, N1179);
or OR2 (N6390, N6384, N6129);
nor NOR2 (N6391, N6373, N6352);
nor NOR4 (N6392, N6383, N4593, N3591, N178);
not NOT1 (N6393, N6367);
not NOT1 (N6394, N6392);
buf BUF1 (N6395, N6371);
and AND3 (N6396, N6386, N1835, N4623);
nor NOR2 (N6397, N6396, N648);
and AND2 (N6398, N6395, N1280);
nand NAND2 (N6399, N6389, N1119);
nor NOR4 (N6400, N6393, N2289, N2991, N3645);
xor XOR2 (N6401, N6394, N3066);
or OR4 (N6402, N6390, N5308, N827, N2394);
buf BUF1 (N6403, N6399);
and AND3 (N6404, N6391, N1243, N4024);
nor NOR2 (N6405, N6397, N4989);
or OR2 (N6406, N6376, N2946);
and AND3 (N6407, N6405, N3939, N4296);
not NOT1 (N6408, N6407);
or OR4 (N6409, N6403, N2966, N5872, N1283);
buf BUF1 (N6410, N6406);
buf BUF1 (N6411, N6402);
and AND3 (N6412, N6401, N3335, N6192);
xor XOR2 (N6413, N6409, N3393);
and AND2 (N6414, N6387, N3703);
and AND4 (N6415, N6411, N1976, N4947, N3443);
xor XOR2 (N6416, N6408, N5833);
or OR4 (N6417, N6388, N1545, N6401, N4888);
buf BUF1 (N6418, N6412);
nand NAND3 (N6419, N6410, N1550, N2257);
xor XOR2 (N6420, N6418, N347);
nor NOR3 (N6421, N6415, N2366, N5933);
buf BUF1 (N6422, N6417);
nor NOR2 (N6423, N6398, N5915);
and AND2 (N6424, N6419, N4186);
buf BUF1 (N6425, N6422);
nor NOR2 (N6426, N6414, N983);
nand NAND2 (N6427, N6421, N3922);
buf BUF1 (N6428, N6424);
and AND4 (N6429, N6413, N3628, N3725, N5411);
and AND3 (N6430, N6427, N5511, N5945);
nand NAND3 (N6431, N6400, N2554, N3620);
nand NAND3 (N6432, N6428, N2665, N1127);
xor XOR2 (N6433, N6429, N6400);
xor XOR2 (N6434, N6425, N3108);
nor NOR3 (N6435, N6426, N4949, N48);
or OR4 (N6436, N6416, N1216, N4981, N1108);
nor NOR3 (N6437, N6430, N2045, N2047);
and AND4 (N6438, N6436, N4496, N5487, N68);
buf BUF1 (N6439, N6420);
buf BUF1 (N6440, N6431);
and AND4 (N6441, N6439, N3309, N4896, N3829);
and AND4 (N6442, N6437, N1244, N4868, N3038);
nand NAND3 (N6443, N6434, N1171, N4438);
buf BUF1 (N6444, N6423);
not NOT1 (N6445, N6438);
or OR2 (N6446, N6435, N3016);
and AND2 (N6447, N6433, N4924);
buf BUF1 (N6448, N6404);
buf BUF1 (N6449, N6445);
not NOT1 (N6450, N6441);
and AND2 (N6451, N6444, N212);
and AND2 (N6452, N6451, N2951);
nor NOR3 (N6453, N6442, N4124, N942);
buf BUF1 (N6454, N6432);
buf BUF1 (N6455, N6443);
and AND4 (N6456, N6455, N1973, N794, N1085);
nor NOR3 (N6457, N6456, N2753, N1016);
nand NAND2 (N6458, N6452, N2345);
or OR3 (N6459, N6446, N3902, N2949);
xor XOR2 (N6460, N6447, N1586);
or OR2 (N6461, N6458, N1090);
nor NOR4 (N6462, N6460, N4209, N2921, N5180);
or OR4 (N6463, N6461, N1125, N2350, N5986);
buf BUF1 (N6464, N6454);
and AND3 (N6465, N6457, N5101, N4137);
buf BUF1 (N6466, N6459);
or OR4 (N6467, N6464, N4354, N586, N1028);
not NOT1 (N6468, N6467);
xor XOR2 (N6469, N6448, N5745);
not NOT1 (N6470, N6463);
nor NOR4 (N6471, N6469, N6336, N2790, N4129);
nand NAND2 (N6472, N6465, N636);
or OR3 (N6473, N6453, N4564, N5833);
and AND2 (N6474, N6450, N2881);
xor XOR2 (N6475, N6449, N3641);
and AND3 (N6476, N6471, N3466, N5696);
or OR2 (N6477, N6474, N699);
and AND4 (N6478, N6475, N6121, N885, N2930);
nor NOR4 (N6479, N6466, N1398, N5103, N6375);
nor NOR4 (N6480, N6479, N2310, N2110, N4747);
xor XOR2 (N6481, N6440, N4722);
buf BUF1 (N6482, N6470);
nand NAND3 (N6483, N6476, N5481, N592);
or OR3 (N6484, N6473, N6359, N1026);
and AND3 (N6485, N6478, N4228, N4005);
not NOT1 (N6486, N6462);
nand NAND4 (N6487, N6484, N1972, N6084, N5016);
nand NAND3 (N6488, N6477, N883, N1110);
nor NOR4 (N6489, N6480, N5445, N2571, N2856);
xor XOR2 (N6490, N6489, N700);
not NOT1 (N6491, N6486);
or OR3 (N6492, N6488, N3671, N1844);
xor XOR2 (N6493, N6472, N2884);
or OR3 (N6494, N6481, N3634, N2386);
nand NAND3 (N6495, N6492, N2581, N5531);
not NOT1 (N6496, N6495);
and AND3 (N6497, N6493, N3817, N3402);
not NOT1 (N6498, N6482);
nand NAND4 (N6499, N6490, N3142, N5817, N1432);
and AND4 (N6500, N6499, N5615, N4625, N3781);
buf BUF1 (N6501, N6496);
nor NOR4 (N6502, N6500, N2861, N3243, N4630);
xor XOR2 (N6503, N6502, N3431);
or OR2 (N6504, N6503, N4152);
buf BUF1 (N6505, N6491);
nand NAND2 (N6506, N6504, N2741);
or OR2 (N6507, N6487, N307);
nor NOR4 (N6508, N6498, N3746, N6188, N2078);
and AND4 (N6509, N6508, N3113, N4803, N1196);
nor NOR2 (N6510, N6509, N1219);
not NOT1 (N6511, N6483);
buf BUF1 (N6512, N6506);
not NOT1 (N6513, N6511);
or OR4 (N6514, N6497, N2918, N1677, N980);
nor NOR2 (N6515, N6468, N1339);
nor NOR4 (N6516, N6515, N4432, N3347, N5748);
not NOT1 (N6517, N6485);
or OR2 (N6518, N6512, N5738);
and AND2 (N6519, N6507, N3864);
nand NAND3 (N6520, N6505, N3346, N1985);
buf BUF1 (N6521, N6513);
and AND2 (N6522, N6514, N832);
buf BUF1 (N6523, N6510);
nand NAND4 (N6524, N6523, N1665, N4859, N2278);
and AND4 (N6525, N6516, N4201, N2118, N1355);
buf BUF1 (N6526, N6522);
nor NOR2 (N6527, N6501, N704);
nor NOR3 (N6528, N6519, N5010, N2166);
or OR2 (N6529, N6517, N4106);
buf BUF1 (N6530, N6529);
and AND2 (N6531, N6527, N1084);
xor XOR2 (N6532, N6520, N3126);
buf BUF1 (N6533, N6531);
and AND3 (N6534, N6524, N5855, N2521);
buf BUF1 (N6535, N6494);
nor NOR2 (N6536, N6532, N6304);
buf BUF1 (N6537, N6533);
or OR4 (N6538, N6536, N1219, N4639, N2450);
or OR3 (N6539, N6525, N3976, N4941);
buf BUF1 (N6540, N6535);
nor NOR4 (N6541, N6539, N1253, N1555, N3848);
buf BUF1 (N6542, N6526);
nor NOR2 (N6543, N6541, N87);
nor NOR3 (N6544, N6542, N4449, N193);
buf BUF1 (N6545, N6530);
and AND4 (N6546, N6544, N6535, N3143, N3779);
or OR2 (N6547, N6537, N276);
xor XOR2 (N6548, N6540, N3866);
xor XOR2 (N6549, N6534, N2656);
or OR2 (N6550, N6546, N2291);
or OR4 (N6551, N6518, N261, N3270, N1995);
not NOT1 (N6552, N6547);
and AND2 (N6553, N6550, N2757);
nor NOR3 (N6554, N6543, N5057, N1492);
buf BUF1 (N6555, N6549);
buf BUF1 (N6556, N6521);
and AND4 (N6557, N6548, N175, N639, N976);
xor XOR2 (N6558, N6545, N3030);
buf BUF1 (N6559, N6553);
not NOT1 (N6560, N6551);
nand NAND2 (N6561, N6555, N3968);
not NOT1 (N6562, N6558);
and AND4 (N6563, N6556, N5804, N2328, N2707);
nor NOR3 (N6564, N6559, N6207, N6013);
not NOT1 (N6565, N6554);
buf BUF1 (N6566, N6565);
and AND3 (N6567, N6528, N3673, N2505);
not NOT1 (N6568, N6563);
and AND3 (N6569, N6557, N122, N6277);
nor NOR2 (N6570, N6560, N2210);
xor XOR2 (N6571, N6564, N2969);
buf BUF1 (N6572, N6571);
xor XOR2 (N6573, N6572, N2477);
xor XOR2 (N6574, N6538, N2599);
nor NOR3 (N6575, N6566, N4890, N4374);
nand NAND3 (N6576, N6552, N1335, N4006);
buf BUF1 (N6577, N6562);
or OR3 (N6578, N6569, N3734, N125);
not NOT1 (N6579, N6575);
or OR2 (N6580, N6573, N3872);
nor NOR3 (N6581, N6576, N5338, N5709);
nand NAND4 (N6582, N6568, N1666, N2023, N5352);
nor NOR2 (N6583, N6577, N769);
nand NAND4 (N6584, N6570, N6235, N2389, N711);
or OR3 (N6585, N6574, N2129, N5763);
xor XOR2 (N6586, N6584, N2444);
not NOT1 (N6587, N6583);
xor XOR2 (N6588, N6581, N150);
nand NAND4 (N6589, N6586, N3028, N3506, N183);
nor NOR3 (N6590, N6582, N3888, N2798);
or OR4 (N6591, N6579, N2587, N4645, N6275);
buf BUF1 (N6592, N6580);
nand NAND4 (N6593, N6567, N4936, N656, N3576);
and AND3 (N6594, N6587, N912, N4527);
nand NAND2 (N6595, N6591, N2464);
nand NAND3 (N6596, N6594, N268, N2008);
or OR3 (N6597, N6592, N524, N2646);
buf BUF1 (N6598, N6590);
nand NAND4 (N6599, N6585, N526, N4102, N2468);
nor NOR4 (N6600, N6578, N5527, N6119, N2232);
nand NAND4 (N6601, N6593, N1067, N5187, N3869);
or OR3 (N6602, N6598, N5509, N1444);
or OR4 (N6603, N6596, N1735, N3292, N1910);
nor NOR2 (N6604, N6603, N1561);
nor NOR4 (N6605, N6600, N586, N5004, N5056);
xor XOR2 (N6606, N6597, N1156);
nor NOR4 (N6607, N6602, N4531, N4716, N5603);
and AND3 (N6608, N6595, N2510, N3534);
and AND4 (N6609, N6561, N4724, N1998, N2852);
or OR3 (N6610, N6605, N3843, N4091);
nor NOR4 (N6611, N6604, N6080, N6008, N6034);
not NOT1 (N6612, N6588);
nor NOR3 (N6613, N6601, N3399, N3620);
or OR4 (N6614, N6589, N6451, N4082, N6365);
or OR2 (N6615, N6606, N475);
xor XOR2 (N6616, N6613, N1761);
nand NAND2 (N6617, N6616, N992);
or OR4 (N6618, N6612, N6203, N394, N6170);
and AND2 (N6619, N6611, N3602);
not NOT1 (N6620, N6608);
nand NAND2 (N6621, N6599, N4941);
nor NOR3 (N6622, N6609, N2896, N5570);
xor XOR2 (N6623, N6607, N1028);
and AND2 (N6624, N6617, N4270);
buf BUF1 (N6625, N6624);
buf BUF1 (N6626, N6620);
buf BUF1 (N6627, N6622);
nor NOR3 (N6628, N6610, N4964, N4482);
not NOT1 (N6629, N6618);
buf BUF1 (N6630, N6627);
buf BUF1 (N6631, N6621);
nor NOR3 (N6632, N6626, N944, N6501);
or OR4 (N6633, N6632, N6299, N5200, N6048);
or OR3 (N6634, N6631, N1184, N1167);
buf BUF1 (N6635, N6619);
buf BUF1 (N6636, N6629);
and AND2 (N6637, N6634, N296);
nor NOR2 (N6638, N6625, N4268);
nand NAND3 (N6639, N6633, N2794, N3322);
and AND3 (N6640, N6637, N3414, N2178);
not NOT1 (N6641, N6639);
or OR4 (N6642, N6623, N2603, N6130, N3992);
and AND2 (N6643, N6638, N1326);
or OR2 (N6644, N6643, N6079);
nand NAND2 (N6645, N6640, N1343);
not NOT1 (N6646, N6636);
nand NAND2 (N6647, N6645, N4453);
xor XOR2 (N6648, N6646, N224);
nor NOR4 (N6649, N6615, N4869, N3924, N3020);
and AND4 (N6650, N6647, N3987, N1949, N5734);
or OR3 (N6651, N6642, N3731, N304);
nand NAND2 (N6652, N6648, N5870);
nor NOR3 (N6653, N6651, N2522, N1574);
buf BUF1 (N6654, N6652);
nor NOR2 (N6655, N6649, N4553);
nand NAND3 (N6656, N6655, N5984, N2296);
nand NAND4 (N6657, N6641, N1185, N6489, N2826);
and AND3 (N6658, N6630, N6024, N5804);
buf BUF1 (N6659, N6658);
nand NAND4 (N6660, N6628, N4071, N3687, N2578);
not NOT1 (N6661, N6657);
buf BUF1 (N6662, N6653);
and AND3 (N6663, N6659, N1271, N3831);
or OR3 (N6664, N6644, N1889, N5177);
nor NOR2 (N6665, N6635, N1157);
or OR3 (N6666, N6661, N2280, N6183);
or OR2 (N6667, N6654, N4427);
xor XOR2 (N6668, N6666, N4722);
nand NAND2 (N6669, N6665, N4727);
xor XOR2 (N6670, N6663, N3892);
buf BUF1 (N6671, N6650);
nor NOR4 (N6672, N6656, N265, N1058, N3517);
nor NOR3 (N6673, N6660, N1073, N4421);
not NOT1 (N6674, N6671);
nor NOR4 (N6675, N6673, N1386, N3021, N3567);
buf BUF1 (N6676, N6672);
nor NOR4 (N6677, N6667, N5071, N5314, N461);
nand NAND4 (N6678, N6664, N2097, N1744, N2323);
buf BUF1 (N6679, N6670);
xor XOR2 (N6680, N6662, N1940);
nand NAND3 (N6681, N6668, N5902, N1268);
nand NAND4 (N6682, N6679, N1333, N3102, N5815);
nor NOR3 (N6683, N6681, N1172, N1861);
or OR2 (N6684, N6676, N826);
xor XOR2 (N6685, N6682, N3746);
or OR2 (N6686, N6678, N2610);
or OR4 (N6687, N6680, N3121, N5026, N1533);
and AND3 (N6688, N6669, N4400, N5621);
nand NAND4 (N6689, N6674, N6604, N3145, N430);
nand NAND4 (N6690, N6675, N22, N188, N4944);
xor XOR2 (N6691, N6690, N5681);
not NOT1 (N6692, N6614);
not NOT1 (N6693, N6691);
and AND3 (N6694, N6683, N2926, N5053);
not NOT1 (N6695, N6687);
not NOT1 (N6696, N6688);
nor NOR4 (N6697, N6684, N3284, N3468, N2316);
xor XOR2 (N6698, N6693, N2048);
xor XOR2 (N6699, N6689, N4176);
and AND3 (N6700, N6685, N6557, N6412);
and AND2 (N6701, N6695, N1617);
not NOT1 (N6702, N6686);
nand NAND2 (N6703, N6701, N3147);
not NOT1 (N6704, N6700);
nor NOR4 (N6705, N6703, N3518, N6169, N803);
buf BUF1 (N6706, N6702);
not NOT1 (N6707, N6697);
or OR3 (N6708, N6692, N1141, N3656);
or OR2 (N6709, N6696, N2498);
not NOT1 (N6710, N6699);
xor XOR2 (N6711, N6694, N1209);
nand NAND2 (N6712, N6707, N6522);
buf BUF1 (N6713, N6708);
or OR4 (N6714, N6710, N1570, N3610, N3442);
nand NAND4 (N6715, N6677, N5395, N3001, N3114);
buf BUF1 (N6716, N6715);
buf BUF1 (N6717, N6714);
buf BUF1 (N6718, N6704);
nand NAND4 (N6719, N6706, N5312, N5013, N102);
buf BUF1 (N6720, N6705);
or OR2 (N6721, N6718, N238);
not NOT1 (N6722, N6713);
xor XOR2 (N6723, N6721, N1572);
nand NAND3 (N6724, N6711, N2902, N1710);
buf BUF1 (N6725, N6712);
or OR3 (N6726, N6722, N4052, N956);
buf BUF1 (N6727, N6717);
and AND3 (N6728, N6709, N587, N5811);
not NOT1 (N6729, N6727);
xor XOR2 (N6730, N6728, N2280);
and AND3 (N6731, N6720, N43, N6607);
not NOT1 (N6732, N6725);
nor NOR3 (N6733, N6716, N3832, N1661);
or OR2 (N6734, N6724, N3823);
not NOT1 (N6735, N6734);
nor NOR4 (N6736, N6719, N1948, N5321, N3707);
nand NAND4 (N6737, N6698, N5240, N683, N4060);
and AND3 (N6738, N6731, N5473, N3218);
and AND4 (N6739, N6738, N55, N3605, N1054);
buf BUF1 (N6740, N6732);
nand NAND3 (N6741, N6730, N212, N704);
nor NOR4 (N6742, N6737, N3645, N6455, N4963);
and AND2 (N6743, N6723, N977);
buf BUF1 (N6744, N6733);
buf BUF1 (N6745, N6729);
xor XOR2 (N6746, N6743, N4054);
buf BUF1 (N6747, N6726);
and AND2 (N6748, N6739, N6559);
or OR3 (N6749, N6747, N4626, N5891);
nor NOR4 (N6750, N6736, N2771, N367, N1718);
and AND2 (N6751, N6744, N5370);
and AND3 (N6752, N6750, N4767, N23);
xor XOR2 (N6753, N6745, N2231);
nand NAND2 (N6754, N6748, N1531);
or OR2 (N6755, N6740, N6067);
buf BUF1 (N6756, N6753);
buf BUF1 (N6757, N6751);
buf BUF1 (N6758, N6746);
nor NOR2 (N6759, N6742, N2182);
not NOT1 (N6760, N6749);
nor NOR4 (N6761, N6760, N2580, N805, N3687);
buf BUF1 (N6762, N6758);
nor NOR4 (N6763, N6741, N4806, N3553, N671);
or OR3 (N6764, N6755, N4096, N3538);
nand NAND3 (N6765, N6759, N1994, N6339);
nand NAND4 (N6766, N6762, N1359, N653, N1897);
or OR3 (N6767, N6757, N5896, N3529);
nand NAND4 (N6768, N6765, N5818, N5441, N3459);
nand NAND4 (N6769, N6763, N966, N4368, N134);
buf BUF1 (N6770, N6756);
not NOT1 (N6771, N6735);
nor NOR2 (N6772, N6770, N1524);
xor XOR2 (N6773, N6766, N2940);
and AND2 (N6774, N6771, N6241);
and AND4 (N6775, N6769, N4389, N2797, N1603);
nand NAND3 (N6776, N6774, N4268, N3591);
nand NAND2 (N6777, N6764, N5628);
nor NOR2 (N6778, N6754, N2453);
or OR2 (N6779, N6752, N1375);
buf BUF1 (N6780, N6775);
xor XOR2 (N6781, N6767, N5591);
and AND4 (N6782, N6780, N1376, N3869, N6651);
nor NOR4 (N6783, N6773, N766, N1124, N2469);
xor XOR2 (N6784, N6777, N4047);
not NOT1 (N6785, N6772);
nand NAND2 (N6786, N6784, N230);
buf BUF1 (N6787, N6778);
and AND2 (N6788, N6782, N2097);
not NOT1 (N6789, N6787);
nand NAND2 (N6790, N6781, N5191);
not NOT1 (N6791, N6790);
and AND2 (N6792, N6779, N624);
nor NOR2 (N6793, N6783, N174);
buf BUF1 (N6794, N6768);
nand NAND4 (N6795, N6794, N6530, N4328, N1733);
buf BUF1 (N6796, N6791);
xor XOR2 (N6797, N6785, N4500);
and AND3 (N6798, N6796, N5028, N2309);
nand NAND3 (N6799, N6761, N4538, N5033);
nand NAND4 (N6800, N6792, N4172, N1479, N4073);
nor NOR4 (N6801, N6776, N5623, N1593, N3365);
nor NOR3 (N6802, N6798, N4397, N3199);
and AND4 (N6803, N6801, N1631, N5151, N14);
and AND2 (N6804, N6788, N6699);
xor XOR2 (N6805, N6803, N3106);
buf BUF1 (N6806, N6789);
nor NOR4 (N6807, N6805, N536, N5364, N3305);
not NOT1 (N6808, N6806);
xor XOR2 (N6809, N6807, N250);
and AND3 (N6810, N6809, N4945, N4229);
or OR4 (N6811, N6786, N3869, N1267, N3618);
not NOT1 (N6812, N6797);
nor NOR3 (N6813, N6795, N4403, N5452);
and AND2 (N6814, N6808, N3752);
nor NOR3 (N6815, N6813, N336, N3834);
nand NAND4 (N6816, N6814, N2778, N896, N4390);
xor XOR2 (N6817, N6812, N3536);
and AND4 (N6818, N6804, N988, N5347, N2869);
nor NOR4 (N6819, N6815, N2762, N954, N6111);
nand NAND2 (N6820, N6811, N2107);
xor XOR2 (N6821, N6802, N132);
and AND4 (N6822, N6799, N3172, N1907, N3997);
nand NAND4 (N6823, N6810, N4239, N3383, N1246);
and AND2 (N6824, N6800, N2708);
buf BUF1 (N6825, N6822);
not NOT1 (N6826, N6824);
nand NAND3 (N6827, N6818, N5131, N4667);
buf BUF1 (N6828, N6820);
nor NOR2 (N6829, N6821, N5645);
and AND3 (N6830, N6825, N394, N3917);
nor NOR4 (N6831, N6827, N5770, N6182, N5668);
or OR3 (N6832, N6823, N29, N5043);
and AND2 (N6833, N6826, N2612);
not NOT1 (N6834, N6832);
or OR4 (N6835, N6828, N6493, N1625, N4594);
nand NAND4 (N6836, N6834, N5368, N3123, N1344);
not NOT1 (N6837, N6833);
nor NOR3 (N6838, N6830, N3084, N710);
nor NOR2 (N6839, N6793, N4696);
nand NAND3 (N6840, N6839, N5218, N1477);
nand NAND3 (N6841, N6838, N5005, N1145);
xor XOR2 (N6842, N6819, N2724);
and AND2 (N6843, N6831, N645);
or OR2 (N6844, N6816, N2665);
not NOT1 (N6845, N6829);
buf BUF1 (N6846, N6843);
buf BUF1 (N6847, N6817);
nand NAND3 (N6848, N6842, N6164, N5923);
or OR2 (N6849, N6841, N2360);
or OR3 (N6850, N6849, N1096, N178);
not NOT1 (N6851, N6846);
or OR4 (N6852, N6848, N1899, N1797, N3727);
or OR4 (N6853, N6840, N4592, N5868, N1243);
and AND2 (N6854, N6837, N477);
xor XOR2 (N6855, N6836, N4703);
nor NOR2 (N6856, N6847, N2221);
nand NAND3 (N6857, N6853, N6780, N2220);
and AND3 (N6858, N6852, N6120, N6075);
not NOT1 (N6859, N6850);
buf BUF1 (N6860, N6845);
nor NOR2 (N6861, N6844, N5769);
not NOT1 (N6862, N6855);
and AND3 (N6863, N6835, N6668, N718);
and AND3 (N6864, N6861, N4428, N363);
or OR4 (N6865, N6858, N6426, N3441, N6045);
or OR3 (N6866, N6864, N4283, N4229);
nor NOR2 (N6867, N6860, N3664);
buf BUF1 (N6868, N6863);
or OR4 (N6869, N6854, N2298, N6379, N5327);
buf BUF1 (N6870, N6865);
buf BUF1 (N6871, N6870);
xor XOR2 (N6872, N6856, N2040);
or OR3 (N6873, N6859, N5949, N861);
xor XOR2 (N6874, N6851, N4715);
and AND3 (N6875, N6867, N4556, N3568);
nand NAND2 (N6876, N6875, N6628);
and AND3 (N6877, N6873, N6183, N4604);
nor NOR3 (N6878, N6874, N3723, N3478);
nand NAND2 (N6879, N6871, N870);
and AND3 (N6880, N6877, N4646, N1905);
not NOT1 (N6881, N6857);
buf BUF1 (N6882, N6879);
nor NOR4 (N6883, N6869, N5082, N6401, N3219);
xor XOR2 (N6884, N6872, N1506);
xor XOR2 (N6885, N6868, N5277);
nor NOR3 (N6886, N6876, N3705, N1453);
nor NOR2 (N6887, N6866, N4605);
and AND4 (N6888, N6880, N4865, N5527, N2874);
and AND4 (N6889, N6883, N6566, N5239, N1154);
buf BUF1 (N6890, N6885);
nand NAND4 (N6891, N6878, N4707, N4658, N1253);
xor XOR2 (N6892, N6862, N5285);
buf BUF1 (N6893, N6889);
buf BUF1 (N6894, N6887);
buf BUF1 (N6895, N6891);
and AND2 (N6896, N6884, N5721);
buf BUF1 (N6897, N6890);
xor XOR2 (N6898, N6882, N682);
not NOT1 (N6899, N6898);
or OR3 (N6900, N6886, N2986, N2175);
or OR3 (N6901, N6892, N4262, N1240);
and AND3 (N6902, N6899, N5934, N1908);
nor NOR2 (N6903, N6902, N2041);
xor XOR2 (N6904, N6894, N6610);
or OR4 (N6905, N6904, N4618, N3817, N5303);
buf BUF1 (N6906, N6896);
buf BUF1 (N6907, N6903);
nor NOR3 (N6908, N6897, N4677, N1170);
nand NAND2 (N6909, N6900, N4095);
or OR4 (N6910, N6905, N1475, N6591, N2623);
and AND4 (N6911, N6901, N6558, N6494, N1023);
not NOT1 (N6912, N6906);
nand NAND3 (N6913, N6910, N1662, N4667);
or OR2 (N6914, N6888, N6313);
xor XOR2 (N6915, N6908, N5617);
buf BUF1 (N6916, N6914);
or OR3 (N6917, N6895, N4014, N908);
nand NAND3 (N6918, N6917, N402, N941);
nand NAND2 (N6919, N6893, N3651);
nor NOR4 (N6920, N6915, N6236, N217, N1771);
not NOT1 (N6921, N6909);
nand NAND2 (N6922, N6912, N3124);
xor XOR2 (N6923, N6918, N3306);
buf BUF1 (N6924, N6881);
not NOT1 (N6925, N6919);
or OR4 (N6926, N6922, N1496, N6658, N2767);
and AND2 (N6927, N6911, N2090);
xor XOR2 (N6928, N6907, N2752);
nor NOR2 (N6929, N6923, N42);
nand NAND3 (N6930, N6920, N5935, N3731);
or OR2 (N6931, N6928, N5991);
nand NAND4 (N6932, N6929, N3505, N1781, N6643);
and AND4 (N6933, N6927, N2648, N3821, N4042);
nand NAND3 (N6934, N6926, N5347, N1342);
not NOT1 (N6935, N6930);
nor NOR4 (N6936, N6913, N5383, N5485, N203);
xor XOR2 (N6937, N6916, N2880);
nand NAND3 (N6938, N6936, N583, N3442);
and AND4 (N6939, N6934, N4062, N2452, N409);
and AND2 (N6940, N6937, N6157);
xor XOR2 (N6941, N6935, N5602);
xor XOR2 (N6942, N6939, N3393);
not NOT1 (N6943, N6941);
nor NOR3 (N6944, N6921, N4005, N1163);
nor NOR3 (N6945, N6942, N1859, N2183);
xor XOR2 (N6946, N6938, N5547);
nand NAND2 (N6947, N6933, N561);
nor NOR2 (N6948, N6945, N1395);
nor NOR3 (N6949, N6925, N2025, N6738);
or OR4 (N6950, N6924, N1395, N4658, N4551);
xor XOR2 (N6951, N6947, N312);
nand NAND3 (N6952, N6948, N3965, N2456);
not NOT1 (N6953, N6932);
or OR4 (N6954, N6931, N5500, N5414, N6058);
or OR4 (N6955, N6954, N4266, N6320, N3781);
or OR4 (N6956, N6940, N2257, N2818, N6457);
or OR2 (N6957, N6949, N4210);
nor NOR4 (N6958, N6952, N1722, N2111, N3270);
nor NOR4 (N6959, N6955, N1478, N2464, N2997);
nor NOR4 (N6960, N6959, N1332, N1626, N4327);
nand NAND4 (N6961, N6953, N5141, N2444, N6045);
buf BUF1 (N6962, N6958);
not NOT1 (N6963, N6962);
and AND2 (N6964, N6961, N4428);
nand NAND3 (N6965, N6963, N3907, N3608);
and AND2 (N6966, N6964, N5602);
not NOT1 (N6967, N6966);
nor NOR2 (N6968, N6965, N3322);
xor XOR2 (N6969, N6951, N1141);
and AND2 (N6970, N6969, N1671);
xor XOR2 (N6971, N6950, N5873);
nand NAND4 (N6972, N6960, N5104, N6891, N1240);
nand NAND2 (N6973, N6972, N4838);
buf BUF1 (N6974, N6946);
xor XOR2 (N6975, N6970, N5838);
and AND4 (N6976, N6967, N881, N4151, N2162);
and AND3 (N6977, N6974, N5961, N4614);
not NOT1 (N6978, N6973);
buf BUF1 (N6979, N6971);
xor XOR2 (N6980, N6976, N3704);
buf BUF1 (N6981, N6979);
or OR2 (N6982, N6957, N313);
nand NAND3 (N6983, N6968, N5482, N2950);
nand NAND4 (N6984, N6975, N5576, N3689, N6135);
nor NOR4 (N6985, N6956, N60, N6082, N488);
or OR2 (N6986, N6944, N1795);
nand NAND4 (N6987, N6982, N6765, N4114, N3192);
or OR2 (N6988, N6986, N2616);
nor NOR2 (N6989, N6987, N3594);
xor XOR2 (N6990, N6983, N4030);
buf BUF1 (N6991, N6990);
nor NOR3 (N6992, N6943, N6146, N2800);
nor NOR4 (N6993, N6978, N1642, N2778, N637);
not NOT1 (N6994, N6981);
nor NOR2 (N6995, N6980, N6624);
buf BUF1 (N6996, N6985);
not NOT1 (N6997, N6989);
nor NOR4 (N6998, N6988, N4304, N6505, N2442);
nor NOR4 (N6999, N6992, N5200, N4038, N1932);
not NOT1 (N7000, N6977);
not NOT1 (N7001, N7000);
nand NAND2 (N7002, N6995, N900);
and AND4 (N7003, N6997, N3282, N258, N5537);
nor NOR3 (N7004, N6994, N6676, N229);
or OR2 (N7005, N7001, N396);
xor XOR2 (N7006, N7002, N3048);
not NOT1 (N7007, N7003);
not NOT1 (N7008, N6998);
or OR2 (N7009, N6991, N5291);
or OR3 (N7010, N6993, N5770, N1222);
or OR4 (N7011, N7009, N3959, N1738, N5429);
xor XOR2 (N7012, N6999, N4608);
or OR2 (N7013, N6984, N4173);
and AND4 (N7014, N7013, N483, N5462, N3827);
nor NOR4 (N7015, N7007, N96, N3907, N3604);
buf BUF1 (N7016, N6996);
xor XOR2 (N7017, N7008, N1442);
xor XOR2 (N7018, N7015, N5376);
xor XOR2 (N7019, N7012, N2859);
buf BUF1 (N7020, N7017);
buf BUF1 (N7021, N7016);
xor XOR2 (N7022, N7019, N6060);
nor NOR4 (N7023, N7005, N4319, N5907, N2840);
xor XOR2 (N7024, N7018, N1397);
buf BUF1 (N7025, N7011);
xor XOR2 (N7026, N7024, N6250);
and AND2 (N7027, N7025, N5812);
xor XOR2 (N7028, N7020, N2202);
nor NOR3 (N7029, N7006, N217, N4479);
nor NOR3 (N7030, N7029, N6472, N6368);
buf BUF1 (N7031, N7030);
or OR4 (N7032, N7004, N4530, N2767, N867);
xor XOR2 (N7033, N7027, N2575);
nor NOR4 (N7034, N7032, N3828, N5660, N3581);
or OR4 (N7035, N7028, N6914, N3023, N4428);
nor NOR4 (N7036, N7035, N6603, N1517, N6129);
nor NOR4 (N7037, N7022, N664, N3095, N6327);
nor NOR2 (N7038, N7026, N4418);
nor NOR2 (N7039, N7033, N3980);
not NOT1 (N7040, N7038);
nand NAND3 (N7041, N7010, N1706, N5773);
xor XOR2 (N7042, N7037, N829);
or OR2 (N7043, N7040, N2029);
or OR4 (N7044, N7021, N3366, N2016, N3759);
not NOT1 (N7045, N7034);
nand NAND3 (N7046, N7023, N4280, N6810);
nor NOR3 (N7047, N7046, N117, N4634);
not NOT1 (N7048, N7044);
xor XOR2 (N7049, N7031, N689);
not NOT1 (N7050, N7045);
or OR2 (N7051, N7049, N4993);
nor NOR3 (N7052, N7042, N2096, N12);
nor NOR4 (N7053, N7047, N6153, N6917, N3171);
nand NAND3 (N7054, N7050, N454, N5437);
buf BUF1 (N7055, N7043);
buf BUF1 (N7056, N7036);
nand NAND4 (N7057, N7052, N2766, N3692, N2051);
not NOT1 (N7058, N7014);
nand NAND3 (N7059, N7055, N475, N511);
and AND2 (N7060, N7051, N6211);
buf BUF1 (N7061, N7048);
nand NAND4 (N7062, N7057, N3259, N3405, N3685);
nor NOR4 (N7063, N7058, N3244, N5836, N1209);
nor NOR4 (N7064, N7062, N1754, N3475, N1772);
nor NOR3 (N7065, N7059, N1305, N1391);
nand NAND3 (N7066, N7060, N6686, N2432);
not NOT1 (N7067, N7041);
buf BUF1 (N7068, N7053);
or OR4 (N7069, N7061, N4007, N5536, N4395);
not NOT1 (N7070, N7056);
nand NAND4 (N7071, N7054, N6341, N6042, N4367);
not NOT1 (N7072, N7067);
not NOT1 (N7073, N7065);
and AND4 (N7074, N7068, N2007, N1538, N3791);
not NOT1 (N7075, N7064);
and AND4 (N7076, N7039, N6353, N3457, N6578);
or OR4 (N7077, N7075, N152, N3569, N644);
or OR4 (N7078, N7070, N6846, N176, N754);
or OR3 (N7079, N7077, N3221, N4029);
nor NOR2 (N7080, N7078, N4175);
or OR4 (N7081, N7076, N2273, N3033, N5132);
not NOT1 (N7082, N7073);
and AND3 (N7083, N7063, N3132, N3673);
xor XOR2 (N7084, N7071, N2979);
nand NAND4 (N7085, N7069, N6310, N3587, N5008);
or OR4 (N7086, N7085, N1186, N2111, N2020);
nand NAND3 (N7087, N7086, N390, N1052);
or OR3 (N7088, N7081, N5804, N1509);
not NOT1 (N7089, N7072);
or OR3 (N7090, N7080, N2822, N3808);
buf BUF1 (N7091, N7089);
nor NOR3 (N7092, N7079, N3976, N412);
and AND3 (N7093, N7092, N416, N5580);
nor NOR3 (N7094, N7066, N5347, N4923);
nor NOR2 (N7095, N7094, N6949);
xor XOR2 (N7096, N7082, N978);
buf BUF1 (N7097, N7084);
not NOT1 (N7098, N7096);
nor NOR4 (N7099, N7088, N53, N5128, N6496);
xor XOR2 (N7100, N7093, N5484);
and AND2 (N7101, N7074, N6628);
and AND3 (N7102, N7095, N6626, N4005);
nand NAND2 (N7103, N7090, N4526);
not NOT1 (N7104, N7100);
or OR2 (N7105, N7102, N2237);
xor XOR2 (N7106, N7087, N1856);
not NOT1 (N7107, N7099);
xor XOR2 (N7108, N7097, N1441);
xor XOR2 (N7109, N7104, N5416);
or OR2 (N7110, N7108, N4607);
xor XOR2 (N7111, N7106, N2665);
nand NAND3 (N7112, N7111, N3197, N561);
xor XOR2 (N7113, N7083, N800);
or OR3 (N7114, N7105, N4844, N6820);
xor XOR2 (N7115, N7103, N2268);
nor NOR3 (N7116, N7112, N1706, N1087);
buf BUF1 (N7117, N7107);
buf BUF1 (N7118, N7117);
nor NOR2 (N7119, N7113, N6197);
and AND3 (N7120, N7114, N719, N377);
and AND4 (N7121, N7110, N2704, N4304, N5630);
buf BUF1 (N7122, N7116);
nand NAND2 (N7123, N7118, N3499);
and AND2 (N7124, N7109, N1317);
nor NOR4 (N7125, N7123, N2205, N1580, N4423);
nand NAND2 (N7126, N7098, N3994);
not NOT1 (N7127, N7125);
not NOT1 (N7128, N7124);
xor XOR2 (N7129, N7128, N3057);
not NOT1 (N7130, N7121);
not NOT1 (N7131, N7130);
nor NOR4 (N7132, N7120, N6926, N7125, N168);
nand NAND2 (N7133, N7101, N1426);
not NOT1 (N7134, N7115);
or OR4 (N7135, N7127, N930, N1714, N4691);
not NOT1 (N7136, N7129);
or OR4 (N7137, N7136, N5771, N2393, N464);
buf BUF1 (N7138, N7119);
xor XOR2 (N7139, N7138, N499);
buf BUF1 (N7140, N7134);
and AND4 (N7141, N7131, N1011, N6359, N5727);
and AND4 (N7142, N7091, N6147, N1937, N2625);
or OR3 (N7143, N7140, N3692, N84);
and AND2 (N7144, N7126, N97);
nor NOR3 (N7145, N7142, N2645, N2701);
buf BUF1 (N7146, N7135);
xor XOR2 (N7147, N7145, N2251);
nor NOR4 (N7148, N7122, N4594, N1442, N5343);
and AND4 (N7149, N7141, N4470, N5135, N671);
not NOT1 (N7150, N7132);
nand NAND4 (N7151, N7146, N1133, N1213, N621);
and AND4 (N7152, N7143, N6258, N2076, N3616);
nand NAND3 (N7153, N7150, N6387, N6030);
or OR4 (N7154, N7139, N5667, N595, N2919);
xor XOR2 (N7155, N7137, N447);
nor NOR2 (N7156, N7155, N3891);
or OR2 (N7157, N7153, N770);
and AND2 (N7158, N7154, N4597);
or OR2 (N7159, N7156, N5614);
not NOT1 (N7160, N7158);
and AND3 (N7161, N7144, N1541, N5767);
and AND2 (N7162, N7159, N333);
nand NAND2 (N7163, N7133, N4687);
and AND4 (N7164, N7148, N6457, N1845, N5206);
and AND3 (N7165, N7152, N4787, N1674);
nand NAND4 (N7166, N7149, N5412, N346, N1510);
not NOT1 (N7167, N7151);
buf BUF1 (N7168, N7166);
xor XOR2 (N7169, N7157, N6664);
buf BUF1 (N7170, N7169);
not NOT1 (N7171, N7147);
or OR2 (N7172, N7168, N4165);
and AND2 (N7173, N7172, N3848);
nand NAND4 (N7174, N7167, N5284, N936, N5086);
nor NOR4 (N7175, N7160, N286, N2762, N1656);
buf BUF1 (N7176, N7164);
or OR4 (N7177, N7176, N3247, N618, N3074);
buf BUF1 (N7178, N7175);
buf BUF1 (N7179, N7177);
xor XOR2 (N7180, N7178, N740);
buf BUF1 (N7181, N7171);
nor NOR3 (N7182, N7181, N96, N2506);
nand NAND4 (N7183, N7179, N6345, N2617, N4576);
not NOT1 (N7184, N7174);
buf BUF1 (N7185, N7182);
xor XOR2 (N7186, N7184, N4463);
nor NOR3 (N7187, N7170, N3684, N6830);
and AND3 (N7188, N7165, N5112, N1665);
or OR4 (N7189, N7173, N47, N3473, N6438);
nor NOR2 (N7190, N7188, N3233);
not NOT1 (N7191, N7185);
buf BUF1 (N7192, N7161);
not NOT1 (N7193, N7163);
nand NAND2 (N7194, N7192, N6391);
nand NAND2 (N7195, N7191, N3896);
nand NAND3 (N7196, N7193, N504, N2584);
nand NAND4 (N7197, N7190, N5101, N6457, N6226);
nand NAND2 (N7198, N7197, N1616);
nor NOR2 (N7199, N7186, N712);
and AND4 (N7200, N7196, N1353, N1869, N5698);
nor NOR4 (N7201, N7195, N5197, N2054, N970);
buf BUF1 (N7202, N7198);
buf BUF1 (N7203, N7194);
buf BUF1 (N7204, N7162);
nand NAND4 (N7205, N7199, N2319, N5122, N4658);
not NOT1 (N7206, N7205);
not NOT1 (N7207, N7206);
buf BUF1 (N7208, N7200);
nand NAND3 (N7209, N7187, N413, N1970);
nor NOR3 (N7210, N7209, N2591, N3238);
or OR3 (N7211, N7210, N1807, N4976);
nor NOR3 (N7212, N7211, N5158, N603);
not NOT1 (N7213, N7180);
or OR4 (N7214, N7212, N7178, N4991, N1562);
xor XOR2 (N7215, N7214, N5216);
nand NAND3 (N7216, N7203, N5751, N661);
not NOT1 (N7217, N7213);
nor NOR3 (N7218, N7183, N875, N3719);
xor XOR2 (N7219, N7215, N7197);
buf BUF1 (N7220, N7202);
or OR3 (N7221, N7220, N4174, N3560);
buf BUF1 (N7222, N7207);
nor NOR3 (N7223, N7222, N6663, N6183);
xor XOR2 (N7224, N7189, N6142);
nand NAND2 (N7225, N7216, N5201);
and AND4 (N7226, N7224, N1669, N1416, N6376);
nor NOR2 (N7227, N7201, N1847);
nand NAND2 (N7228, N7217, N5574);
and AND4 (N7229, N7227, N4414, N6412, N295);
not NOT1 (N7230, N7225);
xor XOR2 (N7231, N7228, N1040);
nor NOR2 (N7232, N7208, N1125);
or OR2 (N7233, N7204, N3644);
nor NOR4 (N7234, N7233, N4806, N1235, N2296);
nor NOR2 (N7235, N7223, N4484);
not NOT1 (N7236, N7221);
and AND3 (N7237, N7226, N492, N5041);
nor NOR2 (N7238, N7231, N6796);
buf BUF1 (N7239, N7232);
or OR4 (N7240, N7230, N3612, N3513, N3985);
xor XOR2 (N7241, N7219, N516);
nand NAND3 (N7242, N7234, N2096, N1906);
buf BUF1 (N7243, N7236);
not NOT1 (N7244, N7238);
and AND2 (N7245, N7235, N7074);
nand NAND3 (N7246, N7240, N5147, N6945);
xor XOR2 (N7247, N7242, N2501);
or OR3 (N7248, N7247, N3787, N820);
buf BUF1 (N7249, N7246);
nor NOR4 (N7250, N7237, N4009, N1523, N6444);
nand NAND3 (N7251, N7243, N2566, N3820);
nand NAND4 (N7252, N7244, N1309, N1127, N2730);
not NOT1 (N7253, N7229);
nor NOR3 (N7254, N7252, N1427, N7177);
and AND3 (N7255, N7218, N3851, N4111);
buf BUF1 (N7256, N7250);
xor XOR2 (N7257, N7256, N5162);
or OR3 (N7258, N7245, N883, N3794);
not NOT1 (N7259, N7257);
buf BUF1 (N7260, N7248);
and AND4 (N7261, N7259, N4262, N624, N2639);
buf BUF1 (N7262, N7249);
buf BUF1 (N7263, N7262);
buf BUF1 (N7264, N7254);
xor XOR2 (N7265, N7251, N6262);
nor NOR4 (N7266, N7253, N946, N7019, N3797);
xor XOR2 (N7267, N7255, N4023);
xor XOR2 (N7268, N7258, N6713);
nor NOR4 (N7269, N7268, N4091, N4536, N6815);
nor NOR4 (N7270, N7269, N4639, N2683, N4771);
and AND2 (N7271, N7260, N6809);
or OR3 (N7272, N7271, N4712, N259);
buf BUF1 (N7273, N7270);
nand NAND4 (N7274, N7264, N4372, N4943, N1474);
and AND4 (N7275, N7267, N5790, N3926, N6671);
xor XOR2 (N7276, N7273, N5928);
nor NOR4 (N7277, N7266, N4334, N1532, N3169);
and AND2 (N7278, N7241, N6754);
and AND4 (N7279, N7277, N3192, N124, N4681);
nor NOR4 (N7280, N7275, N1924, N1558, N2904);
buf BUF1 (N7281, N7276);
nand NAND3 (N7282, N7279, N6267, N714);
nand NAND3 (N7283, N7282, N6815, N6315);
not NOT1 (N7284, N7283);
nor NOR4 (N7285, N7263, N1783, N285, N5617);
and AND4 (N7286, N7274, N3178, N3047, N751);
buf BUF1 (N7287, N7285);
not NOT1 (N7288, N7272);
nor NOR3 (N7289, N7278, N2763, N1983);
nor NOR4 (N7290, N7287, N3054, N488, N580);
not NOT1 (N7291, N7286);
buf BUF1 (N7292, N7239);
not NOT1 (N7293, N7281);
and AND4 (N7294, N7293, N3633, N2935, N393);
not NOT1 (N7295, N7265);
nand NAND2 (N7296, N7288, N1685);
and AND3 (N7297, N7261, N1669, N4119);
and AND2 (N7298, N7290, N2752);
nand NAND3 (N7299, N7297, N4199, N5278);
nand NAND4 (N7300, N7289, N748, N1212, N3073);
buf BUF1 (N7301, N7292);
and AND4 (N7302, N7296, N5220, N889, N6228);
nand NAND3 (N7303, N7284, N7180, N5650);
nor NOR2 (N7304, N7300, N3062);
buf BUF1 (N7305, N7302);
nand NAND2 (N7306, N7303, N675);
buf BUF1 (N7307, N7295);
xor XOR2 (N7308, N7298, N186);
nand NAND3 (N7309, N7307, N6896, N183);
and AND2 (N7310, N7280, N2312);
nand NAND2 (N7311, N7310, N5993);
nor NOR4 (N7312, N7306, N5800, N1791, N4788);
not NOT1 (N7313, N7312);
nor NOR2 (N7314, N7301, N2874);
and AND3 (N7315, N7311, N5237, N718);
and AND4 (N7316, N7314, N2495, N7142, N7287);
xor XOR2 (N7317, N7304, N4278);
not NOT1 (N7318, N7291);
not NOT1 (N7319, N7294);
xor XOR2 (N7320, N7319, N38);
not NOT1 (N7321, N7305);
nand NAND4 (N7322, N7320, N6201, N6050, N6801);
or OR3 (N7323, N7299, N2166, N3946);
not NOT1 (N7324, N7323);
xor XOR2 (N7325, N7318, N5927);
or OR4 (N7326, N7324, N1616, N1540, N7184);
and AND2 (N7327, N7308, N7065);
not NOT1 (N7328, N7316);
nor NOR3 (N7329, N7322, N1726, N2015);
and AND4 (N7330, N7326, N641, N6234, N125);
nand NAND4 (N7331, N7327, N6381, N2794, N6150);
xor XOR2 (N7332, N7317, N4229);
not NOT1 (N7333, N7328);
buf BUF1 (N7334, N7309);
nand NAND2 (N7335, N7329, N5862);
buf BUF1 (N7336, N7321);
or OR2 (N7337, N7325, N6847);
or OR4 (N7338, N7332, N2229, N6440, N4386);
or OR3 (N7339, N7331, N3217, N3967);
nor NOR4 (N7340, N7313, N6046, N493, N2423);
xor XOR2 (N7341, N7335, N3502);
nor NOR2 (N7342, N7330, N5885);
nand NAND3 (N7343, N7315, N4062, N6736);
nand NAND2 (N7344, N7340, N4530);
and AND2 (N7345, N7333, N5506);
and AND3 (N7346, N7341, N6479, N7276);
nand NAND4 (N7347, N7342, N125, N5025, N5155);
or OR4 (N7348, N7346, N2716, N2797, N7033);
or OR3 (N7349, N7343, N5945, N6714);
or OR3 (N7350, N7348, N6490, N3741);
not NOT1 (N7351, N7338);
nand NAND4 (N7352, N7336, N6881, N5428, N6952);
nor NOR4 (N7353, N7339, N5537, N6433, N2550);
nand NAND3 (N7354, N7344, N2485, N188);
buf BUF1 (N7355, N7349);
nor NOR2 (N7356, N7355, N5702);
or OR2 (N7357, N7353, N4594);
nor NOR2 (N7358, N7347, N2351);
and AND3 (N7359, N7350, N730, N6558);
or OR3 (N7360, N7359, N4058, N4282);
and AND3 (N7361, N7345, N7196, N4012);
or OR3 (N7362, N7334, N560, N4029);
not NOT1 (N7363, N7357);
or OR4 (N7364, N7358, N7357, N4226, N3447);
nand NAND2 (N7365, N7361, N5585);
not NOT1 (N7366, N7354);
and AND4 (N7367, N7363, N5757, N1179, N4105);
xor XOR2 (N7368, N7364, N2715);
buf BUF1 (N7369, N7368);
not NOT1 (N7370, N7369);
nor NOR4 (N7371, N7366, N1088, N2668, N1642);
buf BUF1 (N7372, N7352);
buf BUF1 (N7373, N7372);
and AND4 (N7374, N7356, N4744, N1941, N2581);
and AND3 (N7375, N7374, N2949, N4740);
nor NOR4 (N7376, N7373, N6653, N2546, N5022);
xor XOR2 (N7377, N7362, N1701);
not NOT1 (N7378, N7371);
not NOT1 (N7379, N7376);
not NOT1 (N7380, N7375);
xor XOR2 (N7381, N7360, N5647);
xor XOR2 (N7382, N7377, N2959);
and AND4 (N7383, N7381, N688, N4417, N5530);
and AND4 (N7384, N7379, N356, N5959, N6794);
nor NOR4 (N7385, N7383, N2272, N4964, N7263);
buf BUF1 (N7386, N7337);
buf BUF1 (N7387, N7365);
nor NOR4 (N7388, N7387, N5521, N762, N7212);
buf BUF1 (N7389, N7351);
not NOT1 (N7390, N7367);
nand NAND4 (N7391, N7382, N6602, N793, N111);
nor NOR2 (N7392, N7391, N1748);
buf BUF1 (N7393, N7370);
buf BUF1 (N7394, N7392);
not NOT1 (N7395, N7386);
or OR2 (N7396, N7384, N6433);
nand NAND3 (N7397, N7380, N6220, N2827);
xor XOR2 (N7398, N7378, N1366);
nor NOR4 (N7399, N7393, N895, N3143, N3165);
nand NAND4 (N7400, N7399, N2797, N3465, N1138);
or OR3 (N7401, N7397, N6061, N778);
not NOT1 (N7402, N7389);
buf BUF1 (N7403, N7390);
xor XOR2 (N7404, N7394, N6121);
nor NOR2 (N7405, N7401, N6718);
and AND3 (N7406, N7405, N2980, N1425);
nor NOR2 (N7407, N7406, N3635);
not NOT1 (N7408, N7398);
or OR2 (N7409, N7388, N693);
buf BUF1 (N7410, N7385);
nor NOR4 (N7411, N7403, N6149, N264, N1713);
buf BUF1 (N7412, N7395);
nor NOR2 (N7413, N7404, N5100);
nor NOR3 (N7414, N7410, N275, N5101);
not NOT1 (N7415, N7413);
nor NOR2 (N7416, N7414, N2411);
nor NOR3 (N7417, N7412, N2518, N7296);
buf BUF1 (N7418, N7396);
nor NOR2 (N7419, N7418, N5511);
nor NOR3 (N7420, N7416, N4508, N6338);
and AND2 (N7421, N7408, N2119);
xor XOR2 (N7422, N7419, N1153);
or OR2 (N7423, N7417, N5677);
xor XOR2 (N7424, N7421, N1050);
not NOT1 (N7425, N7407);
not NOT1 (N7426, N7420);
and AND4 (N7427, N7426, N7315, N2783, N5230);
nor NOR4 (N7428, N7425, N125, N2479, N1458);
nand NAND2 (N7429, N7427, N173);
not NOT1 (N7430, N7415);
and AND4 (N7431, N7409, N3265, N63, N2324);
nand NAND3 (N7432, N7431, N6852, N5146);
and AND4 (N7433, N7428, N3180, N4943, N6963);
not NOT1 (N7434, N7433);
not NOT1 (N7435, N7411);
nand NAND2 (N7436, N7429, N3200);
and AND3 (N7437, N7435, N4767, N1071);
nand NAND4 (N7438, N7434, N4048, N2664, N1821);
nor NOR4 (N7439, N7437, N1240, N5347, N5656);
xor XOR2 (N7440, N7436, N5157);
or OR2 (N7441, N7423, N4451);
buf BUF1 (N7442, N7400);
or OR2 (N7443, N7442, N2020);
and AND3 (N7444, N7438, N4907, N5913);
not NOT1 (N7445, N7424);
and AND3 (N7446, N7402, N170, N729);
and AND4 (N7447, N7443, N239, N4906, N1517);
nand NAND4 (N7448, N7446, N3214, N3246, N6686);
buf BUF1 (N7449, N7440);
nand NAND4 (N7450, N7445, N4632, N3428, N4230);
not NOT1 (N7451, N7430);
nand NAND2 (N7452, N7451, N3433);
or OR3 (N7453, N7441, N211, N3122);
nand NAND2 (N7454, N7450, N3625);
nand NAND4 (N7455, N7432, N3244, N6573, N3430);
not NOT1 (N7456, N7453);
nand NAND3 (N7457, N7448, N6753, N4554);
and AND3 (N7458, N7439, N1994, N7354);
nor NOR4 (N7459, N7454, N6953, N4008, N860);
and AND2 (N7460, N7459, N6174);
nand NAND4 (N7461, N7452, N3652, N6932, N6009);
or OR2 (N7462, N7444, N7404);
or OR4 (N7463, N7462, N7428, N826, N494);
xor XOR2 (N7464, N7458, N2807);
nor NOR4 (N7465, N7457, N6074, N6781, N920);
buf BUF1 (N7466, N7463);
buf BUF1 (N7467, N7449);
not NOT1 (N7468, N7460);
xor XOR2 (N7469, N7455, N4537);
buf BUF1 (N7470, N7467);
xor XOR2 (N7471, N7464, N5281);
xor XOR2 (N7472, N7461, N5081);
buf BUF1 (N7473, N7469);
buf BUF1 (N7474, N7422);
and AND2 (N7475, N7471, N2452);
nor NOR4 (N7476, N7472, N1628, N476, N3476);
xor XOR2 (N7477, N7474, N6487);
and AND3 (N7478, N7468, N4735, N3730);
buf BUF1 (N7479, N7475);
or OR2 (N7480, N7465, N6173);
not NOT1 (N7481, N7480);
nand NAND2 (N7482, N7466, N5645);
nor NOR3 (N7483, N7470, N1069, N6153);
nand NAND2 (N7484, N7483, N1157);
buf BUF1 (N7485, N7484);
or OR3 (N7486, N7482, N2495, N2784);
not NOT1 (N7487, N7486);
buf BUF1 (N7488, N7478);
and AND2 (N7489, N7479, N3681);
xor XOR2 (N7490, N7473, N1981);
and AND3 (N7491, N7447, N3431, N1348);
nand NAND2 (N7492, N7488, N16);
nand NAND3 (N7493, N7492, N5150, N1586);
nor NOR4 (N7494, N7490, N3777, N5248, N5358);
nor NOR2 (N7495, N7477, N3798);
and AND3 (N7496, N7456, N3106, N2286);
and AND3 (N7497, N7494, N6583, N1714);
nand NAND3 (N7498, N7496, N5561, N1546);
nand NAND3 (N7499, N7489, N6961, N310);
xor XOR2 (N7500, N7476, N893);
nand NAND2 (N7501, N7491, N4622);
nor NOR3 (N7502, N7485, N156, N2028);
buf BUF1 (N7503, N7501);
xor XOR2 (N7504, N7481, N4030);
xor XOR2 (N7505, N7500, N6229);
and AND2 (N7506, N7487, N6903);
nor NOR2 (N7507, N7505, N1958);
xor XOR2 (N7508, N7499, N6884);
nor NOR2 (N7509, N7503, N3100);
buf BUF1 (N7510, N7508);
nand NAND3 (N7511, N7502, N93, N409);
nand NAND2 (N7512, N7509, N185);
xor XOR2 (N7513, N7497, N6465);
nand NAND3 (N7514, N7495, N6811, N3454);
not NOT1 (N7515, N7506);
or OR3 (N7516, N7510, N2719, N7385);
nand NAND4 (N7517, N7504, N268, N5756, N4284);
xor XOR2 (N7518, N7513, N4743);
not NOT1 (N7519, N7516);
nor NOR2 (N7520, N7515, N1417);
and AND4 (N7521, N7520, N1522, N2587, N3787);
and AND2 (N7522, N7514, N1787);
nand NAND4 (N7523, N7511, N3195, N3395, N2694);
not NOT1 (N7524, N7512);
or OR2 (N7525, N7498, N6321);
xor XOR2 (N7526, N7518, N2953);
xor XOR2 (N7527, N7507, N5870);
nor NOR2 (N7528, N7517, N5548);
and AND4 (N7529, N7525, N6403, N6492, N200);
not NOT1 (N7530, N7522);
not NOT1 (N7531, N7493);
xor XOR2 (N7532, N7521, N6673);
nor NOR3 (N7533, N7523, N6955, N6832);
xor XOR2 (N7534, N7527, N4804);
xor XOR2 (N7535, N7531, N5084);
nand NAND4 (N7536, N7524, N5568, N5140, N3231);
or OR2 (N7537, N7528, N5921);
nor NOR3 (N7538, N7530, N3765, N6779);
xor XOR2 (N7539, N7536, N2915);
xor XOR2 (N7540, N7538, N7204);
xor XOR2 (N7541, N7532, N552);
nand NAND4 (N7542, N7539, N129, N4737, N5419);
xor XOR2 (N7543, N7542, N3625);
buf BUF1 (N7544, N7537);
nand NAND2 (N7545, N7529, N5093);
not NOT1 (N7546, N7519);
or OR4 (N7547, N7526, N5551, N1452, N7449);
or OR2 (N7548, N7535, N5628);
nor NOR3 (N7549, N7534, N3626, N3510);
not NOT1 (N7550, N7549);
or OR2 (N7551, N7541, N2966);
and AND3 (N7552, N7544, N3039, N6643);
buf BUF1 (N7553, N7540);
nand NAND4 (N7554, N7547, N6534, N7537, N361);
not NOT1 (N7555, N7553);
xor XOR2 (N7556, N7555, N1497);
buf BUF1 (N7557, N7543);
not NOT1 (N7558, N7545);
and AND4 (N7559, N7548, N1151, N5068, N3921);
not NOT1 (N7560, N7550);
not NOT1 (N7561, N7560);
buf BUF1 (N7562, N7561);
xor XOR2 (N7563, N7552, N860);
nand NAND2 (N7564, N7562, N3241);
not NOT1 (N7565, N7558);
not NOT1 (N7566, N7551);
not NOT1 (N7567, N7559);
buf BUF1 (N7568, N7556);
nor NOR2 (N7569, N7554, N5727);
and AND4 (N7570, N7566, N4220, N1136, N1316);
buf BUF1 (N7571, N7546);
buf BUF1 (N7572, N7570);
buf BUF1 (N7573, N7572);
or OR2 (N7574, N7569, N6784);
and AND3 (N7575, N7563, N2033, N7275);
nor NOR3 (N7576, N7568, N6075, N4026);
buf BUF1 (N7577, N7565);
not NOT1 (N7578, N7576);
buf BUF1 (N7579, N7564);
nor NOR3 (N7580, N7577, N5642, N4258);
not NOT1 (N7581, N7575);
or OR3 (N7582, N7567, N3960, N891);
buf BUF1 (N7583, N7571);
xor XOR2 (N7584, N7533, N4417);
nand NAND3 (N7585, N7580, N1474, N5685);
not NOT1 (N7586, N7557);
not NOT1 (N7587, N7582);
and AND2 (N7588, N7578, N5849);
xor XOR2 (N7589, N7586, N3281);
nor NOR2 (N7590, N7589, N6781);
and AND3 (N7591, N7590, N2030, N7212);
not NOT1 (N7592, N7574);
not NOT1 (N7593, N7579);
not NOT1 (N7594, N7588);
nand NAND2 (N7595, N7592, N3973);
or OR2 (N7596, N7594, N4381);
buf BUF1 (N7597, N7573);
xor XOR2 (N7598, N7585, N7447);
nor NOR3 (N7599, N7584, N5696, N3233);
or OR2 (N7600, N7598, N5726);
not NOT1 (N7601, N7587);
not NOT1 (N7602, N7596);
xor XOR2 (N7603, N7599, N3588);
buf BUF1 (N7604, N7581);
nand NAND4 (N7605, N7603, N6756, N5657, N2039);
buf BUF1 (N7606, N7597);
buf BUF1 (N7607, N7583);
xor XOR2 (N7608, N7600, N2868);
or OR4 (N7609, N7591, N5607, N614, N3095);
and AND3 (N7610, N7604, N3408, N7334);
or OR3 (N7611, N7601, N4171, N5019);
xor XOR2 (N7612, N7608, N682);
nand NAND3 (N7613, N7606, N6092, N5331);
not NOT1 (N7614, N7610);
nor NOR3 (N7615, N7593, N3198, N6972);
not NOT1 (N7616, N7609);
nor NOR2 (N7617, N7607, N1756);
not NOT1 (N7618, N7605);
or OR4 (N7619, N7617, N2863, N6515, N942);
buf BUF1 (N7620, N7611);
not NOT1 (N7621, N7619);
xor XOR2 (N7622, N7595, N1856);
not NOT1 (N7623, N7621);
nand NAND2 (N7624, N7613, N1491);
nand NAND2 (N7625, N7622, N5057);
buf BUF1 (N7626, N7602);
or OR4 (N7627, N7612, N6892, N1775, N3241);
xor XOR2 (N7628, N7625, N3643);
buf BUF1 (N7629, N7615);
not NOT1 (N7630, N7624);
and AND4 (N7631, N7626, N1575, N3797, N7388);
not NOT1 (N7632, N7614);
and AND3 (N7633, N7632, N111, N5325);
or OR2 (N7634, N7628, N6495);
or OR3 (N7635, N7618, N1893, N4213);
nand NAND4 (N7636, N7633, N4514, N4419, N3514);
buf BUF1 (N7637, N7616);
buf BUF1 (N7638, N7620);
buf BUF1 (N7639, N7629);
nand NAND2 (N7640, N7627, N5644);
not NOT1 (N7641, N7640);
nor NOR3 (N7642, N7637, N5043, N1974);
not NOT1 (N7643, N7639);
and AND2 (N7644, N7634, N6885);
buf BUF1 (N7645, N7623);
xor XOR2 (N7646, N7630, N4692);
buf BUF1 (N7647, N7642);
buf BUF1 (N7648, N7635);
nor NOR3 (N7649, N7638, N2338, N4598);
nor NOR2 (N7650, N7643, N3174);
and AND2 (N7651, N7647, N2600);
and AND3 (N7652, N7641, N523, N5712);
nand NAND3 (N7653, N7652, N4707, N7001);
nand NAND4 (N7654, N7631, N2055, N4908, N6592);
or OR4 (N7655, N7650, N3764, N5930, N4679);
not NOT1 (N7656, N7645);
xor XOR2 (N7657, N7651, N124);
or OR4 (N7658, N7636, N5080, N4691, N821);
or OR2 (N7659, N7653, N3640);
or OR4 (N7660, N7649, N4375, N754, N4275);
nand NAND4 (N7661, N7644, N25, N6684, N4169);
not NOT1 (N7662, N7646);
and AND2 (N7663, N7648, N2922);
and AND2 (N7664, N7655, N3057);
buf BUF1 (N7665, N7662);
or OR4 (N7666, N7654, N1256, N5858, N2100);
buf BUF1 (N7667, N7656);
nand NAND2 (N7668, N7658, N3861);
buf BUF1 (N7669, N7660);
or OR4 (N7670, N7667, N3604, N3796, N5454);
nand NAND2 (N7671, N7664, N4582);
nor NOR2 (N7672, N7657, N3449);
buf BUF1 (N7673, N7659);
nor NOR4 (N7674, N7663, N1068, N1606, N6673);
not NOT1 (N7675, N7673);
not NOT1 (N7676, N7666);
nor NOR2 (N7677, N7665, N3619);
xor XOR2 (N7678, N7674, N3924);
nand NAND4 (N7679, N7671, N1393, N5330, N4303);
and AND2 (N7680, N7669, N2960);
not NOT1 (N7681, N7675);
xor XOR2 (N7682, N7681, N5505);
buf BUF1 (N7683, N7670);
not NOT1 (N7684, N7679);
buf BUF1 (N7685, N7676);
nor NOR3 (N7686, N7661, N466, N1428);
xor XOR2 (N7687, N7683, N2014);
buf BUF1 (N7688, N7687);
nor NOR2 (N7689, N7688, N3230);
xor XOR2 (N7690, N7680, N4912);
and AND2 (N7691, N7689, N336);
not NOT1 (N7692, N7677);
buf BUF1 (N7693, N7682);
buf BUF1 (N7694, N7693);
and AND4 (N7695, N7685, N1386, N454, N3828);
xor XOR2 (N7696, N7686, N6430);
and AND4 (N7697, N7668, N449, N3695, N7439);
nor NOR4 (N7698, N7690, N1381, N5407, N6275);
and AND2 (N7699, N7694, N3712);
nand NAND3 (N7700, N7696, N688, N4565);
nand NAND3 (N7701, N7697, N6255, N4892);
xor XOR2 (N7702, N7700, N5192);
nor NOR4 (N7703, N7695, N4769, N7077, N3207);
buf BUF1 (N7704, N7691);
nor NOR3 (N7705, N7699, N3989, N5558);
xor XOR2 (N7706, N7698, N2129);
or OR4 (N7707, N7684, N403, N5511, N2497);
xor XOR2 (N7708, N7704, N2082);
nor NOR3 (N7709, N7707, N2522, N35);
nand NAND4 (N7710, N7678, N7692, N2519, N3610);
nor NOR2 (N7711, N2105, N5152);
xor XOR2 (N7712, N7711, N4656);
or OR4 (N7713, N7672, N2039, N7075, N6926);
and AND2 (N7714, N7701, N459);
nand NAND4 (N7715, N7709, N5410, N1321, N7424);
buf BUF1 (N7716, N7712);
or OR2 (N7717, N7708, N5035);
and AND3 (N7718, N7716, N6314, N5090);
buf BUF1 (N7719, N7714);
and AND4 (N7720, N7719, N858, N7180, N4988);
or OR4 (N7721, N7706, N3472, N4926, N902);
nor NOR2 (N7722, N7705, N5802);
xor XOR2 (N7723, N7722, N975);
xor XOR2 (N7724, N7710, N3361);
buf BUF1 (N7725, N7703);
not NOT1 (N7726, N7721);
nor NOR4 (N7727, N7702, N1677, N361, N1565);
or OR4 (N7728, N7725, N420, N2142, N2027);
not NOT1 (N7729, N7727);
not NOT1 (N7730, N7717);
xor XOR2 (N7731, N7713, N1101);
and AND2 (N7732, N7723, N1733);
nor NOR2 (N7733, N7715, N2238);
xor XOR2 (N7734, N7732, N7569);
not NOT1 (N7735, N7729);
buf BUF1 (N7736, N7726);
not NOT1 (N7737, N7728);
nand NAND3 (N7738, N7736, N6655, N1537);
nand NAND2 (N7739, N7737, N696);
not NOT1 (N7740, N7720);
nor NOR2 (N7741, N7738, N1647);
xor XOR2 (N7742, N7734, N2783);
buf BUF1 (N7743, N7735);
nand NAND3 (N7744, N7731, N4093, N5511);
not NOT1 (N7745, N7739);
buf BUF1 (N7746, N7733);
or OR4 (N7747, N7745, N5639, N3017, N6060);
and AND2 (N7748, N7746, N6785);
buf BUF1 (N7749, N7748);
not NOT1 (N7750, N7740);
nand NAND3 (N7751, N7747, N6918, N6155);
not NOT1 (N7752, N7750);
xor XOR2 (N7753, N7741, N4159);
and AND2 (N7754, N7753, N3442);
buf BUF1 (N7755, N7754);
and AND2 (N7756, N7730, N5394);
nor NOR4 (N7757, N7756, N7250, N4135, N1614);
nor NOR2 (N7758, N7749, N6981);
not NOT1 (N7759, N7752);
nand NAND2 (N7760, N7758, N6104);
nor NOR3 (N7761, N7759, N4225, N5872);
not NOT1 (N7762, N7751);
nand NAND3 (N7763, N7757, N2786, N243);
nand NAND2 (N7764, N7762, N56);
nor NOR2 (N7765, N7743, N2352);
or OR2 (N7766, N7744, N5316);
buf BUF1 (N7767, N7760);
xor XOR2 (N7768, N7724, N3549);
buf BUF1 (N7769, N7768);
nor NOR4 (N7770, N7765, N7001, N2944, N268);
xor XOR2 (N7771, N7755, N7027);
not NOT1 (N7772, N7766);
or OR3 (N7773, N7769, N4008, N3497);
nand NAND3 (N7774, N7763, N5335, N6118);
buf BUF1 (N7775, N7718);
and AND2 (N7776, N7742, N486);
or OR2 (N7777, N7772, N1280);
xor XOR2 (N7778, N7761, N5668);
and AND3 (N7779, N7770, N5714, N4857);
nor NOR3 (N7780, N7775, N2954, N6546);
buf BUF1 (N7781, N7779);
buf BUF1 (N7782, N7774);
not NOT1 (N7783, N7780);
buf BUF1 (N7784, N7781);
or OR4 (N7785, N7771, N7111, N2077, N5278);
nand NAND4 (N7786, N7778, N7434, N5799, N5293);
not NOT1 (N7787, N7773);
nand NAND4 (N7788, N7777, N3123, N5113, N696);
or OR2 (N7789, N7787, N4723);
nor NOR2 (N7790, N7785, N114);
xor XOR2 (N7791, N7782, N2667);
not NOT1 (N7792, N7783);
and AND2 (N7793, N7784, N4222);
not NOT1 (N7794, N7764);
and AND3 (N7795, N7767, N2730, N4243);
xor XOR2 (N7796, N7795, N1919);
or OR4 (N7797, N7794, N3623, N541, N3570);
xor XOR2 (N7798, N7796, N1597);
buf BUF1 (N7799, N7792);
nand NAND4 (N7800, N7786, N2236, N6445, N378);
nor NOR4 (N7801, N7788, N924, N4768, N1534);
or OR4 (N7802, N7790, N3697, N1399, N1293);
and AND4 (N7803, N7789, N1392, N2237, N3244);
nor NOR3 (N7804, N7797, N3087, N6227);
nor NOR2 (N7805, N7801, N5375);
nor NOR2 (N7806, N7802, N2404);
nand NAND2 (N7807, N7798, N2156);
xor XOR2 (N7808, N7806, N538);
not NOT1 (N7809, N7807);
or OR2 (N7810, N7805, N3544);
nand NAND2 (N7811, N7799, N6321);
and AND4 (N7812, N7800, N1843, N7026, N3791);
xor XOR2 (N7813, N7803, N1542);
buf BUF1 (N7814, N7793);
nor NOR3 (N7815, N7811, N754, N3793);
and AND2 (N7816, N7804, N1921);
or OR4 (N7817, N7808, N747, N7107, N4267);
buf BUF1 (N7818, N7813);
nor NOR3 (N7819, N7776, N3127, N2737);
nand NAND2 (N7820, N7810, N4353);
or OR2 (N7821, N7817, N4356);
and AND2 (N7822, N7820, N1941);
and AND2 (N7823, N7821, N7113);
buf BUF1 (N7824, N7818);
xor XOR2 (N7825, N7791, N1088);
or OR2 (N7826, N7809, N4665);
and AND3 (N7827, N7812, N5866, N5467);
nand NAND2 (N7828, N7824, N598);
and AND2 (N7829, N7825, N1413);
xor XOR2 (N7830, N7827, N2073);
not NOT1 (N7831, N7815);
not NOT1 (N7832, N7822);
nor NOR2 (N7833, N7816, N1980);
nand NAND4 (N7834, N7819, N496, N6254, N6821);
nand NAND2 (N7835, N7814, N979);
nor NOR2 (N7836, N7826, N7684);
buf BUF1 (N7837, N7831);
and AND3 (N7838, N7836, N4763, N6824);
not NOT1 (N7839, N7832);
xor XOR2 (N7840, N7838, N2976);
or OR3 (N7841, N7823, N1318, N4541);
and AND3 (N7842, N7841, N4663, N2890);
nor NOR4 (N7843, N7833, N2755, N1122, N6831);
xor XOR2 (N7844, N7840, N276);
or OR3 (N7845, N7837, N4766, N6737);
or OR2 (N7846, N7842, N4169);
nand NAND3 (N7847, N7830, N7722, N3536);
nand NAND3 (N7848, N7845, N5494, N5941);
xor XOR2 (N7849, N7835, N330);
buf BUF1 (N7850, N7828);
not NOT1 (N7851, N7850);
nor NOR3 (N7852, N7843, N5235, N3891);
not NOT1 (N7853, N7852);
xor XOR2 (N7854, N7834, N4481);
nand NAND3 (N7855, N7853, N574, N4994);
or OR4 (N7856, N7849, N6370, N51, N616);
not NOT1 (N7857, N7855);
nand NAND3 (N7858, N7856, N4381, N2175);
not NOT1 (N7859, N7857);
xor XOR2 (N7860, N7847, N1381);
nor NOR2 (N7861, N7846, N3188);
or OR4 (N7862, N7829, N906, N778, N7395);
nand NAND2 (N7863, N7862, N1008);
and AND3 (N7864, N7854, N1771, N619);
and AND2 (N7865, N7839, N5352);
or OR4 (N7866, N7848, N2569, N74, N3328);
or OR2 (N7867, N7864, N1312);
nor NOR3 (N7868, N7865, N6482, N1290);
or OR3 (N7869, N7851, N5289, N6059);
xor XOR2 (N7870, N7863, N2535);
nor NOR4 (N7871, N7870, N3935, N1982, N6004);
nor NOR3 (N7872, N7859, N4554, N4171);
or OR2 (N7873, N7871, N1536);
and AND3 (N7874, N7860, N4548, N6954);
nor NOR2 (N7875, N7873, N3251);
not NOT1 (N7876, N7858);
nand NAND2 (N7877, N7876, N7740);
nor NOR2 (N7878, N7868, N7841);
buf BUF1 (N7879, N7861);
not NOT1 (N7880, N7867);
buf BUF1 (N7881, N7872);
xor XOR2 (N7882, N7881, N7405);
nor NOR2 (N7883, N7878, N1073);
xor XOR2 (N7884, N7883, N2075);
xor XOR2 (N7885, N7869, N514);
buf BUF1 (N7886, N7844);
xor XOR2 (N7887, N7880, N1570);
not NOT1 (N7888, N7886);
buf BUF1 (N7889, N7888);
nor NOR2 (N7890, N7875, N6770);
and AND3 (N7891, N7874, N6852, N1498);
xor XOR2 (N7892, N7891, N1705);
xor XOR2 (N7893, N7890, N3904);
and AND3 (N7894, N7882, N539, N5939);
nor NOR4 (N7895, N7866, N6760, N5156, N2761);
xor XOR2 (N7896, N7893, N151);
or OR2 (N7897, N7895, N912);
xor XOR2 (N7898, N7896, N7728);
not NOT1 (N7899, N7897);
and AND2 (N7900, N7887, N6546);
xor XOR2 (N7901, N7884, N2661);
nand NAND2 (N7902, N7889, N4371);
buf BUF1 (N7903, N7901);
not NOT1 (N7904, N7879);
nand NAND2 (N7905, N7894, N4695);
not NOT1 (N7906, N7902);
nand NAND3 (N7907, N7903, N3775, N3197);
xor XOR2 (N7908, N7877, N6969);
nand NAND4 (N7909, N7905, N7201, N4018, N7089);
buf BUF1 (N7910, N7898);
nor NOR2 (N7911, N7885, N5480);
or OR4 (N7912, N7911, N7824, N5451, N3281);
buf BUF1 (N7913, N7892);
buf BUF1 (N7914, N7906);
nor NOR3 (N7915, N7904, N257, N2124);
not NOT1 (N7916, N7915);
xor XOR2 (N7917, N7909, N4593);
xor XOR2 (N7918, N7914, N6418);
xor XOR2 (N7919, N7916, N4591);
or OR2 (N7920, N7908, N4946);
nor NOR4 (N7921, N7907, N4987, N266, N6326);
buf BUF1 (N7922, N7910);
and AND3 (N7923, N7900, N2192, N4620);
nand NAND3 (N7924, N7913, N2143, N2820);
buf BUF1 (N7925, N7917);
nor NOR2 (N7926, N7925, N547);
xor XOR2 (N7927, N7924, N593);
or OR2 (N7928, N7927, N6609);
buf BUF1 (N7929, N7920);
nor NOR3 (N7930, N7918, N6592, N6645);
xor XOR2 (N7931, N7929, N5861);
buf BUF1 (N7932, N7923);
xor XOR2 (N7933, N7899, N2019);
buf BUF1 (N7934, N7933);
not NOT1 (N7935, N7926);
and AND2 (N7936, N7928, N1160);
nand NAND2 (N7937, N7922, N296);
nand NAND4 (N7938, N7930, N7536, N6194, N6296);
buf BUF1 (N7939, N7931);
nor NOR3 (N7940, N7937, N1499, N4153);
or OR4 (N7941, N7938, N1945, N3889, N1795);
or OR4 (N7942, N7941, N9, N6754, N4448);
buf BUF1 (N7943, N7940);
or OR4 (N7944, N7935, N1380, N3348, N5373);
and AND3 (N7945, N7943, N3420, N2862);
xor XOR2 (N7946, N7944, N6878);
nor NOR2 (N7947, N7946, N5248);
or OR2 (N7948, N7912, N1067);
not NOT1 (N7949, N7921);
buf BUF1 (N7950, N7942);
buf BUF1 (N7951, N7948);
nand NAND3 (N7952, N7949, N5118, N7773);
or OR4 (N7953, N7951, N3864, N5769, N1675);
not NOT1 (N7954, N7953);
nand NAND3 (N7955, N7945, N2689, N7378);
nor NOR3 (N7956, N7936, N2937, N1662);
buf BUF1 (N7957, N7952);
buf BUF1 (N7958, N7950);
and AND4 (N7959, N7957, N1522, N4829, N1421);
not NOT1 (N7960, N7919);
or OR3 (N7961, N7939, N1352, N2338);
not NOT1 (N7962, N7961);
not NOT1 (N7963, N7947);
nor NOR2 (N7964, N7959, N6110);
and AND4 (N7965, N7960, N505, N547, N6217);
or OR3 (N7966, N7962, N5308, N5335);
buf BUF1 (N7967, N7965);
and AND3 (N7968, N7932, N3097, N5896);
nand NAND4 (N7969, N7955, N2601, N4918, N2626);
not NOT1 (N7970, N7958);
buf BUF1 (N7971, N7967);
or OR4 (N7972, N7954, N6288, N4099, N1911);
and AND4 (N7973, N7971, N6384, N1499, N6275);
buf BUF1 (N7974, N7934);
nor NOR2 (N7975, N7973, N3353);
and AND3 (N7976, N7972, N4475, N7333);
nand NAND4 (N7977, N7964, N4357, N6014, N4513);
nor NOR4 (N7978, N7963, N845, N6929, N1222);
not NOT1 (N7979, N7974);
nand NAND2 (N7980, N7966, N6704);
xor XOR2 (N7981, N7980, N4166);
xor XOR2 (N7982, N7970, N2662);
or OR4 (N7983, N7981, N5723, N2886, N1538);
not NOT1 (N7984, N7983);
xor XOR2 (N7985, N7968, N6803);
xor XOR2 (N7986, N7982, N3790);
not NOT1 (N7987, N7975);
or OR4 (N7988, N7979, N1494, N2641, N3575);
or OR2 (N7989, N7986, N3574);
or OR4 (N7990, N7978, N1337, N6393, N229);
not NOT1 (N7991, N7989);
xor XOR2 (N7992, N7988, N1878);
not NOT1 (N7993, N7987);
nand NAND4 (N7994, N7976, N2167, N6738, N5637);
or OR2 (N7995, N7991, N233);
not NOT1 (N7996, N7956);
nor NOR2 (N7997, N7992, N18);
xor XOR2 (N7998, N7990, N3315);
or OR2 (N7999, N7969, N7973);
not NOT1 (N8000, N7996);
not NOT1 (N8001, N7997);
xor XOR2 (N8002, N8001, N1975);
nand NAND3 (N8003, N7977, N5804, N7999);
xor XOR2 (N8004, N3712, N266);
nor NOR4 (N8005, N7995, N6717, N687, N5814);
and AND4 (N8006, N8003, N3910, N4525, N911);
xor XOR2 (N8007, N8006, N1237);
or OR2 (N8008, N8000, N4946);
buf BUF1 (N8009, N8008);
nand NAND3 (N8010, N8009, N3086, N5066);
nor NOR4 (N8011, N7993, N5561, N1976, N924);
nor NOR4 (N8012, N8004, N2485, N1692, N5404);
and AND4 (N8013, N7994, N5685, N5267, N6145);
and AND4 (N8014, N8010, N5960, N7214, N5926);
not NOT1 (N8015, N7984);
not NOT1 (N8016, N8007);
nand NAND3 (N8017, N8011, N1926, N6058);
nand NAND3 (N8018, N8005, N3233, N7630);
nand NAND3 (N8019, N8014, N206, N2335);
and AND3 (N8020, N8017, N6658, N7743);
buf BUF1 (N8021, N8018);
not NOT1 (N8022, N8002);
not NOT1 (N8023, N8013);
and AND2 (N8024, N8019, N7414);
nand NAND3 (N8025, N8023, N2420, N2727);
and AND2 (N8026, N7985, N1693);
xor XOR2 (N8027, N8025, N7715);
not NOT1 (N8028, N8026);
or OR3 (N8029, N8020, N6156, N4659);
nand NAND2 (N8030, N8015, N7236);
buf BUF1 (N8031, N7998);
or OR2 (N8032, N8016, N5226);
buf BUF1 (N8033, N8027);
buf BUF1 (N8034, N8032);
nor NOR3 (N8035, N8028, N1712, N3293);
nor NOR3 (N8036, N8029, N2962, N5854);
buf BUF1 (N8037, N8024);
nor NOR3 (N8038, N8035, N4781, N4435);
buf BUF1 (N8039, N8030);
and AND2 (N8040, N8021, N6053);
xor XOR2 (N8041, N8031, N2460);
nand NAND2 (N8042, N8041, N3901);
nand NAND4 (N8043, N8042, N6037, N96, N4982);
not NOT1 (N8044, N8039);
xor XOR2 (N8045, N8036, N1421);
buf BUF1 (N8046, N8045);
or OR3 (N8047, N8043, N2824, N2720);
buf BUF1 (N8048, N8038);
xor XOR2 (N8049, N8046, N3895);
nor NOR2 (N8050, N8044, N314);
or OR4 (N8051, N8048, N7837, N3746, N5756);
xor XOR2 (N8052, N8034, N4945);
not NOT1 (N8053, N8049);
buf BUF1 (N8054, N8047);
nand NAND3 (N8055, N8050, N1607, N4903);
not NOT1 (N8056, N8053);
nor NOR3 (N8057, N8051, N3755, N5534);
not NOT1 (N8058, N8055);
and AND4 (N8059, N8040, N2515, N5464, N3280);
xor XOR2 (N8060, N8037, N6698);
xor XOR2 (N8061, N8022, N1132);
or OR4 (N8062, N8057, N6590, N7401, N8004);
buf BUF1 (N8063, N8033);
or OR2 (N8064, N8063, N3263);
not NOT1 (N8065, N8058);
and AND4 (N8066, N8052, N6223, N5865, N146);
buf BUF1 (N8067, N8054);
xor XOR2 (N8068, N8066, N7112);
and AND2 (N8069, N8012, N1599);
not NOT1 (N8070, N8056);
nor NOR4 (N8071, N8061, N137, N8002, N7021);
buf BUF1 (N8072, N8071);
and AND4 (N8073, N8059, N5328, N3707, N1401);
buf BUF1 (N8074, N8072);
nor NOR2 (N8075, N8060, N216);
not NOT1 (N8076, N8065);
nand NAND2 (N8077, N8075, N1732);
not NOT1 (N8078, N8076);
buf BUF1 (N8079, N8070);
buf BUF1 (N8080, N8079);
and AND3 (N8081, N8080, N3864, N3890);
buf BUF1 (N8082, N8078);
nor NOR3 (N8083, N8074, N7729, N997);
or OR3 (N8084, N8062, N559, N5224);
and AND4 (N8085, N8068, N5296, N5477, N100);
nor NOR3 (N8086, N8073, N1800, N1910);
buf BUF1 (N8087, N8082);
or OR2 (N8088, N8064, N4134);
xor XOR2 (N8089, N8084, N900);
nor NOR2 (N8090, N8069, N4429);
nand NAND4 (N8091, N8089, N3574, N6596, N6028);
and AND4 (N8092, N8088, N4815, N2858, N2622);
nor NOR2 (N8093, N8083, N1323);
nor NOR4 (N8094, N8087, N6217, N2051, N353);
buf BUF1 (N8095, N8086);
nor NOR4 (N8096, N8091, N2351, N2905, N5720);
nand NAND2 (N8097, N8093, N4285);
not NOT1 (N8098, N8085);
not NOT1 (N8099, N8067);
or OR3 (N8100, N8081, N5905, N4268);
xor XOR2 (N8101, N8092, N7411);
and AND3 (N8102, N8096, N6316, N4489);
and AND4 (N8103, N8090, N2143, N3069, N6889);
buf BUF1 (N8104, N8077);
nor NOR3 (N8105, N8102, N1916, N1646);
buf BUF1 (N8106, N8105);
and AND4 (N8107, N8095, N372, N74, N2018);
and AND2 (N8108, N8104, N7786);
xor XOR2 (N8109, N8099, N116);
nand NAND4 (N8110, N8106, N1533, N47, N7691);
xor XOR2 (N8111, N8103, N5343);
and AND3 (N8112, N8111, N3993, N7460);
nand NAND2 (N8113, N8100, N3427);
nor NOR4 (N8114, N8109, N6070, N5205, N5787);
buf BUF1 (N8115, N8110);
and AND3 (N8116, N8098, N1647, N2258);
and AND2 (N8117, N8115, N3332);
xor XOR2 (N8118, N8117, N1083);
buf BUF1 (N8119, N8114);
buf BUF1 (N8120, N8112);
nand NAND2 (N8121, N8107, N929);
not NOT1 (N8122, N8116);
or OR2 (N8123, N8108, N3229);
and AND4 (N8124, N8113, N5588, N4104, N1620);
xor XOR2 (N8125, N8123, N1157);
nand NAND2 (N8126, N8094, N3455);
nor NOR3 (N8127, N8124, N3661, N7090);
or OR3 (N8128, N8121, N5814, N1205);
nand NAND2 (N8129, N8126, N6136);
not NOT1 (N8130, N8118);
nor NOR3 (N8131, N8122, N4463, N5286);
xor XOR2 (N8132, N8129, N7216);
nor NOR2 (N8133, N8132, N349);
or OR4 (N8134, N8125, N1207, N1310, N5172);
nand NAND4 (N8135, N8134, N4908, N7752, N3510);
not NOT1 (N8136, N8133);
or OR4 (N8137, N8128, N79, N1796, N3205);
or OR3 (N8138, N8101, N8017, N5053);
nor NOR2 (N8139, N8137, N7682);
not NOT1 (N8140, N8130);
buf BUF1 (N8141, N8135);
xor XOR2 (N8142, N8140, N7085);
buf BUF1 (N8143, N8127);
nand NAND3 (N8144, N8139, N573, N3377);
xor XOR2 (N8145, N8120, N4870);
buf BUF1 (N8146, N8145);
not NOT1 (N8147, N8143);
nand NAND3 (N8148, N8119, N2742, N4094);
not NOT1 (N8149, N8138);
xor XOR2 (N8150, N8147, N3707);
buf BUF1 (N8151, N8150);
nand NAND2 (N8152, N8151, N3652);
nor NOR2 (N8153, N8136, N1420);
nand NAND2 (N8154, N8153, N232);
nor NOR2 (N8155, N8141, N2257);
not NOT1 (N8156, N8152);
buf BUF1 (N8157, N8149);
or OR2 (N8158, N8146, N6246);
or OR4 (N8159, N8142, N2628, N7212, N5569);
xor XOR2 (N8160, N8157, N1391);
nand NAND3 (N8161, N8144, N5889, N5297);
nand NAND3 (N8162, N8161, N2557, N2168);
and AND2 (N8163, N8131, N1348);
xor XOR2 (N8164, N8160, N4312);
and AND2 (N8165, N8097, N6416);
xor XOR2 (N8166, N8159, N1291);
xor XOR2 (N8167, N8164, N4917);
nand NAND3 (N8168, N8162, N7543, N7732);
and AND3 (N8169, N8167, N7095, N4140);
xor XOR2 (N8170, N8169, N3088);
nor NOR2 (N8171, N8166, N6806);
or OR2 (N8172, N8155, N5347);
xor XOR2 (N8173, N8172, N6226);
or OR4 (N8174, N8170, N6256, N5296, N5429);
buf BUF1 (N8175, N8168);
or OR3 (N8176, N8154, N5105, N5230);
nand NAND2 (N8177, N8176, N6045);
not NOT1 (N8178, N8163);
xor XOR2 (N8179, N8175, N198);
not NOT1 (N8180, N8173);
nor NOR4 (N8181, N8179, N2160, N6181, N1577);
nor NOR4 (N8182, N8181, N7806, N1930, N4712);
nand NAND4 (N8183, N8180, N6315, N5854, N4299);
and AND4 (N8184, N8178, N5705, N1365, N574);
buf BUF1 (N8185, N8171);
buf BUF1 (N8186, N8165);
xor XOR2 (N8187, N8148, N5102);
xor XOR2 (N8188, N8158, N125);
not NOT1 (N8189, N8188);
or OR3 (N8190, N8184, N2253, N4912);
nand NAND3 (N8191, N8177, N3028, N4806);
nor NOR3 (N8192, N8186, N1144, N3006);
not NOT1 (N8193, N8191);
buf BUF1 (N8194, N8183);
or OR4 (N8195, N8189, N7351, N1645, N6322);
buf BUF1 (N8196, N8190);
nand NAND3 (N8197, N8193, N8081, N6551);
nor NOR2 (N8198, N8195, N6625);
xor XOR2 (N8199, N8198, N4044);
and AND4 (N8200, N8182, N3966, N3829, N5698);
or OR3 (N8201, N8196, N4438, N5516);
xor XOR2 (N8202, N8187, N4145);
buf BUF1 (N8203, N8200);
buf BUF1 (N8204, N8197);
xor XOR2 (N8205, N8202, N5641);
not NOT1 (N8206, N8174);
xor XOR2 (N8207, N8199, N6154);
buf BUF1 (N8208, N8206);
not NOT1 (N8209, N8208);
not NOT1 (N8210, N8204);
nand NAND3 (N8211, N8207, N2895, N4834);
nand NAND4 (N8212, N8205, N4839, N7445, N7731);
xor XOR2 (N8213, N8194, N899);
or OR4 (N8214, N8212, N1584, N6828, N1536);
xor XOR2 (N8215, N8213, N7238);
nand NAND3 (N8216, N8192, N6676, N5175);
nor NOR4 (N8217, N8203, N2991, N2494, N1972);
buf BUF1 (N8218, N8156);
xor XOR2 (N8219, N8215, N615);
and AND3 (N8220, N8210, N3463, N6664);
buf BUF1 (N8221, N8209);
and AND2 (N8222, N8219, N8170);
nor NOR2 (N8223, N8216, N700);
or OR2 (N8224, N8217, N1914);
and AND3 (N8225, N8211, N3680, N8061);
xor XOR2 (N8226, N8223, N4258);
nand NAND4 (N8227, N8225, N5335, N3717, N4505);
nand NAND3 (N8228, N8222, N7087, N5799);
nand NAND2 (N8229, N8185, N7947);
nand NAND3 (N8230, N8229, N2392, N2232);
or OR2 (N8231, N8220, N3799);
or OR3 (N8232, N8228, N96, N2327);
nor NOR3 (N8233, N8221, N3540, N5364);
and AND3 (N8234, N8231, N4422, N4667);
nor NOR4 (N8235, N8201, N327, N6373, N5060);
xor XOR2 (N8236, N8224, N413);
nor NOR2 (N8237, N8226, N8213);
xor XOR2 (N8238, N8227, N6654);
and AND4 (N8239, N8235, N7361, N2349, N7805);
not NOT1 (N8240, N8232);
nor NOR2 (N8241, N8233, N7992);
nand NAND3 (N8242, N8234, N1637, N7371);
nor NOR2 (N8243, N8239, N5544);
or OR3 (N8244, N8242, N883, N75);
or OR4 (N8245, N8240, N3725, N2324, N1537);
nor NOR2 (N8246, N8245, N389);
nand NAND2 (N8247, N8244, N5236);
or OR4 (N8248, N8214, N738, N3795, N1191);
not NOT1 (N8249, N8230);
nor NOR4 (N8250, N8247, N5488, N7405, N2474);
or OR4 (N8251, N8238, N5319, N3359, N5221);
buf BUF1 (N8252, N8246);
or OR2 (N8253, N8250, N3151);
and AND4 (N8254, N8251, N4430, N1659, N7241);
nand NAND4 (N8255, N8236, N2, N1351, N1119);
or OR3 (N8256, N8249, N1168, N1947);
xor XOR2 (N8257, N8243, N3990);
buf BUF1 (N8258, N8253);
or OR4 (N8259, N8248, N4112, N5932, N6889);
xor XOR2 (N8260, N8241, N298);
nand NAND4 (N8261, N8256, N2258, N4218, N1300);
buf BUF1 (N8262, N8258);
and AND2 (N8263, N8260, N355);
not NOT1 (N8264, N8257);
xor XOR2 (N8265, N8255, N8);
xor XOR2 (N8266, N8265, N5598);
nand NAND3 (N8267, N8261, N3885, N6842);
nor NOR4 (N8268, N8267, N3816, N4092, N5275);
not NOT1 (N8269, N8237);
nand NAND4 (N8270, N8264, N5685, N7512, N4447);
buf BUF1 (N8271, N8269);
not NOT1 (N8272, N8270);
nor NOR3 (N8273, N8271, N4359, N4860);
xor XOR2 (N8274, N8218, N3807);
xor XOR2 (N8275, N8252, N7437);
not NOT1 (N8276, N8268);
not NOT1 (N8277, N8276);
or OR2 (N8278, N8274, N7105);
not NOT1 (N8279, N8263);
buf BUF1 (N8280, N8279);
buf BUF1 (N8281, N8259);
and AND4 (N8282, N8281, N219, N7143, N4334);
nor NOR4 (N8283, N8254, N5590, N7344, N2088);
nor NOR3 (N8284, N8277, N7667, N442);
buf BUF1 (N8285, N8284);
buf BUF1 (N8286, N8275);
nand NAND2 (N8287, N8278, N50);
nor NOR4 (N8288, N8262, N5382, N5696, N1045);
or OR3 (N8289, N8285, N2717, N532);
not NOT1 (N8290, N8273);
xor XOR2 (N8291, N8290, N5031);
xor XOR2 (N8292, N8288, N5787);
buf BUF1 (N8293, N8280);
nand NAND4 (N8294, N8291, N7921, N6819, N661);
and AND3 (N8295, N8283, N2931, N5440);
xor XOR2 (N8296, N8282, N4690);
nor NOR4 (N8297, N8286, N7321, N5498, N6457);
nand NAND4 (N8298, N8287, N1231, N7849, N1606);
or OR2 (N8299, N8292, N1040);
nor NOR2 (N8300, N8266, N3029);
nor NOR4 (N8301, N8293, N3327, N597, N1582);
or OR2 (N8302, N8300, N6672);
buf BUF1 (N8303, N8302);
nor NOR3 (N8304, N8272, N7534, N6755);
or OR4 (N8305, N8289, N6594, N3441, N6408);
and AND3 (N8306, N8294, N5284, N6805);
xor XOR2 (N8307, N8304, N1032);
nor NOR3 (N8308, N8305, N1997, N4134);
not NOT1 (N8309, N8297);
xor XOR2 (N8310, N8295, N3115);
xor XOR2 (N8311, N8296, N1829);
nand NAND4 (N8312, N8303, N3732, N2391, N3820);
xor XOR2 (N8313, N8312, N5349);
nand NAND2 (N8314, N8311, N4709);
and AND2 (N8315, N8301, N4082);
nand NAND3 (N8316, N8315, N3673, N4708);
not NOT1 (N8317, N8299);
nor NOR3 (N8318, N8309, N2737, N1235);
nand NAND4 (N8319, N8307, N4010, N3408, N6632);
xor XOR2 (N8320, N8310, N6309);
nand NAND3 (N8321, N8308, N6880, N7327);
not NOT1 (N8322, N8321);
buf BUF1 (N8323, N8318);
buf BUF1 (N8324, N8317);
not NOT1 (N8325, N8324);
nand NAND4 (N8326, N8316, N4574, N3856, N8108);
nor NOR4 (N8327, N8298, N7570, N2752, N2017);
xor XOR2 (N8328, N8322, N2765);
not NOT1 (N8329, N8325);
and AND4 (N8330, N8329, N4041, N626, N6591);
xor XOR2 (N8331, N8328, N4450);
buf BUF1 (N8332, N8331);
and AND3 (N8333, N8319, N2153, N4663);
or OR3 (N8334, N8333, N3461, N5091);
nor NOR3 (N8335, N8330, N3568, N1511);
or OR4 (N8336, N8320, N8120, N1370, N1038);
or OR4 (N8337, N8326, N4574, N2018, N4762);
or OR3 (N8338, N8323, N1015, N7449);
and AND4 (N8339, N8306, N3595, N6682, N7350);
buf BUF1 (N8340, N8335);
nor NOR3 (N8341, N8327, N2590, N7936);
nand NAND3 (N8342, N8314, N7576, N2674);
and AND4 (N8343, N8338, N3916, N4446, N169);
nand NAND3 (N8344, N8339, N4514, N3774);
buf BUF1 (N8345, N8336);
xor XOR2 (N8346, N8313, N6615);
not NOT1 (N8347, N8340);
not NOT1 (N8348, N8334);
xor XOR2 (N8349, N8348, N5271);
not NOT1 (N8350, N8337);
nor NOR4 (N8351, N8346, N2696, N7228, N5327);
not NOT1 (N8352, N8350);
nand NAND3 (N8353, N8341, N1873, N1676);
xor XOR2 (N8354, N8352, N6380);
and AND3 (N8355, N8353, N501, N3328);
and AND3 (N8356, N8347, N5207, N8192);
nor NOR4 (N8357, N8355, N7052, N1664, N7985);
nor NOR3 (N8358, N8357, N340, N5339);
nand NAND2 (N8359, N8349, N3722);
and AND3 (N8360, N8342, N3027, N4553);
xor XOR2 (N8361, N8332, N8196);
not NOT1 (N8362, N8361);
or OR2 (N8363, N8359, N138);
or OR2 (N8364, N8356, N4614);
and AND2 (N8365, N8360, N4020);
not NOT1 (N8366, N8344);
xor XOR2 (N8367, N8366, N1813);
buf BUF1 (N8368, N8351);
or OR2 (N8369, N8364, N4874);
and AND3 (N8370, N8365, N6172, N2533);
not NOT1 (N8371, N8368);
buf BUF1 (N8372, N8369);
nor NOR4 (N8373, N8358, N6952, N4355, N174);
xor XOR2 (N8374, N8345, N6227);
buf BUF1 (N8375, N8371);
and AND4 (N8376, N8363, N7030, N5317, N2588);
nand NAND2 (N8377, N8375, N2251);
xor XOR2 (N8378, N8343, N154);
or OR2 (N8379, N8354, N3807);
buf BUF1 (N8380, N8367);
nor NOR4 (N8381, N8376, N4959, N5891, N2323);
and AND2 (N8382, N8372, N7063);
nand NAND4 (N8383, N8374, N6503, N1965, N4496);
nor NOR2 (N8384, N8362, N1372);
nand NAND3 (N8385, N8381, N2003, N7638);
xor XOR2 (N8386, N8380, N4729);
buf BUF1 (N8387, N8382);
and AND3 (N8388, N8373, N3401, N85);
not NOT1 (N8389, N8379);
or OR3 (N8390, N8386, N4517, N6527);
xor XOR2 (N8391, N8390, N10);
and AND3 (N8392, N8384, N3093, N1638);
buf BUF1 (N8393, N8377);
nand NAND2 (N8394, N8378, N4576);
buf BUF1 (N8395, N8383);
nand NAND3 (N8396, N8370, N6518, N3981);
and AND4 (N8397, N8396, N4416, N6674, N8341);
or OR3 (N8398, N8391, N6435, N3657);
xor XOR2 (N8399, N8387, N1647);
nor NOR4 (N8400, N8395, N6176, N6806, N5884);
not NOT1 (N8401, N8393);
xor XOR2 (N8402, N8389, N6347);
or OR4 (N8403, N8385, N1264, N6736, N537);
nand NAND4 (N8404, N8394, N6089, N2510, N4125);
buf BUF1 (N8405, N8402);
nor NOR4 (N8406, N8400, N2870, N3649, N8329);
and AND3 (N8407, N8405, N5458, N5682);
or OR2 (N8408, N8392, N3589);
xor XOR2 (N8409, N8406, N5494);
buf BUF1 (N8410, N8407);
xor XOR2 (N8411, N8399, N570);
or OR2 (N8412, N8398, N5340);
not NOT1 (N8413, N8411);
and AND4 (N8414, N8401, N1053, N2761, N2524);
and AND3 (N8415, N8408, N2434, N1975);
or OR2 (N8416, N8412, N7055);
xor XOR2 (N8417, N8388, N3514);
and AND2 (N8418, N8410, N3881);
nand NAND2 (N8419, N8403, N174);
or OR4 (N8420, N8413, N8018, N3042, N8009);
buf BUF1 (N8421, N8419);
buf BUF1 (N8422, N8416);
nand NAND4 (N8423, N8404, N4211, N848, N1932);
and AND3 (N8424, N8409, N7759, N312);
buf BUF1 (N8425, N8418);
nand NAND2 (N8426, N8415, N3389);
and AND3 (N8427, N8421, N5545, N5186);
or OR3 (N8428, N8425, N2592, N2749);
nor NOR3 (N8429, N8428, N6644, N1147);
and AND2 (N8430, N8417, N5609);
or OR3 (N8431, N8414, N3955, N6492);
nor NOR3 (N8432, N8427, N2382, N6308);
and AND2 (N8433, N8426, N2491);
or OR2 (N8434, N8433, N5167);
or OR4 (N8435, N8422, N2269, N6654, N4848);
or OR3 (N8436, N8430, N7337, N795);
nor NOR3 (N8437, N8424, N7689, N3245);
or OR4 (N8438, N8397, N2698, N3496, N2522);
xor XOR2 (N8439, N8437, N4963);
or OR2 (N8440, N8436, N4044);
buf BUF1 (N8441, N8429);
nand NAND3 (N8442, N8423, N46, N7778);
nor NOR4 (N8443, N8440, N1709, N1634, N4767);
buf BUF1 (N8444, N8441);
not NOT1 (N8445, N8434);
nand NAND4 (N8446, N8443, N2584, N1260, N7346);
buf BUF1 (N8447, N8438);
or OR4 (N8448, N8444, N2699, N6663, N3376);
or OR2 (N8449, N8439, N442);
and AND2 (N8450, N8432, N5825);
and AND4 (N8451, N8435, N1640, N2, N4834);
or OR4 (N8452, N8445, N7313, N4121, N669);
not NOT1 (N8453, N8451);
nor NOR4 (N8454, N8449, N2349, N7981, N2604);
not NOT1 (N8455, N8453);
nor NOR2 (N8456, N8448, N144);
nand NAND4 (N8457, N8450, N7729, N7008, N4873);
nor NOR3 (N8458, N8452, N7089, N476);
nand NAND3 (N8459, N8446, N7257, N1858);
nor NOR4 (N8460, N8458, N5127, N4129, N6783);
buf BUF1 (N8461, N8420);
or OR4 (N8462, N8454, N8061, N7926, N1885);
not NOT1 (N8463, N8431);
not NOT1 (N8464, N8447);
or OR4 (N8465, N8462, N7840, N5480, N2098);
nor NOR4 (N8466, N8463, N7672, N5956, N7854);
xor XOR2 (N8467, N8442, N7696);
buf BUF1 (N8468, N8461);
nand NAND3 (N8469, N8457, N8012, N413);
nand NAND4 (N8470, N8468, N6173, N6810, N407);
nor NOR4 (N8471, N8459, N2258, N8327, N3034);
or OR3 (N8472, N8471, N3950, N5232);
not NOT1 (N8473, N8460);
nor NOR3 (N8474, N8469, N5507, N2047);
not NOT1 (N8475, N8465);
xor XOR2 (N8476, N8464, N6065);
not NOT1 (N8477, N8470);
and AND3 (N8478, N8475, N3881, N7606);
nand NAND2 (N8479, N8473, N778);
buf BUF1 (N8480, N8455);
nor NOR4 (N8481, N8480, N6429, N3622, N1602);
nor NOR3 (N8482, N8481, N1778, N1955);
and AND2 (N8483, N8479, N5017);
buf BUF1 (N8484, N8476);
xor XOR2 (N8485, N8456, N4526);
or OR3 (N8486, N8477, N332, N2082);
nor NOR2 (N8487, N8474, N1026);
or OR4 (N8488, N8472, N959, N5721, N833);
nor NOR4 (N8489, N8483, N2214, N1269, N1256);
not NOT1 (N8490, N8485);
xor XOR2 (N8491, N8487, N7013);
nand NAND4 (N8492, N8486, N4315, N6434, N7911);
not NOT1 (N8493, N8478);
nor NOR4 (N8494, N8493, N8104, N535, N4635);
buf BUF1 (N8495, N8489);
or OR3 (N8496, N8467, N4441, N165);
not NOT1 (N8497, N8482);
nand NAND4 (N8498, N8491, N303, N6503, N904);
not NOT1 (N8499, N8484);
or OR2 (N8500, N8499, N6525);
nand NAND2 (N8501, N8500, N386);
xor XOR2 (N8502, N8498, N6382);
or OR2 (N8503, N8494, N2073);
nor NOR2 (N8504, N8497, N3100);
xor XOR2 (N8505, N8466, N6603);
and AND2 (N8506, N8488, N7342);
xor XOR2 (N8507, N8490, N1667);
nand NAND4 (N8508, N8501, N4666, N6080, N958);
xor XOR2 (N8509, N8496, N2842);
nor NOR3 (N8510, N8502, N6663, N3458);
nor NOR4 (N8511, N8492, N5431, N1740, N819);
or OR4 (N8512, N8507, N6690, N3137, N923);
nand NAND2 (N8513, N8495, N1248);
nor NOR2 (N8514, N8509, N5898);
and AND4 (N8515, N8505, N5515, N4867, N7755);
nand NAND2 (N8516, N8515, N3449);
and AND4 (N8517, N8510, N1134, N7790, N6889);
nand NAND3 (N8518, N8517, N1202, N771);
buf BUF1 (N8519, N8514);
and AND4 (N8520, N8519, N5672, N1900, N1466);
xor XOR2 (N8521, N8516, N5375);
nor NOR3 (N8522, N8520, N527, N6808);
buf BUF1 (N8523, N8512);
nand NAND2 (N8524, N8506, N1066);
not NOT1 (N8525, N8503);
nand NAND2 (N8526, N8518, N2388);
xor XOR2 (N8527, N8526, N4762);
or OR2 (N8528, N8523, N1994);
or OR3 (N8529, N8513, N2236, N392);
buf BUF1 (N8530, N8504);
and AND4 (N8531, N8525, N2149, N2714, N7619);
nor NOR4 (N8532, N8524, N6220, N4930, N4891);
not NOT1 (N8533, N8508);
or OR4 (N8534, N8530, N8289, N3322, N2323);
and AND4 (N8535, N8531, N4869, N1327, N6572);
buf BUF1 (N8536, N8532);
or OR3 (N8537, N8522, N3710, N3682);
xor XOR2 (N8538, N8535, N1742);
xor XOR2 (N8539, N8533, N5156);
nand NAND4 (N8540, N8534, N7570, N2801, N1370);
or OR4 (N8541, N8536, N3379, N4800, N984);
buf BUF1 (N8542, N8511);
buf BUF1 (N8543, N8542);
not NOT1 (N8544, N8529);
nand NAND2 (N8545, N8538, N6766);
and AND2 (N8546, N8537, N517);
not NOT1 (N8547, N8546);
not NOT1 (N8548, N8545);
xor XOR2 (N8549, N8528, N3798);
or OR4 (N8550, N8549, N5664, N562, N1630);
or OR4 (N8551, N8540, N5944, N5133, N7954);
xor XOR2 (N8552, N8544, N7662);
xor XOR2 (N8553, N8541, N7115);
or OR2 (N8554, N8548, N3974);
xor XOR2 (N8555, N8547, N7748);
not NOT1 (N8556, N8521);
and AND2 (N8557, N8556, N3985);
xor XOR2 (N8558, N8550, N1915);
nor NOR4 (N8559, N8558, N7085, N6864, N7876);
xor XOR2 (N8560, N8559, N5439);
not NOT1 (N8561, N8527);
buf BUF1 (N8562, N8543);
xor XOR2 (N8563, N8562, N7857);
xor XOR2 (N8564, N8539, N6535);
not NOT1 (N8565, N8555);
and AND4 (N8566, N8553, N4114, N179, N7036);
xor XOR2 (N8567, N8554, N258);
nand NAND2 (N8568, N8560, N3926);
buf BUF1 (N8569, N8551);
or OR4 (N8570, N8565, N6410, N828, N1067);
nand NAND2 (N8571, N8563, N7571);
xor XOR2 (N8572, N8570, N5041);
not NOT1 (N8573, N8571);
buf BUF1 (N8574, N8566);
buf BUF1 (N8575, N8567);
or OR3 (N8576, N8561, N7612, N8535);
not NOT1 (N8577, N8552);
xor XOR2 (N8578, N8569, N2765);
or OR4 (N8579, N8574, N3905, N6270, N7396);
and AND2 (N8580, N8575, N5529);
or OR2 (N8581, N8576, N8536);
or OR3 (N8582, N8579, N2952, N2335);
not NOT1 (N8583, N8577);
nand NAND4 (N8584, N8568, N6409, N1000, N2281);
buf BUF1 (N8585, N8564);
buf BUF1 (N8586, N8585);
or OR3 (N8587, N8578, N7141, N350);
or OR2 (N8588, N8557, N8173);
not NOT1 (N8589, N8573);
xor XOR2 (N8590, N8584, N139);
buf BUF1 (N8591, N8587);
xor XOR2 (N8592, N8582, N1290);
not NOT1 (N8593, N8572);
xor XOR2 (N8594, N8589, N7771);
not NOT1 (N8595, N8592);
or OR2 (N8596, N8591, N1805);
buf BUF1 (N8597, N8588);
not NOT1 (N8598, N8597);
or OR4 (N8599, N8583, N2003, N2906, N3754);
buf BUF1 (N8600, N8590);
nor NOR2 (N8601, N8596, N2782);
nor NOR4 (N8602, N8594, N1539, N7132, N3449);
or OR3 (N8603, N8599, N2808, N6043);
buf BUF1 (N8604, N8586);
nand NAND3 (N8605, N8604, N300, N6464);
not NOT1 (N8606, N8581);
not NOT1 (N8607, N8602);
or OR4 (N8608, N8600, N5375, N3928, N5471);
buf BUF1 (N8609, N8607);
buf BUF1 (N8610, N8593);
buf BUF1 (N8611, N8601);
and AND4 (N8612, N8595, N7403, N6324, N3697);
nor NOR3 (N8613, N8605, N2652, N2964);
and AND2 (N8614, N8608, N1019);
xor XOR2 (N8615, N8614, N5833);
and AND3 (N8616, N8610, N1592, N2512);
and AND4 (N8617, N8613, N3385, N7126, N435);
not NOT1 (N8618, N8611);
nand NAND2 (N8619, N8616, N1901);
buf BUF1 (N8620, N8598);
xor XOR2 (N8621, N8620, N918);
nand NAND3 (N8622, N8621, N8579, N6187);
not NOT1 (N8623, N8603);
nand NAND2 (N8624, N8609, N76);
nor NOR4 (N8625, N8624, N940, N5728, N7836);
nand NAND4 (N8626, N8612, N666, N5676, N2606);
not NOT1 (N8627, N8606);
nor NOR4 (N8628, N8580, N6984, N1666, N1753);
and AND2 (N8629, N8625, N3049);
nor NOR2 (N8630, N8615, N8371);
not NOT1 (N8631, N8626);
xor XOR2 (N8632, N8629, N6029);
or OR3 (N8633, N8627, N2076, N3511);
buf BUF1 (N8634, N8630);
xor XOR2 (N8635, N8619, N2057);
buf BUF1 (N8636, N8634);
and AND3 (N8637, N8633, N6416, N8248);
buf BUF1 (N8638, N8636);
and AND4 (N8639, N8618, N5560, N1103, N1483);
or OR4 (N8640, N8631, N4646, N3643, N2157);
or OR3 (N8641, N8640, N24, N2353);
and AND3 (N8642, N8617, N4618, N948);
nand NAND4 (N8643, N8635, N6809, N7558, N8387);
xor XOR2 (N8644, N8639, N3667);
or OR3 (N8645, N8642, N4481, N5459);
xor XOR2 (N8646, N8638, N6504);
or OR3 (N8647, N8643, N4926, N7287);
not NOT1 (N8648, N8632);
or OR3 (N8649, N8641, N2630, N946);
nor NOR4 (N8650, N8647, N1854, N3089, N8166);
xor XOR2 (N8651, N8628, N2434);
and AND4 (N8652, N8644, N7258, N7403, N3462);
nand NAND2 (N8653, N8622, N8324);
not NOT1 (N8654, N8645);
xor XOR2 (N8655, N8637, N6395);
nor NOR2 (N8656, N8623, N3634);
buf BUF1 (N8657, N8653);
not NOT1 (N8658, N8652);
not NOT1 (N8659, N8650);
nand NAND4 (N8660, N8656, N5404, N559, N5660);
nand NAND4 (N8661, N8657, N3352, N8048, N5581);
xor XOR2 (N8662, N8658, N6515);
nor NOR3 (N8663, N8646, N4716, N8425);
nand NAND2 (N8664, N8661, N4334);
nand NAND4 (N8665, N8664, N1380, N8096, N8369);
and AND2 (N8666, N8649, N76);
buf BUF1 (N8667, N8663);
xor XOR2 (N8668, N8665, N3269);
or OR4 (N8669, N8654, N3210, N3089, N5997);
not NOT1 (N8670, N8648);
or OR2 (N8671, N8669, N5347);
or OR4 (N8672, N8670, N1025, N8033, N1104);
xor XOR2 (N8673, N8671, N383);
nand NAND2 (N8674, N8651, N1537);
nand NAND3 (N8675, N8662, N813, N310);
buf BUF1 (N8676, N8673);
or OR3 (N8677, N8660, N8351, N5020);
not NOT1 (N8678, N8668);
not NOT1 (N8679, N8678);
nand NAND2 (N8680, N8679, N3799);
xor XOR2 (N8681, N8667, N1526);
or OR3 (N8682, N8655, N1533, N5103);
or OR3 (N8683, N8674, N4254, N116);
nor NOR2 (N8684, N8672, N5801);
buf BUF1 (N8685, N8683);
or OR4 (N8686, N8680, N5721, N3895, N3901);
nand NAND3 (N8687, N8686, N1478, N3820);
nand NAND4 (N8688, N8684, N2035, N7252, N5707);
not NOT1 (N8689, N8659);
nor NOR3 (N8690, N8675, N5772, N4125);
buf BUF1 (N8691, N8666);
nand NAND4 (N8692, N8676, N3052, N7357, N7328);
nand NAND3 (N8693, N8688, N7010, N3968);
and AND2 (N8694, N8690, N1205);
nor NOR2 (N8695, N8677, N7226);
and AND3 (N8696, N8693, N4792, N403);
not NOT1 (N8697, N8692);
xor XOR2 (N8698, N8695, N5479);
buf BUF1 (N8699, N8689);
buf BUF1 (N8700, N8696);
or OR3 (N8701, N8682, N3145, N1972);
nand NAND3 (N8702, N8691, N673, N5821);
not NOT1 (N8703, N8702);
xor XOR2 (N8704, N8703, N254);
or OR3 (N8705, N8697, N5742, N5984);
not NOT1 (N8706, N8700);
or OR3 (N8707, N8705, N196, N4099);
nand NAND2 (N8708, N8687, N7998);
or OR2 (N8709, N8699, N3809);
and AND3 (N8710, N8706, N6495, N7627);
xor XOR2 (N8711, N8710, N4042);
nor NOR4 (N8712, N8704, N1315, N5008, N2561);
and AND3 (N8713, N8712, N7834, N6255);
not NOT1 (N8714, N8701);
or OR2 (N8715, N8681, N7182);
or OR2 (N8716, N8713, N5153);
and AND4 (N8717, N8694, N6590, N5721, N5877);
nor NOR3 (N8718, N8698, N8635, N828);
nand NAND4 (N8719, N8707, N6900, N7439, N1684);
nor NOR4 (N8720, N8708, N2854, N4906, N5435);
nor NOR2 (N8721, N8685, N5528);
xor XOR2 (N8722, N8719, N8293);
xor XOR2 (N8723, N8722, N2209);
buf BUF1 (N8724, N8723);
nor NOR2 (N8725, N8715, N5531);
nor NOR4 (N8726, N8718, N6874, N2481, N3340);
nor NOR4 (N8727, N8717, N5792, N6395, N3456);
or OR2 (N8728, N8721, N5818);
xor XOR2 (N8729, N8726, N7231);
nor NOR4 (N8730, N8716, N7908, N2538, N1779);
xor XOR2 (N8731, N8728, N6934);
and AND3 (N8732, N8731, N4202, N1306);
not NOT1 (N8733, N8709);
buf BUF1 (N8734, N8733);
xor XOR2 (N8735, N8734, N625);
xor XOR2 (N8736, N8735, N8497);
nand NAND3 (N8737, N8711, N6767, N5004);
nor NOR3 (N8738, N8720, N491, N4375);
nor NOR3 (N8739, N8724, N1679, N5905);
nand NAND2 (N8740, N8732, N7494);
or OR4 (N8741, N8730, N4435, N3559, N6185);
buf BUF1 (N8742, N8727);
buf BUF1 (N8743, N8738);
xor XOR2 (N8744, N8736, N2157);
and AND4 (N8745, N8742, N2575, N1739, N7660);
xor XOR2 (N8746, N8729, N5797);
or OR4 (N8747, N8737, N8205, N7736, N3623);
not NOT1 (N8748, N8725);
xor XOR2 (N8749, N8746, N3054);
not NOT1 (N8750, N8747);
not NOT1 (N8751, N8750);
nand NAND3 (N8752, N8744, N8252, N81);
nand NAND3 (N8753, N8748, N7887, N4105);
or OR2 (N8754, N8739, N7220);
nand NAND2 (N8755, N8753, N2208);
nand NAND4 (N8756, N8755, N3514, N4620, N5877);
not NOT1 (N8757, N8756);
nand NAND4 (N8758, N8751, N5589, N1045, N6031);
buf BUF1 (N8759, N8752);
not NOT1 (N8760, N8749);
xor XOR2 (N8761, N8740, N4254);
xor XOR2 (N8762, N8743, N1919);
not NOT1 (N8763, N8754);
not NOT1 (N8764, N8762);
or OR3 (N8765, N8761, N5458, N2630);
xor XOR2 (N8766, N8741, N671);
and AND3 (N8767, N8764, N3811, N6544);
nand NAND3 (N8768, N8758, N3386, N4946);
or OR3 (N8769, N8745, N1896, N7725);
and AND3 (N8770, N8757, N7078, N4849);
nor NOR2 (N8771, N8765, N1067);
nand NAND4 (N8772, N8759, N8585, N524, N6880);
or OR3 (N8773, N8760, N360, N6558);
xor XOR2 (N8774, N8768, N3706);
not NOT1 (N8775, N8769);
nor NOR3 (N8776, N8767, N4725, N74);
and AND2 (N8777, N8714, N4764);
buf BUF1 (N8778, N8773);
xor XOR2 (N8779, N8776, N4420);
xor XOR2 (N8780, N8763, N3981);
not NOT1 (N8781, N8774);
or OR4 (N8782, N8781, N98, N8301, N4646);
not NOT1 (N8783, N8782);
buf BUF1 (N8784, N8783);
not NOT1 (N8785, N8772);
and AND2 (N8786, N8779, N280);
xor XOR2 (N8787, N8777, N3736);
not NOT1 (N8788, N8785);
nor NOR3 (N8789, N8766, N4678, N7181);
or OR4 (N8790, N8789, N4801, N3698, N7021);
or OR3 (N8791, N8784, N7871, N1319);
xor XOR2 (N8792, N8775, N7886);
or OR4 (N8793, N8790, N8687, N8684, N7355);
nor NOR3 (N8794, N8792, N5442, N7295);
or OR4 (N8795, N8788, N4656, N497, N6519);
nor NOR2 (N8796, N8787, N6842);
nand NAND4 (N8797, N8786, N3189, N3196, N8491);
buf BUF1 (N8798, N8795);
or OR2 (N8799, N8797, N1298);
not NOT1 (N8800, N8799);
and AND2 (N8801, N8794, N1099);
nor NOR2 (N8802, N8800, N2205);
xor XOR2 (N8803, N8793, N400);
not NOT1 (N8804, N8802);
and AND2 (N8805, N8804, N6356);
and AND3 (N8806, N8778, N6296, N3315);
nor NOR4 (N8807, N8796, N7697, N8525, N4162);
or OR2 (N8808, N8770, N3560);
nor NOR3 (N8809, N8806, N6607, N6733);
and AND4 (N8810, N8780, N3977, N8139, N7067);
nor NOR3 (N8811, N8798, N2037, N7071);
and AND4 (N8812, N8810, N1506, N7496, N3786);
nand NAND4 (N8813, N8791, N4403, N4168, N2442);
or OR2 (N8814, N8771, N2230);
nand NAND4 (N8815, N8805, N241, N5664, N5721);
buf BUF1 (N8816, N8814);
not NOT1 (N8817, N8813);
and AND4 (N8818, N8807, N3696, N1307, N1428);
nor NOR4 (N8819, N8816, N6423, N2591, N2080);
buf BUF1 (N8820, N8815);
nand NAND4 (N8821, N8811, N1337, N3075, N2672);
nor NOR4 (N8822, N8820, N5338, N7716, N1970);
xor XOR2 (N8823, N8803, N704);
nor NOR4 (N8824, N8819, N418, N8760, N8400);
buf BUF1 (N8825, N8817);
or OR3 (N8826, N8821, N8821, N4129);
nand NAND2 (N8827, N8809, N2672);
or OR4 (N8828, N8801, N8155, N6455, N6206);
nor NOR4 (N8829, N8823, N76, N5468, N3491);
xor XOR2 (N8830, N8826, N8445);
nand NAND3 (N8831, N8812, N5452, N5712);
nor NOR3 (N8832, N8829, N7695, N5301);
or OR3 (N8833, N8824, N4163, N910);
not NOT1 (N8834, N8833);
nor NOR3 (N8835, N8827, N1473, N864);
nor NOR4 (N8836, N8825, N99, N2432, N7234);
or OR3 (N8837, N8832, N5748, N7618);
buf BUF1 (N8838, N8837);
nand NAND3 (N8839, N8836, N5316, N1175);
nor NOR2 (N8840, N8822, N897);
xor XOR2 (N8841, N8831, N2895);
nor NOR2 (N8842, N8840, N8042);
buf BUF1 (N8843, N8838);
xor XOR2 (N8844, N8818, N1740);
buf BUF1 (N8845, N8841);
xor XOR2 (N8846, N8828, N5308);
xor XOR2 (N8847, N8839, N7493);
or OR4 (N8848, N8835, N4341, N8089, N7298);
and AND4 (N8849, N8848, N4106, N7319, N7065);
xor XOR2 (N8850, N8847, N8074);
not NOT1 (N8851, N8830);
nor NOR3 (N8852, N8834, N5912, N6312);
xor XOR2 (N8853, N8843, N5209);
nand NAND3 (N8854, N8808, N1974, N7240);
nand NAND4 (N8855, N8850, N387, N3785, N5340);
xor XOR2 (N8856, N8851, N2069);
buf BUF1 (N8857, N8856);
buf BUF1 (N8858, N8849);
buf BUF1 (N8859, N8857);
not NOT1 (N8860, N8842);
and AND3 (N8861, N8852, N1073, N5052);
xor XOR2 (N8862, N8860, N7811);
not NOT1 (N8863, N8846);
buf BUF1 (N8864, N8861);
not NOT1 (N8865, N8862);
nand NAND2 (N8866, N8863, N1786);
and AND4 (N8867, N8854, N7466, N4947, N1660);
not NOT1 (N8868, N8845);
not NOT1 (N8869, N8844);
and AND4 (N8870, N8865, N7487, N4148, N4418);
or OR3 (N8871, N8859, N4835, N1015);
buf BUF1 (N8872, N8867);
or OR3 (N8873, N8871, N2016, N892);
xor XOR2 (N8874, N8869, N179);
nor NOR3 (N8875, N8873, N4033, N2384);
nor NOR2 (N8876, N8866, N8021);
not NOT1 (N8877, N8855);
xor XOR2 (N8878, N8876, N1965);
not NOT1 (N8879, N8875);
buf BUF1 (N8880, N8878);
nand NAND3 (N8881, N8880, N5090, N3729);
not NOT1 (N8882, N8858);
nor NOR4 (N8883, N8853, N4, N4275, N5904);
not NOT1 (N8884, N8882);
nor NOR3 (N8885, N8879, N1162, N5758);
xor XOR2 (N8886, N8881, N4911);
not NOT1 (N8887, N8868);
buf BUF1 (N8888, N8870);
nor NOR4 (N8889, N8877, N3281, N6186, N8856);
nand NAND2 (N8890, N8884, N3695);
nand NAND4 (N8891, N8886, N2382, N5577, N7263);
not NOT1 (N8892, N8887);
and AND2 (N8893, N8872, N8853);
not NOT1 (N8894, N8888);
nor NOR3 (N8895, N8883, N7966, N4793);
nor NOR2 (N8896, N8891, N1932);
xor XOR2 (N8897, N8889, N5443);
and AND3 (N8898, N8895, N5321, N8287);
or OR4 (N8899, N8890, N6943, N7639, N8593);
not NOT1 (N8900, N8874);
nand NAND2 (N8901, N8896, N8337);
buf BUF1 (N8902, N8894);
xor XOR2 (N8903, N8893, N8745);
not NOT1 (N8904, N8897);
xor XOR2 (N8905, N8901, N2649);
not NOT1 (N8906, N8905);
nor NOR4 (N8907, N8903, N1297, N4139, N5119);
or OR2 (N8908, N8907, N44);
nor NOR4 (N8909, N8885, N4133, N4382, N3083);
buf BUF1 (N8910, N8906);
not NOT1 (N8911, N8898);
nand NAND4 (N8912, N8908, N4679, N54, N8689);
or OR4 (N8913, N8912, N3436, N1069, N6316);
nor NOR2 (N8914, N8913, N7334);
or OR2 (N8915, N8899, N5660);
xor XOR2 (N8916, N8892, N3945);
xor XOR2 (N8917, N8916, N6978);
not NOT1 (N8918, N8914);
nand NAND3 (N8919, N8902, N4641, N7955);
not NOT1 (N8920, N8917);
not NOT1 (N8921, N8918);
or OR3 (N8922, N8900, N7894, N1103);
xor XOR2 (N8923, N8915, N7554);
not NOT1 (N8924, N8921);
not NOT1 (N8925, N8922);
or OR3 (N8926, N8919, N3794, N7138);
xor XOR2 (N8927, N8925, N5044);
not NOT1 (N8928, N8923);
not NOT1 (N8929, N8926);
and AND3 (N8930, N8911, N976, N27);
nor NOR3 (N8931, N8930, N8534, N8305);
xor XOR2 (N8932, N8909, N2641);
not NOT1 (N8933, N8920);
nor NOR2 (N8934, N8924, N287);
nand NAND4 (N8935, N8934, N6517, N6821, N8677);
buf BUF1 (N8936, N8864);
and AND4 (N8937, N8932, N5356, N3095, N1322);
or OR3 (N8938, N8933, N7893, N1148);
buf BUF1 (N8939, N8929);
nor NOR2 (N8940, N8935, N7244);
not NOT1 (N8941, N8928);
and AND2 (N8942, N8937, N1320);
nor NOR4 (N8943, N8938, N545, N5287, N8224);
buf BUF1 (N8944, N8904);
nand NAND3 (N8945, N8942, N6249, N6901);
not NOT1 (N8946, N8941);
nand NAND4 (N8947, N8931, N1303, N1907, N1117);
not NOT1 (N8948, N8946);
nand NAND4 (N8949, N8939, N2577, N6479, N8109);
or OR4 (N8950, N8949, N1155, N8138, N408);
not NOT1 (N8951, N8945);
or OR2 (N8952, N8944, N2741);
xor XOR2 (N8953, N8927, N7200);
or OR3 (N8954, N8952, N1449, N5073);
or OR3 (N8955, N8910, N5529, N2803);
nor NOR3 (N8956, N8951, N1661, N401);
xor XOR2 (N8957, N8955, N6475);
nand NAND3 (N8958, N8947, N5462, N2329);
xor XOR2 (N8959, N8954, N6294);
and AND3 (N8960, N8943, N841, N7846);
or OR3 (N8961, N8940, N925, N3677);
nor NOR3 (N8962, N8958, N992, N5149);
and AND2 (N8963, N8956, N4698);
xor XOR2 (N8964, N8948, N5872);
and AND3 (N8965, N8953, N4623, N4568);
buf BUF1 (N8966, N8962);
buf BUF1 (N8967, N8965);
not NOT1 (N8968, N8959);
nor NOR2 (N8969, N8950, N7315);
buf BUF1 (N8970, N8967);
and AND4 (N8971, N8961, N8911, N5746, N1980);
nor NOR4 (N8972, N8957, N1631, N7765, N5196);
or OR3 (N8973, N8971, N8047, N47);
not NOT1 (N8974, N8964);
nand NAND4 (N8975, N8968, N458, N5626, N443);
xor XOR2 (N8976, N8960, N2539);
or OR4 (N8977, N8975, N807, N5853, N3253);
buf BUF1 (N8978, N8976);
nor NOR4 (N8979, N8963, N437, N2262, N3986);
xor XOR2 (N8980, N8969, N7230);
nand NAND4 (N8981, N8978, N6627, N3415, N2211);
nor NOR2 (N8982, N8979, N6463);
and AND3 (N8983, N8977, N366, N5159);
nand NAND3 (N8984, N8974, N8886, N2305);
buf BUF1 (N8985, N8973);
nand NAND2 (N8986, N8982, N680);
and AND3 (N8987, N8983, N8435, N1550);
buf BUF1 (N8988, N8970);
not NOT1 (N8989, N8984);
xor XOR2 (N8990, N8972, N6001);
buf BUF1 (N8991, N8986);
xor XOR2 (N8992, N8981, N5222);
or OR4 (N8993, N8991, N638, N2596, N3926);
xor XOR2 (N8994, N8990, N5049);
not NOT1 (N8995, N8989);
and AND2 (N8996, N8966, N3493);
and AND2 (N8997, N8996, N8007);
not NOT1 (N8998, N8980);
not NOT1 (N8999, N8988);
buf BUF1 (N9000, N8995);
or OR2 (N9001, N8998, N4527);
nand NAND4 (N9002, N8992, N4378, N5697, N8064);
and AND3 (N9003, N9002, N1623, N1169);
or OR2 (N9004, N9001, N5391);
not NOT1 (N9005, N8999);
and AND4 (N9006, N9003, N5334, N5604, N4809);
or OR2 (N9007, N9005, N2582);
buf BUF1 (N9008, N9006);
and AND2 (N9009, N9004, N873);
buf BUF1 (N9010, N8997);
nand NAND3 (N9011, N9007, N3046, N1335);
nand NAND2 (N9012, N8936, N5833);
nand NAND4 (N9013, N9009, N4371, N2062, N577);
nand NAND4 (N9014, N9012, N6953, N5046, N6132);
nor NOR3 (N9015, N9000, N3786, N747);
not NOT1 (N9016, N9008);
buf BUF1 (N9017, N8985);
buf BUF1 (N9018, N8994);
xor XOR2 (N9019, N9010, N136);
nor NOR2 (N9020, N9017, N5766);
not NOT1 (N9021, N9013);
xor XOR2 (N9022, N9015, N6876);
not NOT1 (N9023, N8993);
nor NOR2 (N9024, N9018, N710);
nand NAND4 (N9025, N9016, N2552, N4289, N1262);
buf BUF1 (N9026, N9014);
not NOT1 (N9027, N9020);
xor XOR2 (N9028, N9021, N6204);
xor XOR2 (N9029, N9024, N4623);
not NOT1 (N9030, N9028);
nand NAND4 (N9031, N9019, N136, N1578, N1271);
nand NAND2 (N9032, N8987, N3174);
buf BUF1 (N9033, N9025);
or OR3 (N9034, N9027, N7048, N5024);
buf BUF1 (N9035, N9032);
or OR3 (N9036, N9029, N2298, N2857);
nand NAND4 (N9037, N9034, N286, N8366, N7578);
nand NAND2 (N9038, N9033, N2786);
and AND2 (N9039, N9011, N2686);
nor NOR2 (N9040, N9038, N1359);
or OR3 (N9041, N9039, N5569, N8006);
buf BUF1 (N9042, N9040);
buf BUF1 (N9043, N9042);
nor NOR3 (N9044, N9022, N6653, N4378);
not NOT1 (N9045, N9036);
nand NAND2 (N9046, N9037, N4061);
nor NOR4 (N9047, N9026, N6446, N7176, N8297);
xor XOR2 (N9048, N9044, N2732);
and AND4 (N9049, N9047, N4510, N898, N6340);
xor XOR2 (N9050, N9030, N3231);
nand NAND2 (N9051, N9048, N6771);
nor NOR2 (N9052, N9046, N5426);
not NOT1 (N9053, N9035);
buf BUF1 (N9054, N9052);
not NOT1 (N9055, N9041);
or OR4 (N9056, N9049, N2584, N316, N2649);
nor NOR2 (N9057, N9023, N7798);
nor NOR2 (N9058, N9055, N6848);
nor NOR2 (N9059, N9054, N8917);
xor XOR2 (N9060, N9050, N5763);
nand NAND2 (N9061, N9031, N7334);
nor NOR4 (N9062, N9051, N8058, N2569, N4850);
buf BUF1 (N9063, N9053);
or OR4 (N9064, N9063, N362, N5739, N3822);
not NOT1 (N9065, N9059);
nand NAND4 (N9066, N9043, N8073, N7998, N7917);
nor NOR2 (N9067, N9066, N6336);
and AND4 (N9068, N9067, N7702, N6894, N754);
not NOT1 (N9069, N9062);
or OR3 (N9070, N9056, N2845, N2617);
buf BUF1 (N9071, N9069);
nor NOR4 (N9072, N9071, N2638, N4695, N5481);
xor XOR2 (N9073, N9045, N3525);
nor NOR3 (N9074, N9064, N6116, N3358);
and AND4 (N9075, N9061, N6675, N3951, N5178);
not NOT1 (N9076, N9065);
nor NOR3 (N9077, N9068, N6427, N2615);
nand NAND2 (N9078, N9076, N1017);
xor XOR2 (N9079, N9074, N6407);
nor NOR3 (N9080, N9077, N3644, N6888);
xor XOR2 (N9081, N9080, N3555);
and AND3 (N9082, N9060, N2855, N7433);
xor XOR2 (N9083, N9079, N3688);
buf BUF1 (N9084, N9081);
buf BUF1 (N9085, N9084);
and AND3 (N9086, N9057, N6785, N8829);
nand NAND2 (N9087, N9072, N1438);
buf BUF1 (N9088, N9083);
nor NOR4 (N9089, N9073, N7937, N4774, N4264);
nand NAND4 (N9090, N9082, N1004, N8403, N7811);
not NOT1 (N9091, N9087);
nand NAND4 (N9092, N9075, N6502, N3636, N4883);
or OR2 (N9093, N9058, N3737);
nor NOR4 (N9094, N9089, N1105, N7719, N8620);
and AND2 (N9095, N9086, N5012);
or OR4 (N9096, N9095, N3472, N4390, N524);
xor XOR2 (N9097, N9078, N7508);
nor NOR4 (N9098, N9088, N7284, N1458, N6821);
and AND4 (N9099, N9094, N5692, N1024, N1467);
not NOT1 (N9100, N9070);
buf BUF1 (N9101, N9091);
buf BUF1 (N9102, N9101);
nor NOR4 (N9103, N9100, N3421, N8780, N1772);
nor NOR2 (N9104, N9103, N6478);
xor XOR2 (N9105, N9092, N8923);
xor XOR2 (N9106, N9104, N2004);
buf BUF1 (N9107, N9099);
or OR4 (N9108, N9102, N7486, N1285, N8458);
and AND3 (N9109, N9085, N8023, N6113);
nand NAND3 (N9110, N9093, N3305, N3660);
buf BUF1 (N9111, N9106);
nand NAND2 (N9112, N9110, N6457);
not NOT1 (N9113, N9109);
xor XOR2 (N9114, N9105, N3594);
buf BUF1 (N9115, N9113);
buf BUF1 (N9116, N9108);
xor XOR2 (N9117, N9112, N2322);
nand NAND2 (N9118, N9111, N647);
buf BUF1 (N9119, N9096);
or OR2 (N9120, N9114, N2386);
and AND3 (N9121, N9097, N4064, N8386);
and AND2 (N9122, N9118, N8559);
xor XOR2 (N9123, N9122, N4560);
nand NAND2 (N9124, N9123, N5256);
or OR3 (N9125, N9117, N7834, N4);
xor XOR2 (N9126, N9107, N4907);
or OR4 (N9127, N9116, N5617, N4876, N670);
not NOT1 (N9128, N9120);
xor XOR2 (N9129, N9127, N1213);
or OR2 (N9130, N9124, N8870);
nand NAND4 (N9131, N9128, N173, N7708, N352);
xor XOR2 (N9132, N9121, N2927);
buf BUF1 (N9133, N9125);
nor NOR4 (N9134, N9132, N6604, N3402, N4132);
or OR4 (N9135, N9126, N4447, N8092, N6361);
xor XOR2 (N9136, N9130, N5101);
or OR2 (N9137, N9115, N7514);
and AND4 (N9138, N9098, N1988, N5680, N20);
xor XOR2 (N9139, N9129, N4473);
xor XOR2 (N9140, N9133, N6908);
xor XOR2 (N9141, N9138, N8371);
nand NAND4 (N9142, N9119, N634, N3875, N7848);
or OR4 (N9143, N9137, N1308, N420, N3037);
or OR2 (N9144, N9141, N2591);
not NOT1 (N9145, N9142);
buf BUF1 (N9146, N9139);
xor XOR2 (N9147, N9144, N1491);
nor NOR2 (N9148, N9146, N8842);
and AND4 (N9149, N9090, N327, N3256, N223);
buf BUF1 (N9150, N9143);
nand NAND3 (N9151, N9131, N8987, N4020);
and AND3 (N9152, N9151, N3679, N7210);
xor XOR2 (N9153, N9149, N7691);
and AND3 (N9154, N9136, N7502, N1318);
nand NAND4 (N9155, N9145, N6343, N7173, N1841);
nor NOR3 (N9156, N9140, N4171, N6447);
nor NOR3 (N9157, N9153, N3960, N6936);
nand NAND3 (N9158, N9155, N5595, N5773);
xor XOR2 (N9159, N9150, N2095);
nor NOR3 (N9160, N9135, N4724, N3978);
buf BUF1 (N9161, N9148);
or OR4 (N9162, N9161, N548, N660, N8491);
nor NOR2 (N9163, N9157, N7558);
nor NOR4 (N9164, N9152, N8320, N2718, N899);
and AND3 (N9165, N9147, N6937, N4398);
nor NOR3 (N9166, N9156, N2577, N7700);
and AND3 (N9167, N9160, N3504, N3129);
and AND3 (N9168, N9159, N3762, N7396);
and AND4 (N9169, N9154, N959, N1748, N4571);
not NOT1 (N9170, N9158);
buf BUF1 (N9171, N9165);
and AND4 (N9172, N9168, N8585, N8769, N2986);
not NOT1 (N9173, N9172);
buf BUF1 (N9174, N9171);
not NOT1 (N9175, N9164);
xor XOR2 (N9176, N9163, N499);
nand NAND3 (N9177, N9134, N1900, N8906);
nor NOR2 (N9178, N9177, N7935);
not NOT1 (N9179, N9174);
or OR3 (N9180, N9173, N2239, N411);
xor XOR2 (N9181, N9162, N8016);
and AND2 (N9182, N9176, N234);
not NOT1 (N9183, N9180);
or OR3 (N9184, N9169, N7607, N3611);
or OR3 (N9185, N9183, N7543, N226);
and AND4 (N9186, N9179, N6298, N650, N1463);
or OR2 (N9187, N9182, N5347);
nand NAND3 (N9188, N9184, N2474, N7378);
nor NOR3 (N9189, N9178, N5942, N7175);
xor XOR2 (N9190, N9188, N4259);
or OR4 (N9191, N9190, N7229, N2720, N5282);
or OR3 (N9192, N9186, N7985, N4033);
not NOT1 (N9193, N9187);
nor NOR4 (N9194, N9191, N7291, N1683, N2652);
xor XOR2 (N9195, N9181, N2387);
or OR4 (N9196, N9192, N7620, N8132, N5476);
buf BUF1 (N9197, N9185);
not NOT1 (N9198, N9175);
nor NOR4 (N9199, N9166, N6644, N1628, N7820);
xor XOR2 (N9200, N9170, N3641);
buf BUF1 (N9201, N9193);
not NOT1 (N9202, N9194);
buf BUF1 (N9203, N9197);
xor XOR2 (N9204, N9201, N7136);
nor NOR3 (N9205, N9189, N652, N323);
buf BUF1 (N9206, N9203);
not NOT1 (N9207, N9199);
nor NOR2 (N9208, N9167, N2007);
xor XOR2 (N9209, N9205, N1742);
nor NOR3 (N9210, N9196, N20, N5784);
and AND2 (N9211, N9198, N90);
nand NAND3 (N9212, N9195, N296, N3367);
and AND3 (N9213, N9211, N1815, N8998);
not NOT1 (N9214, N9212);
xor XOR2 (N9215, N9209, N8163);
or OR2 (N9216, N9202, N5146);
or OR4 (N9217, N9216, N957, N2473, N506);
and AND3 (N9218, N9215, N3123, N3276);
or OR4 (N9219, N9214, N8615, N1140, N4331);
and AND2 (N9220, N9207, N1283);
buf BUF1 (N9221, N9220);
and AND4 (N9222, N9221, N7825, N8372, N5079);
xor XOR2 (N9223, N9217, N2934);
and AND2 (N9224, N9200, N4894);
or OR3 (N9225, N9224, N1914, N2665);
xor XOR2 (N9226, N9204, N8124);
not NOT1 (N9227, N9206);
xor XOR2 (N9228, N9210, N8189);
not NOT1 (N9229, N9223);
or OR3 (N9230, N9227, N7898, N7533);
xor XOR2 (N9231, N9226, N5368);
xor XOR2 (N9232, N9231, N5369);
and AND2 (N9233, N9222, N2143);
nor NOR3 (N9234, N9228, N3598, N849);
and AND2 (N9235, N9225, N271);
and AND3 (N9236, N9219, N1657, N8645);
nor NOR3 (N9237, N9236, N3386, N6582);
not NOT1 (N9238, N9232);
xor XOR2 (N9239, N9237, N8823);
buf BUF1 (N9240, N9230);
or OR3 (N9241, N9238, N1115, N5641);
or OR4 (N9242, N9234, N1538, N4749, N7799);
or OR3 (N9243, N9240, N167, N7532);
and AND3 (N9244, N9229, N3763, N316);
or OR4 (N9245, N9243, N6055, N8243, N6541);
buf BUF1 (N9246, N9245);
xor XOR2 (N9247, N9241, N6665);
not NOT1 (N9248, N9244);
nor NOR4 (N9249, N9247, N6442, N7185, N8823);
nand NAND2 (N9250, N9208, N4655);
xor XOR2 (N9251, N9218, N6100);
nor NOR4 (N9252, N9248, N8075, N6379, N6225);
not NOT1 (N9253, N9239);
not NOT1 (N9254, N9235);
and AND2 (N9255, N9249, N4854);
nand NAND3 (N9256, N9254, N2431, N4284);
xor XOR2 (N9257, N9253, N5697);
buf BUF1 (N9258, N9256);
and AND3 (N9259, N9233, N8197, N519);
or OR2 (N9260, N9255, N4056);
nand NAND4 (N9261, N9252, N7949, N6941, N7750);
or OR4 (N9262, N9258, N3813, N161, N8505);
and AND4 (N9263, N9250, N5007, N1978, N392);
nand NAND4 (N9264, N9263, N8331, N1102, N3616);
nor NOR4 (N9265, N9257, N8220, N5310, N5799);
not NOT1 (N9266, N9260);
xor XOR2 (N9267, N9264, N3457);
or OR2 (N9268, N9267, N6416);
nor NOR2 (N9269, N9259, N4779);
nand NAND2 (N9270, N9251, N4662);
and AND4 (N9271, N9268, N7727, N798, N8415);
nand NAND2 (N9272, N9266, N6912);
buf BUF1 (N9273, N9269);
and AND2 (N9274, N9265, N8515);
and AND2 (N9275, N9213, N1951);
nand NAND4 (N9276, N9274, N3333, N2952, N1177);
and AND3 (N9277, N9273, N4182, N3216);
xor XOR2 (N9278, N9261, N22);
or OR4 (N9279, N9271, N397, N1909, N1970);
nor NOR4 (N9280, N9279, N3315, N8961, N7907);
and AND2 (N9281, N9280, N4149);
nor NOR4 (N9282, N9275, N1816, N174, N1529);
buf BUF1 (N9283, N9276);
or OR4 (N9284, N9281, N2066, N1611, N8910);
not NOT1 (N9285, N9277);
or OR3 (N9286, N9283, N6016, N5040);
nand NAND3 (N9287, N9286, N3219, N638);
or OR3 (N9288, N9282, N1820, N1110);
not NOT1 (N9289, N9287);
nor NOR4 (N9290, N9285, N4356, N3607, N6340);
or OR4 (N9291, N9289, N4944, N1297, N3059);
nand NAND3 (N9292, N9270, N4937, N8702);
or OR3 (N9293, N9288, N8470, N5418);
and AND3 (N9294, N9242, N896, N785);
not NOT1 (N9295, N9272);
nand NAND4 (N9296, N9262, N7137, N7986, N4740);
nand NAND4 (N9297, N9295, N6052, N3400, N1590);
and AND4 (N9298, N9294, N8340, N4628, N1614);
or OR2 (N9299, N9292, N4564);
nor NOR2 (N9300, N9298, N733);
or OR3 (N9301, N9299, N3973, N6228);
nor NOR2 (N9302, N9284, N6025);
and AND2 (N9303, N9291, N2158);
and AND3 (N9304, N9302, N4749, N8031);
buf BUF1 (N9305, N9278);
nor NOR2 (N9306, N9301, N5095);
nand NAND4 (N9307, N9246, N4256, N5059, N5581);
not NOT1 (N9308, N9296);
nor NOR2 (N9309, N9293, N760);
xor XOR2 (N9310, N9290, N3884);
xor XOR2 (N9311, N9300, N8832);
and AND3 (N9312, N9304, N1045, N5161);
or OR2 (N9313, N9303, N5185);
not NOT1 (N9314, N9312);
or OR2 (N9315, N9313, N411);
or OR3 (N9316, N9314, N7872, N2881);
buf BUF1 (N9317, N9311);
buf BUF1 (N9318, N9309);
nand NAND3 (N9319, N9316, N9092, N4912);
or OR3 (N9320, N9317, N3257, N6278);
nor NOR3 (N9321, N9320, N3963, N2538);
buf BUF1 (N9322, N9318);
buf BUF1 (N9323, N9297);
nand NAND3 (N9324, N9306, N2737, N150);
and AND3 (N9325, N9322, N3461, N4987);
buf BUF1 (N9326, N9305);
not NOT1 (N9327, N9325);
not NOT1 (N9328, N9321);
nand NAND3 (N9329, N9308, N4536, N4750);
nor NOR3 (N9330, N9329, N1202, N8071);
nor NOR2 (N9331, N9307, N5456);
or OR4 (N9332, N9331, N8687, N6239, N5011);
and AND3 (N9333, N9326, N6085, N1309);
and AND3 (N9334, N9324, N9201, N25);
not NOT1 (N9335, N9310);
or OR2 (N9336, N9328, N443);
and AND3 (N9337, N9327, N3283, N2193);
xor XOR2 (N9338, N9330, N1261);
nand NAND4 (N9339, N9334, N561, N3486, N3256);
xor XOR2 (N9340, N9315, N4388);
and AND4 (N9341, N9335, N9313, N3850, N2201);
nand NAND3 (N9342, N9332, N4198, N3197);
nand NAND4 (N9343, N9319, N4359, N542, N2048);
nand NAND2 (N9344, N9338, N2466);
nor NOR3 (N9345, N9342, N1475, N5593);
nor NOR3 (N9346, N9345, N5373, N8230);
buf BUF1 (N9347, N9323);
and AND4 (N9348, N9343, N8477, N7017, N9155);
and AND4 (N9349, N9339, N500, N3934, N4477);
or OR2 (N9350, N9349, N1888);
and AND3 (N9351, N9344, N4230, N3525);
not NOT1 (N9352, N9336);
not NOT1 (N9353, N9352);
nand NAND2 (N9354, N9348, N5707);
not NOT1 (N9355, N9350);
buf BUF1 (N9356, N9353);
nand NAND2 (N9357, N9347, N8893);
not NOT1 (N9358, N9346);
or OR2 (N9359, N9356, N8796);
nor NOR3 (N9360, N9354, N2543, N6374);
nand NAND3 (N9361, N9358, N6396, N2071);
buf BUF1 (N9362, N9337);
nand NAND2 (N9363, N9341, N1198);
nor NOR3 (N9364, N9355, N1914, N897);
not NOT1 (N9365, N9361);
xor XOR2 (N9366, N9340, N5505);
nor NOR4 (N9367, N9351, N6439, N5098, N6861);
or OR4 (N9368, N9360, N2892, N5856, N426);
or OR2 (N9369, N9366, N518);
nand NAND4 (N9370, N9359, N8986, N5730, N2860);
buf BUF1 (N9371, N9368);
not NOT1 (N9372, N9357);
nor NOR4 (N9373, N9367, N7983, N5240, N7195);
or OR4 (N9374, N9370, N4326, N4475, N8898);
nor NOR3 (N9375, N9372, N8264, N1470);
not NOT1 (N9376, N9374);
xor XOR2 (N9377, N9371, N7239);
nand NAND2 (N9378, N9375, N3641);
nor NOR3 (N9379, N9377, N7386, N676);
nand NAND3 (N9380, N9333, N7910, N6450);
or OR4 (N9381, N9365, N475, N3120, N3518);
xor XOR2 (N9382, N9362, N9147);
and AND3 (N9383, N9364, N6448, N6131);
not NOT1 (N9384, N9369);
buf BUF1 (N9385, N9380);
xor XOR2 (N9386, N9385, N8774);
nand NAND2 (N9387, N9376, N4305);
buf BUF1 (N9388, N9378);
or OR2 (N9389, N9384, N5864);
buf BUF1 (N9390, N9389);
or OR3 (N9391, N9382, N6049, N5589);
nor NOR4 (N9392, N9381, N8947, N2532, N2393);
nor NOR4 (N9393, N9392, N1888, N4362, N2847);
or OR2 (N9394, N9391, N1958);
buf BUF1 (N9395, N9388);
buf BUF1 (N9396, N9373);
xor XOR2 (N9397, N9383, N5138);
nor NOR2 (N9398, N9386, N6010);
and AND3 (N9399, N9394, N6931, N3846);
buf BUF1 (N9400, N9379);
and AND4 (N9401, N9393, N2487, N7497, N7594);
nand NAND4 (N9402, N9390, N2680, N8976, N6210);
and AND4 (N9403, N9402, N606, N974, N6287);
buf BUF1 (N9404, N9397);
not NOT1 (N9405, N9401);
xor XOR2 (N9406, N9395, N2430);
nand NAND2 (N9407, N9396, N4109);
or OR2 (N9408, N9387, N2008);
xor XOR2 (N9409, N9399, N8973);
or OR2 (N9410, N9400, N142);
or OR4 (N9411, N9398, N6609, N461, N2790);
xor XOR2 (N9412, N9405, N939);
nor NOR3 (N9413, N9403, N7714, N8997);
xor XOR2 (N9414, N9413, N6397);
buf BUF1 (N9415, N9408);
buf BUF1 (N9416, N9410);
not NOT1 (N9417, N9409);
nor NOR4 (N9418, N9407, N1848, N5298, N7894);
not NOT1 (N9419, N9412);
or OR2 (N9420, N9404, N2076);
buf BUF1 (N9421, N9418);
not NOT1 (N9422, N9419);
xor XOR2 (N9423, N9363, N6612);
xor XOR2 (N9424, N9411, N3272);
not NOT1 (N9425, N9417);
nand NAND2 (N9426, N9420, N8314);
not NOT1 (N9427, N9426);
and AND3 (N9428, N9406, N1060, N4997);
not NOT1 (N9429, N9424);
buf BUF1 (N9430, N9415);
xor XOR2 (N9431, N9423, N5841);
not NOT1 (N9432, N9429);
not NOT1 (N9433, N9431);
and AND3 (N9434, N9427, N647, N8695);
buf BUF1 (N9435, N9428);
buf BUF1 (N9436, N9433);
or OR4 (N9437, N9432, N1859, N852, N4549);
buf BUF1 (N9438, N9430);
and AND3 (N9439, N9422, N6738, N5223);
and AND3 (N9440, N9434, N3971, N380);
nor NOR4 (N9441, N9439, N7334, N6453, N6179);
not NOT1 (N9442, N9421);
buf BUF1 (N9443, N9442);
not NOT1 (N9444, N9441);
xor XOR2 (N9445, N9438, N8319);
buf BUF1 (N9446, N9444);
nor NOR4 (N9447, N9443, N2745, N5292, N2803);
not NOT1 (N9448, N9440);
and AND4 (N9449, N9447, N8707, N9268, N4920);
buf BUF1 (N9450, N9437);
xor XOR2 (N9451, N9449, N7765);
nand NAND3 (N9452, N9448, N5423, N7107);
or OR2 (N9453, N9425, N8258);
not NOT1 (N9454, N9450);
or OR4 (N9455, N9445, N4031, N4509, N6666);
not NOT1 (N9456, N9446);
xor XOR2 (N9457, N9455, N6981);
not NOT1 (N9458, N9414);
xor XOR2 (N9459, N9436, N8487);
nor NOR4 (N9460, N9451, N4702, N1529, N4903);
xor XOR2 (N9461, N9460, N376);
nand NAND3 (N9462, N9453, N5561, N6806);
nand NAND4 (N9463, N9452, N7577, N2789, N4150);
or OR2 (N9464, N9461, N1486);
nor NOR4 (N9465, N9463, N3085, N7613, N8966);
or OR3 (N9466, N9459, N1744, N4933);
nand NAND3 (N9467, N9457, N8640, N4909);
nor NOR4 (N9468, N9467, N3754, N3630, N7148);
nor NOR3 (N9469, N9465, N7996, N6418);
nor NOR3 (N9470, N9416, N1974, N8790);
buf BUF1 (N9471, N9469);
not NOT1 (N9472, N9471);
xor XOR2 (N9473, N9470, N4491);
buf BUF1 (N9474, N9435);
nand NAND3 (N9475, N9468, N2027, N7076);
or OR4 (N9476, N9472, N8892, N8964, N3298);
buf BUF1 (N9477, N9474);
nand NAND4 (N9478, N9464, N39, N4351, N698);
and AND2 (N9479, N9458, N1577);
or OR3 (N9480, N9456, N9395, N3055);
and AND2 (N9481, N9473, N201);
not NOT1 (N9482, N9479);
nand NAND3 (N9483, N9466, N2841, N3999);
buf BUF1 (N9484, N9481);
buf BUF1 (N9485, N9462);
buf BUF1 (N9486, N9483);
xor XOR2 (N9487, N9454, N3069);
buf BUF1 (N9488, N9482);
not NOT1 (N9489, N9487);
not NOT1 (N9490, N9488);
nand NAND3 (N9491, N9480, N4827, N7848);
nand NAND2 (N9492, N9478, N4790);
xor XOR2 (N9493, N9486, N6198);
not NOT1 (N9494, N9493);
and AND3 (N9495, N9494, N6989, N6003);
not NOT1 (N9496, N9489);
nand NAND2 (N9497, N9477, N3526);
buf BUF1 (N9498, N9490);
not NOT1 (N9499, N9495);
not NOT1 (N9500, N9476);
buf BUF1 (N9501, N9497);
nand NAND3 (N9502, N9485, N4655, N8864);
buf BUF1 (N9503, N9491);
xor XOR2 (N9504, N9492, N8527);
xor XOR2 (N9505, N9501, N8202);
and AND2 (N9506, N9475, N240);
not NOT1 (N9507, N9496);
nor NOR3 (N9508, N9498, N6778, N1091);
or OR3 (N9509, N9503, N4037, N6633);
nand NAND4 (N9510, N9504, N7858, N6507, N1615);
nor NOR3 (N9511, N9510, N4252, N7430);
not NOT1 (N9512, N9499);
buf BUF1 (N9513, N9502);
not NOT1 (N9514, N9500);
and AND2 (N9515, N9513, N1859);
not NOT1 (N9516, N9505);
and AND3 (N9517, N9511, N1800, N1527);
and AND4 (N9518, N9512, N7299, N6157, N1982);
buf BUF1 (N9519, N9516);
nand NAND2 (N9520, N9514, N9318);
buf BUF1 (N9521, N9515);
nor NOR4 (N9522, N9508, N6533, N4854, N7215);
and AND4 (N9523, N9518, N4499, N6279, N2056);
nor NOR2 (N9524, N9520, N3737);
not NOT1 (N9525, N9524);
nor NOR4 (N9526, N9509, N8262, N4699, N3178);
nor NOR2 (N9527, N9506, N2544);
not NOT1 (N9528, N9526);
nor NOR3 (N9529, N9517, N5852, N4307);
xor XOR2 (N9530, N9525, N2426);
not NOT1 (N9531, N9519);
xor XOR2 (N9532, N9527, N5736);
not NOT1 (N9533, N9522);
nand NAND4 (N9534, N9533, N8522, N3833, N7809);
not NOT1 (N9535, N9530);
nor NOR2 (N9536, N9529, N4310);
or OR3 (N9537, N9528, N3365, N2);
xor XOR2 (N9538, N9536, N5350);
buf BUF1 (N9539, N9534);
not NOT1 (N9540, N9523);
xor XOR2 (N9541, N9531, N4169);
not NOT1 (N9542, N9537);
and AND2 (N9543, N9538, N6988);
buf BUF1 (N9544, N9507);
buf BUF1 (N9545, N9541);
or OR2 (N9546, N9543, N7640);
xor XOR2 (N9547, N9539, N4205);
and AND4 (N9548, N9545, N3423, N3857, N3301);
and AND3 (N9549, N9540, N1180, N2039);
nor NOR3 (N9550, N9548, N5644, N2962);
or OR4 (N9551, N9544, N23, N6369, N9532);
buf BUF1 (N9552, N7741);
not NOT1 (N9553, N9550);
xor XOR2 (N9554, N9546, N3173);
not NOT1 (N9555, N9535);
not NOT1 (N9556, N9549);
and AND2 (N9557, N9556, N978);
nor NOR2 (N9558, N9553, N9524);
nor NOR2 (N9559, N9547, N319);
buf BUF1 (N9560, N9555);
buf BUF1 (N9561, N9521);
buf BUF1 (N9562, N9542);
not NOT1 (N9563, N9557);
and AND4 (N9564, N9562, N653, N321, N7816);
nor NOR3 (N9565, N9560, N5996, N5673);
not NOT1 (N9566, N9554);
or OR4 (N9567, N9552, N5784, N1853, N8023);
or OR3 (N9568, N9567, N6742, N3255);
or OR4 (N9569, N9561, N6302, N5205, N6711);
nor NOR4 (N9570, N9566, N9145, N5250, N5464);
and AND3 (N9571, N9565, N1704, N9323);
and AND3 (N9572, N9559, N3128, N2269);
and AND3 (N9573, N9568, N9493, N1527);
nor NOR2 (N9574, N9571, N2953);
nand NAND3 (N9575, N9569, N8939, N545);
or OR4 (N9576, N9574, N6089, N5158, N4485);
buf BUF1 (N9577, N9575);
nor NOR4 (N9578, N9577, N1332, N2885, N9502);
xor XOR2 (N9579, N9484, N7565);
nor NOR3 (N9580, N9551, N9063, N5808);
or OR3 (N9581, N9564, N637, N7710);
or OR3 (N9582, N9572, N339, N3109);
nor NOR3 (N9583, N9582, N3887, N8012);
not NOT1 (N9584, N9570);
nor NOR3 (N9585, N9581, N6813, N7);
and AND2 (N9586, N9563, N4978);
and AND4 (N9587, N9585, N8627, N9414, N1510);
nand NAND4 (N9588, N9587, N5658, N8957, N988);
nor NOR4 (N9589, N9583, N6806, N533, N3270);
not NOT1 (N9590, N9580);
nand NAND3 (N9591, N9589, N5693, N1514);
nor NOR4 (N9592, N9588, N3038, N9424, N4085);
and AND3 (N9593, N9578, N5468, N9255);
nor NOR3 (N9594, N9558, N2475, N5349);
nand NAND3 (N9595, N9590, N277, N9464);
buf BUF1 (N9596, N9594);
nor NOR2 (N9597, N9586, N2086);
or OR2 (N9598, N9584, N365);
and AND4 (N9599, N9593, N7388, N7732, N4905);
nand NAND4 (N9600, N9597, N1671, N8702, N7474);
nand NAND4 (N9601, N9595, N3296, N5019, N2793);
nand NAND4 (N9602, N9599, N4564, N4749, N873);
nand NAND4 (N9603, N9592, N730, N9053, N8814);
xor XOR2 (N9604, N9579, N8763);
and AND3 (N9605, N9596, N7233, N52);
xor XOR2 (N9606, N9600, N3452);
not NOT1 (N9607, N9605);
buf BUF1 (N9608, N9602);
not NOT1 (N9609, N9603);
nor NOR4 (N9610, N9608, N8254, N205, N4295);
and AND2 (N9611, N9606, N127);
nand NAND2 (N9612, N9601, N5939);
or OR3 (N9613, N9611, N8684, N7624);
buf BUF1 (N9614, N9609);
xor XOR2 (N9615, N9576, N7497);
nor NOR2 (N9616, N9573, N3993);
xor XOR2 (N9617, N9613, N5443);
nand NAND4 (N9618, N9617, N4950, N102, N5696);
or OR4 (N9619, N9616, N865, N3640, N2040);
nand NAND4 (N9620, N9615, N5606, N4642, N3157);
nor NOR4 (N9621, N9610, N3269, N6693, N271);
buf BUF1 (N9622, N9621);
xor XOR2 (N9623, N9622, N9003);
xor XOR2 (N9624, N9612, N7835);
and AND4 (N9625, N9598, N476, N542, N7867);
buf BUF1 (N9626, N9625);
or OR4 (N9627, N9591, N3502, N7667, N7157);
nand NAND4 (N9628, N9623, N2469, N1530, N3471);
nand NAND2 (N9629, N9619, N8495);
buf BUF1 (N9630, N9614);
buf BUF1 (N9631, N9607);
nor NOR3 (N9632, N9630, N5192, N7260);
and AND2 (N9633, N9631, N9377);
nand NAND4 (N9634, N9632, N4757, N7427, N5098);
not NOT1 (N9635, N9627);
nor NOR3 (N9636, N9624, N4165, N7307);
nor NOR4 (N9637, N9636, N2560, N779, N2254);
not NOT1 (N9638, N9634);
nand NAND3 (N9639, N9637, N9331, N3885);
not NOT1 (N9640, N9635);
not NOT1 (N9641, N9626);
xor XOR2 (N9642, N9641, N6338);
and AND2 (N9643, N9618, N5318);
and AND3 (N9644, N9629, N1327, N3777);
nand NAND4 (N9645, N9638, N6003, N6842, N4148);
nand NAND2 (N9646, N9640, N5670);
buf BUF1 (N9647, N9639);
xor XOR2 (N9648, N9643, N6147);
or OR3 (N9649, N9645, N5809, N7096);
and AND2 (N9650, N9644, N8045);
not NOT1 (N9651, N9633);
buf BUF1 (N9652, N9649);
buf BUF1 (N9653, N9651);
nand NAND3 (N9654, N9642, N7944, N7557);
nor NOR3 (N9655, N9628, N535, N1618);
or OR3 (N9656, N9654, N5652, N1935);
nor NOR2 (N9657, N9653, N3801);
or OR2 (N9658, N9656, N2804);
not NOT1 (N9659, N9604);
nand NAND4 (N9660, N9652, N7200, N2687, N8953);
not NOT1 (N9661, N9646);
not NOT1 (N9662, N9661);
nor NOR4 (N9663, N9660, N7427, N9343, N7632);
xor XOR2 (N9664, N9620, N3479);
nor NOR4 (N9665, N9648, N3181, N7285, N460);
and AND4 (N9666, N9662, N8823, N3473, N331);
nand NAND3 (N9667, N9658, N7351, N6489);
nand NAND4 (N9668, N9664, N6781, N7032, N5246);
buf BUF1 (N9669, N9668);
xor XOR2 (N9670, N9657, N1482);
xor XOR2 (N9671, N9669, N6078);
buf BUF1 (N9672, N9659);
or OR3 (N9673, N9670, N9582, N1233);
not NOT1 (N9674, N9650);
buf BUF1 (N9675, N9674);
buf BUF1 (N9676, N9665);
not NOT1 (N9677, N9663);
xor XOR2 (N9678, N9655, N1595);
not NOT1 (N9679, N9676);
xor XOR2 (N9680, N9671, N1560);
nor NOR2 (N9681, N9673, N6168);
nor NOR4 (N9682, N9675, N8500, N8027, N4126);
nor NOR2 (N9683, N9682, N4308);
nor NOR3 (N9684, N9683, N6921, N1704);
xor XOR2 (N9685, N9667, N234);
nor NOR2 (N9686, N9672, N7658);
buf BUF1 (N9687, N9647);
buf BUF1 (N9688, N9679);
nor NOR2 (N9689, N9680, N5762);
nor NOR4 (N9690, N9666, N7502, N5336, N3396);
buf BUF1 (N9691, N9678);
not NOT1 (N9692, N9691);
nor NOR2 (N9693, N9689, N2845);
nand NAND2 (N9694, N9681, N8957);
and AND2 (N9695, N9693, N1989);
nand NAND3 (N9696, N9694, N2809, N286);
not NOT1 (N9697, N9686);
and AND2 (N9698, N9685, N9427);
or OR2 (N9699, N9697, N7276);
and AND4 (N9700, N9690, N3165, N5109, N171);
nand NAND2 (N9701, N9684, N4203);
not NOT1 (N9702, N9695);
not NOT1 (N9703, N9699);
and AND3 (N9704, N9687, N207, N9339);
not NOT1 (N9705, N9702);
and AND3 (N9706, N9701, N9226, N1573);
nand NAND4 (N9707, N9706, N3431, N9430, N7911);
buf BUF1 (N9708, N9707);
not NOT1 (N9709, N9708);
and AND2 (N9710, N9677, N4841);
not NOT1 (N9711, N9704);
or OR4 (N9712, N9709, N4323, N3659, N2057);
and AND2 (N9713, N9712, N9496);
xor XOR2 (N9714, N9692, N9250);
nand NAND2 (N9715, N9711, N2978);
nor NOR4 (N9716, N9713, N1486, N8832, N2826);
nor NOR4 (N9717, N9696, N9716, N5008, N4762);
buf BUF1 (N9718, N605);
buf BUF1 (N9719, N9705);
and AND2 (N9720, N9719, N7713);
nand NAND4 (N9721, N9688, N2831, N9453, N9676);
buf BUF1 (N9722, N9714);
and AND3 (N9723, N9718, N5045, N9299);
and AND4 (N9724, N9723, N7125, N6785, N6389);
nor NOR3 (N9725, N9700, N2226, N7578);
xor XOR2 (N9726, N9717, N4722);
nor NOR3 (N9727, N9720, N9138, N4683);
nand NAND2 (N9728, N9721, N6077);
and AND4 (N9729, N9703, N7833, N2522, N1122);
xor XOR2 (N9730, N9727, N8300);
and AND4 (N9731, N9698, N4754, N7448, N447);
nand NAND4 (N9732, N9728, N2057, N5258, N3788);
or OR2 (N9733, N9729, N9353);
not NOT1 (N9734, N9730);
nor NOR4 (N9735, N9715, N5459, N1082, N6800);
xor XOR2 (N9736, N9724, N5449);
buf BUF1 (N9737, N9731);
and AND2 (N9738, N9710, N2568);
nor NOR4 (N9739, N9726, N3405, N3168, N8956);
xor XOR2 (N9740, N9722, N504);
or OR4 (N9741, N9736, N4076, N7127, N6147);
nor NOR2 (N9742, N9739, N6057);
or OR3 (N9743, N9741, N2465, N2385);
nor NOR3 (N9744, N9725, N6497, N7678);
nand NAND3 (N9745, N9743, N8703, N8935);
or OR3 (N9746, N9745, N5524, N3662);
buf BUF1 (N9747, N9732);
or OR2 (N9748, N9744, N3316);
buf BUF1 (N9749, N9747);
or OR2 (N9750, N9737, N4443);
nand NAND4 (N9751, N9748, N8451, N8054, N9083);
nand NAND3 (N9752, N9746, N5234, N6982);
not NOT1 (N9753, N9733);
nand NAND2 (N9754, N9753, N2422);
nand NAND4 (N9755, N9738, N5512, N3217, N2596);
nor NOR3 (N9756, N9734, N5943, N1007);
or OR2 (N9757, N9755, N850);
nand NAND3 (N9758, N9749, N8337, N7992);
buf BUF1 (N9759, N9754);
buf BUF1 (N9760, N9742);
buf BUF1 (N9761, N9752);
or OR3 (N9762, N9760, N8892, N5698);
nor NOR4 (N9763, N9757, N5975, N1522, N5449);
xor XOR2 (N9764, N9740, N8786);
nand NAND3 (N9765, N9761, N1428, N1319);
xor XOR2 (N9766, N9762, N7321);
not NOT1 (N9767, N9763);
and AND3 (N9768, N9751, N4892, N6175);
not NOT1 (N9769, N9758);
nand NAND2 (N9770, N9765, N7313);
not NOT1 (N9771, N9764);
nor NOR2 (N9772, N9771, N1115);
buf BUF1 (N9773, N9768);
nor NOR4 (N9774, N9766, N7031, N589, N8384);
buf BUF1 (N9775, N9756);
nand NAND4 (N9776, N9774, N5063, N3832, N2774);
xor XOR2 (N9777, N9735, N1755);
nor NOR4 (N9778, N9767, N3860, N8321, N1746);
and AND3 (N9779, N9759, N7989, N2077);
not NOT1 (N9780, N9772);
buf BUF1 (N9781, N9773);
and AND3 (N9782, N9769, N7721, N689);
or OR2 (N9783, N9777, N2925);
or OR2 (N9784, N9779, N3795);
not NOT1 (N9785, N9778);
buf BUF1 (N9786, N9776);
buf BUF1 (N9787, N9750);
not NOT1 (N9788, N9770);
nand NAND4 (N9789, N9781, N5826, N4231, N6385);
nand NAND3 (N9790, N9787, N4770, N8443);
buf BUF1 (N9791, N9785);
xor XOR2 (N9792, N9791, N633);
not NOT1 (N9793, N9782);
not NOT1 (N9794, N9788);
nor NOR3 (N9795, N9775, N5131, N434);
nor NOR2 (N9796, N9790, N4741);
nand NAND3 (N9797, N9794, N1941, N6592);
or OR4 (N9798, N9784, N9049, N8996, N2808);
or OR3 (N9799, N9795, N9595, N9540);
not NOT1 (N9800, N9793);
nand NAND2 (N9801, N9796, N5434);
not NOT1 (N9802, N9798);
xor XOR2 (N9803, N9786, N1140);
nand NAND2 (N9804, N9802, N2543);
or OR4 (N9805, N9799, N7151, N8933, N9443);
and AND4 (N9806, N9797, N2404, N1212, N1509);
not NOT1 (N9807, N9805);
buf BUF1 (N9808, N9803);
not NOT1 (N9809, N9801);
nor NOR3 (N9810, N9806, N2276, N5425);
not NOT1 (N9811, N9792);
xor XOR2 (N9812, N9808, N5345);
nand NAND2 (N9813, N9783, N1770);
nand NAND2 (N9814, N9807, N6566);
or OR3 (N9815, N9812, N9371, N7125);
not NOT1 (N9816, N9814);
or OR4 (N9817, N9810, N5980, N5135, N5537);
not NOT1 (N9818, N9804);
buf BUF1 (N9819, N9816);
buf BUF1 (N9820, N9811);
buf BUF1 (N9821, N9780);
nor NOR2 (N9822, N9817, N3044);
buf BUF1 (N9823, N9809);
and AND2 (N9824, N9818, N1343);
or OR4 (N9825, N9820, N2736, N2962, N4298);
nand NAND3 (N9826, N9822, N2131, N6131);
xor XOR2 (N9827, N9824, N4820);
or OR3 (N9828, N9813, N6275, N2983);
not NOT1 (N9829, N9823);
or OR4 (N9830, N9815, N2811, N9517, N2808);
buf BUF1 (N9831, N9829);
buf BUF1 (N9832, N9819);
nor NOR2 (N9833, N9827, N3976);
nand NAND2 (N9834, N9826, N3154);
buf BUF1 (N9835, N9828);
not NOT1 (N9836, N9834);
xor XOR2 (N9837, N9833, N2219);
and AND4 (N9838, N9825, N8896, N3896, N9683);
and AND2 (N9839, N9821, N6380);
buf BUF1 (N9840, N9832);
nand NAND2 (N9841, N9840, N6634);
nand NAND3 (N9842, N9831, N3863, N2820);
or OR2 (N9843, N9830, N5685);
and AND4 (N9844, N9789, N6307, N850, N8067);
buf BUF1 (N9845, N9800);
nand NAND3 (N9846, N9835, N5952, N8693);
or OR3 (N9847, N9838, N9003, N8873);
buf BUF1 (N9848, N9841);
buf BUF1 (N9849, N9848);
not NOT1 (N9850, N9843);
or OR2 (N9851, N9849, N3232);
nand NAND3 (N9852, N9847, N9488, N3767);
or OR2 (N9853, N9839, N8724);
nand NAND4 (N9854, N9844, N9057, N575, N927);
or OR2 (N9855, N9837, N1484);
nand NAND4 (N9856, N9851, N7560, N8404, N5452);
buf BUF1 (N9857, N9852);
nand NAND3 (N9858, N9857, N8751, N7731);
nor NOR3 (N9859, N9836, N965, N1761);
and AND2 (N9860, N9855, N2455);
or OR2 (N9861, N9854, N2090);
xor XOR2 (N9862, N9860, N8302);
nand NAND4 (N9863, N9845, N6851, N9252, N2631);
not NOT1 (N9864, N9861);
buf BUF1 (N9865, N9856);
and AND3 (N9866, N9853, N9588, N870);
xor XOR2 (N9867, N9858, N3202);
not NOT1 (N9868, N9865);
and AND2 (N9869, N9859, N655);
nand NAND4 (N9870, N9842, N8210, N530, N3161);
nor NOR4 (N9871, N9862, N3783, N5273, N6420);
or OR4 (N9872, N9869, N534, N6977, N4397);
or OR2 (N9873, N9868, N8092);
and AND4 (N9874, N9873, N9686, N2203, N4345);
nand NAND4 (N9875, N9870, N1361, N7755, N2608);
or OR4 (N9876, N9874, N6015, N5402, N5947);
not NOT1 (N9877, N9867);
buf BUF1 (N9878, N9872);
not NOT1 (N9879, N9846);
nand NAND3 (N9880, N9850, N3068, N7071);
nor NOR4 (N9881, N9877, N6373, N7878, N8081);
xor XOR2 (N9882, N9881, N8207);
and AND3 (N9883, N9875, N5593, N5399);
not NOT1 (N9884, N9879);
xor XOR2 (N9885, N9876, N8187);
xor XOR2 (N9886, N9883, N7059);
nand NAND3 (N9887, N9886, N6397, N2127);
buf BUF1 (N9888, N9864);
or OR3 (N9889, N9885, N835, N4903);
xor XOR2 (N9890, N9878, N2565);
buf BUF1 (N9891, N9866);
and AND2 (N9892, N9889, N7618);
and AND4 (N9893, N9884, N3333, N9725, N3097);
not NOT1 (N9894, N9871);
nand NAND4 (N9895, N9894, N1431, N4983, N7642);
not NOT1 (N9896, N9888);
not NOT1 (N9897, N9882);
not NOT1 (N9898, N9893);
xor XOR2 (N9899, N9863, N3076);
xor XOR2 (N9900, N9887, N4629);
nand NAND4 (N9901, N9892, N1496, N886, N1235);
or OR3 (N9902, N9895, N6485, N4630);
nor NOR4 (N9903, N9891, N4168, N2990, N1674);
and AND4 (N9904, N9903, N5640, N8946, N1462);
nand NAND2 (N9905, N9880, N2135);
nand NAND2 (N9906, N9898, N4641);
buf BUF1 (N9907, N9900);
nand NAND3 (N9908, N9899, N4383, N9336);
nand NAND4 (N9909, N9897, N1978, N7634, N8661);
nand NAND4 (N9910, N9905, N5494, N3528, N5865);
not NOT1 (N9911, N9896);
nand NAND2 (N9912, N9909, N3371);
xor XOR2 (N9913, N9890, N7081);
not NOT1 (N9914, N9912);
buf BUF1 (N9915, N9906);
or OR4 (N9916, N9910, N2946, N3295, N5193);
or OR4 (N9917, N9904, N6523, N1753, N3043);
and AND4 (N9918, N9913, N9789, N3263, N2460);
buf BUF1 (N9919, N9908);
nand NAND3 (N9920, N9917, N674, N4926);
nand NAND3 (N9921, N9901, N8824, N5280);
or OR2 (N9922, N9911, N7183);
xor XOR2 (N9923, N9921, N2327);
nand NAND3 (N9924, N9922, N1712, N178);
or OR4 (N9925, N9923, N2781, N2849, N525);
not NOT1 (N9926, N9902);
and AND2 (N9927, N9924, N5638);
not NOT1 (N9928, N9919);
not NOT1 (N9929, N9925);
and AND2 (N9930, N9918, N5035);
buf BUF1 (N9931, N9926);
or OR3 (N9932, N9929, N8586, N5848);
buf BUF1 (N9933, N9930);
not NOT1 (N9934, N9927);
buf BUF1 (N9935, N9928);
nand NAND4 (N9936, N9907, N3909, N9706, N1810);
and AND4 (N9937, N9920, N3137, N2506, N3281);
buf BUF1 (N9938, N9932);
nand NAND2 (N9939, N9937, N5625);
nand NAND4 (N9940, N9916, N6034, N4697, N3429);
not NOT1 (N9941, N9931);
not NOT1 (N9942, N9933);
xor XOR2 (N9943, N9934, N2779);
not NOT1 (N9944, N9936);
buf BUF1 (N9945, N9914);
not NOT1 (N9946, N9945);
xor XOR2 (N9947, N9941, N4451);
or OR3 (N9948, N9915, N1806, N5121);
not NOT1 (N9949, N9939);
nor NOR4 (N9950, N9944, N9817, N7449, N1299);
xor XOR2 (N9951, N9942, N6108);
buf BUF1 (N9952, N9949);
nor NOR3 (N9953, N9948, N8330, N2242);
nand NAND3 (N9954, N9943, N9880, N8776);
nor NOR3 (N9955, N9950, N3814, N5388);
xor XOR2 (N9956, N9953, N6255);
and AND2 (N9957, N9935, N2450);
or OR3 (N9958, N9954, N2363, N3842);
nor NOR3 (N9959, N9947, N1623, N4090);
xor XOR2 (N9960, N9956, N5637);
and AND2 (N9961, N9940, N3763);
and AND2 (N9962, N9958, N7460);
or OR3 (N9963, N9952, N9577, N9711);
not NOT1 (N9964, N9960);
buf BUF1 (N9965, N9957);
nand NAND4 (N9966, N9955, N4284, N2317, N2601);
and AND2 (N9967, N9961, N2906);
buf BUF1 (N9968, N9951);
nand NAND2 (N9969, N9963, N8337);
nand NAND3 (N9970, N9966, N9749, N6351);
nand NAND3 (N9971, N9970, N2306, N6269);
nor NOR4 (N9972, N9969, N4649, N3672, N19);
xor XOR2 (N9973, N9971, N5782);
nor NOR3 (N9974, N9938, N856, N7777);
xor XOR2 (N9975, N9965, N2712);
not NOT1 (N9976, N9974);
or OR3 (N9977, N9964, N5380, N7977);
and AND2 (N9978, N9977, N9652);
buf BUF1 (N9979, N9976);
and AND4 (N9980, N9972, N8532, N4243, N523);
and AND4 (N9981, N9967, N7915, N2473, N9649);
xor XOR2 (N9982, N9980, N4070);
and AND4 (N9983, N9962, N5247, N1393, N8541);
xor XOR2 (N9984, N9975, N2935);
nor NOR3 (N9985, N9978, N1877, N9416);
and AND2 (N9986, N9983, N1364);
nor NOR3 (N9987, N9985, N1666, N2422);
and AND4 (N9988, N9979, N7904, N5234, N304);
nand NAND4 (N9989, N9987, N140, N7995, N7858);
nor NOR4 (N9990, N9959, N4248, N9488, N523);
nor NOR4 (N9991, N9990, N3091, N7987, N6333);
and AND2 (N9992, N9991, N6688);
nor NOR3 (N9993, N9986, N3553, N1442);
or OR4 (N9994, N9988, N5657, N2265, N5219);
nand NAND4 (N9995, N9946, N7529, N2, N6932);
nand NAND3 (N9996, N9995, N7308, N6670);
not NOT1 (N9997, N9982);
and AND3 (N9998, N9996, N1181, N3939);
xor XOR2 (N9999, N9973, N848);
nor NOR3 (N10000, N9992, N6889, N8164);
buf BUF1 (N10001, N10000);
nand NAND2 (N10002, N9997, N9475);
or OR4 (N10003, N9999, N2941, N2221, N6671);
or OR3 (N10004, N9981, N9703, N509);
not NOT1 (N10005, N10001);
not NOT1 (N10006, N10002);
xor XOR2 (N10007, N9989, N5000);
buf BUF1 (N10008, N9993);
or OR4 (N10009, N10004, N1886, N6114, N576);
nor NOR4 (N10010, N9984, N8372, N7794, N6604);
xor XOR2 (N10011, N10007, N2974);
nand NAND4 (N10012, N10011, N6030, N81, N3325);
nand NAND2 (N10013, N10009, N2040);
xor XOR2 (N10014, N9968, N1432);
nand NAND4 (N10015, N10003, N6596, N9170, N8940);
buf BUF1 (N10016, N10008);
xor XOR2 (N10017, N9998, N3300);
not NOT1 (N10018, N10006);
or OR2 (N10019, N10018, N1338);
nor NOR3 (N10020, N10013, N9358, N6328);
nor NOR4 (N10021, N9994, N1343, N4761, N577);
nand NAND2 (N10022, N10010, N765);
buf BUF1 (N10023, N10020);
nor NOR2 (N10024, N10005, N9404);
and AND3 (N10025, N10015, N725, N8737);
nor NOR2 (N10026, N10016, N1768);
and AND4 (N10027, N10023, N7713, N9156, N6082);
and AND2 (N10028, N10014, N7326);
and AND2 (N10029, N10027, N3057);
nor NOR3 (N10030, N10026, N2534, N9943);
nand NAND3 (N10031, N10029, N3942, N9803);
not NOT1 (N10032, N10031);
and AND2 (N10033, N10030, N7709);
nor NOR3 (N10034, N10012, N1399, N5231);
or OR3 (N10035, N10033, N9046, N2182);
and AND4 (N10036, N10034, N7938, N7056, N7144);
nand NAND3 (N10037, N10035, N4851, N5738);
xor XOR2 (N10038, N10017, N8451);
nand NAND2 (N10039, N10019, N7932);
nor NOR2 (N10040, N10036, N6802);
and AND4 (N10041, N10028, N3985, N7628, N8231);
not NOT1 (N10042, N10040);
nand NAND2 (N10043, N10021, N4336);
nand NAND3 (N10044, N10043, N4376, N4210);
or OR2 (N10045, N10038, N4352);
or OR4 (N10046, N10022, N1332, N7694, N5231);
and AND2 (N10047, N10041, N4873);
and AND3 (N10048, N10032, N4639, N7436);
xor XOR2 (N10049, N10046, N6472);
nand NAND4 (N10050, N10042, N7637, N2733, N6762);
nor NOR4 (N10051, N10024, N2646, N1494, N8774);
nand NAND3 (N10052, N10050, N4186, N8162);
buf BUF1 (N10053, N10051);
and AND4 (N10054, N10039, N2811, N2875, N211);
or OR3 (N10055, N10048, N9957, N4953);
and AND4 (N10056, N10025, N8582, N4927, N4568);
buf BUF1 (N10057, N10054);
xor XOR2 (N10058, N10045, N1474);
xor XOR2 (N10059, N10057, N362);
not NOT1 (N10060, N10059);
not NOT1 (N10061, N10044);
xor XOR2 (N10062, N10049, N7718);
or OR3 (N10063, N10058, N7687, N1077);
nand NAND2 (N10064, N10052, N801);
or OR2 (N10065, N10053, N9832);
nand NAND4 (N10066, N10037, N8587, N4302, N9015);
nor NOR4 (N10067, N10060, N6766, N1096, N7389);
or OR2 (N10068, N10066, N357);
not NOT1 (N10069, N10056);
and AND2 (N10070, N10064, N4218);
not NOT1 (N10071, N10070);
xor XOR2 (N10072, N10068, N9753);
or OR4 (N10073, N10062, N147, N5258, N7359);
buf BUF1 (N10074, N10071);
buf BUF1 (N10075, N10065);
nor NOR3 (N10076, N10069, N5848, N1207);
xor XOR2 (N10077, N10075, N2398);
or OR4 (N10078, N10074, N2344, N7672, N5665);
not NOT1 (N10079, N10047);
nand NAND4 (N10080, N10067, N6998, N7329, N7262);
nand NAND3 (N10081, N10063, N9569, N7054);
buf BUF1 (N10082, N10072);
buf BUF1 (N10083, N10079);
and AND2 (N10084, N10083, N8660);
nand NAND3 (N10085, N10082, N1002, N9810);
nor NOR2 (N10086, N10077, N9733);
and AND3 (N10087, N10055, N9266, N8022);
nor NOR4 (N10088, N10076, N4941, N8174, N5005);
not NOT1 (N10089, N10073);
nor NOR2 (N10090, N10061, N5053);
xor XOR2 (N10091, N10084, N2861);
and AND2 (N10092, N10088, N1648);
or OR3 (N10093, N10081, N2682, N9870);
buf BUF1 (N10094, N10093);
buf BUF1 (N10095, N10078);
nand NAND4 (N10096, N10086, N3485, N6007, N5178);
nand NAND4 (N10097, N10095, N9650, N3069, N4441);
nor NOR2 (N10098, N10091, N698);
nand NAND4 (N10099, N10085, N1209, N1669, N141);
not NOT1 (N10100, N10089);
not NOT1 (N10101, N10098);
not NOT1 (N10102, N10094);
not NOT1 (N10103, N10100);
not NOT1 (N10104, N10103);
nor NOR3 (N10105, N10080, N9664, N26);
nand NAND3 (N10106, N10102, N5530, N1627);
or OR2 (N10107, N10097, N918);
nor NOR2 (N10108, N10096, N5629);
buf BUF1 (N10109, N10101);
not NOT1 (N10110, N10099);
or OR2 (N10111, N10106, N8933);
nor NOR3 (N10112, N10087, N5225, N4069);
buf BUF1 (N10113, N10108);
or OR3 (N10114, N10090, N19, N4540);
or OR4 (N10115, N10114, N8668, N6550, N432);
or OR4 (N10116, N10113, N5033, N4599, N8408);
or OR4 (N10117, N10092, N9060, N4774, N913);
nand NAND3 (N10118, N10115, N6793, N7205);
nand NAND3 (N10119, N10107, N450, N8698);
not NOT1 (N10120, N10119);
and AND2 (N10121, N10116, N4205);
not NOT1 (N10122, N10120);
not NOT1 (N10123, N10118);
nor NOR4 (N10124, N10105, N4888, N6696, N2948);
or OR3 (N10125, N10111, N3198, N5151);
nand NAND4 (N10126, N10104, N4106, N4882, N3152);
nand NAND3 (N10127, N10124, N523, N5034);
and AND3 (N10128, N10127, N4532, N6633);
buf BUF1 (N10129, N10122);
nand NAND2 (N10130, N10129, N3329);
not NOT1 (N10131, N10126);
nor NOR4 (N10132, N10109, N6899, N8502, N4342);
or OR2 (N10133, N10112, N3423);
not NOT1 (N10134, N10123);
or OR2 (N10135, N10130, N6532);
not NOT1 (N10136, N10134);
xor XOR2 (N10137, N10133, N2884);
and AND3 (N10138, N10125, N10119, N4698);
or OR3 (N10139, N10137, N347, N9501);
nor NOR3 (N10140, N10117, N1721, N8702);
or OR4 (N10141, N10121, N2245, N2776, N1912);
or OR4 (N10142, N10135, N4123, N5592, N6690);
not NOT1 (N10143, N10110);
or OR4 (N10144, N10131, N4168, N5538, N9142);
and AND2 (N10145, N10142, N676);
and AND4 (N10146, N10128, N3434, N6632, N904);
and AND4 (N10147, N10139, N5645, N4593, N8603);
nor NOR4 (N10148, N10145, N3179, N5689, N4049);
xor XOR2 (N10149, N10147, N5691);
not NOT1 (N10150, N10141);
and AND2 (N10151, N10143, N2637);
nand NAND3 (N10152, N10148, N4070, N2438);
buf BUF1 (N10153, N10140);
or OR2 (N10154, N10144, N8146);
and AND2 (N10155, N10150, N2461);
xor XOR2 (N10156, N10138, N2283);
or OR2 (N10157, N10153, N1005);
nand NAND3 (N10158, N10132, N7963, N4119);
nor NOR3 (N10159, N10156, N4376, N7561);
xor XOR2 (N10160, N10158, N752);
or OR2 (N10161, N10136, N8971);
nand NAND2 (N10162, N10159, N9283);
nand NAND2 (N10163, N10151, N1313);
nand NAND4 (N10164, N10163, N3947, N10077, N6725);
nand NAND2 (N10165, N10164, N8713);
nand NAND2 (N10166, N10146, N3162);
nand NAND3 (N10167, N10155, N709, N5770);
xor XOR2 (N10168, N10160, N2894);
xor XOR2 (N10169, N10165, N6434);
xor XOR2 (N10170, N10162, N7639);
xor XOR2 (N10171, N10149, N8350);
not NOT1 (N10172, N10152);
xor XOR2 (N10173, N10161, N5237);
buf BUF1 (N10174, N10154);
xor XOR2 (N10175, N10168, N10118);
and AND4 (N10176, N10167, N1890, N6827, N3120);
or OR4 (N10177, N10171, N9707, N7555, N5948);
not NOT1 (N10178, N10173);
nand NAND3 (N10179, N10178, N7748, N8926);
and AND4 (N10180, N10179, N548, N497, N10093);
nand NAND2 (N10181, N10175, N3907);
or OR3 (N10182, N10177, N4788, N1136);
and AND3 (N10183, N10181, N4350, N7147);
buf BUF1 (N10184, N10182);
and AND4 (N10185, N10166, N9581, N4879, N6106);
and AND2 (N10186, N10157, N941);
buf BUF1 (N10187, N10184);
buf BUF1 (N10188, N10186);
xor XOR2 (N10189, N10174, N2670);
nand NAND2 (N10190, N10187, N4185);
not NOT1 (N10191, N10189);
nor NOR2 (N10192, N10170, N8703);
nand NAND4 (N10193, N10183, N10159, N8991, N7317);
or OR4 (N10194, N10191, N9488, N8711, N995);
and AND4 (N10195, N10192, N2705, N6277, N268);
not NOT1 (N10196, N10190);
or OR3 (N10197, N10169, N2169, N7736);
and AND4 (N10198, N10194, N4060, N8353, N9317);
xor XOR2 (N10199, N10197, N4724);
nand NAND2 (N10200, N10198, N6020);
and AND2 (N10201, N10180, N5150);
buf BUF1 (N10202, N10201);
or OR3 (N10203, N10195, N1026, N9516);
not NOT1 (N10204, N10176);
and AND2 (N10205, N10199, N9714);
xor XOR2 (N10206, N10203, N7724);
buf BUF1 (N10207, N10188);
or OR2 (N10208, N10196, N3810);
nor NOR2 (N10209, N10200, N6991);
not NOT1 (N10210, N10193);
xor XOR2 (N10211, N10209, N2595);
buf BUF1 (N10212, N10210);
and AND2 (N10213, N10211, N8571);
not NOT1 (N10214, N10172);
nor NOR3 (N10215, N10202, N8359, N4440);
buf BUF1 (N10216, N10206);
not NOT1 (N10217, N10205);
xor XOR2 (N10218, N10217, N5529);
xor XOR2 (N10219, N10208, N54);
buf BUF1 (N10220, N10213);
buf BUF1 (N10221, N10216);
and AND2 (N10222, N10219, N8158);
or OR4 (N10223, N10207, N397, N4413, N4600);
xor XOR2 (N10224, N10212, N4174);
buf BUF1 (N10225, N10222);
buf BUF1 (N10226, N10218);
nand NAND4 (N10227, N10220, N3565, N7805, N1143);
xor XOR2 (N10228, N10224, N4003);
or OR3 (N10229, N10223, N297, N806);
not NOT1 (N10230, N10214);
buf BUF1 (N10231, N10227);
xor XOR2 (N10232, N10228, N5992);
nand NAND4 (N10233, N10232, N4901, N155, N9551);
or OR4 (N10234, N10233, N2628, N3574, N802);
or OR3 (N10235, N10230, N5007, N1316);
or OR3 (N10236, N10215, N6284, N6899);
nand NAND3 (N10237, N10235, N10065, N8595);
buf BUF1 (N10238, N10231);
not NOT1 (N10239, N10237);
xor XOR2 (N10240, N10229, N250);
and AND3 (N10241, N10226, N2473, N7960);
or OR2 (N10242, N10241, N7885);
nand NAND2 (N10243, N10204, N7426);
nand NAND4 (N10244, N10239, N2422, N6344, N1750);
nor NOR2 (N10245, N10221, N3673);
nand NAND3 (N10246, N10245, N6172, N6735);
or OR2 (N10247, N10234, N10094);
and AND3 (N10248, N10242, N8050, N366);
not NOT1 (N10249, N10238);
nand NAND2 (N10250, N10244, N1700);
or OR4 (N10251, N10250, N5887, N3240, N6302);
nand NAND3 (N10252, N10225, N1853, N4225);
buf BUF1 (N10253, N10236);
and AND4 (N10254, N10247, N8121, N5784, N254);
or OR3 (N10255, N10246, N3811, N7660);
or OR3 (N10256, N10248, N1214, N3064);
xor XOR2 (N10257, N10256, N569);
or OR2 (N10258, N10249, N6233);
nor NOR2 (N10259, N10251, N4668);
nand NAND4 (N10260, N10253, N7386, N9411, N8323);
nor NOR2 (N10261, N10258, N5336);
or OR4 (N10262, N10240, N7649, N117, N9578);
xor XOR2 (N10263, N10257, N6297);
not NOT1 (N10264, N10243);
buf BUF1 (N10265, N10254);
nand NAND4 (N10266, N10264, N4033, N3431, N8100);
nor NOR4 (N10267, N10263, N3861, N2889, N3758);
xor XOR2 (N10268, N10252, N3280);
and AND2 (N10269, N10268, N2499);
nor NOR2 (N10270, N10260, N7512);
xor XOR2 (N10271, N10185, N4319);
and AND4 (N10272, N10266, N4269, N2697, N6730);
and AND2 (N10273, N10261, N2755);
buf BUF1 (N10274, N10273);
not NOT1 (N10275, N10269);
or OR3 (N10276, N10262, N3302, N6753);
nor NOR2 (N10277, N10259, N7362);
nor NOR4 (N10278, N10265, N10223, N7641, N2391);
nand NAND4 (N10279, N10277, N6267, N1852, N5782);
nand NAND3 (N10280, N10278, N3882, N2169);
nor NOR2 (N10281, N10280, N6019);
nand NAND2 (N10282, N10271, N3056);
nand NAND2 (N10283, N10255, N2860);
and AND4 (N10284, N10281, N9549, N8834, N10279);
nand NAND2 (N10285, N7561, N2007);
or OR4 (N10286, N10267, N6053, N9899, N808);
not NOT1 (N10287, N10284);
buf BUF1 (N10288, N10287);
and AND4 (N10289, N10286, N415, N4255, N381);
not NOT1 (N10290, N10282);
nand NAND4 (N10291, N10290, N5798, N5759, N136);
or OR3 (N10292, N10291, N5566, N8957);
nand NAND2 (N10293, N10289, N3439);
and AND3 (N10294, N10274, N6127, N4423);
and AND2 (N10295, N10293, N4772);
nor NOR2 (N10296, N10276, N6348);
nand NAND3 (N10297, N10272, N2126, N6309);
xor XOR2 (N10298, N10297, N9715);
nand NAND3 (N10299, N10283, N3343, N7328);
buf BUF1 (N10300, N10270);
buf BUF1 (N10301, N10288);
not NOT1 (N10302, N10299);
xor XOR2 (N10303, N10298, N9686);
xor XOR2 (N10304, N10301, N9403);
nor NOR4 (N10305, N10295, N3136, N4707, N8875);
xor XOR2 (N10306, N10285, N2357);
not NOT1 (N10307, N10305);
and AND2 (N10308, N10302, N8801);
nor NOR2 (N10309, N10296, N731);
and AND3 (N10310, N10300, N1308, N527);
nor NOR3 (N10311, N10309, N7109, N9879);
xor XOR2 (N10312, N10306, N3397);
or OR2 (N10313, N10304, N7759);
not NOT1 (N10314, N10312);
xor XOR2 (N10315, N10292, N5050);
not NOT1 (N10316, N10311);
xor XOR2 (N10317, N10307, N1762);
nor NOR2 (N10318, N10294, N3043);
xor XOR2 (N10319, N10303, N470);
nor NOR4 (N10320, N10317, N8948, N9481, N5939);
and AND4 (N10321, N10315, N6795, N5809, N6062);
xor XOR2 (N10322, N10321, N2558);
buf BUF1 (N10323, N10308);
nand NAND2 (N10324, N10323, N5840);
not NOT1 (N10325, N10316);
or OR4 (N10326, N10318, N9917, N10081, N521);
nor NOR3 (N10327, N10324, N4833, N5062);
and AND2 (N10328, N10326, N3607);
and AND4 (N10329, N10275, N8229, N9886, N3894);
or OR4 (N10330, N10329, N3142, N987, N6770);
or OR2 (N10331, N10314, N5372);
xor XOR2 (N10332, N10328, N4232);
or OR3 (N10333, N10310, N6478, N8236);
nand NAND4 (N10334, N10333, N7049, N6348, N6663);
or OR3 (N10335, N10320, N3048, N10327);
xor XOR2 (N10336, N4361, N4665);
and AND4 (N10337, N10319, N5131, N6527, N4540);
and AND4 (N10338, N10330, N5524, N6515, N4137);
nand NAND4 (N10339, N10338, N6421, N5668, N9330);
not NOT1 (N10340, N10337);
not NOT1 (N10341, N10340);
nor NOR3 (N10342, N10331, N3993, N5203);
and AND2 (N10343, N10339, N3895);
xor XOR2 (N10344, N10342, N7204);
nand NAND4 (N10345, N10336, N3677, N3284, N3627);
and AND2 (N10346, N10345, N4217);
or OR2 (N10347, N10344, N1226);
or OR2 (N10348, N10343, N9131);
buf BUF1 (N10349, N10348);
and AND2 (N10350, N10332, N8352);
not NOT1 (N10351, N10346);
xor XOR2 (N10352, N10350, N917);
xor XOR2 (N10353, N10322, N3522);
not NOT1 (N10354, N10351);
nor NOR4 (N10355, N10341, N1460, N681, N593);
not NOT1 (N10356, N10355);
buf BUF1 (N10357, N10325);
nand NAND2 (N10358, N10334, N9131);
nor NOR2 (N10359, N10335, N2693);
and AND4 (N10360, N10354, N1080, N7865, N7255);
and AND4 (N10361, N10349, N5329, N2906, N10221);
nor NOR3 (N10362, N10361, N6002, N10078);
nor NOR4 (N10363, N10357, N9120, N3754, N9823);
buf BUF1 (N10364, N10356);
nand NAND2 (N10365, N10347, N8081);
not NOT1 (N10366, N10352);
or OR4 (N10367, N10313, N730, N10066, N409);
buf BUF1 (N10368, N10353);
or OR3 (N10369, N10365, N6003, N8011);
or OR3 (N10370, N10359, N1216, N5140);
nand NAND4 (N10371, N10367, N2091, N3623, N1056);
and AND2 (N10372, N10358, N6913);
not NOT1 (N10373, N10369);
buf BUF1 (N10374, N10373);
nand NAND3 (N10375, N10364, N5847, N7554);
buf BUF1 (N10376, N10360);
nand NAND3 (N10377, N10376, N1177, N9012);
nand NAND2 (N10378, N10370, N9351);
not NOT1 (N10379, N10374);
or OR3 (N10380, N10372, N2332, N8678);
nor NOR4 (N10381, N10362, N7786, N5353, N4992);
not NOT1 (N10382, N10379);
nand NAND2 (N10383, N10371, N7087);
and AND3 (N10384, N10363, N6576, N2153);
or OR2 (N10385, N10383, N3952);
or OR3 (N10386, N10366, N3827, N2937);
not NOT1 (N10387, N10381);
xor XOR2 (N10388, N10385, N5263);
and AND4 (N10389, N10384, N6073, N8065, N2724);
not NOT1 (N10390, N10378);
xor XOR2 (N10391, N10382, N9088);
and AND3 (N10392, N10377, N7816, N714);
xor XOR2 (N10393, N10387, N1514);
and AND2 (N10394, N10388, N10384);
not NOT1 (N10395, N10393);
buf BUF1 (N10396, N10391);
not NOT1 (N10397, N10395);
not NOT1 (N10398, N10390);
and AND2 (N10399, N10396, N260);
or OR4 (N10400, N10375, N2553, N10224, N2273);
buf BUF1 (N10401, N10397);
nor NOR2 (N10402, N10400, N25);
buf BUF1 (N10403, N10401);
or OR4 (N10404, N10402, N293, N7303, N9853);
not NOT1 (N10405, N10386);
and AND2 (N10406, N10389, N5699);
nand NAND3 (N10407, N10403, N3585, N3207);
and AND2 (N10408, N10380, N8281);
nand NAND3 (N10409, N10398, N7978, N7251);
nor NOR4 (N10410, N10408, N7523, N8153, N4800);
and AND3 (N10411, N10406, N3658, N6695);
not NOT1 (N10412, N10404);
not NOT1 (N10413, N10407);
xor XOR2 (N10414, N10410, N6936);
buf BUF1 (N10415, N10411);
and AND4 (N10416, N10405, N4426, N4214, N8827);
xor XOR2 (N10417, N10412, N9547);
nand NAND2 (N10418, N10392, N3884);
xor XOR2 (N10419, N10417, N605);
and AND3 (N10420, N10418, N4735, N5296);
nor NOR2 (N10421, N10399, N8341);
buf BUF1 (N10422, N10368);
nor NOR3 (N10423, N10415, N4985, N4590);
nand NAND4 (N10424, N10409, N4637, N9680, N6419);
nor NOR4 (N10425, N10424, N9141, N10224, N1537);
or OR2 (N10426, N10414, N9925);
or OR3 (N10427, N10422, N6139, N106);
not NOT1 (N10428, N10394);
nand NAND3 (N10429, N10421, N7960, N3401);
nand NAND3 (N10430, N10416, N7021, N448);
not NOT1 (N10431, N10428);
or OR3 (N10432, N10426, N1942, N2563);
and AND2 (N10433, N10420, N8093);
buf BUF1 (N10434, N10431);
not NOT1 (N10435, N10427);
nand NAND2 (N10436, N10419, N7932);
nor NOR2 (N10437, N10436, N1177);
not NOT1 (N10438, N10432);
nor NOR3 (N10439, N10430, N1120, N3754);
buf BUF1 (N10440, N10413);
and AND3 (N10441, N10438, N5659, N983);
not NOT1 (N10442, N10423);
nand NAND2 (N10443, N10435, N4708);
nor NOR3 (N10444, N10440, N8925, N4164);
xor XOR2 (N10445, N10444, N2163);
nor NOR2 (N10446, N10425, N1189);
nor NOR2 (N10447, N10446, N2272);
or OR2 (N10448, N10437, N6127);
and AND4 (N10449, N10442, N10057, N259, N785);
and AND3 (N10450, N10447, N9052, N9257);
xor XOR2 (N10451, N10429, N4061);
or OR4 (N10452, N10441, N10081, N7311, N9162);
or OR3 (N10453, N10452, N4310, N9009);
or OR2 (N10454, N10449, N7643);
buf BUF1 (N10455, N10453);
buf BUF1 (N10456, N10439);
xor XOR2 (N10457, N10455, N1426);
not NOT1 (N10458, N10434);
nand NAND3 (N10459, N10457, N4892, N6226);
xor XOR2 (N10460, N10450, N9490);
and AND3 (N10461, N10433, N4663, N2995);
not NOT1 (N10462, N10448);
nand NAND2 (N10463, N10461, N3564);
nor NOR2 (N10464, N10460, N3988);
not NOT1 (N10465, N10463);
xor XOR2 (N10466, N10445, N8113);
nor NOR4 (N10467, N10459, N1245, N5572, N7748);
or OR2 (N10468, N10464, N10260);
nand NAND2 (N10469, N10467, N9371);
buf BUF1 (N10470, N10451);
or OR2 (N10471, N10456, N8495);
nand NAND3 (N10472, N10468, N2982, N6782);
and AND3 (N10473, N10458, N10283, N9156);
nand NAND4 (N10474, N10454, N3775, N4083, N822);
or OR3 (N10475, N10462, N2850, N8600);
buf BUF1 (N10476, N10469);
and AND4 (N10477, N10476, N5538, N1977, N1869);
xor XOR2 (N10478, N10443, N6951);
nand NAND4 (N10479, N10475, N425, N4523, N5016);
and AND2 (N10480, N10473, N9533);
nor NOR4 (N10481, N10480, N1688, N3234, N3608);
buf BUF1 (N10482, N10471);
nand NAND4 (N10483, N10470, N9619, N6622, N646);
xor XOR2 (N10484, N10477, N9065);
buf BUF1 (N10485, N10484);
xor XOR2 (N10486, N10478, N6444);
xor XOR2 (N10487, N10486, N5547);
buf BUF1 (N10488, N10479);
or OR2 (N10489, N10488, N1327);
or OR4 (N10490, N10485, N1084, N9559, N5009);
not NOT1 (N10491, N10466);
xor XOR2 (N10492, N10489, N10197);
or OR4 (N10493, N10492, N237, N8114, N4461);
buf BUF1 (N10494, N10465);
or OR2 (N10495, N10481, N4656);
xor XOR2 (N10496, N10494, N2158);
not NOT1 (N10497, N10474);
or OR3 (N10498, N10497, N4351, N5521);
buf BUF1 (N10499, N10482);
nand NAND4 (N10500, N10495, N3492, N1664, N131);
not NOT1 (N10501, N10496);
xor XOR2 (N10502, N10500, N5972);
nor NOR3 (N10503, N10491, N7364, N6022);
xor XOR2 (N10504, N10483, N1682);
nor NOR3 (N10505, N10504, N10096, N6996);
and AND3 (N10506, N10503, N4398, N7835);
and AND3 (N10507, N10490, N3052, N8100);
nand NAND3 (N10508, N10501, N10194, N1777);
nand NAND2 (N10509, N10499, N5974);
and AND4 (N10510, N10506, N3096, N6032, N5444);
nand NAND3 (N10511, N10510, N6643, N8626);
nor NOR3 (N10512, N10511, N7352, N2196);
or OR4 (N10513, N10509, N9455, N5095, N7894);
xor XOR2 (N10514, N10487, N7076);
and AND4 (N10515, N10502, N7143, N1739, N1960);
buf BUF1 (N10516, N10514);
xor XOR2 (N10517, N10498, N1342);
or OR3 (N10518, N10515, N8891, N5171);
nor NOR2 (N10519, N10508, N2264);
nor NOR2 (N10520, N10507, N645);
or OR3 (N10521, N10519, N1128, N4910);
or OR2 (N10522, N10521, N3756);
and AND2 (N10523, N10493, N1188);
nor NOR4 (N10524, N10513, N8677, N6663, N1897);
nand NAND4 (N10525, N10522, N6870, N2689, N1999);
xor XOR2 (N10526, N10472, N1807);
and AND4 (N10527, N10523, N2661, N5194, N9220);
buf BUF1 (N10528, N10526);
and AND4 (N10529, N10524, N3688, N1696, N4751);
nand NAND2 (N10530, N10505, N9033);
not NOT1 (N10531, N10512);
xor XOR2 (N10532, N10518, N5649);
xor XOR2 (N10533, N10527, N738);
nand NAND2 (N10534, N10529, N3412);
not NOT1 (N10535, N10533);
or OR3 (N10536, N10534, N2247, N2245);
buf BUF1 (N10537, N10530);
nor NOR4 (N10538, N10517, N7556, N5549, N8847);
buf BUF1 (N10539, N10535);
buf BUF1 (N10540, N10520);
and AND4 (N10541, N10537, N9626, N2770, N7073);
nand NAND4 (N10542, N10538, N1535, N7745, N2140);
or OR3 (N10543, N10528, N4318, N8388);
or OR2 (N10544, N10542, N1905);
nand NAND4 (N10545, N10539, N6252, N238, N1927);
buf BUF1 (N10546, N10532);
buf BUF1 (N10547, N10541);
nor NOR3 (N10548, N10516, N10387, N4122);
buf BUF1 (N10549, N10525);
nor NOR2 (N10550, N10531, N8133);
not NOT1 (N10551, N10544);
xor XOR2 (N10552, N10549, N7141);
nand NAND4 (N10553, N10548, N4239, N2010, N3879);
nor NOR4 (N10554, N10550, N5685, N1377, N2689);
nand NAND4 (N10555, N10540, N5662, N1759, N3216);
not NOT1 (N10556, N10555);
buf BUF1 (N10557, N10553);
and AND4 (N10558, N10546, N4783, N1124, N9271);
buf BUF1 (N10559, N10557);
not NOT1 (N10560, N10556);
and AND3 (N10561, N10552, N3228, N1001);
xor XOR2 (N10562, N10558, N345);
nand NAND3 (N10563, N10554, N171, N1358);
or OR4 (N10564, N10551, N2283, N6077, N5686);
buf BUF1 (N10565, N10564);
buf BUF1 (N10566, N10561);
xor XOR2 (N10567, N10566, N10205);
not NOT1 (N10568, N10563);
nand NAND3 (N10569, N10568, N1181, N6618);
and AND2 (N10570, N10567, N1988);
nand NAND3 (N10571, N10562, N1515, N2761);
and AND4 (N10572, N10545, N4379, N5712, N7624);
or OR2 (N10573, N10571, N308);
nand NAND2 (N10574, N10572, N793);
nand NAND4 (N10575, N10559, N8593, N4369, N1073);
buf BUF1 (N10576, N10569);
buf BUF1 (N10577, N10570);
xor XOR2 (N10578, N10543, N3024);
not NOT1 (N10579, N10576);
nand NAND2 (N10580, N10565, N2459);
buf BUF1 (N10581, N10574);
and AND2 (N10582, N10579, N9394);
nor NOR3 (N10583, N10575, N2948, N9802);
not NOT1 (N10584, N10547);
or OR2 (N10585, N10578, N7143);
and AND3 (N10586, N10536, N5759, N8609);
not NOT1 (N10587, N10560);
xor XOR2 (N10588, N10587, N7907);
nor NOR2 (N10589, N10573, N7939);
not NOT1 (N10590, N10588);
xor XOR2 (N10591, N10577, N1607);
not NOT1 (N10592, N10586);
not NOT1 (N10593, N10583);
and AND4 (N10594, N10584, N6740, N10136, N8080);
buf BUF1 (N10595, N10589);
or OR3 (N10596, N10594, N7846, N4366);
buf BUF1 (N10597, N10581);
buf BUF1 (N10598, N10582);
not NOT1 (N10599, N10598);
or OR2 (N10600, N10593, N8230);
or OR4 (N10601, N10599, N6746, N5879, N41);
nor NOR3 (N10602, N10601, N4425, N3436);
and AND2 (N10603, N10592, N8213);
and AND3 (N10604, N10602, N7661, N6372);
or OR2 (N10605, N10591, N9033);
xor XOR2 (N10606, N10596, N1510);
or OR3 (N10607, N10604, N2618, N4908);
nor NOR3 (N10608, N10597, N1042, N9216);
or OR2 (N10609, N10606, N2951);
nand NAND3 (N10610, N10607, N7176, N5221);
not NOT1 (N10611, N10585);
nor NOR2 (N10612, N10595, N10029);
xor XOR2 (N10613, N10580, N4276);
or OR4 (N10614, N10603, N6931, N7158, N6634);
buf BUF1 (N10615, N10605);
not NOT1 (N10616, N10613);
buf BUF1 (N10617, N10611);
nand NAND3 (N10618, N10612, N4208, N1727);
buf BUF1 (N10619, N10610);
and AND4 (N10620, N10616, N10498, N3980, N1435);
or OR3 (N10621, N10600, N3716, N4314);
or OR2 (N10622, N10615, N10291);
or OR3 (N10623, N10620, N9594, N7281);
and AND2 (N10624, N10618, N6772);
and AND4 (N10625, N10622, N945, N8229, N8470);
buf BUF1 (N10626, N10624);
and AND2 (N10627, N10625, N8586);
nor NOR3 (N10628, N10619, N8860, N7919);
xor XOR2 (N10629, N10608, N6275);
nand NAND2 (N10630, N10627, N10537);
xor XOR2 (N10631, N10614, N6521);
and AND2 (N10632, N10629, N1545);
nor NOR4 (N10633, N10631, N4893, N5441, N2705);
nor NOR2 (N10634, N10633, N2162);
or OR3 (N10635, N10590, N5328, N1850);
and AND3 (N10636, N10634, N5904, N6593);
and AND4 (N10637, N10632, N654, N6682, N7952);
not NOT1 (N10638, N10628);
xor XOR2 (N10639, N10636, N1359);
not NOT1 (N10640, N10635);
or OR3 (N10641, N10639, N9656, N8001);
or OR2 (N10642, N10630, N966);
nor NOR4 (N10643, N10640, N4787, N2977, N7680);
nand NAND3 (N10644, N10621, N4929, N8661);
or OR4 (N10645, N10642, N2048, N2513, N1735);
nor NOR3 (N10646, N10623, N4557, N4978);
nor NOR3 (N10647, N10637, N2867, N6512);
or OR4 (N10648, N10641, N1666, N6945, N9735);
or OR2 (N10649, N10648, N9755);
nand NAND4 (N10650, N10626, N9823, N5152, N955);
nor NOR2 (N10651, N10644, N7993);
not NOT1 (N10652, N10649);
nand NAND2 (N10653, N10645, N3405);
nor NOR3 (N10654, N10646, N1764, N7091);
nor NOR3 (N10655, N10643, N1199, N8838);
and AND2 (N10656, N10652, N9000);
or OR2 (N10657, N10651, N1084);
xor XOR2 (N10658, N10609, N10167);
or OR3 (N10659, N10653, N8041, N9941);
xor XOR2 (N10660, N10647, N10185);
and AND4 (N10661, N10656, N8942, N6693, N355);
or OR3 (N10662, N10658, N4329, N6101);
or OR2 (N10663, N10654, N7808);
nor NOR4 (N10664, N10660, N7273, N8379, N4703);
nand NAND4 (N10665, N10655, N8776, N2921, N6681);
nor NOR4 (N10666, N10663, N10249, N6266, N1565);
nor NOR3 (N10667, N10665, N6764, N2553);
not NOT1 (N10668, N10657);
xor XOR2 (N10669, N10662, N9928);
and AND3 (N10670, N10669, N3261, N2395);
buf BUF1 (N10671, N10668);
and AND3 (N10672, N10670, N6374, N87);
buf BUF1 (N10673, N10666);
or OR2 (N10674, N10659, N2194);
buf BUF1 (N10675, N10671);
nor NOR2 (N10676, N10675, N5321);
nor NOR3 (N10677, N10617, N1094, N3124);
not NOT1 (N10678, N10674);
nor NOR4 (N10679, N10676, N8808, N9978, N4693);
not NOT1 (N10680, N10673);
buf BUF1 (N10681, N10678);
xor XOR2 (N10682, N10679, N5454);
and AND2 (N10683, N10664, N4017);
nor NOR2 (N10684, N10683, N8656);
or OR4 (N10685, N10650, N4769, N156, N1547);
xor XOR2 (N10686, N10677, N3804);
buf BUF1 (N10687, N10685);
xor XOR2 (N10688, N10687, N1051);
or OR2 (N10689, N10672, N1768);
buf BUF1 (N10690, N10681);
or OR2 (N10691, N10690, N265);
nand NAND3 (N10692, N10686, N2535, N7030);
and AND4 (N10693, N10661, N7312, N6726, N821);
buf BUF1 (N10694, N10693);
xor XOR2 (N10695, N10682, N2584);
nand NAND2 (N10696, N10688, N9972);
nor NOR3 (N10697, N10680, N7344, N7822);
buf BUF1 (N10698, N10697);
buf BUF1 (N10699, N10696);
buf BUF1 (N10700, N10698);
nor NOR2 (N10701, N10699, N3115);
not NOT1 (N10702, N10694);
nor NOR2 (N10703, N10692, N7574);
and AND4 (N10704, N10702, N68, N3845, N4742);
nand NAND3 (N10705, N10703, N3150, N5059);
and AND3 (N10706, N10684, N10351, N5862);
nand NAND3 (N10707, N10701, N6266, N8777);
xor XOR2 (N10708, N10667, N507);
and AND4 (N10709, N10704, N1987, N4095, N5598);
or OR4 (N10710, N10706, N6464, N5274, N8386);
and AND3 (N10711, N10689, N7677, N6072);
nor NOR2 (N10712, N10710, N8316);
or OR3 (N10713, N10695, N5559, N9815);
not NOT1 (N10714, N10691);
buf BUF1 (N10715, N10705);
not NOT1 (N10716, N10707);
or OR4 (N10717, N10700, N5878, N7100, N4214);
nor NOR3 (N10718, N10709, N2817, N2208);
nand NAND3 (N10719, N10715, N97, N1903);
nand NAND3 (N10720, N10719, N2983, N10554);
and AND3 (N10721, N10716, N5698, N4354);
and AND2 (N10722, N10712, N8335);
buf BUF1 (N10723, N10708);
not NOT1 (N10724, N10714);
buf BUF1 (N10725, N10711);
and AND3 (N10726, N10713, N10614, N9233);
buf BUF1 (N10727, N10722);
buf BUF1 (N10728, N10727);
or OR2 (N10729, N10717, N4933);
not NOT1 (N10730, N10729);
xor XOR2 (N10731, N10720, N9839);
nand NAND2 (N10732, N10726, N9101);
xor XOR2 (N10733, N10723, N5813);
not NOT1 (N10734, N10730);
nand NAND3 (N10735, N10728, N8777, N6134);
xor XOR2 (N10736, N10734, N4805);
nor NOR2 (N10737, N10732, N7405);
xor XOR2 (N10738, N10725, N7884);
nor NOR2 (N10739, N10731, N36);
or OR3 (N10740, N10724, N3229, N1422);
and AND4 (N10741, N10737, N10591, N4959, N6156);
or OR3 (N10742, N10735, N7856, N5981);
xor XOR2 (N10743, N10638, N9394);
nor NOR3 (N10744, N10742, N3398, N6797);
or OR4 (N10745, N10743, N2224, N145, N10576);
not NOT1 (N10746, N10733);
and AND2 (N10747, N10718, N4716);
buf BUF1 (N10748, N10721);
nand NAND3 (N10749, N10740, N9933, N7118);
and AND4 (N10750, N10748, N6434, N3997, N2550);
or OR4 (N10751, N10747, N6495, N4243, N8027);
nand NAND3 (N10752, N10739, N10269, N6945);
nor NOR2 (N10753, N10744, N629);
and AND4 (N10754, N10746, N7816, N9063, N7562);
xor XOR2 (N10755, N10751, N1833);
and AND2 (N10756, N10749, N8107);
nand NAND4 (N10757, N10750, N8923, N1393, N258);
nand NAND4 (N10758, N10755, N3196, N1198, N5725);
not NOT1 (N10759, N10736);
or OR4 (N10760, N10757, N3435, N1606, N3480);
and AND2 (N10761, N10745, N446);
and AND3 (N10762, N10753, N4287, N321);
nor NOR2 (N10763, N10759, N6674);
xor XOR2 (N10764, N10761, N6500);
not NOT1 (N10765, N10764);
buf BUF1 (N10766, N10738);
or OR4 (N10767, N10765, N511, N9990, N5085);
buf BUF1 (N10768, N10767);
buf BUF1 (N10769, N10763);
or OR4 (N10770, N10756, N5163, N8455, N764);
buf BUF1 (N10771, N10766);
or OR3 (N10772, N10741, N9284, N7505);
not NOT1 (N10773, N10758);
nand NAND2 (N10774, N10769, N8680);
buf BUF1 (N10775, N10754);
nor NOR3 (N10776, N10770, N5602, N8581);
xor XOR2 (N10777, N10762, N4408);
xor XOR2 (N10778, N10772, N1740);
or OR3 (N10779, N10773, N8024, N9251);
not NOT1 (N10780, N10777);
buf BUF1 (N10781, N10768);
and AND3 (N10782, N10771, N3542, N7642);
not NOT1 (N10783, N10776);
and AND3 (N10784, N10779, N10106, N5281);
buf BUF1 (N10785, N10775);
or OR4 (N10786, N10782, N3645, N2309, N1952);
buf BUF1 (N10787, N10752);
buf BUF1 (N10788, N10778);
or OR4 (N10789, N10774, N8062, N6875, N7736);
xor XOR2 (N10790, N10785, N5048);
buf BUF1 (N10791, N10760);
and AND2 (N10792, N10790, N6045);
buf BUF1 (N10793, N10791);
xor XOR2 (N10794, N10792, N9571);
or OR4 (N10795, N10787, N1905, N3253, N2750);
buf BUF1 (N10796, N10781);
nor NOR3 (N10797, N10794, N4644, N3943);
nor NOR4 (N10798, N10786, N10723, N5179, N6228);
xor XOR2 (N10799, N10797, N1565);
xor XOR2 (N10800, N10780, N1586);
or OR3 (N10801, N10796, N9789, N5198);
xor XOR2 (N10802, N10784, N967);
buf BUF1 (N10803, N10795);
nand NAND3 (N10804, N10798, N4825, N4373);
or OR2 (N10805, N10800, N10062);
nand NAND4 (N10806, N10799, N7361, N4478, N2451);
or OR2 (N10807, N10783, N302);
or OR2 (N10808, N10807, N1711);
nor NOR2 (N10809, N10789, N8282);
or OR3 (N10810, N10805, N8436, N2200);
xor XOR2 (N10811, N10802, N2289);
and AND3 (N10812, N10811, N8861, N9957);
xor XOR2 (N10813, N10804, N5338);
or OR4 (N10814, N10810, N1752, N6693, N206);
or OR2 (N10815, N10814, N4784);
xor XOR2 (N10816, N10801, N5512);
buf BUF1 (N10817, N10803);
nor NOR4 (N10818, N10788, N2021, N644, N5545);
or OR3 (N10819, N10816, N1470, N4987);
nand NAND2 (N10820, N10813, N3286);
not NOT1 (N10821, N10808);
and AND4 (N10822, N10812, N10516, N9638, N8766);
or OR4 (N10823, N10815, N3289, N3804, N5206);
nand NAND3 (N10824, N10817, N2400, N9110);
buf BUF1 (N10825, N10821);
or OR2 (N10826, N10820, N4040);
and AND2 (N10827, N10818, N184);
and AND4 (N10828, N10809, N4583, N8911, N3786);
nor NOR4 (N10829, N10793, N9341, N8273, N155);
or OR4 (N10830, N10826, N2335, N8779, N3861);
or OR3 (N10831, N10824, N7411, N7072);
not NOT1 (N10832, N10830);
buf BUF1 (N10833, N10827);
nor NOR4 (N10834, N10833, N2078, N8406, N3277);
xor XOR2 (N10835, N10828, N10378);
nand NAND2 (N10836, N10835, N5047);
and AND4 (N10837, N10829, N5688, N8674, N4788);
xor XOR2 (N10838, N10823, N3237);
nor NOR4 (N10839, N10832, N4152, N1018, N5054);
or OR3 (N10840, N10839, N2364, N9455);
or OR4 (N10841, N10838, N2013, N1765, N2783);
buf BUF1 (N10842, N10840);
xor XOR2 (N10843, N10834, N2832);
not NOT1 (N10844, N10836);
buf BUF1 (N10845, N10822);
or OR3 (N10846, N10844, N2032, N5372);
and AND4 (N10847, N10837, N10552, N8780, N1757);
or OR3 (N10848, N10841, N2773, N9586);
nor NOR3 (N10849, N10848, N6531, N7289);
nor NOR2 (N10850, N10846, N3998);
and AND2 (N10851, N10825, N1769);
xor XOR2 (N10852, N10849, N9339);
and AND4 (N10853, N10851, N3981, N749, N2137);
buf BUF1 (N10854, N10831);
or OR2 (N10855, N10806, N1983);
and AND3 (N10856, N10855, N9764, N5199);
buf BUF1 (N10857, N10852);
buf BUF1 (N10858, N10819);
and AND4 (N10859, N10843, N10099, N3474, N9048);
not NOT1 (N10860, N10857);
and AND4 (N10861, N10856, N5304, N5136, N5362);
buf BUF1 (N10862, N10850);
and AND4 (N10863, N10859, N793, N683, N3989);
and AND4 (N10864, N10863, N4841, N9447, N4625);
and AND3 (N10865, N10864, N6469, N8633);
or OR3 (N10866, N10858, N4957, N1671);
buf BUF1 (N10867, N10861);
or OR4 (N10868, N10853, N8239, N7689, N7239);
nor NOR2 (N10869, N10867, N5082);
xor XOR2 (N10870, N10860, N7418);
nand NAND2 (N10871, N10845, N1706);
nor NOR4 (N10872, N10847, N2056, N5838, N3539);
not NOT1 (N10873, N10872);
and AND4 (N10874, N10873, N32, N10637, N8728);
not NOT1 (N10875, N10854);
not NOT1 (N10876, N10874);
not NOT1 (N10877, N10862);
xor XOR2 (N10878, N10866, N2318);
nand NAND4 (N10879, N10875, N919, N9025, N2868);
and AND3 (N10880, N10842, N9558, N8175);
buf BUF1 (N10881, N10879);
and AND4 (N10882, N10878, N427, N10150, N383);
nand NAND2 (N10883, N10880, N9082);
and AND3 (N10884, N10882, N5790, N6230);
nand NAND3 (N10885, N10876, N7913, N3049);
not NOT1 (N10886, N10883);
xor XOR2 (N10887, N10870, N10711);
nor NOR4 (N10888, N10871, N758, N9145, N10478);
and AND4 (N10889, N10885, N2364, N3053, N1154);
nand NAND2 (N10890, N10887, N7177);
not NOT1 (N10891, N10886);
xor XOR2 (N10892, N10890, N5938);
xor XOR2 (N10893, N10884, N1361);
not NOT1 (N10894, N10891);
or OR3 (N10895, N10888, N4391, N5790);
nand NAND2 (N10896, N10892, N1385);
xor XOR2 (N10897, N10877, N2363);
or OR2 (N10898, N10893, N10465);
nand NAND2 (N10899, N10894, N9542);
not NOT1 (N10900, N10895);
xor XOR2 (N10901, N10899, N6860);
not NOT1 (N10902, N10869);
nand NAND3 (N10903, N10900, N7768, N10692);
xor XOR2 (N10904, N10897, N7152);
and AND4 (N10905, N10896, N10098, N8321, N9085);
or OR3 (N10906, N10889, N3089, N3988);
nor NOR2 (N10907, N10868, N9933);
not NOT1 (N10908, N10865);
not NOT1 (N10909, N10903);
nor NOR3 (N10910, N10906, N4966, N9557);
not NOT1 (N10911, N10908);
not NOT1 (N10912, N10904);
not NOT1 (N10913, N10910);
not NOT1 (N10914, N10905);
nor NOR2 (N10915, N10911, N7812);
buf BUF1 (N10916, N10913);
buf BUF1 (N10917, N10909);
not NOT1 (N10918, N10902);
buf BUF1 (N10919, N10898);
nor NOR3 (N10920, N10914, N8234, N5781);
and AND3 (N10921, N10912, N5766, N7936);
nand NAND4 (N10922, N10901, N3701, N6286, N5384);
nand NAND3 (N10923, N10916, N6677, N8331);
buf BUF1 (N10924, N10918);
or OR4 (N10925, N10920, N9494, N725, N10289);
nand NAND2 (N10926, N10921, N7702);
nor NOR2 (N10927, N10919, N5570);
or OR4 (N10928, N10924, N5099, N10708, N1798);
or OR3 (N10929, N10926, N9365, N4691);
nor NOR3 (N10930, N10917, N5381, N10448);
xor XOR2 (N10931, N10928, N7595);
nor NOR4 (N10932, N10881, N1889, N7886, N3622);
buf BUF1 (N10933, N10922);
buf BUF1 (N10934, N10925);
xor XOR2 (N10935, N10907, N5755);
and AND3 (N10936, N10931, N7997, N4200);
xor XOR2 (N10937, N10927, N6051);
nor NOR3 (N10938, N10930, N5141, N7349);
nor NOR2 (N10939, N10934, N10007);
and AND4 (N10940, N10935, N6308, N767, N2847);
and AND3 (N10941, N10939, N8395, N619);
xor XOR2 (N10942, N10936, N1270);
and AND3 (N10943, N10941, N277, N9156);
xor XOR2 (N10944, N10915, N5206);
nand NAND4 (N10945, N10944, N814, N3173, N6570);
buf BUF1 (N10946, N10940);
not NOT1 (N10947, N10929);
xor XOR2 (N10948, N10932, N1443);
not NOT1 (N10949, N10948);
nand NAND3 (N10950, N10949, N2691, N8967);
xor XOR2 (N10951, N10937, N242);
buf BUF1 (N10952, N10951);
nor NOR4 (N10953, N10945, N10267, N8934, N2242);
xor XOR2 (N10954, N10923, N5737);
buf BUF1 (N10955, N10952);
nor NOR2 (N10956, N10946, N8396);
xor XOR2 (N10957, N10943, N765);
not NOT1 (N10958, N10954);
nor NOR3 (N10959, N10956, N3479, N5029);
nor NOR3 (N10960, N10947, N1219, N6745);
xor XOR2 (N10961, N10955, N918);
not NOT1 (N10962, N10961);
and AND4 (N10963, N10950, N167, N6599, N6861);
not NOT1 (N10964, N10933);
nand NAND3 (N10965, N10964, N1414, N1718);
or OR2 (N10966, N10960, N7519);
not NOT1 (N10967, N10958);
or OR4 (N10968, N10959, N5478, N4830, N7060);
and AND3 (N10969, N10965, N9741, N9527);
and AND2 (N10970, N10938, N2219);
not NOT1 (N10971, N10966);
or OR4 (N10972, N10963, N4409, N7920, N7828);
or OR2 (N10973, N10957, N3403);
xor XOR2 (N10974, N10969, N2459);
nand NAND3 (N10975, N10974, N5887, N8796);
not NOT1 (N10976, N10962);
nand NAND3 (N10977, N10942, N3419, N3196);
buf BUF1 (N10978, N10976);
xor XOR2 (N10979, N10973, N5116);
nor NOR2 (N10980, N10953, N1665);
xor XOR2 (N10981, N10972, N452);
nor NOR4 (N10982, N10980, N1445, N786, N1866);
buf BUF1 (N10983, N10967);
nor NOR3 (N10984, N10982, N3135, N4371);
not NOT1 (N10985, N10970);
not NOT1 (N10986, N10968);
nand NAND4 (N10987, N10971, N1875, N10520, N5768);
xor XOR2 (N10988, N10975, N3411);
nor NOR2 (N10989, N10988, N626);
nor NOR4 (N10990, N10981, N720, N4490, N4921);
not NOT1 (N10991, N10986);
nand NAND4 (N10992, N10991, N9569, N7625, N2487);
xor XOR2 (N10993, N10987, N1379);
nor NOR3 (N10994, N10993, N984, N6862);
and AND4 (N10995, N10983, N10796, N215, N8013);
nor NOR2 (N10996, N10989, N1764);
not NOT1 (N10997, N10977);
not NOT1 (N10998, N10995);
xor XOR2 (N10999, N10994, N4118);
and AND3 (N11000, N10985, N784, N5576);
xor XOR2 (N11001, N10998, N697);
buf BUF1 (N11002, N10990);
xor XOR2 (N11003, N10999, N8304);
buf BUF1 (N11004, N10997);
and AND2 (N11005, N11000, N6974);
nor NOR3 (N11006, N11005, N7908, N583);
buf BUF1 (N11007, N11002);
nand NAND3 (N11008, N10992, N9105, N3885);
buf BUF1 (N11009, N11004);
nor NOR3 (N11010, N11006, N648, N6140);
nand NAND2 (N11011, N11009, N10435);
or OR2 (N11012, N11008, N5472);
xor XOR2 (N11013, N10979, N4427);
not NOT1 (N11014, N10996);
nor NOR4 (N11015, N11013, N33, N4846, N9260);
or OR4 (N11016, N11014, N2743, N4171, N7274);
and AND3 (N11017, N11012, N3123, N3569);
nand NAND2 (N11018, N10984, N847);
nor NOR4 (N11019, N11001, N2425, N7601, N7791);
not NOT1 (N11020, N11010);
or OR2 (N11021, N11003, N4588);
and AND2 (N11022, N11021, N1211);
buf BUF1 (N11023, N11022);
nand NAND2 (N11024, N11023, N8198);
buf BUF1 (N11025, N11019);
and AND3 (N11026, N11007, N8012, N6415);
not NOT1 (N11027, N11011);
xor XOR2 (N11028, N11027, N2109);
nand NAND4 (N11029, N11024, N6646, N374, N4);
buf BUF1 (N11030, N11015);
buf BUF1 (N11031, N11026);
or OR3 (N11032, N11025, N3427, N10262);
or OR2 (N11033, N11031, N7138);
or OR2 (N11034, N11016, N2236);
and AND2 (N11035, N11020, N8867);
not NOT1 (N11036, N11028);
xor XOR2 (N11037, N11029, N1817);
or OR2 (N11038, N11036, N5219);
not NOT1 (N11039, N11037);
buf BUF1 (N11040, N11032);
xor XOR2 (N11041, N11035, N5302);
nor NOR4 (N11042, N11040, N5625, N5741, N4960);
and AND3 (N11043, N11038, N10966, N8417);
nor NOR2 (N11044, N11041, N4177);
nor NOR3 (N11045, N11034, N5309, N7952);
not NOT1 (N11046, N11018);
xor XOR2 (N11047, N11030, N356);
nor NOR3 (N11048, N11047, N7766, N2899);
not NOT1 (N11049, N11033);
and AND2 (N11050, N11046, N6595);
xor XOR2 (N11051, N11042, N586);
and AND3 (N11052, N11045, N99, N7509);
or OR2 (N11053, N11052, N4111);
nand NAND4 (N11054, N11053, N9210, N9047, N9622);
nand NAND4 (N11055, N11048, N9371, N2834, N8436);
xor XOR2 (N11056, N11044, N1903);
or OR4 (N11057, N11049, N10385, N1557, N10318);
buf BUF1 (N11058, N11055);
xor XOR2 (N11059, N11057, N942);
and AND3 (N11060, N10978, N6174, N2940);
nor NOR4 (N11061, N11039, N3200, N8495, N3453);
buf BUF1 (N11062, N11051);
nor NOR4 (N11063, N11058, N7267, N10522, N9333);
or OR4 (N11064, N11056, N10234, N8292, N1731);
nor NOR2 (N11065, N11043, N2427);
nor NOR4 (N11066, N11050, N3855, N6598, N4060);
and AND3 (N11067, N11017, N6774, N8768);
or OR4 (N11068, N11067, N10863, N10672, N10678);
nor NOR3 (N11069, N11059, N162, N4710);
buf BUF1 (N11070, N11054);
and AND3 (N11071, N11070, N10268, N9221);
nor NOR3 (N11072, N11061, N725, N6932);
not NOT1 (N11073, N11072);
not NOT1 (N11074, N11060);
not NOT1 (N11075, N11071);
buf BUF1 (N11076, N11075);
xor XOR2 (N11077, N11073, N4101);
buf BUF1 (N11078, N11064);
or OR2 (N11079, N11066, N1819);
or OR3 (N11080, N11069, N8459, N7256);
buf BUF1 (N11081, N11074);
xor XOR2 (N11082, N11079, N5144);
nand NAND2 (N11083, N11080, N636);
buf BUF1 (N11084, N11083);
nor NOR4 (N11085, N11082, N6902, N9028, N10054);
or OR2 (N11086, N11077, N8033);
nor NOR4 (N11087, N11076, N9786, N3563, N4229);
and AND2 (N11088, N11062, N1974);
not NOT1 (N11089, N11063);
not NOT1 (N11090, N11068);
nor NOR4 (N11091, N11081, N9676, N2549, N2491);
nor NOR3 (N11092, N11065, N6147, N6174);
not NOT1 (N11093, N11089);
or OR3 (N11094, N11085, N8505, N10735);
nor NOR4 (N11095, N11086, N8075, N3995, N3391);
nand NAND3 (N11096, N11092, N7396, N7424);
and AND4 (N11097, N11091, N3020, N3719, N8857);
xor XOR2 (N11098, N11097, N1140);
nand NAND2 (N11099, N11093, N8185);
and AND4 (N11100, N11084, N9403, N2395, N810);
not NOT1 (N11101, N11090);
buf BUF1 (N11102, N11078);
buf BUF1 (N11103, N11087);
xor XOR2 (N11104, N11101, N8397);
not NOT1 (N11105, N11100);
nor NOR4 (N11106, N11096, N10441, N10937, N3424);
nor NOR2 (N11107, N11088, N2306);
and AND4 (N11108, N11103, N4990, N4275, N10715);
buf BUF1 (N11109, N11105);
nor NOR3 (N11110, N11108, N5936, N6707);
or OR4 (N11111, N11099, N10080, N4479, N1674);
not NOT1 (N11112, N11111);
and AND4 (N11113, N11107, N748, N2415, N8678);
buf BUF1 (N11114, N11094);
not NOT1 (N11115, N11109);
nor NOR2 (N11116, N11112, N5355);
nor NOR2 (N11117, N11110, N7185);
not NOT1 (N11118, N11098);
not NOT1 (N11119, N11104);
and AND4 (N11120, N11115, N1236, N7169, N2255);
nand NAND4 (N11121, N11102, N4891, N291, N758);
and AND3 (N11122, N11118, N76, N10359);
xor XOR2 (N11123, N11116, N3683);
not NOT1 (N11124, N11114);
nand NAND3 (N11125, N11119, N1895, N2878);
not NOT1 (N11126, N11113);
or OR2 (N11127, N11117, N718);
buf BUF1 (N11128, N11124);
not NOT1 (N11129, N11123);
and AND2 (N11130, N11122, N8616);
or OR2 (N11131, N11127, N6512);
nand NAND2 (N11132, N11129, N3019);
and AND2 (N11133, N11130, N10697);
nor NOR2 (N11134, N11131, N359);
nor NOR4 (N11135, N11133, N2550, N8106, N937);
and AND4 (N11136, N11135, N1002, N3187, N2463);
and AND2 (N11137, N11095, N166);
nand NAND3 (N11138, N11132, N9464, N2458);
or OR3 (N11139, N11125, N5662, N7516);
nand NAND2 (N11140, N11136, N785);
xor XOR2 (N11141, N11138, N2891);
nand NAND4 (N11142, N11139, N9345, N3090, N6151);
nand NAND2 (N11143, N11126, N3057);
nor NOR2 (N11144, N11142, N1184);
not NOT1 (N11145, N11137);
nor NOR2 (N11146, N11141, N8687);
nand NAND3 (N11147, N11121, N3366, N8364);
nor NOR2 (N11148, N11128, N7432);
xor XOR2 (N11149, N11147, N6693);
nor NOR2 (N11150, N11106, N3818);
nand NAND4 (N11151, N11150, N1925, N2271, N4553);
buf BUF1 (N11152, N11149);
and AND3 (N11153, N11148, N9153, N7746);
not NOT1 (N11154, N11153);
buf BUF1 (N11155, N11134);
or OR3 (N11156, N11152, N1878, N10612);
buf BUF1 (N11157, N11155);
nor NOR4 (N11158, N11143, N3854, N7174, N8889);
nor NOR3 (N11159, N11120, N9192, N5775);
nor NOR4 (N11160, N11151, N280, N236, N353);
xor XOR2 (N11161, N11158, N11129);
buf BUF1 (N11162, N11161);
not NOT1 (N11163, N11144);
xor XOR2 (N11164, N11140, N9015);
buf BUF1 (N11165, N11164);
and AND4 (N11166, N11154, N3818, N3575, N9937);
nand NAND2 (N11167, N11145, N3141);
nand NAND3 (N11168, N11166, N5797, N8890);
not NOT1 (N11169, N11165);
not NOT1 (N11170, N11169);
xor XOR2 (N11171, N11156, N10218);
or OR3 (N11172, N11163, N5318, N1992);
nand NAND3 (N11173, N11157, N2523, N350);
buf BUF1 (N11174, N11162);
nand NAND3 (N11175, N11160, N5788, N7439);
nor NOR4 (N11176, N11146, N770, N5835, N6395);
buf BUF1 (N11177, N11170);
nor NOR3 (N11178, N11168, N2939, N9801);
not NOT1 (N11179, N11167);
nand NAND3 (N11180, N11174, N3724, N5402);
xor XOR2 (N11181, N11175, N1184);
nand NAND2 (N11182, N11181, N1863);
nand NAND3 (N11183, N11179, N7095, N4932);
nand NAND2 (N11184, N11183, N9271);
xor XOR2 (N11185, N11182, N5818);
and AND2 (N11186, N11171, N8564);
nor NOR3 (N11187, N11177, N4290, N4190);
not NOT1 (N11188, N11180);
not NOT1 (N11189, N11188);
buf BUF1 (N11190, N11187);
nand NAND3 (N11191, N11178, N9042, N7151);
nor NOR4 (N11192, N11189, N2633, N9296, N8276);
not NOT1 (N11193, N11159);
or OR3 (N11194, N11184, N5429, N7365);
nand NAND3 (N11195, N11185, N6521, N1188);
xor XOR2 (N11196, N11191, N7337);
xor XOR2 (N11197, N11194, N4764);
buf BUF1 (N11198, N11195);
and AND4 (N11199, N11186, N10965, N85, N7174);
nand NAND2 (N11200, N11196, N6729);
not NOT1 (N11201, N11200);
nor NOR2 (N11202, N11201, N10227);
or OR3 (N11203, N11190, N8303, N3077);
not NOT1 (N11204, N11173);
xor XOR2 (N11205, N11202, N7418);
and AND3 (N11206, N11199, N7049, N3028);
xor XOR2 (N11207, N11197, N5741);
xor XOR2 (N11208, N11205, N9958);
nor NOR4 (N11209, N11204, N8624, N8494, N5307);
or OR4 (N11210, N11193, N2481, N7381, N8814);
nor NOR2 (N11211, N11207, N10357);
buf BUF1 (N11212, N11198);
buf BUF1 (N11213, N11212);
or OR2 (N11214, N11213, N7997);
xor XOR2 (N11215, N11208, N5631);
nor NOR2 (N11216, N11209, N8241);
nor NOR3 (N11217, N11210, N1172, N1945);
nand NAND2 (N11218, N11215, N2549);
xor XOR2 (N11219, N11172, N4207);
xor XOR2 (N11220, N11216, N9494);
or OR3 (N11221, N11220, N6760, N10001);
buf BUF1 (N11222, N11192);
buf BUF1 (N11223, N11221);
nor NOR3 (N11224, N11223, N2266, N9569);
or OR4 (N11225, N11218, N7571, N6917, N10816);
xor XOR2 (N11226, N11219, N4400);
nand NAND2 (N11227, N11214, N9577);
not NOT1 (N11228, N11211);
nand NAND2 (N11229, N11176, N8252);
buf BUF1 (N11230, N11217);
or OR4 (N11231, N11230, N9521, N6796, N10847);
nand NAND4 (N11232, N11229, N1779, N8902, N3128);
not NOT1 (N11233, N11231);
and AND3 (N11234, N11206, N1433, N793);
nor NOR4 (N11235, N11203, N2137, N10634, N3869);
nor NOR2 (N11236, N11235, N10086);
or OR2 (N11237, N11227, N6408);
not NOT1 (N11238, N11226);
nor NOR2 (N11239, N11232, N11030);
nor NOR4 (N11240, N11233, N2730, N72, N10567);
nand NAND3 (N11241, N11236, N1508, N5493);
nor NOR3 (N11242, N11224, N4296, N6283);
xor XOR2 (N11243, N11237, N8648);
nand NAND4 (N11244, N11241, N6166, N364, N5792);
not NOT1 (N11245, N11244);
buf BUF1 (N11246, N11234);
buf BUF1 (N11247, N11225);
not NOT1 (N11248, N11246);
buf BUF1 (N11249, N11222);
xor XOR2 (N11250, N11240, N7281);
nor NOR3 (N11251, N11249, N8874, N1660);
and AND4 (N11252, N11239, N1978, N2020, N3123);
buf BUF1 (N11253, N11238);
nand NAND2 (N11254, N11243, N4686);
nand NAND4 (N11255, N11242, N25, N8422, N9759);
not NOT1 (N11256, N11248);
xor XOR2 (N11257, N11254, N4715);
buf BUF1 (N11258, N11252);
not NOT1 (N11259, N11228);
nor NOR3 (N11260, N11257, N942, N3349);
buf BUF1 (N11261, N11247);
not NOT1 (N11262, N11256);
buf BUF1 (N11263, N11255);
or OR3 (N11264, N11260, N7756, N10484);
and AND4 (N11265, N11261, N1139, N1094, N7982);
xor XOR2 (N11266, N11245, N9875);
nand NAND4 (N11267, N11251, N426, N5701, N7338);
or OR2 (N11268, N11264, N2800);
xor XOR2 (N11269, N11267, N3496);
nand NAND2 (N11270, N11250, N606);
nor NOR3 (N11271, N11266, N6320, N7598);
nand NAND2 (N11272, N11259, N6337);
and AND3 (N11273, N11263, N9895, N1347);
and AND2 (N11274, N11273, N3519);
and AND3 (N11275, N11271, N1962, N121);
buf BUF1 (N11276, N11265);
xor XOR2 (N11277, N11269, N11202);
nand NAND3 (N11278, N11276, N6989, N4732);
and AND2 (N11279, N11258, N10793);
nand NAND4 (N11280, N11262, N4835, N10921, N812);
nor NOR3 (N11281, N11272, N6129, N4590);
not NOT1 (N11282, N11281);
or OR3 (N11283, N11280, N7323, N1854);
nand NAND4 (N11284, N11270, N720, N7812, N449);
or OR3 (N11285, N11253, N4482, N2773);
nand NAND4 (N11286, N11283, N6883, N4386, N1486);
nand NAND2 (N11287, N11275, N3129);
nand NAND2 (N11288, N11278, N9410);
xor XOR2 (N11289, N11274, N5557);
buf BUF1 (N11290, N11268);
xor XOR2 (N11291, N11288, N4470);
buf BUF1 (N11292, N11284);
not NOT1 (N11293, N11292);
xor XOR2 (N11294, N11291, N9142);
nor NOR2 (N11295, N11287, N6425);
not NOT1 (N11296, N11293);
xor XOR2 (N11297, N11282, N7405);
nor NOR4 (N11298, N11277, N1668, N9504, N6733);
nor NOR3 (N11299, N11290, N9743, N1151);
xor XOR2 (N11300, N11285, N6702);
nand NAND3 (N11301, N11279, N6241, N1945);
or OR2 (N11302, N11297, N2136);
and AND2 (N11303, N11296, N9998);
not NOT1 (N11304, N11300);
nor NOR4 (N11305, N11286, N3969, N457, N5416);
not NOT1 (N11306, N11298);
or OR3 (N11307, N11305, N7103, N796);
buf BUF1 (N11308, N11307);
not NOT1 (N11309, N11308);
nand NAND2 (N11310, N11299, N9963);
and AND3 (N11311, N11295, N6593, N9951);
nand NAND2 (N11312, N11311, N4476);
nor NOR4 (N11313, N11301, N4807, N5542, N5698);
or OR3 (N11314, N11313, N3360, N547);
nand NAND3 (N11315, N11306, N9086, N10859);
nor NOR4 (N11316, N11315, N10750, N2735, N4071);
and AND4 (N11317, N11310, N9657, N3265, N10942);
nand NAND2 (N11318, N11316, N5542);
nand NAND4 (N11319, N11294, N10144, N6926, N8063);
nor NOR4 (N11320, N11319, N5218, N6045, N7810);
nor NOR3 (N11321, N11314, N9551, N6821);
xor XOR2 (N11322, N11320, N684);
nand NAND4 (N11323, N11322, N8774, N3539, N5525);
nand NAND2 (N11324, N11289, N8955);
not NOT1 (N11325, N11309);
nand NAND3 (N11326, N11318, N148, N7100);
and AND2 (N11327, N11324, N1242);
not NOT1 (N11328, N11323);
buf BUF1 (N11329, N11303);
xor XOR2 (N11330, N11304, N5619);
not NOT1 (N11331, N11317);
not NOT1 (N11332, N11329);
buf BUF1 (N11333, N11312);
xor XOR2 (N11334, N11330, N2956);
or OR2 (N11335, N11334, N7238);
or OR3 (N11336, N11335, N1103, N5684);
and AND4 (N11337, N11321, N10486, N1134, N9461);
not NOT1 (N11338, N11332);
not NOT1 (N11339, N11325);
and AND4 (N11340, N11336, N10527, N10070, N10133);
and AND3 (N11341, N11333, N9889, N406);
buf BUF1 (N11342, N11339);
nand NAND2 (N11343, N11326, N10173);
not NOT1 (N11344, N11337);
nor NOR4 (N11345, N11343, N1650, N2127, N4269);
nor NOR2 (N11346, N11340, N4113);
nand NAND3 (N11347, N11327, N8651, N4792);
nor NOR4 (N11348, N11341, N7935, N2853, N9513);
xor XOR2 (N11349, N11338, N5359);
nand NAND2 (N11350, N11344, N5972);
nor NOR3 (N11351, N11302, N2979, N4082);
xor XOR2 (N11352, N11342, N712);
xor XOR2 (N11353, N11348, N2716);
nand NAND3 (N11354, N11347, N8236, N4296);
and AND4 (N11355, N11351, N5797, N2996, N7277);
buf BUF1 (N11356, N11349);
nor NOR4 (N11357, N11355, N10838, N1428, N910);
buf BUF1 (N11358, N11346);
nand NAND2 (N11359, N11358, N2136);
and AND3 (N11360, N11356, N7842, N5951);
buf BUF1 (N11361, N11360);
and AND2 (N11362, N11359, N9675);
nand NAND3 (N11363, N11357, N3510, N9636);
or OR4 (N11364, N11353, N9731, N9750, N3295);
not NOT1 (N11365, N11331);
buf BUF1 (N11366, N11354);
or OR2 (N11367, N11361, N6575);
xor XOR2 (N11368, N11365, N11065);
not NOT1 (N11369, N11328);
and AND4 (N11370, N11350, N7395, N6602, N6894);
xor XOR2 (N11371, N11363, N2294);
buf BUF1 (N11372, N11352);
nand NAND3 (N11373, N11368, N7153, N770);
or OR3 (N11374, N11373, N2855, N11117);
not NOT1 (N11375, N11364);
buf BUF1 (N11376, N11374);
nor NOR3 (N11377, N11375, N5523, N4812);
not NOT1 (N11378, N11372);
or OR4 (N11379, N11378, N10457, N5076, N5140);
buf BUF1 (N11380, N11376);
xor XOR2 (N11381, N11370, N3915);
nor NOR3 (N11382, N11345, N9814, N10809);
and AND3 (N11383, N11371, N5263, N3627);
or OR4 (N11384, N11379, N3213, N6257, N3452);
and AND2 (N11385, N11383, N10929);
buf BUF1 (N11386, N11382);
nand NAND3 (N11387, N11386, N10146, N6982);
xor XOR2 (N11388, N11369, N9936);
xor XOR2 (N11389, N11380, N2175);
or OR2 (N11390, N11381, N2316);
or OR3 (N11391, N11385, N10319, N6461);
nor NOR4 (N11392, N11384, N5024, N270, N3826);
or OR4 (N11393, N11387, N990, N2461, N9103);
buf BUF1 (N11394, N11362);
nand NAND4 (N11395, N11367, N7953, N6460, N8586);
or OR4 (N11396, N11377, N5276, N6311, N6994);
nand NAND2 (N11397, N11366, N9987);
buf BUF1 (N11398, N11395);
and AND2 (N11399, N11396, N7598);
buf BUF1 (N11400, N11390);
not NOT1 (N11401, N11398);
not NOT1 (N11402, N11397);
xor XOR2 (N11403, N11389, N4898);
xor XOR2 (N11404, N11391, N3347);
and AND4 (N11405, N11400, N10190, N3096, N8112);
buf BUF1 (N11406, N11393);
and AND2 (N11407, N11403, N1271);
nand NAND2 (N11408, N11394, N10597);
nand NAND2 (N11409, N11406, N4614);
nor NOR2 (N11410, N11401, N3478);
buf BUF1 (N11411, N11399);
nand NAND3 (N11412, N11405, N2807, N2941);
xor XOR2 (N11413, N11404, N8674);
or OR2 (N11414, N11409, N5626);
not NOT1 (N11415, N11412);
not NOT1 (N11416, N11415);
xor XOR2 (N11417, N11416, N3508);
xor XOR2 (N11418, N11407, N1058);
nor NOR2 (N11419, N11417, N3086);
buf BUF1 (N11420, N11402);
nand NAND3 (N11421, N11392, N8999, N9272);
not NOT1 (N11422, N11411);
not NOT1 (N11423, N11422);
nor NOR3 (N11424, N11414, N5590, N3994);
and AND2 (N11425, N11424, N9385);
xor XOR2 (N11426, N11419, N3759);
xor XOR2 (N11427, N11426, N9057);
not NOT1 (N11428, N11427);
or OR4 (N11429, N11420, N9874, N10952, N9981);
and AND4 (N11430, N11388, N2257, N8760, N7953);
xor XOR2 (N11431, N11413, N155);
not NOT1 (N11432, N11425);
nor NOR2 (N11433, N11432, N6934);
not NOT1 (N11434, N11428);
or OR2 (N11435, N11418, N4272);
xor XOR2 (N11436, N11433, N5901);
nor NOR3 (N11437, N11435, N10405, N2807);
nor NOR3 (N11438, N11423, N8984, N1709);
xor XOR2 (N11439, N11436, N7004);
or OR4 (N11440, N11410, N4109, N10818, N8354);
and AND4 (N11441, N11429, N5391, N1397, N3246);
xor XOR2 (N11442, N11431, N7247);
not NOT1 (N11443, N11434);
nand NAND4 (N11444, N11438, N2262, N11334, N2835);
xor XOR2 (N11445, N11430, N7478);
buf BUF1 (N11446, N11437);
or OR4 (N11447, N11440, N7129, N4928, N931);
xor XOR2 (N11448, N11439, N9778);
and AND3 (N11449, N11445, N11210, N42);
buf BUF1 (N11450, N11408);
nand NAND3 (N11451, N11442, N6493, N413);
and AND4 (N11452, N11446, N1495, N6276, N8960);
buf BUF1 (N11453, N11443);
or OR2 (N11454, N11452, N1129);
nand NAND4 (N11455, N11447, N3745, N1317, N4712);
nand NAND2 (N11456, N11421, N8799);
not NOT1 (N11457, N11454);
xor XOR2 (N11458, N11451, N10656);
xor XOR2 (N11459, N11450, N812);
not NOT1 (N11460, N11458);
not NOT1 (N11461, N11441);
buf BUF1 (N11462, N11448);
not NOT1 (N11463, N11461);
not NOT1 (N11464, N11453);
nor NOR3 (N11465, N11463, N6631, N2843);
buf BUF1 (N11466, N11444);
and AND2 (N11467, N11460, N3479);
or OR2 (N11468, N11459, N8500);
not NOT1 (N11469, N11457);
xor XOR2 (N11470, N11464, N4127);
xor XOR2 (N11471, N11462, N10526);
not NOT1 (N11472, N11449);
nor NOR3 (N11473, N11470, N2167, N9607);
nand NAND3 (N11474, N11456, N7460, N6585);
or OR3 (N11475, N11469, N3982, N5999);
buf BUF1 (N11476, N11467);
and AND2 (N11477, N11472, N9478);
buf BUF1 (N11478, N11476);
buf BUF1 (N11479, N11471);
buf BUF1 (N11480, N11465);
nor NOR2 (N11481, N11475, N2979);
not NOT1 (N11482, N11455);
nor NOR3 (N11483, N11468, N5273, N10978);
or OR2 (N11484, N11474, N329);
nand NAND4 (N11485, N11466, N803, N2853, N6696);
not NOT1 (N11486, N11473);
buf BUF1 (N11487, N11480);
nor NOR4 (N11488, N11482, N5247, N488, N1017);
not NOT1 (N11489, N11477);
nor NOR2 (N11490, N11488, N11067);
nor NOR3 (N11491, N11481, N5988, N141);
buf BUF1 (N11492, N11486);
or OR3 (N11493, N11492, N7836, N5050);
and AND3 (N11494, N11483, N6613, N38);
and AND3 (N11495, N11494, N7188, N1236);
nand NAND2 (N11496, N11485, N5589);
and AND4 (N11497, N11489, N5742, N4945, N3359);
nor NOR4 (N11498, N11493, N1328, N4396, N5484);
nor NOR3 (N11499, N11496, N6893, N9872);
xor XOR2 (N11500, N11479, N4852);
nor NOR3 (N11501, N11499, N9702, N7519);
nor NOR3 (N11502, N11495, N10923, N10227);
buf BUF1 (N11503, N11478);
buf BUF1 (N11504, N11500);
nand NAND4 (N11505, N11503, N5264, N10094, N2744);
not NOT1 (N11506, N11501);
xor XOR2 (N11507, N11506, N2667);
xor XOR2 (N11508, N11498, N5102);
or OR2 (N11509, N11502, N9002);
or OR4 (N11510, N11509, N5292, N7076, N2429);
buf BUF1 (N11511, N11510);
not NOT1 (N11512, N11487);
nand NAND3 (N11513, N11484, N549, N10624);
nor NOR4 (N11514, N11491, N4058, N7318, N10396);
nand NAND4 (N11515, N11490, N425, N8249, N3787);
not NOT1 (N11516, N11508);
or OR4 (N11517, N11504, N6640, N1743, N5000);
nand NAND2 (N11518, N11497, N8233);
xor XOR2 (N11519, N11511, N9600);
and AND3 (N11520, N11518, N9497, N1693);
not NOT1 (N11521, N11520);
nand NAND4 (N11522, N11507, N5987, N8616, N9196);
nor NOR3 (N11523, N11512, N5792, N3853);
not NOT1 (N11524, N11515);
and AND2 (N11525, N11514, N8280);
or OR4 (N11526, N11519, N5111, N8352, N5817);
and AND3 (N11527, N11524, N1257, N11412);
not NOT1 (N11528, N11505);
buf BUF1 (N11529, N11523);
xor XOR2 (N11530, N11528, N7312);
and AND2 (N11531, N11522, N706);
xor XOR2 (N11532, N11517, N8028);
nand NAND4 (N11533, N11513, N10886, N10099, N5023);
not NOT1 (N11534, N11525);
or OR3 (N11535, N11530, N3573, N7574);
nand NAND3 (N11536, N11526, N2884, N7676);
nand NAND3 (N11537, N11533, N3957, N9252);
nor NOR3 (N11538, N11536, N5045, N664);
or OR3 (N11539, N11516, N3929, N5646);
not NOT1 (N11540, N11537);
nand NAND3 (N11541, N11531, N889, N4533);
not NOT1 (N11542, N11529);
nand NAND3 (N11543, N11539, N10023, N2790);
nor NOR3 (N11544, N11540, N770, N194);
nor NOR3 (N11545, N11527, N6796, N2685);
or OR3 (N11546, N11543, N7370, N1002);
xor XOR2 (N11547, N11545, N8531);
not NOT1 (N11548, N11521);
xor XOR2 (N11549, N11541, N2374);
and AND2 (N11550, N11532, N11414);
nor NOR3 (N11551, N11542, N1226, N97);
or OR4 (N11552, N11535, N6901, N659, N7918);
not NOT1 (N11553, N11551);
or OR2 (N11554, N11549, N5513);
or OR3 (N11555, N11552, N10040, N257);
not NOT1 (N11556, N11546);
buf BUF1 (N11557, N11548);
and AND3 (N11558, N11556, N5482, N2861);
or OR3 (N11559, N11557, N3214, N1101);
not NOT1 (N11560, N11558);
nor NOR2 (N11561, N11547, N9701);
buf BUF1 (N11562, N11534);
or OR2 (N11563, N11555, N4789);
nand NAND2 (N11564, N11562, N3716);
buf BUF1 (N11565, N11538);
nor NOR3 (N11566, N11563, N9621, N3714);
not NOT1 (N11567, N11550);
or OR2 (N11568, N11561, N1305);
nor NOR3 (N11569, N11553, N4146, N134);
not NOT1 (N11570, N11568);
nand NAND4 (N11571, N11567, N7028, N3899, N8253);
buf BUF1 (N11572, N11564);
nand NAND2 (N11573, N11554, N10213);
xor XOR2 (N11574, N11559, N8787);
buf BUF1 (N11575, N11572);
xor XOR2 (N11576, N11573, N9603);
not NOT1 (N11577, N11565);
not NOT1 (N11578, N11569);
xor XOR2 (N11579, N11574, N7407);
nor NOR3 (N11580, N11544, N933, N8722);
xor XOR2 (N11581, N11566, N3890);
and AND3 (N11582, N11581, N3025, N7261);
nor NOR4 (N11583, N11576, N11522, N2345, N9393);
nor NOR4 (N11584, N11570, N2990, N7475, N6246);
and AND4 (N11585, N11582, N6811, N6932, N4373);
and AND3 (N11586, N11579, N1573, N1646);
buf BUF1 (N11587, N11578);
not NOT1 (N11588, N11580);
and AND2 (N11589, N11585, N2066);
nor NOR4 (N11590, N11586, N6102, N5684, N3340);
buf BUF1 (N11591, N11560);
not NOT1 (N11592, N11583);
or OR2 (N11593, N11591, N6915);
buf BUF1 (N11594, N11590);
nand NAND4 (N11595, N11571, N3990, N10065, N10614);
nand NAND2 (N11596, N11587, N7635);
and AND2 (N11597, N11595, N480);
or OR2 (N11598, N11597, N1063);
not NOT1 (N11599, N11596);
xor XOR2 (N11600, N11584, N5159);
buf BUF1 (N11601, N11588);
xor XOR2 (N11602, N11599, N6868);
not NOT1 (N11603, N11602);
nor NOR4 (N11604, N11577, N6637, N7463, N8447);
or OR3 (N11605, N11598, N5916, N1664);
not NOT1 (N11606, N11575);
or OR4 (N11607, N11593, N3091, N3582, N1974);
nor NOR2 (N11608, N11601, N1982);
buf BUF1 (N11609, N11600);
nand NAND4 (N11610, N11589, N3524, N3564, N9655);
nand NAND2 (N11611, N11608, N9259);
and AND2 (N11612, N11604, N5823);
nor NOR3 (N11613, N11607, N3872, N4865);
nor NOR4 (N11614, N11613, N11526, N6631, N4240);
nor NOR4 (N11615, N11611, N2656, N10871, N4311);
xor XOR2 (N11616, N11610, N1607);
not NOT1 (N11617, N11603);
not NOT1 (N11618, N11616);
nor NOR3 (N11619, N11615, N2474, N3648);
nand NAND3 (N11620, N11612, N6296, N5555);
xor XOR2 (N11621, N11617, N11155);
nor NOR2 (N11622, N11619, N7094);
and AND4 (N11623, N11621, N10474, N5092, N667);
not NOT1 (N11624, N11623);
nand NAND3 (N11625, N11605, N3820, N10935);
nor NOR2 (N11626, N11609, N2396);
nor NOR2 (N11627, N11624, N5305);
nand NAND3 (N11628, N11614, N4979, N11140);
and AND3 (N11629, N11625, N4825, N9194);
and AND3 (N11630, N11627, N4234, N9375);
and AND4 (N11631, N11606, N2570, N10250, N3269);
not NOT1 (N11632, N11622);
not NOT1 (N11633, N11630);
and AND3 (N11634, N11631, N8149, N6636);
xor XOR2 (N11635, N11632, N11065);
xor XOR2 (N11636, N11629, N5728);
nor NOR2 (N11637, N11635, N570);
buf BUF1 (N11638, N11592);
not NOT1 (N11639, N11637);
nor NOR3 (N11640, N11618, N1376, N2863);
nor NOR4 (N11641, N11638, N6910, N10887, N7038);
not NOT1 (N11642, N11633);
and AND4 (N11643, N11628, N8387, N3264, N2366);
or OR4 (N11644, N11620, N1209, N5305, N9506);
and AND4 (N11645, N11643, N6095, N8378, N5608);
buf BUF1 (N11646, N11640);
xor XOR2 (N11647, N11636, N7076);
buf BUF1 (N11648, N11639);
and AND2 (N11649, N11644, N8782);
not NOT1 (N11650, N11646);
nor NOR4 (N11651, N11648, N6280, N7102, N3924);
nor NOR4 (N11652, N11642, N6219, N10980, N10800);
buf BUF1 (N11653, N11647);
nand NAND2 (N11654, N11634, N10561);
buf BUF1 (N11655, N11650);
xor XOR2 (N11656, N11649, N4229);
and AND2 (N11657, N11653, N4976);
buf BUF1 (N11658, N11626);
or OR3 (N11659, N11652, N6512, N10379);
nand NAND4 (N11660, N11657, N10311, N2126, N4482);
not NOT1 (N11661, N11660);
and AND3 (N11662, N11651, N550, N9227);
nor NOR3 (N11663, N11661, N7120, N4296);
not NOT1 (N11664, N11654);
nand NAND3 (N11665, N11664, N4492, N5568);
not NOT1 (N11666, N11645);
nor NOR4 (N11667, N11665, N7960, N4527, N905);
nand NAND4 (N11668, N11658, N982, N600, N9453);
not NOT1 (N11669, N11594);
xor XOR2 (N11670, N11656, N1487);
nor NOR4 (N11671, N11667, N439, N3861, N8543);
nand NAND2 (N11672, N11670, N2263);
buf BUF1 (N11673, N11659);
nor NOR4 (N11674, N11641, N5819, N3883, N5100);
nor NOR3 (N11675, N11666, N3027, N2720);
buf BUF1 (N11676, N11668);
xor XOR2 (N11677, N11655, N11663);
buf BUF1 (N11678, N1364);
or OR4 (N11679, N11673, N7494, N4768, N10584);
not NOT1 (N11680, N11674);
and AND3 (N11681, N11676, N2998, N7130);
xor XOR2 (N11682, N11680, N2044);
or OR3 (N11683, N11669, N6649, N7913);
xor XOR2 (N11684, N11679, N9048);
xor XOR2 (N11685, N11662, N4378);
not NOT1 (N11686, N11685);
nand NAND4 (N11687, N11678, N720, N3959, N2140);
buf BUF1 (N11688, N11683);
or OR2 (N11689, N11686, N4548);
xor XOR2 (N11690, N11682, N1512);
xor XOR2 (N11691, N11690, N5688);
and AND4 (N11692, N11677, N8498, N3896, N8404);
or OR4 (N11693, N11684, N9064, N3623, N5269);
nand NAND3 (N11694, N11675, N7307, N4018);
and AND4 (N11695, N11692, N10916, N7734, N6289);
nor NOR4 (N11696, N11688, N3295, N1358, N4665);
not NOT1 (N11697, N11695);
and AND2 (N11698, N11697, N9920);
buf BUF1 (N11699, N11696);
nor NOR3 (N11700, N11689, N805, N6602);
not NOT1 (N11701, N11687);
not NOT1 (N11702, N11700);
or OR3 (N11703, N11681, N6564, N2827);
or OR2 (N11704, N11698, N7996);
and AND2 (N11705, N11671, N10813);
not NOT1 (N11706, N11694);
xor XOR2 (N11707, N11693, N2582);
xor XOR2 (N11708, N11706, N8041);
not NOT1 (N11709, N11702);
and AND2 (N11710, N11672, N6642);
not NOT1 (N11711, N11709);
nor NOR4 (N11712, N11708, N5881, N11305, N802);
and AND3 (N11713, N11704, N8154, N5096);
nor NOR4 (N11714, N11712, N3291, N8563, N7364);
not NOT1 (N11715, N11699);
nand NAND3 (N11716, N11703, N1804, N4409);
not NOT1 (N11717, N11707);
nand NAND3 (N11718, N11715, N8146, N11288);
not NOT1 (N11719, N11710);
xor XOR2 (N11720, N11716, N2489);
xor XOR2 (N11721, N11718, N3258);
xor XOR2 (N11722, N11721, N5395);
nor NOR2 (N11723, N11713, N3198);
or OR2 (N11724, N11717, N2811);
or OR2 (N11725, N11724, N2081);
and AND4 (N11726, N11701, N2493, N3384, N1752);
or OR3 (N11727, N11705, N923, N6466);
xor XOR2 (N11728, N11722, N6703);
and AND4 (N11729, N11691, N1375, N6442, N3761);
nand NAND3 (N11730, N11726, N1012, N1341);
or OR3 (N11731, N11711, N7725, N4944);
buf BUF1 (N11732, N11725);
and AND3 (N11733, N11732, N677, N4405);
nor NOR2 (N11734, N11729, N3613);
nand NAND3 (N11735, N11731, N4185, N9811);
or OR2 (N11736, N11733, N2522);
and AND3 (N11737, N11728, N596, N9342);
buf BUF1 (N11738, N11735);
buf BUF1 (N11739, N11730);
not NOT1 (N11740, N11736);
xor XOR2 (N11741, N11739, N914);
xor XOR2 (N11742, N11737, N8131);
and AND3 (N11743, N11719, N8687, N10882);
not NOT1 (N11744, N11714);
xor XOR2 (N11745, N11727, N11588);
nand NAND4 (N11746, N11738, N8283, N7645, N3054);
and AND2 (N11747, N11720, N3572);
not NOT1 (N11748, N11740);
nand NAND3 (N11749, N11745, N1347, N6348);
nor NOR2 (N11750, N11741, N3055);
or OR4 (N11751, N11747, N1559, N8194, N1303);
or OR2 (N11752, N11734, N8041);
and AND2 (N11753, N11751, N6722);
nor NOR2 (N11754, N11748, N11680);
xor XOR2 (N11755, N11754, N6845);
nor NOR2 (N11756, N11746, N8396);
nor NOR2 (N11757, N11753, N9976);
buf BUF1 (N11758, N11756);
nor NOR4 (N11759, N11742, N42, N2255, N2626);
buf BUF1 (N11760, N11758);
nand NAND3 (N11761, N11723, N10174, N9159);
nor NOR2 (N11762, N11757, N10520);
buf BUF1 (N11763, N11744);
nor NOR3 (N11764, N11743, N10052, N9360);
and AND4 (N11765, N11750, N8999, N9778, N4613);
and AND3 (N11766, N11764, N7526, N512);
and AND2 (N11767, N11749, N2578);
not NOT1 (N11768, N11767);
xor XOR2 (N11769, N11768, N1253);
or OR2 (N11770, N11755, N5442);
xor XOR2 (N11771, N11769, N4061);
xor XOR2 (N11772, N11761, N9369);
and AND3 (N11773, N11752, N3667, N6415);
or OR3 (N11774, N11759, N489, N9000);
buf BUF1 (N11775, N11770);
not NOT1 (N11776, N11773);
xor XOR2 (N11777, N11775, N5228);
not NOT1 (N11778, N11763);
and AND3 (N11779, N11766, N6101, N2870);
buf BUF1 (N11780, N11771);
and AND4 (N11781, N11776, N3854, N7085, N5245);
nand NAND2 (N11782, N11774, N4094);
and AND4 (N11783, N11772, N120, N3389, N8575);
or OR3 (N11784, N11762, N8622, N11095);
nand NAND3 (N11785, N11783, N1620, N10096);
xor XOR2 (N11786, N11785, N6580);
not NOT1 (N11787, N11784);
and AND4 (N11788, N11777, N1978, N5648, N11128);
or OR3 (N11789, N11788, N8249, N6310);
xor XOR2 (N11790, N11782, N2947);
nor NOR2 (N11791, N11790, N269);
xor XOR2 (N11792, N11779, N7643);
nor NOR2 (N11793, N11791, N10983);
and AND4 (N11794, N11778, N10608, N7743, N3046);
not NOT1 (N11795, N11787);
and AND4 (N11796, N11760, N8007, N11385, N5900);
buf BUF1 (N11797, N11780);
xor XOR2 (N11798, N11781, N5850);
buf BUF1 (N11799, N11798);
and AND3 (N11800, N11797, N7333, N2313);
not NOT1 (N11801, N11765);
or OR3 (N11802, N11794, N7291, N9628);
xor XOR2 (N11803, N11801, N6604);
nand NAND2 (N11804, N11803, N1525);
nor NOR3 (N11805, N11804, N5516, N3952);
nor NOR2 (N11806, N11799, N5325);
not NOT1 (N11807, N11800);
nand NAND3 (N11808, N11789, N6334, N1105);
or OR4 (N11809, N11796, N845, N8918, N8537);
xor XOR2 (N11810, N11795, N7283);
nor NOR2 (N11811, N11786, N3271);
buf BUF1 (N11812, N11809);
nand NAND4 (N11813, N11808, N3477, N6917, N4484);
buf BUF1 (N11814, N11793);
or OR4 (N11815, N11805, N10051, N291, N7335);
nand NAND2 (N11816, N11815, N10052);
nand NAND2 (N11817, N11792, N8917);
nand NAND4 (N11818, N11813, N10691, N8881, N9141);
or OR3 (N11819, N11818, N3895, N5466);
nand NAND3 (N11820, N11810, N5303, N11322);
not NOT1 (N11821, N11819);
buf BUF1 (N11822, N11814);
xor XOR2 (N11823, N11802, N3282);
xor XOR2 (N11824, N11823, N218);
buf BUF1 (N11825, N11811);
xor XOR2 (N11826, N11816, N7248);
buf BUF1 (N11827, N11812);
or OR4 (N11828, N11822, N11133, N3319, N11393);
buf BUF1 (N11829, N11817);
not NOT1 (N11830, N11806);
not NOT1 (N11831, N11825);
and AND4 (N11832, N11807, N2996, N523, N10396);
nand NAND2 (N11833, N11832, N3243);
not NOT1 (N11834, N11830);
and AND2 (N11835, N11820, N9304);
not NOT1 (N11836, N11834);
buf BUF1 (N11837, N11831);
not NOT1 (N11838, N11828);
or OR4 (N11839, N11835, N2779, N7388, N9166);
and AND4 (N11840, N11833, N6225, N7503, N11806);
not NOT1 (N11841, N11821);
not NOT1 (N11842, N11841);
xor XOR2 (N11843, N11840, N10488);
nand NAND3 (N11844, N11824, N10712, N4544);
xor XOR2 (N11845, N11829, N273);
and AND3 (N11846, N11837, N675, N1945);
nor NOR3 (N11847, N11838, N1036, N1072);
and AND2 (N11848, N11836, N3873);
buf BUF1 (N11849, N11827);
xor XOR2 (N11850, N11845, N5075);
or OR3 (N11851, N11847, N11081, N106);
nand NAND4 (N11852, N11826, N4981, N5904, N9779);
buf BUF1 (N11853, N11843);
and AND3 (N11854, N11852, N1116, N4493);
xor XOR2 (N11855, N11851, N8703);
xor XOR2 (N11856, N11842, N3588);
nor NOR4 (N11857, N11855, N544, N6479, N10517);
not NOT1 (N11858, N11850);
not NOT1 (N11859, N11858);
buf BUF1 (N11860, N11857);
not NOT1 (N11861, N11860);
nor NOR3 (N11862, N11853, N5366, N4433);
or OR2 (N11863, N11861, N4348);
or OR2 (N11864, N11854, N9600);
or OR2 (N11865, N11863, N6295);
or OR3 (N11866, N11849, N8564, N11147);
and AND3 (N11867, N11846, N4210, N2027);
nand NAND4 (N11868, N11864, N11675, N5711, N11635);
nand NAND2 (N11869, N11839, N7038);
buf BUF1 (N11870, N11862);
xor XOR2 (N11871, N11848, N4610);
and AND3 (N11872, N11868, N8330, N416);
buf BUF1 (N11873, N11844);
xor XOR2 (N11874, N11865, N4845);
nand NAND2 (N11875, N11856, N4181);
not NOT1 (N11876, N11875);
not NOT1 (N11877, N11866);
not NOT1 (N11878, N11876);
or OR2 (N11879, N11867, N8000);
or OR4 (N11880, N11859, N6824, N3626, N4498);
not NOT1 (N11881, N11870);
buf BUF1 (N11882, N11871);
and AND2 (N11883, N11878, N4391);
not NOT1 (N11884, N11873);
nor NOR4 (N11885, N11872, N8866, N2986, N5473);
xor XOR2 (N11886, N11881, N6144);
xor XOR2 (N11887, N11879, N6369);
or OR2 (N11888, N11883, N4078);
buf BUF1 (N11889, N11869);
buf BUF1 (N11890, N11888);
and AND4 (N11891, N11874, N7553, N10425, N9710);
nor NOR4 (N11892, N11886, N4046, N4353, N2954);
xor XOR2 (N11893, N11889, N4723);
or OR3 (N11894, N11880, N2349, N6037);
not NOT1 (N11895, N11892);
nand NAND4 (N11896, N11885, N6101, N6366, N8882);
xor XOR2 (N11897, N11890, N1938);
xor XOR2 (N11898, N11882, N5430);
not NOT1 (N11899, N11895);
not NOT1 (N11900, N11898);
and AND4 (N11901, N11896, N11396, N2529, N8736);
buf BUF1 (N11902, N11884);
nand NAND2 (N11903, N11893, N8702);
nor NOR3 (N11904, N11902, N1844, N5387);
nand NAND3 (N11905, N11891, N7588, N7847);
and AND3 (N11906, N11887, N661, N7589);
and AND2 (N11907, N11899, N7349);
xor XOR2 (N11908, N11903, N1739);
xor XOR2 (N11909, N11897, N5192);
not NOT1 (N11910, N11877);
not NOT1 (N11911, N11907);
nand NAND4 (N11912, N11910, N3256, N11447, N9402);
xor XOR2 (N11913, N11911, N10927);
xor XOR2 (N11914, N11913, N3191);
and AND3 (N11915, N11914, N4870, N7272);
xor XOR2 (N11916, N11908, N3598);
xor XOR2 (N11917, N11900, N8701);
not NOT1 (N11918, N11915);
and AND3 (N11919, N11906, N6004, N4080);
buf BUF1 (N11920, N11916);
nand NAND3 (N11921, N11919, N5748, N3940);
and AND3 (N11922, N11917, N11066, N5937);
not NOT1 (N11923, N11920);
and AND4 (N11924, N11904, N3608, N9624, N8164);
buf BUF1 (N11925, N11912);
nor NOR2 (N11926, N11894, N4324);
buf BUF1 (N11927, N11924);
not NOT1 (N11928, N11918);
or OR3 (N11929, N11922, N3215, N11362);
xor XOR2 (N11930, N11909, N9928);
nand NAND3 (N11931, N11905, N9232, N5830);
xor XOR2 (N11932, N11926, N3975);
nor NOR3 (N11933, N11930, N6921, N9492);
and AND2 (N11934, N11925, N2194);
or OR4 (N11935, N11901, N9451, N2317, N1274);
and AND2 (N11936, N11927, N11641);
nand NAND2 (N11937, N11936, N11735);
and AND4 (N11938, N11937, N2205, N7455, N1023);
or OR4 (N11939, N11938, N3984, N5466, N1819);
nand NAND4 (N11940, N11935, N617, N9413, N10076);
and AND3 (N11941, N11928, N7760, N5095);
xor XOR2 (N11942, N11939, N10811);
buf BUF1 (N11943, N11931);
and AND3 (N11944, N11940, N6130, N7529);
buf BUF1 (N11945, N11941);
and AND2 (N11946, N11921, N11285);
not NOT1 (N11947, N11933);
nor NOR4 (N11948, N11944, N4375, N11248, N6075);
buf BUF1 (N11949, N11932);
nand NAND4 (N11950, N11947, N3440, N11791, N5305);
and AND2 (N11951, N11923, N10626);
xor XOR2 (N11952, N11945, N4869);
xor XOR2 (N11953, N11950, N11133);
xor XOR2 (N11954, N11953, N1086);
xor XOR2 (N11955, N11942, N4995);
nand NAND3 (N11956, N11952, N11107, N979);
buf BUF1 (N11957, N11946);
nor NOR2 (N11958, N11956, N3016);
nand NAND4 (N11959, N11957, N616, N4846, N3954);
xor XOR2 (N11960, N11934, N5627);
or OR3 (N11961, N11949, N8806, N7894);
and AND4 (N11962, N11951, N7416, N10101, N369);
nand NAND2 (N11963, N11943, N993);
nand NAND2 (N11964, N11963, N4626);
nand NAND3 (N11965, N11959, N4773, N3625);
nor NOR3 (N11966, N11961, N186, N10290);
nand NAND4 (N11967, N11955, N11831, N4558, N9645);
not NOT1 (N11968, N11966);
not NOT1 (N11969, N11948);
and AND3 (N11970, N11968, N10117, N2877);
not NOT1 (N11971, N11954);
not NOT1 (N11972, N11969);
or OR3 (N11973, N11967, N1602, N1369);
or OR4 (N11974, N11964, N8247, N9449, N6161);
buf BUF1 (N11975, N11973);
xor XOR2 (N11976, N11958, N8800);
buf BUF1 (N11977, N11971);
nor NOR3 (N11978, N11962, N10414, N2221);
and AND4 (N11979, N11960, N1155, N9022, N8422);
xor XOR2 (N11980, N11976, N10648);
or OR3 (N11981, N11965, N6974, N4867);
nor NOR2 (N11982, N11972, N11221);
and AND2 (N11983, N11929, N8872);
or OR4 (N11984, N11975, N4084, N1944, N11101);
xor XOR2 (N11985, N11970, N1379);
nor NOR3 (N11986, N11983, N8699, N1176);
not NOT1 (N11987, N11979);
and AND3 (N11988, N11985, N839, N4903);
not NOT1 (N11989, N11987);
and AND3 (N11990, N11986, N1244, N9687);
nand NAND2 (N11991, N11981, N10896);
not NOT1 (N11992, N11977);
xor XOR2 (N11993, N11974, N8187);
or OR4 (N11994, N11993, N9618, N4984, N9946);
or OR3 (N11995, N11984, N10481, N6203);
xor XOR2 (N11996, N11988, N1072);
nand NAND3 (N11997, N11978, N11136, N8011);
not NOT1 (N11998, N11990);
nor NOR3 (N11999, N11997, N5374, N3538);
nand NAND2 (N12000, N11994, N9215);
nor NOR3 (N12001, N11992, N5316, N4739);
not NOT1 (N12002, N11995);
not NOT1 (N12003, N12001);
xor XOR2 (N12004, N11991, N8837);
xor XOR2 (N12005, N12003, N2424);
and AND2 (N12006, N11998, N7392);
not NOT1 (N12007, N11996);
and AND2 (N12008, N12002, N1779);
and AND4 (N12009, N11980, N3091, N10564, N1093);
or OR4 (N12010, N12008, N5072, N4118, N315);
not NOT1 (N12011, N11982);
not NOT1 (N12012, N12000);
or OR2 (N12013, N11999, N7700);
buf BUF1 (N12014, N12005);
buf BUF1 (N12015, N12014);
and AND4 (N12016, N12004, N7535, N611, N727);
or OR4 (N12017, N12010, N11894, N2650, N3630);
not NOT1 (N12018, N12013);
buf BUF1 (N12019, N11989);
buf BUF1 (N12020, N12012);
nor NOR3 (N12021, N12007, N10168, N11363);
not NOT1 (N12022, N12021);
and AND3 (N12023, N12018, N873, N3606);
nor NOR2 (N12024, N12023, N9324);
or OR2 (N12025, N12020, N3140);
and AND2 (N12026, N12022, N5478);
xor XOR2 (N12027, N12024, N6186);
or OR2 (N12028, N12026, N7480);
buf BUF1 (N12029, N12011);
nor NOR3 (N12030, N12009, N4340, N7443);
not NOT1 (N12031, N12029);
and AND3 (N12032, N12025, N9548, N11612);
buf BUF1 (N12033, N12032);
nand NAND3 (N12034, N12006, N10596, N1450);
buf BUF1 (N12035, N12015);
or OR2 (N12036, N12027, N542);
not NOT1 (N12037, N12017);
nand NAND4 (N12038, N12037, N1882, N11350, N7130);
xor XOR2 (N12039, N12035, N11622);
and AND3 (N12040, N12034, N2052, N10277);
buf BUF1 (N12041, N12016);
xor XOR2 (N12042, N12038, N9453);
not NOT1 (N12043, N12039);
nor NOR3 (N12044, N12040, N8969, N3114);
and AND3 (N12045, N12043, N7412, N7704);
or OR2 (N12046, N12030, N5177);
xor XOR2 (N12047, N12042, N4036);
or OR3 (N12048, N12046, N7094, N7904);
and AND4 (N12049, N12041, N6565, N8588, N7591);
and AND2 (N12050, N12048, N8087);
nor NOR4 (N12051, N12019, N9506, N1355, N3073);
nand NAND2 (N12052, N12033, N9941);
not NOT1 (N12053, N12044);
xor XOR2 (N12054, N12051, N4076);
buf BUF1 (N12055, N12028);
not NOT1 (N12056, N12036);
or OR3 (N12057, N12050, N9219, N7459);
not NOT1 (N12058, N12054);
nand NAND4 (N12059, N12058, N1744, N6307, N4071);
nand NAND2 (N12060, N12047, N11753);
buf BUF1 (N12061, N12031);
not NOT1 (N12062, N12052);
not NOT1 (N12063, N12045);
nor NOR4 (N12064, N12053, N1375, N2771, N8106);
and AND3 (N12065, N12063, N10294, N10419);
nor NOR3 (N12066, N12060, N1253, N5347);
nand NAND4 (N12067, N12055, N10218, N2372, N357);
nand NAND2 (N12068, N12062, N11989);
and AND2 (N12069, N12065, N9567);
xor XOR2 (N12070, N12057, N494);
and AND3 (N12071, N12061, N11112, N9229);
nor NOR2 (N12072, N12070, N1880);
xor XOR2 (N12073, N12072, N8943);
xor XOR2 (N12074, N12067, N10887);
buf BUF1 (N12075, N12069);
xor XOR2 (N12076, N12056, N9211);
not NOT1 (N12077, N12068);
buf BUF1 (N12078, N12071);
and AND4 (N12079, N12049, N8827, N9608, N1775);
not NOT1 (N12080, N12064);
nor NOR2 (N12081, N12076, N11402);
buf BUF1 (N12082, N12079);
or OR4 (N12083, N12073, N5939, N1785, N4879);
xor XOR2 (N12084, N12078, N8261);
xor XOR2 (N12085, N12082, N4237);
nand NAND3 (N12086, N12066, N11460, N5988);
xor XOR2 (N12087, N12059, N10648);
not NOT1 (N12088, N12085);
buf BUF1 (N12089, N12084);
buf BUF1 (N12090, N12077);
or OR3 (N12091, N12088, N2303, N9715);
buf BUF1 (N12092, N12089);
xor XOR2 (N12093, N12087, N10384);
nor NOR4 (N12094, N12091, N5706, N4387, N751);
nor NOR4 (N12095, N12081, N10558, N2726, N789);
and AND4 (N12096, N12074, N3229, N9241, N149);
nor NOR4 (N12097, N12094, N10049, N5453, N5936);
or OR4 (N12098, N12080, N1315, N611, N2635);
nor NOR2 (N12099, N12097, N6524);
buf BUF1 (N12100, N12098);
or OR2 (N12101, N12083, N1289);
xor XOR2 (N12102, N12101, N1390);
xor XOR2 (N12103, N12092, N9447);
not NOT1 (N12104, N12102);
nor NOR2 (N12105, N12086, N4802);
xor XOR2 (N12106, N12090, N2767);
nand NAND2 (N12107, N12103, N642);
nand NAND2 (N12108, N12107, N2215);
not NOT1 (N12109, N12075);
nand NAND3 (N12110, N12108, N234, N9427);
nor NOR4 (N12111, N12100, N1412, N9603, N3825);
nor NOR4 (N12112, N12105, N3647, N5117, N7900);
not NOT1 (N12113, N12106);
nand NAND2 (N12114, N12109, N10783);
buf BUF1 (N12115, N12111);
not NOT1 (N12116, N12099);
and AND4 (N12117, N12095, N8744, N11808, N12088);
and AND2 (N12118, N12113, N4393);
not NOT1 (N12119, N12116);
nand NAND2 (N12120, N12093, N9820);
nand NAND2 (N12121, N12114, N564);
or OR4 (N12122, N12096, N7230, N8508, N5071);
buf BUF1 (N12123, N12119);
not NOT1 (N12124, N12112);
or OR4 (N12125, N12120, N4649, N478, N6789);
nand NAND3 (N12126, N12118, N3875, N3282);
not NOT1 (N12127, N12126);
and AND4 (N12128, N12104, N9198, N10723, N3588);
xor XOR2 (N12129, N12124, N10650);
not NOT1 (N12130, N12125);
xor XOR2 (N12131, N12121, N5417);
not NOT1 (N12132, N12115);
nand NAND2 (N12133, N12117, N10865);
xor XOR2 (N12134, N12122, N9155);
and AND4 (N12135, N12128, N11746, N7083, N11242);
and AND2 (N12136, N12131, N6177);
xor XOR2 (N12137, N12132, N6489);
nand NAND4 (N12138, N12136, N8009, N6533, N10570);
and AND3 (N12139, N12123, N11853, N7681);
nand NAND4 (N12140, N12138, N5215, N2980, N6683);
nor NOR2 (N12141, N12129, N5992);
nor NOR4 (N12142, N12130, N6177, N1127, N4941);
and AND3 (N12143, N12142, N5299, N2216);
nor NOR4 (N12144, N12139, N6103, N3081, N8551);
or OR3 (N12145, N12110, N6312, N6621);
buf BUF1 (N12146, N12137);
nand NAND3 (N12147, N12144, N1438, N11068);
nand NAND2 (N12148, N12134, N5804);
buf BUF1 (N12149, N12127);
and AND3 (N12150, N12147, N10943, N3831);
buf BUF1 (N12151, N12146);
or OR4 (N12152, N12141, N9242, N9452, N8393);
nand NAND2 (N12153, N12151, N1875);
not NOT1 (N12154, N12148);
buf BUF1 (N12155, N12135);
and AND2 (N12156, N12143, N9200);
buf BUF1 (N12157, N12153);
xor XOR2 (N12158, N12155, N1590);
or OR3 (N12159, N12149, N10981, N790);
nand NAND3 (N12160, N12150, N8828, N117);
and AND2 (N12161, N12158, N161);
or OR2 (N12162, N12152, N11685);
or OR4 (N12163, N12160, N367, N2846, N987);
and AND3 (N12164, N12161, N10869, N6326);
nor NOR3 (N12165, N12145, N2227, N6125);
nor NOR2 (N12166, N12163, N1026);
and AND2 (N12167, N12166, N11296);
and AND3 (N12168, N12133, N1547, N467);
nand NAND4 (N12169, N12167, N6231, N6598, N2253);
or OR2 (N12170, N12165, N3710);
buf BUF1 (N12171, N12156);
nand NAND2 (N12172, N12168, N2203);
xor XOR2 (N12173, N12172, N7243);
nor NOR4 (N12174, N12154, N8338, N2733, N3033);
nand NAND3 (N12175, N12159, N2298, N6389);
nor NOR4 (N12176, N12171, N7054, N9680, N1649);
nor NOR2 (N12177, N12162, N3076);
and AND3 (N12178, N12169, N2033, N10641);
nand NAND2 (N12179, N12164, N11471);
and AND2 (N12180, N12176, N10868);
nand NAND3 (N12181, N12175, N9032, N58);
nand NAND2 (N12182, N12179, N9247);
xor XOR2 (N12183, N12174, N4637);
xor XOR2 (N12184, N12181, N11388);
not NOT1 (N12185, N12182);
and AND3 (N12186, N12184, N8327, N4680);
xor XOR2 (N12187, N12140, N6439);
nor NOR4 (N12188, N12187, N4937, N4253, N8404);
nor NOR4 (N12189, N12170, N6404, N4456, N3395);
and AND3 (N12190, N12183, N2244, N3561);
nor NOR3 (N12191, N12180, N7427, N640);
nor NOR2 (N12192, N12173, N3079);
nand NAND4 (N12193, N12177, N7525, N8266, N8509);
xor XOR2 (N12194, N12191, N1636);
or OR4 (N12195, N12189, N4031, N4321, N3855);
or OR2 (N12196, N12190, N7857);
and AND2 (N12197, N12186, N7143);
not NOT1 (N12198, N12192);
nor NOR4 (N12199, N12178, N3761, N11921, N2757);
not NOT1 (N12200, N12193);
or OR2 (N12201, N12199, N6712);
buf BUF1 (N12202, N12185);
nor NOR3 (N12203, N12157, N4047, N6146);
nor NOR2 (N12204, N12203, N11182);
or OR2 (N12205, N12197, N6427);
nor NOR4 (N12206, N12196, N4067, N3476, N3152);
and AND4 (N12207, N12201, N11720, N4664, N2216);
not NOT1 (N12208, N12206);
and AND2 (N12209, N12204, N11266);
and AND4 (N12210, N12198, N1091, N4908, N11746);
or OR4 (N12211, N12188, N7769, N7673, N7620);
and AND3 (N12212, N12210, N1537, N3203);
and AND3 (N12213, N12207, N8584, N10280);
and AND3 (N12214, N12211, N6579, N2190);
and AND2 (N12215, N12214, N2525);
nor NOR2 (N12216, N12215, N10678);
or OR4 (N12217, N12213, N3260, N4450, N7292);
nor NOR3 (N12218, N12205, N6758, N7818);
not NOT1 (N12219, N12208);
nor NOR4 (N12220, N12216, N2989, N12001, N5272);
not NOT1 (N12221, N12194);
and AND3 (N12222, N12202, N9628, N8512);
nor NOR3 (N12223, N12200, N2361, N4053);
buf BUF1 (N12224, N12220);
not NOT1 (N12225, N12219);
xor XOR2 (N12226, N12224, N1252);
not NOT1 (N12227, N12209);
and AND3 (N12228, N12212, N10145, N3150);
nand NAND3 (N12229, N12217, N4242, N10243);
not NOT1 (N12230, N12218);
buf BUF1 (N12231, N12221);
nor NOR2 (N12232, N12195, N837);
nor NOR2 (N12233, N12231, N6250);
and AND4 (N12234, N12233, N4483, N8240, N948);
not NOT1 (N12235, N12227);
xor XOR2 (N12236, N12226, N5258);
nand NAND2 (N12237, N12229, N6265);
xor XOR2 (N12238, N12232, N7931);
not NOT1 (N12239, N12225);
xor XOR2 (N12240, N12237, N2395);
nor NOR3 (N12241, N12222, N1685, N6258);
and AND4 (N12242, N12235, N3657, N9632, N8046);
nand NAND2 (N12243, N12234, N849);
buf BUF1 (N12244, N12223);
nor NOR3 (N12245, N12238, N2377, N4457);
xor XOR2 (N12246, N12228, N9825);
or OR3 (N12247, N12236, N11791, N10730);
buf BUF1 (N12248, N12246);
nor NOR2 (N12249, N12241, N4317);
xor XOR2 (N12250, N12239, N11232);
or OR2 (N12251, N12230, N4782);
not NOT1 (N12252, N12251);
and AND3 (N12253, N12244, N2981, N1523);
and AND2 (N12254, N12252, N5408);
or OR2 (N12255, N12242, N4244);
nand NAND2 (N12256, N12250, N3004);
xor XOR2 (N12257, N12253, N7925);
xor XOR2 (N12258, N12257, N11832);
buf BUF1 (N12259, N12258);
not NOT1 (N12260, N12245);
nand NAND2 (N12261, N12254, N5671);
not NOT1 (N12262, N12255);
not NOT1 (N12263, N12243);
nand NAND3 (N12264, N12263, N8779, N3454);
nor NOR3 (N12265, N12261, N11906, N11501);
nor NOR4 (N12266, N12240, N4628, N2661, N7660);
xor XOR2 (N12267, N12249, N5530);
nand NAND2 (N12268, N12259, N3708);
buf BUF1 (N12269, N12260);
not NOT1 (N12270, N12266);
nand NAND2 (N12271, N12256, N1952);
xor XOR2 (N12272, N12269, N1970);
nand NAND4 (N12273, N12262, N9667, N2721, N7453);
not NOT1 (N12274, N12272);
not NOT1 (N12275, N12248);
and AND4 (N12276, N12265, N814, N5718, N2910);
buf BUF1 (N12277, N12275);
nand NAND2 (N12278, N12267, N3825);
nor NOR3 (N12279, N12271, N10006, N8012);
not NOT1 (N12280, N12268);
or OR4 (N12281, N12277, N4143, N6205, N11652);
buf BUF1 (N12282, N12247);
and AND3 (N12283, N12276, N1510, N6644);
nor NOR4 (N12284, N12264, N9479, N7544, N1551);
nand NAND3 (N12285, N12280, N3517, N3063);
nand NAND3 (N12286, N12273, N2480, N4143);
not NOT1 (N12287, N12282);
nor NOR2 (N12288, N12285, N3472);
not NOT1 (N12289, N12288);
not NOT1 (N12290, N12289);
and AND2 (N12291, N12274, N11598);
or OR2 (N12292, N12283, N5663);
or OR2 (N12293, N12291, N1507);
nand NAND2 (N12294, N12284, N3899);
xor XOR2 (N12295, N12279, N1868);
or OR2 (N12296, N12292, N395);
not NOT1 (N12297, N12278);
buf BUF1 (N12298, N12281);
not NOT1 (N12299, N12294);
or OR2 (N12300, N12286, N5344);
buf BUF1 (N12301, N12290);
nand NAND4 (N12302, N12298, N7384, N9592, N8785);
nor NOR4 (N12303, N12302, N9359, N10831, N2051);
xor XOR2 (N12304, N12270, N10322);
nor NOR2 (N12305, N12299, N5528);
or OR2 (N12306, N12304, N507);
nor NOR2 (N12307, N12303, N776);
not NOT1 (N12308, N12296);
nand NAND4 (N12309, N12308, N11060, N3823, N5459);
not NOT1 (N12310, N12295);
and AND4 (N12311, N12287, N11654, N6992, N10645);
and AND4 (N12312, N12293, N767, N9213, N7519);
xor XOR2 (N12313, N12307, N1958);
buf BUF1 (N12314, N12301);
or OR3 (N12315, N12312, N6664, N11605);
xor XOR2 (N12316, N12311, N5147);
or OR4 (N12317, N12305, N9018, N8723, N11805);
nor NOR3 (N12318, N12300, N10634, N7558);
and AND2 (N12319, N12317, N11689);
buf BUF1 (N12320, N12318);
and AND3 (N12321, N12313, N1723, N12293);
buf BUF1 (N12322, N12297);
and AND3 (N12323, N12314, N10289, N551);
and AND3 (N12324, N12315, N526, N11197);
nor NOR4 (N12325, N12310, N180, N3758, N103);
xor XOR2 (N12326, N12322, N3947);
and AND3 (N12327, N12316, N7986, N10970);
buf BUF1 (N12328, N12326);
and AND4 (N12329, N12323, N4127, N7573, N4098);
and AND2 (N12330, N12325, N3223);
nor NOR4 (N12331, N12320, N3278, N5804, N3373);
buf BUF1 (N12332, N12319);
nor NOR2 (N12333, N12306, N2833);
not NOT1 (N12334, N12329);
nand NAND2 (N12335, N12321, N9136);
buf BUF1 (N12336, N12333);
and AND3 (N12337, N12336, N7442, N1697);
not NOT1 (N12338, N12330);
nand NAND4 (N12339, N12324, N6975, N8052, N6329);
or OR2 (N12340, N12334, N11041);
not NOT1 (N12341, N12338);
buf BUF1 (N12342, N12327);
xor XOR2 (N12343, N12342, N3244);
not NOT1 (N12344, N12332);
buf BUF1 (N12345, N12328);
nor NOR3 (N12346, N12344, N8270, N9989);
or OR3 (N12347, N12346, N8129, N8137);
nor NOR4 (N12348, N12341, N10451, N7558, N10576);
and AND2 (N12349, N12340, N4079);
nand NAND2 (N12350, N12339, N11430);
nor NOR3 (N12351, N12343, N10293, N5440);
not NOT1 (N12352, N12337);
nor NOR4 (N12353, N12350, N11508, N5456, N1089);
nand NAND3 (N12354, N12352, N12274, N2456);
buf BUF1 (N12355, N12331);
and AND3 (N12356, N12355, N10607, N3770);
nand NAND4 (N12357, N12351, N8681, N6862, N11743);
nor NOR4 (N12358, N12349, N357, N5061, N9196);
nor NOR3 (N12359, N12335, N11170, N7398);
nand NAND3 (N12360, N12309, N8629, N9430);
or OR3 (N12361, N12353, N7568, N10359);
nand NAND2 (N12362, N12348, N5340);
or OR2 (N12363, N12361, N10649);
nor NOR3 (N12364, N12359, N7976, N3895);
not NOT1 (N12365, N12360);
xor XOR2 (N12366, N12362, N5383);
xor XOR2 (N12367, N12366, N1902);
buf BUF1 (N12368, N12358);
nand NAND4 (N12369, N12368, N4248, N732, N8540);
or OR3 (N12370, N12363, N10797, N5170);
xor XOR2 (N12371, N12367, N4476);
or OR4 (N12372, N12365, N8936, N8097, N4561);
or OR3 (N12373, N12372, N11702, N2675);
xor XOR2 (N12374, N12371, N4422);
or OR2 (N12375, N12347, N1839);
not NOT1 (N12376, N12373);
nand NAND2 (N12377, N12354, N9031);
nand NAND3 (N12378, N12345, N9346, N6691);
nand NAND3 (N12379, N12377, N3326, N9915);
not NOT1 (N12380, N12374);
and AND2 (N12381, N12379, N8251);
buf BUF1 (N12382, N12370);
xor XOR2 (N12383, N12375, N2450);
and AND2 (N12384, N12380, N5383);
xor XOR2 (N12385, N12364, N484);
and AND4 (N12386, N12357, N5421, N8253, N1515);
or OR2 (N12387, N12378, N7377);
nand NAND2 (N12388, N12356, N10448);
xor XOR2 (N12389, N12376, N976);
not NOT1 (N12390, N12383);
buf BUF1 (N12391, N12385);
nand NAND4 (N12392, N12389, N1107, N5007, N8387);
and AND3 (N12393, N12390, N11083, N1852);
xor XOR2 (N12394, N12393, N7475);
xor XOR2 (N12395, N12381, N8751);
not NOT1 (N12396, N12384);
or OR2 (N12397, N12396, N12151);
buf BUF1 (N12398, N12382);
and AND4 (N12399, N12394, N5911, N11069, N10529);
nand NAND4 (N12400, N12388, N105, N4826, N10201);
xor XOR2 (N12401, N12398, N7734);
nor NOR2 (N12402, N12399, N1298);
or OR2 (N12403, N12369, N7580);
and AND3 (N12404, N12392, N2633, N7117);
not NOT1 (N12405, N12404);
nor NOR3 (N12406, N12391, N7745, N12334);
not NOT1 (N12407, N12403);
xor XOR2 (N12408, N12407, N3802);
not NOT1 (N12409, N12406);
xor XOR2 (N12410, N12401, N5211);
or OR3 (N12411, N12402, N1017, N8372);
nor NOR2 (N12412, N12387, N500);
or OR3 (N12413, N12410, N10805, N3693);
nand NAND2 (N12414, N12409, N9061);
nand NAND3 (N12415, N12397, N5296, N3232);
xor XOR2 (N12416, N12400, N9281);
or OR4 (N12417, N12386, N3491, N7421, N2972);
buf BUF1 (N12418, N12412);
nor NOR2 (N12419, N12411, N3459);
nand NAND3 (N12420, N12416, N2334, N5636);
and AND4 (N12421, N12415, N3729, N1599, N10256);
nand NAND2 (N12422, N12421, N8593);
buf BUF1 (N12423, N12395);
and AND4 (N12424, N12414, N8106, N4888, N4699);
buf BUF1 (N12425, N12419);
and AND3 (N12426, N12405, N9751, N11822);
nor NOR2 (N12427, N12425, N7503);
xor XOR2 (N12428, N12427, N1912);
and AND3 (N12429, N12422, N7370, N10181);
and AND3 (N12430, N12420, N9670, N10903);
not NOT1 (N12431, N12429);
or OR3 (N12432, N12417, N5019, N6404);
and AND4 (N12433, N12430, N8849, N287, N1607);
nand NAND2 (N12434, N12431, N391);
nor NOR4 (N12435, N12413, N8158, N4442, N5056);
xor XOR2 (N12436, N12408, N10774);
not NOT1 (N12437, N12434);
nor NOR4 (N12438, N12418, N7592, N5275, N5392);
buf BUF1 (N12439, N12433);
nor NOR4 (N12440, N12432, N7687, N9099, N4199);
or OR3 (N12441, N12426, N8349, N7730);
not NOT1 (N12442, N12424);
not NOT1 (N12443, N12435);
or OR2 (N12444, N12428, N5117);
not NOT1 (N12445, N12441);
nand NAND3 (N12446, N12440, N8947, N8408);
nand NAND2 (N12447, N12444, N380);
nor NOR3 (N12448, N12437, N12137, N10610);
xor XOR2 (N12449, N12442, N8930);
nand NAND4 (N12450, N12446, N3833, N1001, N8081);
nand NAND2 (N12451, N12443, N10179);
and AND2 (N12452, N12450, N11262);
and AND3 (N12453, N12436, N4713, N1651);
not NOT1 (N12454, N12445);
or OR3 (N12455, N12438, N6536, N9673);
and AND4 (N12456, N12452, N5767, N9038, N11128);
buf BUF1 (N12457, N12455);
nand NAND2 (N12458, N12451, N1432);
not NOT1 (N12459, N12453);
nand NAND2 (N12460, N12454, N11046);
nor NOR3 (N12461, N12423, N4196, N7813);
or OR3 (N12462, N12458, N3359, N8759);
or OR4 (N12463, N12461, N4467, N10540, N6906);
not NOT1 (N12464, N12463);
not NOT1 (N12465, N12448);
nor NOR4 (N12466, N12459, N9775, N1956, N6805);
nor NOR2 (N12467, N12462, N3885);
nand NAND3 (N12468, N12467, N11428, N5783);
nand NAND3 (N12469, N12460, N1256, N6541);
or OR3 (N12470, N12457, N10707, N7361);
and AND2 (N12471, N12449, N6190);
and AND2 (N12472, N12468, N419);
or OR2 (N12473, N12472, N3364);
nor NOR4 (N12474, N12471, N9579, N7050, N1131);
or OR2 (N12475, N12464, N1159);
and AND2 (N12476, N12473, N6439);
and AND3 (N12477, N12456, N7843, N5779);
nand NAND2 (N12478, N12470, N1734);
and AND3 (N12479, N12477, N955, N3028);
or OR2 (N12480, N12447, N8142);
buf BUF1 (N12481, N12465);
nor NOR3 (N12482, N12474, N269, N1579);
xor XOR2 (N12483, N12482, N1256);
xor XOR2 (N12484, N12483, N8492);
nor NOR3 (N12485, N12484, N5282, N8780);
xor XOR2 (N12486, N12475, N5155);
not NOT1 (N12487, N12480);
buf BUF1 (N12488, N12466);
nand NAND3 (N12489, N12439, N1918, N681);
or OR2 (N12490, N12485, N3303);
nor NOR3 (N12491, N12469, N10565, N2204);
nand NAND4 (N12492, N12490, N7322, N2794, N2030);
or OR2 (N12493, N12492, N11964);
or OR4 (N12494, N12476, N9254, N6807, N6857);
and AND4 (N12495, N12479, N882, N4017, N1592);
not NOT1 (N12496, N12478);
or OR3 (N12497, N12486, N1502, N31);
not NOT1 (N12498, N12481);
buf BUF1 (N12499, N12491);
nor NOR3 (N12500, N12499, N1552, N6790);
or OR4 (N12501, N12493, N3957, N2479, N3581);
and AND4 (N12502, N12495, N7056, N3815, N11695);
nand NAND4 (N12503, N12496, N788, N7404, N644);
buf BUF1 (N12504, N12487);
or OR3 (N12505, N12488, N497, N2269);
nand NAND3 (N12506, N12498, N7647, N9048);
not NOT1 (N12507, N12504);
not NOT1 (N12508, N12494);
nand NAND2 (N12509, N12507, N5446);
or OR4 (N12510, N12500, N10526, N10952, N6930);
nor NOR3 (N12511, N12501, N10170, N6694);
buf BUF1 (N12512, N12505);
not NOT1 (N12513, N12509);
nand NAND2 (N12514, N12503, N4983);
or OR4 (N12515, N12512, N2168, N5641, N2908);
nor NOR2 (N12516, N12508, N6708);
nor NOR3 (N12517, N12489, N2445, N10651);
nor NOR4 (N12518, N12514, N7837, N7633, N5967);
nor NOR2 (N12519, N12515, N9670);
not NOT1 (N12520, N12497);
or OR2 (N12521, N12510, N9115);
buf BUF1 (N12522, N12517);
nand NAND3 (N12523, N12511, N2857, N71);
and AND4 (N12524, N12516, N6828, N9300, N3490);
and AND2 (N12525, N12502, N2959);
and AND2 (N12526, N12506, N2279);
nor NOR2 (N12527, N12521, N2210);
and AND4 (N12528, N12522, N2835, N5736, N3970);
not NOT1 (N12529, N12527);
nor NOR3 (N12530, N12526, N11174, N2084);
not NOT1 (N12531, N12524);
not NOT1 (N12532, N12523);
buf BUF1 (N12533, N12532);
nand NAND3 (N12534, N12513, N6391, N9302);
xor XOR2 (N12535, N12519, N6949);
nand NAND2 (N12536, N12518, N4020);
nand NAND2 (N12537, N12520, N2368);
nand NAND2 (N12538, N12529, N1928);
buf BUF1 (N12539, N12535);
nor NOR4 (N12540, N12531, N2136, N8689, N11001);
nor NOR2 (N12541, N12533, N12266);
not NOT1 (N12542, N12538);
and AND2 (N12543, N12534, N8710);
nand NAND3 (N12544, N12525, N5387, N12078);
nand NAND4 (N12545, N12537, N6446, N5045, N9401);
xor XOR2 (N12546, N12530, N6269);
or OR2 (N12547, N12539, N4081);
not NOT1 (N12548, N12543);
xor XOR2 (N12549, N12548, N9615);
or OR2 (N12550, N12546, N9457);
nand NAND2 (N12551, N12544, N10662);
buf BUF1 (N12552, N12540);
nand NAND3 (N12553, N12547, N9202, N8776);
nor NOR4 (N12554, N12528, N11832, N10680, N7573);
buf BUF1 (N12555, N12551);
and AND4 (N12556, N12550, N11788, N11337, N7477);
or OR2 (N12557, N12552, N6290);
nor NOR2 (N12558, N12556, N3243);
or OR3 (N12559, N12558, N1634, N2402);
nand NAND4 (N12560, N12536, N3056, N71, N3841);
buf BUF1 (N12561, N12560);
xor XOR2 (N12562, N12559, N10875);
nor NOR4 (N12563, N12561, N2135, N4181, N11318);
xor XOR2 (N12564, N12562, N8911);
xor XOR2 (N12565, N12564, N751);
buf BUF1 (N12566, N12557);
not NOT1 (N12567, N12542);
buf BUF1 (N12568, N12565);
nor NOR3 (N12569, N12549, N9366, N4805);
buf BUF1 (N12570, N12566);
xor XOR2 (N12571, N12567, N2301);
xor XOR2 (N12572, N12554, N9291);
buf BUF1 (N12573, N12569);
not NOT1 (N12574, N12541);
nand NAND3 (N12575, N12555, N221, N1637);
not NOT1 (N12576, N12572);
buf BUF1 (N12577, N12568);
or OR4 (N12578, N12553, N508, N4482, N2527);
or OR4 (N12579, N12573, N4212, N9652, N2921);
nor NOR3 (N12580, N12563, N7817, N4980);
and AND3 (N12581, N12578, N2331, N11633);
xor XOR2 (N12582, N12577, N9513);
buf BUF1 (N12583, N12576);
xor XOR2 (N12584, N12570, N1268);
and AND4 (N12585, N12584, N2037, N11705, N11013);
or OR3 (N12586, N12545, N2278, N2258);
buf BUF1 (N12587, N12583);
and AND4 (N12588, N12575, N4517, N8340, N1347);
buf BUF1 (N12589, N12579);
buf BUF1 (N12590, N12574);
and AND4 (N12591, N12586, N3837, N9518, N3577);
buf BUF1 (N12592, N12587);
nor NOR2 (N12593, N12592, N4236);
nor NOR2 (N12594, N12589, N8320);
nor NOR4 (N12595, N12594, N10217, N533, N5132);
or OR3 (N12596, N12595, N12511, N6195);
and AND3 (N12597, N12585, N4930, N750);
or OR4 (N12598, N12581, N9007, N7230, N5105);
or OR2 (N12599, N12591, N6106);
or OR3 (N12600, N12582, N8386, N2538);
nor NOR2 (N12601, N12588, N1051);
buf BUF1 (N12602, N12598);
not NOT1 (N12603, N12580);
nand NAND3 (N12604, N12602, N2338, N10974);
buf BUF1 (N12605, N12571);
xor XOR2 (N12606, N12600, N7356);
xor XOR2 (N12607, N12599, N3209);
buf BUF1 (N12608, N12605);
and AND2 (N12609, N12603, N2334);
nor NOR2 (N12610, N12596, N5296);
nand NAND3 (N12611, N12597, N3625, N10818);
nand NAND3 (N12612, N12601, N1180, N305);
buf BUF1 (N12613, N12607);
and AND2 (N12614, N12608, N8152);
xor XOR2 (N12615, N12593, N9647);
xor XOR2 (N12616, N12614, N991);
nor NOR2 (N12617, N12616, N8660);
not NOT1 (N12618, N12613);
buf BUF1 (N12619, N12604);
nor NOR2 (N12620, N12611, N9154);
nand NAND3 (N12621, N12609, N9765, N12583);
nor NOR4 (N12622, N12612, N12569, N12377, N3675);
and AND2 (N12623, N12621, N6969);
not NOT1 (N12624, N12590);
and AND4 (N12625, N12606, N12587, N2247, N185);
not NOT1 (N12626, N12617);
nor NOR2 (N12627, N12623, N11914);
nand NAND3 (N12628, N12627, N6958, N7003);
or OR3 (N12629, N12628, N4656, N3399);
buf BUF1 (N12630, N12624);
not NOT1 (N12631, N12615);
nand NAND3 (N12632, N12618, N6446, N5683);
buf BUF1 (N12633, N12619);
nand NAND3 (N12634, N12620, N9698, N12252);
buf BUF1 (N12635, N12626);
not NOT1 (N12636, N12635);
buf BUF1 (N12637, N12631);
and AND2 (N12638, N12630, N11626);
buf BUF1 (N12639, N12622);
not NOT1 (N12640, N12637);
nand NAND2 (N12641, N12632, N8809);
buf BUF1 (N12642, N12634);
not NOT1 (N12643, N12639);
nor NOR3 (N12644, N12641, N7307, N9332);
and AND4 (N12645, N12638, N172, N638, N7834);
or OR4 (N12646, N12636, N5516, N1372, N11999);
nor NOR3 (N12647, N12645, N7480, N3296);
not NOT1 (N12648, N12644);
nor NOR4 (N12649, N12646, N8991, N3684, N9634);
nor NOR4 (N12650, N12610, N11696, N10582, N5336);
nor NOR4 (N12651, N12647, N1403, N3442, N1874);
and AND4 (N12652, N12642, N1356, N354, N8642);
and AND2 (N12653, N12648, N10435);
nand NAND4 (N12654, N12653, N12067, N1076, N11752);
buf BUF1 (N12655, N12649);
xor XOR2 (N12656, N12625, N3979);
not NOT1 (N12657, N12652);
nor NOR3 (N12658, N12656, N2599, N763);
and AND4 (N12659, N12640, N186, N6012, N1161);
xor XOR2 (N12660, N12657, N10655);
and AND3 (N12661, N12660, N10929, N1124);
not NOT1 (N12662, N12658);
and AND2 (N12663, N12633, N3663);
xor XOR2 (N12664, N12629, N5491);
nor NOR3 (N12665, N12650, N3681, N10839);
not NOT1 (N12666, N12654);
nand NAND4 (N12667, N12643, N12453, N7522, N8666);
or OR4 (N12668, N12664, N796, N9313, N10117);
xor XOR2 (N12669, N12659, N2467);
or OR2 (N12670, N12663, N6061);
nor NOR3 (N12671, N12661, N9300, N6026);
nor NOR4 (N12672, N12667, N7326, N7545, N1075);
and AND4 (N12673, N12651, N6324, N11583, N7579);
nand NAND3 (N12674, N12655, N4398, N12593);
buf BUF1 (N12675, N12673);
and AND4 (N12676, N12672, N10604, N3396, N12072);
or OR4 (N12677, N12671, N1047, N11666, N1749);
or OR2 (N12678, N12666, N4471);
nand NAND2 (N12679, N12675, N696);
xor XOR2 (N12680, N12669, N551);
buf BUF1 (N12681, N12668);
or OR3 (N12682, N12681, N4713, N8653);
buf BUF1 (N12683, N12677);
or OR4 (N12684, N12670, N7765, N1255, N2919);
not NOT1 (N12685, N12665);
or OR4 (N12686, N12683, N732, N7352, N9285);
buf BUF1 (N12687, N12678);
nor NOR2 (N12688, N12680, N4891);
buf BUF1 (N12689, N12685);
not NOT1 (N12690, N12679);
and AND4 (N12691, N12688, N12503, N4492, N3063);
buf BUF1 (N12692, N12687);
not NOT1 (N12693, N12690);
nand NAND4 (N12694, N12684, N12318, N5103, N1172);
not NOT1 (N12695, N12662);
nand NAND3 (N12696, N12674, N2267, N7413);
and AND3 (N12697, N12695, N5854, N2473);
nand NAND3 (N12698, N12676, N9286, N9764);
nand NAND2 (N12699, N12697, N8825);
nor NOR3 (N12700, N12686, N1419, N1656);
nor NOR3 (N12701, N12700, N4068, N5451);
not NOT1 (N12702, N12692);
and AND2 (N12703, N12691, N8549);
nor NOR3 (N12704, N12698, N10210, N12271);
nor NOR4 (N12705, N12696, N10680, N5389, N6780);
and AND2 (N12706, N12693, N6182);
or OR2 (N12707, N12706, N12403);
xor XOR2 (N12708, N12707, N11793);
and AND2 (N12709, N12699, N6747);
xor XOR2 (N12710, N12702, N6964);
nand NAND3 (N12711, N12689, N9540, N2588);
nor NOR4 (N12712, N12682, N6292, N2171, N11970);
nand NAND3 (N12713, N12705, N12594, N12210);
not NOT1 (N12714, N12711);
or OR3 (N12715, N12694, N8870, N1830);
xor XOR2 (N12716, N12709, N11170);
and AND3 (N12717, N12701, N1841, N6765);
buf BUF1 (N12718, N12715);
or OR2 (N12719, N12713, N2851);
and AND2 (N12720, N12718, N10145);
or OR4 (N12721, N12703, N6325, N9280, N3642);
xor XOR2 (N12722, N12720, N3939);
or OR4 (N12723, N12712, N2508, N6877, N4603);
or OR3 (N12724, N12716, N124, N12201);
xor XOR2 (N12725, N12717, N5227);
or OR2 (N12726, N12704, N7898);
buf BUF1 (N12727, N12722);
or OR2 (N12728, N12710, N10328);
or OR3 (N12729, N12721, N9055, N10184);
nand NAND3 (N12730, N12728, N10151, N7550);
nand NAND3 (N12731, N12729, N12672, N1851);
nand NAND2 (N12732, N12727, N8885);
nand NAND4 (N12733, N12708, N3941, N8917, N8388);
nor NOR3 (N12734, N12731, N7467, N6627);
nor NOR2 (N12735, N12719, N9805);
nor NOR4 (N12736, N12734, N9900, N10935, N5453);
and AND3 (N12737, N12730, N6568, N9646);
or OR4 (N12738, N12726, N2463, N4875, N8784);
not NOT1 (N12739, N12737);
xor XOR2 (N12740, N12739, N9700);
and AND3 (N12741, N12714, N12293, N7021);
and AND3 (N12742, N12732, N4319, N8374);
not NOT1 (N12743, N12733);
nor NOR4 (N12744, N12743, N4092, N8846, N7520);
not NOT1 (N12745, N12725);
or OR4 (N12746, N12735, N6577, N10777, N12564);
nand NAND2 (N12747, N12741, N8560);
nor NOR2 (N12748, N12724, N12111);
buf BUF1 (N12749, N12723);
buf BUF1 (N12750, N12745);
or OR2 (N12751, N12736, N2326);
nand NAND2 (N12752, N12748, N5920);
buf BUF1 (N12753, N12751);
and AND4 (N12754, N12746, N9394, N7397, N1695);
buf BUF1 (N12755, N12747);
nor NOR4 (N12756, N12752, N12490, N4370, N582);
xor XOR2 (N12757, N12749, N39);
and AND2 (N12758, N12740, N10868);
xor XOR2 (N12759, N12758, N6373);
nor NOR4 (N12760, N12759, N5862, N626, N1674);
or OR3 (N12761, N12757, N10104, N319);
nand NAND2 (N12762, N12738, N6916);
or OR4 (N12763, N12744, N9632, N3870, N4355);
or OR2 (N12764, N12753, N1087);
nor NOR4 (N12765, N12756, N10691, N11656, N8311);
nor NOR2 (N12766, N12764, N5499);
not NOT1 (N12767, N12766);
not NOT1 (N12768, N12755);
not NOT1 (N12769, N12768);
not NOT1 (N12770, N12767);
and AND3 (N12771, N12762, N7354, N10497);
xor XOR2 (N12772, N12761, N5161);
xor XOR2 (N12773, N12742, N8686);
or OR2 (N12774, N12763, N3241);
not NOT1 (N12775, N12773);
and AND3 (N12776, N12771, N911, N10424);
xor XOR2 (N12777, N12775, N2382);
and AND3 (N12778, N12750, N6589, N10681);
nor NOR4 (N12779, N12772, N11849, N12252, N263);
xor XOR2 (N12780, N12777, N3571);
nor NOR3 (N12781, N12778, N11173, N10742);
xor XOR2 (N12782, N12754, N2348);
or OR4 (N12783, N12760, N2756, N5170, N11205);
and AND2 (N12784, N12781, N9758);
not NOT1 (N12785, N12780);
nor NOR3 (N12786, N12765, N10025, N883);
nor NOR4 (N12787, N12774, N5698, N7487, N12351);
nand NAND3 (N12788, N12785, N10687, N7946);
not NOT1 (N12789, N12783);
nor NOR2 (N12790, N12788, N4040);
not NOT1 (N12791, N12786);
buf BUF1 (N12792, N12782);
nor NOR4 (N12793, N12792, N8469, N595, N2548);
and AND4 (N12794, N12784, N89, N6729, N8956);
buf BUF1 (N12795, N12794);
not NOT1 (N12796, N12779);
xor XOR2 (N12797, N12791, N972);
or OR4 (N12798, N12787, N5085, N11857, N6795);
xor XOR2 (N12799, N12793, N7180);
nand NAND4 (N12800, N12789, N388, N4270, N8421);
or OR2 (N12801, N12776, N4357);
or OR2 (N12802, N12795, N83);
nand NAND2 (N12803, N12769, N10951);
and AND4 (N12804, N12790, N8415, N8862, N6833);
or OR2 (N12805, N12801, N859);
not NOT1 (N12806, N12797);
buf BUF1 (N12807, N12800);
nand NAND3 (N12808, N12803, N11881, N11755);
buf BUF1 (N12809, N12802);
not NOT1 (N12810, N12804);
nor NOR2 (N12811, N12810, N5762);
nand NAND4 (N12812, N12808, N11526, N3396, N11498);
or OR4 (N12813, N12796, N8249, N5773, N1148);
or OR3 (N12814, N12806, N9524, N5364);
xor XOR2 (N12815, N12811, N12056);
buf BUF1 (N12816, N12812);
not NOT1 (N12817, N12798);
nor NOR2 (N12818, N12807, N9306);
not NOT1 (N12819, N12815);
not NOT1 (N12820, N12809);
xor XOR2 (N12821, N12818, N10041);
buf BUF1 (N12822, N12821);
buf BUF1 (N12823, N12816);
or OR2 (N12824, N12770, N10116);
nand NAND2 (N12825, N12799, N1713);
buf BUF1 (N12826, N12825);
xor XOR2 (N12827, N12824, N3420);
xor XOR2 (N12828, N12805, N7626);
buf BUF1 (N12829, N12823);
nand NAND4 (N12830, N12827, N5815, N10486, N7895);
nor NOR2 (N12831, N12826, N10087);
and AND3 (N12832, N12814, N10183, N10722);
xor XOR2 (N12833, N12830, N792);
xor XOR2 (N12834, N12828, N3516);
xor XOR2 (N12835, N12813, N10361);
buf BUF1 (N12836, N12829);
nor NOR4 (N12837, N12832, N7931, N311, N9491);
buf BUF1 (N12838, N12834);
buf BUF1 (N12839, N12836);
and AND4 (N12840, N12839, N9569, N4133, N731);
nand NAND4 (N12841, N12835, N2985, N2979, N338);
or OR4 (N12842, N12817, N4281, N2800, N2067);
and AND2 (N12843, N12819, N10497);
nor NOR3 (N12844, N12842, N11354, N3093);
nand NAND4 (N12845, N12837, N1935, N12095, N12331);
xor XOR2 (N12846, N12841, N1143);
buf BUF1 (N12847, N12844);
nor NOR2 (N12848, N12822, N9564);
or OR3 (N12849, N12845, N2115, N11284);
nor NOR3 (N12850, N12831, N9830, N9888);
not NOT1 (N12851, N12846);
nand NAND4 (N12852, N12840, N786, N7082, N4485);
or OR2 (N12853, N12850, N4510);
and AND3 (N12854, N12848, N1557, N7884);
nand NAND3 (N12855, N12847, N7020, N2369);
nand NAND2 (N12856, N12820, N10291);
buf BUF1 (N12857, N12849);
or OR4 (N12858, N12843, N12401, N10823, N11124);
xor XOR2 (N12859, N12851, N5220);
or OR4 (N12860, N12859, N11339, N4171, N4948);
nor NOR4 (N12861, N12854, N8652, N5380, N5533);
nor NOR2 (N12862, N12857, N11845);
nand NAND4 (N12863, N12833, N7359, N1412, N197);
and AND3 (N12864, N12862, N6773, N2352);
or OR3 (N12865, N12856, N2183, N1932);
buf BUF1 (N12866, N12858);
xor XOR2 (N12867, N12860, N3277);
or OR4 (N12868, N12865, N11083, N3815, N11376);
and AND2 (N12869, N12855, N2568);
or OR2 (N12870, N12852, N1990);
xor XOR2 (N12871, N12869, N12512);
and AND4 (N12872, N12867, N11700, N10398, N2385);
buf BUF1 (N12873, N12870);
xor XOR2 (N12874, N12871, N346);
nor NOR4 (N12875, N12864, N5908, N3334, N1558);
nor NOR2 (N12876, N12853, N2144);
xor XOR2 (N12877, N12873, N6985);
not NOT1 (N12878, N12866);
not NOT1 (N12879, N12868);
buf BUF1 (N12880, N12838);
nor NOR4 (N12881, N12872, N2827, N7764, N5402);
nand NAND2 (N12882, N12878, N11565);
buf BUF1 (N12883, N12875);
not NOT1 (N12884, N12881);
or OR2 (N12885, N12874, N4848);
nand NAND2 (N12886, N12880, N3520);
buf BUF1 (N12887, N12877);
nand NAND2 (N12888, N12885, N1646);
buf BUF1 (N12889, N12876);
or OR2 (N12890, N12882, N4515);
and AND4 (N12891, N12888, N9003, N4581, N8301);
or OR3 (N12892, N12884, N2182, N1066);
and AND4 (N12893, N12887, N2437, N11742, N4242);
and AND3 (N12894, N12886, N11282, N8313);
and AND3 (N12895, N12891, N994, N11041);
buf BUF1 (N12896, N12883);
and AND2 (N12897, N12895, N523);
and AND2 (N12898, N12892, N427);
not NOT1 (N12899, N12889);
xor XOR2 (N12900, N12879, N2388);
and AND3 (N12901, N12890, N11081, N208);
nor NOR2 (N12902, N12896, N4064);
xor XOR2 (N12903, N12899, N3761);
xor XOR2 (N12904, N12900, N11565);
or OR2 (N12905, N12863, N9487);
nand NAND4 (N12906, N12901, N517, N1769, N9557);
and AND4 (N12907, N12893, N9077, N2566, N3803);
or OR4 (N12908, N12894, N7950, N2741, N11566);
nor NOR3 (N12909, N12897, N3777, N565);
or OR2 (N12910, N12898, N10996);
nand NAND2 (N12911, N12861, N7789);
buf BUF1 (N12912, N12910);
and AND3 (N12913, N12905, N4472, N4823);
or OR2 (N12914, N12911, N4444);
not NOT1 (N12915, N12908);
nand NAND2 (N12916, N12909, N11541);
nand NAND4 (N12917, N12907, N11676, N5721, N8378);
xor XOR2 (N12918, N12906, N2136);
not NOT1 (N12919, N12904);
not NOT1 (N12920, N12916);
and AND3 (N12921, N12915, N4431, N3769);
or OR2 (N12922, N12914, N12227);
or OR3 (N12923, N12919, N11375, N4771);
xor XOR2 (N12924, N12921, N1222);
and AND2 (N12925, N12917, N3015);
buf BUF1 (N12926, N12924);
and AND2 (N12927, N12918, N3590);
and AND2 (N12928, N12925, N11375);
or OR4 (N12929, N12903, N11039, N7914, N9968);
nand NAND2 (N12930, N12923, N12158);
xor XOR2 (N12931, N12913, N7534);
nand NAND4 (N12932, N12920, N12271, N3916, N9289);
buf BUF1 (N12933, N12922);
not NOT1 (N12934, N12929);
not NOT1 (N12935, N12932);
or OR4 (N12936, N12902, N12774, N8093, N12712);
not NOT1 (N12937, N12926);
xor XOR2 (N12938, N12935, N3811);
or OR2 (N12939, N12912, N125);
buf BUF1 (N12940, N12936);
nor NOR3 (N12941, N12937, N4409, N2595);
or OR4 (N12942, N12930, N1259, N7137, N2760);
buf BUF1 (N12943, N12939);
and AND4 (N12944, N12942, N3570, N11426, N1994);
and AND2 (N12945, N12934, N3715);
not NOT1 (N12946, N12941);
nand NAND3 (N12947, N12927, N430, N7561);
buf BUF1 (N12948, N12938);
nor NOR3 (N12949, N12943, N8359, N7501);
nand NAND2 (N12950, N12945, N12804);
or OR3 (N12951, N12950, N5100, N697);
not NOT1 (N12952, N12946);
xor XOR2 (N12953, N12940, N6437);
not NOT1 (N12954, N12952);
nand NAND3 (N12955, N12933, N9154, N9137);
nand NAND2 (N12956, N12928, N7868);
not NOT1 (N12957, N12956);
and AND2 (N12958, N12947, N12232);
nor NOR2 (N12959, N12949, N10189);
not NOT1 (N12960, N12944);
or OR3 (N12961, N12953, N1436, N6458);
nand NAND3 (N12962, N12958, N5361, N3099);
nand NAND3 (N12963, N12962, N5372, N1545);
buf BUF1 (N12964, N12951);
nand NAND2 (N12965, N12954, N10874);
nor NOR3 (N12966, N12963, N9980, N5193);
xor XOR2 (N12967, N12960, N6524);
xor XOR2 (N12968, N12957, N9283);
xor XOR2 (N12969, N12965, N5121);
or OR4 (N12970, N12948, N3439, N6702, N11650);
nor NOR3 (N12971, N12931, N10933, N3438);
not NOT1 (N12972, N12959);
and AND2 (N12973, N12968, N2793);
not NOT1 (N12974, N12973);
not NOT1 (N12975, N12964);
not NOT1 (N12976, N12955);
nor NOR3 (N12977, N12970, N3275, N12314);
or OR2 (N12978, N12977, N2436);
or OR4 (N12979, N12967, N8199, N12192, N11549);
xor XOR2 (N12980, N12978, N828);
xor XOR2 (N12981, N12975, N6909);
or OR4 (N12982, N12966, N748, N8106, N9506);
nand NAND2 (N12983, N12969, N9830);
or OR3 (N12984, N12976, N6017, N11321);
not NOT1 (N12985, N12979);
nor NOR2 (N12986, N12983, N755);
nor NOR2 (N12987, N12971, N9254);
buf BUF1 (N12988, N12961);
not NOT1 (N12989, N12984);
nand NAND2 (N12990, N12980, N10964);
nor NOR4 (N12991, N12974, N4376, N7925, N8465);
not NOT1 (N12992, N12987);
nor NOR3 (N12993, N12989, N9429, N9636);
nor NOR4 (N12994, N12972, N5515, N85, N9146);
xor XOR2 (N12995, N12990, N2212);
xor XOR2 (N12996, N12985, N1045);
xor XOR2 (N12997, N12992, N2111);
xor XOR2 (N12998, N12991, N2978);
or OR3 (N12999, N12995, N568, N8588);
buf BUF1 (N13000, N12998);
xor XOR2 (N13001, N12982, N629);
buf BUF1 (N13002, N13000);
nor NOR3 (N13003, N12993, N8017, N12504);
buf BUF1 (N13004, N13003);
xor XOR2 (N13005, N12988, N6669);
buf BUF1 (N13006, N13005);
nand NAND3 (N13007, N12997, N1323, N11057);
xor XOR2 (N13008, N13002, N6673);
nor NOR4 (N13009, N13006, N11263, N5666, N8861);
not NOT1 (N13010, N12999);
xor XOR2 (N13011, N13009, N1730);
xor XOR2 (N13012, N13007, N12732);
or OR2 (N13013, N13012, N2237);
nand NAND3 (N13014, N12986, N516, N2794);
not NOT1 (N13015, N12981);
xor XOR2 (N13016, N12994, N10831);
or OR3 (N13017, N13015, N9855, N8869);
or OR3 (N13018, N13001, N1609, N4524);
buf BUF1 (N13019, N13010);
buf BUF1 (N13020, N12996);
or OR4 (N13021, N13013, N5296, N2276, N10719);
buf BUF1 (N13022, N13020);
not NOT1 (N13023, N13016);
or OR4 (N13024, N13019, N4427, N5158, N1718);
buf BUF1 (N13025, N13004);
not NOT1 (N13026, N13025);
buf BUF1 (N13027, N13017);
or OR2 (N13028, N13022, N6717);
nand NAND3 (N13029, N13024, N2407, N12519);
xor XOR2 (N13030, N13027, N2191);
nor NOR4 (N13031, N13008, N5114, N6801, N2353);
buf BUF1 (N13032, N13026);
not NOT1 (N13033, N13021);
xor XOR2 (N13034, N13029, N10550);
buf BUF1 (N13035, N13030);
and AND2 (N13036, N13018, N12628);
buf BUF1 (N13037, N13031);
not NOT1 (N13038, N13035);
xor XOR2 (N13039, N13037, N8038);
or OR2 (N13040, N13011, N4084);
not NOT1 (N13041, N13036);
xor XOR2 (N13042, N13039, N4258);
xor XOR2 (N13043, N13014, N3896);
not NOT1 (N13044, N13033);
xor XOR2 (N13045, N13041, N4961);
and AND2 (N13046, N13043, N4222);
xor XOR2 (N13047, N13045, N4561);
and AND2 (N13048, N13038, N2720);
and AND4 (N13049, N13047, N2498, N5513, N8155);
nand NAND4 (N13050, N13028, N10101, N6591, N1927);
nor NOR2 (N13051, N13034, N4537);
not NOT1 (N13052, N13049);
and AND3 (N13053, N13046, N11652, N495);
and AND4 (N13054, N13044, N3790, N4064, N3492);
xor XOR2 (N13055, N13050, N7252);
nand NAND3 (N13056, N13023, N6884, N3401);
nor NOR2 (N13057, N13056, N11724);
nor NOR3 (N13058, N13052, N6975, N12564);
buf BUF1 (N13059, N13058);
nor NOR2 (N13060, N13042, N3141);
nand NAND3 (N13061, N13060, N2981, N234);
nand NAND4 (N13062, N13061, N11193, N5200, N3916);
nand NAND4 (N13063, N13057, N3111, N4561, N11899);
not NOT1 (N13064, N13059);
or OR3 (N13065, N13064, N3559, N9294);
nor NOR3 (N13066, N13048, N765, N9928);
buf BUF1 (N13067, N13054);
not NOT1 (N13068, N13051);
and AND2 (N13069, N13040, N11087);
and AND4 (N13070, N13066, N10329, N4760, N8941);
or OR2 (N13071, N13063, N8778);
or OR3 (N13072, N13068, N6017, N6470);
not NOT1 (N13073, N13067);
and AND2 (N13074, N13032, N6163);
buf BUF1 (N13075, N13071);
nand NAND3 (N13076, N13074, N6196, N1063);
and AND2 (N13077, N13075, N8008);
or OR4 (N13078, N13073, N9920, N1156, N5677);
or OR4 (N13079, N13069, N10651, N3690, N7105);
or OR2 (N13080, N13078, N9759);
nor NOR3 (N13081, N13055, N5229, N8962);
buf BUF1 (N13082, N13072);
nand NAND2 (N13083, N13053, N621);
nand NAND2 (N13084, N13079, N6428);
buf BUF1 (N13085, N13077);
nand NAND2 (N13086, N13084, N11502);
not NOT1 (N13087, N13083);
nand NAND4 (N13088, N13080, N8910, N7949, N7404);
and AND2 (N13089, N13081, N4741);
xor XOR2 (N13090, N13087, N3447);
nor NOR2 (N13091, N13062, N9108);
buf BUF1 (N13092, N13082);
not NOT1 (N13093, N13088);
not NOT1 (N13094, N13091);
nor NOR4 (N13095, N13086, N10733, N9935, N2890);
nand NAND2 (N13096, N13065, N7707);
xor XOR2 (N13097, N13090, N2888);
nand NAND4 (N13098, N13076, N13093, N4859, N9340);
xor XOR2 (N13099, N9889, N2765);
and AND4 (N13100, N13089, N2476, N12545, N9536);
and AND2 (N13101, N13070, N10293);
not NOT1 (N13102, N13092);
not NOT1 (N13103, N13096);
buf BUF1 (N13104, N13098);
and AND2 (N13105, N13094, N1895);
not NOT1 (N13106, N13102);
nor NOR3 (N13107, N13103, N1973, N7373);
xor XOR2 (N13108, N13085, N1750);
nor NOR3 (N13109, N13099, N10532, N5504);
xor XOR2 (N13110, N13104, N12599);
nor NOR4 (N13111, N13101, N277, N9537, N8116);
nor NOR4 (N13112, N13109, N6422, N6709, N9900);
not NOT1 (N13113, N13107);
and AND4 (N13114, N13111, N12299, N8664, N2063);
or OR3 (N13115, N13100, N4384, N9589);
and AND4 (N13116, N13114, N3296, N542, N264);
nor NOR2 (N13117, N13116, N7776);
and AND2 (N13118, N13108, N13083);
buf BUF1 (N13119, N13117);
xor XOR2 (N13120, N13106, N11821);
nor NOR2 (N13121, N13119, N881);
not NOT1 (N13122, N13118);
nor NOR2 (N13123, N13122, N652);
not NOT1 (N13124, N13110);
buf BUF1 (N13125, N13123);
nand NAND2 (N13126, N13105, N1866);
not NOT1 (N13127, N13095);
xor XOR2 (N13128, N13112, N1677);
nor NOR3 (N13129, N13127, N2980, N1073);
and AND3 (N13130, N13115, N9797, N11520);
nand NAND3 (N13131, N13097, N1410, N8172);
not NOT1 (N13132, N13124);
nand NAND3 (N13133, N13113, N5287, N9200);
nor NOR4 (N13134, N13120, N656, N1130, N10743);
xor XOR2 (N13135, N13121, N12677);
nand NAND2 (N13136, N13126, N8669);
or OR2 (N13137, N13125, N6462);
and AND2 (N13138, N13137, N7568);
nand NAND2 (N13139, N13128, N8869);
buf BUF1 (N13140, N13131);
nand NAND3 (N13141, N13140, N1671, N5485);
xor XOR2 (N13142, N13130, N11048);
not NOT1 (N13143, N13135);
xor XOR2 (N13144, N13143, N1234);
and AND4 (N13145, N13133, N6902, N11396, N787);
and AND3 (N13146, N13145, N12385, N865);
and AND3 (N13147, N13134, N6109, N7049);
buf BUF1 (N13148, N13138);
xor XOR2 (N13149, N13148, N193);
not NOT1 (N13150, N13136);
xor XOR2 (N13151, N13147, N13031);
and AND4 (N13152, N13144, N11354, N10910, N10021);
nor NOR3 (N13153, N13129, N4692, N4957);
nor NOR4 (N13154, N13150, N5736, N8534, N5360);
xor XOR2 (N13155, N13149, N12505);
nand NAND3 (N13156, N13139, N8382, N3120);
or OR2 (N13157, N13152, N3833);
and AND3 (N13158, N13132, N7639, N2458);
nand NAND3 (N13159, N13156, N9133, N8640);
nand NAND4 (N13160, N13154, N9671, N1024, N8157);
not NOT1 (N13161, N13158);
nor NOR2 (N13162, N13142, N11471);
xor XOR2 (N13163, N13141, N9882);
nor NOR3 (N13164, N13153, N4896, N13145);
nand NAND4 (N13165, N13157, N8775, N643, N1454);
or OR2 (N13166, N13146, N8323);
nor NOR2 (N13167, N13161, N11110);
not NOT1 (N13168, N13155);
buf BUF1 (N13169, N13167);
and AND2 (N13170, N13151, N2777);
nand NAND4 (N13171, N13163, N10509, N6556, N4023);
and AND3 (N13172, N13164, N10128, N3710);
xor XOR2 (N13173, N13166, N9275);
and AND4 (N13174, N13165, N12801, N1418, N8738);
and AND4 (N13175, N13174, N12011, N10648, N12417);
and AND3 (N13176, N13169, N3540, N8806);
nor NOR3 (N13177, N13159, N499, N389);
and AND4 (N13178, N13173, N9541, N3590, N1669);
nand NAND3 (N13179, N13171, N4902, N1017);
not NOT1 (N13180, N13179);
nand NAND2 (N13181, N13170, N10569);
nand NAND2 (N13182, N13177, N8558);
xor XOR2 (N13183, N13160, N2361);
xor XOR2 (N13184, N13175, N9866);
nand NAND2 (N13185, N13168, N5845);
and AND3 (N13186, N13172, N4734, N10194);
not NOT1 (N13187, N13183);
or OR4 (N13188, N13178, N9530, N13102, N1618);
xor XOR2 (N13189, N13176, N4776);
nand NAND4 (N13190, N13189, N8645, N2516, N8118);
or OR2 (N13191, N13162, N7801);
nand NAND4 (N13192, N13186, N12016, N7096, N12291);
not NOT1 (N13193, N13192);
nand NAND4 (N13194, N13193, N10726, N12611, N147);
buf BUF1 (N13195, N13191);
or OR2 (N13196, N13182, N12084);
not NOT1 (N13197, N13181);
or OR4 (N13198, N13188, N8321, N7950, N2571);
and AND4 (N13199, N13180, N9417, N11156, N7990);
and AND4 (N13200, N13185, N7302, N12727, N6479);
buf BUF1 (N13201, N13187);
xor XOR2 (N13202, N13197, N11348);
not NOT1 (N13203, N13190);
nor NOR4 (N13204, N13199, N6210, N5986, N11445);
nand NAND3 (N13205, N13184, N394, N3208);
or OR3 (N13206, N13203, N6170, N1808);
and AND4 (N13207, N13198, N1148, N5657, N821);
buf BUF1 (N13208, N13201);
nor NOR4 (N13209, N13204, N5683, N5069, N5160);
nand NAND3 (N13210, N13208, N1246, N2861);
buf BUF1 (N13211, N13205);
buf BUF1 (N13212, N13206);
or OR2 (N13213, N13210, N3709);
buf BUF1 (N13214, N13194);
buf BUF1 (N13215, N13207);
xor XOR2 (N13216, N13202, N12144);
xor XOR2 (N13217, N13216, N5635);
and AND2 (N13218, N13214, N7581);
not NOT1 (N13219, N13212);
nor NOR3 (N13220, N13200, N3933, N4555);
xor XOR2 (N13221, N13218, N11673);
nand NAND3 (N13222, N13220, N5718, N8960);
nand NAND2 (N13223, N13209, N5797);
nand NAND3 (N13224, N13222, N9987, N8571);
xor XOR2 (N13225, N13224, N9171);
nand NAND4 (N13226, N13217, N2997, N11866, N3809);
xor XOR2 (N13227, N13211, N8326);
not NOT1 (N13228, N13226);
nor NOR3 (N13229, N13196, N4107, N7636);
nand NAND3 (N13230, N13223, N7782, N9984);
not NOT1 (N13231, N13230);
or OR4 (N13232, N13219, N43, N4528, N8214);
and AND4 (N13233, N13232, N863, N7457, N5942);
and AND3 (N13234, N13231, N10808, N2266);
buf BUF1 (N13235, N13215);
or OR4 (N13236, N13229, N7868, N2407, N10468);
nor NOR4 (N13237, N13236, N5937, N10103, N8462);
or OR2 (N13238, N13195, N10009);
xor XOR2 (N13239, N13228, N1963);
or OR2 (N13240, N13237, N8330);
or OR2 (N13241, N13239, N6758);
buf BUF1 (N13242, N13213);
or OR2 (N13243, N13238, N3491);
and AND2 (N13244, N13240, N1981);
and AND4 (N13245, N13234, N10891, N11101, N6043);
nor NOR3 (N13246, N13227, N4084, N2985);
not NOT1 (N13247, N13244);
buf BUF1 (N13248, N13225);
and AND3 (N13249, N13235, N3096, N9229);
and AND2 (N13250, N13246, N2291);
or OR3 (N13251, N13241, N7252, N10659);
buf BUF1 (N13252, N13243);
or OR3 (N13253, N13248, N10547, N7978);
not NOT1 (N13254, N13221);
nor NOR3 (N13255, N13247, N13039, N12285);
xor XOR2 (N13256, N13252, N4251);
and AND2 (N13257, N13233, N9398);
or OR3 (N13258, N13257, N2536, N2332);
nor NOR3 (N13259, N13256, N9300, N4741);
not NOT1 (N13260, N13242);
xor XOR2 (N13261, N13258, N1946);
nand NAND2 (N13262, N13254, N12763);
not NOT1 (N13263, N13253);
xor XOR2 (N13264, N13250, N7943);
buf BUF1 (N13265, N13264);
not NOT1 (N13266, N13261);
xor XOR2 (N13267, N13263, N5721);
xor XOR2 (N13268, N13262, N2456);
not NOT1 (N13269, N13249);
xor XOR2 (N13270, N13266, N1380);
buf BUF1 (N13271, N13267);
nand NAND4 (N13272, N13259, N13244, N62, N2515);
and AND3 (N13273, N13270, N1453, N11009);
not NOT1 (N13274, N13273);
nand NAND3 (N13275, N13265, N5581, N162);
nand NAND3 (N13276, N13275, N2501, N4482);
buf BUF1 (N13277, N13269);
or OR2 (N13278, N13274, N2838);
nand NAND3 (N13279, N13268, N1357, N3060);
buf BUF1 (N13280, N13260);
nor NOR2 (N13281, N13278, N420);
buf BUF1 (N13282, N13245);
or OR4 (N13283, N13272, N8764, N10363, N10047);
nand NAND2 (N13284, N13276, N1419);
nand NAND4 (N13285, N13251, N11642, N2633, N2502);
nand NAND4 (N13286, N13271, N11347, N2226, N2327);
nand NAND4 (N13287, N13280, N4657, N1989, N238);
nor NOR2 (N13288, N13281, N12380);
buf BUF1 (N13289, N13284);
or OR2 (N13290, N13282, N11090);
and AND3 (N13291, N13289, N12736, N5962);
xor XOR2 (N13292, N13279, N7421);
not NOT1 (N13293, N13291);
nor NOR3 (N13294, N13255, N1425, N8048);
nor NOR4 (N13295, N13286, N2680, N12907, N7983);
buf BUF1 (N13296, N13292);
buf BUF1 (N13297, N13295);
and AND4 (N13298, N13290, N8678, N2418, N10299);
buf BUF1 (N13299, N13293);
xor XOR2 (N13300, N13294, N12508);
and AND2 (N13301, N13288, N5245);
or OR3 (N13302, N13277, N4433, N5177);
or OR2 (N13303, N13300, N6800);
nor NOR3 (N13304, N13299, N5051, N12848);
xor XOR2 (N13305, N13298, N285);
buf BUF1 (N13306, N13285);
xor XOR2 (N13307, N13287, N1390);
buf BUF1 (N13308, N13296);
nor NOR4 (N13309, N13303, N401, N12278, N4580);
or OR3 (N13310, N13309, N8684, N3652);
and AND3 (N13311, N13301, N5541, N4758);
xor XOR2 (N13312, N13306, N2928);
xor XOR2 (N13313, N13312, N1632);
and AND3 (N13314, N13297, N5269, N314);
nand NAND4 (N13315, N13307, N4663, N9036, N4652);
or OR4 (N13316, N13310, N5540, N9630, N6410);
not NOT1 (N13317, N13315);
nor NOR3 (N13318, N13304, N9354, N414);
nand NAND4 (N13319, N13311, N7605, N9613, N7586);
not NOT1 (N13320, N13302);
or OR3 (N13321, N13314, N2328, N11283);
not NOT1 (N13322, N13317);
and AND3 (N13323, N13322, N9060, N10402);
or OR4 (N13324, N13320, N2264, N8528, N4979);
nor NOR3 (N13325, N13319, N13265, N3293);
nand NAND4 (N13326, N13321, N4569, N12185, N7531);
nand NAND2 (N13327, N13308, N1595);
xor XOR2 (N13328, N13318, N7751);
nor NOR4 (N13329, N13325, N4873, N7288, N12834);
xor XOR2 (N13330, N13316, N2472);
and AND4 (N13331, N13328, N855, N11400, N6809);
buf BUF1 (N13332, N13323);
buf BUF1 (N13333, N13313);
xor XOR2 (N13334, N13329, N8790);
not NOT1 (N13335, N13334);
xor XOR2 (N13336, N13327, N2258);
xor XOR2 (N13337, N13324, N8328);
nand NAND2 (N13338, N13333, N7252);
nand NAND2 (N13339, N13338, N3622);
not NOT1 (N13340, N13335);
xor XOR2 (N13341, N13337, N1177);
or OR4 (N13342, N13336, N8569, N12089, N11429);
or OR4 (N13343, N13340, N11563, N7797, N11237);
and AND4 (N13344, N13326, N13143, N6353, N6980);
and AND3 (N13345, N13283, N4605, N5126);
or OR4 (N13346, N13342, N2804, N9811, N10590);
or OR2 (N13347, N13331, N5036);
xor XOR2 (N13348, N13332, N11573);
or OR3 (N13349, N13344, N8367, N734);
and AND2 (N13350, N13339, N8313);
not NOT1 (N13351, N13330);
nor NOR3 (N13352, N13345, N1895, N9336);
not NOT1 (N13353, N13347);
not NOT1 (N13354, N13348);
not NOT1 (N13355, N13354);
buf BUF1 (N13356, N13349);
xor XOR2 (N13357, N13353, N7402);
xor XOR2 (N13358, N13356, N3686);
and AND2 (N13359, N13346, N5897);
nor NOR3 (N13360, N13352, N1904, N10174);
or OR4 (N13361, N13360, N12909, N132, N10362);
not NOT1 (N13362, N13355);
xor XOR2 (N13363, N13350, N6645);
buf BUF1 (N13364, N13358);
and AND2 (N13365, N13343, N10221);
buf BUF1 (N13366, N13362);
nand NAND4 (N13367, N13351, N5906, N10252, N9648);
not NOT1 (N13368, N13359);
and AND4 (N13369, N13305, N10276, N2821, N2235);
or OR3 (N13370, N13367, N9899, N12698);
xor XOR2 (N13371, N13364, N264);
nand NAND4 (N13372, N13368, N4207, N859, N12061);
nand NAND4 (N13373, N13372, N12763, N11685, N4222);
nand NAND4 (N13374, N13341, N3277, N3897, N2945);
xor XOR2 (N13375, N13369, N1910);
not NOT1 (N13376, N13361);
nor NOR2 (N13377, N13375, N9200);
nand NAND3 (N13378, N13363, N8677, N212);
not NOT1 (N13379, N13365);
nand NAND2 (N13380, N13357, N5669);
buf BUF1 (N13381, N13377);
nand NAND3 (N13382, N13374, N13178, N10599);
not NOT1 (N13383, N13366);
buf BUF1 (N13384, N13378);
or OR2 (N13385, N13379, N8412);
not NOT1 (N13386, N13376);
xor XOR2 (N13387, N13371, N2862);
nor NOR3 (N13388, N13381, N5424, N2933);
nand NAND3 (N13389, N13385, N11535, N6537);
buf BUF1 (N13390, N13388);
xor XOR2 (N13391, N13370, N10393);
not NOT1 (N13392, N13387);
nor NOR2 (N13393, N13373, N12491);
not NOT1 (N13394, N13386);
not NOT1 (N13395, N13393);
nand NAND4 (N13396, N13382, N3359, N12586, N2647);
and AND4 (N13397, N13389, N7781, N2588, N8770);
xor XOR2 (N13398, N13391, N2892);
buf BUF1 (N13399, N13380);
and AND3 (N13400, N13390, N8039, N8118);
not NOT1 (N13401, N13395);
nand NAND4 (N13402, N13392, N3040, N10899, N3627);
nand NAND3 (N13403, N13399, N4615, N6521);
or OR2 (N13404, N13394, N1661);
and AND3 (N13405, N13398, N6447, N11385);
buf BUF1 (N13406, N13384);
not NOT1 (N13407, N13401);
not NOT1 (N13408, N13405);
nor NOR3 (N13409, N13402, N4391, N6717);
nor NOR2 (N13410, N13403, N598);
nor NOR2 (N13411, N13397, N11610);
or OR2 (N13412, N13400, N2306);
nor NOR2 (N13413, N13383, N7972);
nor NOR4 (N13414, N13410, N6385, N7732, N7545);
nor NOR4 (N13415, N13404, N4369, N7097, N1126);
not NOT1 (N13416, N13413);
not NOT1 (N13417, N13416);
not NOT1 (N13418, N13396);
or OR2 (N13419, N13409, N9726);
nand NAND3 (N13420, N13418, N5473, N8012);
not NOT1 (N13421, N13411);
buf BUF1 (N13422, N13407);
nand NAND4 (N13423, N13421, N9162, N5040, N12329);
nand NAND2 (N13424, N13414, N9728);
and AND2 (N13425, N13423, N4940);
xor XOR2 (N13426, N13419, N11000);
not NOT1 (N13427, N13424);
nand NAND4 (N13428, N13422, N7725, N3828, N7517);
buf BUF1 (N13429, N13412);
and AND2 (N13430, N13429, N13293);
or OR4 (N13431, N13420, N9754, N8522, N583);
buf BUF1 (N13432, N13406);
buf BUF1 (N13433, N13430);
and AND2 (N13434, N13427, N5633);
or OR2 (N13435, N13431, N714);
nor NOR2 (N13436, N13435, N6178);
and AND3 (N13437, N13425, N4529, N10986);
buf BUF1 (N13438, N13408);
or OR3 (N13439, N13417, N13234, N9186);
and AND3 (N13440, N13428, N4711, N12232);
and AND3 (N13441, N13426, N10696, N11265);
or OR3 (N13442, N13441, N7886, N12033);
nor NOR4 (N13443, N13436, N10488, N1195, N4777);
or OR4 (N13444, N13443, N134, N5436, N13194);
or OR4 (N13445, N13434, N3944, N391, N11986);
nor NOR2 (N13446, N13445, N13366);
xor XOR2 (N13447, N13433, N6340);
nand NAND3 (N13448, N13432, N797, N9953);
and AND2 (N13449, N13438, N5277);
nand NAND2 (N13450, N13448, N10036);
or OR2 (N13451, N13415, N105);
nand NAND4 (N13452, N13437, N1485, N10771, N3159);
buf BUF1 (N13453, N13439);
xor XOR2 (N13454, N13451, N6392);
and AND4 (N13455, N13447, N7612, N6970, N15);
buf BUF1 (N13456, N13450);
nand NAND2 (N13457, N13455, N8099);
nor NOR2 (N13458, N13440, N6596);
buf BUF1 (N13459, N13457);
buf BUF1 (N13460, N13459);
buf BUF1 (N13461, N13444);
nor NOR4 (N13462, N13442, N3359, N556, N3125);
buf BUF1 (N13463, N13446);
nor NOR2 (N13464, N13452, N3492);
or OR3 (N13465, N13464, N4952, N9554);
nor NOR2 (N13466, N13465, N4300);
or OR2 (N13467, N13456, N2089);
and AND3 (N13468, N13461, N5675, N10856);
nand NAND4 (N13469, N13466, N10611, N12005, N13237);
not NOT1 (N13470, N13454);
and AND3 (N13471, N13469, N2590, N5918);
nor NOR3 (N13472, N13453, N5041, N2738);
not NOT1 (N13473, N13468);
nor NOR3 (N13474, N13471, N10851, N1852);
not NOT1 (N13475, N13460);
or OR3 (N13476, N13467, N110, N9319);
nand NAND4 (N13477, N13474, N13363, N12776, N2715);
nor NOR4 (N13478, N13473, N4117, N2259, N6747);
nand NAND2 (N13479, N13449, N4197);
xor XOR2 (N13480, N13479, N5195);
xor XOR2 (N13481, N13462, N10731);
nand NAND3 (N13482, N13472, N7309, N5941);
nor NOR2 (N13483, N13481, N7089);
or OR3 (N13484, N13475, N3942, N12642);
not NOT1 (N13485, N13483);
nor NOR3 (N13486, N13480, N8901, N6736);
or OR2 (N13487, N13477, N6212);
and AND4 (N13488, N13487, N11477, N7996, N10229);
not NOT1 (N13489, N13458);
nand NAND3 (N13490, N13484, N11290, N8517);
nor NOR4 (N13491, N13486, N9783, N12197, N12868);
or OR2 (N13492, N13470, N1813);
nor NOR3 (N13493, N13489, N11789, N12204);
nor NOR3 (N13494, N13491, N3063, N2525);
xor XOR2 (N13495, N13476, N11187);
nor NOR2 (N13496, N13488, N12182);
not NOT1 (N13497, N13493);
nand NAND2 (N13498, N13497, N10526);
not NOT1 (N13499, N13498);
and AND2 (N13500, N13478, N6541);
not NOT1 (N13501, N13496);
xor XOR2 (N13502, N13499, N8022);
nor NOR2 (N13503, N13492, N414);
or OR4 (N13504, N13490, N1560, N7036, N4694);
nand NAND4 (N13505, N13501, N11545, N6732, N1895);
or OR4 (N13506, N13503, N11243, N144, N7699);
nor NOR4 (N13507, N13494, N2348, N9903, N3075);
or OR3 (N13508, N13504, N6120, N12026);
and AND4 (N13509, N13482, N8871, N13394, N13166);
nor NOR3 (N13510, N13506, N1265, N1519);
nor NOR2 (N13511, N13500, N299);
nand NAND4 (N13512, N13463, N12935, N8336, N525);
buf BUF1 (N13513, N13509);
or OR4 (N13514, N13485, N3281, N2005, N4213);
or OR4 (N13515, N13508, N1135, N6152, N5243);
or OR4 (N13516, N13513, N10220, N9718, N4658);
and AND4 (N13517, N13515, N9731, N6606, N6434);
and AND2 (N13518, N13511, N2638);
and AND3 (N13519, N13495, N1427, N12987);
or OR3 (N13520, N13516, N3634, N5141);
or OR2 (N13521, N13512, N1765);
nor NOR2 (N13522, N13514, N7749);
not NOT1 (N13523, N13510);
xor XOR2 (N13524, N13517, N5975);
nand NAND2 (N13525, N13519, N7956);
nor NOR3 (N13526, N13507, N1227, N13202);
xor XOR2 (N13527, N13522, N8196);
nand NAND3 (N13528, N13505, N11352, N9027);
xor XOR2 (N13529, N13525, N12909);
nor NOR2 (N13530, N13527, N10274);
or OR4 (N13531, N13529, N11381, N8404, N10084);
buf BUF1 (N13532, N13521);
nor NOR4 (N13533, N13518, N12054, N3039, N689);
or OR2 (N13534, N13532, N3406);
nand NAND3 (N13535, N13520, N6382, N965);
xor XOR2 (N13536, N13502, N512);
not NOT1 (N13537, N13535);
not NOT1 (N13538, N13537);
not NOT1 (N13539, N13524);
nand NAND2 (N13540, N13538, N3633);
buf BUF1 (N13541, N13523);
and AND3 (N13542, N13536, N6115, N10728);
nand NAND4 (N13543, N13540, N6005, N2576, N8575);
not NOT1 (N13544, N13534);
nor NOR4 (N13545, N13533, N5648, N4733, N1743);
buf BUF1 (N13546, N13528);
not NOT1 (N13547, N13543);
xor XOR2 (N13548, N13544, N5125);
not NOT1 (N13549, N13539);
nand NAND4 (N13550, N13530, N5221, N4852, N3845);
and AND3 (N13551, N13526, N6757, N12147);
xor XOR2 (N13552, N13542, N8706);
xor XOR2 (N13553, N13550, N8859);
buf BUF1 (N13554, N13541);
xor XOR2 (N13555, N13549, N4283);
not NOT1 (N13556, N13551);
buf BUF1 (N13557, N13556);
xor XOR2 (N13558, N13546, N5267);
buf BUF1 (N13559, N13554);
not NOT1 (N13560, N13558);
and AND4 (N13561, N13559, N5402, N3, N3857);
xor XOR2 (N13562, N13557, N5623);
not NOT1 (N13563, N13552);
not NOT1 (N13564, N13531);
xor XOR2 (N13565, N13562, N13504);
and AND4 (N13566, N13565, N6015, N1175, N554);
nand NAND3 (N13567, N13547, N12389, N8987);
not NOT1 (N13568, N13563);
or OR2 (N13569, N13566, N4994);
nand NAND3 (N13570, N13555, N9077, N2392);
buf BUF1 (N13571, N13560);
not NOT1 (N13572, N13553);
and AND4 (N13573, N13568, N572, N12117, N4178);
nor NOR2 (N13574, N13561, N4406);
nor NOR3 (N13575, N13572, N11943, N9515);
nor NOR4 (N13576, N13564, N5096, N1350, N8047);
xor XOR2 (N13577, N13574, N2361);
not NOT1 (N13578, N13569);
and AND2 (N13579, N13567, N6828);
nor NOR2 (N13580, N13548, N6359);
not NOT1 (N13581, N13575);
nand NAND3 (N13582, N13580, N10258, N12280);
nand NAND2 (N13583, N13582, N13145);
buf BUF1 (N13584, N13578);
buf BUF1 (N13585, N13577);
nand NAND2 (N13586, N13585, N5698);
and AND4 (N13587, N13579, N6494, N12996, N4969);
or OR2 (N13588, N13573, N10698);
or OR2 (N13589, N13570, N4158);
not NOT1 (N13590, N13571);
and AND2 (N13591, N13589, N10285);
not NOT1 (N13592, N13581);
nor NOR3 (N13593, N13591, N13589, N12697);
nand NAND3 (N13594, N13588, N6925, N9100);
or OR4 (N13595, N13592, N10392, N12879, N7332);
nand NAND2 (N13596, N13545, N271);
not NOT1 (N13597, N13583);
buf BUF1 (N13598, N13576);
buf BUF1 (N13599, N13595);
or OR2 (N13600, N13599, N9677);
or OR2 (N13601, N13593, N2959);
or OR3 (N13602, N13600, N3096, N5664);
not NOT1 (N13603, N13598);
and AND3 (N13604, N13587, N1603, N7107);
buf BUF1 (N13605, N13594);
or OR4 (N13606, N13584, N10997, N6115, N13266);
or OR4 (N13607, N13601, N11493, N2701, N7137);
nand NAND2 (N13608, N13602, N2147);
and AND2 (N13609, N13604, N4019);
or OR3 (N13610, N13596, N7908, N5987);
not NOT1 (N13611, N13608);
nand NAND2 (N13612, N13586, N735);
nor NOR2 (N13613, N13612, N11198);
not NOT1 (N13614, N13590);
nor NOR2 (N13615, N13614, N8250);
or OR3 (N13616, N13609, N2073, N12213);
nor NOR3 (N13617, N13611, N3950, N8079);
and AND2 (N13618, N13607, N10549);
nand NAND3 (N13619, N13615, N9976, N1411);
not NOT1 (N13620, N13619);
and AND2 (N13621, N13618, N3116);
and AND2 (N13622, N13617, N4216);
or OR3 (N13623, N13622, N10869, N11422);
or OR2 (N13624, N13603, N4577);
buf BUF1 (N13625, N13616);
buf BUF1 (N13626, N13624);
buf BUF1 (N13627, N13626);
or OR3 (N13628, N13621, N7516, N10161);
nand NAND4 (N13629, N13605, N6138, N148, N10592);
nor NOR4 (N13630, N13628, N950, N92, N13542);
xor XOR2 (N13631, N13597, N7648);
nand NAND3 (N13632, N13620, N9233, N11257);
or OR2 (N13633, N13627, N9923);
xor XOR2 (N13634, N13629, N5677);
and AND4 (N13635, N13625, N11586, N9017, N2296);
or OR2 (N13636, N13633, N9068);
nor NOR3 (N13637, N13636, N10695, N9369);
buf BUF1 (N13638, N13637);
nor NOR2 (N13639, N13632, N12237);
and AND4 (N13640, N13610, N4653, N9114, N3942);
nand NAND3 (N13641, N13640, N10251, N8546);
xor XOR2 (N13642, N13631, N9653);
nand NAND4 (N13643, N13606, N5370, N9171, N2610);
nand NAND4 (N13644, N13638, N4483, N7844, N2313);
xor XOR2 (N13645, N13613, N1589);
buf BUF1 (N13646, N13623);
and AND3 (N13647, N13644, N2883, N111);
and AND2 (N13648, N13646, N8199);
nor NOR4 (N13649, N13630, N267, N5206, N8389);
and AND4 (N13650, N13639, N11679, N4642, N2604);
and AND4 (N13651, N13650, N784, N1499, N739);
nand NAND4 (N13652, N13645, N1492, N8590, N4053);
nand NAND2 (N13653, N13648, N8979);
nor NOR4 (N13654, N13635, N13429, N10970, N12981);
buf BUF1 (N13655, N13641);
nand NAND2 (N13656, N13652, N5426);
nor NOR4 (N13657, N13655, N11241, N4715, N2692);
nor NOR4 (N13658, N13653, N6880, N841, N3919);
xor XOR2 (N13659, N13658, N6938);
and AND2 (N13660, N13657, N9518);
nor NOR2 (N13661, N13643, N4849);
nand NAND2 (N13662, N13654, N228);
xor XOR2 (N13663, N13662, N6398);
nand NAND2 (N13664, N13663, N8827);
nor NOR2 (N13665, N13647, N687);
nand NAND4 (N13666, N13649, N684, N2924, N6477);
or OR4 (N13667, N13660, N7481, N102, N2165);
nor NOR4 (N13668, N13634, N12396, N1030, N3245);
nor NOR2 (N13669, N13666, N10922);
xor XOR2 (N13670, N13661, N13183);
or OR2 (N13671, N13667, N12721);
and AND4 (N13672, N13668, N9762, N6258, N13663);
and AND2 (N13673, N13671, N11086);
nand NAND2 (N13674, N13659, N1145);
and AND2 (N13675, N13672, N11424);
nor NOR2 (N13676, N13651, N9774);
nor NOR2 (N13677, N13674, N11964);
and AND3 (N13678, N13676, N8479, N11142);
nor NOR2 (N13679, N13670, N13343);
buf BUF1 (N13680, N13679);
buf BUF1 (N13681, N13665);
buf BUF1 (N13682, N13675);
nor NOR4 (N13683, N13669, N12877, N1828, N12457);
nand NAND3 (N13684, N13681, N11887, N3366);
buf BUF1 (N13685, N13664);
and AND2 (N13686, N13642, N6913);
not NOT1 (N13687, N13673);
not NOT1 (N13688, N13683);
buf BUF1 (N13689, N13687);
and AND2 (N13690, N13685, N2145);
or OR3 (N13691, N13682, N8347, N5545);
not NOT1 (N13692, N13688);
or OR4 (N13693, N13691, N12844, N8313, N8012);
buf BUF1 (N13694, N13686);
and AND2 (N13695, N13693, N11987);
xor XOR2 (N13696, N13677, N5984);
not NOT1 (N13697, N13684);
or OR2 (N13698, N13697, N13196);
or OR4 (N13699, N13656, N7126, N6519, N9701);
not NOT1 (N13700, N13678);
buf BUF1 (N13701, N13699);
nand NAND2 (N13702, N13694, N2037);
or OR2 (N13703, N13696, N3869);
not NOT1 (N13704, N13702);
not NOT1 (N13705, N13695);
not NOT1 (N13706, N13705);
xor XOR2 (N13707, N13692, N8767);
nor NOR2 (N13708, N13703, N4389);
nor NOR3 (N13709, N13706, N1627, N9818);
xor XOR2 (N13710, N13689, N5856);
and AND2 (N13711, N13709, N3305);
not NOT1 (N13712, N13680);
and AND3 (N13713, N13704, N9912, N12531);
not NOT1 (N13714, N13710);
or OR2 (N13715, N13713, N13400);
nand NAND2 (N13716, N13708, N435);
not NOT1 (N13717, N13715);
buf BUF1 (N13718, N13716);
or OR4 (N13719, N13701, N1882, N5426, N1938);
nand NAND4 (N13720, N13717, N6344, N1671, N4224);
nand NAND4 (N13721, N13712, N13125, N4103, N3729);
xor XOR2 (N13722, N13690, N1046);
buf BUF1 (N13723, N13714);
nor NOR4 (N13724, N13721, N32, N9908, N3878);
nand NAND4 (N13725, N13707, N13690, N3114, N5086);
nand NAND4 (N13726, N13723, N3547, N2325, N13638);
and AND3 (N13727, N13722, N12641, N12020);
nor NOR3 (N13728, N13727, N9899, N10966);
xor XOR2 (N13729, N13720, N12695);
xor XOR2 (N13730, N13700, N12790);
xor XOR2 (N13731, N13728, N582);
nand NAND4 (N13732, N13698, N2782, N2467, N11223);
nor NOR4 (N13733, N13729, N4919, N11428, N7725);
nand NAND4 (N13734, N13724, N6208, N7455, N1477);
xor XOR2 (N13735, N13734, N5878);
nand NAND2 (N13736, N13733, N3059);
or OR3 (N13737, N13732, N7172, N8922);
buf BUF1 (N13738, N13736);
nor NOR2 (N13739, N13711, N7004);
nor NOR4 (N13740, N13725, N2726, N5492, N7965);
or OR2 (N13741, N13740, N10937);
buf BUF1 (N13742, N13737);
xor XOR2 (N13743, N13742, N7187);
nand NAND4 (N13744, N13719, N4251, N8764, N10684);
xor XOR2 (N13745, N13739, N12456);
xor XOR2 (N13746, N13745, N6650);
xor XOR2 (N13747, N13735, N3750);
nand NAND3 (N13748, N13744, N983, N10748);
and AND2 (N13749, N13746, N6266);
and AND3 (N13750, N13741, N9007, N13560);
or OR2 (N13751, N13749, N10953);
not NOT1 (N13752, N13730);
not NOT1 (N13753, N13718);
buf BUF1 (N13754, N13731);
and AND3 (N13755, N13743, N9170, N10707);
or OR3 (N13756, N13738, N7125, N11582);
buf BUF1 (N13757, N13755);
buf BUF1 (N13758, N13757);
not NOT1 (N13759, N13756);
and AND2 (N13760, N13751, N8477);
not NOT1 (N13761, N13752);
nand NAND4 (N13762, N13753, N1428, N4270, N12934);
buf BUF1 (N13763, N13762);
buf BUF1 (N13764, N13763);
buf BUF1 (N13765, N13754);
xor XOR2 (N13766, N13761, N7639);
not NOT1 (N13767, N13747);
and AND3 (N13768, N13748, N13397, N8090);
not NOT1 (N13769, N13768);
nand NAND3 (N13770, N13765, N10832, N6315);
nor NOR2 (N13771, N13766, N12091);
buf BUF1 (N13772, N13771);
or OR4 (N13773, N13767, N10530, N2997, N1534);
or OR4 (N13774, N13726, N13635, N1156, N8224);
nor NOR4 (N13775, N13750, N13458, N7335, N7363);
or OR4 (N13776, N13764, N12104, N10663, N7284);
or OR4 (N13777, N13774, N10037, N13607, N135);
not NOT1 (N13778, N13769);
buf BUF1 (N13779, N13760);
or OR3 (N13780, N13770, N1916, N9885);
nor NOR4 (N13781, N13772, N4062, N4471, N9265);
and AND2 (N13782, N13780, N8654);
nand NAND3 (N13783, N13781, N11566, N8435);
not NOT1 (N13784, N13775);
not NOT1 (N13785, N13784);
or OR3 (N13786, N13777, N5005, N9941);
nand NAND4 (N13787, N13778, N7313, N2006, N11472);
xor XOR2 (N13788, N13773, N9618);
buf BUF1 (N13789, N13783);
or OR3 (N13790, N13787, N6206, N1477);
and AND3 (N13791, N13759, N2456, N286);
nand NAND2 (N13792, N13789, N9570);
nor NOR4 (N13793, N13779, N11997, N6748, N2071);
buf BUF1 (N13794, N13788);
not NOT1 (N13795, N13782);
not NOT1 (N13796, N13785);
buf BUF1 (N13797, N13792);
nor NOR4 (N13798, N13790, N1724, N8192, N6083);
nand NAND2 (N13799, N13797, N8017);
not NOT1 (N13800, N13793);
nand NAND2 (N13801, N13786, N13333);
nor NOR4 (N13802, N13796, N2325, N4191, N579);
nand NAND2 (N13803, N13776, N13775);
not NOT1 (N13804, N13791);
nor NOR3 (N13805, N13758, N13075, N4485);
nor NOR2 (N13806, N13799, N8353);
nand NAND2 (N13807, N13802, N3653);
nor NOR4 (N13808, N13794, N1512, N10371, N12019);
nand NAND4 (N13809, N13801, N10232, N4434, N2130);
nor NOR3 (N13810, N13809, N224, N5916);
and AND3 (N13811, N13803, N9192, N6931);
nor NOR3 (N13812, N13795, N5274, N5214);
or OR2 (N13813, N13806, N9593);
and AND4 (N13814, N13804, N3644, N2712, N13048);
not NOT1 (N13815, N13807);
or OR3 (N13816, N13798, N9783, N11742);
and AND4 (N13817, N13810, N8139, N4659, N7373);
and AND4 (N13818, N13811, N4519, N11318, N12005);
and AND3 (N13819, N13812, N745, N12583);
and AND2 (N13820, N13800, N9297);
nand NAND3 (N13821, N13813, N13786, N11770);
nor NOR4 (N13822, N13820, N5508, N8113, N8310);
or OR2 (N13823, N13816, N9871);
and AND4 (N13824, N13817, N8335, N935, N10822);
buf BUF1 (N13825, N13822);
buf BUF1 (N13826, N13819);
buf BUF1 (N13827, N13815);
buf BUF1 (N13828, N13805);
nor NOR3 (N13829, N13823, N10695, N3389);
nor NOR4 (N13830, N13808, N1032, N3565, N5929);
nand NAND3 (N13831, N13814, N6986, N2074);
nand NAND4 (N13832, N13826, N3623, N6625, N8582);
buf BUF1 (N13833, N13831);
and AND2 (N13834, N13829, N12118);
or OR4 (N13835, N13828, N8939, N7312, N4779);
xor XOR2 (N13836, N13830, N11815);
and AND2 (N13837, N13834, N8727);
nor NOR4 (N13838, N13825, N11583, N822, N13674);
xor XOR2 (N13839, N13821, N9592);
or OR2 (N13840, N13838, N7068);
and AND2 (N13841, N13824, N6046);
nand NAND3 (N13842, N13827, N3828, N7781);
nand NAND4 (N13843, N13836, N1562, N8682, N11307);
or OR2 (N13844, N13835, N7544);
not NOT1 (N13845, N13818);
xor XOR2 (N13846, N13837, N204);
not NOT1 (N13847, N13842);
buf BUF1 (N13848, N13839);
or OR2 (N13849, N13845, N11222);
nor NOR2 (N13850, N13844, N10468);
nand NAND2 (N13851, N13850, N1372);
xor XOR2 (N13852, N13847, N9666);
nor NOR4 (N13853, N13852, N11419, N11967, N9701);
xor XOR2 (N13854, N13848, N8299);
and AND3 (N13855, N13833, N9598, N12621);
not NOT1 (N13856, N13846);
xor XOR2 (N13857, N13843, N6449);
or OR4 (N13858, N13832, N4971, N5334, N6602);
nand NAND3 (N13859, N13858, N1121, N5895);
xor XOR2 (N13860, N13853, N383);
nor NOR3 (N13861, N13840, N6211, N12614);
not NOT1 (N13862, N13860);
nor NOR4 (N13863, N13856, N663, N10470, N3192);
nor NOR4 (N13864, N13855, N10622, N13222, N2126);
nand NAND4 (N13865, N13857, N3848, N8279, N13438);
or OR4 (N13866, N13849, N10749, N13622, N10848);
buf BUF1 (N13867, N13859);
nor NOR4 (N13868, N13841, N10323, N9823, N11171);
nand NAND4 (N13869, N13863, N5432, N2769, N7512);
not NOT1 (N13870, N13865);
not NOT1 (N13871, N13864);
buf BUF1 (N13872, N13851);
or OR3 (N13873, N13867, N13257, N4272);
and AND2 (N13874, N13862, N13635);
nor NOR4 (N13875, N13870, N13339, N5397, N3088);
and AND3 (N13876, N13866, N4375, N3928);
and AND3 (N13877, N13869, N4656, N3964);
and AND3 (N13878, N13873, N6046, N10095);
and AND4 (N13879, N13878, N9007, N9797, N12000);
not NOT1 (N13880, N13861);
not NOT1 (N13881, N13879);
and AND4 (N13882, N13876, N1682, N9972, N3234);
xor XOR2 (N13883, N13882, N9307);
nand NAND2 (N13884, N13854, N9618);
not NOT1 (N13885, N13875);
nand NAND4 (N13886, N13883, N5699, N4839, N10029);
nand NAND4 (N13887, N13886, N8185, N7295, N13260);
not NOT1 (N13888, N13885);
or OR4 (N13889, N13872, N4139, N10264, N11797);
or OR3 (N13890, N13877, N3699, N647);
not NOT1 (N13891, N13871);
not NOT1 (N13892, N13884);
not NOT1 (N13893, N13874);
or OR2 (N13894, N13888, N3001);
not NOT1 (N13895, N13891);
not NOT1 (N13896, N13894);
and AND2 (N13897, N13881, N5190);
nand NAND3 (N13898, N13868, N1725, N1006);
nor NOR3 (N13899, N13897, N11824, N3724);
or OR3 (N13900, N13895, N2571, N13543);
nor NOR4 (N13901, N13890, N10134, N6262, N1841);
xor XOR2 (N13902, N13899, N4998);
and AND3 (N13903, N13900, N2253, N8914);
and AND3 (N13904, N13903, N4146, N5260);
xor XOR2 (N13905, N13887, N7341);
and AND3 (N13906, N13896, N12526, N4093);
xor XOR2 (N13907, N13905, N5450);
nand NAND2 (N13908, N13880, N5268);
or OR3 (N13909, N13898, N5847, N12701);
or OR4 (N13910, N13909, N3633, N9348, N13373);
buf BUF1 (N13911, N13906);
nor NOR3 (N13912, N13893, N8863, N11213);
nand NAND2 (N13913, N13910, N13855);
xor XOR2 (N13914, N13907, N12683);
nand NAND3 (N13915, N13911, N7487, N12928);
nor NOR3 (N13916, N13913, N4637, N9849);
or OR2 (N13917, N13914, N5206);
nor NOR3 (N13918, N13908, N2367, N5654);
and AND3 (N13919, N13912, N4908, N6615);
xor XOR2 (N13920, N13904, N3955);
nor NOR3 (N13921, N13920, N8711, N9295);
nor NOR3 (N13922, N13901, N925, N6748);
not NOT1 (N13923, N13922);
xor XOR2 (N13924, N13919, N6217);
nor NOR4 (N13925, N13923, N7036, N1042, N3717);
not NOT1 (N13926, N13917);
and AND4 (N13927, N13915, N4787, N7452, N131);
not NOT1 (N13928, N13926);
nand NAND4 (N13929, N13928, N336, N9452, N9004);
xor XOR2 (N13930, N13889, N5185);
or OR4 (N13931, N13927, N8107, N3116, N8123);
buf BUF1 (N13932, N13921);
xor XOR2 (N13933, N13930, N6724);
and AND2 (N13934, N13925, N2865);
nor NOR2 (N13935, N13929, N6550);
not NOT1 (N13936, N13924);
nand NAND3 (N13937, N13931, N10406, N6230);
xor XOR2 (N13938, N13916, N13393);
xor XOR2 (N13939, N13892, N2305);
or OR4 (N13940, N13935, N10483, N13097, N5972);
buf BUF1 (N13941, N13940);
not NOT1 (N13942, N13902);
xor XOR2 (N13943, N13932, N10376);
or OR3 (N13944, N13941, N12843, N2803);
and AND2 (N13945, N13939, N11343);
not NOT1 (N13946, N13918);
nand NAND2 (N13947, N13938, N13271);
and AND4 (N13948, N13947, N12850, N7216, N5151);
nand NAND4 (N13949, N13945, N835, N10151, N8394);
nor NOR3 (N13950, N13943, N5585, N4204);
and AND4 (N13951, N13950, N9733, N8444, N10632);
buf BUF1 (N13952, N13942);
nand NAND4 (N13953, N13934, N2474, N3803, N9213);
nor NOR2 (N13954, N13933, N8522);
not NOT1 (N13955, N13952);
not NOT1 (N13956, N13954);
and AND2 (N13957, N13956, N9031);
not NOT1 (N13958, N13936);
and AND2 (N13959, N13946, N5689);
or OR2 (N13960, N13951, N5816);
buf BUF1 (N13961, N13958);
xor XOR2 (N13962, N13955, N9771);
xor XOR2 (N13963, N13957, N8595);
and AND3 (N13964, N13962, N5417, N494);
xor XOR2 (N13965, N13964, N9955);
not NOT1 (N13966, N13960);
buf BUF1 (N13967, N13961);
xor XOR2 (N13968, N13949, N8240);
nor NOR3 (N13969, N13963, N10577, N387);
buf BUF1 (N13970, N13948);
nand NAND2 (N13971, N13965, N4133);
not NOT1 (N13972, N13944);
nand NAND4 (N13973, N13966, N4709, N2795, N10565);
and AND2 (N13974, N13937, N5967);
not NOT1 (N13975, N13967);
nor NOR2 (N13976, N13974, N2969);
and AND4 (N13977, N13972, N8592, N9952, N13621);
or OR4 (N13978, N13970, N13591, N8177, N13557);
or OR2 (N13979, N13975, N2284);
not NOT1 (N13980, N13979);
not NOT1 (N13981, N13968);
not NOT1 (N13982, N13978);
not NOT1 (N13983, N13953);
xor XOR2 (N13984, N13971, N1358);
not NOT1 (N13985, N13982);
or OR3 (N13986, N13959, N2954, N13660);
nand NAND4 (N13987, N13973, N11539, N6019, N6658);
and AND3 (N13988, N13981, N2035, N8947);
nand NAND4 (N13989, N13976, N13199, N9834, N8672);
or OR3 (N13990, N13984, N9461, N11704);
xor XOR2 (N13991, N13980, N1800);
nor NOR4 (N13992, N13977, N1771, N7726, N12102);
not NOT1 (N13993, N13988);
xor XOR2 (N13994, N13992, N5163);
and AND3 (N13995, N13994, N786, N1819);
nor NOR2 (N13996, N13985, N2487);
nor NOR4 (N13997, N13990, N12320, N5574, N5680);
nor NOR2 (N13998, N13997, N13209);
xor XOR2 (N13999, N13995, N5208);
xor XOR2 (N14000, N13987, N4659);
xor XOR2 (N14001, N13986, N11090);
or OR4 (N14002, N14000, N6290, N5528, N11374);
nor NOR2 (N14003, N13999, N2626);
xor XOR2 (N14004, N13993, N6786);
xor XOR2 (N14005, N13983, N12587);
or OR3 (N14006, N13969, N6253, N13086);
and AND3 (N14007, N14005, N4608, N331);
not NOT1 (N14008, N14003);
nor NOR2 (N14009, N14004, N4918);
buf BUF1 (N14010, N14007);
or OR3 (N14011, N13996, N4499, N1320);
or OR3 (N14012, N14011, N3935, N13985);
nand NAND4 (N14013, N14001, N4420, N7257, N8977);
or OR3 (N14014, N14012, N9032, N663);
or OR2 (N14015, N13998, N4642);
buf BUF1 (N14016, N14006);
nor NOR2 (N14017, N14016, N13126);
nand NAND2 (N14018, N14015, N4219);
not NOT1 (N14019, N14008);
or OR2 (N14020, N14018, N5275);
nand NAND3 (N14021, N14014, N9518, N1517);
nand NAND4 (N14022, N14019, N595, N13254, N8768);
buf BUF1 (N14023, N14020);
not NOT1 (N14024, N14022);
buf BUF1 (N14025, N14021);
and AND4 (N14026, N14024, N7471, N9583, N1062);
nor NOR3 (N14027, N13989, N5627, N3726);
nor NOR2 (N14028, N14010, N8752);
not NOT1 (N14029, N13991);
and AND2 (N14030, N14028, N10558);
or OR4 (N14031, N14026, N6889, N5548, N10852);
nand NAND3 (N14032, N14017, N2141, N8234);
buf BUF1 (N14033, N14030);
xor XOR2 (N14034, N14002, N2167);
or OR2 (N14035, N14025, N11987);
and AND3 (N14036, N14029, N11521, N3133);
xor XOR2 (N14037, N14027, N4162);
not NOT1 (N14038, N14023);
nor NOR3 (N14039, N14036, N8293, N12692);
xor XOR2 (N14040, N14039, N6741);
buf BUF1 (N14041, N14031);
or OR2 (N14042, N14041, N13306);
buf BUF1 (N14043, N14042);
buf BUF1 (N14044, N14038);
nand NAND3 (N14045, N14044, N1286, N12202);
buf BUF1 (N14046, N14013);
xor XOR2 (N14047, N14045, N4284);
not NOT1 (N14048, N14047);
buf BUF1 (N14049, N14043);
not NOT1 (N14050, N14034);
buf BUF1 (N14051, N14050);
buf BUF1 (N14052, N14048);
nor NOR4 (N14053, N14032, N3703, N11851, N1660);
not NOT1 (N14054, N14052);
nor NOR2 (N14055, N14051, N1876);
nand NAND4 (N14056, N14054, N10741, N10338, N11252);
nand NAND2 (N14057, N14056, N3377);
or OR4 (N14058, N14049, N11910, N8409, N6083);
nand NAND2 (N14059, N14037, N5024);
nor NOR2 (N14060, N14059, N10578);
and AND2 (N14061, N14046, N8453);
and AND3 (N14062, N14040, N5952, N10394);
buf BUF1 (N14063, N14062);
nor NOR2 (N14064, N14033, N6357);
and AND2 (N14065, N14009, N13231);
buf BUF1 (N14066, N14064);
nand NAND4 (N14067, N14055, N2952, N3601, N9214);
buf BUF1 (N14068, N14053);
nor NOR2 (N14069, N14066, N2452);
not NOT1 (N14070, N14060);
not NOT1 (N14071, N14058);
not NOT1 (N14072, N14068);
nand NAND3 (N14073, N14067, N1674, N12333);
buf BUF1 (N14074, N14063);
nor NOR3 (N14075, N14065, N9313, N6200);
not NOT1 (N14076, N14071);
or OR3 (N14077, N14073, N2541, N5180);
not NOT1 (N14078, N14035);
not NOT1 (N14079, N14074);
or OR4 (N14080, N14079, N527, N3807, N9927);
not NOT1 (N14081, N14061);
xor XOR2 (N14082, N14069, N4989);
and AND3 (N14083, N14078, N12850, N12653);
xor XOR2 (N14084, N14081, N12233);
not NOT1 (N14085, N14070);
and AND4 (N14086, N14085, N11384, N8643, N2065);
buf BUF1 (N14087, N14082);
xor XOR2 (N14088, N14084, N10231);
nand NAND3 (N14089, N14083, N7961, N1231);
nand NAND2 (N14090, N14089, N11151);
and AND2 (N14091, N14076, N11789);
buf BUF1 (N14092, N14086);
xor XOR2 (N14093, N14057, N13110);
nor NOR2 (N14094, N14088, N4741);
not NOT1 (N14095, N14072);
nor NOR3 (N14096, N14090, N13403, N8855);
buf BUF1 (N14097, N14077);
and AND4 (N14098, N14093, N11303, N4707, N12198);
buf BUF1 (N14099, N14098);
and AND4 (N14100, N14099, N4914, N8635, N5576);
buf BUF1 (N14101, N14075);
xor XOR2 (N14102, N14091, N5296);
or OR2 (N14103, N14101, N4558);
nand NAND4 (N14104, N14096, N1461, N1049, N2742);
not NOT1 (N14105, N14094);
buf BUF1 (N14106, N14104);
not NOT1 (N14107, N14100);
buf BUF1 (N14108, N14106);
nor NOR3 (N14109, N14092, N888, N3921);
nand NAND3 (N14110, N14097, N890, N5068);
nor NOR2 (N14111, N14109, N10232);
nor NOR3 (N14112, N14102, N11420, N684);
or OR3 (N14113, N14105, N7113, N9351);
or OR2 (N14114, N14113, N13365);
buf BUF1 (N14115, N14080);
and AND3 (N14116, N14107, N8003, N4070);
nor NOR2 (N14117, N14108, N13408);
xor XOR2 (N14118, N14116, N12384);
nor NOR3 (N14119, N14118, N3675, N1433);
and AND2 (N14120, N14119, N4940);
xor XOR2 (N14121, N14112, N10031);
buf BUF1 (N14122, N14114);
xor XOR2 (N14123, N14111, N22);
not NOT1 (N14124, N14121);
nor NOR2 (N14125, N14110, N13444);
nor NOR4 (N14126, N14123, N4253, N459, N7907);
nor NOR2 (N14127, N14124, N1875);
not NOT1 (N14128, N14095);
not NOT1 (N14129, N14103);
and AND4 (N14130, N14120, N7611, N9706, N6169);
buf BUF1 (N14131, N14122);
not NOT1 (N14132, N14125);
not NOT1 (N14133, N14115);
not NOT1 (N14134, N14133);
and AND4 (N14135, N14131, N1953, N11787, N731);
and AND4 (N14136, N14135, N13295, N1288, N1538);
and AND2 (N14137, N14128, N12719);
nor NOR2 (N14138, N14117, N10814);
nand NAND4 (N14139, N14137, N14131, N6912, N10698);
buf BUF1 (N14140, N14138);
buf BUF1 (N14141, N14127);
nand NAND3 (N14142, N14087, N8177, N7214);
not NOT1 (N14143, N14130);
nand NAND4 (N14144, N14129, N3247, N4068, N10743);
nor NOR4 (N14145, N14143, N6498, N5210, N10691);
buf BUF1 (N14146, N14144);
xor XOR2 (N14147, N14134, N8001);
xor XOR2 (N14148, N14145, N2175);
not NOT1 (N14149, N14126);
or OR2 (N14150, N14148, N4183);
nand NAND2 (N14151, N14146, N10670);
and AND4 (N14152, N14142, N7039, N10062, N7048);
and AND2 (N14153, N14132, N4372);
not NOT1 (N14154, N14153);
nor NOR3 (N14155, N14149, N13378, N6520);
and AND2 (N14156, N14147, N5933);
or OR4 (N14157, N14136, N12878, N1988, N2578);
and AND4 (N14158, N14140, N410, N3040, N6251);
buf BUF1 (N14159, N14150);
nand NAND4 (N14160, N14141, N11685, N1957, N10028);
and AND3 (N14161, N14155, N10919, N13185);
nor NOR3 (N14162, N14154, N13504, N7623);
not NOT1 (N14163, N14157);
or OR3 (N14164, N14159, N13159, N7477);
or OR3 (N14165, N14156, N4190, N8850);
xor XOR2 (N14166, N14164, N6769);
nor NOR4 (N14167, N14161, N8236, N4571, N8692);
nor NOR3 (N14168, N14160, N12835, N4385);
nand NAND4 (N14169, N14162, N13231, N11448, N6908);
nand NAND4 (N14170, N14165, N10196, N12781, N11010);
or OR2 (N14171, N14163, N7990);
xor XOR2 (N14172, N14152, N7032);
nand NAND3 (N14173, N14167, N1809, N3548);
nor NOR2 (N14174, N14158, N4494);
nor NOR4 (N14175, N14170, N211, N10408, N3377);
nand NAND2 (N14176, N14171, N8744);
nand NAND3 (N14177, N14173, N6419, N5445);
or OR2 (N14178, N14177, N7079);
buf BUF1 (N14179, N14172);
not NOT1 (N14180, N14166);
buf BUF1 (N14181, N14139);
buf BUF1 (N14182, N14175);
and AND4 (N14183, N14151, N5501, N10169, N2360);
and AND2 (N14184, N14178, N1606);
not NOT1 (N14185, N14174);
nor NOR4 (N14186, N14184, N11259, N811, N10074);
nand NAND4 (N14187, N14186, N9652, N9592, N3031);
buf BUF1 (N14188, N14183);
not NOT1 (N14189, N14176);
buf BUF1 (N14190, N14182);
nand NAND2 (N14191, N14169, N4481);
and AND3 (N14192, N14185, N4305, N1685);
xor XOR2 (N14193, N14192, N13623);
and AND2 (N14194, N14179, N9095);
xor XOR2 (N14195, N14168, N1201);
and AND4 (N14196, N14191, N4260, N8480, N4332);
xor XOR2 (N14197, N14193, N8643);
or OR2 (N14198, N14181, N10341);
not NOT1 (N14199, N14198);
not NOT1 (N14200, N14194);
nor NOR2 (N14201, N14189, N497);
and AND2 (N14202, N14196, N11487);
not NOT1 (N14203, N14197);
nand NAND4 (N14204, N14195, N1657, N3572, N10418);
nand NAND2 (N14205, N14180, N10347);
nor NOR4 (N14206, N14204, N6150, N2387, N12243);
nor NOR4 (N14207, N14202, N5768, N5252, N10136);
nand NAND2 (N14208, N14201, N8571);
and AND3 (N14209, N14187, N5316, N1718);
not NOT1 (N14210, N14188);
or OR4 (N14211, N14206, N3794, N4270, N10070);
nand NAND4 (N14212, N14208, N538, N11165, N9127);
nor NOR3 (N14213, N14203, N9004, N1900);
nand NAND2 (N14214, N14200, N2750);
or OR2 (N14215, N14212, N10195);
not NOT1 (N14216, N14211);
nand NAND4 (N14217, N14199, N8686, N13037, N11768);
or OR2 (N14218, N14205, N142);
buf BUF1 (N14219, N14216);
not NOT1 (N14220, N14190);
or OR2 (N14221, N14219, N3304);
and AND3 (N14222, N14207, N7869, N6724);
not NOT1 (N14223, N14218);
buf BUF1 (N14224, N14222);
buf BUF1 (N14225, N14214);
nand NAND2 (N14226, N14224, N4620);
nand NAND3 (N14227, N14226, N3694, N10885);
not NOT1 (N14228, N14227);
not NOT1 (N14229, N14223);
nor NOR3 (N14230, N14228, N3095, N7944);
nor NOR2 (N14231, N14225, N6502);
nand NAND2 (N14232, N14210, N267);
nand NAND4 (N14233, N14230, N5939, N5976, N12541);
buf BUF1 (N14234, N14232);
and AND4 (N14235, N14217, N11915, N11178, N788);
buf BUF1 (N14236, N14234);
or OR2 (N14237, N14220, N1167);
and AND4 (N14238, N14237, N24, N7217, N10805);
nand NAND4 (N14239, N14231, N2206, N10136, N8);
nor NOR2 (N14240, N14233, N8519);
xor XOR2 (N14241, N14221, N9431);
or OR3 (N14242, N14213, N7723, N4358);
nand NAND2 (N14243, N14209, N11097);
or OR3 (N14244, N14235, N8722, N1152);
buf BUF1 (N14245, N14229);
nor NOR3 (N14246, N14241, N7306, N4813);
or OR2 (N14247, N14246, N2088);
xor XOR2 (N14248, N14247, N5277);
or OR4 (N14249, N14239, N861, N5455, N7898);
and AND3 (N14250, N14242, N11659, N4996);
not NOT1 (N14251, N14243);
xor XOR2 (N14252, N14245, N8093);
and AND4 (N14253, N14238, N2409, N1769, N13840);
and AND2 (N14254, N14240, N8769);
and AND4 (N14255, N14254, N12341, N13153, N4317);
buf BUF1 (N14256, N14255);
xor XOR2 (N14257, N14236, N13411);
not NOT1 (N14258, N14250);
or OR3 (N14259, N14248, N7602, N8329);
not NOT1 (N14260, N14252);
not NOT1 (N14261, N14260);
buf BUF1 (N14262, N14257);
xor XOR2 (N14263, N14251, N4825);
xor XOR2 (N14264, N14256, N12906);
or OR3 (N14265, N14253, N1329, N7062);
buf BUF1 (N14266, N14215);
or OR3 (N14267, N14265, N5459, N8425);
nand NAND3 (N14268, N14244, N11974, N6735);
and AND3 (N14269, N14266, N10260, N10890);
and AND3 (N14270, N14269, N1573, N10771);
and AND2 (N14271, N14262, N13805);
or OR4 (N14272, N14271, N14035, N6650, N12215);
or OR3 (N14273, N14267, N13339, N9349);
nand NAND3 (N14274, N14268, N3671, N1373);
xor XOR2 (N14275, N14273, N7620);
nand NAND4 (N14276, N14274, N4328, N5408, N6593);
or OR2 (N14277, N14259, N9506);
buf BUF1 (N14278, N14261);
or OR3 (N14279, N14278, N2821, N10837);
buf BUF1 (N14280, N14277);
or OR3 (N14281, N14264, N11402, N2982);
nor NOR4 (N14282, N14275, N13409, N6719, N10549);
or OR2 (N14283, N14258, N6892);
not NOT1 (N14284, N14276);
xor XOR2 (N14285, N14282, N3998);
nand NAND2 (N14286, N14281, N569);
nand NAND2 (N14287, N14283, N5871);
buf BUF1 (N14288, N14284);
xor XOR2 (N14289, N14263, N12110);
not NOT1 (N14290, N14280);
nand NAND3 (N14291, N14286, N4382, N16);
buf BUF1 (N14292, N14249);
nand NAND4 (N14293, N14288, N1252, N10525, N6952);
not NOT1 (N14294, N14279);
nand NAND2 (N14295, N14287, N6656);
xor XOR2 (N14296, N14294, N1428);
or OR4 (N14297, N14272, N1564, N11484, N574);
nand NAND2 (N14298, N14296, N1659);
nor NOR3 (N14299, N14285, N1551, N6920);
buf BUF1 (N14300, N14295);
and AND2 (N14301, N14297, N12951);
buf BUF1 (N14302, N14293);
nor NOR3 (N14303, N14298, N8532, N4435);
xor XOR2 (N14304, N14301, N11332);
and AND2 (N14305, N14270, N7808);
nor NOR3 (N14306, N14303, N471, N848);
xor XOR2 (N14307, N14300, N14298);
nand NAND2 (N14308, N14307, N4710);
buf BUF1 (N14309, N14302);
not NOT1 (N14310, N14289);
and AND4 (N14311, N14299, N3333, N5755, N12872);
nor NOR3 (N14312, N14309, N6992, N6308);
buf BUF1 (N14313, N14305);
nand NAND2 (N14314, N14308, N8801);
or OR3 (N14315, N14314, N421, N6867);
buf BUF1 (N14316, N14310);
nand NAND4 (N14317, N14312, N4103, N12414, N5833);
or OR3 (N14318, N14291, N11998, N8568);
nor NOR2 (N14319, N14317, N8257);
buf BUF1 (N14320, N14319);
and AND3 (N14321, N14304, N10534, N12117);
nor NOR2 (N14322, N14292, N6053);
buf BUF1 (N14323, N14290);
not NOT1 (N14324, N14306);
buf BUF1 (N14325, N14322);
xor XOR2 (N14326, N14316, N13689);
nor NOR3 (N14327, N14311, N8622, N1103);
nor NOR2 (N14328, N14315, N5221);
nor NOR2 (N14329, N14321, N4345);
nor NOR2 (N14330, N14324, N10060);
or OR2 (N14331, N14326, N10685);
buf BUF1 (N14332, N14330);
and AND2 (N14333, N14331, N5637);
nor NOR4 (N14334, N14328, N12836, N10680, N3361);
xor XOR2 (N14335, N14323, N4626);
buf BUF1 (N14336, N14329);
nor NOR2 (N14337, N14332, N8141);
buf BUF1 (N14338, N14325);
and AND2 (N14339, N14313, N8626);
nand NAND2 (N14340, N14318, N13542);
nand NAND2 (N14341, N14320, N11071);
nor NOR2 (N14342, N14340, N12466);
buf BUF1 (N14343, N14341);
xor XOR2 (N14344, N14339, N7046);
nand NAND4 (N14345, N14338, N10618, N208, N11856);
and AND4 (N14346, N14327, N11832, N14046, N11126);
or OR3 (N14347, N14345, N14140, N7614);
and AND2 (N14348, N14342, N8286);
xor XOR2 (N14349, N14336, N13606);
or OR2 (N14350, N14347, N13648);
xor XOR2 (N14351, N14344, N3283);
and AND3 (N14352, N14348, N9561, N6750);
and AND2 (N14353, N14335, N8469);
and AND3 (N14354, N14353, N8477, N12166);
or OR2 (N14355, N14337, N9937);
nor NOR4 (N14356, N14349, N12097, N9817, N6817);
nor NOR2 (N14357, N14356, N4960);
xor XOR2 (N14358, N14343, N5916);
nor NOR2 (N14359, N14351, N9501);
nor NOR4 (N14360, N14355, N11571, N7063, N6225);
and AND4 (N14361, N14354, N2180, N3025, N4078);
nand NAND3 (N14362, N14334, N1149, N11599);
nand NAND2 (N14363, N14352, N2204);
not NOT1 (N14364, N14360);
nand NAND2 (N14365, N14362, N12897);
nand NAND3 (N14366, N14350, N12119, N8099);
not NOT1 (N14367, N14361);
not NOT1 (N14368, N14367);
nor NOR3 (N14369, N14365, N8752, N1066);
nand NAND2 (N14370, N14333, N10135);
xor XOR2 (N14371, N14357, N734);
not NOT1 (N14372, N14369);
or OR2 (N14373, N14364, N12517);
buf BUF1 (N14374, N14368);
not NOT1 (N14375, N14359);
or OR2 (N14376, N14346, N9487);
and AND3 (N14377, N14366, N14282, N3371);
xor XOR2 (N14378, N14374, N12177);
buf BUF1 (N14379, N14373);
not NOT1 (N14380, N14358);
buf BUF1 (N14381, N14377);
not NOT1 (N14382, N14372);
and AND2 (N14383, N14380, N6174);
or OR4 (N14384, N14383, N7842, N1817, N2954);
or OR4 (N14385, N14379, N9683, N7186, N8228);
and AND3 (N14386, N14382, N495, N14181);
or OR3 (N14387, N14363, N12162, N5054);
and AND2 (N14388, N14386, N8379);
nand NAND4 (N14389, N14388, N4379, N5249, N6343);
xor XOR2 (N14390, N14378, N12438);
or OR3 (N14391, N14375, N7203, N6701);
buf BUF1 (N14392, N14387);
nand NAND3 (N14393, N14384, N10218, N4305);
xor XOR2 (N14394, N14376, N6776);
and AND4 (N14395, N14381, N12942, N11843, N2662);
xor XOR2 (N14396, N14370, N5728);
xor XOR2 (N14397, N14391, N8145);
or OR3 (N14398, N14397, N13608, N4354);
or OR2 (N14399, N14396, N14058);
or OR4 (N14400, N14385, N3425, N598, N2257);
nor NOR3 (N14401, N14389, N12571, N9515);
not NOT1 (N14402, N14371);
and AND3 (N14403, N14392, N13733, N9572);
and AND4 (N14404, N14395, N11354, N12171, N11781);
nand NAND3 (N14405, N14399, N13425, N287);
and AND2 (N14406, N14400, N3200);
xor XOR2 (N14407, N14401, N664);
nor NOR3 (N14408, N14393, N922, N1588);
xor XOR2 (N14409, N14407, N11875);
buf BUF1 (N14410, N14398);
not NOT1 (N14411, N14403);
nand NAND3 (N14412, N14390, N3230, N13950);
buf BUF1 (N14413, N14402);
buf BUF1 (N14414, N14413);
or OR4 (N14415, N14414, N10954, N2622, N9741);
xor XOR2 (N14416, N14410, N6173);
nand NAND4 (N14417, N14394, N13243, N1797, N12989);
not NOT1 (N14418, N14412);
nor NOR3 (N14419, N14411, N2998, N8330);
and AND4 (N14420, N14406, N7013, N11643, N9581);
xor XOR2 (N14421, N14416, N12630);
nand NAND2 (N14422, N14421, N14381);
nor NOR2 (N14423, N14419, N7112);
xor XOR2 (N14424, N14409, N11318);
not NOT1 (N14425, N14417);
xor XOR2 (N14426, N14408, N7430);
or OR3 (N14427, N14422, N1744, N2504);
not NOT1 (N14428, N14425);
and AND4 (N14429, N14428, N2721, N7274, N12725);
and AND3 (N14430, N14426, N11186, N8966);
or OR4 (N14431, N14423, N1917, N8814, N11776);
and AND2 (N14432, N14431, N9766);
buf BUF1 (N14433, N14427);
not NOT1 (N14434, N14429);
nor NOR2 (N14435, N14415, N3421);
and AND2 (N14436, N14434, N3261);
not NOT1 (N14437, N14433);
nor NOR4 (N14438, N14424, N5332, N9002, N11290);
buf BUF1 (N14439, N14405);
nor NOR4 (N14440, N14437, N3134, N10159, N7462);
nor NOR3 (N14441, N14436, N10874, N11605);
nand NAND2 (N14442, N14438, N7854);
not NOT1 (N14443, N14420);
xor XOR2 (N14444, N14432, N11912);
nor NOR2 (N14445, N14440, N12404);
or OR3 (N14446, N14435, N11079, N9190);
xor XOR2 (N14447, N14444, N5755);
or OR2 (N14448, N14439, N1142);
xor XOR2 (N14449, N14441, N4953);
xor XOR2 (N14450, N14418, N12607);
xor XOR2 (N14451, N14404, N5567);
nand NAND2 (N14452, N14446, N14162);
nor NOR3 (N14453, N14448, N5467, N2982);
or OR2 (N14454, N14451, N65);
nor NOR4 (N14455, N14430, N3658, N9145, N6762);
not NOT1 (N14456, N14443);
or OR4 (N14457, N14453, N14378, N10688, N7096);
not NOT1 (N14458, N14449);
or OR4 (N14459, N14452, N3616, N8877, N14144);
or OR3 (N14460, N14457, N13634, N10753);
buf BUF1 (N14461, N14450);
and AND3 (N14462, N14447, N12228, N12327);
nand NAND2 (N14463, N14455, N8805);
nor NOR2 (N14464, N14461, N6792);
nor NOR3 (N14465, N14458, N9611, N4663);
nand NAND4 (N14466, N14465, N11405, N7061, N9151);
not NOT1 (N14467, N14460);
or OR3 (N14468, N14463, N7789, N7443);
nand NAND3 (N14469, N14466, N9223, N20);
not NOT1 (N14470, N14454);
not NOT1 (N14471, N14442);
nand NAND4 (N14472, N14469, N13670, N829, N12621);
xor XOR2 (N14473, N14464, N6114);
xor XOR2 (N14474, N14467, N9661);
or OR4 (N14475, N14456, N556, N3405, N7750);
nor NOR3 (N14476, N14468, N990, N7929);
or OR4 (N14477, N14475, N8163, N14455, N6117);
xor XOR2 (N14478, N14445, N10645);
nand NAND4 (N14479, N14470, N8577, N14299, N4417);
xor XOR2 (N14480, N14477, N5037);
and AND2 (N14481, N14459, N9563);
or OR4 (N14482, N14462, N2438, N2222, N10754);
buf BUF1 (N14483, N14476);
buf BUF1 (N14484, N14473);
and AND2 (N14485, N14472, N10527);
and AND3 (N14486, N14485, N2892, N9558);
and AND2 (N14487, N14474, N14390);
buf BUF1 (N14488, N14486);
and AND3 (N14489, N14484, N2932, N12567);
and AND2 (N14490, N14480, N4104);
not NOT1 (N14491, N14487);
and AND3 (N14492, N14483, N11694, N5879);
or OR3 (N14493, N14479, N1155, N11219);
not NOT1 (N14494, N14471);
nor NOR2 (N14495, N14490, N11121);
buf BUF1 (N14496, N14489);
buf BUF1 (N14497, N14478);
not NOT1 (N14498, N14491);
buf BUF1 (N14499, N14497);
buf BUF1 (N14500, N14481);
nand NAND3 (N14501, N14482, N13056, N8675);
nand NAND2 (N14502, N14493, N13405);
nand NAND3 (N14503, N14498, N5755, N11958);
or OR4 (N14504, N14492, N4122, N3251, N7760);
buf BUF1 (N14505, N14488);
nand NAND2 (N14506, N14504, N6489);
xor XOR2 (N14507, N14505, N1443);
nand NAND3 (N14508, N14494, N7501, N6613);
nand NAND4 (N14509, N14507, N13117, N2626, N6144);
buf BUF1 (N14510, N14500);
nor NOR3 (N14511, N14502, N4922, N3670);
and AND2 (N14512, N14495, N8375);
not NOT1 (N14513, N14512);
not NOT1 (N14514, N14511);
nor NOR2 (N14515, N14501, N5632);
not NOT1 (N14516, N14499);
or OR2 (N14517, N14503, N7297);
nand NAND3 (N14518, N14514, N1471, N2794);
xor XOR2 (N14519, N14510, N10549);
xor XOR2 (N14520, N14515, N1600);
xor XOR2 (N14521, N14496, N6891);
or OR3 (N14522, N14517, N9349, N6370);
buf BUF1 (N14523, N14506);
nand NAND3 (N14524, N14508, N1932, N8338);
nor NOR2 (N14525, N14522, N2959);
not NOT1 (N14526, N14520);
or OR2 (N14527, N14518, N12464);
nor NOR3 (N14528, N14527, N2193, N11279);
buf BUF1 (N14529, N14523);
not NOT1 (N14530, N14513);
xor XOR2 (N14531, N14521, N4672);
or OR3 (N14532, N14529, N11794, N5100);
buf BUF1 (N14533, N14526);
not NOT1 (N14534, N14528);
buf BUF1 (N14535, N14516);
not NOT1 (N14536, N14531);
or OR4 (N14537, N14535, N910, N9101, N7579);
not NOT1 (N14538, N14537);
nand NAND3 (N14539, N14534, N6806, N12718);
xor XOR2 (N14540, N14538, N2281);
nand NAND4 (N14541, N14525, N6357, N4123, N12340);
nand NAND2 (N14542, N14532, N10352);
nor NOR4 (N14543, N14530, N10845, N2057, N265);
or OR4 (N14544, N14543, N5794, N4324, N1344);
nor NOR3 (N14545, N14544, N2541, N12619);
or OR4 (N14546, N14539, N5992, N9489, N5017);
or OR3 (N14547, N14542, N144, N7783);
not NOT1 (N14548, N14540);
xor XOR2 (N14549, N14524, N5798);
nor NOR4 (N14550, N14548, N8057, N7276, N14412);
and AND3 (N14551, N14536, N9942, N7648);
buf BUF1 (N14552, N14550);
or OR3 (N14553, N14551, N7497, N148);
xor XOR2 (N14554, N14541, N6636);
buf BUF1 (N14555, N14552);
nor NOR3 (N14556, N14549, N139, N8770);
xor XOR2 (N14557, N14533, N4870);
nor NOR3 (N14558, N14519, N12879, N217);
nor NOR4 (N14559, N14554, N6279, N4636, N1531);
or OR3 (N14560, N14555, N476, N176);
not NOT1 (N14561, N14556);
or OR3 (N14562, N14545, N3035, N3849);
buf BUF1 (N14563, N14547);
xor XOR2 (N14564, N14563, N12928);
and AND2 (N14565, N14558, N5027);
not NOT1 (N14566, N14559);
or OR4 (N14567, N14562, N8601, N12688, N14057);
nor NOR3 (N14568, N14561, N12560, N13695);
or OR2 (N14569, N14564, N13189);
nor NOR3 (N14570, N14569, N9640, N1943);
or OR3 (N14571, N14570, N10941, N9521);
not NOT1 (N14572, N14568);
buf BUF1 (N14573, N14509);
and AND2 (N14574, N14572, N1657);
not NOT1 (N14575, N14566);
xor XOR2 (N14576, N14560, N9110);
or OR2 (N14577, N14576, N10955);
buf BUF1 (N14578, N14574);
nand NAND3 (N14579, N14565, N10916, N3407);
xor XOR2 (N14580, N14577, N6306);
buf BUF1 (N14581, N14580);
buf BUF1 (N14582, N14546);
nand NAND4 (N14583, N14582, N2847, N12884, N5193);
buf BUF1 (N14584, N14578);
or OR3 (N14585, N14571, N10314, N3046);
buf BUF1 (N14586, N14553);
or OR3 (N14587, N14586, N1216, N6880);
and AND2 (N14588, N14585, N10970);
and AND4 (N14589, N14581, N4302, N5906, N3483);
xor XOR2 (N14590, N14589, N13216);
nor NOR3 (N14591, N14584, N9859, N4722);
nand NAND2 (N14592, N14579, N11972);
xor XOR2 (N14593, N14557, N402);
nor NOR4 (N14594, N14587, N10720, N1983, N3524);
nand NAND2 (N14595, N14594, N508);
nand NAND3 (N14596, N14590, N2890, N5552);
not NOT1 (N14597, N14575);
nand NAND2 (N14598, N14595, N13225);
nor NOR4 (N14599, N14592, N14273, N135, N7232);
nor NOR2 (N14600, N14596, N11662);
nor NOR4 (N14601, N14591, N9076, N165, N6274);
not NOT1 (N14602, N14593);
not NOT1 (N14603, N14588);
nand NAND2 (N14604, N14601, N11091);
or OR3 (N14605, N14604, N3008, N10276);
or OR2 (N14606, N14602, N8167);
xor XOR2 (N14607, N14583, N12146);
nor NOR2 (N14608, N14606, N3021);
xor XOR2 (N14609, N14599, N3017);
or OR2 (N14610, N14567, N5868);
xor XOR2 (N14611, N14598, N4202);
nor NOR3 (N14612, N14611, N1928, N12754);
or OR2 (N14613, N14609, N12714);
nor NOR3 (N14614, N14608, N7018, N12978);
nand NAND3 (N14615, N14605, N7849, N12054);
buf BUF1 (N14616, N14573);
or OR4 (N14617, N14610, N5507, N10021, N3878);
nor NOR3 (N14618, N14600, N4927, N10600);
not NOT1 (N14619, N14597);
buf BUF1 (N14620, N14619);
not NOT1 (N14621, N14616);
and AND3 (N14622, N14621, N11310, N3181);
buf BUF1 (N14623, N14613);
not NOT1 (N14624, N14607);
buf BUF1 (N14625, N14623);
not NOT1 (N14626, N14624);
nand NAND2 (N14627, N14622, N7469);
xor XOR2 (N14628, N14618, N14240);
or OR4 (N14629, N14612, N3939, N10411, N2938);
or OR2 (N14630, N14615, N5202);
xor XOR2 (N14631, N14629, N12621);
nor NOR3 (N14632, N14628, N5734, N6512);
xor XOR2 (N14633, N14614, N13413);
buf BUF1 (N14634, N14631);
nor NOR4 (N14635, N14633, N8509, N12068, N13279);
not NOT1 (N14636, N14617);
nand NAND2 (N14637, N14626, N2639);
and AND2 (N14638, N14620, N1820);
nand NAND3 (N14639, N14603, N6884, N2571);
xor XOR2 (N14640, N14635, N5922);
or OR3 (N14641, N14640, N12336, N2377);
buf BUF1 (N14642, N14632);
buf BUF1 (N14643, N14630);
buf BUF1 (N14644, N14642);
xor XOR2 (N14645, N14638, N11727);
xor XOR2 (N14646, N14639, N10439);
nor NOR3 (N14647, N14627, N10200, N32);
and AND2 (N14648, N14636, N5762);
or OR2 (N14649, N14643, N6881);
not NOT1 (N14650, N14648);
buf BUF1 (N14651, N14647);
buf BUF1 (N14652, N14634);
buf BUF1 (N14653, N14637);
or OR3 (N14654, N14651, N13146, N2924);
or OR3 (N14655, N14654, N7522, N10225);
nor NOR3 (N14656, N14644, N1955, N7730);
nand NAND3 (N14657, N14652, N3081, N13111);
or OR2 (N14658, N14649, N10423);
xor XOR2 (N14659, N14645, N13886);
or OR2 (N14660, N14646, N10229);
nand NAND2 (N14661, N14656, N6943);
nor NOR2 (N14662, N14659, N4099);
buf BUF1 (N14663, N14658);
buf BUF1 (N14664, N14655);
xor XOR2 (N14665, N14625, N10929);
nor NOR4 (N14666, N14662, N3779, N7148, N10102);
buf BUF1 (N14667, N14666);
not NOT1 (N14668, N14664);
nand NAND4 (N14669, N14660, N3124, N1431, N10889);
nor NOR4 (N14670, N14668, N2544, N1486, N4378);
not NOT1 (N14671, N14653);
nor NOR2 (N14672, N14661, N4684);
or OR4 (N14673, N14663, N2268, N13130, N753);
or OR2 (N14674, N14667, N1456);
buf BUF1 (N14675, N14650);
and AND2 (N14676, N14671, N9806);
nor NOR3 (N14677, N14641, N2246, N8137);
nor NOR4 (N14678, N14673, N10056, N14452, N8467);
buf BUF1 (N14679, N14669);
xor XOR2 (N14680, N14672, N10368);
not NOT1 (N14681, N14675);
or OR4 (N14682, N14677, N1282, N10887, N14524);
nor NOR2 (N14683, N14680, N10519);
and AND2 (N14684, N14657, N8648);
buf BUF1 (N14685, N14681);
xor XOR2 (N14686, N14674, N3465);
or OR2 (N14687, N14679, N8932);
buf BUF1 (N14688, N14687);
buf BUF1 (N14689, N14670);
buf BUF1 (N14690, N14688);
or OR2 (N14691, N14689, N8763);
or OR2 (N14692, N14682, N1553);
and AND2 (N14693, N14685, N13863);
nor NOR2 (N14694, N14690, N11813);
and AND4 (N14695, N14686, N11544, N2555, N9491);
nand NAND3 (N14696, N14693, N6554, N6008);
buf BUF1 (N14697, N14665);
nand NAND2 (N14698, N14695, N14425);
xor XOR2 (N14699, N14678, N10373);
nand NAND4 (N14700, N14691, N5495, N8421, N8517);
buf BUF1 (N14701, N14676);
and AND2 (N14702, N14683, N13246);
nand NAND3 (N14703, N14700, N14588, N2179);
nand NAND3 (N14704, N14702, N14182, N11435);
nor NOR2 (N14705, N14703, N14271);
nand NAND2 (N14706, N14698, N4803);
or OR4 (N14707, N14692, N1834, N14236, N5369);
and AND4 (N14708, N14697, N6520, N1958, N13777);
not NOT1 (N14709, N14701);
and AND3 (N14710, N14707, N4795, N9933);
nand NAND2 (N14711, N14708, N1821);
or OR3 (N14712, N14710, N2199, N10610);
nand NAND4 (N14713, N14711, N5770, N4556, N3539);
not NOT1 (N14714, N14699);
nand NAND2 (N14715, N14696, N163);
nand NAND3 (N14716, N14706, N7433, N12772);
nand NAND4 (N14717, N14712, N10117, N10923, N335);
buf BUF1 (N14718, N14709);
and AND4 (N14719, N14717, N914, N4213, N9552);
and AND2 (N14720, N14705, N9847);
or OR3 (N14721, N14715, N5989, N4102);
buf BUF1 (N14722, N14694);
xor XOR2 (N14723, N14714, N14244);
not NOT1 (N14724, N14720);
xor XOR2 (N14725, N14724, N7366);
or OR2 (N14726, N14684, N952);
xor XOR2 (N14727, N14722, N3110);
nand NAND2 (N14728, N14704, N12328);
nor NOR3 (N14729, N14723, N10766, N5501);
buf BUF1 (N14730, N14726);
nand NAND4 (N14731, N14727, N5464, N1916, N4853);
and AND4 (N14732, N14721, N13685, N11202, N11482);
and AND4 (N14733, N14725, N5476, N11018, N3675);
nor NOR2 (N14734, N14718, N2788);
nand NAND2 (N14735, N14728, N1058);
nand NAND4 (N14736, N14735, N5768, N11896, N1859);
not NOT1 (N14737, N14733);
nand NAND2 (N14738, N14734, N7533);
xor XOR2 (N14739, N14732, N1227);
not NOT1 (N14740, N14736);
and AND4 (N14741, N14719, N11976, N11882, N11642);
xor XOR2 (N14742, N14737, N8483);
xor XOR2 (N14743, N14731, N6566);
not NOT1 (N14744, N14716);
nand NAND2 (N14745, N14730, N6319);
nor NOR3 (N14746, N14729, N14221, N8821);
not NOT1 (N14747, N14741);
xor XOR2 (N14748, N14745, N4268);
xor XOR2 (N14749, N14746, N14388);
not NOT1 (N14750, N14740);
nand NAND4 (N14751, N14742, N543, N1443, N12300);
nor NOR3 (N14752, N14748, N11214, N13578);
and AND4 (N14753, N14750, N413, N9330, N11841);
nor NOR2 (N14754, N14747, N5300);
or OR3 (N14755, N14749, N9180, N11521);
buf BUF1 (N14756, N14751);
nand NAND3 (N14757, N14713, N9162, N5559);
or OR4 (N14758, N14739, N14131, N13827, N2395);
and AND3 (N14759, N14744, N11702, N13706);
buf BUF1 (N14760, N14756);
xor XOR2 (N14761, N14738, N10802);
not NOT1 (N14762, N14760);
or OR4 (N14763, N14761, N14599, N8720, N4543);
nand NAND4 (N14764, N14763, N4261, N2578, N4375);
nor NOR4 (N14765, N14758, N2498, N11469, N6880);
nand NAND2 (N14766, N14755, N161);
nand NAND3 (N14767, N14743, N6327, N4053);
not NOT1 (N14768, N14762);
not NOT1 (N14769, N14759);
xor XOR2 (N14770, N14752, N11543);
buf BUF1 (N14771, N14754);
or OR3 (N14772, N14765, N7032, N12259);
nand NAND4 (N14773, N14768, N2737, N3486, N6578);
buf BUF1 (N14774, N14753);
or OR3 (N14775, N14769, N12938, N13166);
xor XOR2 (N14776, N14773, N2599);
nor NOR4 (N14777, N14771, N11314, N14059, N2568);
or OR4 (N14778, N14770, N680, N12966, N5350);
or OR3 (N14779, N14764, N3946, N13180);
xor XOR2 (N14780, N14776, N1926);
and AND2 (N14781, N14780, N3460);
not NOT1 (N14782, N14777);
and AND2 (N14783, N14767, N11887);
buf BUF1 (N14784, N14782);
and AND4 (N14785, N14774, N4857, N7785, N11037);
nor NOR3 (N14786, N14778, N3160, N5672);
xor XOR2 (N14787, N14775, N13230);
xor XOR2 (N14788, N14781, N8573);
not NOT1 (N14789, N14779);
or OR3 (N14790, N14783, N12959, N7195);
and AND4 (N14791, N14789, N1349, N2612, N13106);
nand NAND3 (N14792, N14766, N1803, N3003);
or OR3 (N14793, N14786, N6350, N12680);
nor NOR4 (N14794, N14788, N11819, N1510, N6151);
nor NOR3 (N14795, N14793, N5282, N6037);
nor NOR4 (N14796, N14790, N8045, N6731, N345);
and AND2 (N14797, N14787, N2475);
xor XOR2 (N14798, N14791, N6378);
xor XOR2 (N14799, N14795, N7278);
and AND3 (N14800, N14796, N5528, N10146);
buf BUF1 (N14801, N14772);
xor XOR2 (N14802, N14792, N711);
or OR3 (N14803, N14797, N5387, N1202);
buf BUF1 (N14804, N14799);
not NOT1 (N14805, N14801);
buf BUF1 (N14806, N14805);
nand NAND2 (N14807, N14803, N14734);
xor XOR2 (N14808, N14807, N3000);
not NOT1 (N14809, N14808);
nand NAND2 (N14810, N14806, N293);
buf BUF1 (N14811, N14809);
not NOT1 (N14812, N14800);
not NOT1 (N14813, N14785);
nand NAND2 (N14814, N14811, N1272);
not NOT1 (N14815, N14810);
and AND3 (N14816, N14814, N7540, N10372);
nor NOR4 (N14817, N14757, N14217, N3906, N7360);
not NOT1 (N14818, N14813);
buf BUF1 (N14819, N14794);
buf BUF1 (N14820, N14815);
or OR3 (N14821, N14818, N5330, N3424);
or OR2 (N14822, N14819, N13105);
nor NOR3 (N14823, N14821, N2926, N13569);
and AND4 (N14824, N14804, N4945, N3322, N13209);
or OR2 (N14825, N14798, N9853);
and AND3 (N14826, N14825, N2384, N9271);
nand NAND2 (N14827, N14823, N5778);
nor NOR4 (N14828, N14826, N5125, N11625, N12552);
or OR3 (N14829, N14828, N6003, N129);
xor XOR2 (N14830, N14817, N922);
buf BUF1 (N14831, N14824);
not NOT1 (N14832, N14827);
nand NAND3 (N14833, N14816, N4590, N3252);
xor XOR2 (N14834, N14833, N5130);
nand NAND3 (N14835, N14820, N9800, N2669);
nor NOR4 (N14836, N14812, N8719, N1160, N6979);
buf BUF1 (N14837, N14836);
or OR4 (N14838, N14832, N5460, N14485, N2670);
or OR3 (N14839, N14837, N6309, N616);
or OR2 (N14840, N14838, N3531);
buf BUF1 (N14841, N14784);
or OR3 (N14842, N14839, N11713, N8140);
xor XOR2 (N14843, N14841, N8124);
and AND3 (N14844, N14822, N6247, N5526);
or OR3 (N14845, N14829, N11645, N14525);
xor XOR2 (N14846, N14844, N9160);
not NOT1 (N14847, N14831);
nor NOR3 (N14848, N14835, N9368, N8623);
not NOT1 (N14849, N14842);
not NOT1 (N14850, N14840);
or OR3 (N14851, N14834, N8821, N2214);
buf BUF1 (N14852, N14830);
and AND2 (N14853, N14849, N4115);
nand NAND3 (N14854, N14802, N9322, N13939);
buf BUF1 (N14855, N14845);
not NOT1 (N14856, N14853);
not NOT1 (N14857, N14854);
and AND3 (N14858, N14852, N4576, N1657);
not NOT1 (N14859, N14846);
and AND3 (N14860, N14851, N11607, N6003);
nand NAND4 (N14861, N14860, N6966, N1065, N7237);
not NOT1 (N14862, N14855);
nand NAND3 (N14863, N14843, N394, N14421);
nor NOR2 (N14864, N14863, N6467);
not NOT1 (N14865, N14847);
not NOT1 (N14866, N14864);
nand NAND4 (N14867, N14865, N7134, N11095, N8282);
xor XOR2 (N14868, N14862, N4422);
or OR3 (N14869, N14850, N13557, N14581);
buf BUF1 (N14870, N14848);
nor NOR2 (N14871, N14866, N5641);
xor XOR2 (N14872, N14856, N12677);
and AND3 (N14873, N14872, N6766, N2050);
or OR4 (N14874, N14857, N14387, N9923, N1399);
buf BUF1 (N14875, N14861);
nand NAND2 (N14876, N14871, N1160);
buf BUF1 (N14877, N14858);
and AND3 (N14878, N14873, N10349, N3822);
and AND3 (N14879, N14875, N8571, N8915);
or OR4 (N14880, N14879, N6601, N6004, N14823);
buf BUF1 (N14881, N14859);
xor XOR2 (N14882, N14868, N6156);
nand NAND4 (N14883, N14881, N9938, N3953, N2111);
not NOT1 (N14884, N14870);
xor XOR2 (N14885, N14877, N11922);
or OR2 (N14886, N14867, N11469);
or OR4 (N14887, N14880, N10987, N6446, N5299);
buf BUF1 (N14888, N14886);
or OR4 (N14889, N14887, N2401, N14848, N1863);
buf BUF1 (N14890, N14878);
xor XOR2 (N14891, N14876, N13472);
not NOT1 (N14892, N14888);
xor XOR2 (N14893, N14882, N11870);
nor NOR4 (N14894, N14883, N1592, N4985, N2645);
xor XOR2 (N14895, N14889, N13271);
nor NOR4 (N14896, N14892, N7962, N2651, N1124);
or OR4 (N14897, N14894, N3633, N458, N1121);
nor NOR3 (N14898, N14891, N1258, N10124);
xor XOR2 (N14899, N14893, N11438);
xor XOR2 (N14900, N14899, N11372);
nand NAND4 (N14901, N14900, N12803, N5667, N9393);
nand NAND2 (N14902, N14869, N13713);
nand NAND4 (N14903, N14898, N5072, N8115, N7908);
or OR3 (N14904, N14896, N1173, N6739);
not NOT1 (N14905, N14885);
or OR4 (N14906, N14903, N8015, N5327, N11640);
buf BUF1 (N14907, N14895);
not NOT1 (N14908, N14902);
not NOT1 (N14909, N14874);
buf BUF1 (N14910, N14904);
xor XOR2 (N14911, N14890, N7830);
or OR4 (N14912, N14884, N13551, N9724, N6261);
not NOT1 (N14913, N14911);
not NOT1 (N14914, N14909);
xor XOR2 (N14915, N14901, N7062);
nor NOR3 (N14916, N14905, N2641, N1309);
xor XOR2 (N14917, N14913, N10700);
or OR4 (N14918, N14910, N11871, N10331, N10584);
or OR3 (N14919, N14906, N1913, N2856);
xor XOR2 (N14920, N14917, N4543);
not NOT1 (N14921, N14897);
and AND3 (N14922, N14908, N9074, N3663);
nand NAND2 (N14923, N14907, N9498);
nand NAND3 (N14924, N14912, N1721, N11607);
or OR2 (N14925, N14923, N13518);
xor XOR2 (N14926, N14918, N11050);
nand NAND3 (N14927, N14922, N12944, N14779);
buf BUF1 (N14928, N14916);
nand NAND2 (N14929, N14915, N2483);
or OR4 (N14930, N14924, N340, N3410, N141);
and AND3 (N14931, N14927, N6928, N12838);
not NOT1 (N14932, N14925);
buf BUF1 (N14933, N14919);
not NOT1 (N14934, N14929);
nor NOR3 (N14935, N14930, N12030, N8540);
not NOT1 (N14936, N14935);
or OR3 (N14937, N14933, N1084, N11791);
not NOT1 (N14938, N14934);
or OR4 (N14939, N14936, N3939, N9311, N290);
nor NOR3 (N14940, N14926, N7478, N11982);
nand NAND3 (N14941, N14938, N898, N10934);
nand NAND4 (N14942, N14941, N5126, N8805, N7340);
nand NAND4 (N14943, N14939, N13460, N6932, N13926);
and AND2 (N14944, N14931, N3460);
nor NOR4 (N14945, N14914, N6496, N1470, N5381);
buf BUF1 (N14946, N14945);
nand NAND4 (N14947, N14937, N11151, N11970, N11702);
nor NOR3 (N14948, N14928, N10543, N8844);
or OR2 (N14949, N14920, N14814);
buf BUF1 (N14950, N14921);
and AND4 (N14951, N14942, N9639, N13704, N7912);
or OR3 (N14952, N14949, N3416, N13981);
nor NOR2 (N14953, N14940, N11427);
or OR3 (N14954, N14932, N3379, N7183);
xor XOR2 (N14955, N14951, N14035);
buf BUF1 (N14956, N14953);
buf BUF1 (N14957, N14947);
and AND2 (N14958, N14946, N10510);
buf BUF1 (N14959, N14957);
and AND4 (N14960, N14952, N5890, N7262, N5983);
nand NAND3 (N14961, N14950, N698, N2687);
buf BUF1 (N14962, N14959);
buf BUF1 (N14963, N14958);
nand NAND2 (N14964, N14948, N14456);
not NOT1 (N14965, N14956);
not NOT1 (N14966, N14954);
or OR4 (N14967, N14964, N4655, N5621, N7054);
or OR4 (N14968, N14966, N4949, N1395, N10399);
or OR2 (N14969, N14955, N4862);
not NOT1 (N14970, N14944);
xor XOR2 (N14971, N14963, N110);
and AND2 (N14972, N14960, N6145);
xor XOR2 (N14973, N14972, N3392);
buf BUF1 (N14974, N14969);
nand NAND3 (N14975, N14943, N2847, N10566);
not NOT1 (N14976, N14970);
or OR4 (N14977, N14962, N7627, N7071, N334);
or OR3 (N14978, N14967, N11, N6686);
buf BUF1 (N14979, N14977);
buf BUF1 (N14980, N14978);
nand NAND2 (N14981, N14973, N10549);
not NOT1 (N14982, N14975);
or OR3 (N14983, N14979, N8895, N6800);
and AND4 (N14984, N14974, N10765, N3629, N10);
not NOT1 (N14985, N14982);
buf BUF1 (N14986, N14983);
and AND2 (N14987, N14965, N5507);
nor NOR2 (N14988, N14971, N12276);
or OR4 (N14989, N14988, N4080, N5627, N11497);
and AND3 (N14990, N14976, N529, N8383);
and AND3 (N14991, N14989, N6740, N7119);
and AND4 (N14992, N14980, N5770, N12628, N4110);
nor NOR4 (N14993, N14968, N14169, N12754, N6017);
xor XOR2 (N14994, N14991, N9075);
and AND2 (N14995, N14994, N6472);
nor NOR3 (N14996, N14961, N10070, N13477);
and AND4 (N14997, N14985, N7677, N10826, N5867);
nor NOR3 (N14998, N14997, N12796, N6101);
nand NAND2 (N14999, N14996, N10801);
xor XOR2 (N15000, N14995, N10855);
not NOT1 (N15001, N14984);
nor NOR3 (N15002, N14992, N5733, N5063);
buf BUF1 (N15003, N14999);
nor NOR3 (N15004, N14993, N3523, N5620);
xor XOR2 (N15005, N15001, N4166);
xor XOR2 (N15006, N15003, N1169);
nor NOR3 (N15007, N14986, N4025, N9492);
nand NAND2 (N15008, N14990, N7156);
nor NOR3 (N15009, N15006, N2476, N6384);
xor XOR2 (N15010, N15009, N10798);
not NOT1 (N15011, N14981);
nor NOR3 (N15012, N14998, N12764, N5027);
and AND4 (N15013, N15008, N4998, N7535, N14763);
and AND4 (N15014, N15005, N3541, N13022, N2850);
xor XOR2 (N15015, N15002, N9338);
xor XOR2 (N15016, N15004, N1063);
nor NOR4 (N15017, N15015, N7669, N6933, N10921);
not NOT1 (N15018, N15010);
not NOT1 (N15019, N15012);
not NOT1 (N15020, N15011);
nor NOR2 (N15021, N14987, N5725);
not NOT1 (N15022, N15018);
buf BUF1 (N15023, N15014);
nand NAND3 (N15024, N15019, N14448, N12940);
nor NOR3 (N15025, N15020, N6841, N13490);
not NOT1 (N15026, N15024);
and AND2 (N15027, N15016, N11610);
nand NAND3 (N15028, N15026, N2275, N6800);
or OR2 (N15029, N15017, N13853);
xor XOR2 (N15030, N15025, N12905);
nand NAND2 (N15031, N15013, N8567);
not NOT1 (N15032, N15022);
nor NOR3 (N15033, N15029, N14344, N9095);
or OR4 (N15034, N15000, N4186, N3406, N8160);
not NOT1 (N15035, N15028);
buf BUF1 (N15036, N15034);
nor NOR2 (N15037, N15035, N4946);
xor XOR2 (N15038, N15021, N5350);
and AND4 (N15039, N15007, N10232, N8581, N4013);
nor NOR2 (N15040, N15038, N1835);
or OR2 (N15041, N15039, N3126);
nand NAND4 (N15042, N15031, N4957, N8006, N11453);
and AND3 (N15043, N15037, N2670, N5013);
or OR4 (N15044, N15036, N6389, N7864, N9202);
xor XOR2 (N15045, N15023, N4724);
not NOT1 (N15046, N15042);
nor NOR2 (N15047, N15033, N11402);
and AND3 (N15048, N15046, N2238, N6985);
not NOT1 (N15049, N15044);
nor NOR4 (N15050, N15047, N9741, N10873, N14408);
nor NOR3 (N15051, N15027, N4261, N4491);
xor XOR2 (N15052, N15048, N5092);
nand NAND3 (N15053, N15032, N2892, N4419);
or OR2 (N15054, N15045, N10155);
nand NAND3 (N15055, N15030, N4377, N4305);
xor XOR2 (N15056, N15055, N80);
nand NAND2 (N15057, N15054, N5144);
nor NOR3 (N15058, N15040, N2087, N1553);
not NOT1 (N15059, N15052);
nand NAND3 (N15060, N15053, N7420, N1358);
buf BUF1 (N15061, N15043);
not NOT1 (N15062, N15041);
and AND2 (N15063, N15051, N5175);
and AND2 (N15064, N15059, N8682);
nand NAND4 (N15065, N15063, N7847, N12380, N12791);
nand NAND3 (N15066, N15065, N14618, N9798);
and AND3 (N15067, N15061, N7674, N3502);
nand NAND4 (N15068, N15066, N3484, N8599, N10433);
nand NAND4 (N15069, N15060, N7289, N14046, N14699);
nand NAND4 (N15070, N15064, N5165, N5600, N13390);
and AND4 (N15071, N15067, N5267, N13978, N6672);
nand NAND2 (N15072, N15049, N3048);
buf BUF1 (N15073, N15050);
buf BUF1 (N15074, N15058);
buf BUF1 (N15075, N15056);
and AND4 (N15076, N15062, N5375, N4526, N10801);
or OR3 (N15077, N15068, N13701, N7565);
xor XOR2 (N15078, N15073, N3694);
or OR2 (N15079, N15057, N7084);
xor XOR2 (N15080, N15071, N12709);
nor NOR3 (N15081, N15080, N14898, N326);
not NOT1 (N15082, N15074);
not NOT1 (N15083, N15079);
nor NOR3 (N15084, N15069, N393, N1955);
nor NOR4 (N15085, N15076, N7930, N1213, N12669);
not NOT1 (N15086, N15072);
not NOT1 (N15087, N15084);
nor NOR4 (N15088, N15086, N5843, N13394, N14503);
or OR2 (N15089, N15077, N5035);
nand NAND2 (N15090, N15088, N11188);
or OR3 (N15091, N15075, N15034, N14609);
or OR4 (N15092, N15078, N628, N2485, N2931);
buf BUF1 (N15093, N15070);
and AND3 (N15094, N15085, N11362, N13687);
or OR2 (N15095, N15087, N3006);
nor NOR4 (N15096, N15092, N2299, N9986, N10465);
buf BUF1 (N15097, N15096);
or OR2 (N15098, N15089, N12160);
buf BUF1 (N15099, N15098);
xor XOR2 (N15100, N15090, N11547);
nand NAND3 (N15101, N15081, N14544, N11283);
and AND2 (N15102, N15100, N3391);
xor XOR2 (N15103, N15095, N13395);
nor NOR2 (N15104, N15099, N5197);
buf BUF1 (N15105, N15083);
and AND3 (N15106, N15091, N14800, N8817);
nor NOR2 (N15107, N15094, N13307);
nor NOR2 (N15108, N15105, N7599);
or OR3 (N15109, N15108, N14248, N2104);
not NOT1 (N15110, N15093);
not NOT1 (N15111, N15109);
nand NAND4 (N15112, N15102, N10420, N5550, N10584);
nand NAND4 (N15113, N15112, N870, N555, N6573);
buf BUF1 (N15114, N15106);
and AND2 (N15115, N15101, N14107);
buf BUF1 (N15116, N15107);
nor NOR4 (N15117, N15097, N518, N12405, N2663);
xor XOR2 (N15118, N15115, N14818);
xor XOR2 (N15119, N15113, N3316);
or OR4 (N15120, N15082, N8577, N7128, N13103);
buf BUF1 (N15121, N15110);
or OR4 (N15122, N15118, N14260, N3863, N1968);
not NOT1 (N15123, N15104);
and AND2 (N15124, N15116, N14581);
buf BUF1 (N15125, N15114);
nand NAND4 (N15126, N15117, N4533, N6784, N72);
not NOT1 (N15127, N15125);
or OR2 (N15128, N15103, N8152);
nor NOR2 (N15129, N15111, N4198);
buf BUF1 (N15130, N15129);
nand NAND2 (N15131, N15121, N7472);
xor XOR2 (N15132, N15122, N2995);
nor NOR2 (N15133, N15124, N4513);
xor XOR2 (N15134, N15126, N6816);
nor NOR3 (N15135, N15119, N6453, N14583);
buf BUF1 (N15136, N15128);
or OR2 (N15137, N15123, N586);
xor XOR2 (N15138, N15132, N513);
buf BUF1 (N15139, N15120);
nand NAND3 (N15140, N15131, N6779, N9299);
nand NAND2 (N15141, N15130, N4399);
xor XOR2 (N15142, N15136, N11813);
and AND2 (N15143, N15135, N13950);
buf BUF1 (N15144, N15141);
buf BUF1 (N15145, N15127);
xor XOR2 (N15146, N15133, N9240);
buf BUF1 (N15147, N15138);
not NOT1 (N15148, N15143);
nand NAND4 (N15149, N15137, N11642, N1249, N10425);
buf BUF1 (N15150, N15148);
buf BUF1 (N15151, N15140);
not NOT1 (N15152, N15147);
and AND4 (N15153, N15150, N6666, N1188, N5143);
xor XOR2 (N15154, N15153, N936);
or OR2 (N15155, N15152, N2400);
xor XOR2 (N15156, N15139, N14392);
nand NAND4 (N15157, N15146, N1042, N8055, N6036);
xor XOR2 (N15158, N15145, N4407);
nand NAND4 (N15159, N15158, N14516, N657, N3887);
buf BUF1 (N15160, N15149);
or OR2 (N15161, N15134, N9247);
xor XOR2 (N15162, N15142, N11503);
nand NAND3 (N15163, N15144, N5392, N10410);
xor XOR2 (N15164, N15160, N7391);
not NOT1 (N15165, N15154);
nor NOR4 (N15166, N15159, N10856, N11424, N6016);
not NOT1 (N15167, N15164);
not NOT1 (N15168, N15156);
or OR4 (N15169, N15163, N6143, N13207, N2522);
nand NAND2 (N15170, N15161, N2421);
buf BUF1 (N15171, N15157);
or OR4 (N15172, N15166, N10558, N6418, N832);
xor XOR2 (N15173, N15167, N10751);
nor NOR2 (N15174, N15168, N2392);
nor NOR4 (N15175, N15172, N1648, N5327, N2781);
xor XOR2 (N15176, N15169, N13046);
and AND4 (N15177, N15165, N11768, N2550, N12448);
xor XOR2 (N15178, N15171, N8341);
nand NAND4 (N15179, N15151, N2428, N7277, N11359);
buf BUF1 (N15180, N15155);
not NOT1 (N15181, N15162);
nor NOR4 (N15182, N15174, N12289, N10299, N967);
or OR2 (N15183, N15170, N5539);
buf BUF1 (N15184, N15173);
or OR2 (N15185, N15179, N11262);
or OR2 (N15186, N15184, N8290);
nand NAND3 (N15187, N15181, N4436, N12660);
buf BUF1 (N15188, N15178);
xor XOR2 (N15189, N15182, N3602);
nand NAND4 (N15190, N15175, N6767, N1991, N7613);
nand NAND2 (N15191, N15190, N6108);
and AND3 (N15192, N15186, N6433, N4253);
nand NAND4 (N15193, N15177, N10087, N8032, N9079);
not NOT1 (N15194, N15180);
nand NAND3 (N15195, N15194, N9497, N10459);
not NOT1 (N15196, N15188);
or OR2 (N15197, N15185, N12475);
or OR3 (N15198, N15196, N7209, N4974);
and AND4 (N15199, N15187, N9799, N3682, N12443);
buf BUF1 (N15200, N15183);
nor NOR3 (N15201, N15176, N10110, N267);
not NOT1 (N15202, N15193);
buf BUF1 (N15203, N15197);
and AND3 (N15204, N15202, N7222, N1340);
nor NOR3 (N15205, N15199, N2716, N13263);
not NOT1 (N15206, N15192);
xor XOR2 (N15207, N15198, N661);
xor XOR2 (N15208, N15201, N3582);
and AND2 (N15209, N15205, N6242);
or OR2 (N15210, N15206, N12638);
buf BUF1 (N15211, N15209);
not NOT1 (N15212, N15195);
nor NOR4 (N15213, N15212, N1050, N12477, N8193);
xor XOR2 (N15214, N15211, N11553);
nor NOR2 (N15215, N15200, N9125);
xor XOR2 (N15216, N15203, N1999);
and AND2 (N15217, N15208, N1605);
nor NOR2 (N15218, N15204, N7591);
and AND3 (N15219, N15216, N10321, N8164);
and AND4 (N15220, N15207, N12405, N919, N13293);
buf BUF1 (N15221, N15220);
or OR3 (N15222, N15210, N2163, N6530);
or OR2 (N15223, N15213, N14007);
xor XOR2 (N15224, N15221, N473);
nor NOR2 (N15225, N15222, N11996);
xor XOR2 (N15226, N15224, N2316);
or OR4 (N15227, N15219, N1145, N7954, N1240);
buf BUF1 (N15228, N15227);
xor XOR2 (N15229, N15226, N1076);
not NOT1 (N15230, N15218);
buf BUF1 (N15231, N15230);
not NOT1 (N15232, N15189);
not NOT1 (N15233, N15191);
nor NOR3 (N15234, N15214, N3742, N10189);
and AND4 (N15235, N15232, N8381, N15028, N8364);
xor XOR2 (N15236, N15225, N860);
or OR2 (N15237, N15228, N12100);
buf BUF1 (N15238, N15236);
nor NOR2 (N15239, N15215, N1755);
nand NAND2 (N15240, N15229, N13225);
not NOT1 (N15241, N15239);
not NOT1 (N15242, N15238);
buf BUF1 (N15243, N15234);
xor XOR2 (N15244, N15233, N13220);
nand NAND3 (N15245, N15241, N348, N6215);
and AND3 (N15246, N15240, N9488, N5419);
nor NOR4 (N15247, N15231, N15237, N12307, N9857);
buf BUF1 (N15248, N8882);
not NOT1 (N15249, N15248);
xor XOR2 (N15250, N15223, N14788);
nand NAND4 (N15251, N15250, N4455, N4323, N6469);
xor XOR2 (N15252, N15247, N13927);
xor XOR2 (N15253, N15217, N4490);
buf BUF1 (N15254, N15243);
xor XOR2 (N15255, N15249, N8111);
nor NOR2 (N15256, N15235, N8081);
nand NAND2 (N15257, N15252, N9300);
nand NAND4 (N15258, N15245, N14836, N14772, N9433);
buf BUF1 (N15259, N15256);
not NOT1 (N15260, N15259);
or OR3 (N15261, N15242, N6198, N5485);
or OR4 (N15262, N15255, N137, N515, N12136);
and AND3 (N15263, N15262, N6693, N5512);
not NOT1 (N15264, N15261);
not NOT1 (N15265, N15264);
nor NOR4 (N15266, N15258, N4644, N5670, N5114);
nor NOR2 (N15267, N15251, N5248);
or OR4 (N15268, N15267, N14475, N13712, N5979);
not NOT1 (N15269, N15265);
or OR4 (N15270, N15266, N1991, N6104, N7166);
nand NAND3 (N15271, N15257, N1046, N10990);
nor NOR3 (N15272, N15270, N3935, N6584);
buf BUF1 (N15273, N15271);
or OR4 (N15274, N15244, N12026, N2137, N9070);
xor XOR2 (N15275, N15260, N1105);
or OR4 (N15276, N15253, N2739, N1074, N7165);
nand NAND4 (N15277, N15274, N9261, N3471, N14397);
nand NAND3 (N15278, N15246, N2969, N6040);
nand NAND2 (N15279, N15272, N3128);
or OR3 (N15280, N15277, N10608, N2626);
buf BUF1 (N15281, N15279);
nand NAND3 (N15282, N15280, N7661, N7460);
xor XOR2 (N15283, N15273, N1794);
and AND3 (N15284, N15283, N8814, N11525);
not NOT1 (N15285, N15281);
not NOT1 (N15286, N15268);
nor NOR3 (N15287, N15269, N1511, N881);
buf BUF1 (N15288, N15278);
not NOT1 (N15289, N15285);
or OR4 (N15290, N15275, N7430, N1499, N14897);
xor XOR2 (N15291, N15288, N4018);
buf BUF1 (N15292, N15282);
and AND4 (N15293, N15287, N1940, N180, N14654);
xor XOR2 (N15294, N15291, N5970);
buf BUF1 (N15295, N15286);
nor NOR2 (N15296, N15289, N9058);
buf BUF1 (N15297, N15284);
nand NAND3 (N15298, N15296, N9912, N7746);
or OR4 (N15299, N15263, N2423, N4747, N659);
nand NAND3 (N15300, N15276, N11468, N6799);
or OR3 (N15301, N15300, N1844, N11125);
and AND2 (N15302, N15290, N13935);
or OR3 (N15303, N15295, N4820, N2988);
not NOT1 (N15304, N15303);
not NOT1 (N15305, N15254);
xor XOR2 (N15306, N15304, N15258);
or OR4 (N15307, N15293, N4995, N10977, N12015);
and AND4 (N15308, N15305, N1526, N9187, N7803);
xor XOR2 (N15309, N15308, N10892);
buf BUF1 (N15310, N15302);
nand NAND4 (N15311, N15307, N1384, N2908, N4676);
and AND4 (N15312, N15306, N5829, N1158, N8788);
not NOT1 (N15313, N15292);
and AND2 (N15314, N15310, N9647);
nand NAND2 (N15315, N15298, N1700);
xor XOR2 (N15316, N15297, N4909);
nor NOR2 (N15317, N15311, N1241);
and AND3 (N15318, N15309, N11651, N4741);
xor XOR2 (N15319, N15314, N4711);
not NOT1 (N15320, N15315);
nor NOR4 (N15321, N15320, N6262, N3944, N4341);
not NOT1 (N15322, N15299);
nor NOR3 (N15323, N15312, N14352, N14186);
not NOT1 (N15324, N15316);
or OR2 (N15325, N15323, N11904);
and AND4 (N15326, N15294, N6468, N13445, N84);
or OR3 (N15327, N15301, N8242, N2183);
not NOT1 (N15328, N15324);
and AND4 (N15329, N15317, N7070, N6888, N10411);
not NOT1 (N15330, N15313);
nand NAND2 (N15331, N15319, N11871);
nor NOR2 (N15332, N15330, N2518);
not NOT1 (N15333, N15331);
or OR3 (N15334, N15326, N8153, N5902);
buf BUF1 (N15335, N15321);
nand NAND3 (N15336, N15322, N865, N854);
or OR4 (N15337, N15328, N1172, N6358, N3826);
nor NOR4 (N15338, N15335, N8222, N10503, N10596);
nor NOR3 (N15339, N15329, N10698, N11784);
xor XOR2 (N15340, N15339, N14718);
nand NAND4 (N15341, N15327, N7065, N8857, N14781);
buf BUF1 (N15342, N15332);
buf BUF1 (N15343, N15333);
or OR2 (N15344, N15336, N8158);
and AND3 (N15345, N15318, N14511, N9960);
or OR2 (N15346, N15341, N6323);
and AND4 (N15347, N15346, N2800, N14361, N12077);
buf BUF1 (N15348, N15342);
and AND2 (N15349, N15345, N1097);
and AND2 (N15350, N15338, N7802);
nand NAND4 (N15351, N15349, N418, N3237, N6260);
or OR3 (N15352, N15340, N7889, N9362);
and AND4 (N15353, N15344, N12462, N5569, N8778);
and AND3 (N15354, N15325, N11831, N11351);
or OR4 (N15355, N15337, N8441, N12961, N2714);
and AND3 (N15356, N15334, N12822, N13649);
xor XOR2 (N15357, N15355, N325);
or OR2 (N15358, N15354, N8178);
xor XOR2 (N15359, N15348, N8053);
not NOT1 (N15360, N15359);
and AND4 (N15361, N15347, N5249, N2587, N12888);
nand NAND2 (N15362, N15356, N477);
and AND4 (N15363, N15360, N9953, N3364, N12408);
nand NAND3 (N15364, N15353, N4954, N3275);
or OR4 (N15365, N15364, N15333, N13369, N13781);
xor XOR2 (N15366, N15361, N8626);
nand NAND2 (N15367, N15351, N10447);
and AND4 (N15368, N15363, N11740, N15097, N11537);
nor NOR3 (N15369, N15368, N3276, N4108);
not NOT1 (N15370, N15366);
not NOT1 (N15371, N15362);
and AND3 (N15372, N15369, N4420, N14471);
and AND3 (N15373, N15350, N1218, N8621);
nand NAND4 (N15374, N15371, N11718, N9614, N8388);
and AND4 (N15375, N15365, N5081, N12071, N6764);
and AND3 (N15376, N15375, N4045, N12974);
nand NAND3 (N15377, N15343, N1850, N12381);
buf BUF1 (N15378, N15376);
nand NAND2 (N15379, N15370, N4420);
nand NAND4 (N15380, N15379, N12816, N2814, N11440);
and AND4 (N15381, N15372, N13486, N9212, N2010);
buf BUF1 (N15382, N15381);
or OR3 (N15383, N15382, N1880, N1664);
or OR2 (N15384, N15377, N6406);
nor NOR4 (N15385, N15352, N4458, N3485, N6223);
xor XOR2 (N15386, N15373, N2964);
nor NOR4 (N15387, N15358, N12988, N1911, N1705);
nand NAND2 (N15388, N15378, N15042);
not NOT1 (N15389, N15383);
nor NOR3 (N15390, N15385, N7123, N10223);
or OR4 (N15391, N15387, N11732, N8975, N13413);
or OR3 (N15392, N15390, N8169, N12504);
and AND4 (N15393, N15374, N4709, N7983, N13910);
not NOT1 (N15394, N15380);
not NOT1 (N15395, N15393);
or OR2 (N15396, N15391, N5799);
buf BUF1 (N15397, N15392);
buf BUF1 (N15398, N15395);
or OR4 (N15399, N15388, N14741, N10717, N9347);
not NOT1 (N15400, N15367);
buf BUF1 (N15401, N15394);
nor NOR2 (N15402, N15389, N15);
or OR2 (N15403, N15386, N6838);
or OR2 (N15404, N15401, N12533);
not NOT1 (N15405, N15402);
not NOT1 (N15406, N15399);
nand NAND3 (N15407, N15406, N1274, N3301);
and AND4 (N15408, N15405, N3653, N7552, N15097);
buf BUF1 (N15409, N15357);
not NOT1 (N15410, N15400);
and AND4 (N15411, N15396, N11027, N5575, N13095);
not NOT1 (N15412, N15411);
xor XOR2 (N15413, N15404, N10290);
and AND2 (N15414, N15412, N6087);
xor XOR2 (N15415, N15398, N5602);
and AND2 (N15416, N15409, N591);
or OR4 (N15417, N15397, N11314, N3775, N5505);
nor NOR4 (N15418, N15403, N9436, N12506, N2178);
or OR4 (N15419, N15416, N1779, N10288, N7394);
buf BUF1 (N15420, N15414);
nand NAND4 (N15421, N15419, N13685, N26, N912);
and AND2 (N15422, N15420, N1417);
or OR3 (N15423, N15422, N10942, N1850);
not NOT1 (N15424, N15423);
nand NAND2 (N15425, N15421, N10374);
or OR2 (N15426, N15413, N12904);
nor NOR3 (N15427, N15424, N12382, N548);
or OR3 (N15428, N15407, N14372, N13185);
nand NAND3 (N15429, N15408, N11280, N3664);
not NOT1 (N15430, N15425);
buf BUF1 (N15431, N15384);
and AND4 (N15432, N15429, N3619, N7604, N15402);
or OR3 (N15433, N15410, N12870, N3554);
not NOT1 (N15434, N15433);
nor NOR4 (N15435, N15430, N7259, N10410, N7521);
nand NAND4 (N15436, N15428, N8497, N11327, N14925);
xor XOR2 (N15437, N15418, N8285);
nor NOR4 (N15438, N15427, N11016, N4891, N1150);
and AND4 (N15439, N15434, N7969, N8839, N1110);
xor XOR2 (N15440, N15415, N8890);
and AND4 (N15441, N15417, N13638, N2962, N6678);
buf BUF1 (N15442, N15441);
not NOT1 (N15443, N15437);
not NOT1 (N15444, N15435);
nand NAND3 (N15445, N15438, N9053, N10522);
or OR3 (N15446, N15436, N14610, N603);
nand NAND3 (N15447, N15426, N15151, N5188);
buf BUF1 (N15448, N15445);
or OR2 (N15449, N15432, N9324);
xor XOR2 (N15450, N15439, N937);
nor NOR4 (N15451, N15448, N3422, N8613, N12756);
nand NAND4 (N15452, N15431, N4363, N1089, N10789);
not NOT1 (N15453, N15442);
xor XOR2 (N15454, N15440, N10639);
or OR4 (N15455, N15443, N12199, N8109, N12545);
and AND2 (N15456, N15453, N8568);
or OR2 (N15457, N15450, N10828);
and AND2 (N15458, N15452, N7161);
xor XOR2 (N15459, N15454, N15277);
xor XOR2 (N15460, N15459, N4242);
xor XOR2 (N15461, N15444, N1447);
xor XOR2 (N15462, N15449, N8);
nand NAND2 (N15463, N15461, N9954);
nand NAND2 (N15464, N15457, N4689);
nand NAND2 (N15465, N15447, N11288);
nand NAND3 (N15466, N15465, N3794, N1170);
nor NOR3 (N15467, N15463, N10783, N6549);
buf BUF1 (N15468, N15462);
not NOT1 (N15469, N15458);
and AND4 (N15470, N15446, N7247, N9821, N4917);
buf BUF1 (N15471, N15467);
nor NOR2 (N15472, N15451, N9127);
and AND4 (N15473, N15466, N3838, N5029, N7652);
xor XOR2 (N15474, N15472, N9048);
buf BUF1 (N15475, N15460);
or OR2 (N15476, N15470, N14610);
nor NOR2 (N15477, N15464, N10399);
xor XOR2 (N15478, N15471, N14956);
and AND3 (N15479, N15475, N6844, N8235);
buf BUF1 (N15480, N15469);
not NOT1 (N15481, N15468);
xor XOR2 (N15482, N15480, N7366);
and AND3 (N15483, N15479, N12890, N14140);
and AND4 (N15484, N15456, N8294, N9605, N5363);
not NOT1 (N15485, N15483);
nand NAND3 (N15486, N15478, N4471, N11375);
xor XOR2 (N15487, N15455, N2632);
not NOT1 (N15488, N15484);
nand NAND2 (N15489, N15482, N4776);
xor XOR2 (N15490, N15488, N10767);
and AND3 (N15491, N15473, N15395, N15383);
nor NOR4 (N15492, N15485, N15487, N12549, N4384);
xor XOR2 (N15493, N1738, N9900);
not NOT1 (N15494, N15476);
xor XOR2 (N15495, N15481, N5622);
xor XOR2 (N15496, N15486, N7075);
not NOT1 (N15497, N15489);
nor NOR2 (N15498, N15490, N10001);
buf BUF1 (N15499, N15477);
xor XOR2 (N15500, N15498, N10382);
or OR2 (N15501, N15491, N2434);
not NOT1 (N15502, N15494);
xor XOR2 (N15503, N15500, N5103);
nor NOR4 (N15504, N15492, N12867, N3023, N12513);
nand NAND2 (N15505, N15496, N13687);
nor NOR4 (N15506, N15493, N3144, N4813, N12404);
buf BUF1 (N15507, N15499);
xor XOR2 (N15508, N15504, N6445);
xor XOR2 (N15509, N15506, N7799);
buf BUF1 (N15510, N15505);
not NOT1 (N15511, N15503);
nor NOR3 (N15512, N15474, N8638, N5620);
nor NOR2 (N15513, N15497, N11838);
nor NOR4 (N15514, N15508, N6062, N13668, N1949);
buf BUF1 (N15515, N15514);
and AND3 (N15516, N15502, N11537, N4841);
and AND3 (N15517, N15507, N4904, N7084);
nor NOR4 (N15518, N15495, N1221, N8160, N14308);
buf BUF1 (N15519, N15510);
xor XOR2 (N15520, N15509, N2766);
xor XOR2 (N15521, N15515, N13634);
buf BUF1 (N15522, N15519);
xor XOR2 (N15523, N15516, N11816);
xor XOR2 (N15524, N15523, N11951);
nor NOR2 (N15525, N15501, N6136);
and AND2 (N15526, N15512, N8301);
and AND2 (N15527, N15518, N8427);
nand NAND2 (N15528, N15522, N15170);
and AND2 (N15529, N15527, N3118);
or OR3 (N15530, N15520, N1196, N2330);
nand NAND2 (N15531, N15517, N5469);
xor XOR2 (N15532, N15525, N2836);
xor XOR2 (N15533, N15529, N5303);
and AND3 (N15534, N15526, N9898, N5812);
not NOT1 (N15535, N15524);
xor XOR2 (N15536, N15513, N14441);
not NOT1 (N15537, N15532);
nand NAND4 (N15538, N15534, N2502, N7790, N14854);
nand NAND4 (N15539, N15521, N5622, N9441, N4025);
buf BUF1 (N15540, N15531);
and AND2 (N15541, N15528, N5980);
xor XOR2 (N15542, N15511, N12816);
or OR4 (N15543, N15540, N11584, N11098, N2646);
and AND4 (N15544, N15538, N14495, N5785, N13113);
nand NAND2 (N15545, N15539, N1806);
or OR4 (N15546, N15535, N9106, N6504, N681);
and AND2 (N15547, N15536, N826);
nand NAND3 (N15548, N15533, N7733, N9509);
and AND4 (N15549, N15544, N12908, N5852, N127);
xor XOR2 (N15550, N15547, N10564);
xor XOR2 (N15551, N15542, N9845);
nand NAND4 (N15552, N15541, N597, N7360, N3736);
xor XOR2 (N15553, N15543, N296);
nand NAND2 (N15554, N15551, N4476);
or OR4 (N15555, N15549, N15078, N762, N8805);
and AND4 (N15556, N15550, N1455, N13801, N12292);
buf BUF1 (N15557, N15537);
buf BUF1 (N15558, N15553);
nor NOR4 (N15559, N15556, N4873, N10551, N15022);
and AND3 (N15560, N15530, N625, N9846);
nor NOR4 (N15561, N15555, N7276, N3229, N4971);
not NOT1 (N15562, N15560);
not NOT1 (N15563, N15559);
nor NOR2 (N15564, N15546, N5777);
not NOT1 (N15565, N15552);
nand NAND4 (N15566, N15554, N13794, N1006, N4895);
or OR4 (N15567, N15563, N2907, N12624, N4644);
nand NAND4 (N15568, N15567, N13866, N11677, N44);
and AND4 (N15569, N15558, N10626, N10373, N1362);
xor XOR2 (N15570, N15548, N15392);
or OR2 (N15571, N15565, N6728);
and AND2 (N15572, N15564, N11834);
or OR3 (N15573, N15561, N11358, N8242);
buf BUF1 (N15574, N15562);
nor NOR2 (N15575, N15568, N1217);
xor XOR2 (N15576, N15566, N10517);
nand NAND2 (N15577, N15571, N3335);
and AND3 (N15578, N15573, N14964, N8876);
or OR4 (N15579, N15572, N9894, N13139, N2514);
or OR4 (N15580, N15557, N12590, N2575, N5558);
nor NOR4 (N15581, N15545, N946, N12473, N12695);
nor NOR3 (N15582, N15576, N5620, N12501);
nand NAND4 (N15583, N15579, N13011, N10025, N5846);
nor NOR3 (N15584, N15569, N6050, N13490);
buf BUF1 (N15585, N15578);
buf BUF1 (N15586, N15583);
buf BUF1 (N15587, N15581);
and AND4 (N15588, N15570, N6939, N4640, N534);
or OR4 (N15589, N15577, N13877, N13749, N14198);
or OR3 (N15590, N15586, N13341, N14997);
buf BUF1 (N15591, N15575);
not NOT1 (N15592, N15588);
or OR3 (N15593, N15574, N1722, N3548);
buf BUF1 (N15594, N15591);
buf BUF1 (N15595, N15593);
nor NOR3 (N15596, N15587, N6749, N12981);
not NOT1 (N15597, N15580);
or OR3 (N15598, N15597, N12047, N13376);
not NOT1 (N15599, N15589);
or OR4 (N15600, N15584, N4162, N15116, N5283);
not NOT1 (N15601, N15599);
or OR3 (N15602, N15594, N10136, N4371);
not NOT1 (N15603, N15601);
not NOT1 (N15604, N15598);
nand NAND2 (N15605, N15585, N10217);
buf BUF1 (N15606, N15582);
or OR2 (N15607, N15596, N4877);
nor NOR2 (N15608, N15595, N5241);
buf BUF1 (N15609, N15607);
and AND3 (N15610, N15590, N12191, N995);
nand NAND2 (N15611, N15592, N2409);
xor XOR2 (N15612, N15602, N4670);
or OR3 (N15613, N15600, N6851, N12816);
buf BUF1 (N15614, N15611);
buf BUF1 (N15615, N15613);
buf BUF1 (N15616, N15609);
and AND3 (N15617, N15612, N617, N9147);
nor NOR4 (N15618, N15615, N7937, N6575, N2637);
nand NAND2 (N15619, N15610, N7980);
buf BUF1 (N15620, N15614);
not NOT1 (N15621, N15606);
not NOT1 (N15622, N15620);
buf BUF1 (N15623, N15603);
buf BUF1 (N15624, N15608);
and AND2 (N15625, N15624, N2891);
buf BUF1 (N15626, N15605);
buf BUF1 (N15627, N15622);
nor NOR2 (N15628, N15616, N12236);
nor NOR2 (N15629, N15628, N9240);
nand NAND2 (N15630, N15621, N12101);
or OR3 (N15631, N15629, N7373, N7807);
nand NAND4 (N15632, N15625, N6039, N9094, N255);
and AND3 (N15633, N15631, N2630, N11215);
not NOT1 (N15634, N15623);
or OR2 (N15635, N15627, N7449);
nand NAND4 (N15636, N15617, N15294, N12371, N9308);
nand NAND3 (N15637, N15635, N12935, N1184);
buf BUF1 (N15638, N15633);
not NOT1 (N15639, N15636);
xor XOR2 (N15640, N15639, N13282);
xor XOR2 (N15641, N15618, N10046);
or OR3 (N15642, N15619, N8524, N10546);
nor NOR2 (N15643, N15637, N383);
buf BUF1 (N15644, N15604);
nor NOR3 (N15645, N15643, N5698, N2777);
buf BUF1 (N15646, N15642);
buf BUF1 (N15647, N15641);
nand NAND4 (N15648, N15626, N8869, N11562, N10950);
xor XOR2 (N15649, N15638, N14275);
nor NOR2 (N15650, N15632, N3358);
buf BUF1 (N15651, N15650);
nor NOR2 (N15652, N15634, N8817);
xor XOR2 (N15653, N15652, N6815);
nand NAND3 (N15654, N15651, N15032, N8662);
buf BUF1 (N15655, N15646);
and AND3 (N15656, N15649, N3879, N14862);
not NOT1 (N15657, N15653);
nand NAND2 (N15658, N15644, N4372);
not NOT1 (N15659, N15640);
or OR3 (N15660, N15657, N14571, N6740);
and AND3 (N15661, N15630, N12856, N13531);
nand NAND2 (N15662, N15654, N12495);
and AND2 (N15663, N15648, N3341);
or OR3 (N15664, N15663, N3163, N3199);
xor XOR2 (N15665, N15647, N3333);
nand NAND2 (N15666, N15665, N2053);
or OR2 (N15667, N15645, N10635);
nor NOR4 (N15668, N15660, N7876, N3479, N3284);
and AND2 (N15669, N15656, N10430);
or OR4 (N15670, N15664, N10924, N13796, N4167);
or OR2 (N15671, N15662, N1059);
and AND3 (N15672, N15659, N10421, N5348);
or OR4 (N15673, N15669, N8079, N12617, N6833);
or OR3 (N15674, N15661, N12307, N14079);
or OR2 (N15675, N15667, N8054);
and AND4 (N15676, N15671, N2029, N9697, N252);
nor NOR2 (N15677, N15673, N14169);
buf BUF1 (N15678, N15675);
or OR4 (N15679, N15672, N5223, N4276, N13327);
not NOT1 (N15680, N15677);
or OR2 (N15681, N15676, N11815);
nand NAND2 (N15682, N15674, N12184);
buf BUF1 (N15683, N15678);
not NOT1 (N15684, N15680);
xor XOR2 (N15685, N15668, N8032);
or OR2 (N15686, N15682, N9296);
and AND4 (N15687, N15684, N7554, N14488, N14978);
or OR4 (N15688, N15670, N5856, N1100, N12367);
xor XOR2 (N15689, N15666, N10635);
and AND2 (N15690, N15685, N14685);
xor XOR2 (N15691, N15679, N15142);
nand NAND4 (N15692, N15655, N3260, N6366, N7420);
nor NOR4 (N15693, N15689, N14382, N5398, N8880);
xor XOR2 (N15694, N15681, N5698);
and AND4 (N15695, N15688, N1909, N6620, N10516);
and AND3 (N15696, N15686, N6562, N6848);
and AND2 (N15697, N15696, N12539);
and AND2 (N15698, N15691, N8);
and AND3 (N15699, N15695, N14459, N8702);
or OR4 (N15700, N15687, N8070, N5415, N2551);
nand NAND4 (N15701, N15690, N9077, N11188, N15597);
or OR4 (N15702, N15683, N4485, N3920, N15124);
nand NAND2 (N15703, N15694, N15686);
nor NOR2 (N15704, N15703, N1093);
and AND4 (N15705, N15697, N8969, N2052, N5503);
not NOT1 (N15706, N15658);
and AND3 (N15707, N15702, N7442, N4095);
xor XOR2 (N15708, N15700, N3094);
and AND2 (N15709, N15706, N723);
not NOT1 (N15710, N15709);
not NOT1 (N15711, N15707);
nor NOR2 (N15712, N15699, N2969);
not NOT1 (N15713, N15710);
and AND4 (N15714, N15712, N15546, N8682, N12401);
and AND3 (N15715, N15708, N12974, N6633);
nor NOR4 (N15716, N15711, N11735, N2554, N5253);
or OR2 (N15717, N15693, N10581);
nand NAND3 (N15718, N15713, N2427, N14166);
not NOT1 (N15719, N15715);
xor XOR2 (N15720, N15705, N7787);
not NOT1 (N15721, N15714);
xor XOR2 (N15722, N15719, N9989);
or OR3 (N15723, N15716, N7540, N2341);
not NOT1 (N15724, N15692);
nor NOR4 (N15725, N15701, N12985, N203, N9022);
or OR3 (N15726, N15725, N11332, N14142);
not NOT1 (N15727, N15721);
not NOT1 (N15728, N15704);
or OR2 (N15729, N15698, N10327);
buf BUF1 (N15730, N15720);
and AND4 (N15731, N15718, N875, N12889, N9347);
xor XOR2 (N15732, N15731, N12670);
and AND4 (N15733, N15724, N2213, N5695, N5475);
nor NOR4 (N15734, N15727, N15685, N9242, N12883);
xor XOR2 (N15735, N15729, N7567);
xor XOR2 (N15736, N15735, N12350);
nor NOR2 (N15737, N15726, N2690);
and AND4 (N15738, N15733, N2090, N9664, N13293);
nand NAND3 (N15739, N15737, N9045, N15368);
xor XOR2 (N15740, N15738, N7337);
nand NAND3 (N15741, N15734, N6628, N5343);
buf BUF1 (N15742, N15728);
nor NOR4 (N15743, N15742, N12758, N14358, N12905);
and AND2 (N15744, N15741, N10011);
and AND2 (N15745, N15717, N3245);
or OR2 (N15746, N15732, N3316);
or OR2 (N15747, N15744, N1871);
not NOT1 (N15748, N15740);
not NOT1 (N15749, N15722);
nand NAND4 (N15750, N15747, N4879, N4172, N8498);
not NOT1 (N15751, N15739);
not NOT1 (N15752, N15745);
buf BUF1 (N15753, N15736);
or OR3 (N15754, N15751, N3448, N9396);
or OR2 (N15755, N15743, N14376);
buf BUF1 (N15756, N15749);
buf BUF1 (N15757, N15755);
nor NOR4 (N15758, N15754, N13080, N5406, N1504);
buf BUF1 (N15759, N15730);
nand NAND4 (N15760, N15752, N11197, N11406, N7671);
not NOT1 (N15761, N15758);
nor NOR3 (N15762, N15759, N2178, N12209);
or OR2 (N15763, N15757, N5937);
nand NAND2 (N15764, N15756, N13584);
and AND4 (N15765, N15764, N4685, N8103, N6094);
not NOT1 (N15766, N15748);
not NOT1 (N15767, N15746);
buf BUF1 (N15768, N15753);
buf BUF1 (N15769, N15762);
buf BUF1 (N15770, N15763);
nand NAND4 (N15771, N15770, N13774, N7926, N9624);
nor NOR3 (N15772, N15768, N5313, N15485);
and AND3 (N15773, N15723, N15266, N1440);
or OR3 (N15774, N15750, N11917, N8556);
and AND4 (N15775, N15773, N326, N6237, N56);
nand NAND3 (N15776, N15765, N2908, N2541);
nor NOR3 (N15777, N15776, N10767, N10447);
and AND3 (N15778, N15772, N1973, N4142);
or OR2 (N15779, N15767, N1744);
and AND3 (N15780, N15761, N3602, N4039);
buf BUF1 (N15781, N15780);
or OR4 (N15782, N15769, N208, N3570, N5920);
or OR4 (N15783, N15766, N14525, N4960, N9058);
nor NOR4 (N15784, N15778, N15590, N12022, N15155);
not NOT1 (N15785, N15771);
and AND4 (N15786, N15760, N13314, N6409, N13476);
buf BUF1 (N15787, N15784);
xor XOR2 (N15788, N15774, N14018);
buf BUF1 (N15789, N15777);
and AND3 (N15790, N15781, N5693, N3113);
xor XOR2 (N15791, N15788, N14789);
and AND2 (N15792, N15790, N5650);
nor NOR4 (N15793, N15789, N10595, N781, N7825);
not NOT1 (N15794, N15787);
not NOT1 (N15795, N15782);
xor XOR2 (N15796, N15783, N12101);
nand NAND4 (N15797, N15794, N4870, N9187, N703);
or OR4 (N15798, N15795, N10020, N13106, N3464);
nand NAND4 (N15799, N15793, N12216, N389, N6404);
buf BUF1 (N15800, N15779);
and AND4 (N15801, N15799, N13550, N12444, N4914);
not NOT1 (N15802, N15792);
or OR3 (N15803, N15786, N9837, N9314);
xor XOR2 (N15804, N15800, N9026);
buf BUF1 (N15805, N15775);
xor XOR2 (N15806, N15785, N9254);
and AND3 (N15807, N15796, N12065, N13522);
or OR3 (N15808, N15804, N5393, N2784);
and AND3 (N15809, N15808, N12692, N14989);
nor NOR3 (N15810, N15791, N5927, N11847);
or OR3 (N15811, N15809, N7465, N10686);
and AND3 (N15812, N15807, N14590, N8097);
nand NAND3 (N15813, N15806, N14899, N14959);
not NOT1 (N15814, N15802);
and AND2 (N15815, N15798, N7120);
buf BUF1 (N15816, N15803);
buf BUF1 (N15817, N15813);
nand NAND2 (N15818, N15810, N8171);
xor XOR2 (N15819, N15812, N7772);
not NOT1 (N15820, N15818);
xor XOR2 (N15821, N15820, N9841);
nor NOR4 (N15822, N15811, N3533, N2702, N15767);
nand NAND4 (N15823, N15817, N7826, N14758, N4436);
nand NAND2 (N15824, N15822, N10442);
and AND4 (N15825, N15821, N6209, N2718, N1582);
not NOT1 (N15826, N15814);
or OR4 (N15827, N15805, N4031, N8144, N12026);
buf BUF1 (N15828, N15826);
xor XOR2 (N15829, N15824, N12731);
not NOT1 (N15830, N15829);
nor NOR3 (N15831, N15828, N8480, N14479);
xor XOR2 (N15832, N15797, N7355);
buf BUF1 (N15833, N15815);
or OR2 (N15834, N15801, N14269);
nand NAND2 (N15835, N15834, N11103);
buf BUF1 (N15836, N15831);
not NOT1 (N15837, N15835);
nor NOR3 (N15838, N15819, N1015, N7224);
buf BUF1 (N15839, N15836);
or OR3 (N15840, N15838, N8538, N5860);
not NOT1 (N15841, N15823);
buf BUF1 (N15842, N15841);
nand NAND4 (N15843, N15827, N6600, N3021, N15308);
and AND4 (N15844, N15833, N9800, N7373, N7803);
nor NOR2 (N15845, N15843, N8270);
buf BUF1 (N15846, N15832);
not NOT1 (N15847, N15839);
not NOT1 (N15848, N15842);
or OR3 (N15849, N15846, N172, N10289);
not NOT1 (N15850, N15825);
not NOT1 (N15851, N15847);
nor NOR3 (N15852, N15837, N5578, N181);
or OR4 (N15853, N15845, N12085, N10241, N15677);
buf BUF1 (N15854, N15850);
nor NOR2 (N15855, N15853, N12351);
xor XOR2 (N15856, N15816, N14102);
nor NOR3 (N15857, N15849, N6543, N59);
or OR3 (N15858, N15857, N653, N5620);
nor NOR3 (N15859, N15844, N8003, N8954);
or OR3 (N15860, N15851, N13932, N13176);
nor NOR2 (N15861, N15848, N6490);
not NOT1 (N15862, N15859);
or OR2 (N15863, N15861, N5572);
nor NOR4 (N15864, N15860, N40, N4082, N7899);
and AND2 (N15865, N15856, N5183);
or OR3 (N15866, N15840, N11690, N9337);
and AND3 (N15867, N15852, N14862, N2385);
not NOT1 (N15868, N15862);
nand NAND3 (N15869, N15868, N15500, N5845);
xor XOR2 (N15870, N15867, N12185);
or OR4 (N15871, N15870, N6855, N9768, N15864);
not NOT1 (N15872, N2049);
and AND4 (N15873, N15854, N1186, N500, N7547);
buf BUF1 (N15874, N15869);
nor NOR4 (N15875, N15855, N13129, N14261, N4800);
buf BUF1 (N15876, N15874);
and AND4 (N15877, N15872, N14476, N10871, N2105);
nor NOR4 (N15878, N15876, N2963, N11947, N12189);
nor NOR3 (N15879, N15863, N7120, N9474);
nand NAND4 (N15880, N15858, N3071, N4898, N3752);
nor NOR2 (N15881, N15875, N630);
nand NAND3 (N15882, N15873, N11, N3975);
not NOT1 (N15883, N15879);
and AND2 (N15884, N15883, N13502);
nand NAND3 (N15885, N15884, N3728, N7196);
buf BUF1 (N15886, N15871);
xor XOR2 (N15887, N15881, N11631);
nor NOR4 (N15888, N15865, N14094, N13131, N9335);
and AND2 (N15889, N15878, N2170);
nand NAND3 (N15890, N15880, N10762, N6811);
and AND3 (N15891, N15886, N1434, N10795);
buf BUF1 (N15892, N15866);
buf BUF1 (N15893, N15887);
buf BUF1 (N15894, N15882);
nand NAND4 (N15895, N15892, N12160, N2075, N5632);
nand NAND3 (N15896, N15893, N14077, N12602);
nor NOR4 (N15897, N15889, N12988, N13175, N7888);
or OR4 (N15898, N15896, N1885, N189, N5725);
nor NOR4 (N15899, N15891, N15086, N14574, N15693);
nor NOR3 (N15900, N15830, N12513, N13755);
xor XOR2 (N15901, N15877, N5860);
not NOT1 (N15902, N15897);
not NOT1 (N15903, N15888);
xor XOR2 (N15904, N15890, N10752);
not NOT1 (N15905, N15900);
xor XOR2 (N15906, N15904, N9742);
xor XOR2 (N15907, N15894, N11553);
and AND4 (N15908, N15903, N4396, N5229, N11447);
nand NAND2 (N15909, N15898, N9912);
nor NOR4 (N15910, N15885, N2020, N13181, N3313);
or OR3 (N15911, N15909, N12702, N1050);
xor XOR2 (N15912, N15907, N5677);
nor NOR3 (N15913, N15901, N13758, N5953);
nor NOR4 (N15914, N15906, N12480, N894, N5384);
xor XOR2 (N15915, N15911, N13525);
or OR2 (N15916, N15910, N14748);
and AND2 (N15917, N15915, N2722);
nor NOR3 (N15918, N15917, N12256, N6115);
nand NAND3 (N15919, N15913, N13342, N11411);
buf BUF1 (N15920, N15908);
xor XOR2 (N15921, N15914, N5365);
nand NAND4 (N15922, N15905, N6283, N12924, N11757);
nand NAND3 (N15923, N15895, N5260, N1798);
not NOT1 (N15924, N15922);
buf BUF1 (N15925, N15912);
not NOT1 (N15926, N15902);
nand NAND2 (N15927, N15899, N7611);
nor NOR4 (N15928, N15921, N3269, N4436, N11684);
xor XOR2 (N15929, N15923, N5104);
nor NOR3 (N15930, N15925, N5222, N13759);
nor NOR2 (N15931, N15918, N3860);
and AND4 (N15932, N15919, N14310, N6954, N5731);
nand NAND4 (N15933, N15920, N13562, N4780, N1367);
or OR3 (N15934, N15931, N8050, N10626);
xor XOR2 (N15935, N15926, N4825);
nor NOR3 (N15936, N15928, N8969, N1274);
xor XOR2 (N15937, N15932, N7723);
buf BUF1 (N15938, N15916);
nand NAND3 (N15939, N15927, N11315, N4188);
not NOT1 (N15940, N15924);
and AND2 (N15941, N15940, N2032);
nand NAND4 (N15942, N15934, N12372, N13552, N2801);
and AND2 (N15943, N15930, N8807);
or OR3 (N15944, N15929, N8737, N2062);
buf BUF1 (N15945, N15937);
not NOT1 (N15946, N15943);
or OR2 (N15947, N15936, N13215);
not NOT1 (N15948, N15945);
nand NAND3 (N15949, N15938, N9362, N10615);
or OR2 (N15950, N15941, N10468);
nor NOR2 (N15951, N15942, N9216);
or OR4 (N15952, N15946, N12632, N12420, N4239);
or OR4 (N15953, N15952, N12632, N2706, N5600);
not NOT1 (N15954, N15953);
and AND2 (N15955, N15935, N14207);
nand NAND4 (N15956, N15939, N5682, N1271, N3437);
and AND2 (N15957, N15948, N15532);
nand NAND3 (N15958, N15933, N15301, N13203);
nand NAND2 (N15959, N15951, N10189);
and AND2 (N15960, N15955, N2115);
buf BUF1 (N15961, N15944);
or OR2 (N15962, N15956, N8642);
xor XOR2 (N15963, N15960, N5343);
nand NAND2 (N15964, N15963, N4298);
and AND4 (N15965, N15957, N12796, N8664, N10971);
xor XOR2 (N15966, N15958, N10296);
buf BUF1 (N15967, N15964);
nor NOR3 (N15968, N15965, N15209, N14717);
xor XOR2 (N15969, N15961, N5584);
or OR3 (N15970, N15969, N1506, N997);
and AND4 (N15971, N15968, N2801, N3059, N11854);
xor XOR2 (N15972, N15962, N6921);
or OR3 (N15973, N15970, N15714, N10085);
nor NOR4 (N15974, N15949, N2948, N13546, N8532);
buf BUF1 (N15975, N15971);
and AND2 (N15976, N15972, N9372);
xor XOR2 (N15977, N15950, N10001);
nor NOR3 (N15978, N15947, N5253, N6246);
not NOT1 (N15979, N15959);
and AND2 (N15980, N15976, N1890);
xor XOR2 (N15981, N15973, N11674);
nor NOR2 (N15982, N15979, N13032);
not NOT1 (N15983, N15981);
nor NOR3 (N15984, N15974, N5213, N5521);
and AND3 (N15985, N15975, N11706, N9991);
buf BUF1 (N15986, N15967);
and AND3 (N15987, N15986, N5431, N3463);
nor NOR3 (N15988, N15978, N3881, N3794);
buf BUF1 (N15989, N15985);
or OR4 (N15990, N15989, N9057, N13188, N15880);
buf BUF1 (N15991, N15982);
xor XOR2 (N15992, N15988, N3059);
xor XOR2 (N15993, N15954, N7759);
nor NOR4 (N15994, N15990, N8145, N5306, N2374);
not NOT1 (N15995, N15984);
buf BUF1 (N15996, N15992);
or OR4 (N15997, N15983, N2021, N15114, N14286);
xor XOR2 (N15998, N15994, N9329);
buf BUF1 (N15999, N15991);
nor NOR3 (N16000, N15977, N14313, N8146);
nand NAND3 (N16001, N15999, N15103, N885);
and AND3 (N16002, N15987, N4810, N12255);
or OR2 (N16003, N15966, N6457);
not NOT1 (N16004, N16003);
or OR2 (N16005, N16004, N10986);
not NOT1 (N16006, N15996);
nand NAND2 (N16007, N16002, N11254);
nor NOR2 (N16008, N15997, N8509);
xor XOR2 (N16009, N15998, N12683);
xor XOR2 (N16010, N16001, N8779);
buf BUF1 (N16011, N16006);
buf BUF1 (N16012, N16000);
or OR4 (N16013, N16005, N3592, N15297, N5518);
not NOT1 (N16014, N16007);
nand NAND4 (N16015, N16008, N1885, N7885, N4613);
or OR3 (N16016, N16010, N7812, N2878);
xor XOR2 (N16017, N15980, N11331);
nand NAND2 (N16018, N16017, N6938);
nand NAND4 (N16019, N16013, N7939, N5442, N14903);
not NOT1 (N16020, N16009);
buf BUF1 (N16021, N16012);
and AND4 (N16022, N15993, N10205, N6853, N8235);
buf BUF1 (N16023, N15995);
nand NAND4 (N16024, N16019, N2908, N8890, N9405);
and AND3 (N16025, N16018, N519, N13789);
or OR4 (N16026, N16014, N7073, N15084, N9729);
and AND2 (N16027, N16025, N9777);
or OR2 (N16028, N16021, N6053);
buf BUF1 (N16029, N16028);
xor XOR2 (N16030, N16016, N899);
or OR3 (N16031, N16026, N4916, N10403);
nor NOR4 (N16032, N16029, N8573, N14251, N9143);
or OR2 (N16033, N16011, N3405);
or OR2 (N16034, N16027, N6497);
nand NAND2 (N16035, N16032, N15622);
nor NOR4 (N16036, N16015, N8983, N8661, N1121);
nand NAND2 (N16037, N16020, N2512);
nor NOR2 (N16038, N16033, N14890);
buf BUF1 (N16039, N16035);
not NOT1 (N16040, N16023);
and AND3 (N16041, N16031, N11215, N5574);
buf BUF1 (N16042, N16024);
nand NAND4 (N16043, N16038, N6349, N9149, N14305);
or OR4 (N16044, N16022, N4215, N7162, N1504);
and AND4 (N16045, N16034, N13892, N3914, N5843);
and AND3 (N16046, N16040, N10321, N9);
nand NAND3 (N16047, N16043, N9874, N9680);
and AND2 (N16048, N16037, N10598);
nor NOR3 (N16049, N16045, N11934, N2294);
xor XOR2 (N16050, N16047, N642);
xor XOR2 (N16051, N16030, N13139);
or OR3 (N16052, N16048, N1312, N10268);
nand NAND4 (N16053, N16039, N12823, N8394, N12786);
xor XOR2 (N16054, N16041, N16013);
buf BUF1 (N16055, N16042);
buf BUF1 (N16056, N16054);
buf BUF1 (N16057, N16053);
or OR2 (N16058, N16046, N3314);
and AND4 (N16059, N16057, N9068, N8437, N2726);
buf BUF1 (N16060, N16049);
xor XOR2 (N16061, N16056, N3977);
and AND3 (N16062, N16060, N5395, N15908);
nand NAND3 (N16063, N16058, N4995, N14885);
nand NAND3 (N16064, N16061, N4427, N13826);
and AND3 (N16065, N16052, N10274, N15050);
nor NOR4 (N16066, N16036, N11004, N3168, N13103);
and AND4 (N16067, N16055, N7551, N12185, N12054);
or OR4 (N16068, N16064, N4055, N5117, N194);
or OR2 (N16069, N16065, N9248);
buf BUF1 (N16070, N16068);
and AND4 (N16071, N16069, N13940, N9001, N4322);
not NOT1 (N16072, N16051);
nor NOR2 (N16073, N16063, N14426);
not NOT1 (N16074, N16073);
not NOT1 (N16075, N16071);
nor NOR2 (N16076, N16050, N13640);
nor NOR3 (N16077, N16074, N10743, N4659);
xor XOR2 (N16078, N16075, N1169);
or OR3 (N16079, N16059, N5980, N7332);
not NOT1 (N16080, N16077);
or OR3 (N16081, N16076, N12864, N5191);
nor NOR2 (N16082, N16078, N4973);
or OR2 (N16083, N16062, N6374);
buf BUF1 (N16084, N16082);
xor XOR2 (N16085, N16072, N4441);
nor NOR3 (N16086, N16085, N13575, N11554);
or OR2 (N16087, N16080, N10621);
or OR4 (N16088, N16081, N15369, N11612, N3541);
or OR4 (N16089, N16044, N12213, N5634, N1430);
or OR3 (N16090, N16089, N3926, N1172);
nand NAND2 (N16091, N16088, N4990);
nor NOR3 (N16092, N16091, N13584, N47);
not NOT1 (N16093, N16079);
nand NAND4 (N16094, N16067, N3473, N14716, N9596);
xor XOR2 (N16095, N16084, N336);
nor NOR2 (N16096, N16094, N3209);
or OR2 (N16097, N16092, N13547);
not NOT1 (N16098, N16097);
nor NOR3 (N16099, N16087, N9103, N3477);
not NOT1 (N16100, N16098);
nor NOR2 (N16101, N16083, N14148);
and AND4 (N16102, N16100, N3530, N9860, N15385);
not NOT1 (N16103, N16101);
buf BUF1 (N16104, N16070);
xor XOR2 (N16105, N16095, N11603);
xor XOR2 (N16106, N16102, N10665);
or OR2 (N16107, N16099, N3749);
nor NOR3 (N16108, N16066, N7999, N8112);
nand NAND4 (N16109, N16104, N10591, N11563, N13424);
nor NOR2 (N16110, N16103, N2041);
nor NOR2 (N16111, N16090, N7679);
nor NOR2 (N16112, N16105, N14093);
or OR3 (N16113, N16086, N13176, N6163);
and AND3 (N16114, N16096, N5068, N12823);
and AND2 (N16115, N16113, N10815);
nor NOR2 (N16116, N16112, N2820);
nand NAND3 (N16117, N16107, N1738, N13607);
buf BUF1 (N16118, N16108);
and AND2 (N16119, N16109, N11232);
nand NAND4 (N16120, N16093, N6932, N4107, N2448);
nand NAND2 (N16121, N16118, N13398);
not NOT1 (N16122, N16117);
and AND2 (N16123, N16115, N8852);
xor XOR2 (N16124, N16114, N12407);
not NOT1 (N16125, N16121);
nand NAND2 (N16126, N16124, N9966);
xor XOR2 (N16127, N16110, N10190);
xor XOR2 (N16128, N16111, N3526);
nor NOR2 (N16129, N16125, N7185);
xor XOR2 (N16130, N16120, N13580);
not NOT1 (N16131, N16119);
and AND4 (N16132, N16122, N4479, N6480, N14130);
nor NOR3 (N16133, N16116, N2037, N6332);
nor NOR2 (N16134, N16106, N8455);
buf BUF1 (N16135, N16127);
nand NAND2 (N16136, N16133, N8460);
buf BUF1 (N16137, N16136);
buf BUF1 (N16138, N16131);
xor XOR2 (N16139, N16128, N5111);
xor XOR2 (N16140, N16129, N879);
xor XOR2 (N16141, N16139, N1402);
buf BUF1 (N16142, N16140);
and AND4 (N16143, N16137, N952, N4603, N13050);
nor NOR3 (N16144, N16130, N13608, N5531);
nand NAND2 (N16145, N16142, N13250);
not NOT1 (N16146, N16144);
not NOT1 (N16147, N16134);
xor XOR2 (N16148, N16143, N7440);
and AND4 (N16149, N16148, N3082, N585, N826);
nand NAND4 (N16150, N16126, N12194, N14130, N1181);
nor NOR4 (N16151, N16150, N13483, N15209, N15860);
and AND4 (N16152, N16151, N10169, N10877, N10451);
and AND2 (N16153, N16132, N3258);
nand NAND4 (N16154, N16145, N1866, N12792, N15282);
nand NAND3 (N16155, N16123, N5082, N11702);
nand NAND3 (N16156, N16147, N13198, N8575);
nor NOR2 (N16157, N16155, N6983);
not NOT1 (N16158, N16146);
buf BUF1 (N16159, N16141);
buf BUF1 (N16160, N16153);
or OR3 (N16161, N16152, N2122, N15091);
xor XOR2 (N16162, N16161, N1622);
and AND3 (N16163, N16159, N13532, N12698);
buf BUF1 (N16164, N16163);
not NOT1 (N16165, N16160);
not NOT1 (N16166, N16164);
or OR4 (N16167, N16156, N15828, N10884, N15299);
nand NAND3 (N16168, N16154, N10355, N5301);
not NOT1 (N16169, N16138);
nand NAND2 (N16170, N16162, N6840);
or OR3 (N16171, N16169, N7970, N9159);
not NOT1 (N16172, N16157);
not NOT1 (N16173, N16149);
buf BUF1 (N16174, N16172);
nand NAND3 (N16175, N16167, N12909, N2971);
nand NAND2 (N16176, N16173, N4556);
nor NOR2 (N16177, N16170, N10597);
and AND2 (N16178, N16135, N15525);
not NOT1 (N16179, N16165);
and AND2 (N16180, N16158, N15219);
or OR3 (N16181, N16180, N3889, N14556);
nor NOR4 (N16182, N16171, N7800, N1110, N7233);
nor NOR2 (N16183, N16177, N4253);
and AND3 (N16184, N16179, N7438, N13531);
buf BUF1 (N16185, N16166);
not NOT1 (N16186, N16185);
xor XOR2 (N16187, N16168, N9858);
xor XOR2 (N16188, N16182, N7312);
and AND2 (N16189, N16174, N10286);
nor NOR2 (N16190, N16188, N11504);
not NOT1 (N16191, N16175);
nand NAND4 (N16192, N16183, N12750, N8632, N7857);
or OR2 (N16193, N16178, N14373);
not NOT1 (N16194, N16192);
xor XOR2 (N16195, N16186, N8186);
xor XOR2 (N16196, N16176, N15012);
and AND4 (N16197, N16187, N7626, N13029, N7572);
buf BUF1 (N16198, N16196);
xor XOR2 (N16199, N16197, N10848);
buf BUF1 (N16200, N16193);
xor XOR2 (N16201, N16184, N3738);
buf BUF1 (N16202, N16194);
or OR2 (N16203, N16200, N14517);
nand NAND4 (N16204, N16190, N11073, N14084, N15933);
nand NAND4 (N16205, N16199, N3347, N15162, N16185);
and AND3 (N16206, N16189, N10892, N12906);
not NOT1 (N16207, N16198);
xor XOR2 (N16208, N16203, N15718);
nand NAND3 (N16209, N16204, N4347, N9129);
xor XOR2 (N16210, N16206, N5276);
not NOT1 (N16211, N16195);
or OR2 (N16212, N16201, N5219);
xor XOR2 (N16213, N16208, N14972);
nand NAND4 (N16214, N16207, N6626, N15274, N11820);
or OR4 (N16215, N16181, N10966, N4619, N7396);
buf BUF1 (N16216, N16215);
xor XOR2 (N16217, N16213, N16019);
nor NOR2 (N16218, N16216, N12581);
or OR2 (N16219, N16218, N6441);
nor NOR2 (N16220, N16217, N8875);
and AND2 (N16221, N16212, N14355);
xor XOR2 (N16222, N16219, N15563);
not NOT1 (N16223, N16220);
not NOT1 (N16224, N16223);
nor NOR4 (N16225, N16224, N3165, N1587, N6860);
not NOT1 (N16226, N16202);
nor NOR4 (N16227, N16205, N4511, N5736, N11764);
xor XOR2 (N16228, N16222, N8891);
or OR3 (N16229, N16214, N1314, N98);
and AND2 (N16230, N16226, N3553);
or OR3 (N16231, N16227, N11552, N816);
xor XOR2 (N16232, N16229, N4779);
buf BUF1 (N16233, N16211);
nand NAND4 (N16234, N16225, N9387, N176, N13257);
nor NOR4 (N16235, N16210, N12163, N11983, N4580);
not NOT1 (N16236, N16231);
and AND4 (N16237, N16232, N11617, N5399, N10621);
nand NAND3 (N16238, N16209, N5442, N13110);
buf BUF1 (N16239, N16234);
xor XOR2 (N16240, N16238, N2070);
nor NOR2 (N16241, N16233, N2278);
or OR3 (N16242, N16221, N7070, N15064);
nor NOR2 (N16243, N16242, N5172);
xor XOR2 (N16244, N16228, N8212);
xor XOR2 (N16245, N16236, N2706);
buf BUF1 (N16246, N16235);
not NOT1 (N16247, N16246);
and AND2 (N16248, N16239, N2403);
xor XOR2 (N16249, N16240, N2890);
or OR4 (N16250, N16248, N14448, N2176, N13978);
buf BUF1 (N16251, N16250);
buf BUF1 (N16252, N16191);
nor NOR2 (N16253, N16247, N15269);
nor NOR4 (N16254, N16249, N3783, N10753, N1882);
not NOT1 (N16255, N16230);
nor NOR2 (N16256, N16245, N2073);
not NOT1 (N16257, N16251);
not NOT1 (N16258, N16241);
xor XOR2 (N16259, N16257, N10373);
nand NAND4 (N16260, N16258, N1092, N6683, N2402);
nand NAND2 (N16261, N16259, N719);
xor XOR2 (N16262, N16254, N11525);
and AND4 (N16263, N16261, N7684, N3563, N9869);
not NOT1 (N16264, N16262);
not NOT1 (N16265, N16243);
xor XOR2 (N16266, N16264, N4286);
and AND4 (N16267, N16252, N3944, N7045, N8276);
buf BUF1 (N16268, N16253);
and AND2 (N16269, N16255, N994);
or OR3 (N16270, N16268, N619, N6533);
and AND4 (N16271, N16267, N6061, N6847, N15837);
not NOT1 (N16272, N16265);
xor XOR2 (N16273, N16244, N16053);
or OR3 (N16274, N16271, N6044, N11579);
xor XOR2 (N16275, N16266, N12328);
not NOT1 (N16276, N16270);
xor XOR2 (N16277, N16260, N5952);
and AND4 (N16278, N16277, N1732, N3309, N10666);
buf BUF1 (N16279, N16263);
nor NOR2 (N16280, N16269, N6423);
not NOT1 (N16281, N16272);
nand NAND3 (N16282, N16276, N7515, N10773);
nand NAND2 (N16283, N16282, N321);
xor XOR2 (N16284, N16274, N4940);
nor NOR3 (N16285, N16237, N946, N15354);
and AND4 (N16286, N16283, N6639, N764, N13340);
and AND2 (N16287, N16280, N14931);
or OR2 (N16288, N16285, N3784);
and AND4 (N16289, N16275, N6349, N440, N9447);
xor XOR2 (N16290, N16289, N8839);
not NOT1 (N16291, N16288);
nor NOR4 (N16292, N16278, N15551, N11843, N964);
nor NOR2 (N16293, N16286, N15175);
not NOT1 (N16294, N16290);
nand NAND2 (N16295, N16281, N10486);
and AND4 (N16296, N16292, N12552, N6878, N4427);
xor XOR2 (N16297, N16287, N8164);
nand NAND2 (N16298, N16291, N197);
or OR3 (N16299, N16279, N9966, N8823);
or OR3 (N16300, N16298, N8073, N8407);
or OR4 (N16301, N16284, N2891, N12220, N3806);
or OR2 (N16302, N16294, N10011);
not NOT1 (N16303, N16299);
buf BUF1 (N16304, N16273);
and AND2 (N16305, N16295, N13620);
nor NOR2 (N16306, N16302, N4894);
buf BUF1 (N16307, N16293);
or OR2 (N16308, N16256, N10434);
and AND2 (N16309, N16305, N10065);
buf BUF1 (N16310, N16307);
xor XOR2 (N16311, N16301, N8862);
nand NAND2 (N16312, N16309, N3750);
and AND2 (N16313, N16303, N15763);
nor NOR4 (N16314, N16304, N2711, N4236, N12731);
nand NAND3 (N16315, N16297, N8373, N8420);
not NOT1 (N16316, N16311);
not NOT1 (N16317, N16310);
not NOT1 (N16318, N16296);
nor NOR3 (N16319, N16306, N10819, N13213);
nand NAND4 (N16320, N16318, N10177, N13268, N9172);
xor XOR2 (N16321, N16300, N894);
and AND4 (N16322, N16314, N7508, N864, N8769);
not NOT1 (N16323, N16317);
buf BUF1 (N16324, N16323);
nand NAND2 (N16325, N16322, N14081);
or OR4 (N16326, N16325, N9344, N9845, N919);
nor NOR3 (N16327, N16316, N10848, N8550);
or OR2 (N16328, N16308, N2548);
xor XOR2 (N16329, N16324, N6467);
or OR2 (N16330, N16321, N9647);
nor NOR4 (N16331, N16312, N1549, N9914, N10526);
nor NOR3 (N16332, N16313, N13456, N2604);
not NOT1 (N16333, N16328);
or OR2 (N16334, N16327, N15106);
or OR2 (N16335, N16332, N5371);
nand NAND2 (N16336, N16333, N13029);
not NOT1 (N16337, N16315);
nor NOR2 (N16338, N16319, N14871);
and AND2 (N16339, N16338, N69);
nor NOR4 (N16340, N16329, N5641, N15287, N6182);
buf BUF1 (N16341, N16320);
nor NOR4 (N16342, N16330, N12108, N766, N12339);
not NOT1 (N16343, N16326);
nand NAND3 (N16344, N16334, N9742, N14316);
nand NAND2 (N16345, N16336, N16069);
nand NAND3 (N16346, N16331, N12038, N14772);
buf BUF1 (N16347, N16343);
nand NAND2 (N16348, N16339, N12990);
or OR3 (N16349, N16340, N6520, N9006);
or OR2 (N16350, N16349, N9928);
xor XOR2 (N16351, N16342, N14088);
and AND2 (N16352, N16344, N16250);
nand NAND4 (N16353, N16351, N7899, N15421, N4659);
and AND2 (N16354, N16350, N8510);
nor NOR3 (N16355, N16354, N2627, N7370);
or OR3 (N16356, N16355, N15671, N4572);
xor XOR2 (N16357, N16352, N3091);
nor NOR4 (N16358, N16353, N3537, N15886, N12594);
xor XOR2 (N16359, N16337, N1477);
nand NAND2 (N16360, N16335, N6418);
xor XOR2 (N16361, N16360, N11648);
and AND2 (N16362, N16346, N2234);
nand NAND3 (N16363, N16356, N9657, N2847);
nand NAND2 (N16364, N16348, N8541);
nand NAND2 (N16365, N16347, N10659);
buf BUF1 (N16366, N16358);
nor NOR4 (N16367, N16362, N9853, N12263, N5172);
and AND3 (N16368, N16363, N5046, N11047);
and AND4 (N16369, N16359, N9864, N6673, N3596);
not NOT1 (N16370, N16367);
nor NOR4 (N16371, N16368, N1585, N6657, N15645);
and AND3 (N16372, N16364, N14732, N14630);
xor XOR2 (N16373, N16366, N4343);
nor NOR3 (N16374, N16357, N11527, N14811);
xor XOR2 (N16375, N16373, N5255);
nor NOR2 (N16376, N16375, N682);
not NOT1 (N16377, N16361);
or OR2 (N16378, N16370, N14330);
nand NAND2 (N16379, N16365, N8254);
xor XOR2 (N16380, N16341, N11132);
nand NAND4 (N16381, N16377, N10629, N15896, N10339);
not NOT1 (N16382, N16379);
nand NAND2 (N16383, N16369, N6706);
nor NOR2 (N16384, N16372, N4205);
nor NOR4 (N16385, N16376, N14692, N4734, N5245);
and AND3 (N16386, N16380, N7521, N481);
nor NOR4 (N16387, N16386, N3310, N13368, N13073);
xor XOR2 (N16388, N16385, N8673);
buf BUF1 (N16389, N16371);
xor XOR2 (N16390, N16384, N1711);
nor NOR4 (N16391, N16387, N1308, N2887, N15493);
nor NOR3 (N16392, N16388, N4912, N3652);
buf BUF1 (N16393, N16383);
nor NOR3 (N16394, N16391, N8682, N10099);
not NOT1 (N16395, N16390);
not NOT1 (N16396, N16395);
and AND3 (N16397, N16396, N16248, N3485);
or OR3 (N16398, N16374, N9974, N7729);
and AND3 (N16399, N16392, N6656, N4632);
and AND4 (N16400, N16399, N1424, N14717, N9344);
or OR2 (N16401, N16394, N8975);
and AND4 (N16402, N16393, N8235, N5545, N3130);
buf BUF1 (N16403, N16398);
nand NAND4 (N16404, N16381, N4187, N4293, N11869);
nand NAND4 (N16405, N16382, N2976, N14236, N14056);
and AND3 (N16406, N16400, N3539, N13658);
xor XOR2 (N16407, N16405, N9759);
not NOT1 (N16408, N16407);
xor XOR2 (N16409, N16402, N3396);
xor XOR2 (N16410, N16389, N3593);
not NOT1 (N16411, N16406);
nand NAND4 (N16412, N16411, N755, N8395, N6715);
and AND4 (N16413, N16408, N603, N954, N7426);
or OR4 (N16414, N16404, N10288, N12962, N14916);
not NOT1 (N16415, N16401);
not NOT1 (N16416, N16403);
and AND4 (N16417, N16397, N8335, N444, N6091);
buf BUF1 (N16418, N16378);
not NOT1 (N16419, N16409);
xor XOR2 (N16420, N16345, N11153);
xor XOR2 (N16421, N16414, N4258);
nor NOR3 (N16422, N16413, N14235, N15973);
nor NOR4 (N16423, N16421, N396, N16296, N3887);
nor NOR4 (N16424, N16410, N13066, N12662, N8841);
nand NAND4 (N16425, N16416, N13629, N3631, N6587);
and AND2 (N16426, N16415, N10890);
or OR2 (N16427, N16424, N5937);
or OR2 (N16428, N16418, N4289);
buf BUF1 (N16429, N16412);
not NOT1 (N16430, N16425);
or OR2 (N16431, N16423, N10731);
or OR4 (N16432, N16426, N7700, N10433, N11208);
nor NOR2 (N16433, N16431, N8434);
or OR3 (N16434, N16419, N9344, N15659);
xor XOR2 (N16435, N16428, N12081);
nor NOR2 (N16436, N16432, N9515);
and AND4 (N16437, N16427, N11255, N6612, N12297);
or OR4 (N16438, N16417, N10576, N6438, N2308);
buf BUF1 (N16439, N16422);
nand NAND3 (N16440, N16438, N15858, N11354);
not NOT1 (N16441, N16430);
nor NOR2 (N16442, N16439, N13357);
buf BUF1 (N16443, N16436);
not NOT1 (N16444, N16443);
nand NAND4 (N16445, N16435, N10547, N7204, N7088);
not NOT1 (N16446, N16434);
buf BUF1 (N16447, N16429);
buf BUF1 (N16448, N16433);
nor NOR4 (N16449, N16441, N4278, N8175, N1794);
or OR2 (N16450, N16444, N11541);
and AND2 (N16451, N16448, N2011);
nand NAND3 (N16452, N16450, N14592, N3779);
not NOT1 (N16453, N16442);
nand NAND2 (N16454, N16445, N8312);
not NOT1 (N16455, N16449);
or OR2 (N16456, N16446, N2222);
not NOT1 (N16457, N16456);
buf BUF1 (N16458, N16447);
buf BUF1 (N16459, N16454);
or OR4 (N16460, N16437, N14173, N5027, N13057);
or OR2 (N16461, N16457, N7076);
not NOT1 (N16462, N16458);
xor XOR2 (N16463, N16440, N2290);
and AND2 (N16464, N16452, N1779);
and AND3 (N16465, N16453, N9436, N15663);
buf BUF1 (N16466, N16455);
not NOT1 (N16467, N16451);
not NOT1 (N16468, N16463);
or OR3 (N16469, N16466, N16176, N13217);
xor XOR2 (N16470, N16459, N5605);
and AND2 (N16471, N16462, N1566);
buf BUF1 (N16472, N16420);
or OR3 (N16473, N16471, N14841, N6489);
not NOT1 (N16474, N16468);
and AND4 (N16475, N16472, N4093, N10973, N3779);
nor NOR4 (N16476, N16460, N5419, N12835, N863);
buf BUF1 (N16477, N16461);
not NOT1 (N16478, N16469);
xor XOR2 (N16479, N16475, N4093);
buf BUF1 (N16480, N16473);
nand NAND2 (N16481, N16480, N6384);
and AND3 (N16482, N16465, N6527, N4092);
or OR3 (N16483, N16482, N12923, N3709);
not NOT1 (N16484, N16470);
xor XOR2 (N16485, N16478, N5880);
xor XOR2 (N16486, N16467, N13576);
and AND4 (N16487, N16483, N16181, N7900, N5562);
not NOT1 (N16488, N16476);
and AND2 (N16489, N16488, N11497);
buf BUF1 (N16490, N16487);
nand NAND4 (N16491, N16479, N4558, N2871, N3386);
xor XOR2 (N16492, N16491, N7631);
not NOT1 (N16493, N16474);
and AND2 (N16494, N16485, N14494);
xor XOR2 (N16495, N16486, N12487);
and AND4 (N16496, N16477, N10748, N1881, N366);
xor XOR2 (N16497, N16481, N13638);
nand NAND2 (N16498, N16464, N15041);
nand NAND2 (N16499, N16496, N5350);
nor NOR4 (N16500, N16489, N9245, N15006, N9244);
or OR2 (N16501, N16484, N4605);
or OR4 (N16502, N16495, N9720, N5441, N8303);
nand NAND2 (N16503, N16501, N5964);
buf BUF1 (N16504, N16497);
nand NAND3 (N16505, N16504, N12881, N5593);
not NOT1 (N16506, N16493);
not NOT1 (N16507, N16492);
not NOT1 (N16508, N16499);
buf BUF1 (N16509, N16490);
nor NOR4 (N16510, N16509, N8640, N16482, N15798);
xor XOR2 (N16511, N16500, N10918);
and AND3 (N16512, N16503, N15694, N2854);
or OR2 (N16513, N16512, N15861);
and AND4 (N16514, N16502, N13036, N15656, N10610);
buf BUF1 (N16515, N16511);
nor NOR3 (N16516, N16507, N3387, N15854);
not NOT1 (N16517, N16505);
buf BUF1 (N16518, N16517);
buf BUF1 (N16519, N16508);
not NOT1 (N16520, N16510);
xor XOR2 (N16521, N16515, N1792);
not NOT1 (N16522, N16520);
nand NAND3 (N16523, N16521, N14931, N12923);
and AND2 (N16524, N16498, N4852);
xor XOR2 (N16525, N16514, N13480);
nor NOR2 (N16526, N16506, N11177);
xor XOR2 (N16527, N16494, N2908);
and AND2 (N16528, N16523, N13754);
not NOT1 (N16529, N16513);
buf BUF1 (N16530, N16518);
nor NOR3 (N16531, N16524, N14362, N15693);
nand NAND3 (N16532, N16528, N5784, N14193);
and AND2 (N16533, N16532, N9451);
and AND2 (N16534, N16533, N6237);
nor NOR3 (N16535, N16525, N1112, N6967);
nor NOR3 (N16536, N16527, N5856, N10164);
buf BUF1 (N16537, N16531);
not NOT1 (N16538, N16535);
nor NOR3 (N16539, N16530, N3712, N4337);
or OR3 (N16540, N16516, N669, N14037);
not NOT1 (N16541, N16538);
and AND4 (N16542, N16529, N11894, N4031, N1148);
buf BUF1 (N16543, N16542);
nand NAND4 (N16544, N16541, N4551, N10601, N4650);
not NOT1 (N16545, N16544);
xor XOR2 (N16546, N16522, N16282);
or OR2 (N16547, N16543, N12917);
nor NOR3 (N16548, N16539, N4531, N6687);
not NOT1 (N16549, N16534);
not NOT1 (N16550, N16537);
buf BUF1 (N16551, N16540);
or OR3 (N16552, N16536, N1326, N9320);
not NOT1 (N16553, N16519);
nor NOR3 (N16554, N16552, N3819, N15126);
and AND3 (N16555, N16549, N5780, N5446);
not NOT1 (N16556, N16546);
buf BUF1 (N16557, N16548);
nor NOR4 (N16558, N16547, N754, N9868, N12183);
nor NOR4 (N16559, N16556, N4426, N12629, N8301);
and AND4 (N16560, N16545, N7256, N3546, N8858);
not NOT1 (N16561, N16555);
nor NOR2 (N16562, N16558, N6845);
xor XOR2 (N16563, N16557, N14861);
nor NOR4 (N16564, N16553, N961, N8252, N2281);
buf BUF1 (N16565, N16551);
buf BUF1 (N16566, N16564);
or OR2 (N16567, N16559, N14926);
not NOT1 (N16568, N16554);
not NOT1 (N16569, N16526);
buf BUF1 (N16570, N16565);
or OR4 (N16571, N16567, N2402, N15648, N8955);
nand NAND3 (N16572, N16566, N5262, N10892);
or OR3 (N16573, N16550, N5816, N3530);
not NOT1 (N16574, N16560);
nand NAND3 (N16575, N16574, N10645, N11557);
nand NAND3 (N16576, N16563, N1645, N9941);
nor NOR3 (N16577, N16576, N9068, N13679);
buf BUF1 (N16578, N16570);
buf BUF1 (N16579, N16569);
xor XOR2 (N16580, N16568, N7178);
xor XOR2 (N16581, N16575, N16333);
xor XOR2 (N16582, N16572, N10261);
not NOT1 (N16583, N16573);
nand NAND3 (N16584, N16577, N4494, N1005);
nand NAND2 (N16585, N16562, N3591);
nand NAND3 (N16586, N16581, N14788, N8652);
xor XOR2 (N16587, N16571, N14316);
nand NAND2 (N16588, N16585, N3797);
not NOT1 (N16589, N16580);
nand NAND3 (N16590, N16587, N15055, N14695);
and AND4 (N16591, N16586, N13800, N5852, N1180);
and AND3 (N16592, N16561, N3064, N2122);
nor NOR2 (N16593, N16591, N14537);
buf BUF1 (N16594, N16588);
xor XOR2 (N16595, N16593, N15841);
xor XOR2 (N16596, N16579, N2426);
nor NOR2 (N16597, N16578, N10525);
not NOT1 (N16598, N16584);
not NOT1 (N16599, N16590);
or OR2 (N16600, N16582, N4464);
buf BUF1 (N16601, N16598);
nor NOR2 (N16602, N16599, N13196);
not NOT1 (N16603, N16594);
not NOT1 (N16604, N16595);
nor NOR3 (N16605, N16589, N2137, N4850);
buf BUF1 (N16606, N16602);
or OR4 (N16607, N16603, N13640, N736, N1481);
or OR3 (N16608, N16600, N6182, N3214);
or OR2 (N16609, N16601, N13762);
nand NAND2 (N16610, N16583, N2137);
not NOT1 (N16611, N16610);
not NOT1 (N16612, N16604);
not NOT1 (N16613, N16608);
or OR3 (N16614, N16596, N2177, N4981);
not NOT1 (N16615, N16597);
and AND3 (N16616, N16611, N11712, N1819);
nor NOR3 (N16617, N16613, N7255, N12684);
or OR2 (N16618, N16606, N7038);
xor XOR2 (N16619, N16617, N11);
xor XOR2 (N16620, N16609, N689);
not NOT1 (N16621, N16618);
not NOT1 (N16622, N16619);
or OR3 (N16623, N16614, N6695, N14985);
or OR4 (N16624, N16612, N5435, N1835, N1542);
xor XOR2 (N16625, N16620, N9132);
buf BUF1 (N16626, N16624);
buf BUF1 (N16627, N16605);
nor NOR3 (N16628, N16616, N14959, N10601);
nand NAND4 (N16629, N16621, N15302, N7500, N8689);
or OR4 (N16630, N16625, N5815, N12589, N1571);
buf BUF1 (N16631, N16627);
nor NOR3 (N16632, N16631, N3399, N85);
or OR2 (N16633, N16632, N10835);
not NOT1 (N16634, N16630);
and AND2 (N16635, N16629, N12617);
xor XOR2 (N16636, N16592, N12067);
buf BUF1 (N16637, N16622);
and AND2 (N16638, N16626, N14285);
nor NOR4 (N16639, N16633, N10422, N332, N8852);
or OR4 (N16640, N16635, N4140, N5226, N5575);
and AND3 (N16641, N16615, N9230, N15963);
xor XOR2 (N16642, N16640, N9197);
nand NAND3 (N16643, N16628, N15338, N16403);
not NOT1 (N16644, N16639);
or OR3 (N16645, N16637, N2606, N12437);
nor NOR3 (N16646, N16607, N298, N12905);
buf BUF1 (N16647, N16641);
and AND4 (N16648, N16623, N10471, N4108, N1339);
not NOT1 (N16649, N16645);
buf BUF1 (N16650, N16636);
or OR2 (N16651, N16638, N4645);
nor NOR2 (N16652, N16634, N2785);
or OR4 (N16653, N16642, N12686, N13371, N13259);
buf BUF1 (N16654, N16651);
xor XOR2 (N16655, N16644, N8252);
nor NOR4 (N16656, N16646, N3480, N13026, N11774);
or OR3 (N16657, N16650, N1385, N12629);
nand NAND4 (N16658, N16653, N5646, N16525, N11604);
buf BUF1 (N16659, N16647);
or OR3 (N16660, N16656, N15105, N7544);
nor NOR4 (N16661, N16648, N1071, N14901, N7371);
nand NAND4 (N16662, N16657, N10724, N14322, N985);
nor NOR4 (N16663, N16658, N351, N15473, N15814);
and AND2 (N16664, N16661, N4360);
nand NAND2 (N16665, N16643, N1492);
not NOT1 (N16666, N16662);
buf BUF1 (N16667, N16654);
buf BUF1 (N16668, N16655);
not NOT1 (N16669, N16664);
nor NOR3 (N16670, N16660, N16472, N15649);
and AND3 (N16671, N16669, N6957, N16317);
nand NAND3 (N16672, N16649, N13167, N10007);
buf BUF1 (N16673, N16666);
not NOT1 (N16674, N16659);
not NOT1 (N16675, N16673);
nor NOR2 (N16676, N16665, N15240);
xor XOR2 (N16677, N16670, N8326);
buf BUF1 (N16678, N16672);
nor NOR2 (N16679, N16676, N11082);
and AND4 (N16680, N16668, N14926, N16655, N2848);
buf BUF1 (N16681, N16680);
xor XOR2 (N16682, N16677, N12974);
or OR4 (N16683, N16674, N5306, N12161, N6336);
buf BUF1 (N16684, N16678);
buf BUF1 (N16685, N16667);
not NOT1 (N16686, N16683);
not NOT1 (N16687, N16684);
xor XOR2 (N16688, N16652, N796);
not NOT1 (N16689, N16685);
xor XOR2 (N16690, N16689, N9864);
buf BUF1 (N16691, N16687);
xor XOR2 (N16692, N16688, N11589);
not NOT1 (N16693, N16682);
nand NAND4 (N16694, N16692, N9177, N3631, N5107);
nand NAND4 (N16695, N16681, N14732, N4256, N11873);
not NOT1 (N16696, N16690);
and AND4 (N16697, N16675, N3191, N3321, N5550);
and AND2 (N16698, N16697, N2113);
not NOT1 (N16699, N16695);
nor NOR2 (N16700, N16693, N10802);
nand NAND3 (N16701, N16663, N9740, N10819);
and AND4 (N16702, N16679, N16116, N13433, N5452);
xor XOR2 (N16703, N16699, N7866);
nor NOR3 (N16704, N16696, N3550, N1472);
and AND4 (N16705, N16698, N9280, N10503, N7752);
and AND3 (N16706, N16702, N8771, N10873);
buf BUF1 (N16707, N16700);
nand NAND2 (N16708, N16701, N11154);
nand NAND2 (N16709, N16691, N8816);
not NOT1 (N16710, N16703);
nor NOR4 (N16711, N16694, N1837, N15843, N7346);
or OR2 (N16712, N16710, N9641);
and AND3 (N16713, N16705, N2564, N10163);
xor XOR2 (N16714, N16711, N10502);
buf BUF1 (N16715, N16708);
nand NAND3 (N16716, N16707, N6962, N2280);
nor NOR3 (N16717, N16714, N918, N14059);
not NOT1 (N16718, N16709);
nand NAND4 (N16719, N16716, N13621, N9205, N10564);
buf BUF1 (N16720, N16704);
or OR2 (N16721, N16713, N11270);
buf BUF1 (N16722, N16715);
not NOT1 (N16723, N16719);
and AND4 (N16724, N16706, N12321, N1015, N991);
nor NOR3 (N16725, N16721, N16259, N11004);
or OR3 (N16726, N16723, N4328, N13911);
not NOT1 (N16727, N16671);
xor XOR2 (N16728, N16725, N11078);
xor XOR2 (N16729, N16728, N1664);
buf BUF1 (N16730, N16718);
and AND3 (N16731, N16727, N2188, N5234);
not NOT1 (N16732, N16731);
nand NAND2 (N16733, N16712, N8485);
or OR3 (N16734, N16732, N9917, N452);
buf BUF1 (N16735, N16720);
nand NAND2 (N16736, N16735, N11032);
xor XOR2 (N16737, N16730, N3607);
nor NOR3 (N16738, N16724, N6792, N226);
buf BUF1 (N16739, N16717);
nand NAND2 (N16740, N16729, N4677);
not NOT1 (N16741, N16737);
not NOT1 (N16742, N16741);
not NOT1 (N16743, N16738);
xor XOR2 (N16744, N16722, N6171);
nand NAND3 (N16745, N16740, N9769, N6557);
and AND3 (N16746, N16733, N761, N16450);
nor NOR4 (N16747, N16686, N11933, N6289, N554);
nor NOR3 (N16748, N16745, N4834, N7743);
not NOT1 (N16749, N16748);
and AND3 (N16750, N16739, N3048, N6797);
buf BUF1 (N16751, N16726);
xor XOR2 (N16752, N16736, N233);
or OR4 (N16753, N16742, N9063, N217, N12038);
and AND3 (N16754, N16749, N11751, N12173);
xor XOR2 (N16755, N16744, N4466);
not NOT1 (N16756, N16743);
buf BUF1 (N16757, N16756);
or OR3 (N16758, N16751, N302, N6252);
not NOT1 (N16759, N16755);
not NOT1 (N16760, N16752);
or OR4 (N16761, N16760, N16350, N4418, N14834);
not NOT1 (N16762, N16750);
and AND2 (N16763, N16746, N1538);
and AND3 (N16764, N16762, N5726, N2333);
not NOT1 (N16765, N16763);
nand NAND3 (N16766, N16765, N10079, N11712);
or OR3 (N16767, N16758, N16497, N5017);
nor NOR2 (N16768, N16766, N11472);
or OR2 (N16769, N16747, N9958);
xor XOR2 (N16770, N16754, N1522);
nand NAND2 (N16771, N16770, N2375);
nor NOR3 (N16772, N16767, N8800, N15393);
buf BUF1 (N16773, N16753);
nand NAND2 (N16774, N16769, N1903);
xor XOR2 (N16775, N16773, N7853);
and AND3 (N16776, N16775, N2296, N7151);
buf BUF1 (N16777, N16759);
buf BUF1 (N16778, N16764);
or OR4 (N16779, N16777, N6405, N5031, N3040);
or OR2 (N16780, N16771, N8405);
xor XOR2 (N16781, N16780, N7266);
nand NAND2 (N16782, N16774, N3883);
xor XOR2 (N16783, N16776, N11560);
nand NAND2 (N16784, N16783, N12533);
xor XOR2 (N16785, N16784, N2147);
and AND4 (N16786, N16768, N3417, N13025, N15127);
or OR3 (N16787, N16779, N10949, N16422);
buf BUF1 (N16788, N16778);
nor NOR3 (N16789, N16781, N11841, N1392);
and AND4 (N16790, N16757, N3418, N7654, N899);
xor XOR2 (N16791, N16734, N8077);
xor XOR2 (N16792, N16788, N3287);
or OR2 (N16793, N16786, N13607);
or OR3 (N16794, N16772, N13376, N16146);
nand NAND2 (N16795, N16791, N4083);
not NOT1 (N16796, N16793);
xor XOR2 (N16797, N16795, N6186);
nor NOR3 (N16798, N16761, N897, N5360);
not NOT1 (N16799, N16796);
or OR3 (N16800, N16782, N7254, N5266);
not NOT1 (N16801, N16797);
nor NOR2 (N16802, N16792, N2820);
nand NAND2 (N16803, N16794, N7113);
xor XOR2 (N16804, N16801, N5198);
nor NOR4 (N16805, N16790, N12761, N2575, N11627);
or OR3 (N16806, N16805, N3778, N5623);
buf BUF1 (N16807, N16803);
nand NAND3 (N16808, N16806, N14101, N13930);
xor XOR2 (N16809, N16787, N10511);
buf BUF1 (N16810, N16789);
or OR3 (N16811, N16808, N10261, N6922);
xor XOR2 (N16812, N16807, N9608);
not NOT1 (N16813, N16804);
or OR3 (N16814, N16812, N9035, N8777);
nor NOR4 (N16815, N16811, N2030, N5678, N9654);
or OR3 (N16816, N16813, N11659, N10931);
buf BUF1 (N16817, N16814);
or OR2 (N16818, N16785, N11320);
nor NOR2 (N16819, N16798, N15921);
nor NOR2 (N16820, N16800, N12289);
nand NAND4 (N16821, N16820, N5615, N7163, N10786);
nand NAND3 (N16822, N16819, N2658, N15659);
nor NOR4 (N16823, N16799, N9321, N3298, N10000);
nor NOR2 (N16824, N16821, N16227);
buf BUF1 (N16825, N16809);
buf BUF1 (N16826, N16816);
nand NAND3 (N16827, N16825, N81, N1316);
nand NAND2 (N16828, N16822, N1444);
nand NAND4 (N16829, N16827, N16781, N11053, N246);
and AND4 (N16830, N16826, N115, N12221, N11233);
nand NAND4 (N16831, N16818, N10023, N7484, N6762);
or OR4 (N16832, N16802, N10278, N8024, N8576);
and AND4 (N16833, N16828, N10113, N5743, N5074);
and AND3 (N16834, N16831, N2723, N16058);
or OR4 (N16835, N16810, N9916, N8361, N16176);
not NOT1 (N16836, N16833);
nor NOR4 (N16837, N16834, N11586, N8807, N4710);
nor NOR2 (N16838, N16823, N10277);
or OR3 (N16839, N16830, N1075, N4028);
not NOT1 (N16840, N16835);
and AND4 (N16841, N16824, N8070, N8154, N14283);
xor XOR2 (N16842, N16832, N16570);
nand NAND2 (N16843, N16842, N15928);
xor XOR2 (N16844, N16840, N13137);
not NOT1 (N16845, N16839);
nor NOR3 (N16846, N16837, N5708, N1906);
or OR2 (N16847, N16844, N12325);
and AND4 (N16848, N16815, N9869, N8567, N12499);
buf BUF1 (N16849, N16841);
nor NOR2 (N16850, N16848, N9819);
and AND3 (N16851, N16838, N15464, N1712);
buf BUF1 (N16852, N16836);
nor NOR3 (N16853, N16843, N9891, N16841);
and AND2 (N16854, N16845, N8999);
xor XOR2 (N16855, N16846, N11943);
not NOT1 (N16856, N16817);
and AND4 (N16857, N16852, N3984, N7005, N5092);
buf BUF1 (N16858, N16854);
nand NAND3 (N16859, N16849, N4691, N1155);
or OR2 (N16860, N16847, N7182);
or OR3 (N16861, N16857, N5590, N9719);
xor XOR2 (N16862, N16861, N3768);
and AND2 (N16863, N16851, N8646);
buf BUF1 (N16864, N16853);
nand NAND4 (N16865, N16829, N14600, N7637, N16666);
or OR3 (N16866, N16858, N230, N13558);
buf BUF1 (N16867, N16850);
nor NOR2 (N16868, N16866, N7969);
nand NAND3 (N16869, N16868, N14046, N14475);
nor NOR2 (N16870, N16862, N14084);
nand NAND3 (N16871, N16860, N422, N4687);
nand NAND4 (N16872, N16870, N8577, N11417, N534);
nor NOR3 (N16873, N16863, N12411, N9838);
nor NOR3 (N16874, N16873, N8980, N2829);
buf BUF1 (N16875, N16872);
xor XOR2 (N16876, N16869, N4649);
or OR3 (N16877, N16856, N7540, N15751);
and AND4 (N16878, N16859, N13123, N2165, N12532);
and AND2 (N16879, N16871, N11714);
xor XOR2 (N16880, N16874, N6317);
xor XOR2 (N16881, N16877, N15938);
or OR3 (N16882, N16876, N15825, N9820);
nor NOR3 (N16883, N16865, N13420, N4091);
not NOT1 (N16884, N16875);
buf BUF1 (N16885, N16881);
nor NOR3 (N16886, N16879, N700, N3268);
nand NAND4 (N16887, N16882, N9371, N1114, N12385);
not NOT1 (N16888, N16883);
buf BUF1 (N16889, N16887);
nor NOR3 (N16890, N16864, N12484, N12555);
nand NAND4 (N16891, N16885, N7311, N10564, N15632);
buf BUF1 (N16892, N16888);
or OR4 (N16893, N16886, N8535, N9725, N10454);
or OR4 (N16894, N16893, N5305, N7566, N13063);
xor XOR2 (N16895, N16891, N5857);
or OR2 (N16896, N16889, N12967);
or OR2 (N16897, N16890, N10378);
buf BUF1 (N16898, N16894);
xor XOR2 (N16899, N16892, N9956);
buf BUF1 (N16900, N16895);
nand NAND2 (N16901, N16897, N12897);
not NOT1 (N16902, N16855);
nand NAND4 (N16903, N16902, N11415, N4662, N10585);
buf BUF1 (N16904, N16901);
nor NOR2 (N16905, N16880, N7174);
nor NOR4 (N16906, N16904, N321, N13453, N4213);
or OR2 (N16907, N16884, N5810);
xor XOR2 (N16908, N16907, N15285);
buf BUF1 (N16909, N16905);
xor XOR2 (N16910, N16908, N10165);
nor NOR3 (N16911, N16878, N6175, N8108);
buf BUF1 (N16912, N16867);
xor XOR2 (N16913, N16912, N13764);
xor XOR2 (N16914, N16909, N12096);
nor NOR3 (N16915, N16914, N4223, N6791);
buf BUF1 (N16916, N16913);
nor NOR3 (N16917, N16910, N16866, N12073);
not NOT1 (N16918, N16900);
not NOT1 (N16919, N16915);
nor NOR3 (N16920, N16896, N9291, N16291);
and AND2 (N16921, N16898, N15685);
xor XOR2 (N16922, N16903, N14476);
or OR4 (N16923, N16911, N7530, N8239, N1017);
nand NAND3 (N16924, N16919, N13398, N6132);
nor NOR4 (N16925, N16916, N12546, N16209, N16039);
nand NAND3 (N16926, N16922, N12892, N6107);
buf BUF1 (N16927, N16925);
nand NAND3 (N16928, N16920, N13108, N15030);
or OR2 (N16929, N16906, N6779);
or OR4 (N16930, N16923, N8505, N14309, N15943);
nand NAND4 (N16931, N16927, N1165, N14681, N15817);
and AND3 (N16932, N16917, N221, N11409);
buf BUF1 (N16933, N16928);
and AND2 (N16934, N16918, N3577);
xor XOR2 (N16935, N16931, N9107);
buf BUF1 (N16936, N16899);
not NOT1 (N16937, N16934);
buf BUF1 (N16938, N16929);
or OR4 (N16939, N16924, N15333, N3373, N5793);
buf BUF1 (N16940, N16921);
xor XOR2 (N16941, N16937, N6668);
nor NOR4 (N16942, N16936, N9836, N5455, N10939);
buf BUF1 (N16943, N16933);
or OR3 (N16944, N16942, N9800, N1837);
and AND2 (N16945, N16930, N15640);
or OR2 (N16946, N16926, N3865);
not NOT1 (N16947, N16939);
not NOT1 (N16948, N16938);
and AND3 (N16949, N16948, N12860, N11987);
not NOT1 (N16950, N16945);
buf BUF1 (N16951, N16944);
xor XOR2 (N16952, N16940, N6281);
nand NAND2 (N16953, N16951, N176);
or OR2 (N16954, N16949, N7739);
buf BUF1 (N16955, N16954);
nand NAND4 (N16956, N16946, N16477, N13292, N11048);
or OR3 (N16957, N16941, N10467, N15955);
nand NAND2 (N16958, N16935, N9078);
or OR2 (N16959, N16956, N13057);
and AND2 (N16960, N16957, N7511);
or OR4 (N16961, N16955, N12569, N1054, N16111);
xor XOR2 (N16962, N16950, N8413);
and AND3 (N16963, N16953, N237, N9037);
buf BUF1 (N16964, N16952);
not NOT1 (N16965, N16962);
not NOT1 (N16966, N16958);
not NOT1 (N16967, N16947);
or OR2 (N16968, N16963, N11480);
or OR2 (N16969, N16932, N5623);
buf BUF1 (N16970, N16964);
buf BUF1 (N16971, N16959);
and AND2 (N16972, N16971, N606);
and AND2 (N16973, N16967, N1869);
nand NAND4 (N16974, N16961, N5474, N6521, N12898);
xor XOR2 (N16975, N16960, N15632);
xor XOR2 (N16976, N16972, N16642);
xor XOR2 (N16977, N16965, N2903);
xor XOR2 (N16978, N16966, N13658);
buf BUF1 (N16979, N16978);
xor XOR2 (N16980, N16970, N1438);
not NOT1 (N16981, N16979);
buf BUF1 (N16982, N16977);
xor XOR2 (N16983, N16980, N5143);
buf BUF1 (N16984, N16983);
nand NAND3 (N16985, N16975, N9601, N15264);
or OR2 (N16986, N16973, N5191);
or OR4 (N16987, N16974, N6962, N171, N14226);
or OR2 (N16988, N16976, N13673);
xor XOR2 (N16989, N16985, N7912);
or OR2 (N16990, N16987, N14250);
not NOT1 (N16991, N16968);
and AND3 (N16992, N16991, N8998, N5000);
not NOT1 (N16993, N16981);
nor NOR4 (N16994, N16969, N5955, N7143, N988);
or OR4 (N16995, N16988, N4572, N8598, N14737);
and AND3 (N16996, N16995, N15122, N5877);
and AND4 (N16997, N16986, N16457, N4662, N14880);
and AND2 (N16998, N16982, N4580);
buf BUF1 (N16999, N16989);
nand NAND4 (N17000, N16984, N2635, N2076, N11171);
nand NAND4 (N17001, N16992, N12238, N12812, N16413);
xor XOR2 (N17002, N16996, N1217);
buf BUF1 (N17003, N16990);
not NOT1 (N17004, N16998);
buf BUF1 (N17005, N16943);
and AND3 (N17006, N17005, N9605, N11278);
nand NAND4 (N17007, N17003, N9513, N9467, N7816);
and AND4 (N17008, N16994, N13941, N6387, N14267);
xor XOR2 (N17009, N16993, N276);
nor NOR4 (N17010, N17006, N503, N15888, N13807);
and AND4 (N17011, N17000, N412, N9837, N10690);
buf BUF1 (N17012, N17008);
nor NOR4 (N17013, N16997, N16442, N2844, N15444);
not NOT1 (N17014, N17002);
not NOT1 (N17015, N16999);
nor NOR2 (N17016, N17012, N9087);
buf BUF1 (N17017, N17010);
nand NAND2 (N17018, N17009, N16341);
nor NOR4 (N17019, N17011, N12949, N11431, N8043);
not NOT1 (N17020, N17014);
buf BUF1 (N17021, N17019);
or OR2 (N17022, N17020, N546);
nand NAND3 (N17023, N17004, N169, N16702);
or OR4 (N17024, N17018, N7889, N13422, N12908);
buf BUF1 (N17025, N17007);
and AND4 (N17026, N17024, N1278, N13026, N3355);
and AND3 (N17027, N17013, N8848, N2381);
and AND4 (N17028, N17022, N7080, N14668, N15328);
buf BUF1 (N17029, N17021);
buf BUF1 (N17030, N17029);
and AND3 (N17031, N17030, N2199, N14650);
nand NAND4 (N17032, N17023, N4745, N4898, N4504);
or OR4 (N17033, N17016, N4549, N12032, N10556);
nand NAND4 (N17034, N17017, N6890, N8314, N5263);
or OR3 (N17035, N17032, N352, N8356);
xor XOR2 (N17036, N17028, N4768);
xor XOR2 (N17037, N17027, N10855);
nand NAND4 (N17038, N17034, N8362, N4824, N3822);
not NOT1 (N17039, N17026);
buf BUF1 (N17040, N17039);
not NOT1 (N17041, N17001);
or OR4 (N17042, N17035, N6482, N6980, N13931);
nor NOR3 (N17043, N17038, N13503, N14938);
not NOT1 (N17044, N17037);
not NOT1 (N17045, N17025);
or OR2 (N17046, N17036, N4406);
not NOT1 (N17047, N17044);
nand NAND4 (N17048, N17046, N9490, N13569, N5110);
buf BUF1 (N17049, N17042);
not NOT1 (N17050, N17049);
or OR4 (N17051, N17048, N2815, N16717, N15833);
not NOT1 (N17052, N17033);
xor XOR2 (N17053, N17050, N11432);
or OR3 (N17054, N17045, N9811, N11035);
buf BUF1 (N17055, N17054);
xor XOR2 (N17056, N17055, N4481);
nand NAND2 (N17057, N17052, N8285);
or OR4 (N17058, N17056, N12296, N6904, N8737);
nand NAND2 (N17059, N17058, N11771);
and AND4 (N17060, N17059, N14811, N1725, N11209);
buf BUF1 (N17061, N17043);
nor NOR3 (N17062, N17031, N2349, N12325);
and AND3 (N17063, N17047, N4890, N16967);
nor NOR2 (N17064, N17062, N13816);
and AND2 (N17065, N17015, N5428);
and AND4 (N17066, N17060, N7000, N933, N14406);
xor XOR2 (N17067, N17040, N5861);
and AND2 (N17068, N17063, N7348);
nand NAND4 (N17069, N17041, N163, N15641, N4966);
xor XOR2 (N17070, N17068, N15400);
buf BUF1 (N17071, N17065);
nor NOR4 (N17072, N17070, N7052, N5069, N1329);
nand NAND3 (N17073, N17067, N825, N4613);
not NOT1 (N17074, N17073);
xor XOR2 (N17075, N17071, N8412);
and AND2 (N17076, N17057, N14989);
or OR2 (N17077, N17064, N543);
and AND3 (N17078, N17075, N4354, N3124);
not NOT1 (N17079, N17078);
xor XOR2 (N17080, N17077, N7348);
buf BUF1 (N17081, N17051);
xor XOR2 (N17082, N17072, N3445);
buf BUF1 (N17083, N17079);
buf BUF1 (N17084, N17069);
nor NOR4 (N17085, N17066, N16835, N14468, N4502);
and AND2 (N17086, N17053, N7715);
or OR2 (N17087, N17085, N1999);
and AND2 (N17088, N17081, N7210);
or OR2 (N17089, N17086, N8187);
nand NAND3 (N17090, N17087, N8028, N8167);
not NOT1 (N17091, N17088);
buf BUF1 (N17092, N17074);
nand NAND2 (N17093, N17092, N4567);
or OR4 (N17094, N17083, N13784, N6973, N7336);
or OR4 (N17095, N17090, N8026, N12430, N7452);
and AND4 (N17096, N17091, N1325, N12074, N166);
or OR2 (N17097, N17082, N8175);
nor NOR3 (N17098, N17097, N3856, N10729);
nor NOR2 (N17099, N17061, N16400);
not NOT1 (N17100, N17080);
nor NOR3 (N17101, N17093, N7920, N16327);
or OR2 (N17102, N17076, N3402);
or OR2 (N17103, N17101, N8402);
nand NAND4 (N17104, N17094, N15798, N10968, N8726);
and AND3 (N17105, N17103, N9976, N123);
or OR4 (N17106, N17104, N7536, N17024, N5519);
and AND2 (N17107, N17102, N6830);
not NOT1 (N17108, N17100);
xor XOR2 (N17109, N17107, N2267);
buf BUF1 (N17110, N17109);
xor XOR2 (N17111, N17108, N2844);
buf BUF1 (N17112, N17095);
nand NAND3 (N17113, N17084, N3232, N7815);
or OR2 (N17114, N17111, N11889);
not NOT1 (N17115, N17089);
xor XOR2 (N17116, N17115, N6119);
nor NOR2 (N17117, N17096, N1350);
not NOT1 (N17118, N17114);
nand NAND4 (N17119, N17117, N3245, N7906, N16488);
nand NAND2 (N17120, N17116, N2095);
or OR3 (N17121, N17106, N5825, N2789);
or OR2 (N17122, N17105, N5029);
not NOT1 (N17123, N17110);
and AND4 (N17124, N17123, N479, N1637, N8253);
xor XOR2 (N17125, N17098, N6808);
or OR3 (N17126, N17121, N4473, N15899);
xor XOR2 (N17127, N17126, N6698);
not NOT1 (N17128, N17112);
nor NOR4 (N17129, N17120, N15509, N13041, N3408);
and AND4 (N17130, N17124, N6982, N8466, N9571);
not NOT1 (N17131, N17128);
and AND4 (N17132, N17118, N373, N1188, N132);
not NOT1 (N17133, N17129);
not NOT1 (N17134, N17122);
xor XOR2 (N17135, N17127, N8189);
not NOT1 (N17136, N17131);
not NOT1 (N17137, N17130);
nand NAND4 (N17138, N17132, N14959, N16359, N6837);
or OR4 (N17139, N17119, N8709, N5373, N14846);
and AND4 (N17140, N17125, N16157, N8504, N8092);
and AND2 (N17141, N17113, N6610);
nand NAND2 (N17142, N17135, N7769);
xor XOR2 (N17143, N17141, N4246);
nand NAND3 (N17144, N17142, N13397, N9199);
and AND2 (N17145, N17138, N4523);
and AND4 (N17146, N17143, N12870, N8749, N7771);
nand NAND2 (N17147, N17145, N8323);
nor NOR4 (N17148, N17133, N7876, N9249, N12859);
xor XOR2 (N17149, N17136, N5038);
buf BUF1 (N17150, N17144);
and AND3 (N17151, N17137, N5121, N2256);
xor XOR2 (N17152, N17099, N8426);
or OR3 (N17153, N17147, N14695, N7115);
not NOT1 (N17154, N17149);
buf BUF1 (N17155, N17154);
or OR3 (N17156, N17139, N16966, N11600);
not NOT1 (N17157, N17153);
not NOT1 (N17158, N17140);
and AND2 (N17159, N17150, N803);
or OR3 (N17160, N17157, N10529, N3137);
or OR3 (N17161, N17158, N3782, N1880);
or OR4 (N17162, N17161, N9666, N12808, N2460);
not NOT1 (N17163, N17160);
xor XOR2 (N17164, N17151, N14167);
or OR2 (N17165, N17162, N13550);
buf BUF1 (N17166, N17156);
nor NOR2 (N17167, N17165, N14448);
or OR2 (N17168, N17155, N10102);
nand NAND2 (N17169, N17164, N8774);
nor NOR2 (N17170, N17169, N13231);
and AND4 (N17171, N17168, N8117, N4112, N11580);
xor XOR2 (N17172, N17148, N9209);
nand NAND3 (N17173, N17134, N4867, N10763);
xor XOR2 (N17174, N17172, N9660);
or OR2 (N17175, N17173, N2148);
nor NOR2 (N17176, N17170, N13305);
not NOT1 (N17177, N17176);
xor XOR2 (N17178, N17152, N5855);
nand NAND4 (N17179, N17167, N4350, N11478, N14275);
or OR2 (N17180, N17179, N14513);
or OR4 (N17181, N17166, N16894, N9167, N12226);
and AND2 (N17182, N17163, N839);
nor NOR2 (N17183, N17146, N9498);
nand NAND4 (N17184, N17171, N13715, N8230, N3548);
nand NAND2 (N17185, N17184, N5565);
not NOT1 (N17186, N17181);
not NOT1 (N17187, N17186);
or OR2 (N17188, N17180, N14158);
and AND4 (N17189, N17177, N15875, N9912, N10576);
buf BUF1 (N17190, N17182);
nand NAND4 (N17191, N17183, N4597, N3438, N13723);
not NOT1 (N17192, N17191);
nand NAND3 (N17193, N17187, N11116, N8327);
or OR2 (N17194, N17159, N13969);
and AND3 (N17195, N17189, N14242, N12654);
nand NAND2 (N17196, N17175, N6053);
xor XOR2 (N17197, N17188, N2413);
and AND2 (N17198, N17193, N240);
nand NAND2 (N17199, N17192, N10798);
nand NAND4 (N17200, N17199, N14699, N4977, N14364);
nor NOR3 (N17201, N17174, N14951, N13601);
not NOT1 (N17202, N17194);
buf BUF1 (N17203, N17200);
buf BUF1 (N17204, N17202);
nand NAND2 (N17205, N17190, N16080);
nand NAND3 (N17206, N17196, N14368, N3953);
and AND4 (N17207, N17206, N1936, N4316, N3614);
nor NOR2 (N17208, N17195, N9962);
not NOT1 (N17209, N17201);
or OR2 (N17210, N17198, N3794);
or OR2 (N17211, N17210, N12862);
xor XOR2 (N17212, N17203, N16071);
nor NOR4 (N17213, N17211, N15335, N15146, N9820);
nor NOR2 (N17214, N17197, N4568);
nand NAND3 (N17215, N17208, N1470, N2624);
not NOT1 (N17216, N17209);
nor NOR4 (N17217, N17204, N446, N9466, N3407);
xor XOR2 (N17218, N17207, N11970);
nor NOR4 (N17219, N17213, N3449, N7658, N12789);
nor NOR4 (N17220, N17217, N7022, N6310, N7493);
nor NOR2 (N17221, N17185, N5667);
not NOT1 (N17222, N17205);
or OR4 (N17223, N17214, N3163, N13211, N7472);
buf BUF1 (N17224, N17223);
and AND2 (N17225, N17215, N13477);
nor NOR3 (N17226, N17222, N16332, N11986);
nor NOR3 (N17227, N17224, N7065, N11831);
and AND3 (N17228, N17226, N11265, N14544);
and AND2 (N17229, N17218, N14144);
buf BUF1 (N17230, N17219);
and AND3 (N17231, N17221, N6, N11529);
or OR3 (N17232, N17212, N16792, N7063);
xor XOR2 (N17233, N17231, N4789);
not NOT1 (N17234, N17216);
nand NAND3 (N17235, N17233, N5496, N9851);
and AND3 (N17236, N17227, N2081, N16431);
buf BUF1 (N17237, N17234);
buf BUF1 (N17238, N17237);
buf BUF1 (N17239, N17178);
not NOT1 (N17240, N17228);
or OR3 (N17241, N17230, N10801, N6529);
buf BUF1 (N17242, N17229);
nand NAND4 (N17243, N17232, N746, N11849, N15953);
or OR3 (N17244, N17236, N10937, N10556);
nor NOR2 (N17245, N17241, N10778);
buf BUF1 (N17246, N17225);
nor NOR3 (N17247, N17242, N2027, N16938);
nor NOR2 (N17248, N17235, N3667);
buf BUF1 (N17249, N17244);
or OR4 (N17250, N17220, N17076, N8745, N8765);
buf BUF1 (N17251, N17246);
buf BUF1 (N17252, N17238);
and AND2 (N17253, N17243, N967);
nand NAND2 (N17254, N17240, N1251);
and AND3 (N17255, N17248, N11599, N13467);
buf BUF1 (N17256, N17253);
nor NOR2 (N17257, N17249, N16743);
buf BUF1 (N17258, N17252);
and AND3 (N17259, N17256, N826, N8847);
and AND2 (N17260, N17255, N13602);
nor NOR3 (N17261, N17258, N5055, N7541);
buf BUF1 (N17262, N17245);
buf BUF1 (N17263, N17260);
and AND3 (N17264, N17257, N2553, N6416);
nand NAND3 (N17265, N17259, N6952, N16840);
or OR2 (N17266, N17247, N15894);
or OR4 (N17267, N17265, N2157, N6918, N2888);
xor XOR2 (N17268, N17261, N8639);
nand NAND2 (N17269, N17250, N15819);
not NOT1 (N17270, N17268);
nor NOR4 (N17271, N17264, N16021, N11406, N1433);
buf BUF1 (N17272, N17239);
buf BUF1 (N17273, N17267);
nand NAND4 (N17274, N17266, N5289, N6841, N1166);
xor XOR2 (N17275, N17263, N10827);
not NOT1 (N17276, N17272);
nand NAND3 (N17277, N17275, N13208, N6370);
or OR3 (N17278, N17273, N4260, N3185);
xor XOR2 (N17279, N17262, N10177);
xor XOR2 (N17280, N17276, N11427);
buf BUF1 (N17281, N17279);
buf BUF1 (N17282, N17271);
buf BUF1 (N17283, N17274);
not NOT1 (N17284, N17269);
not NOT1 (N17285, N17284);
buf BUF1 (N17286, N17285);
or OR4 (N17287, N17270, N6361, N8281, N10109);
not NOT1 (N17288, N17283);
xor XOR2 (N17289, N17277, N16596);
or OR4 (N17290, N17281, N654, N4442, N10225);
nand NAND2 (N17291, N17288, N13479);
buf BUF1 (N17292, N17286);
or OR3 (N17293, N17280, N13114, N16261);
xor XOR2 (N17294, N17278, N1920);
not NOT1 (N17295, N17291);
or OR3 (N17296, N17294, N4941, N1649);
nand NAND3 (N17297, N17296, N4359, N5454);
buf BUF1 (N17298, N17290);
or OR2 (N17299, N17282, N8802);
xor XOR2 (N17300, N17297, N5967);
and AND4 (N17301, N17289, N1797, N2507, N11939);
buf BUF1 (N17302, N17292);
buf BUF1 (N17303, N17302);
xor XOR2 (N17304, N17298, N14914);
and AND3 (N17305, N17293, N3440, N4617);
not NOT1 (N17306, N17300);
xor XOR2 (N17307, N17305, N13938);
or OR2 (N17308, N17287, N3379);
xor XOR2 (N17309, N17251, N7657);
not NOT1 (N17310, N17295);
not NOT1 (N17311, N17308);
buf BUF1 (N17312, N17301);
nor NOR2 (N17313, N17307, N2934);
not NOT1 (N17314, N17311);
buf BUF1 (N17315, N17306);
or OR2 (N17316, N17299, N16282);
buf BUF1 (N17317, N17310);
not NOT1 (N17318, N17304);
or OR2 (N17319, N17314, N10351);
xor XOR2 (N17320, N17303, N7412);
not NOT1 (N17321, N17319);
nor NOR3 (N17322, N17313, N1068, N17252);
or OR4 (N17323, N17315, N10914, N597, N17007);
nor NOR2 (N17324, N17316, N9482);
buf BUF1 (N17325, N17324);
buf BUF1 (N17326, N17323);
or OR3 (N17327, N17317, N11294, N16656);
not NOT1 (N17328, N17325);
not NOT1 (N17329, N17327);
buf BUF1 (N17330, N17329);
xor XOR2 (N17331, N17318, N10978);
nor NOR3 (N17332, N17328, N15160, N16366);
or OR4 (N17333, N17331, N13170, N4534, N5908);
nor NOR4 (N17334, N17312, N9524, N6932, N12935);
or OR2 (N17335, N17332, N13484);
and AND3 (N17336, N17321, N1360, N3791);
or OR2 (N17337, N17254, N4358);
buf BUF1 (N17338, N17333);
not NOT1 (N17339, N17320);
nand NAND3 (N17340, N17337, N11170, N14428);
buf BUF1 (N17341, N17338);
or OR4 (N17342, N17326, N14601, N11652, N4031);
nand NAND2 (N17343, N17336, N15997);
nand NAND4 (N17344, N17342, N2551, N10824, N12555);
and AND2 (N17345, N17341, N15620);
xor XOR2 (N17346, N17334, N17138);
xor XOR2 (N17347, N17343, N7461);
xor XOR2 (N17348, N17347, N445);
or OR4 (N17349, N17322, N10813, N12400, N1126);
xor XOR2 (N17350, N17340, N15359);
nand NAND3 (N17351, N17330, N14830, N9635);
buf BUF1 (N17352, N17335);
xor XOR2 (N17353, N17344, N13627);
and AND2 (N17354, N17352, N951);
and AND4 (N17355, N17353, N16422, N6292, N5830);
nand NAND3 (N17356, N17351, N9213, N6417);
nor NOR3 (N17357, N17356, N10371, N13335);
not NOT1 (N17358, N17349);
nand NAND4 (N17359, N17339, N3544, N9652, N7856);
and AND2 (N17360, N17350, N8867);
and AND3 (N17361, N17345, N13371, N11338);
not NOT1 (N17362, N17346);
and AND4 (N17363, N17355, N9224, N943, N12020);
nand NAND2 (N17364, N17357, N713);
buf BUF1 (N17365, N17359);
nor NOR3 (N17366, N17309, N9051, N3953);
nor NOR2 (N17367, N17360, N14097);
nor NOR3 (N17368, N17348, N1183, N2710);
or OR4 (N17369, N17358, N9862, N5801, N6197);
and AND4 (N17370, N17369, N14813, N10028, N11644);
xor XOR2 (N17371, N17370, N6563);
not NOT1 (N17372, N17362);
not NOT1 (N17373, N17371);
nand NAND3 (N17374, N17364, N10330, N2335);
and AND3 (N17375, N17367, N269, N10766);
and AND2 (N17376, N17372, N3683);
xor XOR2 (N17377, N17373, N3492);
nand NAND4 (N17378, N17361, N2270, N16122, N4012);
or OR2 (N17379, N17376, N1581);
nand NAND2 (N17380, N17368, N12765);
and AND2 (N17381, N17365, N2310);
or OR2 (N17382, N17378, N16984);
nand NAND3 (N17383, N17382, N14752, N6466);
and AND4 (N17384, N17375, N17341, N5935, N6059);
buf BUF1 (N17385, N17363);
and AND4 (N17386, N17381, N9725, N11605, N8773);
not NOT1 (N17387, N17354);
or OR3 (N17388, N17383, N16534, N859);
nor NOR4 (N17389, N17385, N10865, N8664, N2671);
nor NOR4 (N17390, N17386, N16842, N7184, N11344);
and AND3 (N17391, N17387, N6459, N15046);
buf BUF1 (N17392, N17388);
or OR4 (N17393, N17391, N14088, N8925, N1621);
or OR2 (N17394, N17393, N11981);
nor NOR2 (N17395, N17380, N12961);
and AND2 (N17396, N17392, N15885);
and AND3 (N17397, N17390, N12598, N8560);
not NOT1 (N17398, N17374);
not NOT1 (N17399, N17396);
nor NOR3 (N17400, N17366, N5891, N2640);
and AND4 (N17401, N17395, N12783, N13211, N14224);
nor NOR4 (N17402, N17401, N2737, N6113, N5785);
or OR4 (N17403, N17400, N3144, N11678, N7690);
buf BUF1 (N17404, N17379);
nor NOR4 (N17405, N17402, N474, N11826, N4485);
nor NOR2 (N17406, N17399, N11630);
and AND2 (N17407, N17389, N10531);
buf BUF1 (N17408, N17406);
buf BUF1 (N17409, N17398);
and AND4 (N17410, N17394, N2913, N3209, N8026);
nand NAND2 (N17411, N17410, N3749);
nor NOR3 (N17412, N17409, N6396, N15407);
and AND3 (N17413, N17404, N9061, N15713);
nor NOR4 (N17414, N17377, N10443, N13718, N3740);
and AND4 (N17415, N17384, N16439, N16216, N8179);
nor NOR4 (N17416, N17407, N9869, N15815, N7528);
xor XOR2 (N17417, N17408, N5630);
and AND3 (N17418, N17413, N9165, N10551);
not NOT1 (N17419, N17415);
nor NOR2 (N17420, N17416, N10224);
nand NAND2 (N17421, N17412, N1985);
and AND4 (N17422, N17411, N11412, N14790, N7382);
buf BUF1 (N17423, N17418);
nand NAND2 (N17424, N17397, N8356);
buf BUF1 (N17425, N17405);
xor XOR2 (N17426, N17414, N12563);
buf BUF1 (N17427, N17422);
not NOT1 (N17428, N17417);
xor XOR2 (N17429, N17419, N15711);
or OR4 (N17430, N17420, N14524, N2737, N11736);
or OR4 (N17431, N17426, N12259, N14780, N10435);
nand NAND3 (N17432, N17431, N1582, N10063);
and AND4 (N17433, N17425, N6578, N5158, N3360);
nor NOR3 (N17434, N17428, N15817, N13405);
or OR4 (N17435, N17421, N14217, N9254, N6173);
nand NAND3 (N17436, N17429, N366, N13845);
buf BUF1 (N17437, N17435);
nor NOR4 (N17438, N17403, N11376, N5780, N10229);
and AND3 (N17439, N17424, N11084, N3299);
and AND4 (N17440, N17430, N10047, N15763, N9620);
nand NAND2 (N17441, N17439, N7430);
nor NOR2 (N17442, N17436, N1051);
and AND3 (N17443, N17438, N9293, N13231);
nand NAND3 (N17444, N17441, N12596, N12047);
nand NAND3 (N17445, N17443, N4078, N7743);
or OR3 (N17446, N17445, N8417, N13995);
nand NAND2 (N17447, N17446, N15207);
nand NAND2 (N17448, N17440, N14267);
and AND3 (N17449, N17444, N6636, N10980);
nand NAND2 (N17450, N17433, N707);
buf BUF1 (N17451, N17432);
not NOT1 (N17452, N17437);
and AND3 (N17453, N17423, N9433, N2642);
and AND3 (N17454, N17452, N16989, N4114);
nand NAND4 (N17455, N17434, N2729, N13515, N1199);
xor XOR2 (N17456, N17447, N12154);
buf BUF1 (N17457, N17450);
and AND4 (N17458, N17455, N12255, N8238, N12576);
buf BUF1 (N17459, N17449);
nand NAND2 (N17460, N17453, N3753);
buf BUF1 (N17461, N17427);
and AND2 (N17462, N17459, N17123);
nand NAND4 (N17463, N17448, N4308, N2360, N4967);
or OR2 (N17464, N17462, N390);
not NOT1 (N17465, N17463);
or OR3 (N17466, N17456, N2477, N2301);
or OR3 (N17467, N17461, N3528, N16119);
not NOT1 (N17468, N17457);
or OR4 (N17469, N17465, N12156, N10802, N415);
xor XOR2 (N17470, N17468, N2942);
buf BUF1 (N17471, N17458);
or OR3 (N17472, N17469, N15911, N1310);
nand NAND3 (N17473, N17460, N8677, N3194);
or OR4 (N17474, N17466, N14722, N119, N14302);
or OR2 (N17475, N17473, N4805);
or OR4 (N17476, N17442, N157, N2623, N9048);
nor NOR4 (N17477, N17475, N6955, N11866, N12465);
nand NAND3 (N17478, N17454, N8969, N4939);
not NOT1 (N17479, N17467);
nor NOR3 (N17480, N17477, N8096, N6163);
and AND3 (N17481, N17479, N481, N1959);
or OR3 (N17482, N17464, N956, N5425);
nand NAND2 (N17483, N17481, N9411);
xor XOR2 (N17484, N17474, N2353);
nand NAND4 (N17485, N17471, N4901, N3016, N368);
nand NAND2 (N17486, N17478, N6048);
not NOT1 (N17487, N17472);
not NOT1 (N17488, N17482);
not NOT1 (N17489, N17486);
buf BUF1 (N17490, N17451);
xor XOR2 (N17491, N17485, N7604);
buf BUF1 (N17492, N17483);
nor NOR4 (N17493, N17484, N11745, N17092, N12998);
and AND2 (N17494, N17489, N4602);
not NOT1 (N17495, N17470);
not NOT1 (N17496, N17488);
not NOT1 (N17497, N17491);
or OR3 (N17498, N17496, N8374, N13290);
not NOT1 (N17499, N17495);
not NOT1 (N17500, N17493);
xor XOR2 (N17501, N17497, N15942);
or OR4 (N17502, N17487, N4112, N1188, N493);
not NOT1 (N17503, N17490);
not NOT1 (N17504, N17498);
nand NAND4 (N17505, N17504, N323, N6242, N7206);
and AND2 (N17506, N17476, N5389);
xor XOR2 (N17507, N17505, N14576);
xor XOR2 (N17508, N17492, N13152);
nor NOR2 (N17509, N17494, N2564);
not NOT1 (N17510, N17503);
or OR3 (N17511, N17501, N7970, N15657);
nor NOR3 (N17512, N17502, N14910, N6923);
nand NAND3 (N17513, N17507, N8472, N14447);
not NOT1 (N17514, N17500);
buf BUF1 (N17515, N17510);
and AND4 (N17516, N17508, N9462, N12782, N16321);
nand NAND2 (N17517, N17512, N6446);
xor XOR2 (N17518, N17511, N15254);
and AND3 (N17519, N17518, N9389, N12736);
nand NAND2 (N17520, N17513, N12894);
and AND3 (N17521, N17515, N6663, N699);
buf BUF1 (N17522, N17519);
buf BUF1 (N17523, N17516);
nand NAND3 (N17524, N17522, N2617, N7492);
xor XOR2 (N17525, N17517, N8259);
not NOT1 (N17526, N17509);
nand NAND2 (N17527, N17524, N3916);
not NOT1 (N17528, N17514);
not NOT1 (N17529, N17523);
not NOT1 (N17530, N17520);
or OR2 (N17531, N17521, N6018);
xor XOR2 (N17532, N17499, N10833);
not NOT1 (N17533, N17528);
or OR2 (N17534, N17480, N5610);
and AND3 (N17535, N17526, N16356, N9634);
nand NAND4 (N17536, N17525, N8083, N7100, N8677);
or OR3 (N17537, N17531, N16125, N14750);
not NOT1 (N17538, N17533);
xor XOR2 (N17539, N17532, N2972);
and AND3 (N17540, N17506, N4298, N9828);
and AND4 (N17541, N17530, N7219, N1304, N15901);
buf BUF1 (N17542, N17534);
and AND4 (N17543, N17536, N5594, N7839, N2070);
xor XOR2 (N17544, N17543, N14588);
xor XOR2 (N17545, N17540, N12398);
and AND3 (N17546, N17542, N4057, N5079);
or OR3 (N17547, N17527, N13952, N5988);
xor XOR2 (N17548, N17535, N1273);
xor XOR2 (N17549, N17546, N7240);
and AND2 (N17550, N17544, N13073);
nand NAND4 (N17551, N17550, N7457, N1342, N11267);
and AND3 (N17552, N17538, N8173, N7602);
or OR3 (N17553, N17545, N8909, N3661);
not NOT1 (N17554, N17553);
or OR2 (N17555, N17554, N14658);
nor NOR4 (N17556, N17552, N7329, N10212, N14110);
not NOT1 (N17557, N17539);
not NOT1 (N17558, N17551);
xor XOR2 (N17559, N17541, N10503);
and AND3 (N17560, N17557, N3232, N15531);
and AND4 (N17561, N17549, N493, N16667, N10447);
or OR4 (N17562, N17559, N14562, N16820, N14578);
buf BUF1 (N17563, N17555);
nor NOR2 (N17564, N17548, N1284);
xor XOR2 (N17565, N17562, N16599);
and AND4 (N17566, N17561, N9066, N14488, N6336);
or OR3 (N17567, N17529, N9488, N9502);
or OR3 (N17568, N17563, N17120, N1954);
nor NOR4 (N17569, N17566, N9814, N11382, N1484);
nor NOR4 (N17570, N17537, N6295, N5408, N13583);
or OR3 (N17571, N17568, N15859, N10894);
not NOT1 (N17572, N17558);
and AND4 (N17573, N17572, N7070, N13567, N12133);
buf BUF1 (N17574, N17547);
xor XOR2 (N17575, N17571, N17160);
not NOT1 (N17576, N17570);
buf BUF1 (N17577, N17569);
nand NAND2 (N17578, N17575, N1106);
xor XOR2 (N17579, N17576, N3610);
and AND4 (N17580, N17565, N13439, N15668, N184);
nor NOR2 (N17581, N17560, N2112);
nand NAND4 (N17582, N17556, N7973, N10488, N7918);
buf BUF1 (N17583, N17577);
nor NOR4 (N17584, N17573, N1909, N7697, N11708);
or OR4 (N17585, N17583, N17215, N12908, N10104);
buf BUF1 (N17586, N17564);
xor XOR2 (N17587, N17574, N17143);
xor XOR2 (N17588, N17567, N12209);
or OR2 (N17589, N17585, N9626);
not NOT1 (N17590, N17587);
nor NOR3 (N17591, N17582, N9227, N7062);
or OR2 (N17592, N17588, N12294);
buf BUF1 (N17593, N17590);
xor XOR2 (N17594, N17592, N5148);
nand NAND3 (N17595, N17580, N4548, N7004);
xor XOR2 (N17596, N17593, N6722);
not NOT1 (N17597, N17584);
buf BUF1 (N17598, N17589);
buf BUF1 (N17599, N17578);
nor NOR2 (N17600, N17581, N831);
buf BUF1 (N17601, N17591);
nor NOR4 (N17602, N17586, N11465, N13532, N10184);
buf BUF1 (N17603, N17598);
nand NAND2 (N17604, N17599, N4463);
and AND3 (N17605, N17600, N13472, N14956);
buf BUF1 (N17606, N17596);
buf BUF1 (N17607, N17595);
buf BUF1 (N17608, N17597);
and AND3 (N17609, N17606, N8973, N15651);
xor XOR2 (N17610, N17579, N8872);
or OR3 (N17611, N17607, N7330, N11483);
and AND3 (N17612, N17604, N11685, N11137);
buf BUF1 (N17613, N17602);
and AND2 (N17614, N17608, N9203);
nand NAND3 (N17615, N17594, N1370, N11615);
or OR2 (N17616, N17611, N14322);
and AND3 (N17617, N17613, N5897, N10533);
nor NOR4 (N17618, N17601, N13098, N12588, N2604);
and AND2 (N17619, N17603, N4069);
not NOT1 (N17620, N17616);
not NOT1 (N17621, N17620);
not NOT1 (N17622, N17614);
xor XOR2 (N17623, N17605, N12703);
nand NAND3 (N17624, N17618, N3952, N12785);
nor NOR4 (N17625, N17612, N9182, N14250, N88);
xor XOR2 (N17626, N17610, N1482);
xor XOR2 (N17627, N17624, N9967);
buf BUF1 (N17628, N17617);
or OR3 (N17629, N17619, N7237, N6417);
and AND3 (N17630, N17629, N15543, N2555);
xor XOR2 (N17631, N17615, N5976);
and AND3 (N17632, N17609, N2574, N9956);
not NOT1 (N17633, N17631);
buf BUF1 (N17634, N17621);
not NOT1 (N17635, N17627);
not NOT1 (N17636, N17633);
not NOT1 (N17637, N17628);
xor XOR2 (N17638, N17625, N2321);
xor XOR2 (N17639, N17638, N10499);
buf BUF1 (N17640, N17635);
not NOT1 (N17641, N17634);
buf BUF1 (N17642, N17637);
not NOT1 (N17643, N17622);
and AND2 (N17644, N17636, N2528);
xor XOR2 (N17645, N17623, N5009);
not NOT1 (N17646, N17640);
and AND3 (N17647, N17639, N11983, N14925);
not NOT1 (N17648, N17647);
buf BUF1 (N17649, N17626);
or OR3 (N17650, N17646, N3235, N3332);
not NOT1 (N17651, N17630);
nand NAND2 (N17652, N17650, N9267);
nand NAND3 (N17653, N17651, N10943, N703);
and AND4 (N17654, N17644, N7004, N3051, N10276);
or OR4 (N17655, N17653, N2316, N12764, N897);
xor XOR2 (N17656, N17654, N2496);
nand NAND2 (N17657, N17652, N9075);
or OR2 (N17658, N17641, N3764);
not NOT1 (N17659, N17655);
nor NOR3 (N17660, N17648, N796, N7657);
nand NAND2 (N17661, N17645, N10737);
xor XOR2 (N17662, N17642, N9110);
not NOT1 (N17663, N17657);
xor XOR2 (N17664, N17660, N9903);
buf BUF1 (N17665, N17664);
nor NOR3 (N17666, N17663, N4009, N14973);
or OR4 (N17667, N17662, N1294, N14368, N17251);
and AND2 (N17668, N17666, N8688);
nor NOR3 (N17669, N17632, N8150, N16426);
and AND4 (N17670, N17669, N6431, N8536, N7717);
nand NAND4 (N17671, N17656, N11277, N5466, N4818);
nand NAND4 (N17672, N17649, N17490, N11888, N10840);
buf BUF1 (N17673, N17671);
and AND2 (N17674, N17665, N14552);
and AND2 (N17675, N17674, N110);
nand NAND3 (N17676, N17675, N16925, N7276);
nand NAND2 (N17677, N17676, N13969);
or OR3 (N17678, N17673, N10701, N17495);
and AND4 (N17679, N17668, N16392, N10552, N11641);
nand NAND3 (N17680, N17672, N16923, N5944);
not NOT1 (N17681, N17658);
nand NAND4 (N17682, N17670, N6115, N2935, N1768);
or OR2 (N17683, N17667, N15890);
buf BUF1 (N17684, N17683);
xor XOR2 (N17685, N17677, N134);
or OR2 (N17686, N17679, N7563);
and AND2 (N17687, N17685, N12057);
or OR2 (N17688, N17681, N7288);
and AND4 (N17689, N17678, N8069, N3220, N8732);
buf BUF1 (N17690, N17682);
or OR4 (N17691, N17688, N3741, N7652, N9154);
nand NAND3 (N17692, N17690, N16314, N13505);
or OR3 (N17693, N17684, N1817, N15593);
nand NAND3 (N17694, N17686, N13032, N2084);
nor NOR2 (N17695, N17689, N325);
or OR2 (N17696, N17661, N15843);
nand NAND2 (N17697, N17687, N2970);
nand NAND3 (N17698, N17695, N17681, N13990);
nand NAND2 (N17699, N17659, N13654);
or OR2 (N17700, N17698, N12071);
nand NAND4 (N17701, N17692, N3563, N17272, N5513);
xor XOR2 (N17702, N17696, N507);
xor XOR2 (N17703, N17691, N707);
buf BUF1 (N17704, N17693);
and AND4 (N17705, N17697, N2128, N8523, N11091);
or OR4 (N17706, N17701, N4399, N731, N1885);
not NOT1 (N17707, N17643);
not NOT1 (N17708, N17699);
not NOT1 (N17709, N17680);
buf BUF1 (N17710, N17703);
and AND2 (N17711, N17707, N2871);
buf BUF1 (N17712, N17705);
xor XOR2 (N17713, N17706, N16873);
and AND4 (N17714, N17711, N10035, N16553, N12734);
buf BUF1 (N17715, N17704);
or OR3 (N17716, N17709, N12550, N720);
or OR2 (N17717, N17715, N713);
nor NOR2 (N17718, N17702, N8591);
nand NAND2 (N17719, N17710, N8190);
and AND2 (N17720, N17718, N11789);
nand NAND2 (N17721, N17700, N13509);
nor NOR4 (N17722, N17708, N16055, N6484, N15597);
xor XOR2 (N17723, N17713, N11931);
and AND2 (N17724, N17723, N1301);
xor XOR2 (N17725, N17724, N15625);
and AND2 (N17726, N17717, N3992);
and AND4 (N17727, N17719, N4322, N14332, N1843);
or OR2 (N17728, N17714, N16418);
nor NOR2 (N17729, N17712, N4774);
not NOT1 (N17730, N17720);
and AND4 (N17731, N17729, N7615, N1675, N2852);
not NOT1 (N17732, N17728);
nor NOR3 (N17733, N17722, N4682, N653);
not NOT1 (N17734, N17725);
buf BUF1 (N17735, N17694);
buf BUF1 (N17736, N17733);
and AND4 (N17737, N17721, N1070, N17723, N7313);
xor XOR2 (N17738, N17737, N14659);
or OR4 (N17739, N17734, N510, N6666, N8721);
buf BUF1 (N17740, N17732);
nor NOR3 (N17741, N17716, N14938, N11275);
xor XOR2 (N17742, N17736, N12714);
buf BUF1 (N17743, N17726);
and AND3 (N17744, N17730, N412, N10088);
buf BUF1 (N17745, N17727);
buf BUF1 (N17746, N17735);
nor NOR3 (N17747, N17741, N11950, N11897);
buf BUF1 (N17748, N17743);
nor NOR2 (N17749, N17731, N3441);
and AND2 (N17750, N17747, N15216);
and AND4 (N17751, N17746, N10065, N1768, N3495);
or OR2 (N17752, N17751, N2389);
buf BUF1 (N17753, N17738);
not NOT1 (N17754, N17740);
and AND3 (N17755, N17752, N11753, N11905);
or OR2 (N17756, N17748, N17385);
not NOT1 (N17757, N17753);
and AND4 (N17758, N17745, N3675, N13446, N14368);
or OR4 (N17759, N17754, N9284, N11038, N7855);
or OR2 (N17760, N17744, N1341);
and AND4 (N17761, N17759, N1114, N13300, N3253);
or OR4 (N17762, N17758, N7805, N4170, N7725);
xor XOR2 (N17763, N17762, N177);
nor NOR4 (N17764, N17757, N1523, N7639, N10496);
and AND3 (N17765, N17742, N6640, N15755);
or OR3 (N17766, N17763, N2448, N15411);
buf BUF1 (N17767, N17765);
not NOT1 (N17768, N17764);
xor XOR2 (N17769, N17750, N6661);
nor NOR4 (N17770, N17768, N7491, N4569, N9304);
nand NAND4 (N17771, N17767, N3033, N8410, N5990);
nand NAND3 (N17772, N17769, N8227, N13905);
or OR4 (N17773, N17739, N10199, N4294, N16330);
or OR4 (N17774, N17770, N3444, N15192, N17280);
xor XOR2 (N17775, N17756, N11781);
not NOT1 (N17776, N17760);
xor XOR2 (N17777, N17766, N10214);
or OR4 (N17778, N17755, N17202, N395, N3466);
nand NAND2 (N17779, N17774, N6369);
xor XOR2 (N17780, N17778, N1982);
or OR3 (N17781, N17749, N10472, N13514);
xor XOR2 (N17782, N17771, N9542);
or OR2 (N17783, N17773, N16505);
nor NOR3 (N17784, N17782, N8280, N4531);
nand NAND3 (N17785, N17784, N13185, N10328);
nor NOR2 (N17786, N17783, N9347);
buf BUF1 (N17787, N17777);
xor XOR2 (N17788, N17779, N10245);
xor XOR2 (N17789, N17761, N15644);
buf BUF1 (N17790, N17787);
or OR4 (N17791, N17788, N4942, N5919, N14467);
nor NOR4 (N17792, N17790, N16668, N15100, N16633);
not NOT1 (N17793, N17786);
and AND4 (N17794, N17789, N2003, N14214, N8725);
not NOT1 (N17795, N17791);
or OR4 (N17796, N17780, N7113, N3768, N1874);
nand NAND2 (N17797, N17776, N12491);
buf BUF1 (N17798, N17797);
and AND2 (N17799, N17781, N6530);
or OR4 (N17800, N17796, N7345, N7292, N11772);
xor XOR2 (N17801, N17794, N2447);
or OR4 (N17802, N17798, N8776, N1844, N14720);
not NOT1 (N17803, N17801);
not NOT1 (N17804, N17792);
nor NOR4 (N17805, N17800, N4809, N11954, N6773);
and AND4 (N17806, N17799, N14654, N816, N16197);
not NOT1 (N17807, N17785);
nand NAND3 (N17808, N17806, N6159, N15018);
xor XOR2 (N17809, N17803, N16476);
and AND2 (N17810, N17795, N1451);
or OR4 (N17811, N17793, N10724, N758, N9714);
nand NAND4 (N17812, N17809, N11189, N8522, N3019);
or OR2 (N17813, N17810, N3036);
nand NAND2 (N17814, N17807, N14837);
buf BUF1 (N17815, N17775);
nand NAND2 (N17816, N17772, N9405);
xor XOR2 (N17817, N17804, N10017);
not NOT1 (N17818, N17812);
or OR4 (N17819, N17816, N9433, N5617, N16504);
buf BUF1 (N17820, N17817);
nor NOR4 (N17821, N17813, N16963, N3392, N1162);
or OR4 (N17822, N17818, N14696, N10239, N10815);
or OR2 (N17823, N17821, N6707);
nor NOR3 (N17824, N17822, N11897, N13888);
nor NOR4 (N17825, N17820, N8538, N9030, N14093);
and AND3 (N17826, N17814, N11561, N1764);
buf BUF1 (N17827, N17802);
xor XOR2 (N17828, N17826, N11585);
nand NAND3 (N17829, N17827, N14760, N6096);
and AND3 (N17830, N17805, N9148, N5432);
not NOT1 (N17831, N17825);
not NOT1 (N17832, N17819);
nand NAND4 (N17833, N17830, N13734, N11008, N16405);
nor NOR3 (N17834, N17811, N674, N16044);
or OR4 (N17835, N17824, N7785, N6265, N6590);
and AND2 (N17836, N17833, N7129);
xor XOR2 (N17837, N17828, N15097);
xor XOR2 (N17838, N17836, N14100);
buf BUF1 (N17839, N17837);
nor NOR2 (N17840, N17829, N8332);
or OR3 (N17841, N17840, N5914, N388);
not NOT1 (N17842, N17808);
not NOT1 (N17843, N17835);
not NOT1 (N17844, N17832);
not NOT1 (N17845, N17831);
nor NOR3 (N17846, N17823, N8893, N4341);
or OR4 (N17847, N17815, N17775, N11725, N17781);
nand NAND3 (N17848, N17844, N8531, N4617);
not NOT1 (N17849, N17846);
nand NAND2 (N17850, N17849, N3573);
buf BUF1 (N17851, N17843);
xor XOR2 (N17852, N17847, N7789);
xor XOR2 (N17853, N17848, N7878);
xor XOR2 (N17854, N17834, N8412);
buf BUF1 (N17855, N17838);
and AND3 (N17856, N17845, N13928, N4175);
and AND2 (N17857, N17854, N5119);
nor NOR2 (N17858, N17841, N6472);
not NOT1 (N17859, N17857);
or OR2 (N17860, N17856, N9715);
nand NAND4 (N17861, N17855, N11070, N1197, N7359);
nor NOR4 (N17862, N17850, N2998, N9933, N6369);
and AND3 (N17863, N17839, N4577, N9575);
buf BUF1 (N17864, N17842);
or OR4 (N17865, N17851, N13640, N5645, N8022);
nor NOR2 (N17866, N17858, N11830);
and AND2 (N17867, N17864, N4995);
nand NAND4 (N17868, N17862, N17129, N15703, N5673);
xor XOR2 (N17869, N17865, N2103);
nand NAND4 (N17870, N17863, N15723, N9384, N2525);
nand NAND4 (N17871, N17866, N12925, N2339, N15871);
not NOT1 (N17872, N17868);
xor XOR2 (N17873, N17859, N7769);
nand NAND2 (N17874, N17871, N17293);
not NOT1 (N17875, N17861);
not NOT1 (N17876, N17869);
and AND3 (N17877, N17873, N4085, N13683);
buf BUF1 (N17878, N17853);
and AND3 (N17879, N17860, N10521, N12893);
nand NAND2 (N17880, N17870, N1552);
nor NOR2 (N17881, N17877, N12295);
buf BUF1 (N17882, N17879);
buf BUF1 (N17883, N17852);
nor NOR4 (N17884, N17876, N10094, N15990, N2214);
and AND2 (N17885, N17867, N8229);
xor XOR2 (N17886, N17874, N3230);
and AND4 (N17887, N17880, N10324, N15953, N3802);
not NOT1 (N17888, N17887);
nand NAND3 (N17889, N17878, N4815, N11552);
or OR2 (N17890, N17872, N4367);
xor XOR2 (N17891, N17882, N7283);
xor XOR2 (N17892, N17888, N8512);
nor NOR4 (N17893, N17889, N7899, N8844, N213);
or OR4 (N17894, N17885, N1418, N8870, N17533);
nand NAND3 (N17895, N17893, N16919, N14817);
not NOT1 (N17896, N17884);
nor NOR2 (N17897, N17881, N2298);
or OR2 (N17898, N17896, N15537);
nor NOR3 (N17899, N17883, N13297, N11380);
xor XOR2 (N17900, N17875, N14055);
xor XOR2 (N17901, N17899, N13742);
nand NAND2 (N17902, N17894, N9117);
or OR3 (N17903, N17901, N13673, N12178);
xor XOR2 (N17904, N17903, N15385);
not NOT1 (N17905, N17902);
xor XOR2 (N17906, N17886, N3065);
nor NOR4 (N17907, N17895, N3993, N9638, N3112);
and AND2 (N17908, N17904, N7834);
buf BUF1 (N17909, N17907);
nor NOR4 (N17910, N17898, N171, N15449, N2792);
and AND3 (N17911, N17890, N911, N2444);
nand NAND4 (N17912, N17910, N9894, N17130, N4685);
not NOT1 (N17913, N17911);
nor NOR2 (N17914, N17891, N16512);
or OR4 (N17915, N17892, N8954, N711, N16143);
xor XOR2 (N17916, N17905, N4667);
nand NAND3 (N17917, N17900, N17900, N17622);
not NOT1 (N17918, N17909);
or OR3 (N17919, N17914, N3376, N3129);
xor XOR2 (N17920, N17913, N9188);
buf BUF1 (N17921, N17917);
buf BUF1 (N17922, N17916);
and AND2 (N17923, N17915, N17749);
nand NAND3 (N17924, N17922, N16125, N2553);
or OR4 (N17925, N17906, N11296, N12434, N3311);
xor XOR2 (N17926, N17920, N9538);
nand NAND2 (N17927, N17921, N7516);
nand NAND2 (N17928, N17925, N15163);
and AND4 (N17929, N17927, N1861, N4122, N14473);
xor XOR2 (N17930, N17926, N12487);
or OR4 (N17931, N17908, N10757, N15851, N9828);
xor XOR2 (N17932, N17919, N9764);
nor NOR2 (N17933, N17929, N3915);
not NOT1 (N17934, N17912);
not NOT1 (N17935, N17930);
or OR3 (N17936, N17935, N971, N6745);
and AND3 (N17937, N17933, N10950, N13425);
not NOT1 (N17938, N17928);
nand NAND4 (N17939, N17937, N5164, N4312, N17850);
not NOT1 (N17940, N17931);
xor XOR2 (N17941, N17923, N3288);
not NOT1 (N17942, N17936);
buf BUF1 (N17943, N17942);
buf BUF1 (N17944, N17932);
not NOT1 (N17945, N17924);
nor NOR3 (N17946, N17897, N13786, N3902);
nand NAND3 (N17947, N17938, N9360, N4651);
or OR3 (N17948, N17940, N13537, N12055);
and AND3 (N17949, N17918, N9042, N6929);
nand NAND4 (N17950, N17947, N12550, N4914, N4214);
or OR3 (N17951, N17946, N2848, N9035);
xor XOR2 (N17952, N17948, N14005);
buf BUF1 (N17953, N17949);
not NOT1 (N17954, N17950);
buf BUF1 (N17955, N17952);
nand NAND4 (N17956, N17939, N11914, N1717, N7572);
nor NOR4 (N17957, N17953, N16029, N9704, N2439);
and AND4 (N17958, N17956, N6968, N2565, N13016);
buf BUF1 (N17959, N17957);
and AND3 (N17960, N17943, N4964, N10726);
or OR3 (N17961, N17960, N5913, N17312);
nand NAND2 (N17962, N17954, N4761);
not NOT1 (N17963, N17941);
nor NOR3 (N17964, N17962, N10202, N2794);
not NOT1 (N17965, N17961);
or OR2 (N17966, N17965, N6211);
and AND2 (N17967, N17944, N11504);
and AND4 (N17968, N17955, N8371, N5478, N12934);
not NOT1 (N17969, N17958);
nor NOR3 (N17970, N17967, N772, N13033);
buf BUF1 (N17971, N17963);
xor XOR2 (N17972, N17970, N5121);
not NOT1 (N17973, N17972);
nor NOR3 (N17974, N17971, N10384, N12976);
or OR4 (N17975, N17974, N13408, N6161, N14704);
not NOT1 (N17976, N17973);
nand NAND2 (N17977, N17976, N1918);
nor NOR2 (N17978, N17964, N15233);
or OR3 (N17979, N17969, N9952, N17769);
nand NAND2 (N17980, N17978, N5199);
nor NOR2 (N17981, N17975, N1668);
nand NAND3 (N17982, N17979, N13765, N1414);
and AND2 (N17983, N17945, N10577);
buf BUF1 (N17984, N17977);
and AND3 (N17985, N17959, N15681, N9371);
xor XOR2 (N17986, N17985, N5332);
nor NOR3 (N17987, N17966, N16500, N6627);
nand NAND2 (N17988, N17982, N15903);
nor NOR3 (N17989, N17983, N7096, N5989);
not NOT1 (N17990, N17981);
not NOT1 (N17991, N17988);
xor XOR2 (N17992, N17987, N14721);
xor XOR2 (N17993, N17934, N13626);
xor XOR2 (N17994, N17986, N10354);
not NOT1 (N17995, N17990);
nor NOR3 (N17996, N17995, N15538, N9871);
or OR2 (N17997, N17989, N10680);
or OR3 (N17998, N17951, N8467, N1465);
and AND3 (N17999, N17996, N6532, N17532);
nand NAND2 (N18000, N17980, N973);
and AND3 (N18001, N18000, N2320, N758);
nor NOR3 (N18002, N17984, N4777, N13098);
not NOT1 (N18003, N17998);
nor NOR3 (N18004, N17997, N1744, N9490);
or OR2 (N18005, N17993, N8491);
nor NOR2 (N18006, N18001, N12880);
xor XOR2 (N18007, N17991, N14931);
xor XOR2 (N18008, N18003, N9508);
xor XOR2 (N18009, N18007, N11910);
and AND3 (N18010, N17999, N17244, N3516);
and AND2 (N18011, N18010, N48);
not NOT1 (N18012, N18002);
or OR4 (N18013, N18004, N5196, N7905, N13121);
nand NAND4 (N18014, N18013, N3446, N336, N11616);
buf BUF1 (N18015, N18009);
and AND2 (N18016, N18012, N14002);
and AND2 (N18017, N18014, N7780);
not NOT1 (N18018, N18017);
or OR4 (N18019, N18005, N6438, N16518, N8221);
buf BUF1 (N18020, N18008);
not NOT1 (N18021, N18018);
and AND2 (N18022, N18016, N14378);
not NOT1 (N18023, N18006);
nand NAND2 (N18024, N18021, N3456);
and AND2 (N18025, N18020, N10081);
nand NAND4 (N18026, N18015, N10644, N8996, N17734);
xor XOR2 (N18027, N18022, N10193);
xor XOR2 (N18028, N17992, N10759);
not NOT1 (N18029, N18026);
and AND2 (N18030, N18027, N4408);
and AND2 (N18031, N17968, N219);
not NOT1 (N18032, N18028);
not NOT1 (N18033, N18024);
nor NOR2 (N18034, N18011, N12693);
xor XOR2 (N18035, N18019, N16310);
xor XOR2 (N18036, N18025, N12952);
nand NAND3 (N18037, N18035, N9791, N15538);
nand NAND2 (N18038, N18031, N283);
not NOT1 (N18039, N18029);
nand NAND2 (N18040, N18034, N9939);
nand NAND2 (N18041, N18032, N2946);
and AND3 (N18042, N17994, N8709, N8424);
buf BUF1 (N18043, N18040);
buf BUF1 (N18044, N18038);
not NOT1 (N18045, N18030);
buf BUF1 (N18046, N18023);
or OR2 (N18047, N18044, N17452);
not NOT1 (N18048, N18045);
buf BUF1 (N18049, N18036);
xor XOR2 (N18050, N18041, N11423);
and AND2 (N18051, N18043, N7289);
not NOT1 (N18052, N18037);
buf BUF1 (N18053, N18050);
not NOT1 (N18054, N18052);
xor XOR2 (N18055, N18049, N14982);
not NOT1 (N18056, N18048);
or OR3 (N18057, N18042, N2707, N10538);
nand NAND4 (N18058, N18033, N16423, N6038, N4963);
not NOT1 (N18059, N18046);
or OR4 (N18060, N18055, N12930, N8030, N13964);
xor XOR2 (N18061, N18047, N5675);
not NOT1 (N18062, N18060);
buf BUF1 (N18063, N18053);
xor XOR2 (N18064, N18054, N6593);
and AND4 (N18065, N18039, N10585, N15137, N11441);
or OR3 (N18066, N18058, N9475, N10974);
nand NAND2 (N18067, N18057, N14718);
and AND2 (N18068, N18065, N13718);
nor NOR3 (N18069, N18062, N5659, N742);
not NOT1 (N18070, N18069);
and AND4 (N18071, N18064, N10635, N12792, N14766);
xor XOR2 (N18072, N18070, N5356);
not NOT1 (N18073, N18068);
buf BUF1 (N18074, N18061);
buf BUF1 (N18075, N18066);
nand NAND4 (N18076, N18051, N4266, N13467, N14096);
nand NAND2 (N18077, N18067, N15022);
buf BUF1 (N18078, N18071);
nand NAND2 (N18079, N18074, N9774);
buf BUF1 (N18080, N18073);
and AND2 (N18081, N18063, N14709);
not NOT1 (N18082, N18072);
xor XOR2 (N18083, N18080, N3322);
nand NAND4 (N18084, N18079, N15654, N4521, N14470);
xor XOR2 (N18085, N18081, N14305);
and AND4 (N18086, N18059, N15594, N10376, N13297);
nand NAND3 (N18087, N18082, N14546, N10102);
buf BUF1 (N18088, N18084);
xor XOR2 (N18089, N18075, N11238);
nor NOR2 (N18090, N18083, N13225);
and AND4 (N18091, N18088, N2287, N14972, N3665);
nand NAND3 (N18092, N18078, N8537, N8587);
nand NAND3 (N18093, N18087, N2968, N11543);
or OR3 (N18094, N18077, N4542, N2172);
xor XOR2 (N18095, N18089, N13521);
nor NOR4 (N18096, N18076, N3095, N13269, N7975);
or OR4 (N18097, N18096, N4431, N13106, N2936);
or OR2 (N18098, N18091, N14591);
xor XOR2 (N18099, N18095, N9641);
nand NAND3 (N18100, N18094, N8159, N8505);
and AND4 (N18101, N18090, N12124, N1435, N13335);
not NOT1 (N18102, N18098);
not NOT1 (N18103, N18101);
and AND2 (N18104, N18100, N3537);
and AND3 (N18105, N18093, N2648, N10431);
and AND3 (N18106, N18105, N5717, N2445);
not NOT1 (N18107, N18104);
not NOT1 (N18108, N18107);
buf BUF1 (N18109, N18108);
buf BUF1 (N18110, N18103);
and AND3 (N18111, N18099, N11954, N2251);
xor XOR2 (N18112, N18110, N11552);
nor NOR4 (N18113, N18106, N13685, N6424, N4230);
not NOT1 (N18114, N18097);
nor NOR4 (N18115, N18112, N1287, N15013, N17651);
and AND3 (N18116, N18056, N16310, N581);
and AND4 (N18117, N18102, N17558, N13241, N2698);
not NOT1 (N18118, N18115);
and AND3 (N18119, N18086, N15099, N16491);
not NOT1 (N18120, N18113);
not NOT1 (N18121, N18119);
or OR4 (N18122, N18114, N11959, N5504, N13031);
nor NOR4 (N18123, N18116, N9671, N18036, N15747);
and AND2 (N18124, N18092, N4648);
or OR3 (N18125, N18123, N4205, N17638);
buf BUF1 (N18126, N18125);
and AND3 (N18127, N18117, N14459, N15518);
nand NAND3 (N18128, N18085, N12071, N9393);
xor XOR2 (N18129, N18126, N11604);
nand NAND3 (N18130, N18128, N7663, N14295);
xor XOR2 (N18131, N18129, N2853);
buf BUF1 (N18132, N18130);
nor NOR4 (N18133, N18124, N4356, N54, N17489);
nor NOR3 (N18134, N18109, N17423, N5481);
nor NOR3 (N18135, N18134, N13178, N8413);
buf BUF1 (N18136, N18120);
and AND4 (N18137, N18135, N3561, N4431, N17447);
xor XOR2 (N18138, N18122, N131);
not NOT1 (N18139, N18118);
nand NAND4 (N18140, N18139, N16890, N1593, N16428);
or OR3 (N18141, N18127, N2079, N1526);
xor XOR2 (N18142, N18140, N6052);
nor NOR3 (N18143, N18111, N3562, N9700);
or OR2 (N18144, N18136, N4638);
nor NOR2 (N18145, N18142, N13575);
xor XOR2 (N18146, N18131, N14122);
not NOT1 (N18147, N18144);
nand NAND3 (N18148, N18137, N2014, N11428);
and AND4 (N18149, N18132, N12248, N3255, N3659);
not NOT1 (N18150, N18133);
or OR4 (N18151, N18141, N10385, N1757, N3);
xor XOR2 (N18152, N18147, N3364);
xor XOR2 (N18153, N18152, N15946);
or OR3 (N18154, N18150, N7018, N5194);
buf BUF1 (N18155, N18153);
buf BUF1 (N18156, N18151);
or OR3 (N18157, N18156, N3315, N10735);
nand NAND3 (N18158, N18121, N16225, N15956);
nand NAND3 (N18159, N18154, N11209, N13083);
buf BUF1 (N18160, N18148);
xor XOR2 (N18161, N18143, N1288);
or OR2 (N18162, N18157, N2647);
nor NOR4 (N18163, N18160, N14582, N9605, N3836);
nand NAND3 (N18164, N18161, N16009, N16454);
buf BUF1 (N18165, N18145);
buf BUF1 (N18166, N18163);
nand NAND3 (N18167, N18165, N12523, N8768);
not NOT1 (N18168, N18164);
buf BUF1 (N18169, N18138);
or OR2 (N18170, N18168, N17939);
not NOT1 (N18171, N18158);
and AND4 (N18172, N18155, N14696, N11542, N10459);
or OR2 (N18173, N18172, N5596);
buf BUF1 (N18174, N18171);
buf BUF1 (N18175, N18167);
nand NAND4 (N18176, N18173, N13514, N17799, N13499);
xor XOR2 (N18177, N18174, N9656);
nor NOR2 (N18178, N18162, N2932);
nor NOR2 (N18179, N18169, N2922);
nand NAND3 (N18180, N18146, N13331, N2967);
or OR2 (N18181, N18179, N10012);
and AND3 (N18182, N18175, N758, N3144);
nor NOR2 (N18183, N18178, N13842);
nand NAND2 (N18184, N18181, N6176);
xor XOR2 (N18185, N18183, N13938);
nor NOR3 (N18186, N18184, N14271, N13446);
not NOT1 (N18187, N18182);
xor XOR2 (N18188, N18176, N11028);
and AND2 (N18189, N18159, N16998);
not NOT1 (N18190, N18188);
or OR4 (N18191, N18189, N12101, N53, N16743);
or OR2 (N18192, N18166, N8482);
not NOT1 (N18193, N18191);
buf BUF1 (N18194, N18190);
buf BUF1 (N18195, N18180);
buf BUF1 (N18196, N18185);
nor NOR2 (N18197, N18186, N14833);
nand NAND2 (N18198, N18197, N8951);
nor NOR4 (N18199, N18149, N10552, N10153, N8815);
or OR3 (N18200, N18187, N11216, N16828);
nor NOR3 (N18201, N18192, N11636, N13937);
not NOT1 (N18202, N18193);
xor XOR2 (N18203, N18195, N11764);
buf BUF1 (N18204, N18196);
and AND2 (N18205, N18198, N9327);
xor XOR2 (N18206, N18199, N8422);
nand NAND2 (N18207, N18206, N17206);
and AND4 (N18208, N18177, N1084, N11069, N14293);
nand NAND4 (N18209, N18205, N9417, N4704, N15275);
not NOT1 (N18210, N18209);
not NOT1 (N18211, N18201);
and AND2 (N18212, N18194, N2109);
nand NAND4 (N18213, N18208, N15136, N10978, N9345);
buf BUF1 (N18214, N18204);
nand NAND4 (N18215, N18214, N13639, N7143, N2029);
nand NAND4 (N18216, N18213, N14573, N7078, N8229);
buf BUF1 (N18217, N18211);
xor XOR2 (N18218, N18170, N10172);
nor NOR4 (N18219, N18210, N733, N8850, N12098);
xor XOR2 (N18220, N18212, N1959);
buf BUF1 (N18221, N18218);
and AND2 (N18222, N18221, N8402);
or OR4 (N18223, N18200, N17477, N7307, N6550);
and AND3 (N18224, N18223, N15633, N4397);
nor NOR3 (N18225, N18216, N12501, N3756);
not NOT1 (N18226, N18217);
buf BUF1 (N18227, N18222);
or OR4 (N18228, N18224, N9634, N10040, N15456);
xor XOR2 (N18229, N18228, N7273);
not NOT1 (N18230, N18202);
xor XOR2 (N18231, N18225, N14202);
xor XOR2 (N18232, N18227, N12831);
and AND2 (N18233, N18220, N4728);
xor XOR2 (N18234, N18229, N6086);
and AND2 (N18235, N18232, N8566);
buf BUF1 (N18236, N18207);
or OR3 (N18237, N18231, N16115, N4596);
not NOT1 (N18238, N18234);
nand NAND3 (N18239, N18230, N5749, N5664);
xor XOR2 (N18240, N18215, N372);
nand NAND3 (N18241, N18219, N5082, N6524);
not NOT1 (N18242, N18238);
and AND4 (N18243, N18236, N16220, N16103, N8802);
not NOT1 (N18244, N18226);
buf BUF1 (N18245, N18237);
nand NAND4 (N18246, N18245, N2239, N444, N15628);
and AND4 (N18247, N18233, N10145, N1233, N10611);
nor NOR2 (N18248, N18239, N1876);
nor NOR3 (N18249, N18241, N10966, N7535);
not NOT1 (N18250, N18240);
and AND4 (N18251, N18235, N16376, N16400, N5994);
buf BUF1 (N18252, N18246);
nor NOR3 (N18253, N18243, N16515, N8744);
nor NOR2 (N18254, N18248, N14282);
and AND4 (N18255, N18242, N3478, N14811, N14461);
and AND4 (N18256, N18203, N4916, N5472, N2332);
nor NOR4 (N18257, N18244, N9562, N14991, N11224);
and AND4 (N18258, N18251, N11702, N3947, N3812);
or OR2 (N18259, N18249, N4844);
nand NAND3 (N18260, N18250, N4090, N9612);
nand NAND3 (N18261, N18247, N9942, N16497);
or OR4 (N18262, N18257, N3562, N10484, N234);
buf BUF1 (N18263, N18261);
and AND3 (N18264, N18253, N9900, N16812);
nor NOR2 (N18265, N18263, N2497);
not NOT1 (N18266, N18256);
not NOT1 (N18267, N18259);
buf BUF1 (N18268, N18258);
buf BUF1 (N18269, N18267);
buf BUF1 (N18270, N18252);
or OR3 (N18271, N18264, N8172, N10014);
or OR4 (N18272, N18265, N4898, N16230, N13386);
nor NOR3 (N18273, N18254, N792, N1264);
or OR2 (N18274, N18262, N5833);
xor XOR2 (N18275, N18273, N16906);
xor XOR2 (N18276, N18260, N3760);
buf BUF1 (N18277, N18270);
and AND3 (N18278, N18255, N16623, N15915);
buf BUF1 (N18279, N18276);
xor XOR2 (N18280, N18269, N3788);
nor NOR2 (N18281, N18275, N2041);
nand NAND4 (N18282, N18268, N8831, N13421, N11484);
nor NOR3 (N18283, N18280, N3147, N2468);
or OR2 (N18284, N18266, N14072);
xor XOR2 (N18285, N18272, N10513);
or OR3 (N18286, N18279, N10646, N2781);
nand NAND4 (N18287, N18282, N4842, N3842, N6090);
and AND2 (N18288, N18286, N8263);
nor NOR4 (N18289, N18285, N7053, N17668, N9456);
not NOT1 (N18290, N18287);
xor XOR2 (N18291, N18284, N10495);
not NOT1 (N18292, N18289);
nand NAND4 (N18293, N18278, N16120, N4118, N13163);
buf BUF1 (N18294, N18293);
or OR3 (N18295, N18288, N16749, N5921);
or OR2 (N18296, N18281, N16026);
nor NOR2 (N18297, N18283, N14030);
xor XOR2 (N18298, N18290, N4290);
xor XOR2 (N18299, N18295, N9895);
buf BUF1 (N18300, N18299);
xor XOR2 (N18301, N18274, N5715);
nor NOR2 (N18302, N18294, N2540);
nand NAND3 (N18303, N18298, N5773, N10322);
nand NAND3 (N18304, N18296, N17753, N17815);
not NOT1 (N18305, N18302);
nand NAND4 (N18306, N18291, N11710, N2523, N11135);
not NOT1 (N18307, N18300);
nand NAND3 (N18308, N18304, N9318, N15470);
or OR4 (N18309, N18308, N11730, N16506, N10706);
or OR4 (N18310, N18306, N11133, N3174, N11426);
nand NAND4 (N18311, N18303, N1104, N1283, N205);
or OR3 (N18312, N18307, N3789, N14863);
nand NAND4 (N18313, N18277, N3256, N5000, N14988);
nor NOR3 (N18314, N18301, N2042, N5095);
xor XOR2 (N18315, N18271, N7955);
buf BUF1 (N18316, N18315);
and AND4 (N18317, N18309, N7074, N8660, N16770);
or OR3 (N18318, N18314, N16410, N4240);
xor XOR2 (N18319, N18313, N13756);
xor XOR2 (N18320, N18312, N13874);
xor XOR2 (N18321, N18318, N368);
or OR2 (N18322, N18320, N11766);
and AND2 (N18323, N18292, N3791);
nand NAND2 (N18324, N18311, N13829);
not NOT1 (N18325, N18321);
nor NOR2 (N18326, N18310, N10836);
nor NOR4 (N18327, N18323, N7421, N15723, N44);
buf BUF1 (N18328, N18316);
not NOT1 (N18329, N18328);
not NOT1 (N18330, N18297);
not NOT1 (N18331, N18325);
not NOT1 (N18332, N18329);
and AND2 (N18333, N18332, N14063);
xor XOR2 (N18334, N18317, N7854);
nor NOR2 (N18335, N18333, N1417);
or OR4 (N18336, N18324, N4510, N18075, N8350);
buf BUF1 (N18337, N18336);
xor XOR2 (N18338, N18322, N3099);
nor NOR4 (N18339, N18335, N12514, N16936, N12028);
buf BUF1 (N18340, N18334);
xor XOR2 (N18341, N18326, N18036);
not NOT1 (N18342, N18339);
buf BUF1 (N18343, N18319);
buf BUF1 (N18344, N18340);
nor NOR2 (N18345, N18344, N17022);
and AND3 (N18346, N18342, N10405, N2648);
or OR2 (N18347, N18330, N2180);
not NOT1 (N18348, N18347);
nand NAND2 (N18349, N18327, N9530);
not NOT1 (N18350, N18346);
and AND3 (N18351, N18337, N13358, N16600);
nor NOR4 (N18352, N18345, N6766, N2372, N14397);
xor XOR2 (N18353, N18351, N10301);
and AND2 (N18354, N18352, N12502);
not NOT1 (N18355, N18350);
buf BUF1 (N18356, N18338);
nand NAND4 (N18357, N18305, N12386, N875, N904);
and AND3 (N18358, N18349, N11784, N13257);
nand NAND2 (N18359, N18355, N5755);
or OR4 (N18360, N18354, N18195, N3712, N907);
xor XOR2 (N18361, N18348, N8375);
buf BUF1 (N18362, N18341);
buf BUF1 (N18363, N18331);
and AND3 (N18364, N18356, N2690, N14184);
and AND4 (N18365, N18364, N1500, N12012, N2924);
and AND2 (N18366, N18361, N1990);
nor NOR3 (N18367, N18357, N13809, N3871);
nand NAND2 (N18368, N18365, N15075);
buf BUF1 (N18369, N18367);
nand NAND4 (N18370, N18366, N357, N17404, N6419);
or OR3 (N18371, N18360, N4876, N7554);
and AND3 (N18372, N18359, N15517, N12973);
buf BUF1 (N18373, N18343);
buf BUF1 (N18374, N18363);
nand NAND4 (N18375, N18362, N3580, N17546, N9149);
and AND4 (N18376, N18372, N8891, N1748, N14442);
and AND3 (N18377, N18370, N12842, N13270);
and AND4 (N18378, N18353, N167, N9452, N17485);
nand NAND3 (N18379, N18371, N5368, N9756);
buf BUF1 (N18380, N18368);
and AND3 (N18381, N18376, N10447, N13310);
nor NOR4 (N18382, N18377, N18077, N7478, N9353);
or OR2 (N18383, N18380, N16832);
nand NAND4 (N18384, N18369, N13282, N5321, N4665);
and AND3 (N18385, N18381, N12539, N3530);
not NOT1 (N18386, N18358);
not NOT1 (N18387, N18385);
not NOT1 (N18388, N18379);
nor NOR2 (N18389, N18384, N1579);
nor NOR2 (N18390, N18389, N8794);
or OR2 (N18391, N18375, N13213);
nand NAND3 (N18392, N18391, N611, N8252);
and AND3 (N18393, N18387, N12357, N5322);
or OR3 (N18394, N18390, N9564, N12686);
nor NOR3 (N18395, N18383, N14409, N11233);
not NOT1 (N18396, N18378);
and AND4 (N18397, N18388, N2336, N6769, N4756);
nor NOR3 (N18398, N18386, N10473, N11937);
xor XOR2 (N18399, N18393, N15668);
xor XOR2 (N18400, N18397, N3647);
or OR2 (N18401, N18394, N16396);
buf BUF1 (N18402, N18392);
and AND2 (N18403, N18373, N8899);
nand NAND3 (N18404, N18374, N10451, N5516);
not NOT1 (N18405, N18402);
buf BUF1 (N18406, N18403);
or OR2 (N18407, N18405, N4035);
not NOT1 (N18408, N18401);
not NOT1 (N18409, N18400);
buf BUF1 (N18410, N18407);
not NOT1 (N18411, N18408);
nand NAND3 (N18412, N18409, N12267, N10879);
not NOT1 (N18413, N18398);
not NOT1 (N18414, N18395);
xor XOR2 (N18415, N18413, N18336);
buf BUF1 (N18416, N18410);
and AND3 (N18417, N18382, N1549, N3812);
xor XOR2 (N18418, N18396, N7183);
nor NOR4 (N18419, N18415, N956, N5664, N8038);
xor XOR2 (N18420, N18414, N16840);
nand NAND2 (N18421, N18411, N8566);
nand NAND2 (N18422, N18420, N10178);
or OR2 (N18423, N18399, N5624);
not NOT1 (N18424, N18406);
buf BUF1 (N18425, N18419);
or OR2 (N18426, N18418, N17424);
or OR2 (N18427, N18426, N12842);
buf BUF1 (N18428, N18416);
and AND4 (N18429, N18412, N6737, N14736, N9609);
buf BUF1 (N18430, N18417);
or OR3 (N18431, N18427, N8667, N5796);
not NOT1 (N18432, N18430);
and AND2 (N18433, N18422, N12194);
and AND3 (N18434, N18424, N17849, N221);
nand NAND2 (N18435, N18404, N18288);
xor XOR2 (N18436, N18425, N11222);
buf BUF1 (N18437, N18421);
not NOT1 (N18438, N18431);
buf BUF1 (N18439, N18423);
not NOT1 (N18440, N18432);
nand NAND3 (N18441, N18436, N303, N1477);
nand NAND2 (N18442, N18429, N18224);
nor NOR3 (N18443, N18441, N8903, N274);
nor NOR4 (N18444, N18434, N12479, N14978, N17512);
nor NOR2 (N18445, N18438, N16063);
or OR4 (N18446, N18435, N1732, N6505, N8713);
nand NAND4 (N18447, N18444, N7197, N4552, N5309);
nand NAND3 (N18448, N18439, N17921, N11909);
and AND2 (N18449, N18437, N1058);
buf BUF1 (N18450, N18448);
and AND3 (N18451, N18428, N15168, N11156);
buf BUF1 (N18452, N18445);
not NOT1 (N18453, N18449);
nand NAND2 (N18454, N18442, N3113);
nor NOR2 (N18455, N18453, N13882);
not NOT1 (N18456, N18455);
nor NOR4 (N18457, N18440, N1593, N11707, N9241);
nor NOR3 (N18458, N18446, N4726, N50);
xor XOR2 (N18459, N18456, N10145);
xor XOR2 (N18460, N18452, N6629);
and AND4 (N18461, N18451, N10861, N15181, N4834);
nor NOR4 (N18462, N18457, N1010, N16319, N7657);
not NOT1 (N18463, N18458);
nor NOR4 (N18464, N18461, N8250, N11176, N12935);
nand NAND4 (N18465, N18460, N12559, N6084, N10278);
buf BUF1 (N18466, N18459);
nand NAND2 (N18467, N18454, N15794);
nand NAND4 (N18468, N18450, N5609, N6466, N82);
not NOT1 (N18469, N18462);
not NOT1 (N18470, N18465);
not NOT1 (N18471, N18467);
xor XOR2 (N18472, N18433, N7652);
nand NAND3 (N18473, N18469, N16532, N16858);
buf BUF1 (N18474, N18463);
or OR2 (N18475, N18474, N9127);
nor NOR4 (N18476, N18466, N11919, N10475, N7699);
xor XOR2 (N18477, N18473, N14748);
nand NAND3 (N18478, N18475, N5657, N4789);
nor NOR2 (N18479, N18472, N8592);
nor NOR4 (N18480, N18476, N3522, N17413, N14319);
nand NAND4 (N18481, N18443, N13156, N7305, N17361);
or OR2 (N18482, N18468, N11587);
buf BUF1 (N18483, N18464);
nor NOR2 (N18484, N18480, N8625);
not NOT1 (N18485, N18477);
xor XOR2 (N18486, N18484, N13408);
nand NAND3 (N18487, N18483, N7451, N2152);
nand NAND2 (N18488, N18487, N13766);
xor XOR2 (N18489, N18471, N12202);
or OR3 (N18490, N18485, N8434, N2880);
not NOT1 (N18491, N18481);
buf BUF1 (N18492, N18486);
not NOT1 (N18493, N18492);
nand NAND4 (N18494, N18482, N11776, N1870, N15534);
nor NOR2 (N18495, N18488, N12985);
and AND4 (N18496, N18495, N2718, N989, N12928);
nor NOR2 (N18497, N18470, N7981);
nand NAND4 (N18498, N18497, N7320, N12272, N16801);
xor XOR2 (N18499, N18490, N1746);
nor NOR4 (N18500, N18478, N697, N1391, N10267);
nand NAND2 (N18501, N18447, N12318);
and AND3 (N18502, N18500, N18347, N1651);
not NOT1 (N18503, N18499);
or OR2 (N18504, N18498, N1105);
xor XOR2 (N18505, N18491, N6343);
not NOT1 (N18506, N18501);
or OR4 (N18507, N18506, N17777, N5649, N15553);
not NOT1 (N18508, N18507);
nor NOR2 (N18509, N18493, N168);
and AND4 (N18510, N18508, N3540, N15159, N16434);
and AND2 (N18511, N18494, N2783);
not NOT1 (N18512, N18489);
and AND2 (N18513, N18503, N8904);
nand NAND4 (N18514, N18505, N13608, N4386, N10690);
or OR3 (N18515, N18479, N11913, N13910);
and AND2 (N18516, N18510, N5448);
xor XOR2 (N18517, N18502, N6512);
nand NAND4 (N18518, N18513, N4682, N15264, N13827);
and AND4 (N18519, N18518, N9194, N8451, N574);
nand NAND2 (N18520, N18512, N4611);
nand NAND3 (N18521, N18515, N2838, N14557);
buf BUF1 (N18522, N18509);
nand NAND4 (N18523, N18521, N9698, N5282, N3442);
nor NOR3 (N18524, N18522, N8772, N6961);
xor XOR2 (N18525, N18524, N15741);
buf BUF1 (N18526, N18525);
nor NOR2 (N18527, N18523, N10156);
or OR3 (N18528, N18517, N995, N8380);
not NOT1 (N18529, N18514);
xor XOR2 (N18530, N18520, N18156);
and AND3 (N18531, N18519, N16134, N6918);
xor XOR2 (N18532, N18504, N10804);
nor NOR2 (N18533, N18511, N16555);
or OR3 (N18534, N18526, N14164, N13459);
and AND2 (N18535, N18529, N1644);
xor XOR2 (N18536, N18531, N2778);
xor XOR2 (N18537, N18496, N13354);
nand NAND2 (N18538, N18536, N5020);
nand NAND4 (N18539, N18527, N3938, N996, N16835);
xor XOR2 (N18540, N18537, N1079);
xor XOR2 (N18541, N18532, N4791);
not NOT1 (N18542, N18540);
xor XOR2 (N18543, N18541, N10025);
or OR4 (N18544, N18539, N11395, N15574, N2862);
xor XOR2 (N18545, N18530, N16072);
not NOT1 (N18546, N18542);
and AND4 (N18547, N18543, N3470, N16977, N17367);
xor XOR2 (N18548, N18538, N7518);
nand NAND2 (N18549, N18546, N4284);
buf BUF1 (N18550, N18547);
nor NOR4 (N18551, N18545, N3491, N9700, N2804);
not NOT1 (N18552, N18534);
not NOT1 (N18553, N18549);
nand NAND4 (N18554, N18551, N10315, N3846, N16104);
buf BUF1 (N18555, N18553);
and AND4 (N18556, N18555, N9360, N11058, N10538);
buf BUF1 (N18557, N18556);
and AND2 (N18558, N18550, N1232);
nor NOR2 (N18559, N18557, N6965);
xor XOR2 (N18560, N18516, N10844);
nand NAND2 (N18561, N18548, N16585);
nor NOR4 (N18562, N18544, N15865, N3772, N17960);
not NOT1 (N18563, N18560);
buf BUF1 (N18564, N18561);
buf BUF1 (N18565, N18563);
xor XOR2 (N18566, N18535, N11594);
and AND4 (N18567, N18559, N11768, N613, N13818);
xor XOR2 (N18568, N18565, N11265);
and AND3 (N18569, N18533, N8192, N18050);
buf BUF1 (N18570, N18554);
and AND2 (N18571, N18528, N2444);
xor XOR2 (N18572, N18568, N16994);
not NOT1 (N18573, N18571);
nand NAND2 (N18574, N18573, N5757);
or OR4 (N18575, N18564, N18115, N15516, N6697);
nand NAND3 (N18576, N18569, N9465, N2262);
buf BUF1 (N18577, N18576);
nor NOR3 (N18578, N18575, N2171, N6031);
nand NAND2 (N18579, N18570, N16751);
xor XOR2 (N18580, N18572, N14861);
not NOT1 (N18581, N18577);
or OR4 (N18582, N18552, N14444, N3859, N9932);
buf BUF1 (N18583, N18558);
nand NAND4 (N18584, N18581, N11031, N2689, N8294);
nand NAND3 (N18585, N18580, N6802, N7624);
nand NAND4 (N18586, N18574, N15514, N12046, N12500);
and AND4 (N18587, N18562, N14673, N10755, N9284);
or OR3 (N18588, N18583, N5236, N4634);
and AND3 (N18589, N18587, N11883, N6660);
not NOT1 (N18590, N18579);
or OR2 (N18591, N18589, N17381);
or OR2 (N18592, N18585, N6783);
and AND2 (N18593, N18582, N11227);
or OR2 (N18594, N18592, N7358);
buf BUF1 (N18595, N18591);
not NOT1 (N18596, N18566);
not NOT1 (N18597, N18586);
nand NAND3 (N18598, N18590, N13723, N8808);
nand NAND2 (N18599, N18597, N14292);
nand NAND3 (N18600, N18567, N13053, N8919);
nand NAND3 (N18601, N18594, N17178, N3757);
not NOT1 (N18602, N18584);
and AND4 (N18603, N18598, N125, N10359, N11012);
xor XOR2 (N18604, N18596, N13455);
and AND3 (N18605, N18601, N10489, N11287);
buf BUF1 (N18606, N18600);
or OR4 (N18607, N18603, N6519, N8155, N16777);
nand NAND3 (N18608, N18578, N8963, N13459);
xor XOR2 (N18609, N18604, N16480);
or OR2 (N18610, N18602, N17714);
nand NAND4 (N18611, N18588, N27, N16199, N14277);
not NOT1 (N18612, N18595);
nand NAND2 (N18613, N18610, N7288);
or OR2 (N18614, N18608, N4018);
buf BUF1 (N18615, N18593);
buf BUF1 (N18616, N18611);
nor NOR2 (N18617, N18609, N4725);
nand NAND3 (N18618, N18614, N15239, N5442);
xor XOR2 (N18619, N18607, N18305);
nor NOR4 (N18620, N18605, N14219, N2586, N16711);
nor NOR2 (N18621, N18619, N17375);
nand NAND4 (N18622, N18616, N16819, N17421, N10725);
or OR4 (N18623, N18613, N3295, N1547, N9950);
and AND3 (N18624, N18599, N9988, N11800);
not NOT1 (N18625, N18612);
or OR2 (N18626, N18617, N9854);
xor XOR2 (N18627, N18615, N14950);
nand NAND2 (N18628, N18621, N420);
nor NOR4 (N18629, N18622, N8784, N9665, N13320);
not NOT1 (N18630, N18620);
and AND4 (N18631, N18624, N2972, N12474, N7150);
not NOT1 (N18632, N18618);
nand NAND4 (N18633, N18625, N12423, N12489, N8202);
nor NOR2 (N18634, N18606, N10000);
nand NAND3 (N18635, N18633, N13084, N3990);
or OR2 (N18636, N18629, N12200);
and AND4 (N18637, N18627, N9529, N16729, N3071);
nand NAND3 (N18638, N18634, N9364, N2626);
not NOT1 (N18639, N18628);
and AND2 (N18640, N18631, N5777);
nor NOR2 (N18641, N18632, N5446);
not NOT1 (N18642, N18630);
nor NOR3 (N18643, N18623, N8719, N4716);
xor XOR2 (N18644, N18639, N2524);
xor XOR2 (N18645, N18641, N907);
xor XOR2 (N18646, N18644, N10693);
not NOT1 (N18647, N18636);
or OR4 (N18648, N18647, N14568, N2085, N10785);
nor NOR4 (N18649, N18645, N15002, N1766, N5533);
nand NAND3 (N18650, N18635, N3309, N15000);
xor XOR2 (N18651, N18648, N14025);
buf BUF1 (N18652, N18643);
or OR2 (N18653, N18652, N12867);
buf BUF1 (N18654, N18638);
not NOT1 (N18655, N18626);
xor XOR2 (N18656, N18640, N2865);
not NOT1 (N18657, N18649);
and AND3 (N18658, N18650, N7710, N17918);
nand NAND4 (N18659, N18646, N15420, N4139, N4800);
not NOT1 (N18660, N18656);
nand NAND2 (N18661, N18651, N8865);
nor NOR2 (N18662, N18659, N17898);
nand NAND4 (N18663, N18642, N12155, N3711, N14284);
nand NAND2 (N18664, N18660, N10165);
not NOT1 (N18665, N18664);
not NOT1 (N18666, N18637);
and AND2 (N18667, N18655, N3945);
or OR4 (N18668, N18654, N10337, N5309, N16720);
or OR2 (N18669, N18668, N12346);
not NOT1 (N18670, N18653);
and AND3 (N18671, N18657, N10052, N8332);
nand NAND4 (N18672, N18662, N12904, N7204, N7642);
and AND3 (N18673, N18672, N3298, N6124);
xor XOR2 (N18674, N18663, N4486);
or OR2 (N18675, N18673, N16462);
buf BUF1 (N18676, N18671);
or OR4 (N18677, N18675, N5413, N14068, N15005);
buf BUF1 (N18678, N18661);
nand NAND4 (N18679, N18676, N9372, N17309, N16530);
buf BUF1 (N18680, N18665);
nand NAND2 (N18681, N18678, N7248);
nor NOR2 (N18682, N18669, N3088);
and AND3 (N18683, N18677, N11632, N3190);
xor XOR2 (N18684, N18670, N13731);
and AND4 (N18685, N18658, N16363, N1743, N7009);
or OR2 (N18686, N18680, N2013);
buf BUF1 (N18687, N18682);
xor XOR2 (N18688, N18674, N1715);
nor NOR2 (N18689, N18666, N16279);
or OR3 (N18690, N18689, N9733, N8992);
nand NAND4 (N18691, N18688, N3303, N14876, N9737);
and AND2 (N18692, N18684, N9339);
nor NOR3 (N18693, N18685, N4488, N15968);
xor XOR2 (N18694, N18679, N12584);
and AND2 (N18695, N18667, N13526);
and AND4 (N18696, N18686, N2560, N17184, N9214);
nand NAND4 (N18697, N18681, N16227, N3385, N16410);
and AND3 (N18698, N18694, N1646, N8998);
nor NOR3 (N18699, N18695, N3073, N2493);
nand NAND2 (N18700, N18691, N5496);
nand NAND2 (N18701, N18699, N18604);
buf BUF1 (N18702, N18696);
not NOT1 (N18703, N18697);
not NOT1 (N18704, N18700);
or OR3 (N18705, N18692, N5621, N14381);
xor XOR2 (N18706, N18704, N16330);
xor XOR2 (N18707, N18687, N4250);
not NOT1 (N18708, N18705);
or OR4 (N18709, N18708, N9626, N8930, N18451);
not NOT1 (N18710, N18706);
nand NAND4 (N18711, N18693, N4339, N17534, N13573);
nor NOR3 (N18712, N18701, N13793, N5802);
nand NAND4 (N18713, N18683, N12074, N17882, N11152);
and AND2 (N18714, N18707, N9796);
and AND2 (N18715, N18703, N12696);
nand NAND3 (N18716, N18710, N11879, N14923);
nand NAND3 (N18717, N18716, N18524, N16405);
buf BUF1 (N18718, N18712);
buf BUF1 (N18719, N18709);
nand NAND3 (N18720, N18690, N10764, N7067);
buf BUF1 (N18721, N18718);
or OR2 (N18722, N18713, N1967);
xor XOR2 (N18723, N18715, N9283);
xor XOR2 (N18724, N18714, N11424);
not NOT1 (N18725, N18698);
or OR2 (N18726, N18721, N911);
or OR3 (N18727, N18726, N9675, N14999);
nor NOR2 (N18728, N18727, N7093);
or OR3 (N18729, N18711, N1366, N7175);
xor XOR2 (N18730, N18722, N14753);
buf BUF1 (N18731, N18730);
buf BUF1 (N18732, N18717);
buf BUF1 (N18733, N18702);
nand NAND4 (N18734, N18728, N17395, N12466, N17859);
and AND2 (N18735, N18734, N1066);
and AND2 (N18736, N18731, N6303);
not NOT1 (N18737, N18735);
or OR2 (N18738, N18732, N16161);
not NOT1 (N18739, N18733);
or OR4 (N18740, N18725, N16803, N2295, N10621);
and AND3 (N18741, N18738, N3704, N8313);
and AND4 (N18742, N18740, N7240, N16056, N7641);
buf BUF1 (N18743, N18741);
or OR4 (N18744, N18724, N16754, N8399, N17606);
nand NAND3 (N18745, N18723, N9462, N16731);
xor XOR2 (N18746, N18719, N6458);
xor XOR2 (N18747, N18736, N7931);
nor NOR4 (N18748, N18742, N16797, N6460, N6459);
nand NAND3 (N18749, N18743, N2278, N7618);
not NOT1 (N18750, N18746);
nor NOR2 (N18751, N18749, N7986);
buf BUF1 (N18752, N18739);
xor XOR2 (N18753, N18751, N17591);
nor NOR3 (N18754, N18750, N10106, N9981);
or OR3 (N18755, N18753, N5739, N6357);
nand NAND3 (N18756, N18737, N1028, N11911);
nor NOR2 (N18757, N18744, N4167);
buf BUF1 (N18758, N18720);
nand NAND3 (N18759, N18755, N17882, N4522);
or OR4 (N18760, N18759, N17643, N15971, N11672);
xor XOR2 (N18761, N18754, N12574);
xor XOR2 (N18762, N18729, N2735);
xor XOR2 (N18763, N18760, N12214);
nand NAND2 (N18764, N18752, N10980);
or OR3 (N18765, N18764, N5669, N11855);
not NOT1 (N18766, N18758);
buf BUF1 (N18767, N18765);
nand NAND3 (N18768, N18748, N128, N16451);
or OR3 (N18769, N18745, N13498, N121);
xor XOR2 (N18770, N18756, N17471);
nand NAND4 (N18771, N18761, N18196, N7977, N2859);
nor NOR4 (N18772, N18763, N6626, N14409, N8146);
or OR3 (N18773, N18766, N10421, N18194);
or OR3 (N18774, N18772, N18539, N15459);
nor NOR2 (N18775, N18768, N14620);
not NOT1 (N18776, N18747);
nor NOR3 (N18777, N18773, N5844, N6376);
buf BUF1 (N18778, N18776);
and AND3 (N18779, N18757, N6382, N9903);
xor XOR2 (N18780, N18778, N4667);
or OR2 (N18781, N18769, N12484);
and AND2 (N18782, N18762, N9353);
not NOT1 (N18783, N18777);
xor XOR2 (N18784, N18774, N5820);
or OR3 (N18785, N18767, N17476, N9506);
buf BUF1 (N18786, N18771);
buf BUF1 (N18787, N18770);
or OR2 (N18788, N18787, N15166);
buf BUF1 (N18789, N18775);
not NOT1 (N18790, N18780);
xor XOR2 (N18791, N18786, N2561);
nand NAND4 (N18792, N18783, N16198, N4359, N4216);
buf BUF1 (N18793, N18791);
or OR4 (N18794, N18785, N552, N1924, N17423);
and AND4 (N18795, N18782, N2942, N5760, N13303);
nor NOR4 (N18796, N18789, N9107, N13857, N17724);
xor XOR2 (N18797, N18788, N11521);
or OR4 (N18798, N18779, N15919, N2086, N6708);
nand NAND2 (N18799, N18798, N11335);
buf BUF1 (N18800, N18792);
and AND3 (N18801, N18794, N13226, N350);
and AND4 (N18802, N18781, N4826, N6225, N10156);
nand NAND3 (N18803, N18793, N5224, N5609);
nand NAND2 (N18804, N18795, N14586);
not NOT1 (N18805, N18784);
nor NOR3 (N18806, N18803, N9940, N5201);
or OR3 (N18807, N18799, N13515, N3993);
xor XOR2 (N18808, N18800, N13502);
nor NOR2 (N18809, N18804, N2717);
and AND3 (N18810, N18805, N10373, N4442);
nor NOR2 (N18811, N18806, N8570);
or OR3 (N18812, N18808, N10677, N7257);
nor NOR4 (N18813, N18811, N9355, N12787, N1184);
not NOT1 (N18814, N18813);
not NOT1 (N18815, N18810);
not NOT1 (N18816, N18796);
not NOT1 (N18817, N18816);
nor NOR2 (N18818, N18812, N170);
and AND3 (N18819, N18814, N7316, N6233);
xor XOR2 (N18820, N18801, N3670);
and AND4 (N18821, N18807, N4250, N2833, N15946);
not NOT1 (N18822, N18809);
and AND4 (N18823, N18790, N6913, N11329, N16948);
nor NOR3 (N18824, N18820, N3781, N17038);
nand NAND2 (N18825, N18822, N4514);
xor XOR2 (N18826, N18823, N9793);
buf BUF1 (N18827, N18826);
nand NAND3 (N18828, N18802, N3155, N15370);
and AND3 (N18829, N18817, N15552, N13696);
or OR2 (N18830, N18797, N892);
and AND2 (N18831, N18827, N5230);
nand NAND4 (N18832, N18830, N7055, N2565, N11358);
xor XOR2 (N18833, N18815, N4276);
nand NAND2 (N18834, N18831, N12750);
buf BUF1 (N18835, N18825);
and AND2 (N18836, N18824, N11659);
xor XOR2 (N18837, N18835, N12110);
not NOT1 (N18838, N18818);
nor NOR4 (N18839, N18828, N17820, N16493, N13653);
nor NOR2 (N18840, N18834, N11222);
buf BUF1 (N18841, N18832);
nand NAND2 (N18842, N18833, N14464);
nor NOR4 (N18843, N18829, N18698, N9807, N8160);
and AND4 (N18844, N18836, N786, N17380, N4201);
nand NAND3 (N18845, N18839, N13644, N4073);
not NOT1 (N18846, N18837);
buf BUF1 (N18847, N18838);
nand NAND3 (N18848, N18843, N12734, N4202);
and AND3 (N18849, N18846, N7577, N4956);
not NOT1 (N18850, N18849);
not NOT1 (N18851, N18847);
or OR2 (N18852, N18840, N5584);
xor XOR2 (N18853, N18841, N11827);
and AND4 (N18854, N18844, N9446, N11788, N8925);
nor NOR4 (N18855, N18848, N9193, N11714, N14502);
or OR3 (N18856, N18852, N8797, N9327);
buf BUF1 (N18857, N18854);
nor NOR3 (N18858, N18853, N13013, N12203);
nand NAND2 (N18859, N18851, N17321);
not NOT1 (N18860, N18857);
not NOT1 (N18861, N18821);
or OR4 (N18862, N18858, N12535, N10407, N13025);
nand NAND4 (N18863, N18850, N7144, N3847, N4522);
nor NOR4 (N18864, N18855, N12418, N8016, N18736);
buf BUF1 (N18865, N18845);
xor XOR2 (N18866, N18859, N8382);
nor NOR3 (N18867, N18863, N11293, N5840);
or OR3 (N18868, N18819, N6288, N7220);
buf BUF1 (N18869, N18867);
buf BUF1 (N18870, N18856);
xor XOR2 (N18871, N18860, N472);
not NOT1 (N18872, N18870);
not NOT1 (N18873, N18872);
or OR3 (N18874, N18865, N9305, N15236);
nand NAND2 (N18875, N18873, N9435);
not NOT1 (N18876, N18871);
nand NAND3 (N18877, N18875, N1993, N3653);
nor NOR4 (N18878, N18842, N2423, N12703, N894);
buf BUF1 (N18879, N18876);
and AND4 (N18880, N18879, N17635, N5534, N6157);
nor NOR3 (N18881, N18861, N12942, N16484);
nor NOR4 (N18882, N18881, N17841, N10855, N15793);
not NOT1 (N18883, N18882);
or OR3 (N18884, N18868, N2590, N3947);
not NOT1 (N18885, N18884);
xor XOR2 (N18886, N18869, N17027);
nand NAND2 (N18887, N18885, N8065);
nand NAND2 (N18888, N18877, N6639);
and AND4 (N18889, N18888, N17159, N6278, N12456);
xor XOR2 (N18890, N18862, N966);
nor NOR4 (N18891, N18887, N12676, N9459, N1381);
nor NOR2 (N18892, N18878, N10603);
nor NOR3 (N18893, N18890, N15454, N2256);
not NOT1 (N18894, N18874);
nor NOR2 (N18895, N18883, N18179);
or OR4 (N18896, N18880, N15345, N7787, N6180);
buf BUF1 (N18897, N18894);
nand NAND3 (N18898, N18886, N9343, N16653);
xor XOR2 (N18899, N18889, N14656);
not NOT1 (N18900, N18891);
not NOT1 (N18901, N18893);
xor XOR2 (N18902, N18864, N8846);
or OR3 (N18903, N18898, N13967, N16010);
or OR4 (N18904, N18896, N12681, N1322, N2462);
xor XOR2 (N18905, N18866, N14427);
buf BUF1 (N18906, N18905);
or OR2 (N18907, N18906, N9781);
or OR2 (N18908, N18901, N6827);
nor NOR2 (N18909, N18900, N15837);
buf BUF1 (N18910, N18895);
nor NOR2 (N18911, N18892, N8709);
and AND3 (N18912, N18899, N18036, N7960);
xor XOR2 (N18913, N18910, N14795);
nand NAND4 (N18914, N18904, N15658, N13322, N15463);
nand NAND4 (N18915, N18913, N14044, N14123, N1337);
not NOT1 (N18916, N18902);
and AND3 (N18917, N18897, N1826, N12721);
or OR2 (N18918, N18912, N1715);
nor NOR2 (N18919, N18918, N7622);
or OR4 (N18920, N18908, N10603, N18763, N17377);
buf BUF1 (N18921, N18916);
or OR3 (N18922, N18907, N5914, N9175);
buf BUF1 (N18923, N18922);
nand NAND4 (N18924, N18909, N9297, N8215, N10526);
nand NAND4 (N18925, N18917, N7965, N16094, N7699);
buf BUF1 (N18926, N18914);
xor XOR2 (N18927, N18924, N18434);
xor XOR2 (N18928, N18915, N11608);
not NOT1 (N18929, N18927);
not NOT1 (N18930, N18928);
xor XOR2 (N18931, N18911, N14233);
nand NAND4 (N18932, N18919, N4952, N10917, N3385);
nor NOR4 (N18933, N18926, N11710, N14547, N4835);
buf BUF1 (N18934, N18931);
or OR4 (N18935, N18920, N2617, N5150, N10503);
or OR3 (N18936, N18921, N274, N400);
xor XOR2 (N18937, N18934, N15549);
nand NAND4 (N18938, N18923, N18261, N9865, N10026);
nor NOR2 (N18939, N18933, N7206);
not NOT1 (N18940, N18939);
and AND2 (N18941, N18929, N1339);
xor XOR2 (N18942, N18932, N14525);
xor XOR2 (N18943, N18938, N6827);
xor XOR2 (N18944, N18942, N8459);
not NOT1 (N18945, N18940);
nand NAND2 (N18946, N18935, N8482);
not NOT1 (N18947, N18944);
xor XOR2 (N18948, N18903, N14267);
xor XOR2 (N18949, N18947, N6947);
and AND2 (N18950, N18943, N6246);
buf BUF1 (N18951, N18946);
nor NOR2 (N18952, N18930, N15820);
or OR3 (N18953, N18950, N14644, N3334);
or OR3 (N18954, N18951, N3513, N11827);
and AND4 (N18955, N18953, N18065, N1674, N9327);
nor NOR3 (N18956, N18945, N10405, N5639);
or OR3 (N18957, N18956, N4160, N10638);
or OR2 (N18958, N18949, N2722);
or OR3 (N18959, N18958, N9621, N17086);
and AND2 (N18960, N18948, N11892);
nor NOR3 (N18961, N18937, N196, N13974);
nor NOR2 (N18962, N18954, N12819);
not NOT1 (N18963, N18925);
xor XOR2 (N18964, N18936, N11581);
nor NOR3 (N18965, N18959, N12434, N9668);
nand NAND3 (N18966, N18961, N16711, N14041);
nand NAND4 (N18967, N18960, N14439, N18879, N234);
not NOT1 (N18968, N18963);
nor NOR2 (N18969, N18962, N4343);
or OR4 (N18970, N18966, N8131, N7464, N6385);
or OR2 (N18971, N18941, N4217);
nor NOR3 (N18972, N18970, N3811, N13780);
and AND4 (N18973, N18972, N18790, N13343, N5174);
and AND2 (N18974, N18971, N8498);
buf BUF1 (N18975, N18967);
and AND2 (N18976, N18969, N14797);
nor NOR4 (N18977, N18952, N10005, N13317, N7626);
not NOT1 (N18978, N18975);
xor XOR2 (N18979, N18965, N2762);
xor XOR2 (N18980, N18964, N15007);
and AND3 (N18981, N18955, N4330, N8326);
and AND3 (N18982, N18974, N12518, N5241);
buf BUF1 (N18983, N18982);
not NOT1 (N18984, N18957);
and AND4 (N18985, N18973, N8159, N6469, N13435);
buf BUF1 (N18986, N18976);
xor XOR2 (N18987, N18986, N8788);
and AND2 (N18988, N18978, N10452);
or OR2 (N18989, N18977, N18124);
or OR3 (N18990, N18988, N7315, N3864);
nand NAND3 (N18991, N18984, N18432, N14856);
and AND3 (N18992, N18980, N10445, N5604);
nor NOR4 (N18993, N18989, N207, N18887, N4157);
and AND4 (N18994, N18983, N5385, N16842, N12906);
buf BUF1 (N18995, N18992);
not NOT1 (N18996, N18985);
buf BUF1 (N18997, N18990);
or OR3 (N18998, N18993, N7892, N7942);
buf BUF1 (N18999, N18979);
or OR3 (N19000, N18999, N15040, N15979);
or OR3 (N19001, N18994, N13130, N10265);
xor XOR2 (N19002, N18981, N7521);
buf BUF1 (N19003, N19001);
and AND2 (N19004, N18987, N8391);
buf BUF1 (N19005, N19002);
xor XOR2 (N19006, N18998, N13300);
not NOT1 (N19007, N19005);
buf BUF1 (N19008, N19007);
or OR4 (N19009, N18996, N10428, N14103, N15997);
and AND4 (N19010, N19008, N9141, N14928, N605);
not NOT1 (N19011, N19010);
or OR3 (N19012, N19011, N8032, N1436);
nand NAND3 (N19013, N19009, N1261, N8315);
nand NAND4 (N19014, N19004, N7927, N849, N8071);
not NOT1 (N19015, N19003);
nor NOR4 (N19016, N19013, N15974, N12862, N3135);
not NOT1 (N19017, N19014);
nor NOR4 (N19018, N18968, N10489, N589, N11344);
or OR4 (N19019, N19016, N8383, N17542, N11805);
xor XOR2 (N19020, N19012, N6534);
and AND4 (N19021, N19017, N416, N11755, N3297);
buf BUF1 (N19022, N18997);
xor XOR2 (N19023, N19006, N14531);
nand NAND2 (N19024, N18995, N4437);
xor XOR2 (N19025, N19018, N496);
and AND3 (N19026, N19020, N16668, N285);
nor NOR3 (N19027, N19022, N7319, N3918);
nor NOR2 (N19028, N19024, N12839);
buf BUF1 (N19029, N19026);
nand NAND2 (N19030, N19019, N8316);
buf BUF1 (N19031, N19023);
nand NAND4 (N19032, N19000, N18424, N3771, N11695);
xor XOR2 (N19033, N19021, N8442);
xor XOR2 (N19034, N19031, N3398);
not NOT1 (N19035, N19034);
xor XOR2 (N19036, N19025, N4890);
nand NAND2 (N19037, N19032, N3136);
xor XOR2 (N19038, N19027, N111);
or OR2 (N19039, N19033, N7818);
buf BUF1 (N19040, N19015);
nor NOR4 (N19041, N19037, N15702, N18843, N8671);
xor XOR2 (N19042, N19039, N14960);
buf BUF1 (N19043, N19035);
or OR4 (N19044, N19036, N14935, N2344, N3502);
not NOT1 (N19045, N19043);
buf BUF1 (N19046, N19044);
and AND4 (N19047, N19028, N10426, N5140, N5907);
nand NAND2 (N19048, N19038, N13207);
not NOT1 (N19049, N19048);
buf BUF1 (N19050, N19049);
not NOT1 (N19051, N18991);
not NOT1 (N19052, N19050);
nor NOR3 (N19053, N19042, N9412, N16139);
or OR3 (N19054, N19029, N15723, N18196);
buf BUF1 (N19055, N19030);
nor NOR2 (N19056, N19041, N6029);
nor NOR4 (N19057, N19056, N12668, N14927, N9660);
or OR2 (N19058, N19046, N6585);
or OR2 (N19059, N19047, N1180);
buf BUF1 (N19060, N19040);
xor XOR2 (N19061, N19057, N8324);
buf BUF1 (N19062, N19053);
nor NOR4 (N19063, N19062, N2437, N3440, N18298);
or OR3 (N19064, N19055, N5812, N546);
nand NAND2 (N19065, N19059, N3319);
nor NOR3 (N19066, N19065, N12984, N3397);
not NOT1 (N19067, N19060);
nor NOR2 (N19068, N19064, N14651);
xor XOR2 (N19069, N19054, N3375);
xor XOR2 (N19070, N19052, N1608);
or OR2 (N19071, N19070, N5866);
not NOT1 (N19072, N19066);
buf BUF1 (N19073, N19051);
not NOT1 (N19074, N19045);
buf BUF1 (N19075, N19069);
and AND4 (N19076, N19068, N19029, N5793, N13565);
and AND4 (N19077, N19058, N2228, N9740, N12557);
buf BUF1 (N19078, N19061);
nor NOR2 (N19079, N19076, N2181);
or OR3 (N19080, N19071, N15008, N18999);
buf BUF1 (N19081, N19075);
nand NAND2 (N19082, N19073, N7423);
buf BUF1 (N19083, N19081);
or OR3 (N19084, N19074, N9942, N15800);
not NOT1 (N19085, N19084);
or OR2 (N19086, N19067, N12213);
not NOT1 (N19087, N19077);
not NOT1 (N19088, N19085);
or OR2 (N19089, N19087, N13493);
nand NAND4 (N19090, N19079, N2194, N3130, N7422);
nand NAND2 (N19091, N19089, N3460);
nand NAND2 (N19092, N19072, N17716);
or OR4 (N19093, N19088, N5585, N17375, N8311);
buf BUF1 (N19094, N19082);
nor NOR4 (N19095, N19080, N3730, N18176, N2551);
nand NAND3 (N19096, N19094, N15496, N6419);
xor XOR2 (N19097, N19086, N14323);
nand NAND3 (N19098, N19092, N1832, N5751);
nand NAND3 (N19099, N19063, N3441, N10572);
or OR3 (N19100, N19098, N1686, N4475);
or OR4 (N19101, N19097, N15334, N3431, N8358);
nor NOR2 (N19102, N19095, N711);
not NOT1 (N19103, N19083);
nand NAND4 (N19104, N19096, N11167, N5771, N17217);
nor NOR3 (N19105, N19078, N13663, N2780);
or OR2 (N19106, N19090, N15367);
xor XOR2 (N19107, N19102, N3528);
and AND3 (N19108, N19099, N16392, N13184);
nand NAND4 (N19109, N19105, N7368, N16246, N14337);
nand NAND3 (N19110, N19109, N5773, N16440);
xor XOR2 (N19111, N19107, N13550);
nor NOR3 (N19112, N19091, N666, N7787);
nor NOR2 (N19113, N19103, N11120);
and AND4 (N19114, N19100, N5094, N12770, N9742);
buf BUF1 (N19115, N19104);
nand NAND2 (N19116, N19112, N4828);
xor XOR2 (N19117, N19113, N15711);
nand NAND3 (N19118, N19116, N13766, N13308);
nand NAND3 (N19119, N19093, N2363, N13122);
and AND4 (N19120, N19108, N18132, N10219, N15086);
buf BUF1 (N19121, N19111);
nor NOR3 (N19122, N19106, N17800, N17475);
nand NAND4 (N19123, N19121, N4292, N11762, N7196);
not NOT1 (N19124, N19110);
xor XOR2 (N19125, N19115, N10253);
and AND4 (N19126, N19124, N10362, N15614, N5633);
nor NOR2 (N19127, N19117, N13157);
and AND2 (N19128, N19120, N11062);
and AND4 (N19129, N19122, N9388, N13908, N12621);
or OR4 (N19130, N19126, N6257, N9025, N11141);
buf BUF1 (N19131, N19125);
buf BUF1 (N19132, N19128);
xor XOR2 (N19133, N19130, N7539);
not NOT1 (N19134, N19127);
or OR4 (N19135, N19114, N645, N2280, N8223);
or OR2 (N19136, N19129, N12416);
or OR4 (N19137, N19131, N7448, N11862, N13778);
or OR3 (N19138, N19119, N16932, N17935);
and AND4 (N19139, N19123, N1393, N964, N1901);
nor NOR4 (N19140, N19133, N1341, N2040, N9350);
xor XOR2 (N19141, N19138, N2045);
xor XOR2 (N19142, N19137, N16661);
nand NAND2 (N19143, N19136, N19132);
nand NAND3 (N19144, N15280, N1766, N17786);
buf BUF1 (N19145, N19139);
or OR2 (N19146, N19141, N17925);
buf BUF1 (N19147, N19135);
not NOT1 (N19148, N19144);
nor NOR2 (N19149, N19101, N9093);
nand NAND2 (N19150, N19148, N7405);
xor XOR2 (N19151, N19145, N13119);
nor NOR3 (N19152, N19118, N4056, N370);
nand NAND2 (N19153, N19134, N1885);
not NOT1 (N19154, N19143);
and AND2 (N19155, N19151, N9762);
nor NOR2 (N19156, N19149, N5855);
and AND2 (N19157, N19152, N1368);
nor NOR2 (N19158, N19147, N15515);
and AND3 (N19159, N19150, N2561, N2994);
not NOT1 (N19160, N19142);
nor NOR3 (N19161, N19155, N5829, N1095);
and AND2 (N19162, N19156, N8583);
and AND4 (N19163, N19162, N16132, N15963, N10431);
nand NAND3 (N19164, N19161, N3225, N5983);
xor XOR2 (N19165, N19159, N8544);
nor NOR2 (N19166, N19154, N8777);
nor NOR3 (N19167, N19163, N8991, N5188);
or OR3 (N19168, N19166, N2407, N9053);
not NOT1 (N19169, N19167);
or OR2 (N19170, N19168, N11907);
nand NAND4 (N19171, N19146, N474, N6614, N2424);
and AND2 (N19172, N19160, N6714);
buf BUF1 (N19173, N19171);
or OR2 (N19174, N19140, N10839);
buf BUF1 (N19175, N19170);
not NOT1 (N19176, N19164);
nor NOR4 (N19177, N19175, N15876, N12358, N11274);
nand NAND3 (N19178, N19158, N857, N11277);
and AND3 (N19179, N19176, N4876, N8477);
buf BUF1 (N19180, N19178);
nor NOR2 (N19181, N19179, N10288);
or OR4 (N19182, N19165, N10573, N15603, N3768);
or OR2 (N19183, N19153, N1623);
nor NOR4 (N19184, N19169, N14841, N14618, N12621);
nand NAND2 (N19185, N19184, N16965);
nor NOR4 (N19186, N19181, N9462, N14969, N7725);
xor XOR2 (N19187, N19180, N16655);
or OR2 (N19188, N19174, N12883);
or OR2 (N19189, N19185, N11948);
xor XOR2 (N19190, N19182, N18504);
nor NOR2 (N19191, N19172, N11683);
not NOT1 (N19192, N19191);
and AND4 (N19193, N19177, N19069, N18930, N4972);
nor NOR2 (N19194, N19188, N5747);
or OR2 (N19195, N19183, N3459);
or OR2 (N19196, N19186, N11023);
buf BUF1 (N19197, N19195);
xor XOR2 (N19198, N19194, N8395);
buf BUF1 (N19199, N19189);
or OR4 (N19200, N19190, N9896, N6829, N17978);
or OR3 (N19201, N19187, N7739, N1301);
not NOT1 (N19202, N19173);
or OR2 (N19203, N19201, N2996);
nand NAND3 (N19204, N19157, N10332, N6528);
or OR2 (N19205, N19196, N7225);
nor NOR3 (N19206, N19197, N16161, N5532);
or OR4 (N19207, N19200, N5264, N13257, N10912);
or OR3 (N19208, N19203, N9463, N12600);
buf BUF1 (N19209, N19207);
buf BUF1 (N19210, N19209);
or OR2 (N19211, N19204, N19189);
and AND3 (N19212, N19199, N13001, N16061);
buf BUF1 (N19213, N19202);
and AND3 (N19214, N19213, N13117, N7980);
and AND3 (N19215, N19208, N4299, N8773);
xor XOR2 (N19216, N19193, N11793);
not NOT1 (N19217, N19215);
nor NOR2 (N19218, N19217, N13390);
and AND4 (N19219, N19212, N11270, N1224, N7096);
nor NOR4 (N19220, N19216, N18503, N3230, N7731);
nand NAND4 (N19221, N19219, N9609, N8073, N16117);
not NOT1 (N19222, N19220);
and AND3 (N19223, N19198, N14425, N257);
xor XOR2 (N19224, N19218, N10235);
xor XOR2 (N19225, N19211, N4388);
buf BUF1 (N19226, N19192);
nor NOR2 (N19227, N19223, N1534);
or OR3 (N19228, N19222, N8200, N11365);
nor NOR3 (N19229, N19226, N17603, N16359);
or OR2 (N19230, N19227, N13115);
or OR3 (N19231, N19214, N564, N5533);
or OR3 (N19232, N19230, N18118, N18715);
buf BUF1 (N19233, N19232);
and AND4 (N19234, N19229, N16840, N16425, N2464);
nand NAND4 (N19235, N19228, N16521, N4853, N7123);
nor NOR4 (N19236, N19224, N6703, N1583, N111);
or OR4 (N19237, N19210, N3865, N10705, N5381);
nor NOR3 (N19238, N19205, N6444, N15345);
buf BUF1 (N19239, N19231);
nand NAND4 (N19240, N19239, N11161, N3637, N14422);
or OR4 (N19241, N19225, N12020, N6147, N4244);
not NOT1 (N19242, N19241);
xor XOR2 (N19243, N19233, N448);
not NOT1 (N19244, N19240);
xor XOR2 (N19245, N19244, N497);
nor NOR2 (N19246, N19206, N18245);
xor XOR2 (N19247, N19238, N6838);
nor NOR4 (N19248, N19235, N6248, N1389, N10016);
buf BUF1 (N19249, N19237);
buf BUF1 (N19250, N19242);
xor XOR2 (N19251, N19246, N15317);
nand NAND3 (N19252, N19234, N7258, N13108);
nor NOR4 (N19253, N19243, N7518, N4376, N17081);
not NOT1 (N19254, N19249);
buf BUF1 (N19255, N19253);
not NOT1 (N19256, N19236);
or OR4 (N19257, N19245, N11136, N407, N1873);
nor NOR2 (N19258, N19255, N18798);
not NOT1 (N19259, N19247);
buf BUF1 (N19260, N19221);
xor XOR2 (N19261, N19258, N11739);
or OR2 (N19262, N19254, N3962);
buf BUF1 (N19263, N19260);
xor XOR2 (N19264, N19251, N11756);
buf BUF1 (N19265, N19250);
or OR2 (N19266, N19259, N6126);
not NOT1 (N19267, N19257);
nor NOR4 (N19268, N19263, N11384, N10996, N15690);
nand NAND2 (N19269, N19268, N5381);
or OR3 (N19270, N19265, N1860, N4090);
xor XOR2 (N19271, N19252, N3287);
not NOT1 (N19272, N19262);
nor NOR4 (N19273, N19261, N11077, N18524, N7149);
and AND2 (N19274, N19256, N3262);
xor XOR2 (N19275, N19272, N7468);
xor XOR2 (N19276, N19274, N16474);
not NOT1 (N19277, N19275);
nand NAND4 (N19278, N19266, N16125, N8576, N12593);
xor XOR2 (N19279, N19273, N6589);
buf BUF1 (N19280, N19270);
not NOT1 (N19281, N19271);
nand NAND2 (N19282, N19267, N914);
xor XOR2 (N19283, N19276, N15406);
nor NOR3 (N19284, N19277, N9853, N447);
or OR3 (N19285, N19248, N2465, N9199);
nor NOR4 (N19286, N19281, N15982, N979, N10709);
and AND3 (N19287, N19284, N3814, N2832);
xor XOR2 (N19288, N19280, N12972);
not NOT1 (N19289, N19287);
or OR4 (N19290, N19264, N2146, N13222, N11297);
or OR2 (N19291, N19282, N15233);
buf BUF1 (N19292, N19286);
not NOT1 (N19293, N19288);
or OR3 (N19294, N19289, N5933, N828);
or OR2 (N19295, N19285, N5350);
not NOT1 (N19296, N19290);
or OR4 (N19297, N19278, N10195, N14135, N10130);
and AND3 (N19298, N19297, N1825, N16630);
nor NOR3 (N19299, N19291, N1482, N4234);
nand NAND3 (N19300, N19296, N16193, N16331);
not NOT1 (N19301, N19298);
not NOT1 (N19302, N19299);
xor XOR2 (N19303, N19294, N18742);
nor NOR4 (N19304, N19303, N16345, N9458, N18858);
or OR3 (N19305, N19300, N4299, N5497);
nand NAND4 (N19306, N19295, N19093, N14467, N3617);
and AND2 (N19307, N19292, N4520);
not NOT1 (N19308, N19269);
and AND3 (N19309, N19302, N12149, N10031);
nor NOR2 (N19310, N19304, N16197);
nor NOR3 (N19311, N19306, N6252, N2164);
nand NAND2 (N19312, N19293, N2697);
not NOT1 (N19313, N19301);
and AND4 (N19314, N19308, N3568, N3249, N3218);
or OR3 (N19315, N19314, N8107, N10217);
xor XOR2 (N19316, N19305, N3261);
xor XOR2 (N19317, N19279, N1035);
or OR2 (N19318, N19310, N6913);
not NOT1 (N19319, N19315);
nor NOR2 (N19320, N19311, N2359);
nor NOR4 (N19321, N19319, N13883, N1245, N10939);
nand NAND3 (N19322, N19312, N5785, N3261);
xor XOR2 (N19323, N19320, N18460);
and AND2 (N19324, N19317, N5648);
nor NOR3 (N19325, N19283, N15555, N7801);
and AND4 (N19326, N19321, N14158, N363, N8532);
nand NAND3 (N19327, N19309, N15686, N10848);
nor NOR4 (N19328, N19316, N16742, N18292, N17656);
nand NAND2 (N19329, N19328, N12923);
xor XOR2 (N19330, N19329, N4406);
or OR3 (N19331, N19326, N14518, N12227);
nand NAND4 (N19332, N19325, N9514, N10016, N1791);
or OR2 (N19333, N19322, N18885);
nand NAND2 (N19334, N19307, N14229);
xor XOR2 (N19335, N19327, N10090);
buf BUF1 (N19336, N19324);
xor XOR2 (N19337, N19333, N11283);
nand NAND2 (N19338, N19337, N13624);
not NOT1 (N19339, N19338);
or OR4 (N19340, N19318, N15802, N9237, N7594);
nor NOR2 (N19341, N19332, N10968);
nand NAND2 (N19342, N19331, N8292);
or OR2 (N19343, N19340, N16068);
nand NAND3 (N19344, N19339, N6330, N7768);
or OR3 (N19345, N19342, N16630, N3033);
xor XOR2 (N19346, N19335, N15096);
nor NOR4 (N19347, N19336, N1172, N9951, N13582);
nand NAND4 (N19348, N19330, N18757, N4177, N8999);
not NOT1 (N19349, N19346);
and AND4 (N19350, N19343, N15059, N6892, N7641);
or OR2 (N19351, N19349, N14490);
nand NAND3 (N19352, N19323, N11481, N15325);
nand NAND2 (N19353, N19348, N653);
nor NOR4 (N19354, N19352, N17801, N6833, N5452);
buf BUF1 (N19355, N19347);
buf BUF1 (N19356, N19350);
buf BUF1 (N19357, N19341);
not NOT1 (N19358, N19345);
or OR2 (N19359, N19351, N16592);
nor NOR2 (N19360, N19313, N14137);
not NOT1 (N19361, N19355);
xor XOR2 (N19362, N19353, N5823);
or OR4 (N19363, N19356, N9604, N10913, N18247);
nand NAND2 (N19364, N19359, N17063);
nor NOR3 (N19365, N19360, N4615, N11069);
nand NAND3 (N19366, N19365, N17968, N15571);
and AND3 (N19367, N19357, N8024, N9425);
nand NAND2 (N19368, N19361, N7098);
and AND2 (N19369, N19368, N15279);
or OR4 (N19370, N19344, N12153, N10361, N15431);
buf BUF1 (N19371, N19334);
and AND4 (N19372, N19367, N6182, N8208, N7957);
buf BUF1 (N19373, N19369);
and AND4 (N19374, N19366, N123, N4095, N1242);
xor XOR2 (N19375, N19373, N10860);
nor NOR2 (N19376, N19374, N18325);
not NOT1 (N19377, N19358);
xor XOR2 (N19378, N19371, N12020);
xor XOR2 (N19379, N19363, N7863);
nor NOR3 (N19380, N19377, N13607, N13150);
and AND4 (N19381, N19354, N2373, N906, N112);
buf BUF1 (N19382, N19372);
buf BUF1 (N19383, N19364);
or OR4 (N19384, N19383, N4302, N8976, N14107);
and AND4 (N19385, N19362, N16812, N18207, N5947);
buf BUF1 (N19386, N19378);
nand NAND4 (N19387, N19381, N6512, N19273, N17909);
not NOT1 (N19388, N19385);
nor NOR4 (N19389, N19370, N16176, N6621, N17682);
nor NOR3 (N19390, N19376, N10438, N7823);
and AND3 (N19391, N19380, N1512, N14058);
not NOT1 (N19392, N19379);
buf BUF1 (N19393, N19391);
or OR2 (N19394, N19389, N14595);
nor NOR4 (N19395, N19392, N16043, N18592, N2387);
not NOT1 (N19396, N19388);
xor XOR2 (N19397, N19394, N9350);
not NOT1 (N19398, N19390);
or OR4 (N19399, N19398, N2821, N16184, N9056);
not NOT1 (N19400, N19384);
and AND2 (N19401, N19399, N1809);
or OR2 (N19402, N19386, N14152);
xor XOR2 (N19403, N19382, N3845);
or OR2 (N19404, N19375, N1819);
nand NAND2 (N19405, N19400, N17464);
or OR4 (N19406, N19387, N12986, N12045, N9673);
or OR4 (N19407, N19406, N16846, N6481, N9077);
xor XOR2 (N19408, N19404, N11408);
buf BUF1 (N19409, N19405);
buf BUF1 (N19410, N19402);
not NOT1 (N19411, N19403);
and AND2 (N19412, N19401, N8031);
buf BUF1 (N19413, N19393);
nor NOR2 (N19414, N19410, N16519);
nand NAND4 (N19415, N19395, N2541, N15439, N11725);
nor NOR2 (N19416, N19408, N3833);
nand NAND3 (N19417, N19413, N13793, N7752);
buf BUF1 (N19418, N19417);
nor NOR2 (N19419, N19407, N13608);
nand NAND4 (N19420, N19396, N2957, N18850, N9408);
or OR3 (N19421, N19411, N17244, N5861);
nor NOR4 (N19422, N19420, N13010, N17954, N17669);
nor NOR3 (N19423, N19418, N19315, N10941);
and AND2 (N19424, N19409, N12539);
nor NOR2 (N19425, N19421, N10864);
xor XOR2 (N19426, N19416, N13270);
buf BUF1 (N19427, N19415);
not NOT1 (N19428, N19425);
nor NOR4 (N19429, N19428, N14122, N8756, N16534);
nor NOR4 (N19430, N19422, N13577, N8710, N5885);
buf BUF1 (N19431, N19430);
xor XOR2 (N19432, N19424, N16539);
buf BUF1 (N19433, N19431);
xor XOR2 (N19434, N19414, N9905);
buf BUF1 (N19435, N19423);
xor XOR2 (N19436, N19397, N1170);
or OR2 (N19437, N19433, N2706);
nor NOR4 (N19438, N19437, N843, N8318, N2650);
nor NOR4 (N19439, N19432, N3880, N10389, N6194);
buf BUF1 (N19440, N19429);
not NOT1 (N19441, N19439);
nor NOR4 (N19442, N19441, N18197, N7161, N13267);
buf BUF1 (N19443, N19438);
nand NAND4 (N19444, N19436, N3432, N7889, N5775);
or OR3 (N19445, N19442, N11073, N4206);
or OR2 (N19446, N19443, N7344);
or OR3 (N19447, N19444, N7012, N11400);
xor XOR2 (N19448, N19426, N13974);
or OR2 (N19449, N19447, N18062);
nand NAND3 (N19450, N19427, N15251, N2259);
not NOT1 (N19451, N19448);
buf BUF1 (N19452, N19445);
and AND2 (N19453, N19451, N6553);
xor XOR2 (N19454, N19449, N6065);
xor XOR2 (N19455, N19450, N14731);
xor XOR2 (N19456, N19412, N4896);
nor NOR2 (N19457, N19456, N6330);
xor XOR2 (N19458, N19452, N7606);
and AND2 (N19459, N19419, N10753);
or OR3 (N19460, N19457, N16588, N15673);
xor XOR2 (N19461, N19435, N18714);
nand NAND2 (N19462, N19440, N18621);
xor XOR2 (N19463, N19455, N17730);
xor XOR2 (N19464, N19459, N18963);
or OR3 (N19465, N19453, N4565, N19119);
nor NOR4 (N19466, N19462, N18083, N17732, N3962);
or OR4 (N19467, N19463, N13919, N3781, N7515);
not NOT1 (N19468, N19454);
buf BUF1 (N19469, N19466);
not NOT1 (N19470, N19468);
and AND3 (N19471, N19464, N13177, N11058);
not NOT1 (N19472, N19465);
buf BUF1 (N19473, N19446);
not NOT1 (N19474, N19473);
xor XOR2 (N19475, N19467, N9659);
nand NAND2 (N19476, N19434, N226);
xor XOR2 (N19477, N19472, N19048);
not NOT1 (N19478, N19469);
buf BUF1 (N19479, N19474);
nand NAND3 (N19480, N19479, N3615, N15043);
not NOT1 (N19481, N19460);
not NOT1 (N19482, N19458);
nand NAND4 (N19483, N19480, N2858, N14313, N1153);
nand NAND3 (N19484, N19477, N15234, N1414);
or OR2 (N19485, N19484, N3560);
and AND2 (N19486, N19478, N19351);
nand NAND2 (N19487, N19471, N16154);
or OR4 (N19488, N19487, N18863, N12270, N11922);
or OR3 (N19489, N19475, N18421, N5391);
nor NOR3 (N19490, N19476, N11644, N16890);
nor NOR4 (N19491, N19482, N4003, N19455, N692);
not NOT1 (N19492, N19470);
buf BUF1 (N19493, N19491);
nor NOR3 (N19494, N19490, N19379, N13345);
nor NOR3 (N19495, N19481, N690, N19475);
nand NAND4 (N19496, N19488, N5012, N16359, N5359);
nor NOR3 (N19497, N19495, N17468, N8013);
and AND2 (N19498, N19486, N6824);
buf BUF1 (N19499, N19485);
xor XOR2 (N19500, N19498, N16398);
nor NOR2 (N19501, N19483, N14199);
xor XOR2 (N19502, N19496, N13789);
buf BUF1 (N19503, N19461);
not NOT1 (N19504, N19501);
and AND4 (N19505, N19492, N17420, N12254, N2163);
nor NOR3 (N19506, N19504, N2765, N5606);
and AND4 (N19507, N19502, N8346, N16745, N14804);
nand NAND4 (N19508, N19494, N10281, N2541, N10381);
buf BUF1 (N19509, N19499);
and AND2 (N19510, N19507, N3267);
xor XOR2 (N19511, N19503, N15058);
or OR2 (N19512, N19489, N7949);
and AND3 (N19513, N19512, N731, N11688);
xor XOR2 (N19514, N19513, N11509);
or OR3 (N19515, N19511, N7815, N19101);
and AND3 (N19516, N19505, N4808, N6387);
xor XOR2 (N19517, N19500, N10895);
and AND4 (N19518, N19515, N7710, N5287, N4859);
not NOT1 (N19519, N19518);
buf BUF1 (N19520, N19517);
buf BUF1 (N19521, N19514);
buf BUF1 (N19522, N19493);
nor NOR2 (N19523, N19506, N1302);
or OR2 (N19524, N19509, N2893);
nor NOR3 (N19525, N19523, N3550, N16177);
nor NOR4 (N19526, N19524, N19354, N18401, N14142);
and AND3 (N19527, N19497, N13086, N2444);
or OR3 (N19528, N19519, N6335, N11230);
xor XOR2 (N19529, N19528, N11825);
not NOT1 (N19530, N19510);
nor NOR3 (N19531, N19527, N17341, N17841);
xor XOR2 (N19532, N19525, N3977);
and AND2 (N19533, N19531, N11470);
nor NOR3 (N19534, N19532, N1195, N352);
or OR2 (N19535, N19534, N5221);
not NOT1 (N19536, N19520);
nor NOR2 (N19537, N19530, N5643);
buf BUF1 (N19538, N19521);
nand NAND2 (N19539, N19522, N3560);
not NOT1 (N19540, N19533);
and AND2 (N19541, N19538, N8272);
or OR4 (N19542, N19529, N6652, N5440, N4595);
buf BUF1 (N19543, N19536);
or OR3 (N19544, N19516, N9998, N13154);
buf BUF1 (N19545, N19542);
buf BUF1 (N19546, N19526);
nor NOR2 (N19547, N19540, N10054);
or OR3 (N19548, N19544, N7029, N11860);
and AND2 (N19549, N19545, N10701);
or OR4 (N19550, N19547, N14178, N14031, N16250);
nor NOR2 (N19551, N19508, N19439);
nor NOR4 (N19552, N19543, N3835, N3594, N5696);
nand NAND2 (N19553, N19541, N6260);
nor NOR3 (N19554, N19553, N7854, N5898);
xor XOR2 (N19555, N19535, N2305);
xor XOR2 (N19556, N19550, N14418);
nor NOR3 (N19557, N19549, N11436, N7954);
xor XOR2 (N19558, N19537, N18514);
not NOT1 (N19559, N19548);
buf BUF1 (N19560, N19551);
nor NOR4 (N19561, N19546, N6830, N7483, N4062);
nand NAND4 (N19562, N19539, N8977, N8481, N6055);
nor NOR4 (N19563, N19559, N3257, N1503, N5790);
buf BUF1 (N19564, N19560);
and AND2 (N19565, N19557, N13943);
or OR2 (N19566, N19556, N11278);
not NOT1 (N19567, N19563);
not NOT1 (N19568, N19562);
xor XOR2 (N19569, N19555, N12338);
nand NAND4 (N19570, N19567, N18277, N19142, N8086);
or OR4 (N19571, N19566, N1515, N7171, N6381);
nor NOR4 (N19572, N19569, N8258, N11245, N18696);
nand NAND2 (N19573, N19558, N4600);
or OR4 (N19574, N19572, N8268, N3594, N15078);
or OR3 (N19575, N19565, N14561, N1754);
buf BUF1 (N19576, N19571);
not NOT1 (N19577, N19574);
and AND3 (N19578, N19576, N267, N11368);
buf BUF1 (N19579, N19554);
nand NAND4 (N19580, N19578, N8199, N17053, N7627);
buf BUF1 (N19581, N19561);
xor XOR2 (N19582, N19575, N17305);
nor NOR4 (N19583, N19564, N19133, N14630, N1923);
buf BUF1 (N19584, N19582);
xor XOR2 (N19585, N19552, N7142);
buf BUF1 (N19586, N19568);
and AND4 (N19587, N19577, N15763, N9624, N7194);
and AND4 (N19588, N19583, N17796, N12350, N15381);
nand NAND4 (N19589, N19585, N16427, N14943, N7883);
nor NOR4 (N19590, N19581, N19258, N2828, N13364);
xor XOR2 (N19591, N19580, N12657);
or OR3 (N19592, N19588, N1254, N4718);
nor NOR2 (N19593, N19589, N12616);
and AND2 (N19594, N19586, N2213);
buf BUF1 (N19595, N19587);
or OR2 (N19596, N19595, N17172);
or OR3 (N19597, N19594, N15630, N13542);
buf BUF1 (N19598, N19584);
or OR3 (N19599, N19592, N52, N5044);
buf BUF1 (N19600, N19579);
buf BUF1 (N19601, N19599);
nand NAND4 (N19602, N19591, N519, N14976, N8959);
nand NAND4 (N19603, N19570, N14458, N5070, N3895);
nand NAND3 (N19604, N19593, N15264, N2153);
nand NAND3 (N19605, N19604, N8481, N15541);
not NOT1 (N19606, N19603);
buf BUF1 (N19607, N19597);
and AND3 (N19608, N19602, N10894, N9123);
not NOT1 (N19609, N19596);
and AND3 (N19610, N19590, N4129, N12137);
nor NOR3 (N19611, N19607, N5133, N2735);
nand NAND4 (N19612, N19600, N14719, N17441, N15366);
or OR4 (N19613, N19612, N2294, N9241, N11563);
xor XOR2 (N19614, N19605, N4715);
not NOT1 (N19615, N19601);
xor XOR2 (N19616, N19610, N8054);
and AND3 (N19617, N19609, N12781, N17668);
buf BUF1 (N19618, N19573);
and AND3 (N19619, N19611, N10631, N18042);
xor XOR2 (N19620, N19618, N11067);
xor XOR2 (N19621, N19617, N18578);
and AND3 (N19622, N19608, N14681, N224);
and AND3 (N19623, N19621, N6495, N6740);
xor XOR2 (N19624, N19606, N3322);
nor NOR4 (N19625, N19613, N8308, N17085, N7494);
or OR4 (N19626, N19622, N166, N16821, N8410);
or OR3 (N19627, N19620, N3200, N13602);
nor NOR3 (N19628, N19616, N19431, N12824);
buf BUF1 (N19629, N19624);
nor NOR3 (N19630, N19598, N11169, N8637);
nand NAND4 (N19631, N19628, N15211, N10985, N12658);
or OR3 (N19632, N19615, N14117, N6603);
not NOT1 (N19633, N19619);
or OR3 (N19634, N19627, N1132, N14524);
nand NAND3 (N19635, N19633, N8008, N12340);
buf BUF1 (N19636, N19629);
nand NAND3 (N19637, N19614, N15496, N14138);
not NOT1 (N19638, N19625);
and AND3 (N19639, N19632, N9572, N9370);
not NOT1 (N19640, N19623);
nand NAND3 (N19641, N19636, N3730, N3668);
nand NAND4 (N19642, N19631, N867, N101, N6859);
nand NAND2 (N19643, N19626, N3227);
buf BUF1 (N19644, N19634);
or OR3 (N19645, N19644, N18338, N14453);
buf BUF1 (N19646, N19643);
not NOT1 (N19647, N19630);
xor XOR2 (N19648, N19646, N2207);
xor XOR2 (N19649, N19648, N8745);
and AND3 (N19650, N19649, N14446, N18299);
or OR2 (N19651, N19647, N7192);
nand NAND4 (N19652, N19638, N11430, N12991, N2255);
nand NAND2 (N19653, N19635, N7549);
or OR4 (N19654, N19652, N4507, N8394, N4583);
or OR4 (N19655, N19651, N10393, N14212, N11126);
or OR3 (N19656, N19653, N680, N7779);
nor NOR4 (N19657, N19640, N8867, N2956, N7693);
not NOT1 (N19658, N19650);
nand NAND4 (N19659, N19656, N13104, N794, N14501);
nor NOR4 (N19660, N19639, N9612, N3717, N10634);
xor XOR2 (N19661, N19637, N14271);
buf BUF1 (N19662, N19655);
not NOT1 (N19663, N19654);
xor XOR2 (N19664, N19659, N5680);
buf BUF1 (N19665, N19664);
buf BUF1 (N19666, N19661);
not NOT1 (N19667, N19641);
xor XOR2 (N19668, N19662, N16921);
nor NOR2 (N19669, N19665, N1695);
nand NAND4 (N19670, N19666, N11865, N14854, N12227);
or OR2 (N19671, N19657, N19183);
and AND3 (N19672, N19645, N19337, N140);
nand NAND4 (N19673, N19671, N12542, N7808, N11221);
or OR2 (N19674, N19672, N19501);
nor NOR4 (N19675, N19658, N8418, N10944, N14942);
nor NOR3 (N19676, N19670, N10319, N10472);
nand NAND4 (N19677, N19667, N9773, N1490, N16519);
not NOT1 (N19678, N19669);
or OR3 (N19679, N19677, N17835, N9062);
nand NAND3 (N19680, N19676, N18591, N8727);
buf BUF1 (N19681, N19674);
and AND4 (N19682, N19681, N3519, N13778, N5521);
nand NAND2 (N19683, N19678, N2305);
xor XOR2 (N19684, N19663, N18325);
or OR2 (N19685, N19642, N3802);
nand NAND4 (N19686, N19668, N12164, N6676, N6890);
nor NOR3 (N19687, N19683, N3667, N5426);
nor NOR3 (N19688, N19684, N15535, N456);
or OR2 (N19689, N19687, N6151);
not NOT1 (N19690, N19682);
not NOT1 (N19691, N19675);
or OR2 (N19692, N19679, N16734);
buf BUF1 (N19693, N19680);
buf BUF1 (N19694, N19660);
not NOT1 (N19695, N19694);
nand NAND3 (N19696, N19685, N1501, N2973);
and AND3 (N19697, N19692, N8611, N1900);
not NOT1 (N19698, N19688);
or OR4 (N19699, N19690, N17267, N3920, N5070);
nand NAND4 (N19700, N19698, N18477, N4284, N4588);
xor XOR2 (N19701, N19673, N3413);
buf BUF1 (N19702, N19701);
nand NAND2 (N19703, N19689, N15227);
and AND4 (N19704, N19699, N7864, N10119, N1949);
or OR2 (N19705, N19691, N10193);
nand NAND4 (N19706, N19700, N3238, N9904, N3551);
and AND3 (N19707, N19695, N6726, N6731);
nand NAND3 (N19708, N19706, N9671, N8111);
and AND4 (N19709, N19686, N18217, N11710, N2141);
xor XOR2 (N19710, N19703, N11644);
xor XOR2 (N19711, N19702, N15543);
nand NAND2 (N19712, N19707, N4178);
not NOT1 (N19713, N19710);
or OR4 (N19714, N19693, N12472, N12648, N12767);
or OR2 (N19715, N19714, N17733);
buf BUF1 (N19716, N19713);
and AND3 (N19717, N19704, N13763, N11435);
nand NAND3 (N19718, N19717, N4445, N19331);
not NOT1 (N19719, N19712);
and AND4 (N19720, N19719, N198, N1944, N5698);
nor NOR2 (N19721, N19705, N806);
nand NAND2 (N19722, N19697, N11998);
and AND2 (N19723, N19708, N15838);
buf BUF1 (N19724, N19709);
xor XOR2 (N19725, N19718, N9738);
xor XOR2 (N19726, N19725, N5481);
nor NOR2 (N19727, N19715, N18898);
or OR2 (N19728, N19696, N15428);
xor XOR2 (N19729, N19723, N1129);
buf BUF1 (N19730, N19721);
xor XOR2 (N19731, N19711, N3877);
not NOT1 (N19732, N19729);
nor NOR3 (N19733, N19720, N17353, N4045);
and AND3 (N19734, N19726, N15479, N16000);
nor NOR4 (N19735, N19728, N3202, N1194, N15119);
and AND3 (N19736, N19731, N9277, N6293);
and AND3 (N19737, N19735, N2522, N392);
buf BUF1 (N19738, N19733);
xor XOR2 (N19739, N19724, N3914);
and AND2 (N19740, N19732, N17376);
or OR2 (N19741, N19736, N3800);
xor XOR2 (N19742, N19739, N18377);
buf BUF1 (N19743, N19740);
buf BUF1 (N19744, N19730);
xor XOR2 (N19745, N19727, N11790);
not NOT1 (N19746, N19743);
not NOT1 (N19747, N19744);
buf BUF1 (N19748, N19734);
or OR2 (N19749, N19722, N5258);
and AND4 (N19750, N19749, N7846, N12562, N9652);
buf BUF1 (N19751, N19747);
not NOT1 (N19752, N19737);
xor XOR2 (N19753, N19746, N14720);
xor XOR2 (N19754, N19750, N7768);
xor XOR2 (N19755, N19745, N10454);
buf BUF1 (N19756, N19738);
nor NOR2 (N19757, N19741, N3795);
nor NOR3 (N19758, N19752, N8322, N18384);
xor XOR2 (N19759, N19756, N12571);
nor NOR4 (N19760, N19758, N3045, N4013, N15425);
nor NOR3 (N19761, N19742, N8523, N325);
nor NOR3 (N19762, N19716, N5561, N3962);
xor XOR2 (N19763, N19760, N12703);
nor NOR3 (N19764, N19761, N6106, N5158);
and AND3 (N19765, N19755, N6267, N3753);
and AND4 (N19766, N19757, N18873, N9190, N3796);
buf BUF1 (N19767, N19754);
or OR3 (N19768, N19764, N1888, N5516);
buf BUF1 (N19769, N19765);
not NOT1 (N19770, N19751);
and AND3 (N19771, N19768, N953, N11488);
nor NOR2 (N19772, N19770, N3012);
buf BUF1 (N19773, N19771);
nor NOR3 (N19774, N19759, N11216, N8186);
or OR2 (N19775, N19762, N19216);
and AND4 (N19776, N19767, N2303, N13583, N13870);
buf BUF1 (N19777, N19769);
or OR4 (N19778, N19775, N16358, N353, N2797);
xor XOR2 (N19779, N19778, N3157);
nand NAND4 (N19780, N19763, N7484, N7581, N4250);
nor NOR2 (N19781, N19772, N2826);
nor NOR3 (N19782, N19748, N13358, N6933);
buf BUF1 (N19783, N19773);
or OR2 (N19784, N19781, N13670);
nand NAND4 (N19785, N19783, N19150, N8784, N4433);
or OR3 (N19786, N19774, N7356, N12724);
nor NOR2 (N19787, N19777, N15952);
and AND4 (N19788, N19779, N8471, N135, N8671);
not NOT1 (N19789, N19786);
nand NAND3 (N19790, N19753, N9388, N14211);
nor NOR3 (N19791, N19790, N6941, N17369);
xor XOR2 (N19792, N19766, N4606);
not NOT1 (N19793, N19780);
xor XOR2 (N19794, N19788, N757);
or OR4 (N19795, N19776, N13675, N973, N4615);
buf BUF1 (N19796, N19795);
nand NAND4 (N19797, N19785, N14171, N5059, N26);
and AND3 (N19798, N19789, N12159, N15703);
buf BUF1 (N19799, N19791);
nor NOR2 (N19800, N19793, N948);
xor XOR2 (N19801, N19794, N8517);
and AND2 (N19802, N19800, N6925);
and AND4 (N19803, N19802, N3158, N17713, N2145);
or OR2 (N19804, N19796, N1564);
buf BUF1 (N19805, N19787);
nor NOR4 (N19806, N19782, N10193, N4216, N10892);
nor NOR2 (N19807, N19799, N13415);
nor NOR4 (N19808, N19804, N13438, N13287, N9793);
not NOT1 (N19809, N19805);
and AND4 (N19810, N19809, N17050, N8011, N2291);
and AND3 (N19811, N19792, N4001, N11644);
nor NOR3 (N19812, N19810, N13083, N19056);
nor NOR2 (N19813, N19801, N18958);
nor NOR4 (N19814, N19813, N7517, N1611, N6118);
xor XOR2 (N19815, N19803, N7941);
or OR3 (N19816, N19808, N17419, N11586);
and AND3 (N19817, N19784, N11099, N1245);
not NOT1 (N19818, N19806);
or OR3 (N19819, N19807, N14155, N14004);
or OR2 (N19820, N19818, N1562);
xor XOR2 (N19821, N19798, N16499);
xor XOR2 (N19822, N19814, N3741);
and AND2 (N19823, N19820, N18417);
and AND4 (N19824, N19817, N16154, N8945, N14897);
nor NOR2 (N19825, N19816, N3608);
not NOT1 (N19826, N19819);
and AND3 (N19827, N19797, N3912, N5283);
and AND4 (N19828, N19827, N18051, N18827, N4202);
xor XOR2 (N19829, N19812, N333);
or OR3 (N19830, N19829, N5292, N18910);
nor NOR4 (N19831, N19828, N9853, N16437, N1690);
xor XOR2 (N19832, N19821, N6290);
and AND3 (N19833, N19822, N12267, N9790);
nor NOR3 (N19834, N19831, N3769, N8510);
or OR3 (N19835, N19824, N3132, N5876);
xor XOR2 (N19836, N19823, N17859);
or OR4 (N19837, N19834, N3624, N16743, N11503);
nor NOR2 (N19838, N19815, N3925);
or OR3 (N19839, N19832, N1548, N6256);
buf BUF1 (N19840, N19837);
nor NOR4 (N19841, N19836, N4925, N2753, N10523);
nand NAND4 (N19842, N19826, N14059, N16733, N17255);
not NOT1 (N19843, N19835);
xor XOR2 (N19844, N19842, N2103);
nand NAND2 (N19845, N19844, N10569);
nor NOR4 (N19846, N19838, N7928, N13564, N3097);
and AND4 (N19847, N19839, N15048, N5, N3357);
nor NOR3 (N19848, N19811, N4715, N786);
and AND4 (N19849, N19845, N12310, N4551, N12927);
xor XOR2 (N19850, N19840, N3449);
buf BUF1 (N19851, N19833);
or OR3 (N19852, N19849, N7409, N14038);
xor XOR2 (N19853, N19847, N11010);
nor NOR2 (N19854, N19850, N18085);
nand NAND3 (N19855, N19830, N16209, N12876);
xor XOR2 (N19856, N19855, N15616);
nand NAND2 (N19857, N19848, N4958);
not NOT1 (N19858, N19825);
nand NAND4 (N19859, N19857, N65, N9794, N10902);
buf BUF1 (N19860, N19851);
and AND4 (N19861, N19846, N14219, N13470, N4930);
xor XOR2 (N19862, N19853, N7841);
nor NOR4 (N19863, N19841, N4222, N3408, N7937);
not NOT1 (N19864, N19860);
not NOT1 (N19865, N19862);
or OR4 (N19866, N19859, N12182, N17516, N16102);
nor NOR3 (N19867, N19865, N14152, N12630);
xor XOR2 (N19868, N19854, N6078);
nor NOR3 (N19869, N19863, N12320, N42);
not NOT1 (N19870, N19856);
nor NOR3 (N19871, N19866, N13684, N7771);
xor XOR2 (N19872, N19867, N2369);
buf BUF1 (N19873, N19868);
not NOT1 (N19874, N19870);
buf BUF1 (N19875, N19873);
or OR4 (N19876, N19861, N5301, N11544, N551);
nand NAND4 (N19877, N19852, N17610, N8698, N18065);
and AND2 (N19878, N19872, N849);
xor XOR2 (N19879, N19871, N7582);
nor NOR3 (N19880, N19864, N13284, N19217);
or OR4 (N19881, N19858, N5007, N11461, N15542);
nand NAND3 (N19882, N19874, N12547, N3731);
not NOT1 (N19883, N19875);
xor XOR2 (N19884, N19843, N1072);
or OR3 (N19885, N19883, N5415, N13663);
and AND2 (N19886, N19869, N413);
xor XOR2 (N19887, N19878, N9726);
not NOT1 (N19888, N19882);
or OR3 (N19889, N19880, N3842, N11979);
buf BUF1 (N19890, N19876);
and AND3 (N19891, N19890, N11187, N5237);
buf BUF1 (N19892, N19881);
and AND3 (N19893, N19887, N4354, N3039);
nand NAND2 (N19894, N19889, N627);
buf BUF1 (N19895, N19893);
and AND2 (N19896, N19877, N12898);
not NOT1 (N19897, N19884);
or OR3 (N19898, N19897, N7156, N8540);
and AND2 (N19899, N19891, N15583);
nor NOR4 (N19900, N19894, N15534, N7444, N19124);
xor XOR2 (N19901, N19879, N17243);
or OR3 (N19902, N19892, N8479, N6423);
or OR2 (N19903, N19898, N14469);
not NOT1 (N19904, N19885);
buf BUF1 (N19905, N19903);
or OR4 (N19906, N19896, N15990, N17930, N19744);
xor XOR2 (N19907, N19888, N8375);
nor NOR4 (N19908, N19902, N13276, N2366, N12343);
not NOT1 (N19909, N19901);
nor NOR2 (N19910, N19904, N13541);
buf BUF1 (N19911, N19909);
buf BUF1 (N19912, N19905);
not NOT1 (N19913, N19911);
not NOT1 (N19914, N19907);
nor NOR4 (N19915, N19910, N5733, N6383, N6525);
buf BUF1 (N19916, N19886);
or OR3 (N19917, N19915, N19854, N16416);
nor NOR4 (N19918, N19895, N17135, N17719, N15608);
buf BUF1 (N19919, N19916);
not NOT1 (N19920, N19919);
not NOT1 (N19921, N19913);
buf BUF1 (N19922, N19900);
not NOT1 (N19923, N19906);
and AND4 (N19924, N19922, N479, N5287, N14713);
xor XOR2 (N19925, N19914, N12835);
not NOT1 (N19926, N19923);
and AND2 (N19927, N19917, N7753);
buf BUF1 (N19928, N19925);
not NOT1 (N19929, N19920);
and AND3 (N19930, N19928, N17898, N8465);
and AND2 (N19931, N19924, N18136);
nor NOR3 (N19932, N19912, N14284, N2107);
not NOT1 (N19933, N19921);
and AND4 (N19934, N19927, N767, N9993, N1459);
nand NAND3 (N19935, N19908, N18853, N19149);
buf BUF1 (N19936, N19933);
and AND3 (N19937, N19932, N6250, N5012);
nand NAND3 (N19938, N19931, N15820, N9949);
nand NAND3 (N19939, N19938, N1905, N12170);
not NOT1 (N19940, N19934);
xor XOR2 (N19941, N19935, N17031);
nor NOR2 (N19942, N19899, N13157);
xor XOR2 (N19943, N19918, N15646);
and AND3 (N19944, N19941, N19698, N12911);
nor NOR2 (N19945, N19929, N6996);
buf BUF1 (N19946, N19936);
xor XOR2 (N19947, N19926, N12699);
not NOT1 (N19948, N19944);
buf BUF1 (N19949, N19937);
xor XOR2 (N19950, N19943, N10254);
buf BUF1 (N19951, N19930);
nor NOR3 (N19952, N19950, N16552, N11997);
nor NOR2 (N19953, N19947, N10194);
and AND3 (N19954, N19952, N1499, N15189);
nand NAND4 (N19955, N19939, N17438, N410, N10789);
not NOT1 (N19956, N19948);
xor XOR2 (N19957, N19945, N19438);
xor XOR2 (N19958, N19942, N11575);
nor NOR3 (N19959, N19949, N860, N9865);
nor NOR3 (N19960, N19953, N5334, N17748);
nand NAND4 (N19961, N19958, N14163, N251, N8002);
xor XOR2 (N19962, N19940, N7327);
nand NAND2 (N19963, N19957, N5196);
and AND4 (N19964, N19961, N19694, N14310, N10848);
nand NAND4 (N19965, N19946, N18146, N14899, N4631);
not NOT1 (N19966, N19956);
buf BUF1 (N19967, N19959);
buf BUF1 (N19968, N19964);
nand NAND3 (N19969, N19955, N11902, N16587);
and AND4 (N19970, N19951, N15811, N13512, N14789);
buf BUF1 (N19971, N19969);
nand NAND3 (N19972, N19963, N9161, N3210);
and AND3 (N19973, N19962, N17821, N15071);
buf BUF1 (N19974, N19971);
nand NAND3 (N19975, N19966, N19104, N10908);
nand NAND3 (N19976, N19975, N11115, N18124);
or OR4 (N19977, N19965, N1093, N5864, N5715);
and AND2 (N19978, N19970, N6570);
buf BUF1 (N19979, N19960);
nand NAND3 (N19980, N19972, N17016, N4325);
and AND4 (N19981, N19976, N979, N19357, N13524);
not NOT1 (N19982, N19954);
or OR4 (N19983, N19978, N15440, N10032, N12568);
nor NOR3 (N19984, N19967, N12455, N5228);
nor NOR2 (N19985, N19979, N9752);
nor NOR2 (N19986, N19984, N953);
and AND3 (N19987, N19982, N14361, N17879);
or OR2 (N19988, N19986, N8343);
nand NAND3 (N19989, N19968, N7183, N3316);
and AND3 (N19990, N19977, N16789, N510);
xor XOR2 (N19991, N19973, N67);
nand NAND2 (N19992, N19980, N14017);
or OR2 (N19993, N19983, N9246);
buf BUF1 (N19994, N19988);
not NOT1 (N19995, N19990);
and AND2 (N19996, N19974, N18439);
buf BUF1 (N19997, N19992);
xor XOR2 (N19998, N19987, N6682);
or OR2 (N19999, N19985, N16987);
nor NOR4 (N20000, N19994, N492, N7407, N17397);
or OR4 (N20001, N19998, N17086, N3355, N11130);
nand NAND3 (N20002, N19993, N6112, N12964);
and AND2 (N20003, N20000, N12756);
or OR3 (N20004, N19995, N11462, N9812);
nand NAND3 (N20005, N19989, N9330, N11235);
buf BUF1 (N20006, N19997);
or OR3 (N20007, N20003, N19841, N1692);
or OR2 (N20008, N19991, N9799);
xor XOR2 (N20009, N20007, N4173);
nand NAND3 (N20010, N20005, N14419, N5012);
and AND4 (N20011, N20006, N8881, N3650, N11894);
nor NOR2 (N20012, N20011, N13962);
xor XOR2 (N20013, N20010, N6004);
or OR4 (N20014, N20009, N18662, N17174, N9781);
nor NOR3 (N20015, N19996, N19544, N18593);
nand NAND4 (N20016, N20014, N1375, N19842, N6278);
nand NAND4 (N20017, N20016, N9775, N326, N18460);
not NOT1 (N20018, N20015);
or OR3 (N20019, N19981, N2870, N10006);
nor NOR4 (N20020, N20013, N7952, N348, N18393);
nor NOR4 (N20021, N20017, N3271, N16519, N3166);
not NOT1 (N20022, N20021);
buf BUF1 (N20023, N20012);
nor NOR3 (N20024, N20002, N11822, N3027);
not NOT1 (N20025, N20004);
nand NAND2 (N20026, N20019, N2412);
nand NAND4 (N20027, N20022, N6959, N15333, N14308);
or OR3 (N20028, N20023, N19167, N13003);
or OR2 (N20029, N20020, N5587);
and AND4 (N20030, N20029, N19125, N14424, N5290);
nor NOR2 (N20031, N20024, N745);
xor XOR2 (N20032, N20025, N1100);
nor NOR3 (N20033, N20030, N7835, N15711);
and AND2 (N20034, N20033, N2834);
xor XOR2 (N20035, N20026, N997);
nand NAND4 (N20036, N20034, N9320, N17424, N5596);
nand NAND2 (N20037, N19999, N14387);
and AND3 (N20038, N20037, N5219, N7207);
and AND3 (N20039, N20038, N14692, N583);
xor XOR2 (N20040, N20035, N9440);
nor NOR4 (N20041, N20008, N14537, N13497, N12710);
or OR3 (N20042, N20001, N3576, N7010);
buf BUF1 (N20043, N20018);
nand NAND2 (N20044, N20032, N10636);
nor NOR4 (N20045, N20036, N11114, N6230, N15357);
or OR4 (N20046, N20043, N17154, N19272, N16106);
nand NAND2 (N20047, N20046, N3712);
buf BUF1 (N20048, N20027);
nand NAND2 (N20049, N20031, N5857);
not NOT1 (N20050, N20042);
or OR2 (N20051, N20050, N10390);
xor XOR2 (N20052, N20045, N19032);
xor XOR2 (N20053, N20028, N925);
xor XOR2 (N20054, N20052, N9602);
and AND2 (N20055, N20054, N8415);
buf BUF1 (N20056, N20047);
nand NAND4 (N20057, N20040, N14400, N8643, N11249);
buf BUF1 (N20058, N20053);
xor XOR2 (N20059, N20057, N171);
xor XOR2 (N20060, N20056, N12531);
and AND2 (N20061, N20041, N11806);
nand NAND4 (N20062, N20058, N7548, N16822, N17559);
buf BUF1 (N20063, N20051);
and AND2 (N20064, N20060, N4022);
nand NAND2 (N20065, N20055, N13901);
nand NAND3 (N20066, N20048, N8787, N16800);
nor NOR2 (N20067, N20049, N9814);
xor XOR2 (N20068, N20063, N13332);
or OR3 (N20069, N20061, N18765, N8010);
xor XOR2 (N20070, N20062, N8104);
nand NAND2 (N20071, N20044, N6409);
or OR2 (N20072, N20064, N5957);
and AND4 (N20073, N20039, N17111, N9580, N14970);
buf BUF1 (N20074, N20066);
or OR3 (N20075, N20074, N2173, N3979);
and AND2 (N20076, N20068, N18227);
nor NOR3 (N20077, N20075, N17785, N14722);
nand NAND4 (N20078, N20069, N287, N11623, N15572);
nor NOR4 (N20079, N20072, N12631, N16321, N9667);
xor XOR2 (N20080, N20067, N3584);
or OR2 (N20081, N20065, N17454);
buf BUF1 (N20082, N20079);
and AND4 (N20083, N20078, N8206, N17513, N4215);
not NOT1 (N20084, N20071);
nor NOR2 (N20085, N20083, N3820);
not NOT1 (N20086, N20082);
nand NAND2 (N20087, N20085, N15519);
or OR3 (N20088, N20077, N5489, N17112);
xor XOR2 (N20089, N20084, N4653);
and AND4 (N20090, N20086, N14382, N3349, N8318);
buf BUF1 (N20091, N20076);
and AND4 (N20092, N20091, N10936, N7207, N8578);
and AND3 (N20093, N20059, N11248, N4342);
xor XOR2 (N20094, N20088, N18632);
nand NAND4 (N20095, N20093, N12281, N12641, N8445);
nand NAND4 (N20096, N20092, N18706, N6689, N7340);
nor NOR2 (N20097, N20073, N4803);
xor XOR2 (N20098, N20097, N7164);
not NOT1 (N20099, N20080);
and AND3 (N20100, N20070, N15126, N10602);
or OR2 (N20101, N20099, N4559);
nand NAND4 (N20102, N20095, N9357, N8832, N17110);
nor NOR2 (N20103, N20089, N12644);
buf BUF1 (N20104, N20094);
or OR4 (N20105, N20103, N3471, N499, N7788);
not NOT1 (N20106, N20104);
or OR4 (N20107, N20098, N12767, N10300, N1185);
nor NOR4 (N20108, N20096, N7697, N6065, N3885);
nand NAND3 (N20109, N20107, N8142, N11440);
xor XOR2 (N20110, N20108, N16028);
nor NOR4 (N20111, N20090, N11515, N14000, N9447);
buf BUF1 (N20112, N20111);
xor XOR2 (N20113, N20106, N18618);
nor NOR4 (N20114, N20101, N6969, N19415, N10224);
xor XOR2 (N20115, N20087, N8883);
and AND2 (N20116, N20102, N3653);
xor XOR2 (N20117, N20105, N12991);
nand NAND3 (N20118, N20110, N16862, N964);
or OR2 (N20119, N20081, N7985);
xor XOR2 (N20120, N20116, N10346);
and AND4 (N20121, N20120, N3653, N8314, N15579);
nand NAND4 (N20122, N20112, N15485, N18374, N13454);
and AND2 (N20123, N20115, N12809);
nand NAND3 (N20124, N20121, N9834, N4632);
and AND4 (N20125, N20109, N14626, N3121, N211);
or OR3 (N20126, N20117, N10847, N18969);
nand NAND3 (N20127, N20113, N19709, N7711);
not NOT1 (N20128, N20123);
and AND2 (N20129, N20127, N16795);
nand NAND3 (N20130, N20100, N8529, N8516);
nand NAND4 (N20131, N20130, N18509, N18055, N9625);
nor NOR2 (N20132, N20114, N11435);
buf BUF1 (N20133, N20125);
buf BUF1 (N20134, N20118);
and AND4 (N20135, N20129, N7463, N11362, N4126);
or OR3 (N20136, N20132, N12449, N6171);
nor NOR4 (N20137, N20131, N17275, N1597, N6073);
nand NAND2 (N20138, N20126, N16462);
nand NAND3 (N20139, N20119, N11550, N18545);
nor NOR3 (N20140, N20136, N7936, N1853);
xor XOR2 (N20141, N20139, N19137);
nand NAND3 (N20142, N20135, N8213, N7377);
nor NOR2 (N20143, N20124, N20140);
buf BUF1 (N20144, N12375);
buf BUF1 (N20145, N20141);
buf BUF1 (N20146, N20144);
xor XOR2 (N20147, N20145, N9016);
buf BUF1 (N20148, N20128);
not NOT1 (N20149, N20146);
nor NOR2 (N20150, N20149, N5186);
nor NOR3 (N20151, N20137, N7660, N4058);
not NOT1 (N20152, N20150);
buf BUF1 (N20153, N20122);
nor NOR3 (N20154, N20147, N8132, N5757);
and AND2 (N20155, N20152, N14526);
buf BUF1 (N20156, N20151);
and AND4 (N20157, N20138, N1971, N16741, N5590);
and AND3 (N20158, N20133, N9889, N7588);
xor XOR2 (N20159, N20158, N13233);
and AND3 (N20160, N20156, N10178, N13455);
nor NOR3 (N20161, N20157, N14674, N14956);
nor NOR2 (N20162, N20153, N4614);
or OR3 (N20163, N20161, N17701, N12870);
and AND3 (N20164, N20159, N6279, N449);
buf BUF1 (N20165, N20155);
and AND3 (N20166, N20160, N6229, N16641);
nor NOR2 (N20167, N20134, N2075);
nor NOR3 (N20168, N20167, N8772, N2730);
not NOT1 (N20169, N20165);
buf BUF1 (N20170, N20169);
nand NAND2 (N20171, N20154, N19153);
nor NOR4 (N20172, N20168, N4155, N1057, N14027);
nor NOR3 (N20173, N20142, N6845, N13791);
nor NOR3 (N20174, N20163, N10383, N16844);
xor XOR2 (N20175, N20143, N859);
or OR4 (N20176, N20166, N14602, N14446, N10082);
not NOT1 (N20177, N20170);
and AND2 (N20178, N20175, N18241);
and AND3 (N20179, N20162, N6730, N2173);
nor NOR4 (N20180, N20173, N2130, N589, N7523);
nor NOR3 (N20181, N20164, N9621, N5055);
not NOT1 (N20182, N20148);
nand NAND2 (N20183, N20178, N17401);
nand NAND4 (N20184, N20179, N1390, N17746, N10450);
nor NOR4 (N20185, N20184, N6287, N13974, N15333);
or OR2 (N20186, N20181, N11653);
not NOT1 (N20187, N20185);
buf BUF1 (N20188, N20182);
nand NAND4 (N20189, N20171, N9486, N969, N8944);
nand NAND4 (N20190, N20180, N3987, N11951, N15052);
or OR3 (N20191, N20188, N2962, N12789);
and AND4 (N20192, N20191, N18595, N17339, N16531);
nand NAND3 (N20193, N20176, N18913, N15007);
or OR3 (N20194, N20193, N8037, N6578);
not NOT1 (N20195, N20190);
nand NAND3 (N20196, N20195, N4556, N15356);
buf BUF1 (N20197, N20192);
or OR4 (N20198, N20174, N8241, N16523, N16239);
nand NAND3 (N20199, N20177, N7947, N630);
or OR3 (N20200, N20186, N11725, N4698);
xor XOR2 (N20201, N20200, N12071);
buf BUF1 (N20202, N20194);
nor NOR3 (N20203, N20172, N5083, N4158);
or OR3 (N20204, N20183, N18943, N5414);
nor NOR4 (N20205, N20189, N9822, N7750, N18423);
or OR3 (N20206, N20202, N6076, N17344);
nor NOR4 (N20207, N20203, N12953, N8902, N17552);
nor NOR2 (N20208, N20187, N3577);
nor NOR4 (N20209, N20196, N14024, N17698, N13242);
nor NOR3 (N20210, N20208, N12530, N10976);
nor NOR3 (N20211, N20206, N6607, N845);
or OR4 (N20212, N20198, N18907, N19032, N9913);
nor NOR2 (N20213, N20204, N2472);
xor XOR2 (N20214, N20212, N12407);
nand NAND3 (N20215, N20197, N3136, N11176);
or OR4 (N20216, N20205, N16772, N769, N4983);
nand NAND4 (N20217, N20216, N16085, N2733, N17661);
not NOT1 (N20218, N20209);
not NOT1 (N20219, N20217);
and AND3 (N20220, N20215, N18145, N6573);
xor XOR2 (N20221, N20220, N3755);
xor XOR2 (N20222, N20218, N12691);
xor XOR2 (N20223, N20210, N18467);
xor XOR2 (N20224, N20219, N1171);
not NOT1 (N20225, N20223);
buf BUF1 (N20226, N20222);
xor XOR2 (N20227, N20213, N7728);
not NOT1 (N20228, N20225);
nor NOR4 (N20229, N20214, N2560, N7338, N15527);
xor XOR2 (N20230, N20211, N850);
not NOT1 (N20231, N20229);
buf BUF1 (N20232, N20224);
nand NAND2 (N20233, N20227, N13027);
and AND2 (N20234, N20226, N8398);
xor XOR2 (N20235, N20228, N3708);
or OR2 (N20236, N20199, N747);
buf BUF1 (N20237, N20236);
not NOT1 (N20238, N20207);
nand NAND2 (N20239, N20234, N11564);
or OR3 (N20240, N20201, N10616, N1735);
buf BUF1 (N20241, N20237);
buf BUF1 (N20242, N20235);
not NOT1 (N20243, N20221);
not NOT1 (N20244, N20243);
nand NAND3 (N20245, N20239, N6209, N373);
buf BUF1 (N20246, N20245);
buf BUF1 (N20247, N20241);
xor XOR2 (N20248, N20238, N8762);
not NOT1 (N20249, N20244);
nor NOR4 (N20250, N20232, N15065, N18840, N10479);
or OR4 (N20251, N20248, N9653, N351, N1086);
and AND2 (N20252, N20249, N3988);
xor XOR2 (N20253, N20247, N9547);
not NOT1 (N20254, N20246);
or OR2 (N20255, N20250, N11142);
nor NOR3 (N20256, N20231, N8942, N11060);
or OR4 (N20257, N20252, N13905, N10352, N10558);
nand NAND2 (N20258, N20256, N1613);
not NOT1 (N20259, N20242);
not NOT1 (N20260, N20257);
or OR2 (N20261, N20230, N4665);
or OR3 (N20262, N20258, N6527, N12564);
and AND2 (N20263, N20253, N6897);
not NOT1 (N20264, N20255);
nand NAND4 (N20265, N20263, N10359, N12876, N2429);
or OR2 (N20266, N20264, N12922);
nor NOR2 (N20267, N20259, N792);
nand NAND4 (N20268, N20233, N921, N18717, N570);
nand NAND4 (N20269, N20240, N3798, N13664, N15724);
not NOT1 (N20270, N20268);
and AND4 (N20271, N20262, N13897, N6782, N5141);
nor NOR2 (N20272, N20261, N13760);
or OR4 (N20273, N20270, N4012, N7136, N18183);
not NOT1 (N20274, N20271);
nor NOR2 (N20275, N20251, N18690);
nor NOR2 (N20276, N20265, N10147);
nor NOR3 (N20277, N20269, N2526, N11551);
buf BUF1 (N20278, N20273);
or OR4 (N20279, N20277, N15735, N2649, N18306);
nand NAND3 (N20280, N20279, N6163, N20199);
nand NAND2 (N20281, N20266, N10898);
and AND3 (N20282, N20281, N15153, N6132);
buf BUF1 (N20283, N20254);
nor NOR3 (N20284, N20278, N15187, N2713);
buf BUF1 (N20285, N20280);
or OR4 (N20286, N20276, N10135, N20265, N12963);
not NOT1 (N20287, N20267);
and AND3 (N20288, N20260, N15216, N565);
or OR4 (N20289, N20283, N17261, N10340, N11888);
buf BUF1 (N20290, N20275);
buf BUF1 (N20291, N20285);
buf BUF1 (N20292, N20286);
or OR3 (N20293, N20282, N13310, N3450);
xor XOR2 (N20294, N20293, N9752);
nand NAND2 (N20295, N20294, N754);
xor XOR2 (N20296, N20284, N9053);
and AND3 (N20297, N20291, N211, N4151);
nand NAND4 (N20298, N20274, N11222, N18433, N7695);
nand NAND4 (N20299, N20287, N12318, N9512, N12469);
and AND4 (N20300, N20289, N19974, N20251, N10250);
nand NAND4 (N20301, N20292, N18287, N15696, N6982);
buf BUF1 (N20302, N20299);
or OR3 (N20303, N20288, N20141, N6243);
xor XOR2 (N20304, N20295, N6278);
and AND2 (N20305, N20290, N16311);
and AND4 (N20306, N20298, N17220, N2230, N9928);
nor NOR3 (N20307, N20302, N16083, N14747);
buf BUF1 (N20308, N20301);
not NOT1 (N20309, N20304);
nand NAND2 (N20310, N20303, N7340);
nor NOR2 (N20311, N20305, N2342);
nand NAND2 (N20312, N20309, N16542);
and AND3 (N20313, N20272, N12323, N8159);
nand NAND3 (N20314, N20300, N16303, N12151);
nand NAND2 (N20315, N20308, N8184);
not NOT1 (N20316, N20296);
xor XOR2 (N20317, N20313, N11805);
or OR4 (N20318, N20312, N18451, N9154, N4849);
buf BUF1 (N20319, N20297);
buf BUF1 (N20320, N20319);
not NOT1 (N20321, N20314);
and AND4 (N20322, N20315, N8663, N10380, N7770);
xor XOR2 (N20323, N20310, N7467);
not NOT1 (N20324, N20321);
or OR3 (N20325, N20322, N8552, N7041);
and AND2 (N20326, N20307, N19930);
or OR4 (N20327, N20326, N15948, N10935, N15920);
xor XOR2 (N20328, N20320, N6029);
nand NAND2 (N20329, N20317, N1112);
nand NAND2 (N20330, N20318, N18613);
or OR4 (N20331, N20325, N19785, N17041, N9491);
nor NOR4 (N20332, N20311, N19287, N11298, N11785);
not NOT1 (N20333, N20316);
nor NOR2 (N20334, N20323, N16899);
not NOT1 (N20335, N20329);
nand NAND3 (N20336, N20327, N10678, N4677);
nor NOR3 (N20337, N20330, N1655, N8101);
nand NAND2 (N20338, N20332, N5601);
nand NAND2 (N20339, N20333, N11094);
nand NAND2 (N20340, N20306, N6163);
buf BUF1 (N20341, N20337);
xor XOR2 (N20342, N20331, N8258);
xor XOR2 (N20343, N20336, N10726);
xor XOR2 (N20344, N20341, N9497);
buf BUF1 (N20345, N20344);
buf BUF1 (N20346, N20335);
nor NOR2 (N20347, N20339, N10863);
or OR2 (N20348, N20342, N18976);
or OR2 (N20349, N20338, N604);
nand NAND4 (N20350, N20346, N9643, N18559, N13529);
and AND2 (N20351, N20349, N3637);
xor XOR2 (N20352, N20345, N18287);
xor XOR2 (N20353, N20347, N13465);
xor XOR2 (N20354, N20352, N17041);
or OR2 (N20355, N20324, N11219);
buf BUF1 (N20356, N20334);
not NOT1 (N20357, N20356);
nand NAND4 (N20358, N20340, N13229, N18773, N14903);
buf BUF1 (N20359, N20353);
or OR2 (N20360, N20328, N2373);
nor NOR2 (N20361, N20359, N16276);
and AND3 (N20362, N20357, N9493, N12521);
not NOT1 (N20363, N20354);
or OR3 (N20364, N20358, N19033, N12594);
not NOT1 (N20365, N20355);
nor NOR2 (N20366, N20364, N11906);
and AND3 (N20367, N20362, N6794, N2406);
nand NAND3 (N20368, N20363, N5225, N2762);
buf BUF1 (N20369, N20365);
buf BUF1 (N20370, N20351);
nor NOR3 (N20371, N20350, N3686, N1747);
nor NOR4 (N20372, N20370, N8563, N10934, N14068);
not NOT1 (N20373, N20348);
nand NAND4 (N20374, N20343, N6385, N3657, N12067);
or OR4 (N20375, N20374, N9417, N5450, N12078);
and AND3 (N20376, N20361, N1237, N5157);
and AND3 (N20377, N20372, N6599, N2439);
nor NOR2 (N20378, N20366, N4571);
and AND2 (N20379, N20368, N8472);
not NOT1 (N20380, N20375);
or OR4 (N20381, N20373, N3006, N6148, N4143);
nand NAND3 (N20382, N20376, N2654, N18925);
and AND3 (N20383, N20381, N8230, N20247);
xor XOR2 (N20384, N20360, N5975);
xor XOR2 (N20385, N20384, N19797);
buf BUF1 (N20386, N20383);
buf BUF1 (N20387, N20386);
or OR4 (N20388, N20382, N18870, N10329, N5207);
or OR3 (N20389, N20380, N17123, N18699);
and AND3 (N20390, N20387, N14695, N10475);
and AND2 (N20391, N20377, N19702);
and AND2 (N20392, N20388, N7560);
buf BUF1 (N20393, N20391);
nor NOR3 (N20394, N20393, N992, N13066);
nand NAND3 (N20395, N20379, N2836, N1393);
buf BUF1 (N20396, N20369);
or OR3 (N20397, N20371, N10189, N5566);
and AND2 (N20398, N20394, N5731);
and AND4 (N20399, N20390, N6440, N4140, N3106);
nor NOR3 (N20400, N20397, N11542, N18377);
or OR4 (N20401, N20389, N11903, N14845, N3351);
not NOT1 (N20402, N20392);
or OR2 (N20403, N20401, N19184);
and AND3 (N20404, N20385, N5915, N19662);
and AND3 (N20405, N20395, N8625, N19809);
nor NOR2 (N20406, N20396, N13353);
and AND2 (N20407, N20378, N12007);
and AND2 (N20408, N20398, N14140);
and AND4 (N20409, N20403, N20161, N8207, N8329);
not NOT1 (N20410, N20407);
xor XOR2 (N20411, N20406, N5998);
buf BUF1 (N20412, N20409);
or OR3 (N20413, N20367, N8477, N19721);
xor XOR2 (N20414, N20413, N16554);
nor NOR2 (N20415, N20402, N7284);
nand NAND4 (N20416, N20411, N14310, N11134, N18118);
and AND3 (N20417, N20404, N18686, N17773);
nand NAND4 (N20418, N20415, N14952, N10357, N18342);
xor XOR2 (N20419, N20408, N8818);
buf BUF1 (N20420, N20419);
nand NAND3 (N20421, N20412, N17442, N11780);
or OR2 (N20422, N20421, N3538);
nor NOR2 (N20423, N20420, N4161);
nor NOR4 (N20424, N20417, N3391, N12881, N12832);
or OR2 (N20425, N20424, N1212);
nor NOR2 (N20426, N20422, N5655);
buf BUF1 (N20427, N20416);
nand NAND2 (N20428, N20405, N7485);
nand NAND3 (N20429, N20428, N7426, N1497);
buf BUF1 (N20430, N20399);
nand NAND2 (N20431, N20426, N17627);
and AND3 (N20432, N20400, N1755, N10741);
buf BUF1 (N20433, N20425);
nand NAND2 (N20434, N20423, N8676);
nor NOR3 (N20435, N20429, N15835, N20093);
not NOT1 (N20436, N20434);
not NOT1 (N20437, N20432);
buf BUF1 (N20438, N20436);
and AND3 (N20439, N20437, N18562, N18747);
nand NAND2 (N20440, N20438, N2326);
xor XOR2 (N20441, N20414, N14412);
not NOT1 (N20442, N20430);
xor XOR2 (N20443, N20441, N3346);
nand NAND3 (N20444, N20439, N811, N13889);
not NOT1 (N20445, N20435);
not NOT1 (N20446, N20410);
or OR2 (N20447, N20418, N6039);
or OR2 (N20448, N20433, N13347);
nand NAND4 (N20449, N20446, N19810, N14849, N8897);
not NOT1 (N20450, N20447);
nor NOR2 (N20451, N20450, N15941);
xor XOR2 (N20452, N20431, N10537);
nor NOR4 (N20453, N20452, N14431, N3832, N152);
nand NAND3 (N20454, N20448, N12738, N9060);
not NOT1 (N20455, N20453);
buf BUF1 (N20456, N20455);
buf BUF1 (N20457, N20427);
nand NAND3 (N20458, N20457, N16262, N18350);
xor XOR2 (N20459, N20445, N16950);
nor NOR2 (N20460, N20449, N17806);
buf BUF1 (N20461, N20442);
not NOT1 (N20462, N20454);
xor XOR2 (N20463, N20443, N15401);
nor NOR4 (N20464, N20462, N2485, N8708, N10940);
xor XOR2 (N20465, N20456, N3);
not NOT1 (N20466, N20444);
nor NOR4 (N20467, N20463, N2451, N12526, N4003);
buf BUF1 (N20468, N20466);
nand NAND4 (N20469, N20461, N6478, N7713, N7875);
buf BUF1 (N20470, N20458);
buf BUF1 (N20471, N20460);
not NOT1 (N20472, N20465);
buf BUF1 (N20473, N20469);
buf BUF1 (N20474, N20464);
not NOT1 (N20475, N20473);
nand NAND3 (N20476, N20467, N18193, N19333);
nor NOR3 (N20477, N20459, N17969, N2237);
or OR4 (N20478, N20476, N5262, N12902, N16024);
and AND2 (N20479, N20470, N6707);
not NOT1 (N20480, N20477);
buf BUF1 (N20481, N20475);
buf BUF1 (N20482, N20471);
buf BUF1 (N20483, N20440);
not NOT1 (N20484, N20479);
and AND2 (N20485, N20482, N18698);
or OR4 (N20486, N20451, N17976, N1798, N6237);
nand NAND2 (N20487, N20472, N12816);
or OR4 (N20488, N20480, N12582, N9201, N10673);
nor NOR4 (N20489, N20488, N281, N8067, N13754);
nor NOR4 (N20490, N20468, N1933, N17830, N12827);
nand NAND2 (N20491, N20487, N11862);
buf BUF1 (N20492, N20478);
nor NOR4 (N20493, N20491, N13825, N18845, N701);
not NOT1 (N20494, N20493);
or OR2 (N20495, N20494, N3253);
or OR4 (N20496, N20489, N1319, N19741, N12537);
buf BUF1 (N20497, N20492);
or OR2 (N20498, N20474, N317);
nor NOR2 (N20499, N20498, N8533);
nor NOR2 (N20500, N20495, N2445);
nor NOR4 (N20501, N20486, N19346, N14992, N18912);
nor NOR3 (N20502, N20484, N19624, N17665);
or OR3 (N20503, N20500, N6534, N8132);
nand NAND3 (N20504, N20503, N7132, N17784);
nand NAND3 (N20505, N20501, N17821, N12275);
or OR2 (N20506, N20481, N2966);
xor XOR2 (N20507, N20485, N5195);
buf BUF1 (N20508, N20505);
not NOT1 (N20509, N20496);
nor NOR4 (N20510, N20508, N11672, N16, N3028);
and AND2 (N20511, N20490, N7004);
nor NOR3 (N20512, N20511, N18556, N9993);
xor XOR2 (N20513, N20506, N9937);
not NOT1 (N20514, N20497);
not NOT1 (N20515, N20507);
nor NOR4 (N20516, N20483, N12442, N15572, N7745);
or OR3 (N20517, N20516, N13180, N17663);
or OR3 (N20518, N20513, N6057, N1769);
not NOT1 (N20519, N20512);
nand NAND4 (N20520, N20510, N17202, N20164, N10591);
nand NAND4 (N20521, N20504, N13852, N8228, N18078);
buf BUF1 (N20522, N20515);
and AND3 (N20523, N20519, N18531, N14694);
not NOT1 (N20524, N20499);
nor NOR2 (N20525, N20523, N13385);
buf BUF1 (N20526, N20514);
and AND4 (N20527, N20520, N3303, N11032, N16648);
nor NOR4 (N20528, N20525, N18619, N8747, N98);
nand NAND3 (N20529, N20509, N1282, N11528);
or OR4 (N20530, N20521, N15436, N13061, N12480);
buf BUF1 (N20531, N20517);
buf BUF1 (N20532, N20528);
or OR3 (N20533, N20524, N2658, N284);
or OR3 (N20534, N20532, N19337, N13328);
not NOT1 (N20535, N20527);
and AND2 (N20536, N20533, N13607);
or OR2 (N20537, N20535, N8894);
buf BUF1 (N20538, N20526);
and AND4 (N20539, N20531, N19437, N12968, N4169);
xor XOR2 (N20540, N20534, N17426);
not NOT1 (N20541, N20539);
nand NAND2 (N20542, N20537, N10999);
or OR2 (N20543, N20538, N4686);
nor NOR2 (N20544, N20518, N3538);
nor NOR4 (N20545, N20536, N9147, N6881, N19793);
nor NOR4 (N20546, N20530, N6796, N16580, N1318);
not NOT1 (N20547, N20546);
and AND2 (N20548, N20543, N13549);
or OR4 (N20549, N20547, N2078, N8551, N9971);
nor NOR2 (N20550, N20540, N17009);
not NOT1 (N20551, N20549);
nand NAND3 (N20552, N20551, N15546, N1304);
or OR4 (N20553, N20529, N274, N5800, N11469);
nand NAND3 (N20554, N20545, N912, N3556);
or OR4 (N20555, N20541, N7639, N13385, N15449);
or OR4 (N20556, N20522, N12465, N18035, N4959);
nand NAND3 (N20557, N20554, N5676, N13265);
or OR4 (N20558, N20557, N12020, N16174, N6134);
buf BUF1 (N20559, N20553);
or OR3 (N20560, N20556, N15858, N8880);
xor XOR2 (N20561, N20560, N15814);
buf BUF1 (N20562, N20559);
or OR3 (N20563, N20558, N1167, N8862);
nand NAND3 (N20564, N20544, N3400, N8427);
buf BUF1 (N20565, N20552);
nor NOR3 (N20566, N20542, N6258, N2440);
xor XOR2 (N20567, N20562, N9647);
or OR2 (N20568, N20565, N9145);
or OR3 (N20569, N20563, N7559, N10334);
and AND2 (N20570, N20567, N19227);
not NOT1 (N20571, N20548);
nor NOR4 (N20572, N20555, N4308, N3983, N16920);
nand NAND4 (N20573, N20572, N4864, N16552, N5604);
nand NAND3 (N20574, N20568, N4941, N18944);
not NOT1 (N20575, N20564);
or OR4 (N20576, N20569, N2199, N6730, N8222);
not NOT1 (N20577, N20550);
xor XOR2 (N20578, N20561, N8076);
not NOT1 (N20579, N20566);
nor NOR3 (N20580, N20576, N16918, N10002);
buf BUF1 (N20581, N20578);
xor XOR2 (N20582, N20570, N20048);
or OR4 (N20583, N20577, N19745, N901, N10156);
not NOT1 (N20584, N20579);
nand NAND2 (N20585, N20582, N17367);
nand NAND4 (N20586, N20574, N11879, N20118, N5232);
xor XOR2 (N20587, N20502, N12621);
xor XOR2 (N20588, N20573, N910);
xor XOR2 (N20589, N20575, N3135);
and AND2 (N20590, N20580, N5598);
xor XOR2 (N20591, N20584, N5073);
nand NAND4 (N20592, N20581, N15656, N14141, N18837);
and AND2 (N20593, N20586, N10888);
and AND2 (N20594, N20571, N16996);
nor NOR4 (N20595, N20589, N17738, N9346, N6622);
not NOT1 (N20596, N20588);
not NOT1 (N20597, N20590);
nor NOR4 (N20598, N20593, N11759, N9985, N10563);
nand NAND2 (N20599, N20591, N11225);
xor XOR2 (N20600, N20597, N13582);
nor NOR4 (N20601, N20585, N19561, N18772, N16057);
nor NOR4 (N20602, N20598, N8320, N10239, N16138);
xor XOR2 (N20603, N20600, N8838);
xor XOR2 (N20604, N20596, N18037);
not NOT1 (N20605, N20601);
nand NAND3 (N20606, N20604, N11568, N7847);
nor NOR4 (N20607, N20603, N15698, N2440, N11536);
not NOT1 (N20608, N20594);
or OR4 (N20609, N20592, N2814, N18738, N6675);
or OR4 (N20610, N20605, N12581, N12543, N1601);
buf BUF1 (N20611, N20610);
xor XOR2 (N20612, N20609, N16314);
xor XOR2 (N20613, N20612, N16422);
and AND3 (N20614, N20583, N5408, N13771);
nor NOR4 (N20615, N20587, N16877, N16366, N5576);
buf BUF1 (N20616, N20606);
not NOT1 (N20617, N20602);
nand NAND2 (N20618, N20616, N17628);
buf BUF1 (N20619, N20614);
buf BUF1 (N20620, N20615);
or OR3 (N20621, N20607, N13155, N18550);
nor NOR4 (N20622, N20611, N18922, N13253, N15814);
xor XOR2 (N20623, N20618, N17554);
and AND4 (N20624, N20599, N2094, N20477, N14307);
or OR4 (N20625, N20621, N18338, N5725, N13907);
or OR3 (N20626, N20595, N3556, N20013);
buf BUF1 (N20627, N20620);
nor NOR3 (N20628, N20608, N13612, N18440);
buf BUF1 (N20629, N20619);
or OR4 (N20630, N20622, N17317, N3082, N12728);
buf BUF1 (N20631, N20629);
xor XOR2 (N20632, N20626, N14719);
or OR2 (N20633, N20631, N6733);
nor NOR4 (N20634, N20632, N3972, N6273, N2531);
nand NAND2 (N20635, N20630, N17071);
and AND3 (N20636, N20635, N5910, N15225);
not NOT1 (N20637, N20623);
and AND3 (N20638, N20625, N11645, N16454);
not NOT1 (N20639, N20613);
or OR3 (N20640, N20636, N11363, N12566);
nand NAND4 (N20641, N20624, N13410, N11723, N2005);
nand NAND2 (N20642, N20633, N9710);
nand NAND4 (N20643, N20627, N10827, N9985, N2305);
not NOT1 (N20644, N20628);
and AND4 (N20645, N20643, N7008, N1754, N8865);
or OR3 (N20646, N20642, N11485, N3297);
buf BUF1 (N20647, N20646);
and AND3 (N20648, N20617, N8614, N20221);
and AND3 (N20649, N20639, N20519, N20592);
and AND3 (N20650, N20641, N19649, N12598);
nand NAND4 (N20651, N20634, N3901, N16377, N18420);
or OR4 (N20652, N20644, N6278, N1751, N5988);
and AND4 (N20653, N20640, N13490, N10981, N16784);
and AND3 (N20654, N20638, N8987, N16301);
buf BUF1 (N20655, N20645);
nor NOR4 (N20656, N20650, N15592, N4643, N7854);
not NOT1 (N20657, N20654);
or OR4 (N20658, N20657, N17824, N585, N1994);
and AND3 (N20659, N20647, N11789, N10669);
buf BUF1 (N20660, N20659);
and AND3 (N20661, N20653, N4893, N8759);
nand NAND3 (N20662, N20655, N8079, N19876);
not NOT1 (N20663, N20648);
and AND4 (N20664, N20652, N2811, N15465, N1203);
and AND3 (N20665, N20651, N10997, N4799);
and AND2 (N20666, N20661, N1086);
buf BUF1 (N20667, N20662);
not NOT1 (N20668, N20665);
not NOT1 (N20669, N20637);
nor NOR3 (N20670, N20667, N15778, N14333);
not NOT1 (N20671, N20670);
nor NOR2 (N20672, N20668, N17963);
not NOT1 (N20673, N20656);
buf BUF1 (N20674, N20658);
xor XOR2 (N20675, N20660, N5967);
buf BUF1 (N20676, N20669);
not NOT1 (N20677, N20673);
not NOT1 (N20678, N20675);
nor NOR2 (N20679, N20672, N5096);
and AND2 (N20680, N20649, N10576);
nor NOR3 (N20681, N20666, N17135, N17744);
buf BUF1 (N20682, N20679);
buf BUF1 (N20683, N20677);
nor NOR3 (N20684, N20676, N13998, N14114);
not NOT1 (N20685, N20680);
nor NOR2 (N20686, N20663, N5912);
xor XOR2 (N20687, N20674, N263);
xor XOR2 (N20688, N20683, N2354);
or OR3 (N20689, N20688, N11610, N11347);
nor NOR3 (N20690, N20687, N3005, N11014);
or OR3 (N20691, N20689, N20415, N139);
or OR4 (N20692, N20690, N3077, N2633, N10589);
and AND4 (N20693, N20671, N13361, N18927, N18621);
and AND3 (N20694, N20664, N6196, N9378);
and AND2 (N20695, N20692, N16865);
or OR2 (N20696, N20685, N5559);
nand NAND4 (N20697, N20694, N9028, N7891, N6309);
nor NOR2 (N20698, N20684, N8567);
or OR3 (N20699, N20681, N20698, N15500);
buf BUF1 (N20700, N16429);
xor XOR2 (N20701, N20693, N17650);
nand NAND2 (N20702, N20699, N214);
xor XOR2 (N20703, N20691, N10668);
or OR3 (N20704, N20695, N2617, N13707);
not NOT1 (N20705, N20697);
and AND2 (N20706, N20701, N10876);
nand NAND2 (N20707, N20696, N13771);
xor XOR2 (N20708, N20703, N6588);
and AND3 (N20709, N20702, N7569, N13892);
nand NAND3 (N20710, N20709, N17430, N18412);
nor NOR4 (N20711, N20706, N15675, N2396, N15334);
xor XOR2 (N20712, N20704, N5475);
xor XOR2 (N20713, N20712, N4773);
nand NAND4 (N20714, N20711, N3893, N7612, N17664);
nor NOR4 (N20715, N20713, N15597, N20551, N11971);
nand NAND3 (N20716, N20705, N14905, N10016);
nand NAND4 (N20717, N20686, N10006, N16509, N7972);
nor NOR2 (N20718, N20715, N16556);
xor XOR2 (N20719, N20682, N8127);
buf BUF1 (N20720, N20678);
and AND4 (N20721, N20710, N3267, N13294, N10039);
xor XOR2 (N20722, N20719, N7575);
not NOT1 (N20723, N20721);
not NOT1 (N20724, N20717);
or OR4 (N20725, N20723, N17735, N19587, N14350);
or OR2 (N20726, N20720, N20289);
buf BUF1 (N20727, N20724);
and AND3 (N20728, N20707, N1145, N7574);
nand NAND2 (N20729, N20722, N3859);
buf BUF1 (N20730, N20708);
buf BUF1 (N20731, N20716);
buf BUF1 (N20732, N20729);
not NOT1 (N20733, N20732);
xor XOR2 (N20734, N20714, N6587);
nor NOR4 (N20735, N20734, N4659, N17458, N5124);
xor XOR2 (N20736, N20731, N16240);
nor NOR4 (N20737, N20718, N7217, N14369, N3567);
nor NOR3 (N20738, N20726, N3120, N4131);
and AND2 (N20739, N20727, N4197);
or OR2 (N20740, N20736, N19788);
nand NAND3 (N20741, N20725, N2588, N2605);
not NOT1 (N20742, N20730);
or OR4 (N20743, N20742, N20639, N2735, N19481);
and AND3 (N20744, N20733, N1000, N254);
or OR4 (N20745, N20744, N760, N9448, N10537);
and AND4 (N20746, N20743, N5577, N10550, N10732);
buf BUF1 (N20747, N20746);
or OR2 (N20748, N20700, N13316);
nand NAND3 (N20749, N20748, N14477, N19052);
or OR3 (N20750, N20745, N7450, N2542);
xor XOR2 (N20751, N20735, N8601);
xor XOR2 (N20752, N20741, N651);
and AND3 (N20753, N20737, N337, N12433);
and AND2 (N20754, N20738, N5913);
nor NOR4 (N20755, N20752, N674, N2228, N10220);
and AND3 (N20756, N20755, N9956, N9317);
nand NAND2 (N20757, N20740, N226);
xor XOR2 (N20758, N20753, N12138);
and AND3 (N20759, N20728, N2885, N14144);
or OR3 (N20760, N20747, N10564, N259);
or OR4 (N20761, N20760, N16967, N14915, N19956);
xor XOR2 (N20762, N20759, N5608);
xor XOR2 (N20763, N20758, N3084);
xor XOR2 (N20764, N20754, N12291);
buf BUF1 (N20765, N20763);
or OR3 (N20766, N20757, N18667, N2462);
and AND3 (N20767, N20751, N19671, N1831);
xor XOR2 (N20768, N20765, N20434);
nor NOR4 (N20769, N20761, N15337, N2380, N16246);
not NOT1 (N20770, N20762);
nand NAND2 (N20771, N20750, N15185);
nand NAND2 (N20772, N20766, N14471);
xor XOR2 (N20773, N20739, N1155);
nand NAND3 (N20774, N20767, N9125, N16521);
and AND2 (N20775, N20769, N14985);
or OR4 (N20776, N20756, N14654, N4891, N14503);
xor XOR2 (N20777, N20770, N11582);
or OR2 (N20778, N20768, N16256);
and AND3 (N20779, N20776, N17854, N17985);
nand NAND3 (N20780, N20771, N15666, N18179);
buf BUF1 (N20781, N20774);
not NOT1 (N20782, N20781);
buf BUF1 (N20783, N20779);
and AND3 (N20784, N20778, N5525, N2628);
buf BUF1 (N20785, N20749);
not NOT1 (N20786, N20772);
nand NAND2 (N20787, N20773, N5429);
nor NOR4 (N20788, N20777, N2553, N13975, N20194);
buf BUF1 (N20789, N20783);
buf BUF1 (N20790, N20784);
nand NAND2 (N20791, N20790, N17839);
nor NOR4 (N20792, N20785, N4517, N9777, N1520);
or OR2 (N20793, N20791, N20296);
buf BUF1 (N20794, N20780);
buf BUF1 (N20795, N20775);
nand NAND2 (N20796, N20764, N607);
xor XOR2 (N20797, N20795, N14401);
xor XOR2 (N20798, N20789, N8705);
not NOT1 (N20799, N20786);
nand NAND2 (N20800, N20799, N13311);
or OR3 (N20801, N20798, N10561, N19873);
or OR4 (N20802, N20793, N6056, N7331, N79);
not NOT1 (N20803, N20782);
nor NOR4 (N20804, N20800, N1302, N4285, N2527);
and AND3 (N20805, N20792, N19962, N669);
not NOT1 (N20806, N20796);
xor XOR2 (N20807, N20788, N7282);
xor XOR2 (N20808, N20801, N11936);
or OR2 (N20809, N20808, N9129);
xor XOR2 (N20810, N20802, N19521);
nor NOR4 (N20811, N20787, N19035, N11807, N10293);
or OR2 (N20812, N20810, N12138);
and AND3 (N20813, N20803, N18159, N6102);
xor XOR2 (N20814, N20797, N2521);
buf BUF1 (N20815, N20807);
and AND2 (N20816, N20804, N18560);
nand NAND2 (N20817, N20805, N5773);
not NOT1 (N20818, N20814);
buf BUF1 (N20819, N20815);
xor XOR2 (N20820, N20817, N17694);
nor NOR4 (N20821, N20820, N12865, N3685, N4623);
buf BUF1 (N20822, N20812);
buf BUF1 (N20823, N20821);
nor NOR4 (N20824, N20818, N19562, N7041, N11752);
nor NOR3 (N20825, N20809, N6351, N16984);
or OR3 (N20826, N20813, N7002, N1035);
buf BUF1 (N20827, N20825);
buf BUF1 (N20828, N20794);
xor XOR2 (N20829, N20824, N15092);
not NOT1 (N20830, N20828);
buf BUF1 (N20831, N20819);
buf BUF1 (N20832, N20827);
xor XOR2 (N20833, N20806, N1492);
nand NAND2 (N20834, N20830, N5854);
nor NOR3 (N20835, N20829, N16072, N9264);
not NOT1 (N20836, N20823);
nand NAND3 (N20837, N20826, N18386, N9025);
and AND4 (N20838, N20811, N3337, N24, N1095);
xor XOR2 (N20839, N20837, N7356);
buf BUF1 (N20840, N20836);
and AND3 (N20841, N20839, N20408, N13878);
or OR2 (N20842, N20838, N17146);
buf BUF1 (N20843, N20831);
nand NAND2 (N20844, N20833, N10426);
nor NOR4 (N20845, N20843, N15957, N10444, N7643);
nor NOR4 (N20846, N20841, N18937, N20722, N12020);
nor NOR4 (N20847, N20834, N18951, N748, N3157);
xor XOR2 (N20848, N20816, N16213);
nor NOR3 (N20849, N20822, N11936, N2488);
buf BUF1 (N20850, N20842);
xor XOR2 (N20851, N20845, N20443);
xor XOR2 (N20852, N20832, N11598);
nor NOR3 (N20853, N20835, N18014, N8226);
buf BUF1 (N20854, N20846);
nor NOR3 (N20855, N20850, N3769, N5019);
or OR3 (N20856, N20844, N15655, N19646);
not NOT1 (N20857, N20854);
or OR3 (N20858, N20852, N11858, N10370);
and AND2 (N20859, N20857, N16564);
nand NAND4 (N20860, N20840, N856, N10923, N20647);
not NOT1 (N20861, N20853);
and AND3 (N20862, N20860, N8555, N4719);
or OR3 (N20863, N20859, N3148, N15961);
xor XOR2 (N20864, N20863, N13733);
not NOT1 (N20865, N20856);
buf BUF1 (N20866, N20864);
nor NOR2 (N20867, N20866, N10099);
nand NAND4 (N20868, N20867, N6709, N12744, N9270);
xor XOR2 (N20869, N20848, N6552);
xor XOR2 (N20870, N20849, N4924);
xor XOR2 (N20871, N20855, N3256);
nand NAND3 (N20872, N20869, N17397, N6968);
buf BUF1 (N20873, N20870);
or OR3 (N20874, N20861, N19285, N16220);
not NOT1 (N20875, N20865);
buf BUF1 (N20876, N20873);
and AND2 (N20877, N20851, N3256);
and AND2 (N20878, N20858, N17888);
xor XOR2 (N20879, N20871, N6613);
and AND2 (N20880, N20874, N6877);
or OR4 (N20881, N20862, N9776, N9081, N19160);
xor XOR2 (N20882, N20878, N6109);
not NOT1 (N20883, N20879);
or OR4 (N20884, N20847, N3954, N7206, N88);
or OR4 (N20885, N20875, N5982, N10654, N12191);
or OR2 (N20886, N20882, N4153);
buf BUF1 (N20887, N20885);
buf BUF1 (N20888, N20886);
or OR2 (N20889, N20872, N12183);
and AND2 (N20890, N20880, N12329);
nor NOR4 (N20891, N20877, N10918, N3323, N12039);
nor NOR3 (N20892, N20887, N19976, N15332);
or OR2 (N20893, N20876, N9752);
or OR4 (N20894, N20889, N1366, N8167, N18695);
and AND3 (N20895, N20893, N19279, N5816);
xor XOR2 (N20896, N20884, N16700);
not NOT1 (N20897, N20888);
nor NOR2 (N20898, N20868, N5949);
nand NAND3 (N20899, N20883, N2249, N7278);
nand NAND2 (N20900, N20894, N11790);
and AND2 (N20901, N20891, N10777);
nor NOR4 (N20902, N20899, N3808, N9961, N10406);
and AND3 (N20903, N20896, N9806, N1700);
nand NAND4 (N20904, N20900, N17354, N3365, N12732);
not NOT1 (N20905, N20898);
or OR2 (N20906, N20901, N2885);
not NOT1 (N20907, N20881);
or OR2 (N20908, N20892, N2470);
xor XOR2 (N20909, N20895, N18058);
xor XOR2 (N20910, N20906, N6116);
not NOT1 (N20911, N20903);
xor XOR2 (N20912, N20904, N12391);
not NOT1 (N20913, N20897);
buf BUF1 (N20914, N20910);
not NOT1 (N20915, N20912);
and AND2 (N20916, N20902, N19384);
nand NAND3 (N20917, N20890, N8980, N20507);
xor XOR2 (N20918, N20908, N10387);
or OR3 (N20919, N20914, N1114, N535);
or OR4 (N20920, N20917, N16575, N5830, N15074);
nor NOR3 (N20921, N20916, N15530, N20625);
nor NOR2 (N20922, N20919, N20338);
nand NAND3 (N20923, N20913, N6798, N6747);
and AND4 (N20924, N20921, N16121, N11520, N15966);
and AND4 (N20925, N20905, N17994, N9326, N1053);
nor NOR3 (N20926, N20922, N9383, N1456);
not NOT1 (N20927, N20925);
nor NOR2 (N20928, N20924, N11595);
buf BUF1 (N20929, N20918);
nand NAND2 (N20930, N20927, N18537);
and AND2 (N20931, N20911, N10445);
and AND2 (N20932, N20926, N14331);
not NOT1 (N20933, N20920);
nor NOR3 (N20934, N20930, N19634, N20174);
not NOT1 (N20935, N20915);
nor NOR2 (N20936, N20929, N8831);
buf BUF1 (N20937, N20907);
or OR3 (N20938, N20909, N11892, N13542);
nand NAND4 (N20939, N20936, N2402, N2242, N149);
xor XOR2 (N20940, N20934, N20204);
not NOT1 (N20941, N20937);
xor XOR2 (N20942, N20941, N10636);
xor XOR2 (N20943, N20938, N7201);
nor NOR3 (N20944, N20940, N13476, N17374);
xor XOR2 (N20945, N20928, N833);
not NOT1 (N20946, N20923);
and AND2 (N20947, N20945, N11576);
and AND2 (N20948, N20939, N10769);
buf BUF1 (N20949, N20933);
nand NAND3 (N20950, N20949, N9596, N17833);
and AND3 (N20951, N20942, N11027, N19330);
buf BUF1 (N20952, N20947);
buf BUF1 (N20953, N20946);
not NOT1 (N20954, N20943);
nand NAND2 (N20955, N20932, N3791);
or OR2 (N20956, N20955, N19272);
nor NOR3 (N20957, N20944, N19191, N13657);
xor XOR2 (N20958, N20954, N9145);
nor NOR3 (N20959, N20950, N18916, N11282);
nor NOR4 (N20960, N20935, N19647, N1368, N14331);
and AND3 (N20961, N20953, N7503, N18028);
xor XOR2 (N20962, N20961, N17614);
buf BUF1 (N20963, N20960);
buf BUF1 (N20964, N20931);
xor XOR2 (N20965, N20948, N12656);
not NOT1 (N20966, N20956);
buf BUF1 (N20967, N20957);
or OR3 (N20968, N20952, N15504, N2442);
or OR2 (N20969, N20958, N4816);
xor XOR2 (N20970, N20959, N13075);
nand NAND3 (N20971, N20968, N81, N6321);
buf BUF1 (N20972, N20963);
and AND2 (N20973, N20972, N1815);
nor NOR3 (N20974, N20951, N13024, N12627);
or OR3 (N20975, N20962, N7305, N6702);
nor NOR2 (N20976, N20969, N18302);
and AND3 (N20977, N20967, N9794, N5582);
nor NOR3 (N20978, N20973, N3896, N2351);
buf BUF1 (N20979, N20966);
and AND3 (N20980, N20979, N12446, N20072);
nor NOR2 (N20981, N20974, N7942);
nor NOR4 (N20982, N20978, N20647, N18740, N4294);
or OR2 (N20983, N20964, N2844);
or OR4 (N20984, N20970, N12258, N12913, N13081);
nor NOR3 (N20985, N20977, N17240, N7243);
not NOT1 (N20986, N20981);
not NOT1 (N20987, N20982);
xor XOR2 (N20988, N20987, N17776);
nor NOR4 (N20989, N20984, N19943, N20642, N10736);
nor NOR2 (N20990, N20989, N3549);
buf BUF1 (N20991, N20983);
nand NAND2 (N20992, N20991, N12898);
buf BUF1 (N20993, N20986);
buf BUF1 (N20994, N20990);
xor XOR2 (N20995, N20965, N17537);
or OR3 (N20996, N20975, N14089, N19116);
nor NOR3 (N20997, N20980, N12157, N13550);
xor XOR2 (N20998, N20992, N19059);
buf BUF1 (N20999, N20995);
nand NAND4 (N21000, N20976, N14353, N16878, N7766);
xor XOR2 (N21001, N20971, N10889);
xor XOR2 (N21002, N20998, N11767);
nand NAND3 (N21003, N20997, N8067, N11105);
not NOT1 (N21004, N21003);
not NOT1 (N21005, N20988);
not NOT1 (N21006, N20993);
not NOT1 (N21007, N21001);
not NOT1 (N21008, N21004);
xor XOR2 (N21009, N21007, N13578);
nor NOR2 (N21010, N21006, N8201);
not NOT1 (N21011, N20999);
buf BUF1 (N21012, N21010);
nor NOR4 (N21013, N20996, N12764, N522, N17173);
xor XOR2 (N21014, N21013, N15703);
nor NOR2 (N21015, N21012, N5138);
buf BUF1 (N21016, N20994);
buf BUF1 (N21017, N21014);
nor NOR3 (N21018, N21011, N9526, N4914);
xor XOR2 (N21019, N21017, N2854);
or OR2 (N21020, N21016, N4200);
nor NOR2 (N21021, N21005, N1230);
buf BUF1 (N21022, N21019);
not NOT1 (N21023, N21021);
nand NAND4 (N21024, N21018, N15774, N7721, N14148);
and AND2 (N21025, N21023, N3928);
or OR4 (N21026, N21020, N15643, N16005, N3981);
buf BUF1 (N21027, N21000);
nor NOR2 (N21028, N21009, N17934);
xor XOR2 (N21029, N21015, N17424);
and AND2 (N21030, N21024, N16578);
and AND3 (N21031, N21002, N15487, N5221);
xor XOR2 (N21032, N21031, N2538);
or OR4 (N21033, N21008, N6817, N6398, N10589);
xor XOR2 (N21034, N21033, N918);
nor NOR2 (N21035, N21030, N6247);
not NOT1 (N21036, N21034);
nand NAND3 (N21037, N21025, N12986, N13276);
xor XOR2 (N21038, N21035, N2168);
nor NOR3 (N21039, N21037, N5219, N15174);
xor XOR2 (N21040, N20985, N4347);
not NOT1 (N21041, N21038);
or OR4 (N21042, N21029, N7812, N12879, N7710);
buf BUF1 (N21043, N21036);
or OR2 (N21044, N21040, N9037);
or OR2 (N21045, N21039, N10389);
nand NAND4 (N21046, N21043, N3780, N357, N10399);
not NOT1 (N21047, N21044);
and AND2 (N21048, N21032, N6569);
nand NAND2 (N21049, N21045, N5645);
not NOT1 (N21050, N21026);
and AND2 (N21051, N21048, N8093);
nand NAND4 (N21052, N21051, N11439, N13535, N12532);
and AND3 (N21053, N21046, N20932, N17768);
nand NAND3 (N21054, N21047, N18484, N410);
and AND2 (N21055, N21053, N4403);
or OR4 (N21056, N21027, N18174, N10063, N6220);
not NOT1 (N21057, N21055);
not NOT1 (N21058, N21041);
not NOT1 (N21059, N21049);
and AND2 (N21060, N21042, N16712);
nor NOR4 (N21061, N21056, N2380, N13933, N28);
and AND2 (N21062, N21022, N12595);
nand NAND3 (N21063, N21028, N20962, N11678);
or OR2 (N21064, N21054, N10013);
buf BUF1 (N21065, N21059);
nand NAND2 (N21066, N21060, N182);
or OR2 (N21067, N21066, N3090);
or OR4 (N21068, N21064, N3228, N14184, N14441);
xor XOR2 (N21069, N21062, N4098);
xor XOR2 (N21070, N21063, N17268);
and AND4 (N21071, N21057, N12231, N4266, N10601);
buf BUF1 (N21072, N21061);
and AND3 (N21073, N21072, N7195, N12477);
nand NAND3 (N21074, N21052, N665, N10815);
and AND3 (N21075, N21070, N2662, N13876);
and AND4 (N21076, N21073, N9108, N1955, N11154);
and AND4 (N21077, N21068, N3216, N9784, N18293);
nor NOR2 (N21078, N21058, N10199);
nand NAND3 (N21079, N21075, N15582, N20910);
buf BUF1 (N21080, N21074);
xor XOR2 (N21081, N21071, N10066);
nand NAND3 (N21082, N21079, N19378, N16783);
buf BUF1 (N21083, N21065);
buf BUF1 (N21084, N21077);
not NOT1 (N21085, N21069);
not NOT1 (N21086, N21084);
and AND2 (N21087, N21078, N18594);
nor NOR4 (N21088, N21085, N20725, N12835, N9141);
buf BUF1 (N21089, N21080);
xor XOR2 (N21090, N21076, N2570);
nor NOR4 (N21091, N21088, N870, N16828, N6085);
and AND3 (N21092, N21087, N2221, N6206);
or OR3 (N21093, N21086, N12589, N17099);
not NOT1 (N21094, N21092);
nand NAND4 (N21095, N21067, N8640, N8519, N16808);
buf BUF1 (N21096, N21095);
nor NOR3 (N21097, N21090, N15042, N3478);
and AND4 (N21098, N21050, N14451, N6354, N12371);
nand NAND2 (N21099, N21081, N16288);
and AND2 (N21100, N21097, N8692);
nor NOR2 (N21101, N21094, N15752);
not NOT1 (N21102, N21098);
not NOT1 (N21103, N21083);
nand NAND2 (N21104, N21099, N16299);
nand NAND4 (N21105, N21103, N4566, N8154, N16081);
nor NOR4 (N21106, N21100, N6042, N4367, N9519);
buf BUF1 (N21107, N21082);
or OR4 (N21108, N21106, N19961, N14126, N2376);
xor XOR2 (N21109, N21096, N19404);
or OR2 (N21110, N21108, N5540);
nor NOR4 (N21111, N21091, N5145, N11254, N1477);
and AND4 (N21112, N21107, N12343, N14836, N7598);
nor NOR4 (N21113, N21101, N8450, N6538, N18697);
nor NOR4 (N21114, N21104, N17464, N19247, N1819);
xor XOR2 (N21115, N21089, N9956);
nand NAND3 (N21116, N21105, N2808, N15467);
xor XOR2 (N21117, N21116, N6001);
nor NOR4 (N21118, N21102, N7311, N18037, N4969);
or OR2 (N21119, N21117, N16578);
nor NOR4 (N21120, N21115, N4304, N10833, N15727);
or OR3 (N21121, N21113, N18489, N6230);
nand NAND2 (N21122, N21120, N8775);
nor NOR2 (N21123, N21114, N6221);
nor NOR2 (N21124, N21110, N13558);
not NOT1 (N21125, N21119);
xor XOR2 (N21126, N21112, N11709);
or OR3 (N21127, N21121, N10904, N14779);
and AND4 (N21128, N21125, N7406, N5729, N13411);
not NOT1 (N21129, N21124);
nor NOR3 (N21130, N21126, N13948, N6290);
nand NAND4 (N21131, N21111, N3589, N9532, N14602);
buf BUF1 (N21132, N21131);
and AND2 (N21133, N21093, N18095);
buf BUF1 (N21134, N21109);
nand NAND4 (N21135, N21118, N7522, N9334, N9944);
buf BUF1 (N21136, N21123);
not NOT1 (N21137, N21122);
and AND3 (N21138, N21135, N262, N5351);
nor NOR2 (N21139, N21127, N21004);
xor XOR2 (N21140, N21138, N2859);
or OR3 (N21141, N21139, N6700, N6433);
and AND2 (N21142, N21134, N20182);
xor XOR2 (N21143, N21141, N7809);
nor NOR4 (N21144, N21128, N6763, N21114, N11977);
not NOT1 (N21145, N21142);
or OR2 (N21146, N21132, N10700);
nor NOR3 (N21147, N21145, N20325, N20301);
not NOT1 (N21148, N21133);
and AND3 (N21149, N21129, N2962, N3767);
xor XOR2 (N21150, N21146, N4088);
nor NOR3 (N21151, N21140, N2478, N9873);
or OR4 (N21152, N21144, N1710, N2068, N16423);
and AND3 (N21153, N21151, N11322, N3391);
and AND2 (N21154, N21148, N10590);
nor NOR4 (N21155, N21130, N16691, N1840, N4398);
nor NOR2 (N21156, N21155, N18805);
and AND3 (N21157, N21152, N18811, N7038);
not NOT1 (N21158, N21137);
nand NAND4 (N21159, N21136, N6084, N3043, N15541);
buf BUF1 (N21160, N21149);
and AND2 (N21161, N21154, N6860);
buf BUF1 (N21162, N21160);
nand NAND3 (N21163, N21161, N1256, N15083);
or OR3 (N21164, N21156, N10574, N18591);
nand NAND4 (N21165, N21157, N9595, N10241, N16189);
or OR2 (N21166, N21147, N428);
xor XOR2 (N21167, N21164, N17686);
and AND3 (N21168, N21163, N9640, N8861);
buf BUF1 (N21169, N21166);
xor XOR2 (N21170, N21165, N16272);
nor NOR3 (N21171, N21167, N17527, N18456);
buf BUF1 (N21172, N21143);
nand NAND3 (N21173, N21158, N6924, N7558);
or OR4 (N21174, N21162, N9969, N7085, N6486);
or OR4 (N21175, N21168, N12039, N7481, N20909);
and AND4 (N21176, N21174, N4648, N1346, N6208);
nand NAND4 (N21177, N21169, N10083, N2974, N8247);
and AND4 (N21178, N21159, N15527, N18848, N14867);
not NOT1 (N21179, N21153);
not NOT1 (N21180, N21176);
nand NAND3 (N21181, N21177, N1052, N19383);
or OR4 (N21182, N21178, N240, N19423, N11674);
not NOT1 (N21183, N21181);
xor XOR2 (N21184, N21150, N14950);
buf BUF1 (N21185, N21183);
xor XOR2 (N21186, N21182, N17908);
nor NOR4 (N21187, N21170, N17568, N16094, N5159);
not NOT1 (N21188, N21171);
xor XOR2 (N21189, N21184, N5997);
nand NAND4 (N21190, N21172, N1718, N14346, N9953);
nor NOR2 (N21191, N21185, N4276);
or OR2 (N21192, N21179, N3481);
not NOT1 (N21193, N21188);
not NOT1 (N21194, N21175);
or OR3 (N21195, N21192, N14529, N6372);
nor NOR3 (N21196, N21187, N5627, N548);
or OR3 (N21197, N21186, N15083, N11065);
not NOT1 (N21198, N21194);
and AND4 (N21199, N21195, N2704, N21041, N15939);
nor NOR4 (N21200, N21190, N2370, N20948, N15151);
buf BUF1 (N21201, N21193);
nor NOR3 (N21202, N21189, N1043, N15174);
and AND3 (N21203, N21199, N11498, N8926);
nand NAND4 (N21204, N21200, N10890, N12025, N14250);
nor NOR4 (N21205, N21198, N4042, N16075, N10856);
buf BUF1 (N21206, N21203);
not NOT1 (N21207, N21202);
or OR4 (N21208, N21204, N3750, N13188, N18163);
not NOT1 (N21209, N21180);
not NOT1 (N21210, N21173);
xor XOR2 (N21211, N21197, N5665);
and AND3 (N21212, N21191, N2773, N17353);
buf BUF1 (N21213, N21196);
nor NOR4 (N21214, N21210, N17249, N15576, N19684);
nor NOR2 (N21215, N21209, N11273);
nor NOR2 (N21216, N21207, N14608);
buf BUF1 (N21217, N21208);
buf BUF1 (N21218, N21217);
and AND4 (N21219, N21205, N4931, N2577, N14117);
nor NOR3 (N21220, N21218, N989, N17335);
and AND3 (N21221, N21201, N20549, N12118);
nand NAND2 (N21222, N21212, N9291);
buf BUF1 (N21223, N21211);
nor NOR2 (N21224, N21222, N11544);
and AND4 (N21225, N21224, N5537, N17472, N457);
xor XOR2 (N21226, N21213, N351);
xor XOR2 (N21227, N21220, N1366);
nor NOR2 (N21228, N21221, N2209);
buf BUF1 (N21229, N21206);
xor XOR2 (N21230, N21225, N20933);
and AND4 (N21231, N21228, N5272, N9680, N3749);
nand NAND2 (N21232, N21226, N12450);
buf BUF1 (N21233, N21214);
nand NAND4 (N21234, N21227, N1119, N14249, N7172);
and AND2 (N21235, N21229, N7518);
nor NOR4 (N21236, N21215, N6065, N10032, N17933);
buf BUF1 (N21237, N21232);
or OR3 (N21238, N21216, N6535, N20807);
nand NAND3 (N21239, N21230, N16109, N16356);
nand NAND2 (N21240, N21223, N10103);
or OR2 (N21241, N21237, N6929);
xor XOR2 (N21242, N21234, N14537);
buf BUF1 (N21243, N21238);
xor XOR2 (N21244, N21239, N19390);
not NOT1 (N21245, N21231);
nand NAND3 (N21246, N21244, N1025, N11640);
buf BUF1 (N21247, N21219);
or OR2 (N21248, N21240, N19340);
xor XOR2 (N21249, N21246, N2456);
and AND2 (N21250, N21236, N9312);
xor XOR2 (N21251, N21235, N10042);
nand NAND3 (N21252, N21250, N13547, N15465);
buf BUF1 (N21253, N21251);
xor XOR2 (N21254, N21242, N10911);
buf BUF1 (N21255, N21241);
nand NAND3 (N21256, N21255, N18769, N4885);
buf BUF1 (N21257, N21233);
nand NAND4 (N21258, N21257, N7607, N20418, N9619);
and AND4 (N21259, N21248, N19192, N4652, N21045);
xor XOR2 (N21260, N21258, N4914);
buf BUF1 (N21261, N21243);
or OR2 (N21262, N21249, N1091);
nor NOR4 (N21263, N21247, N8742, N4486, N6395);
not NOT1 (N21264, N21261);
or OR2 (N21265, N21256, N6158);
and AND4 (N21266, N21259, N12504, N16829, N1384);
nor NOR4 (N21267, N21245, N1086, N13786, N2674);
and AND4 (N21268, N21264, N18816, N9716, N11737);
xor XOR2 (N21269, N21262, N18073);
and AND3 (N21270, N21253, N1268, N6319);
xor XOR2 (N21271, N21265, N13948);
nand NAND2 (N21272, N21271, N8438);
or OR3 (N21273, N21260, N15257, N5340);
and AND2 (N21274, N21252, N15761);
nand NAND3 (N21275, N21273, N2909, N12506);
not NOT1 (N21276, N21269);
nand NAND3 (N21277, N21254, N9773, N3915);
or OR2 (N21278, N21272, N747);
and AND2 (N21279, N21270, N13276);
or OR3 (N21280, N21278, N16324, N20474);
xor XOR2 (N21281, N21268, N10250);
buf BUF1 (N21282, N21277);
not NOT1 (N21283, N21274);
buf BUF1 (N21284, N21263);
xor XOR2 (N21285, N21283, N12802);
and AND3 (N21286, N21281, N16903, N18328);
nand NAND4 (N21287, N21279, N1435, N16112, N14855);
nand NAND2 (N21288, N21267, N5437);
not NOT1 (N21289, N21287);
or OR3 (N21290, N21289, N19842, N8983);
nand NAND3 (N21291, N21284, N11115, N18191);
xor XOR2 (N21292, N21290, N9990);
not NOT1 (N21293, N21280);
buf BUF1 (N21294, N21275);
not NOT1 (N21295, N21276);
and AND2 (N21296, N21294, N1563);
or OR2 (N21297, N21296, N517);
and AND3 (N21298, N21291, N9677, N14776);
buf BUF1 (N21299, N21295);
xor XOR2 (N21300, N21288, N21092);
nand NAND3 (N21301, N21300, N10014, N7636);
not NOT1 (N21302, N21285);
xor XOR2 (N21303, N21298, N3533);
or OR4 (N21304, N21282, N9863, N422, N5907);
or OR2 (N21305, N21303, N16943);
or OR3 (N21306, N21293, N20383, N4564);
xor XOR2 (N21307, N21286, N5806);
or OR2 (N21308, N21299, N19255);
nand NAND2 (N21309, N21305, N6128);
nor NOR2 (N21310, N21308, N2160);
and AND2 (N21311, N21301, N6723);
nor NOR3 (N21312, N21304, N930, N8336);
nand NAND2 (N21313, N21311, N3114);
and AND2 (N21314, N21313, N18507);
nand NAND2 (N21315, N21302, N4336);
nor NOR3 (N21316, N21309, N19479, N6671);
or OR3 (N21317, N21312, N13072, N19132);
nor NOR4 (N21318, N21297, N13575, N2899, N17974);
nor NOR2 (N21319, N21318, N7437);
nand NAND4 (N21320, N21292, N2924, N18453, N15372);
or OR3 (N21321, N21317, N687, N1572);
not NOT1 (N21322, N21320);
and AND4 (N21323, N21322, N18546, N16202, N10109);
and AND4 (N21324, N21314, N17028, N17143, N13046);
xor XOR2 (N21325, N21315, N10856);
buf BUF1 (N21326, N21321);
or OR4 (N21327, N21324, N18014, N1515, N4688);
and AND4 (N21328, N21319, N19533, N15865, N176);
nor NOR3 (N21329, N21310, N13239, N11004);
buf BUF1 (N21330, N21266);
nor NOR4 (N21331, N21326, N20103, N9453, N8234);
nor NOR4 (N21332, N21323, N9645, N15452, N9076);
and AND2 (N21333, N21331, N12592);
or OR2 (N21334, N21325, N5121);
nand NAND2 (N21335, N21316, N11166);
or OR2 (N21336, N21307, N7675);
and AND2 (N21337, N21330, N9991);
buf BUF1 (N21338, N21335);
nor NOR3 (N21339, N21338, N17972, N7162);
and AND3 (N21340, N21329, N5756, N20683);
buf BUF1 (N21341, N21328);
nor NOR3 (N21342, N21332, N4064, N12874);
buf BUF1 (N21343, N21337);
nand NAND2 (N21344, N21327, N8183);
or OR3 (N21345, N21342, N19080, N11513);
nor NOR4 (N21346, N21340, N17272, N1545, N18552);
buf BUF1 (N21347, N21339);
nor NOR2 (N21348, N21346, N6567);
nand NAND3 (N21349, N21343, N16055, N10820);
not NOT1 (N21350, N21345);
xor XOR2 (N21351, N21344, N5003);
and AND3 (N21352, N21334, N2981, N2571);
buf BUF1 (N21353, N21349);
nand NAND2 (N21354, N21353, N16248);
nor NOR2 (N21355, N21341, N17354);
buf BUF1 (N21356, N21352);
buf BUF1 (N21357, N21306);
and AND4 (N21358, N21351, N7274, N13244, N7312);
nand NAND4 (N21359, N21358, N2421, N10044, N8484);
nand NAND2 (N21360, N21333, N4781);
buf BUF1 (N21361, N21360);
buf BUF1 (N21362, N21347);
nor NOR3 (N21363, N21355, N2153, N2377);
xor XOR2 (N21364, N21361, N527);
not NOT1 (N21365, N21356);
nor NOR3 (N21366, N21354, N12802, N7019);
buf BUF1 (N21367, N21348);
nand NAND4 (N21368, N21367, N7544, N8798, N16037);
and AND4 (N21369, N21362, N8402, N15518, N5612);
xor XOR2 (N21370, N21336, N3551);
not NOT1 (N21371, N21369);
nand NAND4 (N21372, N21350, N19726, N13674, N6034);
nand NAND3 (N21373, N21357, N13210, N12933);
not NOT1 (N21374, N21364);
not NOT1 (N21375, N21365);
nor NOR4 (N21376, N21359, N1661, N4310, N15079);
xor XOR2 (N21377, N21376, N3068);
or OR4 (N21378, N21370, N16681, N7513, N2966);
not NOT1 (N21379, N21378);
xor XOR2 (N21380, N21363, N2293);
nand NAND3 (N21381, N21371, N4617, N13879);
buf BUF1 (N21382, N21379);
xor XOR2 (N21383, N21366, N13444);
nor NOR3 (N21384, N21375, N486, N14665);
nand NAND4 (N21385, N21380, N17785, N16804, N3316);
not NOT1 (N21386, N21377);
xor XOR2 (N21387, N21373, N12050);
not NOT1 (N21388, N21372);
nand NAND4 (N21389, N21388, N461, N19490, N14318);
nor NOR3 (N21390, N21387, N15682, N15783);
and AND2 (N21391, N21386, N4129);
and AND3 (N21392, N21374, N3058, N15485);
or OR3 (N21393, N21368, N16706, N18401);
buf BUF1 (N21394, N21381);
nor NOR4 (N21395, N21389, N4084, N20546, N6013);
xor XOR2 (N21396, N21394, N2642);
buf BUF1 (N21397, N21390);
xor XOR2 (N21398, N21395, N4744);
and AND3 (N21399, N21398, N18263, N17570);
or OR3 (N21400, N21393, N19759, N10275);
xor XOR2 (N21401, N21397, N5126);
not NOT1 (N21402, N21396);
and AND3 (N21403, N21384, N1626, N17991);
nand NAND3 (N21404, N21400, N13645, N16484);
nor NOR2 (N21405, N21392, N1192);
not NOT1 (N21406, N21385);
not NOT1 (N21407, N21391);
nor NOR4 (N21408, N21407, N16493, N6698, N20936);
or OR3 (N21409, N21404, N6493, N4489);
or OR3 (N21410, N21406, N9232, N3917);
not NOT1 (N21411, N21408);
xor XOR2 (N21412, N21401, N15880);
buf BUF1 (N21413, N21411);
nand NAND3 (N21414, N21409, N19502, N14444);
or OR2 (N21415, N21382, N19523);
nand NAND4 (N21416, N21403, N2231, N13058, N17178);
nand NAND2 (N21417, N21413, N8820);
nor NOR3 (N21418, N21414, N10413, N17744);
and AND3 (N21419, N21416, N10303, N834);
not NOT1 (N21420, N21402);
or OR3 (N21421, N21420, N3880, N606);
or OR3 (N21422, N21417, N9734, N4007);
nor NOR3 (N21423, N21418, N16847, N5165);
buf BUF1 (N21424, N21410);
not NOT1 (N21425, N21412);
xor XOR2 (N21426, N21424, N19259);
or OR4 (N21427, N21425, N17014, N5212, N21133);
or OR3 (N21428, N21422, N10966, N13849);
xor XOR2 (N21429, N21421, N15963);
xor XOR2 (N21430, N21405, N15521);
or OR4 (N21431, N21427, N13154, N1858, N19631);
buf BUF1 (N21432, N21423);
and AND3 (N21433, N21399, N17906, N9615);
or OR3 (N21434, N21433, N12538, N13812);
buf BUF1 (N21435, N21419);
not NOT1 (N21436, N21432);
nor NOR4 (N21437, N21434, N14821, N17074, N14100);
xor XOR2 (N21438, N21428, N783);
or OR4 (N21439, N21437, N12762, N6515, N21405);
and AND4 (N21440, N21435, N3993, N14237, N11774);
xor XOR2 (N21441, N21440, N3955);
nand NAND2 (N21442, N21426, N9913);
nand NAND2 (N21443, N21429, N16993);
not NOT1 (N21444, N21383);
and AND2 (N21445, N21431, N16532);
not NOT1 (N21446, N21415);
nor NOR3 (N21447, N21443, N7610, N18627);
xor XOR2 (N21448, N21436, N6114);
and AND3 (N21449, N21442, N12358, N19337);
xor XOR2 (N21450, N21444, N1604);
not NOT1 (N21451, N21445);
buf BUF1 (N21452, N21450);
xor XOR2 (N21453, N21451, N19482);
and AND3 (N21454, N21441, N1284, N12370);
nand NAND4 (N21455, N21454, N8790, N17926, N16825);
or OR4 (N21456, N21449, N9754, N7428, N9215);
buf BUF1 (N21457, N21453);
nor NOR3 (N21458, N21446, N11952, N9550);
nand NAND2 (N21459, N21457, N12414);
xor XOR2 (N21460, N21456, N21232);
buf BUF1 (N21461, N21430);
or OR2 (N21462, N21438, N18366);
not NOT1 (N21463, N21461);
or OR2 (N21464, N21455, N11239);
nand NAND3 (N21465, N21452, N14804, N18281);
not NOT1 (N21466, N21448);
xor XOR2 (N21467, N21464, N5572);
xor XOR2 (N21468, N21439, N19809);
nor NOR3 (N21469, N21467, N14943, N140);
buf BUF1 (N21470, N21463);
or OR2 (N21471, N21447, N2369);
and AND4 (N21472, N21465, N2950, N13260, N655);
buf BUF1 (N21473, N21462);
buf BUF1 (N21474, N21473);
not NOT1 (N21475, N21468);
not NOT1 (N21476, N21469);
nand NAND2 (N21477, N21459, N18762);
and AND2 (N21478, N21471, N16391);
xor XOR2 (N21479, N21475, N12389);
not NOT1 (N21480, N21470);
nor NOR2 (N21481, N21458, N4114);
and AND3 (N21482, N21479, N1707, N14012);
nor NOR2 (N21483, N21477, N6218);
and AND2 (N21484, N21482, N13977);
buf BUF1 (N21485, N21483);
and AND3 (N21486, N21460, N13997, N10805);
xor XOR2 (N21487, N21472, N16998);
not NOT1 (N21488, N21485);
nor NOR4 (N21489, N21476, N4587, N4779, N19420);
nand NAND3 (N21490, N21488, N9384, N14313);
and AND4 (N21491, N21484, N17003, N1570, N7380);
nor NOR3 (N21492, N21486, N13552, N14671);
or OR3 (N21493, N21466, N5337, N18582);
buf BUF1 (N21494, N21478);
xor XOR2 (N21495, N21493, N19785);
or OR2 (N21496, N21492, N7889);
or OR2 (N21497, N21491, N5282);
or OR3 (N21498, N21481, N8806, N13145);
nor NOR4 (N21499, N21487, N3960, N7223, N17464);
buf BUF1 (N21500, N21499);
nor NOR4 (N21501, N21494, N11173, N17868, N7983);
nand NAND3 (N21502, N21490, N394, N6301);
and AND4 (N21503, N21497, N4799, N11162, N16524);
buf BUF1 (N21504, N21496);
not NOT1 (N21505, N21498);
or OR2 (N21506, N21495, N10348);
buf BUF1 (N21507, N21503);
or OR2 (N21508, N21500, N19929);
xor XOR2 (N21509, N21501, N14633);
nor NOR2 (N21510, N21506, N5275);
nand NAND3 (N21511, N21509, N14867, N20514);
not NOT1 (N21512, N21489);
buf BUF1 (N21513, N21510);
buf BUF1 (N21514, N21505);
buf BUF1 (N21515, N21474);
and AND4 (N21516, N21502, N19683, N9882, N4998);
or OR3 (N21517, N21514, N18740, N19131);
and AND3 (N21518, N21504, N5710, N400);
nor NOR4 (N21519, N21512, N19102, N14988, N13200);
buf BUF1 (N21520, N21516);
nand NAND4 (N21521, N21511, N16397, N20893, N19158);
and AND4 (N21522, N21515, N3634, N2423, N16556);
or OR3 (N21523, N21518, N6187, N4490);
xor XOR2 (N21524, N21480, N20171);
or OR2 (N21525, N21517, N13489);
nor NOR3 (N21526, N21524, N19211, N18179);
or OR4 (N21527, N21508, N17408, N18569, N18547);
or OR3 (N21528, N21523, N6103, N1164);
buf BUF1 (N21529, N21521);
nand NAND2 (N21530, N21528, N15425);
nor NOR4 (N21531, N21519, N15465, N2594, N7477);
buf BUF1 (N21532, N21513);
nor NOR4 (N21533, N21526, N752, N7267, N15773);
and AND4 (N21534, N21520, N12655, N11101, N11896);
and AND3 (N21535, N21527, N20004, N2801);
or OR3 (N21536, N21533, N2648, N10832);
and AND4 (N21537, N21534, N9394, N5139, N10645);
not NOT1 (N21538, N21525);
nor NOR2 (N21539, N21530, N10952);
nand NAND2 (N21540, N21539, N16035);
not NOT1 (N21541, N21532);
xor XOR2 (N21542, N21536, N14464);
buf BUF1 (N21543, N21538);
xor XOR2 (N21544, N21535, N6663);
or OR2 (N21545, N21537, N17908);
nand NAND2 (N21546, N21541, N1557);
nand NAND3 (N21547, N21543, N19886, N169);
buf BUF1 (N21548, N21542);
buf BUF1 (N21549, N21507);
not NOT1 (N21550, N21546);
and AND4 (N21551, N21549, N20667, N4314, N1860);
xor XOR2 (N21552, N21540, N15795);
and AND3 (N21553, N21544, N3126, N18118);
and AND3 (N21554, N21547, N19588, N1511);
nor NOR3 (N21555, N21551, N5965, N14044);
buf BUF1 (N21556, N21531);
buf BUF1 (N21557, N21554);
nor NOR4 (N21558, N21553, N14688, N17959, N15923);
or OR2 (N21559, N21558, N6697);
buf BUF1 (N21560, N21550);
buf BUF1 (N21561, N21556);
nand NAND2 (N21562, N21557, N11128);
xor XOR2 (N21563, N21561, N7190);
nor NOR3 (N21564, N21562, N19261, N8707);
not NOT1 (N21565, N21555);
not NOT1 (N21566, N21559);
nand NAND3 (N21567, N21545, N15475, N722);
not NOT1 (N21568, N21552);
or OR3 (N21569, N21567, N4578, N175);
xor XOR2 (N21570, N21529, N7168);
not NOT1 (N21571, N21522);
and AND2 (N21572, N21569, N5924);
not NOT1 (N21573, N21568);
not NOT1 (N21574, N21560);
not NOT1 (N21575, N21565);
nand NAND4 (N21576, N21548, N5806, N1367, N7840);
and AND3 (N21577, N21574, N3244, N4025);
buf BUF1 (N21578, N21566);
nand NAND3 (N21579, N21571, N18975, N14827);
not NOT1 (N21580, N21575);
or OR2 (N21581, N21564, N4150);
or OR2 (N21582, N21580, N19472);
xor XOR2 (N21583, N21573, N4770);
or OR4 (N21584, N21582, N12479, N1140, N2734);
nand NAND4 (N21585, N21572, N18016, N4953, N9998);
nand NAND3 (N21586, N21579, N8872, N7272);
or OR4 (N21587, N21576, N16693, N18556, N12264);
not NOT1 (N21588, N21570);
nor NOR3 (N21589, N21577, N2490, N8605);
nand NAND3 (N21590, N21586, N5258, N2613);
not NOT1 (N21591, N21581);
not NOT1 (N21592, N21578);
buf BUF1 (N21593, N21587);
nor NOR4 (N21594, N21593, N2317, N17428, N16818);
nand NAND2 (N21595, N21590, N16800);
and AND2 (N21596, N21563, N16627);
buf BUF1 (N21597, N21589);
xor XOR2 (N21598, N21585, N6028);
not NOT1 (N21599, N21592);
xor XOR2 (N21600, N21583, N8670);
or OR3 (N21601, N21591, N3830, N3058);
or OR4 (N21602, N21584, N18448, N19400, N2898);
xor XOR2 (N21603, N21596, N18239);
nor NOR3 (N21604, N21603, N13328, N9522);
and AND2 (N21605, N21602, N13931);
nor NOR3 (N21606, N21588, N911, N8868);
not NOT1 (N21607, N21598);
not NOT1 (N21608, N21604);
and AND4 (N21609, N21606, N9941, N12161, N14608);
nand NAND3 (N21610, N21609, N17414, N10803);
not NOT1 (N21611, N21608);
buf BUF1 (N21612, N21594);
not NOT1 (N21613, N21611);
nor NOR3 (N21614, N21600, N12782, N17842);
xor XOR2 (N21615, N21610, N5623);
nand NAND3 (N21616, N21597, N4921, N9931);
nor NOR2 (N21617, N21615, N19435);
or OR4 (N21618, N21607, N19540, N20069, N14001);
nor NOR2 (N21619, N21616, N19213);
and AND4 (N21620, N21612, N16436, N14781, N4880);
nand NAND4 (N21621, N21620, N9298, N4105, N1014);
nor NOR4 (N21622, N21614, N13924, N13437, N21619);
xor XOR2 (N21623, N17889, N313);
buf BUF1 (N21624, N21617);
nand NAND2 (N21625, N21613, N10586);
and AND2 (N21626, N21605, N9592);
or OR2 (N21627, N21622, N3462);
nor NOR4 (N21628, N21624, N16662, N7630, N17226);
nand NAND3 (N21629, N21621, N20299, N4816);
nand NAND2 (N21630, N21626, N13460);
and AND2 (N21631, N21599, N17059);
xor XOR2 (N21632, N21618, N767);
and AND3 (N21633, N21595, N17513, N1178);
buf BUF1 (N21634, N21628);
nor NOR3 (N21635, N21633, N11364, N11963);
not NOT1 (N21636, N21635);
and AND3 (N21637, N21601, N4987, N3447);
not NOT1 (N21638, N21623);
buf BUF1 (N21639, N21632);
buf BUF1 (N21640, N21637);
or OR3 (N21641, N21634, N14286, N18983);
xor XOR2 (N21642, N21630, N20051);
or OR2 (N21643, N21629, N5258);
xor XOR2 (N21644, N21643, N17344);
and AND2 (N21645, N21642, N8063);
not NOT1 (N21646, N21638);
buf BUF1 (N21647, N21645);
and AND2 (N21648, N21641, N4722);
and AND4 (N21649, N21646, N4935, N3460, N897);
not NOT1 (N21650, N21640);
or OR4 (N21651, N21647, N16091, N19094, N8993);
xor XOR2 (N21652, N21648, N16461);
and AND4 (N21653, N21649, N7133, N11220, N20358);
nand NAND2 (N21654, N21636, N19076);
buf BUF1 (N21655, N21652);
buf BUF1 (N21656, N21625);
xor XOR2 (N21657, N21653, N11275);
xor XOR2 (N21658, N21657, N4724);
nor NOR4 (N21659, N21650, N17363, N6235, N20123);
buf BUF1 (N21660, N21659);
xor XOR2 (N21661, N21639, N642);
nor NOR4 (N21662, N21656, N16277, N5287, N20810);
not NOT1 (N21663, N21627);
nor NOR3 (N21664, N21655, N17888, N13237);
xor XOR2 (N21665, N21654, N11403);
xor XOR2 (N21666, N21664, N13814);
nand NAND2 (N21667, N21662, N9923);
nor NOR2 (N21668, N21665, N13605);
and AND2 (N21669, N21667, N13590);
and AND4 (N21670, N21668, N19191, N12157, N15991);
or OR2 (N21671, N21644, N3803);
xor XOR2 (N21672, N21663, N5214);
not NOT1 (N21673, N21672);
buf BUF1 (N21674, N21661);
nand NAND4 (N21675, N21670, N19643, N18993, N13612);
or OR3 (N21676, N21671, N5652, N11883);
nand NAND3 (N21677, N21631, N20308, N10978);
xor XOR2 (N21678, N21666, N20861);
or OR2 (N21679, N21674, N11516);
or OR3 (N21680, N21676, N6438, N2658);
xor XOR2 (N21681, N21678, N701);
xor XOR2 (N21682, N21658, N16954);
nor NOR3 (N21683, N21669, N15324, N6975);
or OR4 (N21684, N21677, N8816, N13054, N18711);
or OR4 (N21685, N21679, N9364, N18422, N2353);
not NOT1 (N21686, N21685);
or OR2 (N21687, N21682, N8122);
xor XOR2 (N21688, N21687, N4444);
and AND4 (N21689, N21688, N1988, N1677, N1991);
xor XOR2 (N21690, N21689, N2297);
not NOT1 (N21691, N21673);
xor XOR2 (N21692, N21686, N11784);
nand NAND3 (N21693, N21660, N9207, N3624);
or OR2 (N21694, N21675, N9155);
nor NOR3 (N21695, N21693, N3874, N17228);
nor NOR3 (N21696, N21651, N3139, N9600);
nand NAND2 (N21697, N21683, N20916);
or OR2 (N21698, N21696, N2447);
and AND2 (N21699, N21691, N11469);
xor XOR2 (N21700, N21698, N16850);
buf BUF1 (N21701, N21700);
nand NAND4 (N21702, N21690, N1070, N9744, N1904);
and AND4 (N21703, N21681, N11381, N7738, N15327);
xor XOR2 (N21704, N21699, N10000);
and AND3 (N21705, N21703, N8243, N8128);
not NOT1 (N21706, N21702);
buf BUF1 (N21707, N21694);
buf BUF1 (N21708, N21706);
or OR2 (N21709, N21704, N19225);
or OR2 (N21710, N21709, N9218);
nand NAND2 (N21711, N21701, N9529);
nand NAND3 (N21712, N21711, N13292, N16233);
xor XOR2 (N21713, N21684, N14395);
or OR4 (N21714, N21692, N3909, N7131, N14541);
buf BUF1 (N21715, N21697);
buf BUF1 (N21716, N21680);
buf BUF1 (N21717, N21705);
not NOT1 (N21718, N21714);
buf BUF1 (N21719, N21708);
or OR3 (N21720, N21715, N1387, N9905);
not NOT1 (N21721, N21717);
nor NOR2 (N21722, N21719, N4082);
xor XOR2 (N21723, N21722, N14775);
nand NAND3 (N21724, N21695, N13485, N3506);
nand NAND2 (N21725, N21707, N20205);
xor XOR2 (N21726, N21721, N1886);
not NOT1 (N21727, N21720);
nor NOR3 (N21728, N21713, N20873, N9583);
not NOT1 (N21729, N21724);
buf BUF1 (N21730, N21725);
nand NAND2 (N21731, N21710, N16356);
and AND4 (N21732, N21730, N438, N19048, N631);
nor NOR3 (N21733, N21723, N17264, N4138);
or OR2 (N21734, N21729, N10537);
buf BUF1 (N21735, N21726);
or OR4 (N21736, N21731, N11872, N6108, N20367);
nor NOR3 (N21737, N21727, N7221, N5249);
not NOT1 (N21738, N21712);
and AND3 (N21739, N21734, N10975, N12646);
nand NAND2 (N21740, N21737, N12637);
buf BUF1 (N21741, N21716);
not NOT1 (N21742, N21739);
xor XOR2 (N21743, N21728, N12858);
not NOT1 (N21744, N21718);
and AND2 (N21745, N21738, N12127);
nand NAND4 (N21746, N21743, N9926, N5882, N1406);
and AND3 (N21747, N21746, N6043, N13083);
and AND3 (N21748, N21745, N19939, N4665);
buf BUF1 (N21749, N21744);
nor NOR3 (N21750, N21741, N12318, N15720);
xor XOR2 (N21751, N21740, N4011);
or OR3 (N21752, N21733, N11244, N19671);
nor NOR2 (N21753, N21750, N21172);
buf BUF1 (N21754, N21748);
or OR3 (N21755, N21736, N2606, N6072);
not NOT1 (N21756, N21753);
or OR3 (N21757, N21754, N13835, N12440);
nor NOR3 (N21758, N21735, N3159, N5245);
not NOT1 (N21759, N21747);
and AND4 (N21760, N21757, N13359, N12429, N3722);
buf BUF1 (N21761, N21752);
nand NAND4 (N21762, N21759, N3079, N18620, N21457);
nor NOR3 (N21763, N21762, N20570, N12831);
xor XOR2 (N21764, N21732, N13809);
buf BUF1 (N21765, N21755);
buf BUF1 (N21766, N21763);
xor XOR2 (N21767, N21765, N17571);
and AND4 (N21768, N21749, N3045, N986, N20727);
nand NAND4 (N21769, N21767, N11863, N16174, N8985);
or OR2 (N21770, N21768, N250);
nand NAND4 (N21771, N21766, N5938, N17157, N737);
xor XOR2 (N21772, N21758, N5664);
or OR3 (N21773, N21770, N9767, N15010);
nand NAND2 (N21774, N21764, N4686);
nor NOR4 (N21775, N21751, N17493, N20863, N12786);
not NOT1 (N21776, N21774);
or OR4 (N21777, N21760, N18989, N14102, N9260);
or OR2 (N21778, N21742, N9638);
nand NAND4 (N21779, N21773, N14487, N11020, N15885);
or OR2 (N21780, N21776, N7360);
or OR3 (N21781, N21778, N10659, N844);
not NOT1 (N21782, N21771);
xor XOR2 (N21783, N21780, N14147);
and AND3 (N21784, N21761, N347, N5229);
and AND2 (N21785, N21772, N4416);
xor XOR2 (N21786, N21782, N14992);
xor XOR2 (N21787, N21786, N8217);
or OR4 (N21788, N21784, N6824, N13554, N11720);
not NOT1 (N21789, N21777);
not NOT1 (N21790, N21788);
xor XOR2 (N21791, N21775, N329);
nor NOR4 (N21792, N21756, N17534, N6494, N155);
or OR2 (N21793, N21783, N7653);
nand NAND4 (N21794, N21790, N15453, N1718, N17227);
not NOT1 (N21795, N21785);
nand NAND4 (N21796, N21779, N7598, N14714, N21521);
buf BUF1 (N21797, N21789);
and AND4 (N21798, N21794, N4706, N17200, N9534);
not NOT1 (N21799, N21787);
or OR4 (N21800, N21795, N9570, N7366, N2952);
nor NOR3 (N21801, N21791, N14281, N11716);
nand NAND2 (N21802, N21797, N15697);
nand NAND2 (N21803, N21798, N7781);
nand NAND2 (N21804, N21799, N6959);
buf BUF1 (N21805, N21800);
not NOT1 (N21806, N21801);
not NOT1 (N21807, N21805);
xor XOR2 (N21808, N21793, N9227);
nand NAND4 (N21809, N21796, N21207, N18154, N13288);
nor NOR3 (N21810, N21803, N5243, N16499);
xor XOR2 (N21811, N21804, N12406);
not NOT1 (N21812, N21807);
not NOT1 (N21813, N21812);
and AND4 (N21814, N21806, N792, N873, N1360);
and AND3 (N21815, N21813, N4564, N4191);
and AND2 (N21816, N21808, N2005);
buf BUF1 (N21817, N21811);
nand NAND4 (N21818, N21769, N21539, N21083, N21574);
xor XOR2 (N21819, N21810, N7919);
not NOT1 (N21820, N21816);
or OR3 (N21821, N21815, N2310, N21196);
xor XOR2 (N21822, N21802, N8368);
buf BUF1 (N21823, N21818);
not NOT1 (N21824, N21817);
nor NOR3 (N21825, N21814, N19673, N21717);
or OR2 (N21826, N21820, N18095);
not NOT1 (N21827, N21826);
nor NOR2 (N21828, N21821, N19062);
buf BUF1 (N21829, N21822);
nand NAND2 (N21830, N21828, N14688);
nor NOR4 (N21831, N21809, N20930, N82, N8283);
not NOT1 (N21832, N21831);
buf BUF1 (N21833, N21823);
not NOT1 (N21834, N21781);
not NOT1 (N21835, N21834);
nor NOR2 (N21836, N21833, N8366);
xor XOR2 (N21837, N21792, N18766);
nand NAND2 (N21838, N21835, N11943);
nor NOR4 (N21839, N21819, N6608, N10868, N16797);
buf BUF1 (N21840, N21827);
not NOT1 (N21841, N21838);
xor XOR2 (N21842, N21837, N6078);
not NOT1 (N21843, N21839);
and AND2 (N21844, N21832, N11795);
nand NAND3 (N21845, N21825, N5502, N9477);
and AND3 (N21846, N21844, N13706, N6572);
xor XOR2 (N21847, N21830, N7690);
not NOT1 (N21848, N21843);
and AND3 (N21849, N21836, N13009, N9354);
and AND2 (N21850, N21845, N17290);
buf BUF1 (N21851, N21829);
nand NAND2 (N21852, N21841, N7258);
buf BUF1 (N21853, N21847);
xor XOR2 (N21854, N21824, N7519);
or OR4 (N21855, N21854, N9127, N4180, N10517);
nand NAND2 (N21856, N21855, N21748);
xor XOR2 (N21857, N21849, N11248);
buf BUF1 (N21858, N21848);
nand NAND4 (N21859, N21857, N283, N12578, N10177);
nor NOR3 (N21860, N21859, N450, N9117);
or OR3 (N21861, N21853, N5147, N15476);
nor NOR4 (N21862, N21851, N8507, N17361, N13923);
and AND3 (N21863, N21861, N12098, N19137);
and AND4 (N21864, N21863, N13906, N5113, N12657);
xor XOR2 (N21865, N21852, N20359);
not NOT1 (N21866, N21860);
or OR2 (N21867, N21840, N17783);
xor XOR2 (N21868, N21856, N11779);
nand NAND2 (N21869, N21868, N20974);
buf BUF1 (N21870, N21867);
not NOT1 (N21871, N21858);
nor NOR3 (N21872, N21846, N12042, N6139);
xor XOR2 (N21873, N21842, N21064);
nand NAND3 (N21874, N21869, N4066, N7523);
xor XOR2 (N21875, N21866, N18284);
or OR2 (N21876, N21864, N19177);
or OR4 (N21877, N21873, N2545, N1988, N4849);
nor NOR3 (N21878, N21875, N1043, N20779);
xor XOR2 (N21879, N21850, N14103);
and AND4 (N21880, N21878, N3099, N5199, N307);
and AND3 (N21881, N21862, N13034, N19977);
nor NOR3 (N21882, N21870, N19846, N9360);
or OR2 (N21883, N21876, N2306);
nand NAND3 (N21884, N21871, N14123, N21844);
buf BUF1 (N21885, N21879);
or OR2 (N21886, N21877, N13816);
buf BUF1 (N21887, N21883);
and AND2 (N21888, N21885, N20773);
nor NOR4 (N21889, N21880, N11974, N21838, N10560);
not NOT1 (N21890, N21884);
buf BUF1 (N21891, N21890);
not NOT1 (N21892, N21882);
not NOT1 (N21893, N21888);
and AND4 (N21894, N21886, N11299, N18293, N2740);
not NOT1 (N21895, N21881);
buf BUF1 (N21896, N21874);
buf BUF1 (N21897, N21865);
nor NOR3 (N21898, N21872, N18457, N10455);
nor NOR3 (N21899, N21895, N2755, N14848);
xor XOR2 (N21900, N21889, N20237);
or OR3 (N21901, N21892, N16883, N19788);
nor NOR4 (N21902, N21893, N13047, N130, N3258);
not NOT1 (N21903, N21887);
nand NAND2 (N21904, N21901, N14528);
not NOT1 (N21905, N21898);
or OR4 (N21906, N21902, N13460, N11959, N9214);
xor XOR2 (N21907, N21904, N15385);
nand NAND3 (N21908, N21896, N18544, N12212);
not NOT1 (N21909, N21905);
and AND4 (N21910, N21894, N7982, N5558, N18264);
not NOT1 (N21911, N21899);
or OR3 (N21912, N21900, N20167, N12434);
and AND4 (N21913, N21912, N7217, N15816, N9085);
xor XOR2 (N21914, N21913, N17167);
xor XOR2 (N21915, N21910, N11542);
not NOT1 (N21916, N21915);
or OR2 (N21917, N21906, N19918);
buf BUF1 (N21918, N21903);
or OR4 (N21919, N21916, N11064, N4025, N12495);
nand NAND3 (N21920, N21917, N6292, N9145);
and AND2 (N21921, N21920, N8194);
nor NOR2 (N21922, N21914, N4469);
nor NOR2 (N21923, N21908, N13198);
not NOT1 (N21924, N21922);
and AND3 (N21925, N21919, N7412, N8180);
not NOT1 (N21926, N21891);
or OR2 (N21927, N21911, N2757);
nor NOR2 (N21928, N21907, N12496);
or OR2 (N21929, N21926, N15762);
not NOT1 (N21930, N21923);
buf BUF1 (N21931, N21921);
or OR4 (N21932, N21929, N3037, N13830, N14722);
and AND3 (N21933, N21918, N16033, N2769);
not NOT1 (N21934, N21932);
or OR4 (N21935, N21927, N21647, N528, N11324);
nor NOR2 (N21936, N21924, N6586);
not NOT1 (N21937, N21930);
buf BUF1 (N21938, N21931);
buf BUF1 (N21939, N21937);
or OR3 (N21940, N21928, N5857, N829);
not NOT1 (N21941, N21935);
not NOT1 (N21942, N21909);
or OR2 (N21943, N21936, N51);
not NOT1 (N21944, N21933);
nand NAND2 (N21945, N21938, N15157);
xor XOR2 (N21946, N21945, N18941);
nand NAND4 (N21947, N21941, N9229, N12877, N11914);
nor NOR3 (N21948, N21939, N3471, N4802);
nor NOR3 (N21949, N21947, N3001, N16011);
and AND2 (N21950, N21943, N19881);
nand NAND2 (N21951, N21940, N21317);
not NOT1 (N21952, N21951);
and AND3 (N21953, N21934, N1638, N18178);
and AND2 (N21954, N21952, N2444);
nor NOR2 (N21955, N21953, N4507);
not NOT1 (N21956, N21948);
or OR2 (N21957, N21944, N21002);
buf BUF1 (N21958, N21955);
or OR4 (N21959, N21897, N8780, N18664, N378);
not NOT1 (N21960, N21959);
nand NAND2 (N21961, N21956, N4763);
buf BUF1 (N21962, N21961);
not NOT1 (N21963, N21954);
or OR3 (N21964, N21958, N3488, N4697);
or OR2 (N21965, N21957, N1625);
not NOT1 (N21966, N21960);
or OR3 (N21967, N21925, N4, N20235);
buf BUF1 (N21968, N21967);
and AND2 (N21969, N21965, N971);
not NOT1 (N21970, N21964);
xor XOR2 (N21971, N21962, N5839);
or OR2 (N21972, N21946, N17933);
not NOT1 (N21973, N21966);
xor XOR2 (N21974, N21950, N13754);
nand NAND4 (N21975, N21973, N15585, N14272, N3824);
buf BUF1 (N21976, N21968);
or OR2 (N21977, N21942, N17089);
nor NOR3 (N21978, N21972, N14610, N7555);
not NOT1 (N21979, N21949);
nor NOR4 (N21980, N21977, N12958, N15768, N3360);
nor NOR3 (N21981, N21971, N10770, N3614);
or OR4 (N21982, N21963, N4357, N10306, N8744);
nor NOR4 (N21983, N21981, N4086, N15539, N11155);
or OR2 (N21984, N21976, N1831);
or OR2 (N21985, N21969, N21645);
buf BUF1 (N21986, N21982);
or OR4 (N21987, N21986, N4880, N4365, N18370);
nor NOR2 (N21988, N21970, N1757);
and AND2 (N21989, N21974, N13766);
buf BUF1 (N21990, N21989);
xor XOR2 (N21991, N21988, N18607);
and AND3 (N21992, N21979, N2847, N21277);
nor NOR2 (N21993, N21987, N13353);
nand NAND3 (N21994, N21985, N3643, N1607);
nand NAND2 (N21995, N21994, N5441);
or OR3 (N21996, N21984, N17107, N15014);
not NOT1 (N21997, N21992);
or OR4 (N21998, N21993, N6922, N2344, N21483);
and AND4 (N21999, N21997, N6904, N16794, N6530);
buf BUF1 (N22000, N21999);
nor NOR3 (N22001, N21996, N18042, N7583);
or OR2 (N22002, N21998, N17992);
not NOT1 (N22003, N21978);
nand NAND3 (N22004, N21983, N21557, N14080);
xor XOR2 (N22005, N22003, N20305);
xor XOR2 (N22006, N21995, N10372);
xor XOR2 (N22007, N22001, N2982);
and AND4 (N22008, N21991, N6276, N11882, N20313);
or OR3 (N22009, N21990, N17034, N7196);
or OR2 (N22010, N22002, N15639);
not NOT1 (N22011, N22004);
not NOT1 (N22012, N22007);
nand NAND3 (N22013, N22005, N2153, N21341);
or OR2 (N22014, N22009, N12758);
nand NAND2 (N22015, N22008, N4161);
not NOT1 (N22016, N22015);
and AND2 (N22017, N22006, N21374);
nor NOR2 (N22018, N22014, N2854);
and AND4 (N22019, N21980, N223, N17935, N557);
or OR3 (N22020, N22012, N10819, N16844);
nor NOR3 (N22021, N22017, N5505, N6457);
nand NAND2 (N22022, N22018, N18504);
buf BUF1 (N22023, N22011);
not NOT1 (N22024, N22000);
buf BUF1 (N22025, N22013);
and AND4 (N22026, N22025, N5579, N10424, N19391);
nor NOR3 (N22027, N21975, N15298, N12831);
nor NOR3 (N22028, N22026, N14201, N4587);
xor XOR2 (N22029, N22023, N5599);
not NOT1 (N22030, N22029);
nor NOR3 (N22031, N22020, N21452, N1219);
or OR2 (N22032, N22027, N9051);
nand NAND2 (N22033, N22028, N19188);
nor NOR3 (N22034, N22033, N18833, N7861);
buf BUF1 (N22035, N22030);
not NOT1 (N22036, N22010);
not NOT1 (N22037, N22021);
or OR4 (N22038, N22035, N5737, N21401, N4452);
nand NAND3 (N22039, N22031, N20218, N19208);
not NOT1 (N22040, N22034);
and AND4 (N22041, N22037, N1001, N5134, N6787);
nand NAND2 (N22042, N22022, N8657);
buf BUF1 (N22043, N22024);
or OR4 (N22044, N22016, N4753, N15047, N17723);
xor XOR2 (N22045, N22044, N16767);
and AND2 (N22046, N22036, N4774);
not NOT1 (N22047, N22038);
nand NAND3 (N22048, N22039, N17741, N7403);
or OR2 (N22049, N22040, N1097);
nor NOR2 (N22050, N22047, N13575);
nand NAND2 (N22051, N22046, N5585);
nor NOR3 (N22052, N22045, N868, N343);
xor XOR2 (N22053, N22049, N5624);
nand NAND3 (N22054, N22041, N17827, N9699);
buf BUF1 (N22055, N22052);
buf BUF1 (N22056, N22042);
not NOT1 (N22057, N22050);
and AND2 (N22058, N22057, N20435);
not NOT1 (N22059, N22056);
xor XOR2 (N22060, N22053, N18631);
nand NAND4 (N22061, N22060, N2070, N16404, N4819);
and AND3 (N22062, N22058, N16707, N2422);
buf BUF1 (N22063, N22051);
nand NAND2 (N22064, N22032, N17746);
not NOT1 (N22065, N22059);
nand NAND3 (N22066, N22064, N7408, N12390);
nor NOR4 (N22067, N22066, N8855, N15979, N21946);
not NOT1 (N22068, N22043);
buf BUF1 (N22069, N22054);
nand NAND3 (N22070, N22055, N6650, N11582);
nand NAND3 (N22071, N22065, N16112, N14015);
buf BUF1 (N22072, N22067);
nor NOR2 (N22073, N22068, N3154);
nand NAND3 (N22074, N22073, N11262, N13736);
nor NOR2 (N22075, N22070, N1766);
and AND4 (N22076, N22069, N1699, N9575, N16520);
and AND3 (N22077, N22062, N19897, N20234);
nand NAND2 (N22078, N22077, N15894);
xor XOR2 (N22079, N22078, N8878);
not NOT1 (N22080, N22061);
nand NAND2 (N22081, N22048, N12862);
or OR2 (N22082, N22074, N3950);
nor NOR2 (N22083, N22076, N12708);
and AND2 (N22084, N22082, N15352);
xor XOR2 (N22085, N22084, N21664);
nand NAND3 (N22086, N22063, N14449, N17318);
xor XOR2 (N22087, N22075, N4050);
xor XOR2 (N22088, N22081, N18602);
xor XOR2 (N22089, N22086, N4760);
buf BUF1 (N22090, N22079);
buf BUF1 (N22091, N22071);
or OR2 (N22092, N22087, N15348);
nand NAND3 (N22093, N22092, N10555, N930);
xor XOR2 (N22094, N22085, N14397);
nand NAND4 (N22095, N22072, N12865, N21551, N18140);
nand NAND3 (N22096, N22088, N5529, N18398);
and AND4 (N22097, N22080, N3750, N10957, N16271);
and AND4 (N22098, N22094, N18160, N15512, N4947);
not NOT1 (N22099, N22096);
nor NOR4 (N22100, N22083, N4129, N2626, N9000);
nor NOR4 (N22101, N22089, N8624, N3092, N20655);
not NOT1 (N22102, N22091);
not NOT1 (N22103, N22090);
xor XOR2 (N22104, N22101, N2091);
and AND2 (N22105, N22102, N883);
not NOT1 (N22106, N22019);
xor XOR2 (N22107, N22098, N4122);
nor NOR4 (N22108, N22104, N18838, N1225, N9776);
xor XOR2 (N22109, N22103, N7481);
nand NAND3 (N22110, N22107, N10804, N11268);
or OR2 (N22111, N22100, N2323);
nor NOR2 (N22112, N22108, N9362);
not NOT1 (N22113, N22105);
nor NOR3 (N22114, N22093, N12010, N21718);
nor NOR3 (N22115, N22113, N10302, N2726);
nand NAND4 (N22116, N22106, N4005, N20899, N12628);
not NOT1 (N22117, N22095);
not NOT1 (N22118, N22115);
nor NOR2 (N22119, N22110, N8798);
buf BUF1 (N22120, N22117);
nor NOR4 (N22121, N22099, N410, N9076, N1709);
nand NAND2 (N22122, N22114, N6233);
not NOT1 (N22123, N22118);
xor XOR2 (N22124, N22097, N3819);
buf BUF1 (N22125, N22109);
nor NOR4 (N22126, N22121, N7403, N10623, N14779);
and AND4 (N22127, N22120, N4081, N20743, N21442);
xor XOR2 (N22128, N22127, N3833);
xor XOR2 (N22129, N22128, N17040);
or OR4 (N22130, N22129, N16825, N8866, N5321);
not NOT1 (N22131, N22125);
and AND4 (N22132, N22126, N15812, N20022, N11041);
nand NAND3 (N22133, N22130, N5198, N20791);
and AND3 (N22134, N22123, N5912, N1836);
nand NAND3 (N22135, N22116, N16662, N16553);
and AND3 (N22136, N22133, N7600, N20093);
and AND4 (N22137, N22136, N13167, N8018, N13330);
and AND2 (N22138, N22119, N11242);
or OR3 (N22139, N22132, N7028, N5289);
nor NOR2 (N22140, N22138, N9501);
xor XOR2 (N22141, N22112, N4699);
buf BUF1 (N22142, N22140);
or OR4 (N22143, N22141, N8240, N8037, N10151);
xor XOR2 (N22144, N22143, N15657);
xor XOR2 (N22145, N22144, N4408);
buf BUF1 (N22146, N22142);
nand NAND2 (N22147, N22134, N15599);
or OR2 (N22148, N22137, N1025);
not NOT1 (N22149, N22111);
nand NAND3 (N22150, N22122, N14373, N9704);
nand NAND3 (N22151, N22139, N3050, N14508);
buf BUF1 (N22152, N22131);
xor XOR2 (N22153, N22146, N6982);
buf BUF1 (N22154, N22153);
nor NOR2 (N22155, N22135, N6207);
buf BUF1 (N22156, N22147);
and AND4 (N22157, N22155, N17796, N15719, N12125);
and AND2 (N22158, N22124, N7731);
nor NOR3 (N22159, N22158, N698, N4309);
not NOT1 (N22160, N22145);
or OR4 (N22161, N22151, N16120, N21418, N3726);
or OR4 (N22162, N22159, N12616, N12762, N18303);
or OR3 (N22163, N22150, N18030, N3098);
nand NAND4 (N22164, N22162, N877, N17328, N14790);
not NOT1 (N22165, N22164);
not NOT1 (N22166, N22148);
nor NOR4 (N22167, N22160, N9172, N16452, N6327);
or OR2 (N22168, N22167, N1426);
and AND2 (N22169, N22163, N21513);
or OR2 (N22170, N22154, N18307);
nand NAND2 (N22171, N22156, N18131);
not NOT1 (N22172, N22170);
xor XOR2 (N22173, N22149, N12368);
not NOT1 (N22174, N22172);
not NOT1 (N22175, N22171);
and AND4 (N22176, N22157, N2295, N1176, N14538);
and AND2 (N22177, N22169, N17838);
or OR4 (N22178, N22161, N18388, N12430, N7611);
and AND2 (N22179, N22175, N21881);
and AND2 (N22180, N22166, N7671);
and AND2 (N22181, N22178, N17388);
buf BUF1 (N22182, N22168);
xor XOR2 (N22183, N22179, N13406);
xor XOR2 (N22184, N22182, N2252);
not NOT1 (N22185, N22165);
nand NAND3 (N22186, N22177, N22014, N6602);
or OR3 (N22187, N22173, N11684, N1813);
not NOT1 (N22188, N22180);
and AND4 (N22189, N22187, N12688, N2575, N10170);
or OR2 (N22190, N22174, N10895);
xor XOR2 (N22191, N22176, N10005);
and AND4 (N22192, N22181, N8330, N1768, N520);
buf BUF1 (N22193, N22183);
buf BUF1 (N22194, N22185);
and AND2 (N22195, N22190, N15793);
xor XOR2 (N22196, N22192, N1132);
xor XOR2 (N22197, N22188, N11191);
not NOT1 (N22198, N22184);
not NOT1 (N22199, N22197);
nor NOR2 (N22200, N22196, N14245);
not NOT1 (N22201, N22195);
xor XOR2 (N22202, N22200, N11356);
and AND3 (N22203, N22191, N21635, N17946);
or OR2 (N22204, N22202, N4129);
xor XOR2 (N22205, N22203, N7418);
nand NAND4 (N22206, N22198, N16650, N19451, N11748);
buf BUF1 (N22207, N22193);
not NOT1 (N22208, N22152);
nand NAND2 (N22209, N22194, N2549);
nand NAND2 (N22210, N22209, N783);
not NOT1 (N22211, N22205);
xor XOR2 (N22212, N22204, N15354);
and AND3 (N22213, N22206, N9275, N19284);
and AND4 (N22214, N22212, N4349, N6359, N18755);
buf BUF1 (N22215, N22201);
nand NAND2 (N22216, N22189, N11306);
not NOT1 (N22217, N22199);
nand NAND3 (N22218, N22217, N1677, N280);
xor XOR2 (N22219, N22218, N16997);
buf BUF1 (N22220, N22208);
nor NOR4 (N22221, N22215, N13488, N12770, N10538);
not NOT1 (N22222, N22213);
and AND2 (N22223, N22214, N8096);
or OR3 (N22224, N22216, N18626, N13166);
nor NOR4 (N22225, N22221, N20467, N4589, N2833);
nand NAND3 (N22226, N22225, N1396, N482);
or OR4 (N22227, N22211, N1914, N754, N17147);
nand NAND3 (N22228, N22186, N3191, N9137);
nand NAND4 (N22229, N22223, N7189, N11607, N16076);
buf BUF1 (N22230, N22207);
not NOT1 (N22231, N22219);
and AND4 (N22232, N22229, N13980, N4788, N13014);
xor XOR2 (N22233, N22220, N8275);
not NOT1 (N22234, N22231);
and AND3 (N22235, N22210, N20447, N18010);
nor NOR2 (N22236, N22235, N11019);
and AND3 (N22237, N22236, N2844, N22167);
nor NOR3 (N22238, N22234, N8161, N21933);
and AND4 (N22239, N22232, N20756, N8197, N10095);
or OR3 (N22240, N22230, N12006, N21227);
buf BUF1 (N22241, N22227);
buf BUF1 (N22242, N22237);
nor NOR4 (N22243, N22240, N14829, N5118, N1667);
xor XOR2 (N22244, N22224, N16289);
buf BUF1 (N22245, N22233);
buf BUF1 (N22246, N22245);
and AND4 (N22247, N22226, N8867, N21578, N14268);
buf BUF1 (N22248, N22243);
nor NOR2 (N22249, N22246, N6904);
and AND2 (N22250, N22241, N8143);
not NOT1 (N22251, N22249);
buf BUF1 (N22252, N22251);
nor NOR3 (N22253, N22248, N2009, N8363);
nand NAND2 (N22254, N22238, N8287);
nand NAND3 (N22255, N22242, N14987, N9110);
xor XOR2 (N22256, N22255, N495);
buf BUF1 (N22257, N22239);
xor XOR2 (N22258, N22254, N16677);
nor NOR4 (N22259, N22252, N14480, N10087, N11274);
not NOT1 (N22260, N22259);
or OR3 (N22261, N22260, N1016, N3612);
xor XOR2 (N22262, N22258, N12200);
xor XOR2 (N22263, N22244, N11286);
and AND2 (N22264, N22247, N14601);
buf BUF1 (N22265, N22256);
buf BUF1 (N22266, N22264);
buf BUF1 (N22267, N22261);
xor XOR2 (N22268, N22263, N14427);
or OR2 (N22269, N22257, N21870);
nand NAND3 (N22270, N22228, N13461, N12673);
and AND3 (N22271, N22269, N20032, N7792);
or OR2 (N22272, N22268, N17604);
or OR4 (N22273, N22253, N21336, N21785, N532);
nand NAND2 (N22274, N22266, N21785);
or OR4 (N22275, N22272, N1406, N17549, N20627);
or OR3 (N22276, N22274, N17761, N654);
nor NOR4 (N22277, N22271, N12984, N12051, N5434);
nor NOR3 (N22278, N22267, N17288, N9444);
nor NOR4 (N22279, N22278, N10777, N21262, N17296);
buf BUF1 (N22280, N22250);
nor NOR2 (N22281, N22275, N15525);
not NOT1 (N22282, N22222);
nor NOR2 (N22283, N22273, N17888);
xor XOR2 (N22284, N22280, N9282);
not NOT1 (N22285, N22283);
buf BUF1 (N22286, N22285);
or OR3 (N22287, N22281, N2348, N18970);
xor XOR2 (N22288, N22279, N5030);
nor NOR2 (N22289, N22276, N18003);
or OR2 (N22290, N22286, N20202);
buf BUF1 (N22291, N22284);
xor XOR2 (N22292, N22291, N339);
or OR3 (N22293, N22288, N17801, N5726);
xor XOR2 (N22294, N22265, N18215);
nor NOR2 (N22295, N22282, N15305);
or OR3 (N22296, N22270, N7595, N18234);
nand NAND2 (N22297, N22262, N11072);
nor NOR3 (N22298, N22290, N9984, N13007);
buf BUF1 (N22299, N22295);
not NOT1 (N22300, N22293);
buf BUF1 (N22301, N22277);
nor NOR3 (N22302, N22301, N2611, N6027);
not NOT1 (N22303, N22300);
and AND2 (N22304, N22297, N21890);
and AND2 (N22305, N22298, N17927);
and AND2 (N22306, N22289, N21708);
xor XOR2 (N22307, N22287, N8361);
and AND2 (N22308, N22302, N8962);
xor XOR2 (N22309, N22294, N1825);
and AND3 (N22310, N22305, N11433, N20195);
and AND3 (N22311, N22310, N16761, N10721);
buf BUF1 (N22312, N22296);
and AND3 (N22313, N22299, N10487, N10970);
xor XOR2 (N22314, N22308, N3467);
and AND2 (N22315, N22311, N6551);
not NOT1 (N22316, N22307);
nand NAND3 (N22317, N22309, N15113, N20396);
buf BUF1 (N22318, N22313);
and AND3 (N22319, N22315, N16068, N5797);
xor XOR2 (N22320, N22312, N15525);
or OR2 (N22321, N22314, N21559);
or OR2 (N22322, N22321, N10340);
and AND4 (N22323, N22316, N848, N14923, N3083);
xor XOR2 (N22324, N22319, N13229);
or OR3 (N22325, N22306, N4963, N5665);
nand NAND2 (N22326, N22323, N7114);
buf BUF1 (N22327, N22303);
xor XOR2 (N22328, N22292, N4383);
or OR3 (N22329, N22318, N19603, N5865);
not NOT1 (N22330, N22325);
not NOT1 (N22331, N22322);
not NOT1 (N22332, N22326);
or OR2 (N22333, N22317, N5558);
nand NAND4 (N22334, N22329, N19446, N4802, N11379);
xor XOR2 (N22335, N22324, N19358);
not NOT1 (N22336, N22328);
not NOT1 (N22337, N22333);
or OR3 (N22338, N22304, N11477, N16281);
and AND4 (N22339, N22331, N15184, N11049, N5653);
nand NAND3 (N22340, N22337, N11527, N18208);
buf BUF1 (N22341, N22330);
and AND4 (N22342, N22332, N7069, N17520, N3825);
not NOT1 (N22343, N22336);
nor NOR4 (N22344, N22343, N9325, N3379, N17473);
and AND3 (N22345, N22327, N17639, N17548);
and AND3 (N22346, N22340, N13805, N11908);
buf BUF1 (N22347, N22341);
or OR3 (N22348, N22339, N10295, N15241);
and AND3 (N22349, N22346, N16873, N8872);
and AND2 (N22350, N22320, N84);
buf BUF1 (N22351, N22335);
not NOT1 (N22352, N22344);
and AND4 (N22353, N22334, N18315, N20460, N17804);
nand NAND3 (N22354, N22348, N17997, N2586);
and AND4 (N22355, N22354, N19687, N3217, N9594);
or OR3 (N22356, N22342, N276, N15626);
buf BUF1 (N22357, N22351);
or OR2 (N22358, N22338, N10276);
or OR2 (N22359, N22356, N2329);
and AND2 (N22360, N22358, N8207);
xor XOR2 (N22361, N22355, N10603);
xor XOR2 (N22362, N22352, N19715);
nor NOR4 (N22363, N22362, N7106, N21214, N5703);
and AND4 (N22364, N22363, N11635, N10030, N21267);
and AND3 (N22365, N22360, N6860, N11075);
nand NAND4 (N22366, N22349, N16523, N14709, N11791);
not NOT1 (N22367, N22364);
or OR4 (N22368, N22365, N12881, N9745, N7504);
or OR2 (N22369, N22368, N819);
and AND4 (N22370, N22367, N20193, N7338, N17611);
buf BUF1 (N22371, N22350);
nor NOR3 (N22372, N22370, N11996, N12219);
nor NOR2 (N22373, N22347, N11749);
nand NAND3 (N22374, N22353, N885, N1815);
or OR3 (N22375, N22372, N6463, N12073);
nor NOR2 (N22376, N22357, N7892);
nor NOR2 (N22377, N22374, N589);
nor NOR3 (N22378, N22366, N21919, N19297);
and AND2 (N22379, N22373, N20778);
buf BUF1 (N22380, N22369);
xor XOR2 (N22381, N22371, N18761);
nor NOR2 (N22382, N22381, N9423);
xor XOR2 (N22383, N22379, N20702);
xor XOR2 (N22384, N22382, N2020);
xor XOR2 (N22385, N22384, N19563);
nor NOR3 (N22386, N22359, N17361, N13784);
xor XOR2 (N22387, N22378, N1344);
buf BUF1 (N22388, N22375);
and AND3 (N22389, N22388, N2571, N9331);
buf BUF1 (N22390, N22376);
or OR4 (N22391, N22377, N20732, N19358, N15297);
not NOT1 (N22392, N22387);
and AND2 (N22393, N22386, N1941);
and AND4 (N22394, N22361, N17569, N14520, N7911);
or OR2 (N22395, N22390, N19053);
buf BUF1 (N22396, N22393);
nand NAND3 (N22397, N22345, N12292, N1944);
buf BUF1 (N22398, N22391);
nand NAND4 (N22399, N22397, N2491, N8431, N8379);
and AND3 (N22400, N22383, N11972, N7281);
and AND2 (N22401, N22395, N6662);
or OR4 (N22402, N22389, N16143, N6874, N19652);
and AND3 (N22403, N22396, N21985, N17093);
xor XOR2 (N22404, N22398, N13904);
nand NAND3 (N22405, N22385, N11226, N250);
nor NOR2 (N22406, N22399, N16016);
nand NAND3 (N22407, N22392, N17094, N15675);
or OR2 (N22408, N22407, N10975);
nand NAND4 (N22409, N22404, N16639, N14769, N2375);
not NOT1 (N22410, N22405);
nand NAND4 (N22411, N22402, N11658, N521, N21638);
or OR3 (N22412, N22400, N21271, N9436);
xor XOR2 (N22413, N22403, N267);
buf BUF1 (N22414, N22394);
not NOT1 (N22415, N22406);
and AND2 (N22416, N22410, N9595);
and AND2 (N22417, N22411, N17548);
not NOT1 (N22418, N22408);
or OR2 (N22419, N22412, N21341);
nand NAND3 (N22420, N22417, N17679, N6183);
xor XOR2 (N22421, N22380, N15292);
xor XOR2 (N22422, N22420, N9902);
buf BUF1 (N22423, N22415);
nand NAND2 (N22424, N22409, N20042);
or OR4 (N22425, N22422, N13876, N11771, N15145);
nand NAND2 (N22426, N22425, N16021);
and AND3 (N22427, N22413, N7463, N14961);
buf BUF1 (N22428, N22418);
and AND2 (N22429, N22427, N9893);
nor NOR2 (N22430, N22416, N17846);
or OR4 (N22431, N22419, N13420, N17682, N22291);
not NOT1 (N22432, N22401);
nor NOR2 (N22433, N22429, N3469);
not NOT1 (N22434, N22430);
not NOT1 (N22435, N22433);
nand NAND4 (N22436, N22435, N5499, N18625, N12054);
buf BUF1 (N22437, N22426);
nor NOR4 (N22438, N22414, N2871, N2511, N10589);
not NOT1 (N22439, N22437);
and AND3 (N22440, N22439, N1649, N2515);
not NOT1 (N22441, N22432);
or OR2 (N22442, N22434, N1586);
buf BUF1 (N22443, N22428);
xor XOR2 (N22444, N22438, N3326);
nand NAND2 (N22445, N22423, N12504);
nor NOR4 (N22446, N22424, N11146, N81, N8925);
not NOT1 (N22447, N22446);
buf BUF1 (N22448, N22421);
xor XOR2 (N22449, N22443, N6463);
not NOT1 (N22450, N22436);
not NOT1 (N22451, N22431);
not NOT1 (N22452, N22450);
nand NAND2 (N22453, N22449, N10008);
or OR3 (N22454, N22448, N22273, N14620);
xor XOR2 (N22455, N22444, N15313);
nor NOR2 (N22456, N22447, N4495);
not NOT1 (N22457, N22452);
or OR2 (N22458, N22451, N5140);
nand NAND3 (N22459, N22440, N21183, N18612);
nor NOR3 (N22460, N22456, N22291, N12519);
not NOT1 (N22461, N22459);
not NOT1 (N22462, N22457);
and AND2 (N22463, N22454, N12281);
and AND3 (N22464, N22445, N7370, N21104);
not NOT1 (N22465, N22458);
not NOT1 (N22466, N22460);
buf BUF1 (N22467, N22464);
nand NAND2 (N22468, N22461, N13552);
and AND3 (N22469, N22442, N20555, N12620);
and AND2 (N22470, N22466, N11540);
or OR3 (N22471, N22470, N10840, N9864);
nand NAND4 (N22472, N22467, N12987, N2305, N11400);
buf BUF1 (N22473, N22463);
nand NAND2 (N22474, N22471, N18901);
or OR4 (N22475, N22441, N7290, N7961, N5996);
xor XOR2 (N22476, N22465, N10042);
and AND3 (N22477, N22473, N425, N3673);
or OR2 (N22478, N22455, N6428);
and AND4 (N22479, N22474, N7594, N8428, N12617);
and AND2 (N22480, N22477, N12321);
and AND2 (N22481, N22472, N4120);
and AND4 (N22482, N22462, N470, N2847, N17444);
or OR2 (N22483, N22468, N653);
nor NOR3 (N22484, N22483, N19173, N22381);
or OR3 (N22485, N22484, N10411, N12156);
or OR2 (N22486, N22481, N10642);
nand NAND4 (N22487, N22453, N10565, N4546, N13494);
or OR4 (N22488, N22486, N6315, N13883, N3772);
nor NOR2 (N22489, N22482, N13890);
and AND3 (N22490, N22487, N6525, N11227);
buf BUF1 (N22491, N22476);
xor XOR2 (N22492, N22488, N18980);
or OR3 (N22493, N22469, N19583, N10634);
xor XOR2 (N22494, N22491, N19821);
buf BUF1 (N22495, N22475);
and AND4 (N22496, N22490, N12157, N15296, N17595);
not NOT1 (N22497, N22478);
and AND4 (N22498, N22489, N8014, N2853, N5912);
nand NAND2 (N22499, N22496, N94);
nand NAND3 (N22500, N22494, N13132, N19777);
or OR2 (N22501, N22497, N16014);
nand NAND2 (N22502, N22485, N3835);
xor XOR2 (N22503, N22492, N20225);
nor NOR4 (N22504, N22501, N8662, N16437, N20376);
or OR4 (N22505, N22498, N1300, N11543, N16379);
or OR2 (N22506, N22493, N471);
buf BUF1 (N22507, N22504);
or OR4 (N22508, N22506, N21757, N19738, N4844);
buf BUF1 (N22509, N22508);
and AND4 (N22510, N22507, N13886, N19675, N19342);
nor NOR2 (N22511, N22502, N4689);
or OR3 (N22512, N22499, N1638, N9319);
nand NAND2 (N22513, N22495, N20954);
and AND2 (N22514, N22500, N17833);
nor NOR4 (N22515, N22512, N2125, N6845, N5500);
nand NAND2 (N22516, N22505, N6421);
xor XOR2 (N22517, N22515, N16417);
nand NAND4 (N22518, N22480, N21554, N17986, N2742);
and AND4 (N22519, N22503, N21389, N14774, N15042);
xor XOR2 (N22520, N22510, N21301);
nor NOR2 (N22521, N22518, N15869);
buf BUF1 (N22522, N22511);
nand NAND3 (N22523, N22520, N12559, N17318);
xor XOR2 (N22524, N22522, N3259);
nand NAND2 (N22525, N22516, N826);
nor NOR2 (N22526, N22525, N18755);
nand NAND4 (N22527, N22514, N20425, N4497, N10886);
not NOT1 (N22528, N22524);
xor XOR2 (N22529, N22521, N5771);
xor XOR2 (N22530, N22529, N1348);
buf BUF1 (N22531, N22530);
not NOT1 (N22532, N22509);
nand NAND3 (N22533, N22519, N20348, N6009);
nand NAND2 (N22534, N22531, N14663);
xor XOR2 (N22535, N22513, N21308);
nor NOR4 (N22536, N22533, N13056, N21109, N6478);
and AND2 (N22537, N22536, N12852);
nor NOR2 (N22538, N22532, N22118);
or OR4 (N22539, N22537, N6890, N21592, N3895);
or OR3 (N22540, N22527, N16137, N5945);
nand NAND3 (N22541, N22539, N2243, N10376);
and AND2 (N22542, N22540, N2642);
or OR2 (N22543, N22535, N13720);
xor XOR2 (N22544, N22479, N14038);
buf BUF1 (N22545, N22523);
nor NOR2 (N22546, N22545, N8438);
and AND4 (N22547, N22538, N10748, N21426, N11850);
or OR4 (N22548, N22541, N17624, N17669, N6592);
or OR2 (N22549, N22534, N15029);
nand NAND2 (N22550, N22544, N14499);
xor XOR2 (N22551, N22548, N1035);
nor NOR2 (N22552, N22528, N22240);
and AND3 (N22553, N22549, N18680, N11684);
or OR3 (N22554, N22553, N18546, N20302);
buf BUF1 (N22555, N22543);
xor XOR2 (N22556, N22542, N18591);
and AND4 (N22557, N22547, N20526, N977, N6584);
nand NAND4 (N22558, N22551, N7582, N2344, N20435);
nor NOR3 (N22559, N22552, N17936, N12725);
nor NOR4 (N22560, N22555, N13562, N2848, N6079);
or OR4 (N22561, N22556, N3295, N11583, N6748);
or OR3 (N22562, N22561, N19707, N10668);
xor XOR2 (N22563, N22558, N8247);
buf BUF1 (N22564, N22550);
buf BUF1 (N22565, N22564);
xor XOR2 (N22566, N22554, N372);
nor NOR4 (N22567, N22557, N13335, N7442, N6097);
not NOT1 (N22568, N22559);
and AND2 (N22569, N22568, N22371);
buf BUF1 (N22570, N22562);
not NOT1 (N22571, N22567);
buf BUF1 (N22572, N22517);
nand NAND4 (N22573, N22570, N4407, N21846, N22328);
nand NAND4 (N22574, N22569, N4033, N865, N10304);
nor NOR2 (N22575, N22565, N10642);
or OR4 (N22576, N22575, N15751, N14529, N1420);
nand NAND2 (N22577, N22546, N7762);
buf BUF1 (N22578, N22526);
and AND4 (N22579, N22563, N21164, N7482, N18916);
not NOT1 (N22580, N22578);
or OR4 (N22581, N22571, N18931, N15797, N19401);
not NOT1 (N22582, N22560);
not NOT1 (N22583, N22581);
not NOT1 (N22584, N22574);
nand NAND4 (N22585, N22577, N19533, N13653, N1047);
buf BUF1 (N22586, N22582);
and AND2 (N22587, N22566, N5271);
nor NOR3 (N22588, N22572, N6766, N14726);
nor NOR4 (N22589, N22586, N21648, N22524, N3416);
or OR3 (N22590, N22587, N7392, N9094);
or OR2 (N22591, N22589, N12033);
or OR4 (N22592, N22579, N14574, N15409, N1423);
xor XOR2 (N22593, N22580, N19310);
or OR3 (N22594, N22576, N3392, N12228);
buf BUF1 (N22595, N22583);
or OR2 (N22596, N22584, N7581);
not NOT1 (N22597, N22594);
buf BUF1 (N22598, N22590);
not NOT1 (N22599, N22588);
not NOT1 (N22600, N22573);
buf BUF1 (N22601, N22591);
xor XOR2 (N22602, N22601, N14064);
not NOT1 (N22603, N22600);
xor XOR2 (N22604, N22596, N11035);
not NOT1 (N22605, N22598);
nand NAND2 (N22606, N22603, N19748);
nor NOR3 (N22607, N22585, N6779, N13488);
nor NOR4 (N22608, N22599, N8213, N13692, N14450);
nor NOR3 (N22609, N22605, N20165, N21196);
nand NAND2 (N22610, N22592, N19808);
and AND4 (N22611, N22609, N5163, N12343, N18099);
and AND3 (N22612, N22604, N291, N20719);
and AND2 (N22613, N22593, N20219);
buf BUF1 (N22614, N22597);
nand NAND2 (N22615, N22608, N19400);
or OR4 (N22616, N22595, N20945, N13031, N7406);
nor NOR4 (N22617, N22614, N3723, N13040, N19216);
not NOT1 (N22618, N22607);
nor NOR4 (N22619, N22613, N16116, N20586, N3762);
and AND2 (N22620, N22611, N7941);
nand NAND4 (N22621, N22615, N1557, N9266, N18991);
not NOT1 (N22622, N22616);
and AND2 (N22623, N22619, N14969);
not NOT1 (N22624, N22618);
nor NOR3 (N22625, N22617, N2705, N854);
nand NAND2 (N22626, N22612, N20799);
not NOT1 (N22627, N22610);
not NOT1 (N22628, N22621);
or OR3 (N22629, N22606, N11185, N7195);
or OR3 (N22630, N22622, N17389, N21941);
not NOT1 (N22631, N22602);
buf BUF1 (N22632, N22625);
nor NOR4 (N22633, N22627, N5991, N18054, N8675);
buf BUF1 (N22634, N22628);
and AND2 (N22635, N22632, N15475);
not NOT1 (N22636, N22633);
buf BUF1 (N22637, N22635);
or OR3 (N22638, N22629, N13892, N1783);
not NOT1 (N22639, N22620);
buf BUF1 (N22640, N22626);
not NOT1 (N22641, N22636);
nand NAND3 (N22642, N22623, N6581, N4648);
and AND2 (N22643, N22624, N20975);
buf BUF1 (N22644, N22640);
nor NOR3 (N22645, N22630, N2438, N8687);
buf BUF1 (N22646, N22634);
or OR3 (N22647, N22645, N18749, N9032);
nor NOR2 (N22648, N22637, N2410);
nor NOR4 (N22649, N22638, N10624, N1012, N11311);
nand NAND3 (N22650, N22631, N567, N19552);
buf BUF1 (N22651, N22643);
nand NAND3 (N22652, N22644, N8344, N1262);
buf BUF1 (N22653, N22652);
buf BUF1 (N22654, N22649);
not NOT1 (N22655, N22653);
or OR3 (N22656, N22647, N6618, N13090);
and AND3 (N22657, N22651, N9915, N16377);
xor XOR2 (N22658, N22650, N12797);
xor XOR2 (N22659, N22639, N7629);
buf BUF1 (N22660, N22646);
or OR2 (N22661, N22648, N11563);
not NOT1 (N22662, N22661);
buf BUF1 (N22663, N22656);
nand NAND4 (N22664, N22660, N6554, N5537, N3231);
xor XOR2 (N22665, N22664, N17009);
and AND3 (N22666, N22655, N22099, N1085);
nand NAND4 (N22667, N22663, N3242, N20599, N6294);
buf BUF1 (N22668, N22641);
xor XOR2 (N22669, N22665, N1344);
buf BUF1 (N22670, N22668);
buf BUF1 (N22671, N22662);
xor XOR2 (N22672, N22670, N2607);
nand NAND3 (N22673, N22654, N7729, N8823);
nor NOR4 (N22674, N22642, N21413, N7436, N227);
not NOT1 (N22675, N22666);
and AND4 (N22676, N22658, N7588, N6189, N19883);
nand NAND4 (N22677, N22675, N1559, N17703, N6081);
not NOT1 (N22678, N22659);
nor NOR3 (N22679, N22657, N5838, N15539);
and AND2 (N22680, N22669, N20282);
nor NOR2 (N22681, N22673, N11003);
xor XOR2 (N22682, N22676, N12597);
not NOT1 (N22683, N22674);
buf BUF1 (N22684, N22680);
nor NOR2 (N22685, N22684, N21925);
not NOT1 (N22686, N22683);
or OR3 (N22687, N22671, N7858, N16527);
or OR2 (N22688, N22678, N21274);
nand NAND2 (N22689, N22667, N3726);
nor NOR4 (N22690, N22689, N8599, N977, N21961);
not NOT1 (N22691, N22677);
xor XOR2 (N22692, N22681, N22501);
and AND3 (N22693, N22672, N17891, N7352);
nor NOR3 (N22694, N22693, N12363, N12735);
or OR2 (N22695, N22679, N10623);
nand NAND4 (N22696, N22690, N15209, N20958, N6156);
buf BUF1 (N22697, N22694);
buf BUF1 (N22698, N22696);
nand NAND3 (N22699, N22698, N4827, N17283);
nor NOR4 (N22700, N22699, N9335, N4696, N6251);
nand NAND3 (N22701, N22688, N14903, N7220);
buf BUF1 (N22702, N22685);
nor NOR4 (N22703, N22686, N16872, N9807, N21615);
not NOT1 (N22704, N22695);
nand NAND2 (N22705, N22687, N16178);
nor NOR2 (N22706, N22702, N4957);
nand NAND3 (N22707, N22691, N5243, N6889);
buf BUF1 (N22708, N22700);
xor XOR2 (N22709, N22692, N11108);
nor NOR3 (N22710, N22707, N9416, N9328);
or OR4 (N22711, N22682, N15512, N10628, N2798);
and AND3 (N22712, N22708, N8485, N4840);
nand NAND3 (N22713, N22711, N11351, N5169);
or OR3 (N22714, N22701, N21582, N10123);
and AND3 (N22715, N22704, N16982, N13703);
xor XOR2 (N22716, N22712, N10104);
nor NOR4 (N22717, N22706, N15287, N17877, N13462);
not NOT1 (N22718, N22714);
not NOT1 (N22719, N22715);
buf BUF1 (N22720, N22697);
buf BUF1 (N22721, N22710);
nor NOR2 (N22722, N22721, N248);
nor NOR4 (N22723, N22716, N20732, N19552, N5632);
xor XOR2 (N22724, N22723, N21848);
or OR2 (N22725, N22719, N3681);
nand NAND3 (N22726, N22725, N18978, N8445);
and AND2 (N22727, N22709, N16224);
or OR2 (N22728, N22718, N21550);
nor NOR3 (N22729, N22720, N13729, N2315);
buf BUF1 (N22730, N22729);
buf BUF1 (N22731, N22728);
nand NAND3 (N22732, N22731, N4188, N1006);
xor XOR2 (N22733, N22726, N6293);
nand NAND2 (N22734, N22724, N17734);
and AND4 (N22735, N22733, N19888, N4663, N17472);
nor NOR2 (N22736, N22732, N12560);
nand NAND3 (N22737, N22734, N13052, N20850);
not NOT1 (N22738, N22717);
nor NOR2 (N22739, N22722, N17932);
or OR4 (N22740, N22727, N1080, N18493, N2920);
and AND2 (N22741, N22739, N4814);
xor XOR2 (N22742, N22713, N5092);
buf BUF1 (N22743, N22737);
nand NAND3 (N22744, N22740, N20746, N1823);
and AND3 (N22745, N22730, N10119, N4546);
nor NOR4 (N22746, N22735, N14011, N18072, N12884);
nand NAND3 (N22747, N22738, N8970, N11103);
nor NOR3 (N22748, N22743, N8651, N21475);
and AND4 (N22749, N22736, N11458, N15114, N2612);
or OR2 (N22750, N22703, N10541);
buf BUF1 (N22751, N22744);
xor XOR2 (N22752, N22742, N9340);
xor XOR2 (N22753, N22705, N19804);
nand NAND3 (N22754, N22750, N17227, N8165);
buf BUF1 (N22755, N22747);
nor NOR3 (N22756, N22753, N15794, N6207);
or OR2 (N22757, N22751, N1775);
or OR3 (N22758, N22748, N20535, N10174);
nor NOR4 (N22759, N22756, N4996, N18841, N20992);
and AND2 (N22760, N22757, N15156);
buf BUF1 (N22761, N22760);
and AND4 (N22762, N22755, N21439, N14673, N14633);
nand NAND2 (N22763, N22746, N11588);
nor NOR3 (N22764, N22762, N20235, N9453);
buf BUF1 (N22765, N22754);
and AND4 (N22766, N22745, N271, N16921, N1261);
nor NOR3 (N22767, N22749, N10357, N8071);
not NOT1 (N22768, N22741);
nor NOR3 (N22769, N22765, N5542, N17494);
not NOT1 (N22770, N22769);
not NOT1 (N22771, N22763);
xor XOR2 (N22772, N22767, N2681);
nand NAND2 (N22773, N22770, N1851);
buf BUF1 (N22774, N22771);
buf BUF1 (N22775, N22772);
not NOT1 (N22776, N22766);
not NOT1 (N22777, N22759);
not NOT1 (N22778, N22761);
and AND3 (N22779, N22752, N12894, N882);
and AND4 (N22780, N22779, N22472, N14887, N1140);
and AND2 (N22781, N22778, N1613);
buf BUF1 (N22782, N22774);
nand NAND3 (N22783, N22777, N8535, N1989);
buf BUF1 (N22784, N22764);
or OR3 (N22785, N22781, N17305, N17342);
and AND3 (N22786, N22783, N22255, N18516);
xor XOR2 (N22787, N22780, N2105);
or OR4 (N22788, N22773, N10546, N15882, N17994);
nand NAND4 (N22789, N22787, N6285, N11930, N9725);
and AND4 (N22790, N22785, N12762, N8543, N20076);
nand NAND2 (N22791, N22782, N15778);
nand NAND2 (N22792, N22791, N10444);
or OR3 (N22793, N22792, N7215, N11644);
not NOT1 (N22794, N22786);
nand NAND2 (N22795, N22793, N7250);
or OR3 (N22796, N22788, N18087, N5912);
not NOT1 (N22797, N22775);
not NOT1 (N22798, N22794);
nor NOR2 (N22799, N22758, N4095);
nor NOR4 (N22800, N22796, N10792, N8008, N7399);
not NOT1 (N22801, N22789);
xor XOR2 (N22802, N22799, N16562);
and AND4 (N22803, N22784, N2851, N4251, N7201);
and AND2 (N22804, N22802, N17801);
nand NAND3 (N22805, N22800, N19132, N11342);
not NOT1 (N22806, N22801);
xor XOR2 (N22807, N22776, N11919);
nand NAND4 (N22808, N22806, N13970, N9745, N19252);
or OR3 (N22809, N22807, N137, N12151);
nand NAND4 (N22810, N22798, N9332, N19268, N9249);
not NOT1 (N22811, N22805);
xor XOR2 (N22812, N22804, N11397);
and AND4 (N22813, N22790, N10796, N3477, N1494);
xor XOR2 (N22814, N22812, N7127);
not NOT1 (N22815, N22810);
nor NOR3 (N22816, N22811, N174, N18939);
or OR2 (N22817, N22797, N18697);
nor NOR3 (N22818, N22803, N4520, N17186);
or OR2 (N22819, N22813, N9330);
nor NOR2 (N22820, N22818, N18143);
and AND2 (N22821, N22768, N4574);
or OR4 (N22822, N22814, N13807, N2661, N8508);
and AND3 (N22823, N22821, N9558, N16481);
buf BUF1 (N22824, N22817);
buf BUF1 (N22825, N22819);
nor NOR4 (N22826, N22822, N5945, N6794, N960);
xor XOR2 (N22827, N22826, N19002);
not NOT1 (N22828, N22815);
nor NOR4 (N22829, N22808, N5592, N20104, N1600);
xor XOR2 (N22830, N22816, N18746);
or OR2 (N22831, N22828, N738);
nor NOR2 (N22832, N22825, N19261);
and AND3 (N22833, N22827, N16717, N16966);
or OR2 (N22834, N22824, N12056);
nand NAND4 (N22835, N22831, N21040, N10330, N22073);
or OR2 (N22836, N22795, N22543);
buf BUF1 (N22837, N22829);
and AND2 (N22838, N22835, N7364);
and AND4 (N22839, N22820, N724, N11082, N16038);
xor XOR2 (N22840, N22823, N5237);
or OR2 (N22841, N22836, N3552);
nand NAND4 (N22842, N22839, N3924, N4412, N5312);
buf BUF1 (N22843, N22832);
xor XOR2 (N22844, N22842, N5484);
and AND3 (N22845, N22834, N3468, N19150);
not NOT1 (N22846, N22844);
buf BUF1 (N22847, N22846);
buf BUF1 (N22848, N22841);
and AND4 (N22849, N22840, N12528, N15488, N21706);
nor NOR4 (N22850, N22843, N18531, N10919, N13259);
xor XOR2 (N22851, N22837, N11753);
nor NOR2 (N22852, N22845, N7320);
or OR3 (N22853, N22852, N9977, N17814);
buf BUF1 (N22854, N22809);
nand NAND2 (N22855, N22847, N19978);
and AND2 (N22856, N22850, N4178);
nor NOR4 (N22857, N22848, N2569, N7540, N2242);
buf BUF1 (N22858, N22849);
xor XOR2 (N22859, N22856, N14047);
not NOT1 (N22860, N22855);
or OR3 (N22861, N22830, N13134, N15327);
not NOT1 (N22862, N22857);
and AND2 (N22863, N22861, N13411);
buf BUF1 (N22864, N22853);
or OR4 (N22865, N22862, N10422, N2978, N18431);
nor NOR3 (N22866, N22859, N15377, N1573);
buf BUF1 (N22867, N22860);
nor NOR4 (N22868, N22866, N10084, N21413, N3537);
not NOT1 (N22869, N22833);
xor XOR2 (N22870, N22865, N4026);
nor NOR3 (N22871, N22867, N14708, N17684);
nor NOR2 (N22872, N22871, N18567);
or OR3 (N22873, N22868, N9818, N4704);
buf BUF1 (N22874, N22838);
nand NAND3 (N22875, N22873, N12261, N16523);
nor NOR3 (N22876, N22863, N17563, N15905);
xor XOR2 (N22877, N22872, N11208);
xor XOR2 (N22878, N22869, N17501);
and AND2 (N22879, N22878, N3570);
nand NAND2 (N22880, N22879, N12205);
xor XOR2 (N22881, N22874, N5191);
xor XOR2 (N22882, N22876, N2584);
not NOT1 (N22883, N22881);
xor XOR2 (N22884, N22854, N16250);
or OR2 (N22885, N22858, N3116);
xor XOR2 (N22886, N22851, N19107);
and AND3 (N22887, N22884, N5595, N22244);
nor NOR3 (N22888, N22886, N5593, N1744);
nand NAND4 (N22889, N22882, N2370, N21721, N5451);
nor NOR2 (N22890, N22883, N6638);
and AND3 (N22891, N22880, N13286, N8344);
not NOT1 (N22892, N22891);
nor NOR2 (N22893, N22887, N3180);
nor NOR2 (N22894, N22875, N21564);
buf BUF1 (N22895, N22889);
xor XOR2 (N22896, N22892, N803);
nor NOR2 (N22897, N22890, N1351);
xor XOR2 (N22898, N22896, N11830);
buf BUF1 (N22899, N22897);
and AND4 (N22900, N22894, N10792, N1841, N6106);
not NOT1 (N22901, N22899);
buf BUF1 (N22902, N22893);
buf BUF1 (N22903, N22900);
not NOT1 (N22904, N22885);
buf BUF1 (N22905, N22898);
not NOT1 (N22906, N22903);
nor NOR4 (N22907, N22906, N7461, N18272, N20918);
not NOT1 (N22908, N22888);
xor XOR2 (N22909, N22870, N1137);
nor NOR4 (N22910, N22877, N16899, N823, N22267);
and AND2 (N22911, N22864, N11897);
buf BUF1 (N22912, N22904);
nand NAND3 (N22913, N22911, N21738, N19109);
nand NAND3 (N22914, N22895, N22712, N884);
not NOT1 (N22915, N22914);
buf BUF1 (N22916, N22910);
not NOT1 (N22917, N22916);
or OR4 (N22918, N22902, N14141, N2241, N1318);
not NOT1 (N22919, N22907);
and AND3 (N22920, N22912, N12991, N9880);
not NOT1 (N22921, N22919);
buf BUF1 (N22922, N22915);
nand NAND3 (N22923, N22922, N16157, N12283);
not NOT1 (N22924, N22909);
buf BUF1 (N22925, N22905);
not NOT1 (N22926, N22908);
and AND3 (N22927, N22921, N3128, N16317);
and AND2 (N22928, N22927, N2572);
buf BUF1 (N22929, N22923);
not NOT1 (N22930, N22918);
not NOT1 (N22931, N22924);
buf BUF1 (N22932, N22925);
nor NOR4 (N22933, N22932, N8918, N10040, N22329);
not NOT1 (N22934, N22930);
xor XOR2 (N22935, N22926, N11386);
and AND3 (N22936, N22917, N4405, N21525);
nor NOR3 (N22937, N22934, N10972, N3410);
xor XOR2 (N22938, N22937, N5261);
nor NOR3 (N22939, N22931, N612, N9249);
not NOT1 (N22940, N22913);
xor XOR2 (N22941, N22938, N18688);
xor XOR2 (N22942, N22940, N15340);
not NOT1 (N22943, N22935);
nor NOR2 (N22944, N22939, N20844);
or OR2 (N22945, N22941, N12517);
buf BUF1 (N22946, N22929);
nand NAND2 (N22947, N22928, N1158);
and AND3 (N22948, N22945, N10263, N17181);
buf BUF1 (N22949, N22943);
xor XOR2 (N22950, N22947, N1944);
buf BUF1 (N22951, N22950);
and AND2 (N22952, N22936, N17817);
buf BUF1 (N22953, N22942);
xor XOR2 (N22954, N22901, N21417);
not NOT1 (N22955, N22948);
buf BUF1 (N22956, N22955);
buf BUF1 (N22957, N22956);
nand NAND3 (N22958, N22920, N11447, N3177);
not NOT1 (N22959, N22958);
or OR3 (N22960, N22952, N920, N19700);
xor XOR2 (N22961, N22959, N9244);
buf BUF1 (N22962, N22946);
or OR2 (N22963, N22962, N8238);
and AND2 (N22964, N22944, N6121);
nor NOR2 (N22965, N22949, N18614);
nor NOR3 (N22966, N22954, N11283, N14836);
not NOT1 (N22967, N22951);
nand NAND4 (N22968, N22961, N6253, N13101, N3946);
and AND4 (N22969, N22960, N16116, N16599, N14134);
and AND3 (N22970, N22933, N3935, N17289);
buf BUF1 (N22971, N22969);
or OR4 (N22972, N22968, N18667, N5011, N14326);
buf BUF1 (N22973, N22965);
and AND3 (N22974, N22966, N6941, N15061);
not NOT1 (N22975, N22953);
not NOT1 (N22976, N22972);
buf BUF1 (N22977, N22975);
xor XOR2 (N22978, N22964, N12310);
nand NAND4 (N22979, N22973, N1463, N19965, N4949);
nor NOR4 (N22980, N22967, N4807, N13092, N7335);
buf BUF1 (N22981, N22979);
or OR4 (N22982, N22980, N12569, N8107, N19884);
nand NAND2 (N22983, N22974, N6251);
or OR3 (N22984, N22976, N19118, N22717);
buf BUF1 (N22985, N22981);
buf BUF1 (N22986, N22984);
or OR4 (N22987, N22971, N15429, N2089, N21002);
or OR2 (N22988, N22983, N20753);
nor NOR3 (N22989, N22977, N8074, N5699);
buf BUF1 (N22990, N22985);
and AND4 (N22991, N22989, N15872, N3882, N14996);
nor NOR2 (N22992, N22987, N18870);
buf BUF1 (N22993, N22957);
xor XOR2 (N22994, N22963, N18952);
buf BUF1 (N22995, N22970);
and AND4 (N22996, N22995, N374, N1923, N8094);
nor NOR2 (N22997, N22986, N916);
xor XOR2 (N22998, N22997, N1352);
xor XOR2 (N22999, N22991, N19963);
and AND3 (N23000, N22998, N1496, N9484);
or OR4 (N23001, N22990, N7158, N4048, N21130);
nor NOR4 (N23002, N22993, N17971, N13170, N12583);
buf BUF1 (N23003, N22988);
xor XOR2 (N23004, N22996, N12910);
and AND4 (N23005, N22994, N22184, N16347, N13853);
nor NOR4 (N23006, N23004, N16049, N10191, N449);
nand NAND3 (N23007, N22999, N4648, N12281);
nand NAND4 (N23008, N22978, N18327, N3525, N3054);
nor NOR4 (N23009, N23005, N6969, N19057, N21996);
and AND2 (N23010, N22992, N5451);
xor XOR2 (N23011, N23002, N10164);
nand NAND4 (N23012, N22982, N15302, N15882, N18278);
nand NAND2 (N23013, N23001, N3269);
nor NOR2 (N23014, N23008, N3546);
nand NAND2 (N23015, N23006, N17433);
and AND2 (N23016, N23011, N21732);
buf BUF1 (N23017, N23013);
or OR2 (N23018, N23010, N17377);
buf BUF1 (N23019, N23000);
and AND4 (N23020, N23019, N13814, N17452, N18657);
xor XOR2 (N23021, N23018, N3315);
xor XOR2 (N23022, N23012, N17329);
and AND2 (N23023, N23015, N6985);
xor XOR2 (N23024, N23003, N22874);
and AND3 (N23025, N23023, N4746, N20156);
xor XOR2 (N23026, N23022, N11335);
not NOT1 (N23027, N23007);
xor XOR2 (N23028, N23027, N20529);
nand NAND3 (N23029, N23014, N6689, N19325);
nor NOR4 (N23030, N23029, N8382, N19298, N1148);
nor NOR2 (N23031, N23021, N2461);
not NOT1 (N23032, N23028);
buf BUF1 (N23033, N23009);
nand NAND3 (N23034, N23016, N6225, N10551);
and AND3 (N23035, N23030, N15663, N17723);
and AND3 (N23036, N23032, N16074, N19704);
nand NAND3 (N23037, N23034, N5752, N1984);
buf BUF1 (N23038, N23017);
buf BUF1 (N23039, N23031);
buf BUF1 (N23040, N23026);
not NOT1 (N23041, N23025);
nor NOR4 (N23042, N23038, N1035, N668, N18608);
not NOT1 (N23043, N23042);
xor XOR2 (N23044, N23035, N11836);
nand NAND2 (N23045, N23043, N12000);
and AND2 (N23046, N23040, N16035);
nand NAND3 (N23047, N23045, N22906, N4671);
nor NOR4 (N23048, N23024, N1409, N10639, N5455);
xor XOR2 (N23049, N23037, N22515);
nor NOR3 (N23050, N23036, N8116, N22152);
or OR2 (N23051, N23046, N18250);
buf BUF1 (N23052, N23048);
xor XOR2 (N23053, N23041, N20326);
buf BUF1 (N23054, N23051);
nand NAND3 (N23055, N23049, N14534, N613);
nand NAND4 (N23056, N23050, N2163, N14401, N19843);
buf BUF1 (N23057, N23055);
and AND3 (N23058, N23052, N14780, N9162);
nor NOR3 (N23059, N23058, N22868, N10142);
nand NAND4 (N23060, N23053, N1624, N13578, N13775);
and AND4 (N23061, N23060, N7175, N22331, N10649);
or OR2 (N23062, N23033, N15402);
not NOT1 (N23063, N23059);
not NOT1 (N23064, N23044);
not NOT1 (N23065, N23057);
buf BUF1 (N23066, N23061);
buf BUF1 (N23067, N23054);
xor XOR2 (N23068, N23062, N11302);
xor XOR2 (N23069, N23047, N8173);
nand NAND4 (N23070, N23063, N15860, N18797, N10860);
buf BUF1 (N23071, N23065);
xor XOR2 (N23072, N23070, N16254);
nor NOR2 (N23073, N23066, N15785);
xor XOR2 (N23074, N23020, N916);
and AND3 (N23075, N23064, N15553, N20607);
or OR4 (N23076, N23039, N8286, N17468, N5656);
nand NAND4 (N23077, N23071, N15184, N5375, N20792);
buf BUF1 (N23078, N23056);
and AND4 (N23079, N23067, N12650, N4965, N6646);
not NOT1 (N23080, N23078);
nand NAND4 (N23081, N23068, N554, N17643, N20332);
xor XOR2 (N23082, N23069, N790);
not NOT1 (N23083, N23082);
not NOT1 (N23084, N23073);
buf BUF1 (N23085, N23075);
or OR4 (N23086, N23084, N20032, N17200, N669);
nand NAND3 (N23087, N23079, N20646, N2728);
nand NAND4 (N23088, N23081, N21514, N19158, N14381);
nor NOR2 (N23089, N23083, N3041);
xor XOR2 (N23090, N23072, N3201);
or OR2 (N23091, N23080, N10266);
and AND3 (N23092, N23090, N1645, N18693);
nor NOR4 (N23093, N23077, N5464, N2170, N1141);
nand NAND2 (N23094, N23076, N3903);
or OR2 (N23095, N23091, N1153);
and AND3 (N23096, N23093, N12656, N4844);
not NOT1 (N23097, N23092);
nor NOR4 (N23098, N23095, N3073, N12277, N20897);
xor XOR2 (N23099, N23096, N14697);
or OR4 (N23100, N23086, N13596, N11589, N13725);
not NOT1 (N23101, N23099);
buf BUF1 (N23102, N23089);
and AND2 (N23103, N23097, N14775);
nand NAND3 (N23104, N23094, N5490, N1103);
or OR4 (N23105, N23088, N20705, N8485, N23047);
xor XOR2 (N23106, N23101, N12655);
nor NOR3 (N23107, N23103, N20065, N1787);
and AND4 (N23108, N23107, N14332, N6812, N9319);
nor NOR3 (N23109, N23085, N2066, N21567);
xor XOR2 (N23110, N23074, N20436);
xor XOR2 (N23111, N23098, N14389);
not NOT1 (N23112, N23100);
not NOT1 (N23113, N23105);
xor XOR2 (N23114, N23104, N5632);
xor XOR2 (N23115, N23102, N21722);
nor NOR3 (N23116, N23109, N4343, N13887);
nand NAND4 (N23117, N23108, N19115, N10618, N18101);
nand NAND3 (N23118, N23087, N5455, N4896);
not NOT1 (N23119, N23116);
not NOT1 (N23120, N23106);
not NOT1 (N23121, N23110);
or OR2 (N23122, N23114, N255);
buf BUF1 (N23123, N23113);
nand NAND2 (N23124, N23120, N7824);
not NOT1 (N23125, N23117);
not NOT1 (N23126, N23124);
or OR2 (N23127, N23126, N16278);
nor NOR3 (N23128, N23123, N3916, N5692);
not NOT1 (N23129, N23125);
nand NAND3 (N23130, N23118, N22764, N7206);
xor XOR2 (N23131, N23111, N8481);
buf BUF1 (N23132, N23131);
xor XOR2 (N23133, N23130, N12204);
nor NOR4 (N23134, N23133, N6333, N6952, N21962);
nand NAND4 (N23135, N23132, N474, N8096, N9200);
or OR2 (N23136, N23121, N15897);
and AND4 (N23137, N23112, N15867, N10967, N15310);
nor NOR2 (N23138, N23135, N16633);
buf BUF1 (N23139, N23136);
or OR4 (N23140, N23139, N20102, N17783, N16548);
buf BUF1 (N23141, N23127);
and AND4 (N23142, N23115, N4286, N17136, N3514);
not NOT1 (N23143, N23142);
nand NAND3 (N23144, N23119, N8477, N3614);
nand NAND2 (N23145, N23128, N7539);
nand NAND4 (N23146, N23144, N5900, N17481, N13635);
nor NOR4 (N23147, N23145, N23076, N2993, N23130);
buf BUF1 (N23148, N23141);
xor XOR2 (N23149, N23148, N19892);
not NOT1 (N23150, N23147);
and AND3 (N23151, N23150, N6251, N17514);
and AND4 (N23152, N23122, N4742, N20291, N10138);
or OR2 (N23153, N23152, N1931);
or OR3 (N23154, N23149, N21167, N890);
buf BUF1 (N23155, N23129);
and AND2 (N23156, N23137, N10460);
nand NAND2 (N23157, N23155, N10885);
and AND3 (N23158, N23157, N17044, N1666);
xor XOR2 (N23159, N23140, N15650);
not NOT1 (N23160, N23138);
nor NOR3 (N23161, N23151, N9989, N485);
nor NOR2 (N23162, N23160, N4752);
not NOT1 (N23163, N23156);
nor NOR4 (N23164, N23161, N1011, N6109, N5861);
xor XOR2 (N23165, N23162, N7367);
not NOT1 (N23166, N23165);
buf BUF1 (N23167, N23154);
buf BUF1 (N23168, N23146);
and AND3 (N23169, N23134, N17224, N19355);
nand NAND3 (N23170, N23163, N11855, N20557);
and AND2 (N23171, N23153, N8678);
buf BUF1 (N23172, N23168);
xor XOR2 (N23173, N23158, N16039);
buf BUF1 (N23174, N23166);
nand NAND2 (N23175, N23174, N22034);
buf BUF1 (N23176, N23169);
or OR4 (N23177, N23172, N12972, N1358, N2780);
xor XOR2 (N23178, N23159, N5041);
or OR4 (N23179, N23178, N5733, N5973, N10819);
buf BUF1 (N23180, N23170);
and AND3 (N23181, N23175, N3994, N21030);
and AND3 (N23182, N23167, N19177, N16682);
xor XOR2 (N23183, N23181, N20742);
nor NOR4 (N23184, N23183, N3411, N2646, N16813);
xor XOR2 (N23185, N23180, N4568);
buf BUF1 (N23186, N23164);
nor NOR3 (N23187, N23173, N7305, N959);
xor XOR2 (N23188, N23179, N12688);
nor NOR2 (N23189, N23187, N3102);
and AND2 (N23190, N23186, N1511);
or OR3 (N23191, N23188, N1697, N7137);
and AND3 (N23192, N23182, N11800, N20252);
and AND3 (N23193, N23185, N13460, N13928);
nand NAND3 (N23194, N23177, N4387, N23040);
nand NAND2 (N23195, N23176, N22944);
nand NAND3 (N23196, N23193, N6146, N15049);
or OR2 (N23197, N23192, N21435);
nor NOR2 (N23198, N23195, N8768);
not NOT1 (N23199, N23184);
buf BUF1 (N23200, N23191);
not NOT1 (N23201, N23189);
or OR4 (N23202, N23171, N12803, N18094, N15841);
nand NAND4 (N23203, N23194, N19243, N4692, N12473);
or OR3 (N23204, N23143, N4224, N858);
xor XOR2 (N23205, N23203, N16069);
nand NAND2 (N23206, N23197, N15461);
and AND2 (N23207, N23201, N11034);
nand NAND4 (N23208, N23198, N14157, N15935, N2010);
and AND3 (N23209, N23205, N3999, N20736);
nand NAND2 (N23210, N23204, N15176);
nor NOR4 (N23211, N23208, N11905, N9716, N21063);
buf BUF1 (N23212, N23206);
xor XOR2 (N23213, N23211, N14064);
nor NOR4 (N23214, N23212, N13327, N22489, N13875);
xor XOR2 (N23215, N23214, N3959);
and AND4 (N23216, N23190, N6759, N963, N13102);
not NOT1 (N23217, N23209);
or OR2 (N23218, N23200, N13584);
and AND4 (N23219, N23210, N12787, N12548, N1244);
or OR2 (N23220, N23218, N3390);
xor XOR2 (N23221, N23207, N11676);
or OR4 (N23222, N23213, N22956, N1963, N16008);
nor NOR4 (N23223, N23202, N12687, N9315, N18572);
xor XOR2 (N23224, N23220, N18886);
nand NAND3 (N23225, N23221, N688, N3906);
or OR2 (N23226, N23219, N6086);
xor XOR2 (N23227, N23223, N22599);
or OR3 (N23228, N23225, N11853, N21649);
buf BUF1 (N23229, N23199);
and AND4 (N23230, N23226, N3936, N9395, N4543);
or OR3 (N23231, N23222, N13733, N4081);
or OR4 (N23232, N23196, N5899, N2942, N15368);
not NOT1 (N23233, N23228);
nor NOR4 (N23234, N23216, N56, N1637, N7035);
or OR3 (N23235, N23234, N5665, N498);
and AND4 (N23236, N23215, N8792, N9324, N17925);
nor NOR3 (N23237, N23229, N20821, N19856);
and AND2 (N23238, N23230, N8159);
buf BUF1 (N23239, N23235);
and AND2 (N23240, N23233, N9567);
nor NOR4 (N23241, N23237, N8063, N11994, N10946);
nand NAND4 (N23242, N23236, N20869, N1018, N5205);
not NOT1 (N23243, N23217);
nor NOR2 (N23244, N23243, N9080);
xor XOR2 (N23245, N23232, N2471);
not NOT1 (N23246, N23239);
buf BUF1 (N23247, N23231);
nor NOR2 (N23248, N23227, N10781);
buf BUF1 (N23249, N23244);
or OR4 (N23250, N23248, N7329, N1535, N14355);
not NOT1 (N23251, N23247);
buf BUF1 (N23252, N23249);
buf BUF1 (N23253, N23238);
not NOT1 (N23254, N23242);
not NOT1 (N23255, N23254);
or OR3 (N23256, N23240, N3085, N1308);
buf BUF1 (N23257, N23253);
or OR4 (N23258, N23245, N1314, N787, N6246);
and AND4 (N23259, N23251, N4234, N13222, N2864);
xor XOR2 (N23260, N23255, N12830);
and AND2 (N23261, N23250, N8154);
buf BUF1 (N23262, N23246);
and AND3 (N23263, N23261, N11109, N22293);
or OR3 (N23264, N23259, N3959, N22483);
nand NAND2 (N23265, N23258, N17923);
buf BUF1 (N23266, N23262);
not NOT1 (N23267, N23256);
and AND2 (N23268, N23267, N19414);
not NOT1 (N23269, N23263);
not NOT1 (N23270, N23257);
nand NAND3 (N23271, N23270, N18506, N10638);
xor XOR2 (N23272, N23268, N1495);
or OR3 (N23273, N23252, N12009, N16171);
buf BUF1 (N23274, N23260);
not NOT1 (N23275, N23265);
nand NAND2 (N23276, N23264, N7002);
and AND4 (N23277, N23273, N16388, N1330, N19861);
xor XOR2 (N23278, N23277, N18570);
or OR4 (N23279, N23274, N21512, N21763, N8232);
nand NAND3 (N23280, N23266, N19620, N17040);
not NOT1 (N23281, N23275);
or OR3 (N23282, N23224, N15927, N3522);
and AND3 (N23283, N23269, N4638, N552);
nor NOR3 (N23284, N23241, N21948, N18930);
buf BUF1 (N23285, N23271);
xor XOR2 (N23286, N23282, N22545);
xor XOR2 (N23287, N23276, N21588);
and AND4 (N23288, N23280, N2283, N1924, N17090);
buf BUF1 (N23289, N23281);
buf BUF1 (N23290, N23284);
nand NAND4 (N23291, N23283, N9292, N4668, N12297);
buf BUF1 (N23292, N23279);
or OR2 (N23293, N23292, N4237);
buf BUF1 (N23294, N23290);
buf BUF1 (N23295, N23289);
buf BUF1 (N23296, N23288);
buf BUF1 (N23297, N23293);
not NOT1 (N23298, N23285);
not NOT1 (N23299, N23287);
nand NAND3 (N23300, N23297, N9711, N8921);
nor NOR2 (N23301, N23298, N22393);
or OR3 (N23302, N23301, N101, N4484);
xor XOR2 (N23303, N23295, N12820);
or OR4 (N23304, N23299, N1356, N9929, N13116);
buf BUF1 (N23305, N23291);
buf BUF1 (N23306, N23305);
nand NAND2 (N23307, N23304, N7953);
xor XOR2 (N23308, N23272, N3601);
nor NOR3 (N23309, N23306, N6846, N19593);
buf BUF1 (N23310, N23303);
buf BUF1 (N23311, N23302);
or OR4 (N23312, N23296, N15710, N16295, N16726);
nand NAND4 (N23313, N23309, N9887, N6475, N22378);
nor NOR2 (N23314, N23312, N47);
buf BUF1 (N23315, N23300);
not NOT1 (N23316, N23310);
not NOT1 (N23317, N23311);
nor NOR3 (N23318, N23315, N11232, N21172);
or OR4 (N23319, N23294, N2071, N10440, N852);
buf BUF1 (N23320, N23278);
not NOT1 (N23321, N23318);
and AND2 (N23322, N23308, N16314);
and AND2 (N23323, N23317, N951);
nand NAND4 (N23324, N23314, N9398, N16231, N2851);
xor XOR2 (N23325, N23321, N15232);
not NOT1 (N23326, N23325);
nand NAND4 (N23327, N23307, N15696, N10205, N5848);
not NOT1 (N23328, N23323);
nor NOR2 (N23329, N23322, N19637);
or OR4 (N23330, N23324, N4381, N6957, N4009);
not NOT1 (N23331, N23319);
nor NOR4 (N23332, N23329, N8503, N12844, N6221);
buf BUF1 (N23333, N23328);
not NOT1 (N23334, N23316);
buf BUF1 (N23335, N23332);
nand NAND4 (N23336, N23327, N14711, N19672, N4604);
or OR4 (N23337, N23286, N18901, N12130, N12662);
buf BUF1 (N23338, N23320);
nand NAND2 (N23339, N23338, N11646);
nor NOR3 (N23340, N23313, N16938, N8726);
not NOT1 (N23341, N23335);
xor XOR2 (N23342, N23330, N16906);
nor NOR4 (N23343, N23334, N1183, N2629, N5122);
or OR4 (N23344, N23340, N11209, N4549, N1441);
buf BUF1 (N23345, N23331);
not NOT1 (N23346, N23343);
not NOT1 (N23347, N23344);
or OR4 (N23348, N23347, N18248, N22740, N11929);
or OR4 (N23349, N23326, N19265, N12971, N15748);
or OR3 (N23350, N23348, N1423, N4470);
nor NOR2 (N23351, N23341, N2932);
or OR2 (N23352, N23333, N12804);
xor XOR2 (N23353, N23350, N3847);
not NOT1 (N23354, N23342);
buf BUF1 (N23355, N23351);
or OR4 (N23356, N23339, N8516, N22773, N16509);
nand NAND4 (N23357, N23337, N5526, N21925, N10365);
nor NOR4 (N23358, N23353, N20389, N5603, N16411);
not NOT1 (N23359, N23356);
nor NOR2 (N23360, N23336, N20901);
nor NOR2 (N23361, N23354, N1936);
buf BUF1 (N23362, N23359);
or OR4 (N23363, N23349, N12014, N16140, N5370);
nand NAND3 (N23364, N23346, N12947, N14339);
or OR4 (N23365, N23357, N6857, N11241, N11855);
nor NOR4 (N23366, N23363, N15089, N12725, N10904);
xor XOR2 (N23367, N23366, N4468);
xor XOR2 (N23368, N23367, N13290);
nor NOR2 (N23369, N23362, N14523);
nand NAND4 (N23370, N23360, N9290, N9918, N4365);
nand NAND3 (N23371, N23370, N14419, N10470);
xor XOR2 (N23372, N23371, N14017);
or OR2 (N23373, N23355, N19650);
and AND2 (N23374, N23372, N13958);
nand NAND2 (N23375, N23358, N4412);
nand NAND4 (N23376, N23374, N19707, N10241, N8399);
or OR2 (N23377, N23375, N3756);
buf BUF1 (N23378, N23368);
and AND2 (N23379, N23373, N14926);
and AND3 (N23380, N23361, N5859, N14951);
nor NOR3 (N23381, N23379, N13548, N21543);
nand NAND2 (N23382, N23378, N6446);
and AND4 (N23383, N23369, N5540, N10952, N18087);
or OR2 (N23384, N23376, N9276);
xor XOR2 (N23385, N23382, N5933);
nand NAND3 (N23386, N23381, N20135, N7469);
buf BUF1 (N23387, N23345);
or OR4 (N23388, N23383, N3941, N16025, N22309);
and AND2 (N23389, N23385, N6173);
nor NOR2 (N23390, N23365, N11391);
buf BUF1 (N23391, N23388);
buf BUF1 (N23392, N23352);
or OR3 (N23393, N23389, N7642, N4871);
nand NAND2 (N23394, N23380, N12864);
nor NOR4 (N23395, N23390, N13366, N21618, N6844);
nor NOR2 (N23396, N23393, N7428);
nand NAND2 (N23397, N23364, N20399);
not NOT1 (N23398, N23384);
buf BUF1 (N23399, N23387);
nor NOR2 (N23400, N23386, N14646);
nand NAND2 (N23401, N23398, N6910);
buf BUF1 (N23402, N23397);
or OR2 (N23403, N23400, N7085);
buf BUF1 (N23404, N23395);
nand NAND3 (N23405, N23377, N16943, N19423);
xor XOR2 (N23406, N23404, N5802);
not NOT1 (N23407, N23396);
and AND2 (N23408, N23403, N11944);
or OR4 (N23409, N23402, N17940, N14632, N20805);
not NOT1 (N23410, N23409);
or OR4 (N23411, N23410, N22833, N1959, N9566);
or OR2 (N23412, N23405, N22818);
xor XOR2 (N23413, N23391, N20360);
nor NOR4 (N23414, N23394, N22626, N11468, N7209);
nor NOR4 (N23415, N23407, N11708, N382, N4878);
and AND4 (N23416, N23411, N2900, N22972, N3292);
xor XOR2 (N23417, N23416, N22451);
buf BUF1 (N23418, N23399);
and AND4 (N23419, N23413, N20876, N12593, N17607);
xor XOR2 (N23420, N23408, N3119);
and AND3 (N23421, N23417, N1274, N17435);
not NOT1 (N23422, N23406);
and AND4 (N23423, N23392, N22882, N18960, N5153);
nand NAND3 (N23424, N23421, N8565, N21190);
nand NAND2 (N23425, N23420, N12897);
buf BUF1 (N23426, N23401);
nor NOR4 (N23427, N23426, N22255, N5681, N4718);
or OR2 (N23428, N23418, N11709);
or OR3 (N23429, N23415, N9363, N22335);
nor NOR2 (N23430, N23427, N23182);
not NOT1 (N23431, N23412);
not NOT1 (N23432, N23422);
nor NOR4 (N23433, N23424, N11700, N8370, N5443);
nor NOR4 (N23434, N23425, N7156, N11931, N2752);
not NOT1 (N23435, N23432);
and AND2 (N23436, N23429, N23419);
and AND2 (N23437, N19422, N8914);
buf BUF1 (N23438, N23436);
or OR4 (N23439, N23435, N9230, N13248, N9442);
or OR3 (N23440, N23437, N7469, N21911);
nand NAND4 (N23441, N23440, N12572, N1531, N22778);
xor XOR2 (N23442, N23438, N11666);
or OR4 (N23443, N23414, N19093, N11463, N20792);
not NOT1 (N23444, N23431);
xor XOR2 (N23445, N23434, N20736);
buf BUF1 (N23446, N23439);
xor XOR2 (N23447, N23430, N2576);
nand NAND4 (N23448, N23442, N18263, N18399, N17042);
nor NOR2 (N23449, N23444, N4927);
nor NOR4 (N23450, N23447, N20856, N18805, N13496);
nor NOR3 (N23451, N23423, N21717, N4470);
buf BUF1 (N23452, N23445);
buf BUF1 (N23453, N23452);
xor XOR2 (N23454, N23433, N19565);
and AND3 (N23455, N23454, N3763, N5148);
nor NOR3 (N23456, N23455, N18118, N12730);
nand NAND2 (N23457, N23448, N5082);
not NOT1 (N23458, N23451);
nand NAND3 (N23459, N23450, N4702, N541);
nand NAND3 (N23460, N23428, N23074, N4668);
nand NAND2 (N23461, N23456, N10178);
nand NAND2 (N23462, N23457, N1115);
not NOT1 (N23463, N23441);
not NOT1 (N23464, N23462);
not NOT1 (N23465, N23461);
or OR3 (N23466, N23460, N10058, N16180);
not NOT1 (N23467, N23459);
and AND2 (N23468, N23443, N2860);
nor NOR2 (N23469, N23449, N9786);
xor XOR2 (N23470, N23468, N5021);
and AND4 (N23471, N23465, N4448, N12269, N20174);
not NOT1 (N23472, N23453);
nor NOR3 (N23473, N23472, N5059, N9793);
or OR4 (N23474, N23466, N21615, N10998, N6577);
nand NAND3 (N23475, N23471, N8776, N3223);
not NOT1 (N23476, N23473);
nor NOR2 (N23477, N23463, N17148);
nor NOR2 (N23478, N23464, N5755);
not NOT1 (N23479, N23467);
not NOT1 (N23480, N23475);
buf BUF1 (N23481, N23469);
and AND2 (N23482, N23478, N1379);
not NOT1 (N23483, N23458);
or OR4 (N23484, N23479, N8332, N9294, N7618);
not NOT1 (N23485, N23482);
buf BUF1 (N23486, N23485);
nand NAND3 (N23487, N23480, N16259, N6175);
or OR3 (N23488, N23446, N14054, N6672);
nand NAND4 (N23489, N23477, N15500, N17573, N8557);
not NOT1 (N23490, N23488);
not NOT1 (N23491, N23483);
not NOT1 (N23492, N23490);
or OR2 (N23493, N23491, N1930);
nor NOR2 (N23494, N23487, N18737);
and AND2 (N23495, N23470, N8570);
nand NAND2 (N23496, N23493, N8108);
xor XOR2 (N23497, N23474, N15349);
nor NOR2 (N23498, N23489, N5862);
buf BUF1 (N23499, N23484);
buf BUF1 (N23500, N23494);
and AND3 (N23501, N23498, N6255, N22453);
xor XOR2 (N23502, N23496, N15354);
nand NAND4 (N23503, N23481, N10563, N16092, N21300);
buf BUF1 (N23504, N23495);
nor NOR4 (N23505, N23497, N7107, N1710, N21667);
nand NAND4 (N23506, N23504, N6056, N22682, N17217);
not NOT1 (N23507, N23486);
or OR2 (N23508, N23505, N9974);
nand NAND2 (N23509, N23508, N5534);
buf BUF1 (N23510, N23503);
nand NAND3 (N23511, N23507, N6667, N7284);
nor NOR4 (N23512, N23506, N23185, N11365, N10672);
and AND3 (N23513, N23500, N14012, N12390);
nand NAND3 (N23514, N23513, N10859, N11879);
nor NOR4 (N23515, N23501, N14807, N16929, N1601);
and AND3 (N23516, N23510, N6221, N3238);
nor NOR2 (N23517, N23511, N3132);
not NOT1 (N23518, N23515);
and AND2 (N23519, N23517, N19286);
nor NOR2 (N23520, N23519, N21396);
not NOT1 (N23521, N23509);
buf BUF1 (N23522, N23499);
and AND2 (N23523, N23522, N23101);
buf BUF1 (N23524, N23521);
xor XOR2 (N23525, N23524, N17892);
nand NAND4 (N23526, N23514, N2787, N22766, N12173);
or OR3 (N23527, N23512, N17288, N11914);
xor XOR2 (N23528, N23492, N18210);
nand NAND4 (N23529, N23528, N10717, N19331, N15484);
not NOT1 (N23530, N23526);
nor NOR4 (N23531, N23525, N689, N5100, N9523);
nor NOR4 (N23532, N23518, N6514, N5057, N4990);
xor XOR2 (N23533, N23529, N13365);
and AND3 (N23534, N23502, N1262, N13138);
buf BUF1 (N23535, N23476);
nor NOR4 (N23536, N23531, N16821, N7552, N13346);
buf BUF1 (N23537, N23532);
and AND2 (N23538, N23523, N8860);
and AND3 (N23539, N23533, N1601, N7049);
and AND4 (N23540, N23537, N4404, N8155, N14340);
nor NOR4 (N23541, N23520, N240, N20627, N12359);
xor XOR2 (N23542, N23534, N15447);
not NOT1 (N23543, N23539);
buf BUF1 (N23544, N23536);
nand NAND2 (N23545, N23541, N15461);
nor NOR3 (N23546, N23538, N19733, N19978);
xor XOR2 (N23547, N23543, N14889);
not NOT1 (N23548, N23530);
or OR4 (N23549, N23527, N17376, N10160, N4202);
buf BUF1 (N23550, N23549);
nand NAND3 (N23551, N23546, N14748, N57);
nor NOR3 (N23552, N23544, N15375, N17454);
and AND4 (N23553, N23552, N21630, N2264, N21451);
xor XOR2 (N23554, N23547, N18514);
not NOT1 (N23555, N23554);
nor NOR2 (N23556, N23548, N7719);
nand NAND3 (N23557, N23542, N9270, N9422);
xor XOR2 (N23558, N23545, N6404);
or OR4 (N23559, N23551, N4362, N12767, N2663);
not NOT1 (N23560, N23516);
nand NAND4 (N23561, N23560, N4345, N9679, N23451);
nor NOR3 (N23562, N23558, N13760, N14093);
and AND4 (N23563, N23540, N14196, N10054, N15364);
and AND3 (N23564, N23557, N13404, N10791);
nand NAND3 (N23565, N23555, N15213, N7845);
nand NAND4 (N23566, N23562, N9491, N14748, N8169);
xor XOR2 (N23567, N23565, N11315);
nor NOR2 (N23568, N23564, N14715);
and AND4 (N23569, N23563, N16697, N9299, N8263);
and AND2 (N23570, N23566, N1975);
xor XOR2 (N23571, N23553, N22930);
xor XOR2 (N23572, N23569, N19739);
xor XOR2 (N23573, N23570, N19041);
and AND4 (N23574, N23571, N21970, N17084, N3040);
and AND3 (N23575, N23561, N11390, N6503);
or OR3 (N23576, N23559, N4719, N1839);
and AND3 (N23577, N23575, N11736, N16036);
not NOT1 (N23578, N23568);
not NOT1 (N23579, N23567);
xor XOR2 (N23580, N23579, N13095);
buf BUF1 (N23581, N23550);
or OR3 (N23582, N23572, N18436, N10764);
and AND3 (N23583, N23582, N18599, N18609);
and AND4 (N23584, N23581, N22634, N23342, N209);
xor XOR2 (N23585, N23574, N9317);
or OR2 (N23586, N23585, N21166);
buf BUF1 (N23587, N23576);
nor NOR2 (N23588, N23577, N3399);
xor XOR2 (N23589, N23556, N18173);
nor NOR4 (N23590, N23584, N845, N17266, N5314);
not NOT1 (N23591, N23535);
nor NOR2 (N23592, N23590, N14943);
or OR3 (N23593, N23591, N6891, N9589);
nor NOR3 (N23594, N23589, N20752, N16924);
xor XOR2 (N23595, N23588, N8912);
buf BUF1 (N23596, N23578);
nor NOR3 (N23597, N23573, N8524, N1154);
buf BUF1 (N23598, N23583);
and AND2 (N23599, N23587, N11261);
nor NOR4 (N23600, N23580, N2882, N2162, N21204);
and AND3 (N23601, N23599, N15459, N6110);
xor XOR2 (N23602, N23586, N20736);
xor XOR2 (N23603, N23600, N14078);
nand NAND3 (N23604, N23602, N21849, N6676);
not NOT1 (N23605, N23604);
buf BUF1 (N23606, N23605);
xor XOR2 (N23607, N23603, N13006);
and AND4 (N23608, N23597, N11377, N14363, N12693);
or OR3 (N23609, N23607, N4049, N22260);
buf BUF1 (N23610, N23593);
or OR2 (N23611, N23609, N3309);
nand NAND4 (N23612, N23595, N7598, N20514, N1651);
buf BUF1 (N23613, N23611);
nor NOR4 (N23614, N23601, N4170, N18465, N21208);
or OR4 (N23615, N23594, N18191, N18879, N16857);
and AND2 (N23616, N23606, N20420);
and AND3 (N23617, N23610, N4287, N13426);
not NOT1 (N23618, N23616);
nand NAND2 (N23619, N23613, N17963);
nand NAND2 (N23620, N23618, N13691);
buf BUF1 (N23621, N23614);
xor XOR2 (N23622, N23612, N13709);
and AND2 (N23623, N23596, N9826);
nand NAND3 (N23624, N23592, N12758, N19409);
xor XOR2 (N23625, N23619, N5746);
and AND3 (N23626, N23623, N18883, N18129);
buf BUF1 (N23627, N23626);
not NOT1 (N23628, N23620);
nor NOR2 (N23629, N23624, N15281);
not NOT1 (N23630, N23617);
nor NOR4 (N23631, N23628, N4805, N18382, N21572);
xor XOR2 (N23632, N23598, N13432);
nand NAND2 (N23633, N23627, N5797);
buf BUF1 (N23634, N23631);
nand NAND4 (N23635, N23633, N9059, N5483, N1625);
and AND4 (N23636, N23621, N420, N11553, N3105);
nand NAND2 (N23637, N23608, N239);
not NOT1 (N23638, N23634);
not NOT1 (N23639, N23629);
buf BUF1 (N23640, N23635);
buf BUF1 (N23641, N23639);
or OR3 (N23642, N23615, N15043, N17967);
nor NOR3 (N23643, N23637, N4284, N15897);
or OR2 (N23644, N23630, N16674);
nor NOR2 (N23645, N23644, N10266);
or OR4 (N23646, N23643, N11963, N7961, N6853);
nand NAND3 (N23647, N23632, N22388, N5339);
or OR4 (N23648, N23642, N15238, N5788, N14157);
or OR2 (N23649, N23646, N3077);
xor XOR2 (N23650, N23622, N7402);
nor NOR4 (N23651, N23640, N12294, N11667, N8466);
or OR3 (N23652, N23648, N4913, N3614);
buf BUF1 (N23653, N23638);
and AND2 (N23654, N23649, N9177);
nor NOR2 (N23655, N23645, N9903);
buf BUF1 (N23656, N23641);
and AND2 (N23657, N23647, N6868);
or OR4 (N23658, N23625, N18901, N1406, N2966);
or OR2 (N23659, N23650, N19411);
or OR4 (N23660, N23657, N2851, N7704, N7504);
not NOT1 (N23661, N23660);
nand NAND4 (N23662, N23661, N22068, N14398, N14738);
nor NOR4 (N23663, N23656, N5446, N8080, N4081);
and AND4 (N23664, N23651, N13527, N6902, N17321);
xor XOR2 (N23665, N23654, N5147);
and AND4 (N23666, N23636, N18393, N13806, N16281);
nand NAND3 (N23667, N23662, N18521, N10154);
nand NAND4 (N23668, N23663, N4555, N21303, N5853);
or OR4 (N23669, N23655, N14113, N465, N13158);
not NOT1 (N23670, N23667);
not NOT1 (N23671, N23670);
buf BUF1 (N23672, N23653);
buf BUF1 (N23673, N23665);
or OR3 (N23674, N23658, N5282, N19287);
nand NAND4 (N23675, N23652, N19151, N9881, N15378);
nor NOR2 (N23676, N23675, N22895);
xor XOR2 (N23677, N23673, N11947);
buf BUF1 (N23678, N23666);
nor NOR3 (N23679, N23668, N10657, N23660);
nand NAND2 (N23680, N23676, N44);
or OR4 (N23681, N23671, N4189, N13199, N13949);
or OR3 (N23682, N23678, N22840, N16092);
not NOT1 (N23683, N23682);
or OR3 (N23684, N23677, N9415, N20152);
or OR2 (N23685, N23679, N5903);
not NOT1 (N23686, N23659);
not NOT1 (N23687, N23686);
xor XOR2 (N23688, N23672, N11784);
nand NAND2 (N23689, N23688, N1178);
and AND3 (N23690, N23681, N15300, N1525);
or OR3 (N23691, N23689, N17874, N10302);
or OR4 (N23692, N23664, N7175, N22330, N19715);
or OR4 (N23693, N23684, N18113, N5320, N10486);
nand NAND4 (N23694, N23674, N11174, N10053, N3113);
nand NAND3 (N23695, N23680, N12739, N2898);
and AND2 (N23696, N23694, N9428);
and AND2 (N23697, N23692, N14244);
or OR4 (N23698, N23693, N5708, N5885, N15002);
nand NAND2 (N23699, N23691, N23345);
or OR2 (N23700, N23697, N5270);
or OR3 (N23701, N23700, N23043, N10649);
buf BUF1 (N23702, N23687);
xor XOR2 (N23703, N23695, N18571);
or OR3 (N23704, N23696, N13917, N18325);
nor NOR3 (N23705, N23703, N22581, N8726);
nand NAND3 (N23706, N23685, N17201, N22074);
buf BUF1 (N23707, N23706);
xor XOR2 (N23708, N23698, N15670);
or OR3 (N23709, N23690, N16377, N11361);
and AND3 (N23710, N23702, N15979, N13369);
nand NAND3 (N23711, N23710, N11896, N19752);
nor NOR3 (N23712, N23709, N3125, N17541);
not NOT1 (N23713, N23699);
nand NAND2 (N23714, N23701, N17970);
nand NAND4 (N23715, N23705, N10329, N6390, N12921);
xor XOR2 (N23716, N23683, N4070);
buf BUF1 (N23717, N23715);
nor NOR3 (N23718, N23713, N22723, N22812);
or OR2 (N23719, N23718, N22986);
xor XOR2 (N23720, N23707, N21214);
nor NOR2 (N23721, N23717, N15190);
nand NAND2 (N23722, N23714, N1437);
and AND4 (N23723, N23704, N21398, N13792, N3698);
or OR3 (N23724, N23716, N7216, N9057);
nand NAND2 (N23725, N23708, N12316);
or OR3 (N23726, N23724, N5024, N21074);
not NOT1 (N23727, N23725);
nor NOR3 (N23728, N23669, N9543, N14066);
not NOT1 (N23729, N23720);
and AND3 (N23730, N23727, N17010, N21063);
nand NAND4 (N23731, N23729, N17728, N15760, N6088);
or OR4 (N23732, N23731, N10058, N16766, N4816);
nor NOR4 (N23733, N23723, N22117, N15917, N18493);
nand NAND4 (N23734, N23711, N3328, N17308, N4330);
nand NAND4 (N23735, N23733, N13311, N9354, N6224);
not NOT1 (N23736, N23721);
xor XOR2 (N23737, N23736, N12415);
buf BUF1 (N23738, N23735);
and AND2 (N23739, N23712, N10120);
and AND4 (N23740, N23728, N8418, N2175, N15829);
buf BUF1 (N23741, N23734);
nand NAND4 (N23742, N23741, N4265, N22283, N3311);
nor NOR2 (N23743, N23742, N5960);
nand NAND3 (N23744, N23719, N21489, N18653);
xor XOR2 (N23745, N23739, N22180);
or OR3 (N23746, N23732, N8012, N8978);
nand NAND2 (N23747, N23745, N8118);
nor NOR2 (N23748, N23738, N11581);
nor NOR3 (N23749, N23747, N19687, N19923);
nor NOR4 (N23750, N23749, N15226, N9781, N22566);
nor NOR3 (N23751, N23744, N12073, N15625);
and AND2 (N23752, N23740, N23707);
nor NOR3 (N23753, N23752, N17762, N19234);
nand NAND3 (N23754, N23722, N6845, N7969);
buf BUF1 (N23755, N23730);
and AND4 (N23756, N23754, N11496, N20365, N23520);
or OR4 (N23757, N23746, N9469, N11144, N18496);
buf BUF1 (N23758, N23756);
not NOT1 (N23759, N23757);
and AND3 (N23760, N23755, N6783, N14853);
and AND3 (N23761, N23759, N18325, N11715);
xor XOR2 (N23762, N23761, N16722);
nand NAND4 (N23763, N23737, N16792, N20078, N12524);
or OR4 (N23764, N23726, N9024, N20510, N10452);
xor XOR2 (N23765, N23758, N17211);
nand NAND3 (N23766, N23762, N1870, N11459);
nor NOR4 (N23767, N23753, N18176, N670, N20528);
and AND3 (N23768, N23743, N23327, N2543);
xor XOR2 (N23769, N23766, N982);
xor XOR2 (N23770, N23765, N9047);
nand NAND2 (N23771, N23750, N14767);
buf BUF1 (N23772, N23751);
or OR2 (N23773, N23771, N2576);
xor XOR2 (N23774, N23772, N20265);
or OR2 (N23775, N23763, N3729);
nand NAND3 (N23776, N23767, N6447, N15668);
nor NOR4 (N23777, N23770, N14508, N8395, N16010);
or OR2 (N23778, N23774, N13232);
nand NAND2 (N23779, N23775, N15459);
buf BUF1 (N23780, N23776);
and AND2 (N23781, N23760, N172);
nand NAND4 (N23782, N23764, N5691, N18164, N1927);
buf BUF1 (N23783, N23778);
xor XOR2 (N23784, N23779, N4109);
not NOT1 (N23785, N23773);
nand NAND4 (N23786, N23781, N6745, N22578, N14900);
nand NAND3 (N23787, N23784, N567, N9374);
buf BUF1 (N23788, N23777);
or OR3 (N23789, N23782, N10580, N4921);
nor NOR2 (N23790, N23768, N23603);
or OR4 (N23791, N23786, N9251, N19216, N19839);
nor NOR2 (N23792, N23791, N11216);
or OR3 (N23793, N23748, N530, N15569);
nor NOR2 (N23794, N23789, N17266);
nand NAND3 (N23795, N23792, N1531, N16857);
and AND2 (N23796, N23788, N13825);
buf BUF1 (N23797, N23769);
or OR3 (N23798, N23790, N13838, N23567);
xor XOR2 (N23799, N23793, N22119);
xor XOR2 (N23800, N23799, N23634);
and AND2 (N23801, N23796, N21912);
nor NOR3 (N23802, N23787, N7446, N19215);
or OR4 (N23803, N23783, N19856, N10301, N15040);
xor XOR2 (N23804, N23798, N20207);
nor NOR4 (N23805, N23785, N17928, N13965, N7888);
and AND4 (N23806, N23794, N13054, N14882, N10875);
xor XOR2 (N23807, N23805, N23072);
and AND3 (N23808, N23797, N7309, N18875);
or OR3 (N23809, N23780, N12229, N12548);
and AND4 (N23810, N23808, N9599, N3182, N1292);
buf BUF1 (N23811, N23795);
nand NAND4 (N23812, N23806, N1907, N10508, N4098);
not NOT1 (N23813, N23809);
or OR2 (N23814, N23810, N19324);
and AND2 (N23815, N23802, N9495);
nand NAND4 (N23816, N23812, N1126, N4974, N14899);
nor NOR3 (N23817, N23800, N20984, N20421);
xor XOR2 (N23818, N23816, N22578);
nand NAND3 (N23819, N23803, N9713, N4630);
nand NAND3 (N23820, N23813, N14095, N10340);
and AND2 (N23821, N23811, N21984);
nor NOR4 (N23822, N23818, N7634, N23467, N17071);
nor NOR2 (N23823, N23822, N12259);
buf BUF1 (N23824, N23814);
and AND4 (N23825, N23819, N18705, N19513, N22324);
or OR4 (N23826, N23820, N4499, N15600, N16023);
not NOT1 (N23827, N23817);
nor NOR3 (N23828, N23825, N18354, N14783);
nand NAND3 (N23829, N23807, N19008, N8176);
and AND4 (N23830, N23815, N19029, N22447, N20376);
xor XOR2 (N23831, N23823, N5139);
and AND4 (N23832, N23830, N5199, N15134, N13822);
buf BUF1 (N23833, N23831);
nand NAND3 (N23834, N23827, N10552, N7286);
and AND3 (N23835, N23828, N7830, N19077);
buf BUF1 (N23836, N23834);
not NOT1 (N23837, N23836);
or OR3 (N23838, N23837, N1295, N11149);
nand NAND3 (N23839, N23833, N21155, N19227);
not NOT1 (N23840, N23824);
nand NAND4 (N23841, N23821, N973, N7028, N14372);
nand NAND2 (N23842, N23838, N19662);
nor NOR4 (N23843, N23840, N21848, N3112, N13905);
or OR2 (N23844, N23842, N15768);
and AND3 (N23845, N23843, N16404, N16410);
and AND3 (N23846, N23801, N23335, N22391);
not NOT1 (N23847, N23844);
or OR3 (N23848, N23832, N6342, N13441);
nor NOR2 (N23849, N23845, N7291);
buf BUF1 (N23850, N23826);
buf BUF1 (N23851, N23841);
or OR3 (N23852, N23835, N18867, N10198);
nor NOR4 (N23853, N23851, N4739, N13315, N8635);
and AND4 (N23854, N23804, N17213, N11219, N15509);
not NOT1 (N23855, N23853);
buf BUF1 (N23856, N23852);
not NOT1 (N23857, N23829);
not NOT1 (N23858, N23854);
nand NAND2 (N23859, N23839, N1530);
buf BUF1 (N23860, N23850);
buf BUF1 (N23861, N23849);
xor XOR2 (N23862, N23846, N20049);
nand NAND3 (N23863, N23857, N7565, N23018);
xor XOR2 (N23864, N23855, N6372);
buf BUF1 (N23865, N23860);
buf BUF1 (N23866, N23865);
nor NOR3 (N23867, N23863, N7728, N3426);
and AND3 (N23868, N23856, N18082, N15740);
xor XOR2 (N23869, N23858, N10662);
nor NOR3 (N23870, N23866, N9604, N22228);
nor NOR3 (N23871, N23869, N20928, N5003);
not NOT1 (N23872, N23861);
xor XOR2 (N23873, N23859, N14673);
nor NOR4 (N23874, N23872, N17680, N15349, N11470);
nand NAND4 (N23875, N23873, N17807, N2989, N5154);
nand NAND4 (N23876, N23862, N16139, N972, N13062);
nand NAND2 (N23877, N23871, N630);
or OR3 (N23878, N23868, N12007, N4262);
buf BUF1 (N23879, N23848);
and AND2 (N23880, N23879, N1417);
not NOT1 (N23881, N23878);
nand NAND4 (N23882, N23847, N17637, N3800, N4585);
buf BUF1 (N23883, N23876);
xor XOR2 (N23884, N23864, N23365);
and AND3 (N23885, N23884, N15191, N21279);
buf BUF1 (N23886, N23880);
or OR4 (N23887, N23877, N4896, N20197, N8440);
and AND3 (N23888, N23874, N1117, N21573);
nand NAND3 (N23889, N23886, N21204, N14900);
buf BUF1 (N23890, N23870);
not NOT1 (N23891, N23885);
nand NAND3 (N23892, N23888, N7737, N23239);
and AND3 (N23893, N23881, N6695, N20517);
not NOT1 (N23894, N23882);
nand NAND4 (N23895, N23894, N5402, N11261, N7100);
nand NAND4 (N23896, N23890, N8666, N12556, N7938);
and AND4 (N23897, N23896, N10852, N14663, N5895);
xor XOR2 (N23898, N23897, N10038);
nand NAND4 (N23899, N23892, N17546, N16194, N19889);
buf BUF1 (N23900, N23867);
or OR2 (N23901, N23893, N8738);
nor NOR4 (N23902, N23895, N12618, N23753, N16994);
nor NOR2 (N23903, N23889, N7259);
or OR2 (N23904, N23891, N4080);
buf BUF1 (N23905, N23887);
nand NAND3 (N23906, N23883, N5402, N13104);
or OR4 (N23907, N23875, N152, N2750, N18187);
and AND4 (N23908, N23898, N17629, N21472, N14012);
nor NOR3 (N23909, N23906, N11676, N16029);
xor XOR2 (N23910, N23905, N18191);
nor NOR4 (N23911, N23900, N3594, N20429, N16624);
nand NAND2 (N23912, N23904, N19397);
or OR2 (N23913, N23899, N18216);
buf BUF1 (N23914, N23901);
nor NOR3 (N23915, N23911, N22855, N8789);
not NOT1 (N23916, N23902);
and AND4 (N23917, N23916, N12727, N13761, N3494);
not NOT1 (N23918, N23903);
or OR2 (N23919, N23912, N2807);
or OR4 (N23920, N23914, N1262, N4604, N840);
or OR2 (N23921, N23920, N2625);
nor NOR4 (N23922, N23913, N5816, N22398, N20038);
nand NAND4 (N23923, N23915, N16562, N18553, N5382);
and AND3 (N23924, N23909, N23213, N18657);
buf BUF1 (N23925, N23919);
buf BUF1 (N23926, N23910);
not NOT1 (N23927, N23924);
nand NAND2 (N23928, N23923, N7156);
or OR4 (N23929, N23921, N8567, N19739, N2933);
nor NOR3 (N23930, N23918, N8548, N20568);
nand NAND3 (N23931, N23929, N22631, N9358);
buf BUF1 (N23932, N23926);
buf BUF1 (N23933, N23932);
nand NAND2 (N23934, N23907, N6454);
nor NOR2 (N23935, N23922, N8054);
nor NOR3 (N23936, N23933, N22279, N2461);
nor NOR3 (N23937, N23925, N9191, N174);
buf BUF1 (N23938, N23935);
not NOT1 (N23939, N23927);
xor XOR2 (N23940, N23936, N687);
not NOT1 (N23941, N23938);
and AND4 (N23942, N23908, N3782, N8448, N6308);
or OR3 (N23943, N23940, N882, N21455);
not NOT1 (N23944, N23939);
nand NAND2 (N23945, N23931, N22121);
not NOT1 (N23946, N23937);
and AND3 (N23947, N23944, N9025, N23580);
or OR3 (N23948, N23941, N4108, N11370);
xor XOR2 (N23949, N23930, N21237);
and AND3 (N23950, N23948, N16313, N16688);
nand NAND4 (N23951, N23950, N20197, N15879, N13510);
nand NAND2 (N23952, N23946, N4704);
nand NAND4 (N23953, N23952, N20278, N3713, N1482);
not NOT1 (N23954, N23949);
and AND4 (N23955, N23934, N12927, N12334, N2921);
nand NAND3 (N23956, N23953, N6812, N7798);
buf BUF1 (N23957, N23951);
not NOT1 (N23958, N23928);
or OR4 (N23959, N23957, N790, N18579, N901);
nor NOR3 (N23960, N23945, N6706, N3038);
buf BUF1 (N23961, N23960);
nand NAND2 (N23962, N23954, N21643);
and AND3 (N23963, N23962, N7412, N7632);
or OR3 (N23964, N23943, N5801, N8340);
and AND4 (N23965, N23942, N14401, N854, N20391);
or OR2 (N23966, N23917, N22828);
and AND2 (N23967, N23966, N18117);
nor NOR4 (N23968, N23963, N15416, N21764, N19599);
not NOT1 (N23969, N23967);
and AND4 (N23970, N23964, N12960, N12635, N17692);
not NOT1 (N23971, N23958);
or OR3 (N23972, N23959, N4048, N8713);
or OR4 (N23973, N23965, N17364, N15739, N10222);
nor NOR4 (N23974, N23972, N978, N10696, N11486);
xor XOR2 (N23975, N23970, N14900);
not NOT1 (N23976, N23974);
not NOT1 (N23977, N23961);
or OR4 (N23978, N23971, N6535, N8364, N5710);
nand NAND3 (N23979, N23975, N22683, N19716);
not NOT1 (N23980, N23968);
buf BUF1 (N23981, N23977);
xor XOR2 (N23982, N23976, N13607);
or OR4 (N23983, N23947, N1628, N1927, N19582);
nand NAND4 (N23984, N23983, N16316, N18414, N15643);
or OR4 (N23985, N23973, N7453, N13868, N4908);
buf BUF1 (N23986, N23984);
not NOT1 (N23987, N23982);
not NOT1 (N23988, N23980);
nand NAND2 (N23989, N23988, N11805);
or OR4 (N23990, N23969, N23651, N22523, N13551);
not NOT1 (N23991, N23979);
not NOT1 (N23992, N23989);
not NOT1 (N23993, N23986);
and AND3 (N23994, N23987, N14681, N20030);
or OR3 (N23995, N23956, N12598, N15499);
nor NOR3 (N23996, N23955, N2015, N216);
nor NOR2 (N23997, N23993, N14100);
xor XOR2 (N23998, N23991, N3280);
not NOT1 (N23999, N23994);
nand NAND3 (N24000, N23996, N17953, N971);
or OR3 (N24001, N23999, N2043, N5400);
xor XOR2 (N24002, N23985, N7946);
nand NAND4 (N24003, N23981, N1889, N2762, N14334);
not NOT1 (N24004, N23998);
xor XOR2 (N24005, N23995, N8868);
or OR3 (N24006, N24002, N21599, N14254);
buf BUF1 (N24007, N24006);
nor NOR4 (N24008, N24005, N6754, N9501, N13840);
nand NAND3 (N24009, N23978, N7359, N17579);
and AND2 (N24010, N24000, N13814);
nor NOR3 (N24011, N24001, N19798, N7270);
or OR2 (N24012, N24011, N17111);
and AND3 (N24013, N23990, N13778, N9765);
nor NOR3 (N24014, N24004, N21892, N21443);
xor XOR2 (N24015, N24007, N20553);
nand NAND3 (N24016, N24014, N14759, N5917);
nor NOR4 (N24017, N24008, N19201, N6340, N9622);
not NOT1 (N24018, N24009);
or OR3 (N24019, N24018, N3608, N16842);
or OR4 (N24020, N24003, N22887, N8069, N21357);
xor XOR2 (N24021, N24019, N16029);
nand NAND3 (N24022, N24015, N13148, N18881);
xor XOR2 (N24023, N24021, N9317);
not NOT1 (N24024, N24013);
buf BUF1 (N24025, N24016);
and AND3 (N24026, N24023, N18502, N11822);
xor XOR2 (N24027, N23997, N7985);
nand NAND2 (N24028, N24027, N21185);
xor XOR2 (N24029, N24026, N17203);
and AND2 (N24030, N24025, N703);
buf BUF1 (N24031, N24030);
nor NOR2 (N24032, N24012, N237);
nor NOR4 (N24033, N24017, N14827, N1900, N15374);
nand NAND3 (N24034, N24031, N16800, N5379);
xor XOR2 (N24035, N24028, N11827);
nand NAND4 (N24036, N24035, N21781, N14571, N6498);
or OR2 (N24037, N24024, N19109);
buf BUF1 (N24038, N24022);
xor XOR2 (N24039, N24010, N5065);
nor NOR2 (N24040, N24029, N6575);
and AND3 (N24041, N24038, N14072, N7032);
xor XOR2 (N24042, N24040, N11532);
and AND4 (N24043, N24032, N17856, N17811, N20388);
not NOT1 (N24044, N24042);
nand NAND2 (N24045, N24020, N14630);
nor NOR3 (N24046, N24043, N7300, N8832);
buf BUF1 (N24047, N24045);
nor NOR3 (N24048, N24039, N6999, N2246);
nand NAND2 (N24049, N24036, N22518);
xor XOR2 (N24050, N24034, N14901);
buf BUF1 (N24051, N24047);
or OR2 (N24052, N24048, N14191);
nor NOR3 (N24053, N24050, N22975, N23128);
buf BUF1 (N24054, N24041);
and AND4 (N24055, N24054, N15081, N18861, N12097);
nand NAND3 (N24056, N23992, N15826, N13494);
or OR3 (N24057, N24049, N4367, N23298);
nand NAND2 (N24058, N24055, N2111);
nor NOR2 (N24059, N24051, N11998);
buf BUF1 (N24060, N24058);
and AND2 (N24061, N24060, N1244);
xor XOR2 (N24062, N24056, N8938);
not NOT1 (N24063, N24061);
and AND4 (N24064, N24052, N2513, N12707, N8003);
and AND3 (N24065, N24064, N222, N14489);
buf BUF1 (N24066, N24063);
or OR3 (N24067, N24053, N16967, N1004);
nand NAND3 (N24068, N24062, N2947, N3143);
not NOT1 (N24069, N24066);
and AND4 (N24070, N24069, N11434, N8015, N11825);
xor XOR2 (N24071, N24068, N20013);
nor NOR2 (N24072, N24067, N23068);
buf BUF1 (N24073, N24037);
buf BUF1 (N24074, N24065);
xor XOR2 (N24075, N24057, N22769);
nor NOR2 (N24076, N24059, N9958);
xor XOR2 (N24077, N24033, N22512);
nand NAND4 (N24078, N24071, N3009, N10787, N8919);
buf BUF1 (N24079, N24073);
buf BUF1 (N24080, N24075);
not NOT1 (N24081, N24080);
xor XOR2 (N24082, N24081, N4152);
not NOT1 (N24083, N24072);
or OR2 (N24084, N24070, N15252);
or OR2 (N24085, N24082, N90);
not NOT1 (N24086, N24084);
or OR4 (N24087, N24083, N12622, N2293, N2759);
xor XOR2 (N24088, N24087, N21711);
xor XOR2 (N24089, N24074, N16310);
or OR2 (N24090, N24044, N20002);
and AND3 (N24091, N24086, N11066, N20264);
or OR2 (N24092, N24088, N244);
nand NAND3 (N24093, N24079, N7944, N18211);
nand NAND2 (N24094, N24078, N6307);
xor XOR2 (N24095, N24076, N14307);
buf BUF1 (N24096, N24095);
xor XOR2 (N24097, N24085, N6614);
not NOT1 (N24098, N24046);
nor NOR3 (N24099, N24096, N23481, N16424);
or OR2 (N24100, N24077, N9790);
nor NOR2 (N24101, N24097, N9145);
xor XOR2 (N24102, N24099, N22525);
and AND4 (N24103, N24102, N3665, N14688, N12536);
or OR2 (N24104, N24101, N11951);
nand NAND3 (N24105, N24098, N11545, N21287);
nand NAND3 (N24106, N24094, N18935, N9088);
not NOT1 (N24107, N24104);
nand NAND3 (N24108, N24089, N881, N4989);
nand NAND4 (N24109, N24107, N12539, N8020, N14584);
and AND2 (N24110, N24100, N766);
xor XOR2 (N24111, N24106, N1796);
nor NOR2 (N24112, N24092, N2751);
or OR4 (N24113, N24111, N2205, N15363, N20571);
not NOT1 (N24114, N24113);
buf BUF1 (N24115, N24090);
nand NAND3 (N24116, N24091, N20968, N6010);
nor NOR2 (N24117, N24110, N4051);
or OR4 (N24118, N24117, N14028, N790, N22280);
nor NOR3 (N24119, N24103, N7335, N6996);
buf BUF1 (N24120, N24105);
nand NAND3 (N24121, N24112, N7103, N12642);
nand NAND3 (N24122, N24120, N22950, N12467);
nand NAND4 (N24123, N24116, N20080, N13281, N23463);
xor XOR2 (N24124, N24121, N19860);
nor NOR2 (N24125, N24118, N14327);
xor XOR2 (N24126, N24109, N19412);
and AND4 (N24127, N24122, N18028, N9527, N7242);
xor XOR2 (N24128, N24127, N6265);
xor XOR2 (N24129, N24108, N1952);
and AND4 (N24130, N24119, N21962, N13571, N3389);
not NOT1 (N24131, N24123);
or OR2 (N24132, N24130, N5871);
not NOT1 (N24133, N24126);
not NOT1 (N24134, N24133);
nand NAND4 (N24135, N24125, N4479, N14880, N24052);
nor NOR4 (N24136, N24135, N15580, N21835, N7711);
and AND4 (N24137, N24093, N12545, N19355, N19422);
not NOT1 (N24138, N24115);
and AND3 (N24139, N24114, N15973, N1456);
nand NAND2 (N24140, N24139, N10795);
and AND2 (N24141, N24129, N21400);
buf BUF1 (N24142, N24141);
and AND3 (N24143, N24134, N7142, N7278);
or OR4 (N24144, N24136, N4559, N23917, N1847);
not NOT1 (N24145, N24131);
and AND4 (N24146, N24128, N13917, N7260, N15781);
nand NAND4 (N24147, N24140, N1069, N15268, N20269);
and AND3 (N24148, N24137, N8169, N3634);
not NOT1 (N24149, N24143);
and AND4 (N24150, N24144, N6212, N6893, N13526);
not NOT1 (N24151, N24132);
not NOT1 (N24152, N24138);
and AND3 (N24153, N24147, N10592, N10226);
xor XOR2 (N24154, N24146, N4119);
not NOT1 (N24155, N24145);
and AND4 (N24156, N24124, N608, N16130, N5848);
xor XOR2 (N24157, N24156, N18647);
not NOT1 (N24158, N24142);
and AND4 (N24159, N24149, N721, N5501, N12001);
nand NAND2 (N24160, N24159, N17242);
buf BUF1 (N24161, N24148);
buf BUF1 (N24162, N24153);
not NOT1 (N24163, N24155);
not NOT1 (N24164, N24160);
or OR2 (N24165, N24161, N23988);
not NOT1 (N24166, N24157);
not NOT1 (N24167, N24166);
and AND3 (N24168, N24162, N5616, N23770);
nand NAND2 (N24169, N24151, N17905);
not NOT1 (N24170, N24169);
nor NOR2 (N24171, N24165, N4055);
buf BUF1 (N24172, N24168);
xor XOR2 (N24173, N24158, N4784);
buf BUF1 (N24174, N24150);
and AND2 (N24175, N24154, N19398);
xor XOR2 (N24176, N24152, N12159);
nor NOR2 (N24177, N24173, N3999);
buf BUF1 (N24178, N24164);
not NOT1 (N24179, N24177);
xor XOR2 (N24180, N24174, N13478);
nor NOR2 (N24181, N24176, N7320);
not NOT1 (N24182, N24175);
xor XOR2 (N24183, N24179, N9391);
nand NAND3 (N24184, N24163, N20480, N23775);
not NOT1 (N24185, N24167);
nor NOR2 (N24186, N24171, N11746);
buf BUF1 (N24187, N24170);
and AND4 (N24188, N24182, N14020, N11830, N8842);
and AND3 (N24189, N24178, N9915, N15509);
or OR3 (N24190, N24183, N21970, N15261);
nor NOR2 (N24191, N24187, N5986);
xor XOR2 (N24192, N24186, N17760);
nor NOR3 (N24193, N24181, N18904, N8607);
xor XOR2 (N24194, N24193, N18962);
xor XOR2 (N24195, N24190, N8237);
and AND3 (N24196, N24172, N17554, N3573);
not NOT1 (N24197, N24189);
and AND4 (N24198, N24185, N5863, N19004, N4494);
nor NOR2 (N24199, N24197, N11722);
nor NOR2 (N24200, N24194, N5711);
not NOT1 (N24201, N24191);
buf BUF1 (N24202, N24195);
xor XOR2 (N24203, N24202, N4185);
or OR4 (N24204, N24188, N13150, N11631, N3464);
not NOT1 (N24205, N24203);
nor NOR2 (N24206, N24192, N20972);
or OR2 (N24207, N24198, N12824);
nand NAND2 (N24208, N24201, N5533);
buf BUF1 (N24209, N24196);
nor NOR3 (N24210, N24200, N11260, N22374);
and AND3 (N24211, N24199, N21654, N1072);
nand NAND4 (N24212, N24207, N10321, N6806, N6437);
nor NOR4 (N24213, N24184, N17099, N17641, N912);
nand NAND4 (N24214, N24205, N19483, N19714, N23062);
and AND3 (N24215, N24214, N13093, N15907);
xor XOR2 (N24216, N24180, N9205);
or OR3 (N24217, N24212, N13345, N4228);
not NOT1 (N24218, N24216);
nor NOR2 (N24219, N24213, N4892);
or OR3 (N24220, N24218, N16709, N901);
nand NAND3 (N24221, N24208, N19431, N7045);
not NOT1 (N24222, N24209);
nor NOR4 (N24223, N24210, N12167, N7459, N2172);
or OR3 (N24224, N24215, N1011, N18999);
nor NOR3 (N24225, N24204, N8890, N16223);
and AND4 (N24226, N24225, N1021, N4470, N10941);
not NOT1 (N24227, N24224);
and AND3 (N24228, N24220, N20193, N21931);
and AND2 (N24229, N24217, N21064);
and AND4 (N24230, N24228, N895, N12856, N18682);
not NOT1 (N24231, N24229);
nor NOR4 (N24232, N24211, N11801, N3993, N7263);
nand NAND2 (N24233, N24222, N7051);
nor NOR4 (N24234, N24233, N18633, N17528, N666);
nand NAND4 (N24235, N24223, N16598, N20853, N21423);
nor NOR4 (N24236, N24232, N2727, N22392, N11553);
or OR2 (N24237, N24206, N5957);
not NOT1 (N24238, N24219);
nand NAND4 (N24239, N24235, N23731, N11203, N8263);
nor NOR4 (N24240, N24226, N10467, N17287, N8370);
buf BUF1 (N24241, N24221);
nor NOR2 (N24242, N24236, N17006);
and AND2 (N24243, N24238, N22564);
xor XOR2 (N24244, N24240, N7308);
nand NAND2 (N24245, N24230, N14861);
or OR3 (N24246, N24237, N14982, N19872);
nor NOR2 (N24247, N24231, N20692);
or OR4 (N24248, N24244, N13653, N22017, N14975);
nor NOR3 (N24249, N24239, N19603, N22705);
and AND2 (N24250, N24246, N20629);
xor XOR2 (N24251, N24234, N19205);
or OR4 (N24252, N24245, N7530, N11286, N2866);
nand NAND3 (N24253, N24250, N22044, N10800);
not NOT1 (N24254, N24251);
nor NOR3 (N24255, N24253, N17647, N8082);
and AND4 (N24256, N24248, N21853, N8214, N18593);
or OR3 (N24257, N24243, N9300, N14794);
and AND3 (N24258, N24256, N12200, N17792);
nor NOR2 (N24259, N24242, N23705);
xor XOR2 (N24260, N24249, N21257);
buf BUF1 (N24261, N24259);
nand NAND4 (N24262, N24254, N9797, N7931, N2423);
nor NOR2 (N24263, N24252, N19664);
xor XOR2 (N24264, N24247, N2658);
nand NAND4 (N24265, N24260, N12290, N20240, N16125);
xor XOR2 (N24266, N24258, N15561);
nor NOR4 (N24267, N24255, N3440, N11865, N7425);
xor XOR2 (N24268, N24264, N9461);
and AND2 (N24269, N24241, N6342);
xor XOR2 (N24270, N24263, N19);
nor NOR3 (N24271, N24261, N15502, N18648);
nor NOR4 (N24272, N24257, N8047, N9971, N10297);
not NOT1 (N24273, N24227);
or OR3 (N24274, N24268, N12108, N2872);
and AND4 (N24275, N24267, N1311, N15004, N6293);
xor XOR2 (N24276, N24272, N1427);
nand NAND4 (N24277, N24273, N5146, N22748, N5346);
or OR2 (N24278, N24271, N18277);
not NOT1 (N24279, N24276);
and AND2 (N24280, N24262, N16323);
nand NAND3 (N24281, N24280, N21768, N19192);
nand NAND2 (N24282, N24266, N7395);
nor NOR3 (N24283, N24279, N575, N15837);
xor XOR2 (N24284, N24274, N10438);
nand NAND3 (N24285, N24269, N8549, N18383);
and AND3 (N24286, N24270, N19355, N2981);
not NOT1 (N24287, N24277);
xor XOR2 (N24288, N24275, N16790);
buf BUF1 (N24289, N24287);
nor NOR2 (N24290, N24278, N8123);
not NOT1 (N24291, N24282);
buf BUF1 (N24292, N24265);
nand NAND2 (N24293, N24281, N9918);
xor XOR2 (N24294, N24292, N18239);
buf BUF1 (N24295, N24288);
buf BUF1 (N24296, N24285);
not NOT1 (N24297, N24289);
and AND2 (N24298, N24295, N7602);
or OR4 (N24299, N24283, N4653, N16603, N466);
not NOT1 (N24300, N24293);
or OR4 (N24301, N24294, N21735, N7498, N10093);
buf BUF1 (N24302, N24298);
xor XOR2 (N24303, N24299, N15991);
buf BUF1 (N24304, N24291);
xor XOR2 (N24305, N24296, N5745);
and AND4 (N24306, N24284, N5086, N5089, N6544);
or OR4 (N24307, N24300, N16233, N8379, N9074);
xor XOR2 (N24308, N24301, N21603);
and AND4 (N24309, N24308, N23668, N10357, N4305);
not NOT1 (N24310, N24307);
nand NAND3 (N24311, N24290, N4557, N6035);
or OR4 (N24312, N24302, N9432, N6081, N21080);
not NOT1 (N24313, N24304);
nor NOR2 (N24314, N24309, N17696);
buf BUF1 (N24315, N24297);
buf BUF1 (N24316, N24305);
and AND4 (N24317, N24286, N10685, N3721, N13106);
and AND2 (N24318, N24316, N7153);
nor NOR3 (N24319, N24310, N3003, N21521);
xor XOR2 (N24320, N24319, N23516);
nor NOR4 (N24321, N24306, N21570, N15038, N19208);
or OR4 (N24322, N24320, N17562, N14986, N17660);
nand NAND4 (N24323, N24318, N10638, N19729, N14177);
nand NAND3 (N24324, N24321, N16543, N12964);
buf BUF1 (N24325, N24324);
and AND4 (N24326, N24312, N6190, N22070, N18080);
or OR2 (N24327, N24311, N15809);
nor NOR4 (N24328, N24326, N13513, N15762, N24277);
nand NAND3 (N24329, N24325, N1057, N15155);
nand NAND3 (N24330, N24329, N10442, N5125);
nor NOR3 (N24331, N24323, N18923, N17692);
xor XOR2 (N24332, N24327, N22474);
or OR4 (N24333, N24330, N6325, N5504, N3664);
nor NOR2 (N24334, N24331, N16984);
nor NOR2 (N24335, N24333, N5887);
not NOT1 (N24336, N24332);
xor XOR2 (N24337, N24322, N4005);
or OR4 (N24338, N24317, N10930, N2234, N17156);
nor NOR2 (N24339, N24303, N19930);
buf BUF1 (N24340, N24336);
buf BUF1 (N24341, N24334);
and AND4 (N24342, N24341, N17252, N3106, N9395);
buf BUF1 (N24343, N24339);
nor NOR3 (N24344, N24338, N15584, N11626);
nor NOR2 (N24345, N24314, N18551);
nor NOR3 (N24346, N24335, N13679, N11001);
xor XOR2 (N24347, N24342, N9605);
or OR4 (N24348, N24347, N2157, N22850, N19845);
buf BUF1 (N24349, N24340);
xor XOR2 (N24350, N24349, N10770);
buf BUF1 (N24351, N24343);
nand NAND2 (N24352, N24348, N8063);
not NOT1 (N24353, N24315);
and AND4 (N24354, N24352, N20560, N14973, N17322);
nand NAND3 (N24355, N24313, N6405, N5385);
or OR2 (N24356, N24350, N2798);
or OR4 (N24357, N24328, N3196, N3183, N1582);
not NOT1 (N24358, N24357);
xor XOR2 (N24359, N24346, N10327);
nand NAND2 (N24360, N24356, N17501);
and AND2 (N24361, N24344, N11260);
or OR3 (N24362, N24354, N20496, N7466);
buf BUF1 (N24363, N24358);
buf BUF1 (N24364, N24363);
xor XOR2 (N24365, N24355, N19218);
buf BUF1 (N24366, N24361);
xor XOR2 (N24367, N24360, N16582);
not NOT1 (N24368, N24359);
or OR3 (N24369, N24364, N3536, N20475);
not NOT1 (N24370, N24365);
buf BUF1 (N24371, N24368);
nand NAND3 (N24372, N24351, N8540, N12285);
or OR3 (N24373, N24337, N13180, N22684);
not NOT1 (N24374, N24369);
not NOT1 (N24375, N24366);
or OR2 (N24376, N24345, N8383);
or OR3 (N24377, N24353, N18825, N10507);
nand NAND3 (N24378, N24362, N8393, N5051);
xor XOR2 (N24379, N24375, N21261);
nor NOR4 (N24380, N24367, N1531, N14902, N1100);
nand NAND3 (N24381, N24378, N16709, N8533);
buf BUF1 (N24382, N24370);
nand NAND2 (N24383, N24374, N12577);
not NOT1 (N24384, N24377);
and AND2 (N24385, N24382, N19726);
not NOT1 (N24386, N24371);
not NOT1 (N24387, N24385);
nor NOR3 (N24388, N24387, N13458, N21616);
nor NOR2 (N24389, N24381, N3361);
nand NAND3 (N24390, N24383, N21031, N22201);
and AND4 (N24391, N24390, N16184, N21010, N6114);
not NOT1 (N24392, N24376);
and AND2 (N24393, N24388, N24381);
nor NOR2 (N24394, N24391, N9300);
nand NAND3 (N24395, N24373, N4215, N3331);
not NOT1 (N24396, N24392);
xor XOR2 (N24397, N24386, N19301);
xor XOR2 (N24398, N24389, N17237);
nand NAND3 (N24399, N24379, N4449, N17800);
buf BUF1 (N24400, N24384);
not NOT1 (N24401, N24400);
nand NAND2 (N24402, N24372, N3554);
or OR2 (N24403, N24401, N21380);
not NOT1 (N24404, N24399);
buf BUF1 (N24405, N24396);
nor NOR3 (N24406, N24380, N19010, N5847);
nor NOR4 (N24407, N24398, N18972, N23621, N1499);
xor XOR2 (N24408, N24403, N8521);
and AND2 (N24409, N24405, N19878);
buf BUF1 (N24410, N24395);
not NOT1 (N24411, N24402);
nand NAND2 (N24412, N24397, N1748);
nor NOR2 (N24413, N24408, N16154);
and AND3 (N24414, N24413, N11083, N305);
xor XOR2 (N24415, N24414, N2186);
xor XOR2 (N24416, N24412, N1369);
nand NAND3 (N24417, N24393, N11218, N21895);
buf BUF1 (N24418, N24411);
buf BUF1 (N24419, N24417);
xor XOR2 (N24420, N24416, N17178);
xor XOR2 (N24421, N24418, N20856);
xor XOR2 (N24422, N24420, N5203);
and AND2 (N24423, N24394, N115);
not NOT1 (N24424, N24406);
nor NOR4 (N24425, N24422, N4752, N9957, N10466);
xor XOR2 (N24426, N24424, N11800);
buf BUF1 (N24427, N24415);
nand NAND3 (N24428, N24427, N5622, N16065);
xor XOR2 (N24429, N24421, N20429);
or OR3 (N24430, N24409, N2745, N1980);
buf BUF1 (N24431, N24429);
xor XOR2 (N24432, N24430, N11142);
buf BUF1 (N24433, N24432);
not NOT1 (N24434, N24404);
not NOT1 (N24435, N24434);
or OR3 (N24436, N24435, N7981, N11887);
nand NAND4 (N24437, N24428, N13549, N5746, N15956);
and AND2 (N24438, N24431, N18241);
xor XOR2 (N24439, N24423, N21913);
xor XOR2 (N24440, N24407, N20008);
not NOT1 (N24441, N24436);
buf BUF1 (N24442, N24441);
xor XOR2 (N24443, N24438, N13762);
xor XOR2 (N24444, N24443, N1597);
not NOT1 (N24445, N24440);
nand NAND2 (N24446, N24426, N22198);
not NOT1 (N24447, N24425);
xor XOR2 (N24448, N24439, N11202);
nor NOR3 (N24449, N24433, N10088, N18599);
xor XOR2 (N24450, N24442, N14115);
buf BUF1 (N24451, N24419);
nor NOR4 (N24452, N24410, N5215, N11779, N11879);
buf BUF1 (N24453, N24451);
nor NOR3 (N24454, N24445, N24011, N2127);
not NOT1 (N24455, N24446);
not NOT1 (N24456, N24454);
nor NOR2 (N24457, N24453, N24328);
nand NAND2 (N24458, N24452, N13796);
and AND4 (N24459, N24448, N8360, N434, N14045);
or OR3 (N24460, N24457, N19412, N7964);
nor NOR4 (N24461, N24455, N5846, N11097, N18026);
buf BUF1 (N24462, N24460);
and AND4 (N24463, N24450, N4703, N14141, N8595);
or OR4 (N24464, N24463, N24355, N18749, N7059);
nor NOR4 (N24465, N24462, N14349, N9394, N10858);
or OR4 (N24466, N24461, N10889, N13800, N21384);
nand NAND4 (N24467, N24447, N7541, N16101, N20850);
xor XOR2 (N24468, N24459, N7228);
and AND4 (N24469, N24467, N1481, N658, N1746);
buf BUF1 (N24470, N24456);
and AND2 (N24471, N24469, N1651);
and AND2 (N24472, N24470, N19105);
not NOT1 (N24473, N24464);
nor NOR4 (N24474, N24465, N20718, N6284, N16281);
or OR2 (N24475, N24468, N17243);
nand NAND3 (N24476, N24458, N3957, N13550);
nand NAND4 (N24477, N24444, N4655, N10559, N23579);
nand NAND2 (N24478, N24466, N16816);
nand NAND4 (N24479, N24476, N14124, N10556, N18484);
nand NAND2 (N24480, N24477, N1079);
buf BUF1 (N24481, N24474);
not NOT1 (N24482, N24449);
not NOT1 (N24483, N24437);
xor XOR2 (N24484, N24482, N3613);
and AND4 (N24485, N24478, N23439, N639, N17408);
xor XOR2 (N24486, N24475, N14387);
nand NAND4 (N24487, N24484, N12615, N17092, N3527);
buf BUF1 (N24488, N24479);
xor XOR2 (N24489, N24486, N15914);
xor XOR2 (N24490, N24488, N7996);
xor XOR2 (N24491, N24481, N19220);
xor XOR2 (N24492, N24471, N11916);
and AND4 (N24493, N24485, N7486, N20744, N1143);
nand NAND2 (N24494, N24487, N17628);
buf BUF1 (N24495, N24473);
not NOT1 (N24496, N24491);
xor XOR2 (N24497, N24472, N452);
nor NOR4 (N24498, N24490, N16686, N9880, N6540);
xor XOR2 (N24499, N24480, N5556);
buf BUF1 (N24500, N24493);
buf BUF1 (N24501, N24497);
xor XOR2 (N24502, N24501, N16142);
xor XOR2 (N24503, N24496, N12641);
buf BUF1 (N24504, N24502);
and AND4 (N24505, N24499, N5918, N24332, N20105);
nor NOR3 (N24506, N24495, N5009, N8222);
and AND2 (N24507, N24498, N8439);
nand NAND3 (N24508, N24483, N8665, N17400);
xor XOR2 (N24509, N24508, N17309);
or OR2 (N24510, N24506, N6145);
xor XOR2 (N24511, N24489, N378);
nand NAND3 (N24512, N24500, N187, N13186);
or OR2 (N24513, N24512, N19325);
nand NAND2 (N24514, N24510, N4549);
xor XOR2 (N24515, N24504, N10818);
nor NOR2 (N24516, N24513, N1628);
and AND4 (N24517, N24503, N22916, N1476, N8603);
nand NAND3 (N24518, N24511, N16310, N21501);
and AND2 (N24519, N24517, N20676);
not NOT1 (N24520, N24516);
not NOT1 (N24521, N24514);
xor XOR2 (N24522, N24519, N19530);
or OR3 (N24523, N24505, N1472, N24356);
xor XOR2 (N24524, N24522, N16840);
buf BUF1 (N24525, N24509);
and AND4 (N24526, N24523, N23196, N10980, N699);
or OR4 (N24527, N24525, N2286, N2994, N18626);
buf BUF1 (N24528, N24526);
xor XOR2 (N24529, N24492, N1417);
buf BUF1 (N24530, N24529);
and AND2 (N24531, N24520, N18107);
and AND2 (N24532, N24530, N20529);
nand NAND3 (N24533, N24494, N5822, N15366);
xor XOR2 (N24534, N24521, N18759);
and AND4 (N24535, N24507, N17097, N7337, N4704);
nor NOR2 (N24536, N24527, N7032);
xor XOR2 (N24537, N24534, N15770);
nor NOR3 (N24538, N24531, N1160, N17051);
buf BUF1 (N24539, N24536);
not NOT1 (N24540, N24524);
xor XOR2 (N24541, N24533, N19331);
nor NOR2 (N24542, N24515, N10036);
xor XOR2 (N24543, N24528, N10489);
nor NOR2 (N24544, N24539, N5401);
and AND4 (N24545, N24538, N21919, N6058, N4354);
and AND3 (N24546, N24537, N3963, N9845);
and AND2 (N24547, N24545, N5668);
buf BUF1 (N24548, N24547);
not NOT1 (N24549, N24543);
xor XOR2 (N24550, N24518, N22520);
and AND3 (N24551, N24550, N6413, N23675);
nor NOR3 (N24552, N24540, N4509, N21528);
nand NAND4 (N24553, N24551, N16301, N6162, N11685);
or OR4 (N24554, N24553, N15473, N16039, N1252);
and AND4 (N24555, N24535, N12092, N1732, N11577);
nand NAND4 (N24556, N24548, N6830, N13539, N15623);
or OR4 (N24557, N24542, N3388, N7062, N5491);
or OR3 (N24558, N24544, N9761, N11423);
nor NOR2 (N24559, N24532, N19803);
not NOT1 (N24560, N24557);
and AND4 (N24561, N24560, N1209, N16005, N1743);
not NOT1 (N24562, N24552);
nor NOR2 (N24563, N24558, N22087);
not NOT1 (N24564, N24541);
not NOT1 (N24565, N24562);
nor NOR3 (N24566, N24565, N5120, N19845);
nand NAND4 (N24567, N24555, N10422, N11394, N11611);
not NOT1 (N24568, N24549);
and AND2 (N24569, N24559, N17374);
nand NAND4 (N24570, N24569, N15784, N13088, N10203);
nand NAND3 (N24571, N24561, N22702, N10047);
xor XOR2 (N24572, N24571, N17541);
or OR2 (N24573, N24556, N19470);
buf BUF1 (N24574, N24570);
xor XOR2 (N24575, N24574, N9311);
nor NOR4 (N24576, N24567, N23793, N10985, N5916);
xor XOR2 (N24577, N24576, N23188);
nor NOR4 (N24578, N24566, N12350, N334, N1852);
nor NOR2 (N24579, N24563, N24461);
nor NOR2 (N24580, N24579, N23335);
nand NAND2 (N24581, N24554, N5288);
buf BUF1 (N24582, N24572);
nand NAND2 (N24583, N24575, N12030);
buf BUF1 (N24584, N24581);
xor XOR2 (N24585, N24564, N18349);
nor NOR3 (N24586, N24585, N8822, N3161);
nor NOR3 (N24587, N24546, N19716, N14671);
xor XOR2 (N24588, N24584, N19924);
and AND3 (N24589, N24583, N12307, N8311);
nor NOR2 (N24590, N24589, N20265);
buf BUF1 (N24591, N24587);
and AND2 (N24592, N24578, N15487);
nand NAND4 (N24593, N24592, N9902, N17085, N21573);
xor XOR2 (N24594, N24586, N24042);
or OR3 (N24595, N24590, N23621, N12716);
not NOT1 (N24596, N24588);
or OR2 (N24597, N24577, N16087);
and AND2 (N24598, N24580, N9017);
xor XOR2 (N24599, N24597, N5755);
xor XOR2 (N24600, N24582, N20316);
not NOT1 (N24601, N24594);
nand NAND2 (N24602, N24600, N19593);
buf BUF1 (N24603, N24599);
xor XOR2 (N24604, N24591, N24270);
and AND4 (N24605, N24598, N7755, N13444, N11470);
buf BUF1 (N24606, N24568);
nand NAND3 (N24607, N24596, N8178, N10822);
and AND3 (N24608, N24603, N11932, N13200);
or OR4 (N24609, N24573, N21598, N12800, N6551);
not NOT1 (N24610, N24605);
and AND3 (N24611, N24608, N18660, N13569);
not NOT1 (N24612, N24606);
buf BUF1 (N24613, N24601);
and AND3 (N24614, N24595, N18297, N8785);
xor XOR2 (N24615, N24614, N12327);
nor NOR2 (N24616, N24593, N18694);
nor NOR4 (N24617, N24615, N12447, N4256, N21265);
not NOT1 (N24618, N24613);
buf BUF1 (N24619, N24609);
or OR2 (N24620, N24611, N22173);
nand NAND2 (N24621, N24607, N2600);
nand NAND3 (N24622, N24618, N3731, N1162);
and AND2 (N24623, N24622, N15235);
or OR4 (N24624, N24616, N11877, N9841, N20898);
nand NAND4 (N24625, N24621, N845, N3547, N11327);
nand NAND2 (N24626, N24610, N18667);
nor NOR4 (N24627, N24617, N10752, N1128, N9764);
and AND4 (N24628, N24612, N12410, N11977, N21042);
and AND3 (N24629, N24625, N9533, N18241);
buf BUF1 (N24630, N24624);
xor XOR2 (N24631, N24602, N9646);
xor XOR2 (N24632, N24628, N12426);
nand NAND3 (N24633, N24623, N15320, N731);
buf BUF1 (N24634, N24627);
nor NOR4 (N24635, N24604, N8376, N18914, N7234);
nor NOR3 (N24636, N24630, N15106, N12428);
xor XOR2 (N24637, N24629, N12396);
nand NAND3 (N24638, N24632, N12326, N22674);
nand NAND2 (N24639, N24638, N11536);
buf BUF1 (N24640, N24631);
xor XOR2 (N24641, N24619, N8812);
or OR3 (N24642, N24633, N20430, N18399);
buf BUF1 (N24643, N24640);
buf BUF1 (N24644, N24637);
and AND2 (N24645, N24644, N3413);
not NOT1 (N24646, N24639);
nor NOR2 (N24647, N24646, N21866);
and AND2 (N24648, N24620, N5073);
or OR4 (N24649, N24647, N7365, N20350, N7667);
or OR4 (N24650, N24649, N18597, N3198, N17677);
xor XOR2 (N24651, N24642, N21881);
buf BUF1 (N24652, N24643);
not NOT1 (N24653, N24634);
xor XOR2 (N24654, N24648, N16446);
buf BUF1 (N24655, N24652);
and AND4 (N24656, N24641, N19489, N24168, N23713);
nor NOR2 (N24657, N24645, N1491);
or OR4 (N24658, N24626, N17191, N10892, N21);
and AND3 (N24659, N24658, N7531, N8709);
buf BUF1 (N24660, N24657);
or OR3 (N24661, N24650, N4261, N22070);
and AND3 (N24662, N24660, N3652, N674);
or OR2 (N24663, N24654, N14384);
and AND4 (N24664, N24661, N19619, N21137, N528);
not NOT1 (N24665, N24662);
and AND2 (N24666, N24665, N13161);
and AND4 (N24667, N24656, N9582, N2502, N22822);
or OR2 (N24668, N24663, N14661);
buf BUF1 (N24669, N24635);
buf BUF1 (N24670, N24653);
buf BUF1 (N24671, N24655);
buf BUF1 (N24672, N24671);
nand NAND2 (N24673, N24651, N16610);
or OR2 (N24674, N24673, N9349);
or OR4 (N24675, N24659, N3793, N2222, N17);
not NOT1 (N24676, N24667);
buf BUF1 (N24677, N24675);
xor XOR2 (N24678, N24672, N21137);
not NOT1 (N24679, N24664);
nand NAND4 (N24680, N24674, N9046, N21153, N13487);
not NOT1 (N24681, N24677);
not NOT1 (N24682, N24636);
or OR2 (N24683, N24670, N20015);
and AND4 (N24684, N24676, N8209, N2616, N14110);
xor XOR2 (N24685, N24678, N13312);
or OR2 (N24686, N24680, N10483);
and AND4 (N24687, N24686, N12408, N9066, N4402);
not NOT1 (N24688, N24687);
buf BUF1 (N24689, N24668);
or OR2 (N24690, N24684, N22690);
or OR4 (N24691, N24682, N19775, N24269, N15657);
or OR4 (N24692, N24666, N22035, N19376, N4716);
nor NOR4 (N24693, N24679, N19094, N15072, N24457);
and AND3 (N24694, N24688, N21659, N12726);
xor XOR2 (N24695, N24691, N15718);
not NOT1 (N24696, N24693);
or OR3 (N24697, N24690, N10303, N9175);
and AND4 (N24698, N24695, N13266, N11614, N12170);
buf BUF1 (N24699, N24669);
buf BUF1 (N24700, N24699);
buf BUF1 (N24701, N24700);
nand NAND3 (N24702, N24683, N1255, N6540);
not NOT1 (N24703, N24694);
and AND4 (N24704, N24698, N10677, N10403, N22245);
nand NAND3 (N24705, N24685, N18878, N18974);
nor NOR4 (N24706, N24692, N22133, N18819, N1976);
and AND4 (N24707, N24703, N4221, N14904, N8303);
not NOT1 (N24708, N24707);
nand NAND4 (N24709, N24701, N23549, N11509, N9732);
or OR3 (N24710, N24696, N3527, N11329);
and AND4 (N24711, N24681, N9608, N8620, N10758);
not NOT1 (N24712, N24697);
and AND4 (N24713, N24706, N20459, N23534, N11195);
nor NOR2 (N24714, N24702, N7792);
nand NAND4 (N24715, N24714, N14151, N19325, N22878);
nand NAND4 (N24716, N24709, N515, N16242, N11059);
and AND3 (N24717, N24710, N9490, N11024);
buf BUF1 (N24718, N24716);
xor XOR2 (N24719, N24708, N19718);
not NOT1 (N24720, N24704);
nand NAND3 (N24721, N24717, N19416, N24605);
and AND4 (N24722, N24711, N6363, N22596, N11310);
and AND4 (N24723, N24713, N13013, N6401, N15402);
nand NAND4 (N24724, N24705, N24425, N16806, N4120);
or OR4 (N24725, N24719, N19583, N107, N19052);
nor NOR2 (N24726, N24715, N15056);
and AND4 (N24727, N24720, N9164, N14704, N447);
nand NAND4 (N24728, N24726, N197, N2515, N17386);
and AND3 (N24729, N24724, N7975, N4562);
xor XOR2 (N24730, N24728, N6248);
xor XOR2 (N24731, N24722, N20873);
not NOT1 (N24732, N24730);
or OR2 (N24733, N24689, N4130);
nor NOR3 (N24734, N24718, N1250, N23849);
buf BUF1 (N24735, N24731);
and AND2 (N24736, N24734, N6517);
xor XOR2 (N24737, N24729, N4109);
not NOT1 (N24738, N24712);
not NOT1 (N24739, N24725);
not NOT1 (N24740, N24736);
and AND4 (N24741, N24737, N8687, N22865, N9122);
buf BUF1 (N24742, N24727);
buf BUF1 (N24743, N24738);
nor NOR4 (N24744, N24741, N20960, N24718, N7074);
and AND4 (N24745, N24723, N15449, N5535, N2965);
nand NAND2 (N24746, N24745, N8437);
buf BUF1 (N24747, N24742);
not NOT1 (N24748, N24740);
buf BUF1 (N24749, N24732);
and AND2 (N24750, N24747, N15962);
xor XOR2 (N24751, N24735, N8272);
nor NOR4 (N24752, N24733, N18043, N12651, N9243);
nor NOR3 (N24753, N24752, N9575, N1572);
nand NAND2 (N24754, N24748, N4728);
nand NAND2 (N24755, N24749, N4361);
nand NAND4 (N24756, N24739, N23100, N23911, N10996);
nand NAND2 (N24757, N24751, N5548);
nor NOR2 (N24758, N24757, N3769);
and AND4 (N24759, N24753, N8016, N17578, N17758);
and AND2 (N24760, N24756, N906);
or OR2 (N24761, N24746, N11038);
nor NOR4 (N24762, N24761, N470, N2903, N8530);
buf BUF1 (N24763, N24743);
nand NAND3 (N24764, N24754, N4309, N9944);
nor NOR3 (N24765, N24721, N7796, N20964);
nor NOR4 (N24766, N24763, N7666, N3836, N1919);
or OR4 (N24767, N24755, N20995, N2845, N21037);
nor NOR4 (N24768, N24765, N14721, N18199, N21054);
and AND2 (N24769, N24764, N2373);
nor NOR3 (N24770, N24762, N7889, N20916);
buf BUF1 (N24771, N24769);
nand NAND3 (N24772, N24770, N11102, N3259);
or OR2 (N24773, N24772, N17405);
and AND4 (N24774, N24767, N6711, N12800, N9662);
not NOT1 (N24775, N24771);
nand NAND3 (N24776, N24774, N9408, N15585);
xor XOR2 (N24777, N24773, N726);
nor NOR4 (N24778, N24777, N16827, N16160, N12059);
nand NAND2 (N24779, N24744, N2356);
or OR2 (N24780, N24750, N134);
and AND3 (N24781, N24780, N3195, N24691);
xor XOR2 (N24782, N24768, N201);
and AND2 (N24783, N24781, N3508);
and AND3 (N24784, N24779, N13656, N18660);
and AND3 (N24785, N24783, N1014, N14896);
buf BUF1 (N24786, N24784);
xor XOR2 (N24787, N24778, N2832);
nor NOR2 (N24788, N24760, N19505);
nor NOR2 (N24789, N24758, N9034);
xor XOR2 (N24790, N24788, N9603);
buf BUF1 (N24791, N24789);
and AND3 (N24792, N24791, N6732, N5755);
and AND3 (N24793, N24786, N14205, N14990);
buf BUF1 (N24794, N24776);
or OR2 (N24795, N24792, N21208);
or OR4 (N24796, N24795, N24788, N412, N10566);
not NOT1 (N24797, N24796);
and AND3 (N24798, N24797, N2840, N12904);
xor XOR2 (N24799, N24759, N8137);
nor NOR2 (N24800, N24782, N15957);
or OR4 (N24801, N24785, N13698, N21839, N11356);
not NOT1 (N24802, N24790);
and AND4 (N24803, N24794, N2723, N12564, N7888);
nor NOR4 (N24804, N24799, N21591, N23240, N4367);
or OR4 (N24805, N24787, N6917, N21645, N6283);
not NOT1 (N24806, N24803);
not NOT1 (N24807, N24804);
xor XOR2 (N24808, N24793, N6777);
buf BUF1 (N24809, N24806);
nor NOR4 (N24810, N24766, N19056, N11, N6638);
not NOT1 (N24811, N24807);
buf BUF1 (N24812, N24809);
not NOT1 (N24813, N24810);
or OR3 (N24814, N24800, N15193, N19520);
and AND4 (N24815, N24775, N20601, N21441, N13078);
xor XOR2 (N24816, N24811, N4043);
nor NOR3 (N24817, N24812, N10363, N23525);
or OR2 (N24818, N24813, N24234);
not NOT1 (N24819, N24818);
nor NOR2 (N24820, N24816, N20880);
nand NAND3 (N24821, N24802, N15330, N4029);
buf BUF1 (N24822, N24817);
not NOT1 (N24823, N24808);
and AND2 (N24824, N24801, N6733);
not NOT1 (N24825, N24822);
xor XOR2 (N24826, N24815, N4028);
buf BUF1 (N24827, N24821);
or OR4 (N24828, N24798, N9087, N21212, N4945);
buf BUF1 (N24829, N24825);
nand NAND2 (N24830, N24829, N17570);
buf BUF1 (N24831, N24830);
buf BUF1 (N24832, N24824);
nand NAND2 (N24833, N24819, N23797);
nand NAND2 (N24834, N24805, N22525);
nand NAND4 (N24835, N24814, N22893, N22811, N12030);
xor XOR2 (N24836, N24833, N3326);
nor NOR4 (N24837, N24823, N9205, N21418, N24430);
or OR2 (N24838, N24831, N16555);
or OR4 (N24839, N24832, N3568, N8567, N1601);
not NOT1 (N24840, N24835);
xor XOR2 (N24841, N24839, N17191);
buf BUF1 (N24842, N24828);
nand NAND4 (N24843, N24826, N17450, N9250, N12586);
nor NOR3 (N24844, N24836, N6242, N14264);
nor NOR4 (N24845, N24820, N7138, N1153, N1334);
not NOT1 (N24846, N24834);
or OR4 (N24847, N24846, N9398, N12479, N13075);
buf BUF1 (N24848, N24838);
and AND3 (N24849, N24848, N3233, N4578);
and AND4 (N24850, N24841, N16918, N1941, N13025);
buf BUF1 (N24851, N24844);
buf BUF1 (N24852, N24845);
and AND4 (N24853, N24850, N4215, N11045, N4177);
nand NAND3 (N24854, N24849, N18250, N13853);
and AND2 (N24855, N24843, N23680);
nand NAND2 (N24856, N24854, N4298);
or OR2 (N24857, N24827, N23558);
and AND4 (N24858, N24852, N6322, N15709, N20895);
xor XOR2 (N24859, N24837, N24397);
and AND2 (N24860, N24858, N6068);
xor XOR2 (N24861, N24860, N4496);
and AND2 (N24862, N24861, N7469);
or OR2 (N24863, N24859, N13056);
xor XOR2 (N24864, N24862, N23629);
nor NOR4 (N24865, N24853, N24573, N19780, N938);
buf BUF1 (N24866, N24855);
xor XOR2 (N24867, N24865, N15562);
not NOT1 (N24868, N24864);
and AND3 (N24869, N24856, N2677, N23573);
and AND3 (N24870, N24868, N12685, N2247);
xor XOR2 (N24871, N24866, N11023);
not NOT1 (N24872, N24851);
and AND2 (N24873, N24857, N1382);
or OR4 (N24874, N24842, N21342, N1359, N2969);
and AND3 (N24875, N24840, N19757, N2717);
xor XOR2 (N24876, N24863, N15710);
nand NAND3 (N24877, N24874, N5448, N13437);
or OR4 (N24878, N24873, N559, N24460, N14413);
not NOT1 (N24879, N24867);
or OR3 (N24880, N24876, N949, N15265);
buf BUF1 (N24881, N24880);
nor NOR3 (N24882, N24869, N13901, N24379);
or OR2 (N24883, N24875, N85);
nor NOR3 (N24884, N24870, N19299, N5499);
not NOT1 (N24885, N24877);
and AND4 (N24886, N24885, N12188, N22169, N18899);
xor XOR2 (N24887, N24883, N12578);
not NOT1 (N24888, N24847);
xor XOR2 (N24889, N24871, N5468);
xor XOR2 (N24890, N24884, N8889);
buf BUF1 (N24891, N24879);
or OR2 (N24892, N24878, N24836);
xor XOR2 (N24893, N24872, N20594);
or OR4 (N24894, N24890, N13959, N3675, N20966);
and AND4 (N24895, N24891, N24210, N21127, N21514);
not NOT1 (N24896, N24887);
nand NAND3 (N24897, N24881, N15099, N15914);
nor NOR4 (N24898, N24893, N17320, N11142, N21461);
xor XOR2 (N24899, N24894, N7271);
nand NAND2 (N24900, N24889, N23921);
buf BUF1 (N24901, N24898);
and AND4 (N24902, N24897, N4638, N826, N18359);
nor NOR3 (N24903, N24888, N18496, N1320);
nor NOR2 (N24904, N24900, N4876);
not NOT1 (N24905, N24896);
xor XOR2 (N24906, N24902, N23223);
not NOT1 (N24907, N24906);
nand NAND4 (N24908, N24903, N18821, N11885, N8054);
and AND3 (N24909, N24901, N10113, N23636);
or OR2 (N24910, N24899, N23824);
xor XOR2 (N24911, N24892, N11192);
and AND2 (N24912, N24911, N7642);
or OR2 (N24913, N24895, N6470);
not NOT1 (N24914, N24905);
buf BUF1 (N24915, N24914);
or OR3 (N24916, N24886, N8791, N9329);
or OR2 (N24917, N24882, N8651);
xor XOR2 (N24918, N24917, N14511);
or OR4 (N24919, N24913, N7943, N9368, N19338);
and AND2 (N24920, N24919, N24885);
xor XOR2 (N24921, N24907, N10940);
and AND3 (N24922, N24916, N19835, N16675);
not NOT1 (N24923, N24922);
and AND4 (N24924, N24904, N11454, N4406, N17449);
and AND3 (N24925, N24920, N12148, N19909);
nand NAND3 (N24926, N24908, N19900, N14490);
xor XOR2 (N24927, N24924, N9194);
xor XOR2 (N24928, N24915, N14060);
xor XOR2 (N24929, N24927, N9283);
or OR2 (N24930, N24912, N1900);
buf BUF1 (N24931, N24929);
and AND2 (N24932, N24910, N8351);
buf BUF1 (N24933, N24931);
nor NOR4 (N24934, N24928, N2112, N5454, N22589);
or OR4 (N24935, N24930, N19072, N10172, N9442);
xor XOR2 (N24936, N24921, N5039);
not NOT1 (N24937, N24936);
xor XOR2 (N24938, N24934, N22855);
nand NAND2 (N24939, N24933, N3060);
or OR4 (N24940, N24923, N23031, N7611, N24790);
and AND4 (N24941, N24935, N10262, N12696, N17779);
buf BUF1 (N24942, N24941);
and AND4 (N24943, N24937, N5314, N17048, N5611);
not NOT1 (N24944, N24909);
nor NOR2 (N24945, N24926, N4504);
nand NAND2 (N24946, N24932, N10286);
nand NAND4 (N24947, N24945, N24524, N12760, N19429);
or OR2 (N24948, N24918, N24271);
xor XOR2 (N24949, N24946, N23829);
not NOT1 (N24950, N24939);
buf BUF1 (N24951, N24947);
xor XOR2 (N24952, N24942, N7432);
buf BUF1 (N24953, N24925);
buf BUF1 (N24954, N24938);
or OR3 (N24955, N24950, N9000, N18286);
and AND4 (N24956, N24952, N9885, N11033, N21871);
buf BUF1 (N24957, N24956);
or OR2 (N24958, N24954, N8815);
xor XOR2 (N24959, N24953, N18316);
not NOT1 (N24960, N24955);
xor XOR2 (N24961, N24943, N13691);
nor NOR4 (N24962, N24961, N15282, N3299, N18525);
xor XOR2 (N24963, N24951, N8125);
nand NAND2 (N24964, N24958, N3849);
and AND3 (N24965, N24944, N3315, N7736);
or OR2 (N24966, N24965, N22374);
not NOT1 (N24967, N24962);
xor XOR2 (N24968, N24948, N12797);
not NOT1 (N24969, N24966);
or OR2 (N24970, N24969, N19368);
buf BUF1 (N24971, N24959);
and AND3 (N24972, N24971, N10274, N22716);
nand NAND2 (N24973, N24940, N4435);
or OR4 (N24974, N24967, N14573, N2479, N8726);
buf BUF1 (N24975, N24964);
nor NOR3 (N24976, N24949, N22892, N24335);
and AND4 (N24977, N24963, N4907, N21075, N1336);
xor XOR2 (N24978, N24972, N4326);
xor XOR2 (N24979, N24975, N5483);
or OR2 (N24980, N24978, N5332);
not NOT1 (N24981, N24960);
nand NAND4 (N24982, N24970, N12140, N15174, N11160);
nor NOR4 (N24983, N24981, N22501, N18985, N21588);
buf BUF1 (N24984, N24982);
or OR4 (N24985, N24984, N24886, N24643, N6777);
or OR4 (N24986, N24977, N5481, N11889, N3925);
and AND3 (N24987, N24985, N9307, N9835);
or OR2 (N24988, N24987, N14602);
nand NAND4 (N24989, N24979, N11426, N11791, N7966);
or OR2 (N24990, N24989, N22897);
xor XOR2 (N24991, N24980, N1610);
nand NAND4 (N24992, N24986, N3988, N3174, N1940);
nand NAND4 (N24993, N24974, N2204, N9839, N15789);
nand NAND4 (N24994, N24993, N10423, N13940, N4978);
not NOT1 (N24995, N24992);
nor NOR3 (N24996, N24968, N9805, N16027);
not NOT1 (N24997, N24957);
nand NAND4 (N24998, N24996, N17919, N895, N21825);
or OR2 (N24999, N24998, N12585);
xor XOR2 (N25000, N24997, N3188);
xor XOR2 (N25001, N24995, N16833);
not NOT1 (N25002, N24973);
xor XOR2 (N25003, N24988, N23629);
and AND3 (N25004, N25002, N7634, N10332);
xor XOR2 (N25005, N25001, N4004);
not NOT1 (N25006, N24991);
buf BUF1 (N25007, N25003);
and AND3 (N25008, N25007, N18362, N8162);
buf BUF1 (N25009, N25000);
buf BUF1 (N25010, N25008);
and AND2 (N25011, N24983, N19533);
or OR3 (N25012, N24994, N19647, N16681);
and AND4 (N25013, N25010, N19687, N14405, N12405);
nor NOR2 (N25014, N25005, N19742);
xor XOR2 (N25015, N25014, N21310);
buf BUF1 (N25016, N24976);
nand NAND4 (N25017, N25006, N14994, N8196, N13969);
nor NOR2 (N25018, N25016, N7092);
buf BUF1 (N25019, N25017);
not NOT1 (N25020, N25012);
nor NOR3 (N25021, N25013, N11372, N24898);
and AND3 (N25022, N25021, N23292, N19306);
and AND2 (N25023, N25019, N8102);
nand NAND2 (N25024, N25018, N9656);
xor XOR2 (N25025, N25011, N14340);
or OR4 (N25026, N25022, N22393, N11262, N851);
and AND2 (N25027, N25023, N10956);
xor XOR2 (N25028, N25025, N24730);
or OR2 (N25029, N25015, N13098);
and AND3 (N25030, N24999, N19473, N2261);
xor XOR2 (N25031, N25020, N16396);
buf BUF1 (N25032, N25026);
buf BUF1 (N25033, N25024);
not NOT1 (N25034, N25032);
nand NAND4 (N25035, N25004, N20064, N23514, N10867);
nor NOR4 (N25036, N25035, N21940, N2706, N22638);
nor NOR4 (N25037, N25027, N8857, N20197, N22995);
nor NOR3 (N25038, N25036, N2888, N6904);
not NOT1 (N25039, N25034);
or OR4 (N25040, N25030, N19827, N23063, N14030);
nand NAND3 (N25041, N25029, N24842, N20145);
nand NAND2 (N25042, N24990, N14154);
or OR2 (N25043, N25037, N4904);
buf BUF1 (N25044, N25042);
buf BUF1 (N25045, N25039);
buf BUF1 (N25046, N25045);
or OR4 (N25047, N25033, N22849, N7442, N5379);
buf BUF1 (N25048, N25046);
nor NOR3 (N25049, N25041, N16981, N3974);
and AND2 (N25050, N25038, N14747);
buf BUF1 (N25051, N25043);
xor XOR2 (N25052, N25051, N9981);
xor XOR2 (N25053, N25044, N21495);
buf BUF1 (N25054, N25049);
nor NOR3 (N25055, N25053, N16217, N21119);
xor XOR2 (N25056, N25048, N11414);
buf BUF1 (N25057, N25054);
xor XOR2 (N25058, N25031, N6941);
xor XOR2 (N25059, N25056, N21767);
or OR2 (N25060, N25047, N17244);
not NOT1 (N25061, N25009);
buf BUF1 (N25062, N25060);
nor NOR4 (N25063, N25052, N11769, N24306, N22847);
nor NOR2 (N25064, N25028, N15433);
buf BUF1 (N25065, N25064);
buf BUF1 (N25066, N25040);
nand NAND3 (N25067, N25059, N24854, N18508);
nor NOR3 (N25068, N25061, N20177, N6077);
not NOT1 (N25069, N25062);
nand NAND3 (N25070, N25069, N11521, N8457);
xor XOR2 (N25071, N25050, N5350);
nand NAND3 (N25072, N25058, N18782, N923);
nor NOR3 (N25073, N25067, N20171, N7508);
nor NOR2 (N25074, N25063, N10772);
buf BUF1 (N25075, N25072);
nand NAND4 (N25076, N25066, N490, N18759, N9842);
nand NAND2 (N25077, N25074, N21158);
or OR2 (N25078, N25073, N24681);
buf BUF1 (N25079, N25078);
nand NAND4 (N25080, N25057, N13480, N1406, N2595);
xor XOR2 (N25081, N25070, N17882);
and AND4 (N25082, N25081, N24779, N12739, N775);
buf BUF1 (N25083, N25065);
or OR4 (N25084, N25082, N4053, N24672, N18419);
nor NOR4 (N25085, N25080, N16384, N2058, N11982);
or OR3 (N25086, N25055, N18752, N1937);
and AND2 (N25087, N25084, N4441);
and AND2 (N25088, N25071, N4914);
nor NOR3 (N25089, N25075, N24407, N387);
not NOT1 (N25090, N25077);
and AND2 (N25091, N25079, N4858);
and AND2 (N25092, N25076, N11085);
nand NAND3 (N25093, N25068, N5080, N14839);
buf BUF1 (N25094, N25090);
nor NOR3 (N25095, N25087, N13022, N9219);
nand NAND3 (N25096, N25089, N12456, N17823);
buf BUF1 (N25097, N25095);
nor NOR3 (N25098, N25083, N2012, N8527);
not NOT1 (N25099, N25085);
nor NOR2 (N25100, N25094, N23767);
buf BUF1 (N25101, N25088);
buf BUF1 (N25102, N25100);
buf BUF1 (N25103, N25096);
buf BUF1 (N25104, N25097);
and AND3 (N25105, N25093, N10829, N21423);
xor XOR2 (N25106, N25105, N9960);
buf BUF1 (N25107, N25099);
nor NOR2 (N25108, N25091, N20634);
nand NAND3 (N25109, N25102, N18610, N8390);
or OR4 (N25110, N25107, N12047, N22868, N24845);
nor NOR2 (N25111, N25101, N12541);
buf BUF1 (N25112, N25111);
nand NAND2 (N25113, N25109, N3502);
or OR3 (N25114, N25113, N302, N8493);
and AND4 (N25115, N25092, N23564, N10117, N2468);
not NOT1 (N25116, N25112);
and AND4 (N25117, N25086, N14275, N15517, N13473);
not NOT1 (N25118, N25116);
or OR2 (N25119, N25098, N19576);
or OR3 (N25120, N25119, N22464, N23986);
nand NAND4 (N25121, N25118, N15311, N2220, N7490);
nand NAND3 (N25122, N25117, N4223, N2274);
xor XOR2 (N25123, N25115, N12009);
nand NAND3 (N25124, N25106, N13141, N6688);
xor XOR2 (N25125, N25110, N9999);
not NOT1 (N25126, N25125);
or OR2 (N25127, N25108, N18144);
nand NAND3 (N25128, N25104, N19611, N6539);
xor XOR2 (N25129, N25103, N5371);
xor XOR2 (N25130, N25114, N12788);
not NOT1 (N25131, N25120);
nor NOR3 (N25132, N25121, N23127, N7525);
or OR2 (N25133, N25129, N17880);
and AND4 (N25134, N25123, N1952, N21764, N13801);
not NOT1 (N25135, N25133);
nand NAND2 (N25136, N25135, N19675);
buf BUF1 (N25137, N25136);
or OR4 (N25138, N25128, N2019, N5356, N8341);
and AND2 (N25139, N25130, N4626);
xor XOR2 (N25140, N25127, N19902);
buf BUF1 (N25141, N25134);
not NOT1 (N25142, N25132);
nand NAND2 (N25143, N25140, N17282);
nand NAND3 (N25144, N25138, N17354, N11520);
or OR4 (N25145, N25144, N18655, N6532, N16251);
nor NOR2 (N25146, N25139, N6456);
buf BUF1 (N25147, N25142);
or OR3 (N25148, N25145, N22074, N14768);
not NOT1 (N25149, N25131);
nand NAND2 (N25150, N25148, N10072);
and AND4 (N25151, N25141, N8767, N15432, N2793);
xor XOR2 (N25152, N25124, N19845);
or OR4 (N25153, N25147, N7309, N22930, N21294);
and AND3 (N25154, N25146, N24400, N6524);
or OR2 (N25155, N25122, N10508);
nand NAND4 (N25156, N25155, N887, N18001, N18084);
nor NOR4 (N25157, N25152, N11589, N17444, N20092);
not NOT1 (N25158, N25157);
buf BUF1 (N25159, N25149);
buf BUF1 (N25160, N25159);
not NOT1 (N25161, N25160);
nor NOR4 (N25162, N25151, N24949, N1911, N20343);
and AND4 (N25163, N25126, N20502, N5036, N8073);
nor NOR3 (N25164, N25153, N23742, N11599);
or OR2 (N25165, N25150, N14998);
xor XOR2 (N25166, N25158, N10678);
buf BUF1 (N25167, N25162);
nand NAND2 (N25168, N25166, N23773);
xor XOR2 (N25169, N25163, N4392);
nor NOR2 (N25170, N25164, N19221);
or OR4 (N25171, N25161, N2858, N21524, N10992);
nor NOR4 (N25172, N25170, N5435, N23014, N20793);
not NOT1 (N25173, N25165);
and AND4 (N25174, N25168, N6605, N23558, N1240);
and AND4 (N25175, N25169, N19932, N2311, N2880);
or OR2 (N25176, N25173, N947);
or OR3 (N25177, N25137, N17921, N8638);
or OR2 (N25178, N25154, N14793);
not NOT1 (N25179, N25175);
buf BUF1 (N25180, N25156);
not NOT1 (N25181, N25176);
nor NOR2 (N25182, N25171, N21090);
or OR2 (N25183, N25180, N20158);
nor NOR3 (N25184, N25174, N5056, N1981);
nand NAND3 (N25185, N25183, N22643, N18125);
or OR4 (N25186, N25178, N6197, N6898, N2386);
not NOT1 (N25187, N25184);
not NOT1 (N25188, N25177);
not NOT1 (N25189, N25186);
nand NAND4 (N25190, N25167, N12296, N17550, N19097);
nand NAND4 (N25191, N25188, N16242, N13062, N16918);
not NOT1 (N25192, N25187);
or OR2 (N25193, N25181, N23021);
or OR3 (N25194, N25190, N18696, N16173);
nand NAND4 (N25195, N25189, N3634, N1120, N6667);
nand NAND3 (N25196, N25191, N23743, N7362);
nor NOR3 (N25197, N25194, N17019, N16902);
and AND4 (N25198, N25143, N18125, N19292, N10878);
not NOT1 (N25199, N25182);
nand NAND3 (N25200, N25185, N4372, N4008);
or OR4 (N25201, N25192, N20698, N14156, N8462);
not NOT1 (N25202, N25196);
nor NOR4 (N25203, N25202, N24129, N16826, N6255);
nor NOR3 (N25204, N25195, N18981, N10422);
xor XOR2 (N25205, N25200, N14327);
buf BUF1 (N25206, N25198);
or OR3 (N25207, N25205, N10629, N19925);
xor XOR2 (N25208, N25179, N761);
nand NAND3 (N25209, N25172, N7111, N6535);
buf BUF1 (N25210, N25207);
nand NAND2 (N25211, N25204, N24628);
xor XOR2 (N25212, N25206, N17900);
buf BUF1 (N25213, N25201);
nor NOR2 (N25214, N25212, N17209);
xor XOR2 (N25215, N25199, N8829);
nor NOR2 (N25216, N25197, N15999);
not NOT1 (N25217, N25213);
nand NAND3 (N25218, N25216, N21737, N9679);
buf BUF1 (N25219, N25218);
buf BUF1 (N25220, N25217);
and AND3 (N25221, N25211, N22527, N20998);
buf BUF1 (N25222, N25220);
xor XOR2 (N25223, N25219, N21493);
not NOT1 (N25224, N25221);
nor NOR3 (N25225, N25209, N21030, N15586);
not NOT1 (N25226, N25208);
not NOT1 (N25227, N25210);
or OR4 (N25228, N25214, N12060, N2982, N24750);
xor XOR2 (N25229, N25215, N22582);
or OR4 (N25230, N25203, N4877, N3970, N12415);
nor NOR3 (N25231, N25229, N8626, N20517);
buf BUF1 (N25232, N25228);
and AND4 (N25233, N25226, N21132, N486, N24434);
xor XOR2 (N25234, N25222, N8578);
nand NAND4 (N25235, N25231, N24511, N17835, N18926);
not NOT1 (N25236, N25235);
buf BUF1 (N25237, N25236);
nor NOR2 (N25238, N25237, N10331);
nand NAND4 (N25239, N25227, N6790, N10281, N10676);
or OR2 (N25240, N25238, N13438);
nand NAND3 (N25241, N25224, N1300, N15231);
xor XOR2 (N25242, N25193, N2459);
buf BUF1 (N25243, N25223);
nor NOR2 (N25244, N25239, N10276);
nand NAND3 (N25245, N25225, N6102, N7337);
nand NAND3 (N25246, N25234, N22512, N5960);
nor NOR2 (N25247, N25232, N8664);
not NOT1 (N25248, N25243);
or OR3 (N25249, N25242, N9516, N23285);
buf BUF1 (N25250, N25249);
nand NAND3 (N25251, N25247, N8239, N5556);
nand NAND2 (N25252, N25248, N10878);
xor XOR2 (N25253, N25251, N12564);
nand NAND3 (N25254, N25246, N6771, N6229);
buf BUF1 (N25255, N25245);
nor NOR2 (N25256, N25244, N9112);
buf BUF1 (N25257, N25240);
not NOT1 (N25258, N25254);
not NOT1 (N25259, N25233);
buf BUF1 (N25260, N25259);
or OR4 (N25261, N25257, N11308, N9516, N24884);
nor NOR2 (N25262, N25253, N21943);
buf BUF1 (N25263, N25250);
buf BUF1 (N25264, N25260);
nand NAND3 (N25265, N25230, N5615, N7203);
buf BUF1 (N25266, N25255);
nor NOR3 (N25267, N25262, N83, N11719);
or OR4 (N25268, N25258, N6402, N24330, N3489);
xor XOR2 (N25269, N25266, N10543);
nor NOR4 (N25270, N25261, N4825, N22614, N19195);
buf BUF1 (N25271, N25268);
nand NAND4 (N25272, N25263, N18296, N1037, N3671);
or OR4 (N25273, N25241, N8311, N18955, N9202);
xor XOR2 (N25274, N25273, N1956);
nand NAND2 (N25275, N25270, N12324);
nand NAND4 (N25276, N25271, N11228, N12305, N2078);
nand NAND3 (N25277, N25265, N24484, N3897);
xor XOR2 (N25278, N25256, N17995);
or OR2 (N25279, N25272, N1367);
and AND3 (N25280, N25275, N11827, N12161);
buf BUF1 (N25281, N25280);
nor NOR3 (N25282, N25278, N3450, N7962);
or OR3 (N25283, N25252, N3712, N4118);
xor XOR2 (N25284, N25276, N15334);
not NOT1 (N25285, N25281);
buf BUF1 (N25286, N25267);
xor XOR2 (N25287, N25285, N8758);
not NOT1 (N25288, N25279);
xor XOR2 (N25289, N25283, N15633);
and AND3 (N25290, N25277, N5661, N6070);
not NOT1 (N25291, N25286);
nand NAND4 (N25292, N25282, N22257, N21816, N1568);
xor XOR2 (N25293, N25264, N20089);
nand NAND2 (N25294, N25274, N2331);
xor XOR2 (N25295, N25289, N12467);
or OR3 (N25296, N25292, N23174, N18331);
nand NAND2 (N25297, N25291, N23815);
xor XOR2 (N25298, N25287, N5236);
and AND2 (N25299, N25290, N9946);
xor XOR2 (N25300, N25284, N2522);
xor XOR2 (N25301, N25293, N18778);
and AND3 (N25302, N25294, N11320, N24310);
or OR4 (N25303, N25269, N19418, N3918, N8428);
nor NOR4 (N25304, N25302, N7098, N8921, N9328);
buf BUF1 (N25305, N25299);
or OR4 (N25306, N25288, N9312, N21111, N4873);
nand NAND2 (N25307, N25301, N1476);
nand NAND2 (N25308, N25298, N19692);
or OR3 (N25309, N25308, N6679, N10882);
not NOT1 (N25310, N25303);
nand NAND2 (N25311, N25297, N15803);
and AND2 (N25312, N25306, N8550);
nor NOR2 (N25313, N25311, N12137);
and AND4 (N25314, N25307, N16445, N23517, N8924);
nor NOR2 (N25315, N25304, N21644);
xor XOR2 (N25316, N25312, N6204);
not NOT1 (N25317, N25296);
nor NOR3 (N25318, N25310, N19132, N767);
xor XOR2 (N25319, N25317, N8601);
not NOT1 (N25320, N25313);
xor XOR2 (N25321, N25309, N18436);
xor XOR2 (N25322, N25319, N15518);
xor XOR2 (N25323, N25305, N14689);
nand NAND2 (N25324, N25322, N22034);
and AND3 (N25325, N25314, N10356, N15577);
and AND2 (N25326, N25323, N24330);
nor NOR2 (N25327, N25321, N12741);
not NOT1 (N25328, N25325);
nor NOR2 (N25329, N25295, N11972);
buf BUF1 (N25330, N25329);
nand NAND2 (N25331, N25330, N19533);
nor NOR3 (N25332, N25320, N9358, N786);
buf BUF1 (N25333, N25316);
and AND3 (N25334, N25331, N144, N9435);
nor NOR4 (N25335, N25315, N4546, N1197, N1657);
buf BUF1 (N25336, N25328);
xor XOR2 (N25337, N25326, N4210);
not NOT1 (N25338, N25337);
nor NOR2 (N25339, N25334, N19479);
nand NAND4 (N25340, N25339, N22098, N10326, N10024);
not NOT1 (N25341, N25333);
buf BUF1 (N25342, N25318);
buf BUF1 (N25343, N25327);
nand NAND4 (N25344, N25342, N13511, N11958, N9786);
or OR3 (N25345, N25332, N21662, N4711);
not NOT1 (N25346, N25300);
and AND2 (N25347, N25324, N22351);
or OR4 (N25348, N25344, N10662, N9547, N14332);
nand NAND3 (N25349, N25335, N2263, N6845);
nor NOR2 (N25350, N25341, N14174);
buf BUF1 (N25351, N25348);
or OR2 (N25352, N25346, N14499);
xor XOR2 (N25353, N25336, N21698);
buf BUF1 (N25354, N25338);
nor NOR4 (N25355, N25351, N18897, N11479, N15222);
buf BUF1 (N25356, N25345);
buf BUF1 (N25357, N25356);
xor XOR2 (N25358, N25352, N15607);
nor NOR3 (N25359, N25343, N18923, N17934);
or OR3 (N25360, N25347, N13312, N21964);
or OR3 (N25361, N25355, N1691, N17233);
nand NAND2 (N25362, N25357, N17232);
and AND4 (N25363, N25350, N11869, N12541, N10837);
nor NOR2 (N25364, N25359, N17224);
and AND2 (N25365, N25349, N24423);
or OR2 (N25366, N25362, N8366);
nor NOR2 (N25367, N25353, N1950);
nor NOR4 (N25368, N25340, N3922, N18091, N9474);
or OR4 (N25369, N25363, N14576, N22237, N23315);
xor XOR2 (N25370, N25361, N19832);
and AND3 (N25371, N25369, N11718, N18719);
nand NAND2 (N25372, N25365, N17435);
xor XOR2 (N25373, N25371, N19233);
not NOT1 (N25374, N25364);
and AND2 (N25375, N25358, N8181);
xor XOR2 (N25376, N25354, N21843);
not NOT1 (N25377, N25374);
buf BUF1 (N25378, N25372);
nand NAND3 (N25379, N25373, N403, N18702);
or OR4 (N25380, N25367, N11185, N5578, N10897);
nor NOR2 (N25381, N25368, N2100);
buf BUF1 (N25382, N25380);
or OR4 (N25383, N25378, N4256, N5007, N21708);
and AND4 (N25384, N25366, N13624, N13139, N13403);
buf BUF1 (N25385, N25384);
or OR3 (N25386, N25381, N23714, N14141);
and AND4 (N25387, N25379, N6136, N22261, N24504);
nand NAND2 (N25388, N25386, N6816);
and AND4 (N25389, N25360, N3041, N72, N9877);
buf BUF1 (N25390, N25375);
or OR2 (N25391, N25376, N12023);
nand NAND2 (N25392, N25370, N3447);
and AND2 (N25393, N25392, N23916);
buf BUF1 (N25394, N25383);
buf BUF1 (N25395, N25382);
xor XOR2 (N25396, N25377, N3343);
and AND2 (N25397, N25385, N1453);
nor NOR2 (N25398, N25395, N21407);
and AND4 (N25399, N25396, N23761, N13293, N21092);
nand NAND2 (N25400, N25397, N21723);
or OR2 (N25401, N25394, N22769);
nand NAND3 (N25402, N25393, N17720, N21639);
nor NOR2 (N25403, N25402, N22382);
nor NOR2 (N25404, N25390, N15951);
or OR3 (N25405, N25387, N13288, N17757);
not NOT1 (N25406, N25389);
and AND4 (N25407, N25401, N6516, N22129, N24823);
and AND2 (N25408, N25399, N24789);
nand NAND3 (N25409, N25388, N2997, N4095);
and AND2 (N25410, N25403, N16468);
and AND2 (N25411, N25406, N19578);
or OR3 (N25412, N25391, N17448, N12749);
not NOT1 (N25413, N25405);
not NOT1 (N25414, N25400);
nor NOR2 (N25415, N25409, N18540);
buf BUF1 (N25416, N25408);
or OR4 (N25417, N25411, N14211, N11019, N9266);
nand NAND4 (N25418, N25412, N21446, N7364, N22188);
xor XOR2 (N25419, N25415, N561);
and AND2 (N25420, N25407, N15219);
or OR3 (N25421, N25417, N13343, N17225);
not NOT1 (N25422, N25410);
nor NOR2 (N25423, N25413, N7359);
not NOT1 (N25424, N25420);
nor NOR4 (N25425, N25421, N20381, N4298, N16644);
buf BUF1 (N25426, N25414);
buf BUF1 (N25427, N25425);
buf BUF1 (N25428, N25419);
and AND2 (N25429, N25422, N20772);
nor NOR2 (N25430, N25398, N7616);
or OR4 (N25431, N25426, N17784, N10006, N20836);
nor NOR3 (N25432, N25431, N22598, N2903);
xor XOR2 (N25433, N25429, N21049);
or OR2 (N25434, N25416, N6036);
buf BUF1 (N25435, N25432);
buf BUF1 (N25436, N25424);
xor XOR2 (N25437, N25433, N7556);
not NOT1 (N25438, N25435);
not NOT1 (N25439, N25437);
or OR2 (N25440, N25427, N12587);
xor XOR2 (N25441, N25418, N13809);
nor NOR4 (N25442, N25436, N9438, N21753, N25226);
and AND3 (N25443, N25440, N4343, N14269);
nand NAND2 (N25444, N25441, N12477);
or OR3 (N25445, N25444, N23576, N22605);
not NOT1 (N25446, N25434);
nor NOR2 (N25447, N25428, N20204);
not NOT1 (N25448, N25447);
xor XOR2 (N25449, N25404, N1863);
or OR2 (N25450, N25423, N20857);
buf BUF1 (N25451, N25450);
nor NOR2 (N25452, N25446, N69);
or OR4 (N25453, N25442, N15207, N4132, N10965);
not NOT1 (N25454, N25452);
buf BUF1 (N25455, N25439);
buf BUF1 (N25456, N25443);
or OR2 (N25457, N25438, N25015);
xor XOR2 (N25458, N25445, N869);
not NOT1 (N25459, N25448);
or OR3 (N25460, N25449, N23642, N24474);
buf BUF1 (N25461, N25459);
nand NAND3 (N25462, N25454, N15565, N12194);
and AND2 (N25463, N25457, N11597);
and AND3 (N25464, N25458, N5313, N18168);
nor NOR4 (N25465, N25451, N24168, N15109, N19423);
xor XOR2 (N25466, N25462, N18570);
buf BUF1 (N25467, N25456);
or OR2 (N25468, N25463, N23627);
not NOT1 (N25469, N25464);
xor XOR2 (N25470, N25461, N9145);
nand NAND2 (N25471, N25469, N17376);
nand NAND4 (N25472, N25470, N934, N20650, N1439);
xor XOR2 (N25473, N25467, N3969);
xor XOR2 (N25474, N25466, N12177);
nor NOR2 (N25475, N25474, N8753);
or OR4 (N25476, N25430, N17839, N15798, N22985);
nand NAND2 (N25477, N25473, N15969);
and AND3 (N25478, N25465, N2157, N3502);
nor NOR3 (N25479, N25460, N6210, N12894);
or OR2 (N25480, N25472, N1824);
or OR2 (N25481, N25453, N2444);
buf BUF1 (N25482, N25479);
or OR3 (N25483, N25482, N18834, N555);
and AND4 (N25484, N25468, N23873, N19422, N8947);
nand NAND3 (N25485, N25478, N14157, N25172);
and AND4 (N25486, N25483, N19358, N18633, N19303);
or OR4 (N25487, N25486, N22531, N3570, N700);
buf BUF1 (N25488, N25471);
xor XOR2 (N25489, N25477, N2817);
xor XOR2 (N25490, N25481, N15102);
nor NOR3 (N25491, N25489, N24936, N6833);
buf BUF1 (N25492, N25455);
not NOT1 (N25493, N25484);
and AND4 (N25494, N25491, N2457, N21823, N1770);
not NOT1 (N25495, N25480);
xor XOR2 (N25496, N25476, N11611);
or OR2 (N25497, N25495, N24307);
not NOT1 (N25498, N25494);
not NOT1 (N25499, N25497);
buf BUF1 (N25500, N25485);
buf BUF1 (N25501, N25499);
or OR3 (N25502, N25487, N17148, N24352);
nand NAND3 (N25503, N25496, N22510, N13518);
and AND3 (N25504, N25500, N8734, N8995);
and AND2 (N25505, N25502, N3281);
not NOT1 (N25506, N25488);
buf BUF1 (N25507, N25503);
nor NOR3 (N25508, N25490, N24493, N6253);
buf BUF1 (N25509, N25493);
not NOT1 (N25510, N25508);
nor NOR2 (N25511, N25510, N5179);
not NOT1 (N25512, N25511);
buf BUF1 (N25513, N25509);
nor NOR4 (N25514, N25504, N2339, N19987, N1989);
and AND3 (N25515, N25501, N2240, N2062);
buf BUF1 (N25516, N25514);
not NOT1 (N25517, N25506);
not NOT1 (N25518, N25513);
and AND3 (N25519, N25475, N22316, N20993);
and AND2 (N25520, N25518, N505);
xor XOR2 (N25521, N25516, N23326);
buf BUF1 (N25522, N25519);
or OR2 (N25523, N25521, N839);
nor NOR2 (N25524, N25515, N11723);
or OR2 (N25525, N25517, N14319);
nor NOR3 (N25526, N25520, N8430, N8345);
not NOT1 (N25527, N25526);
and AND2 (N25528, N25505, N10919);
nand NAND2 (N25529, N25498, N10402);
and AND4 (N25530, N25507, N3541, N20453, N16638);
and AND4 (N25531, N25525, N12187, N10335, N3213);
xor XOR2 (N25532, N25531, N11261);
buf BUF1 (N25533, N25527);
and AND4 (N25534, N25533, N6669, N7446, N3273);
nor NOR2 (N25535, N25530, N10127);
buf BUF1 (N25536, N25529);
or OR4 (N25537, N25522, N7044, N14868, N18854);
nand NAND3 (N25538, N25534, N1144, N25393);
not NOT1 (N25539, N25524);
and AND3 (N25540, N25538, N5367, N21725);
and AND3 (N25541, N25492, N22278, N14107);
xor XOR2 (N25542, N25528, N1877);
nand NAND3 (N25543, N25536, N7328, N5529);
and AND3 (N25544, N25535, N15828, N11596);
nand NAND4 (N25545, N25532, N14147, N17151, N11277);
nor NOR3 (N25546, N25537, N10802, N19847);
nand NAND3 (N25547, N25546, N15242, N11744);
not NOT1 (N25548, N25547);
and AND2 (N25549, N25548, N6638);
buf BUF1 (N25550, N25540);
not NOT1 (N25551, N25523);
buf BUF1 (N25552, N25543);
or OR2 (N25553, N25545, N4381);
xor XOR2 (N25554, N25512, N19251);
nor NOR2 (N25555, N25539, N9520);
buf BUF1 (N25556, N25555);
nand NAND4 (N25557, N25542, N20651, N21538, N13250);
buf BUF1 (N25558, N25556);
nand NAND3 (N25559, N25552, N4195, N21531);
or OR4 (N25560, N25558, N14823, N7740, N22321);
nor NOR3 (N25561, N25541, N18433, N20818);
xor XOR2 (N25562, N25559, N2172);
nor NOR4 (N25563, N25562, N20950, N11566, N8790);
nand NAND2 (N25564, N25561, N1595);
nor NOR4 (N25565, N25544, N97, N7698, N24001);
nand NAND2 (N25566, N25560, N16628);
buf BUF1 (N25567, N25550);
nand NAND3 (N25568, N25563, N4183, N5212);
buf BUF1 (N25569, N25557);
buf BUF1 (N25570, N25567);
nor NOR3 (N25571, N25569, N9954, N12583);
and AND4 (N25572, N25553, N15034, N22554, N9376);
and AND4 (N25573, N25554, N14310, N21028, N24434);
not NOT1 (N25574, N25551);
not NOT1 (N25575, N25549);
and AND4 (N25576, N25574, N21541, N8921, N13815);
not NOT1 (N25577, N25575);
and AND2 (N25578, N25576, N7238);
nand NAND3 (N25579, N25564, N3576, N17927);
xor XOR2 (N25580, N25573, N25082);
buf BUF1 (N25581, N25578);
xor XOR2 (N25582, N25568, N19245);
not NOT1 (N25583, N25580);
or OR2 (N25584, N25572, N10395);
nand NAND3 (N25585, N25571, N4458, N18086);
xor XOR2 (N25586, N25566, N9661);
or OR4 (N25587, N25579, N477, N4386, N3719);
buf BUF1 (N25588, N25570);
and AND4 (N25589, N25585, N13847, N10960, N21552);
xor XOR2 (N25590, N25586, N6202);
nor NOR2 (N25591, N25589, N8989);
nor NOR3 (N25592, N25587, N13493, N11741);
or OR3 (N25593, N25581, N24989, N6180);
buf BUF1 (N25594, N25583);
nor NOR2 (N25595, N25593, N17945);
not NOT1 (N25596, N25588);
nand NAND4 (N25597, N25565, N15705, N13946, N17627);
nor NOR2 (N25598, N25596, N14218);
or OR3 (N25599, N25594, N16067, N18584);
nand NAND4 (N25600, N25577, N13289, N18682, N8119);
and AND2 (N25601, N25598, N10803);
buf BUF1 (N25602, N25592);
xor XOR2 (N25603, N25601, N17983);
or OR3 (N25604, N25582, N18758, N2820);
not NOT1 (N25605, N25591);
and AND3 (N25606, N25590, N18067, N8514);
or OR2 (N25607, N25599, N18121);
or OR4 (N25608, N25605, N5701, N11497, N13846);
nand NAND3 (N25609, N25604, N5156, N3830);
xor XOR2 (N25610, N25600, N20081);
and AND2 (N25611, N25584, N18703);
not NOT1 (N25612, N25602);
not NOT1 (N25613, N25607);
buf BUF1 (N25614, N25609);
not NOT1 (N25615, N25597);
endmodule