// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16;

output N3206,N3212,N3204,N3209,N3205,N3215,N3213,N3214,N3207,N3216;

xor XOR2 (N17, N2, N13);
and AND4 (N18, N15, N7, N1, N13);
xor XOR2 (N19, N13, N13);
not NOT1 (N20, N15);
buf BUF1 (N21, N6);
and AND4 (N22, N12, N19, N7, N7);
not NOT1 (N23, N3);
nor NOR3 (N24, N17, N18, N18);
nand NAND3 (N25, N11, N19, N19);
xor XOR2 (N26, N2, N20);
nor NOR3 (N27, N20, N22, N6);
not NOT1 (N28, N17);
buf BUF1 (N29, N21);
nand NAND2 (N30, N20, N5);
buf BUF1 (N31, N7);
not NOT1 (N32, N7);
xor XOR2 (N33, N27, N21);
and AND2 (N34, N30, N2);
nand NAND4 (N35, N34, N3, N7, N19);
xor XOR2 (N36, N29, N16);
not NOT1 (N37, N35);
and AND4 (N38, N26, N26, N27, N14);
or OR3 (N39, N31, N1, N21);
and AND2 (N40, N33, N33);
and AND2 (N41, N24, N21);
or OR4 (N42, N28, N20, N18, N41);
nand NAND2 (N43, N6, N30);
nor NOR3 (N44, N43, N22, N35);
buf BUF1 (N45, N32);
nand NAND4 (N46, N38, N7, N40, N9);
and AND2 (N47, N6, N28);
not NOT1 (N48, N47);
nor NOR2 (N49, N23, N24);
buf BUF1 (N50, N48);
or OR3 (N51, N50, N28, N5);
or OR3 (N52, N44, N9, N48);
buf BUF1 (N53, N36);
buf BUF1 (N54, N45);
nor NOR2 (N55, N25, N34);
and AND4 (N56, N37, N26, N48, N14);
xor XOR2 (N57, N49, N32);
nand NAND2 (N58, N51, N36);
or OR2 (N59, N54, N11);
or OR2 (N60, N42, N40);
not NOT1 (N61, N58);
buf BUF1 (N62, N53);
not NOT1 (N63, N46);
nor NOR3 (N64, N62, N12, N12);
buf BUF1 (N65, N63);
xor XOR2 (N66, N57, N27);
nor NOR2 (N67, N56, N36);
nor NOR3 (N68, N39, N45, N37);
xor XOR2 (N69, N55, N3);
nand NAND2 (N70, N65, N2);
and AND3 (N71, N52, N36, N37);
xor XOR2 (N72, N60, N37);
nor NOR2 (N73, N68, N7);
nand NAND2 (N74, N70, N31);
and AND3 (N75, N72, N38, N46);
or OR4 (N76, N59, N72, N66, N49);
and AND3 (N77, N19, N73, N65);
or OR2 (N78, N6, N65);
nand NAND4 (N79, N67, N58, N4, N78);
buf BUF1 (N80, N72);
nand NAND4 (N81, N69, N72, N64, N79);
nand NAND2 (N82, N42, N74);
buf BUF1 (N83, N17);
buf BUF1 (N84, N20);
xor XOR2 (N85, N71, N7);
or OR2 (N86, N82, N69);
nor NOR2 (N87, N75, N27);
and AND4 (N88, N85, N1, N45, N82);
nor NOR3 (N89, N76, N31, N27);
not NOT1 (N90, N61);
buf BUF1 (N91, N83);
nor NOR2 (N92, N90, N49);
or OR3 (N93, N80, N16, N55);
or OR4 (N94, N88, N23, N1, N27);
or OR4 (N95, N86, N48, N52, N53);
and AND4 (N96, N89, N85, N43, N46);
buf BUF1 (N97, N93);
nor NOR3 (N98, N95, N14, N6);
not NOT1 (N99, N97);
xor XOR2 (N100, N77, N95);
nor NOR2 (N101, N96, N62);
nand NAND2 (N102, N100, N89);
buf BUF1 (N103, N81);
nand NAND4 (N104, N101, N50, N2, N31);
xor XOR2 (N105, N87, N52);
nor NOR3 (N106, N102, N85, N42);
buf BUF1 (N107, N106);
xor XOR2 (N108, N99, N13);
xor XOR2 (N109, N104, N24);
not NOT1 (N110, N94);
buf BUF1 (N111, N105);
buf BUF1 (N112, N84);
nand NAND2 (N113, N110, N14);
nand NAND2 (N114, N107, N95);
nand NAND2 (N115, N98, N7);
xor XOR2 (N116, N112, N10);
and AND2 (N117, N103, N22);
not NOT1 (N118, N113);
xor XOR2 (N119, N115, N87);
xor XOR2 (N120, N92, N31);
nand NAND4 (N121, N117, N52, N116, N107);
or OR2 (N122, N107, N66);
nand NAND3 (N123, N118, N87, N114);
nand NAND2 (N124, N116, N17);
not NOT1 (N125, N91);
nand NAND2 (N126, N119, N12);
buf BUF1 (N127, N126);
or OR4 (N128, N111, N25, N11, N112);
nand NAND3 (N129, N124, N93, N21);
nor NOR3 (N130, N122, N72, N112);
nand NAND2 (N131, N120, N13);
xor XOR2 (N132, N131, N118);
buf BUF1 (N133, N125);
nor NOR3 (N134, N129, N34, N56);
xor XOR2 (N135, N130, N82);
not NOT1 (N136, N108);
nand NAND4 (N137, N109, N29, N84, N136);
xor XOR2 (N138, N77, N115);
or OR2 (N139, N128, N28);
not NOT1 (N140, N139);
or OR3 (N141, N127, N48, N88);
not NOT1 (N142, N135);
nor NOR4 (N143, N138, N74, N32, N83);
xor XOR2 (N144, N132, N125);
not NOT1 (N145, N143);
nor NOR2 (N146, N121, N41);
buf BUF1 (N147, N123);
nor NOR3 (N148, N144, N91, N59);
buf BUF1 (N149, N133);
or OR3 (N150, N147, N9, N40);
or OR4 (N151, N134, N1, N3, N20);
or OR4 (N152, N140, N49, N19, N140);
buf BUF1 (N153, N145);
not NOT1 (N154, N148);
nand NAND2 (N155, N141, N68);
xor XOR2 (N156, N153, N106);
and AND3 (N157, N142, N12, N78);
xor XOR2 (N158, N137, N143);
and AND3 (N159, N146, N20, N107);
xor XOR2 (N160, N151, N89);
or OR4 (N161, N156, N85, N121, N111);
not NOT1 (N162, N155);
and AND2 (N163, N159, N98);
or OR3 (N164, N154, N30, N24);
nor NOR2 (N165, N161, N62);
nand NAND2 (N166, N157, N71);
or OR4 (N167, N152, N1, N123, N124);
nor NOR2 (N168, N163, N17);
buf BUF1 (N169, N149);
not NOT1 (N170, N168);
nand NAND2 (N171, N170, N162);
or OR2 (N172, N121, N97);
xor XOR2 (N173, N166, N79);
nand NAND2 (N174, N160, N121);
or OR2 (N175, N172, N141);
xor XOR2 (N176, N173, N43);
not NOT1 (N177, N158);
nor NOR3 (N178, N164, N7, N153);
buf BUF1 (N179, N176);
and AND3 (N180, N165, N89, N151);
nand NAND4 (N181, N169, N6, N47, N84);
or OR4 (N182, N167, N57, N152, N5);
or OR2 (N183, N175, N163);
not NOT1 (N184, N174);
nand NAND3 (N185, N171, N141, N179);
nor NOR3 (N186, N38, N148, N70);
or OR2 (N187, N177, N82);
or OR4 (N188, N187, N121, N147, N112);
not NOT1 (N189, N180);
nor NOR3 (N190, N188, N186, N154);
nand NAND2 (N191, N106, N61);
nand NAND3 (N192, N185, N166, N155);
or OR4 (N193, N191, N21, N68, N24);
nand NAND4 (N194, N189, N12, N48, N170);
nand NAND3 (N195, N193, N35, N163);
or OR4 (N196, N150, N149, N98, N58);
nand NAND4 (N197, N192, N110, N53, N84);
or OR2 (N198, N184, N65);
or OR2 (N199, N195, N121);
not NOT1 (N200, N198);
nand NAND3 (N201, N190, N33, N149);
xor XOR2 (N202, N183, N125);
nor NOR2 (N203, N196, N119);
xor XOR2 (N204, N182, N151);
xor XOR2 (N205, N202, N167);
or OR4 (N206, N197, N168, N95, N172);
nand NAND3 (N207, N200, N59, N189);
not NOT1 (N208, N203);
not NOT1 (N209, N207);
not NOT1 (N210, N208);
buf BUF1 (N211, N209);
buf BUF1 (N212, N206);
and AND3 (N213, N204, N40, N170);
nor NOR2 (N214, N181, N44);
xor XOR2 (N215, N178, N140);
and AND2 (N216, N214, N59);
nor NOR4 (N217, N210, N143, N73, N187);
nand NAND4 (N218, N205, N158, N41, N133);
nand NAND3 (N219, N201, N35, N70);
nand NAND4 (N220, N218, N7, N10, N218);
nor NOR2 (N221, N216, N212);
xor XOR2 (N222, N48, N3);
xor XOR2 (N223, N221, N215);
nand NAND3 (N224, N66, N15, N161);
or OR3 (N225, N217, N50, N140);
xor XOR2 (N226, N199, N25);
or OR4 (N227, N213, N4, N213, N5);
and AND4 (N228, N222, N183, N166, N115);
not NOT1 (N229, N220);
not NOT1 (N230, N228);
xor XOR2 (N231, N223, N188);
not NOT1 (N232, N231);
xor XOR2 (N233, N229, N26);
nand NAND2 (N234, N225, N24);
buf BUF1 (N235, N234);
and AND3 (N236, N211, N163, N196);
nand NAND2 (N237, N235, N176);
nor NOR4 (N238, N230, N125, N77, N168);
and AND4 (N239, N232, N25, N92, N135);
or OR3 (N240, N219, N123, N124);
and AND2 (N241, N240, N194);
nor NOR2 (N242, N88, N141);
nand NAND3 (N243, N242, N137, N59);
nand NAND4 (N244, N241, N70, N194, N66);
or OR4 (N245, N237, N32, N197, N186);
nand NAND3 (N246, N245, N170, N97);
buf BUF1 (N247, N239);
or OR2 (N248, N243, N243);
or OR3 (N249, N246, N47, N236);
buf BUF1 (N250, N19);
xor XOR2 (N251, N227, N181);
nand NAND3 (N252, N233, N29, N28);
buf BUF1 (N253, N250);
not NOT1 (N254, N251);
and AND3 (N255, N238, N220, N59);
or OR3 (N256, N252, N80, N29);
not NOT1 (N257, N247);
or OR3 (N258, N244, N8, N156);
xor XOR2 (N259, N255, N22);
not NOT1 (N260, N224);
and AND3 (N261, N254, N18, N197);
or OR2 (N262, N226, N232);
nand NAND2 (N263, N253, N107);
nand NAND4 (N264, N257, N137, N88, N228);
or OR2 (N265, N264, N253);
and AND2 (N266, N248, N170);
or OR3 (N267, N263, N88, N241);
nand NAND2 (N268, N249, N2);
nor NOR2 (N269, N266, N20);
nor NOR4 (N270, N256, N169, N166, N51);
and AND4 (N271, N261, N112, N200, N265);
and AND4 (N272, N42, N259, N107, N110);
xor XOR2 (N273, N243, N17);
buf BUF1 (N274, N262);
and AND2 (N275, N267, N123);
or OR4 (N276, N271, N164, N195, N68);
buf BUF1 (N277, N275);
not NOT1 (N278, N258);
or OR3 (N279, N260, N257, N132);
xor XOR2 (N280, N272, N229);
not NOT1 (N281, N270);
not NOT1 (N282, N279);
or OR4 (N283, N281, N216, N84, N159);
not NOT1 (N284, N283);
not NOT1 (N285, N268);
xor XOR2 (N286, N278, N9);
not NOT1 (N287, N286);
or OR4 (N288, N277, N272, N232, N10);
xor XOR2 (N289, N287, N178);
nor NOR4 (N290, N289, N167, N27, N3);
buf BUF1 (N291, N290);
nand NAND2 (N292, N282, N288);
buf BUF1 (N293, N69);
or OR2 (N294, N274, N170);
not NOT1 (N295, N276);
not NOT1 (N296, N285);
nand NAND4 (N297, N269, N285, N149, N143);
nand NAND4 (N298, N294, N113, N135, N159);
xor XOR2 (N299, N284, N76);
or OR2 (N300, N295, N37);
nand NAND4 (N301, N299, N227, N46, N36);
xor XOR2 (N302, N296, N270);
nand NAND3 (N303, N301, N13, N100);
nor NOR3 (N304, N280, N260, N250);
buf BUF1 (N305, N300);
and AND4 (N306, N273, N39, N189, N292);
not NOT1 (N307, N133);
and AND2 (N308, N291, N106);
xor XOR2 (N309, N303, N128);
and AND4 (N310, N304, N223, N167, N55);
and AND3 (N311, N297, N130, N116);
and AND2 (N312, N310, N299);
nor NOR3 (N313, N302, N111, N290);
not NOT1 (N314, N313);
xor XOR2 (N315, N308, N174);
not NOT1 (N316, N298);
nor NOR3 (N317, N314, N228, N270);
nand NAND4 (N318, N311, N28, N296, N216);
or OR2 (N319, N293, N263);
nor NOR4 (N320, N306, N161, N302, N86);
and AND2 (N321, N305, N65);
buf BUF1 (N322, N318);
not NOT1 (N323, N315);
buf BUF1 (N324, N316);
buf BUF1 (N325, N324);
buf BUF1 (N326, N323);
nand NAND3 (N327, N317, N179, N47);
or OR4 (N328, N312, N275, N184, N11);
not NOT1 (N329, N328);
or OR2 (N330, N325, N8);
xor XOR2 (N331, N319, N276);
nor NOR4 (N332, N322, N286, N115, N305);
xor XOR2 (N333, N320, N146);
nor NOR3 (N334, N332, N299, N76);
buf BUF1 (N335, N307);
or OR4 (N336, N326, N319, N217, N95);
or OR2 (N337, N330, N206);
or OR2 (N338, N309, N296);
and AND2 (N339, N321, N69);
or OR2 (N340, N336, N44);
or OR3 (N341, N333, N216, N192);
not NOT1 (N342, N329);
nor NOR2 (N343, N331, N233);
and AND3 (N344, N338, N124, N249);
nor NOR3 (N345, N339, N189, N7);
buf BUF1 (N346, N344);
not NOT1 (N347, N334);
and AND2 (N348, N337, N121);
or OR4 (N349, N348, N143, N246, N265);
and AND2 (N350, N349, N173);
buf BUF1 (N351, N340);
xor XOR2 (N352, N347, N11);
not NOT1 (N353, N342);
xor XOR2 (N354, N353, N246);
xor XOR2 (N355, N354, N41);
or OR4 (N356, N341, N23, N258, N234);
xor XOR2 (N357, N346, N322);
xor XOR2 (N358, N345, N134);
buf BUF1 (N359, N343);
nor NOR4 (N360, N350, N288, N57, N85);
not NOT1 (N361, N327);
or OR4 (N362, N352, N248, N41, N255);
nor NOR4 (N363, N357, N95, N157, N159);
and AND3 (N364, N360, N219, N119);
or OR3 (N365, N363, N297, N110);
or OR2 (N366, N365, N223);
or OR3 (N367, N361, N254, N110);
nand NAND4 (N368, N335, N303, N347, N182);
nor NOR2 (N369, N362, N253);
nand NAND2 (N370, N359, N286);
or OR4 (N371, N368, N16, N198, N308);
not NOT1 (N372, N356);
or OR2 (N373, N369, N146);
nand NAND3 (N374, N358, N257, N219);
nand NAND4 (N375, N373, N365, N169, N78);
not NOT1 (N376, N367);
and AND4 (N377, N372, N376, N27, N64);
not NOT1 (N378, N90);
and AND3 (N379, N366, N347, N104);
nand NAND2 (N380, N364, N10);
or OR2 (N381, N377, N111);
and AND3 (N382, N370, N26, N312);
not NOT1 (N383, N379);
nor NOR4 (N384, N374, N72, N294, N301);
xor XOR2 (N385, N355, N285);
xor XOR2 (N386, N383, N179);
buf BUF1 (N387, N384);
xor XOR2 (N388, N382, N133);
and AND4 (N389, N378, N91, N122, N128);
buf BUF1 (N390, N385);
xor XOR2 (N391, N390, N10);
xor XOR2 (N392, N351, N165);
xor XOR2 (N393, N386, N195);
xor XOR2 (N394, N375, N165);
xor XOR2 (N395, N381, N142);
not NOT1 (N396, N393);
buf BUF1 (N397, N388);
xor XOR2 (N398, N392, N65);
and AND2 (N399, N387, N280);
nor NOR2 (N400, N395, N391);
or OR2 (N401, N170, N393);
or OR3 (N402, N397, N307, N45);
nor NOR3 (N403, N401, N377, N59);
xor XOR2 (N404, N402, N258);
or OR4 (N405, N389, N178, N24, N62);
nand NAND2 (N406, N399, N36);
nor NOR4 (N407, N396, N63, N248, N28);
nand NAND4 (N408, N398, N303, N78, N299);
xor XOR2 (N409, N403, N199);
not NOT1 (N410, N404);
nor NOR4 (N411, N405, N260, N365, N165);
xor XOR2 (N412, N406, N345);
or OR3 (N413, N412, N50, N354);
and AND3 (N414, N400, N166, N140);
buf BUF1 (N415, N408);
nand NAND4 (N416, N411, N23, N372, N360);
not NOT1 (N417, N414);
nand NAND2 (N418, N413, N3);
or OR2 (N419, N409, N202);
buf BUF1 (N420, N371);
xor XOR2 (N421, N410, N50);
xor XOR2 (N422, N407, N43);
buf BUF1 (N423, N421);
buf BUF1 (N424, N380);
nand NAND4 (N425, N416, N369, N280, N163);
and AND3 (N426, N425, N72, N91);
nand NAND3 (N427, N423, N321, N202);
buf BUF1 (N428, N420);
not NOT1 (N429, N424);
buf BUF1 (N430, N428);
and AND3 (N431, N418, N419, N40);
not NOT1 (N432, N104);
not NOT1 (N433, N431);
nand NAND3 (N434, N426, N311, N187);
buf BUF1 (N435, N422);
or OR3 (N436, N433, N385, N228);
nand NAND4 (N437, N432, N83, N7, N292);
xor XOR2 (N438, N437, N334);
buf BUF1 (N439, N436);
buf BUF1 (N440, N438);
and AND3 (N441, N430, N220, N188);
and AND2 (N442, N427, N8);
nand NAND3 (N443, N394, N24, N402);
xor XOR2 (N444, N415, N48);
nand NAND4 (N445, N429, N310, N353, N237);
not NOT1 (N446, N444);
nor NOR4 (N447, N442, N254, N248, N146);
xor XOR2 (N448, N417, N90);
and AND4 (N449, N435, N18, N91, N416);
not NOT1 (N450, N440);
nand NAND2 (N451, N446, N183);
xor XOR2 (N452, N447, N102);
and AND3 (N453, N449, N363, N447);
xor XOR2 (N454, N443, N396);
nand NAND4 (N455, N450, N180, N67, N252);
not NOT1 (N456, N455);
xor XOR2 (N457, N434, N46);
or OR4 (N458, N451, N191, N222, N357);
or OR3 (N459, N453, N456, N369);
and AND3 (N460, N23, N218, N81);
not NOT1 (N461, N445);
buf BUF1 (N462, N441);
and AND2 (N463, N454, N125);
xor XOR2 (N464, N452, N321);
buf BUF1 (N465, N457);
and AND4 (N466, N459, N229, N285, N106);
or OR4 (N467, N463, N81, N397, N111);
nand NAND2 (N468, N460, N128);
not NOT1 (N469, N439);
and AND4 (N470, N466, N5, N105, N149);
xor XOR2 (N471, N469, N437);
or OR2 (N472, N471, N184);
not NOT1 (N473, N464);
nor NOR4 (N474, N462, N376, N12, N283);
not NOT1 (N475, N461);
or OR4 (N476, N465, N369, N409, N467);
xor XOR2 (N477, N228, N410);
nand NAND3 (N478, N458, N144, N372);
nor NOR2 (N479, N473, N435);
not NOT1 (N480, N476);
buf BUF1 (N481, N479);
nor NOR3 (N482, N472, N189, N199);
xor XOR2 (N483, N470, N176);
and AND3 (N484, N475, N54, N457);
and AND3 (N485, N474, N445, N444);
nor NOR3 (N486, N468, N257, N224);
or OR2 (N487, N486, N337);
and AND2 (N488, N482, N264);
and AND3 (N489, N480, N95, N232);
nor NOR3 (N490, N448, N340, N65);
nand NAND3 (N491, N488, N347, N279);
buf BUF1 (N492, N489);
not NOT1 (N493, N485);
xor XOR2 (N494, N491, N328);
buf BUF1 (N495, N478);
nor NOR4 (N496, N483, N229, N174, N4);
not NOT1 (N497, N492);
nor NOR4 (N498, N481, N160, N235, N283);
not NOT1 (N499, N497);
buf BUF1 (N500, N484);
buf BUF1 (N501, N494);
nor NOR3 (N502, N498, N424, N30);
not NOT1 (N503, N495);
nor NOR3 (N504, N500, N276, N134);
or OR4 (N505, N504, N476, N227, N150);
buf BUF1 (N506, N496);
nand NAND3 (N507, N505, N457, N352);
not NOT1 (N508, N493);
nor NOR2 (N509, N487, N251);
buf BUF1 (N510, N506);
xor XOR2 (N511, N507, N135);
nor NOR2 (N512, N509, N229);
nor NOR4 (N513, N511, N18, N98, N151);
not NOT1 (N514, N513);
xor XOR2 (N515, N490, N306);
or OR4 (N516, N508, N466, N278, N184);
xor XOR2 (N517, N499, N144);
nor NOR2 (N518, N503, N90);
buf BUF1 (N519, N515);
or OR2 (N520, N514, N49);
nand NAND2 (N521, N519, N5);
not NOT1 (N522, N518);
nor NOR3 (N523, N522, N225, N118);
nand NAND3 (N524, N521, N302, N489);
and AND4 (N525, N502, N504, N42, N377);
not NOT1 (N526, N517);
buf BUF1 (N527, N526);
xor XOR2 (N528, N510, N7);
and AND2 (N529, N528, N130);
nor NOR4 (N530, N523, N474, N223, N442);
not NOT1 (N531, N512);
or OR3 (N532, N531, N471, N300);
buf BUF1 (N533, N516);
nand NAND2 (N534, N530, N22);
nand NAND2 (N535, N533, N480);
not NOT1 (N536, N527);
and AND3 (N537, N535, N86, N498);
not NOT1 (N538, N525);
not NOT1 (N539, N477);
nor NOR2 (N540, N534, N438);
not NOT1 (N541, N520);
xor XOR2 (N542, N532, N357);
not NOT1 (N543, N542);
not NOT1 (N544, N538);
nand NAND2 (N545, N524, N188);
nor NOR3 (N546, N501, N241, N222);
not NOT1 (N547, N529);
nand NAND2 (N548, N543, N458);
xor XOR2 (N549, N546, N382);
or OR3 (N550, N537, N175, N230);
nor NOR3 (N551, N536, N239, N138);
and AND4 (N552, N544, N208, N22, N299);
nor NOR4 (N553, N545, N38, N254, N460);
and AND2 (N554, N548, N414);
xor XOR2 (N555, N553, N386);
nor NOR2 (N556, N541, N536);
xor XOR2 (N557, N539, N523);
nor NOR3 (N558, N555, N3, N315);
nand NAND2 (N559, N549, N343);
buf BUF1 (N560, N540);
xor XOR2 (N561, N560, N254);
xor XOR2 (N562, N557, N349);
nand NAND2 (N563, N554, N66);
and AND3 (N564, N563, N158, N468);
xor XOR2 (N565, N550, N507);
buf BUF1 (N566, N547);
and AND2 (N567, N556, N224);
nand NAND3 (N568, N565, N20, N359);
not NOT1 (N569, N566);
not NOT1 (N570, N552);
buf BUF1 (N571, N559);
or OR3 (N572, N570, N368, N61);
buf BUF1 (N573, N569);
nor NOR3 (N574, N568, N478, N238);
xor XOR2 (N575, N574, N238);
xor XOR2 (N576, N562, N30);
buf BUF1 (N577, N571);
and AND2 (N578, N567, N396);
nor NOR4 (N579, N576, N178, N308, N528);
not NOT1 (N580, N577);
buf BUF1 (N581, N558);
buf BUF1 (N582, N572);
not NOT1 (N583, N581);
nor NOR3 (N584, N573, N485, N244);
or OR2 (N585, N579, N16);
and AND2 (N586, N580, N319);
or OR2 (N587, N582, N399);
buf BUF1 (N588, N561);
nor NOR4 (N589, N551, N521, N158, N436);
xor XOR2 (N590, N589, N365);
and AND4 (N591, N587, N52, N240, N533);
xor XOR2 (N592, N583, N581);
xor XOR2 (N593, N592, N462);
not NOT1 (N594, N585);
nor NOR3 (N595, N593, N496, N371);
xor XOR2 (N596, N588, N517);
not NOT1 (N597, N564);
nand NAND2 (N598, N597, N52);
not NOT1 (N599, N596);
buf BUF1 (N600, N594);
not NOT1 (N601, N586);
and AND3 (N602, N601, N374, N121);
or OR4 (N603, N578, N457, N31, N462);
and AND4 (N604, N599, N468, N315, N541);
xor XOR2 (N605, N604, N151);
nor NOR2 (N606, N595, N164);
and AND2 (N607, N602, N47);
or OR3 (N608, N605, N75, N199);
not NOT1 (N609, N584);
or OR4 (N610, N591, N72, N192, N401);
nand NAND3 (N611, N575, N400, N71);
xor XOR2 (N612, N600, N528);
and AND3 (N613, N608, N105, N183);
not NOT1 (N614, N606);
xor XOR2 (N615, N613, N135);
buf BUF1 (N616, N609);
nor NOR3 (N617, N607, N43, N588);
and AND2 (N618, N590, N31);
not NOT1 (N619, N617);
not NOT1 (N620, N598);
xor XOR2 (N621, N614, N39);
nand NAND3 (N622, N616, N448, N207);
buf BUF1 (N623, N621);
or OR3 (N624, N618, N340, N613);
nand NAND2 (N625, N610, N404);
nand NAND4 (N626, N620, N534, N129, N623);
nor NOR4 (N627, N56, N573, N486, N68);
nand NAND2 (N628, N627, N284);
or OR3 (N629, N619, N1, N225);
and AND2 (N630, N622, N210);
buf BUF1 (N631, N612);
xor XOR2 (N632, N615, N56);
xor XOR2 (N633, N624, N131);
nand NAND3 (N634, N626, N495, N549);
not NOT1 (N635, N625);
buf BUF1 (N636, N628);
and AND3 (N637, N631, N267, N375);
xor XOR2 (N638, N629, N509);
not NOT1 (N639, N603);
nand NAND3 (N640, N630, N475, N59);
nand NAND4 (N641, N633, N552, N99, N158);
xor XOR2 (N642, N640, N83);
buf BUF1 (N643, N611);
not NOT1 (N644, N638);
xor XOR2 (N645, N636, N287);
xor XOR2 (N646, N645, N110);
or OR4 (N647, N646, N548, N610, N44);
nand NAND4 (N648, N639, N600, N166, N536);
xor XOR2 (N649, N648, N335);
not NOT1 (N650, N643);
and AND3 (N651, N637, N641, N40);
and AND3 (N652, N187, N41, N245);
and AND4 (N653, N647, N334, N622, N86);
xor XOR2 (N654, N653, N190);
and AND3 (N655, N654, N567, N263);
or OR3 (N656, N634, N91, N435);
not NOT1 (N657, N652);
nand NAND4 (N658, N650, N99, N499, N224);
nand NAND2 (N659, N656, N348);
nand NAND3 (N660, N655, N494, N327);
or OR4 (N661, N632, N194, N239, N260);
buf BUF1 (N662, N659);
nand NAND3 (N663, N658, N632, N379);
or OR3 (N664, N661, N218, N63);
not NOT1 (N665, N642);
and AND4 (N666, N662, N612, N368, N314);
xor XOR2 (N667, N644, N573);
xor XOR2 (N668, N649, N304);
or OR4 (N669, N663, N421, N48, N634);
buf BUF1 (N670, N668);
buf BUF1 (N671, N670);
nor NOR4 (N672, N664, N493, N281, N528);
and AND4 (N673, N665, N73, N149, N175);
not NOT1 (N674, N671);
or OR3 (N675, N674, N540, N223);
buf BUF1 (N676, N669);
xor XOR2 (N677, N667, N353);
xor XOR2 (N678, N672, N559);
buf BUF1 (N679, N673);
or OR4 (N680, N660, N78, N450, N388);
xor XOR2 (N681, N679, N102);
and AND4 (N682, N651, N628, N330, N429);
buf BUF1 (N683, N677);
nor NOR2 (N684, N675, N592);
or OR4 (N685, N680, N368, N350, N136);
and AND3 (N686, N676, N591, N601);
or OR4 (N687, N684, N137, N51, N222);
nor NOR4 (N688, N678, N112, N405, N329);
or OR2 (N689, N681, N556);
xor XOR2 (N690, N687, N118);
buf BUF1 (N691, N690);
buf BUF1 (N692, N686);
nor NOR2 (N693, N685, N200);
or OR3 (N694, N689, N397, N273);
and AND2 (N695, N694, N243);
not NOT1 (N696, N657);
not NOT1 (N697, N693);
and AND4 (N698, N683, N370, N446, N693);
buf BUF1 (N699, N696);
nor NOR2 (N700, N688, N533);
and AND4 (N701, N691, N589, N614, N43);
and AND2 (N702, N682, N491);
xor XOR2 (N703, N699, N497);
and AND2 (N704, N697, N402);
or OR4 (N705, N702, N663, N457, N2);
nor NOR4 (N706, N701, N344, N278, N424);
nor NOR2 (N707, N706, N18);
nand NAND3 (N708, N695, N604, N424);
xor XOR2 (N709, N698, N229);
nor NOR2 (N710, N692, N623);
nor NOR4 (N711, N707, N21, N469, N314);
nor NOR4 (N712, N711, N630, N607, N64);
and AND2 (N713, N712, N369);
xor XOR2 (N714, N666, N527);
not NOT1 (N715, N713);
buf BUF1 (N716, N710);
nand NAND4 (N717, N715, N516, N640, N450);
and AND4 (N718, N709, N555, N394, N445);
not NOT1 (N719, N703);
and AND4 (N720, N708, N484, N377, N158);
buf BUF1 (N721, N635);
not NOT1 (N722, N716);
xor XOR2 (N723, N705, N116);
and AND4 (N724, N714, N515, N678, N416);
and AND4 (N725, N720, N322, N623, N297);
buf BUF1 (N726, N723);
buf BUF1 (N727, N717);
buf BUF1 (N728, N700);
buf BUF1 (N729, N718);
nand NAND3 (N730, N719, N215, N59);
nand NAND4 (N731, N724, N133, N457, N67);
or OR2 (N732, N729, N4);
or OR4 (N733, N730, N360, N209, N184);
nor NOR3 (N734, N733, N33, N567);
nor NOR2 (N735, N734, N504);
or OR3 (N736, N721, N614, N585);
or OR3 (N737, N728, N594, N576);
nor NOR3 (N738, N731, N289, N626);
not NOT1 (N739, N737);
xor XOR2 (N740, N725, N343);
xor XOR2 (N741, N726, N371);
buf BUF1 (N742, N732);
or OR3 (N743, N742, N329, N206);
nand NAND4 (N744, N743, N625, N262, N140);
nor NOR4 (N745, N744, N31, N321, N1);
nor NOR2 (N746, N740, N526);
nor NOR2 (N747, N727, N583);
not NOT1 (N748, N722);
xor XOR2 (N749, N747, N313);
nor NOR2 (N750, N745, N339);
nor NOR4 (N751, N748, N348, N490, N443);
xor XOR2 (N752, N739, N620);
nand NAND4 (N753, N746, N474, N551, N374);
or OR4 (N754, N749, N321, N54, N513);
nor NOR4 (N755, N735, N665, N83, N457);
or OR3 (N756, N738, N343, N87);
and AND3 (N757, N754, N343, N41);
and AND2 (N758, N736, N472);
buf BUF1 (N759, N758);
not NOT1 (N760, N755);
not NOT1 (N761, N741);
nand NAND4 (N762, N704, N452, N296, N742);
or OR4 (N763, N757, N477, N20, N425);
nand NAND3 (N764, N751, N248, N574);
and AND2 (N765, N759, N481);
buf BUF1 (N766, N763);
and AND4 (N767, N766, N27, N331, N641);
or OR2 (N768, N765, N391);
not NOT1 (N769, N767);
and AND2 (N770, N769, N417);
buf BUF1 (N771, N752);
nand NAND2 (N772, N761, N433);
and AND3 (N773, N764, N396, N338);
or OR4 (N774, N768, N500, N539, N81);
or OR4 (N775, N756, N731, N206, N22);
xor XOR2 (N776, N760, N522);
xor XOR2 (N777, N775, N221);
not NOT1 (N778, N774);
and AND4 (N779, N771, N557, N114, N746);
xor XOR2 (N780, N777, N191);
not NOT1 (N781, N773);
xor XOR2 (N782, N762, N254);
not NOT1 (N783, N770);
and AND3 (N784, N783, N440, N234);
or OR4 (N785, N782, N641, N269, N446);
or OR2 (N786, N781, N640);
nand NAND2 (N787, N785, N438);
xor XOR2 (N788, N778, N420);
xor XOR2 (N789, N780, N537);
nand NAND3 (N790, N786, N771, N125);
nand NAND4 (N791, N779, N20, N586, N309);
nor NOR3 (N792, N776, N8, N686);
xor XOR2 (N793, N790, N540);
buf BUF1 (N794, N793);
and AND2 (N795, N791, N197);
buf BUF1 (N796, N794);
nor NOR4 (N797, N772, N717, N228, N162);
nor NOR2 (N798, N787, N122);
buf BUF1 (N799, N792);
buf BUF1 (N800, N753);
nand NAND2 (N801, N788, N695);
nand NAND4 (N802, N750, N433, N571, N361);
and AND2 (N803, N800, N339);
buf BUF1 (N804, N784);
nor NOR4 (N805, N798, N630, N272, N424);
buf BUF1 (N806, N801);
nand NAND2 (N807, N797, N282);
xor XOR2 (N808, N799, N534);
not NOT1 (N809, N806);
and AND4 (N810, N795, N688, N54, N707);
nor NOR2 (N811, N796, N85);
buf BUF1 (N812, N811);
or OR2 (N813, N803, N811);
buf BUF1 (N814, N804);
not NOT1 (N815, N789);
buf BUF1 (N816, N810);
buf BUF1 (N817, N805);
xor XOR2 (N818, N816, N686);
not NOT1 (N819, N807);
buf BUF1 (N820, N819);
or OR4 (N821, N808, N33, N288, N380);
or OR2 (N822, N809, N640);
nand NAND3 (N823, N820, N517, N526);
or OR2 (N824, N814, N32);
buf BUF1 (N825, N821);
xor XOR2 (N826, N802, N473);
not NOT1 (N827, N824);
and AND2 (N828, N818, N245);
or OR4 (N829, N813, N69, N167, N662);
nor NOR3 (N830, N822, N110, N14);
nor NOR3 (N831, N823, N5, N586);
xor XOR2 (N832, N828, N479);
nand NAND4 (N833, N832, N423, N83, N442);
nor NOR4 (N834, N827, N597, N704, N192);
or OR3 (N835, N833, N501, N260);
buf BUF1 (N836, N829);
xor XOR2 (N837, N830, N68);
nor NOR2 (N838, N837, N537);
xor XOR2 (N839, N815, N559);
nand NAND4 (N840, N826, N688, N494, N299);
not NOT1 (N841, N838);
nand NAND2 (N842, N839, N606);
nand NAND3 (N843, N835, N274, N801);
not NOT1 (N844, N825);
nor NOR2 (N845, N841, N613);
nand NAND4 (N846, N844, N201, N747, N256);
nand NAND2 (N847, N812, N191);
or OR4 (N848, N836, N544, N801, N499);
nor NOR2 (N849, N845, N133);
and AND4 (N850, N843, N84, N54, N171);
xor XOR2 (N851, N846, N762);
xor XOR2 (N852, N842, N794);
not NOT1 (N853, N847);
xor XOR2 (N854, N831, N777);
and AND2 (N855, N840, N30);
or OR3 (N856, N849, N272, N358);
and AND2 (N857, N817, N555);
or OR3 (N858, N854, N73, N221);
nor NOR3 (N859, N850, N335, N126);
buf BUF1 (N860, N834);
nand NAND2 (N861, N855, N292);
or OR2 (N862, N858, N803);
xor XOR2 (N863, N861, N285);
nand NAND4 (N864, N852, N227, N457, N341);
or OR2 (N865, N857, N703);
or OR3 (N866, N865, N576, N52);
nor NOR3 (N867, N866, N16, N356);
xor XOR2 (N868, N859, N6);
buf BUF1 (N869, N867);
not NOT1 (N870, N862);
xor XOR2 (N871, N863, N479);
nor NOR4 (N872, N856, N261, N254, N865);
buf BUF1 (N873, N871);
and AND3 (N874, N870, N276, N235);
and AND3 (N875, N851, N688, N308);
nand NAND4 (N876, N860, N63, N363, N710);
or OR3 (N877, N872, N142, N612);
or OR3 (N878, N864, N871, N128);
not NOT1 (N879, N873);
nand NAND3 (N880, N874, N699, N860);
xor XOR2 (N881, N878, N226);
nor NOR4 (N882, N848, N77, N252, N731);
buf BUF1 (N883, N868);
not NOT1 (N884, N853);
xor XOR2 (N885, N879, N12);
not NOT1 (N886, N877);
buf BUF1 (N887, N880);
buf BUF1 (N888, N883);
not NOT1 (N889, N884);
nand NAND4 (N890, N869, N430, N810, N652);
nand NAND4 (N891, N886, N392, N115, N766);
or OR2 (N892, N889, N196);
nor NOR4 (N893, N892, N634, N109, N814);
and AND3 (N894, N881, N874, N854);
not NOT1 (N895, N882);
nor NOR4 (N896, N891, N590, N185, N115);
and AND3 (N897, N896, N333, N887);
not NOT1 (N898, N506);
xor XOR2 (N899, N898, N120);
or OR2 (N900, N895, N884);
and AND4 (N901, N894, N522, N330, N665);
xor XOR2 (N902, N888, N142);
xor XOR2 (N903, N897, N346);
xor XOR2 (N904, N885, N351);
nor NOR3 (N905, N899, N713, N588);
not NOT1 (N906, N904);
nand NAND2 (N907, N900, N508);
not NOT1 (N908, N876);
xor XOR2 (N909, N893, N360);
nand NAND4 (N910, N903, N276, N427, N188);
or OR4 (N911, N875, N603, N785, N441);
or OR2 (N912, N908, N883);
buf BUF1 (N913, N912);
not NOT1 (N914, N911);
or OR3 (N915, N905, N569, N417);
buf BUF1 (N916, N909);
nand NAND3 (N917, N910, N537, N290);
and AND2 (N918, N902, N392);
not NOT1 (N919, N906);
and AND4 (N920, N913, N634, N220, N871);
xor XOR2 (N921, N920, N311);
nand NAND4 (N922, N901, N291, N396, N437);
nor NOR2 (N923, N921, N63);
xor XOR2 (N924, N914, N582);
buf BUF1 (N925, N916);
nand NAND2 (N926, N915, N458);
and AND2 (N927, N919, N153);
nor NOR2 (N928, N890, N383);
nor NOR2 (N929, N924, N246);
or OR4 (N930, N928, N879, N64, N868);
nor NOR4 (N931, N929, N278, N851, N268);
nor NOR2 (N932, N927, N874);
not NOT1 (N933, N922);
or OR2 (N934, N933, N766);
nand NAND2 (N935, N907, N106);
not NOT1 (N936, N934);
buf BUF1 (N937, N931);
buf BUF1 (N938, N932);
buf BUF1 (N939, N930);
or OR2 (N940, N935, N758);
and AND4 (N941, N923, N360, N865, N101);
xor XOR2 (N942, N917, N377);
buf BUF1 (N943, N941);
and AND2 (N944, N936, N73);
or OR4 (N945, N937, N770, N816, N91);
nand NAND4 (N946, N945, N546, N220, N677);
and AND3 (N947, N942, N408, N76);
xor XOR2 (N948, N944, N817);
xor XOR2 (N949, N918, N231);
nand NAND4 (N950, N925, N100, N312, N261);
xor XOR2 (N951, N949, N670);
or OR4 (N952, N951, N510, N710, N464);
and AND3 (N953, N950, N708, N838);
or OR3 (N954, N943, N96, N65);
buf BUF1 (N955, N952);
nor NOR3 (N956, N947, N899, N596);
and AND3 (N957, N954, N882, N70);
and AND3 (N958, N939, N729, N833);
and AND3 (N959, N956, N88, N8);
and AND2 (N960, N948, N601);
or OR2 (N961, N957, N916);
nor NOR2 (N962, N959, N280);
or OR3 (N963, N961, N896, N548);
buf BUF1 (N964, N963);
nor NOR2 (N965, N964, N21);
buf BUF1 (N966, N926);
nand NAND4 (N967, N955, N963, N785, N833);
or OR3 (N968, N940, N835, N123);
nand NAND4 (N969, N968, N964, N637, N540);
nor NOR2 (N970, N958, N309);
and AND2 (N971, N953, N73);
xor XOR2 (N972, N970, N860);
nor NOR2 (N973, N971, N338);
and AND2 (N974, N966, N141);
or OR3 (N975, N946, N189, N154);
and AND3 (N976, N969, N860, N510);
or OR4 (N977, N973, N136, N63, N234);
not NOT1 (N978, N960);
not NOT1 (N979, N977);
nor NOR3 (N980, N979, N24, N580);
nand NAND3 (N981, N976, N806, N490);
xor XOR2 (N982, N962, N789);
or OR4 (N983, N981, N127, N473, N546);
buf BUF1 (N984, N982);
nor NOR3 (N985, N967, N751, N763);
or OR4 (N986, N984, N654, N398, N493);
xor XOR2 (N987, N983, N545);
or OR4 (N988, N965, N368, N6, N869);
not NOT1 (N989, N978);
not NOT1 (N990, N972);
or OR2 (N991, N938, N730);
not NOT1 (N992, N987);
nand NAND3 (N993, N992, N935, N276);
or OR2 (N994, N974, N557);
buf BUF1 (N995, N994);
or OR3 (N996, N990, N666, N55);
and AND3 (N997, N986, N158, N845);
buf BUF1 (N998, N988);
and AND4 (N999, N991, N593, N510, N878);
nor NOR3 (N1000, N993, N628, N5);
not NOT1 (N1001, N997);
and AND2 (N1002, N980, N433);
nor NOR4 (N1003, N998, N906, N169, N686);
xor XOR2 (N1004, N1003, N647);
or OR4 (N1005, N1004, N80, N454, N407);
nor NOR4 (N1006, N1002, N954, N841, N653);
and AND4 (N1007, N999, N162, N341, N895);
nor NOR2 (N1008, N975, N286);
not NOT1 (N1009, N1005);
nand NAND2 (N1010, N989, N260);
xor XOR2 (N1011, N1008, N954);
nand NAND2 (N1012, N1001, N157);
not NOT1 (N1013, N1011);
not NOT1 (N1014, N1010);
xor XOR2 (N1015, N1012, N950);
or OR4 (N1016, N1000, N886, N541, N396);
or OR2 (N1017, N1013, N82);
buf BUF1 (N1018, N985);
nand NAND4 (N1019, N1015, N889, N231, N444);
not NOT1 (N1020, N1014);
not NOT1 (N1021, N996);
and AND4 (N1022, N1019, N203, N689, N291);
nand NAND2 (N1023, N1017, N902);
not NOT1 (N1024, N1009);
or OR4 (N1025, N1007, N275, N587, N373);
xor XOR2 (N1026, N1020, N248);
nor NOR3 (N1027, N1026, N525, N752);
xor XOR2 (N1028, N1024, N306);
not NOT1 (N1029, N995);
buf BUF1 (N1030, N1029);
buf BUF1 (N1031, N1016);
and AND2 (N1032, N1025, N787);
xor XOR2 (N1033, N1027, N706);
or OR4 (N1034, N1028, N596, N852, N276);
nor NOR3 (N1035, N1030, N186, N791);
nor NOR3 (N1036, N1018, N26, N709);
and AND2 (N1037, N1034, N933);
not NOT1 (N1038, N1022);
or OR2 (N1039, N1021, N160);
xor XOR2 (N1040, N1033, N539);
nor NOR3 (N1041, N1035, N309, N682);
and AND2 (N1042, N1006, N796);
nor NOR4 (N1043, N1036, N534, N767, N783);
not NOT1 (N1044, N1041);
xor XOR2 (N1045, N1031, N864);
nand NAND2 (N1046, N1044, N770);
not NOT1 (N1047, N1046);
and AND2 (N1048, N1040, N156);
buf BUF1 (N1049, N1045);
xor XOR2 (N1050, N1043, N1020);
not NOT1 (N1051, N1049);
nor NOR2 (N1052, N1042, N641);
and AND3 (N1053, N1048, N222, N753);
not NOT1 (N1054, N1047);
xor XOR2 (N1055, N1023, N296);
or OR3 (N1056, N1037, N367, N99);
and AND3 (N1057, N1053, N565, N285);
not NOT1 (N1058, N1039);
buf BUF1 (N1059, N1056);
buf BUF1 (N1060, N1051);
or OR3 (N1061, N1055, N423, N83);
buf BUF1 (N1062, N1054);
nor NOR3 (N1063, N1059, N116, N901);
nand NAND4 (N1064, N1038, N76, N22, N384);
or OR4 (N1065, N1062, N808, N209, N162);
and AND4 (N1066, N1057, N925, N36, N679);
buf BUF1 (N1067, N1050);
nor NOR4 (N1068, N1061, N859, N112, N881);
nor NOR3 (N1069, N1065, N928, N633);
not NOT1 (N1070, N1064);
xor XOR2 (N1071, N1058, N415);
xor XOR2 (N1072, N1069, N858);
xor XOR2 (N1073, N1052, N658);
buf BUF1 (N1074, N1063);
nor NOR4 (N1075, N1070, N150, N327, N488);
nor NOR3 (N1076, N1074, N659, N173);
and AND4 (N1077, N1032, N498, N747, N840);
buf BUF1 (N1078, N1068);
nor NOR4 (N1079, N1066, N1046, N57, N842);
xor XOR2 (N1080, N1075, N1009);
buf BUF1 (N1081, N1080);
or OR3 (N1082, N1071, N1029, N432);
not NOT1 (N1083, N1081);
nor NOR3 (N1084, N1082, N207, N265);
buf BUF1 (N1085, N1073);
not NOT1 (N1086, N1079);
or OR2 (N1087, N1076, N357);
or OR3 (N1088, N1087, N814, N1020);
nor NOR2 (N1089, N1072, N956);
or OR3 (N1090, N1060, N365, N752);
nor NOR2 (N1091, N1083, N359);
nor NOR2 (N1092, N1086, N1013);
buf BUF1 (N1093, N1077);
nand NAND4 (N1094, N1078, N979, N95, N998);
or OR3 (N1095, N1089, N686, N357);
nor NOR3 (N1096, N1084, N505, N141);
not NOT1 (N1097, N1067);
not NOT1 (N1098, N1093);
buf BUF1 (N1099, N1085);
not NOT1 (N1100, N1095);
nand NAND3 (N1101, N1099, N725, N934);
not NOT1 (N1102, N1091);
or OR3 (N1103, N1090, N733, N33);
or OR3 (N1104, N1101, N414, N202);
not NOT1 (N1105, N1097);
and AND2 (N1106, N1094, N698);
nand NAND2 (N1107, N1096, N302);
buf BUF1 (N1108, N1105);
not NOT1 (N1109, N1102);
or OR4 (N1110, N1100, N46, N315, N869);
and AND2 (N1111, N1109, N576);
nor NOR2 (N1112, N1111, N180);
or OR3 (N1113, N1107, N637, N112);
nor NOR3 (N1114, N1112, N224, N45);
not NOT1 (N1115, N1108);
or OR3 (N1116, N1106, N170, N437);
nand NAND2 (N1117, N1104, N156);
nor NOR4 (N1118, N1092, N723, N351, N234);
nor NOR4 (N1119, N1117, N585, N866, N1073);
buf BUF1 (N1120, N1115);
nand NAND4 (N1121, N1098, N160, N211, N627);
nor NOR3 (N1122, N1110, N674, N253);
nor NOR3 (N1123, N1113, N582, N804);
not NOT1 (N1124, N1121);
nand NAND3 (N1125, N1119, N994, N571);
nand NAND3 (N1126, N1116, N559, N654);
and AND3 (N1127, N1088, N609, N1064);
nor NOR2 (N1128, N1123, N615);
buf BUF1 (N1129, N1126);
not NOT1 (N1130, N1120);
not NOT1 (N1131, N1129);
xor XOR2 (N1132, N1122, N1054);
not NOT1 (N1133, N1118);
not NOT1 (N1134, N1114);
not NOT1 (N1135, N1124);
nor NOR2 (N1136, N1135, N1073);
buf BUF1 (N1137, N1134);
buf BUF1 (N1138, N1130);
nand NAND4 (N1139, N1132, N663, N110, N120);
and AND3 (N1140, N1131, N225, N203);
and AND4 (N1141, N1136, N1095, N842, N908);
nand NAND4 (N1142, N1133, N286, N736, N138);
xor XOR2 (N1143, N1141, N670);
or OR3 (N1144, N1143, N581, N297);
or OR4 (N1145, N1103, N684, N723, N949);
nand NAND2 (N1146, N1144, N180);
buf BUF1 (N1147, N1146);
not NOT1 (N1148, N1137);
nor NOR3 (N1149, N1147, N864, N160);
buf BUF1 (N1150, N1140);
not NOT1 (N1151, N1148);
not NOT1 (N1152, N1151);
not NOT1 (N1153, N1149);
and AND3 (N1154, N1127, N645, N526);
or OR2 (N1155, N1154, N230);
and AND2 (N1156, N1153, N38);
nor NOR4 (N1157, N1156, N8, N916, N1074);
not NOT1 (N1158, N1138);
and AND2 (N1159, N1128, N359);
nand NAND2 (N1160, N1152, N794);
nand NAND2 (N1161, N1157, N1052);
nor NOR3 (N1162, N1139, N994, N85);
xor XOR2 (N1163, N1145, N1106);
not NOT1 (N1164, N1159);
nor NOR3 (N1165, N1162, N1025, N414);
or OR3 (N1166, N1158, N45, N918);
or OR2 (N1167, N1125, N235);
buf BUF1 (N1168, N1166);
buf BUF1 (N1169, N1150);
nor NOR4 (N1170, N1165, N978, N132, N1041);
and AND3 (N1171, N1161, N967, N1155);
nor NOR2 (N1172, N569, N984);
xor XOR2 (N1173, N1160, N377);
not NOT1 (N1174, N1170);
and AND4 (N1175, N1167, N157, N205, N267);
not NOT1 (N1176, N1171);
not NOT1 (N1177, N1172);
xor XOR2 (N1178, N1168, N847);
nand NAND2 (N1179, N1163, N855);
or OR3 (N1180, N1174, N64, N630);
nor NOR4 (N1181, N1173, N757, N1128, N41);
xor XOR2 (N1182, N1181, N1022);
buf BUF1 (N1183, N1169);
buf BUF1 (N1184, N1175);
nand NAND4 (N1185, N1176, N88, N586, N362);
nand NAND3 (N1186, N1179, N805, N739);
not NOT1 (N1187, N1183);
and AND3 (N1188, N1186, N750, N1146);
nand NAND2 (N1189, N1185, N658);
or OR2 (N1190, N1182, N395);
not NOT1 (N1191, N1190);
not NOT1 (N1192, N1188);
not NOT1 (N1193, N1142);
not NOT1 (N1194, N1193);
nand NAND3 (N1195, N1187, N104, N1151);
or OR4 (N1196, N1164, N1139, N1052, N763);
and AND2 (N1197, N1192, N835);
nor NOR4 (N1198, N1197, N768, N203, N805);
and AND2 (N1199, N1180, N888);
or OR2 (N1200, N1196, N929);
xor XOR2 (N1201, N1184, N798);
nand NAND3 (N1202, N1178, N878, N1100);
xor XOR2 (N1203, N1198, N126);
buf BUF1 (N1204, N1203);
nand NAND4 (N1205, N1200, N839, N975, N485);
or OR3 (N1206, N1177, N656, N968);
not NOT1 (N1207, N1202);
buf BUF1 (N1208, N1194);
not NOT1 (N1209, N1191);
and AND2 (N1210, N1199, N993);
or OR4 (N1211, N1195, N1119, N1116, N473);
buf BUF1 (N1212, N1210);
nor NOR4 (N1213, N1208, N1062, N432, N627);
xor XOR2 (N1214, N1189, N69);
and AND2 (N1215, N1201, N113);
nand NAND2 (N1216, N1207, N219);
nor NOR2 (N1217, N1213, N833);
xor XOR2 (N1218, N1206, N772);
or OR2 (N1219, N1216, N513);
and AND4 (N1220, N1214, N642, N419, N527);
or OR3 (N1221, N1211, N958, N55);
and AND3 (N1222, N1204, N122, N920);
nand NAND2 (N1223, N1222, N530);
not NOT1 (N1224, N1221);
or OR2 (N1225, N1219, N428);
xor XOR2 (N1226, N1215, N112);
or OR4 (N1227, N1220, N842, N715, N302);
or OR3 (N1228, N1205, N96, N215);
nand NAND2 (N1229, N1209, N721);
nor NOR4 (N1230, N1212, N357, N759, N516);
buf BUF1 (N1231, N1228);
nor NOR4 (N1232, N1227, N92, N888, N1044);
and AND3 (N1233, N1229, N773, N392);
xor XOR2 (N1234, N1226, N598);
nand NAND3 (N1235, N1234, N459, N867);
nand NAND4 (N1236, N1218, N347, N889, N1175);
and AND4 (N1237, N1217, N963, N960, N831);
nand NAND2 (N1238, N1223, N36);
xor XOR2 (N1239, N1230, N145);
and AND4 (N1240, N1232, N365, N528, N682);
nor NOR4 (N1241, N1236, N755, N728, N554);
and AND2 (N1242, N1224, N1101);
xor XOR2 (N1243, N1242, N499);
and AND4 (N1244, N1240, N383, N1161, N912);
not NOT1 (N1245, N1231);
nor NOR2 (N1246, N1244, N440);
or OR3 (N1247, N1237, N710, N790);
buf BUF1 (N1248, N1243);
and AND3 (N1249, N1235, N160, N131);
nand NAND4 (N1250, N1239, N599, N1207, N558);
not NOT1 (N1251, N1241);
not NOT1 (N1252, N1251);
and AND2 (N1253, N1233, N637);
nor NOR4 (N1254, N1225, N410, N1159, N1166);
buf BUF1 (N1255, N1247);
not NOT1 (N1256, N1245);
xor XOR2 (N1257, N1246, N706);
or OR4 (N1258, N1250, N1172, N582, N576);
nor NOR3 (N1259, N1238, N711, N575);
nand NAND4 (N1260, N1252, N1171, N1113, N1166);
or OR4 (N1261, N1255, N430, N888, N345);
or OR4 (N1262, N1258, N897, N606, N277);
buf BUF1 (N1263, N1248);
buf BUF1 (N1264, N1259);
or OR2 (N1265, N1264, N812);
or OR4 (N1266, N1262, N378, N353, N1157);
nand NAND2 (N1267, N1249, N601);
nand NAND3 (N1268, N1257, N621, N947);
not NOT1 (N1269, N1265);
or OR2 (N1270, N1266, N61);
or OR4 (N1271, N1256, N426, N580, N272);
buf BUF1 (N1272, N1263);
nand NAND3 (N1273, N1270, N777, N1167);
nand NAND3 (N1274, N1267, N23, N1094);
xor XOR2 (N1275, N1254, N945);
nand NAND4 (N1276, N1261, N770, N807, N1046);
not NOT1 (N1277, N1275);
not NOT1 (N1278, N1277);
xor XOR2 (N1279, N1278, N1146);
not NOT1 (N1280, N1271);
nor NOR2 (N1281, N1272, N763);
and AND3 (N1282, N1260, N282, N810);
buf BUF1 (N1283, N1276);
nor NOR2 (N1284, N1279, N382);
nand NAND2 (N1285, N1284, N1122);
xor XOR2 (N1286, N1274, N93);
not NOT1 (N1287, N1268);
not NOT1 (N1288, N1283);
xor XOR2 (N1289, N1281, N936);
nor NOR2 (N1290, N1286, N1235);
nor NOR2 (N1291, N1269, N149);
xor XOR2 (N1292, N1291, N771);
nand NAND4 (N1293, N1288, N995, N718, N999);
xor XOR2 (N1294, N1285, N16);
buf BUF1 (N1295, N1253);
or OR4 (N1296, N1295, N370, N961, N146);
or OR3 (N1297, N1292, N978, N788);
xor XOR2 (N1298, N1294, N1);
not NOT1 (N1299, N1293);
nand NAND4 (N1300, N1289, N919, N325, N444);
buf BUF1 (N1301, N1300);
xor XOR2 (N1302, N1301, N378);
buf BUF1 (N1303, N1282);
nor NOR3 (N1304, N1280, N35, N600);
xor XOR2 (N1305, N1302, N1234);
not NOT1 (N1306, N1298);
not NOT1 (N1307, N1273);
xor XOR2 (N1308, N1287, N52);
not NOT1 (N1309, N1303);
buf BUF1 (N1310, N1290);
not NOT1 (N1311, N1308);
nand NAND3 (N1312, N1304, N622, N972);
buf BUF1 (N1313, N1311);
nor NOR4 (N1314, N1307, N1181, N253, N1239);
nor NOR2 (N1315, N1313, N731);
nor NOR3 (N1316, N1314, N966, N351);
buf BUF1 (N1317, N1305);
buf BUF1 (N1318, N1312);
xor XOR2 (N1319, N1309, N1117);
and AND3 (N1320, N1319, N680, N687);
not NOT1 (N1321, N1306);
nand NAND2 (N1322, N1315, N1319);
nand NAND3 (N1323, N1318, N937, N46);
buf BUF1 (N1324, N1323);
and AND3 (N1325, N1296, N319, N312);
or OR4 (N1326, N1324, N721, N293, N777);
not NOT1 (N1327, N1326);
or OR2 (N1328, N1316, N1091);
buf BUF1 (N1329, N1320);
not NOT1 (N1330, N1322);
and AND2 (N1331, N1327, N217);
nor NOR2 (N1332, N1331, N271);
or OR2 (N1333, N1332, N1037);
nor NOR3 (N1334, N1310, N1282, N820);
xor XOR2 (N1335, N1321, N336);
nand NAND4 (N1336, N1317, N1012, N1167, N806);
xor XOR2 (N1337, N1328, N923);
xor XOR2 (N1338, N1329, N10);
buf BUF1 (N1339, N1299);
nand NAND3 (N1340, N1325, N1106, N573);
not NOT1 (N1341, N1333);
nand NAND4 (N1342, N1341, N743, N691, N328);
xor XOR2 (N1343, N1338, N20);
nor NOR2 (N1344, N1335, N461);
or OR2 (N1345, N1344, N80);
nand NAND4 (N1346, N1336, N407, N128, N564);
xor XOR2 (N1347, N1339, N1255);
and AND4 (N1348, N1330, N32, N1264, N90);
nand NAND2 (N1349, N1297, N1267);
nand NAND4 (N1350, N1343, N654, N1001, N1112);
not NOT1 (N1351, N1347);
not NOT1 (N1352, N1346);
and AND4 (N1353, N1334, N543, N787, N1034);
nor NOR2 (N1354, N1348, N942);
not NOT1 (N1355, N1353);
or OR3 (N1356, N1355, N1129, N910);
and AND2 (N1357, N1349, N1306);
or OR3 (N1358, N1340, N1356, N22);
xor XOR2 (N1359, N1277, N1076);
or OR4 (N1360, N1351, N353, N216, N762);
xor XOR2 (N1361, N1360, N744);
xor XOR2 (N1362, N1352, N857);
not NOT1 (N1363, N1337);
buf BUF1 (N1364, N1342);
and AND2 (N1365, N1361, N696);
not NOT1 (N1366, N1365);
xor XOR2 (N1367, N1357, N944);
xor XOR2 (N1368, N1345, N906);
xor XOR2 (N1369, N1368, N671);
xor XOR2 (N1370, N1367, N512);
buf BUF1 (N1371, N1354);
buf BUF1 (N1372, N1370);
nand NAND2 (N1373, N1363, N1230);
or OR3 (N1374, N1358, N277, N168);
buf BUF1 (N1375, N1359);
nor NOR4 (N1376, N1375, N1333, N1130, N1205);
not NOT1 (N1377, N1374);
nand NAND3 (N1378, N1371, N558, N1283);
buf BUF1 (N1379, N1377);
and AND3 (N1380, N1364, N1205, N512);
buf BUF1 (N1381, N1372);
nand NAND2 (N1382, N1381, N1170);
not NOT1 (N1383, N1379);
and AND3 (N1384, N1378, N943, N1181);
not NOT1 (N1385, N1366);
and AND2 (N1386, N1385, N704);
xor XOR2 (N1387, N1350, N1323);
or OR4 (N1388, N1386, N1153, N354, N855);
or OR3 (N1389, N1383, N1043, N866);
nor NOR4 (N1390, N1369, N1374, N841, N671);
nand NAND2 (N1391, N1388, N1354);
nor NOR3 (N1392, N1376, N1214, N422);
nor NOR3 (N1393, N1373, N1341, N1263);
nor NOR3 (N1394, N1387, N719, N1373);
xor XOR2 (N1395, N1390, N1251);
or OR2 (N1396, N1384, N893);
nor NOR3 (N1397, N1396, N897, N1233);
or OR2 (N1398, N1393, N465);
xor XOR2 (N1399, N1389, N1079);
nand NAND4 (N1400, N1395, N999, N557, N1092);
or OR3 (N1401, N1391, N621, N143);
nor NOR4 (N1402, N1392, N110, N756, N732);
nor NOR3 (N1403, N1362, N988, N24);
buf BUF1 (N1404, N1394);
nand NAND3 (N1405, N1400, N1334, N804);
nand NAND2 (N1406, N1404, N1261);
nor NOR4 (N1407, N1406, N841, N1252, N630);
and AND4 (N1408, N1402, N391, N619, N601);
buf BUF1 (N1409, N1382);
not NOT1 (N1410, N1407);
buf BUF1 (N1411, N1401);
nand NAND3 (N1412, N1408, N763, N397);
or OR3 (N1413, N1405, N526, N350);
xor XOR2 (N1414, N1413, N1162);
nor NOR4 (N1415, N1414, N279, N745, N678);
or OR2 (N1416, N1403, N1248);
and AND2 (N1417, N1415, N602);
buf BUF1 (N1418, N1380);
nor NOR2 (N1419, N1411, N936);
nor NOR3 (N1420, N1409, N7, N398);
not NOT1 (N1421, N1398);
and AND4 (N1422, N1420, N628, N235, N625);
buf BUF1 (N1423, N1412);
not NOT1 (N1424, N1397);
and AND3 (N1425, N1417, N516, N995);
not NOT1 (N1426, N1422);
not NOT1 (N1427, N1425);
nor NOR4 (N1428, N1399, N609, N85, N410);
not NOT1 (N1429, N1427);
or OR4 (N1430, N1418, N1229, N672, N264);
not NOT1 (N1431, N1426);
buf BUF1 (N1432, N1428);
nand NAND4 (N1433, N1431, N685, N641, N545);
buf BUF1 (N1434, N1410);
nor NOR3 (N1435, N1432, N1303, N490);
or OR3 (N1436, N1429, N940, N415);
and AND4 (N1437, N1433, N352, N854, N1294);
nor NOR3 (N1438, N1430, N760, N382);
nor NOR3 (N1439, N1423, N1433, N840);
nor NOR3 (N1440, N1435, N88, N557);
nor NOR3 (N1441, N1421, N334, N329);
or OR4 (N1442, N1424, N107, N954, N583);
and AND4 (N1443, N1434, N266, N1013, N531);
or OR4 (N1444, N1440, N1443, N157, N422);
not NOT1 (N1445, N897);
xor XOR2 (N1446, N1437, N952);
and AND3 (N1447, N1436, N1309, N204);
nor NOR3 (N1448, N1441, N652, N973);
nand NAND4 (N1449, N1444, N534, N1151, N1321);
or OR2 (N1450, N1447, N1165);
buf BUF1 (N1451, N1448);
not NOT1 (N1452, N1446);
not NOT1 (N1453, N1419);
nand NAND2 (N1454, N1450, N1006);
not NOT1 (N1455, N1451);
buf BUF1 (N1456, N1454);
nor NOR3 (N1457, N1445, N189, N955);
or OR2 (N1458, N1453, N885);
nand NAND4 (N1459, N1449, N892, N386, N161);
nor NOR3 (N1460, N1455, N1305, N201);
or OR2 (N1461, N1458, N333);
nand NAND4 (N1462, N1456, N942, N29, N1042);
and AND3 (N1463, N1452, N966, N584);
or OR3 (N1464, N1459, N718, N695);
buf BUF1 (N1465, N1442);
nor NOR3 (N1466, N1464, N205, N471);
nor NOR3 (N1467, N1457, N921, N1385);
or OR4 (N1468, N1463, N139, N877, N1241);
xor XOR2 (N1469, N1468, N828);
buf BUF1 (N1470, N1439);
not NOT1 (N1471, N1438);
not NOT1 (N1472, N1462);
nand NAND2 (N1473, N1466, N359);
nand NAND3 (N1474, N1469, N36, N1077);
nand NAND3 (N1475, N1460, N1404, N1117);
xor XOR2 (N1476, N1467, N373);
and AND2 (N1477, N1474, N377);
buf BUF1 (N1478, N1471);
or OR2 (N1479, N1476, N842);
or OR4 (N1480, N1473, N842, N128, N139);
and AND4 (N1481, N1475, N1310, N1054, N175);
nand NAND4 (N1482, N1465, N775, N1444, N252);
nor NOR4 (N1483, N1416, N662, N1350, N563);
or OR4 (N1484, N1470, N1455, N1187, N283);
not NOT1 (N1485, N1478);
nand NAND4 (N1486, N1480, N253, N1041, N1094);
nor NOR4 (N1487, N1477, N991, N159, N1208);
nand NAND3 (N1488, N1487, N1474, N597);
and AND3 (N1489, N1461, N1222, N1243);
not NOT1 (N1490, N1486);
and AND3 (N1491, N1483, N1095, N865);
buf BUF1 (N1492, N1484);
and AND2 (N1493, N1472, N1413);
or OR2 (N1494, N1491, N544);
not NOT1 (N1495, N1489);
xor XOR2 (N1496, N1482, N335);
buf BUF1 (N1497, N1496);
buf BUF1 (N1498, N1481);
xor XOR2 (N1499, N1497, N566);
buf BUF1 (N1500, N1492);
and AND4 (N1501, N1498, N735, N939, N237);
not NOT1 (N1502, N1479);
not NOT1 (N1503, N1494);
or OR4 (N1504, N1503, N921, N40, N289);
and AND4 (N1505, N1499, N374, N1267, N112);
and AND3 (N1506, N1504, N553, N236);
not NOT1 (N1507, N1485);
and AND2 (N1508, N1502, N413);
nand NAND2 (N1509, N1488, N1478);
buf BUF1 (N1510, N1495);
buf BUF1 (N1511, N1505);
buf BUF1 (N1512, N1501);
not NOT1 (N1513, N1507);
xor XOR2 (N1514, N1510, N1193);
nand NAND4 (N1515, N1513, N544, N209, N1254);
xor XOR2 (N1516, N1514, N1352);
xor XOR2 (N1517, N1493, N245);
not NOT1 (N1518, N1516);
xor XOR2 (N1519, N1511, N1390);
xor XOR2 (N1520, N1490, N637);
xor XOR2 (N1521, N1509, N24);
or OR4 (N1522, N1515, N388, N1371, N34);
xor XOR2 (N1523, N1512, N774);
buf BUF1 (N1524, N1506);
nand NAND2 (N1525, N1520, N30);
and AND3 (N1526, N1517, N645, N997);
nand NAND4 (N1527, N1522, N605, N933, N102);
buf BUF1 (N1528, N1508);
and AND2 (N1529, N1519, N107);
xor XOR2 (N1530, N1525, N200);
buf BUF1 (N1531, N1524);
nor NOR3 (N1532, N1518, N569, N945);
or OR2 (N1533, N1526, N896);
nor NOR2 (N1534, N1532, N413);
not NOT1 (N1535, N1523);
nor NOR4 (N1536, N1534, N367, N130, N954);
nand NAND4 (N1537, N1529, N742, N1531, N197);
buf BUF1 (N1538, N425);
buf BUF1 (N1539, N1530);
and AND3 (N1540, N1538, N1073, N1131);
or OR4 (N1541, N1539, N478, N1155, N1168);
buf BUF1 (N1542, N1500);
and AND3 (N1543, N1527, N513, N2);
buf BUF1 (N1544, N1540);
nand NAND4 (N1545, N1537, N137, N863, N184);
nand NAND2 (N1546, N1533, N1342);
xor XOR2 (N1547, N1545, N1522);
not NOT1 (N1548, N1544);
xor XOR2 (N1549, N1548, N344);
or OR2 (N1550, N1542, N1162);
xor XOR2 (N1551, N1521, N921);
not NOT1 (N1552, N1541);
nand NAND4 (N1553, N1546, N728, N1163, N375);
buf BUF1 (N1554, N1553);
not NOT1 (N1555, N1551);
buf BUF1 (N1556, N1536);
xor XOR2 (N1557, N1556, N62);
or OR4 (N1558, N1557, N303, N571, N771);
buf BUF1 (N1559, N1558);
nand NAND4 (N1560, N1550, N1105, N1288, N431);
not NOT1 (N1561, N1543);
not NOT1 (N1562, N1535);
buf BUF1 (N1563, N1528);
xor XOR2 (N1564, N1563, N207);
and AND4 (N1565, N1552, N1469, N83, N76);
nand NAND4 (N1566, N1560, N546, N345, N1200);
nor NOR2 (N1567, N1559, N1137);
nand NAND4 (N1568, N1561, N676, N1446, N127);
and AND4 (N1569, N1565, N1407, N134, N617);
buf BUF1 (N1570, N1564);
nor NOR2 (N1571, N1554, N1077);
not NOT1 (N1572, N1566);
buf BUF1 (N1573, N1549);
not NOT1 (N1574, N1569);
xor XOR2 (N1575, N1570, N832);
buf BUF1 (N1576, N1573);
buf BUF1 (N1577, N1568);
nand NAND3 (N1578, N1575, N1379, N616);
xor XOR2 (N1579, N1574, N1008);
or OR3 (N1580, N1567, N1304, N41);
or OR4 (N1581, N1547, N1201, N278, N1409);
or OR2 (N1582, N1581, N496);
or OR2 (N1583, N1572, N1268);
not NOT1 (N1584, N1576);
nor NOR4 (N1585, N1577, N994, N1175, N978);
or OR2 (N1586, N1583, N464);
nor NOR2 (N1587, N1582, N810);
or OR2 (N1588, N1586, N801);
or OR4 (N1589, N1588, N115, N148, N534);
not NOT1 (N1590, N1562);
buf BUF1 (N1591, N1585);
or OR4 (N1592, N1571, N1336, N1093, N1228);
buf BUF1 (N1593, N1589);
or OR3 (N1594, N1590, N881, N108);
or OR4 (N1595, N1584, N1388, N618, N761);
buf BUF1 (N1596, N1592);
and AND3 (N1597, N1587, N744, N1446);
nor NOR2 (N1598, N1580, N217);
buf BUF1 (N1599, N1593);
buf BUF1 (N1600, N1594);
buf BUF1 (N1601, N1591);
nor NOR2 (N1602, N1598, N1335);
and AND2 (N1603, N1599, N1390);
and AND3 (N1604, N1597, N164, N1386);
not NOT1 (N1605, N1579);
not NOT1 (N1606, N1601);
and AND3 (N1607, N1603, N763, N861);
buf BUF1 (N1608, N1605);
not NOT1 (N1609, N1604);
buf BUF1 (N1610, N1596);
or OR4 (N1611, N1600, N178, N1258, N1136);
buf BUF1 (N1612, N1595);
nor NOR2 (N1613, N1610, N1385);
buf BUF1 (N1614, N1611);
not NOT1 (N1615, N1578);
or OR4 (N1616, N1607, N610, N253, N145);
or OR4 (N1617, N1616, N1443, N1075, N1049);
xor XOR2 (N1618, N1613, N946);
and AND3 (N1619, N1606, N1575, N391);
buf BUF1 (N1620, N1615);
or OR3 (N1621, N1617, N1414, N583);
or OR3 (N1622, N1620, N758, N1579);
or OR2 (N1623, N1608, N504);
xor XOR2 (N1624, N1622, N1475);
and AND2 (N1625, N1612, N1100);
or OR4 (N1626, N1555, N1609, N1621, N1319);
nor NOR3 (N1627, N905, N155, N1436);
and AND4 (N1628, N1266, N971, N887, N655);
buf BUF1 (N1629, N1628);
xor XOR2 (N1630, N1602, N696);
buf BUF1 (N1631, N1624);
or OR3 (N1632, N1625, N113, N413);
xor XOR2 (N1633, N1614, N197);
xor XOR2 (N1634, N1619, N372);
xor XOR2 (N1635, N1634, N264);
xor XOR2 (N1636, N1630, N1252);
nor NOR3 (N1637, N1629, N849, N1018);
not NOT1 (N1638, N1623);
nor NOR3 (N1639, N1632, N379, N1007);
not NOT1 (N1640, N1636);
nor NOR4 (N1641, N1638, N507, N212, N96);
nand NAND4 (N1642, N1639, N38, N1607, N1354);
xor XOR2 (N1643, N1637, N600);
nor NOR3 (N1644, N1627, N951, N1303);
xor XOR2 (N1645, N1641, N775);
not NOT1 (N1646, N1642);
nand NAND3 (N1647, N1645, N1389, N1444);
nor NOR4 (N1648, N1640, N567, N1582, N1402);
or OR3 (N1649, N1647, N1388, N871);
or OR2 (N1650, N1618, N804);
nor NOR2 (N1651, N1648, N1612);
nand NAND3 (N1652, N1643, N687, N342);
nor NOR3 (N1653, N1626, N419, N204);
nand NAND4 (N1654, N1635, N1634, N1200, N595);
nand NAND3 (N1655, N1653, N1448, N430);
and AND4 (N1656, N1633, N1414, N237, N990);
nor NOR2 (N1657, N1650, N197);
nor NOR3 (N1658, N1657, N670, N1510);
xor XOR2 (N1659, N1655, N1346);
and AND2 (N1660, N1654, N551);
not NOT1 (N1661, N1660);
and AND2 (N1662, N1631, N1494);
not NOT1 (N1663, N1661);
and AND4 (N1664, N1644, N1447, N1032, N527);
nand NAND4 (N1665, N1658, N1239, N1061, N488);
not NOT1 (N1666, N1646);
or OR4 (N1667, N1659, N1139, N1470, N511);
not NOT1 (N1668, N1662);
nor NOR2 (N1669, N1656, N387);
xor XOR2 (N1670, N1664, N1387);
or OR2 (N1671, N1665, N632);
not NOT1 (N1672, N1666);
xor XOR2 (N1673, N1668, N889);
buf BUF1 (N1674, N1667);
nor NOR4 (N1675, N1669, N948, N285, N323);
xor XOR2 (N1676, N1670, N448);
or OR4 (N1677, N1663, N1655, N1084, N1593);
buf BUF1 (N1678, N1677);
and AND2 (N1679, N1651, N1483);
nand NAND4 (N1680, N1675, N126, N1601, N225);
not NOT1 (N1681, N1671);
xor XOR2 (N1682, N1674, N1369);
xor XOR2 (N1683, N1652, N478);
buf BUF1 (N1684, N1679);
not NOT1 (N1685, N1673);
buf BUF1 (N1686, N1682);
nand NAND3 (N1687, N1686, N521, N1029);
xor XOR2 (N1688, N1680, N1057);
not NOT1 (N1689, N1678);
or OR2 (N1690, N1683, N619);
buf BUF1 (N1691, N1689);
not NOT1 (N1692, N1688);
xor XOR2 (N1693, N1681, N337);
nand NAND2 (N1694, N1685, N1060);
not NOT1 (N1695, N1672);
or OR4 (N1696, N1695, N704, N949, N418);
not NOT1 (N1697, N1691);
nor NOR3 (N1698, N1690, N973, N1311);
and AND4 (N1699, N1698, N691, N712, N1258);
nand NAND2 (N1700, N1692, N322);
nor NOR2 (N1701, N1700, N1175);
nand NAND3 (N1702, N1693, N765, N804);
xor XOR2 (N1703, N1702, N241);
not NOT1 (N1704, N1694);
or OR2 (N1705, N1697, N1208);
not NOT1 (N1706, N1696);
xor XOR2 (N1707, N1699, N754);
not NOT1 (N1708, N1701);
buf BUF1 (N1709, N1676);
not NOT1 (N1710, N1706);
nand NAND4 (N1711, N1705, N171, N1203, N388);
not NOT1 (N1712, N1703);
or OR2 (N1713, N1708, N332);
not NOT1 (N1714, N1710);
not NOT1 (N1715, N1712);
xor XOR2 (N1716, N1713, N1351);
nand NAND4 (N1717, N1711, N237, N393, N216);
xor XOR2 (N1718, N1717, N1523);
buf BUF1 (N1719, N1715);
nand NAND3 (N1720, N1649, N1364, N315);
nor NOR2 (N1721, N1716, N1159);
not NOT1 (N1722, N1719);
nor NOR2 (N1723, N1721, N563);
nand NAND3 (N1724, N1704, N885, N1112);
nor NOR2 (N1725, N1723, N311);
and AND3 (N1726, N1687, N1203, N1070);
buf BUF1 (N1727, N1725);
or OR4 (N1728, N1718, N80, N200, N461);
nand NAND4 (N1729, N1722, N402, N1638, N1592);
or OR2 (N1730, N1726, N1461);
and AND2 (N1731, N1707, N138);
and AND3 (N1732, N1720, N608, N1668);
not NOT1 (N1733, N1730);
buf BUF1 (N1734, N1732);
buf BUF1 (N1735, N1684);
nand NAND2 (N1736, N1727, N1184);
not NOT1 (N1737, N1736);
xor XOR2 (N1738, N1729, N605);
buf BUF1 (N1739, N1735);
nand NAND2 (N1740, N1737, N1201);
nor NOR3 (N1741, N1740, N1252, N735);
xor XOR2 (N1742, N1741, N590);
xor XOR2 (N1743, N1728, N1601);
nand NAND2 (N1744, N1714, N177);
buf BUF1 (N1745, N1742);
and AND2 (N1746, N1724, N1161);
not NOT1 (N1747, N1743);
nand NAND3 (N1748, N1734, N749, N184);
and AND2 (N1749, N1748, N1521);
and AND2 (N1750, N1733, N1190);
buf BUF1 (N1751, N1731);
or OR2 (N1752, N1745, N1184);
and AND3 (N1753, N1746, N248, N1544);
and AND3 (N1754, N1744, N695, N1132);
xor XOR2 (N1755, N1751, N1085);
xor XOR2 (N1756, N1747, N158);
and AND2 (N1757, N1738, N172);
xor XOR2 (N1758, N1739, N887);
and AND2 (N1759, N1757, N501);
and AND4 (N1760, N1752, N154, N719, N1720);
and AND3 (N1761, N1709, N1734, N717);
buf BUF1 (N1762, N1749);
nand NAND2 (N1763, N1761, N1244);
buf BUF1 (N1764, N1759);
buf BUF1 (N1765, N1755);
and AND4 (N1766, N1760, N1116, N256, N1260);
xor XOR2 (N1767, N1766, N195);
xor XOR2 (N1768, N1753, N1417);
or OR3 (N1769, N1756, N1494, N1440);
not NOT1 (N1770, N1765);
and AND4 (N1771, N1770, N471, N1004, N772);
not NOT1 (N1772, N1758);
nor NOR2 (N1773, N1764, N1051);
not NOT1 (N1774, N1769);
buf BUF1 (N1775, N1754);
or OR4 (N1776, N1774, N1720, N22, N1457);
nor NOR2 (N1777, N1775, N567);
and AND2 (N1778, N1777, N1202);
nand NAND4 (N1779, N1778, N958, N144, N1649);
xor XOR2 (N1780, N1762, N1415);
nand NAND4 (N1781, N1773, N717, N575, N871);
and AND2 (N1782, N1780, N197);
not NOT1 (N1783, N1771);
or OR3 (N1784, N1763, N341, N11);
or OR4 (N1785, N1768, N807, N1013, N1747);
and AND3 (N1786, N1767, N370, N1241);
or OR4 (N1787, N1779, N248, N1448, N995);
nand NAND4 (N1788, N1782, N1010, N142, N1609);
nor NOR2 (N1789, N1772, N458);
nand NAND2 (N1790, N1789, N1378);
or OR3 (N1791, N1776, N1257, N1766);
or OR2 (N1792, N1785, N157);
nor NOR2 (N1793, N1750, N1466);
or OR4 (N1794, N1783, N781, N424, N1090);
and AND4 (N1795, N1790, N136, N669, N622);
nor NOR3 (N1796, N1794, N779, N433);
nor NOR2 (N1797, N1781, N534);
and AND2 (N1798, N1784, N562);
xor XOR2 (N1799, N1793, N1492);
buf BUF1 (N1800, N1791);
and AND4 (N1801, N1797, N1601, N32, N929);
nand NAND4 (N1802, N1788, N545, N1620, N1095);
nand NAND3 (N1803, N1801, N762, N1422);
and AND3 (N1804, N1787, N77, N221);
xor XOR2 (N1805, N1798, N646);
nor NOR4 (N1806, N1803, N1317, N82, N1071);
nor NOR2 (N1807, N1804, N298);
nor NOR2 (N1808, N1807, N547);
nand NAND3 (N1809, N1808, N113, N1214);
or OR3 (N1810, N1809, N395, N1775);
nand NAND3 (N1811, N1796, N1479, N285);
not NOT1 (N1812, N1786);
and AND4 (N1813, N1811, N1385, N424, N1313);
buf BUF1 (N1814, N1810);
not NOT1 (N1815, N1800);
nand NAND2 (N1816, N1805, N1654);
and AND4 (N1817, N1806, N1650, N1419, N974);
or OR4 (N1818, N1813, N836, N1366, N722);
and AND4 (N1819, N1812, N1724, N641, N1544);
and AND3 (N1820, N1815, N821, N260);
or OR2 (N1821, N1817, N333);
or OR3 (N1822, N1802, N1295, N722);
buf BUF1 (N1823, N1792);
not NOT1 (N1824, N1823);
nor NOR3 (N1825, N1819, N250, N1120);
xor XOR2 (N1826, N1820, N1538);
nor NOR3 (N1827, N1818, N1443, N1273);
nand NAND3 (N1828, N1825, N1640, N1303);
nor NOR2 (N1829, N1816, N322);
or OR2 (N1830, N1824, N342);
and AND3 (N1831, N1822, N577, N346);
and AND3 (N1832, N1795, N1056, N188);
nor NOR3 (N1833, N1830, N200, N505);
not NOT1 (N1834, N1829);
nor NOR3 (N1835, N1814, N652, N500);
nor NOR4 (N1836, N1831, N63, N1556, N149);
nor NOR3 (N1837, N1828, N1441, N586);
or OR2 (N1838, N1837, N1809);
or OR3 (N1839, N1834, N1795, N826);
buf BUF1 (N1840, N1839);
and AND3 (N1841, N1821, N1798, N499);
or OR4 (N1842, N1836, N389, N1133, N95);
and AND2 (N1843, N1826, N669);
nor NOR2 (N1844, N1835, N777);
and AND4 (N1845, N1843, N147, N315, N141);
not NOT1 (N1846, N1838);
not NOT1 (N1847, N1840);
or OR2 (N1848, N1844, N1521);
not NOT1 (N1849, N1799);
not NOT1 (N1850, N1846);
or OR4 (N1851, N1848, N1021, N28, N1087);
and AND2 (N1852, N1850, N31);
xor XOR2 (N1853, N1851, N770);
buf BUF1 (N1854, N1827);
buf BUF1 (N1855, N1842);
not NOT1 (N1856, N1853);
and AND3 (N1857, N1855, N807, N247);
not NOT1 (N1858, N1845);
nand NAND2 (N1859, N1852, N1519);
buf BUF1 (N1860, N1859);
and AND4 (N1861, N1856, N1153, N1471, N1840);
buf BUF1 (N1862, N1847);
nor NOR2 (N1863, N1833, N1477);
buf BUF1 (N1864, N1849);
not NOT1 (N1865, N1854);
and AND3 (N1866, N1860, N606, N1001);
xor XOR2 (N1867, N1862, N257);
xor XOR2 (N1868, N1861, N1205);
not NOT1 (N1869, N1867);
nand NAND2 (N1870, N1865, N1172);
or OR3 (N1871, N1869, N1126, N1335);
not NOT1 (N1872, N1870);
and AND4 (N1873, N1858, N1175, N1047, N142);
and AND2 (N1874, N1863, N1250);
and AND4 (N1875, N1864, N301, N1444, N477);
buf BUF1 (N1876, N1872);
xor XOR2 (N1877, N1873, N1184);
buf BUF1 (N1878, N1874);
nand NAND3 (N1879, N1868, N1311, N1079);
xor XOR2 (N1880, N1879, N1322);
and AND4 (N1881, N1875, N57, N1143, N1850);
nand NAND2 (N1882, N1871, N181);
and AND3 (N1883, N1882, N802, N877);
not NOT1 (N1884, N1876);
and AND4 (N1885, N1880, N1468, N1044, N1300);
buf BUF1 (N1886, N1878);
or OR3 (N1887, N1886, N1451, N927);
nor NOR4 (N1888, N1832, N1205, N1261, N1793);
nand NAND2 (N1889, N1877, N1189);
not NOT1 (N1890, N1881);
and AND4 (N1891, N1866, N83, N1802, N372);
not NOT1 (N1892, N1857);
xor XOR2 (N1893, N1841, N444);
xor XOR2 (N1894, N1884, N94);
nand NAND2 (N1895, N1892, N355);
nand NAND4 (N1896, N1889, N1012, N407, N317);
nor NOR3 (N1897, N1890, N689, N386);
nor NOR4 (N1898, N1885, N977, N1624, N1060);
and AND3 (N1899, N1888, N1665, N906);
nand NAND3 (N1900, N1883, N1588, N152);
nand NAND4 (N1901, N1895, N1764, N1421, N764);
nand NAND2 (N1902, N1894, N1721);
not NOT1 (N1903, N1900);
nor NOR4 (N1904, N1887, N318, N1754, N306);
nor NOR4 (N1905, N1893, N1446, N10, N1153);
or OR4 (N1906, N1891, N756, N1388, N330);
not NOT1 (N1907, N1898);
nor NOR2 (N1908, N1905, N1758);
xor XOR2 (N1909, N1899, N1537);
buf BUF1 (N1910, N1904);
not NOT1 (N1911, N1906);
xor XOR2 (N1912, N1903, N795);
buf BUF1 (N1913, N1902);
not NOT1 (N1914, N1896);
or OR2 (N1915, N1908, N721);
or OR3 (N1916, N1901, N1039, N1204);
and AND4 (N1917, N1910, N1326, N1716, N94);
nand NAND3 (N1918, N1911, N1202, N1432);
not NOT1 (N1919, N1916);
nor NOR4 (N1920, N1915, N495, N54, N2);
buf BUF1 (N1921, N1912);
buf BUF1 (N1922, N1913);
not NOT1 (N1923, N1897);
nand NAND3 (N1924, N1918, N521, N886);
xor XOR2 (N1925, N1907, N1567);
buf BUF1 (N1926, N1914);
nand NAND2 (N1927, N1921, N1896);
buf BUF1 (N1928, N1926);
nand NAND4 (N1929, N1922, N28, N1899, N364);
xor XOR2 (N1930, N1928, N1821);
xor XOR2 (N1931, N1917, N461);
xor XOR2 (N1932, N1919, N755);
or OR4 (N1933, N1923, N656, N119, N1119);
nand NAND4 (N1934, N1931, N263, N1228, N211);
xor XOR2 (N1935, N1929, N974);
not NOT1 (N1936, N1932);
and AND2 (N1937, N1924, N373);
nor NOR4 (N1938, N1925, N849, N246, N918);
and AND3 (N1939, N1927, N199, N753);
or OR3 (N1940, N1937, N1801, N781);
buf BUF1 (N1941, N1936);
nand NAND4 (N1942, N1940, N1416, N15, N490);
not NOT1 (N1943, N1941);
not NOT1 (N1944, N1934);
and AND4 (N1945, N1909, N1814, N534, N1195);
buf BUF1 (N1946, N1935);
buf BUF1 (N1947, N1938);
and AND2 (N1948, N1947, N1253);
not NOT1 (N1949, N1939);
or OR4 (N1950, N1948, N586, N1467, N1718);
buf BUF1 (N1951, N1945);
and AND4 (N1952, N1943, N952, N304, N1381);
and AND3 (N1953, N1952, N684, N1200);
and AND3 (N1954, N1920, N1306, N879);
or OR2 (N1955, N1930, N1574);
or OR3 (N1956, N1949, N1760, N1507);
and AND2 (N1957, N1933, N1166);
buf BUF1 (N1958, N1944);
nor NOR2 (N1959, N1951, N511);
nor NOR4 (N1960, N1953, N1862, N733, N1521);
xor XOR2 (N1961, N1950, N1897);
buf BUF1 (N1962, N1942);
nand NAND2 (N1963, N1958, N47);
xor XOR2 (N1964, N1955, N957);
xor XOR2 (N1965, N1964, N248);
nand NAND2 (N1966, N1961, N550);
and AND3 (N1967, N1956, N1328, N1146);
nand NAND2 (N1968, N1959, N1873);
nand NAND3 (N1969, N1946, N1430, N1848);
or OR2 (N1970, N1962, N243);
buf BUF1 (N1971, N1967);
not NOT1 (N1972, N1966);
and AND3 (N1973, N1968, N476, N324);
buf BUF1 (N1974, N1972);
buf BUF1 (N1975, N1973);
nand NAND3 (N1976, N1975, N648, N1065);
nor NOR4 (N1977, N1960, N934, N182, N1755);
nand NAND2 (N1978, N1976, N308);
not NOT1 (N1979, N1970);
buf BUF1 (N1980, N1957);
buf BUF1 (N1981, N1977);
nor NOR4 (N1982, N1974, N1237, N489, N960);
xor XOR2 (N1983, N1979, N160);
not NOT1 (N1984, N1954);
xor XOR2 (N1985, N1980, N27);
and AND2 (N1986, N1965, N478);
not NOT1 (N1987, N1984);
xor XOR2 (N1988, N1983, N260);
xor XOR2 (N1989, N1987, N1233);
or OR2 (N1990, N1981, N774);
not NOT1 (N1991, N1986);
nand NAND3 (N1992, N1985, N643, N430);
and AND4 (N1993, N1963, N1936, N1788, N1598);
nor NOR2 (N1994, N1982, N1986);
and AND2 (N1995, N1994, N1409);
and AND2 (N1996, N1993, N513);
xor XOR2 (N1997, N1989, N229);
or OR4 (N1998, N1995, N1474, N1289, N1970);
buf BUF1 (N1999, N1991);
xor XOR2 (N2000, N1969, N205);
xor XOR2 (N2001, N1998, N529);
nor NOR2 (N2002, N1999, N1176);
nand NAND2 (N2003, N1971, N988);
nand NAND3 (N2004, N2003, N1374, N2000);
and AND3 (N2005, N1486, N1629, N1805);
nor NOR4 (N2006, N1990, N151, N1084, N748);
nor NOR2 (N2007, N2002, N1720);
nor NOR3 (N2008, N2005, N1284, N1613);
and AND2 (N2009, N2008, N775);
nor NOR3 (N2010, N1996, N1675, N825);
and AND4 (N2011, N2007, N1497, N292, N342);
buf BUF1 (N2012, N2006);
not NOT1 (N2013, N2001);
not NOT1 (N2014, N1997);
nand NAND2 (N2015, N2011, N1372);
buf BUF1 (N2016, N2015);
not NOT1 (N2017, N2012);
or OR3 (N2018, N1992, N1138, N586);
not NOT1 (N2019, N2010);
xor XOR2 (N2020, N2009, N903);
not NOT1 (N2021, N2004);
nand NAND2 (N2022, N2018, N1795);
nand NAND3 (N2023, N2022, N1554, N1903);
xor XOR2 (N2024, N2021, N886);
nand NAND3 (N2025, N2024, N1000, N57);
or OR2 (N2026, N2023, N314);
and AND2 (N2027, N2026, N1652);
nor NOR4 (N2028, N1988, N655, N211, N1364);
not NOT1 (N2029, N2025);
nand NAND2 (N2030, N2017, N879);
or OR3 (N2031, N2028, N529, N1730);
or OR3 (N2032, N2019, N269, N1960);
buf BUF1 (N2033, N2016);
buf BUF1 (N2034, N1978);
nand NAND2 (N2035, N2029, N755);
nor NOR3 (N2036, N2013, N1120, N1934);
and AND4 (N2037, N2031, N827, N1306, N1717);
buf BUF1 (N2038, N2037);
or OR4 (N2039, N2014, N1455, N625, N1387);
buf BUF1 (N2040, N2039);
not NOT1 (N2041, N2033);
not NOT1 (N2042, N2035);
and AND4 (N2043, N2032, N939, N1141, N1448);
nor NOR3 (N2044, N2042, N423, N531);
buf BUF1 (N2045, N2027);
and AND3 (N2046, N2038, N1655, N827);
and AND4 (N2047, N2036, N1394, N1276, N1204);
nor NOR2 (N2048, N2030, N117);
nand NAND4 (N2049, N2040, N1837, N1035, N1447);
nand NAND3 (N2050, N2020, N1377, N1170);
nand NAND4 (N2051, N2047, N822, N319, N1351);
xor XOR2 (N2052, N2049, N239);
buf BUF1 (N2053, N2043);
xor XOR2 (N2054, N2034, N1836);
and AND4 (N2055, N2048, N1968, N1938, N259);
nand NAND4 (N2056, N2041, N1546, N622, N972);
nor NOR2 (N2057, N2051, N1069);
and AND4 (N2058, N2055, N139, N1238, N1537);
nor NOR4 (N2059, N2054, N840, N1791, N963);
or OR2 (N2060, N2056, N957);
nor NOR3 (N2061, N2058, N1923, N1232);
xor XOR2 (N2062, N2045, N144);
xor XOR2 (N2063, N2050, N1485);
or OR4 (N2064, N2044, N270, N86, N325);
xor XOR2 (N2065, N2063, N1634);
buf BUF1 (N2066, N2064);
and AND4 (N2067, N2066, N1356, N1534, N369);
xor XOR2 (N2068, N2052, N1441);
not NOT1 (N2069, N2062);
or OR4 (N2070, N2061, N1383, N1043, N12);
or OR2 (N2071, N2065, N436);
and AND4 (N2072, N2070, N2068, N1010, N436);
and AND4 (N2073, N1491, N392, N1781, N1003);
xor XOR2 (N2074, N2053, N1714);
and AND4 (N2075, N2069, N1234, N1746, N1271);
or OR2 (N2076, N2057, N255);
or OR2 (N2077, N2075, N1398);
buf BUF1 (N2078, N2046);
xor XOR2 (N2079, N2077, N227);
and AND2 (N2080, N2073, N651);
nor NOR3 (N2081, N2080, N43, N1265);
nor NOR3 (N2082, N2067, N1094, N812);
buf BUF1 (N2083, N2076);
nand NAND2 (N2084, N2082, N498);
not NOT1 (N2085, N2059);
buf BUF1 (N2086, N2081);
buf BUF1 (N2087, N2083);
nor NOR3 (N2088, N2072, N588, N1269);
not NOT1 (N2089, N2088);
nor NOR3 (N2090, N2074, N184, N1494);
nand NAND3 (N2091, N2085, N1862, N728);
nor NOR3 (N2092, N2060, N402, N225);
buf BUF1 (N2093, N2079);
not NOT1 (N2094, N2071);
and AND3 (N2095, N2084, N1163, N1876);
and AND4 (N2096, N2093, N1213, N1158, N2048);
xor XOR2 (N2097, N2086, N105);
and AND4 (N2098, N2097, N1885, N1938, N1300);
xor XOR2 (N2099, N2078, N1210);
not NOT1 (N2100, N2087);
xor XOR2 (N2101, N2099, N946);
nand NAND3 (N2102, N2092, N231, N349);
xor XOR2 (N2103, N2101, N1401);
and AND4 (N2104, N2095, N418, N1295, N604);
not NOT1 (N2105, N2102);
not NOT1 (N2106, N2089);
nand NAND2 (N2107, N2103, N1216);
or OR4 (N2108, N2096, N886, N1618, N717);
nor NOR3 (N2109, N2098, N741, N604);
or OR3 (N2110, N2109, N1437, N2043);
nand NAND2 (N2111, N2107, N598);
xor XOR2 (N2112, N2091, N1806);
or OR2 (N2113, N2104, N809);
xor XOR2 (N2114, N2105, N688);
nor NOR3 (N2115, N2112, N1409, N1784);
or OR2 (N2116, N2115, N991);
and AND4 (N2117, N2110, N2029, N1595, N874);
nand NAND2 (N2118, N2108, N1786);
or OR4 (N2119, N2118, N887, N2094, N498);
buf BUF1 (N2120, N437);
nand NAND4 (N2121, N2106, N252, N1623, N1749);
or OR4 (N2122, N2119, N168, N994, N1465);
nor NOR3 (N2123, N2114, N153, N1030);
nor NOR4 (N2124, N2090, N1808, N1137, N1727);
buf BUF1 (N2125, N2111);
or OR2 (N2126, N2125, N1989);
or OR4 (N2127, N2117, N630, N1782, N2076);
xor XOR2 (N2128, N2124, N858);
or OR2 (N2129, N2120, N898);
not NOT1 (N2130, N2113);
not NOT1 (N2131, N2116);
or OR4 (N2132, N2130, N1577, N196, N1464);
or OR4 (N2133, N2127, N2104, N1414, N1512);
xor XOR2 (N2134, N2122, N2109);
xor XOR2 (N2135, N2128, N660);
nor NOR2 (N2136, N2129, N217);
and AND3 (N2137, N2136, N1818, N1319);
nand NAND2 (N2138, N2132, N1768);
or OR4 (N2139, N2126, N44, N564, N1383);
not NOT1 (N2140, N2133);
or OR3 (N2141, N2138, N977, N1637);
nor NOR3 (N2142, N2137, N1546, N1862);
buf BUF1 (N2143, N2139);
or OR3 (N2144, N2121, N446, N1922);
or OR2 (N2145, N2141, N243);
buf BUF1 (N2146, N2134);
buf BUF1 (N2147, N2145);
or OR3 (N2148, N2135, N1857, N1952);
and AND2 (N2149, N2131, N786);
xor XOR2 (N2150, N2140, N1482);
nor NOR4 (N2151, N2100, N611, N939, N1830);
buf BUF1 (N2152, N2150);
buf BUF1 (N2153, N2147);
or OR2 (N2154, N2149, N647);
buf BUF1 (N2155, N2123);
and AND2 (N2156, N2148, N271);
and AND4 (N2157, N2154, N1987, N606, N2016);
xor XOR2 (N2158, N2146, N1924);
xor XOR2 (N2159, N2155, N272);
xor XOR2 (N2160, N2158, N1388);
and AND3 (N2161, N2142, N769, N622);
buf BUF1 (N2162, N2157);
xor XOR2 (N2163, N2152, N731);
xor XOR2 (N2164, N2156, N814);
nor NOR4 (N2165, N2161, N812, N320, N1861);
nor NOR4 (N2166, N2164, N1606, N1212, N138);
nor NOR3 (N2167, N2166, N518, N2046);
or OR4 (N2168, N2143, N794, N998, N619);
not NOT1 (N2169, N2160);
nand NAND2 (N2170, N2165, N70);
not NOT1 (N2171, N2163);
or OR4 (N2172, N2169, N958, N1576, N643);
xor XOR2 (N2173, N2167, N509);
nor NOR4 (N2174, N2172, N626, N1667, N1521);
xor XOR2 (N2175, N2171, N713);
xor XOR2 (N2176, N2174, N1234);
not NOT1 (N2177, N2168);
xor XOR2 (N2178, N2176, N880);
or OR4 (N2179, N2153, N1383, N139, N758);
xor XOR2 (N2180, N2178, N2076);
and AND4 (N2181, N2173, N1733, N2178, N1749);
not NOT1 (N2182, N2159);
xor XOR2 (N2183, N2179, N1212);
xor XOR2 (N2184, N2180, N142);
nor NOR3 (N2185, N2177, N1890, N1557);
xor XOR2 (N2186, N2162, N410);
xor XOR2 (N2187, N2175, N1490);
not NOT1 (N2188, N2170);
not NOT1 (N2189, N2184);
nand NAND2 (N2190, N2181, N998);
nor NOR4 (N2191, N2187, N1207, N632, N1758);
nor NOR3 (N2192, N2151, N430, N255);
nand NAND2 (N2193, N2186, N1593);
xor XOR2 (N2194, N2191, N1875);
nand NAND3 (N2195, N2189, N1953, N978);
and AND3 (N2196, N2185, N249, N1065);
xor XOR2 (N2197, N2196, N833);
buf BUF1 (N2198, N2144);
nor NOR3 (N2199, N2183, N1673, N1658);
nand NAND4 (N2200, N2194, N201, N1937, N1785);
or OR3 (N2201, N2199, N398, N546);
buf BUF1 (N2202, N2201);
buf BUF1 (N2203, N2190);
buf BUF1 (N2204, N2188);
nand NAND2 (N2205, N2197, N1051);
or OR2 (N2206, N2198, N1528);
or OR3 (N2207, N2195, N1515, N834);
not NOT1 (N2208, N2192);
not NOT1 (N2209, N2208);
nor NOR4 (N2210, N2205, N853, N1632, N1557);
nand NAND3 (N2211, N2207, N1005, N1866);
nand NAND2 (N2212, N2202, N1882);
not NOT1 (N2213, N2204);
xor XOR2 (N2214, N2213, N1198);
buf BUF1 (N2215, N2200);
nor NOR4 (N2216, N2203, N319, N1861, N697);
not NOT1 (N2217, N2216);
and AND4 (N2218, N2182, N1345, N622, N156);
buf BUF1 (N2219, N2212);
xor XOR2 (N2220, N2219, N367);
nand NAND4 (N2221, N2218, N1837, N2087, N1894);
nand NAND2 (N2222, N2206, N218);
and AND2 (N2223, N2217, N81);
buf BUF1 (N2224, N2222);
nand NAND2 (N2225, N2220, N1910);
xor XOR2 (N2226, N2224, N1685);
and AND4 (N2227, N2209, N38, N139, N1590);
nor NOR2 (N2228, N2211, N1331);
nand NAND4 (N2229, N2210, N1457, N1051, N646);
buf BUF1 (N2230, N2223);
nor NOR4 (N2231, N2221, N1843, N1932, N1626);
nand NAND3 (N2232, N2227, N1166, N1696);
nor NOR3 (N2233, N2215, N1793, N1085);
xor XOR2 (N2234, N2225, N556);
or OR2 (N2235, N2230, N1253);
xor XOR2 (N2236, N2232, N136);
and AND4 (N2237, N2193, N1826, N905, N1359);
or OR4 (N2238, N2228, N1610, N1599, N1570);
and AND3 (N2239, N2231, N770, N441);
nor NOR2 (N2240, N2226, N1893);
not NOT1 (N2241, N2214);
not NOT1 (N2242, N2229);
buf BUF1 (N2243, N2234);
or OR2 (N2244, N2241, N1662);
not NOT1 (N2245, N2235);
or OR2 (N2246, N2244, N2229);
nand NAND4 (N2247, N2239, N341, N1487, N278);
xor XOR2 (N2248, N2233, N1823);
and AND3 (N2249, N2236, N1742, N586);
and AND2 (N2250, N2237, N1192);
or OR3 (N2251, N2242, N1316, N325);
or OR4 (N2252, N2238, N394, N2018, N1951);
nor NOR3 (N2253, N2247, N933, N734);
nor NOR4 (N2254, N2249, N883, N29, N481);
nor NOR2 (N2255, N2253, N1496);
nand NAND4 (N2256, N2243, N1027, N1467, N1433);
or OR2 (N2257, N2240, N1906);
or OR3 (N2258, N2245, N1895, N603);
and AND4 (N2259, N2246, N1708, N605, N278);
nand NAND4 (N2260, N2254, N1793, N1116, N2219);
nor NOR4 (N2261, N2255, N1836, N1483, N1483);
nand NAND3 (N2262, N2261, N84, N1670);
nor NOR2 (N2263, N2262, N224);
xor XOR2 (N2264, N2257, N1793);
and AND2 (N2265, N2251, N1022);
buf BUF1 (N2266, N2263);
nor NOR4 (N2267, N2259, N468, N757, N967);
nand NAND2 (N2268, N2266, N409);
xor XOR2 (N2269, N2260, N1307);
xor XOR2 (N2270, N2258, N908);
buf BUF1 (N2271, N2252);
or OR4 (N2272, N2248, N932, N2203, N2263);
not NOT1 (N2273, N2268);
xor XOR2 (N2274, N2267, N1097);
nor NOR3 (N2275, N2269, N1817, N1223);
not NOT1 (N2276, N2250);
nor NOR4 (N2277, N2275, N202, N1418, N455);
and AND4 (N2278, N2272, N1487, N1832, N129);
xor XOR2 (N2279, N2271, N866);
xor XOR2 (N2280, N2270, N158);
buf BUF1 (N2281, N2264);
buf BUF1 (N2282, N2280);
buf BUF1 (N2283, N2277);
buf BUF1 (N2284, N2276);
not NOT1 (N2285, N2256);
buf BUF1 (N2286, N2282);
not NOT1 (N2287, N2279);
nand NAND2 (N2288, N2278, N943);
xor XOR2 (N2289, N2286, N319);
xor XOR2 (N2290, N2274, N978);
or OR2 (N2291, N2265, N1558);
nand NAND2 (N2292, N2283, N1539);
and AND3 (N2293, N2285, N800, N1006);
nand NAND2 (N2294, N2284, N239);
buf BUF1 (N2295, N2273);
nand NAND4 (N2296, N2290, N635, N1942, N800);
not NOT1 (N2297, N2289);
nand NAND2 (N2298, N2293, N1479);
nand NAND3 (N2299, N2298, N926, N1485);
buf BUF1 (N2300, N2287);
buf BUF1 (N2301, N2294);
and AND2 (N2302, N2300, N581);
nand NAND2 (N2303, N2301, N647);
xor XOR2 (N2304, N2303, N1911);
not NOT1 (N2305, N2296);
nor NOR2 (N2306, N2302, N1038);
nor NOR4 (N2307, N2299, N2184, N957, N1958);
nand NAND4 (N2308, N2291, N152, N2207, N1429);
not NOT1 (N2309, N2308);
or OR2 (N2310, N2292, N146);
not NOT1 (N2311, N2305);
or OR4 (N2312, N2306, N1781, N1981, N2028);
nand NAND4 (N2313, N2295, N1373, N645, N1311);
and AND2 (N2314, N2281, N839);
xor XOR2 (N2315, N2304, N2308);
xor XOR2 (N2316, N2311, N759);
nor NOR2 (N2317, N2297, N2245);
buf BUF1 (N2318, N2314);
xor XOR2 (N2319, N2307, N664);
or OR4 (N2320, N2319, N632, N863, N1010);
nand NAND4 (N2321, N2316, N1740, N593, N834);
xor XOR2 (N2322, N2321, N487);
nand NAND2 (N2323, N2312, N1268);
buf BUF1 (N2324, N2317);
or OR2 (N2325, N2318, N797);
nor NOR3 (N2326, N2310, N2236, N821);
not NOT1 (N2327, N2322);
buf BUF1 (N2328, N2315);
buf BUF1 (N2329, N2323);
not NOT1 (N2330, N2328);
nor NOR2 (N2331, N2326, N2075);
nor NOR2 (N2332, N2330, N994);
not NOT1 (N2333, N2329);
or OR2 (N2334, N2288, N978);
xor XOR2 (N2335, N2325, N1845);
nor NOR3 (N2336, N2331, N820, N131);
nor NOR2 (N2337, N2320, N2310);
nor NOR3 (N2338, N2327, N2247, N2006);
not NOT1 (N2339, N2309);
buf BUF1 (N2340, N2337);
nand NAND2 (N2341, N2340, N873);
nor NOR4 (N2342, N2335, N1207, N50, N2231);
and AND2 (N2343, N2333, N1301);
or OR4 (N2344, N2338, N1400, N737, N1359);
buf BUF1 (N2345, N2324);
xor XOR2 (N2346, N2345, N722);
nor NOR2 (N2347, N2339, N778);
nand NAND2 (N2348, N2342, N217);
nand NAND2 (N2349, N2341, N2075);
not NOT1 (N2350, N2334);
and AND2 (N2351, N2348, N1286);
and AND2 (N2352, N2351, N467);
xor XOR2 (N2353, N2347, N1154);
nor NOR2 (N2354, N2332, N542);
xor XOR2 (N2355, N2346, N1348);
nor NOR3 (N2356, N2349, N1302, N1661);
nor NOR3 (N2357, N2355, N1772, N142);
nor NOR4 (N2358, N2313, N388, N522, N1509);
nand NAND4 (N2359, N2358, N1398, N337, N234);
xor XOR2 (N2360, N2343, N1229);
nor NOR4 (N2361, N2344, N1310, N236, N2111);
buf BUF1 (N2362, N2356);
or OR2 (N2363, N2354, N222);
not NOT1 (N2364, N2360);
nand NAND2 (N2365, N2352, N342);
not NOT1 (N2366, N2336);
and AND3 (N2367, N2357, N1332, N239);
nand NAND4 (N2368, N2353, N1284, N51, N1388);
not NOT1 (N2369, N2350);
nand NAND2 (N2370, N2368, N1626);
xor XOR2 (N2371, N2366, N256);
and AND4 (N2372, N2364, N488, N1609, N1349);
or OR2 (N2373, N2370, N1052);
not NOT1 (N2374, N2359);
nand NAND3 (N2375, N2371, N1447, N1895);
xor XOR2 (N2376, N2365, N385);
nand NAND4 (N2377, N2373, N2275, N1661, N1959);
nor NOR4 (N2378, N2377, N2296, N1700, N122);
nand NAND2 (N2379, N2376, N2159);
buf BUF1 (N2380, N2372);
nand NAND2 (N2381, N2374, N2356);
buf BUF1 (N2382, N2378);
buf BUF1 (N2383, N2369);
not NOT1 (N2384, N2361);
buf BUF1 (N2385, N2383);
nor NOR2 (N2386, N2384, N2114);
buf BUF1 (N2387, N2379);
buf BUF1 (N2388, N2375);
buf BUF1 (N2389, N2363);
buf BUF1 (N2390, N2381);
xor XOR2 (N2391, N2386, N1376);
or OR2 (N2392, N2391, N457);
or OR4 (N2393, N2385, N1525, N1641, N470);
nor NOR3 (N2394, N2382, N158, N1471);
xor XOR2 (N2395, N2389, N564);
xor XOR2 (N2396, N2394, N1924);
xor XOR2 (N2397, N2367, N564);
nor NOR4 (N2398, N2388, N912, N2353, N310);
or OR3 (N2399, N2380, N997, N374);
nand NAND2 (N2400, N2362, N1608);
nand NAND3 (N2401, N2399, N258, N1269);
buf BUF1 (N2402, N2396);
nor NOR2 (N2403, N2401, N161);
nor NOR3 (N2404, N2402, N1892, N906);
buf BUF1 (N2405, N2400);
xor XOR2 (N2406, N2403, N2312);
or OR3 (N2407, N2393, N532, N2126);
not NOT1 (N2408, N2392);
nor NOR4 (N2409, N2387, N192, N559, N769);
or OR3 (N2410, N2407, N1131, N1226);
xor XOR2 (N2411, N2408, N2138);
nor NOR2 (N2412, N2405, N1872);
or OR4 (N2413, N2398, N1980, N1761, N1644);
nand NAND3 (N2414, N2404, N1449, N2158);
and AND3 (N2415, N2410, N1890, N1380);
nor NOR2 (N2416, N2412, N2167);
nor NOR2 (N2417, N2397, N1214);
and AND2 (N2418, N2414, N926);
nand NAND2 (N2419, N2409, N1949);
nor NOR3 (N2420, N2416, N2223, N763);
or OR3 (N2421, N2420, N556, N937);
xor XOR2 (N2422, N2413, N769);
nor NOR4 (N2423, N2411, N2280, N467, N2415);
xor XOR2 (N2424, N1020, N905);
buf BUF1 (N2425, N2418);
nor NOR4 (N2426, N2425, N546, N639, N2303);
buf BUF1 (N2427, N2423);
not NOT1 (N2428, N2390);
and AND2 (N2429, N2422, N1316);
xor XOR2 (N2430, N2428, N1520);
xor XOR2 (N2431, N2417, N1953);
nand NAND4 (N2432, N2406, N181, N1775, N68);
buf BUF1 (N2433, N2427);
or OR3 (N2434, N2433, N405, N614);
nand NAND4 (N2435, N2421, N1370, N2142, N539);
buf BUF1 (N2436, N2395);
xor XOR2 (N2437, N2435, N899);
not NOT1 (N2438, N2419);
and AND2 (N2439, N2426, N224);
not NOT1 (N2440, N2438);
nor NOR4 (N2441, N2440, N592, N1480, N1742);
xor XOR2 (N2442, N2441, N1875);
or OR2 (N2443, N2429, N223);
buf BUF1 (N2444, N2424);
nor NOR4 (N2445, N2432, N2100, N277, N794);
not NOT1 (N2446, N2431);
xor XOR2 (N2447, N2443, N2399);
buf BUF1 (N2448, N2446);
buf BUF1 (N2449, N2437);
nand NAND2 (N2450, N2430, N356);
or OR3 (N2451, N2434, N618, N188);
xor XOR2 (N2452, N2436, N2132);
buf BUF1 (N2453, N2452);
buf BUF1 (N2454, N2450);
or OR4 (N2455, N2454, N1585, N53, N950);
and AND3 (N2456, N2439, N118, N1827);
nand NAND4 (N2457, N2444, N2283, N100, N271);
xor XOR2 (N2458, N2453, N603);
xor XOR2 (N2459, N2447, N622);
xor XOR2 (N2460, N2456, N1054);
nand NAND4 (N2461, N2445, N367, N1242, N713);
and AND3 (N2462, N2458, N171, N1699);
nand NAND2 (N2463, N2448, N1574);
and AND4 (N2464, N2442, N729, N1244, N571);
not NOT1 (N2465, N2462);
or OR4 (N2466, N2459, N438, N160, N2290);
nand NAND2 (N2467, N2463, N1439);
not NOT1 (N2468, N2461);
or OR3 (N2469, N2464, N1465, N823);
or OR4 (N2470, N2451, N1675, N2281, N599);
buf BUF1 (N2471, N2466);
nand NAND2 (N2472, N2469, N2310);
nor NOR3 (N2473, N2471, N203, N699);
nor NOR2 (N2474, N2473, N1321);
or OR4 (N2475, N2472, N1562, N1671, N915);
nand NAND4 (N2476, N2470, N1450, N750, N1632);
buf BUF1 (N2477, N2455);
and AND2 (N2478, N2449, N647);
and AND3 (N2479, N2477, N1461, N702);
not NOT1 (N2480, N2460);
xor XOR2 (N2481, N2467, N1920);
and AND3 (N2482, N2475, N2431, N2021);
and AND2 (N2483, N2474, N1208);
or OR2 (N2484, N2478, N1352);
and AND2 (N2485, N2479, N118);
nand NAND2 (N2486, N2468, N352);
nand NAND3 (N2487, N2481, N2149, N648);
or OR4 (N2488, N2465, N1841, N1870, N1084);
or OR4 (N2489, N2487, N950, N2103, N1751);
xor XOR2 (N2490, N2483, N2079);
not NOT1 (N2491, N2476);
xor XOR2 (N2492, N2490, N764);
nand NAND4 (N2493, N2482, N97, N315, N1540);
and AND4 (N2494, N2457, N2372, N1705, N2024);
xor XOR2 (N2495, N2489, N482);
not NOT1 (N2496, N2485);
xor XOR2 (N2497, N2486, N624);
xor XOR2 (N2498, N2480, N1229);
nand NAND3 (N2499, N2494, N189, N248);
nand NAND3 (N2500, N2496, N374, N400);
not NOT1 (N2501, N2491);
or OR3 (N2502, N2484, N350, N2306);
or OR2 (N2503, N2492, N2437);
not NOT1 (N2504, N2488);
or OR2 (N2505, N2499, N1801);
and AND3 (N2506, N2502, N260, N1932);
or OR3 (N2507, N2495, N945, N176);
nor NOR3 (N2508, N2507, N564, N255);
buf BUF1 (N2509, N2503);
nand NAND2 (N2510, N2505, N637);
buf BUF1 (N2511, N2509);
nand NAND3 (N2512, N2501, N2384, N918);
nor NOR2 (N2513, N2498, N1059);
xor XOR2 (N2514, N2493, N1333);
nand NAND2 (N2515, N2506, N1199);
xor XOR2 (N2516, N2508, N1008);
xor XOR2 (N2517, N2514, N1544);
and AND3 (N2518, N2500, N1703, N1885);
not NOT1 (N2519, N2511);
or OR4 (N2520, N2512, N1975, N2358, N2303);
and AND4 (N2521, N2515, N290, N2304, N1379);
not NOT1 (N2522, N2516);
nand NAND3 (N2523, N2519, N123, N41);
not NOT1 (N2524, N2522);
not NOT1 (N2525, N2504);
buf BUF1 (N2526, N2497);
nand NAND4 (N2527, N2520, N1976, N2073, N2065);
nor NOR4 (N2528, N2524, N1621, N1122, N1857);
xor XOR2 (N2529, N2513, N1400);
nand NAND3 (N2530, N2527, N35, N2421);
and AND4 (N2531, N2529, N1354, N232, N2239);
not NOT1 (N2532, N2517);
nand NAND2 (N2533, N2532, N1351);
not NOT1 (N2534, N2523);
nor NOR3 (N2535, N2526, N1186, N273);
and AND4 (N2536, N2533, N551, N1928, N1963);
or OR2 (N2537, N2534, N2279);
or OR4 (N2538, N2525, N2392, N1119, N764);
nand NAND3 (N2539, N2528, N1929, N1283);
and AND3 (N2540, N2521, N1745, N883);
buf BUF1 (N2541, N2510);
or OR4 (N2542, N2541, N1800, N1140, N870);
buf BUF1 (N2543, N2542);
or OR3 (N2544, N2530, N2071, N1860);
or OR2 (N2545, N2537, N1875);
nand NAND3 (N2546, N2540, N1242, N759);
or OR3 (N2547, N2539, N1451, N1687);
not NOT1 (N2548, N2531);
nand NAND2 (N2549, N2544, N1722);
buf BUF1 (N2550, N2535);
buf BUF1 (N2551, N2548);
not NOT1 (N2552, N2551);
nand NAND2 (N2553, N2538, N1782);
or OR3 (N2554, N2543, N1483, N764);
and AND4 (N2555, N2550, N74, N1514, N1150);
buf BUF1 (N2556, N2547);
nand NAND3 (N2557, N2556, N1193, N1927);
or OR4 (N2558, N2552, N797, N774, N2113);
xor XOR2 (N2559, N2546, N1300);
xor XOR2 (N2560, N2545, N2307);
buf BUF1 (N2561, N2549);
xor XOR2 (N2562, N2518, N2379);
nand NAND3 (N2563, N2553, N198, N2150);
not NOT1 (N2564, N2536);
buf BUF1 (N2565, N2564);
nand NAND2 (N2566, N2560, N851);
xor XOR2 (N2567, N2566, N2395);
xor XOR2 (N2568, N2554, N2192);
xor XOR2 (N2569, N2567, N497);
xor XOR2 (N2570, N2559, N755);
and AND3 (N2571, N2561, N64, N1501);
xor XOR2 (N2572, N2565, N1858);
nand NAND2 (N2573, N2572, N1268);
not NOT1 (N2574, N2562);
nand NAND2 (N2575, N2558, N1049);
buf BUF1 (N2576, N2573);
nor NOR3 (N2577, N2571, N2006, N1693);
not NOT1 (N2578, N2574);
buf BUF1 (N2579, N2575);
and AND3 (N2580, N2569, N1369, N1896);
nor NOR4 (N2581, N2555, N425, N2195, N1540);
or OR4 (N2582, N2579, N301, N1894, N1520);
xor XOR2 (N2583, N2557, N1307);
and AND3 (N2584, N2577, N2041, N2156);
not NOT1 (N2585, N2582);
or OR2 (N2586, N2563, N1386);
xor XOR2 (N2587, N2583, N704);
and AND4 (N2588, N2585, N2351, N130, N74);
and AND2 (N2589, N2581, N1527);
and AND3 (N2590, N2586, N407, N971);
and AND2 (N2591, N2578, N821);
and AND4 (N2592, N2570, N1793, N283, N2282);
xor XOR2 (N2593, N2592, N339);
buf BUF1 (N2594, N2588);
nor NOR2 (N2595, N2580, N113);
nand NAND2 (N2596, N2595, N2503);
buf BUF1 (N2597, N2584);
xor XOR2 (N2598, N2596, N1404);
nand NAND4 (N2599, N2593, N2359, N1288, N2126);
xor XOR2 (N2600, N2589, N2074);
buf BUF1 (N2601, N2568);
xor XOR2 (N2602, N2591, N1880);
and AND2 (N2603, N2601, N2188);
and AND4 (N2604, N2590, N228, N593, N1827);
nor NOR2 (N2605, N2604, N1858);
nand NAND3 (N2606, N2600, N2190, N1169);
or OR3 (N2607, N2598, N811, N1939);
xor XOR2 (N2608, N2606, N1502);
nand NAND3 (N2609, N2603, N831, N45);
nand NAND2 (N2610, N2605, N2270);
not NOT1 (N2611, N2597);
buf BUF1 (N2612, N2594);
xor XOR2 (N2613, N2608, N2064);
not NOT1 (N2614, N2610);
xor XOR2 (N2615, N2599, N33);
or OR4 (N2616, N2587, N323, N679, N614);
not NOT1 (N2617, N2612);
nor NOR3 (N2618, N2609, N729, N2257);
and AND2 (N2619, N2602, N496);
nor NOR3 (N2620, N2616, N4, N1222);
nand NAND3 (N2621, N2615, N1820, N2392);
or OR2 (N2622, N2576, N504);
nor NOR2 (N2623, N2618, N491);
and AND2 (N2624, N2623, N854);
not NOT1 (N2625, N2607);
and AND4 (N2626, N2614, N2607, N1421, N1083);
or OR4 (N2627, N2620, N879, N1450, N1044);
not NOT1 (N2628, N2622);
buf BUF1 (N2629, N2611);
and AND4 (N2630, N2625, N1773, N636, N1683);
or OR2 (N2631, N2629, N203);
nor NOR4 (N2632, N2613, N1041, N410, N2513);
not NOT1 (N2633, N2619);
nor NOR4 (N2634, N2624, N1067, N1452, N2076);
buf BUF1 (N2635, N2631);
not NOT1 (N2636, N2634);
or OR3 (N2637, N2626, N791, N1317);
not NOT1 (N2638, N2621);
or OR4 (N2639, N2630, N2435, N652, N398);
buf BUF1 (N2640, N2627);
or OR3 (N2641, N2637, N2352, N1915);
buf BUF1 (N2642, N2639);
xor XOR2 (N2643, N2617, N2006);
nand NAND3 (N2644, N2636, N575, N200);
or OR2 (N2645, N2642, N1221);
or OR2 (N2646, N2632, N446);
not NOT1 (N2647, N2640);
buf BUF1 (N2648, N2641);
nand NAND3 (N2649, N2635, N671, N238);
not NOT1 (N2650, N2638);
or OR2 (N2651, N2645, N1618);
xor XOR2 (N2652, N2650, N2031);
not NOT1 (N2653, N2648);
xor XOR2 (N2654, N2628, N2126);
nand NAND3 (N2655, N2646, N2532, N656);
not NOT1 (N2656, N2644);
xor XOR2 (N2657, N2656, N709);
nor NOR2 (N2658, N2651, N1416);
buf BUF1 (N2659, N2643);
or OR4 (N2660, N2655, N585, N1085, N1368);
nand NAND4 (N2661, N2658, N93, N1407, N2389);
nand NAND4 (N2662, N2660, N271, N1920, N1150);
buf BUF1 (N2663, N2647);
nor NOR3 (N2664, N2633, N328, N1458);
nor NOR4 (N2665, N2662, N1831, N1468, N2042);
nand NAND2 (N2666, N2649, N2043);
and AND2 (N2667, N2654, N52);
not NOT1 (N2668, N2653);
nor NOR4 (N2669, N2657, N2632, N1479, N2334);
xor XOR2 (N2670, N2667, N672);
nor NOR4 (N2671, N2659, N660, N2341, N172);
or OR2 (N2672, N2664, N592);
not NOT1 (N2673, N2670);
buf BUF1 (N2674, N2673);
nand NAND4 (N2675, N2661, N83, N1540, N1200);
not NOT1 (N2676, N2671);
and AND4 (N2677, N2666, N99, N1293, N2414);
not NOT1 (N2678, N2665);
xor XOR2 (N2679, N2677, N2417);
nor NOR3 (N2680, N2669, N1805, N2515);
and AND3 (N2681, N2675, N1925, N2038);
nand NAND3 (N2682, N2674, N577, N1931);
and AND2 (N2683, N2676, N856);
and AND3 (N2684, N2668, N856, N897);
or OR4 (N2685, N2682, N373, N1828, N1782);
and AND4 (N2686, N2678, N916, N231, N1741);
or OR4 (N2687, N2686, N1434, N519, N1733);
xor XOR2 (N2688, N2684, N550);
nand NAND3 (N2689, N2687, N1760, N1195);
not NOT1 (N2690, N2672);
xor XOR2 (N2691, N2680, N1564);
xor XOR2 (N2692, N2691, N1086);
nand NAND4 (N2693, N2689, N1627, N1139, N392);
or OR3 (N2694, N2663, N1089, N1796);
buf BUF1 (N2695, N2681);
and AND2 (N2696, N2694, N537);
xor XOR2 (N2697, N2679, N1269);
and AND2 (N2698, N2693, N2122);
or OR4 (N2699, N2688, N1380, N2661, N903);
and AND3 (N2700, N2683, N2030, N2629);
not NOT1 (N2701, N2698);
or OR2 (N2702, N2690, N73);
and AND3 (N2703, N2692, N1222, N1704);
not NOT1 (N2704, N2685);
not NOT1 (N2705, N2703);
or OR3 (N2706, N2700, N1117, N2159);
nand NAND3 (N2707, N2652, N1315, N1573);
and AND2 (N2708, N2697, N1344);
buf BUF1 (N2709, N2699);
or OR2 (N2710, N2704, N1656);
and AND4 (N2711, N2695, N1930, N2661, N200);
nand NAND4 (N2712, N2709, N308, N837, N1263);
or OR3 (N2713, N2707, N122, N1705);
xor XOR2 (N2714, N2696, N148);
nor NOR3 (N2715, N2714, N2089, N620);
and AND2 (N2716, N2712, N1686);
not NOT1 (N2717, N2705);
nand NAND4 (N2718, N2706, N2004, N1558, N377);
buf BUF1 (N2719, N2718);
xor XOR2 (N2720, N2711, N642);
nor NOR3 (N2721, N2715, N1934, N388);
nor NOR4 (N2722, N2721, N787, N610, N1180);
and AND4 (N2723, N2716, N2340, N1537, N693);
nor NOR3 (N2724, N2719, N1430, N2543);
xor XOR2 (N2725, N2724, N924);
xor XOR2 (N2726, N2702, N1676);
and AND2 (N2727, N2710, N146);
and AND4 (N2728, N2722, N344, N1255, N2625);
xor XOR2 (N2729, N2701, N678);
nor NOR4 (N2730, N2723, N1369, N2160, N1780);
nor NOR2 (N2731, N2728, N1361);
or OR2 (N2732, N2727, N2286);
not NOT1 (N2733, N2725);
nand NAND2 (N2734, N2726, N1627);
not NOT1 (N2735, N2731);
nor NOR2 (N2736, N2730, N1380);
and AND2 (N2737, N2717, N3);
buf BUF1 (N2738, N2734);
nor NOR3 (N2739, N2713, N1557, N1492);
or OR3 (N2740, N2733, N488, N2530);
nand NAND3 (N2741, N2737, N2364, N1530);
not NOT1 (N2742, N2739);
xor XOR2 (N2743, N2729, N2062);
not NOT1 (N2744, N2742);
and AND3 (N2745, N2735, N858, N1206);
xor XOR2 (N2746, N2744, N128);
buf BUF1 (N2747, N2746);
nor NOR4 (N2748, N2732, N1884, N1662, N2052);
and AND2 (N2749, N2741, N2632);
nor NOR4 (N2750, N2743, N2328, N2086, N1885);
and AND4 (N2751, N2738, N357, N2567, N651);
or OR4 (N2752, N2748, N66, N618, N326);
and AND4 (N2753, N2752, N54, N2444, N160);
and AND2 (N2754, N2747, N1855);
not NOT1 (N2755, N2708);
xor XOR2 (N2756, N2751, N1277);
and AND3 (N2757, N2736, N2258, N1902);
nor NOR2 (N2758, N2749, N2420);
not NOT1 (N2759, N2745);
buf BUF1 (N2760, N2720);
or OR2 (N2761, N2753, N948);
and AND3 (N2762, N2759, N475, N1443);
buf BUF1 (N2763, N2754);
buf BUF1 (N2764, N2762);
not NOT1 (N2765, N2758);
xor XOR2 (N2766, N2764, N1835);
and AND3 (N2767, N2750, N498, N2678);
not NOT1 (N2768, N2763);
or OR3 (N2769, N2767, N2094, N2187);
buf BUF1 (N2770, N2740);
nand NAND4 (N2771, N2766, N1418, N1092, N1465);
nor NOR3 (N2772, N2771, N1969, N2077);
buf BUF1 (N2773, N2761);
xor XOR2 (N2774, N2773, N2722);
xor XOR2 (N2775, N2760, N70);
not NOT1 (N2776, N2774);
nor NOR2 (N2777, N2756, N765);
buf BUF1 (N2778, N2770);
or OR4 (N2779, N2775, N2700, N1013, N2184);
not NOT1 (N2780, N2765);
and AND4 (N2781, N2772, N643, N129, N917);
or OR2 (N2782, N2768, N960);
or OR3 (N2783, N2780, N1640, N2593);
nand NAND4 (N2784, N2778, N912, N55, N134);
not NOT1 (N2785, N2776);
xor XOR2 (N2786, N2782, N1023);
nand NAND4 (N2787, N2769, N1798, N1483, N2282);
buf BUF1 (N2788, N2757);
xor XOR2 (N2789, N2788, N1951);
buf BUF1 (N2790, N2755);
xor XOR2 (N2791, N2785, N2380);
xor XOR2 (N2792, N2784, N769);
buf BUF1 (N2793, N2781);
buf BUF1 (N2794, N2786);
not NOT1 (N2795, N2792);
xor XOR2 (N2796, N2783, N2434);
buf BUF1 (N2797, N2793);
xor XOR2 (N2798, N2791, N1382);
nor NOR2 (N2799, N2790, N1048);
nand NAND4 (N2800, N2795, N2176, N2221, N196);
not NOT1 (N2801, N2798);
nand NAND4 (N2802, N2789, N2410, N632, N2017);
xor XOR2 (N2803, N2802, N1908);
buf BUF1 (N2804, N2787);
and AND2 (N2805, N2803, N982);
and AND3 (N2806, N2779, N1223, N752);
buf BUF1 (N2807, N2797);
or OR3 (N2808, N2800, N2477, N957);
buf BUF1 (N2809, N2796);
nor NOR3 (N2810, N2805, N805, N1276);
buf BUF1 (N2811, N2801);
and AND3 (N2812, N2799, N1428, N2240);
not NOT1 (N2813, N2810);
xor XOR2 (N2814, N2812, N704);
nor NOR4 (N2815, N2807, N1495, N2743, N1835);
and AND3 (N2816, N2815, N886, N1201);
xor XOR2 (N2817, N2806, N154);
nand NAND3 (N2818, N2817, N1627, N2807);
not NOT1 (N2819, N2814);
nand NAND3 (N2820, N2816, N1112, N1399);
nand NAND4 (N2821, N2820, N1475, N1095, N148);
nor NOR4 (N2822, N2819, N1307, N171, N2720);
xor XOR2 (N2823, N2809, N1027);
not NOT1 (N2824, N2818);
not NOT1 (N2825, N2824);
and AND2 (N2826, N2822, N97);
not NOT1 (N2827, N2813);
and AND2 (N2828, N2825, N1903);
and AND3 (N2829, N2794, N1647, N2589);
and AND4 (N2830, N2804, N879, N379, N1482);
xor XOR2 (N2831, N2777, N856);
nand NAND2 (N2832, N2811, N239);
xor XOR2 (N2833, N2832, N1789);
nand NAND4 (N2834, N2833, N156, N2275, N2672);
not NOT1 (N2835, N2830);
xor XOR2 (N2836, N2827, N616);
not NOT1 (N2837, N2823);
and AND4 (N2838, N2836, N1779, N567, N2152);
and AND3 (N2839, N2837, N443, N1347);
or OR3 (N2840, N2839, N2193, N89);
and AND3 (N2841, N2834, N580, N393);
and AND3 (N2842, N2840, N1352, N2561);
xor XOR2 (N2843, N2835, N1908);
buf BUF1 (N2844, N2828);
nor NOR3 (N2845, N2826, N2273, N2760);
and AND2 (N2846, N2838, N2543);
xor XOR2 (N2847, N2831, N1074);
or OR2 (N2848, N2844, N2005);
not NOT1 (N2849, N2847);
not NOT1 (N2850, N2849);
nand NAND3 (N2851, N2848, N156, N1846);
and AND4 (N2852, N2845, N20, N1304, N141);
buf BUF1 (N2853, N2821);
not NOT1 (N2854, N2852);
buf BUF1 (N2855, N2851);
and AND2 (N2856, N2842, N1917);
or OR2 (N2857, N2853, N1145);
and AND2 (N2858, N2850, N2504);
nand NAND2 (N2859, N2855, N2262);
nand NAND4 (N2860, N2859, N1387, N2425, N377);
or OR4 (N2861, N2854, N778, N1622, N797);
and AND3 (N2862, N2858, N2550, N1796);
or OR2 (N2863, N2843, N448);
buf BUF1 (N2864, N2841);
and AND3 (N2865, N2864, N448, N2049);
and AND3 (N2866, N2865, N1261, N2820);
not NOT1 (N2867, N2866);
not NOT1 (N2868, N2863);
and AND4 (N2869, N2861, N1415, N593, N172);
xor XOR2 (N2870, N2808, N827);
not NOT1 (N2871, N2857);
nand NAND4 (N2872, N2846, N599, N631, N1746);
nor NOR3 (N2873, N2868, N271, N1936);
or OR3 (N2874, N2856, N656, N841);
nand NAND2 (N2875, N2860, N1191);
or OR4 (N2876, N2873, N1179, N1533, N1845);
not NOT1 (N2877, N2871);
nor NOR4 (N2878, N2862, N141, N1306, N1057);
nor NOR3 (N2879, N2878, N1458, N2455);
nor NOR2 (N2880, N2872, N759);
not NOT1 (N2881, N2880);
xor XOR2 (N2882, N2877, N1667);
not NOT1 (N2883, N2881);
buf BUF1 (N2884, N2867);
and AND4 (N2885, N2870, N668, N2080, N668);
nor NOR4 (N2886, N2884, N2188, N1990, N2804);
buf BUF1 (N2887, N2882);
not NOT1 (N2888, N2886);
not NOT1 (N2889, N2869);
nor NOR2 (N2890, N2875, N2331);
nor NOR4 (N2891, N2887, N2427, N2029, N185);
nor NOR2 (N2892, N2829, N1366);
not NOT1 (N2893, N2883);
xor XOR2 (N2894, N2876, N627);
xor XOR2 (N2895, N2891, N1137);
or OR4 (N2896, N2895, N2639, N1615, N1379);
nor NOR3 (N2897, N2874, N1150, N2496);
nand NAND3 (N2898, N2889, N1097, N2764);
not NOT1 (N2899, N2897);
and AND4 (N2900, N2899, N1983, N2118, N1538);
or OR2 (N2901, N2892, N2591);
or OR3 (N2902, N2894, N191, N1758);
xor XOR2 (N2903, N2890, N471);
nand NAND2 (N2904, N2888, N1586);
nand NAND4 (N2905, N2901, N2563, N2381, N863);
or OR2 (N2906, N2896, N992);
nor NOR4 (N2907, N2903, N2185, N2625, N1713);
or OR2 (N2908, N2905, N2762);
xor XOR2 (N2909, N2908, N530);
buf BUF1 (N2910, N2907);
or OR2 (N2911, N2893, N2419);
nor NOR2 (N2912, N2879, N1165);
or OR2 (N2913, N2911, N897);
xor XOR2 (N2914, N2885, N1842);
and AND3 (N2915, N2898, N2695, N2842);
nand NAND2 (N2916, N2914, N2712);
nand NAND4 (N2917, N2904, N2587, N624, N2531);
nand NAND2 (N2918, N2917, N2429);
nand NAND2 (N2919, N2918, N200);
not NOT1 (N2920, N2906);
buf BUF1 (N2921, N2900);
xor XOR2 (N2922, N2921, N332);
buf BUF1 (N2923, N2909);
buf BUF1 (N2924, N2912);
nand NAND2 (N2925, N2913, N2166);
or OR2 (N2926, N2924, N502);
not NOT1 (N2927, N2926);
and AND4 (N2928, N2910, N2610, N1792, N1425);
not NOT1 (N2929, N2922);
and AND3 (N2930, N2929, N1204, N2519);
nor NOR2 (N2931, N2928, N834);
not NOT1 (N2932, N2920);
and AND4 (N2933, N2930, N788, N1282, N1942);
and AND4 (N2934, N2925, N1957, N2295, N2667);
and AND2 (N2935, N2923, N1302);
or OR2 (N2936, N2934, N2638);
or OR4 (N2937, N2932, N165, N1743, N2661);
or OR4 (N2938, N2936, N678, N1021, N2604);
not NOT1 (N2939, N2919);
nand NAND4 (N2940, N2939, N1644, N143, N1740);
xor XOR2 (N2941, N2940, N1519);
or OR3 (N2942, N2933, N2835, N2635);
not NOT1 (N2943, N2935);
not NOT1 (N2944, N2927);
not NOT1 (N2945, N2902);
nand NAND3 (N2946, N2931, N465, N26);
and AND3 (N2947, N2941, N233, N428);
not NOT1 (N2948, N2916);
nand NAND2 (N2949, N2938, N2502);
buf BUF1 (N2950, N2949);
nor NOR4 (N2951, N2942, N585, N72, N759);
nor NOR4 (N2952, N2951, N1226, N806, N2524);
not NOT1 (N2953, N2948);
not NOT1 (N2954, N2937);
not NOT1 (N2955, N2945);
nand NAND2 (N2956, N2952, N1371);
not NOT1 (N2957, N2954);
nand NAND4 (N2958, N2944, N1190, N657, N1864);
buf BUF1 (N2959, N2956);
or OR4 (N2960, N2953, N2563, N2118, N47);
nand NAND4 (N2961, N2915, N820, N2168, N2813);
nor NOR4 (N2962, N2947, N199, N1743, N314);
or OR3 (N2963, N2961, N1287, N1082);
or OR3 (N2964, N2946, N703, N2110);
buf BUF1 (N2965, N2963);
buf BUF1 (N2966, N2962);
buf BUF1 (N2967, N2965);
buf BUF1 (N2968, N2964);
and AND4 (N2969, N2958, N831, N1630, N405);
and AND2 (N2970, N2957, N1605);
nand NAND4 (N2971, N2959, N1593, N2400, N1067);
not NOT1 (N2972, N2950);
buf BUF1 (N2973, N2972);
not NOT1 (N2974, N2969);
and AND4 (N2975, N2955, N372, N2941, N96);
buf BUF1 (N2976, N2975);
nand NAND4 (N2977, N2971, N188, N892, N1025);
buf BUF1 (N2978, N2977);
nor NOR3 (N2979, N2976, N2388, N665);
not NOT1 (N2980, N2943);
and AND2 (N2981, N2978, N1538);
not NOT1 (N2982, N2974);
xor XOR2 (N2983, N2966, N614);
buf BUF1 (N2984, N2979);
buf BUF1 (N2985, N2967);
nand NAND3 (N2986, N2980, N576, N2214);
xor XOR2 (N2987, N2981, N2869);
not NOT1 (N2988, N2985);
not NOT1 (N2989, N2968);
nand NAND4 (N2990, N2984, N290, N2771, N1219);
nand NAND2 (N2991, N2986, N984);
and AND3 (N2992, N2989, N2485, N2446);
not NOT1 (N2993, N2991);
not NOT1 (N2994, N2992);
not NOT1 (N2995, N2987);
buf BUF1 (N2996, N2970);
buf BUF1 (N2997, N2995);
nand NAND3 (N2998, N2993, N1707, N1567);
nor NOR3 (N2999, N2960, N2734, N1610);
and AND3 (N3000, N2999, N703, N1449);
not NOT1 (N3001, N2982);
or OR4 (N3002, N2988, N692, N535, N246);
nand NAND3 (N3003, N2983, N385, N941);
not NOT1 (N3004, N2997);
xor XOR2 (N3005, N2998, N2269);
and AND4 (N3006, N3002, N183, N132, N1218);
xor XOR2 (N3007, N3000, N1154);
buf BUF1 (N3008, N3004);
not NOT1 (N3009, N3007);
or OR3 (N3010, N3001, N939, N1188);
nand NAND2 (N3011, N3010, N2943);
nand NAND3 (N3012, N3008, N1871, N2055);
not NOT1 (N3013, N3009);
and AND4 (N3014, N3011, N1133, N2630, N2980);
nor NOR3 (N3015, N3012, N2405, N2270);
and AND3 (N3016, N3013, N2188, N1495);
buf BUF1 (N3017, N2973);
or OR4 (N3018, N2990, N1511, N2130, N965);
nor NOR3 (N3019, N2996, N2343, N2661);
nand NAND3 (N3020, N3006, N835, N1567);
not NOT1 (N3021, N3005);
or OR2 (N3022, N3014, N1799);
or OR3 (N3023, N3019, N2957, N265);
xor XOR2 (N3024, N3003, N292);
and AND3 (N3025, N3023, N1147, N440);
and AND2 (N3026, N3025, N938);
nor NOR2 (N3027, N3015, N116);
nor NOR4 (N3028, N2994, N1165, N1558, N1430);
buf BUF1 (N3029, N3026);
xor XOR2 (N3030, N3022, N2368);
and AND4 (N3031, N3017, N491, N2773, N2582);
nor NOR4 (N3032, N3031, N642, N1709, N1346);
not NOT1 (N3033, N3020);
and AND2 (N3034, N3032, N1718);
nand NAND4 (N3035, N3033, N738, N1150, N539);
or OR4 (N3036, N3034, N1643, N583, N158);
xor XOR2 (N3037, N3036, N83);
or OR4 (N3038, N3037, N2173, N1371, N911);
buf BUF1 (N3039, N3018);
xor XOR2 (N3040, N3016, N1916);
nor NOR4 (N3041, N3030, N1416, N1040, N1729);
buf BUF1 (N3042, N3024);
and AND4 (N3043, N3027, N2932, N104, N43);
nand NAND3 (N3044, N3038, N2658, N2171);
and AND3 (N3045, N3028, N2938, N3036);
and AND4 (N3046, N3042, N355, N2610, N1297);
not NOT1 (N3047, N3046);
xor XOR2 (N3048, N3045, N1562);
and AND3 (N3049, N3040, N1770, N533);
not NOT1 (N3050, N3029);
xor XOR2 (N3051, N3021, N1136);
xor XOR2 (N3052, N3035, N2535);
nand NAND4 (N3053, N3050, N1200, N858, N2995);
nand NAND4 (N3054, N3043, N2553, N825, N1231);
or OR2 (N3055, N3047, N1765);
nor NOR4 (N3056, N3039, N95, N2574, N701);
nor NOR3 (N3057, N3041, N1838, N1790);
nand NAND2 (N3058, N3051, N2143);
xor XOR2 (N3059, N3055, N2706);
buf BUF1 (N3060, N3059);
nand NAND2 (N3061, N3044, N2275);
xor XOR2 (N3062, N3052, N860);
or OR4 (N3063, N3049, N1945, N2794, N779);
and AND3 (N3064, N3062, N1114, N996);
xor XOR2 (N3065, N3053, N2395);
not NOT1 (N3066, N3058);
nand NAND2 (N3067, N3057, N1213);
buf BUF1 (N3068, N3060);
nand NAND3 (N3069, N3067, N2192, N2435);
nor NOR4 (N3070, N3061, N1373, N2337, N618);
nor NOR4 (N3071, N3065, N2166, N506, N151);
or OR3 (N3072, N3070, N505, N1810);
buf BUF1 (N3073, N3071);
buf BUF1 (N3074, N3064);
nand NAND2 (N3075, N3069, N1029);
nor NOR4 (N3076, N3056, N226, N686, N2336);
buf BUF1 (N3077, N3063);
nor NOR3 (N3078, N3076, N2806, N1182);
buf BUF1 (N3079, N3048);
buf BUF1 (N3080, N3075);
or OR4 (N3081, N3080, N104, N1687, N1435);
xor XOR2 (N3082, N3081, N1967);
not NOT1 (N3083, N3079);
nor NOR2 (N3084, N3082, N2047);
nor NOR2 (N3085, N3077, N1502);
nand NAND3 (N3086, N3066, N2844, N790);
or OR2 (N3087, N3085, N55);
xor XOR2 (N3088, N3072, N643);
not NOT1 (N3089, N3073);
and AND2 (N3090, N3088, N2139);
or OR4 (N3091, N3090, N2082, N136, N159);
xor XOR2 (N3092, N3054, N2112);
buf BUF1 (N3093, N3086);
and AND2 (N3094, N3091, N1914);
nor NOR3 (N3095, N3092, N2700, N2782);
nor NOR2 (N3096, N3078, N1588);
xor XOR2 (N3097, N3096, N133);
xor XOR2 (N3098, N3083, N1708);
or OR2 (N3099, N3068, N138);
nor NOR4 (N3100, N3094, N2611, N2868, N1427);
buf BUF1 (N3101, N3074);
nor NOR2 (N3102, N3089, N2867);
nor NOR4 (N3103, N3102, N1352, N1339, N581);
not NOT1 (N3104, N3101);
buf BUF1 (N3105, N3100);
nor NOR4 (N3106, N3105, N1377, N221, N888);
and AND4 (N3107, N3098, N1877, N455, N2478);
nand NAND4 (N3108, N3107, N864, N1844, N1789);
not NOT1 (N3109, N3087);
buf BUF1 (N3110, N3097);
or OR4 (N3111, N3104, N1363, N1941, N1296);
or OR3 (N3112, N3103, N1553, N2450);
nor NOR3 (N3113, N3093, N1201, N1904);
xor XOR2 (N3114, N3110, N2643);
buf BUF1 (N3115, N3114);
nor NOR3 (N3116, N3115, N272, N2851);
nand NAND4 (N3117, N3099, N1316, N1353, N2821);
xor XOR2 (N3118, N3084, N2209);
or OR2 (N3119, N3112, N117);
buf BUF1 (N3120, N3109);
and AND2 (N3121, N3113, N1813);
and AND3 (N3122, N3119, N754, N2925);
not NOT1 (N3123, N3108);
or OR3 (N3124, N3111, N2016, N1285);
nand NAND4 (N3125, N3122, N2035, N1147, N2075);
buf BUF1 (N3126, N3124);
nand NAND2 (N3127, N3095, N1951);
and AND3 (N3128, N3126, N1399, N1233);
buf BUF1 (N3129, N3120);
or OR2 (N3130, N3125, N3078);
nand NAND4 (N3131, N3116, N286, N2912, N154);
and AND4 (N3132, N3130, N1878, N2199, N1815);
not NOT1 (N3133, N3121);
buf BUF1 (N3134, N3132);
nor NOR2 (N3135, N3133, N1230);
buf BUF1 (N3136, N3127);
buf BUF1 (N3137, N3106);
and AND3 (N3138, N3129, N230, N764);
nand NAND4 (N3139, N3117, N2459, N2223, N1863);
buf BUF1 (N3140, N3137);
and AND2 (N3141, N3140, N2344);
nand NAND4 (N3142, N3131, N452, N1079, N713);
or OR2 (N3143, N3142, N1246);
or OR2 (N3144, N3134, N1470);
nor NOR2 (N3145, N3118, N1296);
buf BUF1 (N3146, N3123);
xor XOR2 (N3147, N3138, N675);
not NOT1 (N3148, N3141);
or OR2 (N3149, N3147, N1499);
nand NAND3 (N3150, N3145, N1577, N2523);
and AND2 (N3151, N3128, N132);
and AND2 (N3152, N3146, N2692);
nor NOR4 (N3153, N3139, N1618, N2404, N2682);
or OR4 (N3154, N3150, N843, N2683, N895);
and AND3 (N3155, N3143, N2641, N1827);
xor XOR2 (N3156, N3144, N2134);
or OR3 (N3157, N3136, N1154, N1620);
nor NOR2 (N3158, N3151, N625);
nand NAND4 (N3159, N3148, N573, N1333, N139);
xor XOR2 (N3160, N3135, N1509);
xor XOR2 (N3161, N3156, N2634);
buf BUF1 (N3162, N3161);
or OR3 (N3163, N3153, N983, N2724);
not NOT1 (N3164, N3162);
not NOT1 (N3165, N3158);
buf BUF1 (N3166, N3160);
not NOT1 (N3167, N3157);
not NOT1 (N3168, N3159);
nor NOR4 (N3169, N3152, N2674, N1794, N1868);
nand NAND4 (N3170, N3154, N2472, N2312, N883);
and AND3 (N3171, N3165, N58, N1402);
nor NOR3 (N3172, N3163, N1923, N1748);
or OR2 (N3173, N3155, N300);
nand NAND4 (N3174, N3164, N2359, N2887, N2959);
or OR4 (N3175, N3174, N2556, N35, N273);
and AND2 (N3176, N3173, N1046);
and AND2 (N3177, N3149, N2882);
not NOT1 (N3178, N3169);
or OR3 (N3179, N3176, N147, N183);
and AND3 (N3180, N3171, N907, N1934);
nand NAND3 (N3181, N3179, N2973, N3040);
xor XOR2 (N3182, N3168, N1380);
and AND4 (N3183, N3178, N2520, N2994, N2183);
or OR4 (N3184, N3180, N2612, N548, N1871);
xor XOR2 (N3185, N3181, N791);
or OR4 (N3186, N3172, N1379, N3131, N291);
or OR4 (N3187, N3184, N1456, N3153, N2627);
and AND3 (N3188, N3177, N860, N218);
and AND4 (N3189, N3166, N1291, N1813, N2732);
nor NOR2 (N3190, N3170, N1992);
xor XOR2 (N3191, N3183, N1329);
buf BUF1 (N3192, N3175);
xor XOR2 (N3193, N3192, N31);
or OR3 (N3194, N3167, N443, N1562);
or OR3 (N3195, N3194, N1645, N958);
not NOT1 (N3196, N3187);
buf BUF1 (N3197, N3196);
xor XOR2 (N3198, N3182, N420);
nor NOR4 (N3199, N3185, N820, N2746, N1820);
not NOT1 (N3200, N3198);
or OR3 (N3201, N3189, N2137, N2525);
nand NAND3 (N3202, N3199, N1583, N192);
and AND4 (N3203, N3195, N2072, N3148, N2799);
nor NOR3 (N3204, N3190, N1271, N3087);
nand NAND4 (N3205, N3200, N2645, N320, N1846);
xor XOR2 (N3206, N3191, N1506);
and AND2 (N3207, N3186, N2265);
buf BUF1 (N3208, N3193);
not NOT1 (N3209, N3208);
xor XOR2 (N3210, N3202, N1375);
or OR4 (N3211, N3188, N2955, N1176, N935);
nor NOR4 (N3212, N3203, N2648, N2931, N1299);
nor NOR4 (N3213, N3197, N2528, N2246, N2072);
buf BUF1 (N3214, N3211);
nor NOR4 (N3215, N3201, N1208, N3124, N2426);
xor XOR2 (N3216, N3210, N495);
endmodule