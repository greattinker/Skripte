// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17;

output N2008,N1993,N2010,N2000,N1998,N2007,N2014,N2009,N2012,N2017;

xor XOR2 (N18, N15, N2);
buf BUF1 (N19, N11);
or OR3 (N20, N17, N13, N15);
and AND2 (N21, N18, N3);
buf BUF1 (N22, N13);
or OR3 (N23, N10, N12, N13);
nor NOR2 (N24, N18, N7);
buf BUF1 (N25, N1);
xor XOR2 (N26, N19, N24);
not NOT1 (N27, N16);
not NOT1 (N28, N16);
not NOT1 (N29, N6);
nand NAND4 (N30, N4, N27, N29, N16);
not NOT1 (N31, N1);
buf BUF1 (N32, N10);
nor NOR2 (N33, N30, N26);
nor NOR4 (N34, N25, N15, N19, N22);
or OR4 (N35, N22, N30, N32, N23);
nand NAND3 (N36, N29, N34, N12);
xor XOR2 (N37, N10, N30);
xor XOR2 (N38, N36, N23);
xor XOR2 (N39, N36, N12);
nor NOR3 (N40, N5, N11, N3);
or OR4 (N41, N31, N17, N10, N32);
and AND3 (N42, N20, N30, N1);
buf BUF1 (N43, N38);
buf BUF1 (N44, N40);
and AND4 (N45, N33, N39, N7, N7);
xor XOR2 (N46, N38, N38);
buf BUF1 (N47, N35);
or OR2 (N48, N41, N23);
buf BUF1 (N49, N48);
xor XOR2 (N50, N44, N1);
and AND3 (N51, N21, N35, N46);
or OR4 (N52, N6, N19, N15, N10);
or OR3 (N53, N49, N45, N29);
buf BUF1 (N54, N5);
xor XOR2 (N55, N28, N15);
not NOT1 (N56, N37);
nand NAND3 (N57, N55, N35, N38);
or OR3 (N58, N42, N1, N7);
xor XOR2 (N59, N51, N49);
nor NOR4 (N60, N53, N39, N26, N18);
not NOT1 (N61, N50);
not NOT1 (N62, N52);
buf BUF1 (N63, N56);
or OR2 (N64, N60, N7);
and AND4 (N65, N47, N43, N19, N62);
or OR4 (N66, N57, N13, N47, N19);
nand NAND4 (N67, N22, N5, N13, N32);
nand NAND3 (N68, N60, N51, N50);
nand NAND3 (N69, N68, N42, N20);
and AND2 (N70, N67, N36);
nand NAND2 (N71, N64, N17);
nor NOR3 (N72, N71, N56, N26);
xor XOR2 (N73, N63, N19);
nor NOR2 (N74, N66, N5);
nand NAND2 (N75, N59, N69);
nand NAND4 (N76, N42, N2, N46, N60);
or OR3 (N77, N58, N60, N17);
and AND2 (N78, N54, N17);
or OR2 (N79, N72, N57);
and AND2 (N80, N65, N62);
buf BUF1 (N81, N70);
and AND2 (N82, N73, N70);
and AND3 (N83, N82, N76, N30);
not NOT1 (N84, N79);
nand NAND3 (N85, N46, N14, N64);
nand NAND2 (N86, N85, N78);
nor NOR4 (N87, N46, N71, N17, N71);
nor NOR4 (N88, N84, N9, N34, N87);
or OR2 (N89, N56, N74);
nor NOR2 (N90, N8, N60);
or OR4 (N91, N83, N73, N77, N56);
or OR2 (N92, N40, N16);
or OR3 (N93, N88, N45, N58);
xor XOR2 (N94, N61, N9);
nand NAND2 (N95, N91, N22);
xor XOR2 (N96, N89, N92);
buf BUF1 (N97, N6);
nor NOR3 (N98, N94, N62, N91);
buf BUF1 (N99, N75);
and AND2 (N100, N86, N9);
or OR4 (N101, N80, N95, N62, N23);
and AND2 (N102, N19, N15);
xor XOR2 (N103, N93, N20);
nand NAND2 (N104, N102, N61);
not NOT1 (N105, N101);
nand NAND3 (N106, N96, N76, N100);
and AND3 (N107, N101, N74, N1);
nand NAND2 (N108, N103, N83);
buf BUF1 (N109, N99);
buf BUF1 (N110, N81);
buf BUF1 (N111, N97);
buf BUF1 (N112, N109);
not NOT1 (N113, N112);
nor NOR4 (N114, N105, N89, N32, N22);
nand NAND2 (N115, N98, N55);
or OR3 (N116, N115, N31, N76);
xor XOR2 (N117, N106, N4);
nor NOR3 (N118, N116, N14, N112);
or OR2 (N119, N113, N28);
or OR3 (N120, N107, N46, N37);
nor NOR2 (N121, N90, N51);
buf BUF1 (N122, N120);
not NOT1 (N123, N119);
and AND3 (N124, N104, N59, N118);
nor NOR3 (N125, N52, N118, N65);
nand NAND3 (N126, N123, N28, N77);
nand NAND2 (N127, N114, N85);
or OR4 (N128, N117, N123, N15, N125);
nand NAND4 (N129, N123, N85, N66, N80);
xor XOR2 (N130, N126, N90);
not NOT1 (N131, N124);
nor NOR2 (N132, N108, N4);
nor NOR2 (N133, N110, N77);
nor NOR2 (N134, N133, N104);
xor XOR2 (N135, N129, N87);
not NOT1 (N136, N111);
not NOT1 (N137, N132);
xor XOR2 (N138, N131, N124);
buf BUF1 (N139, N136);
xor XOR2 (N140, N137, N21);
and AND2 (N141, N128, N55);
nor NOR2 (N142, N140, N9);
buf BUF1 (N143, N134);
xor XOR2 (N144, N142, N112);
nor NOR4 (N145, N144, N97, N61, N65);
or OR3 (N146, N121, N69, N97);
not NOT1 (N147, N139);
xor XOR2 (N148, N146, N140);
and AND3 (N149, N130, N50, N38);
nor NOR4 (N150, N141, N30, N136, N101);
buf BUF1 (N151, N147);
nor NOR3 (N152, N150, N51, N80);
and AND4 (N153, N135, N5, N90, N120);
not NOT1 (N154, N145);
or OR4 (N155, N122, N140, N109, N63);
or OR3 (N156, N143, N65, N41);
and AND3 (N157, N151, N128, N13);
buf BUF1 (N158, N127);
and AND4 (N159, N154, N2, N119, N46);
nor NOR2 (N160, N153, N57);
not NOT1 (N161, N138);
buf BUF1 (N162, N155);
xor XOR2 (N163, N152, N134);
nor NOR2 (N164, N157, N136);
and AND3 (N165, N156, N71, N37);
nand NAND3 (N166, N158, N25, N72);
nand NAND4 (N167, N148, N112, N35, N64);
or OR3 (N168, N164, N155, N5);
and AND2 (N169, N166, N86);
xor XOR2 (N170, N165, N38);
not NOT1 (N171, N149);
buf BUF1 (N172, N160);
nor NOR2 (N173, N163, N150);
or OR2 (N174, N170, N119);
nor NOR3 (N175, N171, N123, N113);
and AND3 (N176, N172, N152, N170);
and AND4 (N177, N173, N143, N144, N117);
not NOT1 (N178, N167);
nand NAND3 (N179, N168, N120, N111);
and AND4 (N180, N179, N82, N154, N124);
xor XOR2 (N181, N178, N178);
and AND4 (N182, N159, N69, N77, N163);
not NOT1 (N183, N169);
or OR2 (N184, N177, N118);
xor XOR2 (N185, N176, N117);
and AND3 (N186, N162, N3, N13);
and AND3 (N187, N186, N9, N30);
nor NOR3 (N188, N184, N33, N21);
and AND4 (N189, N175, N156, N134, N182);
and AND4 (N190, N109, N85, N182, N134);
not NOT1 (N191, N180);
buf BUF1 (N192, N191);
buf BUF1 (N193, N190);
buf BUF1 (N194, N187);
or OR3 (N195, N161, N13, N81);
nand NAND3 (N196, N188, N182, N119);
not NOT1 (N197, N189);
not NOT1 (N198, N193);
or OR3 (N199, N174, N134, N43);
not NOT1 (N200, N183);
and AND4 (N201, N192, N194, N65, N144);
buf BUF1 (N202, N87);
buf BUF1 (N203, N196);
or OR2 (N204, N199, N190);
not NOT1 (N205, N201);
nand NAND3 (N206, N202, N92, N46);
nand NAND4 (N207, N198, N94, N68, N122);
not NOT1 (N208, N205);
nand NAND2 (N209, N207, N82);
xor XOR2 (N210, N204, N139);
buf BUF1 (N211, N208);
nor NOR3 (N212, N200, N144, N190);
not NOT1 (N213, N197);
nand NAND2 (N214, N210, N19);
nand NAND2 (N215, N211, N70);
not NOT1 (N216, N213);
nor NOR4 (N217, N203, N109, N35, N135);
or OR2 (N218, N209, N32);
buf BUF1 (N219, N185);
buf BUF1 (N220, N181);
or OR2 (N221, N217, N17);
or OR2 (N222, N218, N28);
or OR4 (N223, N214, N68, N200, N144);
or OR2 (N224, N219, N177);
or OR3 (N225, N220, N13, N11);
nor NOR4 (N226, N223, N29, N182, N170);
or OR4 (N227, N216, N122, N69, N163);
buf BUF1 (N228, N224);
or OR2 (N229, N228, N208);
or OR3 (N230, N212, N150, N154);
xor XOR2 (N231, N226, N56);
xor XOR2 (N232, N230, N131);
and AND4 (N233, N222, N220, N118, N88);
xor XOR2 (N234, N232, N179);
xor XOR2 (N235, N229, N4);
nand NAND3 (N236, N231, N127, N110);
buf BUF1 (N237, N235);
buf BUF1 (N238, N233);
nand NAND4 (N239, N215, N139, N217, N182);
nor NOR4 (N240, N237, N165, N120, N154);
not NOT1 (N241, N234);
or OR3 (N242, N241, N177, N19);
xor XOR2 (N243, N206, N124);
not NOT1 (N244, N239);
xor XOR2 (N245, N225, N12);
or OR3 (N246, N221, N131, N158);
nor NOR3 (N247, N240, N44, N131);
or OR2 (N248, N236, N49);
buf BUF1 (N249, N246);
and AND2 (N250, N195, N132);
not NOT1 (N251, N250);
nor NOR3 (N252, N245, N132, N97);
not NOT1 (N253, N242);
nor NOR4 (N254, N253, N29, N110, N217);
nor NOR4 (N255, N249, N57, N215, N104);
buf BUF1 (N256, N251);
buf BUF1 (N257, N238);
not NOT1 (N258, N244);
nor NOR3 (N259, N227, N217, N63);
xor XOR2 (N260, N248, N71);
nor NOR4 (N261, N254, N69, N165, N109);
nand NAND2 (N262, N247, N123);
nor NOR4 (N263, N261, N44, N48, N63);
not NOT1 (N264, N255);
or OR4 (N265, N259, N109, N162, N85);
not NOT1 (N266, N252);
nor NOR4 (N267, N243, N41, N197, N255);
or OR3 (N268, N256, N26, N63);
and AND2 (N269, N264, N239);
or OR3 (N270, N268, N194, N12);
or OR4 (N271, N260, N132, N36, N260);
or OR2 (N272, N270, N261);
not NOT1 (N273, N265);
and AND3 (N274, N257, N37, N267);
not NOT1 (N275, N184);
not NOT1 (N276, N274);
xor XOR2 (N277, N273, N79);
or OR4 (N278, N262, N142, N44, N245);
buf BUF1 (N279, N263);
xor XOR2 (N280, N269, N28);
not NOT1 (N281, N280);
or OR3 (N282, N277, N171, N114);
xor XOR2 (N283, N275, N186);
nand NAND2 (N284, N276, N221);
not NOT1 (N285, N272);
nor NOR2 (N286, N266, N178);
and AND2 (N287, N279, N124);
and AND4 (N288, N285, N216, N280, N8);
not NOT1 (N289, N258);
buf BUF1 (N290, N286);
not NOT1 (N291, N281);
xor XOR2 (N292, N289, N10);
nand NAND3 (N293, N284, N46, N225);
nand NAND4 (N294, N291, N179, N175, N74);
xor XOR2 (N295, N287, N227);
buf BUF1 (N296, N290);
not NOT1 (N297, N283);
nor NOR3 (N298, N295, N156, N152);
not NOT1 (N299, N296);
buf BUF1 (N300, N271);
and AND4 (N301, N297, N56, N239, N166);
buf BUF1 (N302, N282);
nand NAND2 (N303, N301, N191);
not NOT1 (N304, N293);
not NOT1 (N305, N292);
nor NOR4 (N306, N288, N145, N282, N219);
or OR3 (N307, N303, N176, N169);
nor NOR4 (N308, N305, N184, N206, N34);
not NOT1 (N309, N308);
nand NAND2 (N310, N304, N280);
or OR4 (N311, N300, N82, N104, N43);
nor NOR4 (N312, N311, N218, N294, N226);
xor XOR2 (N313, N309, N216);
buf BUF1 (N314, N162);
and AND3 (N315, N307, N253, N26);
nor NOR3 (N316, N312, N212, N50);
nand NAND4 (N317, N314, N34, N51, N275);
buf BUF1 (N318, N278);
and AND2 (N319, N302, N7);
buf BUF1 (N320, N298);
and AND2 (N321, N306, N182);
not NOT1 (N322, N321);
or OR4 (N323, N310, N72, N199, N35);
xor XOR2 (N324, N318, N293);
nor NOR3 (N325, N316, N166, N276);
not NOT1 (N326, N319);
xor XOR2 (N327, N315, N267);
not NOT1 (N328, N317);
or OR2 (N329, N313, N54);
buf BUF1 (N330, N327);
xor XOR2 (N331, N325, N200);
nand NAND3 (N332, N299, N9, N88);
or OR2 (N333, N326, N13);
and AND2 (N334, N331, N115);
buf BUF1 (N335, N330);
buf BUF1 (N336, N322);
nand NAND2 (N337, N323, N76);
nand NAND3 (N338, N328, N227, N198);
not NOT1 (N339, N320);
buf BUF1 (N340, N336);
and AND4 (N341, N329, N16, N214, N82);
xor XOR2 (N342, N341, N24);
not NOT1 (N343, N332);
nand NAND2 (N344, N340, N259);
not NOT1 (N345, N343);
or OR4 (N346, N338, N49, N67, N78);
or OR3 (N347, N342, N292, N164);
nor NOR3 (N348, N346, N51, N340);
nand NAND3 (N349, N337, N321, N114);
buf BUF1 (N350, N348);
buf BUF1 (N351, N333);
xor XOR2 (N352, N334, N3);
not NOT1 (N353, N324);
buf BUF1 (N354, N351);
or OR3 (N355, N335, N23, N90);
not NOT1 (N356, N355);
or OR3 (N357, N339, N345, N355);
xor XOR2 (N358, N217, N111);
or OR4 (N359, N344, N304, N55, N335);
xor XOR2 (N360, N347, N26);
not NOT1 (N361, N360);
nor NOR4 (N362, N353, N181, N328, N236);
buf BUF1 (N363, N354);
or OR2 (N364, N362, N6);
xor XOR2 (N365, N361, N228);
xor XOR2 (N366, N364, N187);
buf BUF1 (N367, N365);
or OR2 (N368, N356, N75);
and AND4 (N369, N366, N134, N253, N312);
xor XOR2 (N370, N352, N105);
xor XOR2 (N371, N367, N322);
or OR3 (N372, N357, N72, N177);
not NOT1 (N373, N363);
nor NOR3 (N374, N369, N60, N269);
not NOT1 (N375, N368);
or OR2 (N376, N350, N108);
buf BUF1 (N377, N371);
not NOT1 (N378, N377);
or OR3 (N379, N359, N115, N349);
and AND3 (N380, N188, N124, N6);
not NOT1 (N381, N373);
not NOT1 (N382, N374);
or OR4 (N383, N370, N75, N9, N358);
buf BUF1 (N384, N87);
nand NAND4 (N385, N378, N57, N139, N136);
xor XOR2 (N386, N380, N255);
nand NAND4 (N387, N381, N256, N227, N274);
and AND3 (N388, N376, N99, N196);
and AND3 (N389, N372, N68, N229);
nor NOR4 (N390, N384, N76, N32, N246);
nor NOR2 (N391, N382, N332);
nor NOR3 (N392, N391, N245, N183);
nand NAND2 (N393, N375, N86);
nand NAND4 (N394, N388, N195, N307, N362);
and AND2 (N395, N394, N188);
and AND2 (N396, N383, N274);
not NOT1 (N397, N389);
nor NOR4 (N398, N386, N360, N299, N242);
or OR2 (N399, N385, N303);
not NOT1 (N400, N387);
nor NOR2 (N401, N393, N234);
buf BUF1 (N402, N390);
xor XOR2 (N403, N395, N266);
not NOT1 (N404, N397);
not NOT1 (N405, N402);
not NOT1 (N406, N405);
xor XOR2 (N407, N406, N6);
or OR2 (N408, N398, N181);
buf BUF1 (N409, N404);
or OR2 (N410, N409, N389);
and AND2 (N411, N401, N101);
buf BUF1 (N412, N407);
nand NAND3 (N413, N412, N245, N68);
xor XOR2 (N414, N400, N121);
not NOT1 (N415, N411);
buf BUF1 (N416, N379);
or OR4 (N417, N413, N88, N263, N397);
or OR4 (N418, N396, N47, N394, N148);
and AND2 (N419, N392, N53);
nand NAND3 (N420, N418, N184, N148);
xor XOR2 (N421, N410, N92);
and AND2 (N422, N399, N228);
nand NAND2 (N423, N417, N76);
buf BUF1 (N424, N414);
nand NAND3 (N425, N423, N261, N169);
nor NOR2 (N426, N416, N177);
buf BUF1 (N427, N420);
or OR2 (N428, N425, N148);
buf BUF1 (N429, N426);
xor XOR2 (N430, N424, N93);
xor XOR2 (N431, N419, N124);
and AND4 (N432, N408, N136, N64, N311);
and AND3 (N433, N422, N139, N425);
buf BUF1 (N434, N427);
nor NOR3 (N435, N421, N215, N309);
not NOT1 (N436, N433);
not NOT1 (N437, N415);
not NOT1 (N438, N428);
or OR3 (N439, N403, N393, N383);
and AND2 (N440, N434, N294);
nand NAND4 (N441, N429, N417, N190, N193);
and AND4 (N442, N437, N217, N413, N314);
xor XOR2 (N443, N440, N370);
nor NOR4 (N444, N443, N36, N260, N215);
nor NOR3 (N445, N435, N275, N183);
and AND4 (N446, N441, N212, N8, N42);
xor XOR2 (N447, N431, N368);
and AND2 (N448, N430, N374);
and AND3 (N449, N442, N382, N46);
nor NOR2 (N450, N448, N205);
nor NOR3 (N451, N444, N198, N185);
buf BUF1 (N452, N447);
and AND2 (N453, N439, N268);
and AND3 (N454, N450, N67, N189);
nand NAND3 (N455, N436, N297, N372);
or OR4 (N456, N445, N327, N135, N368);
not NOT1 (N457, N456);
or OR3 (N458, N453, N314, N2);
nand NAND2 (N459, N457, N113);
nand NAND3 (N460, N455, N288, N58);
not NOT1 (N461, N459);
not NOT1 (N462, N458);
nand NAND4 (N463, N452, N401, N399, N281);
and AND3 (N464, N438, N169, N174);
not NOT1 (N465, N461);
nand NAND3 (N466, N446, N223, N428);
buf BUF1 (N467, N463);
xor XOR2 (N468, N464, N456);
not NOT1 (N469, N466);
not NOT1 (N470, N460);
nand NAND4 (N471, N468, N8, N317, N381);
xor XOR2 (N472, N462, N430);
not NOT1 (N473, N469);
not NOT1 (N474, N473);
nor NOR3 (N475, N432, N344, N113);
nor NOR2 (N476, N451, N363);
and AND2 (N477, N449, N274);
nor NOR4 (N478, N454, N161, N272, N30);
xor XOR2 (N479, N475, N397);
nor NOR4 (N480, N476, N277, N138, N312);
not NOT1 (N481, N472);
and AND2 (N482, N467, N242);
xor XOR2 (N483, N465, N94);
buf BUF1 (N484, N479);
or OR4 (N485, N470, N389, N189, N390);
buf BUF1 (N486, N478);
xor XOR2 (N487, N486, N80);
xor XOR2 (N488, N477, N258);
not NOT1 (N489, N471);
not NOT1 (N490, N485);
xor XOR2 (N491, N482, N76);
and AND2 (N492, N481, N421);
xor XOR2 (N493, N487, N239);
nor NOR3 (N494, N493, N435, N162);
not NOT1 (N495, N483);
and AND3 (N496, N490, N197, N153);
and AND3 (N497, N496, N423, N320);
not NOT1 (N498, N497);
and AND3 (N499, N474, N248, N11);
and AND4 (N500, N492, N395, N125, N486);
and AND2 (N501, N489, N42);
or OR4 (N502, N495, N208, N200, N384);
not NOT1 (N503, N501);
and AND2 (N504, N502, N31);
or OR2 (N505, N491, N214);
or OR2 (N506, N494, N131);
and AND4 (N507, N506, N501, N419, N133);
or OR2 (N508, N484, N101);
buf BUF1 (N509, N508);
nor NOR3 (N510, N509, N259, N486);
not NOT1 (N511, N500);
not NOT1 (N512, N488);
nor NOR4 (N513, N512, N364, N115, N56);
and AND3 (N514, N505, N159, N188);
not NOT1 (N515, N514);
nor NOR2 (N516, N504, N145);
nor NOR4 (N517, N480, N309, N511, N447);
and AND2 (N518, N128, N149);
xor XOR2 (N519, N507, N44);
or OR4 (N520, N510, N121, N279, N450);
or OR2 (N521, N520, N332);
nand NAND3 (N522, N516, N72, N385);
nand NAND3 (N523, N521, N402, N65);
nand NAND3 (N524, N519, N472, N89);
not NOT1 (N525, N513);
or OR4 (N526, N498, N382, N493, N333);
buf BUF1 (N527, N524);
not NOT1 (N528, N499);
buf BUF1 (N529, N503);
and AND2 (N530, N529, N353);
buf BUF1 (N531, N527);
or OR3 (N532, N515, N176, N48);
not NOT1 (N533, N523);
nand NAND2 (N534, N518, N206);
nand NAND2 (N535, N517, N334);
and AND3 (N536, N532, N123, N102);
nor NOR4 (N537, N525, N382, N185, N418);
and AND4 (N538, N533, N454, N384, N383);
xor XOR2 (N539, N538, N263);
or OR2 (N540, N530, N312);
nand NAND3 (N541, N522, N24, N381);
not NOT1 (N542, N539);
nor NOR4 (N543, N534, N298, N235, N446);
nand NAND4 (N544, N540, N540, N444, N248);
buf BUF1 (N545, N537);
nor NOR2 (N546, N526, N319);
nand NAND3 (N547, N536, N113, N77);
and AND2 (N548, N531, N315);
or OR3 (N549, N544, N447, N32);
buf BUF1 (N550, N549);
xor XOR2 (N551, N547, N272);
nand NAND2 (N552, N545, N380);
nand NAND4 (N553, N541, N489, N90, N270);
xor XOR2 (N554, N543, N376);
or OR2 (N555, N535, N439);
not NOT1 (N556, N548);
not NOT1 (N557, N546);
xor XOR2 (N558, N556, N1);
nor NOR4 (N559, N553, N112, N238, N320);
nand NAND2 (N560, N557, N347);
and AND4 (N561, N552, N475, N508, N545);
xor XOR2 (N562, N555, N210);
nor NOR3 (N563, N559, N460, N248);
nand NAND3 (N564, N550, N87, N75);
nor NOR2 (N565, N561, N246);
xor XOR2 (N566, N563, N530);
nand NAND3 (N567, N565, N178, N201);
not NOT1 (N568, N542);
nand NAND2 (N569, N564, N416);
or OR2 (N570, N568, N288);
buf BUF1 (N571, N528);
nand NAND2 (N572, N571, N328);
nand NAND3 (N573, N558, N223, N427);
nor NOR2 (N574, N567, N516);
not NOT1 (N575, N562);
nand NAND4 (N576, N554, N221, N11, N403);
nand NAND2 (N577, N569, N70);
buf BUF1 (N578, N575);
nand NAND4 (N579, N566, N257, N71, N539);
buf BUF1 (N580, N574);
buf BUF1 (N581, N572);
nand NAND3 (N582, N576, N358, N49);
not NOT1 (N583, N580);
xor XOR2 (N584, N577, N140);
xor XOR2 (N585, N582, N513);
and AND3 (N586, N560, N382, N394);
or OR4 (N587, N579, N357, N8, N109);
nor NOR4 (N588, N585, N110, N147, N482);
nor NOR2 (N589, N588, N486);
nand NAND3 (N590, N570, N136, N56);
nand NAND4 (N591, N583, N473, N14, N210);
buf BUF1 (N592, N590);
nand NAND4 (N593, N581, N144, N320, N31);
or OR2 (N594, N578, N325);
or OR3 (N595, N592, N559, N458);
xor XOR2 (N596, N551, N267);
or OR4 (N597, N593, N442, N201, N231);
and AND2 (N598, N597, N470);
buf BUF1 (N599, N591);
xor XOR2 (N600, N589, N325);
not NOT1 (N601, N596);
or OR2 (N602, N587, N551);
not NOT1 (N603, N599);
or OR2 (N604, N602, N602);
xor XOR2 (N605, N573, N195);
not NOT1 (N606, N604);
nor NOR3 (N607, N606, N411, N135);
buf BUF1 (N608, N605);
not NOT1 (N609, N608);
nor NOR2 (N610, N594, N486);
xor XOR2 (N611, N607, N394);
or OR4 (N612, N609, N299, N425, N386);
nor NOR2 (N613, N611, N492);
nor NOR3 (N614, N595, N118, N431);
not NOT1 (N615, N613);
and AND2 (N616, N610, N209);
or OR3 (N617, N598, N89, N406);
xor XOR2 (N618, N601, N296);
nor NOR3 (N619, N584, N73, N370);
buf BUF1 (N620, N618);
nand NAND2 (N621, N614, N30);
and AND2 (N622, N620, N302);
or OR3 (N623, N617, N177, N337);
nor NOR2 (N624, N615, N327);
or OR2 (N625, N586, N484);
xor XOR2 (N626, N612, N59);
nand NAND4 (N627, N623, N497, N419, N236);
and AND4 (N628, N619, N81, N559, N564);
nor NOR4 (N629, N627, N215, N419, N95);
xor XOR2 (N630, N600, N245);
nand NAND3 (N631, N616, N268, N335);
nand NAND3 (N632, N621, N276, N309);
or OR2 (N633, N630, N45);
or OR2 (N634, N628, N208);
nor NOR3 (N635, N633, N420, N616);
and AND3 (N636, N629, N532, N192);
not NOT1 (N637, N626);
buf BUF1 (N638, N634);
xor XOR2 (N639, N635, N49);
nor NOR4 (N640, N624, N498, N308, N539);
not NOT1 (N641, N639);
and AND4 (N642, N637, N316, N320, N176);
or OR2 (N643, N603, N9);
and AND2 (N644, N641, N405);
nor NOR2 (N645, N642, N531);
not NOT1 (N646, N622);
buf BUF1 (N647, N636);
xor XOR2 (N648, N625, N293);
nor NOR3 (N649, N632, N148, N496);
or OR3 (N650, N649, N593, N331);
and AND3 (N651, N640, N639, N273);
nand NAND4 (N652, N646, N622, N462, N481);
or OR2 (N653, N648, N417);
buf BUF1 (N654, N647);
xor XOR2 (N655, N631, N80);
or OR3 (N656, N650, N540, N395);
or OR4 (N657, N656, N632, N432, N374);
nand NAND2 (N658, N643, N307);
xor XOR2 (N659, N652, N277);
or OR3 (N660, N657, N612, N94);
nor NOR4 (N661, N655, N333, N584, N27);
nand NAND3 (N662, N654, N51, N308);
or OR4 (N663, N638, N192, N268, N163);
xor XOR2 (N664, N662, N456);
nor NOR3 (N665, N660, N453, N169);
or OR4 (N666, N664, N159, N69, N311);
xor XOR2 (N667, N653, N345);
xor XOR2 (N668, N666, N456);
xor XOR2 (N669, N651, N238);
and AND3 (N670, N659, N159, N190);
and AND3 (N671, N669, N76, N164);
buf BUF1 (N672, N665);
nor NOR3 (N673, N672, N50, N522);
nand NAND2 (N674, N670, N347);
and AND3 (N675, N661, N135, N76);
nand NAND4 (N676, N674, N49, N581, N596);
nor NOR3 (N677, N671, N172, N185);
nor NOR4 (N678, N675, N156, N108, N247);
buf BUF1 (N679, N663);
and AND2 (N680, N667, N333);
not NOT1 (N681, N658);
or OR2 (N682, N678, N438);
nor NOR4 (N683, N645, N653, N272, N88);
nor NOR4 (N684, N679, N262, N505, N73);
nand NAND4 (N685, N676, N305, N125, N626);
nand NAND2 (N686, N682, N102);
nand NAND4 (N687, N673, N116, N82, N642);
nor NOR2 (N688, N644, N78);
not NOT1 (N689, N681);
nand NAND4 (N690, N686, N400, N514, N206);
and AND4 (N691, N688, N280, N682, N11);
nand NAND2 (N692, N677, N147);
or OR3 (N693, N692, N657, N353);
not NOT1 (N694, N691);
not NOT1 (N695, N680);
not NOT1 (N696, N690);
and AND4 (N697, N684, N678, N132, N409);
or OR4 (N698, N683, N212, N164, N418);
xor XOR2 (N699, N685, N381);
xor XOR2 (N700, N699, N148);
not NOT1 (N701, N697);
and AND4 (N702, N687, N389, N162, N80);
buf BUF1 (N703, N700);
buf BUF1 (N704, N668);
nand NAND4 (N705, N694, N24, N261, N232);
and AND4 (N706, N703, N346, N69, N523);
or OR2 (N707, N705, N355);
and AND4 (N708, N693, N81, N455, N651);
or OR4 (N709, N702, N301, N707, N345);
not NOT1 (N710, N289);
and AND4 (N711, N689, N149, N649, N239);
buf BUF1 (N712, N701);
nor NOR3 (N713, N708, N49, N561);
nor NOR3 (N714, N712, N164, N562);
not NOT1 (N715, N704);
buf BUF1 (N716, N713);
or OR3 (N717, N716, N711, N524);
xor XOR2 (N718, N622, N64);
nand NAND4 (N719, N710, N539, N324, N52);
buf BUF1 (N720, N696);
and AND4 (N721, N706, N188, N159, N348);
nor NOR3 (N722, N709, N195, N563);
nand NAND3 (N723, N722, N388, N19);
and AND2 (N724, N714, N577);
xor XOR2 (N725, N721, N180);
or OR4 (N726, N724, N681, N468, N207);
or OR3 (N727, N698, N490, N689);
buf BUF1 (N728, N695);
xor XOR2 (N729, N720, N654);
xor XOR2 (N730, N728, N27);
buf BUF1 (N731, N726);
xor XOR2 (N732, N715, N426);
xor XOR2 (N733, N717, N458);
not NOT1 (N734, N731);
or OR4 (N735, N719, N492, N628, N667);
nor NOR2 (N736, N735, N735);
buf BUF1 (N737, N730);
not NOT1 (N738, N718);
and AND2 (N739, N725, N355);
xor XOR2 (N740, N736, N421);
nor NOR2 (N741, N734, N275);
not NOT1 (N742, N733);
buf BUF1 (N743, N740);
xor XOR2 (N744, N727, N435);
or OR3 (N745, N744, N235, N208);
or OR4 (N746, N737, N631, N477, N351);
xor XOR2 (N747, N739, N15);
buf BUF1 (N748, N732);
buf BUF1 (N749, N742);
nand NAND4 (N750, N723, N80, N171, N417);
buf BUF1 (N751, N745);
or OR2 (N752, N746, N131);
not NOT1 (N753, N743);
buf BUF1 (N754, N738);
and AND3 (N755, N754, N116, N679);
nor NOR2 (N756, N755, N661);
nor NOR2 (N757, N749, N580);
nand NAND2 (N758, N752, N483);
nor NOR2 (N759, N758, N727);
not NOT1 (N760, N756);
nand NAND4 (N761, N757, N118, N291, N187);
nor NOR2 (N762, N759, N372);
or OR4 (N763, N760, N717, N369, N22);
nand NAND4 (N764, N747, N501, N109, N419);
xor XOR2 (N765, N764, N726);
nor NOR4 (N766, N763, N538, N78, N439);
not NOT1 (N767, N729);
not NOT1 (N768, N761);
or OR2 (N769, N748, N720);
nand NAND4 (N770, N766, N46, N15, N623);
buf BUF1 (N771, N750);
nor NOR4 (N772, N771, N32, N611, N283);
nor NOR2 (N773, N765, N250);
buf BUF1 (N774, N773);
nor NOR3 (N775, N753, N620, N303);
buf BUF1 (N776, N770);
not NOT1 (N777, N767);
xor XOR2 (N778, N774, N230);
nand NAND2 (N779, N762, N715);
nand NAND2 (N780, N776, N445);
xor XOR2 (N781, N772, N633);
nor NOR2 (N782, N741, N63);
buf BUF1 (N783, N768);
buf BUF1 (N784, N775);
not NOT1 (N785, N783);
not NOT1 (N786, N779);
not NOT1 (N787, N751);
xor XOR2 (N788, N781, N710);
buf BUF1 (N789, N788);
or OR3 (N790, N778, N685, N643);
not NOT1 (N791, N785);
or OR3 (N792, N784, N2, N151);
xor XOR2 (N793, N791, N298);
buf BUF1 (N794, N787);
or OR4 (N795, N780, N395, N357, N534);
nand NAND2 (N796, N792, N548);
not NOT1 (N797, N777);
not NOT1 (N798, N793);
not NOT1 (N799, N769);
and AND2 (N800, N789, N772);
and AND2 (N801, N796, N606);
xor XOR2 (N802, N786, N733);
nor NOR4 (N803, N802, N244, N475, N695);
or OR4 (N804, N799, N60, N338, N586);
xor XOR2 (N805, N795, N404);
nor NOR3 (N806, N794, N10, N3);
buf BUF1 (N807, N803);
or OR3 (N808, N800, N704, N137);
buf BUF1 (N809, N805);
not NOT1 (N810, N790);
not NOT1 (N811, N808);
not NOT1 (N812, N782);
nand NAND4 (N813, N806, N255, N635, N199);
and AND2 (N814, N810, N86);
xor XOR2 (N815, N798, N34);
or OR3 (N816, N797, N615, N333);
nand NAND4 (N817, N816, N107, N438, N437);
or OR4 (N818, N804, N601, N605, N655);
nand NAND4 (N819, N811, N532, N216, N107);
not NOT1 (N820, N819);
nor NOR4 (N821, N817, N1, N325, N50);
buf BUF1 (N822, N815);
and AND2 (N823, N818, N675);
not NOT1 (N824, N809);
xor XOR2 (N825, N820, N344);
xor XOR2 (N826, N824, N144);
nand NAND3 (N827, N812, N119, N197);
or OR3 (N828, N821, N494, N14);
or OR2 (N829, N828, N133);
buf BUF1 (N830, N825);
buf BUF1 (N831, N813);
buf BUF1 (N832, N807);
and AND2 (N833, N829, N260);
buf BUF1 (N834, N823);
nand NAND3 (N835, N827, N369, N478);
and AND3 (N836, N822, N38, N523);
not NOT1 (N837, N814);
buf BUF1 (N838, N801);
and AND2 (N839, N826, N382);
nor NOR4 (N840, N837, N368, N744, N793);
and AND2 (N841, N834, N31);
xor XOR2 (N842, N839, N190);
nor NOR4 (N843, N832, N814, N505, N94);
nand NAND3 (N844, N830, N93, N748);
buf BUF1 (N845, N835);
nand NAND4 (N846, N843, N469, N427, N600);
xor XOR2 (N847, N846, N73);
and AND3 (N848, N836, N567, N247);
and AND3 (N849, N838, N96, N79);
or OR4 (N850, N842, N410, N574, N458);
or OR3 (N851, N833, N149, N299);
or OR3 (N852, N849, N481, N243);
not NOT1 (N853, N844);
buf BUF1 (N854, N831);
not NOT1 (N855, N841);
nand NAND4 (N856, N848, N381, N628, N596);
nand NAND2 (N857, N856, N655);
or OR2 (N858, N850, N3);
buf BUF1 (N859, N852);
not NOT1 (N860, N845);
not NOT1 (N861, N840);
xor XOR2 (N862, N858, N333);
nand NAND4 (N863, N860, N475, N827, N415);
xor XOR2 (N864, N861, N84);
xor XOR2 (N865, N862, N713);
nand NAND3 (N866, N853, N455, N729);
buf BUF1 (N867, N859);
xor XOR2 (N868, N857, N781);
or OR3 (N869, N867, N537, N743);
xor XOR2 (N870, N864, N216);
nor NOR4 (N871, N863, N184, N592, N172);
and AND4 (N872, N868, N566, N248, N713);
buf BUF1 (N873, N847);
xor XOR2 (N874, N854, N592);
and AND2 (N875, N872, N246);
nand NAND2 (N876, N874, N848);
not NOT1 (N877, N871);
and AND3 (N878, N869, N622, N238);
nor NOR3 (N879, N876, N360, N92);
nand NAND4 (N880, N870, N296, N425, N423);
xor XOR2 (N881, N875, N676);
not NOT1 (N882, N880);
nand NAND4 (N883, N879, N449, N58, N560);
not NOT1 (N884, N881);
xor XOR2 (N885, N851, N276);
not NOT1 (N886, N866);
buf BUF1 (N887, N885);
or OR3 (N888, N887, N463, N170);
xor XOR2 (N889, N878, N748);
not NOT1 (N890, N877);
xor XOR2 (N891, N883, N154);
nand NAND3 (N892, N889, N201, N146);
nor NOR4 (N893, N886, N604, N72, N305);
buf BUF1 (N894, N891);
buf BUF1 (N895, N855);
not NOT1 (N896, N882);
xor XOR2 (N897, N873, N392);
xor XOR2 (N898, N893, N552);
and AND2 (N899, N896, N844);
nand NAND3 (N900, N898, N231, N845);
or OR2 (N901, N890, N403);
buf BUF1 (N902, N901);
not NOT1 (N903, N865);
and AND2 (N904, N903, N64);
nand NAND2 (N905, N884, N4);
buf BUF1 (N906, N897);
xor XOR2 (N907, N904, N464);
nor NOR2 (N908, N902, N543);
nand NAND3 (N909, N908, N898, N576);
and AND3 (N910, N907, N611, N725);
buf BUF1 (N911, N905);
not NOT1 (N912, N910);
nand NAND2 (N913, N911, N854);
not NOT1 (N914, N894);
buf BUF1 (N915, N900);
nor NOR3 (N916, N895, N32, N812);
nand NAND4 (N917, N916, N868, N425, N278);
xor XOR2 (N918, N906, N716);
buf BUF1 (N919, N912);
xor XOR2 (N920, N918, N146);
nor NOR4 (N921, N919, N494, N9, N439);
nor NOR2 (N922, N899, N892);
nand NAND3 (N923, N123, N711, N316);
and AND3 (N924, N922, N907, N29);
buf BUF1 (N925, N921);
and AND3 (N926, N924, N324, N790);
or OR2 (N927, N888, N333);
nor NOR4 (N928, N927, N484, N144, N568);
nor NOR4 (N929, N926, N27, N31, N627);
and AND3 (N930, N920, N162, N748);
and AND3 (N931, N913, N816, N815);
buf BUF1 (N932, N915);
nor NOR2 (N933, N930, N366);
and AND3 (N934, N923, N259, N570);
nor NOR3 (N935, N931, N552, N490);
buf BUF1 (N936, N928);
and AND2 (N937, N933, N313);
not NOT1 (N938, N937);
not NOT1 (N939, N938);
buf BUF1 (N940, N914);
xor XOR2 (N941, N940, N262);
or OR2 (N942, N917, N25);
or OR4 (N943, N909, N380, N482, N681);
and AND4 (N944, N925, N744, N33, N159);
xor XOR2 (N945, N934, N102);
xor XOR2 (N946, N945, N733);
nor NOR3 (N947, N929, N167, N267);
or OR2 (N948, N946, N676);
and AND4 (N949, N942, N402, N361, N220);
not NOT1 (N950, N932);
nor NOR4 (N951, N936, N613, N832, N175);
nand NAND2 (N952, N947, N442);
xor XOR2 (N953, N944, N949);
nor NOR2 (N954, N763, N398);
xor XOR2 (N955, N943, N347);
not NOT1 (N956, N955);
not NOT1 (N957, N941);
nand NAND3 (N958, N950, N740, N681);
and AND2 (N959, N956, N419);
nand NAND3 (N960, N951, N18, N392);
xor XOR2 (N961, N960, N843);
buf BUF1 (N962, N952);
xor XOR2 (N963, N954, N104);
and AND2 (N964, N948, N474);
nor NOR4 (N965, N959, N553, N835, N197);
nor NOR4 (N966, N962, N716, N592, N200);
buf BUF1 (N967, N963);
buf BUF1 (N968, N965);
nor NOR4 (N969, N953, N912, N415, N295);
or OR3 (N970, N939, N203, N673);
not NOT1 (N971, N961);
buf BUF1 (N972, N968);
nor NOR2 (N973, N967, N961);
xor XOR2 (N974, N969, N836);
nor NOR2 (N975, N973, N950);
not NOT1 (N976, N966);
and AND3 (N977, N975, N282, N924);
not NOT1 (N978, N974);
or OR3 (N979, N957, N569, N670);
nand NAND3 (N980, N935, N286, N546);
xor XOR2 (N981, N976, N826);
nor NOR2 (N982, N978, N29);
nand NAND3 (N983, N972, N536, N12);
nor NOR4 (N984, N970, N716, N878, N818);
nand NAND3 (N985, N984, N978, N512);
nand NAND3 (N986, N958, N494, N79);
and AND3 (N987, N982, N508, N386);
buf BUF1 (N988, N980);
not NOT1 (N989, N964);
buf BUF1 (N990, N988);
nor NOR2 (N991, N986, N468);
and AND2 (N992, N977, N36);
xor XOR2 (N993, N991, N66);
nand NAND4 (N994, N971, N518, N373, N752);
and AND2 (N995, N992, N752);
nor NOR4 (N996, N989, N189, N652, N76);
nand NAND3 (N997, N983, N800, N57);
xor XOR2 (N998, N994, N539);
and AND3 (N999, N981, N432, N773);
nand NAND3 (N1000, N985, N773, N240);
or OR4 (N1001, N998, N149, N592, N279);
nor NOR3 (N1002, N990, N495, N894);
buf BUF1 (N1003, N979);
or OR2 (N1004, N1003, N414);
and AND2 (N1005, N987, N328);
or OR3 (N1006, N995, N283, N410);
and AND3 (N1007, N1006, N543, N156);
buf BUF1 (N1008, N1007);
not NOT1 (N1009, N1000);
buf BUF1 (N1010, N993);
nand NAND2 (N1011, N1008, N631);
nand NAND4 (N1012, N999, N504, N706, N411);
buf BUF1 (N1013, N1011);
nor NOR4 (N1014, N1012, N512, N492, N323);
or OR4 (N1015, N1009, N884, N917, N696);
nand NAND2 (N1016, N1004, N532);
or OR3 (N1017, N1013, N932, N343);
buf BUF1 (N1018, N997);
nor NOR4 (N1019, N1005, N989, N832, N659);
or OR4 (N1020, N1016, N3, N223, N848);
nand NAND4 (N1021, N1018, N43, N616, N862);
nand NAND2 (N1022, N1010, N430);
nand NAND3 (N1023, N1019, N868, N751);
and AND3 (N1024, N1021, N852, N153);
or OR2 (N1025, N1023, N167);
not NOT1 (N1026, N1024);
not NOT1 (N1027, N1015);
not NOT1 (N1028, N1022);
nand NAND4 (N1029, N1027, N936, N614, N320);
nand NAND4 (N1030, N1002, N935, N24, N428);
not NOT1 (N1031, N1030);
or OR4 (N1032, N1031, N152, N816, N938);
or OR3 (N1033, N1017, N945, N649);
and AND4 (N1034, N1029, N632, N411, N553);
or OR3 (N1035, N1020, N618, N341);
buf BUF1 (N1036, N1026);
and AND2 (N1037, N996, N756);
nor NOR2 (N1038, N1032, N272);
not NOT1 (N1039, N1037);
nand NAND3 (N1040, N1014, N486, N43);
not NOT1 (N1041, N1028);
nand NAND3 (N1042, N1001, N253, N387);
buf BUF1 (N1043, N1034);
nand NAND3 (N1044, N1041, N476, N1009);
buf BUF1 (N1045, N1035);
buf BUF1 (N1046, N1045);
xor XOR2 (N1047, N1039, N264);
not NOT1 (N1048, N1043);
xor XOR2 (N1049, N1025, N339);
buf BUF1 (N1050, N1046);
or OR2 (N1051, N1038, N275);
nand NAND2 (N1052, N1040, N156);
buf BUF1 (N1053, N1050);
or OR4 (N1054, N1048, N356, N1000, N650);
nor NOR4 (N1055, N1053, N258, N700, N624);
and AND3 (N1056, N1036, N77, N121);
xor XOR2 (N1057, N1047, N133);
nand NAND2 (N1058, N1057, N862);
buf BUF1 (N1059, N1042);
nand NAND2 (N1060, N1054, N291);
not NOT1 (N1061, N1058);
nor NOR4 (N1062, N1061, N727, N461, N778);
or OR4 (N1063, N1060, N818, N690, N24);
or OR3 (N1064, N1033, N1011, N74);
nor NOR3 (N1065, N1049, N307, N40);
not NOT1 (N1066, N1059);
not NOT1 (N1067, N1062);
and AND2 (N1068, N1051, N905);
or OR4 (N1069, N1056, N459, N769, N827);
nand NAND3 (N1070, N1067, N772, N346);
not NOT1 (N1071, N1064);
nand NAND4 (N1072, N1063, N818, N905, N230);
not NOT1 (N1073, N1071);
nand NAND2 (N1074, N1065, N556);
nor NOR4 (N1075, N1072, N860, N461, N1023);
buf BUF1 (N1076, N1044);
or OR4 (N1077, N1074, N351, N163, N541);
nand NAND3 (N1078, N1069, N832, N53);
and AND4 (N1079, N1070, N582, N552, N133);
and AND2 (N1080, N1066, N480);
not NOT1 (N1081, N1068);
nor NOR4 (N1082, N1077, N125, N236, N978);
not NOT1 (N1083, N1078);
nor NOR2 (N1084, N1055, N347);
and AND3 (N1085, N1076, N879, N888);
or OR2 (N1086, N1082, N190);
and AND3 (N1087, N1073, N706, N349);
xor XOR2 (N1088, N1079, N690);
or OR2 (N1089, N1084, N443);
not NOT1 (N1090, N1086);
xor XOR2 (N1091, N1085, N877);
xor XOR2 (N1092, N1075, N833);
and AND2 (N1093, N1090, N957);
nor NOR3 (N1094, N1052, N750, N302);
nor NOR2 (N1095, N1083, N151);
nand NAND3 (N1096, N1095, N157, N269);
and AND2 (N1097, N1096, N153);
or OR2 (N1098, N1087, N194);
nand NAND3 (N1099, N1097, N325, N493);
nor NOR3 (N1100, N1092, N943, N719);
nand NAND2 (N1101, N1080, N523);
nand NAND2 (N1102, N1089, N59);
nand NAND4 (N1103, N1093, N1003, N410, N411);
and AND2 (N1104, N1100, N1044);
xor XOR2 (N1105, N1088, N128);
buf BUF1 (N1106, N1091);
nand NAND4 (N1107, N1101, N497, N89, N358);
not NOT1 (N1108, N1105);
or OR2 (N1109, N1107, N602);
not NOT1 (N1110, N1094);
or OR2 (N1111, N1081, N409);
or OR3 (N1112, N1110, N1090, N69);
not NOT1 (N1113, N1098);
and AND2 (N1114, N1113, N455);
xor XOR2 (N1115, N1108, N990);
xor XOR2 (N1116, N1102, N794);
nor NOR4 (N1117, N1103, N971, N994, N301);
or OR3 (N1118, N1111, N82, N165);
buf BUF1 (N1119, N1115);
and AND2 (N1120, N1114, N388);
nand NAND4 (N1121, N1106, N925, N1078, N642);
or OR3 (N1122, N1116, N225, N171);
or OR2 (N1123, N1117, N503);
nor NOR3 (N1124, N1121, N884, N153);
and AND4 (N1125, N1122, N884, N70, N587);
and AND4 (N1126, N1099, N269, N183, N645);
buf BUF1 (N1127, N1119);
xor XOR2 (N1128, N1104, N619);
not NOT1 (N1129, N1118);
xor XOR2 (N1130, N1127, N609);
buf BUF1 (N1131, N1120);
xor XOR2 (N1132, N1112, N722);
or OR4 (N1133, N1131, N70, N367, N848);
not NOT1 (N1134, N1124);
and AND2 (N1135, N1134, N220);
xor XOR2 (N1136, N1133, N576);
nor NOR4 (N1137, N1109, N481, N1064, N706);
not NOT1 (N1138, N1128);
xor XOR2 (N1139, N1129, N839);
or OR4 (N1140, N1139, N1111, N613, N350);
buf BUF1 (N1141, N1136);
nor NOR4 (N1142, N1126, N478, N1130, N170);
not NOT1 (N1143, N191);
or OR3 (N1144, N1141, N202, N469);
buf BUF1 (N1145, N1143);
xor XOR2 (N1146, N1132, N1137);
and AND2 (N1147, N451, N100);
nor NOR3 (N1148, N1145, N343, N221);
nor NOR2 (N1149, N1146, N210);
nand NAND2 (N1150, N1144, N711);
nor NOR4 (N1151, N1138, N75, N245, N465);
nor NOR3 (N1152, N1148, N683, N1137);
nor NOR4 (N1153, N1123, N976, N840, N204);
xor XOR2 (N1154, N1140, N1022);
not NOT1 (N1155, N1153);
nor NOR2 (N1156, N1149, N110);
xor XOR2 (N1157, N1154, N77);
or OR3 (N1158, N1151, N738, N188);
nand NAND2 (N1159, N1147, N1151);
or OR3 (N1160, N1150, N33, N14);
xor XOR2 (N1161, N1156, N1055);
not NOT1 (N1162, N1158);
or OR4 (N1163, N1161, N837, N866, N598);
and AND2 (N1164, N1155, N972);
not NOT1 (N1165, N1142);
xor XOR2 (N1166, N1164, N51);
not NOT1 (N1167, N1160);
buf BUF1 (N1168, N1159);
and AND2 (N1169, N1125, N457);
or OR3 (N1170, N1168, N760, N672);
nand NAND2 (N1171, N1135, N399);
not NOT1 (N1172, N1169);
xor XOR2 (N1173, N1165, N940);
not NOT1 (N1174, N1173);
not NOT1 (N1175, N1157);
buf BUF1 (N1176, N1175);
nand NAND2 (N1177, N1167, N363);
nand NAND3 (N1178, N1170, N94, N341);
xor XOR2 (N1179, N1174, N64);
not NOT1 (N1180, N1178);
and AND3 (N1181, N1179, N1060, N53);
and AND4 (N1182, N1181, N551, N423, N171);
not NOT1 (N1183, N1163);
not NOT1 (N1184, N1171);
not NOT1 (N1185, N1183);
nor NOR4 (N1186, N1162, N301, N1015, N845);
nor NOR2 (N1187, N1182, N624);
and AND4 (N1188, N1184, N771, N345, N421);
buf BUF1 (N1189, N1188);
xor XOR2 (N1190, N1189, N485);
xor XOR2 (N1191, N1186, N255);
and AND2 (N1192, N1180, N950);
or OR3 (N1193, N1192, N397, N399);
nor NOR2 (N1194, N1187, N500);
buf BUF1 (N1195, N1191);
and AND3 (N1196, N1185, N1118, N898);
nand NAND3 (N1197, N1177, N856, N327);
buf BUF1 (N1198, N1193);
buf BUF1 (N1199, N1152);
nand NAND4 (N1200, N1176, N1015, N841, N998);
buf BUF1 (N1201, N1196);
nor NOR4 (N1202, N1201, N951, N98, N40);
nand NAND2 (N1203, N1194, N906);
xor XOR2 (N1204, N1198, N918);
or OR3 (N1205, N1166, N975, N175);
nor NOR2 (N1206, N1203, N712);
or OR3 (N1207, N1206, N729, N212);
buf BUF1 (N1208, N1172);
nand NAND3 (N1209, N1200, N716, N785);
and AND3 (N1210, N1195, N617, N1006);
xor XOR2 (N1211, N1208, N588);
nand NAND3 (N1212, N1209, N256, N249);
not NOT1 (N1213, N1197);
xor XOR2 (N1214, N1204, N111);
and AND2 (N1215, N1190, N700);
not NOT1 (N1216, N1212);
not NOT1 (N1217, N1207);
nand NAND3 (N1218, N1217, N726, N1046);
and AND3 (N1219, N1218, N841, N529);
xor XOR2 (N1220, N1210, N146);
or OR2 (N1221, N1199, N1175);
nor NOR4 (N1222, N1213, N92, N1125, N187);
buf BUF1 (N1223, N1222);
and AND2 (N1224, N1221, N363);
not NOT1 (N1225, N1215);
not NOT1 (N1226, N1225);
not NOT1 (N1227, N1211);
nor NOR4 (N1228, N1216, N373, N480, N1095);
or OR2 (N1229, N1219, N1153);
nand NAND4 (N1230, N1227, N564, N1035, N1064);
buf BUF1 (N1231, N1223);
xor XOR2 (N1232, N1205, N1167);
nand NAND4 (N1233, N1226, N917, N1075, N278);
buf BUF1 (N1234, N1229);
xor XOR2 (N1235, N1234, N73);
not NOT1 (N1236, N1202);
not NOT1 (N1237, N1214);
xor XOR2 (N1238, N1235, N810);
nand NAND2 (N1239, N1232, N853);
xor XOR2 (N1240, N1237, N1159);
or OR3 (N1241, N1224, N1224, N133);
not NOT1 (N1242, N1241);
nand NAND4 (N1243, N1240, N959, N992, N972);
or OR4 (N1244, N1230, N77, N154, N4);
nor NOR3 (N1245, N1244, N279, N1132);
buf BUF1 (N1246, N1242);
nor NOR3 (N1247, N1245, N1030, N450);
buf BUF1 (N1248, N1228);
nor NOR2 (N1249, N1238, N1207);
nor NOR3 (N1250, N1220, N320, N776);
buf BUF1 (N1251, N1233);
buf BUF1 (N1252, N1249);
and AND4 (N1253, N1251, N890, N225, N132);
buf BUF1 (N1254, N1253);
and AND4 (N1255, N1248, N715, N427, N660);
buf BUF1 (N1256, N1231);
buf BUF1 (N1257, N1247);
or OR3 (N1258, N1256, N234, N29);
nand NAND3 (N1259, N1243, N240, N417);
not NOT1 (N1260, N1250);
nor NOR2 (N1261, N1239, N920);
or OR3 (N1262, N1260, N560, N48);
xor XOR2 (N1263, N1252, N1162);
nand NAND3 (N1264, N1263, N455, N369);
buf BUF1 (N1265, N1262);
nor NOR2 (N1266, N1257, N1164);
or OR3 (N1267, N1266, N691, N486);
or OR4 (N1268, N1265, N826, N379, N620);
nand NAND4 (N1269, N1261, N709, N998, N995);
nor NOR2 (N1270, N1267, N869);
nand NAND2 (N1271, N1254, N945);
not NOT1 (N1272, N1264);
not NOT1 (N1273, N1258);
xor XOR2 (N1274, N1272, N539);
nor NOR3 (N1275, N1255, N580, N342);
and AND4 (N1276, N1236, N998, N847, N719);
or OR4 (N1277, N1271, N724, N195, N1019);
nor NOR4 (N1278, N1246, N1153, N654, N158);
not NOT1 (N1279, N1273);
and AND4 (N1280, N1274, N1087, N19, N1158);
nand NAND4 (N1281, N1259, N537, N861, N287);
nor NOR3 (N1282, N1269, N627, N230);
nor NOR4 (N1283, N1275, N1056, N494, N1158);
or OR2 (N1284, N1280, N880);
not NOT1 (N1285, N1281);
nor NOR3 (N1286, N1278, N987, N179);
nor NOR4 (N1287, N1284, N13, N225, N566);
nand NAND2 (N1288, N1276, N990);
or OR4 (N1289, N1286, N416, N720, N305);
nand NAND4 (N1290, N1277, N1135, N84, N540);
not NOT1 (N1291, N1289);
or OR3 (N1292, N1288, N1016, N1256);
not NOT1 (N1293, N1282);
and AND3 (N1294, N1287, N638, N1153);
nand NAND2 (N1295, N1270, N291);
buf BUF1 (N1296, N1285);
not NOT1 (N1297, N1290);
nor NOR4 (N1298, N1297, N862, N1017, N1245);
and AND3 (N1299, N1298, N791, N1009);
or OR3 (N1300, N1291, N1131, N1049);
not NOT1 (N1301, N1299);
nand NAND4 (N1302, N1292, N291, N145, N778);
nand NAND2 (N1303, N1295, N713);
not NOT1 (N1304, N1300);
and AND3 (N1305, N1304, N295, N529);
or OR2 (N1306, N1302, N970);
or OR4 (N1307, N1294, N898, N1059, N57);
xor XOR2 (N1308, N1301, N738);
buf BUF1 (N1309, N1307);
nand NAND3 (N1310, N1293, N496, N1124);
buf BUF1 (N1311, N1268);
and AND3 (N1312, N1311, N887, N323);
or OR3 (N1313, N1308, N21, N587);
and AND3 (N1314, N1296, N439, N845);
xor XOR2 (N1315, N1312, N843);
not NOT1 (N1316, N1315);
not NOT1 (N1317, N1303);
nor NOR2 (N1318, N1313, N715);
or OR4 (N1319, N1318, N725, N398, N537);
buf BUF1 (N1320, N1309);
nor NOR4 (N1321, N1310, N1310, N544, N512);
nand NAND3 (N1322, N1314, N976, N1139);
xor XOR2 (N1323, N1321, N130);
buf BUF1 (N1324, N1283);
and AND4 (N1325, N1316, N84, N422, N681);
buf BUF1 (N1326, N1305);
xor XOR2 (N1327, N1322, N1010);
nand NAND3 (N1328, N1317, N389, N995);
nand NAND4 (N1329, N1326, N595, N1141, N1088);
buf BUF1 (N1330, N1324);
or OR4 (N1331, N1323, N820, N1148, N1312);
and AND3 (N1332, N1328, N614, N361);
xor XOR2 (N1333, N1279, N54);
or OR2 (N1334, N1306, N1264);
xor XOR2 (N1335, N1334, N361);
xor XOR2 (N1336, N1319, N1281);
buf BUF1 (N1337, N1335);
nor NOR2 (N1338, N1336, N932);
not NOT1 (N1339, N1337);
buf BUF1 (N1340, N1325);
buf BUF1 (N1341, N1338);
nor NOR4 (N1342, N1332, N358, N691, N1328);
nor NOR4 (N1343, N1340, N114, N252, N438);
xor XOR2 (N1344, N1320, N35);
xor XOR2 (N1345, N1342, N208);
buf BUF1 (N1346, N1339);
nor NOR3 (N1347, N1330, N943, N4);
or OR4 (N1348, N1331, N311, N516, N407);
nand NAND3 (N1349, N1333, N988, N78);
or OR3 (N1350, N1345, N1045, N809);
xor XOR2 (N1351, N1344, N646);
nor NOR2 (N1352, N1346, N536);
not NOT1 (N1353, N1341);
not NOT1 (N1354, N1353);
or OR2 (N1355, N1347, N333);
nand NAND3 (N1356, N1355, N664, N530);
nand NAND2 (N1357, N1356, N1176);
xor XOR2 (N1358, N1351, N564);
or OR2 (N1359, N1350, N957);
nor NOR4 (N1360, N1359, N794, N365, N631);
or OR2 (N1361, N1329, N967);
nand NAND4 (N1362, N1348, N1176, N159, N1304);
nor NOR2 (N1363, N1358, N1209);
buf BUF1 (N1364, N1352);
nor NOR3 (N1365, N1343, N532, N647);
buf BUF1 (N1366, N1360);
not NOT1 (N1367, N1365);
nand NAND4 (N1368, N1366, N402, N1095, N1068);
and AND4 (N1369, N1361, N482, N279, N1025);
or OR3 (N1370, N1367, N885, N788);
not NOT1 (N1371, N1357);
buf BUF1 (N1372, N1349);
or OR2 (N1373, N1363, N848);
xor XOR2 (N1374, N1362, N1271);
or OR4 (N1375, N1369, N251, N318, N1324);
nand NAND3 (N1376, N1373, N466, N336);
nor NOR4 (N1377, N1368, N1094, N1000, N776);
nand NAND2 (N1378, N1364, N620);
nor NOR2 (N1379, N1376, N571);
xor XOR2 (N1380, N1372, N338);
xor XOR2 (N1381, N1378, N555);
not NOT1 (N1382, N1374);
nand NAND4 (N1383, N1380, N717, N490, N1071);
and AND3 (N1384, N1371, N462, N743);
nand NAND2 (N1385, N1383, N300);
nor NOR2 (N1386, N1375, N1318);
and AND2 (N1387, N1354, N1343);
or OR3 (N1388, N1385, N240, N729);
nor NOR3 (N1389, N1382, N625, N629);
or OR3 (N1390, N1327, N1192, N1030);
buf BUF1 (N1391, N1377);
nand NAND2 (N1392, N1388, N873);
buf BUF1 (N1393, N1384);
nand NAND3 (N1394, N1386, N1024, N556);
buf BUF1 (N1395, N1391);
and AND3 (N1396, N1395, N776, N986);
nand NAND2 (N1397, N1379, N393);
nor NOR2 (N1398, N1370, N196);
nand NAND2 (N1399, N1392, N22);
buf BUF1 (N1400, N1389);
buf BUF1 (N1401, N1397);
not NOT1 (N1402, N1401);
and AND3 (N1403, N1396, N545, N256);
not NOT1 (N1404, N1381);
not NOT1 (N1405, N1390);
and AND4 (N1406, N1404, N924, N1133, N1019);
nor NOR3 (N1407, N1405, N312, N939);
nor NOR3 (N1408, N1400, N960, N367);
buf BUF1 (N1409, N1403);
buf BUF1 (N1410, N1406);
buf BUF1 (N1411, N1402);
and AND3 (N1412, N1399, N700, N523);
xor XOR2 (N1413, N1408, N568);
xor XOR2 (N1414, N1410, N1070);
not NOT1 (N1415, N1393);
or OR2 (N1416, N1394, N1349);
xor XOR2 (N1417, N1409, N1275);
and AND3 (N1418, N1413, N1304, N264);
or OR4 (N1419, N1414, N982, N1381, N984);
nor NOR3 (N1420, N1411, N262, N876);
buf BUF1 (N1421, N1415);
and AND4 (N1422, N1417, N279, N827, N1260);
xor XOR2 (N1423, N1412, N176);
xor XOR2 (N1424, N1419, N1015);
buf BUF1 (N1425, N1423);
xor XOR2 (N1426, N1424, N544);
and AND4 (N1427, N1416, N1410, N13, N1377);
not NOT1 (N1428, N1387);
buf BUF1 (N1429, N1427);
not NOT1 (N1430, N1425);
buf BUF1 (N1431, N1426);
nor NOR2 (N1432, N1407, N796);
not NOT1 (N1433, N1420);
buf BUF1 (N1434, N1421);
nand NAND2 (N1435, N1431, N88);
and AND3 (N1436, N1418, N917, N745);
not NOT1 (N1437, N1432);
xor XOR2 (N1438, N1398, N815);
buf BUF1 (N1439, N1422);
and AND2 (N1440, N1429, N93);
and AND3 (N1441, N1437, N365, N935);
xor XOR2 (N1442, N1436, N600);
and AND2 (N1443, N1440, N602);
buf BUF1 (N1444, N1433);
xor XOR2 (N1445, N1442, N604);
nand NAND4 (N1446, N1428, N94, N787, N432);
nor NOR2 (N1447, N1438, N1435);
xor XOR2 (N1448, N26, N550);
not NOT1 (N1449, N1439);
or OR2 (N1450, N1446, N428);
not NOT1 (N1451, N1434);
and AND3 (N1452, N1450, N1086, N738);
xor XOR2 (N1453, N1448, N428);
buf BUF1 (N1454, N1449);
and AND3 (N1455, N1441, N110, N38);
nand NAND2 (N1456, N1445, N515);
and AND3 (N1457, N1451, N674, N669);
xor XOR2 (N1458, N1457, N165);
nor NOR2 (N1459, N1444, N1138);
or OR3 (N1460, N1458, N928, N224);
or OR3 (N1461, N1443, N236, N1166);
or OR2 (N1462, N1452, N595);
nand NAND3 (N1463, N1460, N686, N943);
xor XOR2 (N1464, N1454, N34);
nand NAND3 (N1465, N1455, N805, N699);
nor NOR3 (N1466, N1462, N247, N890);
xor XOR2 (N1467, N1453, N332);
buf BUF1 (N1468, N1456);
buf BUF1 (N1469, N1465);
xor XOR2 (N1470, N1468, N1076);
xor XOR2 (N1471, N1469, N1133);
and AND4 (N1472, N1467, N1028, N1082, N879);
not NOT1 (N1473, N1447);
nand NAND4 (N1474, N1470, N902, N940, N178);
nor NOR4 (N1475, N1430, N1382, N599, N361);
nor NOR4 (N1476, N1472, N619, N1018, N1072);
not NOT1 (N1477, N1474);
nand NAND2 (N1478, N1473, N1415);
xor XOR2 (N1479, N1459, N1062);
not NOT1 (N1480, N1464);
not NOT1 (N1481, N1475);
buf BUF1 (N1482, N1471);
not NOT1 (N1483, N1482);
not NOT1 (N1484, N1481);
not NOT1 (N1485, N1478);
not NOT1 (N1486, N1461);
nand NAND3 (N1487, N1466, N472, N1417);
buf BUF1 (N1488, N1484);
and AND4 (N1489, N1485, N1167, N559, N1083);
or OR2 (N1490, N1480, N1302);
buf BUF1 (N1491, N1487);
buf BUF1 (N1492, N1491);
not NOT1 (N1493, N1488);
xor XOR2 (N1494, N1463, N1207);
or OR2 (N1495, N1494, N788);
and AND4 (N1496, N1492, N203, N459, N1357);
and AND4 (N1497, N1493, N523, N711, N987);
xor XOR2 (N1498, N1496, N1190);
nor NOR3 (N1499, N1498, N645, N1049);
not NOT1 (N1500, N1477);
xor XOR2 (N1501, N1495, N1139);
nand NAND2 (N1502, N1476, N1302);
xor XOR2 (N1503, N1490, N265);
and AND3 (N1504, N1499, N773, N359);
nor NOR4 (N1505, N1483, N160, N1418, N762);
buf BUF1 (N1506, N1500);
not NOT1 (N1507, N1501);
nor NOR4 (N1508, N1503, N567, N1446, N403);
and AND4 (N1509, N1504, N1299, N133, N592);
nor NOR2 (N1510, N1505, N413);
buf BUF1 (N1511, N1508);
or OR4 (N1512, N1489, N720, N1055, N735);
nor NOR4 (N1513, N1511, N867, N532, N924);
buf BUF1 (N1514, N1497);
and AND3 (N1515, N1507, N944, N1176);
not NOT1 (N1516, N1514);
nor NOR3 (N1517, N1512, N1159, N806);
not NOT1 (N1518, N1513);
nand NAND3 (N1519, N1515, N1040, N586);
not NOT1 (N1520, N1519);
xor XOR2 (N1521, N1510, N757);
and AND3 (N1522, N1517, N994, N464);
buf BUF1 (N1523, N1520);
not NOT1 (N1524, N1521);
and AND3 (N1525, N1506, N1406, N1179);
and AND2 (N1526, N1525, N399);
or OR3 (N1527, N1509, N1342, N454);
or OR4 (N1528, N1479, N349, N1298, N433);
and AND4 (N1529, N1518, N671, N819, N60);
xor XOR2 (N1530, N1528, N383);
and AND4 (N1531, N1527, N637, N1145, N1203);
nor NOR3 (N1532, N1516, N1354, N255);
not NOT1 (N1533, N1502);
nor NOR2 (N1534, N1531, N1366);
nor NOR2 (N1535, N1522, N822);
and AND3 (N1536, N1530, N409, N151);
and AND3 (N1537, N1536, N731, N561);
nor NOR4 (N1538, N1486, N1209, N188, N774);
or OR2 (N1539, N1532, N1006);
and AND2 (N1540, N1537, N209);
or OR3 (N1541, N1540, N77, N133);
and AND3 (N1542, N1533, N1057, N789);
nor NOR2 (N1543, N1529, N1040);
not NOT1 (N1544, N1542);
nand NAND3 (N1545, N1543, N1494, N32);
not NOT1 (N1546, N1544);
nor NOR3 (N1547, N1546, N1361, N291);
xor XOR2 (N1548, N1523, N703);
nand NAND2 (N1549, N1526, N811);
buf BUF1 (N1550, N1541);
not NOT1 (N1551, N1534);
nand NAND4 (N1552, N1538, N773, N1098, N1458);
not NOT1 (N1553, N1545);
buf BUF1 (N1554, N1548);
nand NAND3 (N1555, N1539, N87, N217);
and AND4 (N1556, N1524, N1064, N1058, N57);
and AND3 (N1557, N1550, N1187, N202);
buf BUF1 (N1558, N1557);
not NOT1 (N1559, N1552);
nand NAND3 (N1560, N1559, N967, N1370);
nand NAND3 (N1561, N1558, N1260, N1144);
and AND4 (N1562, N1555, N1522, N166, N176);
or OR2 (N1563, N1562, N19);
and AND4 (N1564, N1535, N1231, N1188, N1248);
not NOT1 (N1565, N1564);
nor NOR2 (N1566, N1549, N1366);
or OR4 (N1567, N1563, N1458, N102, N977);
and AND3 (N1568, N1567, N496, N1183);
or OR3 (N1569, N1568, N1380, N1082);
nor NOR2 (N1570, N1565, N720);
xor XOR2 (N1571, N1553, N386);
nand NAND3 (N1572, N1570, N1491, N121);
buf BUF1 (N1573, N1554);
not NOT1 (N1574, N1556);
or OR3 (N1575, N1551, N157, N800);
and AND4 (N1576, N1561, N1381, N506, N677);
or OR3 (N1577, N1575, N905, N263);
not NOT1 (N1578, N1576);
and AND2 (N1579, N1547, N975);
or OR3 (N1580, N1569, N1461, N1006);
nor NOR3 (N1581, N1578, N405, N1353);
xor XOR2 (N1582, N1577, N976);
nor NOR4 (N1583, N1574, N1161, N1157, N1216);
and AND3 (N1584, N1579, N1144, N717);
buf BUF1 (N1585, N1573);
nor NOR4 (N1586, N1560, N620, N310, N492);
buf BUF1 (N1587, N1584);
buf BUF1 (N1588, N1580);
nand NAND3 (N1589, N1588, N157, N1423);
xor XOR2 (N1590, N1572, N298);
xor XOR2 (N1591, N1587, N55);
not NOT1 (N1592, N1583);
nor NOR3 (N1593, N1589, N321, N266);
xor XOR2 (N1594, N1591, N1349);
xor XOR2 (N1595, N1593, N1212);
nor NOR3 (N1596, N1571, N573, N661);
and AND2 (N1597, N1566, N601);
xor XOR2 (N1598, N1582, N891);
xor XOR2 (N1599, N1590, N1180);
buf BUF1 (N1600, N1581);
not NOT1 (N1601, N1594);
nor NOR2 (N1602, N1585, N209);
and AND2 (N1603, N1601, N569);
buf BUF1 (N1604, N1596);
buf BUF1 (N1605, N1586);
not NOT1 (N1606, N1603);
and AND4 (N1607, N1600, N624, N886, N551);
xor XOR2 (N1608, N1598, N323);
xor XOR2 (N1609, N1599, N454);
nor NOR2 (N1610, N1608, N1374);
nand NAND3 (N1611, N1595, N1433, N205);
nand NAND4 (N1612, N1606, N1450, N1201, N1218);
not NOT1 (N1613, N1604);
or OR2 (N1614, N1602, N625);
not NOT1 (N1615, N1607);
nor NOR3 (N1616, N1597, N441, N328);
or OR4 (N1617, N1610, N1533, N1071, N666);
nor NOR2 (N1618, N1592, N1152);
and AND3 (N1619, N1617, N1430, N224);
nor NOR4 (N1620, N1611, N821, N1041, N1440);
nor NOR4 (N1621, N1609, N1561, N1313, N266);
nand NAND2 (N1622, N1619, N589);
nor NOR4 (N1623, N1613, N1386, N1109, N745);
buf BUF1 (N1624, N1605);
or OR4 (N1625, N1620, N946, N991, N850);
or OR2 (N1626, N1612, N725);
nand NAND2 (N1627, N1626, N488);
nor NOR4 (N1628, N1615, N1223, N198, N404);
and AND4 (N1629, N1621, N152, N201, N236);
not NOT1 (N1630, N1623);
not NOT1 (N1631, N1627);
xor XOR2 (N1632, N1628, N1162);
and AND2 (N1633, N1632, N774);
nor NOR2 (N1634, N1625, N371);
and AND2 (N1635, N1622, N1115);
or OR3 (N1636, N1631, N776, N775);
nand NAND4 (N1637, N1634, N1043, N196, N1630);
or OR4 (N1638, N651, N215, N1399, N754);
nor NOR2 (N1639, N1637, N797);
xor XOR2 (N1640, N1635, N800);
nor NOR2 (N1641, N1640, N504);
xor XOR2 (N1642, N1616, N1509);
not NOT1 (N1643, N1614);
and AND3 (N1644, N1643, N1265, N1554);
nand NAND3 (N1645, N1644, N1245, N1224);
not NOT1 (N1646, N1624);
buf BUF1 (N1647, N1641);
nand NAND2 (N1648, N1645, N427);
and AND3 (N1649, N1646, N1643, N1500);
nand NAND3 (N1650, N1629, N1294, N138);
nand NAND4 (N1651, N1650, N294, N270, N976);
and AND2 (N1652, N1639, N1111);
nand NAND3 (N1653, N1651, N1494, N1132);
xor XOR2 (N1654, N1653, N546);
and AND4 (N1655, N1633, N1176, N1256, N168);
nor NOR3 (N1656, N1649, N468, N1239);
buf BUF1 (N1657, N1636);
and AND4 (N1658, N1655, N729, N1177, N1595);
or OR3 (N1659, N1656, N1105, N235);
buf BUF1 (N1660, N1654);
nor NOR3 (N1661, N1618, N509, N1147);
buf BUF1 (N1662, N1659);
buf BUF1 (N1663, N1652);
buf BUF1 (N1664, N1657);
nand NAND2 (N1665, N1642, N843);
buf BUF1 (N1666, N1647);
buf BUF1 (N1667, N1663);
or OR2 (N1668, N1665, N524);
not NOT1 (N1669, N1660);
nor NOR2 (N1670, N1668, N873);
buf BUF1 (N1671, N1667);
and AND4 (N1672, N1669, N1465, N604, N926);
or OR3 (N1673, N1661, N935, N1382);
buf BUF1 (N1674, N1672);
buf BUF1 (N1675, N1638);
nor NOR2 (N1676, N1664, N489);
buf BUF1 (N1677, N1662);
and AND3 (N1678, N1673, N1508, N1198);
buf BUF1 (N1679, N1676);
or OR4 (N1680, N1666, N1113, N350, N544);
and AND2 (N1681, N1678, N40);
nand NAND4 (N1682, N1677, N278, N71, N885);
xor XOR2 (N1683, N1674, N701);
buf BUF1 (N1684, N1683);
and AND2 (N1685, N1684, N228);
nor NOR4 (N1686, N1675, N542, N1138, N876);
and AND4 (N1687, N1671, N1104, N373, N301);
nand NAND2 (N1688, N1648, N224);
buf BUF1 (N1689, N1686);
and AND3 (N1690, N1688, N1528, N341);
xor XOR2 (N1691, N1670, N1653);
and AND2 (N1692, N1682, N1361);
and AND3 (N1693, N1658, N4, N191);
nand NAND4 (N1694, N1692, N457, N198, N1449);
nand NAND2 (N1695, N1689, N1210);
and AND3 (N1696, N1691, N1062, N510);
and AND3 (N1697, N1685, N1193, N1606);
nand NAND3 (N1698, N1695, N837, N1183);
xor XOR2 (N1699, N1698, N1237);
nand NAND4 (N1700, N1697, N1627, N755, N1129);
and AND3 (N1701, N1696, N301, N580);
not NOT1 (N1702, N1693);
nand NAND4 (N1703, N1702, N738, N234, N184);
nand NAND3 (N1704, N1680, N1138, N1572);
not NOT1 (N1705, N1690);
buf BUF1 (N1706, N1687);
buf BUF1 (N1707, N1681);
or OR2 (N1708, N1700, N142);
xor XOR2 (N1709, N1703, N24);
nand NAND4 (N1710, N1701, N1473, N1690, N56);
nor NOR4 (N1711, N1699, N1106, N606, N854);
buf BUF1 (N1712, N1679);
nor NOR2 (N1713, N1706, N594);
nand NAND2 (N1714, N1709, N33);
buf BUF1 (N1715, N1711);
buf BUF1 (N1716, N1714);
xor XOR2 (N1717, N1716, N906);
xor XOR2 (N1718, N1704, N542);
or OR2 (N1719, N1694, N1333);
or OR2 (N1720, N1715, N1352);
not NOT1 (N1721, N1718);
not NOT1 (N1722, N1713);
nand NAND2 (N1723, N1717, N286);
nand NAND4 (N1724, N1708, N18, N1534, N538);
not NOT1 (N1725, N1723);
and AND3 (N1726, N1719, N127, N877);
nand NAND3 (N1727, N1705, N634, N168);
and AND3 (N1728, N1724, N1264, N1336);
or OR4 (N1729, N1728, N1098, N199, N1724);
or OR4 (N1730, N1712, N604, N532, N1169);
and AND4 (N1731, N1707, N270, N205, N99);
not NOT1 (N1732, N1722);
buf BUF1 (N1733, N1726);
nor NOR2 (N1734, N1727, N8);
buf BUF1 (N1735, N1725);
nand NAND3 (N1736, N1732, N81, N525);
and AND3 (N1737, N1730, N1604, N140);
xor XOR2 (N1738, N1735, N1688);
nor NOR3 (N1739, N1736, N516, N1408);
nand NAND3 (N1740, N1721, N835, N733);
nand NAND4 (N1741, N1729, N387, N1161, N1635);
xor XOR2 (N1742, N1720, N627);
nand NAND2 (N1743, N1710, N1657);
xor XOR2 (N1744, N1742, N756);
and AND3 (N1745, N1733, N1628, N1312);
not NOT1 (N1746, N1737);
nand NAND3 (N1747, N1743, N1742, N1256);
nand NAND4 (N1748, N1739, N1264, N243, N1467);
and AND2 (N1749, N1746, N234);
and AND2 (N1750, N1734, N761);
buf BUF1 (N1751, N1740);
or OR4 (N1752, N1731, N1499, N939, N444);
xor XOR2 (N1753, N1744, N427);
or OR2 (N1754, N1751, N337);
or OR3 (N1755, N1750, N321, N636);
or OR2 (N1756, N1752, N619);
or OR4 (N1757, N1738, N1472, N9, N969);
nand NAND2 (N1758, N1745, N1503);
nand NAND3 (N1759, N1758, N1568, N1060);
not NOT1 (N1760, N1741);
nor NOR2 (N1761, N1760, N1446);
nand NAND2 (N1762, N1753, N1178);
xor XOR2 (N1763, N1756, N323);
xor XOR2 (N1764, N1759, N464);
nand NAND3 (N1765, N1754, N693, N1533);
nor NOR3 (N1766, N1764, N331, N1288);
buf BUF1 (N1767, N1755);
nor NOR3 (N1768, N1765, N1605, N789);
nor NOR3 (N1769, N1749, N1534, N308);
not NOT1 (N1770, N1767);
buf BUF1 (N1771, N1762);
nor NOR4 (N1772, N1757, N737, N537, N1099);
nor NOR2 (N1773, N1771, N717);
and AND2 (N1774, N1768, N1443);
nor NOR2 (N1775, N1761, N424);
xor XOR2 (N1776, N1748, N1548);
xor XOR2 (N1777, N1773, N439);
nand NAND2 (N1778, N1769, N483);
not NOT1 (N1779, N1778);
not NOT1 (N1780, N1766);
xor XOR2 (N1781, N1763, N1587);
nand NAND2 (N1782, N1774, N1617);
nand NAND4 (N1783, N1775, N899, N1213, N960);
xor XOR2 (N1784, N1781, N580);
nor NOR4 (N1785, N1776, N4, N89, N675);
and AND3 (N1786, N1784, N913, N1741);
or OR4 (N1787, N1770, N1719, N387, N1577);
nor NOR3 (N1788, N1783, N931, N516);
xor XOR2 (N1789, N1782, N1489);
and AND3 (N1790, N1785, N1532, N1681);
buf BUF1 (N1791, N1780);
buf BUF1 (N1792, N1789);
buf BUF1 (N1793, N1786);
buf BUF1 (N1794, N1779);
not NOT1 (N1795, N1794);
or OR2 (N1796, N1747, N531);
nand NAND4 (N1797, N1788, N964, N128, N1108);
not NOT1 (N1798, N1792);
xor XOR2 (N1799, N1791, N1497);
not NOT1 (N1800, N1787);
or OR4 (N1801, N1797, N593, N86, N266);
nor NOR2 (N1802, N1772, N1082);
nor NOR4 (N1803, N1801, N1270, N98, N373);
nand NAND4 (N1804, N1795, N643, N469, N217);
not NOT1 (N1805, N1802);
nor NOR3 (N1806, N1777, N944, N1543);
not NOT1 (N1807, N1796);
buf BUF1 (N1808, N1790);
nand NAND2 (N1809, N1800, N1042);
nand NAND4 (N1810, N1808, N1632, N171, N1460);
or OR4 (N1811, N1810, N1218, N472, N116);
and AND2 (N1812, N1807, N797);
xor XOR2 (N1813, N1803, N1675);
and AND2 (N1814, N1804, N1256);
buf BUF1 (N1815, N1814);
xor XOR2 (N1816, N1806, N375);
nor NOR2 (N1817, N1798, N1485);
nand NAND4 (N1818, N1817, N660, N664, N247);
buf BUF1 (N1819, N1816);
nor NOR2 (N1820, N1793, N140);
and AND3 (N1821, N1820, N1026, N1641);
nand NAND3 (N1822, N1818, N1231, N707);
not NOT1 (N1823, N1809);
or OR4 (N1824, N1805, N866, N776, N1063);
nand NAND2 (N1825, N1821, N1773);
nand NAND2 (N1826, N1823, N433);
xor XOR2 (N1827, N1826, N628);
buf BUF1 (N1828, N1813);
nand NAND3 (N1829, N1822, N782, N687);
not NOT1 (N1830, N1827);
and AND4 (N1831, N1830, N530, N864, N77);
xor XOR2 (N1832, N1829, N204);
buf BUF1 (N1833, N1819);
not NOT1 (N1834, N1815);
buf BUF1 (N1835, N1828);
nand NAND2 (N1836, N1811, N401);
nor NOR2 (N1837, N1832, N1095);
xor XOR2 (N1838, N1831, N492);
nand NAND2 (N1839, N1836, N793);
not NOT1 (N1840, N1835);
or OR2 (N1841, N1840, N783);
nor NOR4 (N1842, N1833, N1831, N1446, N111);
nand NAND3 (N1843, N1838, N1026, N370);
buf BUF1 (N1844, N1824);
nor NOR2 (N1845, N1834, N720);
buf BUF1 (N1846, N1839);
or OR2 (N1847, N1843, N1099);
nor NOR4 (N1848, N1844, N49, N698, N624);
nor NOR2 (N1849, N1847, N1481);
not NOT1 (N1850, N1845);
xor XOR2 (N1851, N1825, N825);
xor XOR2 (N1852, N1848, N565);
and AND3 (N1853, N1837, N973, N1256);
nor NOR4 (N1854, N1846, N1122, N1213, N1449);
nand NAND3 (N1855, N1841, N1026, N669);
xor XOR2 (N1856, N1842, N48);
xor XOR2 (N1857, N1849, N190);
nor NOR4 (N1858, N1856, N1819, N250, N1857);
or OR3 (N1859, N355, N703, N1105);
and AND4 (N1860, N1859, N938, N1049, N1755);
nor NOR4 (N1861, N1852, N489, N59, N467);
nor NOR4 (N1862, N1851, N1023, N1316, N1616);
or OR3 (N1863, N1858, N1357, N872);
or OR2 (N1864, N1862, N645);
buf BUF1 (N1865, N1855);
nor NOR4 (N1866, N1854, N1848, N1790, N673);
nor NOR4 (N1867, N1866, N294, N1565, N1655);
or OR2 (N1868, N1812, N747);
xor XOR2 (N1869, N1861, N838);
or OR4 (N1870, N1869, N742, N128, N99);
and AND3 (N1871, N1860, N1581, N596);
nor NOR3 (N1872, N1799, N711, N856);
buf BUF1 (N1873, N1872);
nand NAND4 (N1874, N1865, N298, N1220, N58);
buf BUF1 (N1875, N1853);
nand NAND3 (N1876, N1873, N988, N664);
buf BUF1 (N1877, N1875);
not NOT1 (N1878, N1871);
not NOT1 (N1879, N1863);
nand NAND2 (N1880, N1864, N432);
not NOT1 (N1881, N1874);
and AND2 (N1882, N1870, N220);
and AND3 (N1883, N1879, N1799, N681);
not NOT1 (N1884, N1868);
nand NAND4 (N1885, N1882, N1088, N1221, N646);
not NOT1 (N1886, N1884);
not NOT1 (N1887, N1878);
xor XOR2 (N1888, N1885, N508);
nor NOR4 (N1889, N1876, N1606, N407, N1685);
xor XOR2 (N1890, N1881, N2);
nand NAND2 (N1891, N1880, N1114);
xor XOR2 (N1892, N1867, N840);
buf BUF1 (N1893, N1890);
and AND4 (N1894, N1883, N1068, N798, N78);
xor XOR2 (N1895, N1877, N588);
buf BUF1 (N1896, N1850);
and AND4 (N1897, N1896, N1866, N1438, N63);
nand NAND2 (N1898, N1891, N1432);
or OR4 (N1899, N1894, N737, N1588, N458);
and AND3 (N1900, N1888, N233, N192);
and AND2 (N1901, N1889, N1426);
buf BUF1 (N1902, N1897);
and AND4 (N1903, N1895, N1318, N1135, N546);
xor XOR2 (N1904, N1887, N1058);
or OR3 (N1905, N1893, N1013, N995);
not NOT1 (N1906, N1899);
and AND4 (N1907, N1902, N29, N1517, N1171);
xor XOR2 (N1908, N1886, N1523);
buf BUF1 (N1909, N1905);
buf BUF1 (N1910, N1901);
xor XOR2 (N1911, N1903, N719);
and AND4 (N1912, N1910, N1504, N1801, N989);
and AND2 (N1913, N1904, N1173);
not NOT1 (N1914, N1909);
xor XOR2 (N1915, N1912, N774);
nor NOR4 (N1916, N1906, N619, N1192, N1400);
and AND4 (N1917, N1913, N125, N213, N647);
and AND4 (N1918, N1917, N1651, N192, N392);
xor XOR2 (N1919, N1914, N1186);
not NOT1 (N1920, N1898);
xor XOR2 (N1921, N1916, N819);
buf BUF1 (N1922, N1919);
and AND4 (N1923, N1892, N552, N1613, N1569);
or OR2 (N1924, N1907, N1478);
or OR3 (N1925, N1922, N42, N857);
not NOT1 (N1926, N1908);
xor XOR2 (N1927, N1915, N995);
or OR4 (N1928, N1923, N545, N1128, N1023);
and AND3 (N1929, N1918, N245, N1447);
or OR3 (N1930, N1926, N80, N1320);
buf BUF1 (N1931, N1928);
or OR3 (N1932, N1927, N1083, N699);
and AND4 (N1933, N1921, N857, N1658, N1426);
or OR4 (N1934, N1925, N789, N1918, N1238);
nand NAND3 (N1935, N1931, N1248, N1021);
and AND4 (N1936, N1934, N256, N699, N803);
buf BUF1 (N1937, N1929);
not NOT1 (N1938, N1911);
buf BUF1 (N1939, N1935);
and AND4 (N1940, N1939, N1861, N1238, N163);
or OR3 (N1941, N1933, N1864, N914);
not NOT1 (N1942, N1920);
or OR2 (N1943, N1940, N1148);
buf BUF1 (N1944, N1941);
xor XOR2 (N1945, N1937, N1760);
or OR3 (N1946, N1932, N587, N1199);
xor XOR2 (N1947, N1946, N1548);
nand NAND3 (N1948, N1924, N1238, N10);
nor NOR3 (N1949, N1900, N1664, N983);
and AND2 (N1950, N1944, N596);
nand NAND4 (N1951, N1938, N1716, N168, N901);
or OR4 (N1952, N1947, N1814, N358, N1470);
buf BUF1 (N1953, N1950);
not NOT1 (N1954, N1951);
and AND2 (N1955, N1948, N707);
and AND2 (N1956, N1930, N690);
not NOT1 (N1957, N1956);
xor XOR2 (N1958, N1955, N191);
or OR3 (N1959, N1954, N884, N1464);
not NOT1 (N1960, N1957);
buf BUF1 (N1961, N1936);
xor XOR2 (N1962, N1960, N1218);
or OR2 (N1963, N1949, N943);
xor XOR2 (N1964, N1962, N1373);
nor NOR2 (N1965, N1942, N274);
nand NAND2 (N1966, N1953, N1480);
nor NOR3 (N1967, N1945, N1908, N1845);
and AND4 (N1968, N1966, N902, N843, N1587);
or OR3 (N1969, N1963, N1003, N310);
not NOT1 (N1970, N1965);
xor XOR2 (N1971, N1968, N762);
buf BUF1 (N1972, N1964);
nand NAND4 (N1973, N1967, N722, N1045, N1240);
not NOT1 (N1974, N1961);
xor XOR2 (N1975, N1959, N1767);
or OR2 (N1976, N1975, N1651);
xor XOR2 (N1977, N1973, N365);
buf BUF1 (N1978, N1976);
xor XOR2 (N1979, N1974, N106);
nor NOR4 (N1980, N1971, N460, N535, N1456);
or OR2 (N1981, N1977, N117);
and AND4 (N1982, N1969, N333, N37, N1336);
buf BUF1 (N1983, N1970);
nand NAND3 (N1984, N1972, N698, N37);
not NOT1 (N1985, N1982);
xor XOR2 (N1986, N1952, N1219);
and AND4 (N1987, N1943, N739, N1947, N872);
nand NAND2 (N1988, N1985, N1756);
nor NOR3 (N1989, N1988, N884, N838);
nand NAND4 (N1990, N1989, N1935, N47, N793);
buf BUF1 (N1991, N1981);
xor XOR2 (N1992, N1979, N970);
or OR3 (N1993, N1991, N1917, N1120);
xor XOR2 (N1994, N1980, N349);
buf BUF1 (N1995, N1978);
nor NOR4 (N1996, N1986, N765, N792, N1780);
nand NAND2 (N1997, N1996, N1618);
and AND3 (N1998, N1987, N330, N1290);
nand NAND4 (N1999, N1992, N344, N1253, N663);
xor XOR2 (N2000, N1995, N1396);
buf BUF1 (N2001, N1994);
not NOT1 (N2002, N1997);
not NOT1 (N2003, N1984);
and AND4 (N2004, N1990, N1131, N1773, N1282);
and AND3 (N2005, N2002, N1573, N209);
or OR4 (N2006, N1983, N1065, N1545, N138);
nand NAND2 (N2007, N2003, N1166);
or OR2 (N2008, N2001, N1972);
buf BUF1 (N2009, N1958);
or OR3 (N2010, N2006, N1515, N1132);
or OR4 (N2011, N1999, N1758, N593, N84);
not NOT1 (N2012, N2011);
buf BUF1 (N2013, N2005);
nand NAND4 (N2014, N2013, N1996, N1079, N1951);
and AND2 (N2015, N2004, N1241);
buf BUF1 (N2016, N2015);
buf BUF1 (N2017, N2016);
endmodule