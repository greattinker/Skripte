// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11;

output N85,N92,N106,N110,N108,N109,N101,N98,N102,N111;

nor NOR3 (N12, N6, N10, N1);
not NOT1 (N13, N3);
xor XOR2 (N14, N2, N2);
nor NOR2 (N15, N6, N5);
or OR3 (N16, N13, N11, N6);
or OR2 (N17, N5, N12);
and AND2 (N18, N1, N5);
or OR3 (N19, N1, N7, N3);
xor XOR2 (N20, N1, N7);
nand NAND4 (N21, N16, N9, N14, N4);
xor XOR2 (N22, N2, N6);
nor NOR3 (N23, N5, N20, N9);
buf BUF1 (N24, N20);
nand NAND3 (N25, N24, N5, N14);
buf BUF1 (N26, N11);
not NOT1 (N27, N24);
nand NAND2 (N28, N18, N24);
or OR4 (N29, N21, N24, N18, N11);
nor NOR3 (N30, N27, N25, N16);
nand NAND3 (N31, N13, N26, N28);
not NOT1 (N32, N10);
buf BUF1 (N33, N28);
buf BUF1 (N34, N23);
or OR4 (N35, N31, N22, N29, N32);
not NOT1 (N36, N16);
nand NAND4 (N37, N1, N26, N3, N28);
buf BUF1 (N38, N20);
nor NOR2 (N39, N17, N8);
nor NOR3 (N40, N34, N33, N33);
or OR3 (N41, N19, N19, N1);
not NOT1 (N42, N40);
nor NOR3 (N43, N40, N26, N21);
or OR3 (N44, N30, N34, N12);
buf BUF1 (N45, N43);
or OR4 (N46, N44, N11, N25, N25);
not NOT1 (N47, N42);
buf BUF1 (N48, N46);
nor NOR3 (N49, N45, N25, N47);
nand NAND4 (N50, N38, N23, N5, N1);
or OR3 (N51, N35, N23, N30);
or OR2 (N52, N51, N40);
xor XOR2 (N53, N42, N4);
xor XOR2 (N54, N53, N31);
or OR4 (N55, N48, N11, N29, N51);
not NOT1 (N56, N52);
and AND4 (N57, N41, N52, N23, N39);
not NOT1 (N58, N1);
nand NAND4 (N59, N56, N20, N7, N13);
nor NOR4 (N60, N57, N55, N20, N45);
not NOT1 (N61, N42);
xor XOR2 (N62, N58, N53);
buf BUF1 (N63, N36);
nand NAND2 (N64, N62, N49);
and AND4 (N65, N31, N42, N60, N2);
or OR2 (N66, N27, N23);
or OR3 (N67, N65, N61, N28);
or OR4 (N68, N65, N59, N13, N35);
nor NOR2 (N69, N54, N18);
xor XOR2 (N70, N69, N45);
not NOT1 (N71, N14);
buf BUF1 (N72, N66);
nand NAND2 (N73, N64, N60);
buf BUF1 (N74, N37);
nor NOR2 (N75, N71, N55);
or OR4 (N76, N50, N6, N66, N70);
nand NAND4 (N77, N43, N25, N69, N23);
nand NAND3 (N78, N75, N21, N20);
nand NAND3 (N79, N63, N77, N65);
and AND4 (N80, N63, N70, N19, N14);
nand NAND4 (N81, N78, N63, N52, N10);
nor NOR4 (N82, N67, N5, N81, N11);
or OR2 (N83, N62, N2);
nor NOR2 (N84, N80, N58);
xor XOR2 (N85, N76, N10);
nand NAND2 (N86, N72, N15);
and AND3 (N87, N54, N32, N10);
not NOT1 (N88, N86);
and AND2 (N89, N88, N15);
buf BUF1 (N90, N68);
nor NOR3 (N91, N87, N10, N61);
and AND4 (N92, N84, N23, N52, N75);
buf BUF1 (N93, N82);
buf BUF1 (N94, N89);
buf BUF1 (N95, N90);
nor NOR2 (N96, N91, N34);
or OR4 (N97, N83, N19, N24, N3);
xor XOR2 (N98, N97, N21);
and AND2 (N99, N93, N57);
and AND3 (N100, N73, N17, N91);
or OR4 (N101, N100, N100, N18, N19);
not NOT1 (N102, N95);
nor NOR2 (N103, N79, N90);
xor XOR2 (N104, N103, N68);
nand NAND4 (N105, N104, N42, N43, N8);
nand NAND4 (N106, N74, N67, N7, N54);
or OR4 (N107, N96, N97, N48, N50);
xor XOR2 (N108, N94, N68);
buf BUF1 (N109, N107);
not NOT1 (N110, N105);
and AND3 (N111, N99, N45, N74);
endmodule