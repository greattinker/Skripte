// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17;

output N708,N700,N704,N713,N702,N716,N701,N715,N709,N717;

nor NOR2 (N18, N5, N7);
xor XOR2 (N19, N10, N5);
and AND3 (N20, N13, N12, N6);
buf BUF1 (N21, N17);
or OR2 (N22, N7, N11);
xor XOR2 (N23, N1, N2);
or OR3 (N24, N18, N23, N14);
or OR4 (N25, N19, N19, N22, N23);
xor XOR2 (N26, N21, N10);
buf BUF1 (N27, N22);
or OR4 (N28, N16, N19, N3, N3);
nand NAND2 (N29, N8, N24);
nand NAND3 (N30, N11, N20, N23);
and AND2 (N31, N25, N7);
and AND4 (N32, N19, N29, N28, N1);
or OR2 (N33, N24, N4);
not NOT1 (N34, N21);
xor XOR2 (N35, N8, N3);
xor XOR2 (N36, N13, N4);
xor XOR2 (N37, N10, N17);
xor XOR2 (N38, N34, N35);
buf BUF1 (N39, N31);
xor XOR2 (N40, N12, N22);
nor NOR4 (N41, N26, N5, N32, N14);
buf BUF1 (N42, N39);
nor NOR3 (N43, N33, N10, N29);
or OR3 (N44, N43, N13, N40);
or OR3 (N45, N4, N9, N25);
not NOT1 (N46, N23);
nor NOR4 (N47, N46, N11, N37, N3);
buf BUF1 (N48, N7);
buf BUF1 (N49, N27);
not NOT1 (N50, N38);
xor XOR2 (N51, N44, N5);
buf BUF1 (N52, N48);
nor NOR2 (N53, N30, N46);
nand NAND4 (N54, N50, N1, N33, N38);
nand NAND3 (N55, N36, N3, N54);
nor NOR4 (N56, N18, N20, N44, N28);
xor XOR2 (N57, N45, N55);
nand NAND2 (N58, N19, N7);
xor XOR2 (N59, N41, N54);
nand NAND3 (N60, N52, N50, N3);
not NOT1 (N61, N57);
and AND4 (N62, N56, N12, N52, N49);
nor NOR4 (N63, N37, N40, N20, N11);
buf BUF1 (N64, N62);
nor NOR2 (N65, N53, N41);
nand NAND4 (N66, N63, N20, N6, N5);
and AND3 (N67, N51, N32, N45);
nand NAND2 (N68, N61, N60);
nand NAND2 (N69, N21, N26);
nand NAND3 (N70, N65, N63, N19);
and AND2 (N71, N64, N56);
and AND2 (N72, N70, N64);
not NOT1 (N73, N68);
xor XOR2 (N74, N69, N18);
or OR4 (N75, N59, N29, N45, N33);
and AND3 (N76, N66, N26, N22);
nand NAND3 (N77, N58, N30, N71);
not NOT1 (N78, N70);
nor NOR4 (N79, N78, N53, N20, N49);
xor XOR2 (N80, N73, N50);
and AND2 (N81, N76, N13);
and AND4 (N82, N47, N57, N5, N36);
or OR3 (N83, N67, N48, N29);
and AND4 (N84, N77, N12, N35, N44);
nor NOR3 (N85, N82, N32, N12);
nand NAND2 (N86, N83, N75);
nor NOR3 (N87, N18, N34, N73);
nand NAND2 (N88, N87, N72);
nand NAND3 (N89, N25, N61, N31);
buf BUF1 (N90, N84);
or OR3 (N91, N90, N58, N58);
not NOT1 (N92, N89);
buf BUF1 (N93, N88);
xor XOR2 (N94, N86, N29);
buf BUF1 (N95, N80);
buf BUF1 (N96, N79);
nor NOR2 (N97, N95, N8);
nor NOR4 (N98, N92, N44, N75, N14);
nand NAND3 (N99, N81, N21, N40);
or OR2 (N100, N97, N75);
xor XOR2 (N101, N42, N44);
and AND4 (N102, N100, N85, N54, N96);
xor XOR2 (N103, N72, N73);
nand NAND3 (N104, N99, N98, N19);
or OR4 (N105, N61, N19, N18, N60);
nor NOR4 (N106, N42, N32, N28, N49);
buf BUF1 (N107, N103);
buf BUF1 (N108, N91);
or OR2 (N109, N107, N87);
nor NOR2 (N110, N109, N41);
xor XOR2 (N111, N101, N104);
xor XOR2 (N112, N103, N97);
buf BUF1 (N113, N111);
xor XOR2 (N114, N106, N37);
or OR3 (N115, N112, N69, N50);
and AND4 (N116, N94, N115, N25, N97);
not NOT1 (N117, N64);
or OR3 (N118, N116, N13, N106);
buf BUF1 (N119, N110);
nor NOR2 (N120, N74, N83);
not NOT1 (N121, N108);
or OR4 (N122, N120, N59, N34, N17);
and AND4 (N123, N93, N43, N16, N54);
nor NOR3 (N124, N117, N10, N33);
buf BUF1 (N125, N124);
or OR3 (N126, N119, N101, N49);
or OR3 (N127, N121, N63, N30);
nand NAND2 (N128, N123, N121);
not NOT1 (N129, N102);
and AND3 (N130, N114, N19, N16);
xor XOR2 (N131, N125, N116);
nor NOR3 (N132, N113, N35, N108);
and AND3 (N133, N105, N13, N78);
nor NOR4 (N134, N129, N16, N89, N70);
xor XOR2 (N135, N127, N10);
nand NAND2 (N136, N122, N54);
nand NAND4 (N137, N135, N20, N83, N11);
buf BUF1 (N138, N133);
xor XOR2 (N139, N126, N26);
nor NOR4 (N140, N132, N28, N87, N18);
nor NOR2 (N141, N130, N115);
or OR2 (N142, N138, N25);
and AND2 (N143, N118, N33);
nor NOR4 (N144, N131, N19, N136, N128);
not NOT1 (N145, N123);
xor XOR2 (N146, N96, N20);
or OR2 (N147, N145, N3);
not NOT1 (N148, N139);
nand NAND4 (N149, N144, N104, N148, N79);
or OR4 (N150, N25, N119, N24, N143);
nand NAND3 (N151, N38, N117, N51);
and AND2 (N152, N150, N30);
nor NOR4 (N153, N147, N110, N114, N47);
xor XOR2 (N154, N152, N98);
or OR2 (N155, N142, N72);
or OR3 (N156, N155, N135, N76);
not NOT1 (N157, N154);
xor XOR2 (N158, N156, N120);
or OR2 (N159, N151, N129);
not NOT1 (N160, N137);
nand NAND3 (N161, N146, N5, N89);
buf BUF1 (N162, N158);
or OR2 (N163, N159, N79);
and AND2 (N164, N163, N38);
and AND4 (N165, N161, N9, N78, N4);
or OR4 (N166, N164, N40, N127, N70);
not NOT1 (N167, N165);
nor NOR2 (N168, N141, N140);
xor XOR2 (N169, N142, N21);
or OR4 (N170, N153, N82, N6, N118);
nand NAND2 (N171, N149, N11);
buf BUF1 (N172, N170);
nand NAND2 (N173, N166, N95);
buf BUF1 (N174, N169);
and AND2 (N175, N173, N2);
or OR4 (N176, N174, N12, N87, N121);
not NOT1 (N177, N157);
nand NAND3 (N178, N172, N3, N82);
buf BUF1 (N179, N162);
not NOT1 (N180, N171);
or OR4 (N181, N167, N169, N178, N95);
and AND4 (N182, N124, N103, N75, N148);
not NOT1 (N183, N182);
nand NAND3 (N184, N180, N53, N25);
nor NOR2 (N185, N175, N41);
buf BUF1 (N186, N185);
nand NAND2 (N187, N134, N16);
buf BUF1 (N188, N168);
nand NAND3 (N189, N184, N78, N26);
or OR3 (N190, N186, N116, N22);
not NOT1 (N191, N177);
xor XOR2 (N192, N179, N86);
and AND3 (N193, N183, N116, N127);
nand NAND4 (N194, N181, N20, N49, N93);
nor NOR4 (N195, N190, N129, N157, N57);
buf BUF1 (N196, N195);
nand NAND2 (N197, N189, N129);
and AND2 (N198, N193, N33);
buf BUF1 (N199, N194);
xor XOR2 (N200, N199, N19);
nand NAND3 (N201, N187, N30, N131);
buf BUF1 (N202, N192);
and AND4 (N203, N198, N13, N181, N29);
not NOT1 (N204, N202);
buf BUF1 (N205, N191);
nand NAND4 (N206, N205, N154, N117, N135);
and AND4 (N207, N197, N124, N187, N8);
nand NAND3 (N208, N176, N202, N63);
or OR4 (N209, N204, N48, N75, N10);
and AND3 (N210, N203, N116, N60);
nor NOR3 (N211, N210, N178, N187);
and AND3 (N212, N196, N116, N84);
buf BUF1 (N213, N160);
nor NOR4 (N214, N211, N53, N128, N122);
or OR3 (N215, N212, N60, N100);
and AND2 (N216, N188, N48);
nand NAND3 (N217, N206, N147, N129);
not NOT1 (N218, N216);
or OR2 (N219, N214, N46);
or OR2 (N220, N215, N21);
and AND4 (N221, N219, N47, N190, N39);
and AND3 (N222, N217, N131, N221);
not NOT1 (N223, N145);
buf BUF1 (N224, N208);
or OR3 (N225, N223, N151, N20);
buf BUF1 (N226, N201);
or OR3 (N227, N209, N49, N219);
xor XOR2 (N228, N222, N169);
not NOT1 (N229, N227);
and AND2 (N230, N225, N95);
buf BUF1 (N231, N207);
or OR4 (N232, N218, N115, N216, N34);
nand NAND2 (N233, N226, N175);
nand NAND3 (N234, N200, N104, N120);
or OR4 (N235, N213, N98, N221, N61);
buf BUF1 (N236, N228);
nand NAND2 (N237, N224, N210);
nand NAND2 (N238, N229, N70);
not NOT1 (N239, N238);
nor NOR4 (N240, N230, N42, N139, N191);
nor NOR4 (N241, N235, N187, N236, N46);
and AND3 (N242, N178, N154, N11);
or OR3 (N243, N220, N60, N45);
or OR3 (N244, N240, N170, N220);
and AND2 (N245, N243, N100);
or OR4 (N246, N233, N11, N227, N67);
xor XOR2 (N247, N246, N196);
nor NOR3 (N248, N244, N16, N187);
buf BUF1 (N249, N247);
nor NOR2 (N250, N231, N239);
and AND4 (N251, N124, N93, N149, N178);
xor XOR2 (N252, N234, N23);
nor NOR2 (N253, N245, N95);
and AND4 (N254, N253, N66, N246, N32);
not NOT1 (N255, N241);
nor NOR4 (N256, N251, N250, N196, N220);
nor NOR2 (N257, N140, N20);
xor XOR2 (N258, N249, N214);
and AND4 (N259, N232, N89, N139, N182);
nor NOR2 (N260, N258, N196);
not NOT1 (N261, N260);
xor XOR2 (N262, N242, N205);
or OR2 (N263, N237, N124);
buf BUF1 (N264, N254);
not NOT1 (N265, N257);
not NOT1 (N266, N263);
xor XOR2 (N267, N252, N242);
or OR2 (N268, N255, N45);
buf BUF1 (N269, N264);
xor XOR2 (N270, N256, N123);
buf BUF1 (N271, N270);
nand NAND4 (N272, N259, N176, N32, N145);
or OR3 (N273, N268, N92, N100);
and AND3 (N274, N248, N99, N10);
or OR3 (N275, N261, N164, N148);
nand NAND3 (N276, N272, N272, N167);
nand NAND2 (N277, N273, N224);
and AND2 (N278, N266, N263);
nor NOR2 (N279, N276, N90);
nor NOR2 (N280, N274, N194);
and AND2 (N281, N277, N54);
not NOT1 (N282, N281);
and AND4 (N283, N279, N48, N147, N150);
xor XOR2 (N284, N271, N147);
or OR4 (N285, N267, N257, N21, N94);
nand NAND3 (N286, N275, N121, N77);
or OR4 (N287, N285, N36, N137, N184);
nor NOR3 (N288, N262, N4, N186);
nand NAND4 (N289, N269, N233, N221, N71);
not NOT1 (N290, N288);
not NOT1 (N291, N284);
buf BUF1 (N292, N283);
buf BUF1 (N293, N286);
xor XOR2 (N294, N290, N68);
buf BUF1 (N295, N280);
and AND2 (N296, N265, N47);
not NOT1 (N297, N296);
nor NOR3 (N298, N278, N126, N49);
or OR4 (N299, N287, N34, N225, N37);
nand NAND4 (N300, N299, N58, N12, N1);
not NOT1 (N301, N297);
and AND4 (N302, N289, N214, N116, N155);
or OR2 (N303, N282, N284);
nor NOR2 (N304, N303, N219);
buf BUF1 (N305, N298);
nand NAND4 (N306, N292, N76, N56, N2);
buf BUF1 (N307, N293);
not NOT1 (N308, N307);
or OR4 (N309, N306, N15, N184, N55);
or OR2 (N310, N294, N245);
xor XOR2 (N311, N295, N46);
nand NAND3 (N312, N308, N171, N148);
buf BUF1 (N313, N291);
or OR2 (N314, N300, N18);
or OR3 (N315, N314, N58, N158);
nand NAND3 (N316, N311, N263, N185);
xor XOR2 (N317, N302, N309);
xor XOR2 (N318, N217, N89);
nand NAND4 (N319, N316, N208, N289, N15);
not NOT1 (N320, N319);
nor NOR2 (N321, N310, N11);
buf BUF1 (N322, N321);
or OR2 (N323, N312, N4);
buf BUF1 (N324, N304);
or OR2 (N325, N323, N148);
nor NOR2 (N326, N320, N132);
and AND2 (N327, N305, N186);
and AND2 (N328, N313, N54);
not NOT1 (N329, N322);
xor XOR2 (N330, N317, N326);
nand NAND2 (N331, N88, N330);
and AND2 (N332, N138, N70);
nor NOR4 (N333, N332, N90, N297, N138);
nand NAND3 (N334, N328, N258, N48);
buf BUF1 (N335, N327);
xor XOR2 (N336, N325, N300);
and AND4 (N337, N324, N229, N333, N160);
nor NOR4 (N338, N186, N335, N223, N112);
and AND3 (N339, N5, N242, N251);
xor XOR2 (N340, N334, N268);
nand NAND2 (N341, N337, N160);
nand NAND4 (N342, N331, N254, N128, N77);
and AND3 (N343, N315, N264, N30);
or OR4 (N344, N339, N258, N13, N309);
buf BUF1 (N345, N336);
nor NOR3 (N346, N301, N324, N190);
nor NOR3 (N347, N341, N209, N213);
and AND2 (N348, N340, N171);
and AND4 (N349, N348, N206, N80, N184);
xor XOR2 (N350, N347, N46);
or OR4 (N351, N345, N283, N301, N49);
buf BUF1 (N352, N344);
nor NOR2 (N353, N338, N174);
xor XOR2 (N354, N352, N181);
not NOT1 (N355, N351);
nor NOR4 (N356, N343, N141, N19, N153);
nand NAND2 (N357, N355, N121);
nor NOR3 (N358, N350, N171, N272);
or OR3 (N359, N357, N308, N289);
xor XOR2 (N360, N358, N145);
xor XOR2 (N361, N329, N347);
nand NAND4 (N362, N349, N233, N222, N292);
xor XOR2 (N363, N362, N163);
not NOT1 (N364, N361);
buf BUF1 (N365, N342);
and AND2 (N366, N353, N35);
not NOT1 (N367, N346);
buf BUF1 (N368, N354);
and AND2 (N369, N366, N305);
buf BUF1 (N370, N356);
and AND3 (N371, N365, N349, N109);
nor NOR2 (N372, N360, N61);
nand NAND3 (N373, N359, N202, N114);
buf BUF1 (N374, N363);
buf BUF1 (N375, N318);
and AND3 (N376, N368, N163, N180);
nor NOR4 (N377, N369, N69, N49, N111);
or OR3 (N378, N373, N104, N376);
nand NAND4 (N379, N59, N356, N120, N213);
or OR3 (N380, N372, N96, N289);
nand NAND2 (N381, N374, N41);
buf BUF1 (N382, N378);
buf BUF1 (N383, N375);
nand NAND3 (N384, N381, N343, N353);
xor XOR2 (N385, N379, N171);
nand NAND4 (N386, N371, N127, N172, N44);
not NOT1 (N387, N384);
buf BUF1 (N388, N367);
buf BUF1 (N389, N385);
nor NOR4 (N390, N388, N127, N49, N290);
not NOT1 (N391, N364);
and AND3 (N392, N377, N248, N134);
or OR3 (N393, N382, N369, N46);
not NOT1 (N394, N370);
buf BUF1 (N395, N383);
not NOT1 (N396, N395);
xor XOR2 (N397, N391, N334);
nor NOR2 (N398, N386, N342);
and AND2 (N399, N397, N121);
nor NOR3 (N400, N387, N78, N68);
not NOT1 (N401, N399);
and AND2 (N402, N394, N93);
xor XOR2 (N403, N393, N76);
buf BUF1 (N404, N398);
and AND3 (N405, N392, N339, N306);
nor NOR4 (N406, N403, N362, N301, N142);
nand NAND3 (N407, N380, N243, N46);
nand NAND2 (N408, N396, N293);
and AND4 (N409, N389, N197, N204, N79);
not NOT1 (N410, N405);
and AND3 (N411, N401, N380, N253);
nor NOR4 (N412, N406, N407, N180, N190);
xor XOR2 (N413, N212, N262);
nand NAND2 (N414, N390, N305);
nand NAND4 (N415, N408, N241, N12, N289);
buf BUF1 (N416, N411);
not NOT1 (N417, N415);
buf BUF1 (N418, N402);
nor NOR3 (N419, N404, N34, N346);
nand NAND4 (N420, N417, N37, N3, N203);
buf BUF1 (N421, N409);
nor NOR2 (N422, N410, N39);
nor NOR3 (N423, N419, N234, N397);
nand NAND3 (N424, N418, N44, N318);
or OR4 (N425, N420, N349, N78, N311);
or OR2 (N426, N400, N323);
not NOT1 (N427, N414);
buf BUF1 (N428, N425);
or OR3 (N429, N423, N92, N364);
and AND2 (N430, N428, N363);
nand NAND3 (N431, N424, N268, N294);
nor NOR2 (N432, N416, N13);
xor XOR2 (N433, N427, N123);
not NOT1 (N434, N421);
buf BUF1 (N435, N412);
buf BUF1 (N436, N435);
xor XOR2 (N437, N431, N60);
or OR4 (N438, N434, N68, N144, N281);
and AND3 (N439, N433, N350, N109);
and AND3 (N440, N436, N136, N339);
xor XOR2 (N441, N439, N247);
or OR3 (N442, N430, N333, N79);
nor NOR3 (N443, N426, N421, N379);
not NOT1 (N444, N429);
not NOT1 (N445, N444);
and AND4 (N446, N422, N245, N155, N259);
not NOT1 (N447, N443);
nand NAND3 (N448, N440, N224, N376);
not NOT1 (N449, N432);
not NOT1 (N450, N449);
xor XOR2 (N451, N445, N324);
and AND3 (N452, N441, N36, N285);
nand NAND2 (N453, N448, N43);
or OR3 (N454, N413, N55, N181);
nor NOR3 (N455, N452, N289, N209);
not NOT1 (N456, N454);
not NOT1 (N457, N446);
xor XOR2 (N458, N453, N406);
or OR2 (N459, N456, N59);
not NOT1 (N460, N451);
or OR4 (N461, N457, N39, N120, N191);
nor NOR3 (N462, N460, N126, N244);
xor XOR2 (N463, N461, N277);
buf BUF1 (N464, N462);
nand NAND3 (N465, N437, N315, N85);
not NOT1 (N466, N463);
nand NAND3 (N467, N464, N356, N107);
buf BUF1 (N468, N459);
nor NOR2 (N469, N468, N63);
nand NAND4 (N470, N442, N79, N109, N3);
nor NOR2 (N471, N470, N370);
xor XOR2 (N472, N450, N362);
nor NOR4 (N473, N472, N215, N425, N30);
and AND2 (N474, N458, N252);
buf BUF1 (N475, N447);
buf BUF1 (N476, N469);
nor NOR2 (N477, N465, N119);
and AND3 (N478, N466, N372, N347);
xor XOR2 (N479, N476, N96);
not NOT1 (N480, N479);
or OR3 (N481, N480, N354, N45);
nor NOR4 (N482, N473, N363, N461, N334);
xor XOR2 (N483, N475, N163);
nor NOR2 (N484, N477, N363);
xor XOR2 (N485, N471, N235);
not NOT1 (N486, N455);
buf BUF1 (N487, N484);
or OR3 (N488, N483, N165, N337);
nand NAND2 (N489, N482, N387);
or OR4 (N490, N438, N18, N360, N175);
not NOT1 (N491, N490);
not NOT1 (N492, N474);
buf BUF1 (N493, N485);
nor NOR2 (N494, N487, N449);
nand NAND3 (N495, N494, N78, N309);
xor XOR2 (N496, N489, N237);
xor XOR2 (N497, N491, N264);
nor NOR3 (N498, N492, N472, N243);
or OR3 (N499, N481, N147, N64);
and AND3 (N500, N497, N49, N199);
and AND2 (N501, N499, N358);
nor NOR3 (N502, N498, N491, N293);
buf BUF1 (N503, N478);
or OR4 (N504, N503, N66, N154, N143);
not NOT1 (N505, N496);
xor XOR2 (N506, N505, N276);
or OR2 (N507, N488, N328);
not NOT1 (N508, N506);
nor NOR3 (N509, N504, N63, N38);
xor XOR2 (N510, N509, N131);
nand NAND3 (N511, N502, N171, N355);
nor NOR4 (N512, N486, N299, N79, N390);
buf BUF1 (N513, N507);
or OR2 (N514, N510, N358);
nor NOR4 (N515, N467, N454, N223, N11);
not NOT1 (N516, N512);
not NOT1 (N517, N493);
nor NOR2 (N518, N501, N72);
nand NAND3 (N519, N513, N466, N59);
or OR3 (N520, N518, N130, N127);
xor XOR2 (N521, N495, N475);
nand NAND4 (N522, N521, N466, N303, N110);
xor XOR2 (N523, N517, N249);
nor NOR3 (N524, N511, N226, N391);
not NOT1 (N525, N514);
buf BUF1 (N526, N525);
not NOT1 (N527, N526);
xor XOR2 (N528, N500, N496);
nor NOR2 (N529, N515, N497);
nor NOR2 (N530, N524, N339);
nor NOR3 (N531, N529, N135, N392);
xor XOR2 (N532, N516, N266);
xor XOR2 (N533, N520, N366);
nand NAND2 (N534, N527, N317);
or OR2 (N535, N522, N56);
buf BUF1 (N536, N533);
and AND4 (N537, N519, N239, N484, N210);
buf BUF1 (N538, N535);
buf BUF1 (N539, N531);
nor NOR2 (N540, N537, N241);
not NOT1 (N541, N534);
not NOT1 (N542, N523);
not NOT1 (N543, N532);
nand NAND2 (N544, N508, N184);
nand NAND3 (N545, N540, N368, N351);
or OR2 (N546, N541, N27);
nor NOR2 (N547, N542, N99);
buf BUF1 (N548, N546);
and AND3 (N549, N538, N375, N320);
buf BUF1 (N550, N536);
or OR3 (N551, N544, N454, N185);
and AND4 (N552, N548, N36, N349, N115);
xor XOR2 (N553, N547, N527);
not NOT1 (N554, N530);
nand NAND3 (N555, N554, N173, N190);
nor NOR2 (N556, N539, N165);
not NOT1 (N557, N543);
nor NOR3 (N558, N550, N360, N238);
nand NAND4 (N559, N552, N235, N143, N543);
or OR4 (N560, N553, N295, N40, N48);
not NOT1 (N561, N528);
nand NAND4 (N562, N551, N296, N325, N451);
or OR3 (N563, N555, N222, N543);
or OR3 (N564, N559, N506, N520);
not NOT1 (N565, N545);
not NOT1 (N566, N562);
or OR4 (N567, N566, N320, N555, N138);
or OR3 (N568, N565, N452, N162);
nand NAND2 (N569, N549, N194);
nand NAND3 (N570, N563, N129, N385);
buf BUF1 (N571, N567);
buf BUF1 (N572, N556);
buf BUF1 (N573, N558);
not NOT1 (N574, N561);
not NOT1 (N575, N569);
buf BUF1 (N576, N564);
and AND4 (N577, N574, N476, N322, N403);
xor XOR2 (N578, N576, N83);
xor XOR2 (N579, N557, N328);
and AND3 (N580, N568, N228, N116);
not NOT1 (N581, N570);
not NOT1 (N582, N577);
xor XOR2 (N583, N580, N324);
xor XOR2 (N584, N572, N143);
or OR4 (N585, N575, N473, N328, N395);
and AND3 (N586, N573, N536, N242);
xor XOR2 (N587, N583, N396);
or OR3 (N588, N578, N473, N407);
not NOT1 (N589, N585);
or OR4 (N590, N588, N181, N499, N351);
nand NAND4 (N591, N579, N504, N100, N30);
xor XOR2 (N592, N581, N397);
or OR2 (N593, N571, N210);
xor XOR2 (N594, N591, N34);
xor XOR2 (N595, N594, N294);
xor XOR2 (N596, N589, N592);
or OR2 (N597, N262, N221);
nand NAND3 (N598, N597, N242, N373);
not NOT1 (N599, N598);
buf BUF1 (N600, N584);
buf BUF1 (N601, N587);
buf BUF1 (N602, N599);
and AND2 (N603, N602, N104);
nand NAND4 (N604, N586, N132, N329, N41);
xor XOR2 (N605, N596, N560);
or OR4 (N606, N22, N81, N47, N511);
and AND3 (N607, N603, N384, N390);
xor XOR2 (N608, N582, N483);
nor NOR2 (N609, N600, N535);
or OR4 (N610, N601, N19, N149, N239);
nor NOR2 (N611, N610, N280);
or OR3 (N612, N595, N191, N511);
nor NOR2 (N613, N612, N30);
xor XOR2 (N614, N607, N426);
xor XOR2 (N615, N606, N452);
not NOT1 (N616, N614);
and AND3 (N617, N613, N366, N117);
nor NOR4 (N618, N605, N462, N116, N153);
buf BUF1 (N619, N593);
nor NOR3 (N620, N617, N115, N264);
nor NOR2 (N621, N615, N345);
nand NAND2 (N622, N608, N513);
nand NAND3 (N623, N621, N246, N266);
nand NAND3 (N624, N619, N52, N447);
xor XOR2 (N625, N618, N435);
buf BUF1 (N626, N622);
buf BUF1 (N627, N626);
nand NAND2 (N628, N627, N446);
buf BUF1 (N629, N624);
not NOT1 (N630, N629);
and AND4 (N631, N609, N335, N518, N215);
xor XOR2 (N632, N628, N82);
or OR4 (N633, N620, N541, N80, N503);
nand NAND2 (N634, N611, N411);
not NOT1 (N635, N604);
nand NAND2 (N636, N630, N522);
xor XOR2 (N637, N634, N69);
and AND4 (N638, N633, N213, N149, N256);
buf BUF1 (N639, N625);
nand NAND3 (N640, N632, N263, N580);
nand NAND2 (N641, N616, N437);
or OR3 (N642, N639, N602, N257);
and AND2 (N643, N637, N234);
xor XOR2 (N644, N638, N486);
and AND4 (N645, N644, N73, N167, N302);
not NOT1 (N646, N623);
nand NAND4 (N647, N642, N117, N637, N28);
buf BUF1 (N648, N636);
nand NAND3 (N649, N640, N241, N180);
not NOT1 (N650, N649);
nor NOR2 (N651, N647, N624);
not NOT1 (N652, N651);
nor NOR2 (N653, N635, N563);
xor XOR2 (N654, N631, N650);
nor NOR2 (N655, N432, N468);
nor NOR3 (N656, N648, N336, N533);
nand NAND4 (N657, N653, N91, N621, N75);
not NOT1 (N658, N655);
nand NAND2 (N659, N646, N561);
nand NAND3 (N660, N654, N7, N73);
buf BUF1 (N661, N656);
nand NAND2 (N662, N657, N235);
nor NOR3 (N663, N645, N36, N320);
not NOT1 (N664, N663);
nor NOR4 (N665, N658, N60, N237, N14);
or OR3 (N666, N652, N132, N184);
and AND3 (N667, N659, N188, N121);
and AND2 (N668, N666, N205);
buf BUF1 (N669, N664);
nand NAND2 (N670, N590, N545);
nor NOR4 (N671, N641, N613, N641, N549);
not NOT1 (N672, N669);
not NOT1 (N673, N661);
or OR2 (N674, N665, N659);
not NOT1 (N675, N660);
xor XOR2 (N676, N643, N529);
nand NAND4 (N677, N673, N386, N327, N450);
nor NOR3 (N678, N675, N381, N441);
or OR4 (N679, N676, N41, N536, N253);
nand NAND3 (N680, N679, N535, N587);
not NOT1 (N681, N674);
nand NAND2 (N682, N672, N591);
buf BUF1 (N683, N667);
buf BUF1 (N684, N678);
and AND2 (N685, N670, N188);
and AND2 (N686, N662, N311);
nand NAND3 (N687, N682, N385, N595);
xor XOR2 (N688, N683, N417);
xor XOR2 (N689, N680, N440);
and AND2 (N690, N681, N616);
not NOT1 (N691, N668);
or OR2 (N692, N688, N363);
and AND3 (N693, N686, N163, N154);
buf BUF1 (N694, N690);
and AND3 (N695, N691, N536, N246);
or OR3 (N696, N684, N666, N418);
nand NAND3 (N697, N693, N590, N533);
nor NOR2 (N698, N694, N351);
nor NOR3 (N699, N695, N401, N241);
nor NOR3 (N700, N699, N349, N169);
xor XOR2 (N701, N671, N119);
and AND3 (N702, N697, N131, N518);
xor XOR2 (N703, N698, N606);
buf BUF1 (N704, N689);
nand NAND2 (N705, N685, N598);
nor NOR2 (N706, N696, N699);
or OR4 (N707, N706, N134, N326, N255);
nand NAND3 (N708, N705, N42, N705);
not NOT1 (N709, N703);
and AND4 (N710, N692, N153, N384, N136);
xor XOR2 (N711, N677, N164);
or OR3 (N712, N711, N79, N566);
xor XOR2 (N713, N707, N124);
not NOT1 (N714, N710);
nand NAND2 (N715, N712, N30);
xor XOR2 (N716, N714, N278);
xor XOR2 (N717, N687, N79);
endmodule