// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21;

output N1015,N1019,N1013,N1017,N1009,N1016,N988,N1014,N1020,N1021;

nor NOR2 (N22, N18, N18);
and AND2 (N23, N13, N21);
xor XOR2 (N24, N6, N1);
or OR2 (N25, N11, N4);
nor NOR3 (N26, N7, N23, N7);
not NOT1 (N27, N14);
and AND2 (N28, N22, N1);
nand NAND2 (N29, N25, N25);
xor XOR2 (N30, N11, N10);
buf BUF1 (N31, N24);
nand NAND2 (N32, N19, N30);
and AND3 (N33, N25, N10, N20);
not NOT1 (N34, N31);
and AND3 (N35, N29, N10, N6);
nand NAND2 (N36, N31, N6);
or OR2 (N37, N14, N17);
xor XOR2 (N38, N19, N34);
not NOT1 (N39, N23);
or OR4 (N40, N35, N18, N18, N3);
and AND2 (N41, N40, N27);
xor XOR2 (N42, N28, N35);
nand NAND3 (N43, N15, N15, N22);
and AND3 (N44, N32, N24, N41);
buf BUF1 (N45, N37);
nor NOR3 (N46, N37, N21, N12);
not NOT1 (N47, N39);
or OR4 (N48, N26, N27, N43, N19);
buf BUF1 (N49, N18);
nand NAND2 (N50, N48, N38);
and AND3 (N51, N41, N26, N24);
buf BUF1 (N52, N42);
buf BUF1 (N53, N36);
buf BUF1 (N54, N52);
xor XOR2 (N55, N51, N54);
buf BUF1 (N56, N49);
nand NAND4 (N57, N32, N46, N29, N33);
nor NOR2 (N58, N47, N27);
buf BUF1 (N59, N7);
nand NAND4 (N60, N51, N30, N49, N29);
or OR3 (N61, N56, N17, N34);
or OR3 (N62, N55, N40, N41);
or OR3 (N63, N61, N53, N15);
buf BUF1 (N64, N30);
and AND2 (N65, N63, N40);
nand NAND2 (N66, N44, N60);
nor NOR4 (N67, N23, N10, N7, N55);
and AND3 (N68, N64, N66, N31);
buf BUF1 (N69, N51);
and AND2 (N70, N58, N42);
not NOT1 (N71, N70);
or OR4 (N72, N59, N23, N17, N17);
and AND2 (N73, N50, N42);
and AND2 (N74, N57, N29);
and AND4 (N75, N65, N70, N32, N15);
nor NOR3 (N76, N71, N34, N2);
buf BUF1 (N77, N72);
and AND3 (N78, N75, N4, N6);
and AND4 (N79, N45, N15, N43, N18);
and AND2 (N80, N62, N56);
or OR4 (N81, N78, N54, N53, N11);
buf BUF1 (N82, N80);
nand NAND4 (N83, N73, N59, N27, N30);
buf BUF1 (N84, N74);
and AND3 (N85, N68, N46, N38);
xor XOR2 (N86, N84, N26);
nand NAND3 (N87, N86, N45, N33);
not NOT1 (N88, N81);
not NOT1 (N89, N85);
and AND3 (N90, N67, N8, N36);
nor NOR4 (N91, N88, N30, N40, N38);
xor XOR2 (N92, N83, N26);
and AND2 (N93, N87, N73);
and AND3 (N94, N92, N90, N73);
nor NOR2 (N95, N59, N23);
nand NAND2 (N96, N94, N94);
buf BUF1 (N97, N91);
nand NAND3 (N98, N79, N9, N79);
nand NAND4 (N99, N77, N33, N11, N58);
nand NAND4 (N100, N82, N40, N61, N32);
buf BUF1 (N101, N96);
nor NOR4 (N102, N98, N50, N27, N39);
nor NOR3 (N103, N95, N91, N73);
nand NAND4 (N104, N89, N48, N47, N62);
buf BUF1 (N105, N69);
xor XOR2 (N106, N105, N87);
and AND4 (N107, N103, N65, N44, N31);
xor XOR2 (N108, N99, N107);
buf BUF1 (N109, N80);
or OR4 (N110, N97, N2, N39, N104);
buf BUF1 (N111, N44);
not NOT1 (N112, N102);
nand NAND4 (N113, N108, N108, N77, N31);
buf BUF1 (N114, N112);
not NOT1 (N115, N111);
and AND3 (N116, N100, N30, N90);
nand NAND3 (N117, N93, N3, N17);
xor XOR2 (N118, N106, N44);
or OR4 (N119, N117, N55, N36, N8);
and AND3 (N120, N113, N7, N119);
buf BUF1 (N121, N101);
xor XOR2 (N122, N48, N20);
nor NOR2 (N123, N116, N9);
nand NAND2 (N124, N76, N104);
xor XOR2 (N125, N118, N67);
and AND3 (N126, N123, N86, N50);
not NOT1 (N127, N114);
and AND3 (N128, N127, N101, N126);
buf BUF1 (N129, N120);
and AND2 (N130, N89, N88);
nand NAND2 (N131, N115, N45);
and AND4 (N132, N121, N7, N50, N65);
xor XOR2 (N133, N110, N85);
buf BUF1 (N134, N125);
nand NAND2 (N135, N122, N94);
nor NOR4 (N136, N132, N74, N128, N105);
nor NOR4 (N137, N89, N122, N96, N134);
buf BUF1 (N138, N93);
nand NAND2 (N139, N136, N2);
not NOT1 (N140, N131);
buf BUF1 (N141, N138);
buf BUF1 (N142, N140);
and AND3 (N143, N130, N113, N81);
xor XOR2 (N144, N109, N78);
nor NOR3 (N145, N124, N90, N32);
and AND3 (N146, N143, N53, N108);
buf BUF1 (N147, N144);
nor NOR4 (N148, N137, N73, N104, N14);
not NOT1 (N149, N148);
xor XOR2 (N150, N142, N121);
xor XOR2 (N151, N147, N127);
and AND2 (N152, N135, N100);
not NOT1 (N153, N152);
nand NAND2 (N154, N133, N18);
or OR2 (N155, N141, N4);
and AND2 (N156, N150, N90);
or OR3 (N157, N156, N142, N106);
and AND2 (N158, N129, N117);
or OR2 (N159, N155, N121);
and AND3 (N160, N145, N84, N34);
not NOT1 (N161, N158);
or OR3 (N162, N159, N36, N57);
buf BUF1 (N163, N153);
not NOT1 (N164, N151);
nand NAND3 (N165, N157, N95, N142);
not NOT1 (N166, N146);
not NOT1 (N167, N149);
buf BUF1 (N168, N164);
xor XOR2 (N169, N168, N145);
and AND3 (N170, N154, N61, N89);
or OR4 (N171, N170, N60, N112, N166);
nor NOR2 (N172, N102, N158);
or OR2 (N173, N172, N54);
nand NAND3 (N174, N139, N107, N173);
nor NOR4 (N175, N15, N41, N155, N167);
not NOT1 (N176, N37);
nor NOR4 (N177, N174, N149, N142, N154);
buf BUF1 (N178, N163);
buf BUF1 (N179, N175);
and AND3 (N180, N177, N43, N17);
or OR4 (N181, N160, N87, N57, N143);
or OR2 (N182, N181, N111);
buf BUF1 (N183, N165);
nand NAND3 (N184, N161, N1, N168);
not NOT1 (N185, N179);
xor XOR2 (N186, N184, N61);
not NOT1 (N187, N183);
and AND2 (N188, N185, N103);
or OR2 (N189, N186, N50);
xor XOR2 (N190, N182, N144);
and AND3 (N191, N162, N82, N125);
and AND2 (N192, N187, N174);
nor NOR2 (N193, N171, N170);
nor NOR3 (N194, N188, N135, N190);
nand NAND2 (N195, N174, N179);
nand NAND4 (N196, N180, N142, N103, N148);
not NOT1 (N197, N176);
and AND2 (N198, N178, N176);
or OR4 (N199, N198, N69, N86, N2);
or OR3 (N200, N197, N184, N107);
not NOT1 (N201, N194);
and AND3 (N202, N191, N180, N147);
and AND2 (N203, N201, N179);
not NOT1 (N204, N169);
or OR2 (N205, N193, N18);
buf BUF1 (N206, N204);
not NOT1 (N207, N202);
nand NAND3 (N208, N203, N178, N71);
or OR3 (N209, N195, N18, N182);
xor XOR2 (N210, N199, N1);
or OR2 (N211, N207, N167);
and AND4 (N212, N211, N51, N117, N97);
buf BUF1 (N213, N189);
or OR2 (N214, N200, N1);
nand NAND4 (N215, N212, N163, N160, N193);
or OR2 (N216, N192, N166);
not NOT1 (N217, N208);
nand NAND4 (N218, N217, N152, N206, N116);
buf BUF1 (N219, N27);
nor NOR3 (N220, N216, N203, N32);
buf BUF1 (N221, N196);
nor NOR4 (N222, N214, N101, N86, N32);
nor NOR4 (N223, N218, N141, N100, N26);
nor NOR4 (N224, N205, N128, N48, N23);
buf BUF1 (N225, N224);
nor NOR3 (N226, N225, N94, N193);
buf BUF1 (N227, N210);
not NOT1 (N228, N226);
nand NAND2 (N229, N221, N187);
or OR2 (N230, N220, N88);
xor XOR2 (N231, N223, N219);
not NOT1 (N232, N141);
or OR4 (N233, N229, N137, N27, N179);
not NOT1 (N234, N231);
buf BUF1 (N235, N222);
and AND4 (N236, N233, N157, N1, N79);
nand NAND2 (N237, N235, N226);
buf BUF1 (N238, N213);
buf BUF1 (N239, N237);
and AND4 (N240, N238, N131, N85, N31);
nor NOR3 (N241, N215, N171, N186);
and AND2 (N242, N209, N124);
not NOT1 (N243, N239);
nor NOR3 (N244, N243, N25, N90);
buf BUF1 (N245, N234);
xor XOR2 (N246, N227, N162);
nor NOR4 (N247, N242, N129, N32, N50);
nor NOR3 (N248, N240, N202, N107);
nor NOR3 (N249, N248, N49, N119);
xor XOR2 (N250, N232, N80);
buf BUF1 (N251, N228);
buf BUF1 (N252, N245);
or OR3 (N253, N246, N135, N214);
buf BUF1 (N254, N236);
or OR2 (N255, N251, N61);
xor XOR2 (N256, N244, N75);
nor NOR4 (N257, N241, N88, N211, N141);
xor XOR2 (N258, N230, N7);
xor XOR2 (N259, N247, N86);
nand NAND4 (N260, N252, N156, N14, N75);
not NOT1 (N261, N253);
and AND3 (N262, N255, N181, N195);
buf BUF1 (N263, N259);
not NOT1 (N264, N254);
nor NOR3 (N265, N263, N196, N15);
xor XOR2 (N266, N260, N85);
buf BUF1 (N267, N250);
or OR4 (N268, N261, N185, N74, N174);
or OR4 (N269, N268, N84, N157, N91);
not NOT1 (N270, N262);
not NOT1 (N271, N258);
or OR3 (N272, N270, N235, N26);
not NOT1 (N273, N264);
not NOT1 (N274, N269);
nand NAND2 (N275, N267, N228);
or OR2 (N276, N266, N79);
nor NOR4 (N277, N272, N183, N93, N216);
and AND4 (N278, N274, N227, N270, N127);
xor XOR2 (N279, N265, N41);
xor XOR2 (N280, N277, N156);
xor XOR2 (N281, N273, N248);
and AND4 (N282, N256, N155, N227, N83);
not NOT1 (N283, N281);
nand NAND4 (N284, N278, N97, N182, N267);
nand NAND2 (N285, N257, N195);
nor NOR3 (N286, N285, N241, N262);
nand NAND2 (N287, N276, N140);
buf BUF1 (N288, N280);
or OR2 (N289, N279, N38);
nor NOR2 (N290, N287, N104);
nand NAND4 (N291, N271, N114, N134, N47);
nand NAND2 (N292, N283, N121);
xor XOR2 (N293, N275, N218);
nor NOR4 (N294, N291, N114, N170, N144);
or OR3 (N295, N288, N238, N125);
or OR4 (N296, N282, N78, N50, N140);
buf BUF1 (N297, N295);
or OR3 (N298, N290, N207, N57);
nand NAND4 (N299, N297, N102, N121, N64);
not NOT1 (N300, N292);
and AND4 (N301, N293, N98, N94, N9);
or OR3 (N302, N294, N208, N272);
buf BUF1 (N303, N286);
not NOT1 (N304, N299);
xor XOR2 (N305, N296, N210);
and AND2 (N306, N305, N99);
xor XOR2 (N307, N289, N143);
not NOT1 (N308, N303);
nand NAND4 (N309, N301, N296, N237, N161);
buf BUF1 (N310, N307);
xor XOR2 (N311, N249, N220);
buf BUF1 (N312, N298);
or OR3 (N313, N310, N60, N173);
not NOT1 (N314, N313);
buf BUF1 (N315, N306);
not NOT1 (N316, N302);
nor NOR4 (N317, N300, N49, N294, N58);
and AND4 (N318, N315, N107, N31, N252);
not NOT1 (N319, N309);
not NOT1 (N320, N304);
or OR4 (N321, N308, N18, N42, N259);
or OR3 (N322, N317, N34, N138);
xor XOR2 (N323, N316, N260);
nand NAND4 (N324, N319, N259, N212, N20);
nand NAND4 (N325, N324, N41, N243, N181);
not NOT1 (N326, N322);
and AND3 (N327, N312, N320, N117);
buf BUF1 (N328, N133);
buf BUF1 (N329, N325);
and AND3 (N330, N327, N1, N14);
xor XOR2 (N331, N318, N150);
nand NAND2 (N332, N321, N197);
xor XOR2 (N333, N329, N288);
nor NOR3 (N334, N284, N206, N314);
and AND2 (N335, N3, N181);
not NOT1 (N336, N323);
nor NOR3 (N337, N328, N90, N17);
and AND2 (N338, N332, N109);
and AND4 (N339, N331, N233, N76, N69);
and AND2 (N340, N326, N153);
or OR4 (N341, N340, N67, N36, N330);
not NOT1 (N342, N271);
or OR2 (N343, N336, N309);
or OR4 (N344, N342, N5, N308, N82);
nor NOR4 (N345, N337, N4, N32, N185);
and AND2 (N346, N335, N60);
and AND2 (N347, N339, N246);
xor XOR2 (N348, N338, N241);
and AND3 (N349, N345, N93, N273);
buf BUF1 (N350, N347);
buf BUF1 (N351, N344);
not NOT1 (N352, N346);
and AND2 (N353, N348, N217);
xor XOR2 (N354, N352, N16);
or OR3 (N355, N350, N98, N315);
nand NAND2 (N356, N343, N313);
nand NAND4 (N357, N355, N59, N132, N253);
nand NAND4 (N358, N351, N163, N343, N19);
xor XOR2 (N359, N358, N193);
nand NAND4 (N360, N334, N72, N223, N56);
buf BUF1 (N361, N341);
nor NOR4 (N362, N359, N204, N39, N89);
nor NOR3 (N363, N353, N198, N208);
xor XOR2 (N364, N333, N50);
not NOT1 (N365, N357);
nand NAND2 (N366, N361, N339);
xor XOR2 (N367, N363, N350);
buf BUF1 (N368, N354);
or OR3 (N369, N366, N204, N298);
and AND3 (N370, N369, N153, N365);
xor XOR2 (N371, N220, N26);
buf BUF1 (N372, N368);
nand NAND3 (N373, N349, N193, N65);
buf BUF1 (N374, N360);
buf BUF1 (N375, N374);
nand NAND3 (N376, N372, N325, N305);
xor XOR2 (N377, N311, N175);
buf BUF1 (N378, N376);
and AND4 (N379, N362, N66, N152, N196);
nand NAND2 (N380, N364, N217);
not NOT1 (N381, N377);
nor NOR3 (N382, N381, N321, N381);
nand NAND4 (N383, N379, N228, N33, N1);
xor XOR2 (N384, N371, N24);
nor NOR3 (N385, N383, N220, N154);
nor NOR3 (N386, N380, N275, N169);
nand NAND3 (N387, N384, N159, N162);
not NOT1 (N388, N367);
xor XOR2 (N389, N388, N314);
xor XOR2 (N390, N382, N139);
nor NOR4 (N391, N386, N60, N305, N206);
not NOT1 (N392, N389);
not NOT1 (N393, N356);
and AND4 (N394, N385, N126, N249, N225);
and AND3 (N395, N375, N118, N334);
buf BUF1 (N396, N392);
buf BUF1 (N397, N390);
and AND2 (N398, N395, N335);
buf BUF1 (N399, N387);
or OR3 (N400, N394, N163, N15);
or OR2 (N401, N398, N303);
or OR3 (N402, N393, N288, N268);
xor XOR2 (N403, N391, N223);
and AND4 (N404, N378, N255, N277, N300);
not NOT1 (N405, N403);
buf BUF1 (N406, N405);
xor XOR2 (N407, N401, N186);
buf BUF1 (N408, N396);
nor NOR4 (N409, N407, N123, N203, N338);
nand NAND4 (N410, N399, N408, N332, N182);
nand NAND2 (N411, N117, N261);
and AND3 (N412, N406, N8, N130);
or OR2 (N413, N397, N245);
and AND3 (N414, N413, N232, N301);
xor XOR2 (N415, N370, N332);
nor NOR3 (N416, N373, N56, N393);
buf BUF1 (N417, N402);
not NOT1 (N418, N409);
not NOT1 (N419, N416);
and AND2 (N420, N410, N220);
not NOT1 (N421, N414);
nand NAND4 (N422, N412, N261, N188, N332);
and AND3 (N423, N422, N349, N120);
xor XOR2 (N424, N400, N356);
xor XOR2 (N425, N421, N4);
and AND2 (N426, N420, N325);
and AND3 (N427, N415, N9, N169);
buf BUF1 (N428, N418);
buf BUF1 (N429, N419);
nand NAND2 (N430, N411, N300);
and AND3 (N431, N427, N388, N41);
and AND2 (N432, N425, N20);
or OR3 (N433, N424, N118, N171);
nand NAND3 (N434, N429, N156, N224);
and AND4 (N435, N404, N340, N270, N198);
and AND3 (N436, N417, N353, N315);
or OR4 (N437, N428, N252, N330, N337);
buf BUF1 (N438, N430);
buf BUF1 (N439, N426);
or OR4 (N440, N436, N114, N213, N70);
buf BUF1 (N441, N423);
nand NAND4 (N442, N441, N70, N303, N360);
nor NOR2 (N443, N442, N363);
and AND3 (N444, N438, N367, N148);
nor NOR2 (N445, N431, N80);
buf BUF1 (N446, N434);
and AND3 (N447, N439, N246, N137);
or OR3 (N448, N447, N430, N182);
and AND3 (N449, N444, N78, N442);
nor NOR3 (N450, N446, N257, N28);
and AND4 (N451, N450, N103, N446, N235);
xor XOR2 (N452, N448, N217);
nor NOR3 (N453, N435, N439, N274);
nand NAND4 (N454, N453, N210, N6, N155);
buf BUF1 (N455, N454);
xor XOR2 (N456, N449, N355);
not NOT1 (N457, N437);
nor NOR2 (N458, N432, N58);
and AND4 (N459, N440, N331, N299, N159);
nor NOR2 (N460, N445, N406);
or OR3 (N461, N433, N147, N323);
nand NAND4 (N462, N458, N33, N127, N38);
or OR2 (N463, N459, N15);
xor XOR2 (N464, N456, N266);
nor NOR2 (N465, N457, N72);
nor NOR4 (N466, N461, N144, N280, N346);
buf BUF1 (N467, N464);
buf BUF1 (N468, N466);
or OR4 (N469, N455, N201, N70, N447);
and AND2 (N470, N451, N258);
and AND2 (N471, N463, N208);
and AND2 (N472, N465, N4);
nor NOR2 (N473, N468, N372);
not NOT1 (N474, N443);
nor NOR3 (N475, N452, N35, N381);
and AND4 (N476, N460, N218, N142, N119);
nor NOR3 (N477, N462, N16, N422);
not NOT1 (N478, N467);
nor NOR4 (N479, N473, N91, N12, N232);
or OR4 (N480, N477, N280, N452, N53);
xor XOR2 (N481, N478, N371);
not NOT1 (N482, N470);
or OR4 (N483, N476, N255, N103, N175);
not NOT1 (N484, N475);
nor NOR4 (N485, N483, N223, N216, N237);
nand NAND3 (N486, N479, N100, N51);
and AND4 (N487, N482, N83, N143, N227);
not NOT1 (N488, N480);
buf BUF1 (N489, N472);
xor XOR2 (N490, N474, N208);
buf BUF1 (N491, N481);
nor NOR2 (N492, N471, N155);
not NOT1 (N493, N469);
not NOT1 (N494, N485);
and AND4 (N495, N491, N334, N376, N137);
and AND2 (N496, N484, N238);
buf BUF1 (N497, N494);
buf BUF1 (N498, N490);
and AND4 (N499, N492, N115, N302, N247);
or OR2 (N500, N498, N485);
or OR3 (N501, N495, N102, N485);
xor XOR2 (N502, N493, N392);
buf BUF1 (N503, N502);
not NOT1 (N504, N503);
xor XOR2 (N505, N487, N460);
nor NOR4 (N506, N499, N172, N338, N406);
not NOT1 (N507, N486);
buf BUF1 (N508, N488);
nor NOR2 (N509, N489, N210);
nor NOR4 (N510, N504, N320, N400, N354);
nor NOR3 (N511, N508, N433, N250);
nand NAND3 (N512, N496, N184, N269);
or OR4 (N513, N500, N291, N256, N365);
nor NOR2 (N514, N507, N473);
or OR4 (N515, N509, N505, N258, N378);
nand NAND2 (N516, N99, N88);
nand NAND2 (N517, N501, N147);
xor XOR2 (N518, N512, N267);
and AND3 (N519, N513, N225, N290);
nor NOR4 (N520, N518, N17, N431, N256);
and AND2 (N521, N497, N511);
and AND3 (N522, N490, N232, N497);
or OR4 (N523, N521, N284, N231, N339);
buf BUF1 (N524, N514);
and AND4 (N525, N519, N92, N350, N312);
not NOT1 (N526, N522);
nor NOR4 (N527, N520, N222, N440, N310);
and AND3 (N528, N523, N448, N76);
not NOT1 (N529, N528);
not NOT1 (N530, N506);
nor NOR3 (N531, N530, N45, N463);
nor NOR2 (N532, N531, N516);
xor XOR2 (N533, N292, N214);
buf BUF1 (N534, N529);
xor XOR2 (N535, N526, N517);
and AND2 (N536, N444, N226);
or OR3 (N537, N532, N306, N386);
not NOT1 (N538, N535);
and AND4 (N539, N524, N331, N211, N3);
xor XOR2 (N540, N527, N381);
not NOT1 (N541, N525);
nor NOR3 (N542, N533, N408, N106);
xor XOR2 (N543, N542, N53);
nand NAND4 (N544, N537, N7, N349, N269);
nand NAND3 (N545, N544, N215, N147);
not NOT1 (N546, N510);
nor NOR2 (N547, N545, N41);
nand NAND3 (N548, N547, N379, N263);
nor NOR4 (N549, N515, N119, N140, N119);
not NOT1 (N550, N540);
and AND2 (N551, N550, N95);
nor NOR3 (N552, N539, N258, N30);
and AND4 (N553, N534, N254, N496, N404);
xor XOR2 (N554, N552, N368);
nor NOR2 (N555, N551, N406);
or OR2 (N556, N554, N436);
not NOT1 (N557, N541);
nand NAND2 (N558, N538, N347);
nand NAND4 (N559, N546, N398, N406, N245);
xor XOR2 (N560, N556, N195);
nand NAND4 (N561, N557, N150, N94, N376);
xor XOR2 (N562, N553, N452);
xor XOR2 (N563, N559, N159);
buf BUF1 (N564, N555);
nor NOR3 (N565, N558, N421, N523);
or OR3 (N566, N536, N67, N268);
not NOT1 (N567, N561);
or OR4 (N568, N566, N489, N79, N516);
xor XOR2 (N569, N565, N302);
buf BUF1 (N570, N549);
xor XOR2 (N571, N563, N392);
and AND2 (N572, N569, N417);
not NOT1 (N573, N572);
not NOT1 (N574, N571);
buf BUF1 (N575, N567);
or OR4 (N576, N570, N478, N275, N528);
not NOT1 (N577, N543);
or OR4 (N578, N577, N6, N290, N15);
nor NOR4 (N579, N575, N26, N266, N261);
nor NOR2 (N580, N574, N214);
xor XOR2 (N581, N562, N436);
buf BUF1 (N582, N578);
xor XOR2 (N583, N576, N226);
and AND3 (N584, N579, N6, N7);
and AND3 (N585, N580, N333, N211);
nor NOR2 (N586, N568, N459);
nor NOR4 (N587, N584, N30, N138, N379);
not NOT1 (N588, N573);
and AND3 (N589, N585, N452, N514);
not NOT1 (N590, N589);
not NOT1 (N591, N548);
not NOT1 (N592, N587);
buf BUF1 (N593, N583);
nand NAND3 (N594, N588, N217, N198);
and AND4 (N595, N593, N580, N108, N553);
nand NAND4 (N596, N591, N172, N360, N251);
buf BUF1 (N597, N586);
buf BUF1 (N598, N595);
not NOT1 (N599, N592);
nor NOR2 (N600, N582, N464);
or OR2 (N601, N590, N285);
not NOT1 (N602, N581);
and AND2 (N603, N560, N86);
or OR4 (N604, N597, N268, N337, N211);
xor XOR2 (N605, N564, N313);
nor NOR2 (N606, N601, N588);
buf BUF1 (N607, N606);
buf BUF1 (N608, N605);
and AND2 (N609, N603, N26);
or OR2 (N610, N598, N59);
nand NAND4 (N611, N596, N222, N176, N527);
nand NAND2 (N612, N594, N323);
or OR2 (N613, N602, N266);
xor XOR2 (N614, N610, N197);
xor XOR2 (N615, N611, N530);
nor NOR3 (N616, N609, N326, N266);
nor NOR4 (N617, N614, N30, N4, N272);
and AND3 (N618, N607, N371, N467);
and AND3 (N619, N617, N507, N196);
not NOT1 (N620, N615);
or OR3 (N621, N616, N21, N460);
nand NAND4 (N622, N612, N115, N613, N475);
xor XOR2 (N623, N477, N466);
and AND3 (N624, N621, N240, N141);
and AND3 (N625, N622, N394, N526);
xor XOR2 (N626, N624, N212);
nand NAND2 (N627, N618, N29);
nand NAND4 (N628, N600, N549, N614, N9);
xor XOR2 (N629, N623, N151);
buf BUF1 (N630, N629);
or OR4 (N631, N599, N621, N4, N27);
nand NAND4 (N632, N604, N347, N464, N213);
nand NAND2 (N633, N608, N126);
or OR3 (N634, N619, N487, N585);
or OR2 (N635, N627, N350);
nor NOR3 (N636, N626, N129, N446);
and AND3 (N637, N625, N583, N129);
and AND3 (N638, N630, N277, N54);
nand NAND3 (N639, N628, N338, N421);
nor NOR2 (N640, N633, N410);
xor XOR2 (N641, N636, N133);
not NOT1 (N642, N635);
and AND4 (N643, N637, N501, N409, N477);
xor XOR2 (N644, N641, N386);
not NOT1 (N645, N631);
and AND4 (N646, N632, N366, N550, N499);
buf BUF1 (N647, N642);
nor NOR4 (N648, N644, N128, N36, N216);
or OR4 (N649, N646, N344, N92, N291);
and AND2 (N650, N647, N225);
and AND4 (N651, N645, N470, N488, N628);
and AND3 (N652, N634, N527, N179);
or OR4 (N653, N649, N589, N27, N545);
and AND3 (N654, N653, N642, N221);
and AND2 (N655, N638, N252);
and AND2 (N656, N654, N388);
nor NOR4 (N657, N648, N540, N608, N6);
and AND3 (N658, N656, N637, N189);
xor XOR2 (N659, N655, N107);
not NOT1 (N660, N652);
nor NOR3 (N661, N659, N134, N552);
nor NOR3 (N662, N643, N630, N402);
or OR2 (N663, N639, N119);
nor NOR3 (N664, N650, N255, N261);
or OR3 (N665, N662, N61, N303);
or OR2 (N666, N664, N469);
buf BUF1 (N667, N657);
nand NAND3 (N668, N667, N382, N1);
or OR4 (N669, N661, N512, N127, N191);
or OR3 (N670, N668, N582, N525);
nor NOR4 (N671, N658, N445, N642, N350);
and AND2 (N672, N665, N124);
or OR2 (N673, N670, N26);
xor XOR2 (N674, N660, N631);
nand NAND2 (N675, N671, N256);
not NOT1 (N676, N640);
nor NOR2 (N677, N663, N289);
xor XOR2 (N678, N666, N597);
nor NOR4 (N679, N651, N151, N130, N274);
buf BUF1 (N680, N673);
xor XOR2 (N681, N677, N341);
not NOT1 (N682, N680);
or OR4 (N683, N675, N243, N175, N124);
xor XOR2 (N684, N676, N666);
and AND4 (N685, N679, N210, N627, N489);
nand NAND2 (N686, N672, N230);
or OR2 (N687, N685, N320);
buf BUF1 (N688, N686);
not NOT1 (N689, N678);
nor NOR3 (N690, N689, N565, N335);
nand NAND2 (N691, N669, N438);
not NOT1 (N692, N690);
or OR3 (N693, N681, N305, N126);
buf BUF1 (N694, N691);
xor XOR2 (N695, N687, N552);
nor NOR2 (N696, N693, N306);
nor NOR4 (N697, N694, N423, N450, N5);
nor NOR2 (N698, N620, N309);
not NOT1 (N699, N684);
buf BUF1 (N700, N699);
xor XOR2 (N701, N674, N414);
nand NAND2 (N702, N688, N59);
nand NAND2 (N703, N692, N692);
buf BUF1 (N704, N703);
nand NAND2 (N705, N700, N679);
nand NAND4 (N706, N704, N195, N576, N281);
or OR4 (N707, N702, N72, N287, N454);
and AND3 (N708, N695, N12, N94);
xor XOR2 (N709, N698, N223);
buf BUF1 (N710, N708);
nand NAND4 (N711, N710, N174, N69, N251);
buf BUF1 (N712, N705);
buf BUF1 (N713, N696);
buf BUF1 (N714, N709);
xor XOR2 (N715, N683, N373);
xor XOR2 (N716, N713, N239);
or OR4 (N717, N716, N69, N629, N471);
nand NAND2 (N718, N682, N89);
and AND3 (N719, N714, N713, N369);
or OR4 (N720, N711, N692, N72, N6);
nor NOR3 (N721, N697, N436, N324);
xor XOR2 (N722, N715, N669);
buf BUF1 (N723, N707);
nor NOR3 (N724, N721, N681, N412);
xor XOR2 (N725, N717, N96);
or OR4 (N726, N725, N104, N563, N418);
nor NOR2 (N727, N701, N57);
not NOT1 (N728, N726);
nand NAND3 (N729, N706, N619, N129);
nor NOR3 (N730, N724, N112, N87);
xor XOR2 (N731, N727, N364);
or OR4 (N732, N712, N143, N294, N527);
not NOT1 (N733, N722);
buf BUF1 (N734, N731);
or OR2 (N735, N732, N207);
nor NOR2 (N736, N729, N501);
and AND3 (N737, N734, N81, N419);
and AND2 (N738, N718, N109);
nand NAND4 (N739, N736, N348, N58, N626);
not NOT1 (N740, N728);
xor XOR2 (N741, N720, N352);
and AND3 (N742, N723, N356, N189);
buf BUF1 (N743, N730);
nor NOR4 (N744, N739, N115, N357, N37);
xor XOR2 (N745, N742, N105);
and AND3 (N746, N738, N551, N367);
buf BUF1 (N747, N743);
and AND4 (N748, N747, N426, N587, N572);
xor XOR2 (N749, N744, N332);
nand NAND2 (N750, N735, N683);
xor XOR2 (N751, N745, N88);
xor XOR2 (N752, N748, N325);
buf BUF1 (N753, N733);
nor NOR2 (N754, N752, N334);
not NOT1 (N755, N740);
buf BUF1 (N756, N753);
nand NAND3 (N757, N719, N304, N367);
nor NOR4 (N758, N749, N580, N430, N447);
or OR4 (N759, N746, N292, N669, N553);
or OR3 (N760, N754, N621, N79);
not NOT1 (N761, N759);
and AND3 (N762, N760, N709, N208);
xor XOR2 (N763, N751, N188);
xor XOR2 (N764, N761, N672);
nand NAND4 (N765, N758, N524, N583, N542);
buf BUF1 (N766, N762);
not NOT1 (N767, N766);
buf BUF1 (N768, N764);
nand NAND3 (N769, N755, N521, N380);
not NOT1 (N770, N757);
buf BUF1 (N771, N763);
buf BUF1 (N772, N741);
buf BUF1 (N773, N772);
buf BUF1 (N774, N756);
or OR4 (N775, N769, N612, N622, N412);
and AND4 (N776, N773, N614, N347, N39);
not NOT1 (N777, N767);
nand NAND2 (N778, N768, N723);
nand NAND4 (N779, N774, N159, N490, N486);
not NOT1 (N780, N776);
buf BUF1 (N781, N775);
xor XOR2 (N782, N779, N705);
buf BUF1 (N783, N782);
buf BUF1 (N784, N765);
and AND2 (N785, N750, N705);
nor NOR3 (N786, N771, N422, N311);
nand NAND3 (N787, N778, N690, N467);
nand NAND4 (N788, N781, N429, N468, N574);
nor NOR3 (N789, N783, N670, N682);
nor NOR2 (N790, N770, N372);
and AND3 (N791, N784, N305, N559);
xor XOR2 (N792, N777, N172);
xor XOR2 (N793, N792, N218);
buf BUF1 (N794, N793);
nor NOR3 (N795, N790, N10, N112);
not NOT1 (N796, N737);
xor XOR2 (N797, N786, N243);
or OR2 (N798, N789, N671);
not NOT1 (N799, N785);
xor XOR2 (N800, N798, N169);
not NOT1 (N801, N795);
or OR2 (N802, N796, N257);
not NOT1 (N803, N791);
and AND4 (N804, N780, N179, N410, N494);
xor XOR2 (N805, N797, N797);
or OR4 (N806, N787, N114, N332, N256);
or OR3 (N807, N800, N633, N47);
nand NAND3 (N808, N802, N787, N489);
buf BUF1 (N809, N788);
xor XOR2 (N810, N809, N403);
and AND3 (N811, N794, N208, N76);
nor NOR4 (N812, N810, N305, N505, N120);
xor XOR2 (N813, N803, N775);
buf BUF1 (N814, N807);
xor XOR2 (N815, N806, N528);
xor XOR2 (N816, N804, N561);
or OR4 (N817, N813, N567, N808, N280);
buf BUF1 (N818, N56);
nor NOR2 (N819, N799, N703);
or OR4 (N820, N812, N719, N209, N277);
nor NOR3 (N821, N819, N615, N752);
and AND3 (N822, N818, N487, N106);
nand NAND2 (N823, N820, N801);
nand NAND3 (N824, N60, N623, N411);
xor XOR2 (N825, N817, N198);
or OR3 (N826, N815, N693, N748);
buf BUF1 (N827, N826);
or OR3 (N828, N805, N432, N331);
nand NAND2 (N829, N811, N84);
and AND2 (N830, N816, N333);
xor XOR2 (N831, N830, N127);
and AND3 (N832, N821, N746, N628);
nand NAND2 (N833, N829, N264);
nor NOR2 (N834, N814, N377);
xor XOR2 (N835, N823, N415);
nand NAND2 (N836, N822, N686);
nand NAND4 (N837, N825, N195, N633, N525);
buf BUF1 (N838, N837);
and AND2 (N839, N831, N609);
nand NAND3 (N840, N834, N116, N376);
nor NOR4 (N841, N827, N653, N556, N736);
xor XOR2 (N842, N841, N103);
not NOT1 (N843, N835);
buf BUF1 (N844, N840);
and AND4 (N845, N844, N321, N316, N378);
nor NOR4 (N846, N824, N407, N804, N379);
and AND2 (N847, N828, N846);
or OR3 (N848, N831, N834, N356);
buf BUF1 (N849, N839);
or OR4 (N850, N845, N135, N549, N164);
not NOT1 (N851, N850);
xor XOR2 (N852, N843, N773);
nand NAND4 (N853, N848, N378, N238, N54);
or OR4 (N854, N836, N289, N217, N691);
not NOT1 (N855, N838);
and AND4 (N856, N832, N595, N661, N244);
nand NAND2 (N857, N852, N295);
nand NAND2 (N858, N847, N682);
nand NAND4 (N859, N833, N654, N694, N259);
buf BUF1 (N860, N858);
nor NOR4 (N861, N854, N6, N549, N676);
buf BUF1 (N862, N855);
nor NOR4 (N863, N856, N763, N101, N698);
xor XOR2 (N864, N853, N221);
not NOT1 (N865, N863);
not NOT1 (N866, N857);
or OR2 (N867, N860, N230);
nand NAND2 (N868, N867, N346);
and AND2 (N869, N851, N791);
and AND3 (N870, N862, N794, N534);
xor XOR2 (N871, N870, N833);
not NOT1 (N872, N864);
and AND4 (N873, N865, N234, N568, N452);
nand NAND2 (N874, N868, N96);
not NOT1 (N875, N842);
buf BUF1 (N876, N859);
xor XOR2 (N877, N869, N485);
xor XOR2 (N878, N871, N544);
and AND2 (N879, N872, N770);
nor NOR3 (N880, N874, N392, N752);
not NOT1 (N881, N873);
nor NOR3 (N882, N877, N383, N507);
buf BUF1 (N883, N881);
nor NOR3 (N884, N883, N863, N774);
buf BUF1 (N885, N884);
xor XOR2 (N886, N875, N422);
nor NOR3 (N887, N886, N784, N656);
not NOT1 (N888, N861);
nor NOR2 (N889, N849, N109);
nor NOR4 (N890, N866, N172, N162, N831);
not NOT1 (N891, N882);
and AND4 (N892, N888, N346, N695, N85);
buf BUF1 (N893, N876);
and AND4 (N894, N891, N714, N19, N767);
nand NAND4 (N895, N878, N161, N501, N684);
not NOT1 (N896, N885);
nor NOR2 (N897, N887, N799);
nor NOR4 (N898, N880, N37, N809, N331);
nand NAND4 (N899, N889, N237, N565, N392);
xor XOR2 (N900, N896, N108);
or OR4 (N901, N899, N641, N444, N512);
and AND3 (N902, N894, N458, N270);
nor NOR3 (N903, N895, N642, N554);
xor XOR2 (N904, N893, N448);
nor NOR4 (N905, N898, N210, N594, N199);
and AND2 (N906, N901, N834);
nor NOR2 (N907, N897, N88);
buf BUF1 (N908, N879);
nand NAND2 (N909, N906, N267);
and AND4 (N910, N909, N859, N516, N715);
or OR2 (N911, N910, N348);
not NOT1 (N912, N890);
nor NOR2 (N913, N892, N187);
nor NOR2 (N914, N904, N168);
nand NAND3 (N915, N905, N134, N676);
nand NAND2 (N916, N902, N176);
or OR3 (N917, N900, N125, N275);
nor NOR4 (N918, N907, N206, N62, N31);
not NOT1 (N919, N915);
not NOT1 (N920, N919);
xor XOR2 (N921, N913, N447);
nor NOR3 (N922, N908, N584, N173);
nand NAND3 (N923, N916, N56, N717);
nor NOR2 (N924, N923, N175);
not NOT1 (N925, N911);
not NOT1 (N926, N917);
not NOT1 (N927, N918);
and AND3 (N928, N927, N795, N285);
or OR4 (N929, N928, N913, N925, N732);
buf BUF1 (N930, N659);
or OR3 (N931, N922, N245, N904);
and AND3 (N932, N921, N114, N294);
buf BUF1 (N933, N924);
not NOT1 (N934, N914);
not NOT1 (N935, N903);
nor NOR4 (N936, N920, N830, N700, N777);
not NOT1 (N937, N936);
or OR4 (N938, N932, N377, N398, N845);
and AND2 (N939, N912, N326);
and AND2 (N940, N934, N768);
and AND4 (N941, N929, N195, N390, N41);
xor XOR2 (N942, N939, N717);
and AND2 (N943, N935, N344);
xor XOR2 (N944, N931, N839);
and AND2 (N945, N943, N811);
xor XOR2 (N946, N933, N114);
nand NAND3 (N947, N944, N769, N539);
buf BUF1 (N948, N938);
nor NOR2 (N949, N946, N890);
buf BUF1 (N950, N937);
not NOT1 (N951, N950);
or OR2 (N952, N942, N563);
nor NOR2 (N953, N926, N319);
nor NOR3 (N954, N948, N942, N111);
nand NAND2 (N955, N954, N102);
or OR4 (N956, N940, N74, N329, N203);
xor XOR2 (N957, N949, N828);
nor NOR3 (N958, N957, N2, N588);
xor XOR2 (N959, N952, N743);
buf BUF1 (N960, N945);
nand NAND4 (N961, N959, N866, N882, N684);
not NOT1 (N962, N961);
nand NAND2 (N963, N947, N203);
and AND4 (N964, N962, N288, N472, N402);
or OR2 (N965, N930, N676);
buf BUF1 (N966, N958);
not NOT1 (N967, N964);
buf BUF1 (N968, N953);
and AND3 (N969, N960, N378, N763);
and AND2 (N970, N963, N405);
and AND2 (N971, N956, N362);
and AND3 (N972, N967, N231, N843);
buf BUF1 (N973, N965);
and AND4 (N974, N971, N230, N267, N671);
or OR2 (N975, N974, N372);
and AND3 (N976, N975, N820, N544);
or OR2 (N977, N970, N915);
or OR4 (N978, N966, N588, N322, N716);
and AND2 (N979, N977, N64);
not NOT1 (N980, N973);
buf BUF1 (N981, N969);
nor NOR4 (N982, N981, N894, N207, N808);
nand NAND4 (N983, N980, N230, N549, N446);
buf BUF1 (N984, N979);
not NOT1 (N985, N968);
and AND2 (N986, N972, N972);
nand NAND3 (N987, N983, N968, N220);
or OR2 (N988, N984, N465);
xor XOR2 (N989, N987, N497);
xor XOR2 (N990, N955, N543);
buf BUF1 (N991, N978);
or OR2 (N992, N989, N283);
and AND4 (N993, N986, N916, N785, N884);
and AND4 (N994, N992, N214, N805, N663);
or OR4 (N995, N990, N346, N222, N430);
or OR4 (N996, N993, N351, N199, N599);
and AND2 (N997, N994, N876);
and AND3 (N998, N976, N990, N451);
nor NOR4 (N999, N941, N397, N641, N617);
not NOT1 (N1000, N995);
not NOT1 (N1001, N951);
and AND4 (N1002, N999, N956, N701, N820);
or OR4 (N1003, N998, N70, N996, N487);
or OR3 (N1004, N331, N130, N489);
not NOT1 (N1005, N1004);
buf BUF1 (N1006, N1002);
not NOT1 (N1007, N1003);
buf BUF1 (N1008, N1006);
and AND4 (N1009, N1000, N552, N537, N868);
or OR4 (N1010, N991, N332, N756, N428);
not NOT1 (N1011, N982);
not NOT1 (N1012, N1010);
not NOT1 (N1013, N1005);
nor NOR3 (N1014, N1012, N356, N693);
not NOT1 (N1015, N1001);
nor NOR3 (N1016, N1011, N61, N400);
buf BUF1 (N1017, N997);
not NOT1 (N1018, N1008);
or OR2 (N1019, N1007, N848);
and AND3 (N1020, N985, N747, N416);
and AND2 (N1021, N1018, N824);
endmodule