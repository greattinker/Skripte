// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16;

output N1015,N1011,N1009,N1014,N1010,N1007,N1012,N1008,N1013,N1016;

nor NOR4 (N17, N7, N9, N3, N5);
not NOT1 (N18, N3);
not NOT1 (N19, N4);
xor XOR2 (N20, N18, N2);
and AND3 (N21, N3, N3, N15);
buf BUF1 (N22, N8);
not NOT1 (N23, N7);
or OR2 (N24, N18, N1);
xor XOR2 (N25, N23, N18);
nand NAND2 (N26, N13, N12);
and AND3 (N27, N8, N4, N3);
or OR3 (N28, N27, N13, N11);
buf BUF1 (N29, N8);
nor NOR4 (N30, N19, N28, N9, N18);
not NOT1 (N31, N27);
buf BUF1 (N32, N17);
buf BUF1 (N33, N30);
buf BUF1 (N34, N29);
nor NOR4 (N35, N25, N27, N12, N19);
and AND4 (N36, N31, N26, N28, N2);
nand NAND4 (N37, N16, N26, N33, N5);
nand NAND2 (N38, N14, N7);
nor NOR3 (N39, N22, N27, N2);
and AND3 (N40, N37, N2, N30);
nand NAND4 (N41, N39, N19, N19, N7);
or OR2 (N42, N34, N36);
nor NOR4 (N43, N25, N15, N7, N7);
xor XOR2 (N44, N43, N42);
xor XOR2 (N45, N7, N13);
buf BUF1 (N46, N24);
nor NOR2 (N47, N40, N4);
not NOT1 (N48, N45);
buf BUF1 (N49, N48);
and AND4 (N50, N21, N27, N14, N49);
nand NAND4 (N51, N31, N13, N23, N12);
and AND2 (N52, N41, N31);
not NOT1 (N53, N50);
buf BUF1 (N54, N35);
and AND2 (N55, N38, N35);
nand NAND4 (N56, N44, N50, N53, N38);
not NOT1 (N57, N6);
buf BUF1 (N58, N57);
xor XOR2 (N59, N51, N26);
buf BUF1 (N60, N59);
not NOT1 (N61, N55);
xor XOR2 (N62, N58, N48);
nand NAND2 (N63, N54, N33);
nand NAND2 (N64, N20, N15);
xor XOR2 (N65, N60, N45);
or OR2 (N66, N65, N12);
or OR2 (N67, N61, N13);
buf BUF1 (N68, N52);
not NOT1 (N69, N47);
buf BUF1 (N70, N62);
nand NAND4 (N71, N67, N28, N2, N56);
nor NOR2 (N72, N25, N50);
nand NAND4 (N73, N68, N36, N46, N38);
or OR2 (N74, N44, N5);
nor NOR4 (N75, N69, N68, N50, N15);
or OR4 (N76, N75, N31, N18, N53);
xor XOR2 (N77, N32, N57);
nor NOR4 (N78, N64, N21, N61, N7);
nor NOR2 (N79, N76, N64);
buf BUF1 (N80, N74);
xor XOR2 (N81, N66, N74);
or OR3 (N82, N73, N43, N48);
buf BUF1 (N83, N82);
buf BUF1 (N84, N71);
not NOT1 (N85, N72);
and AND4 (N86, N78, N47, N82, N9);
nor NOR2 (N87, N84, N41);
nand NAND2 (N88, N86, N18);
not NOT1 (N89, N63);
not NOT1 (N90, N80);
nor NOR3 (N91, N77, N13, N67);
not NOT1 (N92, N70);
not NOT1 (N93, N83);
not NOT1 (N94, N91);
nand NAND3 (N95, N85, N5, N65);
nor NOR3 (N96, N95, N64, N35);
not NOT1 (N97, N93);
nand NAND2 (N98, N94, N57);
or OR4 (N99, N79, N48, N81, N98);
nor NOR4 (N100, N66, N97, N55, N78);
or OR4 (N101, N88, N67, N8, N13);
nand NAND4 (N102, N62, N25, N88, N22);
or OR4 (N103, N95, N73, N72, N4);
or OR3 (N104, N101, N81, N33);
nand NAND2 (N105, N96, N64);
nand NAND2 (N106, N87, N39);
nor NOR3 (N107, N106, N14, N22);
buf BUF1 (N108, N99);
nand NAND2 (N109, N100, N91);
xor XOR2 (N110, N109, N30);
or OR3 (N111, N103, N93, N86);
xor XOR2 (N112, N92, N101);
or OR4 (N113, N90, N52, N49, N46);
nand NAND2 (N114, N102, N55);
and AND3 (N115, N104, N72, N12);
nor NOR3 (N116, N113, N114, N69);
buf BUF1 (N117, N23);
xor XOR2 (N118, N89, N102);
and AND4 (N119, N108, N74, N75, N30);
xor XOR2 (N120, N115, N73);
or OR3 (N121, N119, N53, N41);
not NOT1 (N122, N121);
or OR3 (N123, N120, N121, N62);
nor NOR4 (N124, N105, N55, N41, N72);
nand NAND3 (N125, N110, N50, N14);
not NOT1 (N126, N117);
nor NOR4 (N127, N116, N61, N71, N13);
buf BUF1 (N128, N125);
buf BUF1 (N129, N112);
or OR4 (N130, N111, N128, N70, N128);
or OR2 (N131, N37, N103);
nor NOR3 (N132, N123, N101, N31);
not NOT1 (N133, N122);
or OR4 (N134, N130, N53, N57, N124);
xor XOR2 (N135, N131, N47);
or OR3 (N136, N87, N44, N38);
nor NOR3 (N137, N118, N66, N132);
buf BUF1 (N138, N127);
buf BUF1 (N139, N86);
buf BUF1 (N140, N126);
nand NAND2 (N141, N134, N108);
xor XOR2 (N142, N107, N104);
and AND3 (N143, N137, N86, N31);
nor NOR3 (N144, N136, N137, N37);
not NOT1 (N145, N141);
nand NAND3 (N146, N129, N5, N90);
buf BUF1 (N147, N138);
or OR4 (N148, N139, N63, N71, N14);
not NOT1 (N149, N148);
nor NOR2 (N150, N140, N32);
and AND3 (N151, N146, N87, N3);
nand NAND2 (N152, N150, N68);
nor NOR4 (N153, N133, N131, N97, N144);
xor XOR2 (N154, N24, N51);
xor XOR2 (N155, N153, N44);
not NOT1 (N156, N154);
or OR3 (N157, N149, N70, N128);
nor NOR4 (N158, N152, N53, N120, N132);
nor NOR4 (N159, N145, N134, N18, N16);
xor XOR2 (N160, N151, N138);
nand NAND2 (N161, N155, N30);
nand NAND4 (N162, N135, N88, N132, N16);
nand NAND2 (N163, N142, N127);
or OR2 (N164, N158, N161);
or OR3 (N165, N24, N117, N21);
and AND3 (N166, N159, N62, N165);
not NOT1 (N167, N18);
buf BUF1 (N168, N164);
nand NAND2 (N169, N166, N14);
buf BUF1 (N170, N147);
not NOT1 (N171, N170);
not NOT1 (N172, N169);
xor XOR2 (N173, N171, N59);
nor NOR4 (N174, N157, N128, N95, N54);
and AND4 (N175, N163, N4, N68, N47);
not NOT1 (N176, N143);
or OR3 (N177, N162, N82, N141);
nand NAND4 (N178, N176, N130, N87, N156);
and AND4 (N179, N79, N97, N143, N124);
nor NOR4 (N180, N172, N94, N27, N72);
nor NOR4 (N181, N180, N75, N18, N153);
xor XOR2 (N182, N160, N145);
or OR4 (N183, N177, N146, N6, N136);
buf BUF1 (N184, N168);
buf BUF1 (N185, N174);
and AND2 (N186, N167, N167);
not NOT1 (N187, N182);
nor NOR4 (N188, N173, N66, N65, N106);
xor XOR2 (N189, N188, N58);
nor NOR3 (N190, N179, N44, N153);
nand NAND4 (N191, N190, N175, N138, N33);
xor XOR2 (N192, N70, N178);
xor XOR2 (N193, N160, N174);
or OR3 (N194, N192, N83, N155);
or OR2 (N195, N181, N54);
nand NAND2 (N196, N194, N29);
buf BUF1 (N197, N187);
or OR2 (N198, N197, N26);
and AND2 (N199, N189, N180);
or OR2 (N200, N186, N57);
and AND2 (N201, N196, N11);
buf BUF1 (N202, N185);
nor NOR2 (N203, N201, N90);
or OR3 (N204, N193, N124, N36);
buf BUF1 (N205, N200);
buf BUF1 (N206, N205);
not NOT1 (N207, N206);
or OR3 (N208, N204, N115, N204);
and AND3 (N209, N191, N190, N10);
or OR3 (N210, N183, N39, N142);
nor NOR4 (N211, N199, N205, N158, N133);
nand NAND4 (N212, N209, N114, N199, N202);
or OR2 (N213, N75, N201);
nor NOR3 (N214, N208, N173, N7);
buf BUF1 (N215, N212);
or OR4 (N216, N203, N56, N57, N88);
nor NOR2 (N217, N198, N199);
nor NOR2 (N218, N210, N149);
not NOT1 (N219, N218);
or OR3 (N220, N215, N62, N21);
not NOT1 (N221, N220);
or OR3 (N222, N213, N118, N44);
not NOT1 (N223, N221);
not NOT1 (N224, N211);
nand NAND2 (N225, N207, N221);
buf BUF1 (N226, N214);
nand NAND3 (N227, N223, N3, N113);
xor XOR2 (N228, N184, N135);
xor XOR2 (N229, N219, N92);
nor NOR2 (N230, N229, N118);
nor NOR3 (N231, N225, N158, N221);
buf BUF1 (N232, N226);
buf BUF1 (N233, N228);
nand NAND2 (N234, N217, N41);
not NOT1 (N235, N224);
nand NAND3 (N236, N235, N209, N120);
not NOT1 (N237, N236);
nor NOR2 (N238, N195, N227);
buf BUF1 (N239, N56);
and AND3 (N240, N233, N176, N49);
or OR3 (N241, N216, N33, N11);
and AND3 (N242, N237, N197, N137);
buf BUF1 (N243, N239);
nand NAND2 (N244, N234, N25);
nand NAND2 (N245, N222, N56);
not NOT1 (N246, N240);
xor XOR2 (N247, N241, N112);
and AND3 (N248, N244, N8, N136);
and AND2 (N249, N247, N41);
and AND4 (N250, N232, N223, N164, N107);
buf BUF1 (N251, N248);
or OR4 (N252, N249, N123, N117, N155);
or OR3 (N253, N245, N211, N110);
not NOT1 (N254, N230);
xor XOR2 (N255, N231, N8);
nand NAND4 (N256, N246, N253, N157, N74);
buf BUF1 (N257, N113);
not NOT1 (N258, N242);
xor XOR2 (N259, N256, N145);
buf BUF1 (N260, N251);
buf BUF1 (N261, N260);
nand NAND3 (N262, N252, N80, N163);
not NOT1 (N263, N255);
not NOT1 (N264, N262);
nand NAND4 (N265, N243, N230, N12, N171);
xor XOR2 (N266, N258, N54);
nor NOR3 (N267, N266, N28, N193);
not NOT1 (N268, N259);
or OR3 (N269, N264, N135, N99);
xor XOR2 (N270, N257, N21);
and AND2 (N271, N267, N41);
or OR2 (N272, N270, N219);
not NOT1 (N273, N272);
or OR2 (N274, N261, N199);
buf BUF1 (N275, N250);
not NOT1 (N276, N274);
not NOT1 (N277, N275);
and AND2 (N278, N238, N207);
nor NOR4 (N279, N265, N66, N240, N261);
nor NOR4 (N280, N277, N184, N190, N243);
buf BUF1 (N281, N254);
and AND3 (N282, N278, N11, N119);
nor NOR2 (N283, N276, N85);
xor XOR2 (N284, N269, N27);
buf BUF1 (N285, N284);
not NOT1 (N286, N271);
nor NOR2 (N287, N286, N146);
buf BUF1 (N288, N273);
not NOT1 (N289, N288);
buf BUF1 (N290, N283);
or OR3 (N291, N280, N13, N196);
nand NAND2 (N292, N279, N74);
xor XOR2 (N293, N263, N184);
or OR2 (N294, N282, N261);
and AND3 (N295, N281, N187, N40);
not NOT1 (N296, N289);
nor NOR2 (N297, N294, N31);
or OR2 (N298, N287, N218);
xor XOR2 (N299, N295, N127);
nor NOR2 (N300, N299, N225);
or OR2 (N301, N296, N175);
nor NOR4 (N302, N301, N218, N244, N253);
nand NAND3 (N303, N298, N152, N188);
buf BUF1 (N304, N285);
and AND3 (N305, N293, N248, N299);
xor XOR2 (N306, N305, N205);
or OR2 (N307, N292, N142);
or OR4 (N308, N304, N271, N26, N127);
buf BUF1 (N309, N308);
xor XOR2 (N310, N307, N143);
nor NOR3 (N311, N291, N152, N157);
nand NAND4 (N312, N311, N62, N11, N149);
nand NAND4 (N313, N309, N69, N168, N132);
buf BUF1 (N314, N300);
or OR4 (N315, N312, N133, N230, N299);
nor NOR2 (N316, N290, N179);
not NOT1 (N317, N314);
nor NOR3 (N318, N317, N309, N107);
xor XOR2 (N319, N268, N157);
or OR3 (N320, N316, N137, N128);
not NOT1 (N321, N315);
nand NAND2 (N322, N321, N220);
xor XOR2 (N323, N303, N146);
nand NAND3 (N324, N306, N297, N119);
or OR4 (N325, N43, N197, N311, N315);
or OR2 (N326, N323, N30);
xor XOR2 (N327, N324, N245);
not NOT1 (N328, N313);
nand NAND2 (N329, N320, N139);
nor NOR3 (N330, N310, N126, N108);
nand NAND3 (N331, N302, N230, N22);
buf BUF1 (N332, N325);
nand NAND2 (N333, N330, N161);
xor XOR2 (N334, N333, N92);
and AND2 (N335, N318, N181);
buf BUF1 (N336, N326);
nor NOR3 (N337, N336, N168, N331);
nand NAND3 (N338, N305, N25, N13);
xor XOR2 (N339, N337, N164);
nand NAND4 (N340, N332, N161, N282, N99);
or OR3 (N341, N329, N198, N274);
nor NOR4 (N342, N335, N109, N74, N135);
and AND4 (N343, N341, N210, N197, N306);
or OR4 (N344, N322, N273, N319, N47);
nor NOR3 (N345, N85, N131, N23);
and AND2 (N346, N345, N224);
buf BUF1 (N347, N328);
or OR4 (N348, N339, N311, N152, N64);
buf BUF1 (N349, N338);
not NOT1 (N350, N348);
and AND4 (N351, N346, N176, N152, N208);
or OR4 (N352, N342, N122, N46, N243);
buf BUF1 (N353, N352);
or OR2 (N354, N334, N260);
and AND2 (N355, N354, N208);
buf BUF1 (N356, N349);
not NOT1 (N357, N343);
nand NAND4 (N358, N355, N305, N350, N32);
not NOT1 (N359, N282);
nor NOR3 (N360, N327, N332, N214);
nor NOR2 (N361, N353, N358);
xor XOR2 (N362, N61, N12);
xor XOR2 (N363, N360, N22);
not NOT1 (N364, N359);
buf BUF1 (N365, N361);
nor NOR4 (N366, N362, N201, N16, N88);
and AND4 (N367, N366, N167, N340, N202);
nor NOR4 (N368, N130, N284, N180, N174);
or OR3 (N369, N368, N87, N266);
and AND3 (N370, N356, N295, N21);
xor XOR2 (N371, N363, N166);
xor XOR2 (N372, N369, N350);
xor XOR2 (N373, N364, N173);
nor NOR2 (N374, N351, N365);
nand NAND2 (N375, N204, N263);
and AND4 (N376, N344, N217, N296, N288);
buf BUF1 (N377, N371);
buf BUF1 (N378, N367);
or OR4 (N379, N378, N25, N133, N286);
or OR2 (N380, N370, N341);
or OR4 (N381, N380, N134, N97, N69);
buf BUF1 (N382, N381);
buf BUF1 (N383, N372);
or OR2 (N384, N376, N225);
nor NOR2 (N385, N383, N193);
buf BUF1 (N386, N347);
and AND4 (N387, N374, N367, N114, N129);
nand NAND4 (N388, N382, N128, N316, N105);
not NOT1 (N389, N373);
xor XOR2 (N390, N386, N139);
or OR4 (N391, N357, N276, N364, N148);
xor XOR2 (N392, N385, N261);
or OR3 (N393, N384, N91, N369);
not NOT1 (N394, N387);
nor NOR4 (N395, N388, N357, N7, N353);
not NOT1 (N396, N389);
or OR3 (N397, N375, N124, N345);
and AND3 (N398, N393, N217, N361);
not NOT1 (N399, N390);
nand NAND4 (N400, N395, N57, N238, N203);
and AND4 (N401, N396, N114, N146, N351);
or OR2 (N402, N397, N114);
nand NAND3 (N403, N379, N164, N127);
xor XOR2 (N404, N399, N275);
nand NAND4 (N405, N398, N39, N85, N37);
nand NAND3 (N406, N377, N162, N188);
xor XOR2 (N407, N392, N372);
buf BUF1 (N408, N406);
not NOT1 (N409, N407);
nor NOR2 (N410, N400, N70);
or OR2 (N411, N402, N65);
buf BUF1 (N412, N405);
xor XOR2 (N413, N411, N328);
or OR2 (N414, N404, N371);
buf BUF1 (N415, N401);
xor XOR2 (N416, N413, N349);
or OR4 (N417, N415, N4, N104, N35);
xor XOR2 (N418, N403, N200);
and AND3 (N419, N408, N171, N109);
nand NAND3 (N420, N414, N175, N404);
nor NOR2 (N421, N412, N238);
buf BUF1 (N422, N410);
buf BUF1 (N423, N391);
nor NOR4 (N424, N418, N316, N52, N421);
nor NOR3 (N425, N363, N266, N293);
or OR3 (N426, N417, N354, N52);
nor NOR3 (N427, N419, N278, N337);
xor XOR2 (N428, N394, N134);
buf BUF1 (N429, N409);
nand NAND4 (N430, N422, N304, N190, N122);
buf BUF1 (N431, N423);
not NOT1 (N432, N429);
not NOT1 (N433, N426);
and AND4 (N434, N428, N374, N57, N205);
not NOT1 (N435, N434);
nand NAND3 (N436, N425, N244, N32);
or OR3 (N437, N424, N379, N71);
and AND3 (N438, N432, N354, N339);
nor NOR4 (N439, N437, N325, N52, N204);
buf BUF1 (N440, N427);
not NOT1 (N441, N440);
buf BUF1 (N442, N439);
xor XOR2 (N443, N436, N181);
not NOT1 (N444, N441);
and AND3 (N445, N438, N109, N155);
nand NAND4 (N446, N435, N40, N280, N392);
not NOT1 (N447, N420);
buf BUF1 (N448, N444);
nand NAND2 (N449, N445, N11);
or OR2 (N450, N433, N322);
nor NOR4 (N451, N446, N33, N390, N324);
not NOT1 (N452, N430);
and AND3 (N453, N452, N56, N19);
nand NAND4 (N454, N449, N319, N22, N182);
nand NAND2 (N455, N416, N333);
xor XOR2 (N456, N442, N270);
buf BUF1 (N457, N455);
xor XOR2 (N458, N450, N387);
buf BUF1 (N459, N451);
nor NOR2 (N460, N431, N80);
buf BUF1 (N461, N459);
nand NAND3 (N462, N447, N358, N447);
and AND2 (N463, N462, N177);
nand NAND4 (N464, N454, N86, N293, N357);
not NOT1 (N465, N463);
or OR3 (N466, N461, N407, N199);
buf BUF1 (N467, N448);
nand NAND4 (N468, N465, N227, N395, N176);
xor XOR2 (N469, N466, N279);
not NOT1 (N470, N456);
and AND4 (N471, N468, N219, N217, N364);
not NOT1 (N472, N467);
or OR3 (N473, N458, N229, N436);
not NOT1 (N474, N460);
not NOT1 (N475, N474);
nor NOR2 (N476, N457, N256);
not NOT1 (N477, N473);
and AND4 (N478, N471, N173, N403, N356);
not NOT1 (N479, N472);
buf BUF1 (N480, N453);
not NOT1 (N481, N443);
and AND4 (N482, N470, N454, N271, N54);
xor XOR2 (N483, N475, N110);
nor NOR3 (N484, N478, N352, N228);
nor NOR3 (N485, N480, N464, N120);
nand NAND3 (N486, N335, N195, N150);
nand NAND2 (N487, N483, N159);
or OR2 (N488, N482, N182);
not NOT1 (N489, N481);
buf BUF1 (N490, N484);
xor XOR2 (N491, N477, N232);
or OR2 (N492, N488, N489);
and AND4 (N493, N237, N262, N413, N328);
nor NOR2 (N494, N485, N444);
not NOT1 (N495, N491);
buf BUF1 (N496, N493);
nor NOR2 (N497, N496, N84);
or OR4 (N498, N494, N120, N103, N20);
xor XOR2 (N499, N469, N242);
nand NAND2 (N500, N476, N328);
xor XOR2 (N501, N500, N56);
nand NAND4 (N502, N495, N203, N280, N14);
nor NOR2 (N503, N498, N292);
buf BUF1 (N504, N486);
or OR4 (N505, N479, N17, N83, N472);
or OR3 (N506, N502, N39, N279);
not NOT1 (N507, N504);
buf BUF1 (N508, N507);
nor NOR3 (N509, N497, N81, N228);
not NOT1 (N510, N487);
xor XOR2 (N511, N503, N192);
not NOT1 (N512, N509);
xor XOR2 (N513, N512, N461);
nor NOR4 (N514, N508, N473, N458, N466);
buf BUF1 (N515, N490);
nor NOR4 (N516, N501, N67, N157, N172);
nand NAND3 (N517, N499, N364, N377);
buf BUF1 (N518, N514);
not NOT1 (N519, N515);
not NOT1 (N520, N513);
or OR4 (N521, N511, N169, N168, N13);
nand NAND2 (N522, N506, N146);
not NOT1 (N523, N517);
buf BUF1 (N524, N520);
and AND4 (N525, N521, N522, N174, N246);
nor NOR3 (N526, N452, N247, N342);
nand NAND2 (N527, N518, N288);
nand NAND4 (N528, N519, N197, N13, N406);
xor XOR2 (N529, N505, N447);
buf BUF1 (N530, N527);
nand NAND3 (N531, N524, N406, N501);
nand NAND4 (N532, N525, N450, N479, N155);
and AND2 (N533, N532, N218);
nor NOR3 (N534, N531, N63, N416);
xor XOR2 (N535, N523, N446);
or OR2 (N536, N528, N373);
and AND3 (N537, N535, N516, N56);
nor NOR3 (N538, N110, N222, N90);
or OR2 (N539, N529, N201);
nand NAND4 (N540, N510, N217, N420, N126);
not NOT1 (N541, N538);
nor NOR2 (N542, N537, N500);
or OR4 (N543, N542, N268, N430, N58);
or OR3 (N544, N539, N11, N104);
xor XOR2 (N545, N534, N143);
not NOT1 (N546, N492);
nor NOR3 (N547, N546, N472, N298);
xor XOR2 (N548, N536, N452);
nand NAND2 (N549, N543, N98);
nand NAND4 (N550, N545, N121, N211, N58);
not NOT1 (N551, N541);
not NOT1 (N552, N549);
buf BUF1 (N553, N551);
buf BUF1 (N554, N553);
nand NAND4 (N555, N548, N46, N413, N166);
not NOT1 (N556, N530);
nand NAND3 (N557, N540, N518, N68);
not NOT1 (N558, N547);
nor NOR4 (N559, N556, N31, N221, N170);
buf BUF1 (N560, N557);
or OR3 (N561, N550, N552, N230);
or OR2 (N562, N441, N425);
nor NOR4 (N563, N559, N263, N302, N416);
nor NOR3 (N564, N563, N156, N98);
xor XOR2 (N565, N562, N63);
or OR4 (N566, N561, N535, N412, N356);
nor NOR4 (N567, N558, N182, N505, N431);
and AND4 (N568, N526, N507, N109, N34);
nand NAND2 (N569, N554, N171);
and AND2 (N570, N569, N296);
buf BUF1 (N571, N555);
or OR2 (N572, N568, N523);
xor XOR2 (N573, N572, N32);
or OR2 (N574, N544, N426);
buf BUF1 (N575, N574);
not NOT1 (N576, N533);
not NOT1 (N577, N560);
or OR3 (N578, N573, N367, N305);
and AND4 (N579, N566, N4, N244, N75);
and AND4 (N580, N570, N152, N250, N579);
not NOT1 (N581, N273);
not NOT1 (N582, N580);
and AND2 (N583, N576, N375);
or OR4 (N584, N581, N529, N403, N261);
not NOT1 (N585, N571);
buf BUF1 (N586, N584);
buf BUF1 (N587, N567);
and AND4 (N588, N586, N173, N280, N486);
not NOT1 (N589, N577);
nor NOR4 (N590, N578, N389, N487, N47);
nand NAND2 (N591, N575, N152);
buf BUF1 (N592, N588);
not NOT1 (N593, N587);
nand NAND4 (N594, N583, N101, N593, N468);
or OR4 (N595, N82, N400, N493, N454);
xor XOR2 (N596, N564, N577);
nor NOR3 (N597, N585, N240, N466);
xor XOR2 (N598, N592, N426);
nor NOR4 (N599, N582, N329, N263, N11);
buf BUF1 (N600, N596);
buf BUF1 (N601, N594);
nand NAND3 (N602, N590, N590, N459);
not NOT1 (N603, N599);
xor XOR2 (N604, N601, N227);
buf BUF1 (N605, N595);
buf BUF1 (N606, N600);
nor NOR4 (N607, N606, N383, N215, N14);
or OR4 (N608, N607, N264, N425, N201);
or OR2 (N609, N598, N202);
not NOT1 (N610, N605);
xor XOR2 (N611, N565, N67);
nor NOR3 (N612, N604, N226, N157);
and AND3 (N613, N603, N98, N508);
and AND3 (N614, N591, N357, N521);
nor NOR2 (N615, N612, N385);
nor NOR2 (N616, N589, N498);
buf BUF1 (N617, N614);
buf BUF1 (N618, N617);
not NOT1 (N619, N602);
nand NAND3 (N620, N613, N7, N124);
xor XOR2 (N621, N609, N153);
xor XOR2 (N622, N611, N254);
not NOT1 (N623, N620);
nor NOR4 (N624, N623, N378, N3, N394);
not NOT1 (N625, N610);
xor XOR2 (N626, N622, N151);
xor XOR2 (N627, N619, N159);
nand NAND3 (N628, N608, N63, N393);
not NOT1 (N629, N624);
not NOT1 (N630, N615);
and AND3 (N631, N625, N215, N350);
xor XOR2 (N632, N626, N157);
xor XOR2 (N633, N632, N503);
not NOT1 (N634, N618);
nand NAND4 (N635, N634, N347, N255, N198);
xor XOR2 (N636, N616, N180);
not NOT1 (N637, N635);
nand NAND2 (N638, N627, N511);
nor NOR3 (N639, N630, N379, N506);
and AND4 (N640, N621, N391, N24, N120);
not NOT1 (N641, N640);
not NOT1 (N642, N641);
not NOT1 (N643, N642);
buf BUF1 (N644, N597);
xor XOR2 (N645, N633, N454);
xor XOR2 (N646, N645, N244);
not NOT1 (N647, N644);
or OR3 (N648, N639, N600, N31);
nand NAND2 (N649, N631, N364);
nand NAND4 (N650, N648, N302, N111, N179);
xor XOR2 (N651, N643, N31);
xor XOR2 (N652, N649, N161);
and AND4 (N653, N651, N482, N633, N18);
buf BUF1 (N654, N629);
and AND2 (N655, N637, N506);
buf BUF1 (N656, N650);
and AND4 (N657, N646, N461, N265, N268);
or OR3 (N658, N653, N335, N258);
xor XOR2 (N659, N654, N65);
not NOT1 (N660, N657);
nand NAND3 (N661, N628, N73, N209);
nand NAND3 (N662, N658, N78, N13);
and AND4 (N663, N647, N121, N442, N361);
xor XOR2 (N664, N655, N325);
xor XOR2 (N665, N661, N179);
nor NOR4 (N666, N638, N646, N545, N533);
and AND4 (N667, N652, N414, N620, N281);
buf BUF1 (N668, N660);
buf BUF1 (N669, N668);
or OR3 (N670, N664, N515, N328);
nor NOR4 (N671, N666, N418, N564, N178);
not NOT1 (N672, N663);
nand NAND3 (N673, N672, N435, N450);
nor NOR4 (N674, N669, N281, N55, N130);
nand NAND4 (N675, N674, N540, N64, N168);
buf BUF1 (N676, N675);
buf BUF1 (N677, N656);
not NOT1 (N678, N665);
xor XOR2 (N679, N670, N459);
nor NOR3 (N680, N636, N559, N220);
buf BUF1 (N681, N659);
xor XOR2 (N682, N677, N234);
and AND3 (N683, N673, N555, N18);
nor NOR4 (N684, N667, N354, N185, N18);
not NOT1 (N685, N683);
or OR3 (N686, N682, N115, N525);
buf BUF1 (N687, N681);
or OR4 (N688, N686, N604, N138, N138);
buf BUF1 (N689, N684);
nand NAND3 (N690, N685, N152, N598);
or OR4 (N691, N689, N657, N275, N585);
nand NAND3 (N692, N671, N94, N176);
not NOT1 (N693, N691);
nor NOR4 (N694, N662, N243, N370, N56);
nand NAND4 (N695, N693, N544, N459, N624);
nand NAND3 (N696, N680, N271, N642);
nand NAND2 (N697, N696, N176);
not NOT1 (N698, N678);
or OR2 (N699, N695, N578);
or OR3 (N700, N699, N377, N271);
nor NOR2 (N701, N676, N672);
not NOT1 (N702, N698);
nand NAND2 (N703, N687, N373);
and AND4 (N704, N697, N494, N409, N482);
not NOT1 (N705, N694);
nor NOR2 (N706, N692, N565);
and AND2 (N707, N706, N434);
nor NOR4 (N708, N700, N338, N536, N197);
and AND2 (N709, N705, N454);
nor NOR3 (N710, N709, N146, N389);
nand NAND3 (N711, N690, N526, N132);
xor XOR2 (N712, N701, N89);
and AND2 (N713, N703, N75);
and AND3 (N714, N679, N7, N109);
nand NAND3 (N715, N704, N217, N265);
and AND4 (N716, N712, N428, N671, N200);
buf BUF1 (N717, N714);
nor NOR4 (N718, N688, N497, N710, N190);
not NOT1 (N719, N279);
nor NOR4 (N720, N718, N170, N362, N378);
xor XOR2 (N721, N716, N702);
or OR2 (N722, N445, N505);
or OR2 (N723, N708, N720);
xor XOR2 (N724, N194, N450);
buf BUF1 (N725, N707);
not NOT1 (N726, N715);
nand NAND2 (N727, N725, N145);
and AND3 (N728, N723, N86, N366);
buf BUF1 (N729, N724);
and AND3 (N730, N727, N534, N541);
buf BUF1 (N731, N713);
nand NAND4 (N732, N730, N238, N225, N50);
nor NOR3 (N733, N732, N676, N47);
xor XOR2 (N734, N728, N321);
not NOT1 (N735, N719);
xor XOR2 (N736, N722, N317);
nor NOR4 (N737, N733, N121, N604, N538);
not NOT1 (N738, N736);
buf BUF1 (N739, N721);
xor XOR2 (N740, N738, N107);
and AND3 (N741, N735, N254, N85);
xor XOR2 (N742, N734, N467);
not NOT1 (N743, N737);
nand NAND3 (N744, N739, N223, N672);
xor XOR2 (N745, N731, N389);
and AND4 (N746, N744, N616, N451, N134);
nor NOR4 (N747, N743, N394, N586, N417);
and AND4 (N748, N729, N247, N42, N178);
or OR4 (N749, N748, N546, N165, N323);
xor XOR2 (N750, N717, N202);
buf BUF1 (N751, N745);
and AND2 (N752, N741, N311);
xor XOR2 (N753, N747, N565);
nand NAND3 (N754, N746, N228, N511);
nand NAND2 (N755, N726, N506);
buf BUF1 (N756, N751);
xor XOR2 (N757, N752, N635);
nand NAND3 (N758, N757, N26, N290);
nor NOR3 (N759, N756, N339, N28);
and AND3 (N760, N754, N413, N37);
not NOT1 (N761, N759);
or OR3 (N762, N749, N523, N637);
nand NAND3 (N763, N760, N392, N499);
and AND3 (N764, N742, N116, N584);
nor NOR2 (N765, N755, N467);
xor XOR2 (N766, N763, N196);
nand NAND4 (N767, N750, N578, N597, N413);
buf BUF1 (N768, N758);
xor XOR2 (N769, N761, N602);
and AND3 (N770, N766, N498, N212);
or OR2 (N771, N753, N563);
or OR2 (N772, N771, N645);
not NOT1 (N773, N762);
and AND3 (N774, N772, N557, N217);
or OR2 (N775, N773, N733);
xor XOR2 (N776, N765, N507);
and AND3 (N777, N740, N25, N310);
buf BUF1 (N778, N764);
buf BUF1 (N779, N777);
xor XOR2 (N780, N774, N550);
or OR2 (N781, N779, N116);
nor NOR4 (N782, N780, N470, N539, N457);
buf BUF1 (N783, N769);
not NOT1 (N784, N767);
nor NOR4 (N785, N778, N207, N585, N48);
and AND3 (N786, N776, N364, N486);
nor NOR2 (N787, N781, N57);
or OR4 (N788, N782, N511, N309, N531);
buf BUF1 (N789, N770);
buf BUF1 (N790, N787);
xor XOR2 (N791, N790, N556);
and AND4 (N792, N791, N309, N551, N34);
not NOT1 (N793, N768);
buf BUF1 (N794, N792);
and AND3 (N795, N794, N378, N780);
or OR4 (N796, N788, N488, N200, N351);
buf BUF1 (N797, N793);
not NOT1 (N798, N786);
buf BUF1 (N799, N784);
buf BUF1 (N800, N795);
nand NAND2 (N801, N785, N448);
nor NOR3 (N802, N789, N358, N510);
nand NAND2 (N803, N799, N98);
xor XOR2 (N804, N783, N519);
xor XOR2 (N805, N711, N488);
or OR3 (N806, N796, N336, N747);
buf BUF1 (N807, N802);
xor XOR2 (N808, N797, N689);
not NOT1 (N809, N806);
and AND3 (N810, N805, N529, N126);
buf BUF1 (N811, N775);
or OR2 (N812, N804, N324);
and AND2 (N813, N811, N747);
buf BUF1 (N814, N798);
xor XOR2 (N815, N801, N128);
xor XOR2 (N816, N807, N769);
nand NAND3 (N817, N812, N486, N182);
nand NAND2 (N818, N814, N117);
nor NOR4 (N819, N816, N8, N659, N752);
nor NOR4 (N820, N803, N485, N373, N679);
buf BUF1 (N821, N815);
and AND2 (N822, N800, N3);
not NOT1 (N823, N822);
not NOT1 (N824, N818);
not NOT1 (N825, N823);
and AND4 (N826, N810, N408, N695, N52);
or OR2 (N827, N821, N581);
or OR3 (N828, N824, N335, N607);
or OR4 (N829, N827, N383, N637, N304);
and AND2 (N830, N808, N408);
xor XOR2 (N831, N826, N640);
buf BUF1 (N832, N831);
nor NOR2 (N833, N828, N510);
nor NOR4 (N834, N829, N704, N535, N74);
nand NAND2 (N835, N817, N771);
xor XOR2 (N836, N835, N647);
xor XOR2 (N837, N825, N29);
or OR4 (N838, N832, N189, N30, N498);
or OR2 (N839, N833, N504);
or OR3 (N840, N820, N808, N105);
nor NOR4 (N841, N813, N500, N756, N7);
nand NAND4 (N842, N819, N502, N127, N598);
and AND3 (N843, N839, N329, N776);
and AND4 (N844, N834, N45, N408, N371);
or OR4 (N845, N842, N814, N623, N581);
and AND3 (N846, N841, N622, N570);
buf BUF1 (N847, N830);
xor XOR2 (N848, N840, N548);
and AND4 (N849, N843, N811, N596, N756);
or OR2 (N850, N846, N246);
nor NOR2 (N851, N847, N123);
buf BUF1 (N852, N845);
nor NOR4 (N853, N848, N168, N714, N40);
or OR4 (N854, N850, N543, N90, N183);
buf BUF1 (N855, N837);
nand NAND2 (N856, N844, N476);
xor XOR2 (N857, N838, N676);
nor NOR2 (N858, N854, N247);
buf BUF1 (N859, N851);
nand NAND4 (N860, N857, N498, N339, N592);
and AND3 (N861, N856, N535, N525);
nand NAND3 (N862, N809, N614, N493);
not NOT1 (N863, N855);
or OR2 (N864, N859, N462);
xor XOR2 (N865, N853, N624);
and AND4 (N866, N865, N714, N751, N31);
buf BUF1 (N867, N861);
not NOT1 (N868, N866);
not NOT1 (N869, N860);
nor NOR2 (N870, N849, N866);
and AND4 (N871, N836, N197, N251, N529);
not NOT1 (N872, N863);
xor XOR2 (N873, N871, N851);
buf BUF1 (N874, N872);
and AND4 (N875, N873, N414, N283, N161);
or OR3 (N876, N869, N88, N174);
and AND3 (N877, N867, N527, N188);
not NOT1 (N878, N864);
not NOT1 (N879, N870);
not NOT1 (N880, N858);
or OR4 (N881, N874, N116, N462, N246);
not NOT1 (N882, N875);
not NOT1 (N883, N852);
and AND4 (N884, N883, N658, N42, N344);
nor NOR4 (N885, N882, N21, N425, N464);
buf BUF1 (N886, N877);
buf BUF1 (N887, N881);
not NOT1 (N888, N878);
buf BUF1 (N889, N880);
nor NOR2 (N890, N886, N38);
and AND3 (N891, N885, N384, N838);
or OR2 (N892, N876, N365);
buf BUF1 (N893, N862);
buf BUF1 (N894, N891);
and AND3 (N895, N892, N659, N647);
or OR3 (N896, N888, N206, N801);
not NOT1 (N897, N890);
xor XOR2 (N898, N896, N429);
xor XOR2 (N899, N884, N470);
and AND3 (N900, N889, N507, N195);
nor NOR2 (N901, N897, N568);
or OR4 (N902, N895, N803, N286, N610);
and AND2 (N903, N900, N458);
not NOT1 (N904, N902);
not NOT1 (N905, N903);
xor XOR2 (N906, N879, N422);
or OR4 (N907, N898, N186, N874, N790);
nand NAND3 (N908, N899, N112, N202);
nor NOR2 (N909, N887, N116);
xor XOR2 (N910, N906, N683);
nand NAND4 (N911, N893, N202, N230, N590);
not NOT1 (N912, N901);
nor NOR3 (N913, N908, N297, N490);
nand NAND2 (N914, N912, N737);
buf BUF1 (N915, N913);
nor NOR4 (N916, N914, N505, N158, N341);
nand NAND3 (N917, N909, N763, N566);
not NOT1 (N918, N917);
nand NAND4 (N919, N916, N202, N236, N179);
buf BUF1 (N920, N915);
nor NOR3 (N921, N919, N98, N418);
xor XOR2 (N922, N905, N626);
nand NAND4 (N923, N918, N543, N732, N322);
nor NOR4 (N924, N911, N100, N569, N18);
and AND2 (N925, N894, N538);
nor NOR2 (N926, N868, N631);
xor XOR2 (N927, N926, N640);
and AND3 (N928, N925, N847, N507);
and AND2 (N929, N907, N149);
xor XOR2 (N930, N927, N655);
xor XOR2 (N931, N923, N597);
xor XOR2 (N932, N931, N544);
not NOT1 (N933, N932);
or OR2 (N934, N904, N558);
nand NAND4 (N935, N929, N835, N113, N585);
and AND3 (N936, N924, N371, N358);
and AND4 (N937, N928, N462, N787, N62);
or OR4 (N938, N936, N882, N309, N369);
nor NOR4 (N939, N935, N524, N189, N657);
or OR3 (N940, N934, N158, N162);
not NOT1 (N941, N938);
or OR3 (N942, N922, N306, N445);
nand NAND4 (N943, N942, N499, N899, N225);
nand NAND3 (N944, N940, N112, N202);
or OR2 (N945, N930, N378);
or OR4 (N946, N937, N740, N24, N763);
nand NAND4 (N947, N920, N875, N561, N841);
and AND2 (N948, N945, N475);
nor NOR3 (N949, N921, N941, N856);
nand NAND2 (N950, N734, N157);
or OR3 (N951, N943, N463, N564);
xor XOR2 (N952, N949, N89);
nor NOR3 (N953, N910, N228, N524);
buf BUF1 (N954, N947);
and AND2 (N955, N948, N709);
buf BUF1 (N956, N955);
buf BUF1 (N957, N944);
xor XOR2 (N958, N956, N487);
or OR4 (N959, N933, N663, N552, N274);
xor XOR2 (N960, N946, N365);
and AND4 (N961, N958, N493, N366, N280);
xor XOR2 (N962, N950, N30);
nand NAND2 (N963, N957, N63);
nor NOR3 (N964, N961, N950, N317);
and AND4 (N965, N964, N705, N1, N446);
or OR2 (N966, N954, N851);
nand NAND4 (N967, N963, N710, N8, N211);
buf BUF1 (N968, N966);
and AND2 (N969, N951, N226);
xor XOR2 (N970, N965, N234);
nand NAND4 (N971, N952, N756, N843, N150);
xor XOR2 (N972, N969, N926);
xor XOR2 (N973, N971, N58);
xor XOR2 (N974, N962, N709);
nor NOR2 (N975, N972, N228);
xor XOR2 (N976, N973, N915);
buf BUF1 (N977, N976);
xor XOR2 (N978, N960, N79);
nand NAND3 (N979, N970, N768, N84);
buf BUF1 (N980, N953);
nand NAND3 (N981, N978, N735, N186);
and AND3 (N982, N977, N636, N554);
xor XOR2 (N983, N975, N566);
or OR4 (N984, N982, N476, N778, N950);
buf BUF1 (N985, N968);
not NOT1 (N986, N959);
nor NOR4 (N987, N979, N367, N561, N217);
or OR4 (N988, N980, N409, N158, N885);
or OR3 (N989, N974, N522, N344);
nor NOR4 (N990, N981, N437, N804, N217);
buf BUF1 (N991, N990);
nor NOR3 (N992, N967, N848, N337);
or OR3 (N993, N983, N222, N637);
and AND3 (N994, N984, N492, N457);
xor XOR2 (N995, N989, N66);
not NOT1 (N996, N993);
nor NOR3 (N997, N992, N614, N710);
xor XOR2 (N998, N995, N463);
xor XOR2 (N999, N987, N478);
xor XOR2 (N1000, N985, N507);
or OR3 (N1001, N991, N87, N108);
and AND4 (N1002, N998, N631, N807, N937);
not NOT1 (N1003, N994);
and AND4 (N1004, N986, N366, N525, N2);
and AND3 (N1005, N999, N901, N149);
buf BUF1 (N1006, N939);
not NOT1 (N1007, N1002);
xor XOR2 (N1008, N1001, N512);
or OR3 (N1009, N997, N440, N687);
nand NAND2 (N1010, N1005, N87);
nand NAND3 (N1011, N988, N76, N718);
and AND2 (N1012, N1006, N826);
xor XOR2 (N1013, N1004, N557);
or OR4 (N1014, N1000, N782, N660, N72);
nor NOR2 (N1015, N996, N683);
nand NAND4 (N1016, N1003, N830, N219, N130);
endmodule